module s38584(blif_clk_net, blif_reset_net, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972, d_out_1, q_in_1, d_out_2, qn_in_2, d_out_3, q_in_3, d_out_4, q_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, q_in_7, d_out_8, q_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, d_out_12, q_in_12, d_out_13, qn_in_13, d_out_14, qn_in_14, d_out_15, qn_in_15, d_out_16, qn_in_16, d_out_17, q_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, qn_in_20, d_out_21, q_in_21, d_out_22, qn_in_22, d_out_23, q_in_23, d_out_24, q_in_24, d_out_25, q_in_25, d_out_26, qn_in_26, d_out_27, q_in_27, d_out_28, q_in_28, d_out_29, qn_in_29, d_out_30, qn_in_30, d_out_31, qn_in_31, d_out_32, qn_in_32, d_out_33, q_in_33, d_out_34, qn_in_34, d_out_35, q_in_35, d_out_36, qn_in_36, d_out_37, qn_in_37, d_out_38, q_in_38, d_out_39, q_in_39, d_out_40, qn_in_40, d_out_41, qn_in_41, d_out_42, qn_in_42, d_out_43, qn_in_43, d_out_44, q_in_44, d_out_45, qn_in_45, d_out_46, q_in_46, d_out_47, qn_in_47, d_out_48, q_in_48, d_out_49, q_in_49, d_out_50, qn_in_50, d_out_51, qn_in_51, d_out_52, qn_in_52, d_out_53, qn_in_53, d_out_54, qn_in_54, d_out_55, qn_in_55, d_out_56, qn_in_56, d_out_57, q_in_57, d_out_58, q_in_58, d_out_59, qn_in_59, d_out_60, q_in_60, d_out_61, q_in_61, d_out_62, q_in_62, d_out_63, qn_in_63, d_out_64, q_in_64, d_out_65, qn_in_65, d_out_66, q_in_66, d_out_67, qn_in_67, d_out_68, q_in_68, d_out_69, qn_in_69, d_out_70, q_in_70, d_out_71, qn_in_71, d_out_72, q_in_72, d_out_73, qn_in_73, d_out_74, qn_in_74, d_out_75, q_in_75, d_out_76, q_in_76, d_out_77, qn_in_77, d_out_78, q_in_78, d_out_79, qn_in_79, d_out_80, q_in_80, d_out_81, qn_in_81, d_out_82, q_in_82, d_out_83, q_in_83, d_out_84, qn_in_84, d_out_85, q_in_85, d_out_86, q_in_86, d_out_87, q_in_87, d_out_88, qn_in_88, d_out_89, q_in_89, d_out_90, qn_in_90, d_out_91, q_in_91, d_out_92, qn_in_92, d_out_93, q_in_93, d_out_94, qn_in_94, d_out_95, q_in_95, d_out_96, q_in_96, d_out_97, qn_in_97, d_out_98, q_in_98, d_out_99, q_in_99, d_out_100, qn_in_100, d_out_101, q_in_101, d_out_102, q_in_102, d_out_103, q_in_103, d_out_104, q_in_104, d_out_105, q_in_105, d_out_106, qn_in_106, d_out_107, q_in_107, d_out_108, q_in_108, d_out_109, qn_in_109, d_out_110, qn_in_110, d_out_111, qn_in_111, d_out_112, q_in_112, d_out_113, qn_in_113, d_out_114, qn_in_114, d_out_115, qn_in_115, d_out_116, q_in_116, d_out_117, q_in_117, d_out_118, q_in_118, d_out_119, q_in_119, d_out_120, q_in_120, d_out_121, q_in_121, d_out_122, q_in_122, d_out_123, q_in_123, d_out_124, q_in_124, d_out_125, q_in_125, d_out_126, q_in_126, d_out_127, q_in_127, d_out_128, q_in_128, d_out_129, q_in_129, d_out_130, q_in_130, d_out_131, q_in_131, d_out_132, q_in_132, d_out_133, q_in_133, d_out_134, q_in_134, d_out_135, q_in_135, d_out_136, q_in_136, d_out_137, qn_in_137, d_out_138, q_in_138, d_out_139, q_in_139, d_out_140, qn_in_140, d_out_141, qn_in_141, d_out_142, q_in_142, d_out_143, q_in_143, d_out_144, qn_in_144, d_out_145, q_in_145, d_out_146, qn_in_146, d_out_147, qn_in_147, d_out_148, q_in_148, d_out_149, q_in_149, d_out_150, q_in_150, d_out_151, q_in_151, d_out_152, qn_in_152, d_out_153, qn_in_153, d_out_154, q_in_154, d_out_155, q_in_155, d_out_156, q_in_156, d_out_157, q_in_157, d_out_158, q_in_158, d_out_159, q_in_159, d_out_160, q_in_160, d_out_161, q_in_161, d_out_162, q_in_162, d_out_163, q_in_163, d_out_164, q_in_164, d_out_165, q_in_165, d_out_166, q_in_166, d_out_167, q_in_167, d_out_168, q_in_168, d_out_169, qn_in_169, d_out_170, qn_in_170, d_out_171, q_in_171, d_out_172, q_in_172, d_out_173, q_in_173, d_out_174, q_in_174, d_out_175, q_in_175, d_out_176, q_in_176, d_out_177, q_in_177, d_out_178, q_in_178, d_out_179, q_in_179, d_out_180, q_in_180, d_out_181, q_in_181, d_out_182, q_in_182, d_out_183, q_in_183, d_out_184, q_in_184, d_out_185, q_in_185, d_out_186, q_in_186, d_out_187, q_in_187, d_out_188, q_in_188, d_out_189, q_in_189, d_out_190, q_in_190, d_out_191, q_in_191, d_out_192, q_in_192, d_out_193, q_in_193, d_out_194, q_in_194, d_out_195, q_in_195, d_out_196, q_in_196, d_out_197, q_in_197, d_out_198, q_in_198, d_out_199, q_in_199, d_out_200, q_in_200, d_out_201, q_in_201, d_out_202, qn_in_202, d_out_203, q_in_203, d_out_204, q_in_204, d_out_205, q_in_205, d_out_206, q_in_206, d_out_207, qn_in_207, d_out_208, q_in_208, d_out_209, q_in_209, d_out_210, qn_in_210, d_out_211, q_in_211, d_out_212, q_in_212, d_out_213, q_in_213, d_out_214, qn_in_214, d_out_215, qn_in_215, d_out_216, q_in_216, d_out_217, q_in_217, d_out_218, q_in_218, d_out_219, q_in_219, d_out_220, q_in_220, d_out_221, q_in_221, d_out_222, q_in_222, d_out_223, q_in_223, d_out_224, qn_in_224, d_out_225, qn_in_225, d_out_226, q_in_226, d_out_227, q_in_227, d_out_228, q_in_228, d_out_229, q_in_229, d_out_230, q_in_230, d_out_231, qn_in_231, d_out_232, qn_in_232, d_out_233, qn_in_233, d_out_234, qn_in_234, d_out_235, q_in_235, d_out_236, q_in_236, d_out_237, q_in_237, d_out_238, q_in_238, d_out_239, qn_in_239, d_out_240, q_in_240, d_out_241, q_in_241, d_out_242, qn_in_242, d_out_243, qn_in_243, d_out_244, qn_in_244, d_out_245, qn_in_245, d_out_246, qn_in_246, d_out_247, qn_in_247, d_out_248, qn_in_248, d_out_249, qn_in_249, d_out_250, qn_in_250, d_out_251, qn_in_251, d_out_252, qn_in_252, d_out_253, qn_in_253, d_out_254, qn_in_254, d_out_255, qn_in_255, d_out_256, qn_in_256, d_out_257, qn_in_257, d_out_258, qn_in_258, d_out_259, qn_in_259, d_out_260, qn_in_260, d_out_261, q_in_261, d_out_262, q_in_262, d_out_263, qn_in_263, d_out_264, q_in_264, d_out_265, q_in_265, d_out_266, q_in_266, d_out_267, q_in_267, d_out_268, q_in_268, d_out_269, qn_in_269, d_out_270, q_in_270, d_out_271, q_in_271, d_out_272, qn_in_272, d_out_273, q_in_273, d_out_274, q_in_274, d_out_275, qn_in_275, d_out_276, qn_in_276, d_out_277, qn_in_277, d_out_278, qn_in_278, d_out_279, qn_in_279, d_out_280, qn_in_280, d_out_281, qn_in_281, d_out_282, qn_in_282, d_out_283, qn_in_283, d_out_284, qn_in_284, d_out_285, qn_in_285, d_out_286, qn_in_286, d_out_287, qn_in_287, d_out_288, qn_in_288, d_out_289, qn_in_289, d_out_290, qn_in_290, d_out_291, qn_in_291, d_out_292, q_in_292, d_out_293, q_in_293, d_out_294, q_in_294, d_out_295, q_in_295, d_out_296, q_in_296, d_out_297, qn_in_297, d_out_298, qn_in_298, d_out_299, q_in_299, d_out_300, qn_in_300, d_out_301, q_in_301, d_out_302, qn_in_302, d_out_303, q_in_303, d_out_304, q_in_304, d_out_305, q_in_305, d_out_306, q_in_306, d_out_307, qn_in_307, d_out_308, qn_in_308, d_out_309, qn_in_309, d_out_310, qn_in_310, d_out_311, qn_in_311, d_out_312, qn_in_312, d_out_313, qn_in_313, d_out_314, q_in_314, d_out_315, q_in_315, d_out_316, qn_in_316, d_out_317, qn_in_317, d_out_318, qn_in_318, d_out_319, qn_in_319, d_out_320, qn_in_320, d_out_321, qn_in_321, d_out_322, qn_in_322, d_out_323, qn_in_323, d_out_324, qn_in_324, d_out_325, qn_in_325, d_out_326, qn_in_326, d_out_327, qn_in_327, d_out_328, qn_in_328, d_out_329, qn_in_329, d_out_330, q_in_330, d_out_331, q_in_331, d_out_332, q_in_332, d_out_333, q_in_333, d_out_334, q_in_334, d_out_335, q_in_335, d_out_336, qn_in_336, d_out_337, q_in_337, d_out_338, q_in_338, d_out_339, qn_in_339, d_out_340, q_in_340, d_out_341, qn_in_341, d_out_342, qn_in_342, d_out_343, q_in_343, d_out_344, qn_in_344, d_out_345, q_in_345, d_out_346, qn_in_346, d_out_347, qn_in_347, d_out_348, q_in_348, d_out_349, qn_in_349, d_out_350, qn_in_350, d_out_351, q_in_351, d_out_352, q_in_352, d_out_353, q_in_353, d_out_354, q_in_354, d_out_355, q_in_355, d_out_356, q_in_356, d_out_357, q_in_357, d_out_358, q_in_358, d_out_359, q_in_359, d_out_360, q_in_360, d_out_361, q_in_361, d_out_362, q_in_362, d_out_363, q_in_363, d_out_364, qn_in_364, d_out_365, q_in_365, d_out_366, q_in_366, d_out_367, q_in_367, d_out_368, q_in_368, d_out_369, q_in_369, d_out_370, q_in_370, d_out_371, q_in_371, d_out_372, qn_in_372, d_out_373, q_in_373, d_out_374, q_in_374, d_out_375, q_in_375, d_out_376, q_in_376, d_out_377, q_in_377, d_out_378, q_in_378, d_out_379, q_in_379, d_out_380, q_in_380, d_out_381, q_in_381, d_out_382, q_in_382, d_out_383, q_in_383, d_out_384, q_in_384, d_out_385, qn_in_385, d_out_386, q_in_386, d_out_387, q_in_387, d_out_388, q_in_388, d_out_389, q_in_389, d_out_390, q_in_390, d_out_391, q_in_391, d_out_392, q_in_392, d_out_393, q_in_393, d_out_394, q_in_394, d_out_395, q_in_395, d_out_396, q_in_396, d_out_397, q_in_397, d_out_398, q_in_398, d_out_399, q_in_399, d_out_400, q_in_400, d_out_401, q_in_401, d_out_402, qn_in_402, d_out_403, q_in_403, d_out_404, q_in_404, d_out_405, q_in_405, d_out_406, q_in_406, d_out_407, q_in_407, d_out_408, q_in_408, d_out_409, q_in_409, d_out_410, q_in_410, d_out_411, q_in_411, d_out_412, q_in_412, d_out_413, q_in_413, d_out_414, q_in_414, d_out_415, q_in_415, d_out_416, q_in_416, d_out_417, q_in_417, d_out_418, qn_in_418, d_out_419, qn_in_419, d_out_420, qn_in_420, d_out_421, qn_in_421, d_out_422, qn_in_422, d_out_423, qn_in_423, d_out_424, qn_in_424, d_out_425, qn_in_425, d_out_426, qn_in_426, d_out_427, q_in_427, d_out_428, q_in_428, d_out_429, q_in_429, d_out_430, q_in_430, d_out_431, q_in_431, d_out_432, q_in_432, d_out_433, q_in_433, d_out_434, q_in_434, d_out_435, q_in_435, d_out_436, q_in_436, d_out_437, q_in_437, d_out_438, q_in_438, d_out_439, q_in_439, d_out_440, q_in_440, d_out_441, q_in_441, d_out_442, q_in_442, d_out_443, q_in_443, d_out_444, q_in_444, d_out_445, q_in_445, d_out_446, q_in_446, d_out_447, q_in_447, d_out_448, q_in_448, d_out_449, q_in_449, d_out_450, q_in_450, d_out_451, q_in_451, d_out_452, q_in_452, d_out_453, q_in_453, d_out_454, q_in_454, d_out_455, q_in_455, d_out_456, q_in_456, d_out_457, q_in_457, d_out_458, q_in_458, d_out_459, q_in_459, d_out_460, q_in_460, d_out_461, q_in_461, d_out_462, q_in_462, d_out_463, q_in_463, d_out_464, q_in_464, d_out_465, q_in_465, d_out_466, q_in_466, d_out_467, q_in_467, d_out_468, q_in_468, d_out_469, q_in_469, d_out_470, qn_in_470, d_out_471, q_in_471, d_out_472, q_in_472, d_out_473, q_in_473, d_out_474, q_in_474, d_out_475, q_in_475, d_out_476, q_in_476, d_out_477, q_in_477, d_out_478, q_in_478, d_out_479, q_in_479, d_out_480, q_in_480, d_out_481, q_in_481, d_out_482, q_in_482, d_out_483, q_in_483, d_out_484, q_in_484, d_out_485, q_in_485, d_out_486, q_in_486, d_out_487, q_in_487, d_out_488, q_in_488, d_out_489, q_in_489, d_out_490, q_in_490, d_out_491, q_in_491, d_out_492, q_in_492, d_out_493, q_in_493, d_out_494, q_in_494, d_out_495, q_in_495, d_out_496, q_in_496, d_out_497, q_in_497, d_out_498, q_in_498, d_out_499, q_in_499, d_out_500, q_in_500, d_out_501, q_in_501, d_out_502, q_in_502, d_out_503, q_in_503, d_out_504, q_in_504, d_out_505, q_in_505, d_out_506, q_in_506, d_out_507, q_in_507, d_out_508, q_in_508, d_out_509, q_in_509, d_out_510, q_in_510, d_out_511, q_in_511, d_out_512, q_in_512, d_out_513, q_in_513, d_out_514, q_in_514, d_out_515, q_in_515, d_out_516, qn_in_516, d_out_517, q_in_517, d_out_518, q_in_518, d_out_519, q_in_519, d_out_520, q_in_520, d_out_521, q_in_521, d_out_522, q_in_522, d_out_523, q_in_523, d_out_524, q_in_524, d_out_525, q_in_525, d_out_526, q_in_526, d_out_527, q_in_527, d_out_528, q_in_528, d_out_529, q_in_529, d_out_530, q_in_530, d_out_531, q_in_531, d_out_532, q_in_532, d_out_533, q_in_533, d_out_534, q_in_534, d_out_535, q_in_535, d_out_536, q_in_536, d_out_537, q_in_537, d_out_538, q_in_538, d_out_539, q_in_539, d_out_540, q_in_540, d_out_541, q_in_541, d_out_542, q_in_542, d_out_543, q_in_543, d_out_544, q_in_544, d_out_545, q_in_545, d_out_546, q_in_546, d_out_547, q_in_547, d_out_548, q_in_548, d_out_549, q_in_549, d_out_550, qn_in_550, d_out_551, qn_in_551, d_out_552, q_in_552, d_out_553, qn_in_553, d_out_554, qn_in_554, d_out_555, qn_in_555, d_out_556, qn_in_556, d_out_557, q_in_557, d_out_558, qn_in_558, d_out_559, q_in_559, d_out_560, q_in_560, d_out_561, q_in_561, d_out_562, q_in_562, d_out_563, q_in_563, d_out_564, q_in_564, d_out_565, q_in_565, d_out_566, qn_in_566, d_out_567, q_in_567, d_out_568, qn_in_568, d_out_569, q_in_569, d_out_570, q_in_570, d_out_571, q_in_571, d_out_572, qn_in_572, d_out_573, q_in_573, d_out_574, q_in_574, d_out_575, qn_in_575, d_out_576, qn_in_576, d_out_577, qn_in_577, d_out_578, qn_in_578, d_out_579, q_in_579, d_out_580, q_in_580, d_out_581, qn_in_581, d_out_582, qn_in_582, d_out_583, qn_in_583, d_out_584, q_in_584, d_out_585, qn_in_585, d_out_586, qn_in_586, d_out_587, q_in_587, d_out_588, q_in_588, d_out_589, q_in_589, d_out_590, q_in_590, d_out_591, q_in_591, d_out_592, q_in_592, d_out_593, q_in_593, d_out_594, q_in_594, d_out_595, qn_in_595, d_out_596, q_in_596, d_out_597, q_in_597, d_out_598, q_in_598, d_out_599, q_in_599, d_out_600, qn_in_600, d_out_601, q_in_601, d_out_602, qn_in_602, d_out_603, q_in_603, d_out_604, q_in_604, d_out_605, q_in_605, d_out_606, q_in_606, d_out_607, q_in_607, d_out_608, q_in_608, d_out_609, q_in_609, d_out_610, q_in_610, d_out_611, q_in_611, d_out_612, q_in_612, d_out_613, q_in_613, d_out_614, q_in_614, d_out_615, q_in_615, d_out_616, q_in_616, d_out_617, q_in_617, d_out_618, q_in_618, d_out_619, q_in_619, d_out_620, q_in_620, d_out_621, q_in_621, d_out_622, q_in_622, d_out_623, q_in_623, d_out_624, q_in_624, d_out_625, q_in_625, d_out_626, q_in_626, d_out_627, q_in_627, d_out_628, qn_in_628, d_out_629, q_in_629, d_out_630, qn_in_630, d_out_631, qn_in_631, d_out_632, q_in_632, d_out_633, q_in_633, d_out_634, q_in_634, d_out_635, q_in_635, d_out_636, q_in_636, d_out_637, q_in_637, d_out_638, q_in_638, d_out_639, q_in_639, d_out_640, q_in_640, d_out_641, q_in_641, d_out_642, q_in_642, d_out_643, q_in_643, d_out_644, q_in_644, d_out_645, q_in_645, d_out_646, q_in_646, d_out_647, qn_in_647, d_out_648, q_in_648, d_out_649, q_in_649, d_out_650, q_in_650, d_out_651, q_in_651, d_out_652, q_in_652, d_out_653, q_in_653, d_out_654, q_in_654, d_out_655, q_in_655, d_out_656, q_in_656, d_out_657, q_in_657, d_out_658, q_in_658, d_out_659, q_in_659, d_out_660, q_in_660, d_out_661, q_in_661, d_out_662, q_in_662, d_out_663, q_in_663, d_out_664, q_in_664, d_out_665, q_in_665, d_out_666, q_in_666, d_out_667, q_in_667, d_out_668, q_in_668, d_out_669, q_in_669, d_out_670, q_in_670, d_out_671, qn_in_671, d_out_672, q_in_672, d_out_673, q_in_673, d_out_674, qn_in_674, d_out_675, q_in_675, d_out_676, q_in_676, d_out_677, q_in_677, d_out_678, q_in_678, d_out_679, q_in_679, d_out_680, q_in_680, d_out_681, q_in_681, d_out_682, q_in_682, d_out_683, q_in_683, d_out_684, q_in_684, d_out_685, q_in_685, d_out_686, q_in_686, d_out_687, q_in_687, d_out_688, q_in_688, d_out_689, q_in_689, d_out_690, q_in_690, d_out_691, q_in_691, d_out_692, q_in_692, d_out_693, q_in_693, d_out_694, q_in_694, d_out_695, q_in_695, d_out_696, q_in_696, d_out_697, q_in_697, d_out_698, q_in_698, d_out_699, q_in_699, d_out_700, q_in_700, d_out_701, q_in_701, d_out_702, q_in_702, d_out_703, qn_in_703, d_out_704, q_in_704, d_out_705, q_in_705, d_out_706, qn_in_706, d_out_707, qn_in_707, d_out_708, qn_in_708, d_out_709, q_in_709, d_out_710, q_in_710, d_out_711, q_in_711, d_out_712, q_in_712, d_out_713, q_in_713, d_out_714, q_in_714, d_out_715, q_in_715, d_out_716, qn_in_716, d_out_717, q_in_717, d_out_718, q_in_718, d_out_719, q_in_719, d_out_720, q_in_720, d_out_721, q_in_721, d_out_722, q_in_722, d_out_723, q_in_723, d_out_724, q_in_724, d_out_725, qn_in_725, d_out_726, q_in_726, d_out_727, q_in_727, d_out_728, q_in_728, d_out_729, q_in_729, d_out_730, q_in_730, d_out_731, q_in_731, d_out_732, q_in_732, d_out_733, q_in_733, d_out_734, q_in_734, d_out_735, q_in_735, d_out_736, q_in_736, d_out_737, q_in_737, d_out_738, q_in_738, d_out_739, q_in_739, d_out_740, q_in_740, d_out_741, q_in_741, d_out_742, q_in_742, d_out_743, q_in_743, d_out_744, q_in_744, d_out_745, q_in_745, d_out_746, q_in_746, d_out_747, q_in_747, d_out_748, q_in_748, d_out_749, q_in_749, d_out_750, q_in_750, d_out_751, q_in_751, d_out_752, q_in_752, d_out_753, q_in_753, d_out_754, q_in_754, d_out_755, q_in_755, d_out_756, q_in_756, d_out_757, q_in_757, d_out_758, q_in_758, d_out_759, q_in_759, d_out_760, q_in_760, d_out_761, q_in_761, d_out_762, q_in_762, d_out_763, qn_in_763, d_out_764, q_in_764, d_out_765, qn_in_765, d_out_766, q_in_766, d_out_767, q_in_767, d_out_768, q_in_768, d_out_769, q_in_769, d_out_770, q_in_770, d_out_771, q_in_771, d_out_772, q_in_772, d_out_773, q_in_773, d_out_774, q_in_774, d_out_775, q_in_775, d_out_776, qn_in_776, d_out_777, qn_in_777, d_out_778, q_in_778, d_out_779, q_in_779, d_out_780, q_in_780, d_out_781, q_in_781, d_out_782, q_in_782, d_out_783, q_in_783, d_out_784, q_in_784, d_out_785, q_in_785, d_out_786, q_in_786, d_out_787, q_in_787, d_out_788, q_in_788, d_out_789, q_in_789, d_out_790, q_in_790, d_out_791, q_in_791, d_out_792, q_in_792, d_out_793, q_in_793, d_out_794, q_in_794, d_out_795, q_in_795, d_out_796, q_in_796, d_out_797, q_in_797, d_out_798, q_in_798, d_out_799, q_in_799, d_out_800, q_in_800, d_out_801, q_in_801, d_out_802, q_in_802, d_out_803, q_in_803, d_out_804, q_in_804, d_out_805, q_in_805, d_out_806, q_in_806, d_out_807, q_in_807, d_out_808, q_in_808, d_out_809, q_in_809, d_out_810, q_in_810, d_out_811, q_in_811, d_out_812, q_in_812, d_out_813, qn_in_813, d_out_814, qn_in_814, d_out_815, qn_in_815, d_out_816, q_in_816, d_out_817, qn_in_817, d_out_818, qn_in_818, d_out_819, qn_in_819, d_out_820, q_in_820, d_out_821, q_in_821, d_out_822, q_in_822, d_out_823, q_in_823, d_out_824, q_in_824, d_out_825, q_in_825, d_out_826, q_in_826, d_out_827, qn_in_827, d_out_828, qn_in_828, d_out_829, qn_in_829, d_out_830, qn_in_830, d_out_831, q_in_831, d_out_832, q_in_832, d_out_833, q_in_833, d_out_834, q_in_834, d_out_835, q_in_835, d_out_836, q_in_836, d_out_837, q_in_837, d_out_838, q_in_838, d_out_839, q_in_839, d_out_840, q_in_840, d_out_841, q_in_841, d_out_842, q_in_842, d_out_843, q_in_843, d_out_844, q_in_844, d_out_845, q_in_845, d_out_846, q_in_846, d_out_847, q_in_847, d_out_848, q_in_848, d_out_849, q_in_849, d_out_850, q_in_850, d_out_851, q_in_851, d_out_852, q_in_852, d_out_853, q_in_853, d_out_854, q_in_854, d_out_855, q_in_855, d_out_856, q_in_856, d_out_857, q_in_857, d_out_858, q_in_858, d_out_859, q_in_859, d_out_860, q_in_860, d_out_861, qn_in_861, d_out_862, qn_in_862, d_out_863, qn_in_863, d_out_864, q_in_864, d_out_865, q_in_865, d_out_866, q_in_866, d_out_867, q_in_867, d_out_868, q_in_868, d_out_869, q_in_869, d_out_870, q_in_870, d_out_871, q_in_871, d_out_872, q_in_872, d_out_873, q_in_873, d_out_874, q_in_874, d_out_875, q_in_875, d_out_876, q_in_876, d_out_877, q_in_877, d_out_878, q_in_878, d_out_879, q_in_879, d_out_880, qn_in_880, d_out_881, q_in_881, d_out_882, q_in_882, d_out_883, q_in_883, d_out_884, qn_in_884, d_out_885, qn_in_885, d_out_886, q_in_886, d_out_887, q_in_887, d_out_888, q_in_888, d_out_889, q_in_889, d_out_890, q_in_890, d_out_891, q_in_891, d_out_892, q_in_892, d_out_893, q_in_893, d_out_894, q_in_894, d_out_895, q_in_895, d_out_896, q_in_896, d_out_897, q_in_897, d_out_898, q_in_898, d_out_899, q_in_899, d_out_900, q_in_900, d_out_901, q_in_901, d_out_902, q_in_902, d_out_903, q_in_903, d_out_904, q_in_904, d_out_905, q_in_905, d_out_906, q_in_906, d_out_907, q_in_907, d_out_908, q_in_908, d_out_909, q_in_909, d_out_910, q_in_910, d_out_911, q_in_911, d_out_912, q_in_912, d_out_913, q_in_913, d_out_914, q_in_914, d_out_915, q_in_915, d_out_916, q_in_916, d_out_917, q_in_917, d_out_918, q_in_918, d_out_919, q_in_919, d_out_920, q_in_920, d_out_921, q_in_921, d_out_922, q_in_922, d_out_923, q_in_923, d_out_924, q_in_924, d_out_925, q_in_925, d_out_926, q_in_926, d_out_927, qn_in_927, d_out_928, q_in_928, d_out_929, q_in_929, d_out_930, q_in_930, d_out_931, q_in_931, d_out_932, q_in_932, d_out_933, qn_in_933, d_out_934, q_in_934, d_out_935, q_in_935, d_out_936, q_in_936, d_out_937, q_in_937, d_out_938, q_in_938, d_out_939, q_in_939, d_out_940, qn_in_940, d_out_941, qn_in_941, d_out_942, qn_in_942, d_out_943, qn_in_943, d_out_944, qn_in_944, d_out_945, qn_in_945, d_out_946, q_in_946, d_out_947, q_in_947, d_out_948, q_in_948, d_out_949, q_in_949, d_out_950, q_in_950, d_out_951, q_in_951, d_out_952, qn_in_952, d_out_953, qn_in_953, d_out_954, q_in_954, d_out_955, q_in_955, d_out_956, q_in_956, d_out_957, q_in_957, d_out_958, q_in_958, d_out_959, qn_in_959, d_out_960, q_in_960, d_out_961, q_in_961, d_out_962, qn_in_962, d_out_963, q_in_963, d_out_964, qn_in_964, d_out_965, q_in_965, d_out_966, q_in_966, d_out_967, qn_in_967, d_out_968, qn_in_968, d_out_969, q_in_969, d_out_970, q_in_970, d_out_971, q_in_971, d_out_972, q_in_972, d_out_973, q_in_973, d_out_974, q_in_974, d_out_975, q_in_975, d_out_976, qn_in_976, d_out_977, qn_in_977, d_out_978, q_in_978, d_out_979, q_in_979, d_out_980, q_in_980, d_out_981, q_in_981, d_out_982, q_in_982, d_out_983, q_in_983, d_out_984, q_in_984, d_out_985, q_in_985, d_out_986, q_in_986, d_out_987, q_in_987, d_out_988, q_in_988, d_out_989, q_in_989, d_out_990, q_in_990, d_out_991, q_in_991, d_out_992, q_in_992, d_out_993, q_in_993, d_out_994, q_in_994, d_out_995, q_in_995, d_out_996, q_in_996, d_out_997, q_in_997, d_out_998, q_in_998, d_out_999, q_in_999, d_out_1000, q_in_1000, d_out_1001, q_in_1001, d_out_1002, q_in_1002, d_out_1003, q_in_1003, d_out_1004, q_in_1004, d_out_1005, q_in_1005, d_out_1006, q_in_1006, d_out_1007, q_in_1007, d_out_1008, q_in_1008, d_out_1009, q_in_1009, d_out_1010, q_in_1010, d_out_1011, q_in_1011, d_out_1012, q_in_1012, d_out_1013, q_in_1013, d_out_1014, q_in_1014, d_out_1015, q_in_1015, d_out_1016, q_in_1016, d_out_1017, q_in_1017, d_out_1018, q_in_1018, d_out_1019, q_in_1019, d_out_1020, q_in_1020, d_out_1021, q_in_1021, d_out_1022, q_in_1022, d_out_1023, q_in_1023, d_out_1024, q_in_1024, d_out_1025, q_in_1025, d_out_1026, q_in_1026, d_out_1027, q_in_1027, d_out_1028, q_in_1028, d_out_1029, q_in_1029, d_out_1030, q_in_1030, d_out_1031, q_in_1031, d_out_1032, q_in_1032, d_out_1033, q_in_1033, d_out_1034, q_in_1034, d_out_1035, q_in_1035, d_out_1036, q_in_1036, d_out_1037, q_in_1037, d_out_1038, q_in_1038, d_out_1039, q_in_1039, d_out_1040, q_in_1040, d_out_1041, q_in_1041, d_out_1042, q_in_1042, d_out_1043, q_in_1043, d_out_1044, qn_in_1044, d_out_1045, q_in_1045, d_out_1046, q_in_1046, d_out_1047, q_in_1047, d_out_1048, qn_in_1048, d_out_1049, qn_in_1049, d_out_1050, q_in_1050, d_out_1051, q_in_1051, d_out_1052, q_in_1052, d_out_1053, q_in_1053, d_out_1054, q_in_1054, d_out_1055, q_in_1055, d_out_1056, qn_in_1056, d_out_1057, q_in_1057, d_out_1058, q_in_1058, d_out_1059, q_in_1059, d_out_1060, qn_in_1060, d_out_1061, q_in_1061, d_out_1062, q_in_1062, d_out_1063, q_in_1063, d_out_1064, q_in_1064, d_out_1065, q_in_1065, d_out_1066, q_in_1066, d_out_1067, qn_in_1067, d_out_1068, q_in_1068, d_out_1069, q_in_1069, d_out_1070, q_in_1070, d_out_1071, q_in_1071, d_out_1072, q_in_1072, d_out_1073, q_in_1073, d_out_1074, qn_in_1074, d_out_1075, q_in_1075, d_out_1076, q_in_1076, d_out_1077, q_in_1077, d_out_1078, q_in_1078, d_out_1079, q_in_1079, d_out_1080, q_in_1080, d_out_1081, q_in_1081, d_out_1082, q_in_1082, d_out_1083, q_in_1083, d_out_1084, q_in_1084, d_out_1085, q_in_1085, d_out_1086, q_in_1086, d_out_1087, q_in_1087, d_out_1088, q_in_1088, d_out_1089, q_in_1089, d_out_1090, q_in_1090, d_out_1091, q_in_1091, d_out_1092, q_in_1092, d_out_1093, q_in_1093, d_out_1094, q_in_1094, d_out_1095, q_in_1095, d_out_1096, q_in_1096, d_out_1097, q_in_1097, d_out_1098, q_in_1098, d_out_1099, q_in_1099, d_out_1100, q_in_1100, d_out_1101, q_in_1101, d_out_1102, q_in_1102, d_out_1103, q_in_1103, d_out_1104, q_in_1104, d_out_1105, q_in_1105, d_out_1106, q_in_1106, d_out_1107, q_in_1107, d_out_1108, q_in_1108, d_out_1109, q_in_1109, d_out_1110, q_in_1110, d_out_1111, q_in_1111, d_out_1112, q_in_1112, d_out_1113, q_in_1113, d_out_1114, q_in_1114, d_out_1115, qn_in_1115, d_out_1116, q_in_1116, d_out_1117, q_in_1117, d_out_1118, q_in_1118, d_out_1119, q_in_1119, d_out_1120, q_in_1120, d_out_1121, q_in_1121, d_out_1122, q_in_1122, d_out_1123, q_in_1123, d_out_1124, q_in_1124, d_out_1125, q_in_1125, d_out_1126, q_in_1126, d_out_1127, q_in_1127, d_out_1128, q_in_1128, d_out_1129, q_in_1129, d_out_1130, q_in_1130, d_out_1131, q_in_1131, d_out_1132, q_in_1132, d_out_1133, qn_in_1133, d_out_1134, q_in_1134, d_out_1135, q_in_1135, d_out_1136, q_in_1136, d_out_1137, q_in_1137, d_out_1138, qn_in_1138, d_out_1139, q_in_1139, d_out_1140, q_in_1140, d_out_1141, q_in_1141, d_out_1142, qn_in_1142, d_out_1143, q_in_1143, d_out_1144, q_in_1144, d_out_1145, q_in_1145, d_out_1146, q_in_1146, d_out_1147, q_in_1147, d_out_1148, q_in_1148, d_out_1149, q_in_1149, d_out_1150, q_in_1150, d_out_1151, q_in_1151, d_out_1152, q_in_1152, d_out_1153, qn_in_1153, d_out_1154, q_in_1154, d_out_1155, q_in_1155, d_out_1156, q_in_1156, d_out_1157, q_in_1157, d_out_1158, q_in_1158, d_out_1159, q_in_1159, d_out_1160, q_in_1160, d_out_1161, q_in_1161, d_out_1162, q_in_1162, d_out_1163, q_in_1163, d_out_1164, q_in_1164, d_out_1165, q_in_1165, d_out_1166, q_in_1166, d_out_1167, q_in_1167, d_out_1168, q_in_1168, d_out_1169, qn_in_1169, d_out_1170, q_in_1170, d_out_1171, q_in_1171, d_out_1172, q_in_1172, d_out_1173, q_in_1173, d_out_1174, q_in_1174, d_out_1175, q_in_1175, d_out_1176, q_in_1176, d_out_1177, q_in_1177, d_out_1178, q_in_1178);
input qn_in_418;
input q_in_417;
input q_in_416;
input q_in_415;
input q_in_414;
input q_in_413;
input q_in_412;
input q_in_411;
input q_in_410;
input q_in_409;
input q_in_408;
input q_in_407;
input q_in_406;
input q_in_405;
input q_in_404;
input q_in_403;
input qn_in_402;
input q_in_401;
input q_in_400;
input q_in_926;
input q_in_399;
input q_in_978;
input q_in_398;
input q_in_889;
input qn_in_976;
input q_in_975;
input q_in_397;
input q_in_1154;
input q_in_973;
input qn_in_1153;
input q_in_972;
input q_in_396;
input q_in_395;
input q_in_969;
input qn_in_968;
input q_in_1161;
input qn_in_967;
input q_in_966;
input q_in_965;
input qn_in_964;
input q_in_963;
input qn_in_962;
input q_in_961;
input q_in_1146;
input q_in_960;
input qn_in_959;
input q_in_1144;
input q_in_888;
input q_in_957;
input q_in_394;
input q_in_955;
input q_in_954;
input qn_in_953;
input q_in_393;
input q_in_392;
input q_in_391;
input q_in_390;
input q_in_389;
input q_in_388;
input q_in_387;
input q_in_951;
input q_in_950;
input q_in_386;
input qn_in_385;
input q_in_947;
input q_in_807;
input q_in_384;
input qn_in_944;
input qn_in_943;
input q_in_383;
input qn_in_941;
input q_in_382;
input q_in_381;
input q_in_380;
input q_in_379;
input q_in_378;
input q_in_377;
input q_in_376;
input q_in_375;
input q_in_374;
input q_in_373;
input qn_in_372;
input q_in_371;
input q_in_370;
input q_in_369;
input q_in_368;
input q_in_367;
input q_in_366;
input q_in_365;
input qn_in_364;
input q_in_363;
input q_in_362;
input q_in_361;
input q_in_360;
input q_in_359;
input q_in_358;
input q_in_357;
input q_in_356;
input q_in_355;
input q_in_354;
input q_in_353;
input q_in_352;
input q_in_351;
input qn_in_350;
input qn_in_349;
input q_in_348;
input qn_in_347;
input qn_in_346;
input q_in_345;
input qn_in_344;
input q_in_343;
input qn_in_342;
input qn_in_341;
input q_in_340;
input qn_in_339;
input q_in_338;
input q_in_337;
input qn_in_336;
input q_in_335;
input q_in_334;
input q_in_333;
input q_in_332;
input q_in_331;
input q_in_330;
input qn_in_329;
input qn_in_328;
input qn_in_327;
input qn_in_326;
input qn_in_325;
input qn_in_324;
input qn_in_323;
input qn_in_322;
input qn_in_321;
input qn_in_320;
input qn_in_319;
input qn_in_318;
input qn_in_317;
input qn_in_316;
input q_in_315;
input q_in_1137;
input q_in_1136;
input q_in_1135;
input q_in_1134;
input qn_in_1133;
input q_in_1132;
input q_in_1131;
input q_in_1130;
input q_in_314;
input q_in_841;
input q_in_1129;
input q_in_1128;
input qn_in_313;
input q_in_924;
input q_in_923;
input q_in_922;
input qn_in_312;
input q_in_920;
input q_in_919;
input q_in_918;
input q_in_917;
input qn_in_311;
input qn_in_310;
input q_in_914;
input qn_in_309;
input q_in_912;
input qn_in_308;
input q_in_910;
input q_in_909;
input qn_in_307;
input q_in_907;
input q_in_906;
input q_in_905;
input q_in_904;
input q_in_903;
input q_in_902;
input q_in_901;
input q_in_900;
input q_in_899;
input q_in_898;
input q_in_897;
input q_in_896;
input q_in_306;
input q_in_305;
input q_in_304;
input q_in_303;
input qn_in_302;
input q_in_301;
input qn_in_300;
input q_in_299;
input qn_in_298;
input qn_in_297;
input q_in_296;
input q_in_295;
input q_in_294;
input q_in_293;
input q_in_292;
input qn_in_291;
input qn_in_290;
input qn_in_289;
input qn_in_288;
input qn_in_287;
input qn_in_286;
input qn_in_285;
input qn_in_284;
input qn_in_283;
input qn_in_282;
input qn_in_281;
input qn_in_280;
input qn_in_279;
input qn_in_278;
input qn_in_277;
input qn_in_276;
input qn_in_275;
input q_in_274;
input q_in_874;
input q_in_873;
input q_in_273;
input q_in_871;
input q_in_870;
input q_in_1165;
input q_in_869;
input qn_in_272;
input q_in_937;
input q_in_271;
input q_in_1116;
input q_in_971;
input q_in_868;
input q_in_867;
input q_in_970;
input q_in_270;
input q_in_866;
input qn_in_1115;
input qn_in_269;
input q_in_268;
input q_in_267;
input q_in_266;
input q_in_265;
input q_in_264;
input qn_in_263;
input q_in_262;
input q_in_261;
input qn_in_260;
input qn_in_259;
input qn_in_258;
input qn_in_257;
input qn_in_256;
input qn_in_255;
input qn_in_254;
input qn_in_253;
input qn_in_252;
input qn_in_251;
input qn_in_250;
input qn_in_249;
input qn_in_248;
input qn_in_247;
input qn_in_246;
input qn_in_245;
input qn_in_244;
input qn_in_243;
input qn_in_242;
input q_in_241;
input qn_in_1138;
input q_in_1150;
input q_in_1041;
input q_in_1061;
input qn_in_942;
input q_in_1073;
input q_in_240;
input q_in_1148;
input q_in_1114;
input q_in_1147;
input qn_in_239;
input qn_in_1049;
input q_in_238;
input q_in_237;
input q_in_236;
input q_in_235;
input qn_in_234;
input qn_in_233;
input qn_in_232;
input qn_in_231;
input q_in_230;
input q_in_859;
input q_in_858;
input q_in_857;
input q_in_856;
input q_in_855;
input q_in_854;
input q_in_958;
input q_in_853;
input q_in_852;
input q_in_851;
input q_in_850;
input q_in_849;
input q_in_229;
input q_in_228;
input q_in_846;
input q_in_845;
input q_in_844;
input q_in_843;
input q_in_842;
input qn_in_827;
input q_in_840;
input q_in_839;
input q_in_838;
input q_in_837;
input q_in_836;
input q_in_227;
input q_in_226;
input qn_in_225;
input qn_in_224;
input q_in_223;
input qn_in_1142;
input q_in_832;
input q_in_831;
input q_in_1112;
input qn_in_830;
input qn_in_829;
input qn_in_828;
input q_in_222;
input q_in_826;
input q_in_221;
input q_in_220;
input q_in_1156;
input q_in_219;
input q_in_218;
input q_in_217;
input q_in_216;
input qn_in_215;
input qn_in_214;
input q_in_213;
input q_in_212;
input q_in_825;
input q_in_1140;
input q_in_211;
input q_in_824;
input q_in_823;
input q_in_822;
input q_in_821;
input q_in_938;
input q_in_820;
input qn_in_210;
input qn_in_818;
input q_in_979;
input q_in_209;
input q_in_816;
input qn_in_815;
input q_in_208;
input qn_in_207;
input q_in_206;
input q_in_205;
input q_in_204;
input q_in_203;
input qn_in_202;
input q_in_949;
input q_in_1111;
input q_in_1110;
input q_in_948;
input q_in_806;
input q_in_1066;
input q_in_1106;
input q_in_1105;
input q_in_1104;
input q_in_810;
input q_in_1009;
input q_in_1006;
input q_in_201;
input q_in_200;
input q_in_946;
input q_in_847;
input q_in_809;
input q_in_808;
input q_in_1101;
input qn_in_945;
input q_in_1100;
input q_in_835;
input q_in_1099;
input q_in_1098;
input q_in_1062;
input q_in_199;
input q_in_198;
input q_in_197;
input q_in_196;
input q_in_195;
input q_in_805;
input q_in_804;
input q_in_803;
input q_in_802;
input q_in_801;
input q_in_800;
input q_in_799;
input q_in_798;
input q_in_797;
input q_in_796;
input q_in_795;
input q_in_794;
input q_in_793;
input q_in_792;
input q_in_791;
input q_in_790;
input q_in_789;
input q_in_788;
input q_in_787;
input q_in_786;
input q_in_785;
input q_in_784;
input q_in_783;
input q_in_782;
input q_in_781;
input q_in_780;
input q_in_779;
input q_in_778;
input qn_in_777;
input qn_in_776;
input q_in_775;
input q_in_774;
input q_in_773;
input q_in_194;
input q_in_193;
input q_in_192;
input q_in_191;
input q_in_190;
input q_in_189;
input q_in_188;
input q_in_187;
input q_in_186;
input q_in_185;
input q_in_184;
input q_in_183;
input q_in_182;
input q_in_181;
input q_in_180;
input q_in_936;
input q_in_179;
input qn_in_819;
input q_in_934;
input q_in_768;
input q_in_767;
input qn_in_817;
input qn_in_977;
input q_in_178;
input q_in_177;
input q_in_176;
input q_in_175;
input q_in_174;
input q_in_173;
input q_in_172;
input qn_in_814;
input q_in_171;
input qn_in_813;
input qn_in_765;
input q_in_764;
input q_in_935;
input qn_in_763;
input q_in_762;
input q_in_761;
input q_in_760;
input q_in_812;
input q_in_811;
input q_in_1097;
input q_in_1096;
input q_in_1095;
input q_in_834;
input q_in_932;
input q_in_1046;
input qn_in_170;
input qn_in_169;
input q_in_758;
input q_in_757;
input q_in_756;
input q_in_755;
input q_in_754;
input q_in_753;
input q_in_752;
input q_in_751;
input q_in_750;
input q_in_694;
input q_in_168;
input q_in_748;
input q_in_747;
input q_in_746;
input q_in_745;
input q_in_744;
input q_in_167;
input q_in_166;
input q_in_165;
input q_in_164;
input q_in_163;
input q_in_162;
input q_in_161;
input q_in_160;
input q_in_159;
input q_in_736;
input q_in_735;
input q_in_734;
input q_in_158;
input q_in_1091;
input q_in_1090;
input q_in_1109;
input q_in_733;
input q_in_1108;
input q_in_848;
input q_in_1089;
input q_in_1159;
input q_in_1002;
input q_in_1103;
input q_in_157;
input q_in_156;
input q_in_155;
input q_in_154;
input qn_in_153;
input q_in_1102;
input q_in_930;
input q_in_731;
input q_in_730;
input q_in_729;
input q_in_929;
input q_in_928;
input qn_in_152;
input q_in_151;
input qn_in_927;
input q_in_150;
input q_in_149;
input q_in_148;
input q_in_728;
input q_in_1007;
input q_in_1155;
input qn_in_147;
input q_in_727;
input q_in_726;
input qn_in_725;
input q_in_1081;
input q_in_1000;
input q_in_1160;
input q_in_1059;
input q_in_724;
input q_in_833;
input qn_in_933;
input q_in_723;
input qn_in_146;
input q_in_999;
input q_in_145;
input q_in_759;
input q_in_980;
input q_in_722;
input q_in_721;
input q_in_720;
input q_in_719;
input q_in_718;
input q_in_717;
input qn_in_716;
input q_in_715;
input q_in_714;
input q_in_713;
input q_in_712;
input q_in_1094;
input q_in_998;
input q_in_711;
input q_in_1139;
input q_in_1164;
input qn_in_144;
input q_in_143;
input q_in_142;
input qn_in_141;
input qn_in_140;
input q_in_139;
input q_in_138;
input qn_in_137;
input q_in_136;
input q_in_135;
input q_in_134;
input q_in_133;
input q_in_132;
input q_in_131;
input q_in_130;
input q_in_129;
input q_in_128;
input q_in_127;
input q_in_126;
input q_in_125;
input q_in_124;
input q_in_123;
input q_in_122;
input q_in_121;
input q_in_120;
input q_in_119;
input q_in_118;
input q_in_117;
input q_in_116;
input qn_in_115;
input qn_in_114;
input qn_in_113;
input q_in_112;
input qn_in_111;
input q_in_925;
input q_in_1076;
input q_in_890;
input qn_in_707;
input qn_in_110;
input qn_in_109;
input q_in_108;
input q_in_107;
input qn_in_106;
input q_in_105;
input q_in_104;
input q_in_103;
input q_in_102;
input q_in_101;
input qn_in_100;
input q_in_99;
input q_in_98;
input qn_in_97;
input q_in_96;
input q_in_95;
input qn_in_94;
input q_in_93;
input qn_in_92;
input q_in_91;
input qn_in_90;
input q_in_89;
input qn_in_88;
input q_in_87;
input q_in_86;
input q_in_85;
input qn_in_84;
input q_in_83;
input q_in_82;
input qn_in_81;
input q_in_80;
input qn_in_79;
input q_in_78;
input qn_in_77;
input q_in_76;
input q_in_75;
input qn_in_74;
input q_in_1069;
input q_in_1088;
input q_in_1087;
input q_in_1086;
input q_in_1085;
input qn_in_73;
input q_in_72;
input qn_in_71;
input q_in_70;
input qn_in_69;
input q_in_68;
input qn_in_67;
input q_in_66;
input qn_in_65;
input q_in_64;
input qn_in_63;
input q_in_62;
input q_in_61;
input q_in_60;
input qn_in_59;
input q_in_58;
input q_in_57;
input qn_in_56;
input qn_in_55;
input qn_in_54;
input qn_in_53;
input qn_in_52;
input qn_in_51;
input q_in_702;
input q_in_701;
input q_in_700;
input q_in_699;
input q_in_698;
input q_in_697;
input q_in_696;
input qn_in_50;
input q_in_49;
input q_in_693;
input q_in_692;
input q_in_691;
input q_in_690;
input q_in_689;
input q_in_48;
input qn_in_47;
input q_in_686;
input q_in_685;
input q_in_684;
input q_in_683;
input q_in_682;
input q_in_46;
input q_in_709;
input q_in_1118;
input qn_in_45;
input q_in_44;
input qn_in_43;
input qn_in_42;
input qn_in_41;
input qn_in_40;
input q_in_39;
input q_in_38;
input qn_in_37;
input qn_in_36;
input q_in_35;
input qn_in_34;
input q_in_33;
input qn_in_32;
input qn_in_31;
input q_in_732;
input qn_in_30;
input q_in_1082;
input qn_in_29;
input q_in_28;
input q_in_27;
input qn_in_26;
input q_in_25;
input q_in_24;
input q_in_23;
input qn_in_22;
input q_in_21;
input qn_in_20;
input q_in_19;
input q_in_18;
input q_in_921;
input q_in_17;
input qn_in_16;
input qn_in_15;
input qn_in_14;
input qn_in_13;
input q_in_12;
input q_in_11;
input q_in_10;
input q_in_9;
input q_in_8;
input q_in_7;
input q_in_6;
input q_in_931;
input q_in_5;
input q_in_1152;
input q_in_916;
input q_in_4;
input q_in_3;
input q_in_915;
input q_in_913;
input q_in_1125;
input q_in_1151;
input q_in_911;
input qn_in_2;
input q_in_1;
input qn_in_952;
input qn_in_708;
input q_in_908;
input q_in_1075;
input q_in_772;
input q_in_680;
input q_in_771;
input q_in_738;
input q_in_770;
input q_in_1124;
input q_in_769;
input q_in_939;
input q_in_1176;
input q_in_974;
input q_in_1123;
input q_in_1122;
input q_in_679;
input q_in_678;
input q_in_1121;
input q_in_677;
input q_in_1168;
input q_in_676;
input qn_in_940;
input q_in_1120;
input q_in_895;
input q_in_989;
input q_in_894;
input q_in_675;
input q_in_1126;
input qn_in_674;
input q_in_893;
input q_in_673;
input q_in_1107;
input q_in_892;
input q_in_891;
input q_in_672;
input qn_in_671;
input q_in_670;
input q_in_669;
input q_in_668;
input q_in_667;
input q_in_666;
input q_in_665;
input q_in_664;
input q_in_663;
input q_in_662;
input q_in_661;
input q_in_660;
input q_in_659;
input q_in_658;
input q_in_887;
input q_in_1052;
input q_in_886;
input q_in_657;
input q_in_1174;
input q_in_1093;
input qn_in_885;
input qn_in_884;
input q_in_1051;
input q_in_883;
input q_in_656;
input q_in_1157;
input q_in_704;
input q_in_882;
input q_in_1092;
input q_in_988;
input q_in_743;
input q_in_881;
input qn_in_706;
input qn_in_880;
input q_in_655;
input q_in_654;
input q_in_653;
input q_in_652;
input q_in_1079;
input q_in_1078;
input q_in_1077;
input q_in_1047;
input q_in_705;
input q_in_742;
input q_in_1127;
input q_in_879;
input q_in_1167;
input q_in_651;
input q_in_1149;
input q_in_650;
input q_in_1045;
input q_in_741;
input q_in_878;
input q_in_1178;
input q_in_649;
input qn_in_1044;
input q_in_1175;
input q_in_648;
input q_in_877;
input q_in_740;
input q_in_876;
input q_in_875;
input qn_in_647;
input q_in_646;
input q_in_739;
input q_in_872;
input q_in_645;
input q_in_644;
input q_in_643;
input q_in_642;
input q_in_641;
input q_in_640;
input q_in_639;
input q_in_638;
input q_in_637;
input q_in_636;
input q_in_635;
input q_in_634;
input q_in_633;
input q_in_632;
input qn_in_631;
input qn_in_630;
input q_in_629;
input qn_in_628;
input q_in_627;
input q_in_626;
input q_in_625;
input q_in_624;
input q_in_1162;
input q_in_623;
input q_in_622;
input q_in_621;
input q_in_1050;
input q_in_1166;
input q_in_766;
input q_in_1117;
input q_in_1145;
input q_in_620;
input q_in_1043;
input q_in_619;
input q_in_618;
input q_in_617;
input q_in_616;
input q_in_615;
input q_in_614;
input q_in_613;
input q_in_612;
input q_in_611;
input q_in_610;
input q_in_609;
input q_in_608;
input q_in_607;
input q_in_606;
input q_in_605;
input q_in_604;
input q_in_603;
input qn_in_602;
input q_in_601;
input qn_in_600;
input q_in_1042;
input q_in_599;
input q_in_598;
input q_in_597;
input q_in_596;
input qn_in_595;
input q_in_594;
input q_in_593;
input q_in_592;
input q_in_591;
input q_in_590;
input q_in_589;
input q_in_1040;
input q_in_588;
input q_in_1039;
input q_in_986;
input q_in_1038;
input q_in_587;
input q_in_1037;
input q_in_1163;
input q_in_1036;
input q_in_1173;
input q_in_1035;
input q_in_1143;
input q_in_1034;
input q_in_1172;
input q_in_985;
input qn_in_703;
input q_in_987;
input q_in_737;
input q_in_1030;
input q_in_865;
input q_in_1029;
input q_in_1084;
input q_in_984;
input q_in_1028;
input q_in_1005;
input q_in_864;
input q_in_1158;
input q_in_1027;
input qn_in_863;
input q_in_1026;
input q_in_1001;
input q_in_1025;
input qn_in_862;
input q_in_1024;
input q_in_1171;
input q_in_983;
input q_in_1023;
input q_in_1022;
input qn_in_586;
input q_in_1021;
input qn_in_861;
input q_in_1020;
input q_in_956;
input q_in_1019;
input q_in_1170;
input q_in_1018;
input q_in_1017;
input q_in_1016;
input q_in_1015;
input q_in_710;
input q_in_1014;
input q_in_1013;
input q_in_1012;
input q_in_1011;
input q_in_1141;
input qn_in_1074;
input q_in_1010;
input q_in_1072;
input q_in_1071;
input q_in_1070;
input q_in_860;
input qn_in_585;
input q_in_584;
input q_in_1068;
input q_in_1008;
input qn_in_583;
input qn_in_582;
input q_in_1119;
input qn_in_1067;
input q_in_695;
input q_in_1065;
input q_in_1064;
input q_in_1063;
input q_in_462;
input qn_in_1048;
input q_in_982;
input q_in_1004;
input q_in_1033;
input q_in_1003;
input qn_in_581;
input q_in_1177;
input q_in_580;
input q_in_579;
input qn_in_578;
input qn_in_577;
input qn_in_576;
input qn_in_575;
input q_in_574;
input q_in_573;
input qn_in_572;
input q_in_571;
input q_in_570;
input q_in_569;
input qn_in_568;
input q_in_567;
input qn_in_566;
input q_in_565;
input q_in_981;
input q_in_688;
input q_in_564;
input q_in_1080;
input q_in_1032;
input q_in_687;
input q_in_1113;
input qn_in_1060;
input q_in_997;
input q_in_1058;
input q_in_1057;
input qn_in_1056;
input q_in_996;
input q_in_563;
input q_in_995;
input qn_in_1169;
input q_in_562;
input q_in_561;
input q_in_994;
input q_in_560;
input q_in_1031;
input q_in_993;
input q_in_1055;
input q_in_992;
input q_in_991;
input q_in_681;
input q_in_749;
input q_in_1083;
input q_in_1054;
input q_in_1053;
input q_in_990;
input q_in_559;
input qn_in_558;
input q_in_557;
input qn_in_556;
input qn_in_555;
input qn_in_554;
input qn_in_553;
input q_in_552;
input qn_in_551;
input qn_in_550;
input q_in_549;
input q_in_548;
input q_in_547;
input q_in_546;
input q_in_545;
input q_in_544;
input q_in_543;
input q_in_542;
input q_in_541;
input q_in_540;
input q_in_539;
input q_in_538;
input q_in_537;
input q_in_536;
input q_in_535;
input q_in_534;
input q_in_533;
input q_in_532;
input q_in_531;
input q_in_530;
input q_in_529;
input q_in_528;
input q_in_527;
input q_in_526;
input q_in_525;
input q_in_524;
input q_in_523;
input q_in_522;
input q_in_521;
input q_in_520;
input q_in_519;
input q_in_518;
input q_in_517;
input qn_in_516;
input q_in_515;
input q_in_514;
input q_in_513;
input q_in_512;
input q_in_511;
input q_in_510;
input q_in_509;
input q_in_508;
input q_in_507;
input q_in_506;
input q_in_505;
input q_in_504;
input q_in_503;
input q_in_502;
input q_in_501;
input q_in_500;
input q_in_499;
input q_in_498;
input q_in_497;
input q_in_496;
input q_in_495;
input q_in_494;
input q_in_493;
input q_in_492;
input q_in_491;
input q_in_490;
input q_in_489;
input q_in_488;
input q_in_487;
input q_in_486;
input q_in_485;
input q_in_484;
input q_in_483;
input q_in_482;
input q_in_481;
input q_in_480;
input q_in_479;
input q_in_478;
input q_in_477;
input q_in_476;
input q_in_475;
input q_in_474;
input q_in_473;
input q_in_472;
input q_in_471;
input qn_in_470;
input q_in_469;
input q_in_468;
input q_in_467;
input q_in_466;
input q_in_465;
input q_in_464;
input q_in_463;
input qn_in_426;
input q_in_461;
input q_in_460;
input q_in_459;
input q_in_458;
input q_in_457;
input q_in_456;
input q_in_455;
input q_in_454;
input q_in_453;
input q_in_452;
input q_in_451;
input q_in_450;
input q_in_449;
input q_in_448;
input q_in_447;
input q_in_446;
input q_in_445;
input q_in_444;
input q_in_443;
input q_in_442;
input q_in_441;
input q_in_440;
input q_in_439;
input q_in_438;
input q_in_437;
input q_in_436;
input q_in_435;
input q_in_434;
input q_in_433;
input q_in_432;
input q_in_431;
input q_in_430;
input q_in_429;
input q_in_428;
input q_in_427;
input qn_in_420;
input qn_in_425;
input qn_in_424;
input qn_in_423;
input qn_in_422;
input qn_in_421;
input blif_clk_net, blif_reset_net, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753;
input qn_in_419;
output d_out_418;
output d_out_417;
output d_out_416;
output d_out_415;
output d_out_414;
output d_out_413;
output d_out_412;
output d_out_411;
output d_out_410;
output d_out_409;
output d_out_408;
output d_out_407;
output d_out_406;
output d_out_405;
output d_out_404;
output d_out_403;
output d_out_402;
output d_out_401;
output d_out_400;
output d_out_926;
output d_out_399;
output d_out_978;
output d_out_398;
output d_out_889;
output d_out_976;
output d_out_975;
output d_out_397;
output d_out_1154;
output d_out_973;
output d_out_1153;
output d_out_972;
output d_out_396;
output d_out_395;
output d_out_969;
output d_out_968;
output d_out_1161;
output d_out_967;
output d_out_966;
output d_out_965;
output d_out_964;
output d_out_963;
output d_out_962;
output d_out_961;
output d_out_1146;
output d_out_960;
output d_out_959;
output d_out_1144;
output d_out_888;
output d_out_957;
output d_out_394;
output d_out_955;
output d_out_954;
output d_out_953;
output d_out_393;
output d_out_392;
output d_out_391;
output d_out_390;
output d_out_389;
output d_out_388;
output d_out_387;
output d_out_951;
output d_out_950;
output d_out_386;
output d_out_385;
output d_out_947;
output d_out_807;
output d_out_384;
output d_out_944;
output d_out_943;
output d_out_383;
output d_out_941;
output d_out_382;
output d_out_381;
output d_out_380;
output d_out_379;
output d_out_378;
output d_out_377;
output d_out_376;
output d_out_375;
output d_out_374;
output d_out_373;
output d_out_372;
output d_out_371;
output d_out_370;
output d_out_369;
output d_out_368;
output d_out_367;
output d_out_366;
output d_out_365;
output d_out_364;
output d_out_363;
output d_out_362;
output d_out_361;
output d_out_360;
output d_out_359;
output d_out_358;
output d_out_357;
output d_out_356;
output d_out_355;
output d_out_354;
output d_out_353;
output d_out_352;
output d_out_351;
output d_out_350;
output d_out_349;
output d_out_348;
output d_out_347;
output d_out_346;
output d_out_345;
output d_out_344;
output d_out_343;
output d_out_342;
output d_out_341;
output d_out_340;
output d_out_339;
output d_out_338;
output d_out_337;
output d_out_336;
output d_out_335;
output d_out_334;
output d_out_333;
output d_out_332;
output d_out_331;
output d_out_330;
output d_out_329;
output d_out_328;
output d_out_327;
output d_out_326;
output d_out_325;
output d_out_324;
output d_out_323;
output d_out_322;
output d_out_321;
output d_out_320;
output d_out_319;
output d_out_318;
output d_out_317;
output d_out_316;
output d_out_315;
output d_out_1137;
output d_out_1136;
output d_out_1135;
output d_out_1134;
output d_out_1133;
output d_out_1132;
output d_out_1131;
output d_out_1130;
output d_out_314;
output d_out_841;
output d_out_1129;
output d_out_1128;
output d_out_313;
output d_out_924;
output d_out_923;
output d_out_922;
output d_out_312;
output d_out_920;
output d_out_919;
output d_out_918;
output d_out_917;
output d_out_311;
output d_out_310;
output d_out_914;
output d_out_309;
output d_out_912;
output d_out_308;
output d_out_910;
output d_out_909;
output d_out_307;
output d_out_907;
output d_out_906;
output d_out_905;
output d_out_904;
output d_out_903;
output d_out_902;
output d_out_901;
output d_out_900;
output d_out_899;
output d_out_898;
output d_out_897;
output d_out_896;
output d_out_306;
output d_out_305;
output d_out_304;
output d_out_303;
output d_out_302;
output d_out_301;
output d_out_300;
output d_out_299;
output d_out_298;
output d_out_297;
output d_out_296;
output d_out_295;
output d_out_294;
output d_out_293;
output d_out_292;
output d_out_291;
output d_out_290;
output d_out_289;
output d_out_288;
output d_out_287;
output d_out_286;
output d_out_285;
output d_out_284;
output d_out_283;
output d_out_282;
output d_out_281;
output d_out_280;
output d_out_279;
output d_out_278;
output d_out_277;
output d_out_276;
output d_out_275;
output d_out_274;
output d_out_874;
output d_out_873;
output d_out_273;
output d_out_871;
output d_out_870;
output d_out_1165;
output d_out_869;
output d_out_272;
output d_out_937;
output d_out_271;
output d_out_1116;
output d_out_971;
output d_out_868;
output d_out_867;
output d_out_970;
output d_out_270;
output d_out_866;
output d_out_1115;
output d_out_269;
output d_out_268;
output d_out_267;
output d_out_266;
output d_out_265;
output d_out_264;
output d_out_263;
output d_out_262;
output d_out_261;
output d_out_260;
output d_out_259;
output d_out_258;
output d_out_257;
output d_out_256;
output d_out_255;
output d_out_254;
output d_out_253;
output d_out_252;
output d_out_251;
output d_out_250;
output d_out_249;
output d_out_248;
output d_out_247;
output d_out_246;
output d_out_245;
output d_out_244;
output d_out_243;
output d_out_242;
output d_out_241;
output d_out_1138;
output d_out_1150;
output d_out_1041;
output d_out_1061;
output d_out_942;
output d_out_1073;
output d_out_240;
output d_out_1148;
output d_out_1114;
output d_out_1147;
output d_out_239;
output d_out_1049;
output d_out_238;
output d_out_237;
output d_out_236;
output d_out_235;
output d_out_234;
output d_out_233;
output d_out_232;
output d_out_231;
output d_out_230;
output d_out_859;
output d_out_858;
output d_out_857;
output d_out_856;
output d_out_855;
output d_out_854;
output d_out_958;
output d_out_853;
output d_out_852;
output d_out_851;
output d_out_850;
output d_out_849;
output d_out_229;
output d_out_228;
output d_out_846;
output d_out_845;
output d_out_844;
output d_out_843;
output d_out_842;
output d_out_827;
output d_out_840;
output d_out_839;
output d_out_838;
output d_out_837;
output d_out_836;
output d_out_227;
output d_out_226;
output d_out_225;
output d_out_224;
output d_out_223;
output d_out_1142;
output d_out_832;
output d_out_831;
output d_out_1112;
output d_out_830;
output d_out_829;
output d_out_828;
output d_out_222;
output d_out_826;
output d_out_221;
output d_out_220;
output d_out_1156;
output d_out_219;
output d_out_218;
output d_out_217;
output d_out_216;
output d_out_215;
output d_out_214;
output d_out_213;
output d_out_212;
output d_out_825;
output d_out_1140;
output d_out_211;
output d_out_824;
output d_out_823;
output d_out_822;
output d_out_821;
output d_out_938;
output d_out_820;
output d_out_210;
output d_out_818;
output d_out_979;
output d_out_209;
output d_out_816;
output d_out_815;
output d_out_208;
output d_out_207;
output d_out_206;
output d_out_205;
output d_out_204;
output d_out_203;
output d_out_202;
output d_out_949;
output d_out_1111;
output d_out_1110;
output d_out_948;
output d_out_806;
output d_out_1066;
output d_out_1106;
output d_out_1105;
output d_out_1104;
output d_out_810;
output d_out_1009;
output d_out_1006;
output d_out_201;
output d_out_200;
output d_out_946;
output d_out_847;
output d_out_809;
output d_out_808;
output d_out_1101;
output d_out_945;
output d_out_1100;
output d_out_835;
output d_out_1099;
output d_out_1098;
output d_out_1062;
output d_out_199;
output d_out_198;
output d_out_197;
output d_out_196;
output d_out_195;
output d_out_805;
output d_out_804;
output d_out_803;
output d_out_802;
output d_out_801;
output d_out_800;
output d_out_799;
output d_out_798;
output d_out_797;
output d_out_796;
output d_out_795;
output d_out_794;
output d_out_793;
output d_out_792;
output d_out_791;
output d_out_790;
output d_out_789;
output d_out_788;
output d_out_787;
output d_out_786;
output d_out_785;
output d_out_784;
output d_out_783;
output d_out_782;
output d_out_781;
output d_out_780;
output d_out_779;
output d_out_778;
output d_out_777;
output d_out_776;
output d_out_775;
output d_out_774;
output d_out_773;
output d_out_194;
output d_out_193;
output d_out_192;
output d_out_191;
output d_out_190;
output d_out_189;
output d_out_188;
output d_out_187;
output d_out_186;
output d_out_185;
output d_out_184;
output d_out_183;
output d_out_182;
output d_out_181;
output d_out_180;
output d_out_936;
output d_out_179;
output d_out_819;
output d_out_934;
output d_out_768;
output d_out_767;
output d_out_817;
output d_out_977;
output d_out_178;
output d_out_177;
output d_out_176;
output d_out_175;
output d_out_174;
output d_out_173;
output d_out_172;
output d_out_814;
output d_out_171;
output d_out_813;
output d_out_765;
output d_out_764;
output d_out_935;
output d_out_763;
output d_out_762;
output d_out_761;
output d_out_760;
output d_out_812;
output d_out_811;
output d_out_1097;
output d_out_1096;
output d_out_1095;
output d_out_834;
output d_out_932;
output d_out_1046;
output d_out_170;
output d_out_169;
output d_out_758;
output d_out_757;
output d_out_756;
output d_out_755;
output d_out_754;
output d_out_753;
output d_out_752;
output d_out_751;
output d_out_750;
output d_out_749;
output d_out_168;
output d_out_748;
output d_out_747;
output d_out_746;
output d_out_745;
output d_out_744;
output d_out_167;
output d_out_166;
output d_out_165;
output d_out_164;
output d_out_163;
output d_out_162;
output d_out_161;
output d_out_160;
output d_out_159;
output d_out_736;
output d_out_735;
output d_out_734;
output d_out_158;
output d_out_1091;
output d_out_1090;
output d_out_1109;
output d_out_733;
output d_out_1108;
output d_out_848;
output d_out_1089;
output d_out_1159;
output d_out_1002;
output d_out_1103;
output d_out_157;
output d_out_156;
output d_out_155;
output d_out_154;
output d_out_153;
output d_out_1102;
output d_out_930;
output d_out_731;
output d_out_730;
output d_out_729;
output d_out_929;
output d_out_928;
output d_out_152;
output d_out_151;
output d_out_927;
output d_out_150;
output d_out_149;
output d_out_148;
output d_out_728;
output d_out_1007;
output d_out_1155;
output d_out_147;
output d_out_727;
output d_out_726;
output d_out_725;
output d_out_1081;
output d_out_1000;
output d_out_1160;
output d_out_1059;
output d_out_724;
output d_out_833;
output d_out_933;
output d_out_723;
output d_out_146;
output d_out_999;
output d_out_145;
output d_out_759;
output d_out_980;
output d_out_1040;
output d_out_722;
output d_out_721;
output d_out_720;
output d_out_719;
output d_out_718;
output d_out_717;
output d_out_716;
output d_out_715;
output d_out_714;
output d_out_713;
output d_out_712;
output d_out_1094;
output d_out_998;
output d_out_711;
output d_out_1139;
output d_out_1164;
output d_out_144;
output d_out_143;
output d_out_142;
output d_out_141;
output d_out_140;
output d_out_139;
output d_out_138;
output d_out_137;
output d_out_136;
output d_out_135;
output d_out_134;
output d_out_133;
output d_out_132;
output d_out_131;
output d_out_130;
output d_out_129;
output d_out_128;
output d_out_127;
output d_out_126;
output d_out_125;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_121;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_116;
output d_out_115;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_111;
output d_out_925;
output d_out_1076;
output d_out_890;
output d_out_707;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_83;
output d_out_82;
output d_out_81;
output d_out_80;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_76;
output d_out_75;
output d_out_74;
output d_out_1069;
output d_out_1088;
output d_out_1087;
output d_out_1086;
output d_out_1085;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_64;
output d_out_63;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_702;
output d_out_701;
output d_out_700;
output d_out_699;
output d_out_698;
output d_out_697;
output d_out_696;
output d_out_50;
output d_out_49;
output d_out_693;
output d_out_692;
output d_out_691;
output d_out_690;
output d_out_689;
output d_out_48;
output d_out_47;
output d_out_686;
output d_out_685;
output d_out_684;
output d_out_683;
output d_out_682;
output d_out_46;
output d_out_709;
output d_out_1118;
output d_out_45;
output d_out_44;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_732;
output d_out_30;
output d_out_1082;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_921;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_931;
output d_out_5;
output d_out_1152;
output d_out_916;
output d_out_4;
output d_out_3;
output d_out_915;
output d_out_913;
output d_out_1125;
output d_out_1151;
output d_out_911;
output d_out_2;
output d_out_1;
output d_out_952;
output d_out_708;
output d_out_908;
output d_out_1075;
output d_out_772;
output d_out_680;
output d_out_771;
output d_out_738;
output d_out_770;
output d_out_1124;
output d_out_769;
output d_out_939;
output d_out_1176;
output d_out_974;
output d_out_1123;
output d_out_1122;
output d_out_679;
output d_out_678;
output d_out_1121;
output d_out_677;
output d_out_676;
output d_out_940;
output d_out_1120;
output d_out_895;
output d_out_989;
output d_out_894;
output d_out_675;
output d_out_1126;
output d_out_674;
output d_out_893;
output d_out_673;
output d_out_1107;
output d_out_892;
output d_out_891;
output d_out_672;
output d_out_671;
output d_out_670;
output d_out_669;
output d_out_668;
output d_out_667;
output d_out_666;
output d_out_665;
output d_out_664;
output d_out_663;
output d_out_662;
output d_out_661;
output d_out_660;
output d_out_659;
output d_out_658;
output d_out_887;
output d_out_1052;
output d_out_886;
output d_out_657;
output d_out_1174;
output d_out_1093;
output d_out_885;
output d_out_884;
output d_out_1051;
output d_out_883;
output d_out_656;
output d_out_1157;
output d_out_704;
output d_out_882;
output d_out_1092;
output d_out_988;
output d_out_743;
output d_out_881;
output d_out_706;
output d_out_880;
output d_out_655;
output d_out_654;
output d_out_653;
output d_out_652;
output d_out_1079;
output d_out_1078;
output d_out_1077;
output d_out_1047;
output d_out_705;
output d_out_742;
output d_out_1127;
output d_out_879;
output d_out_1167;
output d_out_651;
output d_out_1149;
output d_out_650;
output d_out_1045;
output d_out_741;
output d_out_878;
output d_out_1178;
output d_out_649;
output d_out_1044;
output d_out_1175;
output d_out_648;
output d_out_877;
output d_out_740;
output d_out_876;
output d_out_875;
output d_out_647;
output d_out_646;
output d_out_739;
output d_out_872;
output d_out_645;
output d_out_644;
output d_out_643;
output d_out_642;
output d_out_641;
output d_out_640;
output d_out_639;
output d_out_638;
output d_out_637;
output d_out_636;
output d_out_635;
output d_out_634;
output d_out_633;
output d_out_632;
output d_out_631;
output d_out_630;
output d_out_629;
output d_out_628;
output d_out_627;
output d_out_626;
output d_out_625;
output d_out_624;
output d_out_1162;
output d_out_623;
output d_out_622;
output d_out_621;
output d_out_1050;
output d_out_1166;
output d_out_766;
output d_out_1117;
output d_out_1145;
output d_out_620;
output d_out_1043;
output d_out_619;
output d_out_618;
output d_out_617;
output d_out_616;
output d_out_615;
output d_out_614;
output d_out_613;
output d_out_612;
output d_out_611;
output d_out_610;
output d_out_609;
output d_out_608;
output d_out_607;
output d_out_606;
output d_out_605;
output d_out_604;
output d_out_603;
output d_out_602;
output d_out_601;
output d_out_600;
output d_out_1042;
output d_out_599;
output d_out_598;
output d_out_597;
output d_out_596;
output d_out_595;
output d_out_594;
output d_out_593;
output d_out_592;
output d_out_591;
output d_out_590;
output d_out_589;
output d_out_498;
output d_out_588;
output d_out_1039;
output d_out_986;
output d_out_1038;
output d_out_587;
output d_out_1037;
output d_out_1163;
output d_out_1036;
output d_out_1173;
output d_out_1035;
output d_out_1143;
output d_out_1034;
output d_out_1172;
output d_out_985;
output d_out_703;
output d_out_987;
output d_out_737;
output d_out_1030;
output d_out_865;
output d_out_1029;
output d_out_1084;
output d_out_984;
output d_out_1028;
output d_out_1005;
output d_out_864;
output d_out_1158;
output d_out_1027;
output d_out_863;
output d_out_1026;
output d_out_1001;
output d_out_1025;
output d_out_862;
output d_out_1024;
output d_out_1171;
output d_out_983;
output d_out_1023;
output d_out_1022;
output d_out_586;
output d_out_1021;
output d_out_861;
output d_out_1020;
output d_out_956;
output d_out_1019;
output d_out_1170;
output d_out_1018;
output d_out_1017;
output d_out_1016;
output d_out_1015;
output d_out_710;
output d_out_1014;
output d_out_1013;
output d_out_1012;
output d_out_1011;
output d_out_1141;
output d_out_1074;
output d_out_1010;
output d_out_1072;
output d_out_1071;
output d_out_1070;
output d_out_860;
output d_out_585;
output d_out_584;
output d_out_1068;
output d_out_1008;
output d_out_583;
output d_out_582;
output d_out_1119;
output d_out_1067;
output d_out_695;
output d_out_1065;
output d_out_1064;
output d_out_1063;
output d_out_694;
output d_out_1048;
output d_out_982;
output d_out_1004;
output d_out_1033;
output d_out_1003;
output d_out_581;
output d_out_1177;
output d_out_580;
output d_out_579;
output d_out_578;
output d_out_577;
output d_out_576;
output d_out_575;
output d_out_574;
output d_out_573;
output d_out_572;
output d_out_571;
output d_out_570;
output d_out_569;
output d_out_568;
output d_out_567;
output d_out_566;
output d_out_565;
output d_out_981;
output d_out_688;
output d_out_564;
output d_out_1080;
output d_out_1032;
output d_out_687;
output d_out_1113;
output d_out_1060;
output d_out_997;
output d_out_1058;
output d_out_1057;
output d_out_1056;
output d_out_996;
output d_out_563;
output d_out_995;
output d_out_1169;
output d_out_562;
output d_out_561;
output d_out_994;
output d_out_560;
output d_out_1031;
output d_out_993;
output d_out_1055;
output d_out_992;
output d_out_991;
output d_out_681;
output d_out_1168;
output d_out_1083;
output d_out_1054;
output d_out_1053;
output d_out_990;
output d_out_559;
output d_out_558;
output d_out_557;
output d_out_556;
output d_out_555;
output d_out_554;
output d_out_553;
output d_out_552;
output d_out_551;
output d_out_550;
output d_out_549;
output d_out_548;
output d_out_547;
output d_out_546;
output d_out_545;
output d_out_544;
output d_out_543;
output d_out_542;
output d_out_541;
output d_out_540;
output d_out_539;
output d_out_538;
output d_out_537;
output d_out_536;
output d_out_535;
output d_out_534;
output d_out_533;
output d_out_532;
output d_out_531;
output d_out_530;
output d_out_529;
output d_out_528;
output d_out_527;
output d_out_526;
output d_out_525;
output d_out_524;
output d_out_523;
output d_out_522;
output d_out_521;
output d_out_520;
output d_out_519;
output d_out_518;
output d_out_517;
output d_out_516;
output d_out_515;
output d_out_514;
output d_out_513;
output d_out_512;
output d_out_511;
output d_out_510;
output d_out_509;
output d_out_508;
output d_out_507;
output d_out_506;
output d_out_505;
output d_out_504;
output d_out_503;
output d_out_502;
output d_out_501;
output d_out_500;
output d_out_499;
output d_out_432;
output d_out_497;
output d_out_496;
output d_out_495;
output d_out_494;
output d_out_493;
output d_out_492;
output d_out_491;
output d_out_490;
output d_out_489;
output d_out_488;
output d_out_487;
output d_out_486;
output d_out_485;
output d_out_484;
output d_out_483;
output d_out_482;
output d_out_481;
output d_out_480;
output d_out_479;
output d_out_478;
output d_out_477;
output d_out_476;
output d_out_475;
output d_out_474;
output d_out_473;
output d_out_472;
output d_out_471;
output d_out_470;
output d_out_469;
output d_out_468;
output d_out_467;
output d_out_466;
output d_out_465;
output d_out_464;
output d_out_463;
output d_out_462;
output d_out_461;
output d_out_460;
output d_out_459;
output d_out_458;
output d_out_457;
output d_out_456;
output d_out_455;
output d_out_454;
output d_out_453;
output d_out_452;
output d_out_451;
output d_out_450;
output d_out_449;
output d_out_448;
output d_out_447;
output d_out_446;
output d_out_445;
output d_out_444;
output d_out_443;
output d_out_442;
output d_out_441;
output d_out_440;
output d_out_439;
output d_out_438;
output d_out_437;
output d_out_436;
output d_out_435;
output d_out_434;
output d_out_433;
output d_out_421;
output d_out_431;
output d_out_430;
output d_out_429;
output d_out_428;
output d_out_427;
output d_out_426;
output d_out_425;
output d_out_424;
output d_out_423;
output d_out_422;
output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972;
output d_out_420;
output d_out_419;
wire n_11211, n_11212, n_11216, n_11217, n_11218, n_11219, n_11220, n_11221;
wire n_11201, n_11203, n_11205, n_11206, n_11207, n_11208, n_11209, n_11210;
wire n_11191, n_11192, n_11193, n_11194, n_11195, n_11196, n_11197, n_11198;
wire n_11178, n_11184, n_11185, n_11186, n_11187, n_11188, n_11189, n_11190;
wire n_11157, n_11160, n_11162, n_11163, n_11165, n_11171, n_11173, n_11177;
wire n_11124, n_11126, n_11128, n_11129, n_11133, n_11134, n_11138, n_11150;
wire n_11110, n_11113, n_11116, n_11118, n_11119, n_11120, n_11121, n_11122;
wire n_11094, n_11095, n_11097, n_11099, n_11101, n_11104, n_11105, n_11106;
wire n_11073, n_11076, n_11077, n_11079, n_11080, n_11081, n_11088, n_11091;
wire n_11050, n_11051, n_11055, n_11056, n_11064, n_11065, n_11070, n_11071;
wire n_11036, n_11037, n_11038, n_11039, n_11040, n_11041, n_11042, n_11045;
wire n_11028, n_11029, n_11030, n_11031, n_11032, n_11033, n_11034, n_11035;
wire n_10996, n_10997, n_10998, n_11012, n_11013, n_11025, n_11026, n_11027;
wire n_10987, n_10988, n_10989, n_10991, n_10992, n_10993, n_10994, n_10995;
wire n_10976, n_10978, n_10980, n_10981, n_10982, n_10983, n_10984, n_10986;
wire n_10968, n_10969, n_10970, n_10971, n_10972, n_10973, n_10974, n_10975;
wire n_10960, n_10961, n_10962, n_10963, n_10964, n_10965, n_10966, n_10967;
wire n_10950, n_10951, n_10952, n_10953, n_10954, n_10955, n_10956, n_10959;
wire n_10940, n_10941, n_10942, n_10943, n_10944, n_10947, n_10948, n_10949;
wire n_10917, n_10920, n_10921, n_10932, n_10934, n_10936, n_10937, n_10939;
wire n_10906, n_10907, n_10910, n_10911, n_10912, n_10913, n_10915, n_10916;
wire n_10894, n_10895, n_10897, n_10898, n_10899, n_10901, n_10903, n_10905;
wire n_10871, n_10873, n_10874, n_10877, n_10879, n_10883, n_10889, n_10893;
wire n_10852, n_10853, n_10854, n_10856, n_10857, n_10861, n_10863, n_10867;
wire n_10829, n_10830, n_10831, n_10833, n_10834, n_10839, n_10841, n_10846;
wire n_10808, n_10809, n_10813, n_10814, n_10818, n_10823, n_10826, n_10827;
wire n_10789, n_10790, n_10801, n_10802, n_10803, n_10804, n_10805, n_10806;
wire n_10770, n_10771, n_10772, n_10773, n_10781, n_10782, n_10785, n_10787;
wire n_10762, n_10763, n_10764, n_10765, n_10766, n_10767, n_10768, n_10769;
wire n_10753, n_10754, n_10755, n_10756, n_10758, n_10759, n_10760, n_10761;
wire n_10745, n_10746, n_10747, n_10748, n_10749, n_10750, n_10751, n_10752;
wire n_10715, n_10716, n_10717, n_10718, n_10720, n_10723, n_10724, n_10725;
wire n_10698, n_10699, n_10700, n_10708, n_10709, n_10710, n_10713, n_10714;
wire n_10687, n_10689, n_10690, n_10693, n_10694, n_10695, n_10696, n_10697;
wire n_10674, n_10675, n_10678, n_10682, n_10683, n_10684, n_10685, n_10686;
wire n_10657, n_10660, n_10664, n_10667, n_10669, n_10670, n_10671, n_10672;
wire n_10637, n_10638, n_10639, n_10644, n_10647, n_10649, n_10650, n_10656;
wire n_10625, n_10626, n_10628, n_10630, n_10631, n_10632, n_10633, n_10634;
wire n_10616, n_10617, n_10618, n_10620, n_10621, n_10622, n_10623, n_10624;
wire n_10598, n_10599, n_10600, n_10601, n_10607, n_10609, n_10613, n_10614;
wire n_10582, n_10587, n_10588, n_10589, n_10590, n_10595, n_10596, n_10597;
wire n_10569, n_10573, n_10576, n_10577, n_10578, n_10579, n_10580, n_10581;
wire n_10558, n_10560, n_10563, n_10564, n_10565, n_10566, n_10567, n_10568;
wire n_10548, n_10549, n_10550, n_10551, n_10552, n_10553, n_10554, n_10557;
wire n_10525, n_10526, n_10527, n_10528, n_10529, n_10532, n_10534, n_10535;
wire n_10515, n_10516, n_10517, n_10518, n_10519, n_10520, n_10522, n_10524;
wire n_10503, n_10504, n_10505, n_10506, n_10508, n_10512, n_10513, n_10514;
wire n_10470, n_10472, n_10473, n_10475, n_10494, n_10495, n_10496, n_10499;
wire n_10448, n_10460, n_10461, n_10462, n_10463, n_10464, n_10466, n_10467;
wire n_10429, n_10430, n_10431, n_10443, n_10444, n_10445, n_10446, n_10447;
wire n_10416, n_10422, n_10423, n_10424, n_10425, n_10426, n_10427, n_10428;
wire n_10401, n_10402, n_10404, n_10411, n_10412, n_10413, n_10414, n_10415;
wire n_10392, n_10394, n_10395, n_10396, n_10397, n_10398, n_10399, n_10400;
wire n_10382, n_10383, n_10385, n_10386, n_10387, n_10388, n_10390, n_10391;
wire n_10373, n_10374, n_10376, n_10377, n_10378, n_10379, n_10380, n_10381;
wire n_10357, n_10361, n_10362, n_10363, n_10368, n_10369, n_10371, n_10372;
wire n_10330, n_10341, n_10342, n_10343, n_10344, n_10345, n_10346, n_10347;
wire n_10320, n_10321, n_10322, n_10323, n_10325, n_10327, n_10328, n_10329;
wire n_10312, n_10313, n_10314, n_10315, n_10316, n_10317, n_10318, n_10319;
wire n_10303, n_10304, n_10306, n_10307, n_10308, n_10309, n_10310, n_10311;
wire n_10283, n_10285, n_10286, n_10287, n_10288, n_10289, n_10290, n_10296;
wire n_10263, n_10264, n_10268, n_10270, n_10271, n_10280, n_10281, n_10282;
wire n_10243, n_10245, n_10247, n_10257, n_10259, n_10260, n_10261, n_10262;
wire n_10227, n_10228, n_10229, n_10238, n_10239, n_10240, n_10241, n_10242;
wire n_10206, n_10213, n_10214, n_10216, n_10217, n_10224, n_10225, n_10226;
wire n_10196, n_10197, n_10199, n_10200, n_10201, n_10202, n_10203, n_10205;
wire n_10176, n_10177, n_10180, n_10181, n_10184, n_10185, n_10188, n_10192;
wire n_10125, n_10128, n_10129, n_10134, n_10139, n_10142, n_10173, n_10175;
wire n_10107, n_10108, n_10112, n_10113, n_10115, n_10119, n_10120, n_10123;
wire n_10013, n_10063, n_10078, n_10097, n_10099, n_10100, n_10101, n_10103;
wire n_9903, n_9928, n_9940, n_9952, n_9976, n_9978, n_9992, n_10005;
wire n_9836, n_9856, n_9862, n_9871, n_9874, n_9883, n_9884, n_9894;
wire n_9717, n_9750, n_9772, n_9775, n_9797, n_9811, n_9830, n_9834;
wire n_9630, n_9651, n_9664, n_9672, n_9681, n_9693, n_9697, n_9698;
wire n_9505, n_9521, n_9526, n_9553, n_9558, n_9599, n_9627, n_9628;
wire n_9453, n_9454, n_9461, n_9466, n_9469, n_9491, n_9493, n_9501;
wire n_9398, n_9404, n_9419, n_9422, n_9425, n_9431, n_9443, n_9448;
wire n_9300, n_9311, n_9333, n_9351, n_9353, n_9358, n_9359, n_9371;
wire n_9209, n_9218, n_9234, n_9240, n_9256, n_9269, n_9279, n_9297;
wire n_9129, n_9139, n_9141, n_9156, n_9167, n_9172, n_9176, n_9193;
wire n_8915, n_8917, n_8921, n_8955, n_9000, n_9019, n_9091, n_9107;
wire n_8885, n_8886, n_8895, n_8898, n_8906, n_8908, n_8909, n_8913;
wire n_8848, n_8850, n_8855, n_8864, n_8879, n_8880, n_8882, n_8883;
wire n_8833, n_8834, n_8835, n_8836, n_8837, n_8839, n_8840, n_8846;
wire n_8816, n_8817, n_8818, n_8819, n_8820, n_8821, n_8831, n_8832;
wire n_8793, n_8796, n_8799, n_8800, n_8806, n_8807, n_8809, n_8810;
wire n_8764, n_8768, n_8769, n_8770, n_8776, n_8777, n_8778, n_8792;
wire n_8755, n_8756, n_8757, n_8758, n_8759, n_8761, n_8762, n_8763;
wire n_8706, n_8707, n_8730, n_8731, n_8733, n_8734, n_8735, n_8736;
wire n_8691, n_8693, n_8694, n_8697, n_8702, n_8703, n_8704, n_8705;
wire n_8678, n_8679, n_8680, n_8681, n_8682, n_8686, n_8687, n_8690;
wire n_8633, n_8634, n_8637, n_8638, n_8639, n_8675, n_8676, n_8677;
wire n_8616, n_8618, n_8619, n_8620, n_8627, n_8628, n_8629, n_8632;
wire n_8601, n_8603, n_8604, n_8605, n_8609, n_8610, n_8611, n_8615;
wire n_8586, n_8587, n_8588, n_8589, n_8591, n_8594, n_8599, n_8600;
wire n_8556, n_8557, n_8571, n_8572, n_8582, n_8583, n_8584, n_8585;
wire n_8534, n_8537, n_8540, n_8546, n_8547, n_8548, n_8552, n_8555;
wire n_7353, n_7354, n_7383, n_7395, n_7402, n_8508, n_8509, n_8532;
wire n_7330, n_7331, n_7332, n_7333, n_7343, n_7344, n_7348, n_7352;
wire n_7322, n_7323, n_7324, n_7325, n_7326, n_7327, n_7328, n_7329;
wire n_7243, n_7245, n_7247, n_7260, n_7268, n_7275, n_7320, n_7321;
wire n_7213, n_7214, n_7217, n_7218, n_7219, n_7229, n_7235, n_7242;
wire n_7145, n_7146, n_7150, n_7164, n_7165, n_7167, n_7168, n_7208;
wire n_7131, n_7132, n_7133, n_7140, n_7141, n_7142, n_7143, n_7144;
wire n_7120, n_7121, n_7122, n_7123, n_7124, n_7127, n_7128, n_7130;
wire n_7099, n_7101, n_7102, n_7103, n_7105, n_7116, n_7118, n_7119;
wire n_7086, n_7087, n_7088, n_7089, n_7090, n_7093, n_7094, n_7097;
wire n_7043, n_7044, n_7045, n_7046, n_7047, n_7048, n_7049, n_7085;
wire n_7022, n_7023, n_7024, n_7025, n_7032, n_7039, n_7040, n_7042;
wire n_6972, n_6973, n_6978, n_6979, n_7003, n_7004, n_7010, n_7018;
wire n_6948, n_6951, n_6953, n_6954, n_6956, n_6958, n_6967, n_6970;
wire n_6925, n_6926, n_6927, n_6928, n_6937, n_6938, n_6940, n_6941;
wire n_6897, n_6898, n_6899, n_6903, n_6906, n_6907, n_6922, n_6923;
wire n_6877, n_6878, n_6880, n_6891, n_6892, n_6893, n_6895, n_6896;
wire n_6856, n_6857, n_6858, n_6864, n_6865, n_6866, n_6872, n_6876;
wire n_6823, n_6848, n_6849, n_6850, n_6851, n_6852, n_6853, n_6854;
wire n_6800, n_6801, n_6806, n_6807, n_6808, n_6809, n_6821, n_6822;
wire n_6788, n_6789, n_6790, n_6791, n_6794, n_6796, n_6798, n_6799;
wire n_6765, n_6766, n_6767, n_6781, n_6782, n_6785, n_6786, n_6787;
wire n_6755, n_6756, n_6757, n_6758, n_6759, n_6760, n_6762, n_6764;
wire n_6715, n_6716, n_6734, n_6735, n_6742, n_6746, n_6752, n_6754;
wire n_6693, n_6694, n_6695, n_6696, n_6697, n_6705, n_6707, n_6714;
wire n_6684, n_6685, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692;
wire n_6669, n_6670, n_6673, n_6676, n_6677, n_6679, n_6680, n_6683;
wire n_6621, n_6631, n_6639, n_6655, n_6663, n_6664, n_6666, n_6668;
wire n_6577, n_6578, n_6582, n_6584, n_6610, n_6612, n_6618, n_6620;
wire n_6552, n_6553, n_6562, n_6564, n_6565, n_6570, n_6572, n_6574;
wire n_6524, n_6527, n_6539, n_6545, n_6547, n_6548, n_6549, n_6551;
wire n_6503, n_6504, n_6506, n_6507, n_6508, n_6517, n_6522, n_6523;
wire n_6457, n_6460, n_6464, n_6468, n_6479, n_6488, n_6490, n_6501;
wire n_6415, n_6416, n_6417, n_6418, n_6419, n_6421, n_6422, n_6454;
wire n_6407, n_6408, n_6409, n_6410, n_6411, n_6412, n_6413, n_6414;
wire n_6399, n_6400, n_6401, n_6402, n_6403, n_6404, n_6405, n_6406;
wire n_6390, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397, n_6398;
wire n_6381, n_6382, n_6383, n_6384, n_6385, n_6386, n_6388, n_6389;
wire n_6372, n_6373, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380;
wire n_6364, n_6365, n_6366, n_6367, n_6368, n_6369, n_6370, n_6371;
wire n_6355, n_6356, n_6357, n_6359, n_6360, n_6361, n_6362, n_6363;
wire n_6342, n_6345, n_6346, n_6347, n_6348, n_6351, n_6352, n_6353;
wire n_6331, n_6332, n_6334, n_6335, n_6336, n_6337, n_6338, n_6339;
wire n_6320, n_6321, n_6323, n_6324, n_6326, n_6327, n_6328, n_6330;
wire n_6310, n_6311, n_6312, n_6313, n_6315, n_6316, n_6317, n_6318;
wire n_6301, n_6302, n_6303, n_6304, n_6305, n_6306, n_6308, n_6309;
wire n_6288, n_6290, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300;
wire n_6279, n_6280, n_6281, n_6282, n_6283, n_6285, n_6286, n_6287;
wire n_6262, n_6264, n_6265, n_6266, n_6267, n_6271, n_6274, n_6275;
wire n_6253, n_6254, n_6255, n_6256, n_6257, n_6258, n_6259, n_6260;
wire n_6240, n_6241, n_6243, n_6246, n_6247, n_6248, n_6250, n_6252;
wire n_6232, n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239;
wire n_6222, n_6223, n_6224, n_6225, n_6226, n_6228, n_6229, n_6230;
wire n_6210, n_6211, n_6214, n_6216, n_6217, n_6218, n_6220, n_6221;
wire n_6201, n_6202, n_6203, n_6204, n_6206, n_6207, n_6208, n_6209;
wire n_6188, n_6189, n_6190, n_6192, n_6194, n_6197, n_6198, n_6199;
wire n_6176, n_6178, n_6180, n_6182, n_6183, n_6184, n_6185, n_6186;
wire n_6164, n_6165, n_6166, n_6167, n_6168, n_6169, n_6171, n_6174;
wire n_6153, n_6154, n_6155, n_6156, n_6157, n_6160, n_6161, n_6162;
wire n_6140, n_6141, n_6142, n_6143, n_6145, n_6146, n_6149, n_6150;
wire n_6129, n_6130, n_6132, n_6133, n_6134, n_6136, n_6137, n_6138;
wire n_6117, n_6118, n_6120, n_6121, n_6123, n_6125, n_6126, n_6128;
wire n_6107, n_6108, n_6109, n_6110, n_6111, n_6112, n_6114, n_6116;
wire n_6096, n_6098, n_6100, n_6101, n_6102, n_6103, n_6104, n_6105;
wire n_6086, n_6087, n_6089, n_6091, n_6092, n_6093, n_6094, n_6095;
wire n_6074, n_6076, n_6078, n_6079, n_6080, n_6081, n_6082, n_6084;
wire n_6065, n_6066, n_6067, n_6068, n_6070, n_6071, n_6072, n_6073;
wire n_6055, n_6057, n_6058, n_6059, n_6060, n_6061, n_6062, n_6064;
wire n_6045, n_6046, n_6048, n_6049, n_6050, n_6051, n_6052, n_6054;
wire n_6037, n_6038, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044;
wire n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035, n_6036;
wire n_6019, n_6020, n_6021, n_6024, n_6025, n_6026, n_6027, n_6028;
wire n_6011, n_6012, n_6013, n_6014, n_6015, n_6016, n_6017, n_6018;
wire n_6002, n_6003, n_6004, n_6005, n_6006, n_6008, n_6009, n_6010;
wire n_5993, n_5994, n_5995, n_5996, n_5997, n_5999, n_6000, n_6001;
wire n_5982, n_5983, n_5984, n_5985, n_5986, n_5988, n_5991, n_5992;
wire n_5973, n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5981;
wire n_5964, n_5965, n_5967, n_5968, n_5969, n_5970, n_5971, n_5972;
wire n_5954, n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962;
wire n_5945, n_5947, n_5948, n_5949, n_5950, n_5951, n_5952, n_5953;
wire n_5936, n_5937, n_5939, n_5940, n_5941, n_5942, n_5943, n_5944;
wire n_5928, n_5929, n_5930, n_5931, n_5932, n_5933, n_5934, n_5935;
wire n_5918, n_5920, n_5921, n_5922, n_5924, n_5925, n_5926, n_5927;
wire n_5907, n_5908, n_5909, n_5910, n_5913, n_5914, n_5916, n_5917;
wire n_5889, n_5891, n_5896, n_5899, n_5901, n_5904, n_5905, n_5906;
wire n_5881, n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888;
wire n_5873, n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880;
wire n_5863, n_5865, n_5866, n_5868, n_5869, n_5870, n_5871, n_5872;
wire n_5844, n_5849, n_5852, n_5854, n_5857, n_5859, n_5860, n_5862;
wire n_5824, n_5825, n_5828, n_5830, n_5831, n_5833, n_5837, n_5839;
wire n_5815, n_5816, n_5817, n_5818, n_5819, n_5820, n_5821, n_5822;
wire n_5806, n_5807, n_5808, n_5809, n_5810, n_5811, n_5813, n_5814;
wire n_5797, n_5798, n_5799, n_5800, n_5801, n_5803, n_5804, n_5805;
wire n_5784, n_5786, n_5788, n_5790, n_5792, n_5794, n_5795, n_5796;
wire n_5774, n_5775, n_5776, n_5777, n_5779, n_5780, n_5781, n_5782;
wire n_5760, n_5761, n_5762, n_5765, n_5767, n_5768, n_5769, n_5772;
wire n_5745, n_5746, n_5749, n_5755, n_5756, n_5757, n_5758, n_5759;
wire n_5736, n_5737, n_5738, n_5740, n_5741, n_5742, n_5743, n_5744;
wire n_5728, n_5729, n_5730, n_5731, n_5732, n_5733, n_5734, n_5735;
wire n_5718, n_5719, n_5720, n_5723, n_5724, n_5725, n_5726, n_5727;
wire n_5705, n_5707, n_5709, n_5711, n_5712, n_5714, n_5715, n_5716;
wire n_5693, n_5694, n_5695, n_5700, n_5701, n_5702, n_5703, n_5704;
wire n_5680, n_5681, n_5683, n_5686, n_5688, n_5689, n_5690, n_5692;
wire n_5669, n_5671, n_5672, n_5674, n_5675, n_5676, n_5677, n_5678;
wire n_5661, n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668;
wire n_5652, n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660;
wire n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646, n_5650;
wire n_5627, n_5629, n_5630, n_5631, n_5633, n_5634, n_5637, n_5639;
wire n_5614, n_5615, n_5617, n_5619, n_5622, n_5624, n_5625, n_5626;
wire n_5602, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613;
wire n_5587, n_5590, n_5591, n_5592, n_5593, n_5596, n_5599, n_5600;
wire n_5576, n_5578, n_5579, n_5580, n_5581, n_5582, n_5583, n_5584;
wire n_5567, n_5568, n_5569, n_5570, n_5571, n_5573, n_5574, n_5575;
wire n_5557, n_5559, n_5560, n_5562, n_5563, n_5564, n_5565, n_5566;
wire n_5541, n_5542, n_5543, n_5544, n_5547, n_5549, n_5553, n_5556;
wire n_5531, n_5532, n_5534, n_5536, n_5537, n_5538, n_5539, n_5540;
wire n_5520, n_5521, n_5522, n_5524, n_5526, n_5527, n_5529, n_5530;
wire n_5506, n_5508, n_5513, n_5514, n_5515, n_5517, n_5518, n_5519;
wire n_5495, n_5497, n_5499, n_5500, n_5501, n_5502, n_5504, n_5505;
wire n_5481, n_5483, n_5485, n_5486, n_5487, n_5489, n_5490, n_5492;
wire n_5464, n_5465, n_5466, n_5467, n_5468, n_5471, n_5474, n_5476;
wire n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462;
wire n_5445, n_5447, n_5448, n_5449, n_5450, n_5451, n_5453, n_5454;
wire n_5430, n_5431, n_5432, n_5436, n_5437, n_5440, n_5442, n_5444;
wire n_5414, n_5415, n_5420, n_5422, n_5423, n_5424, n_5425, n_5428;
wire n_5405, n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412;
wire n_5395, n_5396, n_5397, n_5398, n_5400, n_5402, n_5403, n_5404;
wire n_5385, n_5386, n_5387, n_5388, n_5391, n_5392, n_5393, n_5394;
wire n_5375, n_5377, n_5378, n_5379, n_5380, n_5382, n_5383, n_5384;
wire n_5363, n_5364, n_5365, n_5369, n_5370, n_5372, n_5373, n_5374;
wire n_5354, n_5355, n_5356, n_5357, n_5358, n_5359, n_5361, n_5362;
wire n_5345, n_5346, n_5347, n_5348, n_5349, n_5350, n_5352, n_5353;
wire n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342, n_5344;
wire n_5326, n_5327, n_5328, n_5329, n_5330, n_5331, n_5333, n_5335;
wire n_5315, n_5317, n_5318, n_5319, n_5321, n_5323, n_5324, n_5325;
wire n_5306, n_5307, n_5308, n_5309, n_5310, n_5311, n_5312, n_5313;
wire n_5293, n_5294, n_5296, n_5297, n_5299, n_5300, n_5302, n_5304;
wire n_5282, n_5283, n_5284, n_5287, n_5288, n_5289, n_5290, n_5291;
wire n_5270, n_5271, n_5272, n_5273, n_5275, n_5276, n_5278, n_5279;
wire n_5253, n_5254, n_5258, n_5259, n_5265, n_5266, n_5267, n_5268;
wire n_5244, n_5245, n_5246, n_5247, n_5248, n_5249, n_5251, n_5252;
wire n_5233, n_5235, n_5236, n_5238, n_5239, n_5240, n_5241, n_5242;
wire n_5224, n_5225, n_5226, n_5227, n_5229, n_5230, n_5231, n_5232;
wire n_5213, n_5214, n_5215, n_5218, n_5219, n_5221, n_5222, n_5223;
wire n_5202, n_5204, n_5205, n_5206, n_5207, n_5209, n_5210, n_5212;
wire n_5190, n_5192, n_5193, n_5195, n_5197, n_5199, n_5200, n_5201;
wire n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5189;
wire n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5177, n_5179;
wire n_5159, n_5160, n_5161, n_5163, n_5164, n_5165, n_5167, n_5168;
wire n_5149, n_5150, n_5151, n_5152, n_5154, n_5155, n_5156, n_5158;
wire n_5136, n_5137, n_5139, n_5141, n_5143, n_5144, n_5146, n_5148;
wire n_5127, n_5128, n_5129, n_5130, n_5131, n_5133, n_5134, n_5135;
wire n_5118, n_5119, n_5121, n_5122, n_5123, n_5124, n_5125, n_5126;
wire n_5107, n_5109, n_5110, n_5111, n_5112, n_5113, n_5115, n_5116;
wire n_5095, n_5097, n_5098, n_5100, n_5101, n_5103, n_5104, n_5106;
wire n_5086, n_5087, n_5088, n_5090, n_5091, n_5092, n_5093, n_5094;
wire n_5076, n_5077, n_5079, n_5081, n_5082, n_5083, n_5084, n_5085;
wire n_5065, n_5067, n_5068, n_5069, n_5071, n_5072, n_5073, n_5075;
wire n_5056, n_5057, n_5058, n_5059, n_5060, n_5062, n_5063, n_5064;
wire n_5046, n_5047, n_5048, n_5050, n_5051, n_5052, n_5053, n_5055;
wire n_5038, n_5039, n_5040, n_5041, n_5042, n_5043, n_5044, n_5045;
wire n_5028, n_5029, n_5030, n_5032, n_5033, n_5034, n_5035, n_5037;
wire n_5019, n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026;
wire n_5009, n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018;
wire n_5001, n_5002, n_5003, n_5004, n_5005, n_5006, n_5007, n_5008;
wire n_4986, n_4987, n_4988, n_4990, n_4991, n_4996, n_4999, n_5000;
wire n_4978, n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985;
wire n_4969, n_4970, n_4971, n_4972, n_4974, n_4975, n_4976, n_4977;
wire n_4961, n_4962, n_4963, n_4964, n_4965, n_4966, n_4967, n_4968;
wire n_4952, n_4953, n_4954, n_4955, n_4956, n_4957, n_4959, n_4960;
wire n_4944, n_4945, n_4946, n_4947, n_4948, n_4949, n_4950, n_4951;
wire n_4931, n_4934, n_4935, n_4936, n_4939, n_4940, n_4942, n_4943;
wire n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930;
wire n_4913, n_4915, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922;
wire n_4899, n_4900, n_4904, n_4905, n_4906, n_4907, n_4911, n_4912;
wire n_4887, n_4888, n_4889, n_4891, n_4893, n_4896, n_4897, n_4898;
wire n_4876, n_4877, n_4878, n_4879, n_4881, n_4884, n_4885, n_4886;
wire n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4874, n_4875;
wire n_4854, n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4864;
wire n_4845, n_4846, n_4847, n_4849, n_4850, n_4851, n_4852, n_4853;
wire n_4836, n_4838, n_4839, n_4840, n_4841, n_4842, n_4843, n_4844;
wire n_4827, n_4828, n_4829, n_4830, n_4832, n_4833, n_4834, n_4835;
wire n_4812, n_4813, n_4815, n_4820, n_4821, n_4822, n_4823, n_4824;
wire n_4800, n_4803, n_4804, n_4805, n_4806, n_4809, n_4810, n_4811;
wire n_4791, n_4792, n_4794, n_4795, n_4796, n_4797, n_4798, n_4799;
wire n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790;
wire n_4774, n_4775, n_4776, n_4777, n_4779, n_4780, n_4781, n_4782;
wire n_4765, n_4766, n_4767, n_4768, n_4769, n_4770, n_4772, n_4773;
wire n_4757, n_4758, n_4759, n_4760, n_4761, n_4762, n_4763, n_4764;
wire n_4747, n_4750, n_4751, n_4752, n_4753, n_4754, n_4755, n_4756;
wire n_4738, n_4739, n_4740, n_4741, n_4742, n_4743, n_4744, n_4746;
wire n_4727, n_4730, n_4731, n_4732, n_4734, n_4735, n_4736, n_4737;
wire n_4715, n_4716, n_4717, n_4719, n_4721, n_4723, n_4725, n_4726;
wire n_4707, n_4708, n_4709, n_4710, n_4711, n_4712, n_4713, n_4714;
wire n_4690, n_4693, n_4695, n_4699, n_4700, n_4704, n_4705, n_4706;
wire n_4678, n_4679, n_4680, n_4682, n_4683, n_4684, n_4688, n_4689;
wire n_4668, n_4669, n_4670, n_4671, n_4672, n_4673, n_4676, n_4677;
wire n_4659, n_4660, n_4661, n_4662, n_4663, n_4665, n_4666, n_4667;
wire n_4651, n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658;
wire n_4638, n_4639, n_4640, n_4642, n_4645, n_4647, n_4649, n_4650;
wire n_4629, n_4630, n_4631, n_4632, n_4633, n_4634, n_4636, n_4637;
wire n_4621, n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628;
wire n_4611, n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620;
wire n_4593, n_4594, n_4597, n_4598, n_4600, n_4603, n_4605, n_4607;
wire n_4584, n_4585, n_4586, n_4587, n_4589, n_4590, n_4591, n_4592;
wire n_4575, n_4576, n_4577, n_4578, n_4579, n_4581, n_4582, n_4583;
wire n_4566, n_4567, n_4568, n_4569, n_4570, n_4572, n_4573, n_4574;
wire n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565;
wire n_4546, n_4547, n_4550, n_4553, n_4554, n_4555, n_4556, n_4557;
wire n_4535, n_4537, n_4538, n_4539, n_4540, n_4541, n_4542, n_4545;
wire n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533, n_4534;
wire n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525, n_4526;
wire n_4508, n_4510, n_4512, n_4513, n_4514, n_4515, n_4516, n_4518;
wire n_4499, n_4500, n_4501, n_4502, n_4503, n_4504, n_4506, n_4507;
wire n_4490, n_4492, n_4493, n_4494, n_4495, n_4496, n_4497, n_4498;
wire n_4481, n_4482, n_4483, n_4485, n_4486, n_4487, n_4488, n_4489;
wire n_4471, n_4472, n_4473, n_4474, n_4475, n_4477, n_4478, n_4479;
wire n_4462, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470;
wire n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461;
wire n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453;
wire n_4437, n_4438, n_4439, n_4440, n_4441, n_4442, n_4444, n_4445;
wire n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4434, n_4436;
wire n_4420, n_4421, n_4422, n_4423, n_4424, n_4425, n_4426, n_4427;
wire n_4412, n_4413, n_4414, n_4415, n_4416, n_4417, n_4418, n_4419;
wire n_4404, n_4405, n_4406, n_4407, n_4408, n_4409, n_4410, n_4411;
wire n_4396, n_4397, n_4398, n_4399, n_4400, n_4401, n_4402, n_4403;
wire n_4388, n_4389, n_4390, n_4391, n_4392, n_4393, n_4394, n_4395;
wire n_4380, n_4381, n_4382, n_4383, n_4384, n_4385, n_4386, n_4387;
wire n_4372, n_4373, n_4374, n_4375, n_4376, n_4377, n_4378, n_4379;
wire n_4364, n_4365, n_4366, n_4367, n_4368, n_4369, n_4370, n_4371;
wire n_4356, n_4357, n_4358, n_4359, n_4360, n_4361, n_4362, n_4363;
wire n_4348, n_4349, n_4350, n_4351, n_4352, n_4353, n_4354, n_4355;
wire n_4338, n_4339, n_4340, n_4343, n_4344, n_4345, n_4346, n_4347;
wire n_4325, n_4327, n_4328, n_4329, n_4330, n_4331, n_4333, n_4336;
wire n_4317, n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324;
wire n_4304, n_4305, n_4306, n_4308, n_4313, n_4314, n_4315, n_4316;
wire n_4293, n_4296, n_4297, n_4298, n_4299, n_4301, n_4302, n_4303;
wire n_4282, n_4283, n_4284, n_4285, n_4286, n_4288, n_4290, n_4291;
wire n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281;
wire n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273;
wire n_4254, n_4255, n_4257, n_4260, n_4262, n_4263, n_4264, n_4265;
wire n_4243, n_4246, n_4247, n_4248, n_4250, n_4251, n_4252, n_4253;
wire n_4232, n_4233, n_4235, n_4237, n_4238, n_4239, n_4241, n_4242;
wire n_4221, n_4223, n_4224, n_4225, n_4226, n_4227, n_4230, n_4231;
wire n_4213, n_4214, n_4215, n_4216, n_4217, n_4218, n_4219, n_4220;
wire n_4205, n_4206, n_4207, n_4208, n_4209, n_4210, n_4211, n_4212;
wire n_4196, n_4198, n_4199, n_4200, n_4201, n_4202, n_4203, n_4204;
wire n_4186, n_4187, n_4188, n_4189, n_4190, n_4192, n_4193, n_4194;
wire n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185;
wire n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177;
wire n_4159, n_4160, n_4161, n_4163, n_4165, n_4167, n_4168, n_4169;
wire n_4149, n_4150, n_4151, n_4152, n_4154, n_4155, n_4156, n_4157;
wire n_4136, n_4137, n_4139, n_4140, n_4142, n_4145, n_4147, n_4148;
wire n_4123, n_4124, n_4125, n_4126, n_4131, n_4133, n_4134, n_4135;
wire n_4111, n_4113, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122;
wire n_4101, n_4102, n_4103, n_4105, n_4107, n_4108, n_4109, n_4110;
wire n_4086, n_4087, n_4088, n_4090, n_4091, n_4092, n_4096, n_4098;
wire n_4074, n_4076, n_4080, n_4081, n_4082, n_4083, n_4084, n_4085;
wire n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073;
wire n_4053, n_4054, n_4055, n_4056, n_4059, n_4060, n_4062, n_4065;
wire n_4042, n_4043, n_4044, n_4045, n_4046, n_4048, n_4049, n_4050;
wire n_4031, n_4032, n_4033, n_4034, n_4035, n_4037, n_4038, n_4040;
wire n_4020, n_4021, n_4022, n_4024, n_4025, n_4028, n_4029, n_4030;
wire n_4012, n_4013, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019;
wire n_4000, n_4002, n_4005, n_4006, n_4008, n_4009, n_4010, n_4011;
wire n_3990, n_3991, n_3992, n_3993, n_3995, n_3996, n_3997, n_3998;
wire n_3977, n_3978, n_3979, n_3981, n_3982, n_3983, n_3984, n_3985;
wire n_3966, n_3968, n_3969, n_3970, n_3971, n_3972, n_3973, n_3974;
wire n_3956, n_3957, n_3958, n_3959, n_3960, n_3962, n_3963, n_3964;
wire n_3946, n_3947, n_3948, n_3949, n_3951, n_3952, n_3953, n_3955;
wire n_3937, n_3938, n_3939, n_3941, n_3942, n_3943, n_3944, n_3945;
wire n_3916, n_3922, n_3925, n_3929, n_3932, n_3933, n_3934, n_3936;
wire n_3905, n_3906, n_3907, n_3910, n_3911, n_3913, n_3914, n_3915;
wire n_3895, n_3896, n_3897, n_3898, n_3900, n_3902, n_3903, n_3904;
wire n_3881, n_3882, n_3883, n_3885, n_3886, n_3891, n_3893, n_3894;
wire n_3866, n_3868, n_3869, n_3870, n_3873, n_3877, n_3878, n_3879;
wire n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, n_3861, n_3863;
wire n_3845, n_3846, n_3847, n_3848, n_3849, n_3851, n_3852, n_3854;
wire n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3843, n_3844;
wire n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835;
wire n_3817, n_3819, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826;
wire n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816;
wire n_3797, n_3798, n_3800, n_3801, n_3802, n_3803, n_3807, n_3808;
wire n_3784, n_3785, n_3786, n_3788, n_3789, n_3792, n_3793, n_3795;
wire n_3775, n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782;
wire n_3764, n_3765, n_3766, n_3767, n_3769, n_3770, n_3771, n_3774;
wire n_3744, n_3745, n_3746, n_3752, n_3753, n_3755, n_3758, n_3761;
wire n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3740, n_3742;
wire n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732;
wire n_3716, n_3717, n_3718, n_3720, n_3721, n_3722, n_3723, n_3724;
wire n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3715;
wire n_3693, n_3695, n_3697, n_3700, n_3701, n_3702, n_3703, n_3706;
wire n_3685, n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692;
wire n_3673, n_3674, n_3675, n_3677, n_3679, n_3680, n_3681, n_3683;
wire n_3659, n_3660, n_3661, n_3662, n_3666, n_3670, n_3671, n_3672;
wire n_3648, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3658;
wire n_3638, n_3639, n_3640, n_3641, n_3642, n_3645, n_3646, n_3647;
wire n_3627, n_3628, n_3629, n_3631, n_3633, n_3634, n_3636, n_3637;
wire n_3616, n_3618, n_3620, n_3621, n_3622, n_3624, n_3625, n_3626;
wire n_3605, n_3606, n_3609, n_3611, n_3612, n_3613, n_3614, n_3615;
wire n_3592, n_3593, n_3596, n_3598, n_3599, n_3601, n_3603, n_3604;
wire n_3580, n_3581, n_3582, n_3585, n_3588, n_3589, n_3590, n_3591;
wire n_3567, n_3569, n_3570, n_3571, n_3572, n_3574, n_3577, n_3578;
wire n_3555, n_3557, n_3559, n_3560, n_3561, n_3563, n_3564, n_3566;
wire n_3543, n_3546, n_3547, n_3549, n_3550, n_3551, n_3552, n_3554;
wire n_3533, n_3534, n_3535, n_3537, n_3538, n_3540, n_3541, n_3542;
wire n_3520, n_3521, n_3522, n_3523, n_3529, n_3530, n_3531, n_3532;
wire n_3510, n_3511, n_3512, n_3514, n_3516, n_3517, n_3518, n_3519;
wire n_3500, n_3501, n_3502, n_3503, n_3505, n_3506, n_3507, n_3508;
wire n_3491, n_3492, n_3493, n_3494, n_3496, n_3497, n_3498, n_3499;
wire n_3482, n_3483, n_3484, n_3486, n_3487, n_3488, n_3489, n_3490;
wire n_3471, n_3473, n_3475, n_3477, n_3478, n_3479, n_3480, n_3481;
wire n_3461, n_3463, n_3464, n_3465, n_3466, n_3468, n_3469, n_3470;
wire n_3447, n_3448, n_3449, n_3454, n_3455, n_3458, n_3459, n_3460;
wire n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442;
wire n_3426, n_3427, n_3429, n_3430, n_3431, n_3432, n_3433, n_3434;
wire n_3416, n_3417, n_3418, n_3420, n_3422, n_3423, n_3424, n_3425;
wire n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415;
wire n_3398, n_3399, n_3400, n_3402, n_3403, n_3404, n_3406, n_3407;
wire n_3385, n_3387, n_3388, n_3389, n_3390, n_3391, n_3394, n_3395;
wire n_3372, n_3373, n_3376, n_3377, n_3381, n_3382, n_3383, n_3384;
wire n_3363, n_3364, n_3365, n_3366, n_3368, n_3369, n_3370, n_3371;
wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362;
wire n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353;
wire n_3336, n_3337, n_3339, n_3340, n_3341, n_3343, n_3344, n_3345;
wire n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, n_3335;
wire n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327;
wire n_3310, n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3319;
wire n_3300, n_3301, n_3302, n_3303, n_3305, n_3307, n_3308, n_3309;
wire n_3288, n_3289, n_3290, n_3291, n_3292, n_3296, n_3298, n_3299;
wire n_3278, n_3279, n_3281, n_3282, n_3283, n_3285, n_3286, n_3287;
wire n_3269, n_3270, n_3271, n_3273, n_3274, n_3275, n_3276, n_3277;
wire n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, n_3267, n_3268;
wire n_3249, n_3253, n_3254, n_3255, n_3257, n_3258, n_3259, n_3260;
wire n_3234, n_3236, n_3239, n_3241, n_3242, n_3243, n_3244, n_3247;
wire n_3222, n_3223, n_3224, n_3225, n_3226, n_3228, n_3229, n_3233;
wire n_3212, n_3213, n_3214, n_3216, n_3217, n_3218, n_3219, n_3221;
wire n_3202, n_3204, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211;
wire n_3191, n_3192, n_3193, n_3194, n_3196, n_3197, n_3200, n_3201;
wire n_3181, n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3189;
wire n_3171, n_3172, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179;
wire n_3158, n_3160, n_3161, n_3162, n_3164, n_3165, n_3167, n_3170;
wire n_3147, n_3148, n_3149, n_3152, n_3153, n_3154, n_3156, n_3157;
wire n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146;
wire n_3130, n_3131, n_3132, n_3133, n_3135, n_3136, n_3137, n_3138;
wire n_3117, n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3127;
wire n_3108, n_3109, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116;
wire n_3098, n_3099, n_3100, n_3102, n_3103, n_3104, n_3105, n_3106;
wire n_3088, n_3090, n_3091, n_3092, n_3094, n_3095, n_3096, n_3097;
wire n_3079, n_3080, n_3081, n_3082, n_3084, n_3085, n_3086, n_3087;
wire n_3066, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3077;
wire n_3055, n_3056, n_3057, n_3058, n_3059, n_3062, n_3063, n_3065;
wire n_3043, n_3044, n_3047, n_3048, n_3049, n_3050, n_3052, n_3053;
wire n_3033, n_3034, n_3035, n_3036, n_3038, n_3040, n_3041, n_3042;
wire n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032;
wire n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022;
wire n_3005, n_3007, n_3008, n_3010, n_3011, n_3012, n_3013, n_3014;
wire n_2986, n_2987, n_2988, n_2989, n_2996, n_3001, n_3003, n_3004;
wire n_2974, n_2975, n_2977, n_2979, n_2980, n_2981, n_2983, n_2985;
wire n_2965, n_2966, n_2967, n_2968, n_2969, n_2971, n_2972, n_2973;
wire n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964;
wire n_2947, n_2948, n_2949, n_2951, n_2953, n_2954, n_2955, n_2956;
wire n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946;
wire n_2929, n_2930, n_2931, n_2933, n_2934, n_2936, n_2937, n_2938;
wire n_2917, n_2918, n_2920, n_2923, n_2924, n_2925, n_2926, n_2928;
wire n_2907, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915;
wire n_2897, n_2898, n_2900, n_2902, n_2903, n_2904, n_2905, n_2906;
wire n_2888, n_2889, n_2890, n_2891, n_2892, n_2894, n_2895, n_2896;
wire n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887;
wire n_2868, n_2869, n_2870, n_2871, n_2872, n_2875, n_2878, n_2879;
wire n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2866, n_2867;
wire n_2850, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, n_2858;
wire n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, n_2849;
wire n_2833, n_2834, n_2835, n_2837, n_2838, n_2839, n_2840, n_2841;
wire n_2824, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832;
wire n_2815, n_2816, n_2817, n_2819, n_2820, n_2821, n_2822, n_2823;
wire n_2806, n_2807, n_2808, n_2809, n_2810, n_2812, n_2813, n_2814;
wire n_2797, n_2798, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805;
wire n_2788, n_2789, n_2790, n_2791, n_2793, n_2794, n_2795, n_2796;
wire n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, n_2787;
wire n_2770, n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778;
wire n_2761, n_2762, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769;
wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
wire n_2742, n_2743, n_2744, n_2746, n_2747, n_2748, n_2749, n_2751;
wire n_2733, n_2734, n_2735, n_2736, n_2738, n_2739, n_2740, n_2741;
wire n_2720, n_2722, n_2723, n_2725, n_2727, n_2729, n_2730, n_2732;
wire n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2718, n_2719;
wire n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2709, n_2710;
wire n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2699, n_2700;
wire n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691;
wire n_2672, n_2673, n_2675, n_2677, n_2678, n_2679, n_2680, n_2682;
wire n_2663, n_2664, n_2665, n_2666, n_2668, n_2669, n_2670, n_2671;
wire n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662;
wire n_2645, n_2646, n_2647, n_2648, n_2651, n_2652, n_2653, n_2654;
wire n_2634, n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2644;
wire n_2616, n_2619, n_2624, n_2625, n_2628, n_2629, n_2630, n_2632;
wire n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615;
wire n_2598, n_2600, n_2601, n_2602, n_2603, n_2604, n_2606, n_2607;
wire n_2588, n_2589, n_2590, n_2592, n_2593, n_2594, n_2595, n_2597;
wire n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587;
wire n_2567, n_2572, n_2573, n_2574, n_2575, n_2577, n_2578, n_2579;
wire n_2557, n_2558, n_2559, n_2560, n_2562, n_2563, n_2564, n_2566;
wire n_2545, n_2546, n_2548, n_2550, n_2551, n_2554, n_2555, n_2556;
wire n_2533, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2543;
wire n_2522, n_2523, n_2524, n_2526, n_2528, n_2529, n_2530, n_2531;
wire n_2512, n_2514, n_2515, n_2517, n_2518, n_2519, n_2520, n_2521;
wire n_2501, n_2502, n_2503, n_2504, n_2506, n_2507, n_2509, n_2510;
wire n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500;
wire n_2481, n_2483, n_2484, n_2485, n_2486, n_2488, n_2491, n_2492;
wire n_2468, n_2469, n_2471, n_2472, n_2474, n_2475, n_2479, n_2480;
wire n_2458, n_2459, n_2460, n_2461, n_2463, n_2464, n_2465, n_2466;
wire n_2448, n_2449, n_2451, n_2452, n_2453, n_2454, n_2456, n_2457;
wire n_2437, n_2438, n_2439, n_2441, n_2442, n_2443, n_2444, n_2447;
wire n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436;
wire n_2416, n_2419, n_2421, n_2423, n_2425, n_2426, n_2427, n_2428;
wire n_2403, n_2406, n_2408, n_2409, n_2410, n_2413, n_2414, n_2415;
wire n_2387, n_2388, n_2389, n_2391, n_2392, n_2397, n_2398, n_2400;
wire n_2373, n_2374, n_2375, n_2376, n_2378, n_2379, n_2382, n_2385;
wire n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2370, n_2372;
wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2356, n_2361;
wire n_2340, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
wire n_2327, n_2329, n_2331, n_2332, n_2334, n_2336, n_2338, n_2339;
wire n_2316, n_2319, n_2320, n_2321, n_2323, n_2324, n_2325, n_2326;
wire n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312;
wire n_2293, n_2294, n_2296, n_2298, n_2301, n_2302, n_2303, n_2304;
wire n_2283, n_2284, n_2285, n_2286, n_2288, n_2289, n_2290, n_2291;
wire n_2271, n_2272, n_2274, n_2276, n_2277, n_2278, n_2280, n_2281;
wire n_2260, n_2263, n_2264, n_2265, n_2266, n_2268, n_2269, n_2270;
wire n_2250, n_2252, n_2253, n_2254, n_2255, n_2256, n_2258, n_2259;
wire n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249;
wire n_2229, n_2230, n_2231, n_2233, n_2234, n_2237, n_2239, n_2241;
wire n_2218, n_2219, n_2221, n_2223, n_2224, n_2225, n_2227, n_2228;
wire n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2215, n_2216;
wire n_2180, n_2181, n_2182, n_2192, n_2203, n_2204, n_2205, n_2206;
wire n_2167, n_2168, n_2172, n_2173, n_2174, n_2176, n_2177, n_2178;
wire n_2156, n_2157, n_2159, n_2160, n_2161, n_2163, n_2165, n_2166;
wire n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155;
wire n_2137, n_2138, n_2140, n_2141, n_2143, n_2144, n_2145, n_2146;
wire n_2128, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135;
wire n_2116, n_2118, n_2119, n_2120, n_2121, n_2122, n_2126, n_2127;
wire n_2106, n_2107, n_2108, n_2110, n_2111, n_2113, n_2114, n_2115;
wire n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2103;
wire n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094;
wire n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086;
wire n_2065, n_2067, n_2068, n_2069, n_2070, n_2072, n_2077, n_2078;
wire n_2055, n_2056, n_2057, n_2060, n_2061, n_2062, n_2063, n_2064;
wire n_2044, n_2045, n_2046, n_2048, n_2049, n_2051, n_2053, n_2054;
wire n_2030, n_2031, n_2032, n_2034, n_2038, n_2039, n_2042, n_2043;
wire n_2018, n_2019, n_2020, n_2023, n_2024, n_2025, n_2027, n_2029;
wire n_2007, n_2008, n_2009, n_2011, n_2014, n_2015, n_2016, n_2017;
wire n_1997, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006;
wire n_1986, n_1989, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996;
wire n_1972, n_1975, n_1976, n_1977, n_1979, n_1980, n_1982, n_1985;
wire n_1882, n_1883, n_1884, n_1885, n_1887, n_1968, n_1969, n_1971;
wire n_1859, n_1860, n_1861, n_1862, n_1863, n_1865, n_1869, n_1875;
wire n_1848, n_1849, n_1850, n_1851, n_1854, n_1855, n_1857, n_1858;
wire n_1839, n_1840, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847;
wire n_1822, n_1826, n_1827, n_1830, n_1831, n_1832, n_1833, n_1838;
wire n_1812, n_1813, n_1814, n_1817, n_1818, n_1819, n_1820, n_1821;
wire n_1804, n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811;
wire n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803;
wire n_1787, n_1788, n_1789, n_1791, n_1792, n_1793, n_1794, n_1795;
wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1783, n_1785, n_1786;
wire n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1775;
wire n_1758, n_1759, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766;
wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757;
wire n_1741, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
wire n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1740;
wire n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731;
wire n_1715, n_1716, n_1717, n_1718, n_1719, n_1721, n_1722, n_1723;
wire n_1706, n_1707, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714;
wire n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705;
wire n_1686, n_1687, n_1688, n_1689, n_1691, n_1694, n_1695, n_1696;
wire n_1674, n_1675, n_1676, n_1677, n_1678, n_1680, n_1681, n_1682;
wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672;
wire n_1649, n_1650, n_1652, n_1655, n_1656, n_1657, n_1658, n_1662;
wire n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647;
wire n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1636;
wire n_1590, n_1591, n_1592, n_1597, n_1599, n_1605, n_1625, n_1626;
wire n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587;
wire n_1568, n_1569, n_1570, n_1571, n_1574, n_1575, n_1576, n_1578;
wire n_1557, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1567;
wire n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556;
wire n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548;
wire n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540;
wire n_1524, n_1525, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532;
wire n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523;
wire n_1505, n_1506, n_1507, n_1509, n_1510, n_1511, n_1514, n_1515;
wire n_1488, n_1491, n_1493, n_1494, n_1499, n_1500, n_1502, n_1503;
wire n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1486, n_1487;
wire n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478;
wire n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470;
wire n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462;
wire n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454;
wire n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446;
wire n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438;
wire n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429;
wire n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419;
wire n_1402, n_1403, n_1404, n_1405, n_1407, n_1408, n_1409, n_1411;
wire n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401;
wire n_1381, n_1382, n_1384, n_1388, n_1390, n_1391, n_1392, n_1393;
wire n_1366, n_1367, n_1369, n_1370, n_1373, n_1375, n_1377, n_1380;
wire n_1349, n_1351, n_1352, n_1353, n_1354, n_1356, n_1363, n_1364;
wire n_1322, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
wire n_1307, n_1308, n_1310, n_1311, n_1312, n_1313, n_1315, n_1321;
wire n_1292, n_1293, n_1295, n_1296, n_1298, n_1299, n_1300, n_1304;
wire n_1278, n_1279, n_1282, n_1283, n_1285, n_1286, n_1290, n_1291;
wire n_1269, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
wire n_1260, n_1261, n_1262, n_1263, n_1264, n_1266, n_1267, n_1268;
wire n_1246, n_1247, n_1248, n_1250, n_1251, n_1252, n_1255, n_1257;
wire n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245;
wire n_1228, n_1230, n_1231, n_1232, n_1234, n_1235, n_1236, n_1237;
wire n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227;
wire n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1219;
wire n_1201, n_1202, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210;
wire n_1191, n_1192, n_1193, n_1194, n_1195, n_1198, n_1199, n_1200;
wire n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189;
wire n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181;
wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1173;
wire n_1154, n_1155, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163;
wire n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1152, n_1153;
wire n_1133, n_1135, n_1136, n_1137, n_1138, n_1139, n_1143, n_1144;
wire n_1121, n_1122, n_1123, n_1124, n_1127, n_1128, n_1130, n_1131;
wire n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120;
wire n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112;
wire n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104;
wire n_1083, n_1084, n_1085, n_1090, n_1093, n_1094, n_1095, n_1096;
wire n_1071, n_1072, n_1074, n_1075, n_1077, n_1079, n_1081, n_1082;
wire n_1058, n_1059, n_1060, n_1062, n_1063, n_1064, n_1065, n_1069;
wire n_1040, n_1043, n_1044, n_1046, n_1052, n_1053, n_1054, n_1055;
wire n_1013, n_1014, n_1015, n_1016, n_1017, n_1021, n_1023, n_1024;
wire n_992, n_993, n_994, n_995, n_998, n_999, n_1002, n_1011;
wire n_981, n_982, n_983, n_986, n_987, n_988, n_989, n_991;
wire n_971, n_973, n_974, n_975, n_976, n_977, n_978, n_980;
wire n_957, n_958, n_961, n_963, n_965, n_967, n_969, n_970;
wire n_946, n_947, n_948, n_950, n_952, n_954, n_955, n_956;
wire n_932, n_933, n_934, n_937, n_938, n_940, n_942, n_943;
wire n_923, n_924, n_925, n_926, n_927, n_928, n_929, n_931;
wire n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921;
wire n_904, n_905, n_906, n_908, n_909, n_910, n_911, n_912;
wire n_896, n_897, n_898, n_899, n_900, n_901, n_902, n_903;
wire n_886, n_887, n_888, n_890, n_891, n_893, n_894, n_895;
wire n_877, n_878, n_880, n_881, n_882, n_883, n_884, n_885;
wire n_863, n_864, n_866, n_867, n_868, n_871, n_872, n_876;
wire n_855, n_856, n_857, n_858, n_859, n_860, n_861, n_862;
wire n_845, n_846, n_847, n_848, n_849, n_851, n_852, n_854;
wire n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844;
wire n_829, n_830, n_831, n_832, n_833, n_834, n_835, n_836;
wire n_820, n_821, n_822, n_823, n_824, n_826, n_827, n_828;
wire n_808, n_810, n_812, n_814, n_816, n_817, n_818, n_819;
wire n_800, n_801, n_802, n_803, n_804, n_805, n_806, n_807;
wire n_790, n_791, n_793, n_794, n_795, n_797, n_798, n_799;
wire n_778, n_779, n_780, n_782, n_783, n_784, n_786, n_789;
wire n_748, n_765, n_769, n_771, n_772, n_775, n_776, n_777;
wire n_730, n_739, n_740, n_741, n_744, n_745, n_746, n_747;
wire n_716, n_717, n_718, n_719, n_720, n_722, n_723, n_724;
wire n_702, n_704, n_705, n_707, n_708, n_709, n_714, n_715;
wire n_691, n_692, n_693, n_694, n_695, n_696, n_697, n_698;
wire n_677, n_678, n_680, n_684, n_685, n_686, n_688, n_690;
wire n_664, n_667, n_669, n_670, n_673, n_674, n_675, n_676;
wire n_650, n_652, n_653, n_659, n_660, n_661, n_662, n_663;
wire n_638, n_639, n_640, n_643, n_644, n_647, n_648, n_649;
wire n_624, n_626, n_627, n_628, n_629, n_635, n_636, n_637;
wire n_615, n_616, n_617, n_618, n_619, n_620, n_621, n_623;
wire n_600, n_603, n_607, n_608, n_609, n_610, n_611, n_612;
wire n_591, n_592, n_594, n_595, n_596, n_597, n_598, n_599;
wire n_580, n_581, n_584, n_585, n_587, n_588, n_589, n_590;
wire n_565, n_566, n_568, n_571, n_572, n_575, n_578, n_579;
wire n_553, n_556, n_557, n_558, n_561, n_562, n_563, n_564;
wire n_524, n_527, n_538, n_540, n_546, n_549, n_551, n_552;
wire n_511, n_512, n_515, n_518, n_519, n_521, n_522, n_523;
wire n_487, n_488, n_490, n_491, n_493, n_496, n_503, n_504;
wire n_469, n_470, n_471, n_474, n_477, n_479, n_482, n_486;
wire n_456, n_458, n_459, n_460, n_461, n_463, n_464, n_465;
wire n_442, n_444, n_446, n_447, n_448, n_450, n_453, n_455;
wire n_424, n_425, n_428, n_429, n_433, n_436, n_437, n_441;
wire n_411, n_412, n_413, n_415, n_416, n_417, n_418, n_423;
wire n_392, n_397, n_399, n_401, n_404, n_406, n_408, n_409;
wire n_377, n_379, n_380, n_382, n_383, n_386, n_388, n_389;
wire n_364, n_365, n_367, n_368, n_370, n_371, n_374, n_376;
wire n_343, n_344, n_347, n_351, n_353, n_356, n_360, n_362;
wire n_332, n_334, n_335, n_336, n_338, n_339, n_340, n_342;
wire n_317, n_322, n_323, n_325, n_326, n_327, n_328, n_330;
wire n_298, n_302, n_303, n_307, n_308, n_309, n_311, n_316;
wire n_284, n_286, n_287, n_290, n_291, n_294, n_295, n_297;
wire n_268, n_269, n_271, n_273, n_276, n_278, n_281, n_282;
wire n_245, n_247, n_248, n_251, n_259, n_261, n_262, n_263;
wire n_227, n_234, n_235, n_238, n_240, n_241, n_242, n_243;
wire n_209, n_213, n_215, n_218, n_220, n_221, n_223, n_224;
wire n_187, n_188, n_191, n_194, n_196, n_202, n_204, n_205;
wire n_153, n_157, n_158, n_162, n_165, n_168, n_169, n_172;
wire n_128, n_129, n_134, n_136, n_143, n_144, n_150, n_151;
wire n_105, n_107, n_110, n_117, n_118, n_125, n_126, n_127;
wire n_92, n_93, n_94, n_95, n_96, n_98, n_101, n_103;
wire n_74, n_75, n_79, n_83, n_85, n_86, n_87, n_89;
wire n_57, n_59, n_60, n_64, n_65, n_67, n_69, n_70;
wire n_38, n_39, n_40, n_43, n_46, n_50, n_52, n_54;
wire n_23, n_26, n_27, n_28, n_29, n_30, n_32, n_35;
wire n_12, n_13, n_16, n_17, n_19, n_20, n_21, n_22;
wire g_22639, gbuf1, gbuf3, n_0, n_1, n_2, n_5, n_11;
wire g_22328, g_22349, g_22371, g_22379, g_22464, g_22552, g_22600, g_22605;
wire g_21806, g_21813, g_22021, g_22034, g_22038, g_22070, g_22236, g_22306;
wire g_21318, g_21447, g_21576, g_21651, g_21720, g_21778, g_21792, g_21799;
wire g_20268, g_20563, g_20614, g_20837, g_20839, g_20909, g_20951, g_20952;
wire g_19659, g_19789, g_19911, g_19913, g_20073, g_20159, g_20208, g_20244;
wire g_19233, g_19241, g_19289, g_19304, g_19414, g_19459, g_19492, g_19515;
wire g_18869, g_18902, g_18980, g_18996, g_19113, g_19136, g_19172, g_19187;
wire g_18308, g_18330, g_18488, g_18590, g_18635, g_18739, g_18793, g_18795;
wire g_17426, g_17653, g_17934, g_18015, g_18112, g_18200, g_18220, g_18238;
wire g_16571, g_16677, g_16769, g_16792, g_16958, g_16983, g_17065, g_17086;
wire g_15879, g_16063, g_16296, g_16311, g_16404, g_16456, g_16464, g_16475;
wire g_15287, g_15380, g_15381, g_15691, g_15740, g_15758, g_15801, g_15838;
wire g_14265, g_14342, g_14535, g_14587, g_14843, g_14965, g_15016, g_15127;
wire g_12922, g_13091, g_13255, g_13278, g_13758, g_13838, g_13871, g_13901;
wire g_11037, g_11293, g_11413, g_12275, g_12276, g_12433, g_12465, g_12791;
wire g_9338, g_9584, g_10092, g_10233, g_10278, g_10556, g_10715, g_10903;
wire g_7220, g_7563, g_8657, g_8864, g_8896, g_9174, g_9176, g_9298;
wire g_5508, g_6131, g_6165, g_6192, g_6283, g_6579, g_6701, g_7062;
wire g_4050, g_4409, g_4449, g_5029, g_5156, g_5313, g_5342, g_5450;
wire g34027, g34028, g34034, g34035, g34036, g_3381, g_3861, g_3974;
wire g6649, g6653, g6657, g6723, g6732, g6736, g6741, g34026;
wire g6617, g6621, g6625, g6629, g6633, g6637, g6641, g6645;
wire g6585, g6589, g6593, g6597, g6601, g6605, g6609, g6613;
wire g6533, g6537, g6541, g6549, g6555, g6565, g6573, g6581;
wire g6444, g6494, g6505, g6509, g6513, g6519, g6523, g6527;
wire g6307, g6311, g6336, g6377, g6381, g6386, g6390, g6395;
wire g6275, g6279, g6283, g6287, g6291, g6295, g6299, g6303;
wire g6243, g6247, g6251, g6255, g6259, g6263, g6267, g6271;
wire g6191, g6195, g6203, g6209, g6219, g6227, g6235, g6239;
wire g6148, g6159, g6163, g6167, g6173, g6177, g6181, g6187;
wire g5961, g5965, g5990, g6031, g6035, g6040, g6044, g6098;
wire g5929, g5933, g5937, g5941, g5945, g5949, g5953, g5957;
wire g5897, g5901, g5905, g5909, g5913, g5917, g5921, g5925;
wire g5845, g5849, g5857, g5863, g5873, g5881, g5889, g5893;
wire g5802, g5813, g5817, g5821, g5827, g5831, g5835, g5841;
wire g5615, g5619, g5644, g5685, g5689, g5694, g5698, g5752;
wire g5583, g5587, g5591, g5595, g5599, g5603, g5607, g5611;
wire g5551, g5555, g5559, g5563, g5567, g5571, g5575, g5579;
wire g5499, g5503, g5511, g5517, g5527, g5535, g5543, g5547;
wire g5456, g5467, g5471, g5475, g5481, g5485, g5489, g5495;
wire g5268, g5272, g5297, g5339, g5343, g5348, g5352, g5406;
wire g5236, g5240, g5244, g5248, g5252, g5256, g5260, g5264;
wire g5204, g5208, g5212, g5216, g5220, g5224, g5228, g5232;
wire g5152, g5156, g5164, g5170, g5180, g5188, g5196, g5200;
wire g5112, g5120, g5124, g5128, g5134, g5138, g5142, g5148;
wire g5069, g5073, g5077, g5080, g5084, g5092, g5097, g5109;
wire g5016, g5029, g5033, g5037, g5041, g5046, g5052, g5057;
wire g4944, g4950, g4955, g4961, g4966, g4983, g4991, g5011;
wire g4899, g4907, g4912, g4917, g4922, g4927, g4933, g4939;
wire g4826, g4831, g4843, g4849, g4854, g4878, g4888, g4894;
wire g4754, g4760, g4765, g4771, g4776, g4785, g4793, g4821;
wire g4709, g4717, g4722, g4727, g4732, g4737, g4743, g4749;
wire g4633, g4653, g4659, g4664, g4669, g4688, g4698, g4704;
wire g4581, g4584, g4593, g4601, g4608, g4616, g4621, g4628;
wire g4558, g4561, g4564, g4567, g4570, g4572, g4575, g4578;
wire g4531, g4534, g4540, g4543, g4546, g4549, g4552, g4555;
wire g4498, g4501, g4504, g4512, g4515, g4519, g4521, g4527;
wire g4474, g4477, g4480, g4483, g4486, g4489, g4492, g4495;
wire g4443, g4452, g4455, g4456, g4459, g4462, g4467, g4473;
wire g4411, g4417, g4420, g4423, g4427, g4430, g4434, g4438;
wire g4369, g4372, g4375, g4382, g4388, g4392, g4401, g4405;
wire g4291, g4297, g4300, g4308, g4311, g4332, g4349, g4366;
wire g4249, g4253, g4258, g4264, g4269, g4273, g4281, g4284;
wire g4157, g4164, g4172, g4176, g4235, g4239, g4242, g4245;
wire g4112, g4116, g4119, g4122, g4141, g4145, g4146, g4153;
wire g4072, g4076, g4082, g4087, g4093, g4098, g4104, g4108;
wire g4031, g4035, g4040, g4045, g4049, g4054, g4057, g4064;
wire g3941, g3945, g3949, g3953, g3957, g3961, g3965, g3990;
wire g3909, g3913, g3917, g3921, g3925, g3929, g3933, g3937;
wire g3863, g3873, g3881, g3889, g3893, g3897, g3901, g3905;
wire g3821, g3827, g3831, g3835, g3841, g3845, g3849, g3857;
wire g3689, g3694, g3698, g3752, g3802, g3808, g3813, g3817;
wire g3598, g3602, g3606, g3610, g3614, g3639, g3680, g3684;
wire g3566, g3570, g3574, g3578, g3582, g3586, g3590, g3594;
wire g3530, g3538, g3542, g3546, g3550, g3554, g3558, g3562;
wire g3480, g3484, g3490, g3494, g3498, g3506, g3512, g3522;
wire g3347, g3401, g3451, g3457, g3462, g3466, g3470, g3476;
wire g3255, g3259, g3263, g3288, g3329, g3333, g3338, g3343;
wire g3223, g3227, g3231, g3235, g3239, g3243, g3247, g3251;
wire g3191, g3195, g3199, g3203, g3207, g3211, g3215, g3219;
wire g3139, g3143, g3147, g3155, g3161, g3171, g3179, g3187;
wire g3100, g3106, g3111, g3115, g3119, g3125, g3129, g3133;
wire g2975, g2980, g2984, g2988, g2994, g2999, g3003, g3050;
wire g2936, g2941, g2946, g2950, g2955, g2960, g2965, g2970;
wire g2898, g2902, g2907, g2912, g2917, g2922, g2927, g2932;
wire g2864, g2868, g2873, g2878, g2882, g2886, g2890, g2894;
wire g2819, g2823, g2827, g2844, g2848, g2852, g2856, g2860;
wire g2787, g2791, g2795, g2799, g2803, g2807, g2811, g2815;
wire g2756, g2759, g2763, g2767, g2771, g2775, g2779, g2783;
wire g2681, g2685, g2697, g2704, g2715, g2724, g2735, g2748;
wire g2643, g2648, g2652, g2657, g2661, g2667, g2671, g2675;
wire g2587, g2595, g2599, g2606, g2619, g2625, g2629, g2638;
wire g2551, g2555, g2563, g2567, g2571, g2575, g2579, g2583;
wire g2514, g2518, g2523, g2527, g2533, g2537, g2541, g2547;
wire g2453, g2461, g2465, g2472, g2485, g2491, g2504, g2509;
wire g2417, g2421, g2429, g2433, g2437, g2441, g2445, g2449;
wire g2380, g2384, g2389, g2393, g2399, g2403, g2407, g2413;
wire g2327, g2331, g2338, g2351, g2357, g2361, g2370, g2375;
wire g2287, g2295, g2299, g2303, g2307, g2311, g2315, g2319;
wire g2250, g2255, g2259, g2265, g2269, g2273, g2279, g2283;
wire g2197, g2204, g2217, g2223, g2227, g2236, g2241, g2246;
wire g2161, g2165, g2169, g2173, g2177, g2181, g2185, g2193;
wire g2112, g2116, g2122, g2126, g2130, g2138, g2145, g2153;
wire g2070, g2079, g2084, g2089, g2093, g2098, g2102, g2108;
wire g2020, g2024, g2028, g2036, g2040, g2047, g2060, g2066;
wire g1982, g1988, g1992, g1996, g2004, g2008, g2012, g2016;
wire g1945, g1950, g1955, g1959, g1964, g1968, g1974, g1978;
wire g1890, g1894, g1902, g1906, g1913, g1926, g1932, g1936;
wire g1854, g1858, g1862, g1870, g1874, g1878, g1882, g1886;
wire g1816, g1821, g1825, g1830, g1834, g1840, g1844, g1848;
wire g1756, g1760, g1768, g1772, g1779, g1792, g1798, g1811;
wire g1720, g1724, g1728, g1736, g1740, g1744, g1748, g1752;
wire g1682, g1687, g1691, g1696, g1700, g1706, g1710, g1714;
wire g1620, g1624, g1632, g1636, g1644, g1657, g1664, g1677;
wire g1585, g1589, g1592, g1600, g1604, g1608, g1612, g1616;
wire g1526, g1532, g1536, g1542, g1548, g1554, g1564, g1579;
wire g1448, g1454, g1467, g1472, g1478, g1484, g1489, g1521;
wire g1384, g1389, g1395, g1404, g1413, g1430, g1437, g1442;
wire g1333, g1339, g1345, g1351, g1361, g1367, g1373, g1379;
wire g1242, g1246, g1291, g1300, g1306, g1312, g1319, g1322;
wire g55, g1171, g1178, g1183, g1189, g1199, g1221, g1236;
wire g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972;
wire blif_clk_net, blif_reset_net, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753;
assign g34972 = 1'b1;
assign g34956 = g34839;
assign g34927 = 1'b1;
assign g34925 = 1'b1;
assign g34923 = 1'b1;
assign g34921 = 1'b1;
assign g34919 = 1'b1;
assign g34917 = 1'b1;
assign g34915 = 1'b1;
assign g34913 = 1'b1;
assign g34788 = g33894;
assign g34597 = 1'b0;
assign g34437 = 1'b1;
assign g34436 = 1'b1;
assign g34435 = g31521;
assign g34425 = 1'b1;
assign g34383 = 1'b1;
assign g34240 = 1'b1;
assign g34239 = 1'b1;
assign g34238 = 1'b1;
assign g34237 = 1'b1;
assign g34236 = 1'b1;
assign g34235 = 1'b1;
assign g34234 = 1'b1;
assign g34233 = 1'b1;
assign g34232 = 1'b1;
assign g34221 = 1'b1;
assign g34201 = 1'b1;
assign g33959 = g28753;
assign g33950 = 1'b1;
assign g33949 = 1'b1;
assign g33948 = 1'b1;
assign g33947 = 1'b1;
assign g33946 = 1'b1;
assign g33945 = 1'b1;
assign g33935 = 1'b1;
assign g33874 = 1'b1;
assign g33659 = 1'b1;
assign g33636 = 1'b1;
assign g33533 = g27831;
assign g32975 = g26801;
assign g32454 = 1'b1;
assign g32429 = 1'b1;
assign g31863 = g25167;
assign g31862 = g25259;
assign g31861 = g25219;
assign g31860 = g25114;
assign g31665 = 1'b1;
assign g31656 = 1'b1;
assign g30332 = g23683;
assign g30331 = g23759;
assign g30330 = g23652;
assign g30329 = g23612;
assign g30327 = g23002;
assign g29221 = g21292;
assign g29220 = g21245;
assign g29219 = g20654;
assign g29218 = g18881;
assign g29217 = g21270;
assign g29216 = g21176;
assign g29215 = g20901;
assign g29214 = g20652;
assign g29213 = g20557;
assign g29212 = g20899;
assign g29211 = g20763;
assign g29210 = g20049;
assign g25590 = 1'b1;
assign g25589 = 1'b1;
assign g25588 = 1'b1;
assign g25587 = 1'b1;
assign g25586 = 1'b1;
assign g25585 = 1'b1;
assign g25584 = 1'b1;
assign g25583 = 1'b1;
assign g25582 = 1'b1;
assign g24151 = 1'b1;
assign g23190 = 1'b1;
assign g21698 = g36;
assign g18101 = g6746;
assign g18100 = g6751;
assign g18099 = g6745;
assign g18098 = g6744;
assign g18097 = g6747;
assign g18096 = g6750;
assign g18095 = g6749;
assign g18094 = g6748;
assign g18092 = g6753;
assign g12368 = 1'b0;
assign g9048 = 1'b0;
assign g8403 = 1'b0;
assign g8353 = 1'b0;
assign g8283 = 1'b0;
assign g8235 = 1'b0;
assign g8178 = 1'b0;
assign g8132 = 1'b0;
CLKBUFX1 gbuf_d_1(.A(n_6422), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(g2955));
MX2X1 g60853(.A (g2941), .B (n_6417), .S0 (n_8955), .Y (n_6422));
CLKBUFX1 gbuf_d_2(.A(n_6419), .Y(d_out_2));
CLKBUFX1 gbuf_qn_2(.A(qn_in_2), .Y(g2864));
NAND3X1 g60850(.A (n_6418), .B (n_6408), .C (n_6416), .Y (g31793));
MX2X1 g60856(.A (n_3499), .B (n_6415), .S0 (n_9000), .Y (n_6419));
NOR2X1 g60852(.A (n_6411), .B (n_6412), .Y (n_6418));
NAND4X1 g60857(.A (n_6414), .B (n_2449), .C (n_3614), .D (n_3498), .Y(n_6417));
AOI21X1 g60855(.A0 (n_6394), .A1 (n_6401), .B0 (n_6410), .Y (n_6416));
OR2X1 g60860(.A (n_6413), .B (n_271), .Y (n_6415));
NOR2X1 g60861(.A (n_3502), .B (n_6413), .Y (n_6414));
OAI33X1 g60854(.A0 (n_1414), .A1 (n_6409), .A2 (n_901), .B0 (n_1454),.B1 (n_6397), .B2 (n_3812), .Y (n_6412));
NAND3X1 g60858(.A (n_6405), .B (n_6386), .C (n_6403), .Y (n_6411));
OAI33X1 g60859(.A0 (n_3376), .A1 (n_1537), .A2 (n_6390), .B0(n_6409), .B1 (n_6402), .B2 (n_6406), .Y (n_6410));
NAND3X1 g60863(.A (n_6407), .B (n_6404), .C (n_2019), .Y (n_6408));
NAND4X1 g60864(.A (n_6407), .B (n_6406), .C (n_1321), .D (n_6398), .Y(n_6413));
NAND4X1 g60865(.A (n_6393), .B (n_1543), .C (n_1321), .D (n_6404), .Y(n_6405));
OR4X1 g60866(.A (n_6390), .B (n_6402), .C (n_6400), .D (n_6399), .Y(n_6403));
OAI21X1 g60862(.A0 (n_6388), .A1 (n_6400), .B0 (n_6389), .Y (n_6401));
NAND4X1 g60867(.A (n_6396), .B (n_6399), .C (n_6395), .D (n_6398), .Y(n_6409));
NAND4X1 g60868(.A (n_6396), .B (n_1212), .C (n_6395), .D (n_6406), .Y(n_6397));
AND2X1 g60869(.A (n_6394), .B (n_6392), .Y (n_6407));
AND2X1 g60871(.A (n_1213), .B (n_6392), .Y (n_6393));
INVX1 g60875(.A (n_6396), .Y (n_6390));
NAND4X1 g60872(.A (n_6388), .B (n_6404), .C (n_4878), .D (n_1321), .Y(n_6389));
AND2X1 g60873(.A (n_6388), .B (n_1055), .Y (n_6392));
AND2X1 g60876(.A (n_6388), .B (n_3641), .Y (n_6396));
NAND4X1 g60870(.A (n_6388), .B (n_1536), .C (n_6399), .D (n_3211), .Y(n_6386));
OAI21X1 g60877(.A0 (g4420), .A1 (g4427), .B0 (g35), .Y (n_6388));
CLKBUFX1 gbuf_d_3(.A(n_6385), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(g4420));
MX2X1 g60879(.A (g4534), .B (n_6384), .S0 (n_10005), .Y (n_6385));
XOR2X1 g60880(.A (g4534), .B (g10306), .Y (n_6384));
CLKBUFX1 gbuf_d_4(.A(n_6383), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(g4534));
OAI21X1 g60882(.A0 (n_6379), .A1 (n_9627), .B0 (n_6382), .Y (n_6383));
OAI21X1 g60883(.A0 (n_6381), .A1 (g2988), .B0 (n_9091), .Y (n_6382));
INVX1 g60884(.A (n_6380), .Y (n_6381));
NAND4X1 g60885(.A (g4564), .B (g4555), .C (g4561), .D (g4558), .Y(n_6380));
INVX1 g60886(.A (g4564), .Y (n_6379));
CLKBUFX1 gbuf_d_5(.A(n_6378), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(g4564));
NAND2X1 g60888(.A (n_6377), .B (n_3113), .Y (n_6378));
NAND2X1 g60889(.A (g4561), .B (n_10078), .Y (n_6377));
CLKBUFX1 gbuf_d_6(.A(n_6376), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(g4561));
NAND2X1 g60891(.A (n_6375), .B (n_3115), .Y (n_6376));
NAND2X1 g60892(.A (g4558), .B (n_10078), .Y (n_6375));
CLKBUFX1 gbuf_d_7(.A(n_6373), .Y(d_out_7));
CLKBUFX1 gbuf_q_7(.A(q_in_7), .Y(g4558));
NAND2X1 g60896(.A (n_6372), .B (n_3117), .Y (n_6373));
NAND2X1 g60898(.A (g4555), .B (n_10078), .Y (n_6372));
CLKBUFX1 gbuf_d_8(.A(gbuf3), .Y(d_out_8));
CLKBUFX1 gbuf_q_8(.A(q_in_8), .Y(g4555));
CLKBUFX1 gbuf_d_9(.A(g4570), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(gbuf3));
CLKBUFX1 gbuf_d_10(.A(n_6370), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(g20763));
CLKBUFX1 gbuf_d_11(.A(n_6371), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(g4570));
CLKBUFX1 gbuf_d_12(.A(n_6369), .Y(d_out_12));
CLKBUFX1 gbuf_q_12(.A(q_in_12), .Y(g_12276));
OAI21X1 g60911(.A0 (n_6364), .A1 (g4552), .B0 (n_6060), .Y (n_6371));
MX2X1 g60962(.A (g_12276), .B (n_6367), .S0 (n_8955), .Y (n_6370));
OAI21X1 g60984(.A0 (g_21792), .A1 (n_9422), .B0 (n_6368), .Y(n_6369));
CLKBUFX1 gbuf_d_13(.A(n_6365), .Y(d_out_13));
CLKBUFX1 gbuf_qn_13(.A(qn_in_13), .Y(g4552));
NAND3X1 g61012(.A (n_6366), .B (g_21792), .C (n_9681), .Y (n_6368));
MX2X1 g61019(.A (n_6366), .B (g20763), .S0 (g_21792), .Y (n_6367));
OAI21X1 g60929(.A0 (g4549), .A1 (n_6364), .B0 (n_6055), .Y (n_6365));
CLKBUFX1 gbuf_d_14(.A(n_6363), .Y(d_out_14));
CLKBUFX1 gbuf_qn_14(.A(qn_in_14), .Y(g_21792));
CLKBUFX1 gbuf_d_15(.A(n_6362), .Y(d_out_15));
CLKBUFX1 gbuf_qn_15(.A(qn_in_15), .Y(g4512));
MX2X1 g61142(.A (n_6359), .B (n_9772), .S0 (g_8657), .Y (n_6363));
CLKBUFX1 gbuf_d_16(.A(n_6361), .Y(d_out_16));
CLKBUFX1 gbuf_qn_16(.A(qn_in_16), .Y(g4549));
CLKBUFX1 gbuf_d_17(.A(n_6360), .Y(d_out_17));
CLKBUFX1 gbuf_q_17(.A(q_in_17), .Y(g4300));
OAI21X1 g60944(.A0 (g4504), .A1 (n_6364), .B0 (n_5821), .Y (n_6362));
OAI21X1 g60986(.A0 (g4546), .A1 (n_6364), .B0 (n_6320), .Y (n_6361));
MX2X1 g61143(.A (g4297), .B (n_6357), .S0 (n_9750), .Y (n_6360));
CLKBUFX1 gbuf_d_18(.A(n_6508), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(g_9338));
AND2X1 g61205(.A (n_9553), .B (g7540), .Y (n_6359));
CLKBUFX1 gbuf_d_19(.A(g7540), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(g_8657));
CLKBUFX1 gbuf_d_20(.A(n_6356), .Y(d_out_20));
CLKBUFX1 gbuf_qn_20(.A(qn_in_20), .Y(g4504));
CLKBUFX1 gbuf_d_21(.A(n_6355), .Y(d_out_21));
CLKBUFX1 gbuf_q_21(.A(q_in_21), .Y(g_10233));
CLKBUFX1 gbuf_d_22(.A(n_6351), .Y(d_out_22));
CLKBUFX1 gbuf_qn_22(.A(qn_in_22), .Y(g4546));
OR2X1 g61211(.A (g4242), .B (g4300), .Y (n_6357));
CLKBUFX1 gbuf_d_23(.A(n_6348), .Y(d_out_23));
CLKBUFX1 gbuf_q_23(.A(q_in_23), .Y(g7540));
CLKBUFX1 gbuf_d_24(.A(n_6353), .Y(d_out_24));
CLKBUFX1 gbuf_q_24(.A(q_in_24), .Y(g8358));
CLKBUFX1 gbuf_d_25(.A(n_6352), .Y(d_out_25));
CLKBUFX1 gbuf_q_25(.A(q_in_25), .Y(g2902));
OAI21X1 g61017(.A0 (g4501), .A1 (n_6334), .B0 (n_6299), .Y (n_6356));
CLKBUFX1 gbuf_d_26(.A(n_6347), .Y(d_out_26));
CLKBUFX1 gbuf_qn_26(.A(qn_in_26), .Y(g_5342));
NAND2X1 g61308(.A (n_6345), .B (n_6346), .Y (n_6355));
MX2X1 g61137(.A (g_10092), .B (n_2648), .S0 (n_9000), .Y (n_6353));
MX2X1 g61168(.A (g2970), .B (n_6336), .S0 (n_9359), .Y (n_6352));
CLKBUFX1 gbuf_d_27(.A(n_6342), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(g4242));
OAI21X1 g61078(.A0 (g4567), .A1 (n_6364), .B0 (n_6297), .Y (n_6351));
OAI22X1 g61330(.A0 (g_8657), .A1 (n_9269), .B0 (g_12275), .B1(n_9830), .Y (n_6348));
NAND2X1 g61367(.A (n_6338), .B (n_6332), .Y (n_6347));
NAND2X1 g61368(.A (g_12275), .B (n_30), .Y (n_6366));
NAND3X1 g61384(.A (n_2221), .B (n_6454), .C (n_10310), .Y (n_6346));
CLKBUFX1 gbuf_d_28(.A(n_6337), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(g_15801));
CLKBUFX1 gbuf_d_29(.A(n_6339), .Y(d_out_29));
CLKBUFX1 gbuf_qn_29(.A(qn_in_29), .Y(g_20909));
AOI22X1 g61383(.A0 (n_2554), .A1 (n_10306), .B0 (n_6331), .B1(n_9526), .Y (n_6345));
CLKBUFX1 gbuf_d_30(.A(n_6335), .Y(d_out_30));
CLKBUFX1 gbuf_qn_30(.A(qn_in_30), .Y(g4501));
OAI22X1 g61329(.A0 (n_6330), .A1 (n_9599), .B0 (g4235), .B1 (n_9862),.Y (n_6342));
CLKBUFX1 gbuf_d_31(.A(n_6323), .Y(d_out_31));
CLKBUFX1 gbuf_qn_31(.A(qn_in_31), .Y(g_12275));
NAND2X1 g61400(.A (n_6317), .B (n_6326), .Y (n_6339));
CLKBUFX1 gbuf_d_32(.A(n_6321), .Y(d_out_32));
CLKBUFX1 gbuf_qn_32(.A(qn_in_32), .Y(g4567));
AOI21X1 g61432(.A0 (n_6324), .A1 (n_9856), .B0 (n_6328), .Y (n_6338));
CLKBUFX1 gbuf_d_33(.A(n_10715), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(g_10092));
MX2X1 g61224(.A (g_19459), .B (n_6316), .S0 (n_9834), .Y (n_6337));
NAND3X1 g61259(.A (n_6318), .B (n_11055), .C (n_3765), .Y (n_6336));
CLKBUFX1 gbuf_d_34(.A(n_6327), .Y(d_out_34));
CLKBUFX1 gbuf_qn_34(.A(qn_in_34), .Y(g_17086));
OAI21X1 g61131(.A0 (g4498), .A1 (n_6334), .B0 (n_6254), .Y (n_6335));
NAND4X1 g61431(.A (n_10315), .B (n_10310), .C (n_9651), .D (n_6331),.Y (n_6332));
XOR2X1 g61434(.A (n_4247), .B (n_6310), .Y (n_6330));
NOR2X1 g61465(.A (n_1865), .B (n_10315), .Y (n_6328));
NAND2X1 g61475(.A (n_6312), .B (n_6309), .Y (n_6327));
NAND3X1 g61477(.A (n_7395), .B (n_6468), .C (n_6324), .Y (n_6326));
OAI22X1 g61483(.A0 (n_6306), .A1 (n_9193), .B0 (g_18980), .B1(n_9698), .Y (n_6323));
OAI21X1 g61221(.A0 (g4543), .A1 (n_6364), .B0 (n_6320), .Y (n_6321));
CLKBUFX1 gbuf_d_35(.A(n_6313), .Y(d_out_35));
CLKBUFX1 gbuf_q_35(.A(q_in_35), .Y(g_16464));
NOR2X1 g61306(.A (n_6315), .B (n_6958), .Y (n_6318));
AOI22X1 g61481(.A0 (n_2311), .A1 (n_6621), .B0 (n_6308), .B1(n_9697), .Y (n_6317));
CLKBUFX1 gbuf_d_36(.A(n_6311), .Y(d_out_36));
CLKBUFX1 gbuf_qn_36(.A(qn_in_36), .Y(g_16769));
NAND2X1 g61305(.A (g_19913), .B (n_32), .Y (n_6316));
INVX1 g61363(.A (g_19913), .Y (n_6315));
NAND2X1 g61497(.A (n_6290), .B (n_6302), .Y (n_6313));
AOI21X1 g61518(.A0 (g_16464), .A1 (n_9019), .B0 (n_6305), .Y(n_6312));
CLKBUFX1 gbuf_d_37(.A(n_6300), .Y(d_out_37));
CLKBUFX1 gbuf_qn_37(.A(qn_in_37), .Y(g4498));
CLKBUFX1 gbuf_d_38(.A(n_6303), .Y(d_out_38));
CLKBUFX1 gbuf_q_38(.A(q_in_38), .Y(g_21799));
CLKBUFX1 gbuf_d_39(.A(n_6301), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(g21176));
CLKBUFX1 gbuf_d_40(.A(n_6295), .Y(d_out_40));
CLKBUFX1 gbuf_qn_40(.A(qn_in_40), .Y(g_19913));
NAND2X2 g61373(.A (n_6285), .B (n_6296), .Y (n_6311));
NAND2X1 g61504(.A (n_6258), .B (n_6288), .Y (n_6310));
NAND3X1 g61512(.A (n_7402), .B (n_6304), .C (n_6308), .Y (n_6309));
AOI21X1 g61547(.A0 (n_6208), .A1 (n_6280), .B0 (n_6286), .Y (n_6306));
CLKBUFX1 gbuf_d_41(.A(n_8605), .Y(d_out_41));
CLKBUFX1 gbuf_qn_41(.A(qn_in_41), .Y(g3106));
CLKBUFX1 gbuf_d_42(.A(n_7133), .Y(d_out_42));
CLKBUFX1 gbuf_qn_42(.A(qn_in_42), .Y(g3457));
CLKBUFX1 gbuf_d_43(.A(n_6878), .Y(d_out_43));
CLKBUFX1 gbuf_qn_43(.A(qn_in_43), .Y(g3808));
CLKBUFX1 gbuf_d_44(.A(n_6287), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(g2799));
CLKBUFX1 gbuf_d_45(.A(n_6298), .Y(d_out_45));
CLKBUFX1 gbuf_qn_45(.A(qn_in_45), .Y(g4543));
NOR3X1 g61536(.A (n_6304), .B (n_6308), .C (n_10078), .Y (n_6305));
NAND2X1 g61544(.A (n_6282), .B (n_6271), .Y (n_6303));
NAND3X1 g61546(.A (n_7395), .B (n_8819), .C (g_16464), .Y (n_6302));
OAI21X1 g61587(.A0 (n_9501), .A1 (n_101), .B0 (n_6281), .Y (n_6301));
OAI21X1 g61261(.A0 (g4495), .A1 (n_6334), .B0 (n_6299), .Y (n_6300));
CLKBUFX1 gbuf_d_46(.A(n_6283), .Y(d_out_46));
CLKBUFX1 gbuf_q_46(.A(q_in_46), .Y(g_15879));
OAI21X1 g61382(.A0 (g4540), .A1 (n_6364), .B0 (n_6297), .Y (n_6298));
NAND3X1 g61401(.A (n_6274), .B (n_2290), .C (n_9398), .Y (n_6296));
AOI21X1 g61402(.A0 (n_6264), .A1 (n_10005), .B0 (g_16769), .Y(n_6295));
AOI22X1 g61549(.A0 (n_2248), .A1 (n_11138), .B0 (g_21799), .B1(n_9193), .Y (n_6290));
OR4X1 g61552(.A (n_6267), .B (g8917), .C (g8915), .D (g8916), .Y(n_6288));
OAI21X1 g61567(.A0 (n_5610), .A1 (n_5761), .B0 (n_6266), .Y (n_6287));
NAND2X1 g61573(.A (n_5520), .B (n_6265), .Y (n_6286));
CLKBUFX1 gbuf_d_47(.A(n_6275), .Y(d_out_47));
CLKBUFX1 gbuf_qn_47(.A(qn_in_47), .Y(g_18590));
CLKBUFX1 gbuf_d_48(.A(n_6279), .Y(d_out_48));
CLKBUFX1 gbuf_q_48(.A(q_in_48), .Y(g_18793));
AOI22X1 g61427(.A0 (n_2291), .A1 (n_6798), .B0 (n_6252), .B1(n_9193), .Y (n_6285));
INVX1 g61569(.A (n_6620), .Y (n_6304));
NAND2X1 g61574(.A (n_6240), .B (n_6259), .Y (n_6283));
AOI21X1 g61591(.A0 (g_15879), .A1 (n_9431), .B0 (n_6262), .Y(n_6282));
OR4X1 g61649(.A (n_6280), .B (g_6192), .C (n_9599), .D (g_18980), .Y(n_6281));
CLKBUFX1 gbuf_d_49(.A(n_6260), .Y(d_out_49));
CLKBUFX1 gbuf_q_49(.A(q_in_49), .Y(g_10903));
CLKBUFX1 gbuf_d_50(.A(n_6255), .Y(d_out_50));
CLKBUFX1 gbuf_qn_50(.A(qn_in_50), .Y(g4495));
NAND3X1 g61449(.A (n_4252), .B (n_6218), .C (n_4025), .Y (n_6279));
NAND2X1 g61468(.A (n_6220), .B (n_6253), .Y (n_6275));
NOR2X1 g61471(.A (n_6153), .B (n_6798), .Y (n_6274));
NAND3X1 g61585(.A (n_7395), .B (n_8821), .C (g_21799), .Y (n_6271));
OR2X1 g61642(.A (n_6239), .B (n_6093), .Y (n_6267));
AOI22X1 g61645(.A0 (g2799), .A1 (n_5675), .B0 (n_9599), .B1 (g20654),.Y (n_6266));
NAND4X1 g61648(.A (g_19187), .B (g_18980), .C (g_16983), .D (n_3519),.Y (n_6265));
CLKBUFX1 gbuf_d_51(.A(n_6257), .Y(d_out_51));
CLKBUFX1 gbuf_qn_51(.A(qn_in_51), .Y(g_22605));
CLKBUFX1 gbuf_d_52(.A(n_6247), .Y(d_out_52));
CLKBUFX1 gbuf_qn_52(.A(qn_in_52), .Y(g3333));
CLKBUFX1 gbuf_d_53(.A(n_6246), .Y(d_out_53));
CLKBUFX1 gbuf_qn_53(.A(qn_in_53), .Y(g3684));
CLKBUFX1 gbuf_d_54(.A(n_6241), .Y(d_out_54));
CLKBUFX1 gbuf_qn_54(.A(qn_in_54), .Y(g4035));
CLKBUFX1 gbuf_d_55(.A(n_6256), .Y(d_out_55));
CLKBUFX1 gbuf_qn_55(.A(qn_in_55), .Y(g1768));
CLKBUFX1 gbuf_d_56(.A(n_6221), .Y(d_out_56));
CLKBUFX1 gbuf_qn_56(.A(qn_in_56), .Y(g4540));
INVX1 g61506(.A (n_6798), .Y (n_6264));
NOR3X1 g61627(.A (n_8821), .B (g_21799), .C (n_9772), .Y (n_6262));
NAND2X1 g61639(.A (n_6214), .B (n_6149), .Y (n_6260));
NAND3X1 g61641(.A (n_7402), .B (n_8820), .C (g_15879), .Y (n_6259));
XOR2X1 g61651(.A (g8870), .B (g4235), .Y (n_6258));
CLKBUFX1 gbuf_d_57(.A(gbuf1), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(g4483));
CLKBUFX1 gbuf_d_58(.A(n_6217), .Y(d_out_58));
CLKBUFX1 gbuf_q_58(.A(q_in_58), .Y(g12923));
CLKBUFX1 gbuf_d_59(.A(n_6235), .Y(d_out_59));
CLKBUFX1 gbuf_qn_59(.A(qn_in_59), .Y(g2661));
CLKBUFX1 gbuf_d_60(.A(n_6234), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(g2685));
CLKBUFX1 gbuf_d_61(.A(n_6232), .Y(d_out_61));
CLKBUFX1 gbuf_q_61(.A(q_in_61), .Y(g1724));
CLKBUFX1 gbuf_d_62(.A(n_6230), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(g1830));
CLKBUFX1 gbuf_d_63(.A(n_6238), .Y(d_out_63));
CLKBUFX1 gbuf_qn_63(.A(qn_in_63), .Y(g1902));
CLKBUFX1 gbuf_d_64(.A(n_6229), .Y(d_out_64));
CLKBUFX1 gbuf_q_64(.A(q_in_64), .Y(g1964));
CLKBUFX1 gbuf_d_65(.A(n_6228), .Y(d_out_65));
CLKBUFX1 gbuf_qn_65(.A(qn_in_65), .Y(g2102));
CLKBUFX1 gbuf_d_66(.A(n_6226), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(g2126));
CLKBUFX1 gbuf_d_67(.A(n_6225), .Y(d_out_67));
CLKBUFX1 gbuf_qn_67(.A(qn_in_67), .Y(g2259));
CLKBUFX1 gbuf_d_68(.A(n_6224), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(g2283));
CLKBUFX1 gbuf_d_69(.A(n_6237), .Y(d_out_69));
CLKBUFX1 gbuf_qn_69(.A(qn_in_69), .Y(g2327));
CLKBUFX1 gbuf_d_70(.A(n_6223), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(g2389));
CLKBUFX1 gbuf_d_71(.A(n_6233), .Y(d_out_71));
CLKBUFX1 gbuf_qn_71(.A(qn_in_71), .Y(g1700));
CLKBUFX1 gbuf_d_72(.A(n_6222), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(g2523));
CLKBUFX1 gbuf_d_73(.A(n_6236), .Y(d_out_73));
CLKBUFX1 gbuf_qn_73(.A(qn_in_73), .Y(g2461));
NAND2X2 g61375(.A (n_6091), .B (n_6927), .Y (n_6257));
NAND3X1 g61922(.A (n_6156), .B (n_2551), .C (n_6066), .Y (n_6256));
OAI21X1 g61405(.A0 (g4480), .A1 (n_6364), .B0 (n_6254), .Y (n_6255));
NAND3X1 g61505(.A (n_6154), .B (n_6252), .C (n_9425), .Y (n_6253));
MX2X1 g61519(.A (g3263), .B (n_6100), .S0 (n_9218), .Y (n_6247));
MX2X1 g61520(.A (g3614), .B (n_6098), .S0 (n_9000), .Y (n_6246));
MX2X1 g61556(.A (g3965), .B (n_6096), .S0 (n_9000), .Y (n_6241));
AOI22X1 g61647(.A0 (n_2250), .A1 (n_6211), .B0 (g_10903), .B1(n_9491), .Y (n_6240));
CLKBUFX1 gbuf_d_74(.A(n_6155), .Y(d_out_74));
CLKBUFX1 gbuf_qn_74(.A(qn_in_74), .Y(g_9176));
CLKBUFX1 gbuf_d_75(.A(n_6150), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(g_18112));
CLKBUFX1 gbuf_d_76(.A(n_6206), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(g2657));
CLKBUFX1 gbuf_d_77(.A(n_6203), .Y(d_out_77));
CLKBUFX1 gbuf_qn_77(.A(qn_in_77), .Y(g2681));
CLKBUFX1 gbuf_d_78(.A(n_6204), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(g1696));
CLKBUFX1 gbuf_d_79(.A(n_6202), .Y(d_out_79));
CLKBUFX1 gbuf_qn_79(.A(qn_in_79), .Y(g1720));
CLKBUFX1 gbuf_d_80(.A(n_6201), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(g1760));
CLKBUFX1 gbuf_d_81(.A(n_6199), .Y(d_out_81));
CLKBUFX1 gbuf_qn_81(.A(qn_in_81), .Y(g1834));
CLKBUFX1 gbuf_d_82(.A(n_6198), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(g1858));
CLKBUFX1 gbuf_d_83(.A(n_6197), .Y(d_out_83));
CLKBUFX1 gbuf_q_83(.A(q_in_83), .Y(g1894));
CLKBUFX1 gbuf_d_84(.A(n_6194), .Y(d_out_84));
CLKBUFX1 gbuf_qn_84(.A(qn_in_84), .Y(g1968));
CLKBUFX1 gbuf_d_85(.A(n_6176), .Y(d_out_85));
CLKBUFX1 gbuf_q_85(.A(q_in_85), .Y(g2028));
CLKBUFX1 gbuf_d_86(.A(n_6190), .Y(d_out_86));
CLKBUFX1 gbuf_q_86(.A(q_in_86), .Y(g2098));
CLKBUFX1 gbuf_d_87(.A(n_6192), .Y(d_out_87));
CLKBUFX1 gbuf_q_87(.A(q_in_87), .Y(g1992));
CLKBUFX1 gbuf_d_88(.A(n_6189), .Y(d_out_88));
CLKBUFX1 gbuf_qn_88(.A(qn_in_88), .Y(g2122));
CLKBUFX1 gbuf_d_89(.A(n_6174), .Y(d_out_89));
CLKBUFX1 gbuf_q_89(.A(q_in_89), .Y(g2185));
CLKBUFX1 gbuf_d_90(.A(n_6210), .Y(d_out_90));
CLKBUFX1 gbuf_qn_90(.A(qn_in_90), .Y(g2193));
CLKBUFX1 gbuf_d_91(.A(n_6188), .Y(d_out_91));
CLKBUFX1 gbuf_q_91(.A(q_in_91), .Y(g2255));
CLKBUFX1 gbuf_d_92(.A(n_6186), .Y(d_out_92));
CLKBUFX1 gbuf_qn_92(.A(qn_in_92), .Y(g2279));
CLKBUFX1 gbuf_d_93(.A(n_6185), .Y(d_out_93));
CLKBUFX1 gbuf_q_93(.A(q_in_93), .Y(g2319));
CLKBUFX1 gbuf_d_94(.A(n_6184), .Y(d_out_94));
CLKBUFX1 gbuf_qn_94(.A(qn_in_94), .Y(g2393));
CLKBUFX1 gbuf_d_95(.A(n_6183), .Y(d_out_95));
CLKBUFX1 gbuf_q_95(.A(q_in_95), .Y(g2417));
CLKBUFX1 gbuf_d_96(.A(n_6182), .Y(d_out_96));
CLKBUFX1 gbuf_q_96(.A(q_in_96), .Y(g2453));
CLKBUFX1 gbuf_d_97(.A(n_6180), .Y(d_out_97));
CLKBUFX1 gbuf_qn_97(.A(qn_in_97), .Y(g2527));
CLKBUFX1 gbuf_d_98(.A(n_6178), .Y(d_out_98));
CLKBUFX1 gbuf_q_98(.A(q_in_98), .Y(g2551));
CLKBUFX1 gbuf_d_99(.A(n_6171), .Y(d_out_99));
CLKBUFX1 gbuf_q_99(.A(q_in_99), .Y(g1624));
CLKBUFX1 gbuf_d_100(.A(n_6209), .Y(d_out_100));
CLKBUFX1 gbuf_qn_100(.A(qn_in_100), .Y(g1632));
CLKBUFX1 gbuf_d_101(.A(n_6169), .Y(d_out_101));
CLKBUFX1 gbuf_q_101(.A(q_in_101), .Y(g2587));
CLKBUFX1 gbuf_d_102(.A(n_6165), .Y(d_out_102));
CLKBUFX1 gbuf_q_102(.A(q_in_102), .Y(n_5996));
CLKBUFX1 gbuf_d_103(.A(n_6166), .Y(d_out_103));
CLKBUFX1 gbuf_q_103(.A(q_in_103), .Y(g1792));
CLKBUFX1 gbuf_d_104(.A(n_6164), .Y(d_out_104));
CLKBUFX1 gbuf_q_104(.A(q_in_104), .Y(g1811));
CLKBUFX1 gbuf_d_105(.A(n_6162), .Y(d_out_105));
CLKBUFX1 gbuf_q_105(.A(q_in_105), .Y(n_5925));
CLKBUFX1 gbuf_d_106(.A(n_6168), .Y(d_out_106));
CLKBUFX1 gbuf_qn_106(.A(qn_in_106), .Y(g2036));
CLKBUFX1 gbuf_d_107(.A(n_6161), .Y(d_out_107));
CLKBUFX1 gbuf_q_107(.A(q_in_107), .Y(n_5917));
CLKBUFX1 gbuf_d_108(.A(n_6160), .Y(d_out_108));
CLKBUFX1 gbuf_q_108(.A(q_in_108), .Y(n_5921));
CLKBUFX1 gbuf_d_109(.A(n_6167), .Y(d_out_109));
CLKBUFX1 gbuf_qn_109(.A(qn_in_109), .Y(g2595));
CLKBUFX1 gbuf_d_110(.A(n_6157), .Y(d_out_110));
CLKBUFX1 gbuf_qn_110(.A(qn_in_110), .Y(g1825));
NAND2X1 g61732(.A (n_6207), .B (g4235), .Y (n_6239));
NAND3X1 g61802(.A (n_6065), .B (n_2307), .C (n_6092), .Y (n_6238));
NAND3X1 g61811(.A (n_6064), .B (n_2294), .C (n_6087), .Y (n_6237));
NAND3X1 g61818(.A (n_6062), .B (n_2781), .C (n_6086), .Y (n_6236));
MX2X1 g61845(.A (g2657), .B (n_6078), .S0 (n_8955), .Y (n_6235));
OAI22X1 g61848(.A0 (n_6082), .A1 (n_9976), .B0 (g2681), .B1 (n_9992),.Y (n_6234));
MX2X1 g61849(.A (g1696), .B (n_6070), .S0 (n_9172), .Y (n_6233));
OAI22X1 g61850(.A0 (n_6080), .A1 (n_9976), .B0 (g1720), .B1 (n_9992),.Y (n_6232));
MX2X1 g61853(.A (n_827), .B (n_6074), .S0 (n_8955), .Y (n_6230));
MX2X1 g61858(.A (n_836), .B (n_6073), .S0 (n_9240), .Y (n_6229));
MX2X1 g61863(.A (g2098), .B (n_6076), .S0 (n_9240), .Y (n_6228));
OAI22X1 g61865(.A0 (n_6081), .A1 (n_9269), .B0 (g2122), .B1 (n_9209),.Y (n_6226));
MX2X1 g61867(.A (g2255), .B (n_6068), .S0 (n_9750), .Y (n_6225));
OAI22X1 g61869(.A0 (n_6079), .A1 (n_9193), .B0 (g2279), .B1 (n_9830),.Y (n_6224));
MX2X1 g61871(.A (n_831), .B (n_6072), .S0 (n_9256), .Y (n_6223));
MX2X1 g61877(.A (n_839), .B (n_6071), .S0 (n_9359), .Y (n_6222));
NAND3X1 g61514(.A (n_6320), .B (n_3996), .C (n_6011), .Y (n_6221));
AOI22X1 g61516(.A0 (n_2308), .A1 (n_6562), .B0 (n_6057), .B1(n_9193), .Y (n_6220));
OR2X1 g61535(.A (n_6216), .B (n_10687), .Y (n_6218));
OAI21X1 g61551(.A0 (n_392), .A1 (n_9425), .B0 (n_6216), .Y (n_6217));
CLKBUFX1 gbuf_d_111(.A(n_6142), .Y(d_out_111));
CLKBUFX1 gbuf_qn_111(.A(qn_in_111), .Y(g1854));
CLKBUFX1 gbuf_d_112(.A(n_6143), .Y(d_out_112));
CLKBUFX1 gbuf_q_112(.A(q_in_112), .Y(g_13871));
CLKBUFX1 gbuf_d_113(.A(n_6141), .Y(d_out_113));
CLKBUFX1 gbuf_qn_113(.A(qn_in_113), .Y(g1988));
CLKBUFX1 gbuf_d_114(.A(n_6140), .Y(d_out_114));
CLKBUFX1 gbuf_qn_114(.A(qn_in_114), .Y(g2413));
CLKBUFX1 gbuf_d_115(.A(n_6138), .Y(d_out_115));
CLKBUFX1 gbuf_qn_115(.A(qn_in_115), .Y(g2547));
CLKBUFX1 gbuf_d_116(.A(n_6133), .Y(d_out_116));
CLKBUFX1 gbuf_q_116(.A(q_in_116), .Y(g1926));
CLKBUFX1 gbuf_d_117(.A(n_6132), .Y(d_out_117));
CLKBUFX1 gbuf_q_117(.A(q_in_117), .Y(g1945));
CLKBUFX1 gbuf_d_118(.A(n_6134), .Y(d_out_118));
CLKBUFX1 gbuf_q_118(.A(q_in_118), .Y(g21270));
CLKBUFX1 gbuf_d_119(.A(n_6130), .Y(d_out_119));
CLKBUFX1 gbuf_q_119(.A(q_in_119), .Y(n_5932));
CLKBUFX1 gbuf_d_120(.A(n_6126), .Y(d_out_120));
CLKBUFX1 gbuf_q_120(.A(q_in_120), .Y(n_5941));
CLKBUFX1 gbuf_d_121(.A(n_6125), .Y(d_out_121));
CLKBUFX1 gbuf_q_121(.A(q_in_121), .Y(g2217));
CLKBUFX1 gbuf_d_122(.A(n_6123), .Y(d_out_122));
CLKBUFX1 gbuf_q_122(.A(q_in_122), .Y(g2236));
CLKBUFX1 gbuf_d_123(.A(n_6129), .Y(d_out_123));
CLKBUFX1 gbuf_q_123(.A(q_in_123), .Y(g2060));
CLKBUFX1 gbuf_d_124(.A(n_6121), .Y(d_out_124));
CLKBUFX1 gbuf_q_124(.A(q_in_124), .Y(g2351));
CLKBUFX1 gbuf_d_125(.A(n_6120), .Y(d_out_125));
CLKBUFX1 gbuf_q_125(.A(q_in_125), .Y(g2370));
CLKBUFX1 gbuf_d_126(.A(n_6128), .Y(d_out_126));
CLKBUFX1 gbuf_q_126(.A(q_in_126), .Y(g2079));
CLKBUFX1 gbuf_d_127(.A(n_6118), .Y(d_out_127));
CLKBUFX1 gbuf_q_127(.A(q_in_127), .Y(g2485));
CLKBUFX1 gbuf_d_128(.A(n_6117), .Y(d_out_128));
CLKBUFX1 gbuf_q_128(.A(q_in_128), .Y(g2504));
CLKBUFX1 gbuf_d_129(.A(n_6116), .Y(d_out_129));
CLKBUFX1 gbuf_q_129(.A(q_in_129), .Y(n_5936));
CLKBUFX1 gbuf_d_130(.A(n_6114), .Y(d_out_130));
CLKBUFX1 gbuf_q_130(.A(q_in_130), .Y(g1657));
CLKBUFX1 gbuf_d_131(.A(n_6112), .Y(d_out_131));
CLKBUFX1 gbuf_q_131(.A(q_in_131), .Y(n_5928));
CLKBUFX1 gbuf_d_132(.A(n_6110), .Y(d_out_132));
CLKBUFX1 gbuf_q_132(.A(q_in_132), .Y(g2619));
CLKBUFX1 gbuf_d_133(.A(n_6109), .Y(d_out_133));
CLKBUFX1 gbuf_q_133(.A(q_in_133), .Y(g2638));
CLKBUFX1 gbuf_d_134(.A(n_6111), .Y(d_out_134));
CLKBUFX1 gbuf_q_134(.A(q_in_134), .Y(g1677));
CLKBUFX1 gbuf_d_135(.A(n_6101), .Y(d_out_135));
CLKBUFX1 gbuf_q_135(.A(q_in_135), .Y(g2652));
CLKBUFX1 gbuf_d_136(.A(n_6108), .Y(d_out_136));
CLKBUFX1 gbuf_q_136(.A(q_in_136), .Y(g1691));
CLKBUFX1 gbuf_d_137(.A(n_6107), .Y(d_out_137));
CLKBUFX1 gbuf_qn_137(.A(qn_in_137), .Y(g1959));
CLKBUFX1 gbuf_d_138(.A(n_6102), .Y(d_out_138));
CLKBUFX1 gbuf_q_138(.A(q_in_138), .Y(g2093));
CLKBUFX1 gbuf_d_139(.A(n_6105), .Y(d_out_139));
CLKBUFX1 gbuf_q_139(.A(q_in_139), .Y(g2250));
CLKBUFX1 gbuf_d_140(.A(n_6104), .Y(d_out_140));
CLKBUFX1 gbuf_qn_140(.A(qn_in_140), .Y(g2384));
CLKBUFX1 gbuf_d_141(.A(n_6103), .Y(d_out_141));
CLKBUFX1 gbuf_qn_141(.A(qn_in_141), .Y(g2518));
CLKBUFX1 gbuf_d_142(.A(g4519), .Y(d_out_142));
CLKBUFX1 gbuf_q_142(.A(q_in_142), .Y(gbuf1));
AOI21X1 g61743(.A0 (g_18112), .A1 (n_9419), .B0 (n_6146), .Y(n_6214));
CLKBUFX1 gbuf_d_143(.A(n_6136), .Y(d_out_143));
CLKBUFX1 gbuf_q_143(.A(q_in_143), .Y(g20654));
CLKBUFX1 gbuf_d_144(.A(n_6137), .Y(d_out_144));
CLKBUFX1 gbuf_qn_144(.A(qn_in_144), .Y(g_18980));
NAND3X1 g61808(.A (n_6010), .B (n_2259), .C (n_6044), .Y (n_6210));
NAND3X1 g61820(.A (n_6009), .B (n_2522), .C (n_6043), .Y (n_6209));
OAI21X1 g61832(.A0 (g_19304), .A1 (g_16983), .B0 (g_19187), .Y(n_6208));
NOR2X1 g61835(.A (g11770), .B (g8920), .Y (n_6207));
MX2X1 g61844(.A (g2652), .B (n_6024), .S0 (n_9311), .Y (n_6206));
MX2X1 g61846(.A (g1691), .B (n_6030), .S0 (n_9156), .Y (n_6204));
MX2X1 g61847(.A (n_6020), .B (n_6021), .S0 (n_9172), .Y (n_6203));
MX2X1 g61851(.A (n_6027), .B (n_6028), .S0 (n_9000), .Y (n_6202));
OAI22X1 g61852(.A0 (n_6042), .A1 (n_9269), .B0 (g1768), .B1 (n_9627),.Y (n_6201));
MX2X1 g61854(.A (g1830), .B (n_6016), .S0 (n_9234), .Y (n_6199));
OAI22X1 g61855(.A0 (n_6038), .A1 (n_10952), .B0 (g1854), .B1(n_9311), .Y (n_6198));
OAI22X1 g61857(.A0 (n_6041), .A1 (n_9599), .B0 (g1902), .B1(n_10063), .Y (n_6197));
MX2X1 g61859(.A (g1964), .B (n_6015), .S0 (n_9834), .Y (n_6194));
OAI22X1 g61861(.A0 (n_6037), .A1 (n_9976), .B0 (g1988), .B1 (n_9862),.Y (n_6192));
MX2X1 g61862(.A (g2093), .B (n_6019), .S0 (n_9172), .Y (n_6190));
MX2X1 g61864(.A (n_6017), .B (n_6018), .S0 (n_9091), .Y (n_6189));
MX2X1 g61866(.A (g2250), .B (n_6029), .S0 (n_9256), .Y (n_6188));
MX2X1 g61868(.A (n_6025), .B (n_6026), .S0 (n_9000), .Y (n_6186));
OAI22X1 g61870(.A0 (n_6040), .A1 (n_9884), .B0 (g2327), .B1 (n_9830),.Y (n_6185));
MX2X1 g61872(.A (g2389), .B (n_6014), .S0 (n_9156), .Y (n_6184));
OAI22X1 g61874(.A0 (n_6034), .A1 (n_9461), .B0 (g2413), .B1(n_10063), .Y (n_6183));
OAI22X1 g61875(.A0 (n_6039), .A1 (n_9772), .B0 (g2461), .B1(n_10005), .Y (n_6182));
MX2X1 g61878(.A (g2523), .B (n_6013), .S0 (n_9797), .Y (n_6180));
OAI22X1 g61880(.A0 (n_6033), .A1 (n_9431), .B0 (g2547), .B1 (n_9811),.Y (n_6178));
OAI22X1 g61881(.A0 (n_6036), .A1 (n_9976), .B0 (g2036), .B1 (n_9627),.Y (n_6176));
OAI22X1 g61882(.A0 (n_6035), .A1 (n_9976), .B0 (g2193), .B1 (n_9651),.Y (n_6174));
OAI22X1 g61883(.A0 (n_6032), .A1 (n_9772), .B0 (g1632), .B1 (n_9862),.Y (n_6171));
OAI22X1 g61884(.A0 (n_6031), .A1 (n_9772), .B0 (g2595), .B1 (n_9811),.Y (n_6169));
NAND3X1 g61924(.A (n_6089), .B (n_2795), .C (n_5956), .Y (n_6168));
NAND3X1 g61936(.A (n_6084), .B (n_2254), .C (n_5951), .Y (n_6167));
MX2X1 g61973(.A (g1798), .B (n_5997), .S0 (n_9894), .Y (n_6166));
MX2X1 g61974(.A (g1760), .B (n_5999), .S0 (n_9469), .Y (n_6165));
MX2X1 g61975(.A (g1792), .B (n_6000), .S0 (n_9425), .Y (n_6164));
MX2X1 g61976(.A (g1894), .B (n_6002), .S0 (n_9091), .Y (n_6162));
MX2X1 g61986(.A (g2319), .B (n_5995), .S0 (n_9469), .Y (n_6161));
MX2X1 g61989(.A (g2453), .B (n_6001), .S0 (n_9091), .Y (n_6160));
OAI21X1 g62028(.A0 (n_2464), .A1 (n_5849), .B0 (n_6061), .Y (n_6157));
NAND3X1 g62054(.A (n_3948), .B (n_5993), .C (n_9501), .Y (n_6156));
NAND2X1 g61541(.A (n_6003), .B (n_6058), .Y (n_6155));
NOR2X1 g61542(.A (n_6153), .B (n_6562), .Y (n_6154));
CLKBUFX1 gbuf_d_145(.A(n_6050), .Y(d_out_145));
CLKBUFX1 gbuf_q_145(.A(q_in_145), .Y(g4527));
NAND2X1 g61720(.A (n_6094), .B (n_6048), .Y (n_6150));
NAND3X1 g61731(.A (n_7395), .B (n_6145), .C (g_10903), .Y (n_6149));
CLKBUFX1 gbuf_d_146(.A(g8920), .Y(d_out_146));
CLKBUFX1 gbuf_qn_146(.A(qn_in_146), .Y(g4235));
INVX1 g61798(.A (n_8820), .Y (n_6211));
NOR3X1 g61803(.A (n_6145), .B (g_10903), .C (n_9772), .Y (n_6146));
NAND2X1 g61824(.A (n_6045), .B (n_5988), .Y (n_6143));
MX2X1 g61856(.A (n_5978), .B (n_5979), .S0 (n_8955), .Y (n_6142));
MX2X1 g61860(.A (n_5975), .B (n_5976), .S0 (n_8955), .Y (n_6141));
MX2X1 g61873(.A (n_5972), .B (n_5973), .S0 (n_9091), .Y (n_6140));
MX2X1 g61879(.A (n_5969), .B (n_5970), .S0 (n_9000), .Y (n_6138));
INVX1 g61904(.A (g_19187), .Y (n_6137));
OAI21X1 g61917(.A0 (g23759), .A1 (n_9425), .B0 (n_5795), .Y (n_6136));
OAI21X1 g61932(.A0 (g23652), .A1 (n_9681), .B0 (n_5792), .Y (n_6134));
MX2X1 g61977(.A (g1932), .B (n_5926), .S0 (n_9797), .Y (n_6133));
MX2X1 g61978(.A (g1926), .B (n_5924), .S0 (n_9558), .Y (n_6132));
MX2X1 g61979(.A (g2028), .B (n_5934), .S0 (n_9681), .Y (n_6130));
MX2X1 g61980(.A (g2066), .B (n_5933), .S0 (n_8955), .Y (n_6129));
MX2X1 g61981(.A (g2060), .B (n_5931), .S0 (n_9425), .Y (n_6128));
MX2X1 g61983(.A (g2185), .B (n_5943), .S0 (n_9558), .Y (n_6126));
MX2X1 g61984(.A (g2223), .B (n_5942), .S0 (n_9234), .Y (n_6125));
MX2X1 g61985(.A (g2217), .B (n_5940), .S0 (n_9139), .Y (n_6123));
MX2X1 g61987(.A (g2357), .B (n_5918), .S0 (n_8955), .Y (n_6121));
MX2X1 g61988(.A (g2351), .B (n_5916), .S0 (n_9558), .Y (n_6120));
MX2X1 g61990(.A (g2491), .B (n_5922), .S0 (n_9091), .Y (n_6118));
MX2X1 g61991(.A (g2485), .B (n_5920), .S0 (n_9558), .Y (n_6117));
MX2X1 g61992(.A (g1624), .B (n_5939), .S0 (n_9558), .Y (n_6116));
MX2X1 g61993(.A (g1664), .B (n_5937), .S0 (n_9091), .Y (n_6114));
MX2X1 g61994(.A (g2587), .B (n_5930), .S0 (n_10063), .Y (n_6112));
MX2X1 g61995(.A (g1657), .B (n_5935), .S0 (n_9558), .Y (n_6111));
MX2X1 g61996(.A (g2625), .B (n_5929), .S0 (n_9992), .Y (n_6110));
MX2X1 g61997(.A (g2619), .B (n_5927), .S0 (n_10063), .Y (n_6109));
NAND3X1 g62022(.A (n_5875), .B (n_2523), .C (n_5904), .Y (n_6108));
OAI21X1 g62033(.A0 (n_2463), .A1 (n_5839), .B0 (n_6008), .Y (n_6107));
NAND3X1 g62038(.A (n_5948), .B (n_2537), .C (n_5899), .Y (n_6105));
OAI21X1 g62042(.A0 (n_2461), .A1 (n_5844), .B0 (n_6006), .Y (n_6104));
OAI21X1 g62046(.A0 (n_2460), .A1 (n_5833), .B0 (n_6004), .Y (n_6103));
NAND3X1 g62049(.A (n_5950), .B (n_2419), .C (n_5901), .Y (n_6102));
NAND3X1 g62051(.A (n_5945), .B (n_2524), .C (n_5896), .Y (n_6101));
CLKBUFX1 gbuf_d_147(.A(n_6012), .Y(d_out_147));
CLKBUFX1 gbuf_qn_147(.A(qn_in_147), .Y(g4480));
NOR2X1 g61539(.A (n_6059), .B (n_6005), .Y (n_6320));
NOR2X1 g61540(.A (n_6054), .B (n_6334), .Y (n_6297));
NAND2X1 g61581(.A (g_19492), .B (n_9894), .Y (n_6216));
OAI21X1 g61593(.A0 (n_3775), .A1 (n_7235), .B0 (n_3603), .Y (n_6100));
OAI21X1 g61594(.A0 (n_3779), .A1 (n_8908), .B0 (n_3599), .Y (n_6098));
OAI21X1 g61650(.A0 (n_6243), .A1 (n_6095), .B0 (n_3593), .Y (n_6096));
CLKBUFX1 gbuf_d_148(.A(n_5994), .Y(d_out_148));
CLKBUFX1 gbuf_q_148(.A(q_in_148), .Y(g4515));
CLKBUFX1 gbuf_d_149(.A(n_6046), .Y(d_out_149));
CLKBUFX1 gbuf_q_149(.A(q_in_149), .Y(n_8793));
CLKBUFX1 gbuf_d_150(.A(n_5991), .Y(d_out_150));
CLKBUFX1 gbuf_q_150(.A(q_in_150), .Y(g4519));
AOI22X1 g61840(.A0 (n_2546), .A1 (n_6457), .B0 (g_13871), .B1(n_9193), .Y (n_6094));
CLKBUFX1 gbuf_d_151(.A(g8919), .Y(d_out_151));
CLKBUFX1 gbuf_q_151(.A(q_in_151), .Y(g8920));
CLKBUFX1 gbuf_d_152(.A(n_5986), .Y(d_out_152));
CLKBUFX1 gbuf_qn_152(.A(qn_in_152), .Y(g_19187));
OR2X1 g61944(.A (n_5984), .B (g8919), .Y (n_6093));
NAND3X1 g62055(.A (n_3945), .B (n_5909), .C (n_9811), .Y (n_6092));
NAND3X1 g61466(.A (n_5981), .B (n_10713), .C (n_10063), .Y (n_6091));
NAND3X1 g62057(.A (n_4318), .B (n_5882), .C (n_9425), .Y (n_6089));
NAND3X1 g62067(.A (n_4124), .B (n_5907), .C (n_9698), .Y (n_6087));
NAND3X1 g62070(.A (n_4122), .B (n_5905), .C (n_9698), .Y (n_6086));
NAND3X1 g62072(.A (n_4118), .B (n_5877), .C (n_9359), .Y (n_6084));
AOI21X1 g62081(.A0 (n_10790), .A1 (g2685), .B0 (n_5957), .Y (n_6082));
AOI21X1 g62087(.A0 (n_10995), .A1 (g2126), .B0 (n_5952), .Y (n_6081));
AOI21X1 g62090(.A0 (n_10617), .A1 (g1724), .B0 (n_10618), .Y(n_6080));
AOI21X1 g62091(.A0 (n_6067), .A1 (g2283), .B0 (n_5960), .Y (n_6079));
OAI21X1 g62106(.A0 (n_5958), .A1 (n_10790), .B0 (n_5959), .Y(n_6078));
OAI21X1 g62109(.A0 (n_5953), .A1 (n_10995), .B0 (n_5954), .Y(n_6076));
MX2X1 g62119(.A (g1830), .B (n_828), .S0 (n_5884), .Y (n_6074));
MX2X1 g62121(.A (g1964), .B (n_837), .S0 (n_5883), .Y (n_6073));
MX2X1 g62125(.A (g2389), .B (n_832), .S0 (n_5880), .Y (n_6072));
MX2X1 g62128(.A (g2523), .B (n_840), .S0 (n_5878), .Y (n_6071));
OAI21X1 g62130(.A0 (n_5964), .A1 (n_10617), .B0 (n_5965), .Y(n_6070));
OAI21X1 g62131(.A0 (n_5961), .A1 (n_6067), .B0 (n_5962), .Y (n_6068));
NAND3X1 g62255(.A (n_5992), .B (n_136), .C (n_9750), .Y (n_6066));
NAND3X1 g62256(.A (n_5910), .B (n_67), .C (n_9139), .Y (n_6065));
NAND3X1 g62264(.A (n_5908), .B (n_57), .C (n_9139), .Y (n_6064));
NAND3X1 g62265(.A (n_5906), .B (n_12), .C (n_10063), .Y (n_6062));
AOI22X1 g62270(.A0 (n_2168), .A1 (n_5849), .B0 (g1811), .B1(n_10376), .Y (n_6061));
INVX1 g61576(.A (n_6059), .Y (n_6060));
NAND3X1 g61580(.A (n_5913), .B (n_6057), .C (n_10063), .Y (n_6058));
INVX1 g61578(.A (n_6054), .Y (n_6055));
NOR2X1 g61622(.A (n_6052), .B (n_8908), .Y (n_6248));
NOR2X1 g61621(.A (n_6051), .B (n_6956), .Y (n_6250));
OAI22X1 g60899(.A0 (n_5869), .A1 (n_9976), .B0 (g4521), .B1 (n_9830),.Y (n_6050));
CLKBUFX1 gbuf_d_153(.A(n_5982), .Y(d_out_153));
CLKBUFX1 gbuf_qn_153(.A(qn_in_153), .Y(g_22070));
CLKBUFX1 gbuf_d_154(.A(n_5914), .Y(d_out_154));
CLKBUFX1 gbuf_q_154(.A(q_in_154), .Y(g_16311));
CLKBUFX1 gbuf_d_155(.A(n_5983), .Y(d_out_155));
CLKBUFX1 gbuf_q_155(.A(q_in_155), .Y(g_10556));
CLKBUFX1 gbuf_d_156(.A(n_5985), .Y(d_out_156));
CLKBUFX1 gbuf_q_156(.A(q_in_156), .Y(g_16296));
CLKBUFX1 gbuf_d_157(.A(n_5967), .Y(d_out_157));
CLKBUFX1 gbuf_q_157(.A(q_in_157), .Y(g_19459));
NOR2X1 g61707(.A (n_6049), .B (n_6095), .Y (n_8883));
NAND3X1 g61833(.A (n_7402), .B (n_6715), .C (g_18112), .Y (n_6048));
INVX1 g61919(.A (n_6716), .Y (n_6145));
NAND2X1 g61923(.A (n_5830), .B (n_5889), .Y (n_6046));
AOI21X1 g61961(.A0 (n_8793), .A1 (n_9141), .B0 (n_5891), .Y (n_6045));
NAND3X1 g62059(.A (n_4109), .B (n_5872), .C (n_9091), .Y (n_6044));
NAND3X1 g62071(.A (n_3938), .B (n_5870), .C (n_9811), .Y (n_6043));
AOI22X1 g62083(.A0 (n_1040), .A1 (n_5788), .B0 (n_5818), .B1 (g1760),.Y (n_6042));
AOI22X1 g62084(.A0 (n_1044), .A1 (n_5784), .B0 (n_5816), .B1 (g1894),.Y (n_6041));
AOI22X1 g62088(.A0 (n_1053), .A1 (n_5786), .B0 (n_5817), .B1 (g2319),.Y (n_6040));
AOI22X1 g62089(.A0 (n_1052), .A1 (n_5782), .B0 (n_5815), .B1 (g2453),.Y (n_6039));
AOI21X1 g62092(.A0 (n_5977), .A1 (g1858), .B0 (n_5888), .Y (n_6038));
AOI21X1 g62093(.A0 (n_5974), .A1 (g1992), .B0 (n_5887), .Y (n_6037));
AOI22X1 g62094(.A0 (n_765), .A1 (n_5949), .B0 (n_5809), .B1 (g2028),.Y (n_6036));
AOI22X1 g62095(.A0 (n_775), .A1 (n_5947), .B0 (n_5806), .B1 (g2185),.Y (n_6035));
AOI21X1 g62096(.A0 (n_5971), .A1 (g2417), .B0 (n_5886), .Y (n_6034));
AOI21X1 g62098(.A0 (n_5968), .A1 (g2551), .B0 (n_5885), .Y (n_6033));
AOI22X1 g62099(.A0 (n_769), .A1 (n_5799), .B0 (n_5801), .B1 (g1624),.Y (n_6032));
AOI22X1 g62100(.A0 (n_782), .A1 (n_5944), .B0 (n_5803), .B1 (g2587),.Y (n_6031));
MX2X1 g62107(.A (n_841), .B (g1696), .S0 (n_5800), .Y (n_6030));
MX2X1 g62110(.A (n_833), .B (g2255), .S0 (n_5797), .Y (n_6029));
MX2X1 g62115(.A (n_6027), .B (n_878), .S0 (n_10617), .Y (n_6028));
MX2X1 g62116(.A (n_6025), .B (n_975), .S0 (n_6067), .Y (n_6026));
MX2X1 g62117(.A (n_829), .B (g2657), .S0 (n_5814), .Y (n_6024));
MX2X1 g62118(.A (n_6020), .B (n_852), .S0 (n_10790), .Y (n_6021));
MX2X1 g62123(.A (n_834), .B (g2098), .S0 (n_5807), .Y (n_6019));
MX2X1 g62124(.A (n_6017), .B (n_860), .S0 (n_10995), .Y (n_6018));
XOR2X1 g62133(.A (n_4948), .B (n_5811), .Y (n_6016));
XOR2X1 g62134(.A (n_4946), .B (n_5810), .Y (n_6015));
XOR2X1 g62135(.A (n_4942), .B (n_5805), .Y (n_6014));
XOR2X1 g62136(.A (n_5229), .B (n_5804), .Y (n_6013));
NAND3X1 g61527(.A (n_6011), .B (n_2356), .C (n_6299), .Y (n_6012));
NAND3X1 g62250(.A (n_5873), .B (n_96), .C (n_9139), .Y (n_6010));
NAND3X1 g62252(.A (n_5871), .B (n_105), .C (n_10063), .Y (n_6009));
AOI22X1 g62271(.A0 (n_2212), .A1 (n_5839), .B0 (g1945), .B1 (n_9193),.Y (n_6008));
AOI22X1 g62275(.A0 (n_2229), .A1 (n_5844), .B0 (g2370), .B1 (n_9404),.Y (n_6006));
AND2X1 g61577(.A (g4575), .B (n_6005), .Y (n_6059));
AOI22X1 g62276(.A0 (n_2230), .A1 (n_5833), .B0 (g2504), .B1 (n_9599),.Y (n_6004));
AND2X1 g61579(.A (g4578), .B (n_6005), .Y (n_6054));
AOI22X1 g61589(.A0 (n_2270), .A1 (n_10261), .B0 (g_16311), .B1(n_10376), .Y (n_6003));
MX2X1 g62310(.A (n_5925), .B (g1894), .S0 (n_5784), .Y (n_6002));
CLKBUFX1 gbuf_d_158(.A(n_5879), .Y(d_out_158));
CLKBUFX1 gbuf_q_158(.A(q_in_158), .Y(g_19492));
MX2X1 g62313(.A (n_5921), .B (g2453), .S0 (n_5782), .Y (n_6001));
MX2X1 g62316(.A (g1811), .B (n_2975), .S0 (n_5788), .Y (n_6000));
MX2X1 g62317(.A (n_5996), .B (g1760), .S0 (n_5788), .Y (n_5999));
MX2X1 g62318(.A (g1792), .B (n_5996), .S0 (n_5788), .Y (n_5997));
MX2X1 g62319(.A (n_5917), .B (g2319), .S0 (n_5786), .Y (n_5995));
CLKBUFX1 gbuf_d_159(.A(n_5874), .Y(d_out_159));
CLKBUFX1 gbuf_q_159(.A(q_in_159), .Y(g12919));
CLKBUFX1 gbuf_d_160(.A(n_5868), .Y(d_out_160));
CLKBUFX1 gbuf_q_160(.A(q_in_160), .Y(g2771));
CLKBUFX1 gbuf_d_161(.A(n_5866), .Y(d_out_161));
CLKBUFX1 gbuf_q_161(.A(q_in_161), .Y(g2775));
CLKBUFX1 gbuf_d_162(.A(n_5865), .Y(d_out_162));
CLKBUFX1 gbuf_q_162(.A(q_in_162), .Y(g2783));
CLKBUFX1 gbuf_d_163(.A(n_5863), .Y(d_out_163));
CLKBUFX1 gbuf_q_163(.A(q_in_163), .Y(g2787));
CLKBUFX1 gbuf_d_164(.A(n_5862), .Y(d_out_164));
CLKBUFX1 gbuf_q_164(.A(q_in_164), .Y(g2803));
CLKBUFX1 gbuf_d_165(.A(n_5860), .Y(d_out_165));
CLKBUFX1 gbuf_q_165(.A(q_in_165), .Y(g2807));
CLKBUFX1 gbuf_d_166(.A(n_5859), .Y(d_out_166));
CLKBUFX1 gbuf_q_166(.A(q_in_166), .Y(g2815));
CLKBUFX1 gbuf_d_167(.A(n_5857), .Y(d_out_167));
CLKBUFX1 gbuf_q_167(.A(q_in_167), .Y(g2819));
MX2X1 g60900(.A (g4527), .B (n_5813), .S0 (n_9000), .Y (n_5994));
INVX1 g62591(.A (n_5992), .Y (n_5993));
MX2X1 g60909(.A (g4515), .B (n_5837), .S0 (n_8955), .Y (n_5991));
AND2X1 g61806(.A (n_5781), .B (n_5831), .Y (n_6095));
NAND3X1 g61942(.A (n_7395), .B (n_6524), .C (g_13871), .Y (n_5988));
CLKBUFX1 gbuf_d_168(.A(g8918), .Y(d_out_168));
CLKBUFX1 gbuf_q_168(.A(q_in_168), .Y(g8919));
NAND2X1 g62029(.A (n_5822), .B (n_5573), .Y (n_5986));
NAND2X1 g62048(.A (n_5775), .B (n_5824), .Y (n_5985));
OR2X1 g62060(.A (g8918), .B (g8870), .Y (n_5984));
OAI21X1 g62085(.A0 (n_7094), .A1 (n_9797), .B0 (n_5825), .Y (n_5983));
NAND2X1 g61496(.A (n_5779), .B (n_5828), .Y (n_5982));
NOR2X1 g61501(.A (n_5723), .B (n_7144), .Y (n_5981));
MX2X1 g62120(.A (n_5978), .B (n_883), .S0 (n_5977), .Y (n_5979));
MX2X1 g62122(.A (n_5975), .B (n_885), .S0 (n_5974), .Y (n_5976));
MX2X1 g62126(.A (n_5972), .B (n_866), .S0 (n_5971), .Y (n_5973));
MX2X1 g62129(.A (n_5969), .B (n_858), .S0 (n_5968), .Y (n_5970));
CLKBUFX1 gbuf_d_169(.A(n_5794), .Y(d_out_169));
CLKBUFX1 gbuf_qn_169(.A(qn_in_169), .Y(g23652));
CLKBUFX1 gbuf_d_170(.A(n_5796), .Y(d_out_170));
CLKBUFX1 gbuf_qn_170(.A(qn_in_170), .Y(g23759));
OAI21X1 g63520(.A0 (n_35), .A1 (n_9493), .B0 (n_5820), .Y (n_5967));
NAND2X1 g62218(.A (n_5964), .B (n_10617), .Y (n_5965));
NAND2X1 g62220(.A (n_5961), .B (n_6067), .Y (n_5962));
NOR2X1 g62221(.A (n_976), .B (n_6067), .Y (n_5960));
NAND2X1 g62223(.A (n_5958), .B (n_10790), .Y (n_5959));
NOR2X1 g62224(.A (n_10790), .B (n_10554), .Y (n_5957));
NAND3X1 g62231(.A (n_5881), .B (n_54), .C (n_9425), .Y (n_5956));
NAND2X1 g62232(.A (n_5953), .B (n_10995), .Y (n_5954));
NOR2X1 g62233(.A (n_861), .B (n_10995), .Y (n_5952));
NAND3X1 g62249(.A (n_5876), .B (n_52), .C (n_9811), .Y (n_5951));
NAND3X1 g62258(.A (n_2080), .B (n_5949), .C (n_9501), .Y (n_5950));
NAND3X1 g62261(.A (n_2079), .B (n_5947), .C (n_9698), .Y (n_5948));
NAND3X1 g62266(.A (n_2081), .B (n_5944), .C (n_9425), .Y (n_5945));
MX2X1 g62295(.A (n_5941), .B (g2185), .S0 (n_5947), .Y (n_5943));
MX2X1 g62296(.A (g2217), .B (n_5941), .S0 (n_5947), .Y (n_5942));
MX2X1 g62297(.A (g2236), .B (n_2651), .S0 (n_5947), .Y (n_5940));
MX2X1 g62299(.A (n_5936), .B (g1624), .S0 (n_5799), .Y (n_5939));
MX2X1 g62300(.A (g1657), .B (n_5936), .S0 (n_5799), .Y (n_5937));
MX2X1 g62301(.A (g1677), .B (n_2469), .S0 (n_5799), .Y (n_5935));
MX2X1 g62304(.A (n_5932), .B (g2028), .S0 (n_5949), .Y (n_5934));
MX2X1 g62305(.A (g2060), .B (n_5932), .S0 (n_5949), .Y (n_5933));
MX2X1 g62306(.A (g2079), .B (n_2472), .S0 (n_5949), .Y (n_5931));
MX2X1 g62307(.A (n_5928), .B (g2587), .S0 (n_5944), .Y (n_5930));
MX2X1 g62308(.A (g2619), .B (n_5928), .S0 (n_5944), .Y (n_5929));
MX2X1 g62309(.A (g2638), .B (n_2466), .S0 (n_5944), .Y (n_5927));
MX2X1 g62311(.A (g1926), .B (n_5925), .S0 (n_5784), .Y (n_5926));
MX2X1 g62312(.A (g1945), .B (n_2738), .S0 (n_5784), .Y (n_5924));
MX2X1 g62314(.A (g2485), .B (n_5921), .S0 (n_5782), .Y (n_5922));
MX2X1 g62315(.A (g2504), .B (n_2969), .S0 (n_5782), .Y (n_5920));
MX2X1 g62320(.A (g2351), .B (n_5917), .S0 (n_5786), .Y (n_5918));
MX2X1 g62321(.A (g2370), .B (n_2967), .S0 (n_5786), .Y (n_5916));
NAND2X1 g61632(.A (n_5769), .B (n_5819), .Y (n_5914));
NOR2X1 g61633(.A (n_6153), .B (n_10261), .Y (n_5913));
NAND2X1 g62592(.A (n_5788), .B (n_1667), .Y (n_5992));
INVX1 g62596(.A (n_5909), .Y (n_5910));
INVX1 g62619(.A (n_5907), .Y (n_5908));
INVX1 g62626(.A (n_5905), .Y (n_5906));
NAND3X1 g62647(.A (n_10614), .B (g1691), .C (n_9894), .Y (n_5904));
NAND3X1 g62653(.A (n_5854), .B (g2093), .C (n_9894), .Y (n_5901));
NAND3X1 g62655(.A (n_5852), .B (g2250), .C (n_9139), .Y (n_5899));
NAND3X1 g62661(.A (n_10787), .B (g2652), .C (n_9811), .Y (n_5896));
CLKBUFX1 gbuf_d_171(.A(n_5774), .Y(d_out_171));
CLKBUFX1 gbuf_q_171(.A(q_in_171), .Y(g_6192));
NOR3X1 g62032(.A (n_9461), .B (g_13871), .C (n_6524), .Y (n_5891));
NAND3X1 g62056(.A (n_7395), .B (n_6523), .C (n_8793), .Y (n_5889));
NOR2X1 g62208(.A (n_884), .B (n_5977), .Y (n_5888));
NOR2X1 g62210(.A (n_886), .B (n_5974), .Y (n_5887));
NOR2X1 g62212(.A (n_867), .B (n_5971), .Y (n_5886));
NOR2X1 g62216(.A (n_859), .B (n_5968), .Y (n_5885));
CLKBUFX1 gbuf_d_172(.A(n_10388), .Y(d_out_172));
CLKBUFX1 gbuf_q_172(.A(q_in_172), .Y(g4575));
CLKBUFX1 gbuf_d_173(.A(n_5772), .Y(d_out_173));
CLKBUFX1 gbuf_q_173(.A(q_in_173), .Y(g4578));
CLKBUFX1 gbuf_d_174(.A(n_5777), .Y(d_out_174));
CLKBUFX1 gbuf_q_174(.A(q_in_174), .Y(g4388));
CLKBUFX1 gbuf_d_175(.A(n_5776), .Y(d_out_175));
CLKBUFX1 gbuf_q_175(.A(q_in_175), .Y(g4401));
CLKBUFX1 gbuf_d_176(.A(n_5790), .Y(d_out_176));
CLKBUFX1 gbuf_q_176(.A(q_in_176), .Y(g_11293));
CLKBUFX1 gbuf_d_177(.A(n_5780), .Y(d_out_177));
CLKBUFX1 gbuf_q_177(.A(q_in_177), .Y(g_21576));
CLKBUFX1 gbuf_d_178(.A(n_5768), .Y(d_out_178));
CLKBUFX1 gbuf_q_178(.A(q_in_178), .Y(g_19304));
NOR2X1 g62593(.A (n_5849), .B (n_1236), .Y (n_5884));
NOR2X1 g62597(.A (n_5839), .B (n_1063), .Y (n_5909));
NOR2X1 g62602(.A (n_5839), .B (n_1230), .Y (n_5883));
INVX1 g62607(.A (n_5881), .Y (n_5882));
NOR2X1 g62620(.A (n_5844), .B (n_1060), .Y (n_5907));
NOR2X1 g62623(.A (n_5844), .B (n_1160), .Y (n_5880));
NOR2X1 g62627(.A (n_5833), .B (n_1065), .Y (n_5905));
MX2X1 g61746(.A (g20901), .B (g_20208), .S0 (n_9359), .Y (n_5879));
NOR2X1 g62629(.A (n_5833), .B (n_1138), .Y (n_5878));
INVX1 g62634(.A (n_5876), .Y (n_5877));
NAND3X1 g62637(.A (n_5799), .B (n_2099), .C (n_9698), .Y (n_5875));
MX2X1 g61748(.A (g20901), .B (n_8799), .S0 (n_9019), .Y (n_5874));
INVX1 g62639(.A (n_5872), .Y (n_5873));
INVX1 g62642(.A (n_5870), .Y (n_5871));
AOI21X1 g60906(.A0 (n_3493), .A1 (g4521), .B0 (n_5767), .Y (n_5869));
MX2X1 g62694(.A (g2775), .B (n_5737), .S0 (n_9091), .Y (n_5868));
MX2X1 g62695(.A (g2783), .B (n_5736), .S0 (n_9797), .Y (n_5866));
MX2X1 g62696(.A (g2787), .B (n_5735), .S0 (n_9797), .Y (n_5865));
MX2X1 g62697(.A (g2795), .B (n_5734), .S0 (n_9834), .Y (n_5863));
MX2X1 g62699(.A (g2807), .B (n_5733), .S0 (n_9448), .Y (n_5862));
MX2X1 g62700(.A (g2815), .B (n_5731), .S0 (n_9797), .Y (n_5860));
MX2X1 g62701(.A (g2819), .B (n_5729), .S0 (n_9750), .Y (n_5859));
MX2X1 g62702(.A (g2827), .B (n_5727), .S0 (n_9000), .Y (n_5857));
INVX1 g62811(.A (n_5949), .Y (n_5854));
INVX1 g62841(.A (n_5947), .Y (n_5852));
INVX4 g62874(.A (n_5786), .Y (n_5844));
INVX2 g62883(.A (n_5784), .Y (n_5839));
OAI21X1 g60914(.A0 (g4512), .A1 (n_5711), .B0 (n_5756), .Y (n_5837));
INVX2 g62892(.A (n_5782), .Y (n_5833));
NOR2X1 g61937(.A (n_10416), .B (n_5506), .Y (n_5831));
AOI22X1 g62086(.A0 (n_2246), .A1 (n_5709), .B0 (g_16296), .B1(n_9599), .Y (n_5830));
CLKBUFX1 gbuf_d_179(.A(g8870), .Y(d_out_179));
CLKBUFX1 gbuf_q_179(.A(q_in_179), .Y(g8918));
NAND3X1 g61534(.A (n_5724), .B (n_6928), .C (n_9630), .Y (n_5828));
NAND2X1 g62209(.A (n_5508), .B (n_7395), .Y (n_5825));
NAND3X1 g62257(.A (n_7402), .B (n_10861), .C (g_16296), .Y (n_5824));
MX2X1 g62292(.A (g_16983), .B (n_5707), .S0 (n_9871), .Y (n_5822));
AND2X1 g61631(.A (n_5821), .B (n_3900), .Y (n_6254));
AOI21X1 g61643(.A0 (n_5755), .A1 (n_9351), .B0 (n_6005), .Y (n_6299));
CLKBUFX1 gbuf_d_180(.A(n_5738), .Y(d_out_180));
CLKBUFX1 gbuf_q_180(.A(q_in_180), .Y(g4382));
CLKBUFX1 gbuf_d_181(.A(n_5714), .Y(d_out_181));
CLKBUFX1 gbuf_q_181(.A(q_in_181), .Y(g7243));
CLKBUFX1 gbuf_d_182(.A(n_5716), .Y(d_out_182));
CLKBUFX1 gbuf_q_182(.A(q_in_182), .Y(g4392));
CLKBUFX1 gbuf_d_183(.A(n_5718), .Y(d_out_183));
CLKBUFX1 gbuf_q_183(.A(q_in_183), .Y(g12832));
CLKBUFX1 gbuf_d_184(.A(n_5720), .Y(d_out_184));
CLKBUFX1 gbuf_q_184(.A(q_in_184), .Y(g7257));
CLKBUFX1 gbuf_d_185(.A(n_5725), .Y(d_out_185));
CLKBUFX1 gbuf_q_185(.A(q_in_185), .Y(g_18308));
CLKBUFX1 gbuf_d_186(.A(n_5719), .Y(d_out_186));
CLKBUFX1 gbuf_q_186(.A(q_in_186), .Y(g4961));
OAI21X1 g64026(.A0 (g_19459), .A1 (n_11056), .B0 (n_7395), .Y(n_5820));
CLKBUFX1 gbuf_d_187(.A(n_5740), .Y(d_out_187));
CLKBUFX1 gbuf_q_187(.A(q_in_187), .Y(g_15691));
CLKBUFX1 gbuf_d_188(.A(n_5762), .Y(d_out_188));
CLKBUFX1 gbuf_q_188(.A(q_in_188), .Y(g2767));
CLKBUFX1 gbuf_d_189(.A(n_5760), .Y(d_out_189));
CLKBUFX1 gbuf_q_189(.A(q_in_189), .Y(g2779));
CLKBUFX1 gbuf_d_190(.A(n_5759), .Y(d_out_190));
CLKBUFX1 gbuf_q_190(.A(q_in_190), .Y(g2791));
CLKBUFX1 gbuf_d_191(.A(n_5758), .Y(d_out_191));
CLKBUFX1 gbuf_q_191(.A(q_in_191), .Y(g2795));
CLKBUFX1 gbuf_d_192(.A(n_5757), .Y(d_out_192));
CLKBUFX1 gbuf_q_192(.A(q_in_192), .Y(g2811));
CLKBUFX1 gbuf_d_193(.A(n_5746), .Y(d_out_193));
CLKBUFX1 gbuf_q_193(.A(q_in_193), .Y(g2823));
CLKBUFX1 gbuf_d_194(.A(n_5745), .Y(d_out_194));
CLKBUFX1 gbuf_q_194(.A(q_in_194), .Y(g2827));
NAND3X1 g61724(.A (n_5765), .B (g_16311), .C (n_10385), .Y (n_5819));
NAND2X1 g62563(.A (n_5788), .B (g1792), .Y (n_5818));
NAND2X1 g62566(.A (n_5786), .B (g2351), .Y (n_5817));
NAND2X1 g62567(.A (n_5784), .B (g1926), .Y (n_5816));
NAND2X1 g62568(.A (n_5782), .B (g2485), .Y (n_5815));
NAND2X1 g62586(.A (n_5944), .B (n_1522), .Y (n_5814));
MX2X1 g60905(.A (g4515), .B (n_2101), .S0 (g4521), .Y (n_5813));
INVX1 g62594(.A (n_5977), .Y (n_5811));
INVX1 g62603(.A (n_5974), .Y (n_5810));
NAND2X1 g62606(.A (n_5808), .B (g2060), .Y (n_5809));
NAND2X1 g62608(.A (n_5808), .B (n_1515), .Y (n_5881));
NAND2X1 g62610(.A (n_5808), .B (n_1524), .Y (n_5807));
NAND2X1 g62611(.A (n_5798), .B (g2217), .Y (n_5806));
NAND2X1 g62612(.A (n_5798), .B (n_1517), .Y (n_6067));
INVX1 g62624(.A (n_5971), .Y (n_5805));
INVX1 g62630(.A (n_5968), .Y (n_5804));
NAND2X1 g62633(.A (n_5944), .B (g2619), .Y (n_5803));
NAND2X1 g62632(.A (n_5799), .B (g1657), .Y (n_5801));
NAND2X1 g62635(.A (n_5944), .B (n_1506), .Y (n_5876));
NAND2X1 g62638(.A (n_5799), .B (n_1531), .Y (n_5800));
AND2X1 g62640(.A (n_5798), .B (n_1520), .Y (n_5872));
NAND2X1 g62641(.A (n_5798), .B (n_1527), .Y (n_5797));
AND2X1 g62643(.A (n_5799), .B (g25167), .Y (n_5870));
OAI21X1 g62663(.A0 (n_326), .A1 (n_9333), .B0 (n_5795), .Y (n_5796));
OAI21X1 g62664(.A0 (n_317), .A1 (n_9797), .B0 (n_5792), .Y (n_5794));
NAND2X1 g61823(.A (n_5624), .B (n_5700), .Y (n_5790));
CLKBUFX1 g62812(.A (n_5808), .Y (n_5949));
CLKBUFX1 g62842(.A (n_5798), .Y (n_5947));
INVX2 g62867(.A (n_5788), .Y (n_5849));
NOR2X1 g62036(.A (n_5695), .B (n_5284), .Y (n_5781));
MX2X1 g62137(.A (n_5663), .B (n_5639), .S0 (n_9218), .Y (n_5780));
AOI22X1 g61548(.A0 (n_2271), .A1 (n_7146), .B0 (g_18308), .B1(n_9193), .Y (n_5779));
MX2X1 g61026(.A (g4401), .B (n_5645), .S0 (n_9311), .Y (n_5777));
MX2X1 g61027(.A (g4405), .B (n_5644), .S0 (n_8955), .Y (n_5776));
AOI21X1 g62294(.A0 (g_10556), .A1 (n_9141), .B0 (n_5688), .Y(n_5775));
MX2X1 g62323(.A (g_22328), .B (g21176), .S0 (n_9599), .Y (n_5774));
CLKBUFX1 gbuf_d_195(.A(n_5693), .Y(d_out_195));
CLKBUFX1 gbuf_q_195(.A(q_in_195), .Y(g4749));
CLKBUFX1 gbuf_d_196(.A(n_5690), .Y(d_out_196));
CLKBUFX1 gbuf_q_196(.A(q_in_196), .Y(g4894));
CLKBUFX1 gbuf_d_197(.A(n_5692), .Y(d_out_197));
CLKBUFX1 gbuf_q_197(.A(q_in_197), .Y(g4771));
CLKBUFX1 gbuf_d_198(.A(n_5689), .Y(d_out_198));
CLKBUFX1 gbuf_q_198(.A(q_in_198), .Y(g4760));
CLKBUFX1 gbuf_d_199(.A(n_5694), .Y(d_out_199));
CLKBUFX1 gbuf_q_199(.A(q_in_199), .Y(g_21813));
AOI21X1 g61939(.A0 (n_5654), .A1 (n_816), .B0 (n_364), .Y (g33894));
OAI21X1 g61708(.A0 (n_5681), .A1 (n_9422), .B0 (n_10601), .Y(n_5772));
OR2X1 g62595(.A (n_5744), .B (n_561), .Y (n_5977));
AOI22X1 g61740(.A0 (n_2249), .A1 (n_8583), .B0 (g_11293), .B1(n_9772), .Y (n_5769));
OR2X1 g62604(.A (n_5742), .B (n_647), .Y (n_5974));
OR2X1 g62625(.A (n_5743), .B (n_592), .Y (n_5971));
OR2X1 g62631(.A (n_5741), .B (n_487), .Y (n_5968));
OAI22X1 g62676(.A0 (n_5668), .A1 (n_10952), .B0 (g_16983), .B1(n_9830), .Y (n_5768));
NOR2X1 g60908(.A (n_2100), .B (g4521), .Y (n_5767));
NOR2X1 g61810(.A (n_6153), .B (n_8583), .Y (n_5765));
OAI21X1 g62793(.A0 (n_5614), .A1 (n_5761), .B0 (n_5676), .Y (n_5762));
OAI21X1 g62794(.A0 (n_5613), .A1 (n_5761), .B0 (n_5674), .Y (n_5760));
OAI21X1 g62795(.A0 (n_5612), .A1 (n_5761), .B0 (n_5672), .Y (n_5759));
OAI21X1 g62796(.A0 (n_5611), .A1 (n_5761), .B0 (n_5671), .Y (n_5758));
OAI21X1 g62797(.A0 (n_5609), .A1 (n_5761), .B0 (n_5669), .Y (n_5757));
NAND2X1 g62800(.A (n_5667), .B (n_9091), .Y (n_5795));
NAND2X1 g62801(.A (n_5666), .B (n_9091), .Y (n_5792));
INVX1 g61836(.A (n_5755), .Y (n_5756));
INVX1 g62813(.A (n_10994), .Y (n_5808));
INVX4 g62830(.A (n_10787), .Y (n_5944));
INVX2 g62843(.A (n_5749), .Y (n_5798));
INVX4 g62855(.A (n_10614), .Y (n_5799));
OAI21X1 g62859(.A0 (n_5608), .A1 (n_5761), .B0 (n_5564), .Y (n_5746));
OAI21X1 g62860(.A0 (n_5607), .A1 (n_5761), .B0 (n_5563), .Y (n_5745));
INVX2 g62868(.A (n_5744), .Y (n_5788));
INVX2 g62877(.A (n_5743), .Y (n_5786));
INVX2 g62886(.A (n_5742), .Y (n_5784));
INVX2 g62895(.A (n_5741), .Y (n_5782));
CLKBUFX1 gbuf_d_200(.A(n_5642), .Y(d_out_200));
CLKBUFX1 gbuf_q_200(.A(q_in_200), .Y(g_19515));
CLKBUFX1 gbuf_d_201(.A(n_5664), .Y(d_out_201));
CLKBUFX1 gbuf_q_201(.A(q_in_201), .Y(g20901));
OAI21X1 g61945(.A0 (g_22605), .A1 (n_10013), .B0 (n_5678), .Y(n_5740));
NAND3X1 g61008(.A (n_5631), .B (n_2269), .C (n_5592), .Y (n_5738));
OAI21X1 g63287(.A0 (g2767), .A1 (n_5732), .B0 (n_5662), .Y (n_5737));
OAI21X1 g63288(.A0 (n_5730), .A1 (g2779), .B0 (n_5661), .Y (n_5736));
OAI21X1 g63289(.A0 (n_5728), .A1 (g2791), .B0 (n_5660), .Y (n_5735));
OAI21X1 g63290(.A0 (n_5726), .A1 (g2795), .B0 (n_5659), .Y (n_5734));
OAI21X1 g63291(.A0 (n_5732), .A1 (g2799), .B0 (n_5658), .Y (n_5733));
OAI21X1 g63292(.A0 (n_5730), .A1 (g2811), .B0 (n_5657), .Y (n_5731));
OAI21X1 g63293(.A0 (n_5728), .A1 (g2823), .B0 (n_5655), .Y (n_5729));
OAI21X1 g63294(.A0 (n_5726), .A1 (g2827), .B0 (n_5656), .Y (n_5727));
NAND2X1 g61571(.A (n_5602), .B (n_5652), .Y (n_5725));
NOR2X1 g61572(.A (n_5723), .B (n_7146), .Y (n_5724));
NAND3X1 g61030(.A (n_5641), .B (n_5273), .C (n_5578), .Y (n_5720));
NAND2X1 g61583(.A (n_3752), .B (n_5650), .Y (n_5719));
OAI21X1 g61031(.A0 (g4455), .A1 (n_9627), .B0 (n_5715), .Y (n_5718));
OAI21X1 g61050(.A0 (n_74), .A1 (n_9681), .B0 (n_5715), .Y (n_5716));
CLKBUFX1 gbuf_d_202(.A(n_6858), .Y(d_out_202));
CLKBUFX1 gbuf_qn_202(.A(qn_in_202), .Y(g1682));
CLKBUFX1 gbuf_d_203(.A(n_5677), .Y(d_out_203));
CLKBUFX1 gbuf_q_203(.A(q_in_203), .Y(g4430));
CLKBUFX1 gbuf_d_204(.A(n_8706), .Y(d_out_204));
CLKBUFX1 gbuf_q_204(.A(q_in_204), .Y(n_3618));
CLKBUFX1 gbuf_d_205(.A(n_5646), .Y(d_out_205));
CLKBUFX1 gbuf_q_205(.A(q_in_205), .Y(n_3589));
CLKBUFX1 gbuf_d_206(.A(n_5686), .Y(d_out_206));
CLKBUFX1 gbuf_q_206(.A(q_in_206), .Y(n_3611));
CLKBUFX1 gbuf_d_207(.A(n_5683), .Y(d_out_207));
CLKBUFX1 gbuf_qn_207(.A(qn_in_207), .Y(g4434));
CLKBUFX1 gbuf_d_208(.A(n_5680), .Y(d_out_208));
CLKBUFX1 gbuf_q_208(.A(q_in_208), .Y(g5084));
NAND2X1 g61051(.A (n_5643), .B (n_5637), .Y (n_5714));
AND2X1 g64156(.A (n_10310), .B (n_9874), .Y (n_7402));
CLKBUFX1 gbuf_d_209(.A(g8917), .Y(d_out_209));
CLKBUFX1 gbuf_q_209(.A(q_in_209), .Y(g8870));
OR2X1 g64274(.A (n_172), .B (n_10311), .Y (n_5712));
NAND3X1 g61733(.A (n_5711), .B (g4572), .C (n_10687), .Y (n_5821));
CLKBUFX1 gbuf_d_210(.A(n_5629), .Y(d_out_210));
CLKBUFX1 gbuf_qn_210(.A(qn_in_210), .Y(g4521));
INVX1 g62761(.A (g_22328), .Y (n_5707));
AND2X1 g61837(.A (n_5711), .B (g20049), .Y (n_5755));
NAND2X1 g62845(.A (n_5622), .B (n_5705), .Y (n_5749));
AOI21X1 g62869(.A0 (n_5569), .A1 (n_5704), .B0 (n_5703), .Y (n_5744));
AOI21X1 g62878(.A0 (n_5567), .A1 (n_5704), .B0 (n_5703), .Y (n_5743));
AOI21X1 g62887(.A0 (n_5568), .A1 (n_5702), .B0 (n_5701), .Y (n_5742));
AOI21X1 g62896(.A0 (n_5566), .A1 (n_5702), .B0 (n_5701), .Y (n_5741));
NAND3X1 g61935(.A (n_5619), .B (g_11293), .C (n_9797), .Y (n_5700));
CLKBUFX1 gbuf_d_211(.A(n_10690), .Y(d_out_211));
CLKBUFX1 gbuf_q_211(.A(q_in_211), .Y(g21245));
NAND4X1 g62286(.A (n_2448), .B (n_2137), .C (n_5543), .D (n_1686), .Y(n_5695));
MX2X1 g62325(.A (g_20208), .B (n_5583), .S0 (n_9359), .Y (n_5694));
NAND2X1 g61634(.A (n_3582), .B (n_5599), .Y (n_5693));
NAND2X1 g61635(.A (n_3580), .B (n_5596), .Y (n_5692));
CLKBUFX1 gbuf_d_212(.A(n_10955), .Y(d_out_212));
CLKBUFX1 gbuf_q_212(.A(q_in_212), .Y(n_3616));
CLKBUFX1 gbuf_d_213(.A(n_5600), .Y(d_out_213));
CLKBUFX1 gbuf_q_213(.A(q_in_213), .Y(n_3604));
CLKBUFX1 gbuf_d_214(.A(n_5593), .Y(d_out_214));
CLKBUFX1 gbuf_qn_214(.A(qn_in_214), .Y(g4826));
CLKBUFX1 gbuf_d_215(.A(n_5627), .Y(d_out_215));
CLKBUFX1 gbuf_qn_215(.A(qn_in_215), .Y(g4831));
CLKBUFX1 gbuf_d_216(.A(n_5625), .Y(d_out_216));
CLKBUFX1 gbuf_q_216(.A(q_in_216), .Y(g7245));
CLKBUFX1 gbuf_d_217(.A(n_5626), .Y(d_out_217));
CLKBUFX1 gbuf_q_217(.A(q_in_217), .Y(g7260));
CLKBUFX1 gbuf_d_218(.A(n_5615), .Y(d_out_218));
CLKBUFX1 gbuf_q_218(.A(q_in_218), .Y(g5080));
CLKBUFX1 gbuf_d_219(.A(n_5590), .Y(d_out_219));
CLKBUFX1 gbuf_q_219(.A(q_in_219), .Y(g_20208));
INVX1 g62589(.A (n_6523), .Y (n_5709));
NAND2X1 g61735(.A (n_5633), .B (n_3578), .Y (n_5690));
NAND2X1 g61734(.A (n_5634), .B (n_3581), .Y (n_5689));
NOR3X1 g62613(.A (n_10861), .B (g_16296), .C (n_9353), .Y (n_5688));
NAND3X1 g61801(.A (n_5576), .B (n_2560), .C (n_3613), .Y (n_5686));
CLKBUFX1 gbuf_d_220(.A(n_5570), .Y(d_out_220));
CLKBUFX1 gbuf_q_220(.A(q_in_220), .Y(g_22328));
CLKBUFX1 gbuf_d_221(.A(g8916), .Y(d_out_221));
CLKBUFX1 gbuf_q_221(.A(q_in_221), .Y(g8917));
MX2X1 g61842(.A (g4452), .B (n_5532), .S0 (n_8955), .Y (n_5683));
INVX1 g61885(.A (g4572), .Y (n_5681));
OAI21X1 g61915(.A0 (n_5515), .A1 (g5080), .B0 (n_5571), .Y (n_5680));
CLKBUFX1 gbuf_d_222(.A(n_5557), .Y(d_out_222));
CLKBUFX1 gbuf_q_222(.A(q_in_222), .Y(g_12922));
NAND4X1 g62061(.A (n_5547), .B (n_9834), .C (n_4126), .D (n_10264),.Y (n_5678));
OAI22X1 g61482(.A0 (n_5521), .A1 (n_9976), .B0 (g4434), .B1 (n_9627),.Y (n_5677));
AOI22X1 g63305(.A0 (g2763), .A1 (n_10078), .B0 (g2767), .B1 (n_5675),.Y (n_5676));
AOI22X1 g63306(.A0 (g2767), .A1 (n_9871), .B0 (g2779), .B1 (n_5675),.Y (n_5674));
AOI22X1 g63307(.A0 (g2779), .A1 (n_10078), .B0 (g2791), .B1 (n_5675),.Y (n_5672));
AOI22X1 g63308(.A0 (g2795), .A1 (n_5675), .B0 (g2791), .B1 (n_10376),.Y (n_5671));
AOI22X1 g63309(.A0 (g2799), .A1 (n_10078), .B0 (g2811), .B1 (n_5675),.Y (n_5669));
AOI21X1 g63330(.A0 (n_5440), .A1 (g_19304), .B0 (n_5565), .Y(n_5668));
AOI22X1 g63336(.A0 (n_5226), .A1 (n_5513), .B0 (n_5224), .B1(n_5665), .Y (n_5667));
AOI22X1 g63343(.A0 (n_5346), .A1 (n_5665), .B0 (n_5225), .B1(n_5513), .Y (n_5666));
MX2X1 g62108(.A (g_19136), .B (n_5663), .S0 (n_10005), .Y (n_5664));
NAND2X1 g63432(.A (n_5732), .B (g2771), .Y (n_5662));
NAND2X1 g63433(.A (n_5730), .B (g2775), .Y (n_5661));
NAND2X1 g63434(.A (n_5728), .B (g2783), .Y (n_5660));
NAND2X1 g63435(.A (n_5726), .B (g2787), .Y (n_5659));
NAND2X1 g63436(.A (n_5732), .B (g2803), .Y (n_5658));
NAND2X1 g63437(.A (n_5730), .B (g2807), .Y (n_5657));
NAND2X1 g63438(.A (n_5726), .B (g2819), .Y (n_5656));
NAND2X1 g63439(.A (n_5728), .B (g2815), .Y (n_5655));
NOR2X1 g62228(.A (g_8896), .B (n_5560), .Y (n_5654));
NAND3X1 g61626(.A (n_5556), .B (g_18308), .C (n_10063), .Y (n_5652));
NAND4X1 g61640(.A (n_5553), .B (n_2064), .C (n_9279), .D (n_10296),.Y (n_5650));
CLKBUFX1 gbuf_d_223(.A(n_5575), .Y(d_out_223));
CLKBUFX1 gbuf_q_223(.A(q_in_223), .Y(g1950));
CLKBUFX1 gbuf_d_224(.A(n_10363), .Y(d_out_224));
CLKBUFX1 gbuf_qn_224(.A(qn_in_224), .Y(g4821));
CLKBUFX1 gbuf_d_225(.A(n_5549), .Y(d_out_225));
CLKBUFX1 gbuf_qn_225(.A(qn_in_225), .Y(g5011));
CLKBUFX1 gbuf_d_226(.A(n_5587), .Y(d_out_226));
CLKBUFX1 gbuf_q_226(.A(q_in_226), .Y(g4704));
CLKBUFX1 gbuf_d_227(.A(n_5574), .Y(d_out_227));
CLKBUFX1 gbuf_q_227(.A(q_in_227), .Y(g_13255));
NAND3X1 g61717(.A (n_5584), .B (n_2540), .C (n_3590), .Y (n_5646));
OR2X1 g61065(.A (n_5581), .B (g4411), .Y (n_5645));
OR2X1 g61066(.A (n_5580), .B (g4405), .Y (n_5644));
AOI21X1 g61073(.A0 (n_5591), .A1 (n_5453), .B0 (n_5630), .Y (n_5715));
NAND3X1 g61075(.A (n_5640), .B (n_5363), .C (n_10005), .Y (n_5643));
MX2X1 g62678(.A (g_9584), .B (n_3559), .S0 (n_9256), .Y (n_5642));
NAND3X1 g61076(.A (n_5640), .B (g4382), .C (n_9359), .Y (n_5641));
MX2X1 g62681(.A (g_21576), .B (g_9584), .S0 (n_5582), .Y (n_5639));
AOI21X1 g61079(.A0 (g4411), .A1 (n_9856), .B0 (n_5579), .Y (n_5637));
NAND3X1 g61817(.A (n_5540), .B (n_2581), .C (n_2067), .Y (n_5634));
NAND3X1 g61819(.A (n_5539), .B (n_4091), .C (n_1626), .Y (n_5633));
INVX1 g61114(.A (n_5630), .Y (n_5631));
OAI21X1 g60915(.A0 (g4512), .A1 (n_9422), .B0 (n_5530), .Y (n_5629));
MX2X1 g61876(.A (g5965), .B (n_5460), .S0 (n_9218), .Y (n_5627));
CLKBUFX1 gbuf_d_228(.A(n_5536), .Y(d_out_228));
CLKBUFX1 gbuf_q_228(.A(q_in_228), .Y(g4572));
CLKBUFX1 gbuf_d_229(.A(n_5534), .Y(d_out_229));
CLKBUFX1 gbuf_q_229(.A(q_in_229), .Y(g20049));
NAND3X1 g61914(.A (n_5517), .B (n_5221), .C (n_5455), .Y (n_5626));
OAI21X1 g61947(.A0 (n_5365), .A1 (n_5454), .B0 (n_5522), .Y (n_5625));
AOI22X1 g61956(.A0 (n_2260), .A1 (n_6655), .B0 (g_15691), .B1(n_9129), .Y (n_5624));
OAI21X1 g63221(.A0 (n_6892), .A1 (g2803), .B0 (n_8557), .Y (n_5622));
NOR2X1 g62047(.A (n_6153), .B (n_6655), .Y (n_5619));
OAI21X1 g63239(.A0 (n_6893), .A1 (g2771), .B0 (n_8557), .Y (n_5617));
OAI21X1 g62105(.A0 (g5077), .A1 (n_9422), .B0 (n_5519), .Y (n_5615));
NAND2X1 g63462(.A (g1632), .B (n_5675), .Y (n_5614));
NAND2X1 g63464(.A (g1768), .B (n_5675), .Y (n_5613));
NAND2X1 g63466(.A (g1902), .B (n_5675), .Y (n_5612));
NAND2X1 g63467(.A (g2036), .B (n_5675), .Y (n_5611));
NAND2X1 g63468(.A (g2193), .B (n_5675), .Y (n_5610));
NAND2X1 g63469(.A (g2327), .B (n_5675), .Y (n_5609));
NAND2X1 g63471(.A (g2461), .B (n_5675), .Y (n_5608));
NAND2X1 g63472(.A (n_5675), .B (g2595), .Y (n_5607));
AOI22X1 g61646(.A0 (n_2296), .A1 (n_11104), .B0 (g_12922), .B1(n_9903), .Y (n_5602));
CLKBUFX1 gbuf_d_230(.A(n_5538), .Y(d_out_230));
CLKBUFX1 gbuf_q_230(.A(q_in_230), .Y(g1816));
CLKBUFX1 gbuf_d_231(.A(n_5529), .Y(d_out_231));
CLKBUFX1 gbuf_qn_231(.A(qn_in_231), .Y(g2161));
CLKBUFX1 gbuf_d_232(.A(n_5527), .Y(d_out_232));
CLKBUFX1 gbuf_qn_232(.A(qn_in_232), .Y(g2169));
CLKBUFX1 gbuf_d_233(.A(n_5526), .Y(d_out_233));
CLKBUFX1 gbuf_qn_233(.A(qn_in_233), .Y(g2173));
CLKBUFX1 gbuf_d_234(.A(n_5524), .Y(d_out_234));
CLKBUFX1 gbuf_qn_234(.A(qn_in_234), .Y(g2181));
CLKBUFX1 gbuf_d_235(.A(n_5531), .Y(d_out_235));
CLKBUFX1 gbuf_q_235(.A(q_in_235), .Y(g2084));
CLKBUFX1 gbuf_d_236(.A(n_6664), .Y(d_out_236));
CLKBUFX1 gbuf_q_236(.A(q_in_236), .Y(g2555));
CLKBUFX1 gbuf_d_237(.A(n_10377), .Y(d_out_237));
CLKBUFX1 gbuf_q_237(.A(q_in_237), .Y(g2153));
CLKBUFX1 gbuf_d_238(.A(n_5537), .Y(d_out_238));
CLKBUFX1 gbuf_q_238(.A(q_in_238), .Y(g_22371));
NAND3X1 g61718(.A (n_5544), .B (n_2298), .C (n_3606), .Y (n_5600));
NAND4X1 g61741(.A (n_5542), .B (n_8906), .C (n_9279), .D (n_2067), .Y(n_5599));
NAND4X1 g61742(.A (n_5541), .B (n_2067), .C (n_9139), .D (n_8694), .Y(n_5596));
MX2X1 g61752(.A (g6311), .B (n_5481), .S0 (n_8955), .Y (n_5593));
NAND3X1 g61074(.A (n_5409), .B (n_5591), .C (n_9453), .Y (n_5592));
MX2X1 g62691(.A (g_22371), .B (n_5465), .S0 (n_9558), .Y (n_5590));
NAND2X1 g61816(.A (n_3588), .B (n_5483), .Y (n_5587));
NAND3X1 g61830(.A (n_7093), .B (n_3394), .C (n_9425), .Y (n_5584));
CLKBUFX1 gbuf_d_239(.A(n_5489), .Y(d_out_239));
CLKBUFX1 gbuf_qn_239(.A(qn_in_239), .Y(g1612));
NOR2X1 g61115(.A (n_1657), .B (n_5591), .Y (n_5630));
MX2X1 g62937(.A (n_5663), .B (g14167), .S0 (n_5582), .Y (n_5583));
NOR2X1 g61124(.A (n_784), .B (n_5591), .Y (n_5581));
NOR2X1 g61125(.A (n_597), .B (n_5591), .Y (n_5580));
AND2X1 g61126(.A (n_5591), .B (g4375), .Y (n_5640));
NOR2X1 g61127(.A (n_5591), .B (n_5378), .Y (n_5579));
OR2X1 g61128(.A (n_5591), .B (n_1980), .Y (n_5578));
NAND3X1 g61940(.A (n_5458), .B (n_5459), .C (n_10385), .Y (n_5576));
NAND3X1 g61152(.A (n_5450), .B (n_2266), .C (n_4131), .Y (n_5575));
CLKBUFX1 gbuf_d_240(.A(g8915), .Y(d_out_240));
CLKBUFX1 gbuf_q_240(.A(q_in_240), .Y(g8916));
NAND3X1 g63208(.A (n_5573), .B (n_2531), .C (n_5370), .Y (n_5574));
AOI22X1 g62080(.A0 (n_5518), .A1 (g5073), .B0 (n_5514), .B1 (g5080),.Y (n_5571));
MX2X1 g63368(.A (g_13255), .B (n_6280), .S0 (n_9681), .Y (n_5570));
NOR2X1 g63476(.A (n_6895), .B (g2775), .Y (n_5569));
NOR2X1 g63486(.A (n_6895), .B (g2783), .Y (n_5568));
NOR2X1 g63504(.A (n_6892), .B (g2807), .Y (n_5567));
NOR2X1 g63508(.A (n_6895), .B (g2815), .Y (n_5566));
NOR2X1 g63518(.A (n_5440), .B (n_3519), .Y (n_5565));
AOI22X1 g63543(.A0 (n_2231), .A1 (n_5562), .B0 (g2811), .B1(n_10376), .Y (n_5564));
AOI22X1 g63544(.A0 (n_1968), .A1 (n_5562), .B0 (g2823), .B1 (n_9129),.Y (n_5563));
INVX1 g62335(.A (g_19136), .Y (n_5560));
NAND2X1 g63878(.A (n_5559), .B (n_8557), .Y (n_5732));
NAND2X1 g63879(.A (n_3866), .B (n_5559), .Y (n_5730));
NAND3X1 g63910(.A (n_5559), .B (n_10650), .C (n_3868), .Y (n_5728));
NAND3X1 g63911(.A (n_5559), .B (n_10650), .C (g2724), .Y (n_5726));
CLKBUFX1 gbuf_d_241(.A(n_5485), .Y(d_out_241));
CLKBUFX1 gbuf_q_241(.A(q_in_241), .Y(g1526));
CLKBUFX1 gbuf_d_242(.A(n_5449), .Y(d_out_242));
CLKBUFX1 gbuf_qn_242(.A(qn_in_242), .Y(g1454));
CLKBUFX1 gbuf_d_243(.A(n_5448), .Y(d_out_243));
CLKBUFX1 gbuf_qn_243(.A(qn_in_243), .Y(g1467));
CLKBUFX1 gbuf_d_244(.A(n_5447), .Y(d_out_244));
CLKBUFX1 gbuf_qn_244(.A(qn_in_244), .Y(g1484));
CLKBUFX1 gbuf_d_245(.A(n_5451), .Y(d_out_245));
CLKBUFX1 gbuf_qn_245(.A(qn_in_245), .Y(g1437));
CLKBUFX1 gbuf_d_246(.A(n_5462), .Y(d_out_246));
CLKBUFX1 gbuf_qn_246(.A(qn_in_246), .Y(g_20839));
CLKBUFX1 gbuf_d_247(.A(n_5461), .Y(d_out_247));
CLKBUFX1 gbuf_qn_247(.A(qn_in_247), .Y(g_18200));
CLKBUFX1 gbuf_d_248(.A(n_5464), .Y(d_out_248));
CLKBUFX1 gbuf_qn_248(.A(qn_in_248), .Y(g_18220));
CLKBUFX1 gbuf_d_249(.A(n_5466), .Y(d_out_249));
CLKBUFX1 gbuf_qn_249(.A(qn_in_249), .Y(g_22236));
CLKBUFX1 gbuf_d_250(.A(n_5445), .Y(d_out_250));
CLKBUFX1 gbuf_qn_250(.A(qn_in_250), .Y(g2241));
CLKBUFX1 gbuf_d_251(.A(n_5444), .Y(d_out_251));
CLKBUFX1 gbuf_qn_251(.A(qn_in_251), .Y(g2375));
CLKBUFX1 gbuf_d_252(.A(n_5442), .Y(d_out_252));
CLKBUFX1 gbuf_qn_252(.A(qn_in_252), .Y(g2643));
CLKBUFX1 gbuf_d_253(.A(n_5467), .Y(d_out_253));
CLKBUFX1 gbuf_qn_253(.A(qn_in_253), .Y(g2177));
CLKBUFX1 gbuf_d_254(.A(n_5502), .Y(d_out_254));
CLKBUFX1 gbuf_qn_254(.A(qn_in_254), .Y(g2004));
CLKBUFX1 gbuf_d_255(.A(n_5499), .Y(d_out_255));
CLKBUFX1 gbuf_qn_255(.A(qn_in_255), .Y(g2020));
CLKBUFX1 gbuf_d_256(.A(n_5495), .Y(d_out_256));
CLKBUFX1 gbuf_qn_256(.A(qn_in_256), .Y(g2024));
CLKBUFX1 gbuf_d_257(.A(n_5492), .Y(d_out_257));
CLKBUFX1 gbuf_qn_257(.A(qn_in_257), .Y(g1600));
CLKBUFX1 gbuf_d_258(.A(n_5490), .Y(d_out_258));
CLKBUFX1 gbuf_qn_258(.A(qn_in_258), .Y(g1608));
CLKBUFX1 gbuf_d_259(.A(n_5487), .Y(d_out_259));
CLKBUFX1 gbuf_qn_259(.A(qn_in_259), .Y(g1620));
CLKBUFX1 gbuf_d_260(.A(n_5497), .Y(d_out_260));
CLKBUFX1 gbuf_qn_260(.A(qn_in_260), .Y(g2016));
CLKBUFX1 gbuf_d_261(.A(n_5468), .Y(d_out_261));
CLKBUFX1 gbuf_q_261(.A(q_in_261), .Y(g4616));
CLKBUFX1 gbuf_d_262(.A(n_5456), .Y(d_out_262));
CLKBUFX1 gbuf_q_262(.A(q_in_262), .Y(g4608));
CLKBUFX1 gbuf_d_263(.A(n_5437), .Y(d_out_263));
CLKBUFX1 gbuf_qn_263(.A(qn_in_263), .Y(g_4449));
CLKBUFX1 gbuf_d_264(.A(n_5504), .Y(d_out_264));
CLKBUFX1 gbuf_q_264(.A(q_in_264), .Y(g_16571));
CLKBUFX1 gbuf_d_265(.A(n_10590), .Y(d_out_265));
CLKBUFX1 gbuf_q_265(.A(q_in_265), .Y(n_11065));
CLKBUFX1 gbuf_d_266(.A(n_6757), .Y(d_out_266));
CLKBUFX1 gbuf_q_266(.A(q_in_266), .Y(g1996));
CLKBUFX1 gbuf_d_267(.A(n_5486), .Y(d_out_267));
CLKBUFX1 gbuf_q_267(.A(q_in_267), .Y(g4040));
CLKBUFX1 gbuf_d_268(.A(n_5476), .Y(d_out_268));
CLKBUFX1 gbuf_q_268(.A(q_in_268), .Y(g3831));
CLKBUFX1 gbuf_d_269(.A(n_5474), .Y(d_out_269));
CLKBUFX1 gbuf_qn_269(.A(qn_in_269), .Y(g3835));
NAND2X1 g61714(.A (n_5431), .B (n_5505), .Y (n_5557));
NOR2X1 g61715(.A (n_5723), .B (n_11104), .Y (n_5556));
AOI21X1 g61736(.A0 (n_5422), .A1 (n_2024), .B0 (n_6243), .Y (n_5553));
MX2X1 g61753(.A (g6657), .B (n_5420), .S0 (n_9234), .Y (n_5549));
INVX1 g62682(.A (n_6153), .Y (n_5547));
NAND3X1 g61831(.A (n_7333), .B (n_3547), .C (n_9558), .Y (n_5544));
CLKBUFX1 gbuf_d_270(.A(n_6631), .Y(d_out_270));
CLKBUFX1 gbuf_q_270(.A(q_in_270), .Y(g2421));
NAND4X1 g62915(.A (g3897), .B (n_4988), .C (n_5402), .D (g4031), .Y(n_5543));
NOR2X1 g61928(.A (n_5408), .B (n_10947), .Y (n_5542));
NOR2X1 g61931(.A (n_5406), .B (n_3784), .Y (n_5541));
NOR2X1 g61930(.A (n_5407), .B (n_3612), .Y (n_5540));
NOR2X1 g61933(.A (n_5405), .B (n_3605), .Y (n_5539));
NAND3X1 g61151(.A (n_5377), .B (n_2242), .C (n_4133), .Y (n_5538));
MX2X1 g63138(.A (g_22600), .B (n_5271), .S0 (n_9091), .Y (n_5537));
INVX1 g62015(.A (n_10601), .Y (n_5536));
INVX1 g62017(.A (n_10386), .Y (n_5534));
OR2X1 g62020(.A (n_5375), .B (g4452), .Y (n_5532));
CLKBUFX1 gbuf_d_271(.A(g14167), .Y(d_out_271));
CLKBUFX1 gbuf_q_271(.A(q_in_271), .Y(g_9584));
NAND3X1 g61161(.A (n_5373), .B (n_2272), .C (n_4614), .Y (n_5531));
CLKBUFX1 gbuf_d_272(.A(n_5369), .Y(d_out_272));
CLKBUFX1 gbuf_qn_272(.A(qn_in_272), .Y(g2509));
OAI21X1 g62066(.A0 (g4531), .A1 (g4581), .B0 (n_10005), .Y (n_5530));
OAI22X1 g61170(.A0 (n_5268), .A1 (n_9884), .B0 (g2165), .B1 (n_9992),.Y (n_5529));
OAI22X1 g61172(.A0 (n_5267), .A1 (n_10952), .B0 (g2161), .B1(n_9627), .Y (n_5527));
OAI22X1 g61173(.A0 (n_5266), .A1 (n_9772), .B0 (g2177), .B1 (n_9651),.Y (n_5526));
OAI22X1 g61175(.A0 (n_5265), .A1 (n_9928), .B0 (g2169), .B1(n_10063), .Y (n_5524));
AOI21X1 g62111(.A0 (g4443), .A1 (n_9772), .B0 (n_5379), .Y (n_5522));
AOI21X1 g61529(.A0 (n_1015), .A1 (n_5454), .B0 (g4443), .Y (n_5521));
NAND3X1 g63532(.A (n_6280), .B (g_19304), .C (g_13901), .Y (n_5520));
NAND2X1 g62222(.A (n_5518), .B (n_5215), .Y (n_5519));
NAND3X1 g62242(.A (n_5374), .B (n_5364), .C (g4382), .Y (n_5517));
OR2X1 g62269(.A (n_5361), .B (n_5514), .Y (n_5515));
CLKBUFX1 gbuf_d_273(.A(n_5430), .Y(d_out_273));
CLKBUFX1 gbuf_q_273(.A(q_in_273), .Y(g_19136));
AND2X1 g63877(.A (n_5562), .B (n_9358), .Y (n_5675));
OAI21X1 g63884(.A0 (n_10841), .A1 (n_5362), .B0 (n_5436), .Y(n_5761));
INVX1 g63959(.A (n_5665), .Y (n_5513));
CLKBUFX1 gbuf_d_274(.A(n_5424), .Y(d_out_274));
CLKBUFX1 gbuf_q_274(.A(q_in_274), .Y(g1379));
CLKBUFX1 gbuf_d_275(.A(n_5404), .Y(d_out_275));
CLKBUFX1 gbuf_qn_275(.A(qn_in_275), .Y(g2165));
CLKBUFX1 gbuf_d_276(.A(n_5400), .Y(d_out_276));
CLKBUFX1 gbuf_qn_276(.A(qn_in_276), .Y(g2295));
CLKBUFX1 gbuf_d_277(.A(n_5398), .Y(d_out_277));
CLKBUFX1 gbuf_qn_277(.A(qn_in_277), .Y(g2303));
CLKBUFX1 gbuf_d_278(.A(n_5396), .Y(d_out_278));
CLKBUFX1 gbuf_qn_278(.A(qn_in_278), .Y(g2307));
CLKBUFX1 gbuf_d_279(.A(n_5395), .Y(d_out_279));
CLKBUFX1 gbuf_qn_279(.A(qn_in_279), .Y(g2311));
CLKBUFX1 gbuf_d_280(.A(n_5394), .Y(d_out_280));
CLKBUFX1 gbuf_qn_280(.A(qn_in_280), .Y(g2315));
CLKBUFX1 gbuf_d_281(.A(n_5392), .Y(d_out_281));
CLKBUFX1 gbuf_qn_281(.A(qn_in_281), .Y(g2429));
CLKBUFX1 gbuf_d_282(.A(n_5388), .Y(d_out_282));
CLKBUFX1 gbuf_qn_282(.A(qn_in_282), .Y(g2441));
CLKBUFX1 gbuf_d_283(.A(n_5387), .Y(d_out_283));
CLKBUFX1 gbuf_qn_283(.A(qn_in_283), .Y(g2445));
CLKBUFX1 gbuf_d_284(.A(n_5386), .Y(d_out_284));
CLKBUFX1 gbuf_qn_284(.A(qn_in_284), .Y(g2449));
CLKBUFX1 gbuf_d_285(.A(n_5385), .Y(d_out_285));
CLKBUFX1 gbuf_qn_285(.A(qn_in_285), .Y(g2563));
CLKBUFX1 gbuf_d_286(.A(n_5384), .Y(d_out_286));
CLKBUFX1 gbuf_qn_286(.A(qn_in_286), .Y(g2571));
CLKBUFX1 gbuf_d_287(.A(n_5382), .Y(d_out_287));
CLKBUFX1 gbuf_qn_287(.A(qn_in_287), .Y(g2579));
CLKBUFX1 gbuf_d_288(.A(n_5380), .Y(d_out_288));
CLKBUFX1 gbuf_qn_288(.A(qn_in_288), .Y(g2583));
CLKBUFX1 gbuf_d_289(.A(n_5391), .Y(d_out_289));
CLKBUFX1 gbuf_qn_289(.A(qn_in_289), .Y(g2437));
CLKBUFX1 gbuf_d_290(.A(n_5383), .Y(d_out_290));
CLKBUFX1 gbuf_qn_290(.A(qn_in_290), .Y(g2575));
CLKBUFX1 gbuf_d_291(.A(n_5428), .Y(d_out_291));
CLKBUFX1 gbuf_qn_291(.A(qn_in_291), .Y(g1616));
CLKBUFX1 gbuf_d_292(.A(n_5393), .Y(d_out_292));
CLKBUFX1 gbuf_q_292(.A(q_in_292), .Y(g_15380));
CLKBUFX1 gbuf_d_293(.A(n_5423), .Y(d_out_293));
CLKBUFX1 gbuf_q_293(.A(q_in_293), .Y(g_19659));
CLKBUFX1 gbuf_d_294(.A(n_5411), .Y(d_out_294));
CLKBUFX1 gbuf_q_294(.A(q_in_294), .Y(g_12465));
CLKBUFX1 gbuf_d_295(.A(n_5372), .Y(d_out_295));
CLKBUFX1 gbuf_q_295(.A(q_in_295), .Y(g_21447));
CLKBUFX1 gbuf_d_296(.A(n_6639), .Y(d_out_296));
CLKBUFX1 gbuf_q_296(.A(q_in_296), .Y(g2287));
CLKBUFX1 gbuf_d_297(.A(n_5359), .Y(d_out_297));
CLKBUFX1 gbuf_qn_297(.A(qn_in_297), .Y(g2089));
CLKBUFX1 gbuf_d_298(.A(n_5358), .Y(d_out_298));
CLKBUFX1 gbuf_qn_298(.A(qn_in_298), .Y(g2246));
CLKBUFX1 gbuf_d_299(.A(n_5357), .Y(d_out_299));
CLKBUFX1 gbuf_q_299(.A(q_in_299), .Y(g2269));
CLKBUFX1 gbuf_d_300(.A(n_5356), .Y(d_out_300));
CLKBUFX1 gbuf_qn_300(.A(qn_in_300), .Y(g2273));
CLKBUFX1 gbuf_d_301(.A(n_5432), .Y(d_out_301));
CLKBUFX1 gbuf_q_301(.A(q_in_301), .Y(g5156));
CLKBUFX1 gbuf_d_302(.A(n_5415), .Y(d_out_302));
CLKBUFX1 gbuf_qn_302(.A(qn_in_302), .Y(g3827));
CLKBUFX1 gbuf_d_303(.A(n_5414), .Y(d_out_303));
CLKBUFX1 gbuf_q_303(.A(q_in_303), .Y(g2197));
CLKBUFX1 gbuf_d_304(.A(n_5412), .Y(d_out_304));
CLKBUFX1 gbuf_q_304(.A(q_in_304), .Y(g2227));
CLKBUFX1 gbuf_d_305(.A(n_5410), .Y(d_out_305));
CLKBUFX1 gbuf_q_305(.A(q_in_305), .Y(g3817));
CLKBUFX1 gbuf_d_306(.A(n_5397), .Y(d_out_306));
CLKBUFX1 gbuf_q_306(.A(q_in_306), .Y(g_22600));
XOR2X1 g62665(.A (g_10556), .B (n_5287), .Y (n_5508));
NAND4X1 g62671(.A (n_5403), .B (n_4607), .C (n_4088), .D (n_4984), .Y(n_5506));
CLKBUFX2 g62683(.A (n_6801), .Y (n_6153));
NAND3X1 g61800(.A (n_5323), .B (g_12922), .C (n_9797), .Y (n_5505));
NAND3X1 g61804(.A (n_5311), .B (n_2255), .C (n_2852), .Y (n_5504));
OAI22X1 g61343(.A0 (n_5068), .A1 (n_9371), .B0 (g2008), .B1 (n_9862),.Y (n_5502));
NAND3X1 g62806(.A (n_5290), .B (g3211), .C (n_8586), .Y (n_5501));
NAND3X1 g62809(.A (n_5289), .B (g3562), .C (n_4682), .Y (n_5500));
OAI22X1 g61347(.A0 (n_5045), .A1 (n_9903), .B0 (g2024), .B1 (n_9811),.Y (n_5499));
OAI22X1 g61346(.A0 (n_5058), .A1 (n_9976), .B0 (g2020), .B1 (n_9664),.Y (n_5497));
OAI22X1 g61348(.A0 (n_5044), .A1 (n_10952), .B0 (g2012), .B1(n_9627), .Y (n_5495));
OAI22X1 g61349(.A0 (n_5039), .A1 (n_9431), .B0 (g1604), .B1 (n_9627),.Y (n_5492));
CLKBUFX1 gbuf_d_307(.A(n_5337), .Y(d_out_307));
CLKBUFX1 gbuf_qn_307(.A(qn_in_307), .Y(g2008));
OAI22X1 g61351(.A0 (n_5030), .A1 (n_9772), .B0 (g1600), .B1 (n_9992),.Y (n_5490));
OAI22X1 g61352(.A0 (n_5022), .A1 (n_9836), .B0 (g1616), .B1 (n_9830),.Y (n_5489));
CLKBUFX1 gbuf_d_308(.A(n_5238), .Y(d_out_308));
CLKBUFX1 gbuf_qn_308(.A(qn_in_308), .Y(g2116));
OAI22X1 g61354(.A0 (n_5019), .A1 (n_9976), .B0 (g1608), .B1(n_10063), .Y (n_5487));
CLKBUFX1 gbuf_d_309(.A(n_5246), .Y(d_out_309));
CLKBUFX1 gbuf_qn_309(.A(qn_in_309), .Y(g1821));
MX2X1 g62925(.A (g4031), .B (n_3430), .S0 (n_9218), .Y (n_5486));
CLKBUFX1 gbuf_d_310(.A(n_5340), .Y(d_out_310));
CLKBUFX1 gbuf_qn_310(.A(qn_in_310), .Y(g1886));
CLKBUFX1 gbuf_d_311(.A(n_5345), .Y(d_out_311));
CLKBUFX1 gbuf_qn_311(.A(qn_in_311), .Y(g1870));
OAI21X1 g60919(.A0 (n_4285), .A1 (n_9693), .B0 (n_5283), .Y (n_5485));
NAND4X1 g61938(.A (n_5288), .B (n_2067), .C (n_9940), .D (n_8777), .Y(n_5483));
NAND3X1 g61948(.A (g4372), .B (g4581), .C (n_9466), .Y (n_6011));
MX2X1 g61966(.A (n_19), .B (n_11196), .S0 (n_3626), .Y (n_5481));
CLKBUFX1 gbuf_d_312(.A(n_5278), .Y(d_out_312));
CLKBUFX1 gbuf_qn_312(.A(qn_in_312), .Y(g2567));
OAI22X1 g63110(.A0 (n_4985), .A1 (n_9269), .B0 (g3827), .B1 (n_9651),.Y (n_5476));
MX2X1 g63111(.A (g3831), .B (n_4971), .S0 (n_9894), .Y (n_5474));
OR4X1 g61153(.A (g4411), .B (g4405), .C (g4375), .D (n_316), .Y(n_5591));
CLKBUFX1 gbuf_d_313(.A(n_5282), .Y(d_out_313));
CLKBUFX1 gbuf_qn_313(.A(qn_in_313), .Y(g2299));
NAND3X1 g61484(.A (n_2564), .B (n_4976), .C (n_4844), .Y (n_5468));
OAI22X1 g61174(.A0 (n_4967), .A1 (n_9903), .B0 (g2181), .B1 (n_9992),.Y (n_5467));
OAI21X1 g61013(.A0 (n_4966), .A1 (n_10952), .B0 (n_3164), .Y(n_5466));
MX2X1 g63335(.A (g_20208), .B (g14147), .S0 (n_5582), .Y (n_5465));
OAI21X1 g61014(.A0 (n_4960), .A1 (n_9693), .B0 (n_3162), .Y (n_5464));
OAI21X1 g61015(.A0 (n_4959), .A1 (n_10078), .B0 (n_3161), .Y(n_5462));
OAI21X1 g61016(.A0 (n_4954), .A1 (n_9672), .B0 (n_3363), .Y (n_5461));
MX2X1 g62127(.A (n_1299), .B (n_5457), .S0 (n_5459), .Y (n_5460));
XOR2X1 g62132(.A (n_2072), .B (n_5457), .Y (n_5458));
CLKBUFX1 gbuf_d_314(.A(g11770), .Y(d_out_314));
CLKBUFX1 gbuf_q_314(.A(q_in_314), .Y(g8915));
OAI22X1 g61554(.A0 (n_4955), .A1 (n_4956), .B0 (n_262), .B1 (n_9627),.Y (n_5456));
NAND2X1 g62243(.A (n_5454), .B (n_5453), .Y (n_5455));
OAI21X1 g60940(.A0 (n_5223), .A1 (n_9628), .B0 (n_3197), .Y (n_5451));
NAND3X1 g61203(.A (n_5258), .B (n_6677), .C (n_9834), .Y (n_5450));
OAI21X1 g60941(.A0 (n_5222), .A1 (n_9371), .B0 (n_3196), .Y (n_5449));
OAI21X1 g60942(.A0 (n_5219), .A1 (n_9903), .B0 (n_3191), .Y (n_5448));
OAI21X1 g60943(.A0 (n_5218), .A1 (n_9775), .B0 (n_3384), .Y (n_5447));
NAND3X1 g61042(.A (n_5259), .B (n_2558), .C (n_4864), .Y (n_5445));
NAND3X1 g61044(.A (n_10548), .B (n_2247), .C (n_10549), .Y (n_5444));
NAND3X1 g63961(.A (n_6897), .B (n_8557), .C (n_11), .Y (n_5665));
NAND3X1 g61046(.A (n_5253), .B (n_2284), .C (n_4611), .Y (n_5442));
CLKBUFX1 gbuf_d_315(.A(n_5291), .Y(d_out_315));
CLKBUFX1 gbuf_q_315(.A(q_in_315), .Y(g1373));
CLKBUFX1 gbuf_d_316(.A(n_5279), .Y(d_out_316));
CLKBUFX1 gbuf_qn_316(.A(qn_in_316), .Y(g2433));
CLKBUFX1 gbuf_d_317(.A(n_5349), .Y(d_out_317));
CLKBUFX1 gbuf_qn_317(.A(qn_in_317), .Y(g1744));
CLKBUFX1 gbuf_d_318(.A(n_5354), .Y(d_out_318));
CLKBUFX1 gbuf_qn_318(.A(qn_in_318), .Y(g1748));
CLKBUFX1 gbuf_d_319(.A(n_5348), .Y(d_out_319));
CLKBUFX1 gbuf_qn_319(.A(qn_in_319), .Y(g1752));
CLKBUFX1 gbuf_d_320(.A(n_5347), .Y(d_out_320));
CLKBUFX1 gbuf_qn_320(.A(qn_in_320), .Y(g1756));
CLKBUFX1 gbuf_d_321(.A(n_5235), .Y(d_out_321));
CLKBUFX1 gbuf_qn_321(.A(qn_in_321), .Y(g1736));
CLKBUFX1 gbuf_d_322(.A(n_5342), .Y(d_out_322));
CLKBUFX1 gbuf_qn_322(.A(qn_in_322), .Y(g1878));
CLKBUFX1 gbuf_d_323(.A(n_5341), .Y(d_out_323));
CLKBUFX1 gbuf_qn_323(.A(qn_in_323), .Y(g1882));
CLKBUFX1 gbuf_d_324(.A(n_5233), .Y(d_out_324));
CLKBUFX1 gbuf_qn_324(.A(qn_in_324), .Y(g1740));
CLKBUFX1 gbuf_d_325(.A(n_5338), .Y(d_out_325));
CLKBUFX1 gbuf_qn_325(.A(qn_in_325), .Y(g1890));
CLKBUFX1 gbuf_d_326(.A(n_5344), .Y(d_out_326));
CLKBUFX1 gbuf_qn_326(.A(qn_in_326), .Y(g1874));
CLKBUFX1 gbuf_d_327(.A(n_5336), .Y(d_out_327));
CLKBUFX1 gbuf_qn_327(.A(qn_in_327), .Y(g2012));
CLKBUFX1 gbuf_d_328(.A(n_5335), .Y(d_out_328));
CLKBUFX1 gbuf_qn_328(.A(qn_in_328), .Y(g1604));
CLKBUFX1 gbuf_d_329(.A(n_5310), .Y(d_out_329));
CLKBUFX1 gbuf_qn_329(.A(qn_in_329), .Y(g_16063));
CLKBUFX1 gbuf_d_330(.A(n_8620), .Y(d_out_330));
CLKBUFX1 gbuf_q_330(.A(q_in_330), .Y(g1183));
CLKBUFX1 gbuf_d_331(.A(n_5270), .Y(d_out_331));
CLKBUFX1 gbuf_q_331(.A(q_in_331), .Y(g_17426));
CLKBUFX1 gbuf_d_332(.A(n_5276), .Y(d_out_332));
CLKBUFX1 gbuf_q_332(.A(q_in_332), .Y(g_20159));
CLKBUFX1 gbuf_d_333(.A(n_5272), .Y(d_out_333));
CLKBUFX1 gbuf_q_333(.A(q_in_333), .Y(g5052));
CLKBUFX1 gbuf_d_334(.A(n_6684), .Y(d_out_334));
CLKBUFX1 gbuf_q_334(.A(q_in_334), .Y(g1862));
CLKBUFX1 gbuf_d_335(.A(n_6866), .Y(d_out_335));
CLKBUFX1 gbuf_q_335(.A(q_in_335), .Y(g1728));
CLKBUFX1 gbuf_d_336(.A(n_5251), .Y(d_out_336));
CLKBUFX1 gbuf_qn_336(.A(qn_in_336), .Y(g2675));
CLKBUFX1 gbuf_d_337(.A(n_5252), .Y(d_out_337));
CLKBUFX1 gbuf_q_337(.A(q_in_337), .Y(g2671));
CLKBUFX1 gbuf_d_338(.A(n_5249), .Y(d_out_338));
CLKBUFX1 gbuf_q_338(.A(q_in_338), .Y(g1710));
CLKBUFX1 gbuf_d_339(.A(n_5248), .Y(d_out_339));
CLKBUFX1 gbuf_qn_339(.A(qn_in_339), .Y(g1714));
CLKBUFX1 gbuf_d_340(.A(n_5245), .Y(d_out_340));
CLKBUFX1 gbuf_q_340(.A(q_in_340), .Y(g1844));
CLKBUFX1 gbuf_d_341(.A(n_5244), .Y(d_out_341));
CLKBUFX1 gbuf_qn_341(.A(qn_in_341), .Y(g1848));
CLKBUFX1 gbuf_d_342(.A(n_5242), .Y(d_out_342));
CLKBUFX1 gbuf_qn_342(.A(qn_in_342), .Y(g1955));
CLKBUFX1 gbuf_d_343(.A(n_5241), .Y(d_out_343));
CLKBUFX1 gbuf_q_343(.A(q_in_343), .Y(g1978));
CLKBUFX1 gbuf_d_344(.A(n_5240), .Y(d_out_344));
CLKBUFX1 gbuf_qn_344(.A(qn_in_344), .Y(g1982));
CLKBUFX1 gbuf_d_345(.A(n_5239), .Y(d_out_345));
CLKBUFX1 gbuf_q_345(.A(q_in_345), .Y(g2112));
CLKBUFX1 gbuf_d_346(.A(n_5236), .Y(d_out_346));
CLKBUFX1 gbuf_qn_346(.A(qn_in_346), .Y(g2265));
CLKBUFX1 gbuf_d_347(.A(n_5355), .Y(d_out_347));
CLKBUFX1 gbuf_qn_347(.A(qn_in_347), .Y(g2407));
CLKBUFX1 gbuf_d_348(.A(n_5353), .Y(d_out_348));
CLKBUFX1 gbuf_q_348(.A(q_in_348), .Y(g2537));
CLKBUFX1 gbuf_d_349(.A(n_5352), .Y(d_out_349));
CLKBUFX1 gbuf_qn_349(.A(qn_in_349), .Y(g2541));
CLKBUFX1 gbuf_d_350(.A(n_5350), .Y(d_out_350));
CLKBUFX1 gbuf_qn_350(.A(qn_in_350), .Y(g2648));
CLKBUFX1 gbuf_d_351(.A(n_5254), .Y(d_out_351));
CLKBUFX1 gbuf_q_351(.A(q_in_351), .Y(g5057));
CLKBUFX1 gbuf_d_352(.A(n_5232), .Y(d_out_352));
CLKBUFX1 gbuf_q_352(.A(q_in_352), .Y(g2403));
CLKBUFX1 gbuf_d_353(.A(n_5331), .Y(d_out_353));
CLKBUFX1 gbuf_q_353(.A(q_in_353), .Y(g3689));
CLKBUFX1 gbuf_d_354(.A(n_5333), .Y(d_out_354));
CLKBUFX1 gbuf_q_354(.A(q_in_354), .Y(g3338));
CLKBUFX1 gbuf_d_355(.A(n_5329), .Y(d_out_355));
CLKBUFX1 gbuf_q_355(.A(q_in_355), .Y(g5252));
CLKBUFX1 gbuf_d_356(.A(n_5328), .Y(d_out_356));
CLKBUFX1 gbuf_q_356(.A(q_in_356), .Y(g5260));
CLKBUFX1 gbuf_d_357(.A(n_5330), .Y(d_out_357));
CLKBUFX1 gbuf_q_357(.A(q_in_357), .Y(g5236));
CLKBUFX1 gbuf_d_358(.A(n_5327), .Y(d_out_358));
CLKBUFX1 gbuf_q_358(.A(q_in_358), .Y(g5264));
CLKBUFX1 gbuf_d_359(.A(n_5326), .Y(d_out_359));
CLKBUFX1 gbuf_q_359(.A(q_in_359), .Y(g5583));
CLKBUFX1 gbuf_d_360(.A(n_5325), .Y(d_out_360));
CLKBUFX1 gbuf_q_360(.A(q_in_360), .Y(g5599));
CLKBUFX1 gbuf_d_361(.A(n_5324), .Y(d_out_361));
CLKBUFX1 gbuf_q_361(.A(q_in_361), .Y(g5929));
CLKBUFX1 gbuf_d_362(.A(n_5321), .Y(d_out_362));
CLKBUFX1 gbuf_q_362(.A(q_in_362), .Y(g5957));
CLKBUFX1 gbuf_d_363(.A(n_5319), .Y(d_out_363));
CLKBUFX1 gbuf_q_363(.A(q_in_363), .Y(g3129));
CLKBUFX1 gbuf_d_364(.A(n_5318), .Y(d_out_364));
CLKBUFX1 gbuf_qn_364(.A(qn_in_364), .Y(g3133));
CLKBUFX1 gbuf_d_365(.A(n_5317), .Y(d_out_365));
CLKBUFX1 gbuf_q_365(.A(q_in_365), .Y(g6275));
CLKBUFX1 gbuf_d_366(.A(n_5315), .Y(d_out_366));
CLKBUFX1 gbuf_q_366(.A(q_in_366), .Y(g6299));
CLKBUFX1 gbuf_d_367(.A(n_5313), .Y(d_out_367));
CLKBUFX1 gbuf_q_367(.A(q_in_367), .Y(g6303));
CLKBUFX1 gbuf_d_368(.A(n_5312), .Y(d_out_368));
CLKBUFX1 gbuf_q_368(.A(q_in_368), .Y(g6307));
CLKBUFX1 gbuf_d_369(.A(n_5309), .Y(d_out_369));
CLKBUFX1 gbuf_q_369(.A(q_in_369), .Y(g6637));
CLKBUFX1 gbuf_d_370(.A(n_5308), .Y(d_out_370));
CLKBUFX1 gbuf_q_370(.A(q_in_370), .Y(g6645));
CLKBUFX1 gbuf_d_371(.A(n_5307), .Y(d_out_371));
CLKBUFX1 gbuf_q_371(.A(q_in_371), .Y(g3480));
CLKBUFX1 gbuf_d_372(.A(n_5306), .Y(d_out_372));
CLKBUFX1 gbuf_qn_372(.A(qn_in_372), .Y(g3484));
CLKBUFX1 gbuf_d_373(.A(n_5304), .Y(d_out_373));
CLKBUFX1 gbuf_q_373(.A(q_in_373), .Y(g2040));
CLKBUFX1 gbuf_d_374(.A(n_5302), .Y(d_out_374));
CLKBUFX1 gbuf_q_374(.A(q_in_374), .Y(g2070));
CLKBUFX1 gbuf_d_375(.A(n_5300), .Y(d_out_375));
CLKBUFX1 gbuf_q_375(.A(q_in_375), .Y(g3945));
CLKBUFX1 gbuf_d_376(.A(n_5299), .Y(d_out_376));
CLKBUFX1 gbuf_q_376(.A(q_in_376), .Y(g3953));
CLKBUFX1 gbuf_d_377(.A(n_5339), .Y(d_out_377));
CLKBUFX1 gbuf_q_377(.A(q_in_377), .Y(g1592));
CLKBUFX1 gbuf_d_378(.A(n_5297), .Y(d_out_378));
CLKBUFX1 gbuf_q_378(.A(q_in_378), .Y(g1636));
CLKBUFX1 gbuf_d_379(.A(n_5296), .Y(d_out_379));
CLKBUFX1 gbuf_q_379(.A(q_in_379), .Y(g2599));
CLKBUFX1 gbuf_d_380(.A(n_5294), .Y(d_out_380));
CLKBUFX1 gbuf_q_380(.A(q_in_380), .Y(n_4120));
CLKBUFX1 gbuf_d_381(.A(n_5293), .Y(d_out_381));
CLKBUFX1 gbuf_q_381(.A(q_in_381), .Y(g2629));
CLKBUFX1 gbuf_d_382(.A(n_5275), .Y(d_out_382));
CLKBUFX1 gbuf_q_382(.A(q_in_382), .Y(g4473));
INVX1 g64074(.A (n_6280), .Y (n_5440));
CLKBUFX1 gbuf_d_383(.A(n_5247), .Y(d_out_383));
CLKBUFX1 gbuf_q_383(.A(q_in_383), .Y(g2756));
NAND3X1 g61739(.A (n_2797), .B (n_4921), .C (n_4961), .Y (n_5437));
INVX1 g64379(.A (n_5436), .Y (n_5559));
CLKBUFX1 gbuf_d_384(.A(n_5127), .Y(d_out_384));
CLKBUFX1 gbuf_q_384(.A(q_in_384), .Y(g6287));
OAI21X1 g62792(.A0 (n_4896), .A1 (n_5007), .B0 (n_4990), .Y (n_5432));
AOI22X1 g61839(.A0 (n_2265), .A1 (n_6549), .B0 (g_19659), .B1(n_10376), .Y (n_5431));
NAND2X1 g62824(.A (n_4889), .B (n_4991), .Y (n_5430));
CLKBUFX1 gbuf_d_385(.A(n_4943), .Y(d_out_385));
CLKBUFX1 gbuf_qn_385(.A(qn_in_385), .Y(g2399));
CLKBUFX1 gbuf_d_386(.A(n_5135), .Y(d_out_386));
CLKBUFX1 gbuf_q_386(.A(q_in_386), .Y(g6255));
OAI22X1 g61353(.A0 (n_4913), .A1 (n_9903), .B0 (g1620), .B1 (n_9862),.Y (n_5428));
NAND4X1 g62914(.A (g3546), .B (n_10576), .C (n_10897), .D (g3680), .Y(n_5425));
CLKBUFX1 gbuf_d_387(.A(n_5141), .Y(d_out_387));
CLKBUFX1 gbuf_q_387(.A(q_in_387), .Y(g6239));
CLKBUFX1 gbuf_d_388(.A(n_5050), .Y(d_out_388));
CLKBUFX1 gbuf_q_388(.A(q_in_388), .Y(g3602));
CLKBUFX1 gbuf_d_389(.A(n_5052), .Y(d_out_389));
CLKBUFX1 gbuf_q_389(.A(q_in_389), .Y(g3594));
CLKBUFX1 gbuf_d_390(.A(n_5150), .Y(d_out_390));
CLKBUFX1 gbuf_q_390(.A(q_in_390), .Y(g5949));
CLKBUFX1 gbuf_d_391(.A(n_5155), .Y(d_out_391));
CLKBUFX1 gbuf_q_391(.A(q_in_391), .Y(g5933));
CLKBUFX1 gbuf_d_392(.A(n_5159), .Y(d_out_392));
CLKBUFX1 gbuf_q_392(.A(q_in_392), .Y(g5917));
NAND3X1 g60918(.A (n_5000), .B (n_2288), .C (n_4888), .Y (n_5424));
CLKBUFX1 gbuf_d_393(.A(n_5059), .Y(d_out_393));
CLKBUFX1 gbuf_q_393(.A(q_in_393), .Y(g3578));
NAND2X1 g61918(.A (n_4999), .B (n_4911), .Y (n_5423));
AOI21X1 g61934(.A0 (n_4874), .A1 (n_3769), .B0 (g4961), .Y (n_5422));
MX2X1 g61967(.A (n_843), .B (n_7329), .S0 (n_3547), .Y (n_5420));
CLKBUFX1 gbuf_d_394(.A(n_5173), .Y(d_out_394));
CLKBUFX1 gbuf_q_394(.A(q_in_394), .Y(g5607));
MX2X1 g63109(.A (g3821), .B (n_4886), .S0 (n_9091), .Y (n_5415));
MX2X1 g63132(.A (g2204), .B (n_4884), .S0 (n_10005), .Y (n_5414));
MX2X1 g63133(.A (g2197), .B (n_4881), .S0 (n_9000), .Y (n_5412));
NAND3X1 g62031(.A (n_4974), .B (n_2526), .C (n_4842), .Y (n_5411));
NAND2X1 g63219(.A (n_4879), .B (n_4987), .Y (n_5410));
XOR2X1 g61167(.A (g4382), .B (g4375), .Y (n_5409));
AOI21X1 g62074(.A0 (n_4021), .A1 (n_4982), .B0 (n_4983), .Y (n_5408));
AOI21X1 g62075(.A0 (n_4020), .A1 (n_4980), .B0 (n_4981), .Y (n_5407));
AOI21X1 g62076(.A0 (n_4019), .A1 (n_4978), .B0 (n_4979), .Y (n_5406));
AOI21X1 g62077(.A0 (n_4018), .A1 (n_11070), .B0 (n_4977), .Y(n_5405));
MX2X1 g61171(.A (n_4906), .B (n_4865), .S0 (n_9358), .Y (n_5404));
NAND4X1 g63298(.A (g3949), .B (n_5402), .C (g16748), .D (n_8917), .Y(n_5403));
OAI22X1 g61176(.A0 (n_4861), .A1 (n_9505), .B0 (g2299), .B1 (n_9651),.Y (n_5400));
OAI22X1 g61178(.A0 (n_4860), .A1 (n_9599), .B0 (g2295), .B1 (n_9992),.Y (n_5398));
MX2X1 g63370(.A (n_11106), .B (n_4857), .S0 (n_8955), .Y (n_5397));
OAI22X1 g61179(.A0 (n_4859), .A1 (n_10952), .B0 (g2311), .B1(n_9992), .Y (n_5396));
CLKBUFX1 gbuf_d_395(.A(n_5064), .Y(d_out_395));
CLKBUFX1 gbuf_q_395(.A(q_in_395), .Y(g3562));
CLKBUFX1 gbuf_d_396(.A(g14147), .Y(d_out_396));
CLKBUFX1 gbuf_q_396(.A(q_in_396), .Y(g14167));
OAI22X1 g61180(.A0 (n_4858), .A1 (n_10078), .B0 (g2315), .B1(n_9830), .Y (n_5395));
OAI22X1 g61181(.A0 (n_4856), .A1 (n_9903), .B0 (g2303), .B1 (n_9992),.Y (n_5394));
NAND3X1 g61517(.A (n_2543), .B (n_4820), .C (n_4875), .Y (n_5393));
OAI22X1 g61183(.A0 (n_4930), .A1 (n_9505), .B0 (g2433), .B1 (n_9811),.Y (n_5392));
OAI22X1 g61185(.A0 (n_4854), .A1 (n_9928), .B0 (g2429), .B1 (n_9992),.Y (n_5391));
OAI22X1 g61186(.A0 (n_4853), .A1 (n_9884), .B0 (g2445), .B1 (n_9862),.Y (n_5388));
OAI22X1 g61187(.A0 (n_4852), .A1 (n_9599), .B0 (g2449), .B1 (n_9811),.Y (n_5387));
OAI22X1 g61188(.A0 (n_4851), .A1 (n_9461), .B0 (g2437), .B1 (n_9651),.Y (n_5386));
OAI22X1 g61189(.A0 (n_4850), .A1 (n_9461), .B0 (g2567), .B1 (n_9992),.Y (n_5385));
CLKBUFX1 gbuf_d_397(.A(n_5184), .Y(d_out_397));
CLKBUFX1 gbuf_q_397(.A(q_in_397), .Y(g5567));
OAI22X1 g61191(.A0 (n_4849), .A1 (n_9431), .B0 (g2563), .B1 (n_9862),.Y (n_5384));
OAI22X1 g61192(.A0 (n_4847), .A1 (n_10952), .B0 (g2579), .B1(n_9992), .Y (n_5383));
OAI22X1 g61193(.A0 (n_4846), .A1 (n_9193), .B0 (g2583), .B1 (n_9862),.Y (n_5382));
OAI22X1 g61194(.A0 (n_4845), .A1 (n_9269), .B0 (g2571), .B1 (n_9992),.Y (n_5380));
NOR2X1 g62241(.A (n_5374), .B (n_5378), .Y (n_5379));
NAND3X1 g61200(.A (n_4965), .B (n_10911), .C (n_9558), .Y (n_5377));
NOR2X1 g62263(.A (n_595), .B (n_5374), .Y (n_5375));
NAND3X1 g61210(.A (n_4962), .B (n_4296), .C (n_9209), .Y (n_5373));
CLKBUFX1 gbuf_d_398(.A(n_5015), .Y(d_out_398));
CLKBUFX1 gbuf_q_398(.A(q_in_398), .Y(g2465));
OAI21X1 g62284(.A0 (n_95), .A1 (n_9333), .B0 (n_4964), .Y (n_5372));
CLKBUFX1 gbuf_d_399(.A(n_5021), .Y(d_out_399));
CLKBUFX1 gbuf_q_399(.A(q_in_399), .Y(g3961));
NAND3X1 g63924(.A (g_13255), .B (g_16983), .C (n_9811), .Y (n_5370));
NAND3X1 g61045(.A (n_4953), .B (n_2533), .C (n_4308), .Y (n_5369));
CLKBUFX1 gbuf_d_400(.A(n_5076), .Y(d_out_400));
CLKBUFX1 gbuf_q_400(.A(q_in_400), .Y(g6653));
CLKBUFX1 gbuf_d_401(.A(n_4986), .Y(d_out_401));
CLKBUFX1 gbuf_q_401(.A(q_in_401), .Y(n_10197));
CLKBUFX1 gbuf_d_402(.A(n_4975), .Y(d_out_402));
CLKBUFX1 gbuf_qn_402(.A(qn_in_402), .Y(g1413));
CLKBUFX1 gbuf_d_403(.A(n_4972), .Y(d_out_403));
CLKBUFX1 gbuf_q_403(.A(q_in_403), .Y(g_14342));
CLKBUFX1 gbuf_d_404(.A(n_4957), .Y(d_out_404));
CLKBUFX1 gbuf_q_404(.A(q_in_404), .Y(g4601));
CLKBUFX1 gbuf_d_405(.A(n_5037), .Y(d_out_405));
CLKBUFX1 gbuf_q_405(.A(q_in_405), .Y(g3909));
CLKBUFX1 gbuf_d_406(.A(n_5085), .Y(d_out_406));
CLKBUFX1 gbuf_q_406(.A(q_in_406), .Y(g3259));
CLKBUFX1 gbuf_d_407(.A(n_5025), .Y(d_out_407));
CLKBUFX1 gbuf_q_407(.A(q_in_407), .Y(g3941));
CLKBUFX1 gbuf_d_408(.A(n_5088), .Y(d_out_408));
CLKBUFX1 gbuf_q_408(.A(q_in_408), .Y(g6617));
CLKBUFX1 gbuf_d_409(.A(n_5023), .Y(d_out_409));
CLKBUFX1 gbuf_q_409(.A(q_in_409), .Y(g3957));
CLKBUFX1 gbuf_d_410(.A(n_5093), .Y(d_out_410));
CLKBUFX1 gbuf_q_410(.A(q_in_410), .Y(g6605));
CLKBUFX1 gbuf_d_411(.A(n_5195), .Y(d_out_411));
CLKBUFX1 gbuf_q_411(.A(q_in_411), .Y(g5268));
CLKBUFX1 gbuf_d_412(.A(n_5122), .Y(d_out_412));
CLKBUFX1 gbuf_q_412(.A(q_in_412), .Y(g3191));
CLKBUFX1 gbuf_d_413(.A(n_5106), .Y(d_out_413));
CLKBUFX1 gbuf_q_413(.A(q_in_413), .Y(g6581));
CLKBUFX1 gbuf_d_414(.A(n_5197), .Y(d_out_414));
CLKBUFX1 gbuf_q_414(.A(q_in_414), .Y(g5256));
CLKBUFX1 gbuf_d_415(.A(n_5204), .Y(d_out_415));
CLKBUFX1 gbuf_q_415(.A(q_in_415), .Y(g5228));
CLKBUFX1 gbuf_d_416(.A(n_5009), .Y(d_out_416));
CLKBUFX1 gbuf_q_416(.A(q_in_416), .Y(g_15016));
CLKBUFX1 gbuf_d_417(.A(n_5207), .Y(d_out_417));
CLKBUFX1 gbuf_q_417(.A(q_in_417), .Y(g5216));
CLKBUFX1 gbuf_d_418(.A(n_4952), .Y(d_out_418));
CLKBUFX1 gbuf_qn_418(.A(qn_in_418), .Y(g1687));
CLKBUFX1 gbuf_d_419(.A(n_4951), .Y(d_out_419));
CLKBUFX1 gbuf_qn_419(.A(qn_in_419), .Y(g2667));
CLKBUFX1 gbuf_d_420(.A(n_4950), .Y(d_out_420));
CLKBUFX1 gbuf_qn_420(.A(qn_in_420), .Y(g1706));
CLKBUFX1 gbuf_d_421(.A(n_4949), .Y(d_out_421));
CLKBUFX1 gbuf_qn_421(.A(qn_in_421), .Y(g1840));
CLKBUFX1 gbuf_d_422(.A(n_4947), .Y(d_out_422));
CLKBUFX1 gbuf_qn_422(.A(qn_in_422), .Y(g1974));
CLKBUFX1 gbuf_d_423(.A(n_4945), .Y(d_out_423));
CLKBUFX1 gbuf_qn_423(.A(qn_in_423), .Y(g2108));
CLKBUFX1 gbuf_d_424(.A(n_4944), .Y(d_out_424));
CLKBUFX1 gbuf_qn_424(.A(qn_in_424), .Y(g2380));
CLKBUFX1 gbuf_d_425(.A(n_5231), .Y(d_out_425));
CLKBUFX1 gbuf_qn_425(.A(qn_in_425), .Y(g2514));
CLKBUFX1 gbuf_d_426(.A(n_5230), .Y(d_out_426));
CLKBUFX1 gbuf_qn_426(.A(qn_in_426), .Y(g2533));
CLKBUFX1 gbuf_d_427(.A(n_5214), .Y(d_out_427));
CLKBUFX1 gbuf_q_427(.A(q_in_427), .Y(g5196));
CLKBUFX1 gbuf_d_428(.A(n_5213), .Y(d_out_428));
CLKBUFX1 gbuf_q_428(.A(q_in_428), .Y(g5200));
CLKBUFX1 gbuf_d_429(.A(n_5210), .Y(d_out_429));
CLKBUFX1 gbuf_q_429(.A(q_in_429), .Y(g5208));
CLKBUFX1 gbuf_d_430(.A(n_5209), .Y(d_out_430));
CLKBUFX1 gbuf_q_430(.A(q_in_430), .Y(g5212));
CLKBUFX1 gbuf_d_431(.A(n_5212), .Y(d_out_431));
CLKBUFX1 gbuf_q_431(.A(q_in_431), .Y(g5204));
CLKBUFX1 gbuf_d_432(.A(n_5205), .Y(d_out_432));
CLKBUFX1 gbuf_q_432(.A(q_in_432), .Y(g5224));
CLKBUFX1 gbuf_d_433(.A(n_5206), .Y(d_out_433));
CLKBUFX1 gbuf_q_433(.A(q_in_433), .Y(g5220));
CLKBUFX1 gbuf_d_434(.A(n_5201), .Y(d_out_434));
CLKBUFX1 gbuf_q_434(.A(q_in_434), .Y(g5240));
CLKBUFX1 gbuf_d_435(.A(n_5200), .Y(d_out_435));
CLKBUFX1 gbuf_q_435(.A(q_in_435), .Y(g5244));
CLKBUFX1 gbuf_d_436(.A(n_5199), .Y(d_out_436));
CLKBUFX1 gbuf_q_436(.A(q_in_436), .Y(g5248));
CLKBUFX1 gbuf_d_437(.A(n_5202), .Y(d_out_437));
CLKBUFX1 gbuf_q_437(.A(q_in_437), .Y(g5232));
CLKBUFX1 gbuf_d_438(.A(n_5193), .Y(d_out_438));
CLKBUFX1 gbuf_q_438(.A(q_in_438), .Y(g5272));
CLKBUFX1 gbuf_d_439(.A(n_5190), .Y(d_out_439));
CLKBUFX1 gbuf_q_439(.A(q_in_439), .Y(g5547));
CLKBUFX1 gbuf_d_440(.A(n_5189), .Y(d_out_440));
CLKBUFX1 gbuf_q_440(.A(q_in_440), .Y(g5551));
CLKBUFX1 gbuf_d_441(.A(n_5187), .Y(d_out_441));
CLKBUFX1 gbuf_q_441(.A(q_in_441), .Y(g5555));
CLKBUFX1 gbuf_d_442(.A(n_5186), .Y(d_out_442));
CLKBUFX1 gbuf_q_442(.A(q_in_442), .Y(g5559));
CLKBUFX1 gbuf_d_443(.A(n_5185), .Y(d_out_443));
CLKBUFX1 gbuf_q_443(.A(q_in_443), .Y(g5563));
CLKBUFX1 gbuf_d_444(.A(n_5183), .Y(d_out_444));
CLKBUFX1 gbuf_q_444(.A(q_in_444), .Y(g5571));
CLKBUFX1 gbuf_d_445(.A(n_5182), .Y(d_out_445));
CLKBUFX1 gbuf_q_445(.A(q_in_445), .Y(g5575));
CLKBUFX1 gbuf_d_446(.A(n_5181), .Y(d_out_446));
CLKBUFX1 gbuf_q_446(.A(q_in_446), .Y(g5579));
CLKBUFX1 gbuf_d_447(.A(n_5192), .Y(d_out_447));
CLKBUFX1 gbuf_q_447(.A(q_in_447), .Y(g5543));
CLKBUFX1 gbuf_d_448(.A(n_5177), .Y(d_out_448));
CLKBUFX1 gbuf_q_448(.A(q_in_448), .Y(g5591));
CLKBUFX1 gbuf_d_449(.A(n_5175), .Y(d_out_449));
CLKBUFX1 gbuf_q_449(.A(q_in_449), .Y(g5595));
CLKBUFX1 gbuf_d_450(.A(n_5179), .Y(d_out_450));
CLKBUFX1 gbuf_q_450(.A(q_in_450), .Y(g5587));
CLKBUFX1 gbuf_d_451(.A(n_5174), .Y(d_out_451));
CLKBUFX1 gbuf_q_451(.A(q_in_451), .Y(g5603));
CLKBUFX1 gbuf_d_452(.A(n_5172), .Y(d_out_452));
CLKBUFX1 gbuf_q_452(.A(q_in_452), .Y(g5611));
CLKBUFX1 gbuf_d_453(.A(n_5171), .Y(d_out_453));
CLKBUFX1 gbuf_q_453(.A(q_in_453), .Y(g5615));
CLKBUFX1 gbuf_d_454(.A(n_5170), .Y(d_out_454));
CLKBUFX1 gbuf_q_454(.A(q_in_454), .Y(g5619));
CLKBUFX1 gbuf_d_455(.A(n_5168), .Y(d_out_455));
CLKBUFX1 gbuf_q_455(.A(q_in_455), .Y(g5889));
CLKBUFX1 gbuf_d_456(.A(n_5165), .Y(d_out_456));
CLKBUFX1 gbuf_q_456(.A(q_in_456), .Y(g5897));
CLKBUFX1 gbuf_d_457(.A(n_5164), .Y(d_out_457));
CLKBUFX1 gbuf_q_457(.A(q_in_457), .Y(g5901));
CLKBUFX1 gbuf_d_458(.A(n_5163), .Y(d_out_458));
CLKBUFX1 gbuf_q_458(.A(q_in_458), .Y(g5905));
CLKBUFX1 gbuf_d_459(.A(n_5161), .Y(d_out_459));
CLKBUFX1 gbuf_q_459(.A(q_in_459), .Y(g5909));
CLKBUFX1 gbuf_d_460(.A(n_5160), .Y(d_out_460));
CLKBUFX1 gbuf_q_460(.A(q_in_460), .Y(g5913));
CLKBUFX1 gbuf_d_461(.A(n_5167), .Y(d_out_461));
CLKBUFX1 gbuf_q_461(.A(q_in_461), .Y(g5893));
CLKBUFX1 gbuf_d_462(.A(n_5158), .Y(d_out_462));
CLKBUFX1 gbuf_q_462(.A(q_in_462), .Y(g5921));
CLKBUFX1 gbuf_d_463(.A(n_5156), .Y(d_out_463));
CLKBUFX1 gbuf_q_463(.A(q_in_463), .Y(g5925));
CLKBUFX1 gbuf_d_464(.A(n_5154), .Y(d_out_464));
CLKBUFX1 gbuf_q_464(.A(q_in_464), .Y(g5937));
CLKBUFX1 gbuf_d_465(.A(n_5152), .Y(d_out_465));
CLKBUFX1 gbuf_q_465(.A(q_in_465), .Y(g5941));
CLKBUFX1 gbuf_d_466(.A(n_5151), .Y(d_out_466));
CLKBUFX1 gbuf_q_466(.A(q_in_466), .Y(g5945));
CLKBUFX1 gbuf_d_467(.A(n_5149), .Y(d_out_467));
CLKBUFX1 gbuf_q_467(.A(q_in_467), .Y(g5953));
CLKBUFX1 gbuf_d_468(.A(n_5148), .Y(d_out_468));
CLKBUFX1 gbuf_q_468(.A(q_in_468), .Y(g5961));
CLKBUFX1 gbuf_d_469(.A(n_5146), .Y(d_out_469));
CLKBUFX1 gbuf_q_469(.A(q_in_469), .Y(g5965));
CLKBUFX1 gbuf_d_470(.A(n_5144), .Y(d_out_470));
CLKBUFX1 gbuf_qn_470(.A(qn_in_470), .Y(g3125));
CLKBUFX1 gbuf_d_471(.A(n_5143), .Y(d_out_471));
CLKBUFX1 gbuf_q_471(.A(q_in_471), .Y(g6235));
CLKBUFX1 gbuf_d_472(.A(n_5139), .Y(d_out_472));
CLKBUFX1 gbuf_q_472(.A(q_in_472), .Y(g6243));
CLKBUFX1 gbuf_d_473(.A(n_5137), .Y(d_out_473));
CLKBUFX1 gbuf_q_473(.A(q_in_473), .Y(g6247));
CLKBUFX1 gbuf_d_474(.A(n_5136), .Y(d_out_474));
CLKBUFX1 gbuf_q_474(.A(q_in_474), .Y(g6251));
CLKBUFX1 gbuf_d_475(.A(n_5134), .Y(d_out_475));
CLKBUFX1 gbuf_q_475(.A(q_in_475), .Y(g6259));
CLKBUFX1 gbuf_d_476(.A(n_5131), .Y(d_out_476));
CLKBUFX1 gbuf_q_476(.A(q_in_476), .Y(g6267));
CLKBUFX1 gbuf_d_477(.A(n_5130), .Y(d_out_477));
CLKBUFX1 gbuf_q_477(.A(q_in_477), .Y(g6271));
CLKBUFX1 gbuf_d_478(.A(n_5133), .Y(d_out_478));
CLKBUFX1 gbuf_q_478(.A(q_in_478), .Y(g6263));
CLKBUFX1 gbuf_d_479(.A(n_5129), .Y(d_out_479));
CLKBUFX1 gbuf_q_479(.A(q_in_479), .Y(g6279));
CLKBUFX1 gbuf_d_480(.A(n_5128), .Y(d_out_480));
CLKBUFX1 gbuf_q_480(.A(q_in_480), .Y(g6283));
CLKBUFX1 gbuf_d_481(.A(n_5126), .Y(d_out_481));
CLKBUFX1 gbuf_q_481(.A(q_in_481), .Y(g6291));
CLKBUFX1 gbuf_d_482(.A(n_5125), .Y(d_out_482));
CLKBUFX1 gbuf_q_482(.A(q_in_482), .Y(g6295));
CLKBUFX1 gbuf_d_483(.A(n_5123), .Y(d_out_483));
CLKBUFX1 gbuf_q_483(.A(q_in_483), .Y(g3187));
CLKBUFX1 gbuf_d_484(.A(n_5124), .Y(d_out_484));
CLKBUFX1 gbuf_q_484(.A(q_in_484), .Y(g6311));
CLKBUFX1 gbuf_d_485(.A(n_5121), .Y(d_out_485));
CLKBUFX1 gbuf_q_485(.A(q_in_485), .Y(g3195));
CLKBUFX1 gbuf_d_486(.A(n_5119), .Y(d_out_486));
CLKBUFX1 gbuf_q_486(.A(q_in_486), .Y(g3199));
CLKBUFX1 gbuf_d_487(.A(n_5118), .Y(d_out_487));
CLKBUFX1 gbuf_q_487(.A(q_in_487), .Y(g3203));
CLKBUFX1 gbuf_d_488(.A(n_5116), .Y(d_out_488));
CLKBUFX1 gbuf_q_488(.A(q_in_488), .Y(g3207));
CLKBUFX1 gbuf_d_489(.A(n_5115), .Y(d_out_489));
CLKBUFX1 gbuf_q_489(.A(q_in_489), .Y(g3211));
CLKBUFX1 gbuf_d_490(.A(n_5113), .Y(d_out_490));
CLKBUFX1 gbuf_q_490(.A(q_in_490), .Y(g3215));
CLKBUFX1 gbuf_d_491(.A(n_5112), .Y(d_out_491));
CLKBUFX1 gbuf_q_491(.A(q_in_491), .Y(g3219));
CLKBUFX1 gbuf_d_492(.A(n_5111), .Y(d_out_492));
CLKBUFX1 gbuf_q_492(.A(q_in_492), .Y(g3223));
CLKBUFX1 gbuf_d_493(.A(n_5110), .Y(d_out_493));
CLKBUFX1 gbuf_q_493(.A(q_in_493), .Y(g3227));
CLKBUFX1 gbuf_d_494(.A(n_5109), .Y(d_out_494));
CLKBUFX1 gbuf_q_494(.A(q_in_494), .Y(g3231));
CLKBUFX1 gbuf_d_495(.A(n_5107), .Y(d_out_495));
CLKBUFX1 gbuf_q_495(.A(q_in_495), .Y(g3235));
CLKBUFX1 gbuf_d_496(.A(n_5104), .Y(d_out_496));
CLKBUFX1 gbuf_q_496(.A(q_in_496), .Y(g3239));
CLKBUFX1 gbuf_d_497(.A(n_5103), .Y(d_out_497));
CLKBUFX1 gbuf_q_497(.A(q_in_497), .Y(g6585));
CLKBUFX1 gbuf_d_498(.A(n_5101), .Y(d_out_498));
CLKBUFX1 gbuf_q_498(.A(q_in_498), .Y(g3243));
CLKBUFX1 gbuf_d_499(.A(n_5100), .Y(d_out_499));
CLKBUFX1 gbuf_q_499(.A(q_in_499), .Y(g6589));
CLKBUFX1 gbuf_d_500(.A(n_5098), .Y(d_out_500));
CLKBUFX1 gbuf_q_500(.A(q_in_500), .Y(g6593));
CLKBUFX1 gbuf_d_501(.A(n_5097), .Y(d_out_501));
CLKBUFX1 gbuf_q_501(.A(q_in_501), .Y(g3247));
CLKBUFX1 gbuf_d_502(.A(n_5095), .Y(d_out_502));
CLKBUFX1 gbuf_q_502(.A(q_in_502), .Y(g6597));
CLKBUFX1 gbuf_d_503(.A(n_5094), .Y(d_out_503));
CLKBUFX1 gbuf_q_503(.A(q_in_503), .Y(g6601));
CLKBUFX1 gbuf_d_504(.A(n_5092), .Y(d_out_504));
CLKBUFX1 gbuf_q_504(.A(q_in_504), .Y(g6609));
CLKBUFX1 gbuf_d_505(.A(n_5091), .Y(d_out_505));
CLKBUFX1 gbuf_q_505(.A(q_in_505), .Y(g3251));
CLKBUFX1 gbuf_d_506(.A(n_5090), .Y(d_out_506));
CLKBUFX1 gbuf_q_506(.A(q_in_506), .Y(g6613));
CLKBUFX1 gbuf_d_507(.A(n_5087), .Y(d_out_507));
CLKBUFX1 gbuf_q_507(.A(q_in_507), .Y(g3255));
CLKBUFX1 gbuf_d_508(.A(n_5086), .Y(d_out_508));
CLKBUFX1 gbuf_q_508(.A(q_in_508), .Y(g6621));
CLKBUFX1 gbuf_d_509(.A(n_5084), .Y(d_out_509));
CLKBUFX1 gbuf_q_509(.A(q_in_509), .Y(g6625));
CLKBUFX1 gbuf_d_510(.A(n_5082), .Y(d_out_510));
CLKBUFX1 gbuf_q_510(.A(q_in_510), .Y(g3263));
CLKBUFX1 gbuf_d_511(.A(n_5081), .Y(d_out_511));
CLKBUFX1 gbuf_q_511(.A(q_in_511), .Y(g6633));
CLKBUFX1 gbuf_d_512(.A(n_5083), .Y(d_out_512));
CLKBUFX1 gbuf_q_512(.A(q_in_512), .Y(g6629));
CLKBUFX1 gbuf_d_513(.A(n_5079), .Y(d_out_513));
CLKBUFX1 gbuf_q_513(.A(q_in_513), .Y(g6641));
CLKBUFX1 gbuf_d_514(.A(n_5077), .Y(d_out_514));
CLKBUFX1 gbuf_q_514(.A(q_in_514), .Y(g6649));
CLKBUFX1 gbuf_d_515(.A(n_5075), .Y(d_out_515));
CLKBUFX1 gbuf_q_515(.A(q_in_515), .Y(g6657));
CLKBUFX1 gbuf_d_516(.A(n_5016), .Y(d_out_516));
CLKBUFX1 gbuf_qn_516(.A(qn_in_516), .Y(g3476));
CLKBUFX1 gbuf_d_517(.A(n_5073), .Y(d_out_517));
CLKBUFX1 gbuf_q_517(.A(q_in_517), .Y(g3538));
CLKBUFX1 gbuf_d_518(.A(n_5072), .Y(d_out_518));
CLKBUFX1 gbuf_q_518(.A(q_in_518), .Y(g3542));
CLKBUFX1 gbuf_d_519(.A(n_5071), .Y(d_out_519));
CLKBUFX1 gbuf_q_519(.A(q_in_519), .Y(g3546));
CLKBUFX1 gbuf_d_520(.A(n_5069), .Y(d_out_520));
CLKBUFX1 gbuf_q_520(.A(q_in_520), .Y(g3550));
CLKBUFX1 gbuf_d_521(.A(n_5067), .Y(d_out_521));
CLKBUFX1 gbuf_q_521(.A(q_in_521), .Y(g3554));
CLKBUFX1 gbuf_d_522(.A(n_5065), .Y(d_out_522));
CLKBUFX1 gbuf_q_522(.A(q_in_522), .Y(g3558));
CLKBUFX1 gbuf_d_523(.A(n_5063), .Y(d_out_523));
CLKBUFX1 gbuf_q_523(.A(q_in_523), .Y(g3566));
CLKBUFX1 gbuf_d_524(.A(n_5062), .Y(d_out_524));
CLKBUFX1 gbuf_q_524(.A(q_in_524), .Y(g3570));
CLKBUFX1 gbuf_d_525(.A(n_5060), .Y(d_out_525));
CLKBUFX1 gbuf_q_525(.A(q_in_525), .Y(g3574));
CLKBUFX1 gbuf_d_526(.A(n_5056), .Y(d_out_526));
CLKBUFX1 gbuf_q_526(.A(q_in_526), .Y(g3582));
CLKBUFX1 gbuf_d_527(.A(n_5055), .Y(d_out_527));
CLKBUFX1 gbuf_q_527(.A(q_in_527), .Y(g3586));
CLKBUFX1 gbuf_d_528(.A(n_5053), .Y(d_out_528));
CLKBUFX1 gbuf_q_528(.A(q_in_528), .Y(g3590));
CLKBUFX1 gbuf_d_529(.A(n_5048), .Y(d_out_529));
CLKBUFX1 gbuf_q_529(.A(q_in_529), .Y(g3606));
CLKBUFX1 gbuf_d_530(.A(n_5047), .Y(d_out_530));
CLKBUFX1 gbuf_q_530(.A(q_in_530), .Y(g3610));
CLKBUFX1 gbuf_d_531(.A(n_5046), .Y(d_out_531));
CLKBUFX1 gbuf_q_531(.A(q_in_531), .Y(g3614));
CLKBUFX1 gbuf_d_532(.A(n_5051), .Y(d_out_532));
CLKBUFX1 gbuf_q_532(.A(q_in_532), .Y(g3598));
CLKBUFX1 gbuf_d_533(.A(n_5043), .Y(d_out_533));
CLKBUFX1 gbuf_q_533(.A(q_in_533), .Y(g3889));
CLKBUFX1 gbuf_d_534(.A(n_5042), .Y(d_out_534));
CLKBUFX1 gbuf_q_534(.A(q_in_534), .Y(g3893));
CLKBUFX1 gbuf_d_535(.A(n_5041), .Y(d_out_535));
CLKBUFX1 gbuf_q_535(.A(q_in_535), .Y(g3897));
CLKBUFX1 gbuf_d_536(.A(n_5040), .Y(d_out_536));
CLKBUFX1 gbuf_q_536(.A(q_in_536), .Y(g3901));
CLKBUFX1 gbuf_d_537(.A(n_5038), .Y(d_out_537));
CLKBUFX1 gbuf_q_537(.A(q_in_537), .Y(g3905));
CLKBUFX1 gbuf_d_538(.A(n_5032), .Y(d_out_538));
CLKBUFX1 gbuf_q_538(.A(q_in_538), .Y(g3925));
CLKBUFX1 gbuf_d_539(.A(n_5029), .Y(d_out_539));
CLKBUFX1 gbuf_q_539(.A(q_in_539), .Y(g3929));
CLKBUFX1 gbuf_d_540(.A(n_5028), .Y(d_out_540));
CLKBUFX1 gbuf_q_540(.A(q_in_540), .Y(g3933));
CLKBUFX1 gbuf_d_541(.A(n_5026), .Y(d_out_541));
CLKBUFX1 gbuf_q_541(.A(q_in_541), .Y(g3937));
CLKBUFX1 gbuf_d_542(.A(n_5033), .Y(d_out_542));
CLKBUFX1 gbuf_q_542(.A(q_in_542), .Y(g3921));
CLKBUFX1 gbuf_d_543(.A(n_5024), .Y(d_out_543));
CLKBUFX1 gbuf_q_543(.A(q_in_543), .Y(g3949));
CLKBUFX1 gbuf_d_544(.A(n_5035), .Y(d_out_544));
CLKBUFX1 gbuf_q_544(.A(q_in_544), .Y(g3913));
CLKBUFX1 gbuf_d_545(.A(n_5020), .Y(d_out_545));
CLKBUFX1 gbuf_q_545(.A(q_in_545), .Y(g3965));
CLKBUFX1 gbuf_d_546(.A(n_5034), .Y(d_out_546));
CLKBUFX1 gbuf_q_546(.A(q_in_546), .Y(g3917));
CLKBUFX1 gbuf_d_547(.A(n_5018), .Y(d_out_547));
CLKBUFX1 gbuf_q_547(.A(q_in_547), .Y(g2331));
CLKBUFX1 gbuf_d_548(.A(n_5017), .Y(d_out_548));
CLKBUFX1 gbuf_q_548(.A(q_in_548), .Y(g2361));
CLKBUFX1 gbuf_d_549(.A(n_5014), .Y(d_out_549));
CLKBUFX1 gbuf_q_549(.A(q_in_549), .Y(n_4339));
CLKBUFX1 gbuf_d_550(.A(n_5008), .Y(d_out_550));
CLKBUFX1 gbuf_qn_550(.A(qn_in_550), .Y(g5503));
CLKBUFX1 gbuf_d_551(.A(n_5006), .Y(d_out_551));
CLKBUFX1 gbuf_qn_551(.A(qn_in_551), .Y(g5849));
CLKBUFX1 gbuf_d_552(.A(n_5013), .Y(d_out_552));
CLKBUFX1 gbuf_q_552(.A(q_in_552), .Y(g3115));
CLKBUFX1 gbuf_d_553(.A(n_5005), .Y(d_out_553));
CLKBUFX1 gbuf_qn_553(.A(qn_in_553), .Y(g6195));
CLKBUFX1 gbuf_d_554(.A(n_5004), .Y(d_out_554));
CLKBUFX1 gbuf_qn_554(.A(qn_in_554), .Y(g3147));
CLKBUFX1 gbuf_d_555(.A(n_5002), .Y(d_out_555));
CLKBUFX1 gbuf_qn_555(.A(qn_in_555), .Y(g3498));
CLKBUFX1 gbuf_d_556(.A(n_5001), .Y(d_out_556));
CLKBUFX1 gbuf_qn_556(.A(qn_in_556), .Y(g3849));
CLKBUFX1 gbuf_d_557(.A(n_5012), .Y(d_out_557));
CLKBUFX1 gbuf_q_557(.A(q_in_557), .Y(g3466));
CLKBUFX1 gbuf_d_558(.A(n_5003), .Y(d_out_558));
CLKBUFX1 gbuf_qn_558(.A(qn_in_558), .Y(g6541));
CLKBUFX1 gbuf_d_559(.A(n_4970), .Y(d_out_559));
CLKBUFX1 gbuf_q_559(.A(q_in_559), .Y(g_20244));
OAI21X1 g64075(.A0 (g_13255), .A1 (g_16983), .B0 (n_3522), .Y(n_6280));
OR2X1 g64154(.A (n_5227), .B (n_10841), .Y (n_5562));
NOR2X1 g62585(.A (g5077), .B (n_9856), .Y (n_5518));
NAND2X1 g62618(.A (n_5364), .B (n_5363), .Y (n_5365));
NAND4X1 g64380(.A (n_10841), .B (n_5362), .C (g2735), .D (n_11012),.Y (n_5436));
NOR2X1 g62645(.A (g5069), .B (g5077), .Y (n_5361));
MX2X1 g62711(.A (g2084), .B (n_4905), .S0 (n_9000), .Y (n_5359));
OAI22X1 g62715(.A0 (n_4907), .A1 (n_9371), .B0 (g2241), .B1 (n_9992),.Y (n_5358));
OAI22X1 g62717(.A0 (n_4904), .A1 (n_9903), .B0 (g2265), .B1(n_10063), .Y (n_5357));
MX2X1 g62718(.A (g2269), .B (n_4899), .S0 (n_9279), .Y (n_5356));
MX2X1 g62722(.A (g2403), .B (n_4708), .S0 (n_9167), .Y (n_5355));
OAI22X1 g61333(.A0 (n_4780), .A1 (n_9976), .B0 (g1752), .B1 (n_9664),.Y (n_5354));
OAI22X1 g62725(.A0 (n_4716), .A1 (n_9431), .B0 (g2533), .B1 (n_9698),.Y (n_5353));
MX2X1 g62726(.A (g2537), .B (n_4707), .S0 (n_9218), .Y (n_5352));
OAI22X1 g62728(.A0 (n_4727), .A1 (n_9772), .B0 (g2643), .B1 (n_9651),.Y (n_5350));
OAI22X1 g61334(.A0 (n_4781), .A1 (n_10952), .B0 (g1736), .B1(n_9664), .Y (n_5349));
OAI22X1 g61335(.A0 (n_4779), .A1 (n_9461), .B0 (g1756), .B1 (n_9209),.Y (n_5348));
OAI22X1 g61336(.A0 (n_4777), .A1 (n_10952), .B0 (g1744), .B1(n_9992), .Y (n_5347));
AOI21X1 g64708(.A0 (n_4224), .A1 (n_8895), .B0 (n_4935), .Y (n_5346));
OAI22X1 g61337(.A0 (n_4776), .A1 (n_9129), .B0 (g1874), .B1(n_10005), .Y (n_5345));
MX2X1 g61338(.A (n_4187), .B (n_4775), .S0 (n_8955), .Y (n_5344));
OAI22X1 g61339(.A0 (n_4774), .A1 (n_9431), .B0 (g1870), .B1 (n_9521),.Y (n_5342));
OAI22X1 g61340(.A0 (n_4773), .A1 (n_9976), .B0 (g1886), .B1 (n_9651),.Y (n_5341));
OAI22X1 g61341(.A0 (n_4772), .A1 (n_9431), .B0 (g1890), .B1 (n_9811),.Y (n_5340));
NOR2X1 g62790(.A (n_4900), .B (n_9019), .Y (n_5339));
OAI22X1 g61342(.A0 (n_4770), .A1 (n_9772), .B0 (g1878), .B1 (n_9651),.Y (n_5338));
MX2X1 g61344(.A (n_4183), .B (n_4769), .S0 (n_9156), .Y (n_5337));
OAI22X1 g61345(.A0 (n_4768), .A1 (n_9976), .B0 (g2004), .B1 (n_9627),.Y (n_5336));
MX2X1 g61350(.A (n_4527), .B (n_4767), .S0 (n_9279), .Y (n_5335));
MX2X1 g62922(.A (g3329), .B (n_3020), .S0 (n_9553), .Y (n_5333));
MX2X1 g62924(.A (g3680), .B (n_3019), .S0 (n_8955), .Y (n_5331));
MX2X1 g62954(.A (g5216), .B (n_4670), .S0 (n_9750), .Y (n_5330));
MX2X1 g62958(.A (g5236), .B (n_4669), .S0 (n_9333), .Y (n_5329));
MX2X1 g62960(.A (g5244), .B (n_4656), .S0 (n_9000), .Y (n_5328));
MX2X1 g62961(.A (g5248), .B (n_4667), .S0 (n_8955), .Y (n_5327));
MX2X1 g62977(.A (g5563), .B (n_4666), .S0 (n_9256), .Y (n_5326));
MX2X1 g62981(.A (g5583), .B (n_4665), .S0 (n_9240), .Y (n_5325));
MX2X1 g63002(.A (g5909), .B (n_4662), .S0 (n_9834), .Y (n_5324));
NOR2X1 g61921(.A (n_5723), .B (n_6549), .Y (n_5323));
MX2X1 g63009(.A (g5941), .B (n_4661), .S0 (n_9797), .Y (n_5321));
OAI22X1 g63016(.A0 (n_4689), .A1 (n_10952), .B0 (g3125), .B1(n_9651), .Y (n_5319));
MX2X1 g63019(.A (g3129), .B (n_4651), .S0 (n_9358), .Y (n_5318));
MX2X1 g63028(.A (g6255), .B (n_4660), .S0 (n_8955), .Y (n_5317));
MX2X1 g63034(.A (g6283), .B (n_4659), .S0 (n_9894), .Y (n_5315));
MX2X1 g63035(.A (g6287), .B (n_4658), .S0 (n_10005), .Y (n_5313));
MX2X1 g63036(.A (g6291), .B (n_4657), .S0 (n_8955), .Y (n_5312));
NAND3X1 g61958(.A (n_4912), .B (g_22552), .C (n_10385), .Y (n_5311));
OAI22X1 g61960(.A0 (n_4963), .A1 (n_3916), .B0 (n_3310), .B1(n_9651), .Y (n_5310));
MX2X1 g63075(.A (g6621), .B (n_4653), .S0 (n_9797), .Y (n_5309));
MX2X1 g63077(.A (g6629), .B (n_4652), .S0 (n_9218), .Y (n_5308));
OAI22X1 g63085(.A0 (n_4688), .A1 (n_9976), .B0 (g3476), .B1 (n_9627),.Y (n_5307));
CLKBUFX1 gbuf_d_560(.A(n_4927), .Y(d_out_560));
CLKBUFX1 gbuf_q_560(.A(q_in_560), .Y(g1772));
MX2X1 g63086(.A (g3480), .B (n_4650), .S0 (n_9218), .Y (n_5306));
MX2X1 g63107(.A (g2047), .B (n_4649), .S0 (n_9834), .Y (n_5304));
MX2X1 g63108(.A (g2040), .B (n_4647), .S0 (n_8955), .Y (n_5302));
CLKBUFX1 gbuf_d_561(.A(n_4940), .Y(d_out_561));
CLKBUFX1 gbuf_q_561(.A(q_in_561), .Y(g_15381));
CLKBUFX1 gbuf_d_562(.A(n_4876), .Y(d_out_562));
CLKBUFX1 gbuf_q_562(.A(q_in_562), .Y(g_5450));
MX2X1 g63126(.A (g3929), .B (n_4655), .S0 (n_9256), .Y (n_5300));
MX2X1 g63128(.A (g3937), .B (n_4654), .S0 (n_9750), .Y (n_5299));
CLKBUFX1 gbuf_d_563(.A(n_4887), .Y(d_out_563));
CLKBUFX1 gbuf_q_563(.A(q_in_563), .Y(g4372));
MX2X1 g63143(.A (g1644), .B (n_4676), .S0 (n_9234), .Y (n_5297));
MX2X1 g63144(.A (g2606), .B (n_4645), .S0 (n_9167), .Y (n_5296));
MX2X1 g63145(.A (g1636), .B (n_4673), .S0 (n_10005), .Y (n_5294));
MX2X1 g63146(.A (g2599), .B (n_4640), .S0 (n_10005), .Y (n_5293));
NAND3X1 g60928(.A (n_4867), .B (n_2794), .C (n_4598), .Y (n_5291));
NOR2X1 g63203(.A (n_4898), .B (n_8588), .Y (n_5290));
NOR2X1 g63211(.A (n_4897), .B (n_10895), .Y (n_5289));
AOI21X1 g62050(.A0 (n_4590), .A1 (n_4251), .B0 (n_8707), .Y (n_5288));
INVX1 g63249(.A (n_6570), .Y (n_5287));
NAND4X1 g63316(.A (n_3219), .B (n_4605), .C (n_4098), .D (n_3895), .Y(n_5284));
AOI22X1 g60931(.A0 (n_4600), .A1 (n_9521), .B0 (n_10196), .B1(n_10952), .Y (n_5283));
MX2X1 g61177(.A (n_4529), .B (n_4603), .S0 (n_9894), .Y (n_5282));
MX2X1 g61184(.A (n_4531), .B (n_4597), .S0 (n_9234), .Y (n_5279));
MX2X1 g61190(.A (n_4726), .B (n_4594), .S0 (n_9172), .Y (n_5278));
NAND3X1 g62240(.A (n_4833), .B (n_2783), .C (n_4809), .Y (n_5276));
OAI22X1 g63645(.A0 (n_4049), .A1 (n_9193), .B0 (g4369), .B1 (n_9992),.Y (n_5275));
NAND2X1 g61212(.A (g4375), .B (n_9019), .Y (n_5273));
MX2X1 g62303(.A (g5046), .B (n_4813), .S0 (n_10063), .Y (n_5272));
MX2X1 g63757(.A (g_22371), .B (g14125), .S0 (n_5582), .Y (n_5271));
MX2X1 g62322(.A (n_11055), .B (n_4806), .S0 (n_9167), .Y (n_5270));
CLKBUFX1 gbuf_d_564(.A(n_4824), .Y(d_out_564));
CLKBUFX1 gbuf_q_564(.A(q_in_564), .Y(g11770));
AOI21X1 g61262(.A0 (n_4836), .A1 (n_1528), .B0 (n_4838), .Y (n_5268));
AOI21X1 g61264(.A0 (n_4834), .A1 (n_1529), .B0 (n_4835), .Y (n_5267));
AOI21X1 g61265(.A0 (n_4829), .A1 (n_2258), .B0 (n_4830), .Y (n_5266));
CLKBUFX1 gbuf_d_565(.A(n_4915), .Y(d_out_565));
CLKBUFX1 gbuf_q_565(.A(q_in_565), .Y(g_19113));
AOI21X1 g61267(.A0 (n_4827), .A1 (n_1519), .B0 (n_4828), .Y (n_5265));
CLKBUFX1 gbuf_d_566(.A(n_4929), .Y(d_out_566));
CLKBUFX1 gbuf_qn_566(.A(qn_in_566), .Y(g5481));
CLKBUFX1 gbuf_d_567(.A(n_4928), .Y(d_out_567));
CLKBUFX1 gbuf_q_567(.A(q_in_567), .Y(g5485));
CLKBUFX1 gbuf_d_568(.A(n_4926), .Y(d_out_568));
CLKBUFX1 gbuf_qn_568(.A(qn_in_568), .Y(g5827));
CLKBUFX1 gbuf_d_569(.A(n_4925), .Y(d_out_569));
CLKBUFX1 gbuf_q_569(.A(q_in_569), .Y(g5831));
CLKBUFX1 gbuf_d_570(.A(n_4924), .Y(d_out_570));
CLKBUFX1 gbuf_q_570(.A(q_in_570), .Y(n_4139));
CLKBUFX1 gbuf_d_571(.A(n_4922), .Y(d_out_571));
CLKBUFX1 gbuf_q_571(.A(q_in_571), .Y(g6177));
CLKBUFX1 gbuf_d_572(.A(n_4923), .Y(d_out_572));
CLKBUFX1 gbuf_qn_572(.A(qn_in_572), .Y(g6173));
CLKBUFX1 gbuf_d_573(.A(n_4918), .Y(d_out_573));
CLKBUFX1 gbuf_q_573(.A(q_in_573), .Y(g1906));
CLKBUFX1 gbuf_d_574(.A(n_4917), .Y(d_out_574));
CLKBUFX1 gbuf_q_574(.A(q_in_574), .Y(g1936));
CLKBUFX1 gbuf_d_575(.A(n_4877), .Y(d_out_575));
CLKBUFX1 gbuf_qn_575(.A(qn_in_575), .Y(g4112));
CLKBUFX1 gbuf_d_576(.A(n_4870), .Y(d_out_576));
CLKBUFX1 gbuf_qn_576(.A(qn_in_576), .Y(g4116));
CLKBUFX1 gbuf_d_577(.A(n_4869), .Y(d_out_577));
CLKBUFX1 gbuf_qn_577(.A(qn_in_577), .Y(g4119));
CLKBUFX1 gbuf_d_578(.A(n_4868), .Y(d_out_578));
CLKBUFX1 gbuf_qn_578(.A(qn_in_578), .Y(g4122));
CLKBUFX1 gbuf_d_579(.A(n_4891), .Y(d_out_579));
CLKBUFX1 gbuf_q_579(.A(q_in_579), .Y(g_3974));
CLKBUFX1 gbuf_d_580(.A(n_4841), .Y(d_out_580));
CLKBUFX1 gbuf_q_580(.A(q_in_580), .Y(n_1356));
OAI21X1 g64370(.A0 (n_4803), .A1 (n_10650), .B0 (n_4822), .Y(g33079));
OAI21X1 g64371(.A0 (n_4804), .A1 (n_10650), .B0 (n_4823), .Y(g33435));
CLKBUFX1 gbuf_d_581(.A(n_4934), .Y(d_out_581));
CLKBUFX1 gbuf_qn_581(.A(qn_in_581), .Y(g4531));
NAND3X1 g61064(.A (n_4787), .B (n_10372), .C (n_10949), .Y (n_5259));
XOR2X1 g61289(.A (n_1261), .B (n_4798), .Y (n_5258));
NAND3X1 g61069(.A (n_4920), .B (n_10669), .C (n_9894), .Y (n_10548));
INVX1 g62616(.A (n_5374), .Y (n_5454));
NAND2X1 g62636(.A (n_4931), .B (n_4572), .Y (n_5254));
NAND3X1 g61072(.A (n_4919), .B (n_10978), .C (n_9209), .Y (n_5253));
OAI22X1 g62689(.A0 (n_4725), .A1 (n_9371), .B0 (g2667), .B1 (n_9992),.Y (n_5252));
MX2X1 g62690(.A (g2671), .B (n_4712), .S0 (n_8955), .Y (n_5251));
OAI22X1 g62693(.A0 (n_4730), .A1 (n_10952), .B0 (g1706), .B1(n_9992), .Y (n_5249));
MX2X1 g62698(.A (g1710), .B (n_4715), .S0 (n_9279), .Y (n_5248));
OR2X1 g64528(.A (n_5362), .B (n_9398), .Y (n_5247));
MX2X1 g62703(.A (g1816), .B (n_10467), .S0 (n_9172), .Y (n_5246));
OAI22X1 g62705(.A0 (n_4723), .A1 (n_9976), .B0 (g1840), .B1 (n_9992),.Y (n_5245));
MX2X1 g62706(.A (g1844), .B (n_4711), .S0 (n_9240), .Y (n_5244));
MX2X1 g62707(.A (g1950), .B (n_4731), .S0 (n_9172), .Y (n_5242));
OAI22X1 g62709(.A0 (n_4721), .A1 (n_9193), .B0 (g1974), .B1 (n_9992),.Y (n_5241));
MX2X1 g62710(.A (g1978), .B (n_4710), .S0 (n_8955), .Y (n_5240));
OAI22X1 g62713(.A0 (n_4719), .A1 (n_10952), .B0 (g2108), .B1(n_9830), .Y (n_5239));
MX2X1 g62714(.A (g2112), .B (n_4709), .S0 (n_9750), .Y (n_5238));
MX2X1 g62716(.A (n_5961), .B (n_4713), .S0 (n_9501), .Y (n_5236));
OAI22X1 g61331(.A0 (n_4783), .A1 (n_10952), .B0 (g1740), .B1(n_9651), .Y (n_5235));
MX2X1 g61332(.A (n_4190), .B (n_4782), .S0 (n_8955), .Y (n_5233));
OAI22X1 g62721(.A0 (n_4717), .A1 (n_9599), .B0 (g2399), .B1 (n_9992),.Y (n_5232));
OAI22X1 g62723(.A0 (n_4532), .A1 (n_9772), .B0 (g2509), .B1 (n_9558),.Y (n_5231));
MX2X1 g62724(.A (n_5229), .B (n_4520), .S0 (n_9311), .Y (n_5230));
NAND2X1 g64655(.A (n_4936), .B (n_11012), .Y (n_5227));
CLKBUFX1 gbuf_d_582(.A(n_4587), .Y(d_out_582));
CLKBUFX1 gbuf_qn_582(.A(qn_in_582), .Y(g_6283));
MX2X1 g64698(.A (n_4556), .B (n_4232), .S0 (n_8895), .Y (n_5226));
CLKBUFX1 gbuf_d_583(.A(n_4746), .Y(d_out_583));
CLKBUFX1 gbuf_qn_583(.A(qn_in_583), .Y(g5077));
MX2X1 g64705(.A (n_4555), .B (n_4230), .S0 (n_8895), .Y (n_5225));
AOI21X1 g64706(.A0 (n_4225), .A1 (n_8895), .B0 (n_4812), .Y (n_5224));
AND2X1 g60974(.A (n_4639), .B (n_4690), .Y (n_5223));
AND2X1 g60975(.A (n_4634), .B (n_4680), .Y (n_5222));
AND2X1 g62821(.A (g4438), .B (n_10687), .Y (n_5364));
NAND2X1 g62822(.A (g4438), .B (n_9107), .Y (n_5221));
AND2X1 g60976(.A (n_4630), .B (n_4678), .Y (n_5219));
AND2X1 g60977(.A (n_4619), .B (n_4677), .Y (n_5218));
AOI21X1 g62921(.A0 (g5069), .A1 (g5084), .B0 (n_4753), .Y (n_5215));
CLKBUFX1 gbuf_d_584(.A(n_4589), .Y(d_out_584));
CLKBUFX1 gbuf_q_584(.A(q_in_584), .Y(g_22306));
CLKBUFX1 gbuf_d_585(.A(n_4789), .Y(d_out_585));
CLKBUFX1 gbuf_qn_585(.A(qn_in_585), .Y(g6181));
MX2X1 g62944(.A (g5188), .B (n_4442), .S0 (n_9469), .Y (n_5214));
MX2X1 g62945(.A (g5204), .B (n_4441), .S0 (n_8955), .Y (n_5213));
MX2X1 g62946(.A (g5256), .B (n_4440), .S0 (n_9000), .Y (n_5212));
MX2X1 g62947(.A (g5212), .B (n_4439), .S0 (n_9256), .Y (n_5210));
MX2X1 g62948(.A (g5260), .B (n_4347), .S0 (n_9311), .Y (n_5209));
MX2X1 g62949(.A (g5220), .B (n_4493), .S0 (n_9172), .Y (n_5207));
MX2X1 g62950(.A (g5264), .B (n_4438), .S0 (n_9000), .Y (n_5206));
MX2X1 g62951(.A (g5196), .B (n_4437), .S0 (n_8955), .Y (n_5205));
MX2X1 g62952(.A (g5200), .B (n_4458), .S0 (n_9091), .Y (n_5204));
MX2X1 g62953(.A (g5208), .B (n_4459), .S0 (n_9240), .Y (n_5202));
MX2X1 g62955(.A (g5224), .B (n_4381), .S0 (n_9000), .Y (n_5201));
MX2X1 g62956(.A (g5228), .B (n_4507), .S0 (n_9156), .Y (n_5200));
MX2X1 g62957(.A (g5232), .B (n_4504), .S0 (n_9167), .Y (n_5199));
MX2X1 g62959(.A (g5240), .B (n_4503), .S0 (n_9256), .Y (n_5197));
MX2X1 g62962(.A (g5252), .B (n_4400), .S0 (n_8955), .Y (n_5195));
MX2X1 g62963(.A (g5268), .B (n_4434), .S0 (n_9256), .Y (n_5193));
MX2X1 g62967(.A (g5535), .B (n_4433), .S0 (n_9091), .Y (n_5192));
MX2X1 g62968(.A (g5551), .B (n_4432), .S0 (n_9797), .Y (n_5190));
MX2X1 g62969(.A (g5603), .B (n_4431), .S0 (n_9359), .Y (n_5189));
MX2X1 g62970(.A (g5559), .B (n_4345), .S0 (n_10687), .Y (n_5187));
MX2X1 g62971(.A (g5607), .B (n_4430), .S0 (n_9172), .Y (n_5186));
MX2X1 g62972(.A (g5567), .B (n_4502), .S0 (n_9240), .Y (n_5185));
MX2X1 g62973(.A (g5611), .B (n_4429), .S0 (n_10005), .Y (n_5184));
MX2X1 g62974(.A (g5543), .B (n_4428), .S0 (n_9834), .Y (n_5183));
MX2X1 g62975(.A (g5547), .B (n_4501), .S0 (n_9311), .Y (n_5182));
MX2X1 g62976(.A (g5555), .B (n_4500), .S0 (n_9000), .Y (n_5181));
MX2X1 g62978(.A (g5571), .B (n_4427), .S0 (n_9992), .Y (n_5179));
MX2X1 g62979(.A (g5575), .B (n_4498), .S0 (n_9797), .Y (n_5177));
MX2X1 g62980(.A (g5579), .B (n_4496), .S0 (n_8955), .Y (n_5175));
MX2X1 g62982(.A (g5587), .B (n_4495), .S0 (n_8955), .Y (n_5174));
MX2X1 g62983(.A (g5591), .B (n_4426), .S0 (n_8955), .Y (n_5173));
MX2X1 g62984(.A (g5595), .B (n_4425), .S0 (n_9000), .Y (n_5172));
MX2X1 g62985(.A (g5599), .B (n_4423), .S0 (n_9992), .Y (n_5171));
MX2X1 g62986(.A (g5615), .B (n_4421), .S0 (n_8955), .Y (n_5170));
MX2X1 g62992(.A (g5881), .B (n_4420), .S0 (n_9466), .Y (n_5168));
MX2X1 g62993(.A (g5897), .B (n_4419), .S0 (n_9834), .Y (n_5167));
MX2X1 g62994(.A (g5949), .B (n_4418), .S0 (n_9156), .Y (n_5165));
MX2X1 g62995(.A (g5905), .B (n_4417), .S0 (n_9167), .Y (n_5164));
MX2X1 g62996(.A (g5953), .B (n_4416), .S0 (n_9156), .Y (n_5163));
MX2X1 g62997(.A (g5913), .B (n_4492), .S0 (n_9000), .Y (n_5161));
MX2X1 g62998(.A (g5957), .B (n_4415), .S0 (n_9359), .Y (n_5160));
MX2X1 g62999(.A (g5889), .B (n_4414), .S0 (n_9000), .Y (n_5159));
MX2X1 g63000(.A (g5893), .B (n_4490), .S0 (n_9992), .Y (n_5158));
MX2X1 g63001(.A (g5901), .B (n_4489), .S0 (n_9156), .Y (n_5156));
MX2X1 g63003(.A (g5917), .B (n_4413), .S0 (n_9311), .Y (n_5155));
MX2X1 g63004(.A (g5921), .B (n_4488), .S0 (n_9218), .Y (n_5154));
MX2X1 g63005(.A (g5925), .B (n_4487), .S0 (n_8955), .Y (n_5152));
MX2X1 g63006(.A (g5929), .B (n_4411), .S0 (n_9000), .Y (n_5151));
MX2X1 g63007(.A (g5933), .B (n_4486), .S0 (n_9359), .Y (n_5150));
MX2X1 g63008(.A (g5937), .B (n_4403), .S0 (n_9172), .Y (n_5149));
MX2X1 g63010(.A (g5945), .B (n_4410), .S0 (n_9797), .Y (n_5148));
MX2X1 g63011(.A (g5961), .B (n_4409), .S0 (n_9992), .Y (n_5146));
MX2X1 g63015(.A (g3119), .B (n_4485), .S0 (n_9664), .Y (n_5144));
MX2X1 g63017(.A (g6227), .B (n_4436), .S0 (n_9172), .Y (n_5143));
MX2X1 g63018(.A (g6243), .B (n_4360), .S0 (n_9358), .Y (n_5141));
MX2X1 g63020(.A (g6295), .B (n_4408), .S0 (n_9091), .Y (n_5139));
MX2X1 g63021(.A (g6251), .B (n_4407), .S0 (n_8955), .Y (n_5137));
MX2X1 g63022(.A (g6299), .B (n_4406), .S0 (n_9333), .Y (n_5136));
MX2X1 g63023(.A (g6259), .B (n_4483), .S0 (n_9000), .Y (n_5135));
MX2X1 g63024(.A (g6303), .B (n_4405), .S0 (n_9234), .Y (n_5134));
MX2X1 g63025(.A (g6235), .B (n_4404), .S0 (n_9311), .Y (n_5133));
MX2X1 g63026(.A (g6239), .B (n_4481), .S0 (n_9681), .Y (n_5131));
MX2X1 g63027(.A (g6247), .B (n_4479), .S0 (n_9681), .Y (n_5130));
MX2X1 g63029(.A (g6263), .B (n_4402), .S0 (n_9333), .Y (n_5129));
MX2X1 g63030(.A (g6267), .B (n_4478), .S0 (n_9240), .Y (n_5128));
MX2X1 g63031(.A (g6271), .B (n_4477), .S0 (n_9894), .Y (n_5127));
MX2X1 g63032(.A (g6275), .B (n_4401), .S0 (n_9797), .Y (n_5126));
MX2X1 g63033(.A (g6279), .B (n_4450), .S0 (n_9797), .Y (n_5125));
MX2X1 g63037(.A (g6307), .B (n_4399), .S0 (n_9311), .Y (n_5124));
MX2X1 g63038(.A (g3179), .B (n_4398), .S0 (n_9256), .Y (n_5123));
MX2X1 g63039(.A (g3195), .B (n_4397), .S0 (n_9234), .Y (n_5122));
MX2X1 g63040(.A (g3247), .B (n_4396), .S0 (n_9234), .Y (n_5121));
MX2X1 g63041(.A (g3203), .B (n_4395), .S0 (n_9156), .Y (n_5119));
MX2X1 g63042(.A (g3251), .B (n_4393), .S0 (n_9000), .Y (n_5118));
MX2X1 g63043(.A (g3211), .B (n_4475), .S0 (n_9000), .Y (n_5116));
MX2X1 g63044(.A (g3255), .B (n_4394), .S0 (n_9172), .Y (n_5115));
MX2X1 g63045(.A (g3187), .B (n_4392), .S0 (n_9172), .Y (n_5113));
MX2X1 g63048(.A (g3191), .B (n_4474), .S0 (n_10687), .Y (n_5112));
CLKBUFX1 gbuf_d_586(.A(n_4796), .Y(d_out_586));
CLKBUFX1 gbuf_qn_586(.A(qn_in_586), .Y(g5835));
MX2X1 g63050(.A (g3199), .B (n_4473), .S0 (n_9000), .Y (n_5111));
MX2X1 g63051(.A (g3207), .B (n_4391), .S0 (n_9000), .Y (n_5110));
MX2X1 g63052(.A (g3215), .B (n_4390), .S0 (n_9000), .Y (n_5109));
MX2X1 g63053(.A (g3219), .B (n_4472), .S0 (n_10005), .Y (n_5107));
MX2X1 g63054(.A (g6573), .B (n_4388), .S0 (n_9139), .Y (n_5106));
MX2X1 g63055(.A (g3223), .B (n_4471), .S0 (n_9311), .Y (n_5104));
MX2X1 g63056(.A (g6589), .B (n_4346), .S0 (n_9256), .Y (n_5103));
MX2X1 g63057(.A (g3227), .B (n_4387), .S0 (n_9091), .Y (n_5101));
MX2X1 g63058(.A (g6641), .B (n_4366), .S0 (n_9797), .Y (n_5100));
MX2X1 g63059(.A (g6597), .B (n_4389), .S0 (n_8955), .Y (n_5098));
MX2X1 g63060(.A (g3231), .B (n_4469), .S0 (n_9172), .Y (n_5097));
MX2X1 g63061(.A (g6645), .B (n_4363), .S0 (n_9359), .Y (n_5095));
MX2X1 g63062(.A (g6605), .B (n_4468), .S0 (n_9359), .Y (n_5094));
MX2X1 g63063(.A (g6649), .B (n_4349), .S0 (n_8955), .Y (n_5093));
MX2X1 g63064(.A (g6581), .B (n_4369), .S0 (n_8955), .Y (n_5092));
MX2X1 g63065(.A (g3235), .B (n_4380), .S0 (n_8955), .Y (n_5091));
MX2X1 g63066(.A (g6585), .B (n_4470), .S0 (n_8955), .Y (n_5090));
MX2X1 g63067(.A (g6593), .B (n_4446), .S0 (n_9172), .Y (n_5088));
MX2X1 g63068(.A (g3239), .B (n_4386), .S0 (n_9218), .Y (n_5087));
MX2X1 g63069(.A (g6601), .B (n_4412), .S0 (n_10005), .Y (n_5086));
MX2X1 g63070(.A (g3243), .B (n_4385), .S0 (n_9256), .Y (n_5085));
MX2X1 g63071(.A (g6609), .B (n_4344), .S0 (n_9000), .Y (n_5084));
MX2X1 g63072(.A (g6613), .B (n_4449), .S0 (n_9894), .Y (n_5083));
MX2X1 g63073(.A (g3259), .B (n_4348), .S0 (n_9234), .Y (n_5082));
MX2X1 g63074(.A (g6617), .B (n_4451), .S0 (n_9978), .Y (n_5081));
MX2X1 g63076(.A (g6625), .B (n_4467), .S0 (n_9218), .Y (n_5079));
MX2X1 g63078(.A (g6633), .B (n_4384), .S0 (n_8955), .Y (n_5077));
MX2X1 g63079(.A (g6637), .B (n_4383), .S0 (n_8955), .Y (n_5076));
MX2X1 g63080(.A (g6653), .B (n_4382), .S0 (n_9797), .Y (n_5075));
MX2X1 g63087(.A (g3530), .B (n_4379), .S0 (n_9466), .Y (n_5073));
MX2X1 g63088(.A (g3546), .B (n_4378), .S0 (n_8955), .Y (n_5072));
MX2X1 g63089(.A (g3598), .B (n_4377), .S0 (n_9311), .Y (n_5071));
MX2X1 g63090(.A (g3554), .B (n_4376), .S0 (n_9311), .Y (n_5069));
MX2X1 g61418(.A (g2004), .B (n_5057), .S0 (n_4306), .Y (n_5068));
MX2X1 g63091(.A (g3602), .B (n_4375), .S0 (n_9167), .Y (n_5067));
MX2X1 g63092(.A (g3562), .B (n_4466), .S0 (n_9750), .Y (n_5065));
MX2X1 g63093(.A (g3606), .B (n_4374), .S0 (n_9234), .Y (n_5064));
MX2X1 g63094(.A (g3538), .B (n_4373), .S0 (n_9750), .Y (n_5063));
MX2X1 g63095(.A (g3542), .B (n_4465), .S0 (n_9218), .Y (n_5062));
MX2X1 g63096(.A (g3550), .B (n_4464), .S0 (n_9359), .Y (n_5060));
MX2X1 g63097(.A (g3558), .B (n_4372), .S0 (n_9359), .Y (n_5059));
MX2X1 g61421(.A (g2016), .B (n_5057), .S0 (n_4305), .Y (n_5058));
MX2X1 g63098(.A (g3566), .B (n_4371), .S0 (n_8955), .Y (n_5056));
MX2X1 g63099(.A (g3570), .B (n_4462), .S0 (n_8955), .Y (n_5055));
MX2X1 g63100(.A (g3574), .B (n_4461), .S0 (n_9156), .Y (n_5053));
MX2X1 g63101(.A (g3578), .B (n_4370), .S0 (n_9156), .Y (n_5052));
MX2X1 g63102(.A (g3582), .B (n_4460), .S0 (n_9311), .Y (n_5051));
MX2X1 g63103(.A (g3586), .B (n_4368), .S0 (n_9172), .Y (n_5050));
MX2X1 g63104(.A (g3590), .B (n_4367), .S0 (n_9234), .Y (n_5048));
MX2X1 g63105(.A (g3594), .B (n_4365), .S0 (n_9311), .Y (n_5047));
MX2X1 g63106(.A (g3610), .B (n_4364), .S0 (n_9000), .Y (n_5046));
MX2X1 g61422(.A (g2020), .B (n_5057), .S0 (n_4319), .Y (n_5045));
MX2X1 g61423(.A (g2024), .B (n_5057), .S0 (n_4303), .Y (n_5044));
MX2X1 g63112(.A (g3881), .B (n_4362), .S0 (n_9553), .Y (n_5043));
MX2X1 g63113(.A (g3897), .B (n_4361), .S0 (n_9000), .Y (n_5042));
MX2X1 g63114(.A (g3949), .B (n_4359), .S0 (n_9750), .Y (n_5041));
MX2X1 g63115(.A (g3905), .B (n_4358), .S0 (n_9000), .Y (n_5040));
AOI21X1 g61424(.A0 (n_4742), .A1 (n_1532), .B0 (n_4744), .Y (n_5039));
MX2X1 g63116(.A (g3953), .B (n_4357), .S0 (n_9240), .Y (n_5038));
MX2X1 g63117(.A (g3913), .B (n_4457), .S0 (n_9553), .Y (n_5037));
MX2X1 g63118(.A (g3957), .B (n_4356), .S0 (n_10687), .Y (n_5035));
MX2X1 g63119(.A (g3889), .B (n_4355), .S0 (n_9311), .Y (n_5034));
MX2X1 g63120(.A (g3893), .B (n_4456), .S0 (n_9000), .Y (n_5033));
MX2X1 g63121(.A (g3901), .B (n_4455), .S0 (n_9000), .Y (n_5032));
AOI21X1 g61426(.A0 (n_4740), .A1 (n_1533), .B0 (n_4741), .Y (n_5030));
MX2X1 g63122(.A (g3909), .B (n_4354), .S0 (n_9000), .Y (n_5029));
MX2X1 g63123(.A (g3917), .B (n_4353), .S0 (n_9359), .Y (n_5028));
MX2X1 g63124(.A (g3921), .B (n_4454), .S0 (n_9000), .Y (n_5026));
MX2X1 g63125(.A (g3925), .B (n_4453), .S0 (n_9000), .Y (n_5025));
MX2X1 g63127(.A (g3933), .B (n_4452), .S0 (n_10005), .Y (n_5024));
MX2X1 g63129(.A (g3941), .B (n_4352), .S0 (n_9750), .Y (n_5023));
AOI21X1 g61428(.A0 (n_4738), .A1 (n_2521), .B0 (n_4739), .Y (n_5022));
MX2X1 g63130(.A (g3945), .B (n_4351), .S0 (n_9091), .Y (n_5021));
MX2X1 g63131(.A (g3961), .B (n_4350), .S0 (n_8955), .Y (n_5020));
AOI21X1 g61430(.A0 (n_4736), .A1 (n_1510), .B0 (n_4737), .Y (n_5019));
MX2X1 g63136(.A (g2338), .B (n_4336), .S0 (n_8955), .Y (n_5018));
MX2X1 g63137(.A (g2331), .B (n_4333), .S0 (n_9240), .Y (n_5017));
MX2X1 g63139(.A (g3470), .B (n_4448), .S0 (n_9091), .Y (n_5016));
MX2X1 g63140(.A (g2472), .B (n_4343), .S0 (n_9000), .Y (n_5015));
MX2X1 g63141(.A (g2465), .B (n_4340), .S0 (n_9000), .Y (n_5014));
NAND2X1 g63205(.A (n_4445), .B (n_4700), .Y (n_5013));
NAND2X1 g63215(.A (n_4444), .B (n_4695), .Y (n_5012));
NAND2X1 g62053(.A (n_3774), .B (n_4642), .Y (n_5009));
AOI22X1 g63248(.A0 (n_4330), .A1 (n_2943), .B0 (n_2944), .B1(n_5007), .Y (n_5008));
AOI22X1 g63252(.A0 (n_4328), .A1 (n_2940), .B0 (n_2941), .B1(n_5007), .Y (n_5006));
AOI22X1 g63254(.A0 (n_4325), .A1 (n_2936), .B0 (n_2937), .B1(n_5007), .Y (n_5005));
AOI22X1 g63256(.A0 (n_4317), .A1 (n_3253), .B0 (n_2933), .B1(n_5007), .Y (n_5004));
AOI22X1 g63258(.A0 (n_4323), .A1 (n_2930), .B0 (n_2931), .B1(n_5007), .Y (n_5003));
AOI22X1 g63263(.A0 (n_4321), .A1 (n_2928), .B0 (n_2929), .B1(n_5007), .Y (n_5002));
AOI22X1 g63264(.A0 (n_4315), .A1 (n_2923), .B0 (n_2924), .B1(n_5007), .Y (n_5001));
NAND4X1 g60930(.A (n_4593), .B (n_4866), .C (n_9750), .D (n_263), .Y(n_5000));
AOI21X1 g62082(.A0 (g_5450), .A1 (n_9856), .B0 (n_4672), .Y (n_4999));
NAND4X1 g63297(.A (n_6973), .B (n_10897), .C (g16722), .D (g3598), .Y(n_4996));
NAND3X1 g63325(.A (n_4693), .B (g_22379), .C (n_9351), .Y (n_4991));
CLKBUFX1 gbuf_d_587(.A(g16748), .Y(d_out_587));
CLKBUFX1 gbuf_q_587(.A(q_in_587), .Y(g4031));
NAND3X1 g63461(.A (n_4616), .B (n_2973), .C (g5156), .Y (n_4990));
NAND3X1 g63492(.A (n_868), .B (n_4293), .C (n_9874), .Y (n_4987));
AOI21X1 g60936(.A0 (n_4575), .A1 (n_2309), .B0 (n_9193), .Y (n_4986));
AOI22X1 g63553(.A0 (n_688), .A1 (n_4293), .B0 (n_4885), .B1 (g3831),.Y (n_4985));
NAND4X1 g63561(.A (n_6787), .B (g3933), .C (g13906), .D (n_5402), .Y(n_4984));
OAI21X1 g62213(.A0 (n_4567), .A1 (n_4982), .B0 (n_1283), .Y (n_4983));
OAI21X1 g62214(.A0 (n_4566), .A1 (n_4980), .B0 (n_1561), .Y (n_4981));
OAI21X1 g62215(.A0 (n_4565), .A1 (n_4978), .B0 (n_1282), .Y (n_4979));
OAI21X1 g62217(.A0 (n_4564), .A1 (n_11070), .B0 (n_1560), .Y(n_4977));
NAND4X1 g61553(.A (n_4581), .B (n_4843), .C (n_10013), .D (g4616), .Y(n_4976));
NAND2X1 g60939(.A (n_4586), .B (n_4243), .Y (n_4975));
NAND4X1 g62268(.A (n_4811), .B (n_4832), .C (n_9279), .D (n_287), .Y(n_4974));
OAI22X1 g61592(.A0 (n_4939), .A1 (n_4579), .B0 (n_79), .B1 (n_9862),.Y (n_4972));
XOR2X1 g63769(.A (n_2692), .B (n_4293), .Y (n_4971));
MX2X1 g63804(.A (g_21318), .B (n_4288), .S0 (n_9000), .Y (n_4970));
CLKBUFX1 gbuf_d_588(.A(g14125), .Y(d_out_588));
CLKBUFX1 gbuf_q_588(.A(q_in_588), .Y(g14147));
OR2X1 g61258(.A (n_4968), .B (g1682), .Y (n_4969));
CLKBUFX1 gbuf_d_589(.A(n_4684), .Y(d_out_589));
CLKBUFX1 gbuf_q_589(.A(q_in_589), .Y(g1367));
CLKBUFX1 gbuf_d_590(.A(n_4591), .Y(d_out_590));
CLKBUFX1 gbuf_q_590(.A(q_in_590), .Y(g1542));
CLKBUFX1 gbuf_d_591(.A(n_4821), .Y(d_out_591));
CLKBUFX1 gbuf_q_591(.A(q_in_591), .Y(g1312));
CLKBUFX1 gbuf_d_592(.A(n_4794), .Y(d_out_592));
CLKBUFX1 gbuf_q_592(.A(q_in_592), .Y(g10500));
CLKBUFX1 gbuf_d_593(.A(n_4626), .Y(d_out_593));
CLKBUFX1 gbuf_q_593(.A(q_in_593), .Y(g4950));
CLKBUFX1 gbuf_d_594(.A(n_4627), .Y(d_out_594));
CLKBUFX1 gbuf_q_594(.A(q_in_594), .Y(g4939));
CLKBUFX1 gbuf_d_595(.A(n_4785), .Y(d_out_595));
CLKBUFX1 gbuf_qn_595(.A(qn_in_595), .Y(g6527));
CLKBUFX1 gbuf_d_596(.A(n_4706), .Y(d_out_596));
CLKBUFX1 gbuf_q_596(.A(q_in_596), .Y(g4593));
CLKBUFX1 gbuf_d_597(.A(n_4714), .Y(d_out_597));
CLKBUFX1 gbuf_q_597(.A(q_in_597), .Y(g4332));
CLKBUFX1 gbuf_d_598(.A(n_4663), .Y(d_out_598));
CLKBUFX1 gbuf_q_598(.A(q_in_598), .Y(g_10715));
CLKBUFX1 gbuf_d_599(.A(n_4585), .Y(d_out_599));
CLKBUFX1 gbuf_q_599(.A(q_in_599), .Y(g4049));
AOI21X1 g61266(.A0 (n_4583), .A1 (n_919), .B0 (n_4584), .Y (n_4967));
CLKBUFX1 gbuf_d_600(.A(n_4800), .Y(d_out_600));
CLKBUFX1 gbuf_qn_600(.A(qn_in_600), .Y(g5134));
CLKBUFX1 gbuf_d_601(.A(n_4799), .Y(d_out_601));
CLKBUFX1 gbuf_q_601(.A(q_in_601), .Y(g5138));
CLKBUFX1 gbuf_d_602(.A(n_4797), .Y(d_out_602));
CLKBUFX1 gbuf_qn_602(.A(qn_in_602), .Y(g5489));
CLKBUFX1 gbuf_d_603(.A(n_4786), .Y(d_out_603));
CLKBUFX1 gbuf_q_603(.A(q_in_603), .Y(g6523));
CLKBUFX1 gbuf_d_604(.A(n_4734), .Y(d_out_604));
CLKBUFX1 gbuf_q_604(.A(q_in_604), .Y(g3639));
CLKBUFX1 gbuf_d_605(.A(n_4732), .Y(d_out_605));
CLKBUFX1 gbuf_q_605(.A(q_in_605), .Y(g3990));
CLKBUFX1 gbuf_d_606(.A(n_4752), .Y(d_out_606));
CLKBUFX1 gbuf_q_606(.A(q_in_606), .Y(g5471));
CLKBUFX1 gbuf_d_607(.A(n_4751), .Y(d_out_607));
CLKBUFX1 gbuf_q_607(.A(q_in_607), .Y(g5817));
CLKBUFX1 gbuf_d_608(.A(n_4750), .Y(d_out_608));
CLKBUFX1 gbuf_q_608(.A(q_in_608), .Y(g6163));
CLKBUFX1 gbuf_d_609(.A(n_4735), .Y(d_out_609));
CLKBUFX1 gbuf_q_609(.A(q_in_609), .Y(g3288));
CLKBUFX1 gbuf_d_610(.A(n_4705), .Y(d_out_610));
CLKBUFX1 gbuf_q_610(.A(q_in_610), .Y(n_7004));
CLKBUFX1 gbuf_d_611(.A(n_4704), .Y(d_out_611));
CLKBUFX1 gbuf_q_611(.A(q_in_611), .Y(n_6979));
CLKBUFX1 gbuf_d_612(.A(n_4747), .Y(d_out_612));
CLKBUFX1 gbuf_q_612(.A(q_in_612), .Y(g5046));
CLKBUFX1 gbuf_d_613(.A(n_4636), .Y(d_out_613));
CLKBUFX1 gbuf_q_613(.A(q_in_613), .Y(g_21318));
CLKBUFX1 gbuf_d_614(.A(n_4624), .Y(d_out_614));
CLKBUFX1 gbuf_q_614(.A(q_in_614), .Y(g3050));
CLKBUFX1 gbuf_d_615(.A(n_4623), .Y(d_out_615));
CLKBUFX1 gbuf_q_615(.A(q_in_615), .Y(g6098));
CLKBUFX1 gbuf_d_616(.A(n_4622), .Y(d_out_616));
CLKBUFX1 gbuf_q_616(.A(q_in_616), .Y(g6444));
CLKBUFX1 gbuf_d_617(.A(n_4620), .Y(d_out_617));
CLKBUFX1 gbuf_q_617(.A(q_in_617), .Y(g3401));
CLKBUFX1 gbuf_d_618(.A(n_4621), .Y(d_out_618));
CLKBUFX1 gbuf_q_618(.A(q_in_618), .Y(g3752));
CLKBUFX1 gbuf_d_619(.A(n_4625), .Y(d_out_619));
CLKBUFX1 gbuf_q_619(.A(q_in_619), .Y(g5752));
AOI21X1 g62254(.A0 (n_4262), .A1 (n_1972), .B0 (g4369), .Y (g34839));
AND2X1 g61063(.A (n_4766), .B (n_4795), .Y (n_4966));
XOR2X1 g61287(.A (n_1260), .B (n_4559), .Y (n_4965));
OR2X1 g62584(.A (n_4963), .B (n_3654), .Y (n_4964));
XOR2X1 g61290(.A (n_1257), .B (n_4562), .Y (n_4962));
NAND4X1 g62600(.A (n_4815), .B (g_4449), .C (n_10013), .D (n_3914),.Y (n_4961));
AND2X1 g61067(.A (n_4763), .B (n_4792), .Y (n_4960));
AND2X1 g61068(.A (n_4759), .B (n_4790), .Y (n_4959));
OR4X1 g62617(.A (g4438), .B (g4452), .C (g4443), .D (n_334), .Y(n_5374));
OAI22X1 g61744(.A0 (n_4519), .A1 (n_4956), .B0 (n_512), .B1 (n_9992),.Y (n_4957));
OR4X1 g62628(.A (n_2756), .B (n_11189), .C (n_11188), .D (n_4205), .Y(n_5457));
XOR2X1 g61745(.A (g4608), .B (n_4554), .Y (n_4955));
AND2X1 g61070(.A (n_4756), .B (n_4788), .Y (n_4954));
NAND3X1 g61071(.A (n_4784), .B (n_10853), .C (n_9834), .Y (n_4953));
MX2X1 g62687(.A (n_4893), .B (n_4528), .S0 (n_9000), .Y (n_4952));
MX2X1 g62688(.A (n_5958), .B (n_4526), .S0 (n_9333), .Y (n_4951));
MX2X1 g62692(.A (n_5964), .B (n_4525), .S0 (n_9172), .Y (n_4950));
MX2X1 g62704(.A (n_4948), .B (n_4524), .S0 (n_9172), .Y (n_4949));
MX2X1 g62708(.A (n_4946), .B (n_4523), .S0 (n_9156), .Y (n_4947));
MX2X1 g62712(.A (n_5953), .B (n_4522), .S0 (n_9218), .Y (n_4945));
OAI22X1 g62719(.A0 (n_4530), .A1 (n_9976), .B0 (g2375), .B1 (n_9862),.Y (n_4944));
MX2X1 g62720(.A (n_4942), .B (n_4521), .S0 (n_9553), .Y (n_4943));
OAI22X1 g61841(.A0 (n_4939), .A1 (n_4155), .B0 (n_126), .B1 (n_9651),.Y (n_4940));
CLKBUFX1 gbuf_d_620(.A(g11678), .Y(d_out_620));
CLKBUFX1 gbuf_q_620(.A(q_in_620), .Y(g_15127));
INVX1 g64835(.A (n_4936), .Y (n_5362));
AOI21X1 g64852(.A0 (n_4223), .A1 (n_4032), .B0 (n_8895), .Y (n_4935));
NAND2X1 g62846(.A (n_4546), .B (n_3214), .Y (n_4934));
AOI21X1 g62932(.A0 (g5052), .A1 (n_10078), .B0 (n_4545), .Y (n_4931));
AOI21X1 g61275(.A0 (n_4273), .A1 (n_1713), .B0 (n_4274), .Y (n_4930));
MX2X1 g62964(.A (g5475), .B (n_4163), .S0 (n_9311), .Y (n_4929));
OAI22X1 g62965(.A0 (n_10346), .A1 (n_9599), .B0 (g5481), .B1(n_9992), .Y (n_4928));
MX2X1 g62987(.A (g1779), .B (n_4142), .S0 (n_9000), .Y (n_4927));
MX2X1 g62988(.A (g5821), .B (n_4161), .S0 (n_9091), .Y (n_4926));
OAI22X1 g62989(.A0 (n_4165), .A1 (n_9371), .B0 (g5827), .B1 (n_9698),.Y (n_4925));
MX2X1 g62991(.A (g1772), .B (n_4140), .S0 (n_9311), .Y (n_4924));
MX2X1 g63012(.A (g6167), .B (n_4160), .S0 (n_9664), .Y (n_4923));
OAI22X1 g63013(.A0 (n_10448), .A1 (n_9599), .B0 (g6173), .B1(n_9992), .Y (n_4922));
NAND4X1 g61941(.A (n_3913), .B (n_11079), .C (n_9139), .D (n_284), .Y(n_4921));
XOR2X1 g61139(.A (n_963), .B (n_4150), .Y (n_4920));
XOR2X1 g61141(.A (n_942), .B (n_4151), .Y (n_4919));
MX2X1 g63081(.A (g1913), .B (n_4147), .S0 (n_9992), .Y (n_4918));
MX2X1 g63082(.A (g1906), .B (n_4145), .S0 (n_9834), .Y (n_4917));
MX2X1 g61982(.A (n_640), .B (n_4152), .S0 (n_9167), .Y (n_4915));
AOI21X1 g61429(.A0 (n_4539), .A1 (n_928), .B0 (n_4540), .Y (n_4913));
NAND2X1 g62019(.A (n_4422), .B (g_16404), .Y (n_4912));
NAND4X1 g62023(.A (n_4576), .B (n_4671), .C (n_9209), .D (g_19659),.Y (n_4911));
AOI22X1 g63265(.A0 (n_917), .A1 (n_10378), .B0 (n_10099), .B1(n_4906), .Y (n_4907));
OAI21X1 g63299(.A0 (n_702), .A1 (n_6752), .B0 (n_4184), .Y (n_4905));
AOI21X1 g63300(.A0 (n_10099), .A1 (g2269), .B0 (n_4514), .Y (n_4904));
AOI22X1 g63323(.A0 (n_783), .A1 (n_4108), .B0 (n_4121), .B1 (g1592),.Y (n_4900));
OAI21X1 g63328(.A0 (n_10097), .A1 (n_6025), .B0 (n_4513), .Y(n_4899));
INVX1 g63399(.A (g3329), .Y (n_4898));
INVX1 g63403(.A (g3680), .Y (n_4897));
CLKBUFX1 gbuf_d_621(.A(n_4553), .Y(d_out_621));
CLKBUFX1 gbuf_q_621(.A(q_in_621), .Y(g_16475));
AND2X1 g63431(.A (n_4615), .B (g5156), .Y (n_4896));
AOI21X1 g63525(.A0 (g13966), .A1 (n_491), .B0 (n_4302), .Y (n_4891));
NAND3X1 g63530(.A (n_4313), .B (g_21806), .C (n_9398), .Y (n_4889));
NAND3X1 g60938(.A (n_4592), .B (g1379), .C (n_9894), .Y (n_4888));
CLKBUFX1 gbuf_d_622(.A(n_4547), .Y(d_out_622));
CLKBUFX1 gbuf_q_622(.A(q_in_622), .Y(g6509));
OR2X1 g62239(.A (n_4286), .B (n_4068), .Y (n_4887));
MX2X1 g63616(.A (g3821), .B (n_85), .S0 (n_4885), .Y (n_4886));
MX2X1 g63624(.A (g2197), .B (g2153), .S0 (n_10378), .Y (n_4884));
MX2X1 g63625(.A (g2227), .B (g2197), .S0 (n_10378), .Y (n_4881));
AOI22X1 g63641(.A0 (n_3596), .A1 (n_9461), .B0 (n_4885), .B1(n_4878), .Y (n_4879));
OAI22X1 g63642(.A0 (n_4087), .A1 (n_9772), .B0 (n_3896), .B1(n_9992), .Y (n_4877));
CLKBUFX1 gbuf_d_623(.A(n_4512), .Y(d_out_623));
CLKBUFX1 gbuf_q_623(.A(q_in_623), .Y(g_4050));
OAI22X1 g62291(.A0 (n_2567), .A1 (n_5723), .B0 (n_21), .B1 (n_9862),.Y (n_4876));
NAND4X1 g61590(.A (g_15380), .B (n_9992), .C (n_1124), .D (n_4578),.Y (n_4875));
XOR2X1 g62302(.A (g4045), .B (g3990), .Y (n_4874));
OAI22X1 g63794(.A0 (n_4086), .A1 (n_9431), .B0 (g4112), .B1 (n_9521),.Y (n_4870));
OAI22X1 g63795(.A0 (n_4085), .A1 (n_9269), .B0 (g4116), .B1(n_10005), .Y (n_4869));
OAI22X1 g63796(.A0 (n_4084), .A1 (n_9599), .B0 (g4119), .B1 (n_9862),.Y (n_4868));
CLKBUFX1 gbuf_d_624(.A(n_4577), .Y(d_out_624));
CLKBUFX1 gbuf_q_624(.A(q_in_624), .Y(g_16958));
NAND4X1 g60945(.A (n_4569), .B (n_4866), .C (n_9359), .D (n_406), .Y(n_4867));
CLKBUFX1 gbuf_d_625(.A(n_4283), .Y(d_out_625));
CLKBUFX1 gbuf_q_625(.A(q_in_625), .Y(g4375));
CLKBUFX1 gbuf_d_626(.A(n_4298), .Y(d_out_626));
CLKBUFX1 gbuf_q_626(.A(q_in_626), .Y(g1361));
CLKBUFX1 gbuf_d_627(.A(n_4573), .Y(d_out_627));
CLKBUFX1 gbuf_q_627(.A(q_in_627), .Y(g1351));
OAI21X1 g61263(.A0 (n_10761), .A1 (n_10097), .B0 (n_4515), .Y(n_4865));
NAND3X1 g64008(.A (n_10373), .B (n_916), .C (n_9894), .Y (n_4864));
CLKBUFX1 gbuf_d_628(.A(n_4557), .Y(d_out_628));
CLKBUFX1 gbuf_qn_628(.A(qn_in_628), .Y(g6519));
CLKBUFX1 gbuf_d_629(.A(n_4533), .Y(d_out_629));
CLKBUFX1 gbuf_q_629(.A(q_in_629), .Y(n_11071));
CLKBUFX1 gbuf_d_630(.A(n_4561), .Y(d_out_630));
CLKBUFX1 gbuf_qn_630(.A(qn_in_630), .Y(g5142));
CLKBUFX1 gbuf_d_631(.A(n_4506), .Y(d_out_631));
CLKBUFX1 gbuf_qn_631(.A(qn_in_631), .Y(g_22639));
CLKBUFX1 gbuf_d_632(.A(n_4290), .Y(d_out_632));
CLKBUFX1 gbuf_q_632(.A(q_in_632), .Y(g1171));
CLKBUFX1 gbuf_d_633(.A(n_4574), .Y(d_out_633));
CLKBUFX1 gbuf_q_633(.A(q_in_633), .Y(g2941));
AOI21X1 g61269(.A0 (n_4281), .A1 (n_1702), .B0 (n_4282), .Y (n_4861));
CLKBUFX1 gbuf_d_634(.A(n_4563), .Y(d_out_634));
CLKBUFX1 gbuf_q_634(.A(q_in_634), .Y(g5041));
CLKBUFX1 gbuf_d_635(.A(n_4538), .Y(d_out_635));
CLKBUFX1 gbuf_q_635(.A(q_in_635), .Y(g5297));
CLKBUFX1 gbuf_d_636(.A(n_4537), .Y(d_out_636));
CLKBUFX1 gbuf_q_636(.A(q_in_636), .Y(g5644));
CLKBUFX1 gbuf_d_637(.A(n_4534), .Y(d_out_637));
CLKBUFX1 gbuf_q_637(.A(q_in_637), .Y(g6336));
CLKBUFX1 gbuf_d_638(.A(n_4535), .Y(d_out_638));
CLKBUFX1 gbuf_q_638(.A(q_in_638), .Y(g5990));
CLKBUFX1 gbuf_d_639(.A(n_4550), .Y(d_out_639));
CLKBUFX1 gbuf_q_639(.A(q_in_639), .Y(g5124));
AOI21X1 g61271(.A0 (n_4279), .A1 (n_1703), .B0 (n_4280), .Y (n_4860));
CLKBUFX1 gbuf_d_640(.A(n_4518), .Y(d_out_640));
CLKBUFX1 gbuf_q_640(.A(q_in_640), .Y(g4054));
CLKBUFX1 gbuf_d_641(.A(n_4338), .Y(d_out_641));
CLKBUFX1 gbuf_q_641(.A(q_in_641), .Y(n_1285));
CLKBUFX1 gbuf_d_642(.A(n_4510), .Y(d_out_642));
CLKBUFX1 gbuf_q_642(.A(q_in_642), .Y(g_9298));
CLKBUFX1 gbuf_d_643(.A(n_4508), .Y(d_out_643));
CLKBUFX1 gbuf_q_643(.A(q_in_643), .Y(g2886));
CLKBUFX1 gbuf_d_644(.A(n_4331), .Y(d_out_644));
CLKBUFX1 gbuf_q_644(.A(q_in_644), .Y(g5406));
CLKBUFX1 gbuf_d_645(.A(n_4297), .Y(d_out_645));
CLKBUFX1 gbuf_q_645(.A(q_in_645), .Y(n_6967));
AOI21X1 g61272(.A0 (n_4277), .A1 (n_2293), .B0 (n_4278), .Y (n_4859));
MX2X1 g61273(.A (g2311), .B (n_8761), .S0 (n_4125), .Y (n_4858));
MX2X1 g64090(.A (g_22600), .B (g14096), .S0 (n_5582), .Y (n_4857));
AOI21X1 g61274(.A0 (n_4275), .A1 (n_1677), .B0 (n_4276), .Y (n_4856));
AOI21X1 g64083(.A0 (g2902), .A1 (g2907), .B0 (n_4291), .Y (g32185));
AOI21X1 g61277(.A0 (n_4271), .A1 (n_1714), .B0 (n_4272), .Y (n_4854));
AOI21X1 g61278(.A0 (n_4269), .A1 (n_2780), .B0 (n_4270), .Y (n_4853));
MX2X1 g61279(.A (g2445), .B (n_8763), .S0 (n_4123), .Y (n_4852));
AOI21X1 g61280(.A0 (n_4267), .A1 (n_1671), .B0 (n_4268), .Y (n_4851));
MX2X1 g61281(.A (g2563), .B (n_11190), .S0 (n_4117), .Y (n_4850));
MX2X1 g61283(.A (g2571), .B (n_11190), .S0 (n_6746), .Y (n_4849));
MX2X1 g61284(.A (g2575), .B (n_11190), .S0 (n_4113), .Y (n_4847));
MX2X1 g61285(.A (g2579), .B (n_11191), .S0 (n_4119), .Y (n_4846));
MX2X1 g61286(.A (g2583), .B (n_11191), .S0 (n_4111), .Y (n_4845));
NAND3X1 g61729(.A (n_2582), .B (n_4843), .C (n_8757), .Y (n_4844));
CLKBUFX1 gbuf_d_646(.A(n_4570), .Y(d_out_646));
CLKBUFX1 gbuf_q_646(.A(q_in_646), .Y(g4584));
NAND3X1 g62601(.A (n_4810), .B (g_12465), .C (n_9698), .Y (n_4842));
NAND3X1 g64355(.A (n_4080), .B (n_4255), .C (n_2590), .Y (n_4841));
NOR2X1 g62622(.A (n_4839), .B (n_8879), .Y (n_4840));
NOR2X1 g61310(.A (n_10761), .B (n_4836), .Y (n_4838));
NOR2X1 g61311(.A (n_10761), .B (n_4834), .Y (n_4835));
NAND4X1 g62670(.A (n_4542), .B (n_4832), .C (n_9359), .D (n_251), .Y(n_4833));
NOR2X1 g61312(.A (n_10761), .B (n_4829), .Y (n_4830));
NOR2X1 g61314(.A (n_10761), .B (n_4827), .Y (n_4828));
MX2X1 g64453(.A (n_10867), .B (n_4248), .S0 (n_9359), .Y (n_4824));
CLKBUFX1 gbuf_d_647(.A(n_4560), .Y(d_out_647));
CLKBUFX1 gbuf_qn_647(.A(qn_in_647), .Y(g_16983));
OAI21X1 g64505(.A0 (n_4235), .A1 (n_4042), .B0 (n_10650), .Y(n_4823));
OAI21X1 g64506(.A0 (n_4239), .A1 (n_4043), .B0 (n_10650), .Y(n_4822));
NOR2X1 g60972(.A (n_4180), .B (n_9976), .Y (n_4821));
NAND4X1 g61826(.A (n_1787), .B (n_4045), .C (n_9874), .D (g_14342),.Y (n_4820));
NAND2X1 g62789(.A (n_11079), .B (n_9521), .Y (n_4963));
AND2X1 g62808(.A (n_11079), .B (n_3915), .Y (n_4815));
NAND3X1 g62834(.A (n_10696), .B (n_2985), .C (n_3985), .Y (n_4813));
INVX1 g64836(.A (g2748), .Y (n_4936));
AOI21X1 g64851(.A0 (n_3863), .A1 (n_4035), .B0 (n_8895), .Y (n_4812));
INVX1 g62839(.A (n_4810), .Y (n_4811));
NAND3X1 g62851(.A (n_4541), .B (g_20159), .C (n_9894), .Y (n_4809));
MX2X1 g62910(.A (n_4805), .B (g_17426), .S0 (n_3177), .Y (n_4806));
AOI21X1 g64979(.A0 (n_326), .A1 (n_3868), .B0 (n_4237), .Y (n_4804));
AOI21X1 g64980(.A0 (n_317), .A1 (n_3868), .B0 (n_4238), .Y (n_4803));
MX2X1 g62941(.A (g5128), .B (n_3983), .S0 (n_9091), .Y (n_4800));
OAI22X1 g62942(.A0 (n_3993), .A1 (n_9772), .B0 (g5134), .B1 (n_9501),.Y (n_4799));
AOI21X1 g61377(.A0 (n_10988), .A1 (g1246), .B0 (n_10989), .Y(n_4798));
MX2X1 g62966(.A (g5485), .B (n_3974), .S0 (n_9172), .Y (n_4797));
CLKBUFX1 gbuf_d_648(.A(n_4198), .Y(d_out_648));
CLKBUFX1 gbuf_q_648(.A(q_in_648), .Y(n_10657));
MX2X1 g62990(.A (g5831), .B (n_3973), .S0 (n_8955), .Y (n_4796));
NAND4X1 g61133(.A (n_4765), .B (n_4764), .C (n_4791), .D (n_2529), .Y(n_4795));
MX2X1 g61385(.A (g1246), .B (n_515), .S0 (n_9311), .Y (n_4794));
NAND4X1 g61134(.A (n_4762), .B (n_4761), .C (n_4791), .D (n_2556), .Y(n_4792));
CLKBUFX1 gbuf_d_649(.A(n_4200), .Y(d_out_649));
CLKBUFX1 gbuf_q_649(.A(q_in_649), .Y(g5033));
NAND4X1 g61135(.A (n_4758), .B (n_4757), .C (n_4791), .D (n_2280), .Y(n_4790));
MX2X1 g63014(.A (g6177), .B (n_3972), .S0 (n_9000), .Y (n_4789));
NAND4X1 g61136(.A (n_4755), .B (n_4791), .C (n_2244), .D (n_4754), .Y(n_4788));
XOR2X1 g61138(.A (n_952), .B (n_3977), .Y (n_4787));
OAI22X1 g63047(.A0 (n_3992), .A1 (n_9772), .B0 (g6519), .B1 (n_9664),.Y (n_4786));
MX2X1 g63049(.A (g6523), .B (n_3971), .S0 (n_10005), .Y (n_4785));
XOR2X1 g61140(.A (n_967), .B (n_3978), .Y (n_4784));
AOI21X1 g61406(.A0 (n_4220), .A1 (n_1710), .B0 (n_4221), .Y (n_4783));
OAI21X1 g61407(.A0 (n_6953), .A1 (n_7025), .B0 (n_4174), .Y (n_4782));
AOI21X1 g61408(.A0 (n_4218), .A1 (n_1711), .B0 (n_4219), .Y (n_4781));
AOI21X1 g61409(.A0 (n_4216), .A1 (n_2550), .B0 (n_4217), .Y (n_4780));
MX2X1 g61410(.A (g1752), .B (n_6953), .S0 (n_3949), .Y (n_4779));
AOI21X1 g61411(.A0 (n_4214), .A1 (n_1666), .B0 (n_4215), .Y (n_4777));
AOI21X1 g61412(.A0 (n_4211), .A1 (n_1705), .B0 (n_4212), .Y (n_4776));
OAI21X1 g61413(.A0 (n_11039), .A1 (n_10920), .B0 (n_4181), .Y(n_4775));
AOI21X1 g61414(.A0 (n_4209), .A1 (n_1706), .B0 (n_4210), .Y (n_4774));
AOI21X1 g61415(.A0 (n_4207), .A1 (n_2306), .B0 (n_4208), .Y (n_4773));
MX2X1 g61416(.A (g1886), .B (n_11039), .S0 (n_3946), .Y (n_4772));
AOI21X1 g61417(.A0 (n_4203), .A1 (n_1688), .B0 (n_4204), .Y (n_4770));
OAI21X1 g61419(.A0 (n_5057), .A1 (n_7102), .B0 (n_4185), .Y (n_4769));
MX2X1 g61420(.A (g2012), .B (n_5057), .S0 (n_3944), .Y (n_4768));
OAI21X1 g61425(.A0 (n_4743), .A1 (n_10899), .B0 (n_4167), .Y(n_4767));
NAND3X1 g61157(.A (n_4765), .B (n_4764), .C (n_4760), .Y (n_4766));
NAND3X1 g61158(.A (n_4762), .B (n_4761), .C (n_4760), .Y (n_4763));
CLKBUFX1 gbuf_d_650(.A(n_4171), .Y(d_out_650));
CLKBUFX1 gbuf_q_650(.A(q_in_650), .Y(g4438));
NAND3X1 g61159(.A (n_4758), .B (n_4757), .C (n_4760), .Y (n_4759));
NAND3X1 g61160(.A (n_4755), .B (n_4760), .C (n_4754), .Y (n_4756));
NOR2X1 g63197(.A (g5073), .B (g5084), .Y (n_4753));
CLKBUFX1 gbuf_d_651(.A(n_4257), .Y(d_out_651));
CLKBUFX1 gbuf_q_651(.A(q_in_651), .Y(g1199));
NAND2X1 g63200(.A (n_4159), .B (n_4005), .Y (n_4752));
NAND2X1 g63202(.A (n_4157), .B (n_4002), .Y (n_4751));
NAND2X1 g63204(.A (n_4156), .B (n_4000), .Y (n_4750));
NAND2X1 g63244(.A (n_4154), .B (n_3816), .Y (n_4747));
AOI21X1 g63246(.A0 (n_3411), .A1 (n_10005), .B0 (g5073), .Y (n_4746));
NOR2X1 g61469(.A (n_4743), .B (n_4742), .Y (n_4744));
NOR2X1 g61470(.A (n_4743), .B (n_4740), .Y (n_4741));
NOR2X1 g61472(.A (n_4743), .B (n_4738), .Y (n_4739));
NOR2X1 g61474(.A (n_4743), .B (n_4736), .Y (n_4737));
OAI21X1 g63276(.A0 (n_3776), .A1 (n_9193), .B0 (n_4102), .Y (n_4735));
OAI21X1 g63278(.A0 (n_3780), .A1 (n_9193), .B0 (n_4105), .Y (n_4734));
OAI21X1 g63279(.A0 (n_3777), .A1 (n_9107), .B0 (n_4103), .Y (n_4732));
OAI21X1 g63281(.A0 (n_914), .A1 (n_6685), .B0 (n_4188), .Y (n_4731));
AOI21X1 g63286(.A0 (n_10901), .A1 (g1710), .B0 (n_4173), .Y (n_4730));
AOI22X1 g63303(.A0 (n_903), .A1 (n_10978), .B0 (n_4726), .B1(n_10874), .Y (n_4727));
AOI21X1 g63304(.A0 (n_10874), .A1 (g2671), .B0 (n_4192), .Y (n_4725));
AOI21X1 g63313(.A0 (n_7025), .A1 (g1844), .B0 (n_4189), .Y (n_4723));
AOI21X1 g63315(.A0 (n_10920), .A1 (g1978), .B0 (n_4186), .Y (n_4721));
AOI21X1 g63318(.A0 (n_7102), .A1 (g2112), .B0 (n_4182), .Y (n_4719));
AOI21X1 g63322(.A0 (n_8628), .A1 (g2403), .B0 (n_4178), .Y (n_4717));
AOI21X1 g63324(.A0 (n_8633), .A1 (g2537), .B0 (n_4176), .Y (n_4716));
OAI21X1 g63326(.A0 (n_10899), .A1 (n_6027), .B0 (n_4172), .Y(n_4715));
NAND3X1 g62102(.A (n_2778), .B (n_3904), .C (n_3819), .Y (n_4714));
MX2X1 g63341(.A (n_5961), .B (n_864), .S0 (n_10097), .Y (n_4713));
XOR2X1 g63348(.A (n_6020), .B (n_10873), .Y (n_4712));
XOR2X1 g63349(.A (n_5978), .B (n_3956), .Y (n_4711));
XOR2X1 g63350(.A (n_5975), .B (n_10921), .Y (n_4710));
XOR2X1 g63351(.A (n_6017), .B (n_3953), .Y (n_4709));
XOR2X1 g63352(.A (n_5972), .B (n_3952), .Y (n_4708));
XOR2X1 g63353(.A (n_5969), .B (n_3951), .Y (n_4707));
OAI22X1 g62112(.A0 (n_4050), .A1 (n_4956), .B0 (n_3624), .B1(n_9698), .Y (n_4706));
MX2X1 g63361(.A (g3347), .B (n_3933), .S0 (n_9172), .Y (n_4705));
MX2X1 g63366(.A (g3698), .B (n_3934), .S0 (n_9311), .Y (n_4704));
CLKBUFX1 gbuf_d_652(.A(n_4196), .Y(d_out_652));
CLKBUFX1 gbuf_q_652(.A(q_in_652), .Y(n_11198));
CLKBUFX1 gbuf_d_653(.A(g16686), .Y(d_out_653));
CLKBUFX1 gbuf_q_653(.A(q_in_653), .Y(g3329));
CLKBUFX1 gbuf_d_654(.A(g16722), .Y(d_out_654));
CLKBUFX1 gbuf_q_654(.A(q_in_654), .Y(g3680));
CLKBUFX1 gbuf_d_655(.A(n_4226), .Y(d_out_655));
CLKBUFX1 gbuf_q_655(.A(q_in_655), .Y(g19357));
NAND3X1 g63482(.A (n_937), .B (n_3929), .C (n_10385), .Y (n_4700));
AOI21X1 g63494(.A0 (n_10372), .A1 (n_4301), .B0 (g2153), .Y (n_4699));
NAND3X1 g63503(.A (n_845), .B (n_3922), .C (n_9351), .Y (n_4695));
NAND2X1 g63507(.A (n_6539), .B (n_10626), .Y (n_4693));
NAND4X1 g61022(.A (n_4638), .B (n_4637), .C (n_4679), .D (n_2535), .Y(n_4690));
AOI22X1 g63548(.A0 (n_615), .A1 (n_3929), .B0 (n_10944), .B1 (g3129),.Y (n_4689));
AOI22X1 g63552(.A0 (n_638), .A1 (n_3922), .B0 (n_4447), .B1 (g3480),.Y (n_4688));
NAND3X1 g60937(.A (n_3911), .B (n_2301), .C (n_4070), .Y (n_4684));
NAND4X1 g63560(.A (n_4682), .B (g3582), .C (g13881), .D (n_10894), .Y(n_4683));
NAND4X1 g61023(.A (n_4633), .B (n_4632), .C (n_4679), .D (n_2538), .Y(n_4680));
NAND4X1 g61024(.A (n_4629), .B (n_4628), .C (n_4679), .D (n_2485), .Y(n_4678));
NAND4X1 g61025(.A (n_4618), .B (n_4679), .C (n_4617), .D (n_3383), .Y(n_4677));
MX2X1 g63629(.A (g1636), .B (g1592), .S0 (n_4108), .Y (n_4676));
MX2X1 g63630(.A (n_4120), .B (g1636), .S0 (n_4108), .Y (n_4673));
NOR3X1 g62253(.A (n_4671), .B (g_19659), .C (n_10078), .Y (n_4672));
MX2X1 g63655(.A (g5236), .B (n_4668), .S0 (n_1205), .Y (n_4670));
MX2X1 g63656(.A (g5252), .B (n_4668), .S0 (n_1225), .Y (n_4669));
MX2X1 g63657(.A (g5264), .B (n_4668), .S0 (n_1465), .Y (n_4667));
MX2X1 g63666(.A (g5583), .B (n_4668), .S0 (n_995), .Y (n_4666));
MX2X1 g63668(.A (g5599), .B (n_4668), .S0 (n_1155), .Y (n_4665));
OAI21X1 g62273(.A0 (n_2584), .A1 (n_3690), .B0 (n_4082), .Y (n_4663));
MX2X1 g63680(.A (g5929), .B (n_4668), .S0 (n_1195), .Y (n_4662));
MX2X1 g63684(.A (g5957), .B (n_4668), .S0 (n_1146), .Y (n_4661));
MX2X1 g63692(.A (g6275), .B (n_4668), .S0 (n_1159), .Y (n_4660));
MX2X1 g63696(.A (g6299), .B (n_4668), .S0 (n_1469), .Y (n_4659));
MX2X1 g63697(.A (g6303), .B (n_4668), .S0 (n_1144), .Y (n_4658));
MX2X1 g63698(.A (g6307), .B (n_4668), .S0 (n_1467), .Y (n_4657));
MX2X1 g63709(.A (g5260), .B (n_4668), .S0 (n_1228), .Y (n_4656));
CLKBUFX1 gbuf_d_656(.A(n_4250), .Y(d_out_656));
CLKBUFX1 gbuf_q_656(.A(q_in_656), .Y(g_13278));
MX2X1 g63748(.A (g3945), .B (n_4668), .S0 (n_1182), .Y (n_4655));
MX2X1 g63749(.A (g3953), .B (n_4668), .S0 (n_1176), .Y (n_4654));
MX2X1 g63753(.A (g6637), .B (n_4668), .S0 (n_1423), .Y (n_4653));
MX2X1 g63755(.A (g6645), .B (n_4668), .S0 (n_1428), .Y (n_4652));
XOR2X1 g63766(.A (n_2686), .B (n_3929), .Y (n_4651));
XOR2X1 g63767(.A (n_2699), .B (n_3922), .Y (n_4650));
MX2X1 g63782(.A (g2040), .B (g1996), .S0 (n_6758), .Y (n_4649));
MX2X1 g63783(.A (g2070), .B (g2040), .S0 (n_6758), .Y (n_4647));
MX2X1 g63784(.A (g2599), .B (g2555), .S0 (n_10978), .Y (n_4645));
AOI22X1 g62326(.A0 (n_4067), .A1 (n_9359), .B0 (n_659), .B1 (n_9693),.Y (n_4642));
MX2X1 g63785(.A (g2629), .B (g2599), .S0 (n_10978), .Y (n_4640));
NAND3X1 g61039(.A (n_4638), .B (n_4637), .C (n_4631), .Y (n_4639));
MX2X1 g63808(.A (n_10568), .B (n_3905), .S0 (n_9000), .Y (n_4636));
NAND3X1 g61040(.A (n_4633), .B (n_4632), .C (n_4631), .Y (n_4634));
NAND3X1 g61041(.A (n_4629), .B (n_4628), .C (n_4631), .Y (n_4630));
NAND2X1 g61637(.A (n_3755), .B (n_4090), .Y (n_4627));
NAND2X1 g61638(.A (n_3753), .B (n_4092), .Y (n_4626));
CLKBUFX1 gbuf_d_657(.A(g13906), .Y(d_out_657));
CLKBUFX1 gbuf_q_657(.A(q_in_657), .Y(g16748));
NAND3X1 g63869(.A (n_4265), .B (n_4055), .C (n_3903), .Y (n_4625));
NAND3X1 g63870(.A (n_4072), .B (n_4066), .C (n_3736), .Y (n_4624));
NAND3X1 g63871(.A (n_4074), .B (n_4065), .C (n_3735), .Y (n_4623));
NAND3X1 g63872(.A (n_4073), .B (n_4056), .C (n_3734), .Y (n_4622));
NAND3X1 g63873(.A (n_4071), .B (n_4060), .C (n_3733), .Y (n_4621));
NAND3X1 g63874(.A (n_4264), .B (n_4062), .C (n_3902), .Y (n_4620));
NAND3X1 g61043(.A (n_4618), .B (n_4631), .C (n_4617), .Y (n_4619));
INVX1 g63908(.A (n_4615), .Y (n_4616));
NAND3X1 g63932(.A (n_6754), .B (g2084), .C (n_9558), .Y (n_4614));
NAND3X1 g63967(.A (n_10982), .B (n_902), .C (n_9811), .Y (n_4611));
CLKBUFX1 gbuf_d_658(.A(n_4233), .Y(d_out_658));
CLKBUFX1 gbuf_q_658(.A(q_in_658), .Y(g7946));
NAND4X1 g64052(.A (g3917), .B (n_5402), .C (g16955), .D (n_6808), .Y(n_4607));
CLKBUFX1 gbuf_d_659(.A(n_4227), .Y(d_out_659));
CLKBUFX1 gbuf_q_659(.A(q_in_659), .Y(g4776));
CLKBUFX1 gbuf_d_660(.A(n_4201), .Y(d_out_660));
CLKBUFX1 gbuf_q_660(.A(q_in_660), .Y(g4966));
CLKBUFX1 gbuf_d_661(.A(n_4148), .Y(d_out_661));
CLKBUFX1 gbuf_q_661(.A(q_in_661), .Y(g_19414));
CLKBUFX1 gbuf_d_662(.A(n_4136), .Y(d_out_662));
CLKBUFX1 gbuf_q_662(.A(q_in_662), .Y(g4785));
CLKBUFX1 gbuf_d_663(.A(n_4081), .Y(d_out_663));
CLKBUFX1 gbuf_q_663(.A(q_in_663), .Y(n_662));
CLKBUFX1 gbuf_d_664(.A(n_4083), .Y(d_out_664));
CLKBUFX1 gbuf_q_664(.A(q_in_664), .Y(g4899));
NAND4X1 g64042(.A (g3925), .B (n_3894), .C (g16955), .D (n_8917), .Y(n_4605));
CLKBUFX1 gbuf_d_665(.A(n_4199), .Y(d_out_665));
CLKBUFX1 gbuf_q_665(.A(q_in_665), .Y(n_8807));
CLKBUFX1 gbuf_d_666(.A(n_4193), .Y(d_out_666));
CLKBUFX1 gbuf_q_666(.A(q_in_666), .Y(g6741));
OAI21X1 g61270(.A0 (n_8761), .A1 (n_8628), .B0 (n_4179), .Y (n_4603));
CLKBUFX1 gbuf_d_667(.A(n_4194), .Y(d_out_667));
CLKBUFX1 gbuf_q_667(.A(q_in_667), .Y(g6395));
CLKBUFX1 gbuf_d_668(.A(n_4137), .Y(d_out_668));
CLKBUFX1 gbuf_q_668(.A(q_in_668), .Y(g_14265));
CLKBUFX1 gbuf_d_669(.A(n_4135), .Y(d_out_669));
CLKBUFX1 gbuf_q_669(.A(q_in_669), .Y(g_12791));
CLKBUFX1 gbuf_d_670(.A(n_4110), .Y(d_out_670));
CLKBUFX1 gbuf_q_670(.A(q_in_670), .Y(g_20268));
NAND3X1 g60953(.A (n_4030), .B (n_11220), .C (n_1442), .Y (n_4600));
NAND4X1 g62648(.A (n_4260), .B (n_3442), .C (n_3026), .D (n_3022), .Y(g28030));
CLKBUFX1 gbuf_d_671(.A(n_4263), .Y(d_out_671));
CLKBUFX1 gbuf_qn_671(.A(qn_in_671), .Y(g4369));
NAND3X1 g60955(.A (n_4568), .B (g1373), .C (n_9811), .Y (n_4598));
CLKBUFX1 gbuf_d_672(.A(g14096), .Y(d_out_672));
CLKBUFX1 gbuf_q_672(.A(q_in_672), .Y(g14125));
OAI21X1 g61276(.A0 (n_8763), .A1 (n_8633), .B0 (n_4177), .Y (n_4597));
OAI21X1 g61282(.A0 (n_11191), .A1 (n_10874), .B0 (n_4175), .Y(n_4594));
INVX1 g60956(.A (n_4592), .Y (n_4593));
OAI21X1 g60958(.A0 (n_367), .A1 (n_9425), .B0 (n_4246), .Y (n_4591));
NOR2X1 g62576(.A (n_4253), .B (g4704), .Y (n_4590));
NAND3X1 g62598(.A (n_4054), .B (n_2528), .C (n_4028), .Y (n_4589));
NAND2X1 g62609(.A (n_4254), .B (n_3846), .Y (n_4587));
AOI22X1 g60960(.A0 (n_4017), .A1 (n_2586), .B0 (g1542), .B1 (n_9903),.Y (n_4586));
NOR2X1 g62654(.A (n_3243), .B (g4045), .Y (n_4585));
NOR2X1 g61313(.A (n_10761), .B (n_4583), .Y (n_4584));
NOR2X1 g61325(.A (n_940), .B (n_4582), .Y (n_4968));
CLKBUFX1 gbuf_d_673(.A(n_4266), .Y(d_out_673));
CLKBUFX1 gbuf_q_673(.A(q_in_673), .Y(n_11129));
NAND2X1 g61795(.A (n_8757), .B (g4608), .Y (n_4581));
CLKBUFX1 gbuf_d_674(.A(n_4048), .Y(d_out_674));
CLKBUFX1 gbuf_qn_674(.A(qn_in_674), .Y(g2856));
OAI21X1 g61834(.A0 (n_4045), .A1 (g_14342), .B0 (n_4578), .Y(n_4579));
NAND3X1 g62807(.A (n_3843), .B (n_2286), .C (n_3824), .Y (n_4577));
INVX1 g62816(.A (n_5723), .Y (n_4576));
CLKBUFX1 gbuf_d_675(.A(n_4044), .Y(d_out_675));
CLKBUFX1 gbuf_q_675(.A(q_in_675), .Y(g2748));
OAI21X1 g62840(.A0 (n_4053), .A1 (g_20159), .B0 (n_4202), .Y(n_4810));
NOR2X1 g60978(.A (n_4031), .B (n_4284), .Y (n_4575));
OAI21X1 g62897(.A0 (g2927), .A1 (n_9311), .B0 (n_4029), .Y (n_4574));
OAI21X1 g60980(.A0 (n_10245), .A1 (n_9333), .B0 (n_3995), .Y(n_4573));
NAND4X1 g62918(.A (n_10700), .B (n_3984), .C (n_9359), .D (g5057), .Y(n_4572));
AOI21X1 g62920(.A0 (n_3001), .A1 (n_521), .B0 (n_4022), .Y (n_8879));
OAI22X1 g62927(.A0 (n_3625), .A1 (n_4956), .B0 (n_448), .B1 (n_9862),.Y (n_4570));
INVX1 g60981(.A (n_4568), .Y (n_4569));
MX2X1 g62933(.A (n_3836), .B (g5698), .S0 (n_10660), .Y (n_4567));
MX2X1 g62934(.A (n_3835), .B (g6044), .S0 (n_11201), .Y (n_4566));
MX2X1 g62935(.A (n_3834), .B (g6390), .S0 (g6395), .Y (n_4565));
MX2X1 g62936(.A (n_3833), .B (g6736), .S0 (n_523), .Y (n_4564));
MX2X1 g62939(.A (g5037), .B (n_3825), .S0 (n_9091), .Y (n_4563));
AOI21X1 g61370(.A0 (n_3838), .A1 (n_4558), .B0 (n_3837), .Y (n_4562));
MX2X1 g62943(.A (g5138), .B (n_3809), .S0 (n_8955), .Y (n_4561));
MX2X1 g65047(.A (g6744), .B (g_13901), .S0 (n_9599), .Y (n_4560));
AOI21X1 g61376(.A0 (n_3832), .A1 (n_4558), .B0 (n_3831), .Y (n_4559));
CLKBUFX1 gbuf_d_676(.A(n_3966), .Y(d_out_676));
CLKBUFX1 gbuf_q_676(.A(q_in_676), .Y(g_19233));
INVX1 g65194(.A (n_7097), .Y (g11678));
MX2X1 g63046(.A (g6513), .B (n_3815), .S0 (n_9359), .Y (n_4557));
AOI21X1 g65434(.A0 (n_4231), .A1 (n_326), .B0 (n_4037), .Y (n_4556));
AOI21X1 g65435(.A0 (n_4231), .A1 (n_317), .B0 (n_4033), .Y (n_4555));
INVX1 g61968(.A (n_8758), .Y (n_4554));
CLKBUFX1 gbuf_d_677(.A(n_4011), .Y(d_out_677));
CLKBUFX1 gbuf_q_677(.A(q_in_677), .Y(g6736));
MX2X1 g63142(.A (g_8896), .B (n_3823), .S0 (n_9256), .Y (n_4553));
CLKBUFX1 gbuf_d_678(.A(n_3970), .Y(d_out_678));
CLKBUFX1 gbuf_q_678(.A(q_in_678), .Y(g1389));
NAND2X1 g63198(.A (n_3982), .B (n_3830), .Y (n_4550));
CLKBUFX1 gbuf_d_679(.A(n_4013), .Y(d_out_679));
CLKBUFX1 gbuf_q_679(.A(q_in_679), .Y(g_15838));
NAND2X1 g63207(.A (n_3813), .B (n_3997), .Y (n_4547));
NAND2X1 g63223(.A (n_9129), .B (g18881), .Y (n_4546));
NOR3X1 g63245(.A (n_9505), .B (g5057), .C (n_10700), .Y (n_4545));
INVX1 g63266(.A (n_4541), .Y (n_4542));
NOR2X1 g61473(.A (n_4743), .B (n_4539), .Y (n_4540));
OAI21X1 g63272(.A0 (n_3792), .A1 (n_9129), .B0 (n_3937), .Y (n_4538));
OAI21X1 g63273(.A0 (n_3788), .A1 (n_9599), .B0 (n_4040), .Y (n_4537));
OAI21X1 g63274(.A0 (n_3786), .A1 (n_9672), .B0 (n_3706), .Y (n_4535));
OAI21X1 g63275(.A0 (n_3785), .A1 (n_9107), .B0 (n_3936), .Y (n_4534));
OAI21X1 g63277(.A0 (n_3781), .A1 (n_9443), .B0 (n_4059), .Y (n_4533));
AOI22X1 g63284(.A0 (n_905), .A1 (n_10857), .B0 (n_4531), .B1(n_8633), .Y (n_4532));
AOI22X1 g63301(.A0 (n_912), .A1 (n_10675), .B0 (n_4529), .B1(n_8628), .Y (n_4530));
MX2X1 g63333(.A (n_4893), .B (n_4527), .S0 (n_10899), .Y (n_4528));
MX2X1 g63334(.A (n_5958), .B (n_716), .S0 (n_10874), .Y (n_4526));
MX2X1 g63337(.A (n_5964), .B (n_856), .S0 (n_10899), .Y (n_4525));
MX2X1 g63338(.A (n_4948), .B (n_854), .S0 (n_7025), .Y (n_4524));
MX2X1 g63339(.A (n_4946), .B (n_871), .S0 (n_10920), .Y (n_4523));
MX2X1 g63340(.A (n_5953), .B (n_862), .S0 (n_7102), .Y (n_4522));
MX2X1 g63342(.A (n_4942), .B (n_846), .S0 (n_8628), .Y (n_4521));
MX2X1 g63344(.A (n_5229), .B (n_714), .S0 (n_8633), .Y (n_4520));
XOR2X1 g62113(.A (g4601), .B (n_8885), .Y (n_4519));
MX2X1 g63367(.A (g4049), .B (n_3770), .S0 (n_9311), .Y (n_4518));
AOI21X1 g63490(.A0 (n_6759), .A1 (n_3943), .B0 (g1996), .Y (n_4516));
NAND2X1 g63495(.A (n_1518), .B (n_10097), .Y (n_4515));
NOR2X1 g63497(.A (n_10099), .B (n_8755), .Y (n_4514));
NAND2X1 g63500(.A (n_10097), .B (n_6025), .Y (n_4513));
AOI21X1 g63523(.A0 (g13895), .A1 (n_464), .B0 (n_3942), .Y (n_4512));
AOI21X1 g63524(.A0 (g13926), .A1 (n_11088), .B0 (n_3941), .Y(n_4510));
OAI21X1 g63541(.A0 (g2878), .A1 (n_9992), .B0 (n_3955), .Y (n_4508));
CLKBUFX1 gbuf_d_680(.A(n_3932), .Y(d_out_680));
CLKBUFX1 gbuf_q_680(.A(q_in_680), .Y(g1536));
MX2X1 g63571(.A (n_4497), .B (g5244), .S0 (n_1401), .Y (n_4507));
NOR2X1 g62207(.A (n_3906), .B (n_9836), .Y (n_4506));
MX2X1 g63572(.A (n_4499), .B (g5248), .S0 (n_1404), .Y (n_4504));
MX2X1 g63573(.A (n_4494), .B (g5256), .S0 (n_1463), .Y (n_4503));
MX2X1 g63575(.A (n_4494), .B (g5563), .S0 (n_1761), .Y (n_4502));
MX2X1 g63576(.A (n_4499), .B (g5575), .S0 (n_1322), .Y (n_4501));
MX2X1 g63577(.A (n_4499), .B (g5579), .S0 (n_1413), .Y (n_4500));
MX2X1 g63578(.A (n_4497), .B (g5591), .S0 (n_1397), .Y (n_4498));
MX2X1 g63579(.A (n_4482), .B (g5595), .S0 (n_1408), .Y (n_4496));
MX2X1 g63580(.A (n_4494), .B (g5603), .S0 (n_1477), .Y (n_4495));
MX2X1 g63581(.A (n_4494), .B (g5216), .S0 (n_1738), .Y (n_4493));
MX2X1 g63583(.A (n_4499), .B (g5909), .S0 (n_1728), .Y (n_4492));
MX2X1 g63584(.A (n_4482), .B (g5921), .S0 (n_1108), .Y (n_4490));
MX2X1 g63585(.A (n_4499), .B (g5925), .S0 (n_1114), .Y (n_4489));
MX2X1 g63586(.A (n_4494), .B (g5937), .S0 (n_1120), .Y (n_4488));
MX2X1 g63587(.A (n_4499), .B (g5941), .S0 (n_1104), .Y (n_4487));
MX2X1 g63588(.A (n_4494), .B (g5949), .S0 (n_1452), .Y (n_4486));
MX2X1 g63590(.A (g3119), .B (n_0), .S0 (n_10944), .Y (n_4485));
MX2X1 g63591(.A (n_4482), .B (g6255), .S0 (n_1721), .Y (n_4483));
MX2X1 g63592(.A (n_4494), .B (g6267), .S0 (n_1128), .Y (n_4481));
MX2X1 g63593(.A (n_4499), .B (g6271), .S0 (n_1107), .Y (n_4479));
MX2X1 g63594(.A (n_4497), .B (g6283), .S0 (n_1127), .Y (n_4478));
MX2X1 g63595(.A (n_4482), .B (g6287), .S0 (n_1106), .Y (n_4477));
MX2X1 g63596(.A (n_4494), .B (g3207), .S0 (n_1748), .Y (n_4475));
MX2X1 g63598(.A (n_4482), .B (g3219), .S0 (n_1102), .Y (n_4474));
MX2X1 g63599(.A (n_4499), .B (g3223), .S0 (n_1105), .Y (n_4473));
MX2X1 g63600(.A (n_4482), .B (g3235), .S0 (n_1121), .Y (n_4472));
MX2X1 g63601(.A (n_4482), .B (g3239), .S0 (n_1123), .Y (n_4471));
MX2X1 g63602(.A (n_4494), .B (g6613), .S0 (n_1122), .Y (n_4470));
MX2X1 g63603(.A (n_4497), .B (g3247), .S0 (n_1418), .Y (n_4469));
MX2X1 g63604(.A (n_4497), .B (g6601), .S0 (n_1730), .Y (n_4468));
MX2X1 g63605(.A (n_4494), .B (g6641), .S0 (n_1415), .Y (n_4467));
MX2X1 g63607(.A (n_4497), .B (g3558), .S0 (n_1749), .Y (n_4466));
MX2X1 g63608(.A (n_4499), .B (g3570), .S0 (n_1119), .Y (n_4465));
MX2X1 g63609(.A (n_4494), .B (g3574), .S0 (n_1118), .Y (n_4464));
MX2X1 g63610(.A (n_4494), .B (g3586), .S0 (n_1117), .Y (n_4462));
MX2X1 g63611(.A (n_4482), .B (g3590), .S0 (n_1116), .Y (n_4461));
MX2X1 g63612(.A (n_4494), .B (g3598), .S0 (n_1447), .Y (n_4460));
MX2X1 g63613(.A (n_4482), .B (g5232), .S0 (n_1400), .Y (n_4459));
MX2X1 g63615(.A (n_4482), .B (g5228), .S0 (n_1398), .Y (n_4458));
MX2X1 g63617(.A (n_4499), .B (g3909), .S0 (n_1740), .Y (n_4457));
MX2X1 g63618(.A (n_4497), .B (g3921), .S0 (n_1112), .Y (n_4456));
MX2X1 g63619(.A (n_4494), .B (g3925), .S0 (n_1111), .Y (n_4455));
MX2X1 g63620(.A (n_4494), .B (g3937), .S0 (n_1130), .Y (n_4454));
MX2X1 g63621(.A (n_4482), .B (g3941), .S0 (n_1110), .Y (n_4453));
MX2X1 g63622(.A (n_4482), .B (g3949), .S0 (n_1435), .Y (n_4452));
MX2X1 g63626(.A (n_4497), .B (g6633), .S0 (n_1392), .Y (n_4451));
MX2X1 g63627(.A (n_4494), .B (g6295), .S0 (n_1433), .Y (n_4450));
MX2X1 g63628(.A (n_4482), .B (g6629), .S0 (n_1393), .Y (n_4449));
MX2X1 g63631(.A (g3470), .B (n_60), .S0 (n_4447), .Y (n_4448));
MX2X1 g63632(.A (n_4482), .B (g6617), .S0 (n_1103), .Y (n_4446));
AOI22X1 g63637(.A0 (n_3609), .A1 (n_9443), .B0 (n_10944), .B1(n_901), .Y (n_4445));
AOI22X1 g63639(.A0 (n_3601), .A1 (n_10078), .B0 (n_4447), .B1(n_2019), .Y (n_4444));
MX2X1 g63649(.A (n_4497), .B (g5196), .S0 (n_1775), .Y (n_4442));
MX2X1 g63650(.A (n_4499), .B (g5200), .S0 (n_1764), .Y (n_4441));
MX2X1 g63651(.A (n_4482), .B (g5204), .S0 (n_1481), .Y (n_4440));
MX2X1 g63652(.A (n_4499), .B (g5208), .S0 (n_1605), .Y (n_4439));
MX2X1 g63653(.A (n_4499), .B (g5220), .S0 (n_1178), .Y (n_4438));
MX2X1 g63654(.A (n_4482), .B (g5224), .S0 (n_1438), .Y (n_4437));
MX2X1 g63658(.A (n_4497), .B (g6235), .S0 (n_1779), .Y (n_4436));
MX2X1 g63659(.A (g5272), .B (n_4497), .S0 (g26801), .Y (n_4434));
MX2X1 g63660(.A (n_4497), .B (g5543), .S0 (n_1773), .Y (n_4433));
MX2X1 g63661(.A (n_4497), .B (g5547), .S0 (n_1778), .Y (n_4432));
MX2X1 g63662(.A (n_4499), .B (g5551), .S0 (n_1425), .Y (n_4431));
MX2X1 g63663(.A (n_4499), .B (g5559), .S0 (n_1131), .Y (n_4430));
MX2X1 g63664(.A (n_4499), .B (g5567), .S0 (n_1235), .Y (n_4429));
MX2X1 g63665(.A (n_4482), .B (g5571), .S0 (n_1466), .Y (n_4428));
MX2X1 g63667(.A (n_4482), .B (g5587), .S0 (n_1424), .Y (n_4427));
MX2X1 g63669(.A (g5607), .B (n_4424), .S0 (n_1187), .Y (n_4426));
MX2X1 g63670(.A (g5611), .B (n_4424), .S0 (n_1223), .Y (n_4425));
MX2X1 g63671(.A (g5615), .B (n_4424), .S0 (n_1239), .Y (n_4423));
OAI21X1 g62272(.A0 (n_3885), .A1 (n_1285), .B0 (n_3184), .Y (n_4422));
MX2X1 g63672(.A (n_4482), .B (g5619), .S0 (n_4329), .Y (n_4421));
MX2X1 g63673(.A (n_4497), .B (g5889), .S0 (n_1722), .Y (n_4420));
MX2X1 g63674(.A (n_4482), .B (g5893), .S0 (n_1726), .Y (n_4419));
MX2X1 g63675(.A (n_4482), .B (g5897), .S0 (n_1437), .Y (n_4418));
MX2X1 g63676(.A (n_4494), .B (g5901), .S0 (n_1755), .Y (n_4417));
MX2X1 g63677(.A (n_4499), .B (g5905), .S0 (n_1170), .Y (n_4416));
MX2X1 g63678(.A (n_4499), .B (g5913), .S0 (n_999), .Y (n_4415));
MX2X1 g63679(.A (n_4499), .B (g5917), .S0 (n_1456), .Y (n_4414));
MX2X1 g63681(.A (n_4499), .B (g5933), .S0 (n_1431), .Y (n_4413));
MX2X1 g63682(.A (g6621), .B (n_4424), .S0 (n_1152), .Y (n_4412));
MX2X1 g63683(.A (g5945), .B (n_4497), .S0 (n_1247), .Y (n_4411));
MX2X1 g63685(.A (g5961), .B (n_4497), .S0 (n_910), .Y (n_4410));
MX2X1 g63686(.A (n_4482), .B (g5965), .S0 (n_4327), .Y (n_4409));
MX2X1 g63687(.A (n_4494), .B (g6243), .S0 (n_1419), .Y (n_4408));
MX2X1 g63688(.A (n_4482), .B (g6247), .S0 (n_1771), .Y (n_4407));
MX2X1 g63689(.A (n_4482), .B (g6251), .S0 (n_1215), .Y (n_4406));
MX2X1 g63690(.A (n_4497), .B (g6259), .S0 (n_1153), .Y (n_4405));
MX2X1 g63691(.A (n_4482), .B (g6263), .S0 (n_1472), .Y (n_4404));
MX2X1 g63693(.A (g5953), .B (n_4424), .S0 (n_1460), .Y (n_4403));
MX2X1 g63694(.A (n_4494), .B (g6279), .S0 (n_1470), .Y (n_4402));
MX2X1 g63695(.A (g6291), .B (n_4424), .S0 (n_1150), .Y (n_4401));
MX2X1 g63699(.A (g5268), .B (n_4424), .S0 (n_1232), .Y (n_4400));
MX2X1 g63700(.A (n_4494), .B (g6311), .S0 (n_4324), .Y (n_4399));
MX2X1 g63701(.A (n_4497), .B (g3187), .S0 (n_1769), .Y (n_4398));
MX2X1 g63702(.A (n_4499), .B (g3191), .S0 (n_1759), .Y (n_4397));
MX2X1 g63703(.A (n_4499), .B (g3195), .S0 (n_1427), .Y (n_4396));
MX2X1 g63704(.A (n_4494), .B (g3199), .S0 (n_1768), .Y (n_4395));
MX2X1 g63705(.A (n_4497), .B (g3211), .S0 (n_1136), .Y (n_4394));
MX2X1 g63707(.A (n_4499), .B (g3203), .S0 (n_993), .Y (n_4393));
MX2X1 g63706(.A (n_4482), .B (g3215), .S0 (n_1585), .Y (n_4392));
MX2X1 g63708(.A (g3227), .B (n_4424), .S0 (n_1244), .Y (n_4391));
MX2X1 g63710(.A (n_4499), .B (g3231), .S0 (n_1478), .Y (n_4390));
MX2X1 g63711(.A (n_4499), .B (g6593), .S0 (n_1780), .Y (n_4389));
MX2X1 g63712(.A (n_4497), .B (g6581), .S0 (n_1766), .Y (n_4388));
MX2X1 g63713(.A (g3243), .B (n_4497), .S0 (n_1148), .Y (n_4387));
MX2X1 g63714(.A (g3255), .B (n_4497), .S0 (n_1483), .Y (n_4386));
MX2X1 g63715(.A (g3259), .B (n_4497), .S0 (n_897), .Y (n_4385));
MX2X1 g63716(.A (g6649), .B (n_4424), .S0 (n_1487), .Y (n_4384));
MX2X1 g63717(.A (g6653), .B (n_4424), .S0 (n_1326), .Y (n_4383));
MX2X1 g63718(.A (n_4494), .B (g6657), .S0 (n_4322), .Y (n_4382));
MX2X1 g63719(.A (n_4497), .B (g5240), .S0 (n_1453), .Y (n_4381));
MX2X1 g63720(.A (g3251), .B (n_4497), .S0 (n_1475), .Y (n_4380));
MX2X1 g63721(.A (n_4494), .B (g3538), .S0 (n_1754), .Y (n_4379));
MX2X1 g63722(.A (n_4499), .B (g3542), .S0 (n_1753), .Y (n_4378));
MX2X1 g63723(.A (n_4499), .B (g3546), .S0 (n_1451), .Y (n_4377));
MX2X1 g63724(.A (n_4494), .B (g3550), .S0 (n_1750), .Y (n_4376));
MX2X1 g63725(.A (n_4497), .B (g3554), .S0 (n_1211), .Y (n_4375));
MX2X1 g63726(.A (n_4494), .B (g3562), .S0 (n_1209), .Y (n_4374));
MX2X1 g63727(.A (n_4494), .B (g3566), .S0 (n_1449), .Y (n_4373));
MX2X1 g63728(.A (g3578), .B (n_4424), .S0 (n_1208), .Y (n_4372));
MX2X1 g63729(.A (n_4494), .B (g3582), .S0 (n_1448), .Y (n_4371));
MX2X1 g63730(.A (g3594), .B (n_4424), .S0 (n_1202), .Y (n_4370));
MX2X1 g63731(.A (n_4482), .B (g6609), .S0 (n_1432), .Y (n_4369));
MX2X1 g63732(.A (g3602), .B (n_4424), .S0 (n_1200), .Y (n_4368));
MX2X1 g63733(.A (g3606), .B (n_4424), .S0 (n_1198), .Y (n_4367));
MX2X1 g63734(.A (n_4499), .B (g6589), .S0 (n_1446), .Y (n_4366));
MX2X1 g63735(.A (g3610), .B (n_4424), .S0 (n_931), .Y (n_4365));
MX2X1 g63736(.A (n_4497), .B (g3614), .S0 (n_4320), .Y (n_4364));
MX2X1 g63737(.A (n_4499), .B (g6597), .S0 (n_1217), .Y (n_4363));
MX2X1 g63738(.A (n_4497), .B (g3889), .S0 (n_1746), .Y (n_4362));
MX2X1 g63739(.A (n_4482), .B (g3893), .S0 (n_1745), .Y (n_4361));
MX2X1 g63740(.A (n_4497), .B (g6239), .S0 (n_1724), .Y (n_4360));
MX2X1 g63741(.A (n_4494), .B (g3897), .S0 (n_1441), .Y (n_4359));
MX2X1 g63742(.A (n_4499), .B (g3901), .S0 (n_1741), .Y (n_4358));
MX2X1 g63743(.A (n_4482), .B (g3905), .S0 (n_1192), .Y (n_4357));
MX2X1 g63744(.A (n_4482), .B (g3913), .S0 (n_1189), .Y (n_4356));
MX2X1 g63745(.A (n_4494), .B (g3917), .S0 (n_1439), .Y (n_4355));
MX2X1 g63746(.A (g3929), .B (n_4424), .S0 (n_1186), .Y (n_4354));
MX2X1 g63747(.A (n_4482), .B (g3933), .S0 (n_1436), .Y (n_4353));
MX2X1 g63750(.A (g3957), .B (n_4497), .S0 (n_1174), .Y (n_4352));
MX2X1 g63751(.A (g3961), .B (n_4497), .S0 (n_921), .Y (n_4351));
MX2X1 g63752(.A (n_4499), .B (g3965), .S0 (n_4314), .Y (n_4350));
MX2X1 g63754(.A (n_4499), .B (g6605), .S0 (n_1167), .Y (n_4349));
MX2X1 g63756(.A (n_4494), .B (g3263), .S0 (n_4316), .Y (n_4348));
MX2X1 g63758(.A (n_4482), .B (g5212), .S0 (n_1164), .Y (n_4347));
MX2X1 g63759(.A (n_4494), .B (g6585), .S0 (n_1719), .Y (n_4346));
MX2X1 g63760(.A (n_4497), .B (g5555), .S0 (n_1716), .Y (n_4345));
MX2X1 g63761(.A (n_4494), .B (g6625), .S0 (n_1416), .Y (n_4344));
MX2X1 g63773(.A (g2465), .B (g2421), .S0 (n_10853), .Y (n_4343));
MX2X1 g63774(.A (n_4339), .B (g2465), .S0 (n_10853), .Y (n_4340));
MX2X1 g63778(.A (g_12791), .B (n_3745), .S0 (n_9992), .Y (n_4338));
MX2X1 g63779(.A (g2331), .B (g2287), .S0 (n_10671), .Y (n_4336));
MX2X1 g63780(.A (g2361), .B (g2331), .S0 (n_10671), .Y (n_4333));
NAND3X1 g63868(.A (n_4076), .B (n_3883), .C (n_3737), .Y (n_4331));
AND2X1 g63909(.A (n_4424), .B (n_1812), .Y (n_4615));
AND2X1 g63914(.A (n_4329), .B (n_4668), .Y (n_4330));
AND2X1 g63917(.A (n_4327), .B (n_4668), .Y (n_4328));
AND2X1 g63922(.A (n_4324), .B (n_4668), .Y (n_4325));
AND2X1 g63923(.A (n_4668), .B (n_4322), .Y (n_4323));
AND2X1 g63929(.A (n_4320), .B (n_4668), .Y (n_4321));
NOR2X1 g63930(.A (n_4304), .B (n_4318), .Y (n_4319));
AND2X1 g63931(.A (n_4316), .B (n_4668), .Y (n_4317));
AND2X1 g63933(.A (n_4314), .B (n_4668), .Y (n_4315));
INVX1 g63940(.A (n_10626), .Y (n_4313));
NAND3X1 g63952(.A (n_10670), .B (n_911), .C (n_9091), .Y (n_10549));
NAND3X1 g63958(.A (n_10852), .B (n_904), .C (n_10005), .Y (n_4308));
NOR2X1 g63971(.A (n_670), .B (n_4304), .Y (n_4306));
NOR2X1 g63973(.A (n_290), .B (n_4304), .Y (n_4305));
NOR2X1 g63974(.A (n_667), .B (n_4304), .Y (n_4303));
NAND4X1 g64001(.A (n_3907), .B (n_3371), .C (n_10063), .D (n_3486),.Y (n_4302));
NAND3X1 g64002(.A (n_4299), .B (n_4301), .C (g2153), .Y (n_4836));
NAND3X1 g64004(.A (n_10372), .B (g2197), .C (n_259), .Y (n_4834));
NAND3X1 g64005(.A (n_4299), .B (g2227), .C (g2153), .Y (n_4829));
CLKBUFX1 gbuf_d_681(.A(n_4010), .Y(d_out_681));
CLKBUFX1 gbuf_q_681(.A(q_in_681), .Y(g_16792));
NAND3X1 g64007(.A (n_4299), .B (n_4301), .C (g2227), .Y (n_4827));
CLKBUFX1 gbuf_d_682(.A(n_3969), .Y(d_out_682));
CLKBUFX1 gbuf_q_682(.A(q_in_682), .Y(g10527));
NAND3X1 g60952(.A (n_3702), .B (n_2779), .C (n_3848), .Y (n_4298));
CLKBUFX1 gbuf_d_683(.A(n_3979), .Y(d_out_683));
CLKBUFX1 gbuf_q_683(.A(q_in_683), .Y(g4709));
CLKBUFX1 gbuf_d_684(.A(n_4069), .Y(d_out_684));
CLKBUFX1 gbuf_q_684(.A(q_in_684), .Y(g_13091));
CLKBUFX1 gbuf_d_685(.A(n_4015), .Y(d_out_685));
CLKBUFX1 gbuf_q_685(.A(q_in_685), .Y(g5698));
CLKBUFX1 gbuf_d_686(.A(n_4014), .Y(d_out_686));
CLKBUFX1 gbuf_q_686(.A(q_in_686), .Y(g6044));
CLKBUFX1 gbuf_d_687(.A(n_4012), .Y(d_out_687));
CLKBUFX1 gbuf_q_687(.A(q_in_687), .Y(g6390));
CLKBUFX1 gbuf_d_688(.A(n_4016), .Y(d_out_688));
CLKBUFX1 gbuf_q_688(.A(q_in_688), .Y(g5352));
CLKBUFX1 gbuf_d_689(.A(n_4008), .Y(d_out_689));
CLKBUFX1 gbuf_q_689(.A(q_in_689), .Y(g19334));
CLKBUFX1 gbuf_d_690(.A(n_4009), .Y(d_out_690));
CLKBUFX1 gbuf_q_690(.A(q_in_690), .Y(g4176));
CLKBUFX1 gbuf_d_691(.A(n_3991), .Y(d_out_691));
CLKBUFX1 gbuf_q_691(.A(q_in_691), .Y(g11447));
CLKBUFX1 gbuf_d_692(.A(n_3981), .Y(d_out_692));
CLKBUFX1 gbuf_q_692(.A(q_in_692), .Y(g_8896));
CLKBUFX1 gbuf_d_693(.A(n_3968), .Y(d_out_693));
CLKBUFX1 gbuf_q_693(.A(q_in_693), .Y(g_15740));
CLKBUFX1 gbuf_d_694(.A(n_3964), .Y(d_out_694));
CLKBUFX1 gbuf_q_694(.A(q_in_694), .Y(n_11163));
CLKBUFX1 gbuf_d_695(.A(n_3963), .Y(d_out_695));
CLKBUFX1 gbuf_q_695(.A(q_in_695), .Y(g_21778));
CLKBUFX1 gbuf_d_696(.A(n_3962), .Y(d_out_696));
CLKBUFX1 gbuf_q_696(.A(q_in_696), .Y(g_17065));
CLKBUFX1 gbuf_d_697(.A(n_3960), .Y(d_out_697));
CLKBUFX1 gbuf_q_697(.A(q_in_697), .Y(g_16677));
CLKBUFX1 gbuf_d_698(.A(n_3959), .Y(d_out_698));
CLKBUFX1 gbuf_q_698(.A(q_in_698), .Y(g_21720));
CLKBUFX1 gbuf_d_699(.A(n_3958), .Y(d_out_699));
CLKBUFX1 gbuf_q_699(.A(q_in_699), .Y(g_13758));
CLKBUFX1 gbuf_d_700(.A(n_3957), .Y(d_out_700));
CLKBUFX1 gbuf_q_700(.A(q_in_700), .Y(g_19289));
CLKBUFX1 gbuf_d_701(.A(n_3947), .Y(d_out_701));
CLKBUFX1 gbuf_q_701(.A(q_in_701), .Y(n_640));
CLKBUFX1 gbuf_d_702(.A(n_4034), .Y(d_out_702));
CLKBUFX1 gbuf_q_702(.A(q_in_702), .Y(n_8898));
NAND3X1 g64135(.A (n_4046), .B (n_2589), .C (n_3882), .Y (n_4297));
INVX1 g64188(.A (n_6754), .Y (n_4296));
OAI21X1 g60957(.A0 (n_3910), .A1 (g1373), .B0 (n_10427), .Y (n_4592));
INVX1 g64222(.A (n_4885), .Y (n_4293));
NAND3X1 g64279(.A (n_3878), .B (n_637), .C (n_3879), .Y (n_4291));
AOI21X1 g62583(.A0 (n_3856), .A1 (n_2310), .B0 (n_9772), .Y (n_4290));
MX2X1 g64407(.A (n_11106), .B (g14217), .S0 (n_5582), .Y (n_4288));
OAI22X1 g62656(.A0 (n_3492), .A1 (n_3192), .B0 (g4366), .B1 (n_9874),.Y (n_4286));
AOI22X1 g60961(.A0 (n_4284), .A1 (n_10196), .B0 (n_1179), .B1(g7946), .Y (n_4285));
NAND2X1 g61316(.A (n_2619), .B (n_4170), .Y (n_4283));
NOR2X1 g61317(.A (n_8761), .B (n_4281), .Y (n_4282));
NOR2X1 g61318(.A (n_8762), .B (n_4279), .Y (n_4280));
NOR2X1 g61319(.A (n_8762), .B (n_4277), .Y (n_4278));
NOR2X1 g61320(.A (n_8762), .B (n_4275), .Y (n_4276));
NOR2X1 g61321(.A (n_8763), .B (n_4273), .Y (n_4274));
NOR2X1 g61322(.A (n_8764), .B (n_4271), .Y (n_4272));
NOR2X1 g61323(.A (n_8764), .B (n_4269), .Y (n_4270));
NOR2X1 g61324(.A (n_8764), .B (n_4267), .Y (n_4268));
XOR2X1 g61083(.A (g1300), .B (n_11025), .Y (n_4618));
MX2X1 g62727(.A (n_684), .B (n_3677), .S0 (n_9218), .Y (n_4266));
CLKBUFX1 gbuf_d_703(.A(n_3847), .Y(d_out_703));
CLKBUFX1 gbuf_qn_703(.A(qn_in_703), .Y(g4045));
NAND4X1 g64714(.A (g5802), .B (n_9627), .C (g9617), .D (g_7062), .Y(n_4265));
NAND4X1 g64728(.A (g3451), .B (n_9521), .C (g8279), .D (g_5313), .Y(n_4264));
MX2X1 g64778(.A (g4459), .B (g4473), .S0 (n_9091), .Y (n_4263));
AND2X1 g62805(.A (n_327), .B (g4366), .Y (n_4262));
CLKBUFX1 g62817(.A (n_7145), .Y (n_5723));
AOI21X1 g62836(.A0 (n_3287), .A1 (n_2747), .B0 (n_3852), .Y (n_4260));
OAI21X1 g62898(.A0 (n_10644), .A1 (n_9681), .B0 (n_3851), .Y(n_4257));
OR2X1 g64931(.A (g5109), .B (n_9398), .Y (n_4255));
AOI22X1 g62903(.A0 (n_3659), .A1 (n_2585), .B0 (g1199), .B1 (n_9628),.Y (n_4254));
OAI22X1 g62911(.A0 (n_10830), .A1 (g5348), .B0 (n_1058), .B1 (g5352),.Y (n_4253));
NAND4X1 g62913(.A (n_3661), .B (n_4024), .C (n_9811), .D (g_18793),.Y (n_4252));
AOI22X1 g62916(.A0 (n_10621), .A1 (g5348), .B0 (g5352), .B1 (g25114),.Y (n_4251));
OAI21X1 g62923(.A0 (n_708), .A1 (n_9311), .B0 (n_3858), .Y (n_4250));
INVX1 g60982(.A (n_10427), .Y (n_4568));
INVX1 g65050(.A (n_4247), .Y (n_4248));
NAND4X1 g60985(.A (n_4242), .B (n_9209), .C (n_4241), .D (n_2593), .Y(n_4246));
AOI21X1 g61381(.A0 (n_10323), .A1 (g1246), .B0 (n_10321), .Y(n_4582));
NAND4X1 g60987(.A (n_4242), .B (n_4241), .C (n_9558), .D (n_16), .Y(n_4243));
NOR2X1 g65269(.A (g2819), .B (n_3868), .Y (n_4239));
NOR2X1 g65272(.A (g2807), .B (n_3868), .Y (n_4238));
NOR2X1 g65273(.A (g2775), .B (n_3868), .Y (n_4237));
NAND2X1 g65298(.A (g_13901), .B (n_9717), .Y (n_5573));
NOR2X1 g65350(.A (g2787), .B (n_3868), .Y (n_4235));
OAI22X1 g60989(.A0 (n_3692), .A1 (n_9193), .B0 (n_2474), .B1(n_9992), .Y (n_4233));
CLKBUFX1 gbuf_d_704(.A(n_3808), .Y(d_out_704));
CLKBUFX1 gbuf_q_704(.A(q_in_704), .Y(g5016));
MX2X1 g65433(.A (g2787), .B (g2783), .S0 (n_4231), .Y (n_4232));
MX2X1 g65436(.A (g2819), .B (g2815), .S0 (n_4231), .Y (n_4230));
AOI21X1 g60990(.A0 (n_2773), .A1 (n_3849), .B0 (n_3861), .Y(n_11220));
NAND3X1 g61959(.A (n_2520), .B (n_3652), .C (n_3717), .Y (n_4227));
MX2X1 g60991(.A (g1333), .B (n_3629), .S0 (n_9091), .Y (n_4226));
MX2X1 g65491(.A (g2079), .B (g1945), .S0 (n_4231), .Y (n_4225));
MX2X1 g65492(.A (g2638), .B (g2504), .S0 (n_4231), .Y (n_4224));
NAND2X1 g65934(.A (g2370), .B (n_3679), .Y (n_4223));
AND2X1 g63194(.A (n_3828), .B (n_1285), .Y (n_11079));
NOR2X1 g61451(.A (n_6953), .B (n_4220), .Y (n_4221));
NOR2X1 g61452(.A (n_6954), .B (n_4218), .Y (n_4219));
NOR2X1 g61455(.A (n_6954), .B (n_4216), .Y (n_4217));
NOR2X1 g61456(.A (n_6954), .B (n_4214), .Y (n_4215));
NAND2X1 g63224(.A (n_3821), .B (n_1576), .Y (n_4213));
NOR2X1 g61458(.A (n_11039), .B (n_4211), .Y (n_4212));
NOR2X1 g61459(.A (n_11040), .B (n_4209), .Y (n_4210));
NOR2X1 g61460(.A (n_11040), .B (n_4207), .Y (n_4208));
NOR2X1 g63235(.A (n_3817), .B (n_2163), .Y (n_4206));
NAND3X1 g63236(.A (n_3826), .B (n_2988), .C (n_2423), .Y (n_4205));
NOR2X1 g61461(.A (n_11040), .B (n_4203), .Y (n_4204));
CLKBUFX1 gbuf_d_705(.A(n_3795), .Y(d_out_705));
CLKBUFX1 gbuf_q_705(.A(q_in_705), .Y(g7916));
INVX1 g63267(.A (n_4202), .Y (n_4541));
NAND3X1 g62104(.A (n_2798), .B (n_3564), .C (n_3683), .Y (n_4201));
CLKBUFX1 gbuf_d_706(.A(n_3766), .Y(d_out_706));
CLKBUFX1 gbuf_qn_706(.A(qn_in_706), .Y(g2917));
MX2X1 g63347(.A (g5029), .B (n_3637), .S0 (n_9797), .Y (n_4200));
MX2X1 g63354(.A (g5352), .B (n_3631), .S0 (n_8955), .Y (n_4199));
MX2X1 g63355(.A (g5698), .B (n_3633), .S0 (n_9240), .Y (n_4198));
MX2X1 g63356(.A (g6044), .B (n_3634), .S0 (n_9234), .Y (n_4196));
MX2X1 g63357(.A (g6390), .B (n_3627), .S0 (n_9834), .Y (n_4194));
MX2X1 g63362(.A (g6736), .B (n_3549), .S0 (n_9750), .Y (n_4193));
CLKBUFX1 gbuf_d_707(.A(n_3771), .Y(d_out_707));
CLKBUFX1 gbuf_qn_707(.A(qn_in_707), .Y(g5073));
NOR2X1 g63430(.A (n_717), .B (n_10874), .Y (n_4192));
NOR2X1 g63442(.A (n_855), .B (n_7025), .Y (n_4189));
NAND2X1 g63443(.A (n_4187), .B (n_10920), .Y (n_4188));
NOR2X1 g63444(.A (n_872), .B (n_10920), .Y (n_4186));
NAND2X1 g63445(.A (n_1514), .B (n_7102), .Y (n_4185));
NAND2X1 g63446(.A (n_4183), .B (n_7102), .Y (n_4184));
NOR2X1 g63447(.A (n_863), .B (n_7102), .Y (n_4182));
NAND2X1 g63448(.A (n_1687), .B (n_10920), .Y (n_4181));
AOI21X1 g61018(.A0 (n_3459), .A1 (n_2177), .B0 (n_3811), .Y (n_4180));
NAND2X1 g63449(.A (n_1676), .B (n_8628), .Y (n_4179));
NOR2X1 g63450(.A (n_847), .B (n_8628), .Y (n_4178));
NAND2X1 g63452(.A (n_1670), .B (n_8633), .Y (n_4177));
NOR2X1 g63456(.A (n_715), .B (n_8633), .Y (n_4176));
NAND2X1 g63458(.A (n_1505), .B (n_10874), .Y (n_4175));
NAND2X1 g63459(.A (n_1665), .B (n_7025), .Y (n_4174));
NOR2X1 g63463(.A (n_857), .B (n_10901), .Y (n_4173));
NAND2X1 g63465(.A (n_10901), .B (n_6027), .Y (n_4172));
INVX1 g63498(.A (n_4170), .Y (n_4171));
AOI21X1 g63502(.A0 (n_10672), .A1 (n_4038), .B0 (g2287), .Y (n_4169));
AOI21X1 g63506(.A0 (n_10854), .A1 (n_3939), .B0 (g2421), .Y (n_4168));
NAND2X1 g63510(.A (n_1509), .B (n_10901), .Y (n_4167));
AOI22X1 g63546(.A0 (n_639), .A1 (n_10473), .B0 (n_10472), .B1(g5831), .Y (n_4165));
CLKBUFX1 gbuf_d_708(.A(n_3877), .Y(d_out_708));
CLKBUFX1 gbuf_qn_708(.A(qn_in_708), .Y(g2882));
MX2X1 g63574(.A (g5475), .B (n_94), .S0 (n_10342), .Y (n_4163));
MX2X1 g63582(.A (g5821), .B (n_65), .S0 (n_10472), .Y (n_4161));
MX2X1 g63589(.A (g6167), .B (n_125), .S0 (n_10444), .Y (n_4160));
AOI21X1 g63634(.A0 (n_3616), .A1 (n_9903), .B0 (n_3803), .Y (n_4159));
AOI21X1 g63635(.A0 (n_3611), .A1 (n_9903), .B0 (n_3802), .Y (n_4157));
AOI21X1 g63636(.A0 (n_3589), .A1 (n_9019), .B0 (n_3801), .Y (n_4156));
OAI21X1 g62260(.A0 (n_3447), .A1 (g_15381), .B0 (n_3448), .Y(n_4155));
AOI21X1 g63647(.A0 (g5041), .A1 (n_9856), .B0 (n_3800), .Y (n_4154));
OAI21X1 g62274(.A0 (n_3715), .A1 (n_3569), .B0 (n_3242), .Y (n_4152));
AOI21X1 g61213(.A0 (n_10289), .A1 (n_4149), .B0 (n_10285), .Y(n_4151));
AOI21X1 g61214(.A0 (n_6951), .A1 (n_4149), .B0 (n_3873), .Y (n_4150));
OAI22X1 g62293(.A0 (n_4939), .A1 (n_3686), .B0 (n_10496), .B1(n_9466), .Y (n_4148));
MX2X1 g63770(.A (g1906), .B (g1862), .S0 (n_6677), .Y (n_4147));
MX2X1 g63771(.A (g1936), .B (g1906), .S0 (n_6677), .Y (n_4145));
MX2X1 g63775(.A (g1772), .B (g1728), .S0 (n_10916), .Y (n_4142));
MX2X1 g63776(.A (n_4139), .B (g1772), .S0 (n_10913), .Y (n_4140));
MX2X1 g63777(.A (g_17934), .B (n_3572), .S0 (n_10005), .Y (n_4137));
MX2X1 g62324(.A (n_10818), .B (n_3708), .S0 (n_9240), .Y (n_4136));
OAI22X1 g63781(.A0 (n_3570), .A1 (n_9976), .B0 (g_22639), .B1(n_9830), .Y (n_4135));
XOR2X1 g61225(.A (g_11413), .B (n_4134), .Y (n_4765));
XOR2X1 g61226(.A (g_16456), .B (n_4134), .Y (n_4762));
XOR2X1 g61227(.A (g_20563), .B (n_4134), .Y (n_4758));
XOR2X1 g61228(.A (g_18869), .B (n_4134), .Y (n_4755));
CLKBUFX1 gbuf_d_709(.A(g13881), .Y(d_out_709));
CLKBUFX1 gbuf_q_709(.A(q_in_709), .Y(g16722));
CLKBUFX1 gbuf_d_710(.A(g13865), .Y(d_out_710));
CLKBUFX1 gbuf_q_710(.A(q_in_710), .Y(g16686));
NAND3X1 g63919(.A (n_10912), .B (g1816), .C (n_9698), .Y (n_4133));
NAND3X1 g63928(.A (n_6685), .B (g1950), .C (n_9448), .Y (n_4131));
OR2X1 g63946(.A (n_11094), .B (g_15691), .Y (n_4126));
NOR2X1 g63948(.A (n_4124), .B (n_10674), .Y (n_4125));
NOR2X1 g63954(.A (n_4122), .B (n_10856), .Y (n_4123));
NAND2X1 g63955(.A (n_4108), .B (n_4120), .Y (n_4121));
NOR2X1 g63965(.A (n_6666), .B (n_4118), .Y (n_4119));
NOR2X1 g63975(.A (n_618), .B (n_6666), .Y (n_4117));
NOR2X1 g63977(.A (n_342), .B (n_6666), .Y (n_4113));
NOR2X1 g63978(.A (n_624), .B (n_6666), .Y (n_4111));
NAND3X1 g63999(.A (n_3567), .B (n_2256), .C (n_3551), .Y (n_4110));
OR2X1 g64006(.A (n_10380), .B (n_4109), .Y (n_4583));
CLKBUFX1 gbuf_d_711(.A(n_3798), .Y(d_out_711));
CLKBUFX1 gbuf_q_711(.A(q_in_711), .Y(g4311));
NAND3X1 g64018(.A (n_4108), .B (g1592), .C (n_347), .Y (n_4742));
NAND3X1 g64019(.A (n_4108), .B (g1636), .C (n_629), .Y (n_4740));
NAND3X1 g64020(.A (n_4108), .B (g1592), .C (n_4120), .Y (n_4738));
NAND2X1 g64023(.A (n_4108), .B (g25259), .Y (n_4736));
CLKBUFX1 gbuf_d_712(.A(n_3840), .Y(d_out_712));
CLKBUFX1 gbuf_q_712(.A(q_in_712), .Y(n_8800));
CLKBUFX1 gbuf_d_713(.A(n_3810), .Y(d_out_713));
CLKBUFX1 gbuf_q_713(.A(q_in_713), .Y(n_8915));
CLKBUFX1 gbuf_d_714(.A(n_3738), .Y(d_out_714));
CLKBUFX1 gbuf_q_714(.A(q_in_714), .Y(g4991));
NAND4X1 g64038(.A (g3574), .B (n_10893), .C (g16924), .D (n_6973), .Y(n_4107));
AOI21X1 g64041(.A0 (n_6978), .A1 (n_9019), .B0 (n_3744), .Y (n_4105));
AOI21X1 g64044(.A0 (g4054), .A1 (n_9772), .B0 (n_3742), .Y (n_4103));
AOI21X1 g64045(.A0 (n_7003), .A1 (n_9836), .B0 (n_3746), .Y (n_4102));
NAND4X1 g64049(.A (g3566), .B (n_10895), .C (g16924), .D (n_11128),.Y (n_4101));
CLKBUFX1 gbuf_d_715(.A(n_3886), .Y(d_out_715));
CLKBUFX1 gbuf_q_715(.A(q_in_715), .Y(n_10649));
CLKBUFX1 gbuf_d_716(.A(n_3839), .Y(d_out_716));
CLKBUFX1 gbuf_qn_716(.A(qn_in_716), .Y(g2898));
CLKBUFX1 gbuf_d_717(.A(n_3859), .Y(d_out_717));
CLKBUFX1 gbuf_q_717(.A(q_in_717), .Y(g20899));
CLKBUFX1 gbuf_d_718(.A(n_3807), .Y(d_out_718));
CLKBUFX1 gbuf_q_718(.A(q_in_718), .Y(g2999));
CLKBUFX1 gbuf_d_719(.A(n_3767), .Y(d_out_719));
CLKBUFX1 gbuf_q_719(.A(q_in_719), .Y(g9019));
CLKBUFX1 gbuf_d_720(.A(n_3793), .Y(d_out_720));
CLKBUFX1 gbuf_q_720(.A(q_in_720), .Y(g5037));
CLKBUFX1 gbuf_d_721(.A(n_3869), .Y(d_out_721));
CLKBUFX1 gbuf_q_721(.A(q_in_721), .Y(n_10656));
CLKBUFX1 gbuf_d_722(.A(g16955), .Y(d_out_722));
CLKBUFX1 gbuf_q_722(.A(q_in_722), .Y(g13906));
OR2X1 g64141(.A (g3808), .B (n_4096), .Y (n_6049));
NAND4X1 g64216(.A (g3901), .B (n_6787), .C (g14518), .D (n_3894), .Y(n_4098));
NAND2X1 g64223(.A (n_11208), .B (n_4096), .Y (n_4885));
INVX1 g62564(.A (n_6551), .Y (n_4671));
NAND3X1 g61737(.A (n_3891), .B (n_10184), .C (n_4091), .Y (n_4092));
NAND3X1 g61738(.A (n_3893), .B (n_10205), .C (n_4091), .Y (n_4090));
NAND4X1 g64378(.A (n_4988), .B (g3889), .C (g14518), .D (n_5402), .Y(n_4088));
AOI21X1 g64398(.A0 (n_3897), .A1 (n_245), .B0 (n_3898), .Y (n_4087));
AOI21X1 g64399(.A0 (n_3730), .A1 (n_282), .B0 (n_3731), .Y (n_4086));
AOI21X1 g64400(.A0 (n_3728), .A1 (n_360), .B0 (n_3729), .Y (n_4085));
AOI21X1 g64401(.A0 (n_3726), .A1 (n_3135), .B0 (n_3727), .Y (n_4084));
OAI21X1 g62662(.A0 (n_3514), .A1 (n_9371), .B0 (n_3881), .Y (n_4083));
AOI22X1 g62666(.A0 (n_3691), .A1 (n_3857), .B0 (g_13278), .B1(n_9129), .Y (n_4082));
OAI22X1 g62677(.A0 (n_3648), .A1 (n_3797), .B0 (n_327), .B1(n_10005), .Y (n_4081));
CLKBUFX1 gbuf_d_723(.A(g14217), .Y(d_out_723));
CLKBUFX1 gbuf_q_723(.A(q_in_723), .Y(g14096));
NAND4X1 g64524(.A (g5109), .B (n_9627), .C (g9497), .D (n_107), .Y(n_4080));
XOR2X1 g61080(.A (g1478), .B (n_11025), .Y (n_4638));
XOR2X1 g61081(.A (g1448), .B (n_11026), .Y (n_4633));
XOR2X1 g61082(.A (g1472), .B (n_11026), .Y (n_4629));
NAND4X1 g64711(.A (g5456), .B (n_9627), .C (g9555), .D (g_5508), .Y(n_4076));
NAND4X1 g64720(.A (g6148), .B (n_9627), .C (g9682), .D (g_14965), .Y(n_4074));
NAND4X1 g64722(.A (g6494), .B (n_9627), .C (g9743), .D (g_3861), .Y(n_4073));
NAND4X1 g64726(.A (g3100), .B (n_9627), .C (g8215), .D (g_6579), .Y(n_4072));
NAND4X1 g64729(.A (g3802), .B (n_9627), .C (g8344), .D (g_5156), .Y(n_4071));
NAND3X1 g60973(.A (n_10429), .B (g1367), .C (n_9717), .Y (n_4070));
NOR2X1 g62791(.A (n_3685), .B (n_9775), .Y (n_4069));
AOI21X1 g62799(.A0 (n_1349), .A1 (n_2471), .B0 (n_3680), .Y (n_4068));
CLKBUFX1 gbuf_d_724(.A(n_3703), .Y(d_out_724));
CLKBUFX1 gbuf_q_724(.A(q_in_724), .Y(n_8509));
NAND2X1 g62826(.A (n_3681), .B (n_3822), .Y (n_4067));
NOR2X1 g64854(.A (n_3697), .B (n_8557), .Y (n_5703));
OR2X1 g64861(.A (g3100), .B (n_9398), .Y (n_4066));
OR2X1 g64866(.A (g6148), .B (n_9398), .Y (n_4065));
OR2X1 g64874(.A (g3451), .B (n_10687), .Y (n_4062));
OR2X1 g64880(.A (g3802), .B (n_9091), .Y (n_4060));
AOI22X1 g64037(.A0 (n_2018), .A1 (n_3547), .B0 (n_523), .B1 (n_9693),.Y (n_4059));
NOR2X1 g64896(.A (n_3695), .B (n_8557), .Y (n_5701));
OR2X1 g64911(.A (g6494), .B (n_9398), .Y (n_4056));
OR2X1 g64913(.A (g5802), .B (n_9398), .Y (n_4055));
OR4X1 g62899(.A (n_11080), .B (n_4053), .C (n_9856), .D (g_22306), .Y(n_4054));
XOR2X1 g62928(.A (g4593), .B (n_10395), .Y (n_4050));
AOI21X1 g65011(.A0 (g4473), .A1 (n_2861), .B0 (g4459), .Y (n_4049));
MX2X1 g62938(.A (g2848), .B (n_3500), .S0 (n_8955), .Y (n_4048));
NAND4X1 g65041(.A (g5112), .B (n_9521), .C (g_11037), .D (g9553), .Y(n_4046));
AOI21X1 g65051(.A0 (g4164), .A1 (g4253), .B0 (n_3701), .Y (n_4247));
CLKBUFX1 gbuf_d_725(.A(g4456), .Y(d_out_725));
CLKBUFX1 gbuf_qn_725(.A(qn_in_725), .Y(g4455));
CLKBUFX1 gbuf_d_726(.A(g12184), .Y(d_out_726));
CLKBUFX1 gbuf_q_726(.A(q_in_726), .Y(g_17653));
NAND2X1 g61916(.A (n_4045), .B (g_14342), .Y (n_4578));
CLKBUFX1 gbuf_d_727(.A(n_3671), .Y(d_out_727));
CLKBUFX1 gbuf_q_727(.A(q_in_727), .Y(g_12433));
AND2X1 g65267(.A (n_11012), .B (n_10078), .Y (n_4044));
NOR2X1 g65289(.A (g2815), .B (g2724), .Y (n_4043));
NOR2X1 g65297(.A (g2783), .B (g2724), .Y (n_4042));
AOI22X1 g64033(.A0 (n_2007), .A1 (n_10948), .B0 (n_10660), .B1(n_10078), .Y (n_4040));
NAND3X1 g64010(.A (n_10672), .B (n_4038), .C (g2287), .Y (n_4281));
CLKBUFX1 gbuf_d_728(.A(n_3723), .Y(d_out_728));
CLKBUFX1 gbuf_q_728(.A(q_in_728), .Y(g_14843));
NOR2X1 g65747(.A (n_4231), .B (g2775), .Y (n_4037));
NAND2X1 g65781(.A (g1677), .B (n_4231), .Y (n_4035));
NAND2X1 g65853(.A (n_4231), .B (n_9952), .Y (n_4034));
NOR2X1 g65923(.A (g2715), .B (g2807), .Y (n_4033));
NAND2X1 g65936(.A (g2236), .B (n_4231), .Y (n_4032));
INVX1 g61003(.A (n_4030), .Y (n_4031));
OAI21X1 g63193(.A0 (n_3479), .A1 (g4153), .B0 (n_9627), .Y (n_4029));
NAND3X1 g63209(.A (n_11080), .B (g_22306), .C (n_9698), .Y (n_4028));
NAND3X1 g63210(.A (n_4024), .B (n_3660), .C (n_9651), .Y (n_4025));
NAND2X1 g63225(.A (n_3656), .B (n_1434), .Y (n_4022));
NOR2X1 g63227(.A (g5694), .B (n_10660), .Y (n_4021));
NOR2X1 g63229(.A (g6040), .B (n_11201), .Y (n_4020));
NOR2X1 g63230(.A (g6386), .B (g6395), .Y (n_4019));
NOR2X1 g63237(.A (g6732), .B (n_523), .Y (n_4018));
NOR2X1 g61007(.A (n_3778), .B (n_2172), .Y (n_4017));
AND2X1 g63247(.A (n_3172), .B (g5348), .Y (n_4016));
NOR2X1 g63251(.A (n_2882), .B (g5694), .Y (n_4015));
NOR2X1 g63253(.A (n_2613), .B (g6040), .Y (n_4014));
OAI21X1 g63255(.A0 (n_2150), .A1 (n_9978), .B0 (n_3653), .Y (n_4013));
NOR2X1 g63257(.A (n_2607), .B (g6386), .Y (n_4012));
NOR2X1 g63259(.A (n_2872), .B (g6732), .Y (n_4011));
AOI21X1 g63268(.A0 (n_2987), .A1 (n_286), .B0 (n_11081), .Y (n_4202));
CLKBUFX1 gbuf_d_729(.A(n_3647), .Y(d_out_729));
CLKBUFX1 gbuf_q_729(.A(q_in_729), .Y(g17320));
CLKBUFX1 gbuf_d_730(.A(n_3666), .Y(d_out_730));
CLKBUFX1 gbuf_q_730(.A(q_in_730), .Y(g1384));
OAI22X1 g63327(.A0 (n_4939), .A1 (n_3432), .B0 (n_2583), .B1(n_9627), .Y (n_4010));
MX2X1 g63346(.A (g4172), .B (n_3480), .S0 (n_9091), .Y (n_4009));
MX2X1 g63365(.A (g_15287), .B (n_3521), .S0 (n_9359), .Y (n_4008));
CLKBUFX1 gbuf_d_731(.A(n_3636), .Y(d_out_731));
CLKBUFX1 gbuf_q_731(.A(q_in_731), .Y(g18881));
AOI21X1 g63470(.A0 (n_10915), .A1 (n_3789), .B0 (g1728), .Y (n_4006));
NAND3X1 g63473(.A (n_1097), .B (n_10347), .C (n_10063), .Y (n_4005));
NAND3X1 g63478(.A (n_1098), .B (n_10473), .C (n_9209), .Y (n_4002));
NAND3X1 g63481(.A (n_1269), .B (n_10445), .C (n_9359), .Y (n_4000));
AOI21X1 g63483(.A0 (n_6676), .A1 (n_3782), .B0 (g1862), .Y (n_3998));
NAND3X1 g63485(.A (n_1099), .B (n_3455), .C (n_10385), .Y (n_3997));
NAND3X1 g63488(.A (n_3640), .B (n_1285), .C (n_11056), .Y (n_4805));
NAND2X1 g63499(.A (g4423), .B (n_10385), .Y (n_4170));
NAND2X1 g63505(.A (g4423), .B (n_9952), .Y (n_3996));
AOI22X1 g61021(.A0 (n_3460), .A1 (n_9627), .B0 (n_3372), .B1(n_3459), .Y (n_3995));
AOI22X1 g63542(.A0 (n_540), .A1 (n_7242), .B0 (n_7245), .B1 (g5138),.Y (n_3993));
CLKBUFX1 gbuf_d_732(.A(n_3700), .Y(d_out_732));
CLKBUFX1 gbuf_q_732(.A(q_in_732), .Y(g_22034));
AOI22X1 g63549(.A0 (n_600), .A1 (n_3455), .B0 (n_3814), .B1 (g6523),.Y (n_3992));
OAI22X1 g63555(.A0 (n_2748), .A1 (n_9193), .B0 (n_3410), .B1(n_9627), .Y (n_3991));
NAND4X1 g63557(.A (n_2145), .B (n_2144), .C (n_3269), .D (n_2332), .Y(n_3990));
NAND4X1 g63566(.A (n_2128), .B (n_2126), .C (n_3266), .D (n_2029), .Y(n_11189));
NAND4X1 g63569(.A (n_7018), .B (n_3984), .C (g5052), .D (n_10697), .Y(n_3985));
MX2X1 g63570(.A (g5128), .B (n_168), .S0 (n_7245), .Y (n_3983));
AOI21X1 g63633(.A0 (n_3618), .A1 (n_9193), .B0 (n_3642), .Y (n_3982));
MX2X1 g63648(.A (n_10813), .B (n_3449), .S0 (n_8955), .Y (n_3981));
OAI21X1 g62267(.A0 (n_3537), .A1 (n_9599), .B0 (n_3709), .Y (n_3979));
AOI21X1 g61215(.A0 (n_11211), .A1 (g1589), .B0 (n_3870), .Y (n_3978));
AOI21X1 g61220(.A0 (n_10763), .A1 (g1589), .B0 (n_10762), .Y(n_3977));
XOR2X1 g63763(.A (n_3011), .B (n_10347), .Y (n_3974));
XOR2X1 g63764(.A (n_2684), .B (n_10473), .Y (n_3973));
XOR2X1 g63765(.A (n_2704), .B (n_10445), .Y (n_3972));
XOR2X1 g63768(.A (n_3007), .B (n_3455), .Y (n_3971));
NAND3X1 g61037(.A (n_3369), .B (n_2555), .C (n_3523), .Y (n_3970));
MX2X1 g61223(.A (g1589), .B (n_649), .S0 (n_8955), .Y (n_3969));
MX2X1 g63791(.A (n_1285), .B (n_3429), .S0 (n_8955), .Y (n_3968));
MX2X1 g63792(.A (g_17065), .B (n_3424), .S0 (n_8955), .Y (n_3966));
MX2X1 g63793(.A (n_3550), .B (n_3423), .S0 (n_9156), .Y (n_3964));
MX2X1 g63797(.A (g_19113), .B (n_3422), .S0 (n_9091), .Y (n_3963));
MX2X1 g63799(.A (g_16677), .B (n_3420), .S0 (n_9000), .Y (n_3962));
MX2X1 g63800(.A (g_21720), .B (n_3418), .S0 (n_9000), .Y (n_3960));
MX2X1 g63801(.A (g_13758), .B (n_3417), .S0 (n_9000), .Y (n_3959));
MX2X1 g63802(.A (g_19289), .B (n_3416), .S0 (n_9311), .Y (n_3958));
MX2X1 g63807(.A (g_21778), .B (n_3415), .S0 (n_9797), .Y (n_3957));
INVX1 g63880(.A (n_7025), .Y (n_3956));
OR2X1 g63882(.A (n_3615), .B (n_9775), .Y (n_3955));
INVX1 g63887(.A (n_7102), .Y (n_3953));
INVX1 g63890(.A (n_8628), .Y (n_3952));
INVX1 g63897(.A (n_8633), .Y (n_3951));
NOR2X1 g63915(.A (n_3948), .B (n_10917), .Y (n_3949));
NAND2X1 g63925(.A (n_4424), .B (n_9358), .Y (n_5007));
NOR2X1 g63938(.A (n_3557), .B (n_9193), .Y (n_3947));
NOR2X1 g63956(.A (n_3574), .B (n_3945), .Y (n_3946));
NOR3X1 g63972(.A (n_6752), .B (n_3943), .C (g2070), .Y (n_3944));
NAND4X1 g63983(.A (n_3561), .B (n_2918), .C (n_10063), .D (n_3065),.Y (n_3942));
NAND4X1 g63994(.A (n_3560), .B (n_2917), .C (n_9750), .D (n_3062), .Y(n_3941));
CLKBUFX1 gbuf_d_733(.A(n_3689), .Y(d_out_733));
CLKBUFX1 gbuf_q_733(.A(q_in_733), .Y(g1345));
NAND3X1 g64011(.A (n_10672), .B (g2331), .C (n_386), .Y (n_4279));
NAND3X1 g64012(.A (n_10675), .B (g2361), .C (g2287), .Y (n_4277));
NAND3X1 g64013(.A (n_10672), .B (n_4038), .C (g2361), .Y (n_4275));
NAND3X1 g64014(.A (n_10854), .B (n_3939), .C (g2421), .Y (n_4273));
NAND3X1 g64015(.A (n_10854), .B (g2465), .C (n_437), .Y (n_4271));
NAND3X1 g64016(.A (n_10857), .B (n_4339), .C (g2421), .Y (n_4269));
NAND3X1 g64017(.A (n_10854), .B (n_3939), .C (n_4339), .Y (n_4267));
CLKBUFX1 gbuf_d_734(.A(n_3673), .Y(d_out_734));
CLKBUFX1 gbuf_q_734(.A(q_in_734), .Y(g_20073));
CLKBUFX1 gbuf_d_735(.A(n_3585), .Y(d_out_735));
CLKBUFX1 gbuf_q_735(.A(q_in_735), .Y(g_20563));
CLKBUFX1 gbuf_d_736(.A(n_3620), .Y(d_out_736));
CLKBUFX1 gbuf_q_736(.A(q_in_736), .Y(g4669));
OR2X1 g64022(.A (n_3938), .B (n_5471), .Y (n_4539));
CLKBUFX1 gbuf_d_737(.A(n_3725), .Y(d_out_737));
CLKBUFX1 gbuf_q_737(.A(q_in_737), .Y(n_11216));
AOI22X1 g64032(.A0 (n_2588), .A1 (n_3399), .B0 (n_8806), .B1(n_9193), .Y (n_3937));
AOI22X1 g64036(.A0 (n_2015), .A1 (n_3626), .B0 (g6395), .B1(n_10078), .Y (n_3936));
CLKBUFX1 gbuf_d_738(.A(n_3721), .Y(d_out_738));
CLKBUFX1 gbuf_q_738(.A(q_in_738), .Y(g4793));
CLKBUFX1 gbuf_d_739(.A(n_3675), .Y(d_out_739));
CLKBUFX1 gbuf_q_739(.A(q_in_739), .Y(g_18795));
CLKBUFX1 gbuf_d_740(.A(n_3674), .Y(d_out_740));
CLKBUFX1 gbuf_q_740(.A(q_in_740), .Y(g_22038));
CLKBUFX1 gbuf_d_741(.A(n_3670), .Y(d_out_741));
CLKBUFX1 gbuf_q_741(.A(q_in_741), .Y(g_17934));
CLKBUFX1 gbuf_d_742(.A(n_3672), .Y(d_out_742));
CLKBUFX1 gbuf_q_742(.A(q_in_742), .Y(g_18238));
CLKBUFX1 gbuf_d_743(.A(n_3688), .Y(d_out_743));
CLKBUFX1 gbuf_q_743(.A(q_in_743), .Y(g4983));
CLKBUFX1 gbuf_d_744(.A(n_3662), .Y(d_out_744));
CLKBUFX1 gbuf_q_744(.A(q_in_744), .Y(g_19911));
CLKBUFX1 gbuf_d_745(.A(n_3655), .Y(d_out_745));
CLKBUFX1 gbuf_q_745(.A(q_in_745), .Y(g4633));
CLKBUFX1 gbuf_d_746(.A(n_3638), .Y(d_out_746));
CLKBUFX1 gbuf_q_746(.A(q_in_746), .Y(g_18739));
CLKBUFX1 gbuf_d_747(.A(n_3622), .Y(d_out_747));
CLKBUFX1 gbuf_q_747(.A(q_in_747), .Y(g4888));
CLKBUFX1 gbuf_d_748(.A(n_3621), .Y(d_out_748));
CLKBUFX1 gbuf_q_748(.A(q_in_748), .Y(g_19789));
OAI21X1 g64072(.A0 (n_3779), .A1 (n_6978), .B0 (n_3598), .Y (n_3934));
CLKBUFX1 gbuf_d_749(.A(n_3555), .Y(d_out_749));
CLKBUFX1 gbuf_q_749(.A(q_in_749), .Y(g_5029));
CLKBUFX1 gbuf_d_750(.A(n_3591), .Y(d_out_750));
CLKBUFX1 gbuf_q_750(.A(q_in_750), .Y(g1448));
CLKBUFX1 gbuf_d_751(.A(n_3577), .Y(d_out_751));
CLKBUFX1 gbuf_q_751(.A(q_in_751), .Y(g5029));
CLKBUFX1 gbuf_d_752(.A(n_3554), .Y(d_out_752));
CLKBUFX1 gbuf_q_752(.A(q_in_752), .Y(g_18996));
CLKBUFX1 gbuf_d_753(.A(n_3722), .Y(d_out_753));
CLKBUFX1 gbuf_q_753(.A(q_in_753), .Y(g34034));
CLKBUFX1 gbuf_d_754(.A(n_3552), .Y(d_out_754));
CLKBUFX1 gbuf_q_754(.A(q_in_754), .Y(g_22021));
CLKBUFX1 gbuf_d_755(.A(n_3724), .Y(d_out_755));
CLKBUFX1 gbuf_q_755(.A(q_in_755), .Y(g2975));
CLKBUFX1 gbuf_d_756(.A(n_3546), .Y(d_out_756));
CLKBUFX1 gbuf_q_756(.A(q_in_756), .Y(g4621));
CLKBUFX1 gbuf_d_757(.A(n_3712), .Y(d_out_757));
CLKBUFX1 gbuf_q_757(.A(q_in_757), .Y(g5535));
CLKBUFX1 gbuf_d_758(.A(n_3711), .Y(d_out_758));
CLKBUFX1 gbuf_q_758(.A(q_in_758), .Y(g6573));
CLKBUFX1 gbuf_d_759(.A(n_3710), .Y(d_out_759));
CLKBUFX1 gbuf_q_759(.A(q_in_759), .Y(g3530));
OAI21X1 g64080(.A0 (n_3775), .A1 (n_7003), .B0 (n_3592), .Y (n_3933));
NAND2X1 g60954(.A (n_3658), .B (n_3716), .Y (n_3932));
INVX1 g64177(.A (n_10944), .Y (n_3929));
INVX2 g64187(.A (n_6759), .Y (n_4304));
INVX2 g64199(.A (n_3925), .Y (n_4668));
INVX1 g64240(.A (n_4447), .Y (n_3922));
OAI21X1 g62599(.A0 (n_3915), .A1 (n_3914), .B0 (n_3913), .Y (n_3916));
INVX1 g64330(.A (n_10380), .Y (n_4299));
OR4X1 g60959(.A (n_10429), .B (n_3910), .C (n_9856), .D (g1367), .Y(n_3911));
OAI21X1 g64397(.A0 (g16693), .A1 (g14518), .B0 (n_3535), .Y (n_3907));
AOI21X1 g62650(.A0 (n_3718), .A1 (n_28), .B0 (n_11032), .Y (n_3906));
MX2X1 g64408(.A (g_21318), .B (g14201), .S0 (n_5582), .Y (n_3905));
NAND4X1 g62673(.A (n_3646), .B (n_6577), .C (n_10687), .D (g4332), .Y(n_3904));
NAND3X1 g64532(.A (g5752), .B (n_9521), .C (g_7062), .Y (n_3903));
NAND3X1 g64582(.A (g3401), .B (n_9521), .C (g_5313), .Y (n_3902));
INVX1 g64596(.A (n_3900), .Y (n_6364));
NAND3X1 g64664(.A (n_3732), .B (g3965), .C (n_8917), .Y (n_11219));
NOR2X1 g64679(.A (n_3897), .B (n_3896), .Y (n_3898));
NAND4X1 g64732(.A (g3905), .B (n_3894), .C (g16693), .D (n_6808), .Y(n_3895));
AOI21X1 g61821(.A0 (n_1885), .A1 (n_2845), .B0 (n_3775), .Y (n_3893));
AOI21X1 g61822(.A0 (n_1884), .A1 (n_2844), .B0 (n_3779), .Y (n_3891));
CLKBUFX1 gbuf_d_760(.A(g14201), .Y(d_out_760));
CLKBUFX1 gbuf_q_760(.A(q_in_760), .Y(g14217));
NAND2X1 g62833(.A (n_3321), .B (n_3516), .Y (n_3886));
INVX1 g62837(.A (n_11031), .Y (n_3885));
OR2X1 g64855(.A (g5456), .B (n_9091), .Y (n_3883));
NAND3X1 g64930(.A (n_6967), .B (n_9553), .C (g_11037), .Y (n_3882));
AOI22X1 g62909(.A0 (n_3331), .A1 (n_10184), .B0 (n_11134), .B1(n_9107), .Y (n_3881));
AOI22X1 g65024(.A0 (g2960), .A1 (n_3356), .B0 (g2970), .B1 (g2975),.Y (n_3879));
AOI22X1 g65032(.A0 (g2922), .A1 (n_3357), .B0 (g2912), .B1 (n_3463),.Y (n_3878));
MX2X1 g62940(.A (n_3501), .B (n_3330), .S0 (n_9167), .Y (n_3877));
CLKBUFX1 gbuf_d_761(.A(n_3407), .Y(d_out_761));
CLKBUFX1 gbuf_q_761(.A(q_in_761), .Y(g1395));
CLKBUFX1 gbuf_d_762(.A(n_3412), .Y(d_out_762));
CLKBUFX1 gbuf_q_762(.A(q_in_762), .Y(g4659));
CLKBUFX1 gbuf_d_763(.A(g9497), .Y(d_out_763));
CLKBUFX1 gbuf_qn_763(.A(qn_in_763), .Y(g5109));
NAND2X1 g65266(.A (n_3868), .B (n_9019), .Y (n_3869));
CLKBUFX1 gbuf_d_764(.A(n_3414), .Y(d_out_764));
CLKBUFX1 gbuf_q_764(.A(q_in_764), .Y(n_1627));
NOR2X1 g65336(.A (n_10650), .B (n_3868), .Y (n_3866));
NAND2X1 g65810(.A (g1811), .B (n_3679), .Y (n_3863));
CLKBUFX1 gbuf_d_765(.A(n_3494), .Y(d_out_765));
CLKBUFX1 gbuf_qn_765(.A(qn_in_765), .Y(g4366));
INVX1 g61439(.A (g1246), .Y (n_4558));
OR2X1 g61004(.A (n_3860), .B (g7946), .Y (n_4030));
NOR2X1 g61005(.A (n_3860), .B (n_10196), .Y (n_3861));
OAI21X1 g63212(.A0 (n_2425), .A1 (n_10115), .B0 (n_3488), .Y(n_3859));
NAND2X1 g63214(.A (n_3517), .B (n_3857), .Y (n_3858));
NOR2X1 g63234(.A (n_8836), .B (n_3855), .Y (n_3856));
NOR2X1 g63240(.A (n_8836), .B (n_8832), .Y (n_3854));
NAND4X1 g63261(.A (n_3050), .B (n_3302), .C (n_3049), .D (n_3032), .Y(n_3852));
NAND4X1 g63271(.A (n_3845), .B (n_10063), .C (n_3844), .D (n_2428),.Y (n_3851));
NOR2X1 g61009(.A (n_3860), .B (n_3849), .Y (n_4284));
NAND3X1 g61010(.A (n_3484), .B (g1361), .C (n_9811), .Y (n_3848));
OAI21X1 g63283(.A0 (n_3894), .A1 (n_9940), .B0 (n_3487), .Y (n_3847));
NAND4X1 g63285(.A (n_3845), .B (n_3844), .C (n_9279), .D (n_40), .Y(n_3846));
CLKBUFX1 gbuf_d_766(.A(n_3468), .Y(d_out_766));
CLKBUFX1 gbuf_q_766(.A(q_in_766), .Y(g4933));
NAND4X1 g63314(.A (n_4832), .B (n_6767), .C (n_9279), .D (n_416), .Y(n_3843));
AOI21X1 g63332(.A0 (g1183), .A1 (n_8837), .B0 (n_3505), .Y (n_3841));
NAND3X1 g62101(.A (n_2278), .B (n_2711), .C (n_3327), .Y (n_3840));
OAI21X1 g63345(.A0 (g2864), .A1 (n_9894), .B0 (n_3503), .Y (n_3839));
AOI21X1 g61499(.A0 (n_3838), .A1 (g1242), .B0 (n_3837), .Y (n_5057));
INVX1 g63374(.A (g5694), .Y (n_3836));
INVX1 g63376(.A (g6040), .Y (n_3835));
INVX1 g63378(.A (g6386), .Y (n_3834));
INVX1 g63380(.A (g6732), .Y (n_3833));
NAND3X1 g63460(.A (n_1101), .B (n_7243), .C (n_9894), .Y (n_3830));
OR2X1 g63487(.A (n_10532), .B (n_3639), .Y (n_3828));
NOR2X1 g63511(.A (n_2755), .B (n_3478), .Y (n_3826));
NAND3X1 g63517(.A (n_10768), .B (n_2638), .C (n_3264), .Y (n_3825));
NAND3X1 g63521(.A (n_3482), .B (g_16958), .C (n_9493), .Y (n_3824));
NAND3X1 g63533(.A (n_3426), .B (n_3822), .C (n_3438), .Y (n_3823));
AOI22X1 g63536(.A0 (n_3260), .A1 (n_8676), .B0 (n_599), .B1 (n_3259),.Y (n_3821));
NAND4X1 g63562(.A (n_6577), .B (n_3645), .C (n_662), .D (n_3213), .Y(n_3819));
NAND4X1 g63564(.A (n_1849), .B (n_3278), .C (n_1858), .D (n_1574), .Y(n_3817));
NAND4X1 g63568(.A (n_10770), .B (n_3984), .C (n_9359), .D (g5046), .Y(n_3816));
MX2X1 g63597(.A (g6513), .B (n_158), .S0 (n_3814), .Y (n_3815));
AOI22X1 g63638(.A0 (n_3604), .A1 (n_9772), .B0 (n_3814), .B1(n_3812), .Y (n_3813));
CLKBUFX1 gbuf_d_767(.A(n_3532), .Y(d_out_767));
CLKBUFX1 gbuf_q_767(.A(q_in_767), .Y(g5881));
AOI21X1 g61033(.A0 (n_3366), .A1 (n_2178), .B0 (n_3459), .Y (n_3811));
OAI22X1 g62298(.A0 (n_3346), .A1 (n_3720), .B0 (n_8637), .B1(n_9830), .Y (n_3810));
XOR2X1 g63762(.A (n_2718), .B (n_7242), .Y (n_3809));
CLKBUFX1 gbuf_d_768(.A(n_3408), .Y(d_out_768));
CLKBUFX1 gbuf_q_768(.A(q_in_768), .Y(g5499));
MX2X1 g63809(.A (n_6967), .B (n_3271), .S0 (n_9234), .Y (n_3808));
AOI21X1 g63883(.A0 (g2932), .A1 (n_27), .B0 (n_9976), .Y (n_3807));
NOR2X1 g63912(.A (n_10347), .B (n_6399), .Y (n_3803));
NOR2X1 g63916(.A (n_10473), .B (n_6398), .Y (n_3802));
NOR2X1 g63920(.A (n_10445), .B (n_6406), .Y (n_3801));
NOR3X1 g63921(.A (n_10078), .B (g5046), .C (n_10770), .Y (n_3800));
NOR2X1 g63939(.A (n_3538), .B (n_3797), .Y (n_3798));
NAND2X1 g63953(.A (n_4843), .B (n_9493), .Y (n_4956));
MX2X1 g61652(.A (g_20614), .B (n_10752), .S0 (n_9750), .Y (n_3795));
NAND2X1 g63966(.A (n_3427), .B (n_3017), .Y (n_3793));
AOI21X1 g63980(.A0 (n_3244), .A1 (n_11037), .B0 (n_10621), .Y(n_3792));
NAND3X1 g63981(.A (n_10915), .B (n_3789), .C (g1728), .Y (n_4220));
NAND3X1 g63982(.A (n_10915), .B (g1772), .C (n_446), .Y (n_4218));
NAND3X1 g63984(.A (n_10915), .B (n_4139), .C (g1728), .Y (n_4216));
AOI21X1 g63985(.A0 (n_10947), .A1 (n_4982), .B0 (n_7150), .Y(n_3788));
AOI21X1 g63986(.A0 (n_3612), .A1 (n_4980), .B0 (n_10506), .Y(n_3786));
AOI21X1 g63987(.A0 (n_3784), .A1 (n_4978), .B0 (n_3277), .Y (n_3785));
NAND3X1 g63988(.A (n_6676), .B (n_3782), .C (g1862), .Y (n_4211));
NAND3X1 g63989(.A (n_6676), .B (g1936), .C (g1862), .Y (n_4207));
AOI21X1 g63990(.A0 (n_3605), .A1 (n_11070), .B0 (n_3275), .Y(n_3781));
NAND3X1 g63991(.A (n_6676), .B (n_3782), .C (g1936), .Y (n_4203));
NAND3X1 g63992(.A (n_6676), .B (g1906), .C (n_328), .Y (n_4209));
AOI21X1 g63993(.A0 (n_3779), .A1 (g3639), .B0 (n_1273), .Y (n_3780));
INVX1 g61047(.A (n_3778), .Y (n_4242));
AOI21X1 g64000(.A0 (n_6243), .A1 (g3990), .B0 (n_6787), .Y (n_3777));
AOI21X1 g64003(.A0 (n_3775), .A1 (n_10834), .B0 (n_8586), .Y(n_3776));
NAND3X1 g64009(.A (n_10915), .B (n_3789), .C (n_4139), .Y (n_4214));
CLKBUFX1 gbuf_d_769(.A(n_3483), .Y(d_out_769));
CLKBUFX1 gbuf_q_769(.A(q_in_769), .Y(g1404));
CLKBUFX1 gbuf_d_770(.A(n_3454), .Y(d_out_770));
CLKBUFX1 gbuf_q_770(.A(q_in_770), .Y(g_16456));
CLKBUFX1 gbuf_d_771(.A(n_3458), .Y(d_out_771));
CLKBUFX1 gbuf_q_771(.A(q_in_771), .Y(g_18869));
CLKBUFX1 gbuf_d_772(.A(n_3520), .Y(d_out_772));
CLKBUFX1 gbuf_q_772(.A(q_in_772), .Y(g4664));
NAND3X1 g64031(.A (n_3440), .B (n_659), .C (n_9398), .Y (n_3774));
CLKBUFX1 gbuf_d_773(.A(n_3508), .Y(d_out_773));
CLKBUFX1 gbuf_q_773(.A(q_in_773), .Y(g1554));
CLKBUFX1 gbuf_d_774(.A(n_3507), .Y(d_out_774));
CLKBUFX1 gbuf_q_774(.A(q_in_774), .Y(g4854));
CLKBUFX1 gbuf_d_775(.A(n_3529), .Y(d_out_775));
CLKBUFX1 gbuf_q_775(.A(q_in_775), .Y(g4849));
CLKBUFX1 gbuf_d_776(.A(n_3512), .Y(d_out_776));
CLKBUFX1 gbuf_qn_776(.A(qn_in_776), .Y(g3343));
CLKBUFX1 gbuf_d_777(.A(n_3511), .Y(d_out_777));
CLKBUFX1 gbuf_qn_777(.A(qn_in_777), .Y(g3694));
MX2X1 g64062(.A (g5069), .B (n_2044), .S0 (n_9448), .Y (n_3771));
CLKBUFX1 gbuf_d_778(.A(n_3496), .Y(d_out_778));
CLKBUFX1 gbuf_q_778(.A(q_in_778), .Y(g_22464));
CLKBUFX1 gbuf_d_779(.A(n_3490), .Y(d_out_779));
CLKBUFX1 gbuf_q_779(.A(q_in_779), .Y(g4653));
CLKBUFX1 gbuf_d_780(.A(n_3481), .Y(d_out_780));
CLKBUFX1 gbuf_q_780(.A(q_in_780), .Y(g4064));
CLKBUFX1 gbuf_d_781(.A(n_3473), .Y(d_out_781));
CLKBUFX1 gbuf_q_781(.A(q_in_781), .Y(g2848));
CLKBUFX1 gbuf_d_782(.A(n_3470), .Y(d_out_782));
CLKBUFX1 gbuf_q_782(.A(q_in_782), .Y(g4743));
CLKBUFX1 gbuf_d_783(.A(n_3469), .Y(d_out_783));
CLKBUFX1 gbuf_q_783(.A(q_in_783), .Y(g4754));
CLKBUFX1 gbuf_d_784(.A(n_3471), .Y(d_out_784));
CLKBUFX1 gbuf_q_784(.A(q_in_784), .Y(g4698));
CLKBUFX1 gbuf_d_785(.A(n_3475), .Y(d_out_785));
CLKBUFX1 gbuf_q_785(.A(q_in_785), .Y(g4843));
CLKBUFX1 gbuf_d_786(.A(n_3510), .Y(d_out_786));
CLKBUFX1 gbuf_q_786(.A(q_in_786), .Y(g4765));
CLKBUFX1 gbuf_d_787(.A(n_3465), .Y(d_out_787));
CLKBUFX1 gbuf_q_787(.A(q_in_787), .Y(g4955));
CLKBUFX1 gbuf_d_788(.A(n_3466), .Y(d_out_788));
CLKBUFX1 gbuf_q_788(.A(q_in_788), .Y(g4944));
CLKBUFX1 gbuf_d_789(.A(n_3437), .Y(d_out_789));
CLKBUFX1 gbuf_q_789(.A(q_in_789), .Y(g_4409));
CLKBUFX1 gbuf_d_790(.A(n_3436), .Y(d_out_790));
CLKBUFX1 gbuf_q_790(.A(q_in_790), .Y(g_3381));
CLKBUFX1 gbuf_d_791(.A(n_3435), .Y(d_out_791));
CLKBUFX1 gbuf_q_791(.A(q_in_791), .Y(n_11050));
CLKBUFX1 gbuf_d_792(.A(n_3434), .Y(d_out_792));
CLKBUFX1 gbuf_q_792(.A(q_in_792), .Y(g_6165));
CLKBUFX1 gbuf_d_793(.A(n_3461), .Y(d_out_793));
CLKBUFX1 gbuf_q_793(.A(q_in_793), .Y(g1300));
CLKBUFX1 gbuf_d_794(.A(n_3433), .Y(d_out_794));
CLKBUFX1 gbuf_q_794(.A(q_in_794), .Y(g_8864));
CLKBUFX1 gbuf_d_795(.A(n_3413), .Y(d_out_795));
CLKBUFX1 gbuf_q_795(.A(q_in_795), .Y(g_10278));
CLKBUFX1 gbuf_d_796(.A(n_3402), .Y(d_out_796));
CLKBUFX1 gbuf_q_796(.A(q_in_796), .Y(g3494));
CLKBUFX1 gbuf_d_797(.A(n_3403), .Y(d_out_797));
CLKBUFX1 gbuf_q_797(.A(q_in_797), .Y(g6537));
CLKBUFX1 gbuf_d_798(.A(n_3400), .Y(d_out_798));
CLKBUFX1 gbuf_q_798(.A(q_in_798), .Y(g3845));
XOR2X1 g64076(.A (n_3769), .B (n_6243), .Y (n_3770));
CLKBUFX1 gbuf_d_799(.A(n_3404), .Y(d_out_799));
CLKBUFX1 gbuf_q_799(.A(q_in_799), .Y(g3143));
CLKBUFX1 gbuf_d_800(.A(n_3395), .Y(d_out_800));
CLKBUFX1 gbuf_q_800(.A(q_in_800), .Y(g6191));
CLKBUFX1 gbuf_d_801(.A(n_3534), .Y(d_out_801));
CLKBUFX1 gbuf_q_801(.A(q_in_801), .Y(g5188));
CLKBUFX1 gbuf_d_802(.A(n_3531), .Y(d_out_802));
CLKBUFX1 gbuf_q_802(.A(q_in_802), .Y(g6227));
OAI22X1 g64078(.A0 (n_1557), .A1 (n_9599), .B0 (g4284), .B1 (n_9811),.Y (n_3767));
CLKBUFX1 gbuf_d_803(.A(n_3533), .Y(d_out_803));
CLKBUFX1 gbuf_q_803(.A(q_in_803), .Y(g3179));
CLKBUFX1 gbuf_d_804(.A(n_3530), .Y(d_out_804));
CLKBUFX1 gbuf_q_804(.A(q_in_804), .Y(g3881));
CLKBUFX1 gbuf_d_805(.A(n_3518), .Y(d_out_805));
CLKBUFX1 gbuf_q_805(.A(q_in_805), .Y(g4467));
OAI21X1 g64091(.A0 (n_3765), .A1 (n_9311), .B0 (n_3464), .Y (n_3766));
CLKBUFX1 gbuf_d_806(.A(g16924), .Y(d_out_806));
CLKBUFX1 gbuf_q_806(.A(q_in_806), .Y(g13881));
CLKBUFX1 gbuf_d_807(.A(g16874), .Y(d_out_807));
CLKBUFX1 gbuf_q_807(.A(q_in_807), .Y(g13865));
OR2X1 g64137(.A (g3106), .B (n_10943), .Y (n_6051));
OR2X1 g64148(.A (g3457), .B (n_3758), .Y (n_6052));
NAND2X1 g64170(.A (n_3543), .B (n_2653), .Y (n_3764));
NAND4X1 g64184(.A (g3550), .B (n_4682), .C (g14451), .D (n_10883), .Y(n_3761));
INVX1 g64200(.A (n_4424), .Y (n_3925));
BUFX3 g64203(.A (n_4424), .Y (n_4494));
BUFX3 g64204(.A (n_4424), .Y (n_4499));
BUFX3 g64205(.A (n_4424), .Y (n_4482));
BUFX3 g64209(.A (n_4424), .Y (n_4497));
NAND2X1 g64241(.A (n_2996), .B (n_3758), .Y (n_4447));
NAND3X1 g64271(.A (n_3775), .B (g4939), .C (n_9664), .Y (n_3755));
NAND3X1 g64272(.A (n_3779), .B (g4950), .C (n_9717), .Y (n_3753));
NAND3X1 g64273(.A (n_6243), .B (g4961), .C (n_10063), .Y (n_3752));
NOR2X1 g64317(.A (n_2014), .B (n_3775), .Y (n_3746));
INVX1 g64320(.A (n_3571), .Y (n_3745));
NOR2X1 g64325(.A (n_2016), .B (n_3779), .Y (n_3744));
NOR2X1 g64337(.A (n_2009), .B (n_6243), .Y (n_3742));
INVX4 g64345(.A (n_5471), .Y (n_4108));
NAND4X1 g64377(.A (n_10576), .B (g3538), .C (g14451), .D (n_10894),.Y (n_3740));
OAI22X1 g62680(.A0 (n_3314), .A1 (n_3687), .B0 (n_598), .B1 (n_9627),.Y (n_3738));
CLKBUFX1 gbuf_d_808(.A(g14518), .Y(d_out_808));
CLKBUFX1 gbuf_q_808(.A(q_in_808), .Y(g16955));
NAND3X1 g64529(.A (g5406), .B (n_9091), .C (g_5508), .Y (n_3737));
NAND3X1 g64535(.A (g3050), .B (n_9091), .C (g_6579), .Y (n_3736));
NAND3X1 g64543(.A (g6098), .B (n_9521), .C (g_14965), .Y (n_3735));
NAND3X1 g64545(.A (g6444), .B (n_9553), .C (g_3861), .Y (n_3734));
NAND3X1 g64558(.A (g3752), .B (n_9521), .C (g_5156), .Y (n_3733));
CLKBUFX1 gbuf_d_809(.A(n_3406), .Y(d_out_809));
CLKBUFX1 gbuf_q_809(.A(q_in_809), .Y(g5845));
AND2X1 g64565(.A (n_3732), .B (n_8917), .Y (n_4096));
NOR2X1 g64577(.A (n_3730), .B (n_3896), .Y (n_3731));
NOR2X1 g64578(.A (n_3728), .B (n_3896), .Y (n_3729));
NOR2X1 g64581(.A (n_3726), .B (n_3896), .Y (n_3727));
INVX1 g64597(.A (n_6005), .Y (n_3900));
CLKBUFX1 g64598(.A (n_6005), .Y (n_6334));
NAND3X1 g61796(.A (n_2809), .B (n_2234), .C (n_3074), .Y (n_3725));
CLKBUFX1 gbuf_d_810(.A(n_3255), .Y(d_out_810));
CLKBUFX1 gbuf_q_810(.A(q_in_810), .Y(n_10113));
OAI21X1 g64691(.A0 (g2965), .A1 (n_9311), .B0 (n_3377), .Y (n_3724));
OAI21X1 g64697(.A0 (n_2884), .A1 (n_2497), .B0 (n_3370), .Y (n_3723));
INVX1 g64760(.A (n_3540), .Y (n_3722));
NAND2X1 g62810(.A (n_3915), .B (n_3914), .Y (n_3913));
NOR2X1 g62823(.A (n_3257), .B (n_3720), .Y (n_3721));
NAND4X1 g62849(.A (n_3351), .B (n_8913), .C (n_10013), .D (n_10823),.Y (n_3717));
NAND3X1 g60979(.A (n_10005), .B (n_3059), .C (n_2252), .Y (n_3716));
XOR2X1 g62905(.A (n_640), .B (n_3713), .Y (n_3715));
OAI21X1 g64972(.A0 (n_1388), .A1 (n_9443), .B0 (n_3360), .Y (n_3712));
OAI21X1 g64974(.A0 (n_1375), .A1 (n_9903), .B0 (n_3361), .Y (n_3711));
OAI21X1 g64976(.A0 (n_1369), .A1 (n_9129), .B0 (n_3362), .Y (n_3710));
AOI21X1 g62929(.A0 (n_3707), .A1 (n_9836), .B0 (n_3352), .Y (n_3709));
OAI21X1 g62930(.A0 (n_3651), .A1 (n_3707), .B0 (n_3350), .Y (n_3708));
CLKBUFX1 gbuf_d_811(.A(n_3382), .Y(d_out_811));
CLKBUFX1 gbuf_q_811(.A(q_in_811), .Y(g1489));
CLKBUFX1 gbuf_d_812(.A(n_3263), .Y(d_out_812));
CLKBUFX1 gbuf_q_812(.A(q_in_812), .Y(n_10120));
AOI22X1 g64035(.A0 (n_2011), .A1 (n_5459), .B0 (n_11201), .B1(n_9193), .Y (n_3706));
INVX1 g65122(.A (g_7062), .Y (g9680));
INVX1 g65130(.A (g_5313), .Y (g8342));
CLKBUFX1 gbuf_d_813(.A(g8279), .Y(d_out_813));
CLKBUFX1 gbuf_qn_813(.A(qn_in_813), .Y(g3451));
CLKBUFX1 gbuf_d_814(.A(g9617), .Y(d_out_814));
CLKBUFX1 gbuf_qn_814(.A(qn_in_814), .Y(g5802));
CLKBUFX1 gbuf_d_815(.A(g8344), .Y(d_out_815));
CLKBUFX1 gbuf_qn_815(.A(qn_in_815), .Y(g3802));
CLKBUFX1 gbuf_d_816(.A(n_3353), .Y(d_out_816));
CLKBUFX1 gbuf_q_816(.A(q_in_816), .Y(g4459));
CLKBUFX1 gbuf_d_817(.A(g9743), .Y(d_out_817));
CLKBUFX1 gbuf_qn_817(.A(qn_in_817), .Y(g6494));
OAI22X1 g61386(.A0 (n_3075), .A1 (n_1985), .B0 (n_129), .B1 (n_9466),.Y (n_3703));
CLKBUFX1 gbuf_d_818(.A(g8215), .Y(d_out_818));
CLKBUFX1 gbuf_qn_818(.A(qn_in_818), .Y(g3100));
CLKBUFX1 gbuf_d_819(.A(g9682), .Y(d_out_819));
CLKBUFX1 gbuf_qn_819(.A(qn_in_819), .Y(g6148));
NAND4X1 g60988(.A (n_6735), .B (n_4866), .C (n_9359), .D (n_297), .Y(n_3702));
NOR2X1 g65349(.A (g4145), .B (g4253), .Y (n_3701));
CLKBUFX1 gbuf_d_820(.A(n_3292), .Y(d_out_820));
CLKBUFX1 gbuf_q_820(.A(q_in_820), .Y(n_11186));
MX2X1 g63083(.A (g_18793), .B (n_3058), .S0 (n_9218), .Y (n_3700));
CLKBUFX1 gbuf_d_821(.A(n_3261), .Y(d_out_821));
CLKBUFX1 gbuf_q_821(.A(q_in_821), .Y(g3698));
CLKBUFX1 gbuf_d_822(.A(n_3344), .Y(d_out_822));
CLKBUFX1 gbuf_q_822(.A(q_in_822), .Y(n_11013));
CLKBUFX1 gbuf_d_823(.A(n_3341), .Y(d_out_823));
CLKBUFX1 gbuf_q_823(.A(q_in_823), .Y(g4456));
CLKBUFX1 gbuf_d_824(.A(n_3336), .Y(d_out_824));
CLKBUFX1 gbuf_q_824(.A(q_in_824), .Y(g12184));
INVX1 g65715(.A (n_3697), .Y (n_5704));
NOR2X1 g65755(.A (n_3679), .B (n_8895), .Y (n_5705));
INVX1 g65867(.A (n_3695), .Y (n_5702));
CLKBUFX1 gbuf_d_825(.A(n_3345), .Y(d_out_825));
CLKBUFX1 gbuf_q_825(.A(q_in_825), .Y(g1246));
NOR2X1 g63192(.A (n_3325), .B (n_2437), .Y (n_3693));
XOR2X1 g61053(.A (n_1591), .B (n_3628), .Y (n_3692));
AND2X1 g63213(.A (n_3690), .B (g_10715), .Y (n_3691));
NAND3X1 g61006(.A (n_3312), .B (n_2268), .C (n_2875), .Y (n_3689));
NOR2X1 g63241(.A (n_3381), .B (n_3687), .Y (n_3688));
OAI21X1 g63260(.A0 (n_3431), .A1 (g_19414), .B0 (n_3334), .Y(n_3686));
AOI21X1 g63262(.A0 (n_3323), .A1 (n_1540), .B0 (n_3324), .Y (n_3685));
NAND4X1 g63270(.A (n_3329), .B (n_10188), .C (n_9894), .D (n_551), .Y(n_3683));
AOI21X1 g63302(.A0 (n_3234), .A1 (n_3439), .B0 (n_1417), .Y (n_3681));
AOI22X1 g63320(.A0 (n_2304), .A1 (n_3491), .B0 (n_1734), .B1(n_9627), .Y (n_3680));
INVX1 g66266(.A (n_3679), .Y (n_4231));
OAI21X1 g63331(.A0 (n_3563), .A1 (n_11134), .B0 (n_3328), .Y(n_3677));
MX2X1 g63358(.A (g_14265), .B (n_3175), .S0 (n_9000), .Y (n_3675));
MX2X1 g63359(.A (g_18795), .B (n_3043), .S0 (n_8955), .Y (n_3674));
MX2X1 g63360(.A (n_10103), .B (n_3038), .S0 (n_8955), .Y (n_3673));
MX2X1 g63363(.A (n_3042), .B (n_3040), .S0 (n_8955), .Y (n_3672));
MX2X1 g63364(.A (g_20073), .B (n_3041), .S0 (n_9279), .Y (n_3671));
MX2X1 g63369(.A (g_22464), .B (n_3034), .S0 (n_9156), .Y (n_3670));
CLKBUFX1 gbuf_d_826(.A(n_3300), .Y(d_out_826));
CLKBUFX1 gbuf_q_826(.A(q_in_826), .Y(g5348));
CLKBUFX1 gbuf_d_827(.A(n_3319), .Y(d_out_827));
CLKBUFX1 gbuf_qn_827(.A(qn_in_827), .Y(g5694));
CLKBUFX1 gbuf_d_828(.A(n_3299), .Y(d_out_828));
CLKBUFX1 gbuf_qn_828(.A(qn_in_828), .Y(g6040));
CLKBUFX1 gbuf_d_829(.A(n_3298), .Y(d_out_829));
CLKBUFX1 gbuf_qn_829(.A(qn_in_829), .Y(g6386));
CLKBUFX1 gbuf_d_830(.A(n_3296), .Y(d_out_830));
CLKBUFX1 gbuf_qn_830(.A(qn_in_830), .Y(g6732));
NAND3X1 g61052(.A (n_3373), .B (n_2283), .C (n_3187), .Y (n_3666));
AOI21X1 g61515(.A0 (n_10323), .A1 (g23683), .B0 (n_10321), .Y(n_4743));
NAND3X1 g63479(.A (n_3305), .B (n_2285), .C (n_2885), .Y (n_3662));
NAND3X1 g63489(.A (n_3661), .B (n_3660), .C (g_18793), .Y (n_4024));
NOR2X1 g63493(.A (n_3477), .B (n_2043), .Y (n_3659));
AOI22X1 g61020(.A0 (n_2253), .A1 (n_10330), .B0 (g1532), .B1(n_9772), .Y (n_3658));
AOI22X1 g63537(.A0 (n_3014), .A1 (n_8639), .B0 (n_607), .B1 (n_3013),.Y (n_3656));
NAND3X1 g63539(.A (n_2746), .B (n_2545), .C (n_3027), .Y (n_3655));
OR2X1 g63550(.A (n_3309), .B (n_3915), .Y (n_3654));
AOI22X1 g63559(.A0 (n_3029), .A1 (n_9501), .B0 (n_2657), .B1(n_3323), .Y (n_3653));
CLKBUFX1 gbuf_d_831(.A(n_3320), .Y(d_out_831));
CLKBUFX1 gbuf_q_831(.A(q_in_831), .Y(g_20951));
NAND4X1 g62251(.A (n_3333), .B (n_3651), .C (n_9834), .D (n_10818),.Y (n_3652));
XOR2X1 g63644(.A (n_662), .B (n_3258), .Y (n_3648));
NOR2X1 g61038(.A (n_3288), .B (n_961), .Y (n_3647));
CLKBUFX1 gbuf_d_832(.A(g10306), .Y(d_out_832));
CLKBUFX1 gbuf_q_832(.A(q_in_832), .Y(g4423));
NAND2X1 g63889(.A (n_3645), .B (n_662), .Y (n_3646));
NOR2X1 g63907(.A (n_7243), .B (n_3641), .Y (n_3642));
INVX1 g63950(.A (n_3639), .Y (n_3640));
NAND2X1 g63970(.A (n_3247), .B (n_3015), .Y (n_3638));
NAND3X1 g63979(.A (n_6970), .B (n_2364), .C (n_3218), .Y (n_3637));
INVX1 g61048(.A (n_3860), .Y (n_3778));
CLKBUFX1 gbuf_d_833(.A(n_3359), .Y(d_out_833));
CLKBUFX1 gbuf_q_833(.A(q_in_833), .Y(g10122));
CLKBUFX1 gbuf_d_834(.A(n_3348), .Y(d_out_834));
CLKBUFX1 gbuf_q_834(.A(q_in_834), .Y(g1306));
CLKBUFX1 gbuf_d_835(.A(n_3347), .Y(d_out_835));
CLKBUFX1 gbuf_q_835(.A(q_in_835), .Y(g_18488));
OAI21X1 g64040(.A0 (n_227), .A1 (n_9681), .B0 (n_3285), .Y (n_3636));
CLKBUFX1 gbuf_d_836(.A(n_3322), .Y(d_out_836));
CLKBUFX1 gbuf_q_836(.A(q_in_836), .Y(g5689));
CLKBUFX1 gbuf_d_837(.A(n_3317), .Y(d_out_837));
CLKBUFX1 gbuf_q_837(.A(q_in_837), .Y(g_20614));
CLKBUFX1 gbuf_d_838(.A(n_3308), .Y(d_out_838));
CLKBUFX1 gbuf_q_838(.A(q_in_838), .Y(g_18902));
CLKBUFX1 gbuf_d_839(.A(n_3279), .Y(d_out_839));
CLKBUFX1 gbuf_q_839(.A(q_in_839), .Y(g_11413));
CLKBUFX1 gbuf_d_840(.A(n_3262), .Y(d_out_840));
CLKBUFX1 gbuf_q_840(.A(q_in_840), .Y(g3347));
CLKBUFX1 gbuf_d_841(.A(n_3355), .Y(d_out_841));
CLKBUFX1 gbuf_q_841(.A(q_in_841), .Y(g4349));
CLKBUFX1 gbuf_d_842(.A(n_3303), .Y(d_out_842));
CLKBUFX1 gbuf_q_842(.A(q_in_842), .Y(g17291));
CLKBUFX1 gbuf_d_843(.A(n_3315), .Y(d_out_843));
CLKBUFX1 gbuf_q_843(.A(q_in_843), .Y(g5343));
XOR2X1 g64065(.A (n_11201), .B (n_5459), .Y (n_3634));
CLKBUFX1 gbuf_d_844(.A(n_3313), .Y(d_out_844));
CLKBUFX1 gbuf_q_844(.A(q_in_844), .Y(g6381));
CLKBUFX1 gbuf_d_845(.A(n_3301), .Y(d_out_845));
CLKBUFX1 gbuf_q_845(.A(q_in_845), .Y(g6035));
CLKBUFX1 gbuf_d_846(.A(n_3273), .Y(d_out_846));
CLKBUFX1 gbuf_q_846(.A(q_in_846), .Y(n_2458));
XOR2X1 g64066(.A (n_10660), .B (n_10948), .Y (n_3633));
CLKBUFX1 gbuf_d_847(.A(n_3274), .Y(d_out_847));
CLKBUFX1 gbuf_q_847(.A(q_in_847), .Y(g34026));
CLKBUFX1 gbuf_d_848(.A(n_3290), .Y(d_out_848));
CLKBUFX1 gbuf_q_848(.A(q_in_848), .Y(g5152));
CLKBUFX1 gbuf_d_849(.A(n_3289), .Y(d_out_849));
CLKBUFX1 gbuf_q_849(.A(q_in_849), .Y(g_13838));
XOR2X1 g64069(.A (n_8806), .B (g28753), .Y (n_3631));
CLKBUFX1 gbuf_d_850(.A(n_3254), .Y(d_out_850));
CLKBUFX1 gbuf_q_850(.A(q_in_850), .Y(g3111));
CLKBUFX1 gbuf_d_851(.A(n_3283), .Y(d_out_851));
CLKBUFX1 gbuf_q_851(.A(q_in_851), .Y(g1472));
CLKBUFX1 gbuf_d_852(.A(n_3282), .Y(d_out_852));
CLKBUFX1 gbuf_q_852(.A(q_in_852), .Y(g1478));
CLKBUFX1 gbuf_d_853(.A(n_3270), .Y(d_out_853));
CLKBUFX1 gbuf_q_853(.A(q_in_853), .Y(g4628));
XOR2X1 g61054(.A (g1333), .B (n_3628), .Y (n_3629));
CLKBUFX1 gbuf_d_854(.A(n_3358), .Y(d_out_854));
CLKBUFX1 gbuf_q_854(.A(q_in_854), .Y(g_18015));
XOR2X1 g64081(.A (n_3626), .B (g6395), .Y (n_3627));
CLKBUFX1 gbuf_d_855(.A(n_3335), .Y(d_out_855));
CLKBUFX1 gbuf_q_855(.A(q_in_855), .Y(g2763));
CLKBUFX1 gbuf_d_856(.A(n_3337), .Y(d_out_856));
CLKBUFX1 gbuf_q_856(.A(q_in_856), .Y(g4057));
CLKBUFX1 gbuf_d_857(.A(n_3339), .Y(d_out_857));
CLKBUFX1 gbuf_q_857(.A(q_in_857), .Y(g4087));
CLKBUFX1 gbuf_d_858(.A(n_3340), .Y(d_out_858));
CLKBUFX1 gbuf_q_858(.A(q_in_858), .Y(g4141));
CLKBUFX1 gbuf_d_859(.A(n_3343), .Y(d_out_859));
CLKBUFX1 gbuf_q_859(.A(q_in_859), .Y(g4417));
XOR2X1 g64094(.A (n_3624), .B (n_10398), .Y (n_3625));
NOR2X1 g65313(.A (g3003), .B (n_9453), .Y (g21727));
MX2X1 g64101(.A (g4894), .B (n_3217), .S0 (n_9218), .Y (n_3622));
NOR2X1 g64134(.A (n_3389), .B (n_9775), .Y (n_3621));
NAND3X1 g61709(.A (n_2868), .B (n_2604), .C (n_3153), .Y (n_3620));
NOR2X1 g64161(.A (g2886), .B (g2946), .Y (n_3615));
NOR2X1 g64167(.A (g2946), .B (g2955), .Y (n_3614));
NAND3X1 g64168(.A (n_3612), .B (n_3611), .C (n_9894), .Y (n_3613));
NAND3X1 g64180(.A (n_3605), .B (n_3604), .C (n_9698), .Y (n_3606));
NAND2X1 g64182(.A (n_3775), .B (n_64), .Y (n_3603));
NAND2X2 g64210(.A (g4284), .B (n_10871), .Y (n_4424));
NAND2X1 g64212(.A (n_3779), .B (n_1818), .Y (n_3599));
NAND2X1 g64214(.A (n_3779), .B (n_6978), .Y (n_3598));
NAND2X1 g64227(.A (n_6243), .B (n_151), .Y (n_3593));
NAND2X1 g64228(.A (n_3775), .B (n_7003), .Y (n_3592));
NAND3X1 g64229(.A (n_3241), .B (n_2539), .C (n_2920), .Y (n_3591));
NAND3X1 g64234(.A (n_3784), .B (n_3589), .C (n_9811), .Y (n_3590));
NAND3X1 g64248(.A (n_8707), .B (g4704), .C (n_9448), .Y (n_3588));
NAND3X1 g61725(.A (n_3221), .B (n_2281), .C (n_3170), .Y (n_3585));
NAND3X1 g64252(.A (n_10947), .B (g4749), .C (n_9834), .Y (n_3582));
NAND3X1 g64254(.A (n_3612), .B (g4760), .C (n_9627), .Y (n_3581));
NAND3X1 g64255(.A (n_3784), .B (g4771), .C (n_10063), .Y (n_3580));
NAND3X1 g64270(.A (n_3605), .B (g4894), .C (n_9750), .Y (n_3578));
NAND2X1 g64280(.A (n_3189), .B (n_3387), .Y (n_3577));
INVX1 g62580(.A (n_3448), .Y (n_4045));
INVX1 g64303(.A (n_6676), .Y (n_3574));
INVX1 g64318(.A (n_3441), .Y (n_3572));
AOI21X1 g64321(.A0 (n_3569), .A1 (n_1285), .B0 (n_3390), .Y (n_3571));
AOI21X1 g64322(.A0 (n_3569), .A1 (g_12791), .B0 (n_3566), .Y(n_3570));
NAND3X1 g64329(.A (n_3566), .B (n_456), .C (n_9425), .Y (n_3567));
INVX2 g64347(.A (n_10270), .Y (n_5471));
NAND4X1 g62644(.A (n_3307), .B (n_3563), .C (n_9209), .D (n_684), .Y(n_3564));
OAI21X1 g64395(.A0 (g16624), .A1 (g14421), .B0 (n_3210), .Y (n_3561));
OAI21X1 g64396(.A0 (g16656), .A1 (g14451), .B0 (n_3209), .Y (n_3560));
INVX1 g61302(.A (g1589), .Y (n_4149));
MX2X1 g64406(.A (n_10568), .B (g14189), .S0 (n_5582), .Y (n_3559));
AOI22X1 g64417(.A0 (n_3003), .A1 (g_21576), .B0 (n_3569), .B1(n_640), .Y (n_3557));
MX2X1 g64447(.A (n_11113), .B (n_3185), .S0 (n_10005), .Y (n_3555));
NOR2X1 g61315(.A (g_6701), .B (n_6705), .Y (n_4134));
MX2X1 g64461(.A (n_3388), .B (n_3178), .S0 (n_9333), .Y (n_3554));
NAND2X1 g64527(.A (n_3368), .B (n_3216), .Y (n_3552));
NAND3X1 g64567(.A (n_3569), .B (n_3550), .C (n_9466), .Y (n_3551));
XOR2X1 g64077(.A (n_523), .B (n_3547), .Y (n_3549));
NOR2X1 g64599(.A (g4581), .B (n_10376), .Y (n_6005));
NAND2X1 g64602(.A (n_3182), .B (n_3349), .Y (n_3546));
NAND3X1 g64658(.A (n_10940), .B (g3263), .C (n_10941), .Y (n_3543));
NAND3X1 g64683(.A (n_3398), .B (g3614), .C (n_6973), .Y (n_3542));
NAND4X1 g64739(.A (g3554), .B (n_10889), .C (g16656), .D (n_11128),.Y (n_3541));
NAND4X1 g64761(.A (n_1578), .B (n_3073), .C (n_9398), .D (n_477), .Y(n_3540));
XOR2X1 g64789(.A (g4311), .B (n_10396), .Y (n_3538));
INVX1 g64811(.A (g4581), .Y (n_5711));
CLKBUFX1 gbuf_d_860(.A(g16693), .Y(d_out_860));
CLKBUFX1 gbuf_q_860(.A(q_in_860), .Y(g14518));
AOI21X1 g62847(.A0 (n_3651), .A1 (n_10226), .B0 (n_8694), .Y(n_3537));
AND2X1 g64881(.A (n_5402), .B (g16693), .Y (n_3732));
NAND2X1 g64969(.A (g16693), .B (g16659), .Y (n_3535));
OAI21X1 g64971(.A0 (n_1390), .A1 (n_9129), .B0 (n_3160), .Y (n_3534));
OAI21X1 g64973(.A0 (n_1373), .A1 (n_9193), .B0 (n_3154), .Y (n_3533));
OAI21X1 g64975(.A0 (n_1384), .A1 (n_10952), .B0 (n_3158), .Y(n_3532));
OAI21X1 g64977(.A0 (n_1380), .A1 (n_9193), .B0 (n_3157), .Y (n_3531));
OAI21X1 g64978(.A0 (n_1366), .A1 (n_9628), .B0 (n_3156), .Y (n_3530));
OAI22X1 g62931(.A0 (n_3506), .A1 (n_2587), .B0 (n_1274), .B1(n_9651), .Y (n_3529));
INVX1 g65118(.A (g_5156), .Y (g8398));
INVX1 g65120(.A (g_6579), .Y (g8277));
CLKBUFX1 gbuf_d_861(.A(n_3120), .Y(d_out_861));
CLKBUFX1 gbuf_qn_861(.A(qn_in_861), .Y(g_7062));
INVX1 g65124(.A (g_5508), .Y (g9615));
INVX1 g65126(.A (g_14965), .Y (g9741));
INVX1 g65128(.A (g_3861), .Y (g9817));
CLKBUFX1 gbuf_d_862(.A(n_3112), .Y(d_out_862));
CLKBUFX1 gbuf_qn_862(.A(qn_in_862), .Y(g_5313));
NAND3X1 g61130(.A (n_3124), .B (g1389), .C (n_9811), .Y (n_3523));
CLKBUFX1 gbuf_d_863(.A(g9555), .Y(d_out_863));
CLKBUFX1 gbuf_qn_863(.A(qn_in_863), .Y(g5456));
CLKBUFX1 gbuf_d_864(.A(g14189), .Y(d_out_864));
CLKBUFX1 gbuf_q_864(.A(q_in_864), .Y(g14201));
NAND2X1 g65326(.A (g_13255), .B (g_13901), .Y (n_3522));
CLKBUFX1 gbuf_d_865(.A(n_3116), .Y(d_out_865));
CLKBUFX1 gbuf_q_865(.A(q_in_865), .Y(g4489));
OAI21X1 g64071(.A0 (n_10751), .A1 (g_15287), .B0 (n_3033), .Y(n_3521));
OAI22X1 g61962(.A0 (n_3489), .A1 (n_2161), .B0 (n_143), .B1 (n_9862),.Y (n_3520));
CLKBUFX1 gbuf_d_866(.A(n_3018), .Y(d_out_866));
CLKBUFX1 gbuf_q_866(.A(q_in_866), .Y(n_2429));
INVX1 g65561(.A (g_11037), .Y (g9497));
INVX1 g65574(.A (g2724), .Y (n_3868));
INVX1 g65585(.A (g4145), .Y (n_3896));
NAND2X1 g65701(.A (n_1353), .B (n_3072), .Y (n_3518));
OR2X1 g65716(.A (g2715), .B (n_8898), .Y (n_3697));
XOR2X1 g64070(.A (g_13278), .B (n_3291), .Y (n_3517));
NAND2X1 g65868(.A (g2715), .B (n_8895), .Y (n_3695));
NAND3X1 g63243(.A (n_10005), .B (n_2757), .C (n_10647), .Y (n_3516));
CLKBUFX1 gbuf_d_867(.A(n_3122), .Y(d_out_867));
CLKBUFX1 gbuf_q_867(.A(q_in_867), .Y(g9553));
CLKBUFX1 gbuf_d_868(.A(n_3052), .Y(d_out_868));
CLKBUFX1 gbuf_q_868(.A(q_in_868), .Y(g_6131));
AOI21X1 g63269(.A0 (n_3563), .A1 (n_741), .B0 (n_10296), .Y (n_3514));
OAI21X1 g63280(.A0 (n_7383), .A1 (n_9333), .B0 (n_3066), .Y (n_3512));
OAI21X1 g63282(.A0 (n_10889), .A1 (n_9797), .B0 (n_3063), .Y(n_3511));
MX2X1 g64100(.A (g4771), .B (n_2959), .S0 (n_9000), .Y (n_3510));
NAND3X1 g62103(.A (n_2800), .B (n_2697), .C (n_2764), .Y (n_3508));
OAI22X1 g62114(.A0 (n_3506), .A1 (n_2926), .B0 (n_165), .B1 (n_9992),.Y (n_3507));
NOR2X1 g63426(.A (n_8835), .B (n_8768), .Y (n_3505));
OAI21X1 g63440(.A0 (n_3502), .A1 (n_3501), .B0 (n_9279), .Y (n_3503));
OR2X1 g63474(.A (n_3499), .B (n_3497), .Y (n_3500));
NOR2X1 g63477(.A (n_2677), .B (n_3497), .Y (n_3498));
CLKBUFX1 gbuf_d_869(.A(n_3077), .Y(d_out_869));
CLKBUFX1 gbuf_q_869(.A(q_in_869), .Y(g4239));
AOI21X1 g63484(.A0 (n_2751), .A1 (n_2744), .B0 (n_9976), .Y (n_3496));
NOR2X1 g63509(.A (n_8835), .B (n_8837), .Y (n_3855));
AOI21X1 g63526(.A0 (n_1783), .A1 (n_3493), .B0 (n_9836), .Y (n_3494));
AOI21X1 g63527(.A0 (n_7260), .A1 (g4349), .B0 (n_3491), .Y (n_3492));
OAI22X1 g63538(.A0 (n_3489), .A1 (n_1308), .B0 (g4688), .B1 (n_9830),.Y (n_3490));
AOI22X1 g63551(.A0 (n_2519), .A1 (n_10115), .B0 (g_12433), .B1(n_9693), .Y (n_3488));
CLKBUFX1 gbuf_d_870(.A(n_3055), .Y(d_out_870));
CLKBUFX1 gbuf_q_870(.A(q_in_870), .Y(g_22379));
CLKBUFX1 gbuf_d_871(.A(n_3053), .Y(d_out_871));
CLKBUFX1 gbuf_q_871(.A(q_in_871), .Y(g_19241));
CLKBUFX1 gbuf_d_872(.A(n_3138), .Y(d_out_872));
CLKBUFX1 gbuf_q_872(.A(q_in_872), .Y(g_14587));
OAI21X1 g63623(.A0 (n_3486), .A1 (n_3894), .B0 (n_2239), .Y (n_3487));
CLKBUFX1 gbuf_d_873(.A(n_3114), .Y(d_out_873));
CLKBUFX1 gbuf_q_873(.A(q_in_873), .Y(g4492));
CLKBUFX1 gbuf_d_874(.A(n_3136), .Y(d_out_874));
CLKBUFX1 gbuf_q_874(.A(q_in_874), .Y(g4153));
CLKBUFX1 gbuf_d_875(.A(n_3057), .Y(d_out_875));
CLKBUFX1 gbuf_q_875(.A(q_in_875), .Y(g_20837));
CLKBUFX1 gbuf_d_876(.A(n_3141), .Y(d_out_876));
CLKBUFX1 gbuf_q_876(.A(q_in_876), .Y(n_1191));
CLKBUFX1 gbuf_d_877(.A(n_3139), .Y(d_out_877));
CLKBUFX1 gbuf_q_877(.A(q_in_877), .Y(g2984));
INVX1 g61035(.A (n_6735), .Y (n_3484));
OAI22X1 g61222(.A0 (n_2672), .A1 (n_2562), .B0 (n_26), .B1 (n_9651),.Y (n_3483));
CLKBUFX1 gbuf_d_878(.A(n_3133), .Y(d_out_878));
CLKBUFX1 gbuf_q_878(.A(q_in_878), .Y(g_21651));
INVX1 g63926(.A (n_6767), .Y (n_3482));
NAND2X1 g63936(.A (g4072), .B (n_9952), .Y (n_3481));
NAND2X1 g63937(.A (g4072), .B (n_43), .Y (n_3480));
NAND2X1 g63947(.A (g4072), .B (n_98), .Y (n_3479));
NAND3X1 g63951(.A (n_3028), .B (n_83), .C (g_14265), .Y (n_3639));
CLKBUFX1 gbuf_d_879(.A(n_3131), .Y(d_out_879));
CLKBUFX1 gbuf_q_879(.A(q_in_879), .Y(g4273));
OAI33X1 g63962(.A0 (n_1137), .A1 (n_2642), .A2 (n_546), .B0(n_10180), .B1 (n_1100), .B2 (n_75), .Y (n_3478));
INVX1 g63996(.A (n_3477), .Y (n_3845));
NAND2X2 g61049(.A (n_1444), .B (n_10330), .Y (n_3860));
CLKBUFX1 gbuf_d_880(.A(n_3167), .Y(d_out_880));
CLKBUFX1 gbuf_qn_880(.A(qn_in_880), .Y(g1339));
CLKBUFX1 gbuf_d_881(.A(n_3010), .Y(d_out_881));
CLKBUFX1 gbuf_q_881(.A(q_in_881), .Y(g6167));
OAI22X1 g64024(.A0 (n_3506), .A1 (n_1827), .B0 (g4878), .B1(n_10063), .Y (n_3475));
CLKBUFX1 gbuf_d_882(.A(n_3143), .Y(d_out_882));
CLKBUFX1 gbuf_q_882(.A(q_in_882), .Y(g20557));
NAND4X1 g64059(.A (n_2378), .B (n_2965), .C (n_2025), .D (n_2027), .Y(n_11188));
CLKBUFX1 gbuf_d_883(.A(n_3056), .Y(d_out_883));
CLKBUFX1 gbuf_q_883(.A(q_in_883), .Y(g_21806));
CLKBUFX1 gbuf_d_884(.A(n_3012), .Y(d_out_884));
CLKBUFX1 gbuf_qn_884(.A(qn_in_884), .Y(g5495));
CLKBUFX1 gbuf_d_885(.A(n_3008), .Y(d_out_885));
CLKBUFX1 gbuf_qn_885(.A(qn_in_885), .Y(g6533));
CLKBUFX1 gbuf_d_886(.A(n_3005), .Y(d_out_886));
CLKBUFX1 gbuf_q_886(.A(q_in_886), .Y(g_15758));
CLKBUFX1 gbuf_d_887(.A(n_3212), .Y(d_out_887));
CLKBUFX1 gbuf_q_887(.A(q_in_887), .Y(n_276));
CLKBUFX1 gbuf_d_888(.A(n_3147), .Y(d_out_888));
CLKBUFX1 gbuf_q_888(.A(q_in_888), .Y(n_1177));
CLKBUFX1 gbuf_d_889(.A(n_3146), .Y(d_out_889));
CLKBUFX1 gbuf_q_889(.A(q_in_889), .Y(n_1234));
CLKBUFX1 gbuf_d_890(.A(n_3140), .Y(d_out_890));
CLKBUFX1 gbuf_q_890(.A(q_in_890), .Y(n_1169));
CLKBUFX1 gbuf_d_891(.A(n_3144), .Y(d_out_891));
CLKBUFX1 gbuf_q_891(.A(q_in_891), .Y(n_1216));
CLKBUFX1 gbuf_d_892(.A(n_3145), .Y(d_out_892));
CLKBUFX1 gbuf_q_892(.A(q_in_892), .Y(n_1135));
CLKBUFX1 gbuf_d_893(.A(n_3142), .Y(d_out_893));
CLKBUFX1 gbuf_q_893(.A(q_in_893), .Y(n_1210));
CLKBUFX1 gbuf_d_894(.A(n_3137), .Y(d_out_894));
CLKBUFX1 gbuf_q_894(.A(q_in_894), .Y(g8291));
CLKBUFX1 gbuf_d_895(.A(n_3132), .Y(d_out_895));
CLKBUFX1 gbuf_q_895(.A(q_in_895), .Y(g4172));
CLKBUFX1 gbuf_d_896(.A(n_3119), .Y(d_out_896));
CLKBUFX1 gbuf_q_896(.A(q_in_896), .Y(g4486));
CLKBUFX1 gbuf_d_897(.A(n_3105), .Y(d_out_897));
CLKBUFX1 gbuf_q_897(.A(q_in_897), .Y(g2912));
CLKBUFX1 gbuf_d_898(.A(n_3096), .Y(d_out_898));
CLKBUFX1 gbuf_q_898(.A(q_in_898), .Y(g2868));
CLKBUFX1 gbuf_d_899(.A(n_3090), .Y(d_out_899));
CLKBUFX1 gbuf_q_899(.A(q_in_899), .Y(g2936));
CLKBUFX1 gbuf_d_900(.A(n_3097), .Y(d_out_900));
CLKBUFX1 gbuf_q_900(.A(q_in_900), .Y(g1779));
CLKBUFX1 gbuf_d_901(.A(n_3111), .Y(d_out_901));
CLKBUFX1 gbuf_q_901(.A(q_in_901), .Y(g1798));
CLKBUFX1 gbuf_d_902(.A(n_3106), .Y(d_out_902));
CLKBUFX1 gbuf_q_902(.A(q_in_902), .Y(g1913));
CLKBUFX1 gbuf_d_903(.A(n_3080), .Y(d_out_903));
CLKBUFX1 gbuf_q_903(.A(q_in_903), .Y(g1932));
CLKBUFX1 gbuf_d_904(.A(n_3102), .Y(d_out_904));
CLKBUFX1 gbuf_q_904(.A(q_in_904), .Y(g21292));
CLKBUFX1 gbuf_d_905(.A(n_3127), .Y(d_out_905));
CLKBUFX1 gbuf_q_905(.A(q_in_905), .Y(g8719));
CLKBUFX1 gbuf_d_906(.A(n_3099), .Y(d_out_906));
CLKBUFX1 gbuf_q_906(.A(q_in_906), .Y(g2047));
CLKBUFX1 gbuf_d_907(.A(n_3098), .Y(d_out_907));
CLKBUFX1 gbuf_q_907(.A(q_in_907), .Y(g2066));
CLKBUFX1 gbuf_d_908(.A(n_3095), .Y(d_out_908));
CLKBUFX1 gbuf_q_908(.A(q_in_908), .Y(g4146));
CLKBUFX1 gbuf_d_909(.A(n_3103), .Y(d_out_909));
CLKBUFX1 gbuf_q_909(.A(q_in_909), .Y(g2204));
CLKBUFX1 gbuf_d_910(.A(n_3108), .Y(d_out_910));
CLKBUFX1 gbuf_q_910(.A(q_in_910), .Y(g2223));
CLKBUFX1 gbuf_d_911(.A(n_3094), .Y(d_out_911));
CLKBUFX1 gbuf_q_911(.A(q_in_911), .Y(g4249));
CLKBUFX1 gbuf_d_912(.A(n_3081), .Y(d_out_912));
CLKBUFX1 gbuf_q_912(.A(q_in_912), .Y(g2922));
CLKBUFX1 gbuf_d_913(.A(n_3091), .Y(d_out_913));
CLKBUFX1 gbuf_q_913(.A(q_in_913), .Y(g2338));
CLKBUFX1 gbuf_d_914(.A(n_3085), .Y(d_out_914));
CLKBUFX1 gbuf_q_914(.A(q_in_914), .Y(g2357));
CLKBUFX1 gbuf_d_915(.A(n_3130), .Y(d_out_915));
CLKBUFX1 gbuf_q_915(.A(q_in_915), .Y(n_7247));
CLKBUFX1 gbuf_d_916(.A(n_3088), .Y(d_out_916));
CLKBUFX1 gbuf_q_916(.A(q_in_916), .Y(g4717));
CLKBUFX1 gbuf_d_917(.A(n_3086), .Y(d_out_917));
CLKBUFX1 gbuf_q_917(.A(q_in_917), .Y(g1664));
CLKBUFX1 gbuf_d_918(.A(n_3084), .Y(d_out_918));
CLKBUFX1 gbuf_q_918(.A(q_in_918), .Y(g2472));
CLKBUFX1 gbuf_d_919(.A(n_3082), .Y(d_out_919));
CLKBUFX1 gbuf_q_919(.A(q_in_919), .Y(g2491));
CLKBUFX1 gbuf_d_920(.A(n_3092), .Y(d_out_920));
CLKBUFX1 gbuf_q_920(.A(q_in_920), .Y(g4907));
CLKBUFX1 gbuf_d_921(.A(n_3079), .Y(d_out_921));
CLKBUFX1 gbuf_q_921(.A(q_in_921), .Y(g2606));
CLKBUFX1 gbuf_d_922(.A(n_3109), .Y(d_out_922));
CLKBUFX1 gbuf_q_922(.A(q_in_922), .Y(g1644));
CLKBUFX1 gbuf_d_923(.A(n_3100), .Y(d_out_923));
CLKBUFX1 gbuf_q_923(.A(q_in_923), .Y(g2625));
CLKBUFX1 gbuf_d_924(.A(n_3104), .Y(d_out_924));
CLKBUFX1 gbuf_q_924(.A(q_in_924), .Y(g2994));
CLKBUFX1 gbuf_d_925(.A(n_3070), .Y(d_out_925));
CLKBUFX1 gbuf_q_925(.A(q_in_925), .Y(g1291));
MX2X1 g64095(.A (g20652), .B (n_2678), .S0 (n_8955), .Y (n_3473));
MX2X1 g64097(.A (g4704), .B (n_2961), .S0 (n_9234), .Y (n_3471));
MX2X1 g64098(.A (g4749), .B (n_2962), .S0 (n_8955), .Y (n_3470));
MX2X1 g64099(.A (g4760), .B (n_2960), .S0 (n_9000), .Y (n_3469));
MX2X1 g64102(.A (g4939), .B (n_2963), .S0 (n_9000), .Y (n_3468));
MX2X1 g64103(.A (g4950), .B (n_2958), .S0 (n_9156), .Y (n_3466));
MX2X1 g64104(.A (g4961), .B (n_2957), .S0 (n_9311), .Y (n_3465));
OAI21X1 g64136(.A0 (n_2942), .A1 (n_3463), .B0 (n_9091), .Y (n_3464));
NAND3X1 g64179(.A (n_2989), .B (n_2243), .C (n_2632), .Y (n_3461));
OAI33X1 g61062(.A0 (n_2841), .A1 (n_3365), .A2 (n_3459), .B0(n_11073), .B1 (n_3459), .B2 (n_10245), .Y (n_3460));
NAND3X1 g61721(.A (n_2979), .B (n_2245), .C (n_2870), .Y (n_3458));
INVX2 g64232(.A (n_3814), .Y (n_3455));
NAND3X1 g61723(.A (n_3222), .B (n_2557), .C (n_2350), .Y (n_3454));
NAND3X1 g64244(.A (n_10398), .B (g4616), .C (g4584), .Y (n_4843));
AOI21X1 g64290(.A0 (n_2641), .A1 (n_2934), .B0 (n_3391), .Y (n_3449));
NAND2X1 g62581(.A (n_3447), .B (g_15381), .Y (n_3448));
NAND4X1 g64307(.A (n_3030), .B (n_1262), .C (n_3021), .D (n_2456), .Y(n_3442));
AOI21X1 g64316(.A0 (n_2983), .A1 (n_10867), .B0 (n_3832), .Y(n_3831));
AOI21X1 g64319(.A0 (n_3569), .A1 (g_14265), .B0 (n_3174), .Y(n_3441));
AOI21X1 g64324(.A0 (n_2670), .A1 (n_10871), .B0 (n_3838), .Y(n_3837));
AOI21X1 g64340(.A0 (n_11033), .A1 (n_10867), .B0 (n_8629), .Y(n_3873));
AOI21X1 g64342(.A0 (n_11036), .A1 (n_10867), .B0 (n_8634), .Y(n_3870));
OAI21X1 g64352(.A0 (n_3425), .A1 (n_3439), .B0 (n_3438), .Y (n_3440));
AOI21X1 g64356(.A0 (g14662), .A1 (n_465), .B0 (n_3228), .Y (n_3437));
AOI21X1 g64357(.A0 (g14694), .A1 (n_409), .B0 (n_3229), .Y (n_3436));
AOI21X1 g64358(.A0 (g14738), .A1 (n_11045), .B0 (n_3226), .Y(n_3435));
AOI21X1 g64359(.A0 (g14779), .A1 (n_660), .B0 (n_3225), .Y (n_3434));
AOI21X1 g64360(.A0 (g14828), .A1 (n_322), .B0 (n_3223), .Y (n_3433));
OR2X1 g64367(.A (n_3004), .B (n_3431), .Y (n_3432));
XOR2X1 g64374(.A (n_3894), .B (n_3486), .Y (n_3430));
OAI22X1 g64375(.A0 (n_1568), .A1 (n_3569), .B0 (n_3003), .B1 (n_708),.Y (n_3429));
AOI21X1 g64404(.A0 (g5033), .A1 (n_9193), .B0 (n_3233), .Y (n_3427));
CLKBUFX1 gbuf_d_926(.A(n_3179), .Y(d_out_926));
CLKBUFX1 gbuf_q_926(.A(q_in_926), .Y(g1589));
XOR2X1 g64410(.A (n_659), .B (n_3425), .Y (n_3426));
MX2X1 g64415(.A (g_19233), .B (g_17065), .S0 (n_3003), .Y (n_3424));
MX2X1 g64416(.A (n_11162), .B (n_3550), .S0 (n_3003), .Y (n_3423));
MX2X1 g64418(.A (g_21778), .B (g_19113), .S0 (n_3003), .Y (n_3422));
MX2X1 g64419(.A (g_17065), .B (g_16677), .S0 (n_3003), .Y (n_3420));
MX2X1 g64420(.A (g_16677), .B (g_20208), .S0 (n_3003), .Y (n_3418));
MX2X1 g64421(.A (g_21720), .B (g_13758), .S0 (n_3003), .Y (n_3417));
MX2X1 g64422(.A (g_13758), .B (g_19289), .S0 (n_3003), .Y (n_3416));
MX2X1 g64423(.A (g_19289), .B (n_5663), .S0 (n_3003), .Y (n_3415));
OAI21X1 g62667(.A0 (n_221), .A1 (n_9311), .B0 (n_3193), .Y (n_3414));
MX2X1 g64442(.A (g_17426), .B (n_2891), .S0 (n_9172), .Y (n_3413));
OAI22X1 g62679(.A0 (n_3489), .A1 (n_1989), .B0 (n_294), .B1 (n_9862),.Y (n_3412));
INVX1 g64472(.A (g5069), .Y (n_3411));
INVX1 g64488(.A (g2946), .Y (n_3410));
CLKBUFX1 gbuf_d_927(.A(n_3176), .Y(d_out_927));
CLKBUFX1 gbuf_qn_927(.A(qn_in_927), .Y(g_7563));
CLKBUFX1 gbuf_d_928(.A(g14421), .Y(d_out_928));
CLKBUFX1 gbuf_q_928(.A(q_in_928), .Y(g16874));
CLKBUFX1 gbuf_d_929(.A(g14451), .Y(d_out_929));
CLKBUFX1 gbuf_q_929(.A(q_in_929), .Y(g16924));
NOR2X1 g64522(.A (n_3208), .B (n_653), .Y (n_3409));
CLKBUFX1 gbuf_d_930(.A(n_3087), .Y(d_out_930));
CLKBUFX1 gbuf_q_930(.A(q_in_930), .Y(g4722));
OAI21X1 g64531(.A0 (n_2372), .A1 (n_887), .B0 (n_3194), .Y (n_3408));
AOI21X1 g61327(.A0 (n_2060), .A1 (n_26), .B0 (n_3186), .Y (n_3407));
OAI21X1 g64534(.A0 (n_2370), .A1 (n_882), .B0 (n_3207), .Y (n_3406));
OAI21X1 g64544(.A0 (n_2615), .A1 (n_880), .B0 (n_3204), .Y (n_3404));
OAI21X1 g64546(.A0 (n_2366), .A1 (n_888), .B0 (n_3202), .Y (n_3403));
OAI21X1 g64549(.A0 (n_2368), .A1 (n_977), .B0 (n_3201), .Y (n_3402));
OAI21X1 g64566(.A0 (n_2367), .A1 (n_838), .B0 (n_3200), .Y (n_3400));
INVX1 g64571(.A (n_8707), .Y (n_3399));
AND2X1 g64600(.A (n_3398), .B (n_6972), .Y (n_3758));
OAI21X1 g64613(.A0 (n_2365), .A1 (n_881), .B0 (n_3206), .Y (n_3395));
INVX1 g64620(.A (n_3784), .Y (n_3394));
INVX2 g64641(.A (n_3547), .Y (n_3605));
CLKBUFX1 gbuf_d_931(.A(n_2712), .Y(d_out_931));
CLKBUFX1 gbuf_q_931(.A(q_in_931), .Y(g6159));
NAND2X1 g64660(.A (n_3425), .B (n_3391), .Y (n_3822));
CLKBUFX1 gbuf_d_932(.A(n_2854), .Y(d_out_932));
CLKBUFX1 gbuf_q_932(.A(q_in_932), .Y(g3155));
AOI21X1 g64682(.A0 (n_1090), .A1 (n_1279), .B0 (n_3569), .Y (n_3390));
AOI21X1 g64689(.A0 (n_3177), .A1 (n_3388), .B0 (n_2628), .Y (n_3389));
NAND4X1 g64690(.A (n_1656), .B (n_3984), .C (n_10005), .D (g5029), .Y(n_3387));
NAND4X1 g64048(.A (n_2977), .B (n_2389), .C (n_2344), .D (n_2340), .Y(n_3385));
AOI22X1 g64703(.A0 (n_2610), .A1 (n_3383), .B0 (g1472), .B1 (n_9628),.Y (n_3384));
MX2X1 g64707(.A (n_1629), .B (n_2595), .S0 (n_4617), .Y (n_3382));
AOI22X1 g64787(.A0 (n_2361), .A1 (n_598), .B0 (n_3073), .B1 (n_653),.Y (n_3381));
CLKBUFX1 gbuf_d_933(.A(n_2863), .Y(d_out_933));
CLKBUFX1 gbuf_qn_933(.A(qn_in_933), .Y(g4581));
OAI21X1 g64843(.A0 (n_2575), .A1 (g2975), .B0 (n_9351), .Y (n_3377));
NAND2X1 g64918(.A (n_2880), .B (n_6406), .Y (n_3376));
NAND3X1 g61120(.A (n_3372), .B (n_2), .C (n_11041), .Y (n_3373));
AOI21X1 g65001(.A0 (g16775), .A1 (n_493), .B0 (n_2869), .Y (n_3371));
CLKBUFX1 gbuf_d_934(.A(n_2846), .Y(d_out_934));
CLKBUFX1 gbuf_q_934(.A(q_in_934), .Y(g_6701));
CLKBUFX1 gbuf_d_935(.A(n_2914), .Y(d_out_935));
CLKBUFX1 gbuf_q_935(.A(q_in_935), .Y(g5170));
AOI22X1 g65018(.A0 (n_2215), .A1 (n_3177), .B0 (g_22021), .B1(n_9193), .Y (n_3370));
CLKBUFX1 gbuf_d_936(.A(n_2903), .Y(d_out_936));
CLKBUFX1 gbuf_q_936(.A(q_in_936), .Y(g5527));
NAND3X1 g61122(.A (n_3123), .B (n_3364), .C (n_9664), .Y (n_3369));
AOI22X1 g65034(.A0 (n_2496), .A1 (n_3177), .B0 (g_18996), .B1(n_9599), .Y (n_3368));
CLKBUFX1 gbuf_d_937(.A(n_2709), .Y(d_out_937));
CLKBUFX1 gbuf_q_937(.A(q_in_937), .Y(g3119));
CLKBUFX1 gbuf_d_938(.A(n_2720), .Y(d_out_938));
CLKBUFX1 gbuf_q_938(.A(q_in_938), .Y(g5128));
CLKBUFX1 gbuf_d_939(.A(n_2858), .Y(d_out_939));
CLKBUFX1 gbuf_q_939(.A(q_in_939), .Y(g5857));
CLKBUFX1 gbuf_d_940(.A(n_2829), .Y(d_out_940));
CLKBUFX1 gbuf_qn_940(.A(qn_in_940), .Y(g_5156));
CLKBUFX1 gbuf_d_941(.A(n_2831), .Y(d_out_941));
CLKBUFX1 gbuf_qn_941(.A(qn_in_941), .Y(g_6579));
CLKBUFX1 gbuf_d_942(.A(n_2839), .Y(d_out_942));
CLKBUFX1 gbuf_qn_942(.A(qn_in_942), .Y(g_5508));
CLKBUFX1 gbuf_d_943(.A(n_2833), .Y(d_out_943));
CLKBUFX1 gbuf_qn_943(.A(qn_in_943), .Y(g_14965));
CLKBUFX1 gbuf_d_944(.A(n_2837), .Y(d_out_944));
CLKBUFX1 gbuf_qn_944(.A(qn_in_944), .Y(g_3861));
CLKBUFX1 gbuf_d_945(.A(n_2693), .Y(d_out_945));
CLKBUFX1 gbuf_qn_945(.A(qn_in_945), .Y(g3841));
AOI21X1 g61132(.A0 (n_3365), .A1 (n_3364), .B0 (n_2834), .Y (n_3366));
CLKBUFX1 gbuf_d_946(.A(n_2913), .Y(d_out_946));
CLKBUFX1 gbuf_q_946(.A(q_in_946), .Y(g5517));
CLKBUFX1 gbuf_d_947(.A(n_2955), .Y(d_out_947));
CLKBUFX1 gbuf_q_947(.A(q_in_947), .Y(g4462));
CLKBUFX1 gbuf_d_948(.A(n_2949), .Y(d_out_948));
CLKBUFX1 gbuf_q_948(.A(q_in_948), .Y(g4264));
CLKBUFX1 gbuf_d_949(.A(n_2827), .Y(d_out_949));
CLKBUFX1 gbuf_q_949(.A(q_in_949), .Y(g2704));
CLKBUFX1 gbuf_d_950(.A(n_2954), .Y(d_out_950));
CLKBUFX1 gbuf_q_950(.A(q_in_950), .Y(g5092));
CLKBUFX1 gbuf_d_951(.A(n_2947), .Y(d_out_951));
CLKBUFX1 gbuf_q_951(.A(q_in_951), .Y(g1548));
CLKBUFX1 gbuf_d_952(.A(n_2700), .Y(d_out_952));
CLKBUFX1 gbuf_qn_952(.A(qn_in_952), .Y(g3490));
AOI22X1 g61955(.A0 (n_2495), .A1 (n_2878), .B0 (g_20563), .B1(n_9129), .Y (n_3363));
AOI22X1 g65441(.A0 (n_2506), .A1 (n_1751), .B0 (g3522), .B1 (n_9129),.Y (n_3362));
AOI22X1 g65442(.A0 (n_2494), .A1 (n_1718), .B0 (g6565), .B1 (n_9491),.Y (n_3361));
AOI22X1 g65444(.A0 (n_2500), .A1 (n_1777), .B0 (g5527), .B1 (n_9129),.Y (n_3360));
OAI22X1 g65499(.A0 (n_2559), .A1 (g4297), .B0 (n_150), .B1 (n_9992),.Y (n_3359));
OAI21X1 g65529(.A0 (n_32), .A1 (n_9681), .B0 (n_2840), .Y (n_3358));
INVX1 g65534(.A (g2927), .Y (n_3357));
CLKBUFX1 gbuf_d_953(.A(n_2775), .Y(d_out_953));
CLKBUFX1 gbuf_qn_953(.A(qn_in_953), .Y(g2878));
CLKBUFX1 gbuf_d_954(.A(n_2766), .Y(d_out_954));
CLKBUFX1 gbuf_q_954(.A(q_in_954), .Y(g9617));
CLKBUFX1 gbuf_d_955(.A(n_2776), .Y(d_out_955));
CLKBUFX1 gbuf_q_955(.A(q_in_955), .Y(g8215));
CLKBUFX1 gbuf_d_956(.A(n_2765), .Y(d_out_956));
CLKBUFX1 gbuf_q_956(.A(q_in_956), .Y(g9682));
CLKBUFX1 gbuf_d_957(.A(n_2769), .Y(d_out_957));
CLKBUFX1 gbuf_q_957(.A(q_in_957), .Y(g8279));
CLKBUFX1 gbuf_d_958(.A(n_2772), .Y(d_out_958));
CLKBUFX1 gbuf_q_958(.A(q_in_958), .Y(g9743));
INVX1 g65551(.A (g_13901), .Y (n_3519));
CLKBUFX1 gbuf_d_959(.A(n_2777), .Y(d_out_959));
CLKBUFX1 gbuf_qn_959(.A(qn_in_959), .Y(g_11037));
CLKBUFX1 gbuf_d_960(.A(n_2770), .Y(d_out_960));
CLKBUFX1 gbuf_q_960(.A(q_in_960), .Y(g8344));
INVX1 g65567(.A (g2965), .Y (n_3356));
CLKBUFX1 gbuf_d_961(.A(n_2796), .Y(d_out_961));
CLKBUFX1 gbuf_q_961(.A(q_in_961), .Y(g2724));
CLKBUFX1 gbuf_d_962(.A(n_2789), .Y(d_out_962));
CLKBUFX1 gbuf_qn_962(.A(qn_in_962), .Y(g3003));
CLKBUFX1 gbuf_d_963(.A(n_2788), .Y(d_out_963));
CLKBUFX1 gbuf_q_963(.A(q_in_963), .Y(g4145));
CLKBUFX1 gbuf_d_964(.A(n_2793), .Y(d_out_964));
CLKBUFX1 gbuf_qn_964(.A(qn_in_964), .Y(g4164));
CLKBUFX1 gbuf_d_965(.A(n_2774), .Y(d_out_965));
CLKBUFX1 gbuf_q_965(.A(q_in_965), .Y(g1521));
CLKBUFX1 gbuf_d_966(.A(n_2725), .Y(d_out_966));
CLKBUFX1 gbuf_q_966(.A(q_in_966), .Y(g_19172));
CLKBUFX1 gbuf_d_967(.A(n_2705), .Y(d_out_967));
CLKBUFX1 gbuf_qn_967(.A(qn_in_967), .Y(g6187));
MX2X1 g63135(.A (n_7260), .B (n_2484), .S0 (n_9501), .Y (n_3355));
CLKBUFX1 gbuf_d_968(.A(n_2687), .Y(d_out_968));
CLKBUFX1 gbuf_qn_968(.A(qn_in_968), .Y(g3139));
CLKBUFX1 gbuf_d_969(.A(n_2690), .Y(d_out_969));
CLKBUFX1 gbuf_q_969(.A(q_in_969), .Y(g1442));
CLKBUFX1 gbuf_d_970(.A(n_2716), .Y(d_out_970));
CLKBUFX1 gbuf_q_970(.A(q_in_970), .Y(g5467));
CLKBUFX1 gbuf_d_971(.A(n_2703), .Y(d_out_971));
CLKBUFX1 gbuf_q_971(.A(q_in_971), .Y(g3462));
NAND2X1 g65986(.A (n_3071), .B (n_2862), .Y (n_3353));
CLKBUFX1 gbuf_d_972(.A(n_2759), .Y(d_out_972));
CLKBUFX1 gbuf_q_972(.A(q_in_972), .Y(g4269));
NOR2X1 g63226(.A (n_2580), .B (n_3651), .Y (n_3352));
AND2X1 g63231(.A (n_3651), .B (n_3332), .Y (n_3351));
NAND2X1 g63232(.A (n_3651), .B (n_3707), .Y (n_3350));
NAND2X1 g63233(.A (n_3651), .B (n_9493), .Y (n_3720));
CLKBUFX1 gbuf_d_973(.A(n_2787), .Y(d_out_973));
CLKBUFX1 gbuf_q_973(.A(q_in_973), .Y(g4093));
NAND4X1 g66084(.A (n_3181), .B (n_7247), .C (n_9940), .D (n_23), .Y(n_3349));
MX2X1 g61169(.A (g1521), .B (n_2475), .S0 (n_8955), .Y (n_3348));
CLKBUFX1 gbuf_d_974(.A(n_2707), .Y(d_out_974));
CLKBUFX1 gbuf_q_974(.A(q_in_974), .Y(g6505));
CLKBUFX1 gbuf_d_975(.A(n_2864), .Y(d_out_975));
CLKBUFX1 gbuf_q_975(.A(q_in_975), .Y(n_1214));
CLKBUFX1 gbuf_d_976(.A(n_2819), .Y(d_out_976));
CLKBUFX1 gbuf_qn_976(.A(qn_in_976), .Y(g23002));
AOI21X1 g61480(.A0 (n_2192), .A1 (n_129), .B0 (n_2791), .Y (n_3347));
INVX1 g66272(.A (g2715), .Y (n_3679));
XOR2X1 g63329(.A (n_2754), .B (n_8913), .Y (n_3346));
NAND2X1 g61494(.A (n_2488), .B (n_3316), .Y (n_3345));
NOR2X1 g66362(.A (n_11), .B (n_9359), .Y (n_3344));
NOR2X1 g66369(.A (n_5363), .B (n_9453), .Y (n_3343));
CLKBUFX1 gbuf_d_977(.A(n_2719), .Y(d_out_977));
CLKBUFX1 gbuf_qn_977(.A(qn_in_977), .Y(g5148));
CLKBUFX1 gbuf_d_978(.A(n_2753), .Y(d_out_978));
CLKBUFX1 gbuf_q_978(.A(q_in_978), .Y(n_7260));
NOR2X1 g66409(.A (n_596), .B (n_9398), .Y (n_3341));
NOR2X1 g66471(.A (n_571), .B (n_9453), .Y (n_3340));
NOR2X1 g66512(.A (n_118), .B (n_9398), .Y (n_3339));
CLKBUFX1 gbuf_d_979(.A(n_2894), .Y(d_out_979));
CLKBUFX1 gbuf_q_979(.A(q_in_979), .Y(g3522));
NOR2X1 g66528(.A (n_572), .B (n_9940), .Y (n_3337));
NOR2X1 g66558(.A (n_504), .B (n_9940), .Y (n_3336));
OR2X1 g66644(.A (g2759), .B (n_9359), .Y (n_3335));
INVX1 g63453(.A (n_3447), .Y (n_3334));
NAND2X1 g63455(.A (n_3332), .B (n_8913), .Y (n_3333));
NOR2X1 g63457(.A (n_3563), .B (n_9903), .Y (n_3331));
NAND3X1 g63475(.A (n_3149), .B (n_3148), .C (g2882), .Y (n_3330));
CLKBUFX1 gbuf_d_980(.A(n_2814), .Y(d_out_980));
CLKBUFX1 gbuf_q_980(.A(q_in_980), .Y(g2145));
AND2X1 g63513(.A (n_3563), .B (n_2465), .Y (n_3329));
NAND2X1 g63514(.A (n_3563), .B (n_11134), .Y (n_3328));
NAND2X1 g63515(.A (n_3563), .B (n_9553), .Y (n_3687));
NAND4X1 g63519(.A (n_2945), .B (n_1331), .C (n_10119), .D (n_2303),.Y (n_3327));
NAND4X1 g63531(.A (n_2660), .B (n_2209), .C (n_2135), .D (n_1701), .Y(n_3326));
NAND4X1 g63534(.A (n_2986), .B (n_2408), .C (n_2122), .D (n_1698), .Y(n_3325));
AOI21X1 g63540(.A0 (n_2468), .A1 (n_2451), .B0 (n_3323), .Y (n_3324));
OAI22X1 g64064(.A0 (n_2624), .A1 (n_9599), .B0 (n_2645), .B1(n_9811), .Y (n_3322));
AOI22X1 g63554(.A0 (n_2263), .A1 (n_8840), .B0 (g1189), .B1 (n_9193),.Y (n_3321));
OAI21X1 g64043(.A0 (n_719), .A1 (n_9311), .B0 (n_2740), .Y (n_3320));
OAI21X1 g64030(.A0 (n_2734), .A1 (n_9681), .B0 (n_2735), .Y (n_3319));
OAI21X1 g61550(.A0 (n_92), .A1 (n_9978), .B0 (n_3316), .Y (n_3317));
OAI22X1 g64063(.A0 (n_2398), .A1 (n_9269), .B0 (n_2647), .B1(n_9811), .Y (n_3315));
CLKBUFX1 gbuf_d_981(.A(n_2739), .Y(d_out_981));
CLKBUFX1 gbuf_q_981(.A(q_in_981), .Y(g1319));
CLKBUFX1 gbuf_d_982(.A(n_2822), .Y(d_out_982));
CLKBUFX1 gbuf_q_982(.A(q_in_982), .Y(g2860));
XOR2X1 g63646(.A (n_10188), .B (n_2723), .Y (n_3314));
OAI22X1 g64068(.A0 (n_2392), .A1 (n_9836), .B0 (n_2646), .B1(n_9811), .Y (n_3313));
NAND3X1 g61034(.A (n_6734), .B (n_1043), .C (n_9425), .Y (n_3312));
CLKBUFX1 gbuf_d_983(.A(n_2953), .Y(d_out_983));
CLKBUFX1 gbuf_q_983(.A(q_in_983), .Y(n_10129));
CLKBUFX1 gbuf_d_984(.A(n_2804), .Y(d_out_984));
CLKBUFX1 gbuf_q_984(.A(q_in_984), .Y(g4912));
CLKBUFX1 gbuf_d_985(.A(n_2802), .Y(d_out_985));
CLKBUFX1 gbuf_q_985(.A(q_in_985), .Y(g4927));
CLKBUFX1 gbuf_d_986(.A(n_2805), .Y(d_out_986));
CLKBUFX1 gbuf_q_986(.A(q_in_986), .Y(g2907));
CLKBUFX1 gbuf_d_987(.A(n_2860), .Y(d_out_987));
CLKBUFX1 gbuf_q_987(.A(q_in_987), .Y(g5164));
NOR2X1 g63866(.A (n_10532), .B (n_3310), .Y (n_3915));
AND2X1 g63867(.A (n_10115), .B (n_3310), .Y (n_3309));
NAND2X1 g61644(.A (n_2879), .B (n_2742), .Y (n_3308));
NAND2X1 g63902(.A (n_2465), .B (n_10188), .Y (n_3307));
NAND3X1 g63918(.A (n_6766), .B (n_1541), .C (n_9940), .Y (n_3305));
NOR2X1 g63934(.A (n_2749), .B (n_957), .Y (n_3303));
AOI21X1 g63969(.A0 (n_1789), .A1 (n_3031), .B0 (n_2741), .Y (n_3302));
CLKBUFX1 gbuf_d_988(.A(n_2896), .Y(d_out_988));
CLKBUFX1 gbuf_q_988(.A(q_in_988), .Y(g_22552));
OAI22X1 g64067(.A0 (n_2397), .A1 (n_9193), .B0 (n_2642), .B1(n_9311), .Y (n_3301));
INVX1 g63997(.A (n_8835), .Y (n_3477));
CLKBUFX1 gbuf_d_989(.A(n_2816), .Y(d_out_989));
CLKBUFX1 gbuf_q_989(.A(q_in_989), .Y(g2873));
CLKBUFX1 gbuf_d_990(.A(n_2801), .Y(d_out_990));
CLKBUFX1 gbuf_q_990(.A(q_in_990), .Y(g4427));
OAI21X1 g64025(.A0 (n_1695), .A1 (n_9425), .B0 (n_2736), .Y (n_3300));
OAI21X1 g64027(.A0 (n_2421), .A1 (n_9940), .B0 (n_2733), .Y (n_3299));
OAI21X1 g64028(.A0 (n_11150), .A1 (n_9422), .B0 (n_2730), .Y(n_3298));
OAI21X1 g64029(.A0 (n_11173), .A1 (n_9333), .B0 (n_2727), .Y(n_3296));
CLKBUFX1 gbuf_d_991(.A(n_2886), .Y(d_out_991));
CLKBUFX1 gbuf_q_991(.A(q_in_991), .Y(g1189));
CLKBUFX1 gbuf_d_992(.A(n_2694), .Y(d_out_992));
CLKBUFX1 gbuf_q_992(.A(q_in_992), .Y(g3821));
CLKBUFX1 gbuf_d_993(.A(n_2761), .Y(d_out_993));
CLKBUFX1 gbuf_q_993(.A(q_in_993), .Y(g5097));
CLKBUFX1 gbuf_d_994(.A(n_2760), .Y(d_out_994));
CLKBUFX1 gbuf_q_994(.A(q_in_994), .Y(g1221));
CLKBUFX1 gbuf_d_995(.A(n_2758), .Y(d_out_995));
CLKBUFX1 gbuf_q_995(.A(q_in_995), .Y(g1564));
CLKBUFX1 gbuf_d_996(.A(n_2722), .Y(d_out_996));
CLKBUFX1 gbuf_q_996(.A(q_in_996), .Y(g5120));
CLKBUFX1 gbuf_d_997(.A(n_2715), .Y(d_out_997));
CLKBUFX1 gbuf_q_997(.A(q_in_997), .Y(g5475));
CLKBUFX1 gbuf_d_998(.A(n_2713), .Y(d_out_998));
CLKBUFX1 gbuf_q_998(.A(q_in_998), .Y(g5821));
CLKBUFX1 gbuf_d_999(.A(n_2714), .Y(d_out_999));
CLKBUFX1 gbuf_q_999(.A(q_in_999), .Y(g5813));
CLKBUFX1 gbuf_d_1000(.A(n_2706), .Y(d_out_1000));
CLKBUFX1 gbuf_q_1000(.A(q_in_1000), .Y(g6513));
CLKBUFX1 gbuf_d_1001(.A(n_2695), .Y(d_out_1001));
CLKBUFX1 gbuf_q_1001(.A(q_in_1001), .Y(g3813));
CLKBUFX1 gbuf_d_1002(.A(n_2691), .Y(d_out_1002));
CLKBUFX1 gbuf_q_1002(.A(q_in_1002), .Y(g_18635));
CLKBUFX1 gbuf_d_1003(.A(n_2689), .Y(d_out_1003));
CLKBUFX1 gbuf_q_1003(.A(q_in_1003), .Y(g8839));
CLKBUFX1 gbuf_d_1004(.A(n_2688), .Y(d_out_1004));
CLKBUFX1 gbuf_q_1004(.A(q_in_1004), .Y(n_2005));
CLKBUFX1 gbuf_d_1005(.A(n_2682), .Y(d_out_1005));
CLKBUFX1 gbuf_q_1005(.A(q_in_1005), .Y(g9251));
CLKBUFX1 gbuf_d_1006(.A(n_2951), .Y(d_out_1006));
CLKBUFX1 gbuf_q_1006(.A(q_in_1006), .Y(g_20952));
CLKBUFX1 gbuf_d_1007(.A(n_2904), .Y(d_out_1007));
CLKBUFX1 gbuf_q_1007(.A(q_in_1007), .Y(g5180));
CLKBUFX1 gbuf_d_1008(.A(n_2906), .Y(d_out_1008));
CLKBUFX1 gbuf_q_1008(.A(q_in_1008), .Y(g5863));
CLKBUFX1 gbuf_d_1009(.A(n_2897), .Y(d_out_1009));
CLKBUFX1 gbuf_q_1009(.A(q_in_1009), .Y(g3171));
CLKBUFX1 gbuf_d_1010(.A(n_2898), .Y(d_out_1010));
CLKBUFX1 gbuf_q_1010(.A(q_in_1010), .Y(g6219));
CLKBUFX1 gbuf_d_1011(.A(n_2888), .Y(d_out_1011));
CLKBUFX1 gbuf_q_1011(.A(q_in_1011), .Y(g6565));
CLKBUFX1 gbuf_d_1012(.A(n_2910), .Y(d_out_1012));
CLKBUFX1 gbuf_q_1012(.A(q_in_1012), .Y(g3512));
CLKBUFX1 gbuf_d_1013(.A(n_2907), .Y(d_out_1013));
CLKBUFX1 gbuf_q_1013(.A(q_in_1013), .Y(g3863));
CLKBUFX1 gbuf_d_1014(.A(n_2892), .Y(d_out_1014));
CLKBUFX1 gbuf_q_1014(.A(q_in_1014), .Y(g3873));
CLKBUFX1 gbuf_d_1015(.A(n_2909), .Y(d_out_1015));
CLKBUFX1 gbuf_q_1015(.A(q_in_1015), .Y(g3161));
CLKBUFX1 gbuf_d_1016(.A(n_2889), .Y(d_out_1016));
CLKBUFX1 gbuf_q_1016(.A(q_in_1016), .Y(g1532));
CLKBUFX1 gbuf_d_1017(.A(n_2887), .Y(d_out_1017));
CLKBUFX1 gbuf_q_1017(.A(q_in_1017), .Y(g1178));
CLKBUFX1 gbuf_d_1018(.A(n_2911), .Y(d_out_1018));
CLKBUFX1 gbuf_q_1018(.A(q_in_1018), .Y(g6555));
OAI22X1 g64082(.A0 (n_2625), .A1 (n_10078), .B0 (n_2644), .B1(n_10063), .Y (n_3292));
CLKBUFX1 gbuf_d_1019(.A(n_2821), .Y(d_out_1019));
CLKBUFX1 gbuf_q_1019(.A(q_in_1019), .Y(g2844));
CLKBUFX1 gbuf_d_1020(.A(n_2826), .Y(d_out_1020));
CLKBUFX1 gbuf_q_1020(.A(q_in_1020), .Y(g2852));
CLKBUFX1 gbuf_d_1021(.A(n_2856), .Y(d_out_1021));
CLKBUFX1 gbuf_q_1021(.A(q_in_1021), .Y(g5511));
CLKBUFX1 gbuf_d_1022(.A(n_2820), .Y(d_out_1022));
CLKBUFX1 gbuf_q_1022(.A(q_in_1022), .Y(g2894));
CLKBUFX1 gbuf_d_1023(.A(n_2824), .Y(d_out_1023));
CLKBUFX1 gbuf_q_1023(.A(q_in_1023), .Y(g2950));
CLKBUFX1 gbuf_d_1024(.A(n_2843), .Y(d_out_1024));
CLKBUFX1 gbuf_q_1024(.A(q_in_1024), .Y(g6549));
CLKBUFX1 gbuf_d_1025(.A(n_2810), .Y(d_out_1025));
CLKBUFX1 gbuf_q_1025(.A(q_in_1025), .Y(g20652));
CLKBUFX1 gbuf_d_1026(.A(n_2850), .Y(d_out_1026));
CLKBUFX1 gbuf_q_1026(.A(q_in_1026), .Y(g3506));
CLKBUFX1 gbuf_d_1027(.A(n_2807), .Y(d_out_1027));
CLKBUFX1 gbuf_q_1027(.A(q_in_1027), .Y(g2697));
CLKBUFX1 gbuf_d_1028(.A(n_2762), .Y(d_out_1028));
CLKBUFX1 gbuf_q_1028(.A(q_in_1028), .Y(g2988));
CLKBUFX1 gbuf_d_1029(.A(n_2848), .Y(d_out_1029));
CLKBUFX1 gbuf_q_1029(.A(q_in_1029), .Y(g3857));
CLKBUFX1 gbuf_d_1030(.A(n_2815), .Y(d_out_1030));
CLKBUFX1 gbuf_q_1030(.A(q_in_1030), .Y(g2138));
CLKBUFX1 gbuf_d_1031(.A(n_2832), .Y(d_out_1031));
CLKBUFX1 gbuf_q_1031(.A(q_in_1031), .Y(g4157));
CLKBUFX1 gbuf_d_1032(.A(n_2813), .Y(d_out_1032));
CLKBUFX1 gbuf_q_1032(.A(q_in_1032), .Y(g4245));
CLKBUFX1 gbuf_d_1033(.A(n_2812), .Y(d_out_1033));
CLKBUFX1 gbuf_q_1033(.A(q_in_1033), .Y(g4253));
CLKBUFX1 gbuf_d_1034(.A(n_2808), .Y(d_out_1034));
CLKBUFX1 gbuf_q_1034(.A(q_in_1034), .Y(g2970));
CLKBUFX1 gbuf_d_1035(.A(n_2817), .Y(d_out_1035));
CLKBUFX1 gbuf_q_1035(.A(q_in_1035), .Y(g2960));
CLKBUFX1 gbuf_d_1036(.A(n_2806), .Y(d_out_1036));
CLKBUFX1 gbuf_q_1036(.A(q_in_1036), .Y(g4732));
CLKBUFX1 gbuf_d_1037(.A(n_2823), .Y(d_out_1037));
CLKBUFX1 gbuf_q_1037(.A(q_in_1037), .Y(g4737));
CLKBUFX1 gbuf_d_1038(.A(n_2803), .Y(d_out_1038));
CLKBUFX1 gbuf_q_1038(.A(q_in_1038), .Y(g4922));
CLKBUFX1 gbuf_d_1039(.A(n_2767), .Y(d_out_1039));
CLKBUFX1 gbuf_q_1039(.A(q_in_1039), .Y(g4098));
CLKBUFX1 gbuf_d_1040(.A(n_2768), .Y(d_out_1040));
CLKBUFX1 gbuf_q_1040(.A(q_in_1040), .Y(g_22349));
CLKBUFX1 gbuf_d_1041(.A(n_2782), .Y(d_out_1041));
CLKBUFX1 gbuf_q_1041(.A(q_in_1041), .Y(g4258));
CLKBUFX1 gbuf_d_1042(.A(n_2956), .Y(d_out_1042));
CLKBUFX1 gbuf_q_1042(.A(q_in_1042), .Y(g10306));
NAND2X1 g64149(.A (n_3291), .B (g_13278), .Y (n_3690));
OAI21X1 g64153(.A0 (n_2616), .A1 (n_890), .B0 (n_2974), .Y (n_3290));
NOR2X1 g64155(.A (n_2675), .B (n_6694), .Y (n_3289));
OAI21X1 g61061(.A0 (n_2938), .A1 (n_3183), .B0 (n_10005), .Y(n_3288));
AND2X1 g64158(.A (n_2663), .B (n_3025), .Y (n_3287));
NAND4X1 g64166(.A (g5220), .B (n_10621), .C (n_1695), .D (g5339), .Y(n_3286));
CLKBUFX1 gbuf_d_1043(.A(n_2915), .Y(d_out_1043));
CLKBUFX1 gbuf_q_1043(.A(q_in_1043), .Y(g2980));
NAND4X1 g64181(.A (n_2673), .B (n_512), .C (n_448), .D (n_262), .Y(n_3285));
NAND2X2 g64233(.A (n_3236), .B (n_2039), .Y (n_3814));
NAND3X1 g64235(.A (n_2666), .B (n_2486), .C (n_2400), .Y (n_3283));
NAND3X1 g64236(.A (n_2665), .B (n_2536), .C (n_2634), .Y (n_3282));
NAND4X1 g64256(.A (g5567), .B (n_7150), .C (n_2208), .D (g5685), .Y(n_3281));
NAND3X1 g61726(.A (n_2972), .B (n_2530), .C (n_2603), .Y (n_3279));
NAND4X1 g64257(.A (g6259), .B (n_3277), .C (n_11150), .D (g6377), .Y(n_3278));
NAND4X1 g64275(.A (g6605), .B (n_3275), .C (n_11173), .D (g6723), .Y(n_3276));
AND2X1 g64278(.A (n_10693), .B (n_2077), .Y (n_3829));
NOR2X1 g64315(.A (n_2664), .B (n_2866), .Y (n_3274));
NAND3X1 g64039(.A (n_2658), .B (n_2548), .C (n_2459), .Y (n_3273));
AOI21X1 g64361(.A0 (n_2679), .A1 (n_10134), .B0 (n_2680), .Y(n_3271));
OAI21X1 g64365(.A0 (n_23), .A1 (n_9422), .B0 (n_2981), .Y (n_3270));
NAND4X1 g64376(.A (n_10831), .B (g5204), .C (g25219), .D (g5339), .Y(n_3269));
NAND4X1 g64382(.A (n_2439), .B (g5551), .C (n_1023), .D (g5685), .Y(n_3268));
NAND4X1 g64383(.A (n_2413), .B (g6243), .C (n_11157), .D (g6377), .Y(n_3267));
NAND4X1 g64384(.A (n_10809), .B (g5897), .C (n_546), .D (g6031), .Y(n_3266));
NAND4X1 g64385(.A (n_2435), .B (g6589), .C (n_11177), .D (g6723), .Y(n_3265));
NAND4X1 g64387(.A (n_2042), .B (n_3984), .C (g5041), .D (n_10771), .Y(n_3264));
OAI21X1 g62646(.A0 (n_307), .A1 (n_9333), .B0 (n_2946), .Y (n_3263));
CLKBUFX1 gbuf_d_1044(.A(n_2685), .Y(d_out_1044));
CLKBUFX1 gbuf_qn_1044(.A(qn_in_1044), .Y(g5841));
NOR2X1 g62649(.A (n_2662), .B (g3343), .Y (n_3262));
NOR2X1 g62651(.A (n_2669), .B (g3694), .Y (n_3261));
XOR2X1 g64402(.A (n_2637), .B (n_3259), .Y (n_3260));
CLKBUFX1 gbuf_d_1045(.A(n_2900), .Y(d_out_1045));
CLKBUFX1 gbuf_q_1045(.A(q_in_1045), .Y(g5873));
CLKBUFX1 gbuf_d_1046(.A(n_2702), .Y(d_out_1046));
CLKBUFX1 gbuf_q_1046(.A(q_in_1046), .Y(g3470));
INVX1 g64411(.A (n_3258), .Y (n_3645));
AOI22X1 g64414(.A0 (n_2410), .A1 (n_8637), .B0 (n_3152), .B1 (n_644),.Y (n_3257));
OAI21X1 g62658(.A0 (n_1295), .A1 (n_9940), .B0 (n_2939), .Y (n_3255));
MX2X1 g64437(.A (n_3253), .B (n_1802), .S0 (n_9627), .Y (n_3254));
CLKBUFX1 gbuf_d_1047(.A(n_2905), .Y(d_out_1047));
CLKBUFX1 gbuf_q_1047(.A(q_in_1047), .Y(g5069));
CLKBUFX1 gbuf_d_1048(.A(n_2902), .Y(d_out_1048));
CLKBUFX1 gbuf_qn_1048(.A(qn_in_1048), .Y(g2932));
CLKBUFX1 gbuf_d_1049(.A(n_2890), .Y(d_out_1049));
CLKBUFX1 gbuf_qn_1049(.A(qn_in_1049), .Y(g4284));
CLKBUFX1 gbuf_d_1050(.A(n_2895), .Y(d_out_1050));
CLKBUFX1 gbuf_q_1050(.A(q_in_1050), .Y(g2946));
NOR2X1 g64509(.A (n_3569), .B (g_22639), .Y (n_3566));
INVX2 g64537(.A (n_3249), .Y (n_3775));
NAND3X1 g64551(.A (n_2654), .B (n_10664), .C (n_9717), .Y (n_3247));
CLKBUFX1 gbuf_d_1051(.A(n_2948), .Y(d_out_1051));
CLKBUFX1 gbuf_q_1051(.A(q_in_1051), .Y(g_16404));
INVX2 g64569(.A (g28753), .Y (n_3244));
NOR2X1 g64575(.A (n_3486), .B (n_2828), .Y (n_3243));
CLKBUFX1 gbuf_d_1052(.A(n_2912), .Y(d_out_1052));
CLKBUFX1 gbuf_q_1052(.A(q_in_1052), .Y(g6209));
NAND2X1 g64579(.A (n_3569), .B (g_19113), .Y (n_3242));
NAND3X1 g64580(.A (n_835), .B (n_2609), .C (n_9558), .Y (n_3241));
INVX4 g64587(.A (n_3239), .Y (n_3779));
INVX1 g64634(.A (n_4053), .Y (n_4832));
CLKBUFX1 g64642(.A (n_3236), .Y (n_3547));
NAND2X1 g64645(.A (n_3224), .B (n_659), .Y (n_3234));
NOR3X1 g64648(.A (n_3016), .B (g5037), .C (n_9107), .Y (n_3233));
INVX1 g64650(.A (n_10461), .Y (n_3832));
NAND4X1 g64656(.A (n_1643), .B (n_1084), .C (n_9521), .D (n_2881), .Y(n_3229));
NAND4X1 g64657(.A (n_1642), .B (n_1085), .C (n_9501), .D (n_3171), .Y(n_3228));
NAND4X1 g64659(.A (n_1381), .B (n_842), .C (n_9139), .D (n_2732), .Y(n_3226));
NAND4X1 g64661(.A (n_1641), .B (n_1083), .C (n_9091), .D (n_2729), .Y(n_3225));
NAND2X1 g64686(.A (n_3224), .B (n_3391), .Y (n_3438));
NAND4X1 g64688(.A (n_1640), .B (n_1082), .C (n_9091), .D (n_2871), .Y(n_3223));
NAND3X1 g61809(.A (n_851), .B (n_1996), .C (n_10949), .Y (n_3222));
NAND3X1 g61812(.A (n_722), .B (n_1647), .C (n_10949), .Y (n_3221));
NAND4X1 g64731(.A (n_2447), .B (g3953), .C (g16659), .D (n_4988), .Y(n_3219));
NAND4X1 g64772(.A (n_7010), .B (n_1493), .C (g5033), .D (n_3984), .Y(n_3218));
MX2X1 g64781(.A (g4888), .B (g4894), .S0 (n_2351), .Y (n_3217));
CLKBUFX1 gbuf_d_1053(.A(g16624), .Y(d_out_1053));
CLKBUFX1 gbuf_q_1053(.A(q_in_1053), .Y(g14421));
CLKBUFX1 gbuf_d_1054(.A(g16656), .Y(d_out_1054));
CLKBUFX1 gbuf_q_1054(.A(q_in_1054), .Y(g14451));
NAND3X1 g64853(.A (n_2883), .B (g_18996), .C (n_9681), .Y (n_3216));
AND2X1 g64892(.A (n_10897), .B (g16656), .Y (n_3398));
NAND2X1 g64898(.A (n_10400), .B (g4311), .Y (n_3258));
NAND3X1 g64903(.A (n_2055), .B (n_3213), .C (n_276), .Y (n_3214));
AND2X1 g64912(.A (n_2614), .B (g4633), .Y (n_3212));
NOR2X1 g64924(.A (n_3641), .B (n_6400), .Y (n_3211));
NAND2X1 g64939(.A (g16624), .B (g16603), .Y (n_3210));
NAND2X1 g64941(.A (g16656), .B (g16627), .Y (n_3209));
NOR2X1 g64964(.A (n_2602), .B (n_10296), .Y (n_3208));
INVX1 g61116(.A (n_3910), .Y (n_4866));
AOI22X1 g64986(.A0 (n_2218), .A1 (n_4327), .B0 (n_1807), .B1(n_9193), .Y (n_3207));
AOI22X1 g64988(.A0 (n_2206), .A1 (n_4324), .B0 (n_2084), .B1(n_9599), .Y (n_3206));
AOI22X1 g64989(.A0 (n_2227), .A1 (n_4316), .B0 (n_1805), .B1(n_9193), .Y (n_3204));
AOI22X1 g64992(.A0 (n_2204), .A1 (n_4322), .B0 (n_1794), .B1(n_10376), .Y (n_3202));
AOI22X1 g64995(.A0 (n_2207), .A1 (n_4320), .B0 (n_1799), .B1(n_9526), .Y (n_3201));
AOI22X1 g64998(.A0 (n_2211), .A1 (n_4314), .B0 (n_1796), .B1(n_9193), .Y (n_3200));
AOI22X1 g65002(.A0 (n_2205), .A1 (n_1422), .B0 (g1442), .B1 (n_9300),.Y (n_3197));
AOI22X1 g65004(.A0 (n_2210), .A1 (n_2008), .B0 (g1478), .B1 (n_9672),.Y (n_3196));
AOI22X1 g65005(.A0 (n_2228), .A1 (n_4329), .B0 (n_1810), .B1(n_9193), .Y (n_3194));
MX2X1 g62926(.A (n_2305), .B (n_3192), .S0 (n_2166), .Y (n_3193));
AOI22X1 g65006(.A0 (n_2216), .A1 (n_1252), .B0 (g1448), .B1 (n_9300),.Y (n_3191));
AOI22X1 g65019(.A0 (n_2276), .A1 (n_1655), .B0 (n_10134), .B1(n_9129), .Y (n_3189));
NAND3X1 g61121(.A (g1384), .B (n_2830), .C (n_9558), .Y (n_3187));
NAND2X1 g61369(.A (n_2671), .B (n_2563), .Y (n_3186));
OAI21X1 g65052(.A0 (n_3184), .A1 (n_10524), .B0 (n_2611), .Y(n_3185));
AND2X1 g61123(.A (n_1503), .B (n_3183), .Y (n_3628));
AOI22X1 g65058(.A0 (n_2316), .A1 (n_3181), .B0 (n_7247), .B1(n_9491), .Y (n_3182));
OAI21X1 g61372(.A0 (g1585), .A1 (n_9797), .B0 (n_3165), .Y (n_3179));
AOI22X1 g65084(.A0 (n_1221), .A1 (n_2577), .B0 (n_3177), .B1(n_10528), .Y (n_3178));
MX2X1 g65107(.A (n_2017), .B (n_2320), .S0 (n_9000), .Y (n_3176));
MX2X1 g64084(.A (g_18795), .B (g_17934), .S0 (n_3174), .Y (n_3175));
CLKBUFX1 gbuf_d_1055(.A(g16659), .Y(d_out_1055));
CLKBUFX1 gbuf_q_1055(.A(q_in_1055), .Y(g16693));
OR2X1 g65275(.A (n_3171), .B (n_3121), .Y (n_3172));
NAND3X1 g61927(.A (n_1646), .B (g_20563), .C (n_9698), .Y (n_3170));
OAI21X1 g61399(.A0 (g1579), .A1 (n_9425), .B0 (n_3165), .Y (n_3167));
AOI21X1 g61952(.A0 (g_19172), .A1 (n_9775), .B0 (n_2574), .Y(n_3164));
AOI21X1 g61953(.A0 (g_11413), .A1 (n_9775), .B0 (n_2573), .Y(n_3162));
AOI21X1 g61954(.A0 (g_16456), .A1 (n_9884), .B0 (n_2572), .Y(n_3161));
AOI22X1 g65437(.A0 (n_2233), .A1 (n_1762), .B0 (g5180), .B1 (n_9129),.Y (n_3160));
AOI22X1 g65438(.A0 (n_2223), .A1 (n_1725), .B0 (g5873), .B1(n_10376), .Y (n_3158));
AOI22X1 g65440(.A0 (n_2219), .A1 (n_1723), .B0 (g6219), .B1 (n_9129),.Y (n_3157));
AOI22X1 g65443(.A0 (n_2225), .A1 (n_1743), .B0 (g3873), .B1 (n_9129),.Y (n_3156));
AOI22X1 g65446(.A0 (n_2203), .A1 (n_1758), .B0 (g3171), .B1 (n_9107),.Y (n_3154));
NAND4X1 g61957(.A (n_2867), .B (n_3152), .C (n_9359), .D (g4669), .Y(n_3153));
OR2X1 g63963(.A (n_3149), .B (n_3148), .Y (g26877));
OAI22X1 g65493(.A0 (n_2859), .A1 (n_1464), .B0 (n_621), .B1(n_10063), .Y (n_3147));
OAI22X1 g65494(.A0 (n_2855), .A1 (n_673), .B0 (n_686), .B1 (n_9830),.Y (n_3146));
OAI22X1 g65495(.A0 (n_2853), .A1 (n_1482), .B0 (n_623), .B1 (n_9830),.Y (n_3145));
OAI22X1 g65496(.A0 (n_2842), .A1 (n_1486), .B0 (n_603), .B1 (n_9830),.Y (n_3144));
MX2X1 g63084(.A (g5097), .B (n_2182), .S0 (n_10005), .Y (n_3143));
OAI22X1 g65497(.A0 (n_2849), .A1 (n_463), .B0 (n_664), .B1 (n_9992),.Y (n_3142));
OAI22X1 g65498(.A0 (n_2847), .A1 (n_458), .B0 (n_678), .B1 (n_9830),.Y (n_3141));
OAI22X1 g65501(.A0 (n_2857), .A1 (n_1459), .B0 (n_627), .B1(n_10063), .Y (n_3140));
MX2X1 g65530(.A (n_511), .B (g2980), .S0 (n_9269), .Y (n_3139));
MX2X1 g65531(.A (n_1633), .B (g_21651), .S0 (n_9599), .Y (n_3138));
MX2X1 g65532(.A (n_826), .B (n_6958), .S0 (n_9599), .Y (n_3137));
MX2X1 g65533(.A (n_209), .B (n_3135), .S0 (n_9599), .Y (n_3136));
CLKBUFX1 gbuf_d_1056(.A(n_2509), .Y(d_out_1056));
CLKBUFX1 gbuf_qn_1056(.A(qn_in_1056), .Y(g2927));
CLKBUFX1 gbuf_d_1057(.A(n_2517), .Y(d_out_1057));
CLKBUFX1 gbuf_q_1057(.A(q_in_1057), .Y(g9555));
CLKBUFX1 gbuf_d_1058(.A(n_2507), .Y(d_out_1058));
CLKBUFX1 gbuf_q_1058(.A(q_in_1058), .Y(g_13901));
CLKBUFX1 gbuf_d_1059(.A(n_2501), .Y(d_out_1059));
CLKBUFX1 gbuf_q_1059(.A(q_in_1059), .Y(g14189));
CLKBUFX1 gbuf_d_1060(.A(n_2499), .Y(d_out_1060));
CLKBUFX1 gbuf_qn_1060(.A(qn_in_1060), .Y(g2965));
NOR2X1 g65624(.A (n_205), .B (n_9836), .Y (n_3133));
NOR2X1 g65641(.A (n_311), .B (n_9353), .Y (n_3132));
MX2X1 g63134(.A (g4269), .B (n_2181), .S0 (n_9000), .Y (n_3131));
NOR3X1 g65891(.A (n_276), .B (n_7247), .C (n_9505), .Y (n_3130));
NOR3X1 g65901(.A (n_11113), .B (n_9775), .C (g8719), .Y (n_3127));
INVX1 g61165(.A (n_3123), .Y (n_3124));
OAI21X1 g66057(.A0 (n_379), .A1 (n_9425), .B0 (n_3121), .Y (n_3122));
OAI21X1 g66063(.A0 (n_87), .A1 (n_9333), .B0 (n_2612), .Y (n_3120));
OAI21X1 g66066(.A0 (n_93), .A1 (n_9681), .B0 (n_3117), .Y (n_3119));
OAI21X1 g66067(.A0 (n_89), .A1 (n_9681), .B0 (n_3115), .Y (n_3116));
OAI21X1 g66068(.A0 (n_13), .A1 (n_9311), .B0 (n_3113), .Y (n_3114));
OAI21X1 g66078(.A0 (n_59), .A1 (n_9333), .B0 (n_2668), .Y (n_3112));
MX2X1 g66098(.A (g1798), .B (n_5996), .S0 (n_9269), .Y (n_3111));
MX2X1 g66099(.A (g1644), .B (g1592), .S0 (n_9599), .Y (n_3109));
MX2X1 g66105(.A (g2223), .B (n_5941), .S0 (n_9599), .Y (n_3108));
MX2X1 g66107(.A (g1913), .B (g1862), .S0 (n_9672), .Y (n_3106));
MX2X1 g66108(.A (g2912), .B (g2907), .S0 (n_9628), .Y (n_3105));
MX2X1 g66109(.A (g2994), .B (g2999), .S0 (n_9599), .Y (n_3104));
MX2X1 g66110(.A (g2204), .B (g2153), .S0 (n_9672), .Y (n_3103));
MX2X1 g66111(.A (g21292), .B (g_18015), .S0 (n_9269), .Y (n_3102));
MX2X1 g66112(.A (g2625), .B (n_5928), .S0 (n_9599), .Y (n_3100));
MX2X1 g66115(.A (g2047), .B (g1996), .S0 (n_9672), .Y (n_3099));
MX2X1 g66116(.A (g2066), .B (n_5932), .S0 (n_9628), .Y (n_3098));
MX2X1 g66117(.A (g1779), .B (g1728), .S0 (n_9019), .Y (n_3097));
MX2X1 g66122(.A (g2868), .B (g2988), .S0 (n_9599), .Y (n_3096));
MX2X1 g66123(.A (g4146), .B (g4176), .S0 (n_9269), .Y (n_3095));
MX2X1 g66127(.A (g4249), .B (g4253), .S0 (n_9269), .Y (n_3094));
MX2X1 g66130(.A (g4907), .B (g4922), .S0 (n_9599), .Y (n_3092));
MX2X1 g66132(.A (g2338), .B (g2287), .S0 (n_9672), .Y (n_3091));
MX2X1 g66134(.A (g2936), .B (g2922), .S0 (n_9599), .Y (n_3090));
MX2X1 g66135(.A (g4717), .B (g4732), .S0 (n_9269), .Y (n_3088));
MX2X1 g66136(.A (g4722), .B (g4717), .S0 (n_9269), .Y (n_3087));
MX2X1 g66139(.A (g1664), .B (n_5936), .S0 (n_9599), .Y (n_3086));
MX2X1 g66140(.A (g2357), .B (n_5917), .S0 (n_9599), .Y (n_3085));
MX2X1 g66141(.A (g2472), .B (g2421), .S0 (n_9019), .Y (n_3084));
MX2X1 g66142(.A (g2491), .B (n_5921), .S0 (n_9599), .Y (n_3082));
MX2X1 g66144(.A (g2922), .B (g2912), .S0 (n_9269), .Y (n_3081));
MX2X1 g66146(.A (g1932), .B (n_5925), .S0 (n_9599), .Y (n_3080));
MX2X1 g66149(.A (g2606), .B (g2555), .S0 (n_9628), .Y (n_3079));
MX2X1 g66154(.A (n_150), .B (g4273), .S0 (n_9019), .Y (n_3077));
XOR2X1 g61485(.A (n_8508), .B (n_2790), .Y (n_3075));
NAND4X1 g62097(.A (n_2925), .B (n_3073), .C (n_9139), .D (n_11216),.Y (n_3074));
INVX1 g66410(.A (n_3071), .Y (n_3072));
NOR2X1 g66656(.A (n_10956), .B (n_9353), .Y (n_3070));
AND2X1 g63454(.A (n_3431), .B (g_19414), .Y (n_3447));
CLKBUFX1 gbuf_d_1061(.A(n_2512), .Y(d_out_1061));
CLKBUFX1 gbuf_q_1061(.A(q_in_1061), .Y(g4917));
CLKBUFX1 gbuf_d_1062(.A(n_2493), .Y(d_out_1062));
CLKBUFX1 gbuf_q_1062(.A(q_in_1062), .Y(g2890));
CLKBUFX1 gbuf_d_1063(.A(n_2498), .Y(d_out_1063));
CLKBUFX1 gbuf_q_1063(.A(q_in_1063), .Y(g4108));
CLKBUFX1 gbuf_d_1064(.A(n_2510), .Y(d_out_1064));
CLKBUFX1 gbuf_q_1064(.A(q_in_1064), .Y(g2759));
CLKBUFX1 gbuf_d_1065(.A(n_2503), .Y(d_out_1065));
CLKBUFX1 gbuf_q_1065(.A(q_in_1065), .Y(g4082));
OAI21X1 g63606(.A0 (n_3065), .A1 (n_7383), .B0 (n_2237), .Y (n_3066));
OAI21X1 g63614(.A0 (n_3062), .A1 (n_10889), .B0 (n_2264), .Y(n_3063));
CLKBUFX1 gbuf_d_1066(.A(n_2491), .Y(d_out_1066));
CLKBUFX1 gbuf_q_1066(.A(q_in_1066), .Y(g2735));
CLKBUFX1 gbuf_d_1067(.A(n_9453), .Y(d_out_1067));
CLKBUFX1 gbuf_qn_1067(.A(qn_in_1067), .Y(g2715));
OR2X1 g61032(.A (n_4241), .B (g1413), .Y (n_3059));
MX2X1 g63772(.A (g_18793), .B (n_503), .S0 (n_3661), .Y (n_3058));
MX2X1 g63786(.A (g_21806), .B (n_2160), .S0 (n_9469), .Y (n_3057));
MX2X1 g63789(.A (g_22379), .B (n_2159), .S0 (n_9558), .Y (n_3056));
MX2X1 g63790(.A (n_11162), .B (n_2157), .S0 (n_9091), .Y (n_3055));
MX2X1 g63803(.A (g_6131), .B (n_2156), .S0 (n_9172), .Y (n_3053));
MX2X1 g63805(.A (g_20837), .B (n_2155), .S0 (n_9874), .Y (n_3052));
XOR2X1 g63810(.A (n_640), .B (n_2167), .Y (n_3713));
NOR2X1 g63906(.A (n_2743), .B (n_7260), .Y (n_3491));
NAND2X1 g63913(.A (n_3036), .B (n_3035), .Y (n_3497));
NAND4X1 g63968(.A (n_3048), .B (n_965), .C (n_3047), .D (n_2153), .Y(n_3050));
NAND4X1 g63995(.A (n_3048), .B (n_1630), .C (n_3047), .D (n_1263), .Y(n_3049));
NAND4X1 g64046(.A (n_2121), .B (n_1696), .C (n_2038), .D (n_2031), .Y(n_3044));
MX2X1 g64085(.A (n_3042), .B (g_18795), .S0 (n_3174), .Y (n_3043));
MX2X1 g64087(.A (g_12433), .B (g_20073), .S0 (n_3174), .Y (n_3041));
CLKBUFX1 gbuf_d_1068(.A(n_2579), .Y(d_out_1068));
CLKBUFX1 gbuf_q_1068(.A(q_in_1068), .Y(g6203));
MX2X1 g64088(.A (n_10108), .B (n_3042), .S0 (n_3174), .Y (n_3040));
MX2X1 g64089(.A (g_20073), .B (n_10103), .S0 (n_3174), .Y (n_3038));
CLKBUFX1 gbuf_d_1069(.A(n_2492), .Y(d_out_1069));
CLKBUFX1 gbuf_q_1069(.A(q_in_1069), .Y(g4727));
CLKBUFX1 gbuf_d_1070(.A(n_2515), .Y(d_out_1070));
CLKBUFX1 gbuf_q_1070(.A(q_in_1070), .Y(n_11099));
CLKBUFX1 gbuf_d_1071(.A(n_2502), .Y(d_out_1071));
CLKBUFX1 gbuf_q_1071(.A(q_in_1071), .Y(g4076));
CLKBUFX1 gbuf_d_1072(.A(n_2504), .Y(d_out_1072));
CLKBUFX1 gbuf_q_1072(.A(q_in_1072), .Y(g2130));
CLKBUFX1 gbuf_d_1073(.A(n_2514), .Y(d_out_1073));
CLKBUFX1 gbuf_q_1073(.A(q_in_1073), .Y(g4104));
OR2X1 g63949(.A (n_3036), .B (n_3035), .Y (g26876));
CLKBUFX1 gbuf_d_1074(.A(n_2454), .Y(d_out_1074));
CLKBUFX1 gbuf_qn_1074(.A(qn_in_1074), .Y(g4072));
MX2X1 g64086(.A (g_17934), .B (g_22464), .S0 (n_3174), .Y (n_3034));
NAND2X1 g64211(.A (g_15287), .B (n_10751), .Y (n_3033));
NAND3X1 g64213(.A (n_3031), .B (n_3030), .C (n_1250), .Y (n_3032));
NAND2X1 g64226(.A (n_1542), .B (n_2656), .Y (n_3029));
NOR2X1 g64242(.A (n_2453), .B (g_18795), .Y (n_3028));
NAND4X1 g64314(.A (n_2980), .B (n_3181), .C (n_9209), .D (g4633), .Y(n_3027));
NAND4X1 g64326(.A (n_1788), .B (n_3030), .C (n_3025), .D (n_2114), .Y(n_3026));
NAND4X1 g64368(.A (n_3030), .B (n_1266), .C (n_3021), .D (n_2116), .Y(n_3022));
XOR2X1 g64372(.A (n_3065), .B (n_7383), .Y (n_3020));
XOR2X1 g64373(.A (n_3062), .B (n_10889), .Y (n_3019));
MX2X1 g61747(.A (g_18902), .B (n_2346), .S0 (n_10063), .Y (n_3018));
NAND4X1 g64386(.A (n_3016), .B (n_3984), .C (n_10385), .D (g5037), .Y(n_3017));
AOI21X1 g64394(.A0 (n_2458), .A1 (n_9505), .B0 (n_2655), .Y (n_3015));
XOR2X1 g64403(.A (n_2415), .B (n_3013), .Y (n_3014));
XOR2X1 g64409(.A (n_2082), .B (n_2373), .Y (n_3660));
MX2X1 g64430(.A (n_3011), .B (n_1811), .S0 (n_9894), .Y (n_3012));
MX2X1 g64436(.A (g6163), .B (n_2375), .S0 (n_9359), .Y (n_3010));
MX2X1 g64441(.A (n_3007), .B (n_1795), .S0 (n_9553), .Y (n_3008));
MX2X1 g64460(.A (g1178), .B (n_2374), .S0 (n_9333), .Y (n_3005));
NOR2X1 g64508(.A (n_3003), .B (g_16792), .Y (n_3004));
NOR2X1 g64523(.A (n_2629), .B (n_644), .Y (n_3001));
INVX1 g64552(.A (n_7103), .Y (n_3838));
NAND2X1 g64583(.A (n_6577), .B (n_9448), .Y (n_3797));
CLKBUFX1 g64590(.A (n_2996), .Y (n_3239));
INVX1 g64616(.A (n_3612), .Y (n_5459));
INVX1 g64623(.A (n_3784), .Y (n_3626));
NAND3X1 g64630(.A (n_969), .B (n_2053), .C (n_9425), .Y (n_2989));
NAND4X1 g64632(.A (g5957), .B (n_11101), .C (g17715), .D (n_2421), .Y(n_2988));
INVX1 g64635(.A (n_2987), .Y (n_4053));
AND2X1 g64643(.A (n_2409), .B (g34034), .Y (n_3236));
NAND4X1 g64647(.A (g6649), .B (n_2600), .C (g17764), .D (n_11173), .Y(n_2986));
OR2X1 g64649(.A (n_10697), .B (g5052), .Y (n_2985));
NAND4X1 g64684(.A (n_3181), .B (n_10063), .C (n_2980), .D (n_974), .Y(n_2981));
NAND3X1 g61805(.A (n_830), .B (n_2002), .C (n_9425), .Y (n_2979));
NAND4X1 g64701(.A (g5256), .B (g25219), .C (g17639), .D (g25114), .Y(n_2977));
NAND4X1 g64709(.A (n_1163), .B (n_1668), .C (n_1712), .D (n_938), .Y(n_2975));
AOI22X1 g64710(.A0 (n_1813), .A1 (n_10078), .B0 (n_2973), .B1(g5152), .Y (n_2974));
NAND3X1 g61814(.A (n_848), .B (n_1994), .C (n_9209), .Y (n_2972));
NAND4X1 g64721(.A (n_2352), .B (g6295), .C (g17743), .D (n_11157), .Y(n_2971));
NAND4X1 g64723(.A (n_1226), .B (n_1715), .C (n_1672), .D (n_906), .Y(n_2969));
NAND4X1 g64735(.A (n_6806), .B (g3961), .C (g16659), .D (n_6786), .Y(n_2968));
NAND4X1 g64743(.A (n_1162), .B (n_1704), .C (n_1678), .D (n_915), .Y(n_2967));
NAND4X1 g64749(.A (n_2443), .B (g5603), .C (g17678), .D (n_1023), .Y(n_2966));
NAND4X1 g64759(.A (n_10623), .B (g5949), .C (g17715), .D (n_2376), .Y(n_2965));
NAND4X1 g64771(.A (n_2432), .B (g6641), .C (g17764), .D (n_11184), .Y(n_2964));
MX2X1 g64773(.A (g4939), .B (g4933), .S0 (n_2048), .Y (n_2963));
MX2X1 g64774(.A (g4749), .B (g4743), .S0 (n_2051), .Y (n_2962));
MX2X1 g64782(.A (g4698), .B (g4704), .S0 (n_2068), .Y (n_2961));
MX2X1 g64783(.A (g4754), .B (g4760), .S0 (n_2049), .Y (n_2960));
MX2X1 g64784(.A (g4765), .B (g4771), .S0 (n_2069), .Y (n_2959));
MX2X1 g64785(.A (g4944), .B (g4950), .S0 (n_2065), .Y (n_2958));
MX2X1 g64786(.A (g4955), .B (g4961), .S0 (n_2046), .Y (n_2957));
MX2X1 g64790(.A (g4492), .B (n_1563), .S0 (n_9240), .Y (n_2956));
MX2X1 g64791(.A (g4473), .B (n_1354), .S0 (n_9091), .Y (n_2955));
MX2X1 g64792(.A (g5084), .B (n_696), .S0 (n_9091), .Y (n_2954));
MX2X1 g64793(.A (g_18330), .B (n_469), .S0 (n_9834), .Y (n_2953));
MX2X1 g64794(.A (n_10524), .B (n_10535), .S0 (n_9256), .Y (n_2951));
MX2X1 g64795(.A (g4258), .B (n_695), .S0 (n_9172), .Y (n_2949));
MX2X1 g64796(.A (g_22552), .B (n_1095), .S0 (n_9940), .Y (n_2948));
MX2X1 g64797(.A (g1430), .B (n_652), .S0 (n_9894), .Y (n_2947));
NAND4X1 g62835(.A (n_2945), .B (n_9834), .C (n_2710), .D (n_1330), .Y(n_2946));
NAND2X1 g64850(.A (n_2061), .B (n_9398), .Y (n_3506));
NAND3X1 g64859(.A (n_2943), .B (n_4329), .C (n_10013), .Y (n_2944));
NAND2X1 g64860(.A (n_2785), .B (n_2784), .Y (n_2942));
NAND3X1 g64862(.A (n_2940), .B (n_4327), .C (n_9398), .Y (n_2941));
INVX1 g64864(.A (n_3224), .Y (n_3425));
NAND4X1 g62848(.A (n_2938), .B (n_9651), .C (n_2696), .D (n_1327), .Y(n_2939));
NAND3X1 g64867(.A (n_2936), .B (n_4324), .C (n_9466), .Y (n_2937));
NAND2X1 g64868(.A (n_2363), .B (n_2639), .Y (n_2934));
NAND3X1 g64869(.A (n_3253), .B (n_4316), .C (n_10950), .Y (n_2933));
NAND3X1 g64871(.A (n_2930), .B (n_4322), .C (n_9398), .Y (n_2931));
NAND3X1 g64876(.A (n_2928), .B (n_4320), .C (n_10013), .Y (n_2929));
OAI21X1 g62852(.A0 (n_2312), .A1 (g4854), .B0 (n_2925), .Y (n_2926));
NAND3X1 g64885(.A (n_2923), .B (n_4314), .C (n_9139), .Y (n_2924));
INVX2 g64950(.A (n_3003), .Y (n_3569));
NAND3X1 g64958(.A (n_2608), .B (g1448), .C (n_9698), .Y (n_2920));
INVX1 g61117(.A (n_10431), .Y (n_3910));
AOI21X1 g64993(.A0 (g16718), .A1 (n_238), .B0 (n_2348), .Y (n_2918));
AOI21X1 g64997(.A0 (g16744), .A1 (n_242), .B0 (n_2347), .Y (n_2917));
NAND4X1 g65031(.A (g16775), .B (g16659), .C (g11418), .D (g13966), .Y(n_3486));
MX2X1 g65081(.A (g2886), .B (n_992), .S0 (n_9311), .Y (n_2915));
MX2X1 g65086(.A (g5164), .B (n_1650), .S0 (n_9359), .Y (n_2914));
MX2X1 g65087(.A (g5511), .B (n_1649), .S0 (n_9750), .Y (n_2913));
MX2X1 g65088(.A (g6203), .B (n_1017), .S0 (n_9091), .Y (n_2912));
MX2X1 g65090(.A (g6549), .B (n_1396), .S0 (n_9091), .Y (n_2911));
MX2X1 g65091(.A (g3506), .B (n_1115), .S0 (n_9448), .Y (n_2910));
MX2X1 g65092(.A (g3155), .B (n_1109), .S0 (n_9091), .Y (n_2909));
MX2X1 g65094(.A (g3857), .B (n_1113), .S0 (n_9091), .Y (n_2907));
MX2X1 g65096(.A (g5857), .B (n_1002), .S0 (n_9091), .Y (n_2906));
MX2X1 g65097(.A (g5057), .B (n_2045), .S0 (n_9359), .Y (n_2905));
MX2X1 g65098(.A (n_1177), .B (n_1077), .S0 (n_9256), .Y (n_2904));
MX2X1 g65099(.A (n_1234), .B (n_1079), .S0 (n_9000), .Y (n_2903));
MX2X1 g65100(.A (g4308), .B (n_1570), .S0 (n_9834), .Y (n_2902));
MX2X1 g65101(.A (n_1169), .B (n_1069), .S0 (n_9091), .Y (n_2900));
MX2X1 g65102(.A (n_1214), .B (n_1072), .S0 (n_9000), .Y (n_2898));
MX2X1 g65103(.A (n_1135), .B (n_1075), .S0 (n_9750), .Y (n_2897));
MX2X1 g65104(.A (g_16571), .B (n_1081), .S0 (n_9240), .Y (n_2896));
MX2X1 g65105(.A (g4291), .B (n_1556), .S0 (n_9358), .Y (n_2895));
MX2X1 g65106(.A (n_1210), .B (n_1074), .S0 (n_8955), .Y (n_2894));
MX2X1 g65108(.A (n_1191), .B (n_998), .S0 (n_9167), .Y (n_2892));
MX2X1 g65109(.A (g_17426), .B (g_10278), .S0 (n_3177), .Y (n_2891));
MX2X1 g65110(.A (g4281), .B (n_1820), .S0 (n_9091), .Y (n_2890));
MX2X1 g65111(.A (g1306), .B (n_1997), .S0 (n_9000), .Y (n_2889));
MX2X1 g65112(.A (n_1216), .B (n_1071), .S0 (n_9750), .Y (n_2888));
MX2X1 g65113(.A (g1183), .B (n_1991), .S0 (n_9359), .Y (n_2887));
MX2X1 g65114(.A (g_15758), .B (n_1992), .S0 (n_8955), .Y (n_2886));
NAND3X1 g65260(.A (g_19911), .B (n_3323), .C (n_9501), .Y (n_2885));
INVX1 g65264(.A (n_2883), .Y (n_2884));
NOR2X1 g65276(.A (n_2881), .B (n_2838), .Y (n_2882));
NOR2X1 g65278(.A (n_6398), .B (n_2319), .Y (n_2880));
NAND3X1 g61929(.A (g_18902), .B (n_2878), .C (n_9750), .Y (n_2879));
NAND3X1 g65348(.A (g1345), .B (n_3459), .C (n_10063), .Y (n_2875));
NOR2X1 g65371(.A (n_2871), .B (n_2835), .Y (n_2872));
NAND3X1 g61943(.A (n_2003), .B (g_18869), .C (n_9091), .Y (n_2870));
NOR2X1 g65419(.A (g16775), .B (n_2594), .Y (n_2869));
OR4X1 g61951(.A (n_2867), .B (n_2410), .C (n_9129), .D (g4669), .Y(n_2868));
NAND3X1 g65422(.A (n_987), .B (n_986), .C (n_10005), .Y (n_2866));
OAI22X1 g65500(.A0 (n_2578), .A1 (n_1468), .B0 (n_612), .B1(n_10063), .Y (n_2864));
OAI22X1 g65503(.A0 (n_2862), .A1 (g4473), .B0 (n_2861), .B1 (n_9830),.Y (n_2863));
NOR2X1 g65698(.A (n_2859), .B (g5164), .Y (n_2860));
NOR2X1 g65704(.A (n_2857), .B (g5857), .Y (n_2858));
NOR2X1 g65711(.A (n_2855), .B (g5511), .Y (n_2856));
NOR2X1 g65737(.A (n_2853), .B (g3155), .Y (n_2854));
NAND3X1 g65769(.A (g_16404), .B (g_16571), .C (n_9651), .Y (n_2852));
NOR2X1 g65773(.A (n_2849), .B (g3506), .Y (n_2850));
NOR2X1 g65811(.A (n_2847), .B (g3857), .Y (n_2848));
MX2X1 g61435(.A (n_8508), .B (n_1351), .S0 (n_9000), .Y (n_2846));
NOR2X1 g62013(.A (n_2174), .B (g4939), .Y (n_2845));
NOR2X1 g62014(.A (n_2173), .B (g4950), .Y (n_2844));
NOR2X1 g65874(.A (n_2842), .B (g6549), .Y (n_2843));
NAND2X1 g61162(.A (n_10242), .B (n_2176), .Y (n_2841));
OAI21X1 g65951(.A0 (g_18015), .A1 (n_2518), .B0 (n_9351), .Y(n_2840));
OAI21X1 g66005(.A0 (n_144), .A1 (n_9311), .B0 (n_2838), .Y (n_2839));
OAI21X1 g66007(.A0 (n_1), .A1 (n_9422), .B0 (n_2835), .Y (n_2837));
NAND2X1 g61164(.A (n_2180), .B (n_10243), .Y (n_2834));
OAI21X1 g66019(.A0 (n_127), .A1 (n_9422), .B0 (n_2606), .Y (n_2833));
MX2X1 g66124(.A (g4146), .B (g4157), .S0 (n_9240), .Y (n_2832));
OAI21X1 g66029(.A0 (n_39), .A1 (n_9425), .B0 (n_2661), .Y (n_2831));
AOI21X1 g61166(.A0 (n_2), .A1 (n_1275), .B0 (n_2830), .Y (n_3123));
OAI21X1 g66040(.A0 (n_117), .A1 (n_9425), .B0 (n_2828), .Y (n_2829));
OAI22X1 g66096(.A0 (n_10280), .A1 (n_9627), .B0 (n_169), .B1(n_9672), .Y (n_2827));
MX2X1 g66097(.A (g2844), .B (g2852), .S0 (n_9000), .Y (n_2826));
MX2X1 g66101(.A (g2936), .B (g2950), .S0 (n_10005), .Y (n_2824));
MX2X1 g66102(.A (g4722), .B (g4737), .S0 (n_8955), .Y (n_2823));
MX2X1 g66103(.A (g2852), .B (g2860), .S0 (n_9091), .Y (n_2822));
MX2X1 g66106(.A (g2890), .B (g2844), .S0 (n_9000), .Y (n_2821));
MX2X1 g66113(.A (g2860), .B (g2894), .S0 (n_9000), .Y (n_2820));
MX2X1 g66114(.A (g2894), .B (n_22), .S0 (n_9172), .Y (n_2819));
MX2X1 g66118(.A (g2950), .B (g2960), .S0 (n_9311), .Y (n_2817));
MX2X1 g66119(.A (g2868), .B (g2873), .S0 (n_9234), .Y (n_2816));
MX2X1 g66120(.A (g2130), .B (g2138), .S0 (n_9091), .Y (n_2815));
OAI22X1 g66121(.A0 (n_1240), .A1 (n_10385), .B0 (n_308), .B1(n_9903), .Y (n_2814));
MX2X1 g66126(.A (g4249), .B (g4245), .S0 (n_9333), .Y (n_2813));
MX2X1 g66128(.A (g4300), .B (g4253), .S0 (n_9311), .Y (n_2812));
MX2X1 g66129(.A (n_22), .B (g20652), .S0 (n_9834), .Y (n_2810));
OR4X1 g62078(.A (n_2925), .B (n_2361), .C (n_9404), .D (n_11216), .Y(n_2809));
MX2X1 g66133(.A (g2960), .B (g2970), .S0 (n_9167), .Y (n_2808));
MX2X1 g66137(.A (n_11097), .B (g2697), .S0 (n_9091), .Y (n_2807));
MX2X1 g66138(.A (g4727), .B (g4732), .S0 (n_9172), .Y (n_2806));
MX2X1 g66143(.A (g2984), .B (g2907), .S0 (n_9311), .Y (n_2805));
MX2X1 g66145(.A (g4907), .B (g4912), .S0 (n_9834), .Y (n_2804));
MX2X1 g66147(.A (g4917), .B (g4922), .S0 (n_9234), .Y (n_2803));
MX2X1 g66148(.A (g4912), .B (g4927), .S0 (n_9256), .Y (n_2802));
MX2X1 g61486(.A (g4430), .B (n_1315), .S0 (n_8955), .Y (n_2801));
NAND2X1 g66280(.A (n_10112), .B (n_9431), .Y (n_2800));
NAND2X1 g66322(.A (n_10188), .B (n_9371), .Y (n_2798));
NAND2X1 g66323(.A (n_3914), .B (n_9431), .Y (n_2797));
AND2X1 g66398(.A (n_8895), .B (n_9019), .Y (n_2796));
NAND2X1 g66401(.A (n_926), .B (n_9884), .Y (n_2795));
NAND2X1 g66411(.A (n_2861), .B (n_9940), .Y (n_3071));
NAND2X1 g66412(.A (g1367), .B (n_9772), .Y (n_2794));
AND2X1 g66419(.A (g4153), .B (n_9672), .Y (n_2793));
NAND2X1 g61498(.A (n_2790), .B (n_1986), .Y (n_2791));
AND2X1 g66439(.A (g2975), .B (n_9672), .Y (n_2789));
AND2X1 g66443(.A (g4104), .B (n_9672), .Y (n_2788));
AND2X1 g66464(.A (g4087), .B (n_9672), .Y (n_2787));
OR2X1 g64887(.A (n_2785), .B (n_2784), .Y (g28041));
NAND2X1 g66525(.A (g_22306), .B (n_9419), .Y (n_2783));
NOR2X1 g66541(.A (g4258), .B (n_9772), .Y (n_2782));
NAND2X1 g66543(.A (n_2780), .B (n_9836), .Y (n_2781));
NAND2X1 g66549(.A (g1345), .B (n_9505), .Y (n_2779));
NAND2X1 g66557(.A (n_662), .B (n_9952), .Y (n_2778));
AND2X1 g66611(.A (g5188), .B (n_9448), .Y (n_2777));
NOR2X1 g66698(.A (n_553), .B (n_9353), .Y (n_2776));
NAND2X1 g66715(.A (g2882), .B (n_9952), .Y (n_2775));
NAND2X1 g63451(.A (n_2483), .B (n_10818), .Y (n_3651));
MX2X1 g61182(.A (n_2773), .B (n_1869), .S0 (n_8955), .Y (n_2774));
AND2X1 g66753(.A (g6573), .B (n_9698), .Y (n_2772));
AND2X1 g66807(.A (g3881), .B (n_9448), .Y (n_2770));
AND2X1 g66823(.A (g3530), .B (n_9448), .Y (n_2769));
NOR2X1 g66852(.A (n_10557), .B (n_9775), .Y (n_2768));
NAND2X1 g66853(.A (n_955), .B (n_9952), .Y (n_2767));
AND2X1 g66879(.A (g5881), .B (n_9448), .Y (n_2766));
NOR2X1 g66909(.A (n_617), .B (n_9019), .Y (n_2765));
NAND4X1 g63529(.A (n_1597), .B (n_10112), .C (n_9883), .D (n_392), .Y(n_2764));
NAND2X1 g61568(.A (n_9811), .B (g12919), .Y (n_3316));
MX2X1 g66100(.A (g2994), .B (g2988), .S0 (n_9000), .Y (n_2762));
MX2X1 g63787(.A (g5092), .B (n_1590), .S0 (n_10005), .Y (n_2761));
MX2X1 g63788(.A (n_10128), .B (n_1842), .S0 (n_9797), .Y (n_2760));
MX2X1 g63798(.A (g4264), .B (n_1839), .S0 (n_9000), .Y (n_2759));
MX2X1 g63806(.A (g1548), .B (n_1296), .S0 (n_9358), .Y (n_2758));
NAND2X1 g63899(.A (n_2465), .B (n_684), .Y (n_3563));
OR2X1 g63903(.A (n_3844), .B (g_6283), .Y (n_2757));
NAND4X1 g64057(.A (n_2129), .B (n_1669), .C (n_1717), .D (n_1694), .Y(n_2756));
NAND4X1 g64058(.A (n_1846), .B (n_1857), .C (n_1844), .D (n_1699), .Y(n_2755));
INVX1 g64092(.A (n_2754), .Y (n_3332));
MX2X1 g64096(.A (n_276), .B (n_2090), .S0 (n_8955), .Y (n_2753));
OR2X1 g64139(.A (n_3174), .B (n_83), .Y (n_2751));
OAI21X1 g64143(.A0 (n_2945), .A1 (n_10753), .B0 (n_10005), .Y(n_2749));
AOI21X1 g64150(.A0 (n_2110), .A1 (n_344), .B0 (n_643), .Y (n_2748));
NAND3X1 g64165(.A (n_2457), .B (n_2456), .C (n_2747), .Y (n_3502));
OR4X1 g64247(.A (n_2980), .B (n_276), .C (n_9129), .D (g4633), .Y(n_2746));
NAND2X1 g64259(.A (n_3174), .B (g_21576), .Y (n_2744));
INVX1 g64282(.A (n_2743), .Y (n_3493));
NAND2X1 g61730(.A (n_2430), .B (n_10005), .Y (n_2742));
NOR2X1 g64323(.A (n_1632), .B (n_2154), .Y (n_2741));
NAND3X1 g64327(.A (n_1658), .B (n_1887), .C (n_9209), .Y (n_2740));
MX2X1 g61295(.A (g1404), .B (n_1569), .S0 (n_9091), .Y (n_2739));
NAND4X1 g64362(.A (n_1193), .B (n_1689), .C (n_1707), .D (n_932), .Y(n_2738));
OAI21X1 g64388(.A0 (n_3171), .A1 (n_1695), .B0 (n_2302), .Y (n_2736));
OAI21X1 g64389(.A0 (n_2881), .A1 (n_2734), .B0 (n_2241), .Y (n_2735));
OAI21X1 g64390(.A0 (n_2732), .A1 (n_2421), .B0 (n_2289), .Y (n_2733));
OAI21X1 g64391(.A0 (n_2729), .A1 (n_11150), .B0 (n_2277), .Y(n_2730));
OAI21X1 g64392(.A0 (n_2871), .A1 (n_11173), .B0 (n_2274), .Y(n_2727));
MX2X1 g61750(.A (n_2429), .B (n_2032), .S0 (n_9797), .Y (n_2725));
MX2X1 g64425(.A (g5156), .B (n_1792), .S0 (n_9333), .Y (n_2722));
MX2X1 g64426(.A (g5124), .B (n_2087), .S0 (n_9240), .Y (n_2720));
MX2X1 g64427(.A (n_2718), .B (n_1814), .S0 (n_9797), .Y (n_2719));
MX2X1 g64428(.A (n_2943), .B (n_1798), .S0 (n_9000), .Y (n_2716));
MX2X1 g64429(.A (g5471), .B (n_2098), .S0 (n_9091), .Y (n_2715));
MX2X1 g64432(.A (n_2940), .B (n_1809), .S0 (n_9992), .Y (n_2714));
MX2X1 g64433(.A (g5817), .B (n_2097), .S0 (n_9091), .Y (n_2713));
MX2X1 g64435(.A (n_2936), .B (n_2086), .S0 (n_9091), .Y (n_2712));
NAND4X1 g62668(.A (n_2710), .B (n_2945), .C (n_9664), .D (n_8799), .Y(n_2711));
MX2X1 g64438(.A (g3115), .B (n_2092), .S0 (n_9311), .Y (n_2709));
MX2X1 g64439(.A (n_2930), .B (n_1803), .S0 (n_9156), .Y (n_2707));
MX2X1 g64440(.A (g6509), .B (n_2095), .S0 (n_9091), .Y (n_2706));
MX2X1 g64443(.A (n_2704), .B (n_2085), .S0 (n_9000), .Y (n_2705));
MX2X1 g64444(.A (n_2928), .B (n_1801), .S0 (n_9167), .Y (n_2703));
MX2X1 g64445(.A (g3466), .B (n_2091), .S0 (n_9627), .Y (n_2702));
MX2X1 g64446(.A (n_2699), .B (n_1800), .S0 (n_9000), .Y (n_2700));
NAND4X1 g62674(.A (n_2696), .B (n_2938), .C (n_9992), .D (g1554), .Y(n_2697));
MX2X1 g64448(.A (n_2923), .B (n_1843), .S0 (n_9156), .Y (n_2695));
MX2X1 g64449(.A (g3817), .B (n_2093), .S0 (n_9664), .Y (n_2694));
MX2X1 g64450(.A (n_2692), .B (n_1797), .S0 (n_9000), .Y (n_2693));
MX2X1 g64451(.A (g_14535), .B (n_2083), .S0 (n_9218), .Y (n_2691));
MX2X1 g64452(.A (n_2005), .B (n_1793), .S0 (n_9797), .Y (n_2690));
MX2X1 g64454(.A (g4245), .B (n_1821), .S0 (n_9240), .Y (n_2689));
MX2X1 g64455(.A (g1489), .B (n_1804), .S0 (n_9359), .Y (n_2688));
MX2X1 g64456(.A (n_2686), .B (n_1806), .S0 (n_9256), .Y (n_2687));
MX2X1 g64458(.A (n_2684), .B (n_1808), .S0 (n_8955), .Y (n_2685));
AND2X1 g64507(.A (n_10526), .B (g_12791), .Y (n_3291));
NOR2X1 g64510(.A (n_1571), .B (n_9353), .Y (n_2682));
NAND2X1 g64517(.A (n_3152), .B (n_9209), .Y (n_3489));
AOI21X1 g64526(.A0 (n_2679), .A1 (n_3984), .B0 (n_10134), .Y(n_2680));
OR2X1 g64530(.A (n_2426), .B (n_2677), .Y (n_2678));
NAND2X1 g64547(.A (n_6695), .B (n_9627), .Y (n_2675));
NOR2X1 g64548(.A (n_1268), .B (n_2406), .Y (n_2673));
XOR2X1 g61328(.A (g1404), .B (n_2671), .Y (n_2672));
NOR2X1 g64557(.A (n_3062), .B (n_2668), .Y (n_2669));
INVX2 g64563(.A (n_11207), .Y (n_6243));
NAND3X1 g64584(.A (n_981), .B (n_1756), .C (n_9091), .Y (n_2666));
NAND3X1 g64585(.A (n_849), .B (n_2056), .C (n_9558), .Y (n_2665));
AND2X1 g64591(.A (n_2387), .B (g34036), .Y (n_2996));
NAND2X1 g64603(.A (n_3152), .B (n_988), .Y (n_2664));
NOR2X1 g64606(.A (n_2630), .B (n_1549), .Y (n_2663));
NOR2X1 g64626(.A (n_3065), .B (n_2661), .Y (n_2662));
NAND4X1 g64627(.A (g5611), .B (n_2597), .C (g17678), .D (n_2208), .Y(n_2660));
NAND4X1 g64629(.A (g6303), .B (n_2325), .C (g17743), .D (n_11150), .Y(n_2659));
NAND2X1 g64631(.A (n_2118), .B (n_2657), .Y (n_2658));
INVX1 g64636(.A (n_6765), .Y (n_2987));
NAND4X1 g64662(.A (n_777), .B (n_1541), .C (n_1548), .D (n_2452), .Y(n_2656));
NOR2X1 g64663(.A (n_1976), .B (n_2654), .Y (n_2655));
NAND4X1 g64716(.A (n_8586), .B (g3259), .C (g16603), .D (n_8548), .Y(n_2653));
NAND4X1 g64736(.A (n_10879), .B (g3610), .C (g16627), .D (n_4682), .Y(n_2652));
NAND4X1 g64737(.A (n_920), .B (n_1530), .C (n_1521), .D (n_704), .Y(n_2651));
XOR2X1 g64788(.A (g8358), .B (n_1733), .Y (n_2648));
INVX1 g64817(.A (g5339), .Y (n_2647));
INVX1 g64819(.A (g6377), .Y (n_2646));
INVX1 g64828(.A (g5685), .Y (n_2645));
INVX1 g64830(.A (g6723), .Y (n_2644));
INVX1 g64833(.A (g6031), .Y (n_2642));
NAND2X1 g64841(.A (n_2640), .B (g_8896), .Y (n_2641));
NOR2X1 g64865(.A (n_2640), .B (n_2639), .Y (n_3224));
OR2X1 g64873(.A (n_2042), .B (g5041), .Y (n_2638));
NAND2X2 g64906(.A (n_11192), .B (n_11193), .Y (n_3259));
NAND2X1 g64907(.A (n_2034), .B (n_1682), .Y (n_2637));
NAND3X1 g64937(.A (n_2057), .B (g1478), .C (n_9811), .Y (n_2634));
NAND3X1 g64938(.A (n_2054), .B (g1300), .C (n_9558), .Y (n_2632));
BUFX3 g64951(.A (n_10526), .Y (n_3003));
NOR2X1 g64965(.A (n_1975), .B (n_8694), .Y (n_2629));
AOI21X1 g64967(.A0 (n_1363), .A1 (n_10813), .B0 (n_3177), .Y(n_2628));
AND2X1 g64970(.A (n_2070), .B (n_6970), .Y (n_3016));
XOR2X1 g64982(.A (n_2871), .B (n_11171), .Y (n_2625));
XOR2X1 g64985(.A (n_2881), .B (n_2224), .Y (n_2624));
NAND2X1 g61371(.A (g4427), .B (n_9129), .Y (n_2619));
CLKBUFX1 gbuf_d_1075(.A(g16603), .Y(d_out_1075));
CLKBUFX1 gbuf_q_1075(.A(q_in_1075), .Y(g16624));
CLKBUFX1 gbuf_d_1076(.A(g16627), .Y(d_out_1076));
CLKBUFX1 gbuf_q_1076(.A(q_in_1076), .Y(g16656));
NAND2X1 g65236(.A (g26801), .B (n_9750), .Y (n_2616));
OR2X1 g65241(.A (n_4316), .B (n_9772), .Y (n_2615));
NOR2X1 g65248(.A (n_1576), .B (n_9193), .Y (n_4091));
OAI21X1 g65254(.A0 (n_276), .A1 (n_10402), .B0 (n_9894), .Y (n_2614));
NOR2X1 g65265(.A (n_3177), .B (n_3391), .Y (n_2883));
NOR2X1 g65280(.A (n_2732), .B (n_2612), .Y (n_2613));
NAND2X1 g65292(.A (n_6404), .B (n_6395), .Y (n_6400));
NAND2X1 g65324(.A (n_3184), .B (n_10524), .Y (n_2611));
NOR2X1 g65328(.A (n_4617), .B (n_10078), .Y (n_2610));
INVX1 g65346(.A (n_2608), .Y (n_2609));
NOR2X1 g65351(.A (n_2729), .B (n_2606), .Y (n_2607));
NAND2X1 g66420(.A (g4664), .B (n_9884), .Y (n_2604));
NAND3X1 g61949(.A (n_1993), .B (g_11413), .C (n_9311), .Y (n_2603));
OR2X1 g65430(.A (n_2004), .B (n_10184), .Y (n_2602));
NAND4X1 g65473(.A (g6585), .B (n_2600), .C (g12470), .D (n_11171), .Y(n_2601));
NAND4X1 g65477(.A (g5547), .B (n_2597), .C (g12300), .D (n_1023), .Y(n_2598));
OAI21X1 g65502(.A0 (g1442), .A1 (n_9599), .B0 (n_2006), .Y (n_2595));
NAND2X1 g61149(.A (n_2592), .B (g1542), .Y (n_4241));
OR2X1 g61150(.A (n_2592), .B (g1542), .Y (n_2593));
NAND3X1 g65687(.A (n_1356), .B (n_9811), .C (n_107), .Y (n_2590));
OR2X1 g65690(.A (g5112), .B (n_9398), .Y (n_2589));
NOR2X1 g65700(.A (n_1058), .B (n_9107), .Y (n_2588));
OAI21X1 g64021(.A0 (n_1826), .A1 (g4849), .B0 (n_1875), .Y (n_2587));
AND2X1 g61154(.A (n_6781), .B (n_11042), .Y (n_3183));
NOR2X1 g65803(.A (n_1982), .B (n_16), .Y (n_2586));
NOR2X1 g65823(.A (n_1979), .B (n_40), .Y (n_2585));
NAND2X1 g65876(.A (n_2583), .B (n_3857), .Y (n_2584));
NOR2X1 g65887(.A (n_1971), .B (g4616), .Y (n_2582));
INVX1 g65895(.A (n_2580), .Y (n_2581));
NOR2X1 g65908(.A (n_2578), .B (g6203), .Y (n_2579));
NAND2X1 g65953(.A (n_2481), .B (n_2480), .Y (n_2575));
NAND2X1 g61463(.A (n_9359), .B (g12923), .Y (n_3165));
NOR2X1 g62058(.A (n_1969), .B (n_4764), .Y (n_2574));
NOR2X1 g62064(.A (n_2000), .B (n_4761), .Y (n_2573));
NOR2X1 g62065(.A (n_1977), .B (n_4757), .Y (n_2572));
NAND2X1 g66302(.A (n_2566), .B (n_9466), .Y (n_2567));
NAND2X1 g66306(.A (g4608), .B (n_9431), .Y (n_2564));
INVX1 g66309(.A (n_2562), .Y (n_2563));
NAND2X1 g66318(.A (g5813), .B (n_9775), .Y (n_2560));
OR2X1 g66330(.A (n_9672), .B (g10122), .Y (n_2559));
NAND2X1 g66334(.A (g2227), .B (n_9672), .Y (n_2558));
NAND2X1 g66365(.A (n_2556), .B (n_9107), .Y (n_2557));
NAND2X1 g66374(.A (g1384), .B (n_9505), .Y (n_2555));
NOR2X1 g66393(.A (n_10314), .B (n_10716), .Y (n_2554));
NAND2X1 g66397(.A (n_2550), .B (n_9836), .Y (n_2551));
NAND2X1 g66405(.A (g_12465), .B (n_9976), .Y (n_2548));
NOR2X1 g66406(.A (g_18112), .B (n_10376), .Y (n_2546));
NAND2X1 g66413(.A (g4628), .B (n_9599), .Y (n_2545));
NAND2X1 g66438(.A (g_14342), .B (n_9928), .Y (n_2543));
NAND2X1 g66463(.A (g6159), .B (n_9599), .Y (n_2540));
NAND2X1 g66472(.A (n_2538), .B (n_10952), .Y (n_2539));
NAND2X1 g66482(.A (g2236), .B (n_9300), .Y (n_2537));
NAND2X1 g66495(.A (n_2535), .B (n_9193), .Y (n_2536));
NAND2X1 g66501(.A (n_4339), .B (n_9952), .Y (n_2533));
NAND2X1 g66509(.A (g_19304), .B (n_9300), .Y (n_2531));
NAND2X1 g66510(.A (n_2529), .B (n_9628), .Y (n_2530));
NAND2X1 g66522(.A (g_16958), .B (n_10078), .Y (n_2528));
NAND2X1 g66533(.A (g_20159), .B (n_9836), .Y (n_2526));
NAND2X1 g66540(.A (g2638), .B (n_9300), .Y (n_2524));
NAND2X1 g66555(.A (g1677), .B (n_9505), .Y (n_2523));
NAND2X1 g66561(.A (n_2521), .B (n_10952), .Y (n_2522));
NAND2X1 g66565(.A (n_8913), .B (n_9884), .Y (n_2520));
NOR2X1 g66602(.A (n_9836), .B (n_2518), .Y (n_2519));
AND2X1 g66636(.A (g5535), .B (n_9698), .Y (n_2517));
NAND2X1 g66643(.A (n_9553), .B (g6748), .Y (n_3117));
NAND2X1 g66672(.A (g25219), .B (n_9139), .Y (n_3121));
AND2X1 g66676(.A (n_11097), .B (n_9717), .Y (n_2515));
OR2X1 g66684(.A (g4108), .B (n_9627), .Y (n_2514));
AND2X1 g66695(.A (g4917), .B (n_9501), .Y (n_2512));
OR2X1 g66697(.A (g2756), .B (n_9453), .Y (n_2510));
OR2X1 g66701(.A (n_3463), .B (n_9627), .Y (n_2509));
NAND2X1 g66707(.A (n_9553), .B (g6750), .Y (n_3113));
AND2X1 g66714(.A (n_9501), .B (g6745), .Y (n_2507));
NOR2X1 g66727(.A (n_365), .B (n_9884), .Y (n_2506));
AND2X1 g66744(.A (g2130), .B (n_9717), .Y (n_2504));
OR2X1 g66745(.A (g4141), .B (n_9501), .Y (n_2503));
OR2X1 g66750(.A (g4082), .B (n_9627), .Y (n_2502));
AND2X1 g66751(.A (n_9501), .B (g21176), .Y (n_2501));
NOR2X1 g66763(.A (n_383), .B (n_9107), .Y (n_2500));
OR2X1 g66810(.A (g2955), .B (n_9398), .Y (n_2499));
NAND2X1 g66840(.A (n_9627), .B (g6749), .Y (n_3115));
OR2X1 g66844(.A (g4098), .B (n_9627), .Y (n_2498));
INVX1 g66858(.A (n_2496), .Y (n_2497));
NOR2X1 g66893(.A (g_18200), .B (n_9107), .Y (n_2495));
NOR2X1 g66894(.A (n_261), .B (n_10078), .Y (n_2494));
OR2X1 g66897(.A (g2873), .B (n_9501), .Y (n_2493));
AND2X1 g66903(.A (g4727), .B (n_10005), .Y (n_2492));
OR2X1 g66905(.A (n_10650), .B (n_9501), .Y (n_2491));
NAND2X1 g61530(.A (g23683), .B (n_9772), .Y (n_2488));
NAND2X1 g66544(.A (n_2485), .B (n_9628), .Y (n_2486));
XOR2X1 g64079(.A (n_221), .B (n_2165), .Y (n_2484));
INVX1 g64093(.A (n_2483), .Y (n_2754));
OR2X1 g65969(.A (n_2481), .B (n_2480), .Y (g28042));
NAND2X1 g64151(.A (n_1863), .B (n_10949), .Y (n_3148));
NAND4X1 g64185(.A (n_1567), .B (n_1822), .C (n_11051), .D (n_273), .Y(n_2479));
NAND2X1 g64237(.A (n_1862), .B (n_10687), .Y (n_3036));
NAND2X1 g64253(.A (n_1861), .B (n_10949), .Y (n_3035));
NAND2X1 g64261(.A (n_2152), .B (n_9862), .Y (n_3149));
AOI21X1 g64283(.A0 (n_1429), .A1 (n_1832), .B0 (n_1838), .Y (n_2743));
OAI21X1 g61288(.A0 (n_2062), .A1 (n_2474), .B0 (n_2063), .Y (n_2475));
NAND4X1 g64363(.A (n_925), .B (n_1516), .C (n_1525), .D (n_927), .Y(n_2472));
AOI22X1 g64364(.A0 (n_1791), .A1 (n_448), .B0 (n_797), .B1 (g4311),.Y (n_2471));
NAND4X1 g64366(.A (n_929), .B (n_1511), .C (n_1534), .D (n_894), .Y(n_2469));
AOI21X1 g64393(.A0 (n_10664), .A1 (n_1538), .B0 (n_2151), .Y(n_2468));
NAND4X1 g64405(.A (n_934), .B (n_1507), .C (n_1523), .D (n_895), .Y(n_2466));
INVX1 g64413(.A (n_2465), .Y (n_2723));
NOR2X1 g64511(.A (n_10496), .B (n_10525), .Y (n_3431));
OR2X1 g64513(.A (n_2096), .B (n_10952), .Y (n_2464));
OR2X1 g64514(.A (n_2094), .B (n_9193), .Y (n_2463));
OR2X1 g64516(.A (n_2089), .B (n_9193), .Y (n_2461));
OR2X1 g64518(.A (n_2088), .B (n_9491), .Y (n_2460));
NAND3X1 g64550(.A (n_2458), .B (n_10725), .C (n_10063), .Y (n_2459));
AND2X1 g64554(.A (n_2457), .B (n_2456), .Y (n_3031));
AND2X1 g64576(.A (n_2103), .B (n_10005), .Y (n_2454));
NAND2X1 g64592(.A (n_2107), .B (g_17934), .Y (n_2453));
OR2X1 g64888(.A (n_1736), .B (n_2449), .Y (g26875));
NAND4X1 g64702(.A (n_2447), .B (g3937), .C (g16775), .D (n_8917), .Y(n_2448));
NAND4X1 g64742(.A (n_1494), .B (n_2443), .C (g17711), .D (g5591), .Y(n_2444));
INVX1 g64745(.A (n_2134), .Y (n_2442));
NAND4X1 g64747(.A (n_1494), .B (n_2439), .C (g17580), .D (g5607), .Y(n_2441));
NAND4X1 g64748(.A (n_7150), .B (g5575), .C (g14694), .D (n_1494), .Y(n_2438));
INVX1 g64766(.A (n_2120), .Y (n_2437));
NAND4X1 g64768(.A (n_2433), .B (n_2435), .C (g17688), .D (g6645), .Y(n_2436));
NAND4X1 g64769(.A (n_2433), .B (n_2432), .C (g17778), .D (g6629), .Y(n_2434));
NAND4X1 g64770(.A (n_2433), .B (g6613), .C (g14828), .D (n_3275), .Y(n_2431));
OAI21X1 g61838(.A0 (n_2345), .A1 (n_2429), .B0 (n_1645), .Y (n_2430));
CLKBUFX1 gbuf_d_1077(.A(g17639), .Y(d_out_1077));
CLKBUFX1 gbuf_q_1077(.A(q_in_1077), .Y(g5339));
CLKBUFX1 gbuf_d_1078(.A(g17743), .Y(d_out_1078));
CLKBUFX1 gbuf_q_1078(.A(q_in_1078), .Y(g6377));
CLKBUFX1 gbuf_d_1079(.A(g17678), .Y(d_out_1079));
CLKBUFX1 gbuf_q_1079(.A(q_in_1079), .Y(g5685));
CLKBUFX1 gbuf_d_1080(.A(g17764), .Y(d_out_1080));
CLKBUFX1 gbuf_q_1080(.A(q_in_1080), .Y(g6723));
CLKBUFX1 gbuf_d_1081(.A(g17715), .Y(d_out_1081));
CLKBUFX1 gbuf_q_1081(.A(q_in_1081), .Y(g6031));
NAND2X1 g64838(.A (n_2427), .B (g1199), .Y (n_3844));
OR2X1 g64839(.A (n_2427), .B (g1199), .Y (n_2428));
NAND2X1 g64842(.A (n_2449), .B (n_38), .Y (n_2426));
OR2X1 g64845(.A (n_891), .B (n_9526), .Y (n_2425));
NAND4X1 g64856(.A (n_2421), .B (g5941), .C (g14673), .D (n_10808), .Y(n_2423));
INVX1 g64857(.A (n_10268), .Y (g27831));
NAND2X1 g66449(.A (g2079), .B (n_9371), .Y (n_2419));
NAND4X1 g64893(.A (n_1785), .B (n_946), .C (g4698), .D (n_10225), .Y(n_2416));
NAND2X1 g64909(.A (n_1680), .B (n_1675), .Y (n_2415));
NAND2X1 g64910(.A (n_1674), .B (n_1681), .Y (n_3013));
NAND4X1 g64917(.A (n_2413), .B (g6287), .C (g14705), .D (n_11150), .Y(n_2414));
INVX1 g64921(.A (n_2410), .Y (n_3152));
NAND4X1 g64927(.A (n_1786), .B (n_11133), .C (g4888), .D (n_740), .Y(n_2409));
NOR2X1 g64928(.A (n_2061), .B (n_598), .Y (n_2465));
NAND4X1 g64929(.A (n_2435), .B (g6633), .C (g14749), .D (n_11173), .Y(n_2408));
OR4X1 g64932(.A (n_1735), .B (g4616), .C (n_9019), .D (g4608), .Y(n_2406));
NAND3X1 g64956(.A (n_2403), .B (n_572), .C (g4057), .Y (n_3728));
NAND3X1 g64957(.A (n_2403), .B (g4064), .C (g4057), .Y (n_3726));
NAND3X1 g64959(.A (n_2403), .B (g4064), .C (n_571), .Y (n_3730));
NAND3X1 g64960(.A (n_1757), .B (g1472), .C (n_9698), .Y (n_2400));
INVX1 g64962(.A (n_2456), .Y (n_2630));
AOI21X1 g64983(.A0 (g_16456), .A1 (n_10557), .B0 (n_10560), .Y(n_2983));
XOR2X1 g64984(.A (n_3171), .B (g25219), .Y (n_2398));
XOR2X1 g64987(.A (n_2732), .B (n_2376), .Y (n_2397));
NAND2X1 g66444(.A (n_365), .B (n_9091), .Y (n_2849));
XOR2X1 g64991(.A (n_11157), .B (n_2729), .Y (n_2392));
AOI21X1 g64996(.A0 (n_10557), .A1 (g_18869), .B0 (n_10560), .Y(n_2670));
NAND4X1 g65022(.A (n_10906), .B (g4765), .C (n_8639), .D (n_8777), .Y(n_2391));
NAND4X1 g65023(.A (g5240), .B (n_10621), .C (g14597), .D (g25219), .Y(n_2389));
NAND4X1 g65026(.A (g6625), .B (n_3275), .C (g14749), .D (n_11184), .Y(n_2388));
NAND4X1 g65027(.A (g16744), .B (g16627), .C (g11388), .D (g13926), .Y(n_3062));
NAND4X1 g65028(.A (g16718), .B (g16603), .C (g_4050), .D (g13895), .Y(n_3065));
NOR2X1 g66441(.A (g4332), .B (n_9884), .Y (n_3213));
NAND4X1 g65033(.A (n_8676), .B (g4944), .C (n_10984), .D (n_10998),.Y (n_2387));
NAND4X1 g65035(.A (n_10905), .B (g4743), .C (n_8639), .D (n_8810), .Y(n_2385));
NAND4X1 g65037(.A (g5587), .B (n_7150), .C (g14635), .D (n_1023), .Y(n_2382));
NAND4X1 g65038(.A (n_8676), .B (g4933), .C (n_10185), .D (n_10984),.Y (n_10181));
NAND4X1 g65039(.A (g6279), .B (n_3277), .C (g14705), .D (n_11157), .Y(n_2379));
NAND4X1 g65040(.A (g5933), .B (n_10506), .C (g14673), .D (n_2376), .Y(n_2378));
OAI21X1 g65046(.A0 (g6167), .A1 (n_4324), .B0 (n_1776), .Y (n_2375));
MX2X1 g65072(.A (g_20614), .B (g_15758), .S0 (n_1491), .Y (n_2374));
XOR2X1 g65082(.A (n_1409), .B (n_650), .Y (n_2373));
OR2X1 g65240(.A (n_4329), .B (n_9772), .Y (n_2372));
OR2X1 g65242(.A (n_4327), .B (n_9772), .Y (n_2370));
OR2X1 g65244(.A (n_4320), .B (n_9772), .Y (n_2368));
OR2X1 g65247(.A (n_4314), .B (n_9772), .Y (n_2367));
OR2X1 g65250(.A (n_4322), .B (n_9772), .Y (n_2366));
OR2X1 g65251(.A (n_4324), .B (n_9772), .Y (n_2365));
OR2X1 g65270(.A (n_1493), .B (g5033), .Y (n_2364));
INVX1 g65282(.A (n_2640), .Y (n_2363));
INVX1 g65308(.A (n_2361), .Y (n_3073));
NAND2X1 g65332(.A (n_6705), .B (n_10687), .Y (n_2785));
OR2X1 g65347(.A (n_2008), .B (n_1729), .Y (n_2608));
NAND2X1 g65364(.A (g4477), .B (n_9836), .Y (n_2356));
NAND2X1 g65374(.A (n_1124), .B (n_9521), .Y (n_4939));
NAND4X1 g65385(.A (n_2443), .B (g5579), .C (g17813), .D (n_2208), .Y(n_2354));
NAND4X1 g65388(.A (n_2352), .B (g6271), .C (g17845), .D (n_11150), .Y(n_2353));
AND2X1 g65399(.A (n_2064), .B (n_1626), .Y (n_2351));
NAND3X1 g61946(.A (n_1995), .B (g_16456), .C (n_9311), .Y (n_2350));
NAND4X1 g65403(.A (n_2432), .B (g6617), .C (g17871), .D (n_11178), .Y(n_2349));
NOR2X1 g65409(.A (g16718), .B (n_2020), .Y (n_2348));
NOR2X1 g65413(.A (g16744), .B (n_2023), .Y (n_2347));
NAND2X1 g61950(.A (n_1644), .B (n_2345), .Y (n_2346));
NAND4X1 g65452(.A (n_10831), .B (g5196), .C (g13039), .D (g25219), .Y(n_2344));
NAND4X1 g65453(.A (n_2413), .B (g6235), .C (g13085), .D (n_11157), .Y(n_2343));
NAND4X1 g65454(.A (g6247), .B (n_3277), .C (g13085), .D (n_11150), .Y(n_2342));
NAND4X1 g65456(.A (g5224), .B (n_2339), .C (g17787), .D (g25219), .Y(n_2340));
NAND4X1 g65459(.A (g6609), .B (n_2600), .C (g17871), .D (n_11177), .Y(n_2338));
NAND4X1 g65460(.A (n_2439), .B (g5543), .C (g13049), .D (n_1023), .Y(n_2336));
NAND4X1 g65461(.A (g6597), .B (n_2600), .C (g17722), .D (n_11173), .Y(n_2334));
NAND4X1 g65462(.A (g5200), .B (n_2339), .C (g12238), .D (g25219), .Y(n_2332));
NAND4X1 g65474(.A (n_2597), .B (g5559), .C (g17604), .D (n_2208), .Y(n_2331));
NAND4X1 g65475(.A (g5555), .B (n_7150), .C (g13049), .D (n_2208), .Y(n_2329));
NAND4X1 g65478(.A (g5571), .B (n_2597), .C (g17813), .D (n_1023), .Y(n_2327));
NAND4X1 g65480(.A (g6251), .B (n_2325), .C (g17685), .D (n_11150), .Y(n_2326));
NAND4X1 g65482(.A (g6263), .B (n_2325), .C (g17845), .D (n_11157), .Y(n_2324));
NAND4X1 g65487(.A (g6593), .B (n_3275), .C (g13099), .D (n_11178), .Y(n_2323));
NAND4X1 g65488(.A (n_2435), .B (g6581), .C (g13099), .D (n_11184), .Y(n_2321));
INVX1 g65597(.A (g16659), .Y (n_2594));
INVX1 g65644(.A (n_3184), .Y (n_2320));
INVX1 g65688(.A (n_6395), .Y (n_2319));
NOR2X1 g65889(.A (n_10402), .B (n_9107), .Y (n_2316));
NAND2X1 g65896(.A (n_8809), .B (n_9351), .Y (n_2580));
INVX1 g65915(.A (n_3177), .Y (n_2577));
NAND2X1 g63196(.A (n_2312), .B (g4854), .Y (n_2925));
NOR2X1 g66376(.A (n_6324), .B (n_10078), .Y (n_2311));
XOR2X1 g66173(.A (n_8768), .B (n_8837), .Y (n_2310));
XOR2X1 g66182(.A (n_10196), .B (n_3849), .Y (n_2309));
NOR2X1 g66281(.A (n_6252), .B (n_10716), .Y (n_2308));
NAND2X1 g66286(.A (n_2306), .B (n_10078), .Y (n_2307));
INVX1 g66288(.A (n_2304), .Y (n_2305));
NOR2X1 g66291(.A (n_8799), .B (n_9193), .Y (n_2303));
NOR2X1 g66295(.A (g5352), .B (n_9107), .Y (n_2302));
NAND2X1 g66296(.A (g1361), .B (n_9628), .Y (n_2301));
NAND2X1 g66298(.A (g6505), .B (n_9599), .Y (n_2298));
NAND2X1 g66310(.A (n_1502), .B (n_9874), .Y (n_2562));
NAND2X1 g66317(.A (n_303), .B (n_9894), .Y (n_2847));
NOR2X1 g66321(.A (g_18308), .B (n_10078), .Y (n_2296));
NAND2X1 g66326(.A (n_2293), .B (n_10078), .Y (n_2294));
NOR2X1 g66327(.A (n_2290), .B (n_9129), .Y (n_2291));
NOR2X1 g66335(.A (g6044), .B (n_10078), .Y (n_2289));
NAND2X1 g66338(.A (g1373), .B (n_9599), .Y (n_2288));
NAND2X1 g66340(.A (g_19911), .B (n_9193), .Y (n_2286));
NAND2X1 g66341(.A (n_10499), .B (n_9353), .Y (n_2285));
NAND2X1 g66344(.A (g2629), .B (n_9775), .Y (n_2284));
NAND2X1 g66348(.A (g1379), .B (n_9353), .Y (n_2283));
NAND2X1 g66349(.A (n_2280), .B (n_9884), .Y (n_2281));
NAND2X1 g66351(.A (n_10119), .B (n_9300), .Y (n_2278));
NOR2X1 g66352(.A (g6390), .B (n_9371), .Y (n_2277));
NOR2X1 g66361(.A (g5029), .B (n_9672), .Y (n_2276));
NOR2X1 g66372(.A (g6736), .B (n_9903), .Y (n_2274));
NAND2X1 g66383(.A (g2070), .B (n_9884), .Y (n_2272));
NAND2X1 g66388(.A (n_383), .B (n_9894), .Y (n_2855));
NOR2X1 g66395(.A (n_6928), .B (n_9903), .Y (n_2271));
NOR2X1 g66396(.A (n_6057), .B (n_9129), .Y (n_2270));
NAND2X1 g66399(.A (g4388), .B (n_9884), .Y (n_2269));
NAND2X1 g66400(.A (n_261), .B (n_9894), .Y (n_2842));
NAND2X1 g66402(.A (n_1275), .B (n_9599), .Y (n_2268));
NAND2X1 g66403(.A (g1936), .B (n_9672), .Y (n_2266));
NOR2X1 g66404(.A (g_12922), .B (n_9129), .Y (n_2265));
NAND2X1 g66408(.A (n_388), .B (n_9883), .Y (n_2859));
NOR2X1 g66426(.A (g3698), .B (n_9903), .Y (n_2264));
NOR2X1 g66436(.A (n_10647), .B (n_9129), .Y (n_2263));
NOR2X1 g66466(.A (g_11293), .B (n_10782), .Y (n_2260));
NAND2X1 g66467(.A (n_2258), .B (n_9628), .Y (n_2259));
NAND2X1 g66468(.A (g_19233), .B (n_9599), .Y (n_2256));
NAND2X1 g66474(.A (g_21576), .B (n_10952), .Y (n_2255));
NAND2X1 g66476(.A (n_933), .B (n_10078), .Y (n_2254));
NOR2X1 g66477(.A (n_2252), .B (n_10782), .Y (n_2253));
NOR2X1 g66496(.A (g_15879), .B (n_9129), .Y (n_2250));
NOR2X1 g66514(.A (g_16311), .B (n_10782), .Y (n_2249));
NOR2X1 g66518(.A (g_16464), .B (n_9129), .Y (n_2248));
NAND2X1 g66524(.A (g2361), .B (n_9836), .Y (n_2247));
NOR2X1 g66534(.A (n_8793), .B (n_9129), .Y (n_2246));
NAND2X1 g66537(.A (n_2244), .B (n_9976), .Y (n_2245));
NAND2X1 g66539(.A (n_3383), .B (n_9193), .Y (n_2243));
NAND2X1 g66542(.A (n_4139), .B (n_9371), .Y (n_2242));
NOR2X1 g66546(.A (g5698), .B (n_10078), .Y (n_2241));
NOR2X1 g66554(.A (g4049), .B (n_10376), .Y (n_2239));
NOR2X1 g66556(.A (g3347), .B (n_9903), .Y (n_2237));
NAND2X1 g66562(.A (n_370), .B (n_9894), .Y (n_2853));
NAND2X1 g66574(.A (g4854), .B (n_9884), .Y (n_2234));
NAND2X1 g66581(.A (n_215), .B (n_9139), .Y (n_2857));
NOR2X1 g66594(.A (n_388), .B (n_9107), .Y (n_2233));
AND2X1 g66609(.A (g2823), .B (n_9091), .Y (n_2231));
NOR2X1 g66610(.A (g2518), .B (n_9693), .Y (n_2230));
NOR2X1 g66612(.A (g2384), .B (n_9903), .Y (n_2229));
AND2X1 g66616(.A (g5499), .B (n_9209), .Y (n_2228));
AND2X1 g66640(.A (g3143), .B (n_9521), .Y (n_2227));
NOR2X1 g66650(.A (n_303), .B (n_9903), .Y (n_2225));
NAND2X1 g66662(.A (n_2224), .B (n_9139), .Y (n_2838));
NOR2X1 g66671(.A (n_215), .B (n_9775), .Y (n_2223));
NOR2X1 g66678(.A (n_10307), .B (n_10078), .Y (n_2221));
NOR2X1 g66679(.A (n_330), .B (n_9884), .Y (n_2219));
AND2X1 g66683(.A (g5845), .B (n_9521), .Y (n_2218));
NOR2X1 g66685(.A (g1467), .B (n_9353), .Y (n_2216));
AND2X1 g66689(.A (n_10813), .B (n_9521), .Y (n_2215));
NAND2X1 g66700(.A (n_11171), .B (n_9883), .Y (n_2835));
NOR2X1 g66706(.A (g1959), .B (n_9693), .Y (n_2212));
AND2X1 g66719(.A (g3845), .B (n_9521), .Y (n_2211));
NOR2X1 g66726(.A (g1454), .B (n_9107), .Y (n_2210));
NAND4X1 g64872(.A (n_2439), .B (g5595), .C (g14635), .D (n_2208), .Y(n_2209));
AND2X1 g66776(.A (g3494), .B (n_9139), .Y (n_2207));
AND2X1 g66790(.A (g6191), .B (n_9311), .Y (n_2206));
NOR2X1 g66812(.A (g1437), .B (n_9353), .Y (n_2205));
NOR2X1 g66859(.A (n_6527), .B (n_9599), .Y (n_2496));
NAND2X1 g66882(.A (n_5402), .B (n_9139), .Y (n_2828));
AND2X1 g66888(.A (g6537), .B (n_9521), .Y (n_2204));
NOR2X1 g66900(.A (n_370), .B (n_10078), .Y (n_2203));
OR2X1 g61528(.A (n_2192), .B (n_129), .Y (n_2790));
XOR2X1 g63640(.A (g20557), .B (n_1581), .Y (n_2182));
XOR2X1 g63643(.A (g4273), .B (n_1583), .Y (n_2181));
NAND2X1 g61201(.A (n_1277), .B (n_11073), .Y (n_2180));
NAND2X1 g61202(.A (n_11073), .B (n_2177), .Y (n_2178));
NAND2X1 g61204(.A (n_11073), .B (n_6782), .Y (n_2176));
INVX1 g61207(.A (n_11041), .Y (n_2830));
INVX1 g62287(.A (n_1883), .Y (n_2174));
INVX1 g62289(.A (n_1882), .Y (n_2173));
INVX1 g61218(.A (n_2592), .Y (n_2172));
AOI21X1 g64681(.A0 (n_1546), .A1 (n_1312), .B0 (n_2111), .Y (g31521));
NOR2X1 g66856(.A (g1825), .B (n_10376), .Y (n_2168));
OAI21X1 g64146(.A0 (n_692), .A1 (n_11162), .B0 (n_1860), .Y (n_2167));
OR2X1 g64147(.A (n_2165), .B (n_221), .Y (n_2166));
NAND2X1 g64258(.A (n_1700), .B (n_1847), .Y (n_2163));
OAI21X1 g62657(.A0 (n_1840), .A1 (g4664), .B0 (n_2867), .Y (n_2161));
MX2X1 g64424(.A (g_21806), .B (g_20837), .S0 (n_6460), .Y (n_2160));
MX2X1 g64431(.A (g_22379), .B (g_21806), .S0 (n_6460), .Y (n_2159));
MX2X1 g64434(.A (g_21576), .B (g_22379), .S0 (n_6460), .Y (n_2157));
MX2X1 g64457(.A (g_6131), .B (g_19241), .S0 (n_6460), .Y (n_2156));
MX2X1 g64459(.A (n_5663), .B (g_6131), .S0 (n_6460), .Y (n_2155));
AND2X1 g64512(.A (n_1817), .B (n_6464), .Y (n_3174));
NAND3X1 g64555(.A (n_2153), .B (n_2457), .C (n_2747), .Y (n_2154));
NOR2X1 g64605(.A (n_2106), .B (n_8637), .Y (n_2483));
NAND4X1 g64633(.A (n_335), .B (n_17), .C (n_943), .D (n_353), .Y(n_2152));
AOI21X1 g64646(.A0 (n_1013), .A1 (n_2150), .B0 (n_1559), .Y (n_2151));
NAND4X1 g64693(.A (n_2133), .B (n_2439), .C (g14694), .D (g5583), .Y(n_2149));
NAND4X1 g64696(.A (n_2119), .B (n_2435), .C (g14828), .D (g6621), .Y(n_2148));
NAND4X1 g64700(.A (n_10877), .B (g3586), .C (g16744), .D (n_6973), .Y(n_2146));
NAND4X1 g64717(.A (n_2143), .B (g5244), .C (g17674), .D (g25114), .Y(n_2145));
NAND4X1 g64718(.A (n_2143), .B (g5228), .C (g14662), .D (n_10621), .Y(n_2144));
NAND4X1 g64724(.A (n_2131), .B (n_2352), .C (g17760), .D (g6283), .Y(n_2141));
NAND4X1 g64725(.A (n_10879), .B (g3594), .C (g16744), .D (n_11128),.Y (n_2140));
NAND4X1 g64727(.A (n_10877), .B (g3570), .C (g13926), .D (n_4682), .Y(n_2138));
NAND4X1 g64730(.A (n_2447), .B (g3921), .C (g13966), .D (n_6787), .Y(n_2137));
NAND4X1 g64744(.A (n_2133), .B (g5615), .C (g17580), .D (n_7150), .Y(n_2135));
NAND4X1 g64746(.A (n_2133), .B (g5599), .C (g17711), .D (n_2597), .Y(n_2134));
NAND4X1 g64752(.A (n_2131), .B (g6267), .C (g14779), .D (n_3277), .Y(n_2132));
NAND4X1 g64753(.A (n_2131), .B (n_2413), .C (g17649), .D (g6299), .Y(n_2130));
NAND4X1 g64754(.A (n_2127), .B (n_10809), .C (g17607), .D (g5953), .Y(n_2129));
NAND4X1 g64755(.A (n_2127), .B (g5921), .C (g14738), .D (n_10506), .Y(n_2128));
NAND4X1 g64756(.A (n_2127), .B (n_10622), .C (g17739), .D (g5937), .Y(n_2126));
NAND4X1 g64764(.A (n_2119), .B (g6653), .C (g17688), .D (n_3275), .Y(n_2122));
NAND4X1 g64765(.A (n_2143), .B (n_10831), .C (g17519), .D (g5260), .Y(n_2121));
NAND4X1 g64767(.A (n_2119), .B (g6637), .C (g17778), .D (n_2600), .Y(n_2120));
NOR2X1 g65294(.A (g26801), .B (n_9856), .Y (n_2973));
NOR2X1 g64875(.A (n_2458), .B (n_10725), .Y (n_2118));
AND2X1 g64877(.A (n_3021), .B (n_2115), .Y (n_3047));
AND2X1 g64884(.A (n_2113), .B (n_2115), .Y (n_2116));
AND2X1 g64886(.A (n_3021), .B (n_2113), .Y (n_2114));
OR2X1 g64894(.A (n_1737), .B (n_2111), .Y (n_3897));
NOR2X1 g64895(.A (n_1552), .B (g8788), .Y (n_2110));
NOR2X1 g64902(.A (n_10551), .B (n_10552), .Y (n_2107));
INVX1 g64922(.A (n_2106), .Y (n_2410));
NAND4X1 g64955(.A (n_1544), .B (g4087), .C (g4076), .D (g4098), .Y(n_2103));
AND2X1 g64963(.A (n_1555), .B (n_2113), .Y (n_2456));
AOI21X1 g64981(.A0 (n_397), .A1 (n_10499), .B0 (n_10725), .Y(n_2654));
INVX1 g65012(.A (n_2100), .Y (n_2101));
XOR2X1 g65042(.A (g1677), .B (n_1248), .Y (n_2099));
OAI21X1 g65043(.A0 (g5475), .A1 (n_4329), .B0 (n_1535), .Y (n_2098));
OAI21X1 g65044(.A0 (g5821), .A1 (n_4327), .B0 (n_1545), .Y (n_2097));
XOR2X1 g65045(.A (g1811), .B (n_1237), .Y (n_2096));
OAI21X1 g65048(.A0 (g6513), .A1 (n_4322), .B0 (n_1553), .Y (n_2095));
XOR2X1 g65049(.A (g1945), .B (n_1231), .Y (n_2094));
OAI21X1 g65053(.A0 (g3821), .A1 (n_4314), .B0 (n_1547), .Y (n_2093));
OAI21X1 g65054(.A0 (g3119), .A1 (n_4316), .B0 (n_1539), .Y (n_2092));
OAI21X1 g65055(.A0 (g3470), .A1 (n_4320), .B0 (n_1551), .Y (n_2091));
XOR2X1 g65056(.A (n_7260), .B (n_6582), .Y (n_2090));
XOR2X1 g65057(.A (g2370), .B (n_1161), .Y (n_2089));
XOR2X1 g65059(.A (g2504), .B (n_1139), .Y (n_2088));
XOR2X1 g65060(.A (g5128), .B (g26801), .Y (n_2087));
MX2X1 g65061(.A (n_2936), .B (g6159), .S0 (n_4324), .Y (n_2086));
MX2X1 g65066(.A (n_2704), .B (n_2084), .S0 (n_4324), .Y (n_2085));
MX2X1 g65077(.A (n_1732), .B (n_6958), .S0 (n_1731), .Y (n_2083));
XOR2X1 g65083(.A (n_10550), .B (n_10568), .Y (n_2082));
XOR2X1 g65089(.A (g2638), .B (n_1014), .Y (n_2081));
XOR2X1 g65093(.A (g2079), .B (n_1304), .Y (n_2080));
XOR2X1 g65095(.A (g2236), .B (n_1168), .Y (n_2079));
NOR2X1 g65235(.A (n_389), .B (n_2077), .Y (n_2078));
NOR2X1 g65239(.A (n_202), .B (n_10475), .Y (n_2072));
NAND2X1 g65256(.A (n_1662), .B (g5033), .Y (n_2070));
AND2X1 g65261(.A (n_2067), .B (n_8694), .Y (n_2069));
AND2X1 g65263(.A (n_2067), .B (n_8777), .Y (n_2068));
NOR2X1 g66777(.A (n_708), .B (n_10078), .Y (n_3857));
OR2X1 g65283(.A (n_11027), .B (n_1652), .Y (n_2640));
AND2X1 g65285(.A (n_10184), .B (n_2064), .Y (n_2065));
NAND2X1 g65299(.A (n_2062), .B (g1306), .Y (n_2063));
INVX1 g65309(.A (n_2061), .Y (n_2361));
OR2X1 g61396(.A (n_2060), .B (n_26), .Y (n_2671));
NAND2X1 g65338(.A (n_10200), .B (n_9651), .Y (n_2784));
INVX1 g65359(.A (n_2056), .Y (n_2057));
NOR2X1 g65367(.A (n_1462), .B (n_7260), .Y (n_2055));
INVX1 g65368(.A (n_2053), .Y (n_2054));
NOR2X1 g65390(.A (n_10527), .B (g_8896), .Y (n_2639));
NAND2X1 g65394(.A (n_8906), .B (n_2067), .Y (n_2051));
AND2X1 g65395(.A (n_2067), .B (n_8809), .Y (n_2049));
NAND2X1 g65400(.A (n_10205), .B (n_2064), .Y (n_2048));
AND2X1 g65401(.A (n_2064), .B (n_10296), .Y (n_2046));
AND2X1 g65404(.A (n_2045), .B (n_2044), .Y (n_3984));
INVX1 g65417(.A (n_2427), .Y (n_2043));
INVX1 g65427(.A (n_10765), .Y (n_2042));
NAND4X1 g65449(.A (g5208), .B (n_10621), .C (g13039), .D (n_1695), .Y(n_2038));
AOI22X1 g65464(.A0 (n_10206), .A1 (g4888), .B0 (g4955), .B1(n_10214), .Y (n_11192));
AOI22X1 g65466(.A0 (g4917), .A1 (n_10214), .B0 (g4912), .B1(n_10206), .Y (n_2034));
MX2X1 g61964(.A (n_2429), .B (g_19172), .S0 (n_2878), .Y (n_2032));
NAND4X1 g65476(.A (g5212), .B (n_2339), .C (g17577), .D (n_1695), .Y(n_2031));
NAND4X1 g65479(.A (g6239), .B (n_2325), .C (g12422), .D (n_11157), .Y(n_2030));
NAND4X1 g65484(.A (g5893), .B (n_11101), .C (g12350), .D (n_546), .Y(n_2029));
NAND4X1 g65485(.A (g5917), .B (n_11101), .C (g17819), .D (n_546), .Y(n_2027));
NAND4X1 g65486(.A (n_10808), .B (g5889), .C (g13068), .D (n_546), .Y(n_2025));
AOI21X1 g65504(.A0 (n_8917), .A1 (g4049), .B0 (n_1479), .Y (n_2024));
NOR2X1 g65689(.A (n_2019), .B (n_4878), .Y (n_6395));
AND2X1 g65727(.A (n_2600), .B (n_9091), .Y (n_2018));
NAND2X1 g65645(.A (n_2001), .B (n_2017), .Y (n_3184));
NAND2X1 g65794(.A (n_11126), .B (n_10687), .Y (n_2016));
AND2X1 g65796(.A (n_2325), .B (n_10687), .Y (n_2015));
NAND2X1 g65798(.A (n_8572), .B (n_9311), .Y (n_2014));
CLKBUFX1 gbuf_d_1082(.A(g7946), .Y(d_out_1082));
CLKBUFX1 gbuf_q_1082(.A(q_in_1082), .Y(g8475));
AND2X1 g65838(.A (n_11101), .B (n_9521), .Y (n_2011));
NAND2X1 g65843(.A (n_6808), .B (n_10687), .Y (n_2009));
INVX1 g65847(.A (n_2008), .Y (n_4632));
AND2X1 g65865(.A (n_2597), .B (n_9750), .Y (n_2007));
OR2X1 g65866(.A (n_1628), .B (n_2005), .Y (n_2006));
NOR2X1 g65878(.A (g4927), .B (n_1625), .Y (n_2004));
INVX1 g62034(.A (n_2002), .Y (n_2003));
NAND3X1 g65970(.A (n_2001), .B (n_488), .C (n_10524), .Y (n_3718));
NAND2X1 g66747(.A (n_2556), .B (n_9501), .Y (n_2000));
MX2X1 g66125(.A (g1521), .B (g1532), .S0 (n_3849), .Y (n_1997));
INVX1 g62062(.A (n_1995), .Y (n_1996));
INVX1 g62068(.A (n_1993), .Y (n_1994));
MX2X1 g66104(.A (g1178), .B (g1189), .S0 (n_8837), .Y (n_1992));
MX2X1 g66150(.A (g_20614), .B (g1178), .S0 (n_8837), .Y (n_1991));
OAI21X1 g63528(.A0 (n_1307), .A1 (g4659), .B0 (n_1329), .Y (n_1989));
NOR2X1 g66289(.A (n_1627), .B (n_9884), .Y (n_2304));
NAND2X1 g66324(.A (n_330), .B (n_9521), .Y (n_2578));
OR2X1 g66360(.A (g4467), .B (n_9628), .Y (n_2862));
INVX1 g66363(.A (n_1985), .Y (n_1986));
OR2X1 g66527(.A (g1306), .B (n_10078), .Y (n_2480));
NAND2X1 g66583(.A (n_8588), .B (n_9351), .Y (n_2661));
NAND2X1 g66585(.A (g1542), .B (n_9521), .Y (n_1982));
NAND2X1 g66589(.A (n_11157), .B (n_9139), .Y (n_2606));
INVX1 g66592(.A (n_5453), .Y (n_1980));
NAND2X1 g66623(.A (g1199), .B (n_9894), .Y (n_1979));
NAND2X1 g66628(.A (n_10894), .B (n_9351), .Y (n_2668));
NOR2X1 g66677(.A (n_10503), .B (n_9526), .Y (n_2657));
NAND2X1 g66680(.A (n_2376), .B (n_9883), .Y (n_2612));
NAND2X1 g66705(.A (n_2280), .B (n_9501), .Y (n_1977));
NAND2X1 g66713(.A (g_18739), .B (n_9139), .Y (n_1976));
OR2X1 g65414(.A (n_1426), .B (n_8809), .Y (n_1975));
NOR2X1 g66749(.A (n_6782), .B (n_9856), .Y (n_3372));
NOR2X1 g66773(.A (g4332), .B (n_662), .Y (n_1972));
NAND2X1 g66785(.A (g4608), .B (n_9627), .Y (n_1971));
NAND2X1 g66826(.A (n_2529), .B (n_9521), .Y (n_1969));
AND2X1 g66829(.A (g2827), .B (n_10687), .Y (n_1968));
OR2X1 g64846(.A (n_10520), .B (n_2017), .Y (n_1887));
AOI21X1 g62278(.A0 (n_11029), .A1 (g3343), .B0 (n_1473), .Y (n_1885));
AOI21X1 g62279(.A0 (n_10576), .A1 (g3694), .B0 (n_1474), .Y (n_1884));
INVX1 g68049(.A (n_2224), .Y (n_2734));
AOI21X1 g62288(.A0 (n_10941), .A1 (g3347), .B0 (n_1311), .Y (n_1883));
AOI21X1 g62290(.A0 (n_6972), .A1 (g3698), .B0 (n_1310), .Y (n_1882));
AND2X1 g61219(.A (n_1443), .B (n_10329), .Y (n_2592));
CLKBUFX1 gbuf_d_1083(.A(g7916), .Y(d_out_1083));
CLKBUFX1 gbuf_q_1083(.A(q_in_1083), .Y(g8416));
INVX1 g64144(.A (n_2312), .Y (n_1875));
MX2X1 g61296(.A (n_460), .B (g1521), .S0 (n_3849), .Y (n_1869));
NAND2X1 g66478(.A (g_5342), .B (n_9091), .Y (n_1865));
NAND4X1 g64525(.A (n_235), .B (n_157), .C (n_958), .D (n_194), .Y(n_1863));
NAND4X1 g64594(.A (n_425), .B (n_29), .C (n_950), .D (n_428), .Y(n_1862));
NAND4X1 g64619(.A (n_340), .B (n_5), .C (n_947), .D (n_248), .Y(n_1861));
AOI22X1 g64680(.A0 (n_694), .A1 (g_21720), .B0 (n_693), .B1(g_19233), .Y (n_1860));
NAND4X1 g64692(.A (n_1854), .B (n_10833), .C (g14662), .D (g5236), .Y(n_1859));
NAND4X1 g64694(.A (n_1848), .B (n_2413), .C (g14779), .D (g6275), .Y(n_1858));
NAND4X1 g64695(.A (n_1845), .B (n_10809), .C (g14738), .D (g5929), .Y(n_1857));
NAND4X1 g64712(.A (n_1854), .B (g5252), .C (g17674), .D (n_2339), .Y(n_1855));
NAND4X1 g64713(.A (n_1854), .B (g5268), .C (g17519), .D (n_10621), .Y(n_11194));
NAND4X1 g64715(.A (n_8548), .B (g3227), .C (g13895), .D (n_11029), .Y(n_6948));
NAND4X1 g64733(.A (n_6806), .B (g3929), .C (g13966), .D (n_4988), .Y(n_1851));
NAND4X1 g64738(.A (n_10879), .B (g3578), .C (g13926), .D (n_10576),.Y (n_1850));
NAND4X1 g64750(.A (n_1848), .B (g6291), .C (g17760), .D (n_2325), .Y(n_1849));
NAND4X1 g64751(.A (n_1848), .B (g6307), .C (g17649), .D (n_3277), .Y(n_1847));
NAND4X1 g64757(.A (n_1845), .B (g5945), .C (g17739), .D (n_11101), .Y(n_1846));
NAND4X1 g64758(.A (n_1845), .B (g5961), .C (g17607), .D (n_10508), .Y(n_1844));
MX2X1 g65074(.A (n_2923), .B (g3813), .S0 (n_4314), .Y (n_1843));
XOR2X1 g64775(.A (n_307), .B (n_474), .Y (n_1842));
NAND2X1 g62798(.A (n_1840), .B (g4664), .Y (n_2867));
XOR2X1 g64776(.A (g4269), .B (n_1582), .Y (n_1839));
OAI22X1 g64777(.A0 (n_821), .A1 (n_1831), .B0 (n_747), .B1 (g4593),.Y (n_1838));
NAND3X1 g64889(.A (n_991), .B (n_6762), .C (g7916), .Y (n_1833));
AND2X1 g64900(.A (n_1096), .B (n_1831), .Y (n_1832));
INVX1 g64904(.A (n_10597), .Y (n_1830));
OR2X1 g64923(.A (n_10907), .B (g4688), .Y (n_2106));
OR2X1 g64925(.A (n_1016), .B (n_1826), .Y (n_1827));
AOI22X1 g65465(.A0 (g4933), .A1 (n_10185), .B0 (g4944), .B1(n_10998), .Y (n_11193));
AOI21X1 g64994(.A0 (g_13758), .A1 (n_3550), .B0 (n_1291), .Y(n_1822));
OAI21X1 g65007(.A0 (n_1820), .A1 (g8839), .B0 (n_1278), .Y (n_1821));
XOR2X1 g65013(.A (g4527), .B (n_1562), .Y (n_2100));
AOI21X1 g65014(.A0 (n_1818), .A1 (g34036), .B0 (n_994), .Y (n_1819));
MX2X1 g65020(.A (n_6501), .B (n_924), .S0 (n_11051), .Y (n_1817));
MX2X1 g65062(.A (n_2718), .B (n_1813), .S0 (n_1812), .Y (n_1814));
MX2X1 g65063(.A (n_3011), .B (n_1810), .S0 (n_4329), .Y (n_1811));
MX2X1 g65064(.A (n_2940), .B (g5813), .S0 (n_4327), .Y (n_1809));
MX2X1 g65065(.A (n_2684), .B (n_1807), .S0 (n_4327), .Y (n_1808));
MX2X1 g65067(.A (n_2686), .B (n_1805), .S0 (n_4316), .Y (n_1806));
MX2X1 g65068(.A (n_2005), .B (g1489), .S0 (n_4617), .Y (n_1804));
MX2X1 g65069(.A (n_2930), .B (g6505), .S0 (n_4322), .Y (n_1803));
MX2X1 g65070(.A (n_3253), .B (g3111), .S0 (n_4316), .Y (n_1802));
MX2X1 g65071(.A (n_2928), .B (g3462), .S0 (n_4320), .Y (n_1801));
MX2X1 g65073(.A (n_2699), .B (n_1799), .S0 (n_4320), .Y (n_1800));
MX2X1 g65075(.A (n_2943), .B (g5467), .S0 (n_4329), .Y (n_1798));
MX2X1 g65076(.A (n_2692), .B (n_1796), .S0 (n_4314), .Y (n_1797));
MX2X1 g65078(.A (n_3007), .B (n_1794), .S0 (n_4322), .Y (n_1795));
MX2X1 g65079(.A (g1442), .B (n_2005), .S0 (n_4617), .Y (n_1793));
MX2X1 g65080(.A (g5156), .B (g5120), .S0 (n_1812), .Y (n_1792));
AOI21X1 g65085(.A0 (n_720), .A1 (n_564), .B0 (n_1251), .Y (n_1791));
CLKBUFX1 gbuf_d_1084(.A(g14597), .Y(d_out_1084));
CLKBUFX1 gbuf_q_1084(.A(q_in_1084), .Y(g17639));
CLKBUFX1 gbuf_d_1085(.A(g14635), .Y(d_out_1085));
CLKBUFX1 gbuf_q_1085(.A(q_in_1085), .Y(g17678));
CLKBUFX1 gbuf_d_1086(.A(g14673), .Y(d_out_1086));
CLKBUFX1 gbuf_q_1086(.A(q_in_1086), .Y(g17715));
CLKBUFX1 gbuf_d_1087(.A(g14705), .Y(d_out_1087));
CLKBUFX1 gbuf_q_1087(.A(q_in_1087), .Y(g17743));
CLKBUFX1 gbuf_d_1088(.A(g14749), .Y(d_out_1088));
CLKBUFX1 gbuf_q_1088(.A(q_in_1088), .Y(g17764));
NOR2X1 g65232(.A (n_3030), .B (n_1250), .Y (n_1789));
NOR2X1 g65233(.A (n_1266), .B (n_1631), .Y (n_1788));
NOR2X1 g65234(.A (n_1405), .B (g_15380), .Y (n_1787));
AND2X1 g65246(.A (n_10984), .B (n_8676), .Y (n_1786));
AND2X1 g65249(.A (n_8639), .B (n_10905), .Y (n_1785));
NAND2X1 g65252(.A (n_6582), .B (n_7260), .Y (n_2165));
NOR2X1 g65253(.A (n_6578), .B (n_1220), .Y (n_1783));
OR2X1 g65255(.A (n_7010), .B (g5033), .Y (n_6970));
NAND2X1 g65257(.A (n_1765), .B (n_1391), .Y (n_1780));
NAND2X1 g65258(.A (n_1770), .B (n_1471), .Y (n_1779));
NAND2X1 g65259(.A (n_1772), .B (n_1777), .Y (n_1778));
NAND2X1 g65262(.A (g6167), .B (n_4324), .Y (n_1776));
NAND2X1 g65268(.A (n_1763), .B (n_1480), .Y (n_1775));
NAND2X1 g65274(.A (n_1772), .B (n_1476), .Y (n_1773));
NAND2X1 g65284(.A (n_1770), .B (n_1377), .Y (n_1771));
NAND2X1 g65286(.A (n_1767), .B (n_1584), .Y (n_1769));
NAND2X1 g65287(.A (n_1767), .B (n_1370), .Y (n_1768));
NAND2X1 g65290(.A (n_1765), .B (n_1445), .Y (n_1766));
NAND2X1 g65291(.A (n_1763), .B (n_1762), .Y (n_1764));
NAND2X1 g65295(.A (n_1772), .B (n_973), .Y (n_1761));
NAND2X1 g65300(.A (n_1767), .B (n_1758), .Y (n_1759));
INVX1 g65302(.A (n_1756), .Y (n_1757));
NAND2X1 g65304(.A (n_1727), .B (n_1382), .Y (n_1755));
OR2X1 g65310(.A (n_10983), .B (g4878), .Y (n_2061));
NAND2X1 g65314(.A (n_1752), .B (n_1450), .Y (n_1754));
NAND2X1 g65316(.A (n_1752), .B (n_1751), .Y (n_1753));
NAND2X1 g65317(.A (n_1752), .B (n_1367), .Y (n_1750));
NAND2X1 g65319(.A (n_1752), .B (n_1206), .Y (n_1749));
NAND2X1 g65322(.A (n_1767), .B (n_1242), .Y (n_1748));
AND2X1 g65325(.A (n_10214), .B (n_8676), .Y (n_1747));
NAND2X1 g65330(.A (n_1744), .B (n_1440), .Y (n_1746));
NAND2X1 g65331(.A (n_1744), .B (n_1743), .Y (n_1745));
NAND2X1 g65334(.A (n_1744), .B (n_1364), .Y (n_1741));
NAND2X1 g65335(.A (n_1744), .B (n_1184), .Y (n_1740));
NAND2X1 g65341(.A (n_1763), .B (n_970), .Y (n_1738));
INVX1 g65342(.A (n_1737), .Y (n_2403));
INVX1 g65344(.A (n_2677), .Y (n_1736));
NAND2X1 g65357(.A (n_918), .B (n_10949), .Y (n_2449));
NAND3X1 g65361(.A (n_1219), .B (n_7260), .C (n_1734), .Y (n_1735));
NOR2X1 g65362(.A (n_1732), .B (n_1731), .Y (n_1733));
NAND2X1 g65363(.A (n_1765), .B (n_590), .Y (n_1730));
NOR2X1 g65369(.A (n_1729), .B (n_1238), .Y (n_2053));
NAND2X1 g65376(.A (n_1727), .B (n_1245), .Y (n_1728));
NAND2X1 g65377(.A (n_1727), .B (n_1725), .Y (n_1726));
NAND2X1 g65378(.A (n_1770), .B (n_1723), .Y (n_1724));
NAND2X1 g65382(.A (n_1727), .B (n_1455), .Y (n_1722));
NAND2X1 g65384(.A (n_1770), .B (n_1264), .Y (n_1721));
NAND2X1 g65387(.A (n_1765), .B (n_1718), .Y (n_1719));
NAND4X1 g65392(.A (n_10623), .B (g5925), .C (g17819), .D (n_423), .Y(n_1717));
NAND2X1 g65398(.A (n_1772), .B (n_1411), .Y (n_1716));
AOI22X1 g65408(.A0 (n_790), .A1 (n_1714), .B0 (n_1713), .B1 (n_808),.Y (n_1715));
AOI22X1 g65410(.A0 (n_805), .A1 (n_1711), .B0 (n_1710), .B1 (n_798),.Y (n_1712));
NAND3X1 g65411(.A (n_10827), .B (n_746), .C (n_8796), .Y (n_1709));
AOI22X1 g65415(.A0 (n_697), .A1 (n_1706), .B0 (n_1705), .B1 (n_778),.Y (n_1707));
AOI22X1 g65421(.A0 (n_707), .A1 (n_1703), .B0 (n_1702), .B1 (n_793),.Y (n_1704));
NAND3X1 g65423(.A (n_2443), .B (n_1484), .C (g5619), .Y (n_1701));
NAND3X1 g65424(.A (n_2352), .B (n_1457), .C (g6311), .Y (n_1700));
NAND3X1 g65425(.A (n_10622), .B (n_1458), .C (g5965), .Y (n_1699));
NAND3X1 g65426(.A (n_2432), .B (n_1461), .C (g6657), .Y (n_1698));
NAND4X1 g65439(.A (g5232), .B (n_1695), .C (g17787), .D (g25114), .Y(n_1696));
NAND4X1 g65447(.A (g5905), .B (n_11101), .C (g17646), .D (n_423), .Y(n_1694));
NAND4X1 g65450(.A (g3542), .B (n_10895), .C (g11388), .D (n_11128),.Y (n_1691));
AOI22X1 g65455(.A0 (n_1062), .A1 (n_1688), .B0 (n_1687), .B1 (n_648),.Y (n_1689));
NAND4X1 g65457(.A (g3893), .B (n_5402), .C (g11418), .D (n_6808), .Y(n_1686));
AOI22X1 g65467(.A0 (g4907), .A1 (n_10185), .B0 (g4922), .B1(n_10998), .Y (n_1682));
AOI22X1 g65468(.A0 (g4743), .A1 (n_8810), .B0 (g4754), .B1 (n_8693),.Y (n_1681));
AOI22X1 g65469(.A0 (g4722), .A1 (n_10227), .B0 (g4727), .B1 (n_8778),.Y (n_1680));
AOI22X1 g65470(.A0 (n_1059), .A1 (n_1677), .B0 (n_1676), .B1 (n_591),.Y (n_1678));
AOI22X1 g65471(.A0 (g4717), .A1 (n_8810), .B0 (g4732), .B1 (n_8693),.Y (n_1675));
AOI22X1 g65472(.A0 (n_10227), .A1 (g4698), .B0 (g4765), .B1 (n_8778),.Y (n_1674));
AOI22X1 g65481(.A0 (n_1064), .A1 (n_1671), .B0 (n_1670), .B1 (n_486),.Y (n_1672));
NAND4X1 g65483(.A (g5901), .B (n_10506), .C (g13068), .D (n_423), .Y(n_1669));
INVX1 g65508(.A (n_2119), .Y (n_2433));
AOI22X1 g65448(.A0 (n_1667), .A1 (n_1666), .B0 (n_1665), .B1 (n_562),.Y (n_1668));
INVX1 g65592(.A (g16627), .Y (n_2023));
INVX1 g65610(.A (g16603), .Y (n_2020));
NAND3X1 g65707(.A (n_11113), .B (n_1352), .C (n_2017), .Y (n_1658));
OR2X1 g65784(.A (g4417), .B (n_5378), .Y (n_1657));
NAND2X1 g65848(.A (n_978), .B (g13272), .Y (n_2008));
INVX1 g65871(.A (n_1655), .Y (n_1656));
CLKBUFX1 g65917(.A (n_1652), .Y (n_3177));
NAND2X1 g65948(.A (n_817), .B (n_822), .Y (n_1650));
NAND2X1 g65961(.A (n_983), .B (n_795), .Y (n_1649));
NOR2X1 g62035(.A (n_2878), .B (n_799), .Y (n_2002));
INVX1 g62040(.A (n_1646), .Y (n_1647));
OR2X1 g62043(.A (n_2878), .B (g_19172), .Y (n_1645));
NAND2X1 g62044(.A (n_2878), .B (n_2429), .Y (n_1644));
OAI21X1 g66013(.A0 (g17604), .A1 (g13049), .B0 (n_1054), .Y (n_1643));
OAI21X1 g66015(.A0 (g17577), .A1 (g13039), .B0 (n_1094), .Y (n_1642));
OAI21X1 g66024(.A0 (g17685), .A1 (g13085), .B0 (n_1046), .Y (n_1641));
OAI21X1 g66042(.A0 (g17722), .A1 (g13099), .B0 (n_1021), .Y (n_1640));
NAND2X1 g62063(.A (n_4761), .B (n_1599), .Y (n_1995));
CLKBUFX1 gbuf_d_1089(.A(g16775), .Y(d_out_1089));
CLKBUFX1 gbuf_q_1089(.A(q_in_1089), .Y(g16659));
AND2X1 g65418(.A (n_1188), .B (n_1636), .Y (n_2427));
OR2X1 g66328(.A (g5084), .B (n_9836), .Y (n_5514));
OR2X1 g66364(.A (n_10123), .B (n_10376), .Y (n_1985));
OR2X1 g66462(.A (g_15758), .B (n_9371), .Y (n_2481));
NAND2X1 g66498(.A (n_35), .B (n_11055), .Y (n_1633));
NAND3X1 g64878(.A (n_1554), .B (n_1631), .C (n_1630), .Y (n_1632));
NOR2X1 g66593(.A (n_596), .B (n_9884), .Y (n_5453));
INVX1 g66595(.A (n_1628), .Y (n_1629));
NAND2X1 g66626(.A (n_1627), .B (n_9311), .Y (n_3192));
INVX1 g66631(.A (n_1625), .Y (n_1626));
NAND2X1 g65405(.A (n_1763), .B (n_1402), .Y (n_1605));
OAI21X1 g61588(.A0 (n_705), .A1 (g_15287), .B0 (g12919), .Y (n_2192));
NAND2X1 g62069(.A (n_4764), .B (n_1599), .Y (n_1993));
AND2X1 g63895(.A (n_2938), .B (n_1328), .Y (n_1597));
AND2X1 g64145(.A (n_1826), .B (g4849), .Y (n_2312));
NAND2X1 g64243(.A (n_1300), .B (n_1271), .Y (n_1592));
OR4X1 g65365(.A (g1333), .B (g19357), .C (g13272), .D (n_568), .Y(n_1591));
XOR2X1 g64779(.A (g5097), .B (n_1580), .Y (n_1590));
NOR2X1 g65360(.A (n_1729), .B (n_1422), .Y (n_2056));
CLKBUFX1 g68050(.A (n_1023), .Y (n_2224));
NAND3X1 g64593(.A (n_11217), .B (g3558), .C (n_6973), .Y (n_1587));
NAND3X1 g64628(.A (g3207), .B (n_801), .C (n_10941), .Y (n_1586));
NOR2X1 g65303(.A (n_1252), .B (n_1729), .Y (n_1756));
NAND2X1 g65699(.A (n_1243), .B (n_1584), .Y (n_1585));
AND2X1 g64847(.A (n_1582), .B (g4269), .Y (n_1583));
AND2X1 g64848(.A (n_1580), .B (g5097), .Y (n_1581));
INVX1 g65693(.A (n_1576), .Y (n_2064));
NAND3X1 g64936(.A (n_824), .B (g5216), .C (g25114), .Y (n_1575));
NAND3X1 g64940(.A (n_819), .B (n_2352), .C (g6255), .Y (n_1574));
XOR2X1 g65009(.A (g9251), .B (n_1570), .Y (n_1571));
NAND3X1 g61365(.A (g19357), .B (n_415), .C (n_635), .Y (n_1569));
AOI22X1 g65021(.A0 (n_636), .A1 (g_15740), .B0 (n_588), .B1 (n_708),.Y (n_1568));
AOI22X1 g65025(.A0 (n_1290), .A1 (g_22379), .B0 (n_691), .B1(g_19113), .Y (n_1567));
AND2X1 g65226(.A (n_10984), .B (g4955), .Y (n_1564));
NAND2X1 g65227(.A (n_1562), .B (n_162), .Y (n_1563));
AOI21X1 g65229(.A0 (n_268), .A1 (n_4980), .B0 (g4760), .Y (n_1561));
AOI21X1 g65231(.A0 (n_524), .A1 (n_11070), .B0 (g4894), .Y (n_1560));
XOR2X1 g65008(.A (g9019), .B (n_1556), .Y (n_1557));
AND2X1 g65277(.A (n_1554), .B (n_1631), .Y (n_1555));
NAND2X1 g65281(.A (n_10678), .B (n_10667), .Y (n_2452));
NAND2X1 g65288(.A (g6513), .B (n_4322), .Y (n_1553));
AND2X1 g65296(.A (n_3030), .B (n_1550), .Y (n_2747));
OR4X1 g65301(.A (n_954), .B (g8785), .C (g8783), .D (g8784), .Y(n_1552));
NAND2X1 g65311(.A (g3470), .B (n_4320), .Y (n_1551));
AND2X1 g65312(.A (n_3030), .B (n_1554), .Y (n_3048));
AND2X1 g65315(.A (n_1550), .B (n_1549), .Y (n_3021));
AND2X1 g65318(.A (n_1631), .B (n_3025), .Y (n_2115));
AND2X1 g65321(.A (n_3025), .B (n_1549), .Y (n_2457));
OR2X1 g65323(.A (n_1559), .B (n_10499), .Y (n_1548));
NAND2X1 g65327(.A (g3821), .B (n_4314), .Y (n_1547));
AOI21X1 g65345(.A0 (n_442), .A1 (n_241), .B0 (n_9371), .Y (n_2677));
NAND3X1 g65358(.A (n_1313), .B (g4076), .C (n_245), .Y (n_1546));
NAND2X1 g65366(.A (g5821), .B (n_4327), .Y (n_1545));
NOR2X1 g65373(.A (n_956), .B (n_2111), .Y (n_1544));
AND2X1 g65375(.A (n_1536), .B (n_1543), .Y (n_6394));
NAND3X1 g65379(.A (n_1559), .B (n_1541), .C (n_1540), .Y (n_1542));
NAND2X1 g65380(.A (g3119), .B (n_4316), .Y (n_1539));
NOR2X1 g65381(.A (n_965), .B (n_1263), .Y (n_2113));
NAND3X1 g65383(.A (n_10499), .B (n_1538), .C (n_11221), .Y (n_2451));
NAND2X1 g65391(.A (n_1536), .B (n_6399), .Y (n_1537));
NAND2X1 g65402(.A (g5475), .B (n_4329), .Y (n_1535));
AOI22X1 g65406(.A0 (n_608), .A1 (n_1533), .B0 (n_1532), .B1 (n_1531),.Y (n_1534));
AOI22X1 g65407(.A0 (n_620), .A1 (n_1529), .B0 (n_1528), .B1 (n_1527),.Y (n_1530));
NAND3X1 g65412(.A (n_1488), .B (g5272), .C (g25114), .Y (n_11195));
AOI22X1 g65416(.A0 (n_675), .A1 (n_368), .B0 (n_450), .B1 (n_1524),.Y (n_1525));
AOI22X1 g65431(.A0 (n_611), .A1 (n_362), .B0 (n_380), .B1 (n_1522),.Y (n_1523));
AOI22X1 g65451(.A0 (n_1520), .A1 (n_1519), .B0 (n_1518), .B1(n_1517), .Y (n_1521));
AOI22X1 g65458(.A0 (n_1515), .A1 (n_278), .B0 (n_1514), .B1(n_10996), .Y (n_1516));
AOI22X1 g65489(.A0 (n_1510), .A1 (g25167), .B0 (n_1509), .B1(n_10616), .Y (n_1511));
AOI22X1 g65490(.A0 (n_1506), .A1 (n_213), .B0 (n_1505), .B1(n_10789), .Y (n_1507));
XOR2X1 g65505(.A (g1579), .B (n_1502), .Y (n_1503));
INVX2 g65507(.A (n_1845), .Y (n_2127));
INVX1 g65509(.A (n_1500), .Y (n_2119));
INVX1 g65513(.A (n_1848), .Y (n_2131));
INVX2 g65514(.A (n_1854), .Y (n_2143));
INVX1 g65517(.A (n_6806), .Y (n_2447));
INVX2 g65518(.A (n_8548), .Y (n_1499));
INVX2 g65526(.A (n_1494), .Y (n_2133));
INVX1 g65614(.A (n_1493), .Y (n_1662));
OR2X1 g65630(.A (n_581), .B (n_3849), .Y (n_2062));
NAND2X1 g65635(.A (n_745), .B (g7916), .Y (n_1491));
AND2X1 g65695(.A (n_1488), .B (g25114), .Y (n_2077));
NOR2X1 g65702(.A (n_807), .B (n_1486), .Y (n_1487));
NOR2X1 g65712(.A (n_744), .B (n_1482), .Y (n_1483));
NAND2X1 g65718(.A (n_1480), .B (n_1177), .Y (n_1481));
NOR2X1 g65720(.A (n_786), .B (g4049), .Y (n_1479));
NAND2X1 g65724(.A (n_1147), .B (n_1584), .Y (n_1478));
NAND2X1 g65726(.A (n_1476), .B (n_1222), .Y (n_1477));
NOR2X1 g65729(.A (n_814), .B (n_1482), .Y (n_1475));
NOR2X1 g65732(.A (n_11124), .B (g3698), .Y (n_1474));
NOR2X1 g65734(.A (n_794), .B (g3347), .Y (n_1473));
NAND2X1 g65735(.A (n_1158), .B (n_1471), .Y (n_1472));
NAND2X1 g65738(.A (n_1149), .B (n_1471), .Y (n_1470));
NOR2X1 g65740(.A (n_810), .B (n_1468), .Y (n_1469));
NOR2X1 g65741(.A (n_1468), .B (n_411), .Y (n_1467));
NAND2X1 g65744(.A (n_1412), .B (n_1476), .Y (n_1466));
NOR2X1 g65746(.A (n_718), .B (n_1464), .Y (n_1465));
NAND2X1 g65748(.A (n_1480), .B (n_1227), .Y (n_1463));
NAND2X1 g65752(.A (n_1734), .B (n_1267), .Y (n_1462));
AND2X1 g65757(.A (n_2432), .B (n_1461), .Y (n_2039));
NOR2X1 g65759(.A (n_739), .B (n_1459), .Y (n_1460));
NAND2X1 g65768(.A (n_1194), .B (n_1455), .Y (n_1456));
NAND2X1 g65771(.A (n_6399), .B (n_6398), .Y (n_1454));
NAND2X1 g65772(.A (n_1403), .B (n_1480), .Y (n_1453));
NAND2X1 g65774(.A (n_1455), .B (n_1145), .Y (n_1452));
NAND2X1 g65776(.A (n_1450), .B (n_1210), .Y (n_1451));
NAND2X1 g65780(.A (n_1207), .B (n_1450), .Y (n_1449));
NAND2X1 g65785(.A (n_1201), .B (n_1450), .Y (n_1448));
NAND2X1 g65790(.A (n_1450), .B (n_1199), .Y (n_1447));
NAND2X1 g65795(.A (n_1445), .B (n_1216), .Y (n_1446));
NAND2X1 g65801(.A (n_1442), .B (g1536), .Y (n_1444));
NOR2X1 g65802(.A (n_1442), .B (n_3849), .Y (n_1443));
NAND2X1 g65814(.A (n_1440), .B (n_1191), .Y (n_1441));
NAND2X1 g65820(.A (n_1185), .B (n_1440), .Y (n_1439));
NAND2X1 g65821(.A (n_1399), .B (n_1480), .Y (n_1438));
NAND2X1 g65826(.A (n_1455), .B (n_1169), .Y (n_1437));
NAND2X1 g65828(.A (n_1181), .B (n_1440), .Y (n_1436));
NAND2X1 g65831(.A (n_1440), .B (n_1175), .Y (n_1435));
INVX1 g65836(.A (n_1434), .Y (n_2067));
NAND2X1 g65842(.A (n_1471), .B (n_1143), .Y (n_1433));
NAND2X1 g65844(.A (n_1395), .B (n_1445), .Y (n_1432));
NAND2X1 g65852(.A (n_1246), .B (n_1455), .Y (n_1431));
NOR2X1 g65860(.A (n_748), .B (g4616), .Y (n_1429));
NOR2X1 g65863(.A (n_893), .B (n_1486), .Y (n_1428));
NAND2X1 g65869(.A (n_1584), .B (n_1135), .Y (n_1427));
NAND2X1 g65872(.A (n_772), .B (n_1173), .Y (n_1655));
AND2X1 g65873(.A (n_6406), .B (n_6398), .Y (n_6404));
NOR2X1 g65882(.A (g4737), .B (n_8776), .Y (n_1426));
NAND2X1 g62021(.A (g_18902), .B (n_4754), .Y (n_2345));
NAND2X1 g65894(.A (n_1476), .B (n_1234), .Y (n_1425));
NAND2X1 g65898(.A (n_1407), .B (n_1476), .Y (n_1424));
NOR2X1 g65905(.A (n_791), .B (n_1325), .Y (n_1423));
INVX1 g65910(.A (n_1422), .Y (n_4637));
NAND3X1 g65918(.A (n_11113), .B (n_719), .C (g_20951), .Y (n_1652));
NAND2X1 g65932(.A (n_1471), .B (n_1214), .Y (n_1419));
NAND2X1 g65933(.A (n_1584), .B (n_896), .Y (n_1418));
NOR2X1 g65937(.A (n_789), .B (n_659), .Y (n_1417));
NAND2X1 g65938(.A (n_1394), .B (n_1445), .Y (n_1416));
NAND2X1 g65940(.A (n_1445), .B (n_585), .Y (n_1415));
NAND2X1 g65942(.A (n_3812), .B (n_6406), .Y (n_1414));
NAND2X1 g65947(.A (n_1412), .B (n_1411), .Y (n_1413));
NAND2X1 g65950(.A (n_877), .B (n_6923), .Y (n_1409));
NAND2X1 g65952(.A (n_1407), .B (n_1411), .Y (n_1408));
NAND2X1 g65965(.A (n_1403), .B (n_1402), .Y (n_1404));
NAND2X1 g65967(.A (n_1403), .B (n_1762), .Y (n_1401));
NAND2X1 g65975(.A (n_1399), .B (n_1402), .Y (n_1400));
NAND2X1 g65978(.A (n_1399), .B (n_1762), .Y (n_1398));
NAND2X1 g65983(.A (n_1407), .B (n_1777), .Y (n_1397));
NAND2X1 g62041(.A (n_4757), .B (n_1599), .Y (n_1646));
OR2X1 g65991(.A (n_1395), .B (n_1394), .Y (n_1396));
NAND2X1 g65995(.A (n_1394), .B (n_1718), .Y (n_1393));
NAND2X1 g65996(.A (n_1394), .B (n_1391), .Y (n_1392));
AOI21X1 g66003(.A0 (g5188), .A1 (n_388), .B0 (n_1402), .Y (n_1390));
AOI21X1 g66009(.A0 (g5535), .A1 (n_383), .B0 (n_1411), .Y (n_1388));
AOI21X1 g66017(.A0 (g5881), .A1 (n_215), .B0 (n_1382), .Y (n_1384));
OAI21X1 g66018(.A0 (g17646), .A1 (g13068), .B0 (n_779), .Y (n_1381));
AOI21X1 g66021(.A0 (g6227), .A1 (n_330), .B0 (n_1377), .Y (n_1380));
AOI22X1 g66027(.A0 (n_10107), .A1 (n_723), .B0 (n_10108), .B1(n_552), .Y (n_10551));
AOI21X1 g66028(.A0 (g6573), .A1 (n_261), .B0 (n_1391), .Y (n_1375));
AOI21X1 g66030(.A0 (g3179), .A1 (n_370), .B0 (n_1370), .Y (n_1373));
AOI21X1 g66036(.A0 (g3530), .A1 (n_365), .B0 (n_1367), .Y (n_1369));
AOI21X1 g66046(.A0 (g3881), .A1 (n_303), .B0 (n_1364), .Y (n_1366));
AOI21X1 g66080(.A0 (n_6527), .A1 (n_3388), .B0 (n_3391), .Y (n_1363));
NAND4X1 g66086(.A (g17711), .B (g17580), .C (g12300), .D (g14694), .Y(n_2881));
NAND4X1 g66090(.A (g17778), .B (g17688), .C (g12470), .D (g14828), .Y(n_2871));
NAND4X1 g66095(.A (n_110), .B (g5046), .C (n_1356), .D (g5052), .Y(n_2044));
OAI21X1 g61479(.A0 (n_556), .A1 (g1333), .B0 (g12923), .Y (n_2060));
CLKBUFX1 gbuf_d_1090(.A(g16718), .Y(d_out_1090));
CLKBUFX1 gbuf_q_1090(.A(q_in_1090), .Y(g16603));
NAND2X1 g65420(.A (n_709), .B (n_1353), .Y (n_1354));
CLKBUFX1 gbuf_d_1091(.A(g16744), .Y(d_out_1091));
CLKBUFX1 gbuf_q_1091(.A(q_in_1091), .Y(g16627));
NAND2X1 g66596(.A (g1489), .B (n_9717), .Y (n_1628));
INVX1 g66633(.A (n_10214), .Y (n_1625));
AND2X1 g66661(.A (n_1352), .B (g8719), .Y (n_2001));
NAND3X1 g61513(.A (g19334), .B (n_325), .C (n_496), .Y (n_1351));
NOR2X1 g66878(.A (n_7260), .B (g4349), .Y (n_1349));
NAND2X1 g63875(.A (n_1331), .B (n_10119), .Y (n_2710));
OR2X1 g63876(.A (n_1331), .B (n_10119), .Y (n_1330));
INVX1 g63892(.A (n_1840), .Y (n_1329));
NAND2X1 g63894(.A (n_1328), .B (n_10112), .Y (n_2696));
OR2X1 g63896(.A (n_1328), .B (n_10112), .Y (n_1327));
NOR2X1 g65797(.A (n_1486), .B (n_1325), .Y (n_1326));
NAND2X1 g65962(.A (n_1412), .B (n_1777), .Y (n_1322));
INVX1 g66757(.A (n_1321), .Y (n_2019));
CLKBUFX1 gbuf_d_1092(.A(g12470), .Y(d_out_1092));
CLKBUFX1 gbuf_q_1092(.A(q_in_1092), .Y(g14828));
CLKBUFX1 gbuf_d_1093(.A(g12300), .Y(d_out_1093));
CLKBUFX1 gbuf_q_1093(.A(q_in_1093), .Y(g14694));
OR2X1 g61538(.A (n_470), .B (n_724), .Y (n_1315));
NAND3X1 g65343(.A (n_1313), .B (n_1312), .C (n_118), .Y (n_1737));
NOR2X1 g62659(.A (n_8585), .B (g3343), .Y (n_1311));
NOR2X1 g62660(.A (n_1272), .B (g3694), .Y (n_1310));
OR2X1 g64604(.A (n_980), .B (n_1307), .Y (n_1308));
NOR2X1 g65703(.A (n_1524), .B (n_433), .Y (n_1304));
AOI21X1 g64704(.A0 (n_1299), .A1 (g34028), .B0 (n_680), .Y (n_1300));
NAND2X1 g65897(.A (n_8796), .B (n_8591), .Y (n_1298));
XOR2X1 g64780(.A (n_1295), .B (n_982), .Y (n_1296));
NAND3X1 g64942(.A (n_663), .B (g1564), .C (g1554), .Y (n_2938));
NAND3X1 g64954(.A (n_971), .B (n_518), .C (n_8799), .Y (n_2945));
NAND3X1 g64966(.A (n_1093), .B (n_2443), .C (g5563), .Y (n_1293));
NAND3X1 g64968(.A (n_1011), .B (n_2432), .C (g6601), .Y (n_1292));
NOR2X1 g65279(.A (n_1290), .B (g_22379), .Y (n_1291));
CLKBUFX1 gbuf_d_1094(.A(g11418), .Y(d_out_1094));
CLKBUFX1 gbuf_q_1094(.A(q_in_1094), .Y(g13966));
NAND2X1 g66779(.A (n_1285), .B (n_11055), .Y (n_1286));
AOI21X1 g65228(.A0 (n_374), .A1 (n_4982), .B0 (g4749), .Y (n_1283));
AOI21X1 g65230(.A0 (n_339), .A1 (n_4978), .B0 (g4771), .Y (n_1282));
NAND2X1 g65320(.A (n_471), .B (n_1285), .Y (n_1279));
NAND2X1 g65352(.A (n_1820), .B (g8839), .Y (n_1278));
NOR2X1 g65370(.A (n_1276), .B (n_1275), .Y (n_1277));
NOR2X1 g65397(.A (g4878), .B (n_1274), .Y (n_1826));
INVX1 g66421(.A (n_1272), .Y (n_1273));
AOI21X1 g65445(.A0 (g34026), .A1 (g21245), .B0 (n_676), .Y (n_1271));
NAND2X1 g66414(.A (n_596), .B (n_10013), .Y (n_5378));
XOR2X1 g66025(.A (g6159), .B (n_3589), .Y (n_1269));
CLKBUFX1 gbuf_d_1095(.A(g17819), .Y(d_out_1095));
CLKBUFX1 gbuf_q_1095(.A(q_in_1095), .Y(g14673));
CLKBUFX1 gbuf_d_1096(.A(g17871), .Y(d_out_1096));
CLKBUFX1 gbuf_q_1096(.A(q_in_1096), .Y(g14749));
CLKBUFX1 gbuf_d_1097(.A(g4474), .Y(d_out_1097));
CLKBUFX1 gbuf_q_1097(.A(q_in_1097), .Y(g4477));
NAND2X1 g65615(.A (n_771), .B (g5029), .Y (n_1493));
NAND2X1 g65616(.A (n_1267), .B (n_3624), .Y (n_1268));
NOR2X1 g65617(.A (n_578), .B (g5511), .Y (n_1772));
INVX1 g65618(.A (n_1554), .Y (n_1266));
NAND2X1 g65625(.A (n_1264), .B (n_1214), .Y (n_4324));
NOR2X1 g65626(.A (n_566), .B (g6203), .Y (n_1770));
INVX1 g65633(.A (n_1263), .Y (n_2153));
INVX1 g65636(.A (n_3025), .Y (n_1262));
NOR2X1 g65639(.A (n_580), .B (g3506), .Y (n_1752));
NAND2X1 g65640(.A (g1950), .B (n_579), .Y (n_1261));
NAND2X1 g65642(.A (g1816), .B (n_557), .Y (n_1260));
NAND2X1 g65647(.A (g2084), .B (n_558), .Y (n_1257));
NAND2X1 g65649(.A (n_10724), .B (g7916), .Y (n_1255));
NOR2X1 g65651(.A (n_575), .B (g3857), .Y (n_1744));
INVX1 g65655(.A (n_1812), .Y (g26801));
INVX1 g65666(.A (n_1252), .Y (n_4628));
NOR2X1 g65669(.A (n_587), .B (g6549), .Y (n_1765));
NAND2X1 g65670(.A (n_594), .B (n_662), .Y (n_1251));
NOR2X1 g65674(.A (n_479), .B (g5164), .Y (n_1763));
INVX1 g65675(.A (n_1550), .Y (n_1250));
NOR2X1 g65681(.A (n_565), .B (g3155), .Y (n_1767));
NAND2X1 g65694(.A (n_653), .B (n_8677), .Y (n_1576));
NOR2X1 g65696(.A (n_1531), .B (n_187), .Y (n_1248));
AND2X1 g65697(.A (n_1246), .B (n_1245), .Y (n_1247));
AND2X1 g65709(.A (n_1243), .B (n_1242), .Y (n_1244));
NAND3X1 g65714(.A (g2130), .B (n_1240), .C (g2145), .Y (n_1241));
NOR2X1 g65719(.A (n_673), .B (n_1154), .Y (n_1239));
INVX1 g65722(.A (n_4617), .Y (n_1238));
NAND2X1 g65730(.A (n_1236), .B (n_827), .Y (n_1237));
NAND2X1 g65731(.A (n_1411), .B (n_1234), .Y (n_1235));
NOR2X1 g65742(.A (n_1464), .B (n_1224), .Y (n_1232));
NAND2X1 g65743(.A (n_1230), .B (n_836), .Y (n_1231));
AND2X1 g65751(.A (n_1762), .B (n_1227), .Y (n_1228));
NAND3X1 g65753(.A (n_269), .B (n_812), .C (g2453), .Y (n_1226));
NOR2X1 g65754(.A (n_822), .B (n_1224), .Y (n_1225));
AND2X1 g65756(.A (n_1411), .B (n_1222), .Y (n_1223));
NOR2X1 g65758(.A (n_3391), .B (n_3388), .Y (n_1221));
INVX1 g65761(.A (n_1219), .Y (n_1220));
NAND2X1 g65767(.A (n_1718), .B (n_1216), .Y (n_1217));
NAND2X1 g65770(.A (n_1723), .B (n_1214), .Y (n_1215));
NOR2X1 g65777(.A (n_1212), .B (n_3812), .Y (n_1213));
NAND2X1 g65778(.A (n_1751), .B (n_1210), .Y (n_1211));
NAND2X1 g65779(.A (n_1367), .B (n_1210), .Y (n_1209));
AND2X1 g65782(.A (n_1207), .B (n_1206), .Y (n_1208));
NOR2X1 g65783(.A (n_817), .B (n_1224), .Y (n_1205));
AND2X1 g65788(.A (n_1201), .B (n_1206), .Y (n_1202));
AND2X1 g65791(.A (n_1751), .B (n_1199), .Y (n_1200));
AND2X1 g65792(.A (n_1367), .B (n_1199), .Y (n_1198));
AND2X1 g65808(.A (n_1194), .B (n_1245), .Y (n_1195));
NAND3X1 g65812(.A (n_291), .B (n_806), .C (g1894), .Y (n_1193));
NAND2X1 g65816(.A (n_1743), .B (n_1191), .Y (n_1192));
NAND2X1 g65818(.A (n_1364), .B (n_1191), .Y (n_1189));
AND2X1 g65819(.A (n_8832), .B (g7916), .Y (n_1188));
AND2X1 g65824(.A (n_1777), .B (n_1222), .Y (n_1187));
AND2X1 g65825(.A (n_1185), .B (n_1184), .Y (n_1186));
NAND2X1 g65827(.A (n_1024), .B (n_10563), .Y (n_1183));
AND2X1 g65829(.A (n_1181), .B (n_1184), .Y (n_1182));
NAND2X1 g65830(.A (n_1179), .B (n_1165), .Y (n_1180));
NAND2X1 g65833(.A (n_1402), .B (n_1177), .Y (n_1178));
AND2X1 g65834(.A (n_1743), .B (n_1175), .Y (n_1176));
NAND2X1 g65837(.A (n_644), .B (n_11209), .Y (n_1434));
AND2X1 g65839(.A (n_1364), .B (n_1175), .Y (n_1174));
OR2X1 g65840(.A (n_1173), .B (g5029), .Y (n_7010));
NAND2X1 g65856(.A (n_1725), .B (n_1169), .Y (n_1170));
NOR2X1 g65858(.A (n_1527), .B (n_382), .Y (n_1168));
NAND2X1 g65859(.A (n_1391), .B (n_1216), .Y (n_1167));
NAND2X1 g65864(.A (n_978), .B (n_1165), .Y (n_1166));
NAND2X1 g65870(.A (n_1762), .B (n_1177), .Y (n_1164));
NAND2X1 g65875(.A (g_7220), .B (g8291), .Y (n_1731));
NAND3X1 g65880(.A (n_444), .B (n_804), .C (g1760), .Y (n_1163));
NAND3X1 g65881(.A (n_377), .B (n_730), .C (g2319), .Y (n_1162));
NAND2X1 g65885(.A (n_1160), .B (n_831), .Y (n_1161));
AND2X1 g65886(.A (n_1158), .B (n_1264), .Y (n_1159));
NOR2X1 g65892(.A (n_795), .B (n_1154), .Y (n_1155));
NAND2X1 g65893(.A (n_1377), .B (n_1214), .Y (n_1153));
AND2X1 g65902(.A (n_1395), .B (n_590), .Y (n_1152));
AND2X1 g65903(.A (n_1149), .B (n_1264), .Y (n_1150));
AND2X1 g65904(.A (n_1147), .B (n_1242), .Y (n_1148));
AND2X1 g65906(.A (n_1382), .B (n_1145), .Y (n_1146));
AND2X1 g65907(.A (n_1377), .B (n_1143), .Y (n_1144));
NAND2X1 g65911(.A (n_1179), .B (g13272), .Y (n_1422));
NAND2X1 g65925(.A (n_1138), .B (n_839), .Y (n_1139));
NAND2X1 g65926(.A (g5913), .B (n_10508), .Y (n_1137));
INVX1 g65929(.A (n_1536), .Y (n_6402));
NAND2X1 g65931(.A (n_1370), .B (n_1135), .Y (n_1136));
NAND3X1 g65945(.A (g2130), .B (g2138), .C (g2145), .Y (n_1133));
NAND2X1 g65946(.A (n_1777), .B (n_1234), .Y (n_1131));
NAND2X1 g65949(.A (n_1181), .B (n_1743), .Y (n_1130));
NAND2X1 g65955(.A (n_1158), .B (n_1723), .Y (n_1128));
NAND2X1 g65956(.A (n_1149), .B (n_1723), .Y (n_1127));
INVX1 g65958(.A (n_1124), .Y (n_1405));
NAND2X1 g65960(.A (n_1147), .B (n_1370), .Y (n_1123));
NAND2X1 g65963(.A (n_1395), .B (n_1718), .Y (n_1122));
NAND2X1 g65966(.A (n_1147), .B (n_1758), .Y (n_1121));
NAND2X1 g65968(.A (n_1246), .B (n_1725), .Y (n_1120));
NAND2X1 g65971(.A (n_1207), .B (n_1751), .Y (n_1119));
NAND2X1 g65972(.A (n_1207), .B (n_1367), .Y (n_1118));
NAND2X1 g65973(.A (n_1201), .B (n_1751), .Y (n_1117));
NAND2X1 g65974(.A (n_1201), .B (n_1367), .Y (n_1116));
OR2X1 g65976(.A (n_1207), .B (n_1201), .Y (n_1115));
NAND2X1 g65977(.A (n_1194), .B (n_1382), .Y (n_1114));
OR2X1 g65979(.A (n_1185), .B (n_1181), .Y (n_1113));
NAND2X1 g65980(.A (n_1185), .B (n_1743), .Y (n_1112));
NAND2X1 g65981(.A (n_1185), .B (n_1364), .Y (n_1111));
NAND2X1 g65982(.A (n_1181), .B (n_1364), .Y (n_1110));
OR2X1 g65985(.A (n_1243), .B (n_1147), .Y (n_1109));
NAND2X1 g65988(.A (n_1194), .B (n_1725), .Y (n_1108));
NAND2X1 g65989(.A (n_1158), .B (n_1377), .Y (n_1107));
NAND2X1 g65990(.A (n_1149), .B (n_1377), .Y (n_1106));
NAND2X1 g65993(.A (n_1243), .B (n_1370), .Y (n_1105));
NAND2X1 g65997(.A (n_1246), .B (n_1382), .Y (n_1104));
NAND2X1 g65998(.A (n_1395), .B (n_1391), .Y (n_1103));
NAND2X1 g65999(.A (n_1243), .B (n_1758), .Y (n_1102));
XOR2X1 g66000(.A (g5120), .B (n_3618), .Y (n_1101));
OAI21X1 g66014(.A0 (n_423), .A1 (n_11050), .B0 (n_1100), .Y (n_1845));
XOR2X1 g66031(.A (g6505), .B (n_3604), .Y (n_1099));
XOR2X1 g66032(.A (g5813), .B (n_3611), .Y (n_1098));
OAI21X1 g66037(.A0 (n_11160), .A1 (g_6165), .B0 (n_818), .Y (n_1848));
XOR2X1 g66052(.A (g5467), .B (n_3616), .Y (n_1097));
OAI21X1 g66058(.A0 (n_10369), .A1 (g_4409), .B0 (n_823), .Y (n_1854));
AOI21X1 g66060(.A0 (n_512), .A1 (g4601), .B0 (n_820), .Y (n_1096));
XOR2X1 g66069(.A (n_364), .B (g_22552), .Y (n_1095));
NAND2X1 g66732(.A (g17577), .B (g17519), .Y (n_1094));
AOI21X1 g66075(.A0 (n_776), .A1 (n_409), .B0 (n_1093), .Y (n_1494));
NAND4X1 g66085(.A (g17674), .B (g17519), .C (g12238), .D (g14662), .Y(n_3171));
NAND4X1 g66087(.A (g_15380), .B (g_15381), .C (n_413), .D (g_16792),.Y (n_1090));
NAND4X1 g66093(.A (g17760), .B (g17649), .C (g12422), .D (g14779), .Y(n_2729));
NAND4X1 g66094(.A (g17739), .B (g17607), .C (g12350), .D (g14738), .Y(n_2732));
NOR2X1 g65622(.A (n_589), .B (g5857), .Y (n_1727));
MX2X1 g66151(.A (n_527), .B (g14662), .S0 (g17674), .Y (n_1085));
MX2X1 g66152(.A (n_669), .B (g14694), .S0 (g17711), .Y (n_1084));
MX2X1 g66153(.A (n_549), .B (g14779), .S0 (g17760), .Y (n_1083));
MX2X1 g66155(.A (n_538), .B (g14828), .S0 (g17778), .Y (n_1082));
MX2X1 g66157(.A (g_22552), .B (n_364), .S0 (g_16404), .Y (n_1081));
XOR2X1 g66160(.A (g5527), .B (n_1234), .Y (n_1079));
XOR2X1 g66161(.A (g5180), .B (n_1177), .Y (n_1077));
XOR2X1 g66168(.A (g3171), .B (n_1135), .Y (n_1075));
XOR2X1 g66169(.A (g3522), .B (n_1210), .Y (n_1074));
XOR2X1 g66172(.A (g6219), .B (n_1214), .Y (n_1072));
XOR2X1 g66181(.A (g6565), .B (n_1216), .Y (n_1071));
XOR2X1 g66188(.A (g5873), .B (n_1169), .Y (n_1069));
CLKBUFX1 gbuf_d_1098(.A(g17787), .Y(d_out_1098));
CLKBUFX1 gbuf_q_1098(.A(q_in_1098), .Y(g14597));
CLKBUFX1 gbuf_d_1099(.A(g13966), .Y(d_out_1099));
CLKBUFX1 gbuf_q_1099(.A(q_in_1099), .Y(g16775));
INVX1 g66355(.A (n_1064), .Y (n_1065));
INVX1 g66390(.A (n_1062), .Y (n_1063));
INVX1 g66559(.A (n_1059), .Y (n_1060));
INVX1 g66566(.A (n_2339), .Y (n_1058));
INVX1 g66607(.A (n_1055), .Y (n_4878));
NAND2X1 g66642(.A (g17604), .B (g17580), .Y (n_1054));
NOR2X1 g66693(.A (n_5917), .B (g2351), .Y (n_1053));
NOR2X1 g66743(.A (n_5921), .B (g2485), .Y (n_1052));
NAND2X1 g66758(.A (g3466), .B (n_10950), .Y (n_1321));
CLKBUFX1 gbuf_d_1100(.A(g17845), .Y(d_out_1100));
CLKBUFX1 gbuf_q_1100(.A(q_in_1100), .Y(g14705));
NAND2X1 g66799(.A (g17685), .B (g17649), .Y (n_1046));
NOR2X1 g66843(.A (n_5925), .B (g1926), .Y (n_1044));
INVX1 g66846(.A (n_3459), .Y (n_1043));
NOR2X1 g66904(.A (n_5996), .B (g1792), .Y (n_1040));
CLKBUFX1 gbuf_d_1101(.A(g17813), .Y(d_out_1101));
CLKBUFX1 gbuf_q_1101(.A(q_in_1101), .Y(g14635));
INVX2 g67909(.A (n_5402), .Y (n_3894));
INVX1 g62237(.A (n_4754), .Y (n_2878));
AND2X1 g62259(.A (n_8591), .B (g13259), .Y (n_4764));
AND2X1 g62262(.A (n_8832), .B (g13259), .Y (n_4761));
OR2X1 g65994(.A (n_10567), .B (n_1024), .Y (n_10550));
NAND2X1 g66590(.A (g17722), .B (g17688), .Y (n_1021));
OR2X1 g65992(.A (n_1158), .B (n_1149), .Y (n_1017));
AND2X1 g65396(.A (g4878), .B (n_1274), .Y (n_1016));
NOR2X1 g61630(.A (g4434), .B (n_596), .Y (n_1015));
AND2X1 g63893(.A (n_1307), .B (g4659), .Y (n_1840));
NOR2X1 g65733(.A (n_1522), .B (n_418), .Y (n_1014));
OR2X1 g65389(.A (n_989), .B (n_10499), .Y (n_1013));
AOI21X1 g66081(.A0 (n_11185), .A1 (n_322), .B0 (n_1011), .Y (n_1500));
CLKBUFX1 gbuf_d_1102(.A(g17580), .Y(d_out_1102));
CLKBUFX1 gbuf_q_1102(.A(q_in_1102), .Y(g17604));
CLKBUFX1 gbuf_d_1103(.A(g12238), .Y(d_out_1103));
CLKBUFX1 gbuf_q_1103(.A(q_in_1103), .Y(g14662));
CLKBUFX1 gbuf_d_1104(.A(g34034), .Y(d_out_1104));
CLKBUFX1 gbuf_q_1104(.A(q_in_1104), .Y(g34035));
CLKBUFX1 gbuf_d_1105(.A(g12422), .Y(d_out_1105));
CLKBUFX1 gbuf_q_1105(.A(q_in_1105), .Y(g14779));
CLKBUFX1 gbuf_d_1106(.A(g17688), .Y(d_out_1106));
CLKBUFX1 gbuf_q_1106(.A(q_in_1106), .Y(g17722));
CLKBUFX1 gbuf_d_1107(.A(g12350), .Y(d_out_1107));
CLKBUFX1 gbuf_q_1107(.A(q_in_1107), .Y(g14738));
CLKBUFX1 gbuf_d_1108(.A(g11388), .Y(d_out_1108));
CLKBUFX1 gbuf_q_1108(.A(q_in_1108), .Y(g13926));
CLKBUFX1 gbuf_d_1109(.A(g11349), .Y(d_out_1109));
CLKBUFX1 gbuf_q_1109(.A(q_in_1109), .Y(g13895));
CLKBUFX1 gbuf_d_1110(.A(g17649), .Y(d_out_1110));
CLKBUFX1 gbuf_q_1110(.A(q_in_1110), .Y(g17685));
OR2X1 g65954(.A (n_1194), .B (n_1246), .Y (n_1002));
CLKBUFX1 gbuf_d_1111(.A(g17519), .Y(d_out_1111));
CLKBUFX1 gbuf_q_1111(.A(q_in_1111), .Y(g17577));
NAND2X1 g65765(.A (n_1382), .B (n_1169), .Y (n_999));
XOR2X1 g66174(.A (g3873), .B (n_1191), .Y (n_998));
NOR2X1 g65736(.A (n_983), .B (n_1154), .Y (n_995));
NOR2X1 g65372(.A (n_151), .B (g4878), .Y (n_994));
NAND2X1 g65745(.A (n_1758), .B (n_1135), .Y (n_993));
OR2X1 g65721(.A (g_9174), .B (g2980), .Y (n_992));
NOR2X1 g65329(.A (n_6707), .B (n_989), .Y (n_991));
NAND4X1 g64601(.A (n_988), .B (n_987), .C (n_986), .D (g4688), .Y(n_4839));
INVX2 g68008(.A (g25219), .Y (n_1695));
INVX1 g66416(.A (n_983), .Y (n_1412));
NOR2X1 g64840(.A (n_474), .B (n_307), .Y (n_1331));
NOR2X1 g64849(.A (n_982), .B (n_1295), .Y (n_1328));
NOR3X1 g64899(.A (g_16404), .B (g_22552), .C (n_364), .Y (n_5582));
XOR2X1 g66061(.A (n_2485), .B (g1472), .Y (n_981));
NOR2X1 g64914(.A (n_69), .B (g4653), .Y (n_980));
INVX1 g66447(.A (n_978), .Y (n_1442));
NOR2X1 g66793(.A (g3171), .B (g3179), .Y (n_1584));
OAI21X1 g65677(.A0 (g3480), .A1 (g3494), .B0 (n_10949), .Y (n_1550));
XOR2X1 g66034(.A (n_1799), .B (n_2699), .Y (n_977));
OAI21X1 g65683(.A0 (g5485), .A1 (g5499), .B0 (n_8921), .Y (n_1631));
XOR2X1 g66033(.A (n_975), .B (n_6025), .Y (n_976));
OR2X1 g65679(.A (n_948), .B (g4628), .Y (n_974));
CLKBUFX1 gbuf_d_1112(.A(g34026), .Y(d_out_1112));
CLKBUFX1 gbuf_q_1112(.A(q_in_1112), .Y(g34027));
CLKBUFX1 gbuf_d_1113(.A(g34027), .Y(d_out_1113));
CLKBUFX1 gbuf_q_1113(.A(q_in_1113), .Y(g34028));
NAND2X1 g65667(.A (n_908), .B (g13272), .Y (n_1252));
NAND2X1 g65653(.A (n_973), .B (n_1234), .Y (n_4329));
NAND2X1 g65657(.A (n_970), .B (n_1177), .Y (n_1812));
XOR2X1 g66026(.A (g1300), .B (n_3383), .Y (n_969));
NAND3X1 g65861(.A (n_196), .B (n_6967), .C (g5057), .Y (n_2045));
NAND2X1 g65621(.A (n_1245), .B (n_1169), .Y (n_4327));
OR2X1 g65623(.A (g2509), .B (n_8632), .Y (n_967));
INVX1 g65627(.A (n_1630), .Y (n_965));
OR2X1 g65631(.A (g2375), .B (n_8627), .Y (n_963));
NOR2X1 g65634(.A (n_343), .B (n_9297), .Y (n_1263));
NAND2X1 g65638(.A (n_1206), .B (n_1210), .Y (n_4320));
OR2X1 g65646(.A (n_309), .B (g17423), .Y (n_961));
NOR2X1 g65654(.A (n_429), .B (g2357), .Y (n_958));
OR2X1 g65660(.A (n_295), .B (g17400), .Y (n_957));
NAND2X1 g65661(.A (n_1312), .B (n_955), .Y (n_956));
NAND2X1 g65662(.A (n_1242), .B (n_1135), .Y (n_4316));
OR2X1 g65663(.A (n_220), .B (n_10871), .Y (n_954));
OAI21X1 g65664(.A0 (g3129), .A1 (g3143), .B0 (g35), .Y (n_3030));
OR2X1 g65668(.A (g2241), .B (n_8534), .Y (n_952));
AND2X1 g65671(.A (n_188), .B (n_955), .Y (n_1313));
NAND2X1 g65672(.A (n_590), .B (n_1216), .Y (n_4322));
OAI21X1 g65673(.A0 (g3831), .A1 (g3845), .B0 (n_10949), .Y (n_1549));
NOR2X1 g65678(.A (n_302), .B (g2112), .Y (n_950));
NAND2X1 g65680(.A (n_948), .B (g4628), .Y (n_2980));
NOR2X1 g65682(.A (n_436), .B (g2671), .Y (n_947));
INVX1 g68403(.A (n_946), .Y (n_3707));
NOR2X1 g65684(.A (n_298), .B (g1798), .Y (n_943));
OR2X1 g65685(.A (g2643), .B (n_10720), .Y (n_942));
OR2X1 g65686(.A (g1682), .B (n_10271), .Y (n_940));
AND2X1 g65723(.A (n_899), .B (g13272), .Y (n_4617));
NAND2X1 g65725(.A (n_323), .B (n_2550), .Y (n_938));
XOR2X1 g66038(.A (g3111), .B (n_3609), .Y (n_937));
NAND2X1 g65775(.A (n_336), .B (n_933), .Y (n_934));
NAND2X1 g65789(.A (n_441), .B (n_2306), .Y (n_932));
AND2X1 g65793(.A (n_1199), .B (n_1206), .Y (n_931));
NAND3X1 g65805(.A (n_928), .B (g1624), .C (n_677), .Y (n_929));
NAND2X1 g65807(.A (n_240), .B (n_926), .Y (n_927));
NAND3X1 g65809(.A (n_399), .B (n_674), .C (g2028), .Y (n_925));
NOR3X1 g65822(.A (g_21778), .B (n_273), .C (g_19113), .Y (n_924));
OR4X1 g65832(.A (n_10113), .B (g1564), .C (g1554), .D (g1548), .Y(n_2108));
OR2X1 g66729(.A (g8416), .B (g7916), .Y (n_923));
AND2X1 g65841(.A (n_1175), .B (n_1184), .Y (n_921));
NOR2X1 g65850(.A (n_218), .B (n_143), .Y (n_10905));
NAND3X1 g65854(.A (n_919), .B (n_619), .C (g2185), .Y (n_920));
OR4X1 g65855(.A (g2657), .B (g2523), .C (g2255), .D (g2389), .Y(n_918));
AND2X1 g65857(.A (n_916), .B (n_8534), .Y (n_917));
NAND2X1 g65862(.A (n_376), .B (n_2293), .Y (n_915));
NAND2X1 g65877(.A (g1950), .B (n_6790), .Y (n_914));
AND2X1 g65883(.A (n_911), .B (n_8627), .Y (n_912));
AND2X1 g65884(.A (n_6399), .B (n_3641), .Y (n_1543));
AND2X1 g65888(.A (n_1145), .B (n_1245), .Y (n_910));
NAND2X1 g65899(.A (n_908), .B (n_1165), .Y (n_909));
NAND2X1 g65912(.A (n_408), .B (n_2780), .Y (n_906));
AND2X1 g65924(.A (n_904), .B (n_8632), .Y (n_905));
AND2X1 g65927(.A (n_902), .B (n_10720), .Y (n_903));
NOR2X1 g65930(.A (n_901), .B (n_3812), .Y (n_1536));
NAND2X1 g65935(.A (n_1165), .B (n_899), .Y (n_900));
NAND3X1 g65939(.A (g2130), .B (g2138), .C (n_308), .Y (n_898));
AND2X1 g65941(.A (n_896), .B (n_1242), .Y (n_897));
NAND3X1 g65943(.A (n_351), .B (n_610), .C (g2587), .Y (n_895));
NAND2X1 g65944(.A (n_338), .B (n_2521), .Y (n_894));
INVX1 g66380(.A (n_1718), .Y (n_893));
AOI21X1 g65987(.A0 (g_20073), .A1 (g_12433), .B0 (n_891), .Y(n_10552));
XOR2X1 g66002(.A (n_1813), .B (n_2718), .Y (n_890));
XOR2X1 g66006(.A (n_1794), .B (n_3007), .Y (n_888));
XOR2X1 g66008(.A (n_1810), .B (n_3011), .Y (n_887));
XOR2X1 g66011(.A (n_885), .B (n_5975), .Y (n_886));
XOR2X1 g66012(.A (n_883), .B (n_5978), .Y (n_884));
XOR2X1 g66016(.A (n_1807), .B (n_2684), .Y (n_882));
XOR2X1 g66020(.A (n_2084), .B (n_2704), .Y (n_881));
XOR2X1 g66022(.A (n_1805), .B (n_2686), .Y (n_880));
INVX1 g66451(.A (n_876), .Y (n_877));
AND2X1 g66737(.A (n_11177), .B (g17722), .Y (n_1461));
XOR2X1 g66035(.A (n_871), .B (n_4946), .Y (n_872));
OAI21X1 g65637(.A0 (g5138), .A1 (g5152), .B0 (n_10949), .Y (n_3025));
XOR2X1 g66043(.A (g3813), .B (n_3596), .Y (n_868));
XOR2X1 g66045(.A (n_866), .B (n_5972), .Y (n_867));
XOR2X1 g66047(.A (n_864), .B (n_5961), .Y (n_8755));
XOR2X1 g66048(.A (n_862), .B (n_5953), .Y (n_863));
XOR2X1 g66049(.A (n_860), .B (n_6017), .Y (n_861));
XOR2X1 g66050(.A (n_858), .B (n_5969), .Y (n_859));
XOR2X1 g66051(.A (n_856), .B (n_5964), .Y (n_857));
XOR2X1 g66054(.A (n_854), .B (n_4948), .Y (n_855));
XOR2X1 g66055(.A (n_852), .B (n_6020), .Y (n_10554));
XOR2X1 g66059(.A (n_2556), .B (g_16456), .Y (n_851));
XOR2X1 g66062(.A (n_2535), .B (g1478), .Y (n_849));
XOR2X1 g66070(.A (n_2529), .B (g_11413), .Y (n_848));
XOR2X1 g66072(.A (n_846), .B (n_4942), .Y (n_847));
XOR2X1 g66082(.A (g3462), .B (n_3601), .Y (n_845));
OAI21X1 g65620(.A0 (g5831), .A1 (g5845), .B0 (n_8921), .Y (n_1554));
NAND4X1 g66091(.A (g4489), .B (g4483), .C (g4492), .D (g4486), .Y(n_1562));
AOI22X1 g66092(.A0 (g3333), .A1 (g34035), .B0 (n_843), .B1 (g34034),.Y (n_844));
MX2X1 g66156(.A (n_371), .B (g14738), .S0 (g17739), .Y (n_842));
XOR2X1 g66158(.A (g1691), .B (n_4527), .Y (n_841));
XOR2X1 g66159(.A (n_4531), .B (n_839), .Y (n_840));
XOR2X1 g66163(.A (n_1796), .B (n_2692), .Y (n_838));
XOR2X1 g66166(.A (n_4187), .B (n_836), .Y (n_837));
XOR2X1 g66170(.A (g1448), .B (n_2538), .Y (n_835));
XOR2X1 g66171(.A (g2093), .B (n_4183), .Y (n_834));
XOR2X1 g66177(.A (g2250), .B (n_4906), .Y (n_833));
XOR2X1 g66178(.A (n_4529), .B (n_831), .Y (n_832));
XOR2X1 g66180(.A (g_18869), .B (n_2244), .Y (n_830));
XOR2X1 g66183(.A (g2652), .B (n_4726), .Y (n_829));
XOR2X1 g66184(.A (n_4190), .B (n_827), .Y (n_828));
CLKBUFX1 g66185(.A (n_6707), .Y (n_1559));
INVX1 g66208(.A (g_7220), .Y (n_826));
CLKBUFX1 gbuf_d_1114(.A(g13895), .Y(d_out_1114));
CLKBUFX1 gbuf_q_1114(.A(q_in_1114), .Y(g16718));
INVX1 g66284(.A (n_823), .Y (n_824));
INVX1 g66300(.A (n_822), .Y (n_1403));
INVX1 g66303(.A (n_820), .Y (n_821));
INVX1 g66312(.A (n_818), .Y (n_819));
INVX1 g66332(.A (n_817), .Y (n_1399));
INVX1 g66703(.A (n_6552), .Y (n_816));
INVX1 g66342(.A (n_1758), .Y (n_814));
NOR2X1 g66356(.A (n_812), .B (g2485), .Y (n_1064));
INVX1 g66370(.A (n_1723), .Y (n_810));
INVX1 g66377(.A (n_1138), .Y (n_808));
INVX1 g66386(.A (n_1391), .Y (n_807));
NOR2X1 g66391(.A (n_806), .B (g1926), .Y (n_1062));
AND2X1 g66392(.A (n_804), .B (g1792), .Y (n_805));
INVX1 g66422(.A (n_4682), .Y (n_1272));
INVX1 g66434(.A (n_802), .Y (n_803));
INVX1 g66454(.A (n_800), .Y (n_801));
NOR2X1 g66483(.A (n_804), .B (g1792), .Y (n_1667));
INVX1 g66485(.A (n_799), .Y (n_1599));
INVX1 g66489(.A (n_1236), .Y (n_798));
NOR2X1 g66492(.A (n_448), .B (n_662), .Y (n_797));
INVX1 g66505(.A (n_795), .Y (n_1407));
INVX1 g66516(.A (n_8572), .Y (n_794));
INVX1 g66520(.A (n_1160), .Y (n_793));
INVX1 g66535(.A (n_791), .Y (n_1394));
AND2X1 g66548(.A (n_812), .B (g2485), .Y (n_790));
INVX1 g66550(.A (n_3391), .Y (n_789));
INVX1 g66578(.A (n_6808), .Y (n_786));
NOR2X1 g66598(.A (g6565), .B (g6573), .Y (n_1445));
NOR2X1 g66599(.A (g4349), .B (n_1627), .Y (n_1734));
NAND2X1 g66608(.A (g3817), .B (n_10949), .Y (n_1055));
INVX1 g66613(.A (n_590), .Y (n_1325));
NAND2X1 g66618(.A (g4401), .B (g4392), .Y (n_784));
NOR2X1 g66619(.A (g1636), .B (n_4120), .Y (n_783));
NOR2X1 g66622(.A (g3522), .B (g3530), .Y (n_1450));
NOR2X1 g66625(.A (n_5928), .B (g2619), .Y (n_782));
OR2X1 g66639(.A (n_6967), .B (n_1356), .Y (n_2679));
AND2X1 g66649(.A (n_424), .B (g17646), .Y (n_1458));
NAND2X1 g66654(.A (g5817), .B (n_10950), .Y (n_6398));
NOR2X1 g66659(.A (g3873), .B (g3881), .Y (n_1440));
NOR2X1 g66663(.A (g6219), .B (g6227), .Y (n_1471));
NAND2X1 g66674(.A (n_3439), .B (n_659), .Y (n_780));
NAND2X1 g66682(.A (g17646), .B (g17607), .Y (n_779));
INVX1 g66353(.A (n_1230), .Y (n_778));
INVX1 g66711(.A (n_1538), .Y (n_777));
AND2X1 g66736(.A (n_776), .B (g17604), .Y (n_1484));
NOR2X1 g66759(.A (n_5941), .B (g2217), .Y (n_775));
INVX1 g66774(.A (n_771), .Y (n_772));
NOR2X1 g66784(.A (g1657), .B (n_5936), .Y (n_769));
INVX1 g66458(.A (n_10578), .Y (n_11217));
CLKBUFX1 gbuf_d_1115(.A(g34028), .Y(d_out_1115));
CLKBUFX1 gbuf_qn_1115(.A(qn_in_1115), .Y(g4688));
NOR2X1 g66851(.A (n_10213), .B (n_11129), .Y (n_10206));
NOR2X1 g66867(.A (n_5932), .B (g2060), .Y (n_765));
AND2X1 g66870(.A (g25219), .B (g17577), .Y (n_1488));
NAND2X1 g66891(.A (g6163), .B (n_10949), .Y (n_6406));
NOR2X1 g66720(.A (g5873), .B (g5881), .Y (n_1455));
AND2X1 g66660(.A (n_11157), .B (g17685), .Y (n_1457));
INVX1 g66315(.A (n_747), .Y (n_748));
AND2X1 g62238(.A (n_746), .B (g13259), .Y (n_4754));
AND2X1 g62244(.A (n_745), .B (g13259), .Y (n_4757));
INVX1 g66292(.A (n_1370), .Y (n_744));
INVX1 g68093(.A (n_740), .Y (n_741));
INVX1 g66479(.A (n_1725), .Y (n_739));
NOR2X1 g66560(.A (n_730), .B (g2351), .Y (n_1059));
INVX2 g67032(.A (n_2421), .Y (n_2376));
CLKBUFX1 gbuf_d_1116(.A(g13926), .Y(d_out_1116));
CLKBUFX1 gbuf_q_1116(.A(q_in_1116), .Y(g16744));
OAI21X1 g61595(.A0 (g4401), .A1 (g4434), .B0 (n_243), .Y (n_724));
INVX1 g66918(.A (n_723), .Y (n_3042));
XOR2X1 g66077(.A (n_2280), .B (g_20563), .Y (n_722));
CLKBUFX1 gbuf_d_1117(.A(g17607), .Y(d_out_1117));
CLKBUFX1 gbuf_q_1117(.A(q_in_1117), .Y(g17646));
AOI21X1 g65984(.A0 (n_563), .A1 (g4311), .B0 (n_404), .Y (n_720));
INVX1 g68169(.A (n_719), .Y (n_1352));
INVX1 g66529(.A (n_1402), .Y (n_718));
XOR2X1 g66083(.A (n_716), .B (n_5958), .Y (n_717));
XOR2X1 g66079(.A (n_714), .B (n_5229), .Y (n_715));
INVX1 g66186(.A (n_10678), .Y (n_11221));
NOR2X1 g66508(.A (n_10213), .B (n_11187), .Y (n_10185));
OAI21X1 g65964(.A0 (n_2861), .A1 (n_3181), .B0 (g4473), .Y (n_709));
NOR2X1 g66863(.A (g5180), .B (g5188), .Y (n_1480));
OAI21X1 g65959(.A0 (g_10715), .A1 (n_708), .B0 (g_12791), .Y(n_1124));
NOR2X1 g66860(.A (g5527), .B (g5535), .Y (n_1476));
NOR2X1 g66746(.A (n_490), .B (n_11203), .Y (n_10809));
AND2X1 g66497(.A (n_730), .B (g2351), .Y (n_707));
NAND2X1 g65659(.A (n_1184), .B (n_1191), .Y (n_4314));
NOR2X1 g65762(.A (n_204), .B (n_7247), .Y (n_1219));
OR2X1 g62605(.A (g19334), .B (g7916), .Y (n_705));
INVX1 g66819(.A (n_1541), .Y (n_3323));
NAND2X1 g65728(.A (n_234), .B (n_2258), .Y (n_704));
INVX2 g68056(.A (n_2208), .Y (n_1023));
NAND2X1 g65717(.A (g2084), .B (n_7101), .Y (n_702));
NAND2X1 g65713(.A (n_745), .B (n_8796), .Y (n_698));
AND2X1 g66473(.A (n_806), .B (g1926), .Y (n_697));
XOR2X1 g65515(.A (g5084), .B (g5092), .Y (n_696));
AND2X1 g65515_and(.A (g5084), .B (g5092), .Y (n_1580));
XOR2X1 g65521(.A (g4258), .B (g4264), .Y (n_695));
AND2X1 g65521_and(.A (g4258), .B (g4264), .Y (n_1582));
XOR2X1 g65506(.A (n_11163), .B (g_20268), .Y (n_694));
AND2X1 g65506_and(.A (n_11163), .B (g_20268), .Y (n_693));
NOR2X1 g66394(.A (n_482), .B (g5188), .Y (n_1762));
NAND2X1 g66461(.A (g_21778), .B (n_691), .Y (n_692));
NAND2X1 g66435(.A (n_690), .B (g_3974), .Y (n_802));
INVX1 g68404(.A (n_10224), .Y (n_946));
XOR2X1 g66044(.A (g3827), .B (g3821), .Y (n_688));
CLKBUFX1 gbuf_d_1118(.A(g8719), .Y(d_out_1118));
CLKBUFX1 gbuf_q_1118(.A(q_in_1118), .Y(n_11116));
OR2X1 g66493(.A (n_3789), .B (g1728), .Y (n_3948));
CLKBUFX1 gbuf_d_1119(.A(g8788), .Y(d_out_1119));
CLKBUFX1 gbuf_q_1119(.A(q_in_1119), .Y(g8789));
OR2X1 g66490(.A (n_804), .B (g1760), .Y (n_1236));
AND2X1 g66456(.A (n_11110), .B (g_21318), .Y (n_1024));
NAND2X1 g66417(.A (g5511), .B (n_686), .Y (n_983));
NOR2X1 g66811(.A (g4991), .B (n_684), .Y (n_685));
NOR2X1 g64908(.A (n_19), .B (g4688), .Y (n_680));
NOR2X1 g64915(.A (g4688), .B (n_294), .Y (n_1307));
NOR2X1 g66452(.A (n_6922), .B (g_20208), .Y (n_876));
NOR2X1 g66450(.A (g3857), .B (n_678), .Y (n_1181));
NOR2X1 g66437(.A (g1657), .B (n_677), .Y (g25167));
NOR2X1 g65879(.A (n_20), .B (n_988), .Y (n_676));
AND2X1 g66442(.A (n_674), .B (g2060), .Y (n_675));
AND2X1 g66387(.A (n_661), .B (g6573), .Y (n_1391));
CLKBUFX1 gbuf_d_1120(.A(g7243), .Y(d_out_1120));
CLKBUFX1 gbuf_q_1120(.A(q_in_1120), .Y(g4405));
INVX1 g66781(.A (n_673), .Y (n_1222));
CLKBUFX1 gbuf_d_1121(.A(g17711), .Y(d_out_1121));
CLKBUFX1 gbuf_q_1121(.A(q_in_1121), .Y(g17580));
CLKBUFX1 gbuf_d_1122(.A(g8475), .Y(d_out_1122));
CLKBUFX1 gbuf_q_1122(.A(q_in_1122), .Y(g1333));
CLKBUFX1 gbuf_d_1123(.A(g19357), .Y(d_out_1123));
CLKBUFX1 gbuf_q_1123(.A(q_in_1123), .Y(g13272));
NAND2X1 g66418(.A (n_3943), .B (g1996), .Y (n_670));
CLKBUFX1 gbuf_d_1124(.A(g10500), .Y(d_out_1124));
CLKBUFX1 gbuf_q_1124(.A(q_in_1124), .Y(g1236));
NAND2X1 g66427(.A (n_3943), .B (g2070), .Y (n_667));
AND2X1 g66347(.A (n_626), .B (g3881), .Y (n_1364));
OR2X1 g66425(.A (n_3943), .B (g1996), .Y (n_4318));
NOR2X1 g66423(.A (n_128), .B (n_6979), .Y (n_4682));
NAND2X1 g66313(.A (n_11160), .B (g_6165), .Y (n_818));
NOR2X1 g66448(.A (n_10197), .B (n_224), .Y (n_978));
NOR2X1 g66433(.A (g3506), .B (n_664), .Y (n_1201));
MX2X1 g66131(.A (g_21806), .B (g_19241), .S0 (g_20268), .Y (n_1290));
INVX1 g65516(.A (n_982), .Y (n_663));
CLKBUFX1 gbuf_d_1125(.A(g13259), .Y(d_out_1125));
CLKBUFX1 gbuf_q_1125(.A(q_in_1125), .Y(n_10125));
NOR2X1 g66381(.A (n_661), .B (g6573), .Y (n_1718));
OAI21X1 g65629(.A0 (g6523), .A1 (g6537), .B0 (g35), .Y (n_1630));
CLKBUFX1 gbuf_d_1126(.A(g9251), .Y(d_out_1126));
CLKBUFX1 gbuf_q_1126(.A(q_in_1126), .Y(g4308));
CLKBUFX1 gbuf_d_1127(.A(g4467), .Y(d_out_1127));
CLKBUFX1 gbuf_q_1127(.A(q_in_1127), .Y(g4474));
XOR2X1 g66165(.A (g4308), .B (g9251), .Y (n_1570));
XOR2X1 g66179(.A (g1548), .B (g1430), .Y (n_652));
NAND3X1 g65815(.A (n_50), .B (g1178), .C (g_20614), .Y (n_1636));
XOR2X1 g66175(.A (g_22600), .B (g_22371), .Y (n_650));
NAND3X1 g65845(.A (g1367), .B (g1379), .C (g1345), .Y (n_1276));
MX2X1 g61436(.A (g10527), .B (g12923), .S0 (g17423), .Y (n_649));
INVX1 g66800(.A (n_647), .Y (n_648));
INVX1 g66740(.A (n_10622), .Y (n_10180));
XOR2X1 g66053(.A (g8786), .B (n_10867), .Y (n_643));
CLKBUFX1 gbuf_d_1128(.A(n_628), .Y(d_out_1128));
CLKBUFX1 gbuf_q_1128(.A(q_in_1128), .Y(g55));
INVX1 g66733(.A (n_4760), .Y (n_4791));
XOR2X1 g66074(.A (g5827), .B (g5821), .Y (n_639));
CLKBUFX1 gbuf_d_1129(.A(g17646), .Y(d_out_1129));
CLKBUFX1 gbuf_q_1129(.A(q_in_1129), .Y(g13068));
XOR2X1 g66076(.A (g3476), .B (g3470), .Y (n_638));
AOI22X1 g66088(.A0 (g2936), .A1 (g2941), .B0 (g2950), .B1 (g2955), .Y(n_637));
AOI22X1 g66089(.A0 (g_14342), .A1 (g_19414), .B0 (g_10715), .B1(g_12791), .Y (n_636));
OR2X1 g66378(.A (n_812), .B (g2453), .Y (n_1138));
OAI21X1 g61476(.A0 (g1395), .A1 (g1404), .B0 (g12923), .Y (n_635));
NAND2X1 g66455(.A (n_8587), .B (g_4050), .Y (n_800));
CLKBUFX1 gbuf_d_1130(.A(g8416), .Y(d_out_1130));
CLKBUFX1 gbuf_q_1130(.A(q_in_1130), .Y(g_15287));
XOR2X1 g66164(.A (g4281), .B (g8839), .Y (n_1820));
XOR2X1 g66176(.A (g_14535), .B (g8358), .Y (n_1732));
NOR2X1 g66375(.A (g1636), .B (n_629), .Y (g25259));
CLKBUFX1 gbuf_d_1131(.A(n_628), .Y(d_out_1131));
CLKBUFX1 gbuf_q_1131(.A(q_in_1131), .Y(g_9174));
CLKBUFX1 gbuf_d_1132(.A(g13099), .Y(d_out_1132));
CLKBUFX1 gbuf_q_1132(.A(q_in_1132), .Y(g17871));
CLKBUFX1 gbuf_d_1133(.A(g9553), .Y(d_out_1133));
CLKBUFX1 gbuf_qn_1133(.A(qn_in_1133), .Y(g5112));
CLKBUFX1 gbuf_d_1134(.A(g8291), .Y(d_out_1134));
CLKBUFX1 gbuf_q_1134(.A(q_in_1134), .Y(g_7220));
CLKBUFX1 gbuf_d_1135(.A(g13068), .Y(d_out_1135));
CLKBUFX1 gbuf_q_1135(.A(q_in_1135), .Y(g17819));
CLKBUFX1 gbuf_d_1136(.A(g13039), .Y(d_out_1136));
CLKBUFX1 gbuf_q_1136(.A(q_in_1136), .Y(g17787));
CLKBUFX1 gbuf_d_1137(.A(g13085), .Y(d_out_1137));
CLKBUFX1 gbuf_q_1137(.A(q_in_1137), .Y(g17845));
AND2X1 g66373(.A (g5857), .B (n_627), .Y (n_1194));
CLKBUFX1 gbuf_d_1138(.A(g10527), .Y(d_out_1138));
CLKBUFX1 gbuf_qn_1138(.A(qn_in_1138), .Y(g1579));
NOR2X1 g66712(.A (n_416), .B (n_251), .Y (n_1538));
AND2X1 g66371(.A (g6219), .B (n_617), .Y (n_1723));
NOR2X1 g66277(.A (n_626), .B (g3881), .Y (n_1743));
NOR2X1 g66278(.A (n_609), .B (g6395), .Y (n_3277));
NOR2X1 g66283(.A (n_674), .B (g2060), .Y (n_1515));
NAND2X1 g66285(.A (n_10369), .B (g_4409), .Y (n_823));
NOR2X1 g66293(.A (g3171), .B (n_553), .Y (n_1370));
NAND2X1 g66294(.A (n_6742), .B (g2629), .Y (n_624));
NOR2X1 g66307(.A (g3155), .B (n_623), .Y (n_1147));
NAND2X1 g66316(.A (g4608), .B (n_3624), .Y (n_747));
CLKBUFX1 gbuf_d_1139(.A(g17760), .Y(d_out_1139));
CLKBUFX1 gbuf_q_1139(.A(q_in_1139), .Y(g17649));
AND2X1 g66320(.A (g3506), .B (n_664), .Y (n_1207));
NAND2X1 g66333(.A (g5164), .B (n_621), .Y (n_817));
NOR2X1 g66336(.A (g5857), .B (n_627), .Y (n_1246));
AND2X1 g66345(.A (n_619), .B (g2217), .Y (n_620));
NAND2X1 g66346(.A (n_6742), .B (g2555), .Y (n_618));
OR2X1 g66354(.A (n_806), .B (g1894), .Y (n_1230));
NOR2X1 g66366(.A (n_11071), .B (n_134), .Y (n_2600));
NOR2X1 g66367(.A (g6219), .B (n_617), .Y (n_1377));
NOR2X1 g66368(.A (n_619), .B (g2217), .Y (n_1520));
AND2X1 g66382(.A (n_11165), .B (g_8864), .Y (n_1011));
AND2X1 g66384(.A (g3155), .B (n_623), .Y (n_1243));
AND2X1 g66385(.A (n_11071), .B (n_134), .Y (n_3275));
NOR2X1 g66389(.A (n_616), .B (g3530), .Y (n_1751));
AND2X1 g66407(.A (n_616), .B (g3530), .Y (n_1367));
XOR2X1 g66073(.A (g3125), .B (g3119), .Y (n_615));
AND2X1 g66424(.A (g6203), .B (n_612), .Y (n_1158));
AND2X1 g66428(.A (n_610), .B (g2619), .Y (n_611));
AND2X1 g66460(.A (n_609), .B (g6395), .Y (n_2325));
OR2X1 g66465(.A (n_4301), .B (g2153), .Y (n_4109));
AND2X1 g66469(.A (g1657), .B (n_677), .Y (n_608));
OR2X1 g66487(.A (n_3939), .B (g2421), .Y (n_4122));
NOR2X1 g66494(.A (n_8637), .B (n_10818), .Y (n_607));
AND2X1 g66507(.A (n_10197), .B (n_224), .Y (n_1179));
OR2X1 g66513(.A (g4608), .B (n_3624), .Y (n_1831));
NOR2X1 g66519(.A (n_610), .B (g2619), .Y (n_1506));
AND2X1 g66523(.A (g3857), .B (n_678), .Y (n_1185));
NOR2X1 g66531(.A (n_610), .B (g2587), .Y (n_1522));
OR2X1 g66532(.A (n_3782), .B (g1862), .Y (n_3945));
OR2X1 g66536(.A (g6549), .B (n_603), .Y (n_791));
NOR2X1 g66538(.A (g6203), .B (n_612), .Y (n_1149));
NOR2X1 g66551(.A (n_95), .B (g_17426), .Y (n_3391));
AND2X1 g66553(.A (n_455), .B (n_11198), .Y (n_11101));
XOR2X1 g66010(.A (g6519), .B (g6513), .Y (n_600));
OR2X1 g66357(.A (g1592), .B (n_347), .Y (n_3938));
NOR2X1 g66570(.A (n_598), .B (g4966), .Y (n_599));
AND2X1 g66571(.A (n_191), .B (n_10657), .Y (n_2597));
NAND2X1 g66572(.A (g4388), .B (n_596), .Y (n_597));
NAND2X1 g66573(.A (g4430), .B (n_596), .Y (n_595));
NAND2X1 g66575(.A (n_10139), .B (n_6967), .Y (n_1173));
AND2X1 g66577(.A (n_6979), .B (n_128), .Y (n_11128));
AND2X1 g66582(.A (n_401), .B (g_3381), .Y (n_1093));
INVX1 g66586(.A (n_1267), .Y (n_594));
INVX1 g66603(.A (n_1468), .Y (n_1143));
INVX1 g66605(.A (n_591), .Y (n_592));
NAND2X1 g66617(.A (n_627), .B (n_215), .Y (n_589));
NOR2X1 g66624(.A (n_413), .B (n_456), .Y (n_588));
NAND2X1 g66635(.A (n_603), .B (n_261), .Y (n_587));
INVX1 g66646(.A (n_1486), .Y (n_585));
NOR2X1 g66653(.A (n_10630), .B (n_10634), .Y (n_584));
INVX1 g66666(.A (n_908), .Y (n_581));
NAND2X1 g66675(.A (n_664), .B (n_365), .Y (n_580));
INVX1 g66708(.A (n_6790), .Y (n_579));
NAND2X1 g66717(.A (n_686), .B (n_383), .Y (n_578));
INVX1 g66722(.A (n_970), .Y (n_1224));
NOR2X1 g66350(.A (n_619), .B (g2185), .Y (n_1527));
NAND2X1 g66764(.A (n_678), .B (n_303), .Y (n_575));
NOR2X1 g66768(.A (n_10228), .B (n_10225), .Y (n_8778));
INVX1 g66770(.A (n_411), .Y (n_1264));
NOR2X1 g66775(.A (n_10139), .B (n_379), .Y (n_771));
NAND2X1 g66791(.A (n_572), .B (n_571), .Y (n_2111));
INVX1 g66794(.A (n_1145), .Y (n_1459));
INVX1 g66802(.A (n_1464), .Y (n_1227));
OR2X1 g66806(.A (g8475), .B (g7946), .Y (n_568));
NAND2X1 g66825(.A (n_612), .B (n_330), .Y (n_566));
NAND2X1 g66827(.A (n_623), .B (n_370), .Y (n_565));
NAND2X1 g66830(.A (n_563), .B (n_327), .Y (n_564));
INVX1 g66841(.A (n_561), .Y (n_562));
INVX1 g66854(.A (n_7101), .Y (n_558));
CLKBUFX1 gbuf_d_1140(.A(g19334), .Y(d_out_1140));
CLKBUFX1 gbuf_q_1140(.A(q_in_1140), .Y(g13259));
INVX1 g66868(.A (n_7024), .Y (n_557));
OR2X1 g66874(.A (g19357), .B (g7946), .Y (n_556));
NOR2X1 g66889(.A (n_297), .B (n_406), .Y (n_3365));
AND2X1 g66343(.A (g3171), .B (n_553), .Y (n_1758));
INVX1 g66919(.A (n_552), .Y (n_723));
CLKBUFX1 gbuf_d_1141(.A(g17400), .Y(d_out_1141));
CLKBUFX1 gbuf_q_1141(.A(q_in_1141), .Y(g_18330));
CLKBUFX1 gbuf_d_1142(.A(g34036), .Y(d_out_1142));
CLKBUFX1 gbuf_qn_1142(.A(qn_in_1142), .Y(g4878));
XOR2X1 g66001(.A (g5128), .B (g5134), .Y (n_540));
INVX1 g66664(.A (n_973), .Y (n_1154));
NOR2X1 g66311(.A (n_522), .B (g5535), .Y (n_1777));
CLKBUFX1 gbuf_d_1143(.A(g17604), .Y(d_out_1143));
CLKBUFX1 gbuf_q_1143(.A(q_in_1143), .Y(g13049));
NOR2X1 g66337(.A (g1389), .B (n_6782), .Y (n_3364));
CLKBUFX1 gbuf_d_1144(.A(g14738), .Y(d_out_1144));
CLKBUFX1 gbuf_q_1144(.A(q_in_1144), .Y(g17739));
CLKBUFX1 gbuf_d_1145(.A(g34035), .Y(d_out_1145));
CLKBUFX1 gbuf_q_1145(.A(q_in_1145), .Y(g34036));
INVX1 g66669(.A (n_901), .Y (n_1212));
CLKBUFX1 gbuf_d_1146(.A(g14694), .Y(d_out_1146));
CLKBUFX1 gbuf_q_1146(.A(q_in_1146), .Y(g17711));
CLKBUFX1 gbuf_d_1147(.A(g17404), .Y(d_out_1147));
CLKBUFX1 gbuf_q_1147(.A(q_in_1147), .Y(g17423));
CLKBUFX1 gbuf_d_1148(.A(g17739), .Y(d_out_1148));
CLKBUFX1 gbuf_q_1148(.A(q_in_1148), .Y(g17607));
CLKBUFX1 gbuf_d_1149(.A(g17778), .Y(d_out_1149));
CLKBUFX1 gbuf_q_1149(.A(q_in_1149), .Y(g17688));
CLKBUFX1 gbuf_d_1150(.A(g17577), .Y(d_out_1150));
CLKBUFX1 gbuf_q_1150(.A(q_in_1150), .Y(g13039));
NAND2X1 g66329(.A (n_103), .B (n_11050), .Y (n_1100));
AND2X1 g66658(.A (n_523), .B (g6736), .Y (n_524));
AND2X1 g66325(.A (n_522), .B (g5535), .Y (n_1411));
NOR2X1 g66655(.A (n_8913), .B (n_10818), .Y (n_521));
INVX1 g68267(.A (n_10314), .Y (n_519));
MX2X1 g61555(.A (g10500), .B (g12919), .S0 (g17400), .Y (n_515));
CLKBUFX1 gbuf_d_1151(.A(g7257), .Y(d_out_1151));
CLKBUFX1 gbuf_q_1151(.A(q_in_1151), .Y(g4411));
CLKBUFX1 gbuf_d_1152(.A(g7245), .Y(d_out_1152));
CLKBUFX1 gbuf_q_1152(.A(q_in_1152), .Y(g4452));
INVX1 g67211(.A (g4584), .Y (n_3624));
NOR2X1 g66304(.A (n_512), .B (g4601), .Y (n_820));
CLKBUFX1 gbuf_d_1153(.A(g12919), .Y(d_out_1153));
CLKBUFX1 gbuf_qn_1153(.A(qn_in_1153), .Y(g1242));
OR2X1 g66301(.A (g5164), .B (n_621), .Y (n_822));
OR2X1 g66379(.A (g2984), .B (n_628), .Y (n_511));
NAND3X1 g65813(.A (g_22306), .B (g_12465), .C (g_19911), .Y (n_989));
OR2X1 g66290(.A (n_6742), .B (g2555), .Y (n_4118));
CLKBUFX1 gbuf_d_1154(.A(g17316), .Y(d_out_1154));
CLKBUFX1 gbuf_q_1154(.A(q_in_1154), .Y(g17400));
INVX1 g68012(.A (n_503), .Y (n_504));
INVX2 g68057(.A (n_776), .Y (n_2208));
CLKBUFX1 gbuf_d_1155(.A(g13049), .Y(d_out_1155));
CLKBUFX1 gbuf_q_1155(.A(q_in_1155), .Y(g17813));
INVX1 g68119(.A (n_10245), .Y (n_2177));
OAI21X1 g61586(.A0 (g_18488), .A1 (n_8508), .B0 (g12919), .Y (n_496));
INVX4 g67034(.A (n_546), .Y (n_2421));
CLKBUFX1 g68332(.A (n_490), .Y (n_4980));
AND2X1 g66569(.A (n_11038), .B (n_8807), .Y (n_2339));
INVX1 g66906(.A (n_896), .Y (n_1482));
NAND2X1 g66486(.A (n_453), .B (g_19172), .Y (n_799));
INVX1 g68244(.A (n_488), .Y (n_2017));
CLKBUFX1 gbuf_d_1156(.A(g10122), .Y(d_out_1156));
CLKBUFX1 gbuf_q_1156(.A(q_in_1156), .Y(g4297));
CLKBUFX1 gbuf_d_1157(.A(g17320), .Y(d_out_1157));
CLKBUFX1 gbuf_q_1157(.A(q_in_1157), .Y(g17404));
OR2X1 g66506(.A (g5511), .B (n_686), .Y (n_795));
INVX1 g66872(.A (n_486), .Y (n_487));
INVX1 g68170(.A (g_20952), .Y (n_719));
AND2X1 g66530(.A (n_482), .B (g5188), .Y (n_1402));
CLKBUFX1 gbuf_d_1158(.A(g17685), .Y(d_out_1158));
CLKBUFX1 gbuf_q_1158(.A(q_in_1158), .Y(g13085));
AND2X1 g66526(.A (g6549), .B (n_603), .Y (n_1395));
OR2X1 g66521(.A (n_730), .B (g2319), .Y (n_1160));
NAND2X1 g66883(.A (n_621), .B (n_388), .Y (n_479));
CLKBUFX1 gbuf_d_1159(.A(g9019), .Y(d_out_1159));
CLKBUFX1 gbuf_q_1159(.A(q_in_1159), .Y(g4291));
OR2X1 g66511(.A (n_4038), .B (g2287), .Y (n_4124));
INVX1 g66864(.A (n_4631), .Y (n_4679));
INVX1 g65512(.A (n_474), .Y (n_971));
CLKBUFX1 gbuf_d_1160(.A(g17674), .Y(d_out_1160));
CLKBUFX1 gbuf_q_1160(.A(q_in_1160), .Y(g17519));
CLKBUFX1 gbuf_d_1161(.A(g14662), .Y(d_out_1161));
CLKBUFX1 gbuf_q_1161(.A(q_in_1161), .Y(g17674));
CLKBUFX1 gbuf_d_1162(.A(g13272), .Y(d_out_1162));
CLKBUFX1 gbuf_q_1162(.A(q_in_1162), .Y(g1322));
CLKBUFX1 gbuf_d_1163(.A(g11447), .Y(d_out_1163));
CLKBUFX1 gbuf_q_1163(.A(q_in_1163), .Y(g8783));
CLKBUFX1 gbuf_d_1164(.A(g17423), .Y(d_out_1164));
CLKBUFX1 gbuf_q_1164(.A(q_in_1164), .Y(g1430));
CLKBUFX1 gbuf_d_1165(.A(g8783), .Y(d_out_1165));
CLKBUFX1 gbuf_q_1165(.A(q_in_1165), .Y(g8784));
CLKBUFX1 gbuf_d_1166(.A(g8785), .Y(d_out_1166));
CLKBUFX1 gbuf_q_1166(.A(q_in_1166), .Y(g8786));
CLKBUFX1 gbuf_d_1167(.A(g8358), .Y(d_out_1167));
CLKBUFX1 gbuf_q_1167(.A(q_in_1167), .Y(g_14535));
CLKBUFX1 gbuf_d_1168(.A(g14779), .Y(d_out_1168));
CLKBUFX1 gbuf_q_1168(.A(q_in_1168), .Y(g17760));
CLKBUFX1 gbuf_d_1169(.A(g12923), .Y(d_out_1169));
CLKBUFX1 gbuf_qn_1169(.A(qn_in_1169), .Y(g1585));
NAND3X1 g65763(.A (g_10715), .B (g_15740), .C (g_12791), .Y (n_471));
XOR2X1 g66064(.A (g4388), .B (g4430), .Y (n_470));
XOR2X1 g66167(.A (n_10128), .B (g_18330), .Y (n_469));
INVX2 g66848(.A (n_10426), .Y (n_3459));
CLKBUFX1 gbuf_d_1170(.A(g17291), .Y(d_out_1170));
CLKBUFX1 gbuf_q_1170(.A(q_in_1170), .Y(g17316));
CLKBUFX1 gbuf_d_1171(.A(g7260), .Y(d_out_1171));
CLKBUFX1 gbuf_q_1171(.A(q_in_1171), .Y(g4443));
NOR2X1 g66491(.A (n_674), .B (g2028), .Y (n_1524));
CLKBUFX1 gbuf_d_1172(.A(g17722), .Y(d_out_1172));
CLKBUFX1 gbuf_q_1172(.A(q_in_1172), .Y(g13099));
INVX1 g68094(.A (n_10213), .Y (n_740));
CLKBUFX1 gbuf_d_1173(.A(g8839), .Y(d_out_1173));
CLKBUFX1 gbuf_q_1173(.A(q_in_1173), .Y(g4281));
INVX1 g67943(.A (n_464), .Y (g11349));
NOR2X1 g66488(.A (g1624), .B (n_677), .Y (n_1531));
INVX1 g66600(.A (n_1199), .Y (n_463));
XOR2X1 g66162(.A (g4291), .B (g9019), .Y (n_1556));
AND2X1 g66580(.A (n_459), .B (g5881), .Y (n_1382));
NAND2X1 g61309(.A (g1521), .B (n_460), .Y (n_461));
NOR2X1 g66480(.A (n_459), .B (g5881), .Y (n_1725));
INVX1 g66815(.A (n_1175), .Y (n_458));
CLKBUFX1 gbuf_d_1174(.A(g8784), .Y(d_out_1174));
CLKBUFX1 gbuf_q_1174(.A(q_in_1174), .Y(g8785));
CLKBUFX1 gbuf_d_1175(.A(g8786), .Y(d_out_1175));
CLKBUFX1 gbuf_q_1175(.A(q_in_1175), .Y(g8787));
CLKBUFX1 g66820(.A (n_6762), .Y (n_1541));
CLKBUFX1 gbuf_d_1176(.A(g8789), .Y(d_out_1176));
CLKBUFX1 gbuf_q_1176(.A(q_in_1176), .Y(n_10871));
NAND2X1 g66475(.A (g1442), .B (n_412), .Y (n_1729));
CLKBUFX1 gbuf_d_1177(.A(g8787), .Y(d_out_1177));
CLKBUFX1 gbuf_q_1177(.A(q_in_1177), .Y(g8788));
INVX1 g68017(.A (n_1285), .Y (n_456));
INVX1 g67958(.A (n_2150), .Y (n_1540));
CLKBUFX1 gbuf_d_1178(.A(g14828), .Y(d_out_1178));
CLKBUFX1 gbuf_q_1178(.A(q_in_1178), .Y(g17778));
NOR2X1 g66552(.A (n_455), .B (n_11198), .Y (n_10508));
INVX1 g68333(.A (n_455), .Y (n_490));
NOR2X1 g66641(.A (g6336), .B (g6395), .Y (n_2413));
NOR2X1 g66809(.A (g2098), .B (g1964), .Y (n_442));
INVX1 g68245(.A (g_20951), .Y (n_488));
NOR2X1 g66805(.A (g1894), .B (g1926), .Y (n_441));
NAND2X1 g66804(.A (g_18330), .B (n_10128), .Y (n_474));
NAND2X1 g66801(.A (g1894), .B (g1926), .Y (n_647));
OR2X1 g66786(.A (g2537), .B (g2417), .Y (n_436));
AND2X1 g66816(.A (g3857), .B (g3863), .Y (n_1175));
INVX1 g67902(.A (g34034), .Y (n_477));
NAND2X1 g66760(.A (g1548), .B (g1430), .Y (n_982));
OR2X1 g66778(.A (g2338), .B (g2491), .Y (n_429));
NOR2X1 g66730(.A (g1844), .B (g1710), .Y (n_428));
INVX1 g68229(.A (n_6782), .Y (n_1275));
NOR2X1 g66885(.A (n_11071), .B (g6741), .Y (n_2435));
NOR2X1 g66792(.A (g2126), .B (g1992), .Y (n_425));
INVX1 g61358(.A (n_460), .Y (n_2474));
INVX1 g67026(.A (n_423), .Y (n_424));
INVX1 g67975(.A (n_417), .Y (n_659));
AND2X1 g66795(.A (g5857), .B (g5863), .Y (n_1145));
OR2X1 g61462(.A (g1404), .B (g12923), .Y (n_415));
NAND2X1 g66771(.A (g6219), .B (g6227), .Y (n_411));
INVX2 g67915(.A (n_690), .Y (n_5402));
INVX1 g67886(.A (g12238), .Y (n_465));
INVX1 g67798(.A (n_409), .Y (g12300));
NOR2X1 g66696(.A (g2453), .B (g2485), .Y (n_408));
INVX1 g67783(.A (n_6922), .Y (n_5663));
AND2X1 g66796(.A (g3873), .B (g3881), .Y (n_1184));
INVX1 g68058(.A (n_401), .Y (n_776));
NOR2X1 g65890(.A (g34035), .B (g34036), .Y (n_1578));
AND2X1 g66731(.A (g6336), .B (g6395), .Y (n_2352));
NOR2X1 g66728(.A (g2319), .B (g2351), .Y (n_376));
INVX1 g67169(.A (g17688), .Y (n_538));
NAND2X1 g66716(.A (g5124), .B (g35), .Y (n_3641));
AND2X1 g66718(.A (n_10660), .B (g5698), .Y (n_374));
INVX1 g67984(.A (n_367), .Y (n_2252));
INVX1 g68445(.A (g12422), .Y (n_660));
INVX1 g67009(.A (g17580), .Y (n_669));
NOR2X1 g66721(.A (g1664), .B (g1644), .Y (n_353));
AND2X1 g66723(.A (g5180), .B (g5188), .Y (n_970));
NAND2X1 g66724(.A (g4467), .B (g4473), .Y (n_1353));
NOR2X1 g66584(.A (g4141), .B (g4082), .Y (n_1312));
NOR2X1 g66587(.A (g4311), .B (n_662), .Y (n_1267));
NOR2X1 g66597(.A (g8787), .B (g8786), .Y (n_344));
AND2X1 g66907(.A (g3155), .B (g3161), .Y (n_896));
NOR2X1 g66620(.A (g6177), .B (g6191), .Y (n_343));
NAND2X1 g66627(.A (g2629), .B (g2555), .Y (n_342));
AND2X1 g66629(.A (n_10657), .B (g5644), .Y (n_2443));
AND2X1 g66902(.A (n_7247), .B (g4621), .Y (n_948));
NOR2X1 g66657(.A (g2685), .B (g2551), .Y (n_340));
AND2X1 g66673(.A (g2185), .B (g2217), .Y (n_1517));
AND2X1 g66686(.A (g6395), .B (g6390), .Y (n_339));
AND2X1 g66692(.A (g6509), .B (g35), .Y (n_3812));
NOR2X1 g66739(.A (g1624), .B (g1657), .Y (n_338));
NOR2X1 g66754(.A (g2587), .B (g2619), .Y (n_336));
NAND2X1 g66803(.A (g5164), .B (g5170), .Y (n_1464));
AND2X1 g66813(.A (n_11071), .B (g6741), .Y (n_2432));
NOR2X1 g66834(.A (g2066), .B (g2047), .Y (n_335));
OR2X1 g66838(.A (g7260), .B (g7245), .Y (n_334));
NAND2X1 g66842(.A (g1760), .B (g1792), .Y (n_561));
INVX1 g68439(.A (g11418), .Y (n_491));
AND2X1 g66873(.A (g2453), .B (g2485), .Y (n_486));
NOR2X1 g66886(.A (g1183), .B (n_8769), .Y (n_746));
AND2X1 g66699(.A (g3171), .B (g3179), .Y (n_1242));
INVX2 g67035(.A (n_423), .Y (n_546));
AND2X1 g66742(.A (g5873), .B (g5881), .Y (n_1245));
NOR2X1 g66725(.A (n_10657), .B (g5644), .Y (n_2439));
AND2X1 g66665(.A (g5527), .B (g5535), .Y (n_973));
OR2X1 g61584(.A (n_8508), .B (g12919), .Y (n_325));
AND2X1 g66670(.A (g3115), .B (g35), .Y (n_901));
NOR2X1 g66702(.A (g1760), .B (g1792), .Y (n_323));
INVX1 g68290(.A (n_322), .Y (g12470));
OR2X1 g66824(.A (g7257), .B (g7243), .Y (n_316));
NOR2X1 g66808(.A (g4153), .B (g4172), .Y (n_311));
OR2X1 g66652(.A (g17404), .B (g17320), .Y (n_309));
INVX1 g68232(.A (n_307), .Y (n_518));
NAND2X1 g66647(.A (g6549), .B (g6555), .Y (n_1486));
NOR2X1 g66871(.A (g4054), .B (g3990), .Y (n_4988));
OR2X1 g66861(.A (g1978), .B (g1858), .Y (n_302));
OR2X1 g66630(.A (g1779), .B (g1932), .Y (n_298));
OR2X1 g66831(.A (g17316), .B (g17291), .Y (n_295));
NAND2X1 g66881(.A (g2070), .B (g1996), .Y (n_290));
AND2X1 g66615(.A (g6565), .B (g6573), .Y (n_590));
NAND2X1 g66604(.A (g6203), .B (g6209), .Y (n_1468));
AND2X1 g66601(.A (g3506), .B (g3512), .Y (n_1199));
NAND2X1 g66782(.A (g5511), .B (g5517), .Y (n_673));
NAND2X1 g66691(.A (g5037), .B (g5033), .Y (n_281));
INVX1 g68274(.A (n_598), .Y (n_653));
INVX4 g68390(.A (g7946), .Y (n_3849));
AND2X1 g66772(.A (n_11201), .B (g6044), .Y (n_268));
INVX1 g66986(.A (g17649), .Y (n_549));
INVX1 g66943(.A (n_684), .Y (n_551));
INVX1 g68184(.A (n_276), .Y (n_3181));
NOR2X1 g66908(.A (g2403), .B (g2269), .Y (n_248));
INVX2 g66920(.A (n_10634), .Y (n_552));
NAND2X1 g61629(.A (g4401), .B (g4434), .Y (n_243));
NOR2X1 g66901(.A (g1830), .B (g1696), .Y (n_241));
NOR2X1 g66895(.A (g2028), .B (g2060), .Y (n_240));
NOR2X1 g66896(.A (g_20073), .B (g_12433), .Y (n_891));
INVX1 g68324(.A (g13966), .Y (n_493));
AND2X1 g66690(.A (g3522), .B (g3530), .Y (n_1206));
NOR2X1 g66890(.A (g2625), .B (g2606), .Y (n_235));
NAND2X1 g66880(.A (g5471), .B (g35), .Y (n_6399));
NOR2X1 g66887(.A (g2185), .B (g2217), .Y (n_234));
AND2X1 g66748(.A (g1183), .B (n_8769), .Y (n_745));
INVX1 g67875(.A (g17519), .Y (n_527));
INVX1 g68277(.A (n_1627), .Y (n_227));
INVX1 g68158(.A (n_691), .Y (n_3550));
INVX1 g68147(.A (n_224), .Y (n_2773));
INVX1 g68142(.A (n_223), .Y (n_3439));
NOR2X1 g66875(.A (n_10197), .B (g1526), .Y (n_899));
NOR2X1 g66866(.A (g1442), .B (g1489), .Y (n_4631));
AND2X1 g66857(.A (n_6979), .B (g3639), .Y (n_6973));
OR2X1 g66839(.A (g11447), .B (g8789), .Y (n_220));
NAND2X1 g66862(.A (g4669), .B (g4653), .Y (n_218));
AND2X1 g66667(.A (n_10197), .B (g1526), .Y (n_908));
AND2X1 g66651(.A (g1322), .B (g1404), .Y (n_1165));
NOR2X1 g66735(.A (g_18902), .B (g_19172), .Y (n_4760));
INVX1 g67944(.A (g_4050), .Y (n_464));
NAND2X1 g66694(.A (g4146), .B (g4157), .Y (n_209));
NOR2X1 g66648(.A (n_6958), .B (g_21651), .Y (n_205));
NAND2X1 g66845(.A (g4621), .B (g4633), .Y (n_204));
NOR2X1 g66783(.A (g5046), .B (g5052), .Y (n_196));
NOR2X1 g66835(.A (g2223), .B (g2204), .Y (n_194));
AND2X1 g66606(.A (g2319), .B (g2351), .Y (n_591));
INVX1 g67208(.A (n_191), .Y (n_4982));
NOR2X1 g66833(.A (g4087), .B (g4098), .Y (n_188));
AND2X1 g66828(.A (n_8509), .B (n_10125), .Y (n_8796));
INVX1 g68344(.A (n_8637), .Y (n_644));
INVX1 g68013(.A (n_10630), .Y (n_503));
CLKBUFX1 g67959(.A (n_8594), .Y (n_2150));
INVX1 g67122(.A (g2667), .Y (n_716));
INVX1 g68456(.A (g_16464), .Y (n_172));
INVX1 g66913(.A (n_3604), .Y (n_247));
INVX1 g67920(.A (g2040), .Y (n_3943));
INVX1 g67195(.A (g2295), .Y (n_1702));
INVX1 g68291(.A (g_8864), .Y (n_322));
INVX1 g68248(.A (g1959), .Y (n_836));
INVX1 g68114(.A (g2250), .Y (n_382));
INVX1 g68367(.A (g2303), .Y (n_1703));
INVX1 g68214(.A (g2704), .Y (n_169));
INVX1 g67742(.A (g5134), .Y (n_168));
INVX1 g68315(.A (g3133), .Y (n_2686));
INVX1 g68117(.A (g3490), .Y (n_1799));
INVX1 g67182(.A (g4653), .Y (n_294));
INVX1 g68211(.A (g4849), .Y (n_165));
INVX1 g67827(.A (g2856), .Y (n_3499));
INVX1 g68217(.A (g2177), .Y (n_919));
INVX1 g68338(.A (n_640), .Y (n_273));
INVX1 g68190(.A (g3147), .Y (n_3253));
INVX1 g67177(.A (g4462), .Y (n_2861));
CLKBUFX1 g68440(.A (g_3974), .Y (g11418));
INVX1 g66950(.A (g_20909), .Y (n_6324));
INVX1 g66955(.A (g2246), .Y (n_4906));
INVX1 g68353(.A (g2988), .Y (n_162));
INVX1 g68354(.A (g1564), .Y (n_1295));
INVX1 g68086(.A (n_3611), .Y (n_202));
INVX1 g67830(.A (g2571), .Y (n_362));
INVX1 g67126(.A (g6519), .Y (n_158));
INVX1 g68357(.A (g5517), .Y (n_686));
INVX1 g67846(.A (g2472), .Y (n_157));
INVX1 g68166(.A (g2527), .Y (n_5229));
INVX1 g68213(.A (g_18112), .Y (n_153));
INVX1 g67039(.A (g2864), .Y (n_271));
INVX1 g67752(.A (g13926), .Y (n_242));
INVX1 g68377(.A (g2898), .Y (n_3501));
INVX1 g67862(.A (g6555), .Y (n_603));
INVX1 g67747(.A (g1834), .Y (n_4948));
INVX1 g68327(.A (g2399), .Y (n_846));
INVX1 g68308(.A (g4035), .Y (n_151));
INVX1 g68254(.A (g4239), .Y (n_150));
INVX1 g67025(.A (g5170), .Y (n_621));
INVX1 g67093(.A (n_1234), .Y (n_383));
INVX1 g66916(.A (g1882), .Y (n_2306));
INVX1 g67012(.A (g2380), .Y (n_4529));
INVX1 g68263(.A (g2315), .Y (n_1677));
INVX1 g67925(.A (g2016), .Y (n_926));
INVX1 g68104(.A (g2384), .Y (n_831));
INVX1 g66997(.A (g5503), .Y (n_2943));
INVX1 g68394(.A (g2122), .Y (n_860));
INVX1 g67989(.A (g2648), .Y (n_4726));
INVX1 g68048(.A (g5406), .Y (n_144));
CLKBUFX1 g67842(.A (g6741), .Y (n_523));
INVX1 g67096(.A (g4659), .Y (n_143));
INVX1 g66970(.A (g2563), .Y (n_380));
INVX1 g68154(.A (g4515), .Y (n_563));
INVX1 g67209(.A (g5644), .Y (n_191));
INVX1 g67203(.A (g2197), .Y (n_4301));
INVX1 g67980(.A (g5849), .Y (n_2940));
INVX1 g67869(.A (g3139), .Y (n_1805));
INVX1 g68298(.A (g4382), .Y (n_5363));
INVX1 g67818(.A (g4593), .Y (n_512));
INVX1 g66962(.A (g2116), .Y (n_6017));
INVX1 g68198(.A (n_2005), .Y (n_412));
INVX1 g67215(.A (g1768), .Y (n_136));
INVX1 g68317(.A (g2643), .Y (n_902));
INVX1 g67099(.A (g1714), .Y (n_6027));
INVX1 g68261(.A (g3841), .Y (n_1796));
INVX1 g66959(.A (n_3589), .Y (n_332));
INVX1 g67864(.A (g1454), .Y (n_2538));
INVX1 g68078(.A (g3684), .Y (n_1818));
INVX1 g67843(.A (g6741), .Y (n_134));
INVX1 g67790(.A (g13895), .Y (n_238));
INVX1 g68365(.A (g2449), .Y (n_1671));
INVX1 g66262(.A (g34027), .Y (n_988));
INVX1 g67966(.A (g2008), .Y (n_1514));
INVX1 g68436(.A (g1848), .Y (n_5978));
INVX1 g67108(.A (g2012), .Y (n_368));
INVX1 g67155(.A (n_5936), .Y (n_677));
INVX1 g68016(.A (g1706), .Y (n_856));
INVX1 g68084(.A (g2361), .Y (n_386));
INVX1 g66980(.A (n_5928), .Y (n_610));
INVX1 g67871(.A (g2279), .Y (n_975));
INVX1 g68124(.A (g2024), .Y (n_278));
INVX1 g67780(.A (g3522), .Y (n_616));
INVX1 g68305(.A (g1982), .Y (n_5975));
INVX1 g68304(.A (g2020), .Y (n_399));
INVX1 g67103(.A (g2407), .Y (n_5972));
INVX1 g67083(.A (g_18488), .Y (n_129));
INVX1 g68260(.A (g1604), .Y (n_1509));
INVX1 g61359(.A (g1339), .Y (n_460));
INVX1 g67991(.A (g2413), .Y (n_866));
INVX1 g68027(.A (g3639), .Y (n_128));
INVX1 g67976(.A (g_16475), .Y (n_417));
INVX1 g67097(.A (g6098), .Y (n_127));
INVX1 g68165(.A (g6565), .Y (n_661));
INVX1 g66914(.A (g5863), .Y (n_627));
INVX1 g68143(.A (g_15016), .Y (n_223));
INVX1 g68296(.A (g20899), .Y (n_2518));
INVX1 g68074(.A (g2917), .Y (n_3463));
INVX1 g67897(.A (n_3616), .Y (n_356));
INVX1 g67930(.A (g_16958), .Y (n_416));
INVX1 g68180(.A (g4601), .Y (n_262));
CLKBUFX1 g68031(.A (g6336), .Y (n_4978));
INVX1 g67753(.A (g_19414), .Y (n_126));
INVX1 g67006(.A (g2681), .Y (n_852));
INVX1 g66991(.A (g6173), .Y (n_125));
INVX1 g67824(.A (g6181), .Y (n_2704));
INVX1 g68415(.A (g6527), .Y (n_3007));
INVX1 g68102(.A (g2145), .Y (n_308));
INVX1 g67934(.A (g2004), .Y (n_450));
INVX1 g68041(.A (g_12791), .Y (n_413));
INVX1 g67148(.A (g_22306), .Y (n_286));
INVX1 g66978(.A (n_1214), .Y (n_330));
INVX1 g67956(.A (g6195), .Y (n_2936));
INVX1 g68209(.A (g1906), .Y (n_3782));
INVX1 g68173(.A (g6209), .Y (n_612));
INVX1 g67014(.A (g2299), .Y (n_1676));
INVX1 g68116(.A (g1437), .Y (n_2535));
INVX1 g66941(.A (n_4339), .Y (n_437));
INVX1 g66938(.A (g2181), .Y (n_1519));
INVX1 g68236(.A (n_5921), .Y (n_812));
INVX1 g67811(.A (g2138), .Y (n_1240));
INVX1 g68408(.A (g1691), .Y (n_187));
INVX1 g67765(.A (g6541), .Y (n_2930));
INVX1 g68225(.A (g3498), .Y (n_2928));
INVX1 g68363(.A (g_21447), .Y (n_3310));
INVX1 g67200(.A (g2771), .Y (n_326));
INVX1 g67806(.A (g1608), .Y (n_1533));
INVX1 g67171(.A (g3161), .Y (n_623));
INVX1 g68196(.A (g1600), .Y (n_1532));
INVX1 g68362(.A (g2533), .Y (n_714));
INVX1 g67756(.A (g3457), .Y (n_3601));
INVX1 g67088(.A (g_20839), .Y (n_2280));
INVX1 g68370(.A (g2583), .Y (n_213));
INVX1 g68201(.A (g4076), .Y (n_118));
INVX1 g67011(.A (g3752), .Y (n_117));
INVX1 g68360(.A (g1379), .Y (n_263));
INVX1 g66935(.A (g2331), .Y (n_4038));
INVX1 g67891(.A (g55), .Y (n_628));
INVX1 g67150(.A (g5873), .Y (n_459));
INVX1 g67949(.A (g1467), .Y (n_2485));
INVX1 g67218(.A (g2429), .Y (n_1713));
INVX1 g68218(.A (g5835), .Y (n_2684));
INVX1 g68334(.A (g5990), .Y (n_455));
INVX1 g68109(.A (n_3618), .Y (n_389));
INVX1 g68282(.A (g1720), .Y (n_878));
INVX1 g66964(.A (g3808), .Y (n_3596));
INVX1 g68233(.A (g1221), .Y (n_307));
INVX1 g68356(.A (g5527), .Y (n_522));
INVX1 g67812(.A (g4843), .Y (n_1274));
INVX1 g68379(.A (n_2458), .Y (n_397));
INVX1 g66925(.A (g_20159), .Y (n_251));
INVX2 g67916(.A (g4040), .Y (n_690));
INVX1 g67884(.A (g5057), .Y (n_110));
INVX1 g67947(.A (g1322), .Y (n_1502));
INVX1 g67939(.A (n_1169), .Y (n_215));
INVX1 g68189(.A (g2227), .Y (n_259));
INVX1 g66956(.A (g9553), .Y (n_107));
INVX1 g67023(.A (g1632), .Y (n_105));
INVX1 g68148(.A (g1526), .Y (n_224));
INVX1 g67037(.A (g6035), .Y (n_103));
INVX1 g66998(.A (g2089), .Y (n_4183));
INVX1 g68130(.A (g2108), .Y (n_862));
INVX1 g68152(.A (g20763), .Y (n_101));
INVX1 g68220(.A (g1616), .Y (n_928));
INVX1 g68286(.A (g4392), .Y (n_596));
INVX1 g66932(.A (g2941), .Y (n_98));
INVX1 g68453(.A (n_662), .Y (n_404));
INVX1 g68458(.A (g1612), .Y (n_2521));
INVX1 g67791(.A (g1484), .Y (n_3383));
INVX1 g68237(.A (g1968), .Y (n_4946));
INVX1 g67844(.A (g_16063), .Y (n_3914));
INVX1 g67165(.A (n_4120), .Y (n_629));
INVX1 g67803(.A (g2437), .Y (n_1714));
INVX1 g67942(.A (g2193), .Y (n_96));
INVX1 g67950(.A (g3484), .Y (n_2699));
INVX1 g68421(.A (g1752), .Y (n_444));
INVX1 g68144(.A (g_10278), .Y (n_95));
INVX1 g67833(.A (g5481), .Y (n_94));
INVX1 g67743(.A (g4483), .Y (n_93));
INVX1 g67941(.A (g1736), .Y (n_1710));
INVX1 g67216(.A (g1236), .Y (n_92));
INVX1 g67836(.A (g2311), .Y (n_377));
INVX1 g66996(.A (g4486), .Y (n_89));
INVX1 g67982(.A (g_16769), .Y (n_2290));
INVX1 g66982(.A (g_9176), .Y (n_6057));
INVX1 g68112(.A (g1554), .Y (n_392));
INVX1 g68125(.A (g2273), .Y (n_6025));
INVX1 g67098(.A (g5752), .Y (n_87));
INVX1 g67080(.A (g_4449), .Y (n_284));
INVX1 g67120(.A (g_15879), .Y (n_86));
INVX1 g66954(.A (g_10715), .Y (n_2583));
INVX1 g67102(.A (g1840), .Y (n_854));
CLKBUFX1 g66944(.A (g4966), .Y (n_684));
INVX1 g66917(.A (g5495), .Y (n_1810));
INVX1 g67758(.A (g3827), .Y (n_85));
INVX1 g68412(.A (g3835), .Y (n_2692));
INVX1 g67145(.A (g_12465), .Y (n_287));
INVX1 g67997(.A (blif_reset_net), .Y (n_6421));
INVX1 g67153(.A (g4057), .Y (n_571));
INVX1 g67776(.A (g2575), .Y (n_933));
INVX1 g67750(.A (g_22464), .Y (n_83));
INVX1 g68417(.A (g2093), .Y (n_433));
INVX1 g67187(.A (g_16571), .Y (n_364));
INVX1 g67084(.A (g2675), .Y (n_6020));
INVX1 g68423(.A (g2433), .Y (n_1670));
INVX1 g67176(.A (g1886), .Y (n_291));
INVX1 g67928(.A (n_2429), .Y (n_453));
INVX1 g68224(.A (g1988), .Y (n_885));
INVX1 g67764(.A (g6187), .Y (n_2084));
INVX1 g68090(.A (g_15381), .Y (n_79));
INVX1 g67094(.A (g_22236), .Y (n_2529));
INVX1 g68322(.A (g1854), .Y (n_883));
INVX1 g66966(.A (g1874), .Y (n_1687));
INVX1 g67183(.A (g2514), .Y (n_4531));
INVX1 g66994(.A (g2465), .Y (n_3939));
INVX1 g67087(.A (g4116), .Y (n_282));
INVX1 g67986(.A (g1536), .Y (n_367));
INVX1 g68043(.A (g2652), .Y (n_418));
INVX1 g67754(.A (g2541), .Y (n_5969));
INVX1 g68132(.A (g1870), .Y (n_1705));
INVX1 g68181(.A (g4093), .Y (n_955));
INVX1 g67823(.A (g5909), .Y (n_75));
INVX1 g68081(.A (g2445), .Y (n_269));
INVX1 g67795(.A (g4417), .Y (n_74));
INVX1 g68099(.A (g1878), .Y (n_1706));
INVX1 g68381(.A (g3873), .Y (n_626));
INVX1 g68091(.A (g3106), .Y (n_3609));
INVX1 g68352(.A (g4311), .Y (n_327));
INVX1 g67788(.A (g2567), .Y (n_1505));
INVX1 g67040(.A (g3512), .Y (n_664));
INVX1 g67808(.A (g_22600), .Y (n_70));
INVX1 g65203(.A (g4688), .Y (n_69));
INVX1 g67142(.A (g1902), .Y (n_67));
INVX1 g68060(.A (g_18220), .Y (n_2556));
INVX1 g67119(.A (g3849), .Y (n_2923));
INVX1 g67900(.A (n_4139), .Y (n_446));
INVX1 g68163(.A (n_5996), .Y (n_804));
INVX1 g68077(.A (g5827), .Y (n_65));
INVX1 g67019(.A (n_5941), .Y (n_619));
INVX1 g68159(.A (g_20268), .Y (n_691));
INVX1 g67077(.A (g3333), .Y (n_64));
INVX1 g68314(.A (g_10556), .Y (n_447));
INVX1 g68372(.A (g2518), .Y (n_839));
INVX1 g68411(.A (g6227), .Y (n_617));
INVX1 g68135(.A (g2375), .Y (n_911));
INVX1 g67963(.A (g1772), .Y (n_3789));
INVX1 g67799(.A (g_3381), .Y (n_409));
INVX1 g68222(.A (g2509), .Y (n_904));
INVX1 g68292(.A (g3476), .Y (n_60));
INVX1 g67895(.A (g3401), .Y (n_59));
INVX1 g67978(.A (g2165), .Y (n_1518));
INVX1 g66947(.A (g_18200), .Y (n_2244));
INVX2 g68275(.A (g4983), .Y (n_598));
INVX1 g66929(.A (n_5917), .Y (n_730));
INVX1 g67196(.A (g2327), .Y (n_57));
INVX1 g68358(.A (g2441), .Y (n_2780));
INVX1 g67021(.A (g2393), .Y (n_4942));
INVX1 g67894(.A (g5180), .Y (n_482));
INVX1 g67860(.A (n_5932), .Y (n_674));
INVX1 g68256(.A (g2036), .Y (n_54));
INVX1 g67111(.A (g3179), .Y (n_553));
INVX1 g68294(.A (g2595), .Y (n_52));
INVX1 g67017(.A (g1936), .Y (n_328));
INVX1 g67774(.A (g1756), .Y (n_1666));
INVX1 g66967(.A (g2173), .Y (n_2258));
INVX1 g67190(.A (g1189), .Y (n_50));
INVX1 g67786(.A (g_16792), .Y (n_10496));
INVX1 g67141(.A (n_5925), .Y (n_806));
INVX1 g67146(.A (g1682), .Y (n_4893));
INVX1 g67979(.A (g1687), .Y (n_4527));
INVX1 g67761(.A (g1636), .Y (n_347));
INVX1 g67105(.A (g4628), .Y (n_46));
INVX1 g67745(.A (g1373), .Y (n_406));
INVX1 g68375(.A (g2265), .Y (n_864));
INVX1 g67160(.A (g_5342), .Y (n_6331));
INVX1 g68383(.A (g2547), .Y (n_858));
INVX1 g67800(.A (g_18590), .Y (n_6252));
INVX1 g68312(.A (g4054), .Y (n_3769));
INVX1 g68320(.A (g4176), .Y (n_43));
INVX1 g67162(.A (g2169), .Y (n_1529));
INVX1 g67188(.A (g3863), .Y (n_678));
INVX1 g68030(.A (g1974), .Y (n_871));
INVX1 g67178(.A (g_6283), .Y (n_40));
INVX1 g66931(.A (g3050), .Y (n_39));
INVX1 g68293(.A (g2848), .Y (n_38));
INVX1 g68264(.A (g_14587), .Y (n_35));
INVX1 g67820(.A (g4119), .Y (n_360));
INVX1 g66953(.A (g2902), .Y (n_3765));
INVX1 g68206(.A (n_1191), .Y (n_303));
INVX1 g67057(.A (g34026), .Y (n_986));
INVX1 g68176(.A (g4112), .Y (n_245));
INVX1 g67970(.A (g5011), .Y (n_843));
INVX1 g67118(.A (n_1177), .Y (n_388));
INVX1 g66990(.A (g2579), .Y (n_351));
INVX1 g67112(.A (g_15801), .Y (n_32));
INVX1 g68194(.A (g_12276), .Y (n_30));
INVX1 g68160(.A (g1724), .Y (n_29));
INVX1 g67822(.A (g1620), .Y (n_1510));
INVX1 g67946(.A (g_22639), .Y (n_28));
INVX1 g67868(.A (g2803), .Y (n_317));
INVX1 g68418(.A (g1821), .Y (n_4190));
INVX1 g67763(.A (g2999), .Y (n_27));
INVX1 g68347(.A (g1744), .Y (n_1711));
INVX1 g67782(.A (g1740), .Y (n_1665));
INVX1 g68026(.A (g1395), .Y (n_26));
INVX1 g68149(.A (g4122), .Y (n_3135));
INVX1 g67159(.A (g17607), .Y (n_371));
INVX1 g67851(.A (n_1135), .Y (n_370));
INVX1 g67193(.A (n_1356), .Y (n_379));
INVX1 g67794(.A (g2259), .Y (n_5961));
INVX1 g68155(.A (g4621), .Y (n_23));
INVX1 g67741(.A (g_15740), .Y (n_708));
INVX1 g66972(.A (g1890), .Y (n_1688));
INVX1 g66961(.A (g23002), .Y (n_22));
INVX1 g67206(.A (g1361), .Y (n_297));
INVX1 g67883(.A (g4349), .Y (n_221));
INVX1 g67062(.A (g2102), .Y (n_5953));
CLKBUFX1 g67887(.A (g_4409), .Y (g12238));
INVX1 g67214(.A (g_13838), .Y (n_21));
INVX1 g68402(.A (g4821), .Y (n_20));
INVX1 g68258(.A (g4826), .Y (n_19));
INVX1 g68376(.A (g4831), .Y (n_1299));
INVX1 g68457(.A (g2307), .Y (n_2293));
INVX1 g67757(.A (g21292), .Y (g23612));
INVX1 g68414(.A (g2241), .Y (n_916));
INVX1 g67138(.A (g1913), .Y (n_17));
INVX1 g66910(.A (g1413), .Y (n_16));
INVX1 g67004(.A (g4489), .Y (n_13));
INVX1 g68107(.A (g2161), .Y (n_1528));
INVX1 g67804(.A (g1955), .Y (n_4187));
INVX1 g67926(.A (g2461), .Y (n_12));
INVX1 g67826(.A (g2735), .Y (n_11));
INVX1 g68059(.A (g5689), .Y (n_401));
INVX1 g67918(.A (g2661), .Y (n_5958));
INVX1 g67988(.A (g_5450), .Y (n_2566));
INVX1 g67772(.A (g4332), .Y (n_448));
INVX1 g65604(.A (g34028), .Y (n_987));
INVX2 g67036(.A (g6035), .Y (n_423));
INVX1 g68097(.A (g5489), .Y (n_3011));
INVX1 g67837(.A (g1748), .Y (n_2550));
INVX1 g68133(.A (g2283), .Y (n_5));
INVX1 g68136(.A (g6533), .Y (n_1794));
INVX1 g67055(.A (g5841), .Y (n_1807));
INVX1 g67003(.A (n_1216), .Y (n_261));
INVX1 g67996(.A (n_1210), .Y (n_365));
INVX1 g67024(.A (g5142), .Y (n_2718));
INVX1 g68139(.A (g4064), .Y (n_572));
INVX1 g68128(.A (g1700), .Y (n_5964));
INVX1 g68242(.A (g1384), .Y (n_2));
INVX1 g68299(.A (g6444), .Y (n_1));
INVX1 g67173(.A (g3125), .Y (n_0));
INVX1 g68443(.A (g5148), .Y (n_1813));
INVX1 g68032(.A (g6336), .Y (n_609));
INVX1 g68062(.A (g1825), .Y (n_827));
CLKBUFX1 g68446(.A (g_6165), .Y (g12422));
INVX1 g69642(.A (n_10306), .Y (n_6454));
INVX1 g69644(.A (n_6715), .Y (n_6457));
INVX1 g69646(.A (n_6464), .Y (n_6460));
INVX1 g69652(.A (n_6621), .Y (n_6468));
NOR2X1 g53(.A (n_6503), .B (n_10307), .Y (n_6479));
NAND3X1 g49(.A (n_6464), .B (n_6488), .C (n_6501), .Y (n_3661));
NOR2X1 g54(.A (n_10637), .B (n_7275), .Y (n_6464));
NOR2X1 g69656(.A (g_8896), .B (n_6552), .Y (n_6488));
NAND2X1 g69658(.A (n_10814), .B (n_10529), .Y (n_6490));
INVX1 g69664(.A (n_6490), .Y (n_6501));
OAI21X1 g41(.A0 (n_10313), .A1 (n_6504), .B0 (n_6507), .Y (n_6508));
NAND2X1 g69666(.A (n_9698), .B (n_6503), .Y (n_6504));
INVX1 g47(.A (g_9338), .Y (n_6503));
AOI21X1 g42(.A0 (n_7229), .A1 (n_10313), .B0 (n_6506), .Y (n_6507));
AND2X1 g69667(.A (n_7402), .B (g_9338), .Y (n_7229));
NOR2X1 g69668(.A (n_519), .B (n_9698), .Y (n_6506));
NAND2X1 g69670(.A (n_8793), .B (g_13871), .Y (n_6517));
OR2X1 g31(.A (n_6522), .B (n_6523), .Y (n_6524));
OR2X1 g34(.A (n_10311), .B (n_8792), .Y (n_6522));
NAND2X1 g32(.A (n_6610), .B (n_10863), .Y (n_6523));
INVX1 g12(.A (g_22021), .Y (n_6527));
OAI21X1 g69673(.A0 (g_21806), .A1 (g_22379), .B0 (n_11095), .Y(n_10142));
NAND2X1 g69676(.A (n_11094), .B (g_21806), .Y (n_6539));
AND2X1 g69677(.A (n_6548), .B (g_12922), .Y (n_11105));
INVX1 g26(.A (n_6547), .Y (n_6548));
NAND3X1 g21(.A (n_11120), .B (n_10494), .C (n_6690), .Y (n_6547));
NOR2X1 g24(.A (n_2566), .B (n_6545), .Y (n_10494));
NAND2X1 g25(.A (n_11064), .B (g_19659), .Y (n_6545));
CLKBUFX1 g69681(.A (n_6548), .Y (n_6549));
NOR2X1 g22(.A (n_2566), .B (n_7145), .Y (n_6551));
NOR2X1 g69685(.A (g_8896), .B (n_6552), .Y (n_6553));
NAND2X2 g69686(.A (n_417), .B (n_223), .Y (n_6552));
INVX1 g69693(.A (n_6800), .Y (n_6562));
NOR2X1 g69697(.A (n_447), .B (n_10309), .Y (n_6564));
NAND2X1 g69698(.A (n_7097), .B (g12184), .Y (n_6565));
NAND2X1 g23(.A (n_6565), .B (n_11118), .Y (n_6570));
NAND4X1 g69702(.A (n_6572), .B (n_7260), .C (n_662), .D (g4332), .Y(n_6574));
AND2X1 g69703(.A (g4349), .B (n_1627), .Y (n_6572));
NAND2X1 g69706(.A (n_6572), .B (n_7260), .Y (n_6578));
NOR2X1 g69707(.A (n_10402), .B (n_46), .Y (n_6582));
INVX1 g69713(.A (g1478), .Y (n_6584));
INVX1 g69730(.A (n_8546), .Y (n_6610));
NOR2X1 g69733(.A (g_20909), .B (n_5712), .Y (n_6612));
NOR2X1 g69734(.A (g_17086), .B (n_10311), .Y (n_6618));
AND2X1 g69740(.A (n_6618), .B (n_6620), .Y (n_6621));
NOR2X1 g69741(.A (n_5712), .B (n_8819), .Y (n_6620));
INVX1 g69742(.A (g_17086), .Y (n_6308));
AOI21X1 g69743(.A0 (n_6937), .A1 (n_6938), .B0 (n_9836), .Y (n_6631));
OR2X1 g69744(.A (n_4339), .B (n_4168), .Y (n_6938));
NAND2X1 g29(.A (n_10852), .B (g2421), .Y (n_6937));
AOI21X1 g69750(.A0 (n_6940), .A1 (n_6941), .B0 (n_9775), .Y (n_6639));
OR2X1 g69751(.A (g2361), .B (n_4169), .Y (n_6941));
NAND2X1 g69752(.A (n_10670), .B (g2287), .Y (n_6940));
NOR2X1 g18(.A (n_10264), .B (n_6801), .Y (n_6655));
INVX1 g69772(.A (n_6663), .Y (n_6664));
NAND2X1 g69773(.A (n_10981), .B (n_9453), .Y (n_6663));
INVX2 g69782(.A (n_10976), .Y (n_6666));
AOI21X1 g69786(.A0 (n_6668), .A1 (n_11097), .B0 (n_6669), .Y(n_6670));
NOR2X1 g69787(.A (g2704), .B (g2697), .Y (n_6668));
NOR2X1 g69788(.A (g1291), .B (n_6584), .Y (n_6669));
INVX1 g69790(.A (n_6669), .Y (n_6673));
INVX1 g69791(.A (n_6683), .Y (n_6684));
NAND2X1 g69792(.A (n_6680), .B (n_9717), .Y (n_6683));
OAI21X1 g69793(.A0 (n_3998), .A1 (g1936), .B0 (n_6679), .Y (n_6680));
NAND2X1 g69794(.A (n_6685), .B (g1862), .Y (n_6679));
CLKBUFX3 g69796(.A (n_6676), .Y (n_6677));
CLKBUFX3 g69797(.A (n_6789), .Y (n_6676));
INVX2 g69801(.A (n_6677), .Y (n_6685));
OAI21X1 g69802(.A0 (n_6687), .A1 (n_1183), .B0 (n_6689), .Y (n_6690));
OR4X1 g39(.A (g_22371), .B (g_13838), .C (n_70), .D (n_6923), .Y(n_6687));
NAND3X1 g40(.A (n_10566), .B (n_876), .C (n_6688), .Y (n_6689));
AND2X1 g69803(.A (g_22371), .B (g_13838), .Y (n_6688));
AOI21X1 g69804(.A0 (n_6692), .A1 (n_6693), .B0 (g_13838), .Y(n_6694));
NOR2X1 g69805(.A (n_6923), .B (n_6691), .Y (n_6692));
OR2X1 g69806(.A (g_22371), .B (n_70), .Y (n_6691));
INVX1 g69807(.A (n_1183), .Y (n_6693));
NAND3X1 g69808(.A (n_10566), .B (n_876), .C (g_22371), .Y (n_6695));
NOR2X1 g69812(.A (g2138), .B (g2145), .Y (n_6696));
NAND2X1 g69814(.A (n_10557), .B (g_11413), .Y (n_6697));
INVX1 g69818(.A (n_8846), .Y (n_6705));
CLKBUFX1 g3(.A (n_10678), .Y (n_6707));
NOR2X1 g69826(.A (n_6714), .B (n_6715), .Y (n_6716));
INVX1 g69827(.A (n_7043), .Y (n_6714));
NAND2X1 g69828(.A (n_7042), .B (n_10863), .Y (n_6715));
NAND2X1 g69838(.A (n_10399), .B (n_10401), .Y (n_6577));
NOR2X1 g69843(.A (n_3459), .B (n_6734), .Y (n_6735));
NOR2X1 g69845(.A (g1345), .B (n_10430), .Y (n_6734));
NOR3X1 g69852(.A (g2629), .B (n_6742), .C (n_6666), .Y (n_6746));
INVX1 g69853(.A (g2599), .Y (n_6742));
NOR2X1 g69858(.A (n_9019), .B (n_6756), .Y (n_6757));
AOI21X1 g69860(.A0 (n_6754), .A1 (g1996), .B0 (n_6755), .Y (n_6756));
CLKBUFX1 g69861(.A (n_6752), .Y (n_6754));
INVX1 g69863(.A (n_7099), .Y (n_6752));
NOR2X1 g69867(.A (g2070), .B (n_4516), .Y (n_6755));
INVX1 g69868(.A (n_6752), .Y (n_6758));
CLKBUFX1 g69869(.A (n_7099), .Y (n_6759));
NAND2X1 g69870(.A (n_6762), .B (n_10553), .Y (n_11081));
NAND4X1 g69871(.A (n_2451), .B (n_2452), .C (n_2150), .D (n_6760), .Y(n_10553));
NAND2X1 g69872(.A (g_19911), .B (g_16958), .Y (n_6760));
OR2X1 g69873(.A (n_10123), .B (g_15287), .Y (n_6762));
NOR2X1 g69874(.A (n_6764), .B (n_6766), .Y (n_6767));
INVX1 g69875(.A (n_6762), .Y (n_6764));
NOR2X1 g69876(.A (g_19911), .B (n_6765), .Y (n_6766));
NAND3X1 g69877(.A (n_2451), .B (n_2452), .C (n_2150), .Y (n_6765));
INVX1 g69888(.A (n_10803), .Y (n_6781));
CLKBUFX1 g15(.A (n_10801), .Y (n_6782));
CLKBUFX3 g69889(.A (n_6786), .Y (n_6787));
NOR2X1 g69890(.A (g4054), .B (n_6785), .Y (n_6786));
INVX1 g69891(.A (g3990), .Y (n_6785));
NAND2X1 g69892(.A (n_6789), .B (n_6790), .Y (n_6791));
NAND3X1 g69893(.A (n_898), .B (n_6788), .C (n_10986), .Y (n_6789));
OAI21X1 g69894(.A0 (n_698), .A1 (n_10829), .B0 (g17400), .Y (n_6788));
NOR2X1 g69895(.A (g1862), .B (g1936), .Y (n_6790));
AND2X1 g69897(.A (g3990), .B (g4054), .Y (n_8917));
AND2X1 g69898(.A (n_10495), .B (n_10261), .Y (n_6798));
NOR2X1 g69899(.A (g_18590), .B (n_6796), .Y (n_10495));
NAND3X1 g69900(.A (n_6794), .B (n_10142), .C (n_6057), .Y (n_6796));
AND2X1 g69901(.A (n_11120), .B (n_10628), .Y (n_6794));
NAND2X1 g19(.A (n_10261), .B (n_6799), .Y (n_6800));
INVX1 g69903(.A (n_6796), .Y (n_6799));
NAND2X1 g69904(.A (n_6794), .B (n_10142), .Y (n_6801));
NAND4X1 g69909(.A (n_6806), .B (n_6808), .C (g3945), .D (g16775), .Y(n_6809));
OAI21X1 g69910(.A0 (n_690), .A1 (g_3974), .B0 (n_802), .Y (n_6806));
NOR2X1 g69911(.A (g3990), .B (n_6807), .Y (n_6808));
INVX1 g69912(.A (g4054), .Y (n_6807));
NAND2X1 g63(.A (n_6821), .B (n_6822), .Y (n_6823));
NOR2X1 g66(.A (n_3764), .B (n_7168), .Y (n_6821));
INVX1 g67(.A (n_7354), .Y (n_6822));
OAI21X1 g69938(.A0 (n_6854), .A1 (n_6856), .B0 (n_6857), .Y (n_6858));
AOI21X1 g69939(.A0 (n_6848), .A1 (n_6849), .B0 (n_6853), .Y (n_6854));
INVX1 g69940(.A (n_4969), .Y (n_6848));
NOR2X1 g69941(.A (n_10271), .B (n_5471), .Y (n_6849));
OAI21X1 g69942(.A0 (n_6850), .A1 (n_6851), .B0 (n_6852), .Y (n_6853));
OR2X1 g50(.A (n_4968), .B (n_5471), .Y (n_6850));
CLKBUFX1 g69943(.A (n_4582), .Y (n_6851));
NAND2X1 g69944(.A (n_9693), .B (n_4120), .Y (n_6852));
AND2X1 g69945(.A (n_6852), .B (n_9129), .Y (n_6856));
NAND3X1 g69947(.A (n_5471), .B (n_9553), .C (n_4893), .Y (n_6857));
NOR2X1 g69949(.A (n_9019), .B (n_6865), .Y (n_6866));
AOI21X1 g69951(.A0 (n_10910), .A1 (g1728), .B0 (n_6864), .Y (n_6865));
NOR2X1 g69955(.A (n_4139), .B (n_4006), .Y (n_6864));
OAI21X1 g37(.A0 (n_8882), .A1 (n_8883), .B0 (n_6877), .Y (n_6878));
NAND3X1 g69961(.A (n_6872), .B (n_11207), .C (n_9359), .Y (n_8882));
NAND2X1 g69962(.A (n_6049), .B (n_6095), .Y (n_6872));
AOI22X1 g69965(.A0 (g3813), .A1 (n_9193), .B0 (n_9883), .B1 (n_6876),.Y (n_6877));
AND2X1 g69966(.A (n_6243), .B (n_3596), .Y (n_6876));
NAND2X1 g69970(.A (n_6696), .B (g2130), .Y (n_6880));
INVX2 g69974(.A (n_6891), .Y (n_6892));
INVX2 g7(.A (n_10609), .Y (n_6891));
INVX1 g69978(.A (n_6891), .Y (n_6893));
INVX2 g69980(.A (n_6891), .Y (n_6895));
NOR2X1 g69981(.A (n_10841), .B (n_6896), .Y (n_6897));
INVX1 g69982(.A (n_10607), .Y (n_6896));
NOR2X1 g69984(.A (n_6899), .B (n_6906), .Y (n_6907));
NAND2X1 g69985(.A (n_6553), .B (n_6898), .Y (n_6899));
NAND2X1 g69986(.A (n_584), .B (n_10108), .Y (n_6898));
NAND3X1 g69987(.A (n_6903), .B (n_10805), .C (n_10569), .Y (n_6906));
NOR2X1 g69988(.A (n_10637), .B (n_10639), .Y (n_6903));
NAND2X1 g6(.A (n_6922), .B (g_20208), .Y (n_6923));
INVX1 g70007(.A (g_21813), .Y (n_6922));
AOI21X1 g70008(.A0 (n_6925), .A1 (n_7144), .B0 (n_6926), .Y (n_6927));
AND2X1 g70009(.A (n_9521), .B (g_22605), .Y (n_6925));
NOR2X1 g70010(.A (n_9717), .B (g_22070), .Y (n_6926));
INVX1 g70011(.A (g_22070), .Y (n_6928));
AND2X1 g70021(.A (n_10936), .B (n_11034), .Y (n_6951));
AOI21X1 g70022(.A0 (n_3832), .A1 (g1242), .B0 (n_3831), .Y (n_6953));
AOI21X1 g61508_dup(.A0 (n_3832), .A1 (g1242), .B0 (n_3831), .Y(n_6954));
NOR2X1 g70023(.A (n_6823), .B (n_10974), .Y (n_7235));
NOR2X1 g59_dup(.A (n_10974), .B (n_6823), .Y (n_6956));
INVX1 g70025(.A (n_10708), .Y (n_6958));
CLKBUFX1 g70036(.A (n_6973), .Y (n_6972));
CLKBUFX1 g70039(.A (n_6979), .Y (n_6978));
CLKBUFX1 g70059(.A (n_7004), .Y (n_7003));
OR2X1 g70070(.A (g5046), .B (n_10768), .Y (n_7018));
NAND2X2 g70071(.A (n_7023), .B (n_7024), .Y (n_7025));
INVX1 g70072(.A (n_7022), .Y (n_7023));
NOR2X1 g29_dup(.A (n_10461), .B (n_8759), .Y (n_7022));
NAND3X1 g70075(.A (n_10827), .B (n_8832), .C (n_8796), .Y (n_8756));
NOR2X1 g70076(.A (g1728), .B (n_4139), .Y (n_7024));
INVX1 g71(.A (g_10903), .Y (n_7032));
NAND4X1 g70085(.A (n_7039), .B (n_7116), .C (n_8690), .D (n_10638),.Y (n_7040));
INVX1 g70086(.A (n_8691), .Y (n_7039));
NOR2X1 g70087(.A (n_8546), .B (n_7105), .Y (n_7042));
NOR2X1 g70(.A (n_153), .B (n_10311), .Y (n_7043));
NOR2X1 g70090(.A (n_7045), .B (n_7046), .Y (n_7047));
NAND3X1 g70091(.A (n_10577), .B (n_3740), .C (n_7044), .Y (n_7045));
NAND4X1 g70092(.A (n_10883), .B (n_10576), .C (g3590), .D (g13881),.Y (n_7044));
NAND4X1 g70093(.A (n_4107), .B (n_4683), .C (n_3542), .D (n_4996), .Y(n_7046));
AND2X1 g70094(.A (n_3761), .B (n_3541), .Y (n_7048));
AND2X1 g70095(.A (n_2652), .B (n_4101), .Y (n_7049));
XOR2X1 g70129(.A (n_7085), .B (n_11197), .Y (n_7093));
NOR2X1 g70130(.A (n_10443), .B (n_332), .Y (n_7085));
NOR2X1 g70132(.A (n_7086), .B (n_7087), .Y (n_7088));
NAND4X1 g70133(.A (n_2379), .B (n_2324), .C (n_2343), .D (n_2971), .Y(n_7086));
NAND4X1 g70134(.A (n_2326), .B (n_2659), .C (n_2130), .D (n_2414), .Y(n_7087));
NAND2X1 g70136(.A (n_2353), .B (n_2342), .Y (n_7089));
NAND4X1 g70137(.A (n_2141), .B (n_2030), .C (n_2132), .D (n_3267), .Y(n_7090));
INVX1 g70140(.A (g_15127), .Y (n_7094));
INVX1 g8(.A (g_17653), .Y (n_7097));
NAND2X2 g70141(.A (n_7099), .B (n_7101), .Y (n_7102));
NAND3X1 g70143(.A (n_8880), .B (n_1133), .C (n_2670), .Y (n_7099));
NAND2X1 g70144(.A (n_1709), .B (g_18330), .Y (n_8880));
NOR2X1 g70145(.A (g1996), .B (g2070), .Y (n_7101));
NAND2X1 g70146(.A (n_2670), .B (n_1133), .Y (n_7103));
OR2X1 g70150(.A (n_6517), .B (n_10309), .Y (n_7105));
AND2X1 g70159(.A (n_10569), .B (n_10805), .Y (n_7116));
NOR2X1 g70160(.A (n_10177), .B (n_10176), .Y (n_8909));
NAND3X1 g58(.A (n_7047), .B (n_7048), .C (n_7049), .Y (n_10176));
NAND3X1 g70161(.A (n_7119), .B (n_7120), .C (n_7124), .Y (n_10177));
INVX1 g59(.A (n_7118), .Y (n_7119));
NAND4X1 g70162(.A (n_2140), .B (n_1691), .C (n_5500), .D (n_1850), .Y(n_7118));
AND2X1 g70163(.A (n_2146), .B (n_2138), .Y (n_7120));
AOI21X1 g70164(.A0 (n_11126), .A1 (n_7122), .B0 (n_7123), .Y(n_7124));
INVX1 g70165(.A (n_7121), .Y (n_7122));
NAND3X1 g57(.A (n_10883), .B (g16722), .C (g3606), .Y (n_7121));
NAND2X1 g70166(.A (n_1587), .B (n_5425), .Y (n_7123));
NAND3X1 g70167(.A (n_7130), .B (n_7131), .C (n_7132), .Y (n_7133));
NAND3X1 g70168(.A (n_7127), .B (n_7128), .C (n_9558), .Y (n_7130));
INVX1 g70169(.A (n_6248), .Y (n_7127));
OAI22X1 g70170(.A0 (n_3779), .A1 (n_8909), .B0 (n_3779), .B1(n_6052), .Y (n_7128));
NAND2X1 g70172(.A (n_9300), .B (g3462), .Y (n_7131));
NAND3X1 g70173(.A (n_3779), .B (n_9139), .C (n_3601), .Y (n_7132));
AND2X1 g70179(.A (n_11105), .B (n_7143), .Y (n_7144));
NOR2X1 g70180(.A (n_7140), .B (n_7142), .Y (n_7143));
NAND3X1 g70181(.A (n_11055), .B (n_6928), .C (g_18308), .Y (n_7140));
INVX1 g70182(.A (n_7141), .Y (n_7142));
AND2X1 g70183(.A (n_6690), .B (n_11120), .Y (n_7141));
NAND2X1 g70184(.A (n_7141), .B (n_11055), .Y (n_7145));
AND2X1 g70185(.A (n_11105), .B (g_18308), .Y (n_7146));
NOR2X1 g70187(.A (n_10660), .B (n_191), .Y (n_7150));
NAND4X1 g70199(.A (n_8589), .B (n_7164), .C (n_7165), .D (n_7167), .Y(n_7168));
NAND4X1 g70201(.A (n_10941), .B (n_8588), .C (g16686), .D (g3247), .Y(n_7164));
NAND4X1 g70205(.A (n_11029), .B (n_8588), .C (g3187), .D (g14421), .Y(n_7165));
NAND4X1 g70206(.A (n_8572), .B (n_8588), .C (g3215), .D (g16874), .Y(n_7167));
AND2X1 g75(.A (n_2441), .B (n_2354), .Y (n_7208));
NAND3X1 g70249(.A (n_2966), .B (n_2327), .C (n_2336), .Y (n_7213));
NAND3X1 g72(.A (n_2598), .B (n_1293), .C (n_2149), .Y (n_7214));
NOR2X1 g70250(.A (n_356), .B (n_10341), .Y (n_7217));
NOR2X1 g70251(.A (n_7217), .B (n_7218), .Y (n_7219));
NAND4X1 g67_dup(.A (n_10238), .B (n_10239), .C (n_10240), .D(n_10241), .Y (n_7218));
INVX2 g70266(.A (n_7245), .Y (n_7242));
INVX1 g70267(.A (n_7245), .Y (n_7243));
INVX2 g70269(.A (n_3829), .Y (n_7245));
NOR2X1 g70292(.A (n_7032), .B (n_153), .Y (n_7268));
INVX1 g70296(.A (n_10569), .Y (n_7275));
AOI22X1 g70339(.A0 (n_7330), .A1 (n_7332), .B0 (n_7329), .B1(n_7331), .Y (n_7333));
INVX1 g70340(.A (n_7329), .Y (n_7330));
NAND4X1 g70341(.A (n_7322), .B (n_7325), .C (n_7328), .D (n_3693), .Y(n_7329));
NOR2X1 g70342(.A (n_7320), .B (n_7321), .Y (n_7322));
NAND4X1 g70343(.A (n_2436), .B (n_2334), .C (n_2323), .D (n_2349), .Y(n_7320));
NAND3X1 g70344(.A (n_3265), .B (n_2434), .C (n_2431), .Y (n_7321));
INVX1 g70345(.A (n_7324), .Y (n_7325));
NAND3X1 g70346(.A (n_2601), .B (n_7323), .C (n_3276), .Y (n_7324));
AND2X1 g78(.A (n_1292), .B (n_2148), .Y (n_7323));
NOR2X1 g70347(.A (n_7326), .B (n_7327), .Y (n_7328));
NAND2X1 g70348(.A (n_2388), .B (n_2964), .Y (n_7326));
NAND2X1 g77(.A (n_2338), .B (n_2321), .Y (n_7327));
INVX1 g70349(.A (n_7331), .Y (n_7332));
NOR2X1 g70350(.A (n_247), .B (n_2039), .Y (n_7331));
NAND3X1 g70360(.A (n_7343), .B (n_7344), .C (n_7353), .Y (n_7354));
NAND4X1 g70361(.A (n_1499), .B (n_10941), .C (g3235), .D (g16718), .Y(n_7343));
NAND4X1 g70362(.A (n_1499), .B (n_8586), .C (g3219), .D (g13895), .Y(n_7344));
AND2X1 g70363(.A (n_7348), .B (n_7352), .Y (n_7353));
NAND4X1 g70364(.A (n_11030), .B (n_8588), .C (g3195), .D (g3329), .Y(n_7348));
NAND4X1 g70368(.A (n_8572), .B (n_8588), .C (g_4050), .D (g3191), .Y(n_7352));
INVX4 g70397(.A (n_8588), .Y (n_7383));
CLKBUFX3 g70409(.A (n_7402), .Y (n_7395));
CLKBUFX1 g71109(.A (n_8509), .Y (n_8508));
NAND2X1 g71126(.A (n_10379), .B (n_8534), .Y (n_10101));
OAI21X1 g71130(.A0 (n_1180), .A1 (n_2108), .B0 (g17320), .Y (n_8532));
NOR2X1 g71131(.A (g2153), .B (g2227), .Y (n_8534));
NAND2X2 g71132(.A (n_8864), .B (n_8537), .Y (n_10829));
NOR2X1 g71134(.A (n_10129), .B (n_8800), .Y (n_8537));
NAND3X1 g71137(.A (n_10308), .B (n_7268), .C (n_10806), .Y (n_8540));
NAND2X1 g71139(.A (n_10308), .B (g_16296), .Y (n_8546));
NAND4X1 g71140(.A (n_8548), .B (n_8572), .C (g3243), .D (g16718), .Y(n_8552));
NAND2X2 g71141(.A (n_800), .B (n_8547), .Y (n_8548));
OR2X1 g71142(.A (g_4050), .B (n_8587), .Y (n_8547));
INVX2 g71148(.A (n_8556), .Y (n_8557));
INVX1 g71149(.A (n_8555), .Y (n_8556));
NOR2X1 g71150(.A (g2724), .B (n_10656), .Y (n_8555));
INVX2 g71164(.A (n_8571), .Y (n_8572));
NAND2X1 g71165(.A (n_10839), .B (n_7004), .Y (n_8571));
INVX1 g71172(.A (n_8582), .Y (n_8583));
NAND4X1 g71173(.A (n_10262), .B (n_10263), .C (n_11119), .D(n_10142), .Y (n_8582));
NAND4X1 g71175(.A (n_8586), .B (n_8588), .C (g3231), .D (g13865), .Y(n_8589));
INVX2 g71176(.A (n_8585), .Y (n_8586));
NAND2X1 g71177(.A (n_8584), .B (n_10834), .Y (n_8585));
INVX1 g71178(.A (n_7004), .Y (n_8584));
INVX2 g71179(.A (n_8587), .Y (n_8588));
INVX2 g71180(.A (g3338), .Y (n_8587));
NOR2X1 g71181(.A (n_8770), .B (g1183), .Y (n_8591));
INVX2 g71186(.A (g_13091), .Y (n_8594));
NAND2X1 g71190(.A (n_8601), .B (n_8604), .Y (n_8605));
NAND3X1 g71191(.A (n_8599), .B (n_8600), .C (n_9453), .Y (n_8601));
OAI22X1 g71192(.A0 (n_3775), .A1 (n_7235), .B0 (n_3775), .B1(n_6051), .Y (n_8599));
INVX1 g71193(.A (n_6250), .Y (n_8600));
AOI22X1 g71194(.A0 (g3111), .A1 (n_9772), .B0 (n_3775), .B1 (n_8603),.Y (n_8604));
AND2X1 g43(.A (n_10385), .B (n_3609), .Y (n_8603));
NAND2X2 g71198(.A (n_8615), .B (n_8619), .Y (n_8620));
NAND2X1 g71199(.A (n_8611), .B (n_9717), .Y (n_8615));
INVX1 g71200(.A (n_8610), .Y (n_8611));
AOI21X1 g71201(.A0 (n_8768), .A1 (n_3855), .B0 (n_8609), .Y (n_8610));
AND2X1 g71203(.A (g7916), .B (n_8591), .Y (n_8609));
NAND2X2 g71207(.A (n_8616), .B (n_8618), .Y (n_8619));
OR2X1 g71208(.A (n_9466), .B (n_8768), .Y (n_8616));
NAND3X1 g71209(.A (n_3854), .B (n_3841), .C (n_10005), .Y (n_8618));
NAND2X2 g71214(.A (n_10937), .B (n_8627), .Y (n_8628));
NOR2X1 g71217(.A (g2287), .B (g2361), .Y (n_8627));
AND2X1 g71218(.A (n_10936), .B (n_11034), .Y (n_8629));
NAND2X2 g71219(.A (n_10961), .B (n_8632), .Y (n_8633));
NOR2X1 g71222(.A (g2421), .B (n_4339), .Y (n_8632));
AND2X1 g71223(.A (n_10960), .B (n_11035), .Y (n_8634));
INVX2 g71224(.A (n_8638), .Y (n_8639));
NAND2X1 g71225(.A (n_11210), .B (n_8637), .Y (n_8638));
INVX2 g71228(.A (g4793), .Y (n_8637));
NAND2X1 g71255(.A (n_6880), .B (n_10316), .Y (n_10173));
NOR2X1 g71257(.A (n_10228), .B (n_10175), .Y (n_8810));
INVX2 g71261(.A (n_8675), .Y (n_8676));
NAND3X1 g71262(.A (n_10192), .B (g4966), .C (n_598), .Y (n_8675));
AND2X1 g71265(.A (n_10192), .B (g4966), .Y (n_8677));
NOR2X1 g71267(.A (n_8678), .B (n_7105), .Y (n_8679));
NAND3X1 g71268(.A (n_10638), .B (n_10569), .C (g_16296), .Y (n_8678));
INVX1 g71269(.A (n_8681), .Y (n_8682));
NAND2X1 g71270(.A (n_8680), .B (n_6564), .Y (n_8681));
AND2X1 g56_dup(.A (n_6565), .B (n_6898), .Y (n_8680));
NOR2X1 g71271(.A (n_8686), .B (n_8540), .Y (n_8687));
NAND2X1 g71272(.A (n_6553), .B (n_10308), .Y (n_8686));
AND2X1 g71277(.A (n_6565), .B (n_6898), .Y (n_8690));
NAND2X1 g71278(.A (n_6564), .B (n_6553), .Y (n_8691));
CLKBUFX1 g71279(.A (n_8693), .Y (n_8694));
NOR2X1 g71280(.A (g4785), .B (n_10225), .Y (n_8693));
OAI21X1 g71284(.A0 (n_8702), .A1 (n_8703), .B0 (n_8705), .Y (n_8706));
NAND3X1 g71285(.A (n_8697), .B (g28753), .C (n_9521), .Y (n_8702));
OR2X1 g71286(.A (n_10684), .B (n_2078), .Y (n_8697));
AND2X1 g71289(.A (n_2078), .B (n_10684), .Y (n_8703));
AOI22X1 g71290(.A0 (g5120), .A1 (n_9454), .B0 (n_8704), .B1 (n_3244),.Y (n_8705));
AND2X1 g71291(.A (n_9698), .B (n_3618), .Y (n_8704));
INVX1 g45(.A (g28753), .Y (n_8707));
NAND2X1 g71314(.A (n_8731), .B (n_8735), .Y (n_8736));
INVX1 g71315(.A (n_8730), .Y (n_8731));
NAND4X1 g71316(.A (n_11194), .B (n_1575), .C (n_11195), .D (n_1855),.Y (n_8730));
INVX1 g71317(.A (n_8734), .Y (n_8735));
NAND4X1 g71318(.A (n_3286), .B (n_10368), .C (n_8733), .D (n_1859),.Y (n_8734));
NAND4X1 g71320(.A (n_2339), .B (n_1695), .C (g5264), .D (g17639), .Y(n_8733));
NOR2X1 g71335(.A (n_262), .B (n_8885), .Y (n_8757));
NOR2X1 g62211_dup(.A (n_262), .B (n_8886), .Y (n_8758));
AND2X1 g71336(.A (g17316), .B (n_8756), .Y (n_8759));
AOI21X1 g71337(.A0 (n_6951), .A1 (g1585), .B0 (n_3873), .Y (n_8761));
AOI21X1 g61378_dup(.A0 (n_6951), .A1 (g1585), .B0 (n_3873), .Y(n_8762));
AOI21X1 g71338(.A0 (n_11211), .A1 (n_10764), .B0 (n_3870), .Y(n_8763));
AOI21X1 g61379_dup(.A0 (n_11212), .A1 (n_10764), .B0 (n_3870), .Y(n_8764));
CLKBUFX1 g71342(.A (n_8769), .Y (n_8768));
INVX2 g71343(.A (n_8770), .Y (n_8769));
INVX2 g71344(.A (g1171), .Y (n_8770));
INVX1 g71349(.A (n_8777), .Y (n_8776));
CLKBUFX3 g71350(.A (n_8778), .Y (n_8777));
INVX1 g71363(.A (n_8793), .Y (n_8792));
CLKBUFX1 g71368(.A (n_8800), .Y (n_8799));
CLKBUFX1 g71372(.A (n_8807), .Y (n_8806));
CLKBUFX1 g71374(.A (n_8810), .Y (n_8809));
NAND4X1 g71375(.A (n_8679), .B (n_8682), .C (n_8687), .D (n_8818), .Y(n_8819));
NOR2X1 g71376(.A (n_8816), .B (n_8817), .Y (n_8818));
NAND2X1 g71377(.A (n_10310), .B (g_21799), .Y (n_8816));
OR2X1 g71382(.A (n_86), .B (n_10309), .Y (n_8817));
OR2X1 g71384(.A (n_8817), .B (n_8820), .Y (n_8821));
NAND3X1 g71385(.A (n_8679), .B (n_8682), .C (n_8687), .Y (n_8820));
NOR2X1 g71394(.A (g7916), .B (n_8835), .Y (n_8836));
NAND2X2 g71395(.A (n_8831), .B (n_8834), .Y (n_8835));
NAND2X2 g71396(.A (n_1833), .B (n_1255), .Y (n_8831));
AOI21X1 g71397(.A0 (n_8833), .A1 (n_10647), .B0 (n_1636), .Y(n_8834));
INVX1 g71398(.A (n_8832), .Y (n_8833));
AND2X1 g71399(.A (g1183), .B (n_8770), .Y (n_8832));
INVX1 g71400(.A (g7916), .Y (n_8837));
NOR2X1 g71402(.A (n_1636), .B (n_8839), .Y (n_8840));
INVX1 g71403(.A (n_8831), .Y (n_8839));
AND2X1 g71409(.A (n_10724), .B (n_10647), .Y (n_8846));
NAND2X1 g71414(.A (n_8848), .B (n_10286), .Y (n_8850));
NAND2X1 g71415(.A (n_10956), .B (g1300), .Y (n_8848));
INVX1 g71419(.A (n_8848), .Y (n_8855));
NOR2X1 g71426(.A (n_10120), .B (g1221), .Y (n_8864));
OR2X1 g71439(.A (n_512), .B (n_10395), .Y (n_8885));
OR2X1 g63195_dup(.A (n_512), .B (n_10395), .Y (n_8886));
INVX1 g71440(.A (n_10225), .Y (n_10175));
CLKBUFX3 g71446(.A (n_8898), .Y (n_8895));
CLKBUFX1 g71452(.A (n_10227), .Y (n_8906));
CLKBUFX1 g71453(.A (n_8909), .Y (n_8908));
CLKBUFX1 g71458(.A (n_8915), .Y (n_8913));
CLKBUFX1 g71463(.A (g35), .Y (n_8921));
INVX8 g71489(.A (n_9107), .Y (n_8955));
INVX8 g71515(.A (n_9107), .Y (n_9000));
INVX2 g71522(.A (n_10385), .Y (n_9019));
INVX8 g71571(.A (n_9129), .Y (n_9091));
INVX4 g71584(.A (n_10687), .Y (n_9107));
INVX8 g71600(.A (n_10687), .Y (n_9129));
INVX1 g71609(.A (n_9139), .Y (n_9141));
INVX2 g71610(.A (n_9107), .Y (n_9139));
INVX1 g71618(.A (n_9129), .Y (n_9156));
INVX4 g71628(.A (n_9176), .Y (n_9172));
INVX1 g71630(.A (n_9167), .Y (n_9176));
INVX4 g71640(.A (n_9209), .Y (n_9193));
BUFX3 g71654(.A (n_10687), .Y (n_9209));
INVX4 g71655(.A (n_9269), .Y (n_9218));
INVX4 g71664(.A (n_9269), .Y (n_9234));
INVX4 g71668(.A (n_9269), .Y (n_9240));
INVX4 g71677(.A (n_9269), .Y (n_9256));
INVX4 g71686(.A (n_9279), .Y (n_9269));
INVX4 g71699(.A (n_9129), .Y (n_9279));
INVX1 g71705(.A (g35), .Y (n_9297));
INVX8 g71713(.A (n_9300), .Y (n_9311));
INVX2 g71723(.A (n_9300), .Y (n_9333));
INVX8 g71730(.A (n_9358), .Y (n_9300));
INVX2 g71739(.A (n_9351), .Y (n_9353));
CLKBUFX1 g71740(.A (n_9358), .Y (n_9351));
INVX8 g71747(.A (n_9371), .Y (n_9359));
INVX4 g71767(.A (n_9358), .Y (n_9371));
INVX1 g71770(.A (n_9398), .Y (n_9404));
BUFX3 g71773(.A (n_9358), .Y (n_9398));
BUFX3 g71775(.A (n_10949), .Y (n_9358));
INVX2 g71780(.A (n_9425), .Y (n_9419));
INVX4 g71782(.A (n_9419), .Y (n_9422));
INVX8 g71784(.A (n_9491), .Y (n_9425));
INVX2 g71788(.A (n_9425), .Y (n_9431));
INVX1 g71796(.A (n_9448), .Y (n_9443));
CLKBUFX1 g71799(.A (n_9493), .Y (n_9448));
INVX1 g71802(.A (n_9453), .Y (n_9454));
CLKBUFX3 g71804(.A (n_9493), .Y (n_9453));
INVX1 g71807(.A (n_9466), .Y (n_9461));
BUFX3 g71810(.A (n_9493), .Y (n_9466));
INVX1 g71812(.A (n_10952), .Y (n_9469));
INVX2 g71824(.A (n_9493), .Y (n_9491));
INVX4 g71828(.A (n_10716), .Y (n_9493));
INVX2 g71836(.A (n_9501), .Y (n_9505));
INVX2 g71837(.A (n_10716), .Y (n_9501));
INVX1 g71854(.A (n_9521), .Y (n_9526));
INVX4 g71863(.A (n_10376), .Y (n_9521));
INVX8 g71895(.A (n_9599), .Y (n_9558));
INVX8 g71898(.A (n_9553), .Y (n_9599));
INVX4 g71899(.A (n_10376), .Y (n_9553));
INVX1 g71917(.A (n_9628), .Y (n_9630));
INVX8 g71918(.A (n_9627), .Y (n_9628));
INVX4 g71931(.A (n_10782), .Y (n_9627));
INVX2 g71941(.A (n_10782), .Y (n_9651));
INVX4 g71953(.A (n_9672), .Y (n_9681));
INVX4 g71956(.A (n_9664), .Y (n_9672));
INVX2 g71961(.A (n_9664), .Y (n_9693));
BUFX3 g71962(.A (n_10950), .Y (n_9664));
INVX1 g71964(.A (n_9698), .Y (n_9697));
CLKBUFX1 g71972(.A (n_10949), .Y (n_9698));
INVX8 g72006(.A (n_9772), .Y (n_9750));
INVX4 g72018(.A (n_9717), .Y (n_9772));
CLKBUFX3 g72019(.A (n_10949), .Y (n_9717));
INVX8 g72031(.A (n_9775), .Y (n_9797));
INVX4 g72034(.A (n_9834), .Y (n_9775));
INVX8 g72036(.A (n_9775), .Y (n_9811));
INVX2 g72047(.A (n_9836), .Y (n_9830));
INVX4 g72052(.A (n_9834), .Y (n_9836));
BUFX3 g72060(.A (n_10949), .Y (n_9834));
INVX2 g72068(.A (n_9874), .Y (n_9856));
BUFX3 g72069(.A (n_9874), .Y (n_9862));
INVX1 g72071(.A (n_9862), .Y (n_9871));
INVX2 g72074(.A (n_10376), .Y (n_9874));
INVX1 g72080(.A (n_9884), .Y (n_9883));
CLKBUFX3 g72086(.A (n_10376), .Y (n_9884));
INVX8 g72088(.A (n_9928), .Y (n_9894));
INVX8 g72097(.A (n_9894), .Y (n_9903));
INVX4 g72120(.A (n_9903), .Y (n_9940));
CLKBUFX3 g72129(.A (n_10376), .Y (n_9928));
CLKBUFX1 g72132(.A (n_10376), .Y (n_9952));
INVX2 g72146(.A (n_9664), .Y (n_9976));
INVX1 g72148(.A (n_9952), .Y (n_9978));
INVX8 g72159(.A (n_10078), .Y (n_9992));
INVX8 g72169(.A (n_10078), .Y (n_10005));
INVX4 g72203(.A (n_10078), .Y (n_10063));
INVX8 g72221(.A (n_10013), .Y (n_10078));
BUFX3 g72222(.A (n_10949), .Y (n_10013));
INVX2 g72224(.A (n_10100), .Y (n_10097));
INVX2 g72225(.A (n_10100), .Y (n_10099));
INVX2 g72226(.A (n_10101), .Y (n_10100));
INVX1 g72228(.A (n_10107), .Y (n_10103));
INVX1 g72232(.A (n_10108), .Y (n_10107));
INVX2 g72233(.A (n_10631), .Y (n_10108));
CLKBUFX1 g72237(.A (n_10113), .Y (n_10112));
CLKBUFX1 g72239(.A (n_10532), .Y (n_10115));
CLKBUFX1 g72242(.A (n_10120), .Y (n_10119));
CLKBUFX1 g72245(.A (n_10125), .Y (n_10123));
CLKBUFX1 g72249(.A (n_10129), .Y (n_10128));
INVX1 g72253(.A (n_10139), .Y (n_10134));
INVX1 g72259(.A (g5016), .Y (n_10139));
CLKBUFX1 g72292(.A (n_10185), .Y (n_10184));
INVX1 g72294(.A (n_10192), .Y (n_10188));
INVX1 g72299(.A (g4991), .Y (n_10192));
CLKBUFX1 g72301(.A (n_10197), .Y (n_10196));
INVX1 g72303(.A (n_10200), .Y (n_10199));
CLKBUFX2 g72304(.A (n_10202), .Y (n_10200));
INVX1 g72305(.A (n_10202), .Y (n_10201));
CLKBUFX1 g72306(.A (n_10804), .Y (n_10202));
INVX2 g72307(.A (n_10804), .Y (n_10203));
CLKBUFX1 g72308(.A (n_10206), .Y (n_10205));
AND2X1 g72314(.A (n_10213), .B (n_11129), .Y (n_10214));
INVX2 g72315(.A (n_10997), .Y (n_10213));
INVX1 g72321(.A (n_10771), .Y (n_10216));
INVX1 g72322(.A (g5046), .Y (n_10217));
NOR2X1 g72326(.A (n_10224), .B (n_10226), .Y (n_10227));
CLKBUFX1 g72327(.A (g4785), .Y (n_10224));
INVX1 g72328(.A (n_10225), .Y (n_10226));
INVX2 g72329(.A (g4709), .Y (n_10225));
INVX1 g72330(.A (g4785), .Y (n_10228));
AND2X1 g51(.A (n_2444), .B (n_2331), .Y (n_10229));
NOR2X1 g72337(.A (n_10516), .B (n_10512), .Y (n_10238));
INVX1 g72338(.A (n_10514), .Y (n_10239));
NOR2X1 g72339(.A (n_7213), .B (n_7214), .Y (n_10240));
NOR2X1 g72340(.A (n_2442), .B (n_3326), .Y (n_10241));
OR2X1 g72343(.A (n_3364), .B (n_11077), .Y (n_10242));
NAND3X1 g72344(.A (n_11076), .B (n_1275), .C (n_3365), .Y (n_10243));
AOI21X1 g72345(.A0 (g1345), .A1 (g1361), .B0 (n_2177), .Y (n_10247));
CLKBUFX1 g72347(.A (n_10802), .Y (n_10245));
NOR2X1 g72356(.A (n_10257), .B (n_10260), .Y (n_10261));
NAND2X1 g72357(.A (n_11120), .B (n_10142), .Y (n_10257));
NAND4X1 g72358(.A (n_10628), .B (n_11094), .C (n_10259), .D(g_16311), .Y (n_10260));
AND2X1 g72360(.A (g_11293), .B (g_15691), .Y (n_10259));
AND2X1 g72361(.A (n_10628), .B (g_11293), .Y (n_10262));
AND2X1 g72362(.A (n_11094), .B (g_15691), .Y (n_10263));
INVX1 g72363(.A (n_10263), .Y (n_10264));
NAND2X1 g72367(.A (n_10270), .B (n_10271), .Y (n_10901));
NAND2X1 g72368(.A (n_10268), .B (n_10322), .Y (n_10270));
OAI21X1 g72369(.A0 (n_1298), .A1 (n_10829), .B0 (g17291), .Y(n_10268));
NOR2X1 g72371(.A (n_4120), .B (g1592), .Y (n_10271));
NAND2X1 g72379(.A (n_10283), .B (n_11122), .Y (n_10285));
AOI21X1 g72380(.A0 (n_10281), .A1 (n_10282), .B0 (n_8855), .Y(n_10283));
NOR2X1 g72381(.A (n_10867), .B (n_10280), .Y (n_10281));
INVX1 g72382(.A (g2697), .Y (n_10280));
AND2X1 g72384(.A (g2704), .B (n_11099), .Y (n_10282));
AND2X1 g72386(.A (n_10289), .B (g1585), .Y (n_10290));
AND2X1 g72387(.A (n_10288), .B (n_11122), .Y (n_10289));
NOR2X1 g72388(.A (n_10287), .B (n_8855), .Y (n_10288));
INVX1 g72389(.A (n_10286), .Y (n_10287));
NAND2X1 g72390(.A (n_10282), .B (g2697), .Y (n_10286));
CLKBUFX1 g72391(.A (n_10998), .Y (n_10296));
NAND2X1 g72402(.A (n_10306), .B (n_10312), .Y (n_10313));
NOR2X1 g72403(.A (n_10304), .B (n_8819), .Y (n_10306));
NAND3X1 g72404(.A (n_6612), .B (n_6618), .C (n_10303), .Y (n_10304));
NOR2X1 g72405(.A (n_10311), .B (g_5342), .Y (n_10303));
NOR2X1 g72407(.A (n_10307), .B (n_10311), .Y (n_10312));
INVX2 g72408(.A (g_10233), .Y (n_10307));
INVX2 g72409(.A (n_10310), .Y (n_10311));
INVX2 g72410(.A (n_10309), .Y (n_10310));
INVX2 g44(.A (n_10308), .Y (n_10309));
NAND2X2 g72411(.A (n_7094), .B (g_17653), .Y (n_10308));
INVX1 g72412(.A (n_10307), .Y (n_10314));
NAND3X1 g72413(.A (n_11138), .B (n_6612), .C (n_6618), .Y (n_10315));
AOI21X1 g72414(.A0 (n_10319), .A1 (n_10871), .B0 (n_10320), .Y(n_10321));
NOR2X1 g72415(.A (n_10317), .B (n_10318), .Y (n_10319));
INVX1 g72416(.A (n_10316), .Y (n_10317));
AND2X1 g72417(.A (n_11065), .B (n_10708), .Y (n_10316));
NAND3X1 g72418(.A (n_6697), .B (n_10723), .C (n_10649), .Y (n_10318));
NOR2X1 g72419(.A (n_10318), .B (n_10173), .Y (n_10320));
CLKBUFX1 g72420(.A (n_10322), .Y (n_10323));
NOR2X1 g72421(.A (n_10318), .B (n_10173), .Y (n_10322));
AOI21X1 g72422(.A0 (n_10327), .A1 (n_10328), .B0 (n_10329), .Y(n_10330));
NAND4X1 g72423(.A (n_11076), .B (n_10325), .C (n_10426), .D (g7946),.Y (n_10327));
INVX1 g72425(.A (n_1276), .Y (n_10325));
OR2X1 g72427(.A (n_3849), .B (n_6781), .Y (n_10328));
OR2X1 g72428(.A (g1532), .B (n_461), .Y (n_10329));
AOI21X1 g72436(.A0 (n_10342), .A1 (g5485), .B0 (n_10345), .Y(n_10346));
NAND2X1 g72437(.A (n_10781), .B (n_10341), .Y (n_10342));
AND2X1 g72439(.A (n_1484), .B (n_2443), .Y (n_10341));
NOR2X1 g72440(.A (n_10344), .B (n_10342), .Y (n_10345));
OAI21X1 g72441(.A0 (g5481), .A1 (g5475), .B0 (n_10343), .Y (n_10344));
NAND2X1 g72442(.A (g5481), .B (g5475), .Y (n_10343));
INVX1 g72443(.A (n_10342), .Y (n_10347));
NOR2X1 g72452(.A (n_10357), .B (n_10362), .Y (n_10363));
NOR2X1 g72453(.A (n_10687), .B (g5619), .Y (n_10357));
AOI21X1 g72455(.A0 (n_10948), .A1 (n_10519), .B0 (n_10361), .Y(n_10362));
OAI21X1 g72459(.A0 (n_10948), .A1 (g4821), .B0 (n_10687), .Y(n_10361));
NAND4X1 g72461(.A (g5248), .B (n_1695), .C (n_10833), .D (g14597), .Y(n_10368));
CLKBUFX3 g72463(.A (g5343), .Y (g25219));
INVX1 g72465(.A (g5343), .Y (n_10369));
AOI21X1 g72467(.A0 (n_10371), .A1 (n_10374), .B0 (n_10376), .Y(n_10377));
OR2X1 g72468(.A (g2227), .B (n_4699), .Y (n_10371));
NAND2X1 g72469(.A (g2153), .B (n_10373), .Y (n_10374));
INVX1 g72470(.A (n_10372), .Y (n_10373));
NAND2X1 g35_dup(.A (n_8532), .B (n_10763), .Y (n_10372));
INVX4 g72471(.A (n_10949), .Y (n_10376));
CLKBUFX1 g72473(.A (n_10372), .Y (n_10378));
INVX2 g72474(.A (n_10379), .Y (n_10380));
NAND2X2 g72475(.A (n_10763), .B (n_8532), .Y (n_10379));
NAND2X1 g72476(.A (n_10386), .B (n_10387), .Y (n_10388));
OAI21X1 g72477(.A0 (n_4840), .A1 (n_10383), .B0 (n_10385), .Y(n_10386));
NOR2X1 g72478(.A (n_10381), .B (n_10382), .Y (n_10383));
INVX1 g72479(.A (n_4839), .Y (n_10381));
INVX1 g72480(.A (n_1592), .Y (n_10382));
BUFX3 g72481(.A (n_10687), .Y (n_10385));
NAND2X1 g20(.A (n_10078), .B (g20049), .Y (n_10387));
NAND4X1 g72484(.A (n_10390), .B (n_10391), .C (n_10392), .D(n_10394), .Y (n_10395));
INVX1 g72485(.A (n_6574), .Y (n_10390));
NOR2X1 g72486(.A (n_23), .B (n_6578), .Y (n_10391));
NOR2X1 g72487(.A (n_7247), .B (n_46), .Y (n_10392));
NOR2X1 g72488(.A (n_3624), .B (n_46), .Y (n_10394));
NOR2X1 g72490(.A (n_10396), .B (n_10397), .Y (n_10398));
NAND2X1 g72491(.A (n_10391), .B (n_10392), .Y (n_10396));
OR2X1 g72492(.A (n_46), .B (n_6574), .Y (n_10397));
INVX1 g72493(.A (n_10397), .Y (n_10399));
INVX1 g72494(.A (n_10396), .Y (n_10400));
NOR2X1 g72495(.A (n_7247), .B (n_23), .Y (n_10401));
INVX1 g72496(.A (n_10401), .Y (n_10402));
NOR2X1 g72497(.A (n_10504), .B (g_18739), .Y (n_10404));
OR2X1 g72502(.A (n_10412), .B (n_10415), .Y (n_10416));
NAND4X1 g72503(.A (n_11218), .B (n_11219), .C (n_2968), .D (n_10411),.Y (n_10412));
NAND4X1 g72504(.A (n_6787), .B (n_690), .C (g4031), .D (g3913), .Y(n_11218));
NAND3X1 g73(.A (g3909), .B (n_803), .C (n_8917), .Y (n_10411));
NAND4X1 g72506(.A (n_6809), .B (n_10413), .C (n_10414), .D (n_1851),.Y (n_10415));
NAND4X1 g72507(.A (n_3894), .B (n_6808), .C (g3957), .D (g16748), .Y(n_10413));
NAND4X1 g72508(.A (n_3894), .B (n_4988), .C (g3941), .D (g13906), .Y(n_10414));
AND2X1 g72510(.A (n_11037), .B (n_8807), .Y (g25114));
AND2X1 g72514(.A (n_10425), .B (n_10426), .Y (n_10427));
NAND3X1 g72515(.A (n_10242), .B (n_10424), .C (n_10243), .Y(n_10425));
INVX1 g72516(.A (n_10423), .Y (n_10424));
AOI21X1 g72517(.A0 (n_10245), .A1 (n_10422), .B0 (n_10247), .Y(n_10423));
INVX1 g72518(.A (g1367), .Y (n_10422));
OR2X1 g72519(.A (g1322), .B (g1333), .Y (n_10426));
NAND2X1 g72520(.A (n_10428), .B (n_10426), .Y (n_10429));
NAND3X1 g72521(.A (n_10242), .B (n_10243), .C (n_10247), .Y(n_10428));
INVX1 g72522(.A (n_10430), .Y (n_10431));
NAND3X1 g72523(.A (n_10242), .B (n_10243), .C (n_10245), .Y(n_10430));
AOI21X1 g28(.A0 (n_10445), .A1 (n_10446), .B0 (n_10447), .Y(n_10448));
INVX2 g72533(.A (n_10444), .Y (n_10445));
NAND3X1 g72534(.A (n_2391), .B (n_10443), .C (n_69), .Y (n_10444));
AND2X1 g72535(.A (n_2352), .B (n_1457), .Y (n_10443));
XOR2X1 g72536(.A (g6167), .B (g6173), .Y (n_10446));
AND2X1 g72537(.A (n_10444), .B (g6177), .Y (n_10447));
NAND2X2 g72538(.A (n_2391), .B (n_69), .Y (n_3784));
NAND2X1 g72549(.A (n_10460), .B (n_10466), .Y (n_10467));
NAND2X1 g72550(.A (n_7025), .B (n_4190), .Y (n_10460));
NAND3X1 g72551(.A (n_10913), .B (n_7024), .C (g1816), .Y (n_10466));
NAND2X1 g72553(.A (n_10462), .B (n_10463), .Y (n_10464));
INVX1 g72554(.A (n_10461), .Y (n_10462));
NAND2X2 g72555(.A (n_2983), .B (n_1241), .Y (n_10461));
NAND2X1 g72556(.A (n_8756), .B (g17316), .Y (n_10463));
INVX1 g72559(.A (n_10472), .Y (n_10473));
NAND4X1 g72560(.A (n_10470), .B (n_1458), .C (n_10623), .D (g34028),.Y (n_10472));
NAND4X1 g72561(.A (n_8639), .B (n_8694), .C (n_10905), .D (g4754), .Y(n_10470));
NAND2X2 g72563(.A (n_10470), .B (g34028), .Y (n_3612));
AND2X1 g72564(.A (n_1458), .B (n_10623), .Y (n_10475));
INVX2 g72583(.A (n_10503), .Y (n_10499));
CLKBUFX1 g72586(.A (n_10504), .Y (n_10503));
CLKBUFX1 g72587(.A (n_10505), .Y (n_10504));
INVX2 g72588(.A (g_15838), .Y (n_10505));
CLKBUFX1 g72589(.A (n_10508), .Y (n_10506));
NAND4X1 g72593(.A (n_10513), .B (n_10515), .C (n_10517), .D(n_10518), .Y (n_10519));
NOR2X1 g72594(.A (n_2442), .B (n_10512), .Y (n_10513));
NAND2X1 g72595(.A (n_2438), .B (n_2329), .Y (n_10512));
NOR2X1 g72596(.A (n_3326), .B (n_10514), .Y (n_10515));
NAND2X1 g72597(.A (n_2382), .B (n_3281), .Y (n_10514));
INVX1 g72598(.A (n_10516), .Y (n_10517));
NAND3X1 g72599(.A (n_7208), .B (n_10229), .C (n_3268), .Y (n_10516));
NOR2X1 g72600(.A (n_7213), .B (n_7214), .Y (n_10518));
NAND4X1 g72601(.A (n_10526), .B (n_10527), .C (n_10528), .D (n_3388),.Y (n_10532));
INVX1 g72602(.A (n_10525), .Y (n_10526));
NAND3X1 g72603(.A (n_10520), .B (g_20951), .C (n_10524), .Y(n_10525));
AND2X1 g72604(.A (g_20952), .B (n_11116), .Y (n_10520));
INVX1 g72606(.A (n_10522), .Y (n_10524));
INVX1 g72608(.A (g_5029), .Y (n_10522));
NOR2X1 g72609(.A (g_8896), .B (n_780), .Y (n_10527));
INVX1 g72610(.A (g_18996), .Y (n_10528));
INVX1 g72611(.A (n_10529), .Y (n_3388));
INVX1 g72613(.A (g_19789), .Y (n_10529));
NOR2X1 g72614(.A (n_10534), .B (n_10520), .Y (n_10535));
NOR2X1 g72615(.A (n_11113), .B (g_20952), .Y (n_10534));
NOR2X1 g72628(.A (g_7563), .B (n_11027), .Y (n_11095));
INVX2 g72630(.A (g_22349), .Y (n_10557));
NAND4X1 g72631(.A (n_10558), .B (n_10708), .C (n_11065), .D(n_10649), .Y (n_10560));
NAND2X2 g26_dup(.A (n_10505), .B (n_8594), .Y (n_10558));
NOR2X1 g72634(.A (n_10564), .B (n_10565), .Y (n_10566));
OR2X1 g17(.A (n_11110), .B (n_10563), .Y (n_10564));
INVX1 g72635(.A (g_19515), .Y (n_10563));
OR2X1 g72636(.A (g_22600), .B (g_21318), .Y (n_10565));
NOR2X1 g72637(.A (g_21318), .B (n_11110), .Y (n_10567));
INVX1 g72638(.A (n_10563), .Y (n_10568));
AND2X1 g72639(.A (g_20952), .B (n_11116), .Y (n_10569));
NAND4X1 g72641(.A (n_10573), .B (n_10576), .C (g16627), .D (g3602),.Y (n_10577));
MX2X1 g72644(.A (g_9298), .B (n_11091), .S0 (n_10898), .Y (n_10573));
NOR2X1 g72646(.A (n_6979), .B (g3639), .Y (n_10576));
NAND2X1 g72647(.A (n_10883), .B (g11388), .Y (n_10578));
NAND3X1 g72648(.A (n_10587), .B (n_10588), .C (n_10589), .Y(n_10590));
NAND2X1 g72649(.A (n_10582), .B (n_9091), .Y (n_10587));
OAI21X1 g72650(.A0 (n_4805), .A1 (n_10579), .B0 (n_10581), .Y(n_10582));
OR2X1 g72651(.A (n_11055), .B (n_3177), .Y (n_10579));
OR2X1 g72652(.A (n_1286), .B (n_10580), .Y (n_10581));
OR2X1 g72653(.A (n_284), .B (n_3177), .Y (n_10580));
NAND3X1 g72658(.A (n_9894), .B (n_3177), .C (n_11055), .Y (n_10588));
NAND2X1 g72659(.A (n_9884), .B (g20899), .Y (n_10589));
NAND2X2 g72661(.A (n_9493), .B (n_10600), .Y (n_10601));
OAI21X1 g72665(.A0 (n_10596), .A1 (n_10597), .B0 (n_10599), .Y(n_10600));
NOR2X1 g72666(.A (n_10595), .B (n_4213), .Y (n_10596));
AND2X1 g72667(.A (n_3409), .B (n_685), .Y (n_10595));
NAND3X1 g72668(.A (n_1578), .B (n_477), .C (g4878), .Y (n_10597));
INVX1 g72669(.A (n_10598), .Y (n_10599));
AOI21X1 g72670(.A0 (n_1819), .A1 (n_844), .B0 (n_1830), .Y (n_10598));
NOR2X1 g72671(.A (n_8807), .B (n_11037), .Y (n_10833));
NAND3X1 g72676(.A (n_10607), .B (n_10846), .C (g2735), .Y (n_10609));
NOR2X1 g72677(.A (n_11013), .B (g2748), .Y (n_10607));
NOR2X1 g72682(.A (n_10613), .B (n_10617), .Y (n_10618));
XOR2X1 g72683(.A (n_6027), .B (n_878), .Y (n_10613));
NAND2X2 g72684(.A (n_5799), .B (n_10616), .Y (n_10617));
NAND2X2 g72686(.A (n_5617), .B (n_5705), .Y (n_10614));
AND2X1 g72687(.A (g1657), .B (g1624), .Y (n_10616));
INVX2 g72688(.A (n_10620), .Y (n_10621));
OR2X1 g72689(.A (n_8807), .B (n_11038), .Y (n_10620));
AND2X1 g72691(.A (n_11198), .B (g5990), .Y (n_10622));
CLKBUFX1 g72692(.A (n_10622), .Y (n_10623));
AND2X1 g72693(.A (n_10626), .B (n_11064), .Y (n_10628));
OR2X1 g72694(.A (n_10625), .B (n_11028), .Y (n_10626));
NAND2X1 g72695(.A (n_10624), .B (g_20837), .Y (n_10625));
INVX1 g72696(.A (g_7563), .Y (n_10624));
AOI21X1 g72699(.A0 (n_10633), .A1 (n_10634), .B0 (n_10637), .Y(n_10638));
INVX1 g72700(.A (n_10632), .Y (n_10633));
NAND2X2 g72701(.A (n_10630), .B (n_10631), .Y (n_10632));
INVX2 g72702(.A (g_22034), .Y (n_10630));
INVX2 g72703(.A (g_18238), .Y (n_10631));
INVX2 g72706(.A (g_22038), .Y (n_10634));
NAND2X1 g72707(.A (n_10522), .B (g_20951), .Y (n_10637));
NOR2X1 g72708(.A (n_552), .B (n_10632), .Y (n_10639));
INVX1 g72713(.A (n_10647), .Y (n_10644));
CLKBUFX1 g72717(.A (n_10649), .Y (n_10647));
CLKBUFX1 g72722(.A (n_10656), .Y (n_10650));
CLKBUFX2 g72727(.A (n_10657), .Y (n_10660));
INVX1 g72728(.A (n_10667), .Y (n_10664));
INVX1 g72731(.A (n_10404), .Y (n_10667));
INVX1 g72732(.A (n_10670), .Y (n_10669));
INVX2 g72733(.A (n_10671), .Y (n_10670));
CLKBUFX3 g72734(.A (n_10672), .Y (n_10671));
CLKBUFX3 g72735(.A (n_10937), .Y (n_10672));
INVX1 g72737(.A (n_10675), .Y (n_10674));
CLKBUFX2 g72738(.A (n_10937), .Y (n_10675));
XOR2X1 g72739(.A (g_20614), .B (n_10125), .Y (n_10678));
AOI21X1 g72741(.A0 (n_10686), .A1 (n_9167), .B0 (n_10689), .Y(n_10690));
OAI21X1 g72742(.A0 (g28753), .A1 (g21245), .B0 (n_10685), .Y(n_10686));
AND2X1 g43_dup(.A (n_2416), .B (g34026), .Y (g28753));
OR2X1 g72744(.A (n_3244), .B (n_10684), .Y (n_10685));
NAND2X1 g72746(.A (n_10682), .B (n_10683), .Y (n_10684));
NOR2X1 g72747(.A (n_3990), .B (n_3385), .Y (n_10682));
NOR2X1 g72748(.A (n_8736), .B (n_3044), .Y (n_10683));
BUFX3 g72749(.A (n_10687), .Y (n_9167));
BUFX3 g72750(.A (g35), .Y (n_10687));
NOR2X1 g72751(.A (n_9167), .B (g5272), .Y (n_10689));
AND2X1 g72754(.A (n_2416), .B (g34026), .Y (n_10693));
INVX2 g72755(.A (n_10699), .Y (n_10700));
NAND2X1 g72756(.A (n_10696), .B (n_10698), .Y (n_10699));
NAND3X1 g72757(.A (n_10216), .B (n_10695), .C (n_10217), .Y(n_10696));
AND2X1 g72758(.A (n_10766), .B (n_10694), .Y (n_10695));
INVX1 g72759(.A (g5052), .Y (n_10694));
OR2X1 g72760(.A (n_10694), .B (n_10697), .Y (n_10698));
NAND3X1 g72761(.A (n_10765), .B (g5046), .C (g5041), .Y (n_10697));
CLKBUFX2 g72769(.A (n_10709), .Y (n_10710));
AND2X1 g72770(.A (n_11065), .B (n_10708), .Y (n_10709));
INVX2 g72771(.A (g_18635), .Y (n_10708));
OAI21X1 g72772(.A0 (g_19913), .A1 (n_9664), .B0 (n_10714), .Y(n_10715));
NAND3X1 g72775(.A (n_10713), .B (n_9651), .C (n_7144), .Y (n_10714));
INVX1 g72776(.A (g_22605), .Y (n_10713));
INVX1 g72777(.A (n_10949), .Y (n_10716));
NAND2X2 g72778(.A (n_10720), .B (n_10976), .Y (n_10874));
NOR2X1 g72780(.A (n_11121), .B (n_8850), .Y (n_10717));
OAI21X1 g72781(.A0 (n_900), .A1 (n_2108), .B0 (g1430), .Y (n_10718));
NOR2X1 g72782(.A (g2629), .B (g2555), .Y (n_10720));
XOR2X1 g72783(.A (g1322), .B (g1339), .Y (n_11077));
CLKBUFX1 g72786(.A (n_10723), .Y (n_10724));
NAND2X1 g72787(.A (n_10505), .B (n_8594), .Y (n_10723));
NAND2X2 g72788(.A (n_1559), .B (n_6762), .Y (n_10725));
XOR2X1 g72806(.A (n_10745), .B (n_10751), .Y (n_10752));
OR4X1 g72807(.A (g_15287), .B (g13259), .C (g19334), .D (n_923), .Y(n_10745));
OR2X1 g72808(.A (n_10750), .B (n_10725), .Y (n_10751));
AOI21X1 g72809(.A0 (n_10123), .A1 (n_10746), .B0 (n_10749), .Y(n_10750));
NOR2X1 g72810(.A (n_10724), .B (g1236), .Y (n_10746));
NOR2X1 g72811(.A (n_10748), .B (n_10123), .Y (n_10749));
NAND2X1 g72812(.A (n_10747), .B (g1236), .Y (n_10748));
INVX1 g72813(.A (n_10724), .Y (n_10747));
NOR2X1 g72814(.A (n_10724), .B (n_10725), .Y (n_10753));
INVX2 g72815(.A (n_10760), .Y (n_10761));
OAI21X1 g72816(.A0 (g1585), .A1 (n_10755), .B0 (n_10759), .Y(n_10760));
CLKBUFX1 g72817(.A (n_10754), .Y (n_10755));
NAND3X1 g72818(.A (n_10201), .B (n_6670), .C (n_10710), .Y (n_10754));
NAND2X2 g72819(.A (n_10758), .B (n_10755), .Y (n_10759));
NAND4X1 g72820(.A (n_10199), .B (n_10756), .C (n_6673), .D (n_10871),.Y (n_10758));
CLKBUFX1 g72821(.A (n_10710), .Y (n_10756));
INVX1 g72823(.A (n_10759), .Y (n_10762));
INVX2 g72824(.A (n_10754), .Y (n_10763));
INVX1 g72825(.A (g1585), .Y (n_10764));
AOI21X1 g72826(.A0 (n_10765), .A1 (g5041), .B0 (n_10769), .Y(n_10770));
NOR2X1 g72827(.A (n_281), .B (n_1493), .Y (n_10765));
INVX1 g72828(.A (n_10768), .Y (n_10769));
NAND2X1 g72829(.A (n_10766), .B (n_10767), .Y (n_10768));
INVX1 g72830(.A (g5041), .Y (n_10766));
NOR2X1 g72831(.A (g5037), .B (n_6970), .Y (n_10767));
INVX1 g72832(.A (n_10767), .Y (n_10771));
INVX1 g72835(.A (n_7219), .Y (n_10772));
NAND2X1 g72836(.A (n_10519), .B (n_7217), .Y (n_10773));
AND2X1 g72839(.A (g34027), .B (n_2385), .Y (n_10781));
INVX1 g72840(.A (n_10949), .Y (n_10782));
NAND2X2 g72843(.A (n_5944), .B (n_10789), .Y (n_10790));
NAND2X2 g72845(.A (n_10785), .B (n_10993), .Y (n_10787));
OAI21X1 g72846(.A0 (n_6893), .A1 (g2819), .B0 (n_8557), .Y (n_10785));
AND2X1 g72848(.A (g2619), .B (g2587), .Y (n_10789));
NAND2X2 g72859(.A (n_10803), .B (g1536), .Y (n_10804));
NAND2X2 g72860(.A (n_10801), .B (n_10802), .Y (n_10803));
INVX1 g14(.A (g1351), .Y (n_10801));
INVX2 g72861(.A (g1312), .Y (n_10802));
NOR2X1 g72862(.A (n_6490), .B (n_6479), .Y (n_10805));
NOR2X1 g69657_dup(.A (n_6490), .B (n_6479), .Y (n_10806));
CLKBUFX1 g72864(.A (n_10809), .Y (n_10808));
INVX1 g72867(.A (n_10814), .Y (n_10813));
INVX1 g72868(.A (g_14843), .Y (n_10814));
INVX1 g72872(.A (n_10823), .Y (n_10818));
CLKBUFX1 g72879(.A (n_10826), .Y (n_10823));
INVX1 g72880(.A (g4776), .Y (n_10826));
INVX1 g72881(.A (n_10829), .Y (n_10827));
INVX1 g72883(.A (n_10831), .Y (n_10830));
CLKBUFX1 g72884(.A (n_10833), .Y (n_10831));
INVX1 g72885(.A (n_10839), .Y (n_10834));
INVX1 g72889(.A (g3288), .Y (n_10839));
INVX1 g72891(.A (n_10846), .Y (n_10841));
INVX1 g72899(.A (g2756), .Y (n_10846));
INVX1 g72901(.A (n_10853), .Y (n_10852));
CLKBUFX3 g72902(.A (n_10854), .Y (n_10853));
CLKBUFX3 g72903(.A (n_10961), .Y (n_10854));
INVX1 g72905(.A (n_10857), .Y (n_10856));
CLKBUFX1 g72906(.A (n_10961), .Y (n_10857));
INVX1 g72908(.A (n_10863), .Y (n_10861));
INVX1 g72910(.A (n_7040), .Y (n_10863));
CLKBUFX1 g72915(.A (n_10871), .Y (n_10867));
INVX1 g72916(.A (n_10874), .Y (n_10873));
INVX1 g72918(.A (n_10879), .Y (n_10877));
INVX2 g72920(.A (n_10573), .Y (n_10879));
INVX2 g72930(.A (n_10894), .Y (n_10889));
INVX1 g72932(.A (n_10894), .Y (n_10893));
INVX2 g72933(.A (n_10883), .Y (n_10894));
INVX2 g72934(.A (n_10883), .Y (n_10895));
INVX4 g72935(.A (n_10897), .Y (n_10883));
INVX2 g72936(.A (n_10898), .Y (n_10897));
INVX2 g72937(.A (g3689), .Y (n_10898));
INVX2 g72938(.A (n_10903), .Y (n_10899));
INVX1 g72940(.A (n_10901), .Y (n_10903));
INVX1 g72941(.A (n_10907), .Y (n_10906));
INVX1 g72942(.A (n_10905), .Y (n_10907));
INVX1 g72943(.A (n_10913), .Y (n_10910));
INVX1 g72944(.A (n_10912), .Y (n_10911));
INVX1 g72945(.A (n_10913), .Y (n_10912));
CLKBUFX3 g72946(.A (n_10915), .Y (n_10913));
INVX1 g72947(.A (n_10917), .Y (n_10916));
INVX2 g72948(.A (n_10915), .Y (n_10917));
CLKBUFX3 g72949(.A (n_10464), .Y (n_10915));
INVX1 g72950(.A (n_10920), .Y (n_10921));
CLKBUFX3 g72951(.A (n_6791), .Y (n_10920));
NAND3X1 g72959(.A (n_10932), .B (n_11033), .C (n_10936), .Y(n_10937));
OAI21X1 g33(.A0 (n_1166), .A1 (n_2108), .B0 (g17404), .Y (n_10932));
NAND2X1 g36_dup(.A (n_10709), .B (n_10203), .Y (n_10934));
NAND3X1 g72962(.A (n_10280), .B (g2704), .C (n_11097), .Y (n_10936));
NAND2X1 g72964(.A (n_10939), .B (n_10943), .Y (n_10944));
AND2X1 g16_dup(.A (g34035), .B (n_10181), .Y (n_10939));
INVX1 g13(.A (n_10942), .Y (n_10943));
NAND2X1 g72965(.A (n_10940), .B (n_10941), .Y (n_10942));
AND2X1 g72966(.A (n_8588), .B (g16624), .Y (n_10940));
AND2X1 g72967(.A (g3288), .B (n_7004), .Y (n_10941));
AND2X1 g16(.A (g34035), .B (n_10181), .Y (n_3249));
NAND2X1 g72968(.A (n_10951), .B (n_10954), .Y (n_10955));
NAND4X1 g72969(.A (n_10772), .B (n_10773), .C (n_10948), .D(n_10950), .Y (n_10951));
INVX1 g72970(.A (n_10947), .Y (n_10948));
NAND2X1 g72971(.A (n_2385), .B (g34027), .Y (n_10947));
CLKBUFX3 g72973(.A (n_10949), .Y (n_10950));
BUFX3 g1(.A (g35), .Y (n_10949));
AOI22X1 g72974(.A0 (n_10952), .A1 (g5467), .B0 (n_10953), .B1(n_10947), .Y (n_10954));
INVX2 g72975(.A (n_10950), .Y (n_10952));
AND2X1 g72976(.A (n_3616), .B (n_9862), .Y (n_10953));
NAND3X1 g72977(.A (n_11035), .B (n_10959), .C (n_10960), .Y(n_10961));
INVX1 g72979(.A (g1291), .Y (n_10956));
NAND2X2 g72980(.A (n_10203), .B (n_10709), .Y (n_11121));
OAI21X1 g72981(.A0 (n_909), .A1 (n_2108), .B0 (g17423), .Y (n_10959));
NAND3X1 g72982(.A (n_169), .B (g2697), .C (n_11097), .Y (n_10960));
NAND4X1 g98(.A (n_10968), .B (n_10972), .C (n_10973), .D (n_1586), .Y(n_10974));
NOR2X1 g99(.A (n_10964), .B (n_10967), .Y (n_10968));
NAND2X1 g101(.A (n_10962), .B (n_10963), .Y (n_10964));
NAND4X1 g107(.A (n_1499), .B (n_11030), .C (g3251), .D (g16603), .Y(n_10962));
NAND4X1 g105(.A (n_8586), .B (n_7383), .C (g3199), .D (g14421), .Y(n_10963));
NAND3X1 g100(.A (n_6948), .B (n_10965), .C (n_10966), .Y (n_10967));
NAND4X1 g104(.A (n_7383), .B (n_10941), .C (g16874), .D (g3223), .Y(n_10965));
NAND4X1 g103(.A (n_8572), .B (n_8587), .C (g16624), .D (g3203), .Y(n_10966));
AOI21X1 g102(.A0 (n_10970), .A1 (n_8572), .B0 (n_10971), .Y(n_10972));
INVX1 g108(.A (n_10969), .Y (n_10970));
NAND3X1 g109(.A (n_7383), .B (g16686), .C (g3255), .Y (n_10969));
NAND2X1 g110(.A (n_8552), .B (n_5501), .Y (n_10971));
NAND4X1 g106(.A (n_11029), .B (n_7383), .C (g3239), .D (g13865), .Y(n_10973));
OAI21X1 g72983(.A0 (n_10975), .A1 (g2629), .B0 (n_10980), .Y(n_10981));
AOI21X1 g72984(.A0 (n_10976), .A1 (n_6742), .B0 (g2555), .Y(n_10975));
NAND2X1 g72985(.A (n_10982), .B (g2555), .Y (n_10980));
CLKBUFX1 g72987(.A (n_10976), .Y (n_10978));
NAND2X2 g72989(.A (n_10718), .B (n_10717), .Y (n_10976));
INVX1 g72990(.A (n_10978), .Y (n_10982));
INVX2 g72991(.A (n_10983), .Y (n_10984));
NAND3X1 g72992(.A (g4849), .B (g4843), .C (n_11216), .Y (n_10983));
INVX1 g72994(.A (g1242), .Y (g23683));
AND2X1 g26_dup72995(.A (n_898), .B (n_10986), .Y (n_10987));
AOI21X1 g72996(.A0 (n_10557), .A1 (g_20563), .B0 (n_10560), .Y(n_10986));
AOI21X1 g72997(.A0 (n_10871), .A1 (n_10986), .B0 (n_10988), .Y(n_10989));
AND2X1 g72998(.A (n_10986), .B (n_898), .Y (n_10988));
OR2X1 g72999(.A (n_10991), .B (n_10994), .Y (n_10995));
NAND2X1 g73000(.A (g2060), .B (g2028), .Y (n_10991));
NAND2X1 g73001(.A (n_10992), .B (n_10993), .Y (n_10994));
OAI21X1 g73002(.A0 (g2787), .A1 (n_6892), .B0 (n_8557), .Y (n_10992));
AND2X1 g73003(.A (n_3679), .B (n_8895), .Y (n_10993));
INVX1 g73004(.A (n_10991), .Y (n_10996));
NOR2X1 g73005(.A (n_11129), .B (n_10997), .Y (n_10998));
INVX2 g73006(.A (g4899), .Y (n_10997));
CLKBUFX1 g73019(.A (n_11013), .Y (n_11012));
NOR2X1 g73027(.A (g1319), .B (n_10200), .Y (n_11025));
NOR2X1 g61156_dup(.A (g1319), .B (n_10200), .Y (n_11026));
NAND2X1 g73028(.A (n_10813), .B (n_6527), .Y (n_11027));
NAND2X1 g10_dup(.A (n_10813), .B (n_6527), .Y (n_11028));
NOR2X1 g73029(.A (n_10834), .B (n_7004), .Y (n_11029));
NOR2X1 g71188_dup(.A (n_10834), .B (n_7004), .Y (n_11030));
AOI21X1 g73030(.A0 (n_2479), .A1 (n_3713), .B0 (n_3718), .Y(n_11031));
AOI21X1 g62838_dup(.A0 (n_2479), .A1 (n_3713), .B0 (n_3718), .Y(n_11032));
AOI21X1 g73031(.A0 (n_10956), .A1 (g1448), .B0 (n_10934), .Y(n_11033));
AOI21X1 g72960_dup(.A0 (n_10956), .A1 (g1448), .B0 (n_10934), .Y(n_11034));
AOI21X1 g73032(.A0 (n_10956), .A1 (g1472), .B0 (n_11121), .Y(n_11035));
AOI21X1 g72978_dup(.A0 (n_10956), .A1 (g1472), .B0 (n_11121), .Y(n_11036));
INVX2 g73033(.A (n_11038), .Y (n_11037));
INVX1 g73034(.A (g5297), .Y (n_11038));
AOI21X1 g73035(.A0 (g23683), .A1 (n_10987), .B0 (n_10989), .Y(n_11039));
AOI21X1 g72993_dup(.A0 (g23683), .A1 (n_10987), .B0 (n_10989), .Y(n_11040));
NOR2X1 g73036(.A (n_11073), .B (n_3459), .Y (n_11041));
NOR2X1 g61208_dup(.A (n_11076), .B (n_3459), .Y (n_11042));
INVX1 g73039(.A (g12350), .Y (n_11045));
CLKBUFX1 g73042(.A (n_11050), .Y (g12350));
INVX1 g73044(.A (n_11064), .Y (n_11051));
INVX1 g73048(.A (n_11055), .Y (n_11056));
CLKBUFX3 g73052(.A (n_11064), .Y (n_11055));
CLKBUFX1 g73055(.A (n_11065), .Y (n_11064));
CLKBUFX1 g73058(.A (n_11071), .Y (n_11070));
CLKBUFX1 g73061(.A (n_11076), .Y (n_11073));
CLKBUFX2 g73062(.A (n_11077), .Y (n_11076));
CLKBUFX1 g73064(.A (n_11081), .Y (n_11080));
INVX2 g73070(.A (n_11088), .Y (g11388));
CLKBUFX1 g73073(.A (n_11091), .Y (n_11088));
INVX1 g73074(.A (g_9298), .Y (n_11091));
CLKBUFX1 g73076(.A (n_11095), .Y (n_11094));
CLKBUFX1 g73079(.A (n_11099), .Y (n_11097));
CLKBUFX1 g73082(.A (n_11105), .Y (n_11104));
INVX1 g73083(.A (n_11110), .Y (n_11106));
INVX1 g73088(.A (g_20244), .Y (n_11110));
CLKBUFX1 g73091(.A (n_11116), .Y (n_11113));
INVX1 g73093(.A (n_11119), .Y (n_11118));
CLKBUFX1 g73094(.A (n_11120), .Y (n_11119));
INVX2 g73095(.A (n_6907), .Y (n_11120));
INVX1 g73096(.A (n_11121), .Y (n_11122));
INVX1 g73097(.A (n_11126), .Y (n_11124));
CLKBUFX2 g73099(.A (n_11128), .Y (n_11126));
INVX1 g73103(.A (n_11134), .Y (n_11133));
CLKBUFX1 g73104(.A (n_11129), .Y (n_11134));
INVX1 g73106(.A (n_11129), .Y (n_11187));
INVX1 g73107(.A (n_8819), .Y (n_11138));
INVX4 g73122(.A (n_11150), .Y (n_11157));
BUFX3 g73124(.A (n_11160), .Y (n_11150));
INVX1 g73125(.A (g6381), .Y (n_11160));
CLKBUFX1 g73127(.A (n_11163), .Y (n_11162));
INVX1 g73128(.A (n_11186), .Y (n_11165));
INVX1 g73135(.A (n_11173), .Y (n_11171));
INVX2 g73137(.A (n_11177), .Y (n_11173));
CLKBUFX3 g73139(.A (n_11185), .Y (n_11177));
INVX1 g73140(.A (n_11184), .Y (n_11178));
CLKBUFX1 g73146(.A (n_11185), .Y (n_11184));
CLKBUFX1 g73147(.A (n_11186), .Y (n_11185));
NOR2X1 g73148(.A (n_10285), .B (n_10290), .Y (n_11190));
NOR2X1 g72378_dup(.A (n_10285), .B (n_10290), .Y (n_11191));
NAND3X1 g73149(.A (n_4206), .B (n_7088), .C (n_11205), .Y (n_11196));
NAND3X1 g70131_dup(.A (n_4206), .B (n_7088), .C (n_11206), .Y(n_11197));
CLKBUFX1 g73153(.A (n_11203), .Y (n_11201));
CLKBUFX1 g73154(.A (n_11198), .Y (n_11203));
NOR2X1 g73155(.A (n_7089), .B (n_7090), .Y (n_11205));
NOR2X1 g70135_dup(.A (n_7089), .B (n_7090), .Y (n_11206));
AOI21X1 g73156(.A0 (n_1564), .A1 (n_1747), .B0 (g4878), .Y (n_11207));
AOI21X1 g64564_dup(.A0 (n_1564), .A1 (n_1747), .B0 (g4878), .Y(n_11208));
NOR2X1 g73157(.A (n_8915), .B (n_10826), .Y (n_11209));
NOR2X1 g71226_dup(.A (n_8915), .B (n_10826), .Y (n_11210));
AND2X1 g73158(.A (n_10960), .B (n_11036), .Y (n_11211));
AND2X1 g70020_dup(.A (n_10960), .B (n_11036), .Y (n_11212));
endmodule
