module s27(blif_clk_net, blif_reset_net, G0, G1, G2, G3, G17);
input blif_clk_net, blif_reset_net, G0, G1, G2, G3;
output G17;
wire blif_clk_net, blif_reset_net, G0, G1, G2, G3;
wire G17;
wire G5, G6, G7, n_1, n_3, n_4, n_5, n_7;
wire n_8, n_11, n_12, n_14, n_15, n_16, n_21, n_26;
wire n_27, n_28;
DFFSRX1 G5_reg(.RN (n_15), .SN (1'b1), .CK (blif_clk_net), .D (n_16),.Q (G5), .QN ());
INVX2 g69(.A (n_14), .Y (n_16));
DFFSRX1 G6_reg(.RN (n_15), .SN (1'b1), .CK (blif_clk_net), .D (n_12),.Q (G6), .QN ());
NAND2X2 g70(.A (G17), .B (G0), .Y (n_14));
INVX1 g71(.A (G17), .Y (n_12));
DFFSRX1 G7_reg(.RN (n_15), .SN (1'b1), .CK (blif_clk_net), .D (n_11),.Q (G7), .QN ());
NOR2X1 g74(.A (G2), .B (n_8), .Y (n_11));
INVX1 g79(.A (n_7), .Y (n_8));
NAND2X1 g80(.A (n_3), .B (n_1), .Y (n_7));
OR2X1 g77(.A (G0), .B (n_4), .Y (n_5));
INVX1 g81(.A (G1), .Y (n_3));
INVX1 g86(.A (G7), .Y (n_1));
INVX1 g82(.A (G6), .Y (n_4));
INVX1 g84(.A (blif_reset_net), .Y (n_15));
NOR2X1 g23(.A (G0), .B (n_4), .Y (n_21));
NAND2X2 g17(.A (n_27), .B (n_28), .Y (G17));
NOR2X1 g18(.A (G5), .B (n_26), .Y (n_27));
NOR2X1 g19(.A (G3), .B (n_21), .Y (n_26));
NAND2X2 g90(.A (n_5), .B (n_7), .Y (n_28));
