module s27(blif_clk_net, blif_reset_net, G0, G1, G2, G3, G17, d_out_1, q_in_1, d_out_2, q_in_2, d_out_3, q_in_3);
input q_in_3;
input q_in_2;
input blif_clk_net, blif_reset_net, G0, G1, G2, G3;
input q_in_1;
output d_out_3;
output d_out_2;
output G17;
output d_out_1;
wire n_27, n_28;
wire n_8, n_11, n_12, n_14, n_15, n_16, n_21, n_26;
wire G5, G6, G7, n_1, n_3, n_4, n_5, n_7;
wire G17;
wire blif_clk_net, blif_reset_net, G0, G1, G2, G3;
CLKBUFX1 gbuf_d_1(.A(n_16), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(G5));
INVX2 g69(.A (n_14), .Y (n_16));
CLKBUFX1 gbuf_d_2(.A(n_12), .Y(d_out_2));
CLKBUFX1 gbuf_q_2(.A(q_in_2), .Y(G6));
NAND2X2 g70(.A (G17), .B (G0), .Y (n_14));
INVX1 g71(.A (G17), .Y (n_12));
CLKBUFX1 gbuf_d_3(.A(n_11), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(G7));
NOR2X1 g74(.A (G2), .B (n_8), .Y (n_11));
INVX1 g79(.A (n_7), .Y (n_8));
NAND2X1 g80(.A (n_3), .B (n_1), .Y (n_7));
OR2X1 g77(.A (G0), .B (n_4), .Y (n_5));
INVX1 g81(.A (G1), .Y (n_3));
INVX1 g86(.A (G7), .Y (n_1));
INVX1 g82(.A (G6), .Y (n_4));
INVX1 g84(.A (blif_reset_net), .Y (n_15));
NOR2X1 g23(.A (G0), .B (n_4), .Y (n_21));
NAND2X2 g17(.A (n_27), .B (n_28), .Y (G17));
NOR2X1 g18(.A (G5), .B (n_26), .Y (n_27));
NOR2X1 g19(.A (G3), .B (n_21), .Y (n_26));
NAND2X2 g90(.A (n_5), .B (n_7), .Y (n_28));
