module s38417(blif_clk_net, blif_reset_net, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380, d_out_1, q_in_1, d_out_2, q_in_2, d_out_3, qn_in_3, d_out_4, q_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, qn_in_7, d_out_8, q_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, d_out_12, qn_in_12, d_out_13, q_in_13, d_out_14, q_in_14, d_out_15, qn_in_15, d_out_16, q_in_16, d_out_17, q_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, q_in_20, d_out_21, q_in_21, d_out_22, q_in_22, d_out_23, q_in_23, d_out_24, q_in_24, d_out_25, q_in_25, d_out_26, q_in_26, d_out_27, q_in_27, d_out_28, q_in_28, d_out_29, q_in_29, d_out_30, q_in_30, d_out_31, q_in_31, d_out_32, q_in_32, d_out_33, q_in_33, d_out_34, q_in_34, d_out_35, q_in_35, d_out_36, q_in_36, d_out_37, q_in_37, d_out_38, q_in_38, d_out_39, q_in_39, d_out_40, q_in_40, d_out_41, q_in_41, d_out_42, q_in_42, d_out_43, q_in_43, d_out_44, q_in_44, d_out_45, q_in_45, d_out_46, q_in_46, d_out_47, q_in_47, d_out_48, q_in_48, d_out_49, q_in_49, d_out_50, q_in_50, d_out_51, q_in_51, d_out_52, q_in_52, d_out_53, q_in_53, d_out_54, q_in_54, d_out_55, q_in_55, d_out_56, q_in_56, d_out_57, q_in_57, d_out_58, qn_in_58, d_out_59, q_in_59, d_out_60, q_in_60, d_out_61, q_in_61, d_out_62, q_in_62, d_out_63, q_in_63, d_out_64, q_in_64, d_out_65, q_in_65, d_out_66, q_in_66, d_out_67, q_in_67, d_out_68, q_in_68, d_out_69, q_in_69, d_out_70, q_in_70, d_out_71, q_in_71, d_out_72, q_in_72, d_out_73, q_in_73, d_out_74, q_in_74, d_out_75, q_in_75, d_out_76, q_in_76, d_out_77, q_in_77, d_out_78, q_in_78, d_out_79, q_in_79, d_out_80, q_in_80, d_out_81, q_in_81, d_out_82, q_in_82, d_out_83, q_in_83, d_out_84, q_in_84, d_out_85, q_in_85, d_out_86, q_in_86, d_out_87, q_in_87, d_out_88, q_in_88, d_out_89, q_in_89, d_out_90, q_in_90, d_out_91, q_in_91, d_out_92, q_in_92, d_out_93, q_in_93, d_out_94, q_in_94, d_out_95, q_in_95, d_out_96, q_in_96, d_out_97, q_in_97, d_out_98, q_in_98, d_out_99, q_in_99, d_out_100, q_in_100, d_out_101, q_in_101, d_out_102, q_in_102, d_out_103, q_in_103, d_out_104, q_in_104, d_out_105, q_in_105, d_out_106, q_in_106, d_out_107, q_in_107, d_out_108, q_in_108, d_out_109, q_in_109, d_out_110, q_in_110, d_out_111, q_in_111, d_out_112, q_in_112, d_out_113, q_in_113, d_out_114, q_in_114, d_out_115, q_in_115, d_out_116, q_in_116, d_out_117, q_in_117, d_out_118, q_in_118, d_out_119, q_in_119, d_out_120, q_in_120, d_out_121, q_in_121, d_out_122, q_in_122, d_out_123, q_in_123, d_out_124, q_in_124, d_out_125, q_in_125, d_out_126, q_in_126, d_out_127, q_in_127, d_out_128, q_in_128, d_out_129, q_in_129, d_out_130, q_in_130, d_out_131, q_in_131, d_out_132, q_in_132, d_out_133, q_in_133, d_out_134, q_in_134, d_out_135, q_in_135, d_out_136, q_in_136, d_out_137, q_in_137, d_out_138, q_in_138, d_out_139, q_in_139, d_out_140, q_in_140, d_out_141, q_in_141, d_out_142, q_in_142, d_out_143, q_in_143, d_out_144, q_in_144, d_out_145, q_in_145, d_out_146, q_in_146, d_out_147, q_in_147, d_out_148, q_in_148, d_out_149, q_in_149, d_out_150, q_in_150, d_out_151, q_in_151, d_out_152, q_in_152, d_out_153, q_in_153, d_out_154, q_in_154, d_out_155, q_in_155, d_out_156, q_in_156, d_out_157, q_in_157, d_out_158, q_in_158, d_out_159, q_in_159, d_out_160, q_in_160, d_out_161, q_in_161, d_out_162, q_in_162, d_out_163, q_in_163, d_out_164, q_in_164, d_out_165, q_in_165, d_out_166, q_in_166, d_out_167, q_in_167, d_out_168, q_in_168, d_out_169, q_in_169, d_out_170, q_in_170, d_out_171, q_in_171, d_out_172, q_in_172, d_out_173, q_in_173, d_out_174, q_in_174, d_out_175, q_in_175, d_out_176, q_in_176, d_out_177, qn_in_177, d_out_178, qn_in_178, d_out_179, qn_in_179, d_out_180, q_in_180, d_out_181, q_in_181, d_out_182, q_in_182, d_out_183, q_in_183, d_out_184, q_in_184, d_out_185, q_in_185, d_out_186, q_in_186, d_out_187, q_in_187, d_out_188, q_in_188, d_out_189, q_in_189, d_out_190, q_in_190, d_out_191, q_in_191, d_out_192, q_in_192, d_out_193, q_in_193, d_out_194, q_in_194, d_out_195, q_in_195, d_out_196, q_in_196, d_out_197, q_in_197, d_out_198, q_in_198, d_out_199, q_in_199, d_out_200, q_in_200, d_out_201, q_in_201, d_out_202, q_in_202, d_out_203, q_in_203, d_out_204, q_in_204, d_out_205, q_in_205, d_out_206, q_in_206, d_out_207, q_in_207, d_out_208, q_in_208, d_out_209, q_in_209, d_out_210, q_in_210, d_out_211, q_in_211, d_out_212, q_in_212, d_out_213, q_in_213, d_out_214, q_in_214, d_out_215, q_in_215, d_out_216, q_in_216, d_out_217, q_in_217, d_out_218, q_in_218, d_out_219, q_in_219, d_out_220, q_in_220, d_out_221, q_in_221, d_out_222, qn_in_222, d_out_223, qn_in_223, d_out_224, q_in_224, d_out_225, q_in_225, d_out_226, q_in_226, d_out_227, qn_in_227, d_out_228, q_in_228, d_out_229, qn_in_229, d_out_230, q_in_230, d_out_231, q_in_231, d_out_232, q_in_232, d_out_233, q_in_233, d_out_234, q_in_234, d_out_235, q_in_235, d_out_236, q_in_236, d_out_237, qn_in_237, d_out_238, q_in_238, d_out_239, q_in_239, d_out_240, q_in_240, d_out_241, q_in_241, d_out_242, q_in_242, d_out_243, q_in_243, d_out_244, q_in_244, d_out_245, q_in_245, d_out_246, q_in_246, d_out_247, q_in_247, d_out_248, q_in_248, d_out_249, q_in_249, d_out_250, q_in_250, d_out_251, q_in_251, d_out_252, q_in_252, d_out_253, qn_in_253, d_out_254, q_in_254, d_out_255, q_in_255, d_out_256, q_in_256, d_out_257, q_in_257, d_out_258, q_in_258, d_out_259, q_in_259, d_out_260, q_in_260, d_out_261, q_in_261, d_out_262, q_in_262, d_out_263, q_in_263, d_out_264, q_in_264, d_out_265, q_in_265, d_out_266, q_in_266, d_out_267, q_in_267, d_out_268, q_in_268, d_out_269, q_in_269, d_out_270, q_in_270, d_out_271, q_in_271, d_out_272, q_in_272, d_out_273, q_in_273, d_out_274, q_in_274, d_out_275, q_in_275, d_out_276, q_in_276, d_out_277, q_in_277, d_out_278, q_in_278, d_out_279, q_in_279, d_out_280, q_in_280, d_out_281, q_in_281, d_out_282, q_in_282, d_out_283, q_in_283, d_out_284, q_in_284, d_out_285, q_in_285, d_out_286, q_in_286, d_out_287, q_in_287, d_out_288, q_in_288, d_out_289, q_in_289, d_out_290, q_in_290, d_out_291, q_in_291, d_out_292, q_in_292, d_out_293, q_in_293, d_out_294, qn_in_294, d_out_295, q_in_295, d_out_296, q_in_296, d_out_297, q_in_297, d_out_298, q_in_298, d_out_299, q_in_299, d_out_300, q_in_300, d_out_301, qn_in_301, d_out_302, qn_in_302, d_out_303, q_in_303, d_out_304, q_in_304, d_out_305, q_in_305, d_out_306, q_in_306, d_out_307, q_in_307, d_out_308, q_in_308, d_out_309, q_in_309, d_out_310, q_in_310, d_out_311, q_in_311, d_out_312, q_in_312, d_out_313, q_in_313, d_out_314, q_in_314, d_out_315, q_in_315, d_out_316, q_in_316, d_out_317, q_in_317, d_out_318, q_in_318, d_out_319, q_in_319, d_out_320, q_in_320, d_out_321, q_in_321, d_out_322, q_in_322, d_out_323, q_in_323, d_out_324, q_in_324, d_out_325, q_in_325, d_out_326, q_in_326, d_out_327, q_in_327, d_out_328, q_in_328, d_out_329, q_in_329, d_out_330, q_in_330, d_out_331, q_in_331, d_out_332, q_in_332, d_out_333, q_in_333, d_out_334, q_in_334, d_out_335, q_in_335, d_out_336, q_in_336, d_out_337, q_in_337, d_out_338, q_in_338, d_out_339, q_in_339, d_out_340, q_in_340, d_out_341, q_in_341, d_out_342, q_in_342, d_out_343, q_in_343, d_out_344, q_in_344, d_out_345, q_in_345, d_out_346, q_in_346, d_out_347, q_in_347, d_out_348, q_in_348, d_out_349, q_in_349, d_out_350, q_in_350, d_out_351, q_in_351, d_out_352, q_in_352, d_out_353, q_in_353, d_out_354, q_in_354, d_out_355, q_in_355, d_out_356, q_in_356, d_out_357, q_in_357, d_out_358, q_in_358, d_out_359, q_in_359, d_out_360, q_in_360, d_out_361, q_in_361, d_out_362, q_in_362, d_out_363, q_in_363, d_out_364, q_in_364, d_out_365, q_in_365, d_out_366, q_in_366, d_out_367, q_in_367, d_out_368, q_in_368, d_out_369, q_in_369, d_out_370, q_in_370, d_out_371, q_in_371, d_out_372, q_in_372, d_out_373, q_in_373, d_out_374, q_in_374, d_out_375, q_in_375, d_out_376, q_in_376, d_out_377, q_in_377, d_out_378, q_in_378, d_out_379, q_in_379, d_out_380, q_in_380, d_out_381, q_in_381, d_out_382, q_in_382, d_out_383, q_in_383, d_out_384, q_in_384, d_out_385, q_in_385, d_out_386, q_in_386, d_out_387, q_in_387, d_out_388, q_in_388, d_out_389, q_in_389, d_out_390, q_in_390, d_out_391, q_in_391, d_out_392, q_in_392, d_out_393, q_in_393, d_out_394, q_in_394, d_out_395, qn_in_395, d_out_396, q_in_396, d_out_397, q_in_397, d_out_398, q_in_398, d_out_399, q_in_399, d_out_400, q_in_400, d_out_401, q_in_401, d_out_402, q_in_402, d_out_403, q_in_403, d_out_404, q_in_404, d_out_405, q_in_405, d_out_406, q_in_406, d_out_407, q_in_407, d_out_408, q_in_408, d_out_409, q_in_409, d_out_410, q_in_410, d_out_411, q_in_411, d_out_412, q_in_412, d_out_413, q_in_413, d_out_414, q_in_414, d_out_415, q_in_415, d_out_416, q_in_416, d_out_417, q_in_417, d_out_418, q_in_418, d_out_419, q_in_419, d_out_420, q_in_420, d_out_421, q_in_421, d_out_422, q_in_422, d_out_423, q_in_423, d_out_424, q_in_424, d_out_425, q_in_425, d_out_426, q_in_426, d_out_427, q_in_427, d_out_428, qn_in_428, d_out_429, qn_in_429, d_out_430, qn_in_430, d_out_431, q_in_431, d_out_432, q_in_432, d_out_433, q_in_433, d_out_434, q_in_434, d_out_435, qn_in_435, d_out_436, qn_in_436, d_out_437, qn_in_437, d_out_438, qn_in_438, d_out_439, qn_in_439, d_out_440, qn_in_440, d_out_441, q_in_441, d_out_442, q_in_442, d_out_443, q_in_443, d_out_444, q_in_444, d_out_445, q_in_445, d_out_446, q_in_446, d_out_447, q_in_447, d_out_448, q_in_448, d_out_449, q_in_449, d_out_450, q_in_450, d_out_451, q_in_451, d_out_452, q_in_452, d_out_453, q_in_453, d_out_454, q_in_454, d_out_455, qn_in_455, d_out_456, qn_in_456, d_out_457, qn_in_457, d_out_458, qn_in_458, d_out_459, qn_in_459, d_out_460, qn_in_460, d_out_461, q_in_461, d_out_462, q_in_462, d_out_463, q_in_463, d_out_464, q_in_464, d_out_465, q_in_465, d_out_466, q_in_466, d_out_467, q_in_467, d_out_468, q_in_468, d_out_469, q_in_469, d_out_470, q_in_470, d_out_471, q_in_471, d_out_472, q_in_472, d_out_473, q_in_473, d_out_474, q_in_474, d_out_475, q_in_475, d_out_476, q_in_476, d_out_477, q_in_477, d_out_478, qn_in_478, d_out_479, qn_in_479, d_out_480, qn_in_480, d_out_481, q_in_481, d_out_482, q_in_482, d_out_483, q_in_483, d_out_484, q_in_484, d_out_485, q_in_485, d_out_486, qn_in_486, d_out_487, qn_in_487, d_out_488, q_in_488, d_out_489, q_in_489, d_out_490, q_in_490, d_out_491, q_in_491, d_out_492, q_in_492, d_out_493, q_in_493, d_out_494, q_in_494, d_out_495, q_in_495, d_out_496, q_in_496, d_out_497, q_in_497, d_out_498, q_in_498, d_out_499, q_in_499, d_out_500, q_in_500, d_out_501, q_in_501, d_out_502, qn_in_502, d_out_503, qn_in_503, d_out_504, qn_in_504, d_out_505, qn_in_505, d_out_506, q_in_506, d_out_507, qn_in_507, d_out_508, q_in_508, d_out_509, qn_in_509, d_out_510, qn_in_510, d_out_511, qn_in_511, d_out_512, qn_in_512, d_out_513, qn_in_513, d_out_514, qn_in_514, d_out_515, q_in_515, d_out_516, q_in_516, d_out_517, q_in_517, d_out_518, q_in_518, d_out_519, q_in_519, d_out_520, qn_in_520, d_out_521, q_in_521, d_out_522, q_in_522, d_out_523, q_in_523, d_out_524, q_in_524, d_out_525, q_in_525, d_out_526, q_in_526, d_out_527, q_in_527, d_out_528, q_in_528, d_out_529, q_in_529, d_out_530, q_in_530, d_out_531, q_in_531, d_out_532, q_in_532, d_out_533, qn_in_533, d_out_534, q_in_534, d_out_535, qn_in_535, d_out_536, q_in_536, d_out_537, q_in_537, d_out_538, qn_in_538, d_out_539, q_in_539, d_out_540, q_in_540, d_out_541, qn_in_541, d_out_542, q_in_542, d_out_543, q_in_543, d_out_544, q_in_544, d_out_545, q_in_545, d_out_546, q_in_546, d_out_547, qn_in_547, d_out_548, q_in_548, d_out_549, qn_in_549, d_out_550, q_in_550, d_out_551, qn_in_551, d_out_552, q_in_552, d_out_553, q_in_553, d_out_554, q_in_554, d_out_555, q_in_555, d_out_556, q_in_556, d_out_557, q_in_557, d_out_558, q_in_558, d_out_559, q_in_559, d_out_560, q_in_560, d_out_561, q_in_561, d_out_562, q_in_562, d_out_563, q_in_563, d_out_564, q_in_564, d_out_565, q_in_565, d_out_566, qn_in_566, d_out_567, qn_in_567, d_out_568, qn_in_568, d_out_569, q_in_569, d_out_570, q_in_570, d_out_571, q_in_571, d_out_572, q_in_572, d_out_573, q_in_573, d_out_574, q_in_574, d_out_575, q_in_575, d_out_576, q_in_576, d_out_577, q_in_577, d_out_578, q_in_578, d_out_579, q_in_579, d_out_580, q_in_580, d_out_581, q_in_581, d_out_582, q_in_582, d_out_583, q_in_583, d_out_584, qn_in_584, d_out_585, qn_in_585, d_out_586, q_in_586, d_out_587, q_in_587, d_out_588, qn_in_588, d_out_589, qn_in_589, d_out_590, q_in_590, d_out_591, q_in_591, d_out_592, q_in_592, d_out_593, qn_in_593, d_out_594, q_in_594, d_out_595, q_in_595, d_out_596, q_in_596, d_out_597, qn_in_597, d_out_598, q_in_598, d_out_599, q_in_599, d_out_600, q_in_600, d_out_601, q_in_601, d_out_602, q_in_602, d_out_603, q_in_603, d_out_604, q_in_604, d_out_605, q_in_605, d_out_606, q_in_606, d_out_607, q_in_607, d_out_608, q_in_608, d_out_609, qn_in_609, d_out_610, qn_in_610, d_out_611, q_in_611, d_out_612, q_in_612, d_out_613, q_in_613, d_out_614, q_in_614, d_out_615, q_in_615, d_out_616, q_in_616, d_out_617, q_in_617, d_out_618, q_in_618, d_out_619, q_in_619, d_out_620, q_in_620, d_out_621, q_in_621, d_out_622, q_in_622, d_out_623, q_in_623, d_out_624, q_in_624, d_out_625, q_in_625, d_out_626, q_in_626, d_out_627, q_in_627, d_out_628, q_in_628, d_out_629, q_in_629, d_out_630, q_in_630, d_out_631, q_in_631, d_out_632, q_in_632, d_out_633, q_in_633, d_out_634, q_in_634, d_out_635, q_in_635, d_out_636, q_in_636, d_out_637, qn_in_637, d_out_638, q_in_638, d_out_639, q_in_639, d_out_640, qn_in_640, d_out_641, q_in_641, d_out_642, q_in_642, d_out_643, q_in_643, d_out_644, q_in_644, d_out_645, q_in_645, d_out_646, q_in_646, d_out_647, q_in_647, d_out_648, q_in_648, d_out_649, qn_in_649, d_out_650, qn_in_650, d_out_651, q_in_651, d_out_652, q_in_652, d_out_653, q_in_653, d_out_654, q_in_654, d_out_655, q_in_655, d_out_656, q_in_656, d_out_657, q_in_657, d_out_658, q_in_658, d_out_659, q_in_659, d_out_660, q_in_660, d_out_661, q_in_661, d_out_662, q_in_662, d_out_663, qn_in_663, d_out_664, q_in_664, d_out_665, qn_in_665, d_out_666, q_in_666, d_out_667, q_in_667, d_out_668, q_in_668, d_out_669, q_in_669, d_out_670, qn_in_670, d_out_671, q_in_671, d_out_672, q_in_672, d_out_673, q_in_673, d_out_674, q_in_674, d_out_675, q_in_675, d_out_676, q_in_676, d_out_677, q_in_677, d_out_678, q_in_678, d_out_679, q_in_679, d_out_680, q_in_680, d_out_681, qn_in_681, d_out_682, q_in_682, d_out_683, qn_in_683, d_out_684, q_in_684, d_out_685, q_in_685, d_out_686, q_in_686, d_out_687, q_in_687, d_out_688, q_in_688, d_out_689, q_in_689, d_out_690, q_in_690, d_out_691, q_in_691, d_out_692, q_in_692, d_out_693, q_in_693, d_out_694, q_in_694, d_out_695, q_in_695, d_out_696, q_in_696, d_out_697, q_in_697, d_out_698, q_in_698, d_out_699, q_in_699, d_out_700, q_in_700, d_out_701, q_in_701, d_out_702, q_in_702, d_out_703, q_in_703, d_out_704, q_in_704, d_out_705, qn_in_705, d_out_706, q_in_706, d_out_707, q_in_707, d_out_708, q_in_708, d_out_709, q_in_709, d_out_710, q_in_710, d_out_711, q_in_711, d_out_712, q_in_712, d_out_713, q_in_713, d_out_714, q_in_714, d_out_715, q_in_715, d_out_716, q_in_716, d_out_717, q_in_717, d_out_718, q_in_718, d_out_719, q_in_719, d_out_720, q_in_720, d_out_721, q_in_721, d_out_722, q_in_722, d_out_723, q_in_723, d_out_724, q_in_724, d_out_725, q_in_725, d_out_726, q_in_726, d_out_727, q_in_727, d_out_728, q_in_728, d_out_729, q_in_729, d_out_730, q_in_730, d_out_731, q_in_731, d_out_732, q_in_732, d_out_733, q_in_733, d_out_734, q_in_734, d_out_735, q_in_735, d_out_736, q_in_736, d_out_737, q_in_737, d_out_738, q_in_738, d_out_739, q_in_739, d_out_740, q_in_740, d_out_741, q_in_741, d_out_742, q_in_742, d_out_743, q_in_743, d_out_744, q_in_744, d_out_745, q_in_745, d_out_746, qn_in_746, d_out_747, q_in_747, d_out_748, q_in_748, d_out_749, q_in_749, d_out_750, q_in_750, d_out_751, q_in_751, d_out_752, q_in_752, d_out_753, q_in_753, d_out_754, q_in_754, d_out_755, q_in_755, d_out_756, q_in_756, d_out_757, q_in_757, d_out_758, q_in_758, d_out_759, q_in_759, d_out_760, q_in_760, d_out_761, q_in_761, d_out_762, q_in_762, d_out_763, q_in_763, d_out_764, q_in_764, d_out_765, q_in_765, d_out_766, q_in_766, d_out_767, q_in_767, d_out_768, qn_in_768, d_out_769, q_in_769, d_out_770, q_in_770, d_out_771, q_in_771, d_out_772, q_in_772, d_out_773, q_in_773, d_out_774, q_in_774, d_out_775, q_in_775, d_out_776, q_in_776, d_out_777, q_in_777, d_out_778, q_in_778, d_out_779, q_in_779, d_out_780, q_in_780, d_out_781, q_in_781, d_out_782, q_in_782, d_out_783, q_in_783, d_out_784, q_in_784, d_out_785, q_in_785, d_out_786, qn_in_786, d_out_787, q_in_787, d_out_788, q_in_788, d_out_789, q_in_789, d_out_790, qn_in_790, d_out_791, q_in_791, d_out_792, q_in_792, d_out_793, q_in_793, d_out_794, q_in_794, d_out_795, q_in_795, d_out_796, q_in_796, d_out_797, q_in_797, d_out_798, q_in_798, d_out_799, q_in_799, d_out_800, q_in_800, d_out_801, q_in_801, d_out_802, q_in_802, d_out_803, q_in_803, d_out_804, q_in_804, d_out_805, q_in_805, d_out_806, q_in_806, d_out_807, q_in_807, d_out_808, q_in_808, d_out_809, q_in_809, d_out_810, q_in_810, d_out_811, q_in_811, d_out_812, q_in_812, d_out_813, q_in_813, d_out_814, q_in_814, d_out_815, q_in_815, d_out_816, q_in_816, d_out_817, q_in_817, d_out_818, q_in_818, d_out_819, qn_in_819, d_out_820, q_in_820, d_out_821, q_in_821, d_out_822, q_in_822, d_out_823, q_in_823, d_out_824, q_in_824, d_out_825, q_in_825, d_out_826, q_in_826, d_out_827, q_in_827, d_out_828, q_in_828, d_out_829, q_in_829, d_out_830, q_in_830, d_out_831, q_in_831, d_out_832, q_in_832, d_out_833, q_in_833, d_out_834, q_in_834, d_out_835, q_in_835, d_out_836, q_in_836, d_out_837, q_in_837, d_out_838, q_in_838, d_out_839, q_in_839, d_out_840, q_in_840, d_out_841, q_in_841, d_out_842, q_in_842, d_out_843, q_in_843, d_out_844, q_in_844, d_out_845, q_in_845, d_out_846, q_in_846, d_out_847, q_in_847, d_out_848, q_in_848, d_out_849, q_in_849, d_out_850, q_in_850, d_out_851, q_in_851, d_out_852, q_in_852, d_out_853, q_in_853, d_out_854, q_in_854, d_out_855, q_in_855, d_out_856, q_in_856, d_out_857, q_in_857, d_out_858, q_in_858, d_out_859, q_in_859, d_out_860, q_in_860, d_out_861, q_in_861, d_out_862, q_in_862, d_out_863, q_in_863, d_out_864, q_in_864, d_out_865, q_in_865, d_out_866, q_in_866, d_out_867, q_in_867, d_out_868, q_in_868, d_out_869, q_in_869, d_out_870, q_in_870, d_out_871, q_in_871, d_out_872, q_in_872, d_out_873, q_in_873, d_out_874, q_in_874, d_out_875, q_in_875, d_out_876, q_in_876, d_out_877, q_in_877, d_out_878, q_in_878, d_out_879, q_in_879, d_out_880, q_in_880, d_out_881, q_in_881, d_out_882, q_in_882, d_out_883, q_in_883, d_out_884, q_in_884, d_out_885, q_in_885, d_out_886, q_in_886, d_out_887, q_in_887, d_out_888, q_in_888, d_out_889, q_in_889, d_out_890, q_in_890, d_out_891, q_in_891, d_out_892, q_in_892, d_out_893, q_in_893, d_out_894, q_in_894, d_out_895, q_in_895, d_out_896, q_in_896, d_out_897, q_in_897, d_out_898, q_in_898, d_out_899, q_in_899, d_out_900, q_in_900, d_out_901, q_in_901, d_out_902, q_in_902, d_out_903, q_in_903, d_out_904, q_in_904, d_out_905, q_in_905, d_out_906, q_in_906, d_out_907, q_in_907, d_out_908, q_in_908, d_out_909, q_in_909, d_out_910, q_in_910, d_out_911, q_in_911, d_out_912, q_in_912, d_out_913, q_in_913, d_out_914, q_in_914, d_out_915, q_in_915, d_out_916, q_in_916, d_out_917, q_in_917, d_out_918, q_in_918, d_out_919, q_in_919, d_out_920, qn_in_920, d_out_921, q_in_921, d_out_922, q_in_922, d_out_923, q_in_923, d_out_924, q_in_924, d_out_925, q_in_925, d_out_926, q_in_926, d_out_927, q_in_927, d_out_928, q_in_928, d_out_929, q_in_929, d_out_930, q_in_930, d_out_931, q_in_931, d_out_932, qn_in_932, d_out_933, q_in_933, d_out_934, qn_in_934, d_out_935, q_in_935, d_out_936, q_in_936, d_out_937, q_in_937, d_out_938, q_in_938, d_out_939, q_in_939, d_out_940, q_in_940, d_out_941, q_in_941, d_out_942, q_in_942, d_out_943, q_in_943, d_out_944, q_in_944, d_out_945, q_in_945, d_out_946, q_in_946, d_out_947, q_in_947, d_out_948, q_in_948, d_out_949, q_in_949, d_out_950, q_in_950, d_out_951, q_in_951, d_out_952, q_in_952, d_out_953, q_in_953, d_out_954, q_in_954, d_out_955, q_in_955, d_out_956, q_in_956, d_out_957, q_in_957, d_out_958, q_in_958, d_out_959, q_in_959, d_out_960, q_in_960, d_out_961, q_in_961, d_out_962, q_in_962, d_out_963, q_in_963, d_out_964, q_in_964, d_out_965, q_in_965, d_out_966, q_in_966, d_out_967, q_in_967, d_out_968, q_in_968, d_out_969, q_in_969, d_out_970, q_in_970, d_out_971, q_in_971, d_out_972, q_in_972, d_out_973, q_in_973, d_out_974, q_in_974, d_out_975, q_in_975, d_out_976, q_in_976, d_out_977, q_in_977, d_out_978, q_in_978, d_out_979, q_in_979, d_out_980, q_in_980, d_out_981, q_in_981, d_out_982, q_in_982, d_out_983, q_in_983, d_out_984, q_in_984, d_out_985, q_in_985, d_out_986, q_in_986, d_out_987, q_in_987, d_out_988, q_in_988, d_out_989, q_in_989, d_out_990, q_in_990, d_out_991, q_in_991, d_out_992, q_in_992, d_out_993, q_in_993, d_out_994, q_in_994, d_out_995, q_in_995, d_out_996, q_in_996, d_out_997, q_in_997, d_out_998, q_in_998, d_out_999, q_in_999, d_out_1000, qn_in_1000, d_out_1001, q_in_1001, d_out_1002, q_in_1002, d_out_1003, q_in_1003, d_out_1004, q_in_1004, d_out_1005, q_in_1005, d_out_1006, q_in_1006, d_out_1007, q_in_1007, d_out_1008, q_in_1008, d_out_1009, q_in_1009, d_out_1010, q_in_1010, d_out_1011, q_in_1011, d_out_1012, q_in_1012, d_out_1013, q_in_1013, d_out_1014, q_in_1014, d_out_1015, q_in_1015, d_out_1016, q_in_1016, d_out_1017, q_in_1017, d_out_1018, q_in_1018, d_out_1019, q_in_1019, d_out_1020, q_in_1020, d_out_1021, q_in_1021, d_out_1022, q_in_1022, d_out_1023, q_in_1023, d_out_1024, q_in_1024, d_out_1025, q_in_1025, d_out_1026, q_in_1026, d_out_1027, q_in_1027, d_out_1028, q_in_1028, d_out_1029, q_in_1029, d_out_1030, q_in_1030, d_out_1031, q_in_1031, d_out_1032, q_in_1032, d_out_1033, q_in_1033, d_out_1034, q_in_1034, d_out_1035, q_in_1035, d_out_1036, q_in_1036, d_out_1037, q_in_1037, d_out_1038, q_in_1038, d_out_1039, q_in_1039, d_out_1040, q_in_1040, d_out_1041, q_in_1041, d_out_1042, q_in_1042, d_out_1043, q_in_1043, d_out_1044, q_in_1044, d_out_1045, q_in_1045, d_out_1046, q_in_1046, d_out_1047, q_in_1047, d_out_1048, q_in_1048, d_out_1049, q_in_1049, d_out_1050, q_in_1050, d_out_1051, q_in_1051, d_out_1052, q_in_1052, d_out_1053, q_in_1053, d_out_1054, q_in_1054, d_out_1055, q_in_1055, d_out_1056, qn_in_1056, d_out_1057, qn_in_1057, d_out_1058, q_in_1058, d_out_1059, q_in_1059, d_out_1060, qn_in_1060, d_out_1061, qn_in_1061, d_out_1062, q_in_1062, d_out_1063, q_in_1063, d_out_1064, qn_in_1064, d_out_1065, qn_in_1065, d_out_1066, qn_in_1066, d_out_1067, qn_in_1067, d_out_1068, qn_in_1068, d_out_1069, q_in_1069, d_out_1070, q_in_1070, d_out_1071, q_in_1071, d_out_1072, q_in_1072, d_out_1073, q_in_1073, d_out_1074, q_in_1074, d_out_1075, q_in_1075, d_out_1076, q_in_1076, d_out_1077, q_in_1077, d_out_1078, q_in_1078, d_out_1079, q_in_1079, d_out_1080, q_in_1080, d_out_1081, q_in_1081, d_out_1082, q_in_1082, d_out_1083, q_in_1083, d_out_1084, q_in_1084, d_out_1085, q_in_1085, d_out_1086, q_in_1086, d_out_1087, q_in_1087, d_out_1088, q_in_1088, d_out_1089, q_in_1089, d_out_1090, q_in_1090, d_out_1091, q_in_1091, d_out_1092, q_in_1092, d_out_1093, q_in_1093, d_out_1094, q_in_1094, d_out_1095, q_in_1095, d_out_1096, q_in_1096, d_out_1097, q_in_1097, d_out_1098, q_in_1098, d_out_1099, q_in_1099, d_out_1100, q_in_1100, d_out_1101, q_in_1101, d_out_1102, qn_in_1102, d_out_1103, q_in_1103, d_out_1104, q_in_1104, d_out_1105, qn_in_1105, d_out_1106, q_in_1106, d_out_1107, q_in_1107, d_out_1108, q_in_1108, d_out_1109, q_in_1109, d_out_1110, q_in_1110, d_out_1111, q_in_1111, d_out_1112, q_in_1112, d_out_1113, q_in_1113, d_out_1114, q_in_1114, d_out_1115, q_in_1115, d_out_1116, q_in_1116, d_out_1117, q_in_1117, d_out_1118, q_in_1118, d_out_1119, qn_in_1119, d_out_1120, qn_in_1120, d_out_1121, qn_in_1121, d_out_1122, q_in_1122, d_out_1123, q_in_1123, d_out_1124, q_in_1124, d_out_1125, q_in_1125, d_out_1126, q_in_1126, d_out_1127, q_in_1127, d_out_1128, q_in_1128, d_out_1129, q_in_1129, d_out_1130, q_in_1130, d_out_1131, q_in_1131, d_out_1132, q_in_1132, d_out_1133, q_in_1133, d_out_1134, q_in_1134, d_out_1135, q_in_1135, d_out_1136, q_in_1136, d_out_1137, qn_in_1137, d_out_1138, q_in_1138, d_out_1139, qn_in_1139, d_out_1140, qn_in_1140, d_out_1141, q_in_1141, d_out_1142, q_in_1142, d_out_1143, q_in_1143, d_out_1144, q_in_1144, d_out_1145, q_in_1145, d_out_1146, q_in_1146, d_out_1147, q_in_1147, d_out_1148, q_in_1148, d_out_1149, q_in_1149, d_out_1150, q_in_1150, d_out_1151, q_in_1151, d_out_1152, q_in_1152, d_out_1153, q_in_1153, d_out_1154, q_in_1154, d_out_1155, q_in_1155, d_out_1156, q_in_1156, d_out_1157, q_in_1157, d_out_1158, q_in_1158, d_out_1159, q_in_1159, d_out_1160, q_in_1160, d_out_1161, qn_in_1161, d_out_1162, qn_in_1162, d_out_1163, qn_in_1163, d_out_1164, q_in_1164, d_out_1165, q_in_1165, d_out_1166, q_in_1166, d_out_1167, q_in_1167, d_out_1168, q_in_1168, d_out_1169, q_in_1169, d_out_1170, q_in_1170, d_out_1171, q_in_1171, d_out_1172, q_in_1172, d_out_1173, q_in_1173, d_out_1174, q_in_1174, d_out_1175, qn_in_1175, d_out_1176, q_in_1176, d_out_1177, q_in_1177, d_out_1178, q_in_1178, d_out_1179, q_in_1179, d_out_1180, qn_in_1180, d_out_1181, qn_in_1181, d_out_1182, q_in_1182, d_out_1183, q_in_1183, d_out_1184, qn_in_1184, d_out_1185, qn_in_1185, d_out_1186, q_in_1186, d_out_1187, qn_in_1187, d_out_1188, q_in_1188, d_out_1189, q_in_1189, d_out_1190, qn_in_1190, d_out_1191, qn_in_1191, d_out_1192, q_in_1192, d_out_1193, q_in_1193, d_out_1194, qn_in_1194, d_out_1195, q_in_1195, d_out_1196, qn_in_1196, d_out_1197, q_in_1197, d_out_1198, q_in_1198, d_out_1199, qn_in_1199, d_out_1200, qn_in_1200, d_out_1201, qn_in_1201, d_out_1202, qn_in_1202, d_out_1203, q_in_1203, d_out_1204, qn_in_1204, d_out_1205, qn_in_1205, d_out_1206, q_in_1206, d_out_1207, q_in_1207, d_out_1208, qn_in_1208, d_out_1209, q_in_1209, d_out_1210, q_in_1210, d_out_1211, qn_in_1211, d_out_1212, qn_in_1212, d_out_1213, qn_in_1213, d_out_1214, qn_in_1214, d_out_1215, q_in_1215, d_out_1216, q_in_1216, d_out_1217, q_in_1217, d_out_1218, qn_in_1218, d_out_1219, q_in_1219, d_out_1220, qn_in_1220, d_out_1221, qn_in_1221, d_out_1222, q_in_1222, d_out_1223, q_in_1223, d_out_1224, qn_in_1224, d_out_1225, qn_in_1225, d_out_1226, q_in_1226, d_out_1227, qn_in_1227, d_out_1228, q_in_1228, d_out_1229, qn_in_1229, d_out_1230, q_in_1230, d_out_1231, qn_in_1231, d_out_1232, q_in_1232, d_out_1233, q_in_1233, d_out_1234, qn_in_1234, d_out_1235, qn_in_1235, d_out_1236, q_in_1236, d_out_1237, qn_in_1237, d_out_1238, q_in_1238, d_out_1239, q_in_1239, d_out_1240, q_in_1240, d_out_1241, q_in_1241, d_out_1242, q_in_1242, d_out_1243, q_in_1243, d_out_1244, qn_in_1244, d_out_1245, q_in_1245, d_out_1246, qn_in_1246, d_out_1247, q_in_1247, d_out_1248, qn_in_1248, d_out_1249, qn_in_1249, d_out_1250, qn_in_1250, d_out_1251, qn_in_1251, d_out_1252, q_in_1252, d_out_1253, qn_in_1253, d_out_1254, q_in_1254, d_out_1255, qn_in_1255, d_out_1256, q_in_1256, d_out_1257, q_in_1257, d_out_1258, q_in_1258, d_out_1259, q_in_1259, d_out_1260, q_in_1260, d_out_1261, q_in_1261, d_out_1262, q_in_1262, d_out_1263, qn_in_1263, d_out_1264, qn_in_1264, d_out_1265, q_in_1265, d_out_1266, qn_in_1266, d_out_1267, qn_in_1267, d_out_1268, qn_in_1268, d_out_1269, q_in_1269, d_out_1270, q_in_1270, d_out_1271, q_in_1271, d_out_1272, q_in_1272, d_out_1273, q_in_1273, d_out_1274, q_in_1274, d_out_1275, q_in_1275, d_out_1276, q_in_1276, d_out_1277, q_in_1277, d_out_1278, q_in_1278, d_out_1279, q_in_1279, d_out_1280, q_in_1280, d_out_1281, q_in_1281, d_out_1282, q_in_1282, d_out_1283, q_in_1283, d_out_1284, q_in_1284, d_out_1285, q_in_1285, d_out_1286, q_in_1286, d_out_1287, q_in_1287, d_out_1288, qn_in_1288, d_out_1289, q_in_1289, d_out_1290, q_in_1290, d_out_1291, q_in_1291, d_out_1292, qn_in_1292, d_out_1293, q_in_1293, d_out_1294, q_in_1294, d_out_1295, qn_in_1295, d_out_1296, q_in_1296, d_out_1297, qn_in_1297, d_out_1298, qn_in_1298, d_out_1299, q_in_1299, d_out_1300, q_in_1300, d_out_1301, q_in_1301, d_out_1302, q_in_1302, d_out_1303, q_in_1303, d_out_1304, q_in_1304, d_out_1305, q_in_1305, d_out_1306, q_in_1306, d_out_1307, q_in_1307, d_out_1308, qn_in_1308, d_out_1309, q_in_1309, d_out_1310, q_in_1310, d_out_1311, q_in_1311, d_out_1312, q_in_1312, d_out_1313, q_in_1313, d_out_1314, q_in_1314, d_out_1315, q_in_1315, d_out_1316, qn_in_1316, d_out_1317, q_in_1317, d_out_1318, qn_in_1318, d_out_1319, q_in_1319, d_out_1320, q_in_1320, d_out_1321, qn_in_1321, d_out_1322, q_in_1322, d_out_1323, q_in_1323, d_out_1324, q_in_1324, d_out_1325, q_in_1325, d_out_1326, q_in_1326, d_out_1327, q_in_1327, d_out_1328, qn_in_1328, d_out_1329, q_in_1329, d_out_1330, q_in_1330, d_out_1331, q_in_1331, d_out_1332, qn_in_1332, d_out_1333, qn_in_1333, d_out_1334, qn_in_1334, d_out_1335, q_in_1335, d_out_1336, q_in_1336, d_out_1337, q_in_1337, d_out_1338, q_in_1338, d_out_1339, q_in_1339, d_out_1340, q_in_1340, d_out_1341, qn_in_1341, d_out_1342, q_in_1342, d_out_1343, q_in_1343, d_out_1344, q_in_1344, d_out_1345, q_in_1345, d_out_1346, q_in_1346, d_out_1347, q_in_1347, d_out_1348, q_in_1348, d_out_1349, q_in_1349, d_out_1350, q_in_1350, d_out_1351, q_in_1351, d_out_1352, q_in_1352, d_out_1353, q_in_1353, d_out_1354, q_in_1354, d_out_1355, qn_in_1355, d_out_1356, q_in_1356, d_out_1357, q_in_1357, d_out_1358, q_in_1358, d_out_1359, q_in_1359, d_out_1360, q_in_1360, d_out_1361, q_in_1361, d_out_1362, q_in_1362, d_out_1363, q_in_1363, d_out_1364, q_in_1364, d_out_1365, q_in_1365, d_out_1366, q_in_1366, d_out_1367, q_in_1367, d_out_1368, q_in_1368, d_out_1369, qn_in_1369, d_out_1370, qn_in_1370, d_out_1371, q_in_1371, d_out_1372, qn_in_1372, d_out_1373, qn_in_1373, d_out_1374, q_in_1374, d_out_1375, qn_in_1375, d_out_1376, q_in_1376, d_out_1377, q_in_1377, d_out_1378, q_in_1378, d_out_1379, qn_in_1379, d_out_1380, qn_in_1380, d_out_1381, q_in_1381, d_out_1382, q_in_1382, d_out_1383, q_in_1383, d_out_1384, q_in_1384, d_out_1385, q_in_1385, d_out_1386, q_in_1386, d_out_1387, q_in_1387, d_out_1388, qn_in_1388, d_out_1389, q_in_1389, d_out_1390, qn_in_1390, d_out_1391, qn_in_1391, d_out_1392, q_in_1392, d_out_1393, q_in_1393, d_out_1394, qn_in_1394, d_out_1395, q_in_1395, d_out_1396, q_in_1396, d_out_1397, q_in_1397, d_out_1398, q_in_1398, d_out_1399, q_in_1399, d_out_1400, qn_in_1400, d_out_1401, q_in_1401, d_out_1402, qn_in_1402, d_out_1403, qn_in_1403, d_out_1404, qn_in_1404, d_out_1405, q_in_1405, d_out_1406, q_in_1406, d_out_1407, qn_in_1407, d_out_1408, q_in_1408, d_out_1409, q_in_1409, d_out_1410, qn_in_1410, d_out_1411, qn_in_1411, d_out_1412, q_in_1412, d_out_1413, q_in_1413, d_out_1414, q_in_1414, d_out_1415, qn_in_1415, d_out_1416, qn_in_1416, d_out_1417, q_in_1417, d_out_1418, qn_in_1418, d_out_1419, qn_in_1419, d_out_1420, q_in_1420, d_out_1421, q_in_1421, d_out_1422, qn_in_1422, d_out_1423, qn_in_1423, d_out_1424, q_in_1424, d_out_1425, q_in_1425, d_out_1426, qn_in_1426, d_out_1427, qn_in_1427, d_out_1428, qn_in_1428, d_out_1429, q_in_1429, d_out_1430, qn_in_1430, d_out_1431, q_in_1431, d_out_1432, qn_in_1432, d_out_1433, qn_in_1433, d_out_1434, qn_in_1434, d_out_1435, q_in_1435, d_out_1436, q_in_1436, d_out_1437, q_in_1437, d_out_1438, q_in_1438, d_out_1439, q_in_1439, d_out_1440, q_in_1440, d_out_1441, q_in_1441, d_out_1442, q_in_1442, d_out_1443, q_in_1443, d_out_1444, q_in_1444, d_out_1445, q_in_1445, d_out_1446, qn_in_1446, d_out_1447, q_in_1447, d_out_1448, q_in_1448, d_out_1449, q_in_1449, d_out_1450, q_in_1450, d_out_1451, q_in_1451, d_out_1452, q_in_1452, d_out_1453, q_in_1453, d_out_1454, q_in_1454, d_out_1455, q_in_1455, d_out_1456, q_in_1456, d_out_1457, q_in_1457, d_out_1458, q_in_1458, d_out_1459, qn_in_1459, d_out_1460, q_in_1460, d_out_1461, q_in_1461, d_out_1462, q_in_1462, d_out_1463, q_in_1463, d_out_1464, q_in_1464, d_out_1465, q_in_1465, d_out_1466, q_in_1466, d_out_1467, q_in_1467, d_out_1468, q_in_1468, d_out_1469, q_in_1469, d_out_1470, q_in_1470, d_out_1471, q_in_1471, d_out_1472, q_in_1472, d_out_1473, q_in_1473, d_out_1474, q_in_1474, d_out_1475, q_in_1475, d_out_1476, q_in_1476, d_out_1477, qn_in_1477, d_out_1478, q_in_1478, d_out_1479, q_in_1479, d_out_1480, q_in_1480, d_out_1481, q_in_1481, d_out_1482, q_in_1482, d_out_1483, q_in_1483, d_out_1484, q_in_1484, d_out_1485, q_in_1485, d_out_1486, q_in_1486, d_out_1487, q_in_1487, d_out_1488, q_in_1488, d_out_1489, q_in_1489, d_out_1490, q_in_1490, d_out_1491, q_in_1491, d_out_1492, q_in_1492, d_out_1493, q_in_1493, d_out_1494, q_in_1494, d_out_1495, q_in_1495, d_out_1496, q_in_1496, d_out_1497, q_in_1497, d_out_1498, q_in_1498, d_out_1499, q_in_1499, d_out_1500, qn_in_1500, d_out_1501, q_in_1501, d_out_1502, q_in_1502, d_out_1503, q_in_1503, d_out_1504, q_in_1504, d_out_1505, q_in_1505, d_out_1506, q_in_1506, d_out_1507, q_in_1507, d_out_1508, q_in_1508, d_out_1509, q_in_1509, d_out_1510, q_in_1510, d_out_1511, q_in_1511, d_out_1512, q_in_1512, d_out_1513, qn_in_1513, d_out_1514, q_in_1514, d_out_1515, q_in_1515, d_out_1516, q_in_1516, d_out_1517, q_in_1517, d_out_1518, q_in_1518, d_out_1519, qn_in_1519, d_out_1520, q_in_1520, d_out_1521, q_in_1521, d_out_1522, q_in_1522, d_out_1523, q_in_1523, d_out_1524, q_in_1524, d_out_1525, q_in_1525, d_out_1526, q_in_1526, d_out_1527, q_in_1527, d_out_1528, q_in_1528, d_out_1529, q_in_1529, d_out_1530, q_in_1530, d_out_1531, qn_in_1531, d_out_1532, q_in_1532, d_out_1533, qn_in_1533, d_out_1534, q_in_1534, d_out_1535, q_in_1535, d_out_1536, q_in_1536, d_out_1537, q_in_1537, d_out_1538, q_in_1538, d_out_1539, q_in_1539, d_out_1540, q_in_1540, d_out_1541, q_in_1541, d_out_1542, q_in_1542, d_out_1543, qn_in_1543, d_out_1544, q_in_1544, d_out_1545, q_in_1545, d_out_1546, q_in_1546, d_out_1547, q_in_1547, d_out_1548, q_in_1548, d_out_1549, q_in_1549, d_out_1550, q_in_1550, d_out_1551, q_in_1551, d_out_1552, q_in_1552, d_out_1553, q_in_1553, d_out_1554, q_in_1554, d_out_1555, q_in_1555, d_out_1556, q_in_1556, d_out_1557, q_in_1557, d_out_1558, qn_in_1558, d_out_1559, qn_in_1559, d_out_1560, q_in_1560, d_out_1561, q_in_1561, d_out_1562, q_in_1562, d_out_1563, q_in_1563, d_out_1564, q_in_1564);
input q_in_1436;
input q_in_1435;
input qn_in_1434;
input qn_in_1433;
input qn_in_1432;
input q_in_1431;
input qn_in_1430;
input q_in_1429;
input qn_in_1428;
input qn_in_1427;
input qn_in_1426;
input q_in_1425;
input q_in_1424;
input qn_in_1423;
input qn_in_1422;
input q_in_1421;
input q_in_1420;
input qn_in_1419;
input qn_in_1418;
input q_in_1417;
input qn_in_1416;
input qn_in_1415;
input q_in_1414;
input q_in_1413;
input q_in_1412;
input qn_in_1411;
input qn_in_1410;
input q_in_1409;
input q_in_1408;
input qn_in_1407;
input q_in_1406;
input q_in_1405;
input qn_in_1404;
input qn_in_1403;
input qn_in_1402;
input q_in_1401;
input qn_in_1400;
input q_in_1399;
input q_in_1398;
input q_in_1397;
input q_in_1396;
input q_in_1395;
input qn_in_1394;
input q_in_1393;
input q_in_1392;
input qn_in_1391;
input qn_in_1390;
input q_in_1389;
input qn_in_1388;
input q_in_1387;
input q_in_1386;
input q_in_1385;
input q_in_1384;
input q_in_1383;
input q_in_1382;
input q_in_1381;
input qn_in_1380;
input qn_in_1379;
input q_in_1378;
input q_in_1377;
input q_in_1376;
input qn_in_1375;
input q_in_1374;
input qn_in_1373;
input qn_in_1372;
input q_in_1371;
input qn_in_1370;
input qn_in_1369;
input q_in_1368;
input q_in_1367;
input q_in_1366;
input q_in_1365;
input q_in_1364;
input q_in_1363;
input q_in_1362;
input q_in_1361;
input q_in_1360;
input q_in_1359;
input q_in_1358;
input q_in_1357;
input q_in_1356;
input qn_in_1355;
input q_in_1354;
input q_in_1353;
input q_in_1352;
input q_in_1351;
input q_in_1350;
input q_in_1349;
input q_in_1348;
input q_in_1347;
input q_in_1346;
input q_in_1345;
input q_in_1344;
input q_in_1343;
input q_in_1342;
input qn_in_1341;
input q_in_1340;
input q_in_1339;
input q_in_1338;
input q_in_1337;
input q_in_1336;
input q_in_1335;
input qn_in_1334;
input qn_in_1333;
input qn_in_1332;
input q_in_1331;
input q_in_1330;
input q_in_1329;
input qn_in_1328;
input q_in_1327;
input q_in_1326;
input q_in_1325;
input q_in_1324;
input q_in_1323;
input q_in_1322;
input qn_in_1321;
input q_in_1320;
input q_in_1319;
input qn_in_1318;
input q_in_1317;
input qn_in_1316;
input q_in_1315;
input q_in_1314;
input q_in_1313;
input q_in_1312;
input q_in_1311;
input q_in_1310;
input q_in_1309;
input qn_in_1308;
input q_in_1307;
input q_in_1306;
input q_in_1305;
input q_in_1304;
input q_in_1303;
input q_in_1302;
input q_in_1301;
input q_in_1300;
input q_in_1299;
input qn_in_1298;
input qn_in_1297;
input q_in_1296;
input qn_in_1295;
input q_in_1294;
input q_in_1293;
input qn_in_1292;
input q_in_1291;
input q_in_1290;
input q_in_1289;
input qn_in_1288;
input q_in_1287;
input q_in_1286;
input q_in_1285;
input q_in_1284;
input q_in_1283;
input q_in_1282;
input q_in_1281;
input q_in_1280;
input q_in_1279;
input q_in_1278;
input q_in_1277;
input q_in_1276;
input q_in_1275;
input q_in_1274;
input q_in_1273;
input q_in_1272;
input q_in_1271;
input q_in_1270;
input q_in_1269;
input qn_in_1268;
input qn_in_1267;
input qn_in_1266;
input q_in_1265;
input qn_in_1264;
input qn_in_1263;
input q_in_1262;
input q_in_1261;
input q_in_1260;
input q_in_1259;
input q_in_1258;
input q_in_1257;
input q_in_1256;
input qn_in_1255;
input q_in_1254;
input qn_in_1253;
input q_in_1252;
input qn_in_1251;
input qn_in_1250;
input qn_in_1249;
input qn_in_1248;
input q_in_1247;
input qn_in_1246;
input q_in_1245;
input qn_in_1244;
input q_in_1243;
input q_in_1242;
input q_in_1241;
input q_in_1240;
input q_in_1239;
input q_in_1238;
input qn_in_1237;
input q_in_1236;
input qn_in_1235;
input qn_in_1234;
input q_in_1233;
input q_in_1232;
input qn_in_1231;
input q_in_1230;
input qn_in_1229;
input q_in_1228;
input qn_in_1227;
input q_in_1226;
input qn_in_1225;
input qn_in_1224;
input q_in_1223;
input q_in_1222;
input qn_in_1221;
input qn_in_1220;
input q_in_1219;
input qn_in_1218;
input q_in_1217;
input q_in_1216;
input q_in_1215;
input qn_in_1214;
input qn_in_1213;
input qn_in_1212;
input qn_in_1211;
input q_in_1210;
input q_in_1209;
input qn_in_1208;
input q_in_1207;
input q_in_1206;
input qn_in_1205;
input qn_in_1204;
input q_in_1203;
input qn_in_1202;
input qn_in_1201;
input qn_in_1200;
input qn_in_1199;
input q_in_1198;
input q_in_1197;
input qn_in_1196;
input q_in_1195;
input qn_in_1194;
input q_in_1193;
input q_in_1192;
input qn_in_1191;
input qn_in_1190;
input q_in_1189;
input q_in_1188;
input qn_in_1187;
input q_in_1186;
input qn_in_1185;
input qn_in_1184;
input q_in_1183;
input q_in_1182;
input qn_in_1181;
input qn_in_1180;
input q_in_1179;
input q_in_1178;
input q_in_1177;
input q_in_1176;
input qn_in_1175;
input q_in_1174;
input q_in_1173;
input q_in_1172;
input q_in_1171;
input q_in_1170;
input q_in_1169;
input q_in_1168;
input q_in_1167;
input q_in_1166;
input q_in_1165;
input q_in_1164;
input qn_in_1163;
input qn_in_1162;
input qn_in_1161;
input q_in_1160;
input q_in_1159;
input q_in_1158;
input q_in_1157;
input q_in_1156;
input q_in_1155;
input q_in_1154;
input q_in_1153;
input q_in_1152;
input q_in_1151;
input q_in_1150;
input q_in_1149;
input q_in_1148;
input q_in_1147;
input q_in_1146;
input q_in_1145;
input q_in_1144;
input q_in_1143;
input q_in_1142;
input q_in_1141;
input qn_in_1140;
input qn_in_1139;
input q_in_1138;
input qn_in_1137;
input q_in_1136;
input q_in_1135;
input q_in_1134;
input q_in_1133;
input q_in_1132;
input q_in_1131;
input q_in_1130;
input q_in_1129;
input q_in_1128;
input q_in_1127;
input q_in_1126;
input q_in_1125;
input q_in_1124;
input q_in_1123;
input q_in_1122;
input qn_in_1121;
input qn_in_1120;
input qn_in_1119;
input q_in_1118;
input q_in_1117;
input q_in_1116;
input q_in_1115;
input q_in_1114;
input q_in_1113;
input q_in_1112;
input q_in_1111;
input q_in_1110;
input q_in_1109;
input q_in_1108;
input q_in_1107;
input q_in_1106;
input qn_in_1105;
input q_in_1104;
input q_in_1103;
input qn_in_1102;
input q_in_1101;
input q_in_1100;
input q_in_1099;
input q_in_1098;
input q_in_1097;
input q_in_1096;
input q_in_1095;
input q_in_1094;
input q_in_1093;
input q_in_1092;
input q_in_1091;
input q_in_1090;
input q_in_1089;
input q_in_1088;
input q_in_1087;
input q_in_1086;
input q_in_1085;
input q_in_1084;
input q_in_1083;
input q_in_1082;
input q_in_1081;
input q_in_1080;
input q_in_1079;
input q_in_1078;
input q_in_1077;
input q_in_1076;
input q_in_1075;
input q_in_1074;
input q_in_1073;
input q_in_1072;
input q_in_1071;
input q_in_1070;
input q_in_1069;
input qn_in_1068;
input qn_in_1067;
input qn_in_1066;
input qn_in_1065;
input qn_in_1064;
input q_in_1063;
input q_in_1062;
input qn_in_1061;
input qn_in_1060;
input q_in_1059;
input q_in_1058;
input qn_in_1057;
input qn_in_1056;
input q_in_1055;
input q_in_1054;
input q_in_1053;
input q_in_1052;
input q_in_1051;
input q_in_1050;
input q_in_1049;
input q_in_1048;
input q_in_1047;
input q_in_1046;
input q_in_1045;
input q_in_1044;
input q_in_1043;
input q_in_1042;
input q_in_1041;
input q_in_1040;
input q_in_1039;
input q_in_1038;
input q_in_1037;
input q_in_1036;
input q_in_1035;
input q_in_1034;
input q_in_1033;
input q_in_1032;
input q_in_1031;
input q_in_1030;
input q_in_1029;
input q_in_1028;
input q_in_1027;
input q_in_1026;
input q_in_1025;
input q_in_1024;
input q_in_1023;
input q_in_1022;
input q_in_1021;
input q_in_1020;
input q_in_1019;
input q_in_1018;
input q_in_1017;
input q_in_1016;
input q_in_1015;
input q_in_1014;
input q_in_1013;
input q_in_1012;
input q_in_1011;
input q_in_1010;
input q_in_1009;
input q_in_1008;
input q_in_1007;
input q_in_1006;
input q_in_1005;
input q_in_1004;
input q_in_1003;
input q_in_1002;
input q_in_1001;
input qn_in_1000;
input q_in_999;
input q_in_998;
input q_in_997;
input q_in_996;
input q_in_995;
input q_in_994;
input q_in_993;
input q_in_992;
input q_in_991;
input q_in_990;
input q_in_989;
input q_in_988;
input q_in_987;
input q_in_986;
input q_in_985;
input q_in_984;
input q_in_983;
input q_in_982;
input q_in_981;
input q_in_980;
input q_in_979;
input q_in_978;
input q_in_977;
input q_in_976;
input q_in_975;
input q_in_974;
input q_in_973;
input q_in_972;
input q_in_971;
input q_in_970;
input q_in_969;
input q_in_968;
input q_in_967;
input q_in_966;
input q_in_965;
input q_in_964;
input q_in_963;
input q_in_962;
input q_in_961;
input q_in_960;
input q_in_959;
input q_in_958;
input q_in_957;
input q_in_956;
input q_in_955;
input q_in_954;
input q_in_953;
input q_in_952;
input q_in_951;
input q_in_950;
input q_in_949;
input q_in_948;
input q_in_947;
input q_in_946;
input q_in_945;
input q_in_944;
input q_in_943;
input q_in_942;
input q_in_941;
input q_in_940;
input q_in_939;
input q_in_938;
input q_in_937;
input q_in_936;
input q_in_935;
input qn_in_934;
input q_in_933;
input qn_in_932;
input q_in_931;
input q_in_930;
input q_in_929;
input q_in_928;
input q_in_927;
input q_in_926;
input q_in_925;
input q_in_924;
input q_in_923;
input q_in_922;
input q_in_921;
input qn_in_920;
input q_in_919;
input q_in_918;
input q_in_917;
input q_in_916;
input q_in_915;
input q_in_914;
input q_in_913;
input q_in_912;
input q_in_911;
input q_in_910;
input q_in_909;
input q_in_908;
input q_in_907;
input q_in_906;
input q_in_905;
input q_in_904;
input q_in_903;
input q_in_902;
input q_in_901;
input q_in_900;
input q_in_899;
input q_in_898;
input q_in_897;
input q_in_896;
input q_in_895;
input q_in_894;
input q_in_893;
input q_in_892;
input q_in_891;
input q_in_890;
input q_in_889;
input q_in_888;
input q_in_887;
input q_in_886;
input q_in_885;
input q_in_884;
input q_in_883;
input q_in_882;
input q_in_881;
input q_in_880;
input q_in_879;
input q_in_878;
input q_in_877;
input q_in_876;
input q_in_875;
input q_in_874;
input q_in_873;
input q_in_872;
input q_in_871;
input q_in_870;
input q_in_869;
input q_in_868;
input q_in_867;
input q_in_866;
input q_in_865;
input q_in_864;
input q_in_863;
input q_in_862;
input q_in_861;
input q_in_860;
input q_in_859;
input q_in_858;
input q_in_857;
input q_in_856;
input q_in_855;
input q_in_854;
input q_in_853;
input q_in_852;
input q_in_851;
input q_in_850;
input q_in_849;
input q_in_848;
input q_in_847;
input q_in_846;
input q_in_845;
input q_in_844;
input q_in_843;
input q_in_842;
input q_in_841;
input q_in_840;
input q_in_839;
input q_in_838;
input q_in_837;
input q_in_836;
input q_in_835;
input q_in_834;
input q_in_833;
input q_in_832;
input q_in_831;
input q_in_830;
input q_in_829;
input q_in_828;
input q_in_827;
input q_in_826;
input q_in_825;
input q_in_824;
input q_in_823;
input q_in_822;
input q_in_821;
input q_in_820;
input qn_in_819;
input q_in_818;
input q_in_817;
input q_in_816;
input q_in_815;
input q_in_814;
input q_in_813;
input q_in_812;
input q_in_811;
input q_in_810;
input q_in_809;
input q_in_808;
input q_in_807;
input q_in_806;
input q_in_805;
input q_in_804;
input q_in_803;
input q_in_802;
input q_in_801;
input q_in_800;
input q_in_799;
input q_in_798;
input q_in_797;
input q_in_796;
input q_in_795;
input q_in_794;
input q_in_793;
input q_in_792;
input q_in_791;
input qn_in_790;
input q_in_789;
input q_in_788;
input q_in_787;
input qn_in_786;
input q_in_785;
input q_in_784;
input q_in_783;
input q_in_782;
input q_in_781;
input q_in_780;
input q_in_779;
input q_in_778;
input q_in_777;
input q_in_776;
input q_in_775;
input q_in_774;
input q_in_773;
input q_in_772;
input q_in_771;
input q_in_770;
input q_in_769;
input qn_in_768;
input q_in_767;
input q_in_766;
input q_in_765;
input q_in_764;
input q_in_763;
input q_in_762;
input q_in_761;
input q_in_760;
input q_in_759;
input q_in_758;
input q_in_757;
input q_in_756;
input q_in_755;
input q_in_754;
input q_in_753;
input q_in_752;
input q_in_751;
input q_in_750;
input q_in_749;
input q_in_748;
input q_in_747;
input qn_in_746;
input q_in_745;
input q_in_744;
input q_in_743;
input q_in_742;
input q_in_741;
input q_in_740;
input q_in_739;
input q_in_738;
input q_in_737;
input q_in_736;
input q_in_735;
input q_in_734;
input q_in_733;
input q_in_732;
input q_in_731;
input q_in_730;
input q_in_729;
input q_in_728;
input q_in_727;
input q_in_726;
input q_in_725;
input q_in_724;
input q_in_723;
input q_in_722;
input q_in_721;
input q_in_720;
input q_in_719;
input q_in_718;
input q_in_717;
input q_in_716;
input q_in_715;
input q_in_714;
input q_in_713;
input q_in_712;
input q_in_711;
input q_in_710;
input q_in_709;
input q_in_708;
input q_in_707;
input q_in_706;
input qn_in_705;
input q_in_704;
input q_in_703;
input q_in_702;
input q_in_701;
input q_in_700;
input q_in_699;
input q_in_698;
input q_in_697;
input q_in_696;
input q_in_695;
input q_in_694;
input q_in_693;
input q_in_692;
input q_in_691;
input q_in_690;
input q_in_689;
input q_in_688;
input q_in_687;
input q_in_686;
input q_in_685;
input q_in_684;
input qn_in_683;
input q_in_682;
input qn_in_681;
input q_in_680;
input q_in_679;
input q_in_678;
input q_in_677;
input q_in_676;
input q_in_675;
input q_in_674;
input q_in_673;
input q_in_672;
input q_in_671;
input qn_in_670;
input q_in_669;
input q_in_668;
input q_in_667;
input q_in_666;
input qn_in_665;
input q_in_664;
input qn_in_663;
input q_in_662;
input q_in_661;
input q_in_660;
input q_in_659;
input q_in_658;
input q_in_657;
input q_in_656;
input q_in_655;
input q_in_654;
input q_in_653;
input q_in_652;
input q_in_651;
input qn_in_650;
input qn_in_649;
input q_in_648;
input q_in_647;
input q_in_646;
input q_in_645;
input q_in_644;
input q_in_643;
input q_in_642;
input q_in_641;
input qn_in_640;
input q_in_639;
input q_in_638;
input qn_in_637;
input q_in_636;
input q_in_635;
input q_in_634;
input q_in_633;
input q_in_632;
input q_in_631;
input q_in_630;
input q_in_629;
input q_in_628;
input q_in_627;
input q_in_626;
input q_in_625;
input q_in_624;
input q_in_623;
input q_in_622;
input q_in_621;
input q_in_620;
input q_in_619;
input q_in_618;
input q_in_617;
input q_in_616;
input q_in_615;
input q_in_614;
input q_in_613;
input q_in_612;
input q_in_611;
input qn_in_610;
input qn_in_609;
input q_in_608;
input q_in_607;
input q_in_606;
input q_in_605;
input q_in_604;
input q_in_603;
input q_in_602;
input q_in_601;
input q_in_600;
input q_in_599;
input q_in_598;
input qn_in_597;
input q_in_596;
input q_in_595;
input q_in_594;
input qn_in_593;
input q_in_592;
input q_in_591;
input q_in_590;
input qn_in_589;
input qn_in_588;
input q_in_587;
input q_in_586;
input qn_in_585;
input qn_in_584;
input q_in_583;
input q_in_582;
input q_in_581;
input q_in_580;
input q_in_579;
input q_in_578;
input q_in_577;
input q_in_576;
input q_in_575;
input q_in_574;
input q_in_573;
input q_in_572;
input q_in_571;
input q_in_570;
input q_in_569;
input qn_in_568;
input qn_in_567;
input qn_in_566;
input q_in_565;
input q_in_564;
input q_in_563;
input q_in_562;
input q_in_561;
input q_in_560;
input q_in_559;
input q_in_558;
input q_in_557;
input q_in_556;
input q_in_555;
input q_in_554;
input q_in_553;
input q_in_552;
input qn_in_551;
input q_in_550;
input qn_in_549;
input q_in_548;
input qn_in_547;
input q_in_546;
input q_in_545;
input q_in_544;
input q_in_543;
input q_in_542;
input qn_in_541;
input q_in_540;
input q_in_539;
input qn_in_538;
input q_in_537;
input q_in_536;
input qn_in_535;
input q_in_534;
input qn_in_533;
input q_in_532;
input q_in_531;
input q_in_530;
input q_in_529;
input q_in_528;
input q_in_527;
input q_in_526;
input q_in_525;
input q_in_524;
input q_in_523;
input q_in_522;
input q_in_521;
input qn_in_520;
input q_in_519;
input q_in_518;
input q_in_517;
input q_in_516;
input q_in_515;
input qn_in_514;
input qn_in_513;
input qn_in_512;
input qn_in_511;
input qn_in_510;
input qn_in_509;
input q_in_508;
input qn_in_507;
input q_in_506;
input qn_in_505;
input qn_in_504;
input qn_in_503;
input qn_in_502;
input q_in_501;
input q_in_500;
input q_in_499;
input q_in_498;
input q_in_497;
input q_in_496;
input q_in_495;
input q_in_494;
input q_in_493;
input q_in_492;
input q_in_491;
input q_in_490;
input q_in_489;
input q_in_488;
input qn_in_487;
input qn_in_486;
input q_in_485;
input q_in_484;
input q_in_483;
input q_in_482;
input q_in_481;
input qn_in_480;
input qn_in_479;
input qn_in_478;
input q_in_477;
input q_in_476;
input q_in_475;
input q_in_474;
input q_in_473;
input q_in_472;
input q_in_471;
input q_in_470;
input q_in_469;
input q_in_468;
input q_in_467;
input q_in_466;
input q_in_465;
input q_in_464;
input q_in_463;
input q_in_462;
input q_in_461;
input qn_in_460;
input qn_in_459;
input qn_in_458;
input qn_in_457;
input qn_in_456;
input qn_in_455;
input q_in_454;
input q_in_453;
input q_in_452;
input q_in_451;
input q_in_450;
input q_in_449;
input q_in_448;
input q_in_447;
input q_in_446;
input q_in_445;
input q_in_444;
input q_in_443;
input q_in_442;
input q_in_441;
input qn_in_440;
input qn_in_439;
input qn_in_438;
input qn_in_437;
input qn_in_436;
input qn_in_435;
input q_in_434;
input q_in_433;
input q_in_432;
input q_in_431;
input qn_in_430;
input qn_in_429;
input qn_in_428;
input q_in_427;
input q_in_426;
input q_in_425;
input q_in_424;
input q_in_423;
input q_in_422;
input q_in_421;
input q_in_420;
input q_in_419;
input q_in_418;
input q_in_417;
input q_in_416;
input q_in_415;
input q_in_414;
input q_in_413;
input q_in_412;
input q_in_411;
input q_in_410;
input q_in_409;
input q_in_408;
input q_in_407;
input q_in_406;
input q_in_405;
input q_in_404;
input q_in_403;
input q_in_402;
input q_in_401;
input q_in_400;
input q_in_399;
input q_in_398;
input q_in_397;
input q_in_396;
input qn_in_395;
input q_in_394;
input q_in_393;
input q_in_392;
input q_in_391;
input q_in_390;
input q_in_389;
input q_in_388;
input q_in_387;
input q_in_386;
input q_in_385;
input q_in_384;
input q_in_383;
input q_in_382;
input q_in_381;
input q_in_380;
input q_in_379;
input q_in_378;
input q_in_377;
input q_in_376;
input q_in_375;
input q_in_374;
input q_in_373;
input q_in_372;
input q_in_371;
input q_in_370;
input q_in_369;
input q_in_368;
input q_in_367;
input q_in_366;
input q_in_365;
input q_in_364;
input q_in_363;
input q_in_362;
input q_in_361;
input q_in_360;
input q_in_359;
input q_in_358;
input q_in_357;
input q_in_356;
input q_in_355;
input q_in_354;
input q_in_353;
input q_in_352;
input q_in_351;
input q_in_350;
input q_in_349;
input q_in_348;
input q_in_347;
input q_in_346;
input q_in_345;
input q_in_344;
input q_in_343;
input q_in_342;
input q_in_341;
input q_in_340;
input q_in_339;
input q_in_338;
input q_in_337;
input q_in_336;
input q_in_335;
input q_in_334;
input q_in_333;
input q_in_332;
input q_in_331;
input q_in_330;
input q_in_329;
input q_in_328;
input q_in_327;
input q_in_326;
input q_in_325;
input q_in_324;
input q_in_323;
input q_in_322;
input q_in_321;
input q_in_320;
input q_in_319;
input q_in_318;
input q_in_317;
input q_in_316;
input q_in_315;
input q_in_314;
input q_in_313;
input q_in_312;
input q_in_311;
input q_in_310;
input q_in_309;
input q_in_308;
input q_in_307;
input q_in_306;
input q_in_305;
input q_in_304;
input q_in_303;
input qn_in_302;
input qn_in_301;
input q_in_300;
input q_in_299;
input q_in_298;
input q_in_297;
input q_in_296;
input q_in_295;
input qn_in_294;
input q_in_293;
input q_in_292;
input q_in_291;
input q_in_290;
input q_in_289;
input q_in_288;
input q_in_287;
input q_in_286;
input q_in_285;
input q_in_284;
input q_in_283;
input q_in_282;
input q_in_281;
input q_in_280;
input q_in_279;
input q_in_278;
input q_in_277;
input q_in_276;
input q_in_275;
input q_in_274;
input q_in_273;
input q_in_272;
input q_in_271;
input q_in_270;
input q_in_269;
input q_in_268;
input q_in_267;
input q_in_266;
input q_in_265;
input q_in_264;
input q_in_263;
input q_in_262;
input q_in_261;
input q_in_260;
input q_in_259;
input q_in_258;
input q_in_257;
input q_in_256;
input q_in_255;
input q_in_254;
input qn_in_253;
input q_in_252;
input q_in_251;
input q_in_250;
input q_in_249;
input q_in_248;
input q_in_247;
input q_in_246;
input q_in_245;
input q_in_244;
input q_in_243;
input q_in_242;
input q_in_241;
input q_in_240;
input q_in_239;
input q_in_238;
input qn_in_237;
input q_in_236;
input q_in_235;
input q_in_234;
input q_in_233;
input q_in_232;
input q_in_231;
input q_in_230;
input qn_in_229;
input q_in_228;
input qn_in_227;
input q_in_226;
input q_in_225;
input q_in_224;
input qn_in_223;
input qn_in_222;
input q_in_221;
input q_in_220;
input q_in_219;
input q_in_218;
input q_in_217;
input q_in_216;
input q_in_215;
input q_in_214;
input q_in_213;
input q_in_212;
input q_in_211;
input q_in_210;
input q_in_209;
input q_in_208;
input q_in_207;
input q_in_206;
input q_in_205;
input q_in_204;
input q_in_203;
input q_in_202;
input q_in_201;
input q_in_200;
input q_in_199;
input q_in_198;
input q_in_197;
input q_in_196;
input q_in_195;
input q_in_194;
input q_in_193;
input q_in_192;
input q_in_191;
input q_in_190;
input q_in_189;
input q_in_188;
input q_in_187;
input q_in_186;
input q_in_185;
input q_in_184;
input q_in_183;
input q_in_182;
input q_in_181;
input q_in_180;
input qn_in_179;
input qn_in_178;
input qn_in_177;
input q_in_176;
input q_in_175;
input q_in_174;
input q_in_173;
input q_in_172;
input q_in_171;
input q_in_170;
input q_in_169;
input q_in_168;
input q_in_167;
input q_in_166;
input q_in_165;
input q_in_164;
input q_in_163;
input q_in_162;
input q_in_161;
input q_in_160;
input q_in_159;
input q_in_158;
input q_in_157;
input q_in_156;
input q_in_155;
input q_in_154;
input q_in_153;
input q_in_152;
input q_in_151;
input q_in_150;
input q_in_149;
input q_in_148;
input q_in_147;
input q_in_146;
input q_in_145;
input q_in_144;
input q_in_143;
input q_in_142;
input q_in_141;
input q_in_140;
input q_in_139;
input q_in_138;
input q_in_137;
input q_in_136;
input q_in_135;
input q_in_134;
input q_in_133;
input q_in_132;
input q_in_131;
input q_in_130;
input q_in_129;
input q_in_128;
input q_in_127;
input q_in_126;
input q_in_125;
input q_in_124;
input q_in_123;
input q_in_122;
input q_in_121;
input q_in_120;
input q_in_119;
input q_in_118;
input q_in_117;
input q_in_116;
input q_in_115;
input q_in_114;
input q_in_113;
input q_in_112;
input q_in_111;
input q_in_110;
input q_in_109;
input q_in_108;
input q_in_107;
input q_in_106;
input q_in_105;
input q_in_104;
input q_in_103;
input q_in_102;
input q_in_101;
input q_in_100;
input q_in_99;
input q_in_98;
input q_in_97;
input q_in_96;
input q_in_95;
input q_in_94;
input q_in_93;
input q_in_92;
input q_in_91;
input q_in_90;
input q_in_89;
input q_in_88;
input q_in_87;
input q_in_86;
input q_in_85;
input q_in_84;
input q_in_83;
input q_in_82;
input q_in_81;
input q_in_80;
input q_in_79;
input q_in_78;
input q_in_77;
input q_in_76;
input q_in_75;
input q_in_74;
input q_in_73;
input q_in_72;
input q_in_71;
input q_in_70;
input q_in_69;
input q_in_68;
input q_in_67;
input q_in_66;
input q_in_65;
input q_in_64;
input q_in_63;
input q_in_62;
input q_in_61;
input q_in_60;
input q_in_59;
input qn_in_58;
input q_in_57;
input q_in_56;
input q_in_55;
input q_in_54;
input q_in_53;
input q_in_52;
input q_in_51;
input q_in_50;
input q_in_49;
input q_in_48;
input q_in_47;
input q_in_46;
input q_in_45;
input q_in_44;
input q_in_43;
input q_in_42;
input q_in_41;
input q_in_40;
input q_in_39;
input q_in_38;
input q_in_37;
input q_in_36;
input q_in_35;
input q_in_34;
input q_in_33;
input q_in_32;
input q_in_31;
input q_in_30;
input q_in_29;
input q_in_28;
input q_in_27;
input q_in_26;
input q_in_25;
input q_in_24;
input q_in_23;
input q_in_22;
input q_in_21;
input q_in_20;
input q_in_19;
input q_in_18;
input q_in_17;
input q_in_16;
input qn_in_15;
input q_in_14;
input q_in_13;
input qn_in_12;
input q_in_11;
input q_in_10;
input q_in_9;
input q_in_8;
input qn_in_7;
input q_in_6;
input q_in_5;
input q_in_4;
input qn_in_3;
input q_in_2;
input q_in_1;
input q_in_1564;
input q_in_1563;
input q_in_1562;
input q_in_1561;
input q_in_1560;
input qn_in_1559;
input qn_in_1558;
input q_in_1557;
input q_in_1556;
input q_in_1555;
input q_in_1554;
input q_in_1553;
input q_in_1552;
input q_in_1551;
input q_in_1550;
input q_in_1549;
input q_in_1548;
input q_in_1547;
input q_in_1546;
input q_in_1545;
input q_in_1544;
input qn_in_1543;
input q_in_1542;
input q_in_1541;
input q_in_1540;
input q_in_1539;
input q_in_1538;
input q_in_1537;
input q_in_1536;
input q_in_1535;
input q_in_1534;
input qn_in_1533;
input q_in_1532;
input qn_in_1531;
input q_in_1530;
input q_in_1529;
input q_in_1528;
input q_in_1527;
input q_in_1526;
input q_in_1525;
input q_in_1524;
input q_in_1523;
input q_in_1522;
input q_in_1521;
input q_in_1520;
input qn_in_1519;
input q_in_1518;
input q_in_1517;
input q_in_1516;
input q_in_1515;
input q_in_1514;
input qn_in_1513;
input q_in_1512;
input q_in_1511;
input q_in_1510;
input q_in_1509;
input q_in_1508;
input q_in_1507;
input q_in_1506;
input q_in_1505;
input q_in_1504;
input q_in_1503;
input q_in_1502;
input q_in_1501;
input qn_in_1500;
input q_in_1499;
input q_in_1498;
input q_in_1497;
input q_in_1496;
input q_in_1495;
input q_in_1494;
input q_in_1493;
input q_in_1492;
input q_in_1491;
input q_in_1490;
input q_in_1489;
input q_in_1488;
input q_in_1487;
input q_in_1486;
input q_in_1485;
input q_in_1484;
input q_in_1483;
input q_in_1482;
input q_in_1481;
input q_in_1480;
input q_in_1479;
input q_in_1478;
input qn_in_1477;
input q_in_1476;
input q_in_1475;
input q_in_1474;
input q_in_1473;
input q_in_1472;
input q_in_1471;
input q_in_1470;
input q_in_1469;
input q_in_1468;
input q_in_1467;
input q_in_1466;
input q_in_1465;
input q_in_1464;
input q_in_1463;
input q_in_1462;
input q_in_1461;
input q_in_1460;
input qn_in_1459;
input q_in_1458;
input q_in_1457;
input q_in_1456;
input q_in_1455;
input q_in_1454;
input q_in_1453;
input q_in_1452;
input q_in_1451;
input q_in_1450;
input q_in_1449;
input q_in_1448;
input q_in_1447;
input qn_in_1446;
input q_in_1445;
input q_in_1444;
input q_in_1438;
input q_in_1443;
input q_in_1442;
input q_in_1441;
input q_in_1440;
input q_in_1439;
input blif_clk_net, blif_reset_net, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234;
input q_in_1437;
output d_out_1436;
output d_out_1435;
output d_out_1434;
output d_out_1433;
output d_out_1432;
output d_out_1431;
output d_out_1430;
output d_out_1429;
output d_out_1428;
output d_out_1427;
output d_out_1426;
output d_out_1425;
output d_out_1424;
output d_out_1423;
output d_out_1422;
output d_out_1421;
output d_out_1420;
output d_out_1419;
output d_out_1418;
output d_out_1417;
output d_out_1416;
output d_out_1415;
output d_out_1414;
output d_out_1413;
output d_out_1412;
output d_out_1411;
output d_out_1410;
output d_out_1409;
output d_out_1408;
output d_out_1407;
output d_out_1406;
output d_out_1405;
output d_out_1404;
output d_out_1403;
output d_out_1402;
output d_out_1401;
output d_out_1400;
output d_out_1399;
output d_out_1398;
output d_out_1397;
output d_out_1396;
output d_out_1395;
output d_out_1394;
output d_out_1393;
output d_out_1392;
output d_out_1391;
output d_out_1390;
output d_out_1389;
output d_out_1388;
output d_out_1387;
output d_out_1386;
output d_out_1385;
output d_out_1384;
output d_out_1383;
output d_out_1382;
output d_out_1381;
output d_out_1380;
output d_out_1379;
output d_out_1378;
output d_out_1377;
output d_out_1376;
output d_out_1375;
output d_out_1374;
output d_out_1373;
output d_out_1372;
output d_out_1371;
output d_out_1370;
output d_out_1369;
output d_out_1368;
output d_out_1367;
output d_out_1366;
output d_out_1365;
output d_out_1364;
output d_out_1363;
output d_out_1362;
output d_out_1361;
output d_out_1360;
output d_out_1359;
output d_out_1358;
output d_out_1357;
output d_out_1356;
output d_out_1355;
output d_out_1354;
output d_out_1353;
output d_out_1352;
output d_out_1351;
output d_out_1350;
output d_out_1349;
output d_out_1348;
output d_out_1347;
output d_out_1346;
output d_out_1345;
output d_out_1344;
output d_out_1343;
output d_out_1342;
output d_out_1341;
output d_out_1340;
output d_out_1339;
output d_out_1338;
output d_out_1337;
output d_out_1336;
output d_out_1335;
output d_out_1334;
output d_out_1333;
output d_out_1332;
output d_out_1331;
output d_out_1330;
output d_out_1329;
output d_out_1328;
output d_out_1327;
output d_out_1326;
output d_out_1325;
output d_out_1324;
output d_out_1323;
output d_out_1322;
output d_out_1321;
output d_out_1320;
output d_out_1319;
output d_out_1318;
output d_out_1317;
output d_out_1316;
output d_out_1315;
output d_out_1314;
output d_out_1313;
output d_out_1312;
output d_out_1311;
output d_out_1310;
output d_out_1309;
output d_out_1308;
output d_out_1307;
output d_out_1306;
output d_out_1305;
output d_out_1304;
output d_out_1303;
output d_out_1302;
output d_out_1301;
output d_out_1300;
output d_out_1299;
output d_out_1298;
output d_out_1297;
output d_out_1296;
output d_out_1295;
output d_out_1294;
output d_out_1293;
output d_out_1292;
output d_out_1291;
output d_out_1290;
output d_out_1289;
output d_out_1288;
output d_out_1287;
output d_out_1286;
output d_out_1285;
output d_out_1284;
output d_out_1283;
output d_out_1282;
output d_out_1281;
output d_out_1280;
output d_out_1279;
output d_out_1278;
output d_out_1277;
output d_out_1276;
output d_out_1275;
output d_out_1274;
output d_out_1273;
output d_out_1272;
output d_out_1271;
output d_out_1270;
output d_out_1269;
output d_out_1268;
output d_out_1267;
output d_out_1266;
output d_out_1265;
output d_out_1264;
output d_out_1263;
output d_out_1262;
output d_out_1261;
output d_out_1260;
output d_out_1259;
output d_out_1258;
output d_out_1257;
output d_out_1256;
output d_out_1255;
output d_out_1254;
output d_out_1253;
output d_out_1252;
output d_out_1251;
output d_out_1250;
output d_out_1249;
output d_out_1248;
output d_out_1247;
output d_out_1246;
output d_out_1245;
output d_out_1244;
output d_out_1243;
output d_out_1242;
output d_out_1241;
output d_out_1240;
output d_out_1239;
output d_out_1238;
output d_out_1237;
output d_out_1236;
output d_out_1235;
output d_out_1234;
output d_out_1233;
output d_out_1232;
output d_out_1231;
output d_out_1230;
output d_out_1229;
output d_out_1228;
output d_out_1227;
output d_out_1226;
output d_out_1225;
output d_out_1224;
output d_out_1223;
output d_out_1222;
output d_out_1221;
output d_out_1220;
output d_out_1219;
output d_out_1218;
output d_out_1217;
output d_out_1216;
output d_out_1215;
output d_out_1214;
output d_out_1213;
output d_out_1212;
output d_out_1211;
output d_out_1210;
output d_out_1209;
output d_out_1208;
output d_out_1207;
output d_out_1206;
output d_out_1205;
output d_out_1204;
output d_out_1203;
output d_out_1202;
output d_out_1201;
output d_out_1200;
output d_out_1199;
output d_out_1198;
output d_out_1197;
output d_out_1196;
output d_out_1195;
output d_out_1194;
output d_out_1193;
output d_out_1192;
output d_out_1191;
output d_out_1190;
output d_out_1189;
output d_out_1188;
output d_out_1187;
output d_out_1186;
output d_out_1185;
output d_out_1184;
output d_out_1183;
output d_out_1182;
output d_out_1181;
output d_out_1180;
output d_out_1179;
output d_out_1178;
output d_out_1177;
output d_out_1176;
output d_out_1175;
output d_out_1174;
output d_out_1173;
output d_out_1172;
output d_out_1171;
output d_out_1170;
output d_out_1169;
output d_out_1168;
output d_out_1167;
output d_out_1166;
output d_out_1165;
output d_out_1164;
output d_out_1163;
output d_out_1162;
output d_out_1161;
output d_out_1160;
output d_out_1159;
output d_out_1158;
output d_out_1157;
output d_out_1156;
output d_out_1155;
output d_out_1154;
output d_out_1153;
output d_out_1152;
output d_out_1151;
output d_out_1150;
output d_out_1149;
output d_out_1148;
output d_out_1147;
output d_out_1146;
output d_out_1145;
output d_out_1144;
output d_out_1143;
output d_out_1142;
output d_out_1141;
output d_out_1140;
output d_out_1139;
output d_out_1138;
output d_out_1137;
output d_out_1136;
output d_out_1135;
output d_out_1134;
output d_out_1133;
output d_out_1132;
output d_out_1131;
output d_out_1130;
output d_out_1129;
output d_out_1128;
output d_out_1127;
output d_out_1126;
output d_out_1125;
output d_out_1124;
output d_out_1123;
output d_out_1122;
output d_out_1121;
output d_out_1120;
output d_out_1119;
output d_out_1118;
output d_out_1117;
output d_out_1116;
output d_out_1115;
output d_out_1114;
output d_out_1113;
output d_out_1112;
output d_out_1111;
output d_out_1110;
output d_out_1109;
output d_out_1108;
output d_out_1107;
output d_out_1106;
output d_out_1105;
output d_out_1104;
output d_out_1103;
output d_out_1102;
output d_out_1101;
output d_out_1100;
output d_out_1099;
output d_out_1098;
output d_out_1097;
output d_out_1096;
output d_out_1095;
output d_out_1094;
output d_out_1093;
output d_out_1092;
output d_out_1091;
output d_out_1090;
output d_out_1089;
output d_out_1088;
output d_out_1087;
output d_out_1086;
output d_out_1085;
output d_out_1084;
output d_out_1083;
output d_out_1082;
output d_out_1081;
output d_out_1080;
output d_out_1079;
output d_out_1078;
output d_out_1077;
output d_out_1076;
output d_out_1075;
output d_out_1074;
output d_out_1073;
output d_out_1072;
output d_out_1071;
output d_out_1070;
output d_out_1069;
output d_out_1068;
output d_out_1067;
output d_out_1066;
output d_out_1065;
output d_out_1064;
output d_out_1063;
output d_out_1062;
output d_out_1061;
output d_out_1060;
output d_out_1059;
output d_out_1058;
output d_out_1057;
output d_out_1056;
output d_out_1055;
output d_out_1054;
output d_out_1053;
output d_out_1052;
output d_out_1051;
output d_out_1050;
output d_out_1049;
output d_out_1048;
output d_out_1047;
output d_out_1046;
output d_out_1045;
output d_out_1044;
output d_out_1043;
output d_out_1042;
output d_out_1041;
output d_out_1040;
output d_out_1039;
output d_out_1038;
output d_out_1037;
output d_out_1036;
output d_out_1035;
output d_out_1034;
output d_out_1033;
output d_out_1032;
output d_out_1031;
output d_out_1030;
output d_out_1029;
output d_out_1028;
output d_out_1027;
output d_out_1026;
output d_out_1025;
output d_out_1024;
output d_out_1023;
output d_out_1022;
output d_out_1021;
output d_out_1020;
output d_out_1019;
output d_out_1018;
output d_out_1017;
output d_out_1016;
output d_out_1015;
output d_out_1014;
output d_out_1013;
output d_out_1012;
output d_out_1011;
output d_out_1010;
output d_out_1009;
output d_out_1008;
output d_out_1007;
output d_out_1006;
output d_out_1005;
output d_out_1004;
output d_out_1003;
output d_out_1002;
output d_out_1001;
output d_out_1000;
output d_out_999;
output d_out_998;
output d_out_997;
output d_out_996;
output d_out_995;
output d_out_994;
output d_out_993;
output d_out_992;
output d_out_991;
output d_out_990;
output d_out_989;
output d_out_988;
output d_out_987;
output d_out_986;
output d_out_985;
output d_out_984;
output d_out_983;
output d_out_982;
output d_out_981;
output d_out_980;
output d_out_979;
output d_out_978;
output d_out_977;
output d_out_976;
output d_out_975;
output d_out_974;
output d_out_973;
output d_out_972;
output d_out_971;
output d_out_970;
output d_out_969;
output d_out_968;
output d_out_967;
output d_out_966;
output d_out_965;
output d_out_964;
output d_out_963;
output d_out_962;
output d_out_961;
output d_out_960;
output d_out_959;
output d_out_958;
output d_out_957;
output d_out_956;
output d_out_955;
output d_out_954;
output d_out_953;
output d_out_952;
output d_out_951;
output d_out_950;
output d_out_949;
output d_out_948;
output d_out_947;
output d_out_946;
output d_out_945;
output d_out_944;
output d_out_943;
output d_out_942;
output d_out_941;
output d_out_940;
output d_out_939;
output d_out_938;
output d_out_937;
output d_out_936;
output d_out_935;
output d_out_934;
output d_out_933;
output d_out_932;
output d_out_931;
output d_out_930;
output d_out_929;
output d_out_928;
output d_out_927;
output d_out_926;
output d_out_925;
output d_out_924;
output d_out_923;
output d_out_922;
output d_out_921;
output d_out_920;
output d_out_919;
output d_out_918;
output d_out_917;
output d_out_916;
output d_out_915;
output d_out_914;
output d_out_913;
output d_out_912;
output d_out_911;
output d_out_910;
output d_out_909;
output d_out_908;
output d_out_907;
output d_out_906;
output d_out_905;
output d_out_904;
output d_out_903;
output d_out_902;
output d_out_901;
output d_out_900;
output d_out_899;
output d_out_898;
output d_out_897;
output d_out_896;
output d_out_895;
output d_out_894;
output d_out_893;
output d_out_892;
output d_out_891;
output d_out_890;
output d_out_889;
output d_out_888;
output d_out_887;
output d_out_886;
output d_out_885;
output d_out_884;
output d_out_883;
output d_out_882;
output d_out_881;
output d_out_880;
output d_out_879;
output d_out_878;
output d_out_877;
output d_out_876;
output d_out_875;
output d_out_874;
output d_out_873;
output d_out_872;
output d_out_871;
output d_out_870;
output d_out_869;
output d_out_868;
output d_out_867;
output d_out_866;
output d_out_865;
output d_out_864;
output d_out_863;
output d_out_862;
output d_out_861;
output d_out_860;
output d_out_859;
output d_out_858;
output d_out_857;
output d_out_856;
output d_out_855;
output d_out_854;
output d_out_853;
output d_out_852;
output d_out_851;
output d_out_850;
output d_out_849;
output d_out_848;
output d_out_847;
output d_out_846;
output d_out_845;
output d_out_844;
output d_out_843;
output d_out_842;
output d_out_841;
output d_out_840;
output d_out_839;
output d_out_838;
output d_out_837;
output d_out_836;
output d_out_835;
output d_out_834;
output d_out_833;
output d_out_832;
output d_out_831;
output d_out_830;
output d_out_829;
output d_out_828;
output d_out_827;
output d_out_826;
output d_out_825;
output d_out_824;
output d_out_823;
output d_out_822;
output d_out_821;
output d_out_820;
output d_out_819;
output d_out_818;
output d_out_817;
output d_out_816;
output d_out_815;
output d_out_814;
output d_out_813;
output d_out_812;
output d_out_811;
output d_out_810;
output d_out_809;
output d_out_808;
output d_out_807;
output d_out_806;
output d_out_805;
output d_out_804;
output d_out_803;
output d_out_802;
output d_out_801;
output d_out_800;
output d_out_799;
output d_out_798;
output d_out_797;
output d_out_796;
output d_out_795;
output d_out_794;
output d_out_793;
output d_out_792;
output d_out_791;
output d_out_790;
output d_out_789;
output d_out_788;
output d_out_787;
output d_out_786;
output d_out_785;
output d_out_784;
output d_out_783;
output d_out_782;
output d_out_781;
output d_out_780;
output d_out_779;
output d_out_778;
output d_out_777;
output d_out_776;
output d_out_775;
output d_out_774;
output d_out_773;
output d_out_772;
output d_out_771;
output d_out_770;
output d_out_769;
output d_out_768;
output d_out_767;
output d_out_766;
output d_out_765;
output d_out_764;
output d_out_763;
output d_out_762;
output d_out_761;
output d_out_760;
output d_out_759;
output d_out_758;
output d_out_757;
output d_out_756;
output d_out_755;
output d_out_754;
output d_out_753;
output d_out_752;
output d_out_751;
output d_out_750;
output d_out_749;
output d_out_748;
output d_out_747;
output d_out_746;
output d_out_745;
output d_out_744;
output d_out_743;
output d_out_742;
output d_out_741;
output d_out_740;
output d_out_739;
output d_out_738;
output d_out_737;
output d_out_736;
output d_out_735;
output d_out_734;
output d_out_733;
output d_out_732;
output d_out_731;
output d_out_730;
output d_out_729;
output d_out_728;
output d_out_727;
output d_out_726;
output d_out_725;
output d_out_724;
output d_out_723;
output d_out_722;
output d_out_721;
output d_out_720;
output d_out_719;
output d_out_718;
output d_out_717;
output d_out_716;
output d_out_715;
output d_out_714;
output d_out_713;
output d_out_712;
output d_out_711;
output d_out_710;
output d_out_709;
output d_out_708;
output d_out_707;
output d_out_706;
output d_out_705;
output d_out_704;
output d_out_703;
output d_out_702;
output d_out_701;
output d_out_700;
output d_out_699;
output d_out_698;
output d_out_697;
output d_out_696;
output d_out_695;
output d_out_694;
output d_out_693;
output d_out_692;
output d_out_691;
output d_out_690;
output d_out_689;
output d_out_688;
output d_out_687;
output d_out_686;
output d_out_685;
output d_out_684;
output d_out_683;
output d_out_682;
output d_out_681;
output d_out_680;
output d_out_679;
output d_out_678;
output d_out_677;
output d_out_676;
output d_out_675;
output d_out_674;
output d_out_673;
output d_out_672;
output d_out_671;
output d_out_670;
output d_out_669;
output d_out_668;
output d_out_667;
output d_out_666;
output d_out_665;
output d_out_664;
output d_out_663;
output d_out_662;
output d_out_661;
output d_out_660;
output d_out_659;
output d_out_658;
output d_out_657;
output d_out_656;
output d_out_655;
output d_out_654;
output d_out_653;
output d_out_652;
output d_out_651;
output d_out_650;
output d_out_649;
output d_out_648;
output d_out_647;
output d_out_646;
output d_out_645;
output d_out_644;
output d_out_643;
output d_out_642;
output d_out_641;
output d_out_640;
output d_out_639;
output d_out_638;
output d_out_637;
output d_out_636;
output d_out_635;
output d_out_634;
output d_out_633;
output d_out_632;
output d_out_631;
output d_out_630;
output d_out_629;
output d_out_628;
output d_out_627;
output d_out_626;
output d_out_625;
output d_out_624;
output d_out_623;
output d_out_622;
output d_out_621;
output d_out_620;
output d_out_619;
output d_out_618;
output d_out_617;
output d_out_616;
output d_out_615;
output d_out_614;
output d_out_613;
output d_out_612;
output d_out_611;
output d_out_610;
output d_out_609;
output d_out_608;
output d_out_607;
output d_out_606;
output d_out_605;
output d_out_604;
output d_out_603;
output d_out_602;
output d_out_601;
output d_out_600;
output d_out_599;
output d_out_598;
output d_out_597;
output d_out_596;
output d_out_595;
output d_out_594;
output d_out_593;
output d_out_592;
output d_out_591;
output d_out_590;
output d_out_589;
output d_out_588;
output d_out_587;
output d_out_586;
output d_out_585;
output d_out_584;
output d_out_583;
output d_out_582;
output d_out_581;
output d_out_580;
output d_out_579;
output d_out_578;
output d_out_577;
output d_out_576;
output d_out_575;
output d_out_574;
output d_out_573;
output d_out_572;
output d_out_571;
output d_out_570;
output d_out_569;
output d_out_568;
output d_out_567;
output d_out_566;
output d_out_565;
output d_out_564;
output d_out_563;
output d_out_562;
output d_out_561;
output d_out_560;
output d_out_559;
output d_out_558;
output d_out_557;
output d_out_556;
output d_out_555;
output d_out_554;
output d_out_553;
output d_out_552;
output d_out_551;
output d_out_550;
output d_out_549;
output d_out_548;
output d_out_547;
output d_out_546;
output d_out_545;
output d_out_544;
output d_out_543;
output d_out_542;
output d_out_541;
output d_out_540;
output d_out_539;
output d_out_538;
output d_out_537;
output d_out_536;
output d_out_535;
output d_out_534;
output d_out_533;
output d_out_532;
output d_out_531;
output d_out_530;
output d_out_529;
output d_out_528;
output d_out_527;
output d_out_526;
output d_out_525;
output d_out_524;
output d_out_523;
output d_out_522;
output d_out_521;
output d_out_520;
output d_out_519;
output d_out_518;
output d_out_517;
output d_out_516;
output d_out_515;
output d_out_514;
output d_out_513;
output d_out_512;
output d_out_511;
output d_out_510;
output d_out_509;
output d_out_508;
output d_out_507;
output d_out_506;
output d_out_505;
output d_out_504;
output d_out_503;
output d_out_502;
output d_out_501;
output d_out_500;
output d_out_499;
output d_out_498;
output d_out_497;
output d_out_496;
output d_out_495;
output d_out_494;
output d_out_493;
output d_out_492;
output d_out_491;
output d_out_490;
output d_out_489;
output d_out_488;
output d_out_487;
output d_out_486;
output d_out_485;
output d_out_484;
output d_out_483;
output d_out_482;
output d_out_481;
output d_out_480;
output d_out_479;
output d_out_478;
output d_out_477;
output d_out_476;
output d_out_475;
output d_out_474;
output d_out_473;
output d_out_472;
output d_out_471;
output d_out_470;
output d_out_469;
output d_out_468;
output d_out_467;
output d_out_466;
output d_out_465;
output d_out_464;
output d_out_463;
output d_out_462;
output d_out_461;
output d_out_460;
output d_out_459;
output d_out_458;
output d_out_457;
output d_out_456;
output d_out_455;
output d_out_454;
output d_out_453;
output d_out_452;
output d_out_451;
output d_out_450;
output d_out_449;
output d_out_448;
output d_out_447;
output d_out_446;
output d_out_445;
output d_out_444;
output d_out_443;
output d_out_442;
output d_out_441;
output d_out_440;
output d_out_439;
output d_out_438;
output d_out_437;
output d_out_436;
output d_out_435;
output d_out_434;
output d_out_433;
output d_out_432;
output d_out_431;
output d_out_430;
output d_out_429;
output d_out_428;
output d_out_427;
output d_out_426;
output d_out_425;
output d_out_424;
output d_out_423;
output d_out_422;
output d_out_421;
output d_out_420;
output d_out_419;
output d_out_418;
output d_out_417;
output d_out_416;
output d_out_415;
output d_out_414;
output d_out_413;
output d_out_412;
output d_out_411;
output d_out_410;
output d_out_409;
output d_out_408;
output d_out_407;
output d_out_406;
output d_out_405;
output d_out_404;
output d_out_403;
output d_out_402;
output d_out_401;
output d_out_400;
output d_out_399;
output d_out_398;
output d_out_397;
output d_out_396;
output d_out_395;
output d_out_394;
output d_out_393;
output d_out_392;
output d_out_391;
output d_out_390;
output d_out_389;
output d_out_388;
output d_out_387;
output d_out_386;
output d_out_385;
output d_out_384;
output d_out_383;
output d_out_382;
output d_out_381;
output d_out_380;
output d_out_379;
output d_out_378;
output d_out_377;
output d_out_376;
output d_out_375;
output d_out_374;
output d_out_373;
output d_out_372;
output d_out_371;
output d_out_370;
output d_out_369;
output d_out_368;
output d_out_367;
output d_out_366;
output d_out_365;
output d_out_364;
output d_out_363;
output d_out_362;
output d_out_361;
output d_out_360;
output d_out_359;
output d_out_358;
output d_out_357;
output d_out_356;
output d_out_355;
output d_out_354;
output d_out_353;
output d_out_352;
output d_out_351;
output d_out_350;
output d_out_349;
output d_out_348;
output d_out_347;
output d_out_346;
output d_out_345;
output d_out_344;
output d_out_343;
output d_out_342;
output d_out_341;
output d_out_340;
output d_out_339;
output d_out_338;
output d_out_337;
output d_out_336;
output d_out_335;
output d_out_334;
output d_out_333;
output d_out_332;
output d_out_331;
output d_out_330;
output d_out_329;
output d_out_328;
output d_out_327;
output d_out_326;
output d_out_325;
output d_out_324;
output d_out_323;
output d_out_322;
output d_out_321;
output d_out_320;
output d_out_319;
output d_out_318;
output d_out_317;
output d_out_316;
output d_out_315;
output d_out_314;
output d_out_313;
output d_out_312;
output d_out_311;
output d_out_310;
output d_out_309;
output d_out_308;
output d_out_307;
output d_out_306;
output d_out_305;
output d_out_304;
output d_out_303;
output d_out_302;
output d_out_301;
output d_out_300;
output d_out_299;
output d_out_298;
output d_out_297;
output d_out_296;
output d_out_295;
output d_out_294;
output d_out_293;
output d_out_292;
output d_out_291;
output d_out_290;
output d_out_289;
output d_out_288;
output d_out_287;
output d_out_286;
output d_out_285;
output d_out_284;
output d_out_283;
output d_out_282;
output d_out_281;
output d_out_280;
output d_out_279;
output d_out_278;
output d_out_277;
output d_out_276;
output d_out_275;
output d_out_274;
output d_out_273;
output d_out_272;
output d_out_271;
output d_out_270;
output d_out_269;
output d_out_268;
output d_out_267;
output d_out_266;
output d_out_265;
output d_out_264;
output d_out_263;
output d_out_262;
output d_out_261;
output d_out_260;
output d_out_259;
output d_out_258;
output d_out_257;
output d_out_256;
output d_out_255;
output d_out_254;
output d_out_253;
output d_out_252;
output d_out_251;
output d_out_250;
output d_out_249;
output d_out_248;
output d_out_247;
output d_out_246;
output d_out_245;
output d_out_244;
output d_out_243;
output d_out_242;
output d_out_241;
output d_out_240;
output d_out_239;
output d_out_238;
output d_out_237;
output d_out_236;
output d_out_235;
output d_out_234;
output d_out_233;
output d_out_232;
output d_out_231;
output d_out_230;
output d_out_229;
output d_out_228;
output d_out_227;
output d_out_226;
output d_out_225;
output d_out_224;
output d_out_223;
output d_out_222;
output d_out_221;
output d_out_220;
output d_out_219;
output d_out_218;
output d_out_217;
output d_out_216;
output d_out_215;
output d_out_214;
output d_out_213;
output d_out_212;
output d_out_211;
output d_out_210;
output d_out_209;
output d_out_208;
output d_out_207;
output d_out_206;
output d_out_205;
output d_out_204;
output d_out_203;
output d_out_202;
output d_out_201;
output d_out_200;
output d_out_199;
output d_out_198;
output d_out_197;
output d_out_196;
output d_out_195;
output d_out_194;
output d_out_193;
output d_out_192;
output d_out_191;
output d_out_190;
output d_out_189;
output d_out_188;
output d_out_187;
output d_out_186;
output d_out_185;
output d_out_184;
output d_out_183;
output d_out_182;
output d_out_181;
output d_out_180;
output d_out_179;
output d_out_178;
output d_out_177;
output d_out_176;
output d_out_175;
output d_out_174;
output d_out_173;
output d_out_172;
output d_out_171;
output d_out_170;
output d_out_169;
output d_out_168;
output d_out_167;
output d_out_166;
output d_out_165;
output d_out_164;
output d_out_163;
output d_out_162;
output d_out_161;
output d_out_160;
output d_out_159;
output d_out_158;
output d_out_157;
output d_out_156;
output d_out_155;
output d_out_154;
output d_out_153;
output d_out_152;
output d_out_151;
output d_out_150;
output d_out_149;
output d_out_148;
output d_out_147;
output d_out_146;
output d_out_145;
output d_out_144;
output d_out_143;
output d_out_142;
output d_out_141;
output d_out_140;
output d_out_139;
output d_out_138;
output d_out_137;
output d_out_136;
output d_out_135;
output d_out_134;
output d_out_133;
output d_out_132;
output d_out_131;
output d_out_130;
output d_out_129;
output d_out_128;
output d_out_127;
output d_out_126;
output d_out_125;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_121;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_116;
output d_out_115;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_111;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_83;
output d_out_82;
output d_out_81;
output d_out_80;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_76;
output d_out_75;
output d_out_74;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_64;
output d_out_63;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_50;
output d_out_49;
output d_out_48;
output d_out_47;
output d_out_46;
output d_out_45;
output d_out_44;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_30;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_5;
output d_out_4;
output d_out_3;
output d_out_2;
output d_out_1;
output d_out_1506;
output d_out_1564;
output d_out_1563;
output d_out_1562;
output d_out_1561;
output d_out_1560;
output d_out_1559;
output d_out_1558;
output d_out_1557;
output d_out_1556;
output d_out_1555;
output d_out_1554;
output d_out_1553;
output d_out_1552;
output d_out_1551;
output d_out_1550;
output d_out_1549;
output d_out_1548;
output d_out_1547;
output d_out_1546;
output d_out_1545;
output d_out_1544;
output d_out_1543;
output d_out_1542;
output d_out_1541;
output d_out_1540;
output d_out_1539;
output d_out_1538;
output d_out_1537;
output d_out_1536;
output d_out_1535;
output d_out_1534;
output d_out_1533;
output d_out_1532;
output d_out_1531;
output d_out_1530;
output d_out_1529;
output d_out_1528;
output d_out_1527;
output d_out_1526;
output d_out_1525;
output d_out_1524;
output d_out_1523;
output d_out_1522;
output d_out_1521;
output d_out_1520;
output d_out_1519;
output d_out_1518;
output d_out_1517;
output d_out_1516;
output d_out_1515;
output d_out_1514;
output d_out_1513;
output d_out_1512;
output d_out_1511;
output d_out_1510;
output d_out_1509;
output d_out_1508;
output d_out_1507;
output d_out_1448;
output d_out_1505;
output d_out_1504;
output d_out_1503;
output d_out_1502;
output d_out_1501;
output d_out_1500;
output d_out_1499;
output d_out_1498;
output d_out_1497;
output d_out_1496;
output d_out_1495;
output d_out_1494;
output d_out_1493;
output d_out_1492;
output d_out_1491;
output d_out_1490;
output d_out_1489;
output d_out_1488;
output d_out_1487;
output d_out_1486;
output d_out_1485;
output d_out_1484;
output d_out_1483;
output d_out_1482;
output d_out_1481;
output d_out_1480;
output d_out_1479;
output d_out_1478;
output d_out_1477;
output d_out_1476;
output d_out_1475;
output d_out_1474;
output d_out_1473;
output d_out_1472;
output d_out_1471;
output d_out_1470;
output d_out_1469;
output d_out_1468;
output d_out_1467;
output d_out_1466;
output d_out_1465;
output d_out_1464;
output d_out_1463;
output d_out_1462;
output d_out_1461;
output d_out_1460;
output d_out_1459;
output d_out_1458;
output d_out_1457;
output d_out_1456;
output d_out_1455;
output d_out_1454;
output d_out_1453;
output d_out_1452;
output d_out_1451;
output d_out_1450;
output d_out_1449;
output d_out_1439;
output d_out_1447;
output d_out_1446;
output d_out_1445;
output d_out_1444;
output d_out_1443;
output d_out_1442;
output d_out_1441;
output d_out_1440;
output g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380;
output d_out_1438;
output d_out_1437;
wire n_9696, n_9697, n_9698, n_9699;
wire n_9688, n_9689, n_9690, n_9691, n_9692, n_9693, n_9694, n_9695;
wire n_9679, n_9680, n_9682, n_9683, n_9684, n_9685, n_9686, n_9687;
wire n_9671, n_9672, n_9673, n_9674, n_9675, n_9676, n_9677, n_9678;
wire n_9662, n_9663, n_9664, n_9666, n_9667, n_9668, n_9669, n_9670;
wire n_9654, n_9655, n_9656, n_9657, n_9658, n_9659, n_9660, n_9661;
wire n_9640, n_9641, n_9644, n_9647, n_9648, n_9649, n_9650, n_9651;
wire n_9626, n_9627, n_9629, n_9630, n_9631, n_9632, n_9633, n_9637;
wire n_9618, n_9619, n_9620, n_9621, n_9622, n_9623, n_9624, n_9625;
wire n_9610, n_9611, n_9612, n_9613, n_9614, n_9615, n_9616, n_9617;
wire n_9602, n_9603, n_9604, n_9605, n_9606, n_9607, n_9608, n_9609;
wire n_9593, n_9594, n_9595, n_9596, n_9597, n_9598, n_9600, n_9601;
wire n_9585, n_9586, n_9587, n_9588, n_9589, n_9590, n_9591, n_9592;
wire n_9577, n_9578, n_9579, n_9580, n_9581, n_9582, n_9583, n_9584;
wire n_9569, n_9570, n_9571, n_9572, n_9573, n_9574, n_9575, n_9576;
wire n_9557, n_9559, n_9560, n_9561, n_9562, n_9564, n_9565, n_9566;
wire n_9547, n_9548, n_9549, n_9550, n_9553, n_9554, n_9555, n_9556;
wire n_9539, n_9540, n_9541, n_9542, n_9543, n_9544, n_9545, n_9546;
wire n_9518, n_9529, n_9531, n_9533, n_9534, n_9535, n_9537, n_9538;
wire n_9508, n_9509, n_9510, n_9512, n_9514, n_9515, n_9516, n_9517;
wire n_9498, n_9499, n_9500, n_9501, n_9502, n_9503, n_9505, n_9507;
wire n_9483, n_9484, n_9485, n_9486, n_9487, n_9488, n_9489, n_9490;
wire n_9458, n_9460, n_9461, n_9462, n_9463, n_9475, n_9476, n_9477;
wire n_9441, n_9442, n_9443, n_9444, n_9447, n_9448, n_9449, n_9453;
wire n_9431, n_9432, n_9433, n_9434, n_9437, n_9438, n_9439, n_9440;
wire n_9423, n_9424, n_9425, n_9426, n_9427, n_9428, n_9429, n_9430;
wire n_9402, n_9403, n_9404, n_9418, n_9419, n_9420, n_9421, n_9422;
wire n_9393, n_9394, n_9395, n_9397, n_9398, n_9399, n_9400, n_9401;
wire n_9377, n_9378, n_9379, n_9380, n_9381, n_9382, n_9383, n_9392;
wire n_9367, n_9368, n_9369, n_9370, n_9373, n_9374, n_9375, n_9376;
wire n_9345, n_9346, n_9347, n_9361, n_9362, n_9364, n_9365, n_9366;
wire n_9320, n_9321, n_9322, n_9340, n_9341, n_9342, n_9343, n_9344;
wire n_9308, n_9309, n_9311, n_9312, n_9314, n_9315, n_9316, n_9318;
wire n_9298, n_9300, n_9301, n_9302, n_9303, n_9304, n_9305, n_9307;
wire n_9288, n_9289, n_9290, n_9292, n_9294, n_9295, n_9296, n_9297;
wire n_9271, n_9272, n_9273, n_9283, n_9284, n_9285, n_9286, n_9287;
wire n_9243, n_9254, n_9255, n_9256, n_9257, n_9267, n_9268, n_9270;
wire n_9233, n_9234, n_9235, n_9236, n_9237, n_9238, n_9240, n_9242;
wire n_9224, n_9225, n_9226, n_9227, n_9229, n_9230, n_9231, n_9232;
wire n_9214, n_9215, n_9216, n_9217, n_9219, n_9220, n_9222, n_9223;
wire n_9199, n_9200, n_9202, n_9208, n_9209, n_9210, n_9211, n_9212;
wire n_9144, n_9147, n_9148, n_9188, n_9192, n_9195, n_9196, n_9198;
wire n_9116, n_9119, n_9129, n_9136, n_9137, n_9139, n_9140, n_9141;
wire n_9104, n_9106, n_9109, n_9110, n_9111, n_9112, n_9113, n_9114;
wire n_9086, n_9087, n_9088, n_9089, n_9090, n_9091, n_9093, n_9101;
wire n_9076, n_9077, n_9079, n_9080, n_9081, n_9083, n_9084, n_9085;
wire n_9066, n_9067, n_9070, n_9071, n_9072, n_9073, n_9074, n_9075;
wire n_9057, n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9065;
wire n_9049, n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056;
wire n_9037, n_9038, n_9040, n_9041, n_9042, n_9043, n_9044, n_9048;
wire n_9006, n_9010, n_9011, n_9014, n_9021, n_9024, n_9025, n_9036;
wire n_8995, n_8998, n_8999, n_9000, n_9001, n_9002, n_9003, n_9005;
wire n_8984, n_8985, n_8986, n_8987, n_8988, n_8990, n_8993, n_8994;
wire n_8964, n_8965, n_8967, n_8968, n_8979, n_8980, n_8982, n_8983;
wire n_8954, n_8956, n_8957, n_8958, n_8960, n_8961, n_8962, n_8963;
wire n_8943, n_8944, n_8945, n_8946, n_8948, n_8949, n_8951, n_8953;
wire n_8935, n_8936, n_8937, n_8938, n_8939, n_8940, n_8941, n_8942;
wire n_8911, n_8912, n_8913, n_8924, n_8929, n_8931, n_8933, n_8934;
wire n_8887, n_8888, n_8891, n_8892, n_8894, n_8901, n_8905, n_8909;
wire n_8878, n_8879, n_8880, n_8881, n_8882, n_8884, n_8885, n_8886;
wire n_8865, n_8866, n_8867, n_8868, n_8873, n_8874, n_8876, n_8877;
wire n_8839, n_8841, n_8842, n_8843, n_8844, n_8861, n_8862, n_8863;
wire n_8831, n_8832, n_8833, n_8834, n_8835, n_8836, n_8837, n_8838;
wire n_8806, n_8809, n_8810, n_8823, n_8824, n_8825, n_8829, n_8830;
wire n_8789, n_8790, n_8791, n_8792, n_8793, n_8794, n_8796, n_8805;
wire n_8778, n_8781, n_8782, n_8783, n_8784, n_8785, n_8786, n_8788;
wire n_8767, n_8768, n_8769, n_8770, n_8771, n_8774, n_8775, n_8777;
wire n_8757, n_8758, n_8759, n_8760, n_8761, n_8762, n_8764, n_8766;
wire n_8733, n_8734, n_8736, n_8740, n_8741, n_8743, n_8747, n_8756;
wire n_8723, n_8724, n_8725, n_8726, n_8727, n_8730, n_8731, n_8732;
wire n_8707, n_8708, n_8710, n_8718, n_8719, n_8720, n_8721, n_8722;
wire n_8699, n_8700, n_8701, n_8702, n_8703, n_8704, n_8705, n_8706;
wire n_8687, n_8688, n_8689, n_8690, n_8693, n_8694, n_8697, n_8698;
wire n_8655, n_8656, n_8663, n_8667, n_8678, n_8682, n_8685, n_8686;
wire n_8643, n_8644, n_8646, n_8647, n_8649, n_8650, n_8652, n_8653;
wire n_8632, n_8633, n_8634, n_8635, n_8636, n_8639, n_8640, n_8641;
wire n_8622, n_8623, n_8625, n_8626, n_8628, n_8629, n_8630, n_8631;
wire n_8590, n_8591, n_8597, n_8598, n_8607, n_8608, n_8609, n_8621;
wire n_8574, n_8575, n_8576, n_8578, n_8582, n_8583, n_8584, n_8585;
wire n_8552, n_8557, n_8563, n_8566, n_8567, n_8570, n_8571, n_8573;
wire n_8533, n_8534, n_8540, n_8541, n_8542, n_8548, n_8550, n_8551;
wire n_8494, n_8495, n_8497, n_8498, n_8499, n_8515, n_8517, n_8527;
wire n_8485, n_8486, n_8487, n_8488, n_8489, n_8490, n_8492, n_8493;
wire n_8471, n_8472, n_8476, n_8478, n_8481, n_8482, n_8483, n_8484;
wire n_8456, n_8457, n_8459, n_8460, n_8461, n_8462, n_8463, n_8464;
wire n_8424, n_8427, n_8432, n_8437, n_8445, n_8446, n_8454, n_8455;
wire n_8410, n_8411, n_8413, n_8419, n_8420, n_8421, n_8422, n_8423;
wire n_8398, n_8400, n_8401, n_8402, n_8403, n_8404, n_8408, n_8409;
wire n_8389, n_8391, n_8392, n_8393, n_8394, n_8395, n_8396, n_8397;
wire n_8376, n_8377, n_8379, n_8380, n_8383, n_8386, n_8387, n_8388;
wire n_8353, n_8355, n_8357, n_8362, n_8365, n_8366, n_8367, n_8368;
wire n_8278, n_8280, n_8281, n_8305, n_8326, n_8339, n_8346, n_8351;
wire n_8270, n_8271, n_8272, n_8273, n_8274, n_8275, n_8276, n_8277;
wire n_8262, n_8263, n_8264, n_8265, n_8266, n_8267, n_8268, n_8269;
wire n_8253, n_8254, n_8255, n_8256, n_8257, n_8258, n_8259, n_8260;
wire n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248;
wire n_8225, n_8226, n_8227, n_8228, n_8229, n_8230, n_8234, n_8236;
wire n_8215, n_8216, n_8217, n_8218, n_8219, n_8220, n_8221, n_8222;
wire n_8187, n_8189, n_8191, n_8206, n_8207, n_8208, n_8210, n_8211;
wire n_8172, n_8173, n_8174, n_8175, n_8176, n_8178, n_8180, n_8183;
wire n_8164, n_8165, n_8166, n_8167, n_8168, n_8169, n_8170, n_8171;
wire n_8156, n_8157, n_8158, n_8159, n_8160, n_8161, n_8162, n_8163;
wire n_8148, n_8149, n_8150, n_8151, n_8152, n_8153, n_8154, n_8155;
wire n_8140, n_8141, n_8142, n_8143, n_8144, n_8145, n_8146, n_8147;
wire n_8132, n_8133, n_8134, n_8135, n_8136, n_8137, n_8138, n_8139;
wire n_8124, n_8125, n_8126, n_8127, n_8128, n_8129, n_8130, n_8131;
wire n_8116, n_8117, n_8118, n_8119, n_8120, n_8121, n_8122, n_8123;
wire n_8108, n_8109, n_8110, n_8111, n_8112, n_8113, n_8114, n_8115;
wire n_8100, n_8101, n_8102, n_8103, n_8104, n_8105, n_8106, n_8107;
wire n_8087, n_8088, n_8090, n_8092, n_8096, n_8097, n_8098, n_8099;
wire n_8078, n_8079, n_8080, n_8082, n_8083, n_8084, n_8085, n_8086;
wire n_8070, n_8071, n_8072, n_8073, n_8074, n_8075, n_8076, n_8077;
wire n_8062, n_8063, n_8064, n_8065, n_8066, n_8067, n_8068, n_8069;
wire n_8053, n_8054, n_8055, n_8056, n_8057, n_8058, n_8059, n_8060;
wire n_8044, n_8045, n_8047, n_8048, n_8049, n_8050, n_8051, n_8052;
wire n_8029, n_8034, n_8036, n_8037, n_8038, n_8039, n_8040, n_8043;
wire n_8019, n_8020, n_8021, n_8022, n_8023, n_8024, n_8025, n_8028;
wire n_8008, n_8009, n_8010, n_8011, n_8012, n_8014, n_8017, n_8018;
wire n_8000, n_8001, n_8002, n_8003, n_8004, n_8005, n_8006, n_8007;
wire n_7992, n_7993, n_7994, n_7995, n_7996, n_7997, n_7998, n_7999;
wire n_7982, n_7983, n_7984, n_7985, n_7986, n_7987, n_7988, n_7990;
wire n_7972, n_7973, n_7974, n_7976, n_7977, n_7978, n_7979, n_7981;
wire n_7962, n_7963, n_7965, n_7966, n_7968, n_7969, n_7970, n_7971;
wire n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960, n_7961;
wire n_7946, n_7947, n_7948, n_7949, n_7950, n_7951, n_7952, n_7953;
wire n_7938, n_7939, n_7940, n_7941, n_7942, n_7943, n_7944, n_7945;
wire n_7927, n_7928, n_7929, n_7930, n_7932, n_7935, n_7936, n_7937;
wire n_7919, n_7920, n_7921, n_7922, n_7923, n_7924, n_7925, n_7926;
wire n_7911, n_7912, n_7913, n_7914, n_7915, n_7916, n_7917, n_7918;
wire n_7900, n_7901, n_7902, n_7905, n_7906, n_7908, n_7909, n_7910;
wire n_7892, n_7893, n_7894, n_7895, n_7896, n_7897, n_7898, n_7899;
wire n_7883, n_7884, n_7885, n_7886, n_7888, n_7889, n_7890, n_7891;
wire n_7865, n_7866, n_7868, n_7871, n_7876, n_7880, n_7881, n_7882;
wire n_7856, n_7857, n_7858, n_7860, n_7861, n_7862, n_7863, n_7864;
wire n_7847, n_7848, n_7849, n_7851, n_7852, n_7853, n_7854, n_7855;
wire n_7839, n_7840, n_7841, n_7842, n_7843, n_7844, n_7845, n_7846;
wire n_7831, n_7832, n_7833, n_7834, n_7835, n_7836, n_7837, n_7838;
wire n_7823, n_7824, n_7825, n_7826, n_7827, n_7828, n_7829, n_7830;
wire n_7809, n_7811, n_7812, n_7816, n_7817, n_7819, n_7821, n_7822;
wire n_7797, n_7800, n_7801, n_7802, n_7805, n_7806, n_7807, n_7808;
wire n_7788, n_7789, n_7790, n_7791, n_7792, n_7793, n_7794, n_7795;
wire n_7779, n_7780, n_7781, n_7782, n_7784, n_7785, n_7786, n_7787;
wire n_7762, n_7764, n_7768, n_7769, n_7771, n_7772, n_7773, n_7778;
wire n_7749, n_7750, n_7751, n_7753, n_7756, n_7757, n_7759, n_7760;
wire n_7741, n_7742, n_7743, n_7744, n_7745, n_7746, n_7747, n_7748;
wire n_7733, n_7734, n_7735, n_7736, n_7737, n_7738, n_7739, n_7740;
wire n_7713, n_7714, n_7722, n_7723, n_7724, n_7726, n_7730, n_7732;
wire n_7705, n_7706, n_7707, n_7708, n_7709, n_7710, n_7711, n_7712;
wire n_7696, n_7697, n_7698, n_7700, n_7701, n_7702, n_7703, n_7704;
wire n_7686, n_7687, n_7689, n_7691, n_7692, n_7693, n_7694, n_7695;
wire n_7676, n_7677, n_7678, n_7679, n_7680, n_7682, n_7684, n_7685;
wire n_7665, n_7666, n_7668, n_7669, n_7671, n_7673, n_7674, n_7675;
wire n_7653, n_7654, n_7655, n_7656, n_7657, n_7659, n_7660, n_7663;
wire n_7645, n_7646, n_7647, n_7648, n_7649, n_7650, n_7651, n_7652;
wire n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7642, n_7643;
wire n_7626, n_7627, n_7629, n_7630, n_7631, n_7632, n_7633, n_7634;
wire n_7618, n_7619, n_7620, n_7621, n_7622, n_7623, n_7624, n_7625;
wire n_7609, n_7611, n_7612, n_7613, n_7614, n_7615, n_7616, n_7617;
wire n_7595, n_7596, n_7599, n_7600, n_7601, n_7605, n_7607, n_7608;
wire n_7586, n_7587, n_7588, n_7589, n_7590, n_7591, n_7593, n_7594;
wire n_7575, n_7576, n_7577, n_7578, n_7579, n_7581, n_7582, n_7583;
wire n_7563, n_7564, n_7565, n_7566, n_7567, n_7568, n_7569, n_7571;
wire n_7554, n_7555, n_7556, n_7558, n_7559, n_7560, n_7561, n_7562;
wire n_7540, n_7543, n_7545, n_7546, n_7548, n_7550, n_7552, n_7553;
wire n_7530, n_7531, n_7532, n_7533, n_7536, n_7537, n_7538, n_7539;
wire n_7521, n_7523, n_7524, n_7525, n_7526, n_7527, n_7528, n_7529;
wire n_7505, n_7506, n_7507, n_7508, n_7511, n_7517, n_7518, n_7519;
wire n_7492, n_7493, n_7494, n_7495, n_7496, n_7498, n_7499, n_7504;
wire n_7483, n_7484, n_7485, n_7486, n_7488, n_7489, n_7490, n_7491;
wire n_7471, n_7472, n_7474, n_7475, n_7476, n_7477, n_7478, n_7482;
wire n_7461, n_7462, n_7463, n_7464, n_7465, n_7466, n_7469, n_7470;
wire n_7453, n_7454, n_7455, n_7456, n_7457, n_7458, n_7459, n_7460;
wire n_7441, n_7442, n_7443, n_7444, n_7445, n_7448, n_7451, n_7452;
wire n_7429, n_7430, n_7431, n_7432, n_7433, n_7435, n_7438, n_7439;
wire n_7417, n_7418, n_7419, n_7420, n_7421, n_7422, n_7423, n_7426;
wire n_7407, n_7410, n_7411, n_7412, n_7413, n_7414, n_7415, n_7416;
wire n_7389, n_7392, n_7395, n_7397, n_7398, n_7399, n_7403, n_7406;
wire n_7379, n_7380, n_7381, n_7384, n_7385, n_7386, n_7387, n_7388;
wire n_7370, n_7371, n_7372, n_7373, n_7374, n_7375, n_7376, n_7377;
wire n_7359, n_7360, n_7361, n_7362, n_7363, n_7365, n_7366, n_7369;
wire n_7347, n_7348, n_7349, n_7351, n_7353, n_7354, n_7355, n_7358;
wire n_7338, n_7339, n_7341, n_7342, n_7343, n_7344, n_7345, n_7346;
wire n_7330, n_7331, n_7332, n_7333, n_7334, n_7335, n_7336, n_7337;
wire n_7321, n_7322, n_7324, n_7325, n_7326, n_7327, n_7328, n_7329;
wire n_7312, n_7314, n_7315, n_7316, n_7317, n_7318, n_7319, n_7320;
wire n_7303, n_7304, n_7306, n_7307, n_7308, n_7309, n_7310, n_7311;
wire n_7291, n_7292, n_7293, n_7295, n_7296, n_7297, n_7299, n_7301;
wire n_7282, n_7283, n_7284, n_7285, n_7286, n_7287, n_7288, n_7289;
wire n_7274, n_7275, n_7276, n_7277, n_7278, n_7279, n_7280, n_7281;
wire n_7266, n_7267, n_7268, n_7269, n_7270, n_7271, n_7272, n_7273;
wire n_7256, n_7257, n_7258, n_7260, n_7261, n_7262, n_7263, n_7264;
wire n_7241, n_7242, n_7246, n_7247, n_7249, n_7251, n_7252, n_7253;
wire n_7230, n_7232, n_7233, n_7235, n_7237, n_7238, n_7239, n_7240;
wire n_7222, n_7223, n_7224, n_7225, n_7226, n_7227, n_7228, n_7229;
wire n_7209, n_7212, n_7213, n_7214, n_7215, n_7217, n_7218, n_7221;
wire n_7199, n_7200, n_7201, n_7202, n_7203, n_7204, n_7205, n_7208;
wire n_7189, n_7190, n_7193, n_7194, n_7195, n_7196, n_7197, n_7198;
wire n_7179, n_7182, n_7183, n_7184, n_7185, n_7186, n_7187, n_7188;
wire n_7168, n_7171, n_7172, n_7173, n_7174, n_7176, n_7177, n_7178;
wire n_7156, n_7157, n_7160, n_7162, n_7163, n_7164, n_7165, n_7166;
wire n_7147, n_7148, n_7149, n_7150, n_7152, n_7153, n_7154, n_7155;
wire n_7139, n_7140, n_7141, n_7142, n_7143, n_7144, n_7145, n_7146;
wire n_7130, n_7131, n_7132, n_7134, n_7135, n_7136, n_7137, n_7138;
wire n_7119, n_7120, n_7123, n_7124, n_7125, n_7126, n_7127, n_7129;
wire n_7109, n_7110, n_7112, n_7113, n_7114, n_7115, n_7116, n_7118;
wire n_7101, n_7102, n_7103, n_7104, n_7105, n_7106, n_7107, n_7108;
wire n_7090, n_7091, n_7093, n_7094, n_7095, n_7096, n_7099, n_7100;
wire n_7079, n_7080, n_7082, n_7083, n_7085, n_7087, n_7088, n_7089;
wire n_7068, n_7069, n_7070, n_7072, n_7073, n_7074, n_7077, n_7078;
wire n_7058, n_7060, n_7061, n_7062, n_7064, n_7065, n_7066, n_7067;
wire n_7045, n_7046, n_7047, n_7048, n_7049, n_7050, n_7054, n_7057;
wire n_7031, n_7032, n_7036, n_7038, n_7039, n_7042, n_7043, n_7044;
wire n_7022, n_7023, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030;
wire n_7014, n_7015, n_7016, n_7017, n_7018, n_7019, n_7020, n_7021;
wire n_7005, n_7007, n_7008, n_7009, n_7010, n_7011, n_7012, n_7013;
wire n_6994, n_6995, n_6996, n_6999, n_7000, n_7002, n_7003, n_7004;
wire n_6982, n_6985, n_6986, n_6987, n_6988, n_6989, n_6991, n_6992;
wire n_6969, n_6970, n_6971, n_6972, n_6974, n_6975, n_6978, n_6979;
wire n_6959, n_6960, n_6962, n_6963, n_6965, n_6966, n_6967, n_6968;
wire n_6949, n_6950, n_6951, n_6952, n_6954, n_6955, n_6956, n_6958;
wire n_6941, n_6942, n_6943, n_6944, n_6945, n_6946, n_6947, n_6948;
wire n_6933, n_6934, n_6935, n_6936, n_6937, n_6938, n_6939, n_6940;
wire n_6920, n_6921, n_6924, n_6925, n_6926, n_6929, n_6931, n_6932;
wire n_6909, n_6911, n_6913, n_6914, n_6915, n_6916, n_6917, n_6918;
wire n_6901, n_6902, n_6903, n_6904, n_6905, n_6906, n_6907, n_6908;
wire n_6892, n_6893, n_6894, n_6895, n_6896, n_6897, n_6899, n_6900;
wire n_6884, n_6885, n_6886, n_6887, n_6888, n_6889, n_6890, n_6891;
wire n_6873, n_6874, n_6875, n_6877, n_6880, n_6881, n_6882, n_6883;
wire n_6865, n_6866, n_6867, n_6868, n_6869, n_6870, n_6871, n_6872;
wire n_6853, n_6855, n_6859, n_6860, n_6861, n_6862, n_6863, n_6864;
wire n_6844, n_6845, n_6846, n_6847, n_6848, n_6849, n_6850, n_6851;
wire n_6830, n_6831, n_6832, n_6833, n_6836, n_6837, n_6841, n_6843;
wire n_6820, n_6821, n_6822, n_6823, n_6824, n_6826, n_6827, n_6828;
wire n_6810, n_6811, n_6812, n_6813, n_6814, n_6815, n_6816, n_6818;
wire n_6802, n_6803, n_6804, n_6805, n_6806, n_6807, n_6808, n_6809;
wire n_6794, n_6795, n_6796, n_6797, n_6798, n_6799, n_6800, n_6801;
wire n_6785, n_6786, n_6787, n_6788, n_6790, n_6791, n_6792, n_6793;
wire n_6769, n_6772, n_6773, n_6774, n_6775, n_6776, n_6778, n_6782;
wire n_6753, n_6755, n_6756, n_6759, n_6761, n_6762, n_6763, n_6765;
wire n_6743, n_6744, n_6745, n_6746, n_6747, n_6748, n_6749, n_6752;
wire n_6735, n_6736, n_6737, n_6738, n_6739, n_6740, n_6741, n_6742;
wire n_6724, n_6726, n_6728, n_6729, n_6730, n_6731, n_6732, n_6734;
wire n_6713, n_6715, n_6718, n_6719, n_6720, n_6721, n_6722, n_6723;
wire n_6705, n_6706, n_6707, n_6708, n_6709, n_6710, n_6711, n_6712;
wire n_6693, n_6696, n_6697, n_6698, n_6700, n_6702, n_6703, n_6704;
wire n_6685, n_6686, n_6687, n_6688, n_6689, n_6690, n_6691, n_6692;
wire n_6672, n_6673, n_6674, n_6678, n_6680, n_6682, n_6683, n_6684;
wire n_6664, n_6665, n_6666, n_6667, n_6668, n_6669, n_6670, n_6671;
wire n_6656, n_6657, n_6658, n_6659, n_6660, n_6661, n_6662, n_6663;
wire n_6648, n_6649, n_6650, n_6651, n_6652, n_6653, n_6654, n_6655;
wire n_6640, n_6641, n_6642, n_6643, n_6644, n_6645, n_6646, n_6647;
wire n_6631, n_6632, n_6633, n_6634, n_6635, n_6636, n_6638, n_6639;
wire n_6623, n_6624, n_6625, n_6626, n_6627, n_6628, n_6629, n_6630;
wire n_6611, n_6612, n_6616, n_6618, n_6619, n_6620, n_6621, n_6622;
wire n_6599, n_6600, n_6602, n_6603, n_6606, n_6607, n_6609, n_6610;
wire n_6583, n_6589, n_6592, n_6593, n_6594, n_6595, n_6597, n_6598;
wire n_6574, n_6575, n_6576, n_6577, n_6578, n_6579, n_6581, n_6582;
wire n_6566, n_6567, n_6568, n_6569, n_6570, n_6571, n_6572, n_6573;
wire n_6556, n_6557, n_6558, n_6560, n_6561, n_6562, n_6563, n_6565;
wire n_6547, n_6548, n_6550, n_6551, n_6552, n_6553, n_6554, n_6555;
wire n_6539, n_6540, n_6541, n_6542, n_6543, n_6544, n_6545, n_6546;
wire n_6530, n_6531, n_6532, n_6533, n_6534, n_6535, n_6537, n_6538;
wire n_6520, n_6521, n_6522, n_6525, n_6526, n_6527, n_6528, n_6529;
wire n_6510, n_6511, n_6512, n_6513, n_6516, n_6517, n_6518, n_6519;
wire n_6501, n_6502, n_6503, n_6504, n_6505, n_6507, n_6508, n_6509;
wire n_6493, n_6494, n_6495, n_6496, n_6497, n_6498, n_6499, n_6500;
wire n_6484, n_6485, n_6486, n_6487, n_6488, n_6489, n_6490, n_6492;
wire n_6475, n_6476, n_6478, n_6479, n_6480, n_6481, n_6482, n_6483;
wire n_6465, n_6466, n_6467, n_6469, n_6470, n_6472, n_6473, n_6474;
wire n_6457, n_6458, n_6459, n_6460, n_6461, n_6462, n_6463, n_6464;
wire n_6448, n_6450, n_6451, n_6452, n_6453, n_6454, n_6455, n_6456;
wire n_6437, n_6438, n_6439, n_6440, n_6441, n_6442, n_6443, n_6445;
wire n_6427, n_6429, n_6430, n_6431, n_6432, n_6433, n_6435, n_6436;
wire n_6418, n_6419, n_6420, n_6421, n_6422, n_6423, n_6424, n_6425;
wire n_6407, n_6409, n_6410, n_6412, n_6413, n_6414, n_6416, n_6417;
wire n_6398, n_6399, n_6400, n_6402, n_6403, n_6404, n_6405, n_6406;
wire n_6384, n_6391, n_6392, n_6393, n_6394, n_6395, n_6396, n_6397;
wire n_6374, n_6375, n_6376, n_6377, n_6378, n_6379, n_6380, n_6381;
wire n_6365, n_6366, n_6367, n_6368, n_6370, n_6371, n_6372, n_6373;
wire n_6354, n_6356, n_6357, n_6358, n_6359, n_6361, n_6362, n_6363;
wire n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351, n_6353;
wire n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343, n_6344;
wire n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336;
wire n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327, n_6328;
wire n_6308, n_6310, n_6311, n_6314, n_6315, n_6316, n_6319, n_6320;
wire n_6296, n_6299, n_6300, n_6302, n_6303, n_6304, n_6305, n_6307;
wire n_6279, n_6280, n_6282, n_6284, n_6286, n_6287, n_6288, n_6289;
wire n_6271, n_6272, n_6273, n_6274, n_6275, n_6276, n_6277, n_6278;
wire n_6263, n_6264, n_6265, n_6266, n_6267, n_6268, n_6269, n_6270;
wire n_6252, n_6253, n_6254, n_6255, n_6256, n_6260, n_6261, n_6262;
wire n_6240, n_6241, n_6243, n_6245, n_6246, n_6247, n_6250, n_6251;
wire n_6231, n_6232, n_6233, n_6234, n_6236, n_6237, n_6238, n_6239;
wire n_6220, n_6221, n_6222, n_6223, n_6226, n_6227, n_6228, n_6229;
wire n_6212, n_6213, n_6214, n_6215, n_6216, n_6217, n_6218, n_6219;
wire n_6203, n_6204, n_6205, n_6206, n_6207, n_6208, n_6209, n_6210;
wire n_6195, n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202;
wire n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192, n_6193;
wire n_6174, n_6177, n_6179, n_6180, n_6181, n_6182, n_6183, n_6185;
wire n_6165, n_6166, n_6167, n_6168, n_6170, n_6171, n_6172, n_6173;
wire n_6156, n_6157, n_6158, n_6159, n_6161, n_6162, n_6163, n_6164;
wire n_6148, n_6149, n_6150, n_6151, n_6152, n_6153, n_6154, n_6155;
wire n_6136, n_6137, n_6138, n_6139, n_6140, n_6141, n_6144, n_6145;
wire n_6123, n_6124, n_6127, n_6128, n_6131, n_6132, n_6133, n_6134;
wire n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120;
wire n_6105, n_6106, n_6107, n_6108, n_6109, n_6110, n_6111, n_6112;
wire n_6097, n_6098, n_6099, n_6100, n_6101, n_6102, n_6103, n_6104;
wire n_6083, n_6086, n_6089, n_6091, n_6092, n_6093, n_6094, n_6096;
wire n_6073, n_6074, n_6075, n_6076, n_6077, n_6078, n_6079, n_6080;
wire n_6065, n_6066, n_6067, n_6068, n_6069, n_6070, n_6071, n_6072;
wire n_6053, n_6054, n_6055, n_6056, n_6058, n_6062, n_6063, n_6064;
wire n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052;
wire n_6036, n_6037, n_6039, n_6040, n_6041, n_6042, n_6043, n_6044;
wire n_6025, n_6026, n_6027, n_6028, n_6032, n_6033, n_6034, n_6035;
wire n_6009, n_6010, n_6011, n_6012, n_6013, n_6014, n_6019, n_6023;
wire n_6001, n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008;
wire n_5993, n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000;
wire n_5984, n_5985, n_5987, n_5988, n_5989, n_5990, n_5991, n_5992;
wire n_5973, n_5974, n_5976, n_5979, n_5980, n_5981, n_5982, n_5983;
wire n_5963, n_5964, n_5965, n_5966, n_5967, n_5969, n_5970, n_5972;
wire n_5948, n_5949, n_5950, n_5956, n_5957, n_5958, n_5961, n_5962;
wire n_5937, n_5938, n_5939, n_5940, n_5941, n_5942, n_5943, n_5947;
wire n_5927, n_5929, n_5930, n_5932, n_5933, n_5934, n_5935, n_5936;
wire n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5925, n_5926;
wire n_5901, n_5902, n_5905, n_5906, n_5907, n_5908, n_5913, n_5915;
wire n_5890, n_5891, n_5892, n_5893, n_5894, n_5897, n_5898, n_5900;
wire n_5882, n_5883, n_5884, n_5885, n_5886, n_5887, n_5888, n_5889;
wire n_5874, n_5875, n_5876, n_5877, n_5878, n_5879, n_5880, n_5881;
wire n_5864, n_5865, n_5866, n_5867, n_5868, n_5870, n_5871, n_5872;
wire n_5852, n_5853, n_5854, n_5855, n_5856, n_5857, n_5862, n_5863;
wire n_5843, n_5844, n_5846, n_5847, n_5848, n_5849, n_5850, n_5851;
wire n_5832, n_5834, n_5836, n_5837, n_5838, n_5839, n_5841, n_5842;
wire n_5820, n_5821, n_5822, n_5824, n_5825, n_5826, n_5827, n_5828;
wire n_5806, n_5808, n_5809, n_5810, n_5811, n_5817, n_5818, n_5819;
wire n_5797, n_5798, n_5799, n_5800, n_5801, n_5803, n_5804, n_5805;
wire n_5781, n_5782, n_5783, n_5785, n_5786, n_5787, n_5788, n_5796;
wire n_5770, n_5773, n_5774, n_5775, n_5777, n_5778, n_5779, n_5780;
wire n_5761, n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768;
wire n_5753, n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760;
wire n_5738, n_5741, n_5742, n_5743, n_5748, n_5749, n_5750, n_5751;
wire n_5728, n_5730, n_5731, n_5732, n_5734, n_5735, n_5736, n_5737;
wire n_5715, n_5716, n_5717, n_5719, n_5722, n_5723, n_5725, n_5726;
wire n_5705, n_5706, n_5707, n_5708, n_5709, n_5712, n_5713, n_5714;
wire n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703, n_5704;
wire n_5685, n_5686, n_5687, n_5690, n_5692, n_5693, n_5694, n_5696;
wire n_5668, n_5669, n_5670, n_5673, n_5679, n_5680, n_5681, n_5683;
wire n_5656, n_5658, n_5660, n_5663, n_5664, n_5665, n_5666, n_5667;
wire n_5637, n_5638, n_5644, n_5647, n_5651, n_5653, n_5654, n_5655;
wire n_5616, n_5617, n_5624, n_5625, n_5628, n_5632, n_5633, n_5634;
wire n_5605, n_5606, n_5609, n_5610, n_5612, n_5613, n_5614, n_5615;
wire n_5592, n_5593, n_5594, n_5595, n_5600, n_5602, n_5603, n_5604;
wire n_5583, n_5584, n_5585, n_5586, n_5587, n_5589, n_5590, n_5591;
wire n_5573, n_5574, n_5575, n_5576, n_5577, n_5578, n_5580, n_5581;
wire n_5561, n_5562, n_5565, n_5566, n_5567, n_5568, n_5569, n_5570;
wire n_5552, n_5553, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560;
wire n_5541, n_5543, n_5545, n_5547, n_5548, n_5549, n_5550, n_5551;
wire n_5527, n_5528, n_5529, n_5530, n_5531, n_5532, n_5533, n_5539;
wire n_5515, n_5516, n_5518, n_5521, n_5522, n_5523, n_5524, n_5526;
wire n_5506, n_5507, n_5508, n_5510, n_5511, n_5512, n_5513, n_5514;
wire n_5494, n_5498, n_5500, n_5501, n_5502, n_5503, n_5504, n_5505;
wire n_5481, n_5482, n_5485, n_5486, n_5489, n_5491, n_5492, n_5493;
wire n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5479, n_5480;
wire n_5445, n_5446, n_5460, n_5462, n_5463, n_5465, n_5466, n_5469;
wire n_5429, n_5431, n_5433, n_5434, n_5435, n_5438, n_5439, n_5444;
wire n_5417, n_5418, n_5419, n_5420, n_5422, n_5423, n_5424, n_5425;
wire n_5409, n_5410, n_5411, n_5412, n_5413, n_5414, n_5415, n_5416;
wire n_5384, n_5385, n_5386, n_5387, n_5405, n_5406, n_5407, n_5408;
wire n_5374, n_5376, n_5378, n_5379, n_5380, n_5381, n_5382, n_5383;
wire n_5359, n_5365, n_5367, n_5368, n_5369, n_5371, n_5372, n_5373;
wire n_5350, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358;
wire n_5342, n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5349;
wire n_5331, n_5332, n_5334, n_5335, n_5336, n_5337, n_5338, n_5341;
wire n_5322, n_5323, n_5324, n_5325, n_5326, n_5327, n_5329, n_5330;
wire n_5313, n_5314, n_5316, n_5317, n_5318, n_5319, n_5320, n_5321;
wire n_5299, n_5300, n_5303, n_5307, n_5309, n_5310, n_5311, n_5312;
wire n_5291, n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298;
wire n_5281, n_5282, n_5283, n_5285, n_5286, n_5287, n_5288, n_5290;
wire n_5271, n_5272, n_5274, n_5275, n_5277, n_5278, n_5279, n_5280;
wire n_5261, n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5270;
wire n_5253, n_5254, n_5255, n_5256, n_5257, n_5258, n_5259, n_5260;
wire n_5237, n_5238, n_5239, n_5245, n_5246, n_5247, n_5250, n_5251;
wire n_5226, n_5227, n_5229, n_5230, n_5231, n_5232, n_5233, n_5234;
wire n_5210, n_5211, n_5212, n_5213, n_5214, n_5215, n_5220, n_5223;
wire n_5200, n_5201, n_5202, n_5205, n_5206, n_5207, n_5208, n_5209;
wire n_5189, n_5190, n_5191, n_5192, n_5193, n_5196, n_5198, n_5199;
wire n_5180, n_5181, n_5182, n_5183, n_5184, n_5186, n_5187, n_5188;
wire n_5168, n_5169, n_5171, n_5172, n_5175, n_5176, n_5178, n_5179;
wire n_5156, n_5157, n_5159, n_5162, n_5163, n_5165, n_5166, n_5167;
wire n_5143, n_5145, n_5146, n_5148, n_5149, n_5150, n_5154, n_5155;
wire n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5141;
wire n_5117, n_5118, n_5119, n_5120, n_5122, n_5124, n_5126, n_5129;
wire n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116;
wire n_5098, n_5099, n_5100, n_5101, n_5103, n_5104, n_5106, n_5108;
wire n_5081, n_5082, n_5083, n_5086, n_5087, n_5088, n_5089, n_5097;
wire n_5068, n_5069, n_5071, n_5072, n_5073, n_5076, n_5077, n_5078;
wire n_5044, n_5047, n_5049, n_5051, n_5053, n_5059, n_5064, n_5067;
wire n_5030, n_5031, n_5032, n_5033, n_5034, n_5035, n_5036, n_5037;
wire n_5022, n_5023, n_5024, n_5025, n_5026, n_5027, n_5028, n_5029;
wire n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019, n_5020;
wire n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011, n_5012;
wire n_4985, n_4997, n_4999, n_5000, n_5001, n_5002, n_5003, n_5004;
wire n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978, n_4979;
wire n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4970, n_4971;
wire n_4950, n_4951, n_4952, n_4953, n_4954, n_4955, n_4957, n_4958;
wire n_4939, n_4941, n_4944, n_4945, n_4946, n_4947, n_4948, n_4949;
wire n_4928, n_4929, n_4930, n_4932, n_4934, n_4936, n_4937, n_4938;
wire n_4919, n_4920, n_4921, n_4923, n_4924, n_4925, n_4926, n_4927;
wire n_4901, n_4902, n_4910, n_4912, n_4913, n_4915, n_4917, n_4918;
wire n_4885, n_4894, n_4895, n_4896, n_4897, n_4898, n_4899, n_4900;
wire n_4877, n_4878, n_4879, n_4880, n_4881, n_4882, n_4883, n_4884;
wire n_4869, n_4870, n_4871, n_4872, n_4873, n_4874, n_4875, n_4876;
wire n_4857, n_4859, n_4861, n_4862, n_4863, n_4865, n_4866, n_4867;
wire n_4847, n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4856;
wire n_4831, n_4836, n_4838, n_4840, n_4842, n_4843, n_4844, n_4846;
wire n_4816, n_4817, n_4818, n_4822, n_4825, n_4826, n_4827, n_4828;
wire n_4798, n_4800, n_4801, n_4804, n_4805, n_4809, n_4813, n_4815;
wire n_4787, n_4788, n_4789, n_4790, n_4791, n_4792, n_4796, n_4797;
wire n_4779, n_4780, n_4781, n_4782, n_4783, n_4784, n_4785, n_4786;
wire n_4767, n_4769, n_4770, n_4771, n_4772, n_4773, n_4777, n_4778;
wire n_4751, n_4752, n_4755, n_4756, n_4757, n_4760, n_4763, n_4765;
wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
wire n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742;
wire n_4726, n_4727, n_4728, n_4729, n_4731, n_4732, n_4733, n_4734;
wire n_4713, n_4714, n_4715, n_4716, n_4717, n_4718, n_4722, n_4725;
wire n_4704, n_4706, n_4707, n_4708, n_4709, n_4710, n_4711, n_4712;
wire n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701, n_4703;
wire n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693, n_4694;
wire n_4678, n_4679, n_4681, n_4682, n_4683, n_4684, n_4685, n_4686;
wire n_4669, n_4670, n_4671, n_4672, n_4674, n_4675, n_4676, n_4677;
wire n_4660, n_4661, n_4662, n_4663, n_4664, n_4665, n_4666, n_4667;
wire n_4652, n_4653, n_4654, n_4655, n_4656, n_4657, n_4658, n_4659;
wire n_4640, n_4641, n_4642, n_4644, n_4645, n_4648, n_4649, n_4650;
wire n_4626, n_4627, n_4630, n_4631, n_4635, n_4636, n_4637, n_4639;
wire n_4610, n_4612, n_4613, n_4614, n_4615, n_4618, n_4624, n_4625;
wire n_4597, n_4598, n_4599, n_4601, n_4602, n_4603, n_4604, n_4605;
wire n_4585, n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596;
wire n_4577, n_4578, n_4579, n_4580, n_4581, n_4582, n_4583, n_4584;
wire n_4567, n_4568, n_4569, n_4570, n_4572, n_4573, n_4574, n_4576;
wire n_4551, n_4553, n_4558, n_4559, n_4561, n_4562, n_4563, n_4564;
wire n_4540, n_4542, n_4543, n_4544, n_4545, n_4547, n_4548, n_4550;
wire n_4531, n_4532, n_4533, n_4534, n_4535, n_4537, n_4538, n_4539;
wire n_4522, n_4523, n_4524, n_4525, n_4527, n_4528, n_4529, n_4530;
wire n_4514, n_4515, n_4516, n_4517, n_4518, n_4519, n_4520, n_4521;
wire n_4505, n_4507, n_4508, n_4509, n_4510, n_4511, n_4512, n_4513;
wire n_4486, n_4497, n_4498, n_4500, n_4501, n_4502, n_4503, n_4504;
wire n_4475, n_4476, n_4477, n_4478, n_4479, n_4480, n_4483, n_4484;
wire n_4463, n_4464, n_4465, n_4466, n_4468, n_4469, n_4471, n_4474;
wire n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461, n_4462;
wire n_4441, n_4444, n_4446, n_4448, n_4449, n_4450, n_4451, n_4454;
wire n_4426, n_4428, n_4432, n_4433, n_4434, n_4435, n_4436, n_4439;
wire n_4412, n_4416, n_4418, n_4419, n_4420, n_4423, n_4424, n_4425;
wire n_4399, n_4400, n_4401, n_4402, n_4403, n_4409, n_4410, n_4411;
wire n_4389, n_4390, n_4392, n_4393, n_4394, n_4395, n_4397, n_4398;
wire n_4379, n_4380, n_4381, n_4382, n_4384, n_4385, n_4387, n_4388;
wire n_4367, n_4368, n_4369, n_4374, n_4375, n_4376, n_4377, n_4378;
wire n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365, n_4366;
wire n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357, n_4358;
wire n_4342, n_4343, n_4345, n_4346, n_4347, n_4348, n_4349, n_4350;
wire n_4332, n_4333, n_4334, n_4335, n_4337, n_4338, n_4339, n_4341;
wire n_4323, n_4324, n_4325, n_4326, n_4328, n_4329, n_4330, n_4331;
wire n_4312, n_4315, n_4317, n_4318, n_4319, n_4320, n_4321, n_4322;
wire n_4301, n_4302, n_4304, n_4305, n_4306, n_4308, n_4309, n_4311;
wire n_4290, n_4291, n_4292, n_4295, n_4296, n_4297, n_4298, n_4300;
wire n_4282, n_4283, n_4284, n_4285, n_4286, n_4287, n_4288, n_4289;
wire n_4273, n_4274, n_4275, n_4277, n_4278, n_4279, n_4280, n_4281;
wire n_4261, n_4262, n_4263, n_4264, n_4265, n_4266, n_4267, n_4270;
wire n_4242, n_4244, n_4245, n_4246, n_4253, n_4254, n_4256, n_4259;
wire n_4230, n_4231, n_4233, n_4234, n_4236, n_4237, n_4239, n_4240;
wire n_4219, n_4220, n_4221, n_4223, n_4226, n_4227, n_4228, n_4229;
wire n_4208, n_4209, n_4210, n_4211, n_4213, n_4214, n_4216, n_4218;
wire n_4194, n_4195, n_4201, n_4202, n_4203, n_4205, n_4206, n_4207;
wire n_4181, n_4182, n_4183, n_4185, n_4187, n_4188, n_4192, n_4193;
wire n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4178, n_4179;
wire n_4160, n_4161, n_4162, n_4163, n_4164, n_4168, n_4169, n_4170;
wire n_4145, n_4147, n_4149, n_4151, n_4152, n_4153, n_4155, n_4159;
wire n_4133, n_4135, n_4137, n_4138, n_4139, n_4140, n_4141, n_4143;
wire n_4113, n_4114, n_4115, n_4116, n_4117, n_4125, n_4127, n_4128;
wire n_4105, n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112;
wire n_4097, n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104;
wire n_4089, n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096;
wire n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088;
wire n_4072, n_4073, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080;
wire n_4063, n_4064, n_4065, n_4066, n_4067, n_4068, n_4069, n_4071;
wire n_4054, n_4055, n_4056, n_4058, n_4059, n_4060, n_4061, n_4062;
wire n_4046, n_4047, n_4048, n_4049, n_4050, n_4051, n_4052, n_4053;
wire n_4035, n_4037, n_4038, n_4039, n_4042, n_4043, n_4044, n_4045;
wire n_4021, n_4023, n_4025, n_4027, n_4028, n_4029, n_4031, n_4034;
wire n_4011, n_4014, n_4015, n_4016, n_4017, n_4018, n_4019, n_4020;
wire n_3996, n_3997, n_4000, n_4001, n_4003, n_4004, n_4009, n_4010;
wire n_3986, n_3987, n_3988, n_3989, n_3991, n_3992, n_3993, n_3994;
wire n_3975, n_3977, n_3978, n_3979, n_3980, n_3981, n_3984, n_3985;
wire n_3959, n_3960, n_3966, n_3968, n_3970, n_3971, n_3972, n_3974;
wire n_3948, n_3950, n_3951, n_3952, n_3953, n_3954, n_3955, n_3956;
wire n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3945;
wire n_3919, n_3928, n_3929, n_3930, n_3931, n_3933, n_3935, n_3936;
wire n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3914;
wire n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, n_3902;
wire n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, n_3893;
wire n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, n_3884;
wire n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876;
wire n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867;
wire n_3847, n_3848, n_3849, n_3853, n_3854, n_3855, n_3856, n_3859;
wire n_3836, n_3837, n_3840, n_3841, n_3842, n_3844, n_3845, n_3846;
wire n_3825, n_3827, n_3828, n_3829, n_3830, n_3833, n_3834, n_3835;
wire n_3814, n_3815, n_3816, n_3820, n_3821, n_3822, n_3823, n_3824;
wire n_3795, n_3799, n_3800, n_3804, n_3805, n_3808, n_3810, n_3812;
wire n_3772, n_3773, n_3774, n_3781, n_3790, n_3792, n_3793, n_3794;
wire n_3763, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, n_3771;
wire n_3753, n_3754, n_3755, n_3756, n_3759, n_3760, n_3761, n_3762;
wire n_3737, n_3738, n_3739, n_3741, n_3742, n_3743, n_3744, n_3752;
wire n_3726, n_3728, n_3729, n_3731, n_3732, n_3734, n_3735, n_3736;
wire n_3717, n_3718, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725;
wire n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716;
wire n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3707, n_3708;
wire n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698;
wire n_3682, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, n_3690;
wire n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681;
wire n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, n_3669, n_3671;
wire n_3651, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661;
wire n_3635, n_3636, n_3638, n_3642, n_3643, n_3646, n_3648, n_3650;
wire n_3620, n_3625, n_3628, n_3629, n_3630, n_3632, n_3633, n_3634;
wire n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616;
wire n_3597, n_3601, n_3602, n_3603, n_3605, n_3606, n_3607, n_3608;
wire n_3579, n_3580, n_3581, n_3588, n_3589, n_3592, n_3595, n_3596;
wire n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, n_3578;
wire n_3560, n_3561, n_3562, n_3563, n_3565, n_3567, n_3568, n_3569;
wire n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559;
wire n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, n_3551;
wire n_3534, n_3536, n_3537, n_3539, n_3540, n_3541, n_3542, n_3543;
wire n_3523, n_3524, n_3525, n_3527, n_3529, n_3530, n_3531, n_3533;
wire n_3509, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, n_3521;
wire n_3479, n_3480, n_3482, n_3485, n_3489, n_3498, n_3499, n_3508;
wire n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478;
wire n_3460, n_3461, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468;
wire n_3450, n_3451, n_3452, n_3454, n_3455, n_3457, n_3458, n_3459;
wire n_3440, n_3441, n_3442, n_3443, n_3445, n_3447, n_3448, n_3449;
wire n_3427, n_3428, n_3429, n_3430, n_3431, n_3433, n_3438, n_3439;
wire n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426;
wire n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418;
wire n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410;
wire n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402;
wire n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394;
wire n_3378, n_3379, n_3380, n_3381, n_3382, n_3384, n_3385, n_3386;
wire n_3363, n_3364, n_3367, n_3368, n_3370, n_3372, n_3374, n_3377;
wire n_3352, n_3353, n_3354, n_3355, n_3356, n_3357, n_3359, n_3361;
wire n_3343, n_3344, n_3345, n_3346, n_3347, n_3349, n_3350, n_3351;
wire n_3334, n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3342;
wire n_3319, n_3320, n_3322, n_3324, n_3325, n_3331, n_3332, n_3333;
wire n_3308, n_3310, n_3311, n_3312, n_3313, n_3314, n_3316, n_3317;
wire n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307;
wire n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3298, n_3299;
wire n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290;
wire n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282;
wire n_3256, n_3260, n_3263, n_3264, n_3269, n_3270, n_3271, n_3274;
wire n_3245, n_3247, n_3249, n_3251, n_3252, n_3253, n_3254, n_3255;
wire n_3229, n_3231, n_3232, n_3233, n_3235, n_3236, n_3237, n_3239;
wire n_3217, n_3218, n_3220, n_3221, n_3222, n_3224, n_3225, n_3227;
wire n_3203, n_3204, n_3205, n_3206, n_3207, n_3212, n_3213, n_3216;
wire n_3188, n_3190, n_3194, n_3195, n_3199, n_3200, n_3201, n_3202;
wire n_3172, n_3173, n_3174, n_3175, n_3176, n_3178, n_3180, n_3187;
wire n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171;
wire n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163;
wire n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3155;
wire n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146;
wire n_3129, n_3130, n_3131, n_3133, n_3134, n_3136, n_3137, n_3138;
wire n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, n_3128;
wire n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120;
wire n_3103, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112;
wire n_3081, n_3082, n_3083, n_3085, n_3089, n_3093, n_3094, n_3096;
wire n_3070, n_3072, n_3073, n_3074, n_3075, n_3078, n_3079, n_3080;
wire n_3059, n_3061, n_3063, n_3064, n_3065, n_3066, n_3068, n_3069;
wire n_3047, n_3051, n_3052, n_3053, n_3055, n_3056, n_3057, n_3058;
wire n_3038, n_3039, n_3040, n_3041, n_3042, n_3044, n_3045, n_3046;
wire n_3027, n_3029, n_3031, n_3032, n_3034, n_3035, n_3036, n_3037;
wire n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3022, n_3023;
wire n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005;
wire n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2996;
wire n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987;
wire n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, n_2979;
wire n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2967, n_2969;
wire n_2949, n_2951, n_2952, n_2953, n_2954, n_2956, n_2957, n_2958;
wire n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, n_2948;
wire n_2920, n_2921, n_2922, n_2925, n_2927, n_2929, n_2938, n_2940;
wire n_2907, n_2908, n_2909, n_2910, n_2913, n_2915, n_2916, n_2917;
wire n_2896, n_2898, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905;
wire n_2887, n_2888, n_2889, n_2890, n_2892, n_2893, n_2894, n_2895;
wire n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886;
wire n_2870, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878;
wire n_2857, n_2859, n_2861, n_2862, n_2863, n_2865, n_2867, n_2868;
wire n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854;
wire n_2839, n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846;
wire n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838;
wire n_2821, n_2822, n_2823, n_2824, n_2826, n_2828, n_2829, n_2830;
wire n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820;
wire n_2799, n_2803, n_2805, n_2808, n_2809, n_2810, n_2811, n_2812;
wire n_2784, n_2785, n_2786, n_2788, n_2790, n_2794, n_2795, n_2797;
wire n_2770, n_2772, n_2773, n_2774, n_2776, n_2779, n_2780, n_2783;
wire n_2761, n_2762, n_2763, n_2764, n_2765, n_2767, n_2768, n_2769;
wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
wire n_2736, n_2737, n_2738, n_2739, n_2741, n_2742, n_2743, n_2744;
wire n_2719, n_2720, n_2722, n_2723, n_2724, n_2732, n_2733, n_2735;
wire n_2710, n_2711, n_2712, n_2714, n_2715, n_2716, n_2717, n_2718;
wire n_2693, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2709;
wire n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, n_2691, n_2692;
wire n_2677, n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684;
wire n_2665, n_2667, n_2668, n_2670, n_2672, n_2674, n_2675, n_2676;
wire n_2656, n_2657, n_2658, n_2659, n_2660, n_2662, n_2663, n_2664;
wire n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655;
wire n_2636, n_2637, n_2638, n_2639, n_2641, n_2645, n_2646, n_2647;
wire n_2626, n_2627, n_2629, n_2631, n_2632, n_2633, n_2634, n_2635;
wire n_2615, n_2617, n_2618, n_2619, n_2621, n_2623, n_2624, n_2625;
wire n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614;
wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606;
wire n_2588, n_2589, n_2591, n_2593, n_2594, n_2595, n_2597, n_2598;
wire n_2579, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587;
wire n_2566, n_2568, n_2569, n_2570, n_2571, n_2572, n_2576, n_2578;
wire n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2561, n_2563;
wire n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545;
wire n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537;
wire n_2518, n_2520, n_2524, n_2525, n_2526, n_2527, n_2528, n_2529;
wire n_2506, n_2507, n_2508, n_2509, n_2511, n_2512, n_2516, n_2517;
wire n_2496, n_2497, n_2499, n_2501, n_2502, n_2503, n_2504, n_2505;
wire n_2486, n_2488, n_2489, n_2490, n_2492, n_2493, n_2494, n_2495;
wire n_2477, n_2478, n_2479, n_2480, n_2482, n_2483, n_2484, n_2485;
wire n_2468, n_2469, n_2470, n_2472, n_2473, n_2474, n_2475, n_2476;
wire n_2451, n_2454, n_2456, n_2457, n_2458, n_2463, n_2465, n_2466;
wire n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2449, n_2450;
wire n_2416, n_2418, n_2419, n_2422, n_2433, n_2436, n_2437, n_2439;
wire n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2413;
wire n_2391, n_2393, n_2395, n_2396, n_2397, n_2398, n_2399, n_2403;
wire n_2381, n_2382, n_2383, n_2384, n_2386, n_2388, n_2389, n_2390;
wire n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379;
wire n_2360, n_2361, n_2362, n_2363, n_2365, n_2368, n_2369, n_2370;
wire n_2343, n_2346, n_2353, n_2354, n_2355, n_2356, n_2357, n_2358;
wire n_2322, n_2326, n_2334, n_2336, n_2337, n_2338, n_2339, n_2340;
wire n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2318, n_2320;
wire n_2302, n_2303, n_2304, n_2306, n_2307, n_2308, n_2309, n_2310;
wire n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301;
wire n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293;
wire n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284;
wire n_2267, n_2268, n_2269, n_2270, n_2272, n_2273, n_2275, n_2276;
wire n_2254, n_2256, n_2257, n_2258, n_2259, n_2261, n_2264, n_2266;
wire n_2242, n_2243, n_2245, n_2246, n_2250, n_2251, n_2252, n_2253;
wire n_2221, n_2228, n_2231, n_2232, n_2233, n_2235, n_2237, n_2238;
wire n_2208, n_2210, n_2211, n_2212, n_2215, n_2217, n_2218, n_2220;
wire n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207;
wire n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199;
wire n_2182, n_2183, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191;
wire n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181;
wire n_2164, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172;
wire n_2155, n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2163;
wire n_2143, n_2145, n_2147, n_2148, n_2149, n_2151, n_2153, n_2154;
wire n_2134, n_2135, n_2136, n_2137, n_2138, n_2140, n_2141, n_2142;
wire n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, n_2133;
wire n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125;
wire n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116;
wire n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108;
wire n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100;
wire n_2083, n_2084, n_2086, n_2087, n_2089, n_2090, n_2091, n_2092;
wire n_2072, n_2073, n_2074, n_2075, n_2076, n_2078, n_2080, n_2081;
wire n_2063, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071;
wire n_2048, n_2051, n_2052, n_2053, n_2055, n_2056, n_2058, n_2061;
wire n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2046;
wire n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037;
wire n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025;
wire n_2009, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017;
wire n_2000, n_2001, n_2003, n_2004, n_2005, n_2006, n_2007, n_2008;
wire n_1985, n_1986, n_1989, n_1990, n_1992, n_1997, n_1998, n_1999;
wire n_1976, n_1977, n_1978, n_1979, n_1980, n_1982, n_1983, n_1984;
wire n_1967, n_1968, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975;
wire n_1956, n_1957, n_1959, n_1960, n_1962, n_1963, n_1964, n_1966;
wire n_1944, n_1945, n_1946, n_1949, n_1951, n_1952, n_1954, n_1955;
wire n_1932, n_1933, n_1934, n_1935, n_1936, n_1938, n_1942, n_1943;
wire n_1919, n_1920, n_1921, n_1922, n_1924, n_1926, n_1929, n_1930;
wire n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918;
wire n_1901, n_1902, n_1904, n_1906, n_1907, n_1908, n_1909, n_1910;
wire n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, n_1899, n_1900;
wire n_1879, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888;
wire n_1864, n_1866, n_1868, n_1873, n_1874, n_1875, n_1876, n_1878;
wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1856, n_1861;
wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
wire n_1808, n_1809, n_1810, n_1812, n_1813, n_1814, n_1815, n_1816;
wire n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807;
wire n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799;
wire n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791;
wire n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783;
wire n_1767, n_1768, n_1769, n_1770, n_1772, n_1773, n_1774, n_1775;
wire n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766;
wire n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1758;
wire n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749;
wire n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741;
wire n_1724, n_1725, n_1727, n_1728, n_1730, n_1731, n_1732, n_1733;
wire n_1715, n_1716, n_1717, n_1718, n_1719, n_1721, n_1722, n_1723;
wire n_1703, n_1705, n_1707, n_1708, n_1710, n_1711, n_1712, n_1714;
wire n_1689, n_1691, n_1693, n_1696, n_1697, n_1700, n_1701, n_1702;
wire n_1673, n_1675, n_1676, n_1677, n_1678, n_1679, n_1681, n_1682;
wire n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672;
wire n_1653, n_1655, n_1656, n_1657, n_1658, n_1660, n_1662, n_1663;
wire n_1638, n_1639, n_1641, n_1642, n_1649, n_1650, n_1651, n_1652;
wire n_1627, n_1628, n_1629, n_1631, n_1632, n_1634, n_1635, n_1636;
wire n_1615, n_1616, n_1618, n_1619, n_1621, n_1622, n_1624, n_1626;
wire n_1605, n_1606, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613;
wire n_1594, n_1596, n_1597, n_1598, n_1600, n_1601, n_1603, n_1604;
wire n_1575, n_1576, n_1577, n_1580, n_1581, n_1586, n_1587, n_1593;
wire n_1566, n_1567, n_1568, n_1569, n_1571, n_1572, n_1573, n_1574;
wire n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565;
wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
wire n_1533, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
wire n_1525, n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532;
wire n_1514, n_1515, n_1516, n_1517, n_1518, n_1521, n_1523, n_1524;
wire n_1504, n_1505, n_1506, n_1507, n_1508, n_1510, n_1511, n_1513;
wire n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503;
wire n_1465, n_1466, n_1467, n_1469, n_1470, n_1483, n_1492, n_1494;
wire n_1456, n_1457, n_1458, n_1459, n_1461, n_1462, n_1463, n_1464;
wire n_1446, n_1447, n_1448, n_1449, n_1452, n_1453, n_1454, n_1455;
wire n_1436, n_1437, n_1438, n_1439, n_1441, n_1442, n_1443, n_1445;
wire n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1435;
wire n_1416, n_1418, n_1420, n_1421, n_1422, n_1424, n_1425, n_1426;
wire n_1391, n_1392, n_1396, n_1399, n_1401, n_1402, n_1403, n_1410;
wire n_1381, n_1382, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389;
wire n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380;
wire n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372;
wire n_1352, n_1353, n_1354, n_1355, n_1357, n_1359, n_1363, n_1364;
wire n_1340, n_1342, n_1343, n_1344, n_1346, n_1347, n_1348, n_1349;
wire n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339;
wire n_1323, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331;
wire n_1305, n_1312, n_1313, n_1314, n_1315, n_1320, n_1321, n_1322;
wire n_1290, n_1292, n_1295, n_1299, n_1300, n_1301, n_1302, n_1304;
wire n_1275, n_1277, n_1278, n_1279, n_1280, n_1285, n_1287, n_1288;
wire n_1265, n_1266, n_1268, n_1269, n_1270, n_1271, n_1273, n_1274;
wire n_1256, n_1257, n_1258, n_1259, n_1260, n_1262, n_1263, n_1264;
wire n_1245, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253;
wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1240, n_1241, n_1244;
wire n_1213, n_1214, n_1217, n_1218, n_1219, n_1220, n_1223, n_1225;
wire n_1204, n_1205, n_1206, n_1208, n_1209, n_1210, n_1211, n_1212;
wire n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203;
wire n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195;
wire n_1179, n_1180, n_1181, n_1182, n_1184, n_1185, n_1186, n_1187;
wire n_1170, n_1171, n_1172, n_1173, n_1174, n_1176, n_1177, n_1178;
wire n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169;
wire n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161;
wire n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1150, n_1152;
wire n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1140;
wire n_1121, n_1122, n_1123, n_1125, n_1126, n_1127, n_1129, n_1131;
wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1120;
wire n_1100, n_1101, n_1102, n_1104, n_1105, n_1107, n_1108, n_1109;
wire n_1088, n_1089, n_1090, n_1092, n_1093, n_1094, n_1095, n_1099;
wire n_1077, n_1079, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087;
wire n_1067, n_1068, n_1069, n_1070, n_1073, n_1074, n_1075, n_1076;
wire n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066;
wire n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058;
wire n_1040, n_1041, n_1043, n_1044, n_1046, n_1047, n_1048, n_1049;
wire n_1028, n_1030, n_1031, n_1032, n_1033, n_1034, n_1036, n_1039;
wire n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026;
wire n_1006, n_1007, n_1008, n_1013, n_1014, n_1015, n_1016, n_1017;
wire n_985, n_986, n_987, n_998, n_999, n_1001, n_1003, n_1004;
wire n_976, n_977, n_978, n_980, n_981, n_982, n_983, n_984;
wire n_966, n_967, n_969, n_970, n_971, n_972, n_973, n_975;
wire n_952, n_953, n_955, n_956, n_960, n_963, n_964, n_965;
wire n_941, n_942, n_943, n_944, n_946, n_949, n_950, n_951;
wire n_933, n_934, n_935, n_936, n_937, n_938, n_939, n_940;
wire n_913, n_917, n_918, n_920, n_922, n_923, n_930, n_931;
wire n_903, n_904, n_905, n_908, n_909, n_910, n_911, n_912;
wire n_892, n_893, n_894, n_896, n_899, n_900, n_901, n_902;
wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
wire n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883;
wire n_867, n_868, n_870, n_871, n_872, n_873, n_874, n_875;
wire n_854, n_856, n_857, n_862, n_863, n_864, n_865, n_866;
wire n_843, n_844, n_845, n_846, n_848, n_850, n_852, n_853;
wire n_834, n_835, n_836, n_837, n_839, n_840, n_841, n_842;
wire n_818, n_819, n_820, n_821, n_830, n_831, n_832, n_833;
wire n_806, n_807, n_809, n_810, n_811, n_812, n_814, n_816;
wire n_797, n_798, n_799, n_800, n_801, n_802, n_803, n_805;
wire n_787, n_788, n_789, n_790, n_792, n_793, n_794, n_796;
wire n_776, n_777, n_779, n_781, n_782, n_783, n_785, n_786;
wire n_767, n_769, n_770, n_771, n_772, n_773, n_774, n_775;
wire n_756, n_757, n_758, n_759, n_761, n_762, n_763, n_766;
wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
wire n_734, n_735, n_737, n_739, n_742, n_744, n_745, n_747;
wire n_723, n_726, n_727, n_729, n_730, n_731, n_732, n_733;
wire n_711, n_712, n_713, n_714, n_715, n_718, n_719, n_721;
wire n_701, n_703, n_704, n_705, n_706, n_707, n_709, n_710;
wire n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700;
wire n_682, n_686, n_687, n_688, n_689, n_690, n_691, n_692;
wire n_670, n_671, n_672, n_676, n_677, n_678, n_679, n_680;
wire n_660, n_661, n_662, n_664, n_665, n_666, n_667, n_669;
wire n_650, n_651, n_652, n_654, n_655, n_656, n_657, n_659;
wire n_640, n_642, n_643, n_645, n_646, n_647, n_648, n_649;
wire n_630, n_631, n_632, n_633, n_634, n_636, n_638, n_639;
wire n_608, n_609, n_613, n_614, n_616, n_617, n_619, n_624;
wire n_595, n_597, n_599, n_600, n_601, n_602, n_603, n_605;
wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
wire n_576, n_578, n_579, n_580, n_581, n_583, n_584, n_585;
wire n_562, n_563, n_564, n_565, n_568, n_569, n_570, n_571;
wire n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561;
wire n_546, n_547, n_548, n_549, n_550, n_551, n_552, n_553;
wire n_535, n_536, n_537, n_538, n_539, n_540, n_542, n_545;
wire n_518, n_519, n_521, n_522, n_525, n_527, n_528, n_529;
wire n_487, n_494, n_495, n_496, n_501, n_504, n_505, n_517;
wire n_476, n_477, n_478, n_479, n_482, n_483, n_484, n_485;
wire n_466, n_467, n_468, n_470, n_471, n_473, n_474, n_475;
wire n_454, n_455, n_456, n_458, n_459, n_460, n_461, n_465;
wire n_425, n_431, n_433, n_435, n_436, n_442, n_447, n_448;
wire n_413, n_415, n_416, n_417, n_418, n_419, n_420, n_422;
wire n_384, n_385, n_386, n_389, n_404, n_410, n_411, n_412;
wire n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379;
wire n_363, n_364, n_365, n_366, n_367, n_368, n_369, n_370;
wire n_351, n_352, n_355, n_356, n_357, n_358, n_359, n_360;
wire n_338, n_339, n_342, n_343, n_344, n_348, n_349, n_350;
wire n_324, n_326, n_328, n_330, n_332, n_334, n_336, n_337;
wire n_308, n_310, n_313, n_315, n_317, n_319, n_321, n_322;
wire n_294, n_296, n_297, n_298, n_300, n_301, n_303, n_306;
wire n_276, n_278, n_282, n_283, n_286, n_288, n_289, n_293;
wire n_255, n_260, n_264, n_266, n_268, n_269, n_271, n_275;
wire n_237, n_239, n_241, n_245, n_247, n_249, n_251, n_254;
wire n_222, n_225, n_226, n_228, n_231, n_233, n_234, n_236;
wire n_206, n_207, n_209, n_211, n_213, n_215, n_216, n_220;
wire n_185, n_187, n_189, n_193, n_198, n_200, n_202, n_204;
wire n_167, n_170, n_172, n_174, n_176, n_180, n_182, n_183;
wire n_147, n_149, n_151, n_153, n_155, n_157, n_163, n_166;
wire n_126, n_129, n_131, n_132, n_137, n_139, n_141, n_143;
wire n_116, n_117, n_118, n_120, n_121, n_122, n_123, n_125;
wire n_104, n_105, n_106, n_107, n_108, n_111, n_112, n_113;
wire n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_103;
wire n_84, n_86, n_87, n_88, n_89, n_91, n_93, n_94;
wire n_75, n_76, n_77, n_78, n_79, n_80, n_81, n_83;
wire n_63, n_64, n_66, n_67, n_68, n_69, n_70, n_72;
wire n_54, n_55, n_56, n_58, n_59, n_60, n_61, n_62;
wire n_43, n_44, n_45, n_47, n_48, n_51, n_52, n_53;
wire n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_42;
wire n_24, n_25, n_26, n_27, n_28, n_30, n_31, n_32;
wire n_11, n_12, n_14, n_17, n_18, n_21, n_22, n_23;
wire n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10;
wire gbuf207, gbuf210, gbuf211, gbuf212, gbuf213, gbuf214, n_0, n_2;
wire gbuf195, gbuf200, gbuf201, gbuf202, gbuf203, gbuf204, gbuf205, gbuf206;
wire gbuf187, gbuf188, gbuf189, gbuf190, gbuf191, gbuf192, gbuf193, gbuf194;
wire gbuf179, gbuf180, gbuf181, gbuf182, gbuf183, gbuf184, gbuf185, gbuf186;
wire gbuf163, gbuf164, gbuf165, gbuf171, gbuf175, gbuf176, gbuf177, gbuf178;
wire gbuf153, gbuf154, gbuf155, gbuf156, gbuf157, gbuf158, gbuf161, gbuf162;
wire gbuf141, gbuf142, gbuf143, gbuf144, gbuf145, gbuf146, gbuf151, gbuf152;
wire gbuf133, gbuf134, gbuf135, gbuf136, gbuf137, gbuf138, gbuf139, gbuf140;
wire gbuf122, gbuf126, gbuf127, gbuf128, gbuf129, gbuf130, gbuf131, gbuf132;
wire gbuf107, gbuf108, gbuf109, gbuf112, gbuf113, gbuf114, gbuf115, gbuf116;
wire gbuf95, gbuf96, gbuf97, gbuf102, gbuf103, gbuf104, gbuf105, gbuf106;
wire gbuf87, gbuf88, gbuf89, gbuf90, gbuf91, gbuf92, gbuf93, gbuf94;
wire gbuf79, gbuf80, gbuf81, gbuf82, gbuf83, gbuf84, gbuf85, gbuf86;
wire gbuf63, gbuf64, gbuf65, gbuf66, gbuf67, gbuf73, gbuf77, gbuf78;
wire gbuf53, gbuf54, gbuf55, gbuf56, gbuf57, gbuf58, gbuf59, gbuf60;
wire gbuf41, gbuf42, gbuf43, gbuf44, gbuf45, gbuf46, gbuf47, gbuf48;
wire gbuf33, gbuf34, gbuf35, gbuf36, gbuf37, gbuf38, gbuf39, gbuf40;
wire g_32037, g_32166, gbuf24, gbuf28, gbuf29, gbuf30, gbuf31, gbuf32;
wire g_29316, g_29721, g_30039, g_30213, g_30245, g_30261, g_30665, g_31512;
wire g_28035, g_28142, g_28592, g_28702, g_29016, g_29095, g_29207, g_29227;
wire g_27149, g_27699, g_27738, g_27846, g_27919, g_27924, g_27975, g_28034;
wire g_25958, g_25960, g_26059, g_26067, g_26130, g_26381, g_26529, g_26724;
wire g_25348, g_25350, g_25466, g_25523, g_25781, g_25878, g_25914, g_25929;
wire g_24459, g_24593, g_24632, g_24786, g_24794, g_24889, g_24922, g_25247;
wire g_22696, g_22901, g_23490, g_23514, g_23734, g_23988, g_24187, g_24437;
wire g_21690, g_21829, g_21927, g_22281, g_22340, g_22408, g_22536, g_22538;
wire g_20137, g_20180, g_20789, g_20947, g_20948, g_21144, g_21387, g_21556;
wire g_19223, g_19472, g_19787, g_19959, g_19985, g_19993, g_20059, g_20070;
wire g_18628, g_18792, g_18819, g_19017, g_19064, g_19110, g_19132, g_19162;
wire g_17921, g_18003, g_18059, g_18093, g_18173, g_18364, g_18412, g_18564;
wire g_16936, g_17001, g_17130, g_17170, g_17474, g_17483, g_17832, g_17877;
wire g_15095, g_15404, g_15687, g_15833, g_16164, g_16317, g_16484, g_16638;
wire g_14013, g_14626, g_14632, g_14662, g_14677, g_14726, g_14751, g_14855;
wire g_11807, g_12505, g_12670, g_12763, g_13227, g_13515, g_13546, g_13736;
wire g_9649, g_9980, g_10301, g_10341, g_10841, g_10959, g_11049, g_11640;
wire g_8090, g_8187, g_8360, g_8670, g_9014, g_9172, g_9470, g_9473;
wire g_5550, g_5793, g_5844, g_7108, g_7184, g_7905, g_8008, g_8082;
wire g3201, g3207, g3210, g3211, g_4886, g_5095, g_5159, g_5496;
wire g3176, g3179, g3182, g3185, g3191, g3194, g3197, g3198;
wire g3151, g3155, g3158, g3161, g3164, g3167, g3170, g3173;
wire g3132, g3133, g3134, g3135, g3136, g3139, g3142, g3147;
wire g3114, g3120, g3123, g3124, g3125, g3126, g3127, g3128;
wire g3106, g3107, g3108, g3109, g3110, g3111, g3112, g3113;
wire g3098, g3099, g3100, g3101, g3102, g3103, g3104, g3105;
wire g3088, g3091, g3092, g3093, g3094, g3095, g3096, g3097;
wire g3078, g3079, g3080, g3083, g3084, g3085, g3086, g3087;
wire g3070, g3071, g3072, g3073, g3074, g3075, g3076, g3077;
wire g3062, g3063, g3064, g3065, g3066, g3067, g3068, g3069;
wire g3054, g3055, g3056, g3057, g3058, g3059, g3060, g3061;
wire g3046, g3047, g3048, g3049, g3050, g3051, g3052, g3053;
wire g3018, g3024, g3028, g3032, g3036, g3043, g3044, g3045;
wire g2991, g2992, g2997, g2998, g3002, g3006, g3010, g3013;
wire g2975, g2978, g2981, g2984, g2985, g2986, g2987, g2990;
wire g2953, g2956, g2959, g2962, g2963, g2966, g2969, g2972;
wire g2929, g2933, g2934, g2935, g2938, g2941, g2944, g2947;
wire g2888, g2896, g2900, g2908, g2912, g2917, g2920, g2924;
wire g2817, g2857, g2873, g2874, g2877, g2878, g2879, g2883;
wire g2807, g2808, g2809, g2810, g2811, g2812, g2813, g2814;
wire g2799, g2800, g2801, g2802, g2803, g2804, g2805, g2806;
wire g2791, g2792, g2793, g2794, g2795, g2796, g2797, g2798;
wire g2783, g2784, g2785, g2786, g2787, g2788, g2789, g2790;
wire g2775, g2776, g2777, g2778, g2779, g2780, g2781, g2782;
wire g2734, g2740, g2746, g2760, g2766, g2772, g2773, g2774;
wire g2691, g2694, g2704, g2707, g2714, g2720, g2727, g2733;
wire g2667, g2670, g2673, g2676, g2679, g2682, g2685, g2688;
wire g2655, g2656, g2657, g2658, g2659, g2660, g2661, g2664;
wire g2645, g2647, g2649, g2650, g2651, g2652, g2653, g2654;
wire g2616, g2618, g2622, g2628, g2633, g2639, g2641, g2643;
wire g2605, g2606, g2607, g2608, g2610, g2611, g2612, g2615;
wire g2574, g2580, g2581, g2584, g2598, g2599, g2603, g2604;
wire g2560, g2561, g2562, g2563, g2564, g2565, g2568, g2571;
wire g2540, g2543, g2546, g2552, g2553, g2554, g2555, g2559;
wire g2523, g2524, g2526, g2528, g2530, g2533, g2536, g2539;
wire g2503, g2504, g2507, g2510, g2513, g2516, g2519, g2522;
wire g2483, g2486, g2489, g2492, g2495, g2498, g2501, g2502;
wire g2466, g2469, g2471, g2473, g2476, g2477, g2478, g2479;
wire g2444, g2448, g2451, g2454, g2456, g2458, g2459, g2463;
wire g2426, g2428, g2429, g2433, g2436, g2439, g2441, g2443;
wire g2396, g2397, g2398, g2399, g2412, g2418, g2421, g2424;
wire g2388, g2389, g2390, g2391, g2392, g2393, g2394, g2395;
wire g2362, g2364, g2366, g2373, g2374, g2380, g2384, g2387;
wire g2339, g2342, g2345, g2348, g2354, g2356, g2358, g2360;
wire g2315, g2318, g2321, g2324, g2327, g2330, g2333, g2336;
wire g2291, g2294, g2297, g2300, g2303, g2306, g2309, g2312;
wire g2267, g2270, g2273, g2276, g2279, g2282, g2285, g2288;
wire g2251, g2252, g2253, g2254, g2255, g2257, g2261, g2264;
wire g2241, g2244, g2245, g2246, g2247, g2248, g2249, g2250;
wire g2233, g2234, g2235, g2236, g2237, g2238, g2239, g2240;
wire g2225, g2226, g2227, g2228, g2229, g2230, g2231, g2232;
wire g2217, g2218, g2219, g2220, g2221, g2222, g2223, g2224;
wire g2190, g2195, g2205, g2206, g2207, g2208, g2209, g2210;
wire g2151, g2156, g2160, g2165, g2170, g2175, g2180, g2185;
wire g2119, g2120, g2124, g2129, g2133, g2138, g2142, g2147;
wire g2111, g2112, g2113, g2114, g2115, g2116, g2117, g2118;
wire g2103, g2104, g2105, g2106, g2107, g2108, g2109, g2110;
wire g2095, g2096, g2097, g2098, g2099, g2100, g2101, g2102;
wire g2087, g2088, g2089, g2090, g2091, g2092, g2093, g2094;
wire g2079, g2080, g2081, g2082, g2083, g2084, g2085, g2086;
wire g2033, g2039, g2040, g2046, g2052, g2066, g2072, g2078;
wire g1994, g1997, g2000, g2009, g2010, g2013, g2020, g2026;
wire g1970, g1973, g1976, g1979, g1982, g1985, g1988, g1991;
wire g1960, g1961, g1962, g1963, g1964, g1965, g1966, g1967;
wire g1949, g1951, g1953, g1955, g1956, g1957, g1958, g1959;
wire g1924, g1928, g1930, g1934, g1937, g1939, g1945, g1947;
wire g1912, g1913, g1914, g1916, g1917, g1918, g1921, g1922;
wire g1880, g1886, g1887, g1904, g1905, g1909, g1910, g1911;
wire g1866, g1867, g1868, g1869, g1870, g1871, g1874, g1877;
wire g1846, g1849, g1852, g1858, g1859, g1860, g1861, g1865;
wire g1829, g1830, g1832, g1834, g1836, g1839, g1842, g1845;
wire g1809, g1810, g1813, g1816, g1819, g1822, g1825, g1828;
wire g1789, g1792, g1795, g1798, g1801, g1804, g1807, g1808;
wire g1772, g1775, g1777, g1779, g1782, g1783, g1784, g1785;
wire g1750, g1754, g1757, g1760, g1762, g1764, g1765, g1769;
wire g1732, g1734, g1735, g1739, g1742, g1745, g1747, g1749;
wire g1702, g1703, g1704, g1705, g1718, g1724, g1727, g1730;
wire g1694, g1695, g1696, g1697, g1698, g1699, g1700, g1701;
wire g1666, g1668, g1670, g1672, g1679, g1680, g1686, g1693;
wire g1642, g1645, g1648, g1651, g1654, g1660, g1662, g1664;
wire g1618, g1621, g1624, g1627, g1630, g1633, g1636, g1639;
wire g1594, g1597, g1600, g1603, g1606, g1609, g1612, g1615;
wire g1570, g1573, g1576, g1579, g1582, g1585, g1588, g1591;
wire g1555, g1556, g1557, g1558, g1559, g1560, g1561, g1567;
wire g1545, g1546, g1547, g1550, g1551, g1552, g1553, g1554;
wire g1537, g1538, g1539, g1540, g1541, g1542, g1543, g1544;
wire g1529, g1530, g1531, g1532, g1533, g1534, g1535, g1536;
wire g1515, g1516, g1523, g1524, g1525, g1526, g1527, g1528;
wire g1476, g1481, g1486, g1501, g1511, g1512, g1513, g1514;
wire g1439, g1444, g1448, g1453, g1457, g1462, g1466, g1471;
wire g1420, g1421, g1422, g1423, g1424, g1425, g1430, g1435;
wire g1412, g1413, g1414, g1415, g1416, g1417, g1418, g1419;
wire g1404, g1405, g1406, g1407, g1408, g1409, g1410, g1411;
wire g1396, g1397, g1398, g1399, g1400, g1401, g1402, g1403;
wire g1388, g1389, g1390, g1391, g1392, g1393, g1394, g1395;
wire g1352, g1358, g1372, g1378, g1384, g1385, g1386, g1387;
wire g1315, g1316, g1319, g1326, g1332, g1339, g1345, g1346;
wire g1285, g1288, g1291, g1294, g1297, g1300, g1303, g1306;
wire g1269, g1270, g1271, g1272, g1273, g1276, g1279, g1282;
wire g1261, g1262, g1263, g1264, g1265, g1266, g1267, g1268;
wire g1240, g1243, g1245, g1251, g1253, g1255, g1257, g1259;
wire g1220, g1222, g1223, g1224, g1227, g1228, g1230, g1234;
wire g1193, g1210, g1211, g1215, g1216, g1217, g1218, g1219;
wire g1173, g1174, g1175, g1176, g1177, g1180, g1183, g1192;
wire g1155, g1158, g1164, g1165, g1166, g1167, g1171, g1172;
wire g1136, g1138, g1140, g1142, g1145, g1148, g1151, g1152;
wire g1116, g1119, g1122, g1125, g1128, g1131, g1134, g1135;
wire g1098, g1101, g1104, g1107, g1110, g1113, g1114, g1115;
wire g1081, g1083, g1085, g1088, g1089, g1090, g1091, g1095;
wire g1060, g1063, g1066, g1068, g1070, g1071, g1075, g1078;
wire g1040, g1041, g1045, g1048, g1051, g1053, g1055, g1056;
wire g1009, g1010, g1011, g1024, g1030, g1033, g1036, g1038;
wire g1001, g1002, g1003, g1004, g1005, g1006, g1007, g1008;
wire g976, g978, g985, g986, g992, g996, g999, g1000;
wire g954, g957, g960, g966, g968, g970, g972, g974;
wire g930, g933, g936, g939, g942, g945, g948, g951;
wire g906, g909, g912, g915, g918, g921, g924, g927;
wire g882, g885, g888, g891, g894, g897, g900, g903;
wire g864, g865, g866, g867, g869, g873, g876, g879;
wire g856, g857, g858, g859, g860, g861, g862, g863;
wire g845, g846, g847, g848, g849, g850, g851, g852;
wire g837, g838, g839, g840, g841, g842, g843, g844;
wire g829, g830, g831, g832, g833, g834, g835, g836;
wire g809, g813, g817, g818, g819, g820, g821, g822;
wire g776, g780, g785, g789, g793, g797, g801, g805;
wire g733, g734, g735, g736, g737, g738, g739, g771;
wire g725, g726, g727, g728, g729, g730, g731, g732;
wire g717, g718, g719, g720, g721, g722, g723, g724;
wire g709, g710, g711, g712, g713, g714, g715, g716;
wire g701, g702, g703, g704, g705, g706, g707, g708;
wire g660, g666, g672, g686, g692, g698, g699, g700;
wire g620, g629, g630, g633, g640, g646, g653, g659;
wire g596, g599, g602, g605, g608, g611, g614, g617;
wire g582, g583, g584, g585, g586, g587, g590, g593;
wire g573, g575, g576, g577, g578, g579, g580, g581;
wire g550, g554, g557, g559, g565, g567, g569, g571;
wire g487, g488, g489, g499, g524, g542, g544, g548;
wire g471, g477, g478, g479, g480, g484, g485, g486;
wire g451, g453, g455, g458, g461, g464, g465, g468;
wire g432, g435, g438, g441, g444, g447, g448, g449;
wire g414, g417, g420, g423, g426, g427, g428, g429;
wire g396, g398, g401, g402, g403, g404, g408, g411;
wire g361, g369, g373, g376, g384, g388, g391, g394;
wire g309, g312, g313, g322, g343, g346, g354, g358;
wire g252, g255, g258, g261, g264, g267, g270, g273;
wire g185, g231, g234, g237, g240, g243, g246, g249;
wire g97, g101, g105, g109, g113, g117, g121, g125;
wire g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380;
wire blif_clk_net, blif_reset_net, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234;
CLKBUFX1 gbuf_d_1(.A(n_8180), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(g185));
CLKBUFX1 gbuf_d_2(.A(n_8180), .Y(d_out_2));
CLKBUFX1 gbuf_q_2(.A(q_in_2), .Y(g3133));
CLKBUFX1 gbuf_d_3(.A(n_8178), .Y(d_out_3));
CLKBUFX1 gbuf_qn_3(.A(qn_in_3), .Y(g3128));
CLKBUFX1 gbuf_d_4(.A(g27380), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(g3139));
CLKBUFX1 gbuf_d_5(.A(g27380), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(g3151));
CLKBUFX1 gbuf_d_6(.A(g27380), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(n_411));
CLKBUFX1 gbuf_d_7(.A(g26135), .Y(d_out_7));
CLKBUFX1 gbuf_qn_7(.A(qn_in_7), .Y(g3134));
CLKBUFX1 gbuf_d_8(.A(g26135), .Y(d_out_8));
CLKBUFX1 gbuf_q_8(.A(q_in_8), .Y(g3147));
CLKBUFX1 gbuf_d_9(.A(g26135), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(g3114));
CLKBUFX1 gbuf_d_10(.A(g26135), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(n_344));
INVX1 g59420(.A (g27380), .Y (n_8180));
INVX1 g59422(.A (g26135), .Y (n_8178));
NAND4X1 g59421(.A (n_876), .B (n_8175), .C (n_1455), .D (n_980), .Y(g27380));
NAND3X1 g59423(.A (n_8176), .B (n_1199), .C (n_1172), .Y (g26135));
OAI21X1 g59424(.A0 (n_412), .A1 (n_296), .B0 (n_8174), .Y (g25489));
NOR2X1 g59425(.A (n_1458), .B (n_8173), .Y (n_8176));
AOI22X1 g59426(.A0 (n_519), .A1 (n_744), .B0 (n_696), .B1 (n_8169),.Y (n_8175));
MX2X1 g59427(.A (n_8172), .B (n_495), .S0 (g3147), .Y (n_8174));
NAND4X1 g59428(.A (n_8171), .B (n_1082), .C (n_912), .D (n_1465), .Y(n_8173));
AOI21X1 g59429(.A0 (n_8170), .A1 (n_324), .B0 (n_2326), .Y (n_8172));
AOI22X1 g59430(.A0 (n_7712), .A1 (n_2188), .B0 (n_2187), .B1(n_8170), .Y (n_8171));
AOI22X1 g59431(.A0 (g3114), .A1 (n_8170), .B0 (g3120), .B1 (n_2186),.Y (n_8169));
NAND2X1 g59432(.A (g2992), .B (g2991), .Y (n_8170));
CLKBUFX1 gbuf_d_11(.A(n_8167), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(g8258));
CLKBUFX1 gbuf_d_12(.A(n_8168), .Y(d_out_12));
CLKBUFX1 gbuf_qn_12(.A(qn_in_12), .Y(g2991));
XOR2X1 g59435(.A (g2990), .B (n_8166), .Y (n_8168));
XOR2X1 g59436(.A (n_8163), .B (n_8166), .Y (n_8167));
CLKBUFX1 gbuf_d_13(.A(n_8164), .Y(d_out_13));
CLKBUFX1 gbuf_q_13(.A(q_in_13), .Y(g8267));
XOR2X1 g59437(.A (n_8159), .B (n_8160), .Y (n_8166));
CLKBUFX1 gbuf_d_14(.A(n_8161), .Y(d_out_14));
CLKBUFX1 gbuf_q_14(.A(q_in_14), .Y(g2990));
CLKBUFX1 gbuf_d_15(.A(n_8165), .Y(d_out_15));
CLKBUFX1 gbuf_qn_15(.A(qn_in_15), .Y(g2992));
XOR2X1 g59442(.A (g3083), .B (n_8162), .Y (n_8165));
XOR2X1 g59445(.A (n_8163), .B (n_8162), .Y (n_8164));
MX2X1 g59441(.A (g3061), .B (g2997), .S0 (g2987), .Y (n_8161));
XOR2X1 g59443(.A (n_8155), .B (n_8158), .Y (n_8160));
XOR2X1 g59444(.A (n_8156), .B (n_8157), .Y (n_8159));
CLKBUFX1 gbuf_d_16(.A(n_8154), .Y(d_out_16));
CLKBUFX1 gbuf_q_16(.A(q_in_16), .Y(g2997));
XOR2X1 g59451(.A (n_8151), .B (n_8153), .Y (n_8162));
XOR2X1 g59447(.A (g8260), .B (g8263), .Y (n_8158));
XOR2X1 g59449(.A (g8265), .B (g8266), .Y (n_8157));
XOR2X1 g59450(.A (g8262), .B (g8264), .Y (n_8156));
XOR2X1 g59448(.A (g8259), .B (g8261), .Y (n_8155));
CLKBUFX1 gbuf_d_17(.A(n_8152), .Y(d_out_17));
CLKBUFX1 gbuf_q_17(.A(q_in_17), .Y(g3083));
NAND3X1 g59453(.A (n_7930), .B (n_8099), .C (n_8150), .Y (n_8154));
XOR2X1 g59463(.A (n_8142), .B (n_8147), .Y (n_8153));
CLKBUFX1 gbuf_d_18(.A(n_8143), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(g8262));
CLKBUFX1 gbuf_d_19(.A(n_8145), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(g8260));
CLKBUFX1 gbuf_d_20(.A(n_8146), .Y(d_out_20));
CLKBUFX1 gbuf_q_20(.A(q_in_20), .Y(g8263));
CLKBUFX1 gbuf_d_21(.A(n_8144), .Y(d_out_21));
CLKBUFX1 gbuf_q_21(.A(q_in_21), .Y(g8265));
CLKBUFX1 gbuf_d_22(.A(n_8149), .Y(d_out_22));
CLKBUFX1 gbuf_q_22(.A(q_in_22), .Y(g8266));
CLKBUFX1 gbuf_d_23(.A(n_8148), .Y(d_out_23));
CLKBUFX1 gbuf_q_23(.A(q_in_23), .Y(g8264));
MX2X1 g59462(.A (g3051), .B (g3070), .S0 (g2987), .Y (n_8152));
XOR2X1 g59464(.A (n_8141), .B (n_8140), .Y (n_8151));
CLKBUFX1 gbuf_d_24(.A(n_8138), .Y(d_out_24));
CLKBUFX1 gbuf_q_24(.A(q_in_24), .Y(g8261));
CLKBUFX1 gbuf_d_25(.A(n_8139), .Y(d_out_25));
CLKBUFX1 gbuf_q_25(.A(q_in_25), .Y(g8259));
NAND3X1 g59465(.A (n_4050), .B (n_8137), .C (n_8136), .Y (n_8150));
MX2X1 g59472(.A (g3052), .B (g3071), .S0 (g2987), .Y (n_8149));
MX2X1 g59473(.A (g3055), .B (g3073), .S0 (g2987), .Y (n_8148));
XOR2X1 g59475(.A (g8270), .B (g8271), .Y (n_8147));
MX2X1 g59467(.A (g3057), .B (g3075), .S0 (g2987), .Y (n_8146));
MX2X1 g59468(.A (g3058), .B (g3076), .S0 (g2987), .Y (n_8145));
MX2X1 g59469(.A (g3053), .B (g3072), .S0 (g2987), .Y (n_8144));
MX2X1 g59471(.A (g3056), .B (g3074), .S0 (g2987), .Y (n_8143));
CLKBUFX1 gbuf_d_26(.A(n_8135), .Y(d_out_26));
CLKBUFX1 gbuf_q_26(.A(q_in_26), .Y(g3070));
XOR2X1 g59476(.A (g8268), .B (g8269), .Y (n_8142));
XOR2X1 g59477(.A (g8274), .B (g8275), .Y (n_8141));
XOR2X1 g59478(.A (g8272), .B (g8273), .Y (n_8140));
MX2X1 g59466(.A (g3060), .B (g3078), .S0 (g2987), .Y (n_8139));
MX2X1 g59470(.A (g3059), .B (g3077), .S0 (g2987), .Y (n_8138));
NAND2X1 g59487(.A (n_8134), .B (n_8132), .Y (n_8137));
CLKBUFX1 gbuf_d_27(.A(n_8123), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(g3072));
CLKBUFX1 gbuf_d_28(.A(n_8129), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(g3074));
CLKBUFX1 gbuf_d_29(.A(n_8130), .Y(d_out_29));
CLKBUFX1 gbuf_q_29(.A(q_in_29), .Y(g3071));
CLKBUFX1 gbuf_d_30(.A(n_8126), .Y(d_out_30));
CLKBUFX1 gbuf_q_30(.A(q_in_30), .Y(g3073));
CLKBUFX1 gbuf_d_31(.A(n_8125), .Y(d_out_31));
CLKBUFX1 gbuf_q_31(.A(q_in_31), .Y(g3076));
CLKBUFX1 gbuf_d_32(.A(n_8127), .Y(d_out_32));
CLKBUFX1 gbuf_q_32(.A(q_in_32), .Y(g3075));
NAND2X1 g59488(.A (n_8133), .B (n_8131), .Y (n_8136));
NAND2X1 g59489(.A (n_8122), .B (n_7730), .Y (n_8135));
CLKBUFX1 gbuf_d_33(.A(n_8121), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(g8270));
CLKBUFX1 gbuf_d_34(.A(n_8120), .Y(d_out_34));
CLKBUFX1 gbuf_q_34(.A(q_in_34), .Y(g8271));
CLKBUFX1 gbuf_d_35(.A(n_8119), .Y(d_out_35));
CLKBUFX1 gbuf_q_35(.A(q_in_35), .Y(g_12763));
CLKBUFX1 gbuf_d_36(.A(n_8117), .Y(d_out_36));
CLKBUFX1 gbuf_q_36(.A(q_in_36), .Y(g_14632));
CLKBUFX1 gbuf_d_37(.A(n_8118), .Y(d_out_37));
CLKBUFX1 gbuf_q_37(.A(q_in_37), .Y(g_10841));
CLKBUFX1 gbuf_d_38(.A(n_8112), .Y(d_out_38));
CLKBUFX1 gbuf_q_38(.A(q_in_38), .Y(g3078));
CLKBUFX1 gbuf_d_39(.A(n_8113), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(g3077));
CLKBUFX1 gbuf_d_40(.A(n_8105), .Y(d_out_40));
CLKBUFX1 gbuf_q_40(.A(q_in_40), .Y(g8268));
CLKBUFX1 gbuf_d_41(.A(n_8110), .Y(d_out_41));
CLKBUFX1 gbuf_q_41(.A(q_in_41), .Y(g8269));
CLKBUFX1 gbuf_d_42(.A(n_8109), .Y(d_out_42));
CLKBUFX1 gbuf_q_42(.A(q_in_42), .Y(g8272));
CLKBUFX1 gbuf_d_43(.A(n_8108), .Y(d_out_43));
CLKBUFX1 gbuf_q_43(.A(q_in_43), .Y(g8273));
CLKBUFX1 gbuf_d_44(.A(n_8107), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(g8274));
CLKBUFX1 gbuf_d_45(.A(n_8106), .Y(d_out_45));
CLKBUFX1 gbuf_q_45(.A(q_in_45), .Y(g8275));
INVX1 g59509(.A (n_8133), .Y (n_8134));
INVX1 g59511(.A (n_8131), .Y (n_8132));
NAND2X1 g59498(.A (n_8104), .B (n_8128), .Y (n_8130));
NAND2X1 g59499(.A (n_8102), .B (n_8128), .Y (n_8129));
NAND2X1 g59500(.A (n_8101), .B (n_8124), .Y (n_8127));
INVX1 g59501(.A (n_8116), .Y (n_8126));
NAND2X1 g59503(.A (n_8100), .B (n_8124), .Y (n_8125));
INVX1 g59504(.A (n_8115), .Y (n_8123));
AOI22X1 g59506(.A0 (n_8098), .A1 (n_5322), .B0 (n_7914), .B1 (g1937),.Y (n_8122));
XOR2X1 g59510(.A (n_8097), .B (n_8068), .Y (n_8133));
XOR2X1 g59512(.A (n_8096), .B (n_8067), .Y (n_8131));
MX2X1 g59534(.A (g3049), .B (g3068), .S0 (g2987), .Y (n_8121));
MX2X1 g59535(.A (g3050), .B (g3069), .S0 (g2987), .Y (n_8120));
NAND2X1 g59550(.A (n_9658), .B (n_9659), .Y (n_8119));
NAND2X1 g59551(.A (n_9690), .B (n_9691), .Y (n_8118));
NAND2X1 g59552(.A (n_9688), .B (n_9689), .Y (n_8117));
AOI21X1 g59502(.A0 (n_8086), .A1 (n_8103), .B0 (n_8114), .Y (n_8116));
AOI21X1 g59505(.A0 (n_8087), .A1 (n_8103), .B0 (n_8114), .Y (n_8115));
OAI21X1 g59507(.A0 (n_7979), .A1 (n_8111), .B0 (n_8090), .Y (n_8113));
OAI21X1 g59508(.A0 (n_8072), .A1 (n_8111), .B0 (n_8088), .Y (n_8112));
MX2X1 g59533(.A (g3048), .B (g3067), .S0 (g2987), .Y (n_8110));
MX2X1 g59536(.A (g3046), .B (g3065), .S0 (g2987), .Y (n_8109));
MX2X1 g59537(.A (g3045), .B (g3064), .S0 (g2987), .Y (n_8108));
MX2X1 g59538(.A (g3044), .B (g3063), .S0 (g2987), .Y (n_8107));
MX2X1 g59539(.A (g3043), .B (g3062), .S0 (g2987), .Y (n_8106));
MX2X1 g59540(.A (g3047), .B (g3066), .S0 (g2987), .Y (n_8105));
CLKBUFX1 gbuf_d_46(.A(n_8076), .Y(d_out_46));
CLKBUFX1 gbuf_q_46(.A(q_in_46), .Y(g267));
CLKBUFX1 gbuf_d_47(.A(n_8075), .Y(d_out_47));
CLKBUFX1 gbuf_q_47(.A(q_in_47), .Y(g270));
CLKBUFX1 gbuf_d_48(.A(n_8074), .Y(d_out_48));
CLKBUFX1 gbuf_q_48(.A(q_in_48), .Y(g273));
CLKBUFX1 gbuf_d_49(.A(n_8066), .Y(d_out_49));
CLKBUFX1 gbuf_q_49(.A(q_in_49), .Y(g_20070));
CLKBUFX1 gbuf_d_50(.A(n_8065), .Y(d_out_50));
CLKBUFX1 gbuf_q_50(.A(q_in_50), .Y(g_26724));
CLKBUFX1 gbuf_d_51(.A(n_8063), .Y(d_out_51));
CLKBUFX1 gbuf_q_51(.A(q_in_51), .Y(g_16638));
CLKBUFX1 gbuf_d_52(.A(n_8071), .Y(d_out_52));
CLKBUFX1 gbuf_q_52(.A(q_in_52), .Y(g_24437));
CLKBUFX1 gbuf_d_53(.A(n_8070), .Y(d_out_53));
CLKBUFX1 gbuf_q_53(.A(q_in_53), .Y(g_30665));
CLKBUFX1 gbuf_d_54(.A(n_8069), .Y(d_out_54));
CLKBUFX1 gbuf_q_54(.A(q_in_54), .Y(g_26067));
CLKBUFX1 gbuf_d_55(.A(n_8079), .Y(d_out_55));
CLKBUFX1 gbuf_q_55(.A(q_in_55), .Y(g231));
CLKBUFX1 gbuf_d_56(.A(n_8078), .Y(d_out_56));
CLKBUFX1 gbuf_q_56(.A(q_in_56), .Y(g234));
CLKBUFX1 gbuf_d_57(.A(n_8077), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(g237));
NAND2X1 g59526(.A (n_8064), .B (n_8103), .Y (n_8104));
NAND2X1 g59527(.A (n_8083), .B (n_8103), .Y (n_8102));
NAND2X1 g59528(.A (n_8082), .B (n_8103), .Y (n_8101));
NAND2X1 g59529(.A (n_8080), .B (n_8103), .Y (n_8100));
OR2X1 g59530(.A (n_8073), .B (n_300), .Y (n_8099));
CLKBUFX1 gbuf_d_58(.A(n_8062), .Y(d_out_58));
CLKBUFX1 gbuf_qn_58(.A(qn_in_58), .Y(g2380));
CLKBUFX1 gbuf_d_59(.A(n_9518), .Y(d_out_59));
CLKBUFX1 gbuf_q_59(.A(q_in_59), .Y(g2390));
CLKBUFX1 gbuf_d_60(.A(n_8060), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(g2391));
CLKBUFX1 gbuf_d_61(.A(n_8059), .Y(d_out_61));
CLKBUFX1 gbuf_q_61(.A(q_in_61), .Y(g2392));
CLKBUFX1 gbuf_d_62(.A(n_8058), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(g1696));
CLKBUFX1 gbuf_d_63(.A(n_8056), .Y(d_out_63));
CLKBUFX1 gbuf_q_63(.A(q_in_63), .Y(g1697));
CLKBUFX1 gbuf_d_64(.A(n_8053), .Y(d_out_64));
CLKBUFX1 gbuf_q_64(.A(q_in_64), .Y(g1698));
CLKBUFX1 gbuf_d_65(.A(n_8048), .Y(d_out_65));
CLKBUFX1 gbuf_q_65(.A(q_in_65), .Y(g_18003));
CLKBUFX1 gbuf_d_66(.A(n_8047), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(g_18819));
CLKBUFX1 gbuf_d_67(.A(n_8045), .Y(d_out_67));
CLKBUFX1 gbuf_q_67(.A(q_in_67), .Y(g_22281));
XOR2X1 g59549(.A (n_7995), .B (n_8037), .Y (n_8098));
NAND2X1 g59563(.A (n_8052), .B (n_8051), .Y (n_8097));
NAND2X2 g59565(.A (n_8050), .B (n_8049), .Y (n_8096));
CLKBUFX1 gbuf_d_68(.A(n_8057), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(g3068));
CLKBUFX1 gbuf_d_69(.A(n_8055), .Y(d_out_69));
CLKBUFX1 gbuf_q_69(.A(q_in_69), .Y(g3069));
NAND2X1 g59642(.A (n_8092), .B (g5437), .Y (n_9658));
NAND2X1 g59643(.A (n_8092), .B (g6447), .Y (n_9690));
NAND2X1 g59644(.A (n_8092), .B (g401), .Y (n_9688));
OAI21X1 g59531(.A0 (n_8020), .A1 (n_7909), .B0 (n_8103), .Y (n_8090));
OAI21X1 g59532(.A0 (n_8018), .A1 (n_7908), .B0 (n_8103), .Y (n_8088));
AOI22X1 g59543(.A0 (n_1163), .A1 (n_8085), .B0 (n_7974), .B1(n_8084), .Y (n_8087));
CLKBUFX1 gbuf_d_70(.A(n_8038), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(g1654));
CLKBUFX1 gbuf_d_71(.A(n_8039), .Y(d_out_71));
CLKBUFX1 gbuf_q_71(.A(q_in_71), .Y(g1648));
CLKBUFX1 gbuf_d_72(.A(n_8040), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(g1651));
CLKBUFX1 gbuf_d_73(.A(n_8044), .Y(d_out_73));
CLKBUFX1 gbuf_q_73(.A(q_in_73), .Y(g240));
CLKBUFX1 gbuf_d_74(.A(n_8043), .Y(d_out_74));
CLKBUFX1 gbuf_q_74(.A(q_in_74), .Y(g243));
AOI22X1 g59544(.A0 (n_1049), .A1 (n_8085), .B0 (n_7971), .B1(n_8084), .Y (n_8086));
CLKBUFX1 gbuf_d_75(.A(n_9321), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(g246));
AOI22X1 g59545(.A0 (n_1044), .A1 (n_8085), .B0 (n_7969), .B1(n_8084), .Y (n_8083));
AOI22X1 g59546(.A0 (n_1204), .A1 (n_8085), .B0 (n_7966), .B1(n_8084), .Y (n_8082));
AOI22X1 g59547(.A0 (n_1159), .A1 (n_8085), .B0 (n_7963), .B1(n_8084), .Y (n_8080));
NAND2X1 g59731(.A (n_9618), .B (n_9619), .Y (n_8079));
NAND2X2 g59736(.A (n_9594), .B (n_9595), .Y (n_8078));
NAND2X1 g59737(.A (n_9620), .B (n_9621), .Y (n_8077));
NAND2X2 g59750(.A (n_8225), .B (n_8226), .Y (n_8076));
NAND2X2 g59751(.A (n_8227), .B (n_8228), .Y (n_8075));
NAND2X2 g59752(.A (n_8229), .B (n_8230), .Y (n_8074));
XOR2X1 g59562(.A (n_7978), .B (n_8072), .Y (n_8073));
NAND2X1 g59758(.A (n_1581), .B (n_8025), .Y (n_8071));
NAND2X1 g59759(.A (n_3194), .B (n_8023), .Y (n_8070));
NAND2X1 g59760(.A (n_5199), .B (n_8021), .Y (n_8069));
MX2X1 g59564(.A (n_7969), .B (n_7968), .S0 (n_7970), .Y (n_8068));
MX2X1 g59566(.A (n_7960), .B (n_8017), .S0 (n_8019), .Y (n_8067));
CLKBUFX1 gbuf_d_76(.A(n_8010), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(g3062));
CLKBUFX1 gbuf_d_77(.A(n_8011), .Y(d_out_77));
CLKBUFX1 gbuf_q_77(.A(q_in_77), .Y(g3063));
CLKBUFX1 gbuf_d_78(.A(n_8009), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(g3064));
CLKBUFX1 gbuf_d_79(.A(n_8008), .Y(d_out_79));
CLKBUFX1 gbuf_q_79(.A(q_in_79), .Y(g3065));
CLKBUFX1 gbuf_d_80(.A(n_8005), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(g3067));
CLKBUFX1 gbuf_d_81(.A(n_8006), .Y(d_out_81));
CLKBUFX1 gbuf_q_81(.A(q_in_81), .Y(g3066));
NAND2X1 g59705(.A (n_1586), .B (n_8036), .Y (n_8066));
NAND2X1 g59706(.A (n_8259), .B (n_8260), .Y (n_8065));
AOI22X1 g59542(.A0 (n_1158), .A1 (n_8085), .B0 (n_7977), .B1(n_8084), .Y (n_8064));
NAND2X1 g59707(.A (n_8256), .B (n_8257), .Y (n_8063));
CLKBUFX1 gbuf_d_82(.A(n_7987), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(g_5496));
CLKBUFX1 gbuf_d_83(.A(n_7985), .Y(d_out_83));
CLKBUFX1 gbuf_q_83(.A(q_in_83), .Y(g_10959));
CLKBUFX1 gbuf_d_84(.A(n_7981), .Y(d_out_84));
CLKBUFX1 gbuf_q_84(.A(q_in_84), .Y(g_24632));
CLKBUFX1 gbuf_d_85(.A(n_7996), .Y(d_out_85));
CLKBUFX1 gbuf_q_85(.A(q_in_85), .Y(g264));
CLKBUFX1 gbuf_d_86(.A(n_7955), .Y(d_out_86));
CLKBUFX1 gbuf_q_86(.A(q_in_86), .Y(g_25929));
CLKBUFX1 gbuf_d_87(.A(n_7956), .Y(d_out_87));
CLKBUFX1 gbuf_q_87(.A(q_in_87), .Y(g_30245));
CLKBUFX1 gbuf_d_88(.A(n_7953), .Y(d_out_88));
CLKBUFX1 gbuf_q_88(.A(q_in_88), .Y(g_19223));
CLKBUFX1 gbuf_d_89(.A(n_7952), .Y(d_out_89));
CLKBUFX1 gbuf_q_89(.A(q_in_89), .Y(g_28592));
CLKBUFX1 gbuf_d_90(.A(n_7951), .Y(d_out_90));
CLKBUFX1 gbuf_q_90(.A(q_in_90), .Y(g_13736));
CLKBUFX1 gbuf_d_91(.A(n_7998), .Y(d_out_91));
CLKBUFX1 gbuf_q_91(.A(q_in_91), .Y(g261));
CLKBUFX1 gbuf_d_92(.A(n_7949), .Y(d_out_92));
CLKBUFX1 gbuf_q_92(.A(q_in_92), .Y(g_19110));
CLKBUFX1 gbuf_d_93(.A(n_7999), .Y(d_out_93));
CLKBUFX1 gbuf_q_93(.A(q_in_93), .Y(g258));
CLKBUFX1 gbuf_d_94(.A(n_8003), .Y(d_out_94));
CLKBUFX1 gbuf_q_94(.A(q_in_94), .Y(g249));
CLKBUFX1 gbuf_d_95(.A(n_8002), .Y(d_out_95));
CLKBUFX1 gbuf_q_95(.A(q_in_95), .Y(g252));
CLKBUFX1 gbuf_d_96(.A(n_8000), .Y(d_out_96));
CLKBUFX1 gbuf_q_96(.A(q_in_96), .Y(g255));
OAI21X1 g59548(.A0 (n_7928), .A1 (g2374), .B0 (n_7253), .Y (n_8062));
NAND2X1 g59555(.A (n_3199), .B (n_7990), .Y (n_8060));
NAND2X1 g59556(.A (n_5196), .B (n_7988), .Y (n_8059));
NAND2X1 g59559(.A (n_1587), .B (n_7986), .Y (n_8058));
OAI21X1 g59753(.A0 (n_7913), .A1 (n_8054), .B0 (n_7994), .Y (n_8057));
NAND2X1 g59560(.A (n_3431), .B (n_7983), .Y (n_8056));
OAI21X1 g59754(.A0 (n_7912), .A1 (n_8054), .B0 (n_7993), .Y (n_8055));
NAND2X1 g59561(.A (n_9587), .B (n_9588), .Y (n_8053));
NAND2X1 g59635(.A (n_7976), .B (n_7972), .Y (n_8052));
NAND2X1 g59636(.A (n_7977), .B (n_7973), .Y (n_8051));
NAND2X1 g59637(.A (n_7965), .B (n_7961), .Y (n_8050));
NAND2X1 g59638(.A (n_7966), .B (n_7962), .Y (n_8049));
INVX1 g59686(.A (n_8012), .Y (n_8092));
MX2X1 g59967(.A (g_18003), .B (n_8585), .S0 (n_8024), .Y (n_8048));
MX2X1 g59968(.A (g_18819), .B (n_8585), .S0 (g6313), .Y (n_8047));
MX2X1 g59970(.A (g_22281), .B (n_8585), .S0 (n_9315), .Y (n_8045));
CLKBUFX1 gbuf_d_97(.A(n_7945), .Y(d_out_97));
CLKBUFX1 gbuf_q_97(.A(q_in_97), .Y(g2342));
CLKBUFX1 gbuf_d_98(.A(n_7944), .Y(d_out_98));
CLKBUFX1 gbuf_q_98(.A(q_in_98), .Y(g2345));
CLKBUFX1 gbuf_d_99(.A(n_7943), .Y(d_out_99));
CLKBUFX1 gbuf_q_99(.A(q_in_99), .Y(g2348));
CLKBUFX1 gbuf_d_100(.A(n_7948), .Y(d_out_100));
CLKBUFX1 gbuf_q_100(.A(q_in_100), .Y(g2315));
CLKBUFX1 gbuf_d_101(.A(n_7947), .Y(d_out_101));
CLKBUFX1 gbuf_q_101(.A(q_in_101), .Y(g2318));
CLKBUFX1 gbuf_d_102(.A(n_7946), .Y(d_out_102));
CLKBUFX1 gbuf_q_102(.A(q_in_102), .Y(g2321));
CLKBUFX1 gbuf_d_103(.A(n_7940), .Y(d_out_103));
CLKBUFX1 gbuf_q_103(.A(q_in_103), .Y(g1627));
CLKBUFX1 gbuf_d_104(.A(n_7942), .Y(d_out_104));
CLKBUFX1 gbuf_q_104(.A(q_in_104), .Y(g1621));
CLKBUFX1 gbuf_d_105(.A(n_7941), .Y(d_out_105));
CLKBUFX1 gbuf_q_105(.A(q_in_105), .Y(g1624));
OAI21X1 g59743(.A0 (n_9322), .A1 (n_1382), .B0 (n_1580), .Y (n_8044));
OAI21X1 g59745(.A0 (n_9322), .A1 (n_3195), .B0 (n_3200), .Y (n_8043));
NAND2X2 g59747(.A (n_8219), .B (n_8220), .Y (n_8040));
NAND2X2 g59748(.A (n_8217), .B (n_8218), .Y (n_8039));
NAND2X2 g59749(.A (n_8215), .B (n_8216), .Y (n_8038));
XOR2X1 g59768(.A (n_7897), .B (n_7911), .Y (n_8037));
NAND2X1 g59844(.A (n_8034), .B (g6231), .Y (n_8036));
NAND2X1 g59845(.A (n_8034), .B (n_8028), .Y (n_8259));
NAND2X1 g59846(.A (n_8034), .B (n_9312), .Y (n_8256));
NAND2X1 g59863(.A (n_8029), .B (g6231), .Y (n_9618));
NAND2X1 g59865(.A (n_8029), .B (n_8028), .Y (n_9594));
NAND2X1 g59866(.A (n_8029), .B (n_9312), .Y (n_9620));
NAND2X1 g59875(.A (n_8022), .B (n_8024), .Y (n_8025));
NAND2X1 g59876(.A (n_8022), .B (n_8028), .Y (n_8023));
NAND2X1 g59877(.A (n_8022), .B (n_9312), .Y (n_8021));
AND2X1 g59640(.A (n_8019), .B (n_8084), .Y (n_8020));
AND2X1 g59641(.A (n_8017), .B (n_8084), .Y (n_8018));
NAND2X1 g59888(.A (n_8014), .B (g6231), .Y (n_8225));
NAND2X1 g59889(.A (n_8014), .B (n_8028), .Y (n_8227));
NAND2X1 g59890(.A (n_8014), .B (n_9312), .Y (n_8229));
NAND3X1 g59687(.A (n_7891), .B (n_7865), .C (n_7906), .Y (n_8012));
INVX1 g59693(.A (n_7959), .Y (n_8011));
NAND2X1 g59695(.A (n_7939), .B (n_8007), .Y (n_8010));
INVX1 g59696(.A (n_7958), .Y (n_8009));
NAND2X1 g59698(.A (n_7938), .B (n_8007), .Y (n_8008));
NAND2X1 g59699(.A (n_7937), .B (n_8004), .Y (n_8006));
NAND2X1 g59700(.A (n_7936), .B (n_8004), .Y (n_8005));
CLKBUFX1 gbuf_d_106(.A(n_7935), .Y(d_out_106));
CLKBUFX1 gbuf_q_106(.A(q_in_106), .Y(g3061));
CLKBUFX1 gbuf_d_107(.A(n_7923), .Y(d_out_107));
CLKBUFX1 gbuf_q_107(.A(q_in_107), .Y(g2273));
CLKBUFX1 gbuf_d_108(.A(n_7926), .Y(d_out_108));
CLKBUFX1 gbuf_q_108(.A(q_in_108), .Y(g2270));
CLKBUFX1 gbuf_d_109(.A(n_7925), .Y(d_out_109));
CLKBUFX1 gbuf_q_109(.A(q_in_109), .Y(g2276));
CLKBUFX1 gbuf_d_110(.A(n_7919), .Y(d_out_110));
CLKBUFX1 gbuf_q_110(.A(q_in_110), .Y(g2309));
CLKBUFX1 gbuf_d_111(.A(n_7918), .Y(d_out_111));
CLKBUFX1 gbuf_q_111(.A(q_in_111), .Y(g2312));
CLKBUFX1 gbuf_d_112(.A(n_7921), .Y(d_out_112));
CLKBUFX1 gbuf_q_112(.A(q_in_112), .Y(g2306));
CLKBUFX1 gbuf_d_113(.A(n_7922), .Y(d_out_113));
CLKBUFX1 gbuf_q_113(.A(q_in_113), .Y(g1579));
CLKBUFX1 gbuf_d_114(.A(n_7920), .Y(d_out_114));
CLKBUFX1 gbuf_q_114(.A(q_in_114), .Y(g1582));
CLKBUFX1 gbuf_d_115(.A(n_7927), .Y(d_out_115));
CLKBUFX1 gbuf_q_115(.A(q_in_115), .Y(g1576));
CLKBUFX1 gbuf_d_116(.A(n_7917), .Y(d_out_116));
CLKBUFX1 gbuf_q_116(.A(q_in_116), .Y(g1612));
CLKBUFX1 gbuf_d_117(.A(n_7916), .Y(d_out_117));
CLKBUFX1 gbuf_q_117(.A(q_in_117), .Y(g1615));
CLKBUFX1 gbuf_d_118(.A(n_7915), .Y(d_out_118));
CLKBUFX1 gbuf_q_118(.A(q_in_118), .Y(g1618));
MX2X1 g60016(.A (g249), .B (n_8001), .S0 (n_8024), .Y (n_8003));
MX2X1 g60017(.A (g252), .B (n_8001), .S0 (g6313), .Y (n_8002));
MX2X1 g60018(.A (g255), .B (n_8001), .S0 (n_9315), .Y (n_8000));
MX2X1 g60019(.A (g258), .B (n_7997), .S0 (n_8024), .Y (n_7999));
MX2X1 g60020(.A (g261), .B (n_7997), .S0 (g6313), .Y (n_7998));
MX2X1 g60021(.A (g264), .B (n_7997), .S0 (n_9315), .Y (n_7996));
XOR2X1 g59767(.A (n_7899), .B (n_7898), .Y (n_7995));
OAI21X1 g59842(.A0 (n_7896), .A1 (n_7620), .B0 (n_7992), .Y (n_7994));
OAI21X1 g59843(.A0 (n_7894), .A1 (n_7619), .B0 (n_7992), .Y (n_7993));
NAND2X1 g59646(.A (n_9392), .B (n_3085), .Y (n_7990));
NAND2X1 g59647(.A (n_9392), .B (n_4985), .Y (n_7988));
MX2X1 g59894(.A (g_5496), .B (n_7984), .S0 (n_6914), .Y (n_7987));
NAND2X1 g59648(.A (n_7982), .B (n_1483), .Y (n_7986));
MX2X1 g59895(.A (g_10959), .B (n_7984), .S0 (g6447), .Y (n_7985));
NAND2X1 g59649(.A (n_7982), .B (n_3190), .Y (n_7983));
MX2X1 g59896(.A (g_24632), .B (n_7984), .S0 (n_6917), .Y (n_7981));
NAND2X1 g59650(.A (n_7982), .B (n_6832), .Y (n_9587));
INVX1 g59663(.A (n_7978), .Y (n_7979));
AOI21X1 g59665(.A0 (n_3687), .A1 (n_4894), .B0 (n_7910), .Y (n_8072));
INVX2 g59666(.A (n_7976), .Y (n_7977));
INVX1 g59669(.A (n_7973), .Y (n_7974));
INVX1 g59670(.A (n_7973), .Y (n_7972));
INVX1 g59672(.A (n_7970), .Y (n_7971));
INVX2 g59674(.A (n_7968), .Y (n_7969));
INVX2 g59677(.A (n_7965), .Y (n_7966));
INVX1 g59680(.A (n_7962), .Y (n_7963));
INVX1 g59681(.A (n_7962), .Y (n_7961));
INVX1 g59684(.A (n_8017), .Y (n_7960));
AOI21X1 g59694(.A0 (n_7862), .A1 (n_7992), .B0 (n_7957), .Y (n_7959));
AOI21X1 g59697(.A0 (n_7860), .A1 (n_7992), .B0 (n_7957), .Y (n_7958));
MX2X1 g59959(.A (g_30245), .B (n_7954), .S0 (n_8024), .Y (n_7956));
MX2X1 g59960(.A (g_25929), .B (n_7954), .S0 (g6313), .Y (n_7955));
MX2X1 g59961(.A (g_19223), .B (n_7954), .S0 (n_9315), .Y (n_7953));
MX2X1 g59964(.A (g_28592), .B (n_7950), .S0 (n_8024), .Y (n_7952));
MX2X1 g59965(.A (g_13736), .B (n_7950), .S0 (g6313), .Y (n_7951));
MX2X1 g59966(.A (g_19110), .B (n_7950), .S0 (n_9315), .Y (n_7949));
CLKBUFX1 gbuf_d_119(.A(n_7902), .Y(d_out_119));
CLKBUFX1 gbuf_q_119(.A(q_in_119), .Y(g954));
CLKBUFX1 gbuf_d_120(.A(n_7901), .Y(d_out_120));
CLKBUFX1 gbuf_q_120(.A(q_in_120), .Y(g957));
CLKBUFX1 gbuf_d_121(.A(n_7900), .Y(d_out_121));
CLKBUFX1 gbuf_q_121(.A(q_in_121), .Y(g960));
CLKBUFX1 gbuf_d_122(.A(n_7889), .Y(d_out_122));
CLKBUFX1 gbuf_q_122(.A(q_in_122), .Y(g2297));
CLKBUFX1 gbuf_d_123(.A(n_7888), .Y(d_out_123));
CLKBUFX1 gbuf_q_123(.A(q_in_123), .Y(g2300));
CLKBUFX1 gbuf_d_124(.A(n_7886), .Y(d_out_124));
CLKBUFX1 gbuf_q_124(.A(q_in_124), .Y(g2303));
CLKBUFX1 gbuf_d_125(.A(n_7885), .Y(d_out_125));
CLKBUFX1 gbuf_q_125(.A(q_in_125), .Y(g1603));
CLKBUFX1 gbuf_d_126(.A(n_7884), .Y(d_out_126));
CLKBUFX1 gbuf_q_126(.A(q_in_126), .Y(g1606));
CLKBUFX1 gbuf_d_127(.A(n_7882), .Y(d_out_127));
CLKBUFX1 gbuf_q_127(.A(q_in_127), .Y(g1609));
CLKBUFX1 gbuf_d_128(.A(n_7849), .Y(d_out_128));
CLKBUFX1 gbuf_q_128(.A(q_in_128), .Y(g1686));
INVX1 g59996(.A (n_7924), .Y (n_8029));
NAND2X2 g59729(.A (n_8243), .B (n_8244), .Y (n_7948));
NAND2X2 g59730(.A (n_8245), .B (n_8246), .Y (n_7947));
NAND2X2 g59732(.A (n_8247), .B (n_8248), .Y (n_7946));
NAND2X2 g59733(.A (n_8273), .B (n_8274), .Y (n_7945));
NAND2X1 g59734(.A (n_8275), .B (n_8276), .Y (n_7944));
NAND2X1 g59735(.A (n_8262), .B (n_8263), .Y (n_7943));
NAND2X1 g59741(.A (n_9614), .B (n_9615), .Y (n_7942));
NAND2X1 g59742(.A (n_9573), .B (n_9574), .Y (n_7941));
NAND2X1 g59744(.A (n_4390), .B (n_7871), .Y (n_7940));
NAND2X1 g59834(.A (n_7864), .B (n_7992), .Y (n_7939));
NAND2X1 g59835(.A (n_7857), .B (n_7992), .Y (n_7938));
NAND2X1 g59836(.A (n_7854), .B (n_7992), .Y (n_7937));
NAND2X1 g59837(.A (n_7852), .B (n_7992), .Y (n_7936));
NAND2X2 g59639(.A (n_7846), .B (n_7398), .Y (n_7935));
NAND2X1 g59885(.A (n_7932), .B (n_1077), .Y (n_8217));
NAND2X1 g59886(.A (n_7932), .B (n_2422), .Y (n_8219));
NAND2X1 g59887(.A (n_7932), .B (n_4125), .Y (n_8215));
OR2X1 g59893(.A (n_7866), .B (n_1374), .Y (n_7930));
NAND3X1 g59664(.A (n_5108), .B (n_5343), .C (n_7929), .Y (n_7978));
NAND3X1 g59668(.A (n_4706), .B (n_4750), .C (n_7929), .Y (n_7976));
INVX1 g59927(.A (n_7905), .Y (n_8022));
NAND3X1 g59671(.A (n_4704), .B (n_4749), .C (n_7929), .Y (n_7973));
NAND3X1 g59673(.A (n_4895), .B (n_4748), .C (n_7929), .Y (n_7970));
NAND3X1 g59676(.A (n_4703), .B (n_4747), .C (n_7929), .Y (n_7968));
NAND3X1 g59679(.A (n_4701), .B (n_4746), .C (n_7929), .Y (n_7965));
AOI21X1 g59939(.A0 (n_7569), .A1 (n_8582), .B0 (n_7890), .Y (n_8014));
NAND3X1 g59682(.A (n_4700), .B (n_4745), .C (n_7929), .Y (n_7962));
NAND3X1 g59683(.A (n_4699), .B (n_4744), .C (n_7929), .Y (n_8019));
NAND3X1 g59685(.A (n_4697), .B (n_4743), .C (n_7929), .Y (n_8017));
INVX1 g59962(.A (n_9488), .Y (n_8034));
OR2X1 g59702(.A (n_7881), .B (n_8103), .Y (n_8128));
MX2X1 g59703(.A (g2380), .B (n_7848), .S0 (n_2180), .Y (n_7928));
CLKBUFX1 gbuf_d_129(.A(n_7822), .Y(d_out_129));
CLKBUFX1 gbuf_q_129(.A(q_in_129), .Y(g1003));
CLKBUFX1 gbuf_d_130(.A(n_7821), .Y(d_out_130));
CLKBUFX1 gbuf_q_130(.A(q_in_130), .Y(g1004));
CLKBUFX1 gbuf_d_131(.A(n_7819), .Y(d_out_131));
CLKBUFX1 gbuf_q_131(.A(q_in_131), .Y(g1002));
CLKBUFX1 gbuf_d_132(.A(n_7795), .Y(d_out_132));
CLKBUFX1 gbuf_q_132(.A(q_in_132), .Y(g1699));
CLKBUFX1 gbuf_d_133(.A(n_7792), .Y(d_out_133));
CLKBUFX1 gbuf_q_133(.A(q_in_133), .Y(g1700));
CLKBUFX1 gbuf_d_134(.A(n_7794), .Y(d_out_134));
CLKBUFX1 gbuf_q_134(.A(q_in_134), .Y(g1701));
CLKBUFX1 gbuf_d_135(.A(n_7845), .Y(d_out_135));
CLKBUFX1 gbuf_q_135(.A(q_in_135), .Y(g2261));
CLKBUFX1 gbuf_d_136(.A(n_7844), .Y(d_out_136));
CLKBUFX1 gbuf_q_136(.A(q_in_136), .Y(g2264));
CLKBUFX1 gbuf_d_137(.A(n_7842), .Y(d_out_137));
CLKBUFX1 gbuf_q_137(.A(q_in_137), .Y(g2267));
CLKBUFX1 gbuf_d_138(.A(n_7841), .Y(d_out_138));
CLKBUFX1 gbuf_q_138(.A(q_in_138), .Y(g2279));
CLKBUFX1 gbuf_d_139(.A(n_7840), .Y(d_out_139));
CLKBUFX1 gbuf_q_139(.A(q_in_139), .Y(g2282));
CLKBUFX1 gbuf_d_140(.A(n_7838), .Y(d_out_140));
CLKBUFX1 gbuf_q_140(.A(q_in_140), .Y(g2285));
CLKBUFX1 gbuf_d_141(.A(n_7836), .Y(d_out_141));
CLKBUFX1 gbuf_q_141(.A(q_in_141), .Y(g1573));
CLKBUFX1 gbuf_d_142(.A(n_7837), .Y(d_out_142));
CLKBUFX1 gbuf_q_142(.A(q_in_142), .Y(g2288));
CLKBUFX1 gbuf_d_143(.A(n_7790), .Y(d_out_143));
CLKBUFX1 gbuf_q_143(.A(q_in_143), .Y(g1567));
CLKBUFX1 gbuf_d_144(.A(n_7835), .Y(d_out_144));
CLKBUFX1 gbuf_q_144(.A(q_in_144), .Y(g1570));
CLKBUFX1 gbuf_d_145(.A(n_7830), .Y(d_out_145));
CLKBUFX1 gbuf_q_145(.A(q_in_145), .Y(g1585));
CLKBUFX1 gbuf_d_146(.A(n_7829), .Y(d_out_146));
CLKBUFX1 gbuf_q_146(.A(q_in_146), .Y(g1588));
CLKBUFX1 gbuf_d_147(.A(n_7826), .Y(d_out_147));
CLKBUFX1 gbuf_q_147(.A(q_in_147), .Y(g1591));
CLKBUFX1 gbuf_d_148(.A(n_7827), .Y(d_out_148));
CLKBUFX1 gbuf_q_148(.A(q_in_148), .Y(g1594));
CLKBUFX1 gbuf_d_149(.A(n_7831), .Y(d_out_149));
CLKBUFX1 gbuf_q_149(.A(q_in_149), .Y(g2294));
CLKBUFX1 gbuf_d_150(.A(n_7823), .Y(d_out_150));
CLKBUFX1 gbuf_q_150(.A(q_in_150), .Y(g1600));
CLKBUFX1 gbuf_d_151(.A(n_7825), .Y(d_out_151));
CLKBUFX1 gbuf_q_151(.A(q_in_151), .Y(g1597));
CLKBUFX1 gbuf_d_152(.A(n_7833), .Y(d_out_152));
CLKBUFX1 gbuf_q_152(.A(q_in_152), .Y(g2291));
NAND2X1 g59720(.A (n_1401), .B (n_7808), .Y (n_7927));
NAND2X1 g59721(.A (n_9606), .B (n_9607), .Y (n_7926));
NAND2X1 g59722(.A (n_9602), .B (n_9603), .Y (n_7925));
NAND3X1 g59997(.A (n_9486), .B (n_7764), .C (n_8258), .Y (n_7924));
NAND2X1 g59723(.A (n_9600), .B (n_9601), .Y (n_7923));
NAND2X1 g59724(.A (n_9648), .B (n_9649), .Y (n_7922));
NAND2X1 g59725(.A (n_1403), .B (n_7807), .Y (n_7921));
NAND2X1 g59726(.A (n_4385), .B (n_7801), .Y (n_7920));
NAND2X1 g59727(.A (n_2563), .B (n_7806), .Y (n_7919));
NAND2X1 g59728(.A (n_9604), .B (n_9605), .Y (n_7918));
NAND2X1 g59738(.A (n_9622), .B (n_9623), .Y (n_7917));
NAND2X1 g59739(.A (n_9612), .B (n_9613), .Y (n_7916));
NAND2X1 g59740(.A (n_9624), .B (n_9625), .Y (n_7915));
XOR2X1 g60022(.A (n_7913), .B (n_7912), .Y (n_7914));
XOR2X1 g60025(.A (n_7893), .B (n_7895), .Y (n_7911));
NAND2X1 g59838(.A (n_5157), .B (n_7929), .Y (n_7910));
AOI21X1 g59891(.A0 (n_8085), .A1 (g2610), .B0 (n_8084), .Y (n_7909));
AOI21X1 g59892(.A0 (n_8085), .A1 (g2611), .B0 (n_8084), .Y (n_7908));
NAND2X1 g59918(.A (n_7817), .B (n_5099), .Y (n_7906));
NAND3X1 g59928(.A (n_9626), .B (n_7769), .C (n_9486), .Y (n_7905));
INVX1 g59691(.A (n_7847), .Y (n_7982));
AOI21X1 g59701(.A0 (n_6419), .A1 (n_7880), .B0 (n_8103), .Y (n_8114));
CLKBUFX1 gbuf_d_153(.A(n_7789), .Y(d_out_153));
CLKBUFX1 gbuf_q_153(.A(q_in_153), .Y(g888));
CLKBUFX1 gbuf_d_154(.A(n_7736), .Y(d_out_154));
CLKBUFX1 gbuf_q_154(.A(q_in_154), .Y(g882));
CLKBUFX1 gbuf_d_155(.A(n_7735), .Y(d_out_155));
CLKBUFX1 gbuf_q_155(.A(q_in_155), .Y(g885));
CLKBUFX1 gbuf_d_156(.A(n_7772), .Y(d_out_156));
CLKBUFX1 gbuf_q_156(.A(q_in_156), .Y(g909));
CLKBUFX1 gbuf_d_157(.A(n_7771), .Y(d_out_157));
CLKBUFX1 gbuf_q_157(.A(q_in_157), .Y(g912));
CLKBUFX1 gbuf_d_158(.A(n_7773), .Y(d_out_158));
CLKBUFX1 gbuf_q_158(.A(q_in_158), .Y(g915));
CLKBUFX1 gbuf_d_159(.A(n_7788), .Y(d_out_159));
CLKBUFX1 gbuf_q_159(.A(q_in_159), .Y(g918));
CLKBUFX1 gbuf_d_160(.A(n_7787), .Y(d_out_160));
CLKBUFX1 gbuf_q_160(.A(q_in_160), .Y(g921));
CLKBUFX1 gbuf_d_161(.A(n_7786), .Y(d_out_161));
CLKBUFX1 gbuf_q_161(.A(q_in_161), .Y(g924));
CLKBUFX1 gbuf_d_162(.A(n_7750), .Y(d_out_162));
CLKBUFX1 gbuf_q_162(.A(q_in_162), .Y(g2393));
CLKBUFX1 gbuf_d_163(.A(n_7749), .Y(d_out_163));
CLKBUFX1 gbuf_q_163(.A(q_in_163), .Y(g2394));
CLKBUFX1 gbuf_d_164(.A(n_7747), .Y(d_out_164));
CLKBUFX1 gbuf_q_164(.A(q_in_164), .Y(g2395));
CLKBUFX1 gbuf_d_165(.A(n_7744), .Y(d_out_165));
CLKBUFX1 gbuf_q_165(.A(q_in_165), .Y(g2333));
CLKBUFX1 gbuf_d_166(.A(n_7741), .Y(d_out_166));
CLKBUFX1 gbuf_q_166(.A(q_in_166), .Y(g2339));
CLKBUFX1 gbuf_d_167(.A(n_7743), .Y(d_out_167));
CLKBUFX1 gbuf_q_167(.A(q_in_167), .Y(g2336));
CLKBUFX1 gbuf_d_168(.A(n_7739), .Y(d_out_168));
CLKBUFX1 gbuf_q_168(.A(q_in_168), .Y(g1642));
CLKBUFX1 gbuf_d_169(.A(n_7737), .Y(d_out_169));
CLKBUFX1 gbuf_q_169(.A(q_in_169), .Y(g1645));
CLKBUFX1 gbuf_d_170(.A(n_7740), .Y(d_out_170));
CLKBUFX1 gbuf_q_170(.A(q_in_170), .Y(g1639));
CLKBUFX1 gbuf_d_171(.A(n_7785), .Y(d_out_171));
CLKBUFX1 gbuf_q_171(.A(q_in_171), .Y(g2324));
CLKBUFX1 gbuf_d_172(.A(n_7784), .Y(d_out_172));
CLKBUFX1 gbuf_q_172(.A(q_in_172), .Y(g2327));
CLKBUFX1 gbuf_d_173(.A(n_7782), .Y(d_out_173));
CLKBUFX1 gbuf_q_173(.A(q_in_173), .Y(g2330));
CLKBUFX1 gbuf_d_174(.A(n_7781), .Y(d_out_174));
CLKBUFX1 gbuf_q_174(.A(q_in_174), .Y(g1630));
CLKBUFX1 gbuf_d_175(.A(n_7780), .Y(d_out_175));
CLKBUFX1 gbuf_q_175(.A(q_in_175), .Y(g1633));
CLKBUFX1 gbuf_d_176(.A(n_7778), .Y(d_out_176));
CLKBUFX1 gbuf_q_176(.A(q_in_176), .Y(g1636));
NAND2X1 g59717(.A (n_8267), .B (n_8268), .Y (n_7902));
NAND2X2 g59718(.A (n_8269), .B (n_8270), .Y (n_7901));
NAND2X2 g59719(.A (n_8271), .B (n_8272), .Y (n_7900));
XOR2X1 g60023(.A (n_7855), .B (n_7858), .Y (n_7899));
XOR2X1 g60024(.A (n_7863), .B (n_7861), .Y (n_7898));
XOR2X1 g60026(.A (n_7851), .B (n_7853), .Y (n_7897));
AND2X1 g60044(.A (n_7895), .B (n_7892), .Y (n_7896));
AND2X1 g60045(.A (n_7893), .B (n_7892), .Y (n_7894));
AND2X1 g60046(.A (n_7762), .B (n_7891), .Y (n_7984));
NAND2X1 g60054(.A (n_7768), .B (n_9486), .Y (n_7890));
OAI21X1 g59761(.A0 (n_9010), .A1 (n_1305), .B0 (n_1389), .Y (n_7889));
OAI21X1 g59762(.A0 (n_9010), .A1 (n_7811), .B0 (n_2566), .Y (n_7888));
OAI21X1 g59763(.A0 (n_9011), .A1 (n_7809), .B0 (n_4135), .Y (n_7886));
OAI21X1 g59764(.A0 (n_7883), .A1 (n_1392), .B0 (n_1388), .Y (n_7885));
OAI21X1 g59765(.A0 (n_7883), .A1 (n_2433), .B0 (n_2687), .Y (n_7884));
OAI21X1 g59766(.A0 (n_7883), .A1 (n_7800), .B0 (n_4384), .Y (n_7882));
NOR2X1 g60104(.A (n_7756), .B (n_9196), .Y (n_8001));
AOI21X1 g60120(.A0 (n_6362), .A1 (n_8582), .B0 (n_7759), .Y (n_7954));
AOI21X1 g60121(.A0 (n_7205), .A1 (n_8582), .B0 (n_7757), .Y (n_7950));
OAI21X1 g60139(.A0 (n_7490), .A1 (n_9489), .B0 (n_7760), .Y (n_7997));
AND2X1 g59839(.A (n_6329), .B (n_7880), .Y (n_7881));
OR2X1 g59840(.A (n_8103), .B (n_7880), .Y (n_8124));
NAND2X1 g59859(.A (n_7876), .B (g6837), .Y (n_8243));
NAND2X1 g59862(.A (n_7876), .B (n_2520), .Y (n_8245));
NAND2X1 g59864(.A (n_7876), .B (n_3914), .Y (n_8247));
NAND2X1 g59870(.A (n_8634), .B (n_1077), .Y (n_9614));
NAND2X1 g59871(.A (n_8634), .B (g6782), .Y (n_9573));
NAND2X1 g59872(.A (n_8634), .B (n_4125), .Y (n_7871));
NAND2X1 g59882(.A (n_7868), .B (n_1301), .Y (n_8273));
NAND2X1 g59883(.A (n_7868), .B (n_2520), .Y (n_8275));
NAND2X1 g59884(.A (n_7868), .B (n_3914), .Y (n_8262));
NAND2X1 g59914(.A (n_998), .B (n_8085), .Y (n_7866));
NAND2X1 g59917(.A (n_7816), .B (n_7517), .Y (n_7865));
INVX2 g59937(.A (n_7791), .Y (n_7932));
AOI22X1 g59942(.A0 (n_973), .A1 (n_7856), .B0 (n_7863), .B1 (n_7892),.Y (n_7864));
AOI22X1 g59943(.A0 (n_1048), .A1 (n_7856), .B0 (n_7861), .B1(n_7892), .Y (n_7862));
AOI22X1 g59944(.A0 (n_1160), .A1 (n_7856), .B0 (n_7858), .B1(n_7892), .Y (n_7860));
AOI22X1 g59945(.A0 (n_1047), .A1 (n_7856), .B0 (n_7855), .B1(n_7892), .Y (n_7857));
AOI22X1 g59946(.A0 (n_1161), .A1 (n_7856), .B0 (n_7853), .B1(n_7892), .Y (n_7854));
AOI22X1 g59947(.A0 (n_1162), .A1 (n_7856), .B0 (n_7851), .B1(n_7892), .Y (n_7852));
INVX1 g59951(.A (n_7848), .Y (n_7849));
NAND3X1 g59692(.A (n_8476), .B (n_7659), .C (n_7722), .Y (n_7847));
AOI22X1 g59704(.A0 (n_7734), .A1 (n_3698), .B0 (n_7457), .B1 (g1243),.Y (n_7846));
CLKBUFX1 gbuf_d_177(.A(n_7709), .Y(d_out_177));
CLKBUFX1 gbuf_qn_177(.A(qn_in_177), .Y(g3106));
CLKBUFX1 gbuf_d_178(.A(n_7713), .Y(d_out_178));
CLKBUFX1 gbuf_qn_178(.A(qn_in_178), .Y(g3107));
CLKBUFX1 gbuf_d_179(.A(n_7711), .Y(d_out_179));
CLKBUFX1 gbuf_qn_179(.A(qn_in_179), .Y(g3108));
MX2X1 g59984(.A (g2261), .B (n_7843), .S0 (n_1301), .Y (n_7845));
MX2X1 g59985(.A (g2264), .B (n_7843), .S0 (g7084), .Y (n_7844));
MX2X1 g59986(.A (g2267), .B (n_7843), .S0 (n_3588), .Y (n_7842));
MX2X1 g59987(.A (g2279), .B (n_7839), .S0 (n_1301), .Y (n_7841));
MX2X1 g59988(.A (g2282), .B (n_7839), .S0 (n_2520), .Y (n_7840));
MX2X1 g59989(.A (g2285), .B (n_7839), .S0 (n_3588), .Y (n_7838));
MX2X1 g59990(.A (g2288), .B (n_7832), .S0 (n_1301), .Y (n_7837));
MX2X1 g59991(.A (g1573), .B (n_7834), .S0 (n_4125), .Y (n_7836));
MX2X1 g59992(.A (g1570), .B (n_7834), .S0 (g6782), .Y (n_7835));
MX2X1 g59993(.A (g2291), .B (n_7832), .S0 (n_2339), .Y (n_7833));
MX2X1 g59994(.A (g2294), .B (n_7832), .S0 (n_3914), .Y (n_7831));
MX2X1 g59995(.A (g1585), .B (n_7828), .S0 (n_1077), .Y (n_7830));
MX2X1 g59998(.A (g1588), .B (n_7828), .S0 (g6782), .Y (n_7829));
MX2X1 g59999(.A (g1594), .B (n_7824), .S0 (g6573), .Y (n_7827));
MX2X1 g60000(.A (g1591), .B (n_7828), .S0 (n_4125), .Y (n_7826));
MX2X1 g60001(.A (g1597), .B (n_7824), .S0 (g6782), .Y (n_7825));
MX2X1 g60002(.A (g1600), .B (n_7824), .S0 (n_4125), .Y (n_7823));
OAI21X1 g59554(.A0 (n_9378), .A1 (n_2343), .B0 (n_2670), .Y (n_7822));
OAI21X1 g59557(.A0 (n_9378), .A1 (n_6420), .B0 (n_5202), .Y (n_7821));
OAI21X1 g59558(.A0 (n_9378), .A1 (n_8305), .B0 (n_1396), .Y (n_7819));
INVX1 g60055(.A (n_7816), .Y (n_7817));
OR2X1 g59852(.A (n_7812), .B (n_1305), .Y (n_9606));
OR2X1 g59853(.A (n_7812), .B (n_7811), .Y (n_9600));
OR2X1 g59854(.A (n_7812), .B (n_7809), .Y (n_9602));
OR2X1 g59855(.A (n_7802), .B (n_1285), .Y (n_7808));
OR2X1 g59856(.A (n_7805), .B (n_1305), .Y (n_7807));
OR2X1 g59857(.A (n_7805), .B (n_7811), .Y (n_7806));
OR2X1 g59858(.A (n_7805), .B (n_7809), .Y (n_9604));
OR2X1 g59860(.A (n_7802), .B (n_2433), .Y (n_9648));
OR2X1 g59861(.A (n_7802), .B (n_7800), .Y (n_7801));
OR2X1 g59867(.A (n_7797), .B (n_1285), .Y (n_9622));
OR2X1 g59868(.A (n_7797), .B (n_2433), .Y (n_9612));
OR2X1 g59869(.A (n_7797), .B (n_7800), .Y (n_9624));
MX2X1 g59903(.A (g1699), .B (n_7793), .S0 (n_1483), .Y (n_7795));
MX2X1 g59904(.A (g1701), .B (n_7793), .S0 (n_6832), .Y (n_7794));
MX2X1 g59905(.A (g1700), .B (n_7793), .S0 (n_3190), .Y (n_7792));
INVX4 g59912(.A (n_7746), .Y (n_7929));
NAND3X1 g59938(.A (n_7724), .B (n_7596), .C (n_8632), .Y (n_7791));
AOI21X1 g59952(.A0 (g1680), .A1 (g1679), .B0 (n_7733), .Y (n_7848));
MX2X1 g59971(.A (g1567), .B (n_7834), .S0 (n_1077), .Y (n_7790));
NAND2X1 g59710(.A (n_4143), .B (n_7680), .Y (n_7789));
NAND2X1 g59711(.A (n_1391), .B (n_7677), .Y (n_7788));
NAND2X1 g59712(.A (n_2445), .B (n_7689), .Y (n_7787));
NAND2X1 g59713(.A (n_4141), .B (n_7673), .Y (n_7786));
CLKBUFX1 gbuf_d_180(.A(n_7703), .Y(d_out_180));
CLKBUFX1 gbuf_q_180(.A(q_in_180), .Y(g927));
CLKBUFX1 gbuf_d_181(.A(n_7700), .Y(d_out_181));
CLKBUFX1 gbuf_q_181(.A(q_in_181), .Y(g930));
CLKBUFX1 gbuf_d_182(.A(n_7702), .Y(d_out_182));
CLKBUFX1 gbuf_q_182(.A(q_in_182), .Y(g933));
CLKBUFX1 gbuf_d_183(.A(n_7656), .Y(d_out_183));
CLKBUFX1 gbuf_q_183(.A(q_in_183), .Y(g873));
CLKBUFX1 gbuf_d_184(.A(n_7653), .Y(d_out_184));
CLKBUFX1 gbuf_q_184(.A(q_in_184), .Y(g879));
CLKBUFX1 gbuf_d_185(.A(n_7655), .Y(d_out_185));
CLKBUFX1 gbuf_q_185(.A(q_in_185), .Y(g876));
CLKBUFX1 gbuf_d_186(.A(n_7652), .Y(d_out_186));
CLKBUFX1 gbuf_q_186(.A(q_in_186), .Y(g891));
CLKBUFX1 gbuf_d_187(.A(n_7650), .Y(d_out_187));
CLKBUFX1 gbuf_q_187(.A(q_in_187), .Y(g894));
CLKBUFX1 gbuf_d_188(.A(n_7708), .Y(d_out_188));
CLKBUFX1 gbuf_q_188(.A(q_in_188), .Y(g897));
CLKBUFX1 gbuf_d_189(.A(n_7707), .Y(d_out_189));
CLKBUFX1 gbuf_q_189(.A(q_in_189), .Y(g900));
CLKBUFX1 gbuf_d_190(.A(n_7706), .Y(d_out_190));
CLKBUFX1 gbuf_q_190(.A(q_in_190), .Y(g903));
CLKBUFX1 gbuf_d_191(.A(n_7704), .Y(d_out_191));
CLKBUFX1 gbuf_q_191(.A(q_in_191), .Y(g906));
CLKBUFX1 gbuf_d_192(.A(n_7682), .Y(d_out_192));
CLKBUFX1 gbuf_q_192(.A(q_in_192), .Y(g312));
CLKBUFX1 gbuf_d_193(.A(n_7679), .Y(d_out_193));
CLKBUFX1 gbuf_q_193(.A(q_in_193), .Y(g313));
CLKBUFX1 gbuf_d_194(.A(n_7674), .Y(d_out_194));
CLKBUFX1 gbuf_q_194(.A(q_in_194), .Y(g_18093));
MX2X1 g60010(.A (g2324), .B (n_9081), .S0 (n_1301), .Y (n_7785));
MX2X1 g60011(.A (g2327), .B (n_9081), .S0 (g7084), .Y (n_7784));
MX2X1 g60012(.A (g2330), .B (n_9081), .S0 (n_3588), .Y (n_7782));
MX2X1 g60013(.A (g1630), .B (n_7779), .S0 (n_1077), .Y (n_7781));
MX2X1 g60014(.A (g1633), .B (n_7779), .S0 (g6782), .Y (n_7780));
MX2X1 g60015(.A (g1636), .B (n_7779), .S0 (n_4125), .Y (n_7778));
INVX1 g60038(.A (n_7645), .Y (n_8085));
NAND2X1 g60056(.A (n_7698), .B (n_5898), .Y (n_7816));
NAND2X2 g59755(.A (n_4163), .B (n_7666), .Y (n_7773));
NAND2X2 g59756(.A (n_1452), .B (n_7671), .Y (n_7772));
NAND2X2 g59757(.A (n_2449), .B (n_7669), .Y (n_7771));
AOI21X1 g60087(.A0 (n_3539), .A1 (n_7732), .B0 (n_7695), .Y (n_7913));
NAND2X1 g60088(.A (n_4279), .B (n_7693), .Y (n_7895));
AOI21X1 g60089(.A0 (n_4896), .A1 (n_7732), .B0 (n_7692), .Y (n_7912));
NAND2X1 g60090(.A (n_4474), .B (n_7691), .Y (n_7893));
OR2X1 g60093(.A (n_8747), .B (n_8868), .Y (n_7769));
OR2X1 g60102(.A (n_5974), .B (n_8868), .Y (n_7768));
NAND3X1 g60117(.A (n_8874), .B (n_9557), .C (n_5380), .Y (n_7764));
XOR2X1 g60146(.A (n_9219), .B (n_7617), .Y (n_7762));
NAND3X1 g60183(.A (n_9489), .B (n_7504), .C (g125), .Y (n_7760));
NAND2X1 g60195(.A (n_7665), .B (n_9195), .Y (n_7759));
NAND2X1 g60196(.A (n_7663), .B (n_9195), .Y (n_7757));
AOI22X1 g60203(.A0 (n_7217), .A1 (n_9483), .B0 (n_8874), .B1 (n_733),.Y (n_7756));
NAND2X1 g59879(.A (n_7753), .B (g6518), .Y (n_8269));
NAND2X1 g59880(.A (n_7753), .B (n_7686), .Y (n_8267));
NAND2X1 g59881(.A (n_7753), .B (n_3919), .Y (n_8271));
NAND2X1 g60275(.A (n_7657), .B (g121), .Y (n_7751));
MX2X1 g59897(.A (g2393), .B (n_7748), .S0 (g5555), .Y (n_7750));
MX2X1 g59898(.A (g2394), .B (n_7748), .S0 (g7264), .Y (n_7749));
MX2X1 g59899(.A (g2395), .B (n_7748), .S0 (n_6611), .Y (n_7747));
AOI21X1 g59909(.A0 (n_7469), .A1 (n_7629), .B0 (n_9141), .Y (n_7876));
NAND2X2 g59913(.A (n_7745), .B (n_6553), .Y (n_7746));
OR2X1 g59916(.A (n_7745), .B (n_970), .Y (n_7880));
INVX2 g59935(.A (n_7714), .Y (n_7868));
MX2X1 g59953(.A (g2333), .B (n_7742), .S0 (g6837), .Y (n_7744));
MX2X1 g59954(.A (g2336), .B (n_7742), .S0 (n_2339), .Y (n_7743));
MX2X1 g59955(.A (g2339), .B (n_7742), .S0 (n_3588), .Y (n_7741));
MX2X1 g59956(.A (g1639), .B (n_7738), .S0 (n_1077), .Y (n_7740));
MX2X1 g59957(.A (g1642), .B (n_7738), .S0 (g6782), .Y (n_7739));
MX2X1 g59958(.A (g1645), .B (n_7738), .S0 (n_4125), .Y (n_7737));
NAND2X1 g59708(.A (n_1399), .B (n_7687), .Y (n_7736));
NAND2X1 g59709(.A (n_2442), .B (n_7685), .Y (n_7735));
CLKBUFX1 gbuf_d_195(.A(n_7614), .Y(d_out_195));
CLKBUFX1 gbuf_q_195(.A(q_in_195), .Y(g1005));
CLKBUFX1 gbuf_d_196(.A(n_7613), .Y(d_out_196));
CLKBUFX1 gbuf_q_196(.A(q_in_196), .Y(g1006));
CLKBUFX1 gbuf_d_197(.A(n_7611), .Y(d_out_197));
CLKBUFX1 gbuf_q_197(.A(q_in_197), .Y(g1007));
CLKBUFX1 gbuf_d_198(.A(n_7646), .Y(d_out_198));
CLKBUFX1 gbuf_q_198(.A(q_in_198), .Y(g942));
CLKBUFX1 gbuf_d_199(.A(n_7648), .Y(d_out_199));
CLKBUFX1 gbuf_q_199(.A(q_in_199), .Y(g939));
CLKBUFX1 gbuf_d_200(.A(n_7649), .Y(d_out_200));
CLKBUFX1 gbuf_q_200(.A(q_in_200), .Y(g936));
CLKBUFX1 gbuf_d_201(.A(n_7639), .Y(d_out_201));
CLKBUFX1 gbuf_q_201(.A(q_in_201), .Y(g16437));
XOR2X1 g60003(.A (n_7556), .B (n_7588), .Y (n_7734));
CLKBUFX1 gbuf_d_202(.A(n_7630), .Y(d_out_202));
CLKBUFX1 gbuf_q_202(.A(q_in_202), .Y(g3053));
CLKBUFX1 gbuf_d_203(.A(n_7636), .Y(d_out_203));
CLKBUFX1 gbuf_q_203(.A(q_in_203), .Y(g3056));
CLKBUFX1 gbuf_d_204(.A(n_7638), .Y(d_out_204));
CLKBUFX1 gbuf_q_204(.A(q_in_204), .Y(g3052));
CLKBUFX1 gbuf_d_205(.A(n_7637), .Y(d_out_205));
CLKBUFX1 gbuf_q_205(.A(q_in_205), .Y(g3055));
CLKBUFX1 gbuf_d_206(.A(n_7632), .Y(d_out_206));
CLKBUFX1 gbuf_q_206(.A(q_in_206), .Y(g3058));
CLKBUFX1 gbuf_d_207(.A(n_7633), .Y(d_out_207));
CLKBUFX1 gbuf_q_207(.A(q_in_207), .Y(g3057));
NOR2X1 g60050(.A (n_7627), .B (g1680), .Y (n_7733));
AOI21X1 g60081(.A0 (n_3545), .A1 (n_7732), .B0 (n_7626), .Y (n_7863));
AOI21X1 g60082(.A0 (n_4038), .A1 (n_7732), .B0 (n_7625), .Y (n_7861));
AOI21X1 g60083(.A0 (n_3543), .A1 (n_7732), .B0 (n_7623), .Y (n_7858));
NOR3X1 g60084(.A (n_4035), .B (n_4071), .C (n_7694), .Y (n_7855));
AOI21X1 g60085(.A0 (n_3541), .A1 (n_7732), .B0 (n_7621), .Y (n_7853));
AOI21X1 g60086(.A0 (n_4039), .A1 (n_7732), .B0 (n_7622), .Y (n_7851));
NAND4X1 g60184(.A (n_7618), .B (n_7992), .C (n_485), .D (n_1205), .Y(n_7730));
NAND2X1 g60286(.A (n_7537), .B (n_7726), .Y (n_9626));
NAND2X1 g60311(.A (n_6734), .B (n_7726), .Y (n_8258));
NAND2X1 g60321(.A (n_7608), .B (n_7511), .Y (n_7724));
NAND2X1 g59921(.A (n_7643), .B (n_5239), .Y (n_7723));
NAND2X1 g59924(.A (n_7641), .B (n_7277), .Y (n_7722));
NAND3X1 g59929(.A (n_9139), .B (n_8191), .C (n_9575), .Y (n_7812));
NAND3X1 g59930(.A (n_9616), .B (n_9617), .C (n_8632), .Y (n_7802));
NAND3X1 g59932(.A (n_7615), .B (n_7599), .C (n_8632), .Y (n_7883));
NAND3X1 g59936(.A (n_7616), .B (n_7601), .C (n_9139), .Y (n_7714));
NAND3X1 g59940(.A (n_9139), .B (n_8189), .C (n_9576), .Y (n_7805));
NAND3X1 g59941(.A (n_9596), .B (n_9597), .C (n_8632), .Y (n_7797));
MX2X1 g59948(.A (n_7712), .B (n_7710), .S0 (g8030), .Y (n_7713));
MX2X1 g59949(.A (n_1198), .B (n_7710), .S0 (g3109), .Y (n_7711));
MX2X1 g59950(.A (n_1171), .B (n_7710), .S0 (g8106), .Y (n_7709));
MX2X1 g59978(.A (g897), .B (n_7651), .S0 (n_3589), .Y (n_7708));
MX2X1 g59979(.A (g900), .B (n_7705), .S0 (n_7675), .Y (n_7707));
MX2X1 g59980(.A (g903), .B (n_7705), .S0 (g6518), .Y (n_7706));
MX2X1 g59981(.A (g906), .B (n_7705), .S0 (n_3919), .Y (n_7704));
OAI21X1 g59714(.A0 (n_7701), .A1 (n_1032), .B0 (n_1312), .Y (n_7703));
CLKBUFX1 gbuf_d_208(.A(n_7710), .Y(d_out_208));
CLKBUFX1 gbuf_q_208(.A(q_in_208), .Y(g2622));
OAI21X1 g59715(.A0 (n_4162), .A1 (n_7701), .B0 (n_4168), .Y (n_7702));
OAI21X1 g59716(.A0 (n_7701), .A1 (n_8339), .B0 (n_2355), .Y (n_7700));
INVX1 g60042(.A (n_7645), .Y (n_7745));
AND2X1 g60051(.A (n_7589), .B (n_8476), .Y (n_7793));
NAND2X1 g60078(.A (n_7575), .B (n_7371), .Y (n_7698));
AOI21X1 g60123(.A0 (n_6459), .A1 (n_7696), .B0 (n_7582), .Y (n_7834));
AOI21X1 g60126(.A0 (n_6215), .A1 (n_7697), .B0 (n_7583), .Y (n_7843));
AOI21X1 g60127(.A0 (n_7164), .A1 (n_7697), .B0 (n_7581), .Y (n_7839));
AOI21X1 g60128(.A0 (n_7363), .A1 (n_7697), .B0 (n_7579), .Y (n_7832));
AOI21X1 g60129(.A0 (n_7249), .A1 (n_7696), .B0 (n_7578), .Y (n_7828));
CLKBUFX1 gbuf_d_209(.A(n_7571), .Y(d_out_209));
CLKBUFX1 gbuf_q_209(.A(q_in_209), .Y(g3051));
AOI21X1 g60130(.A0 (n_7435), .A1 (n_7696), .B0 (n_7576), .Y (n_7824));
OR2X1 g60140(.A (n_7586), .B (n_7992), .Y (n_8007));
OR2X1 g60162(.A (n_4318), .B (n_7694), .Y (n_7695));
NOR2X1 g60163(.A (n_4067), .B (n_7694), .Y (n_7693));
OR2X1 g60164(.A (n_4507), .B (n_7694), .Y (n_7692));
NOR2X1 g60165(.A (n_4065), .B (n_7694), .Y (n_7691));
NAND2X1 g59841(.A (n_7676), .B (g6518), .Y (n_7689));
NAND2X1 g59847(.A (n_7684), .B (n_7686), .Y (n_7687));
NAND2X1 g59848(.A (n_7684), .B (g6518), .Y (n_7685));
MX2X1 g60205(.A (g312), .B (n_7678), .S0 (n_6914), .Y (n_7682));
NAND2X1 g59849(.A (n_7684), .B (n_3589), .Y (n_7680));
MX2X1 g60206(.A (g313), .B (n_7678), .S0 (g6447), .Y (n_7679));
NAND2X1 g59850(.A (n_7676), .B (n_7675), .Y (n_7677));
MX2X1 g60207(.A (g_18093), .B (n_7678), .S0 (n_6917), .Y (n_7674));
NAND2X1 g59851(.A (n_7676), .B (n_3919), .Y (n_7673));
NAND2X1 g59873(.A (n_7668), .B (g6368), .Y (n_7671));
NAND2X1 g59874(.A (n_7668), .B (g6518), .Y (n_7669));
NAND2X1 g59878(.A (n_7668), .B (n_3919), .Y (n_7666));
NAND2X1 g60257(.A (n_9562), .B (n_5382), .Y (n_7665));
NAND2X1 g60274(.A (n_9562), .B (n_5247), .Y (n_7663));
NAND2X1 g59920(.A (n_7642), .B (n_7347), .Y (n_7660));
NAND2X1 g59923(.A (n_7640), .B (n_7345), .Y (n_7659));
INVX1 g60380(.A (n_9483), .Y (n_7657));
INVX2 g59933(.A (n_7609), .Y (n_7753));
MX2X1 g59969(.A (g873), .B (n_7654), .S0 (n_7675), .Y (n_7656));
MX2X1 g59972(.A (g876), .B (n_7654), .S0 (g6518), .Y (n_7655));
MX2X1 g59973(.A (g879), .B (n_7654), .S0 (n_3589), .Y (n_7653));
MX2X1 g59976(.A (g891), .B (n_7651), .S0 (n_7675), .Y (n_7652));
MX2X1 g59977(.A (g894), .B (n_7651), .S0 (g6518), .Y (n_7650));
CLKBUFX1 gbuf_d_210(.A(n_7564), .Y(d_out_210));
CLKBUFX1 gbuf_q_210(.A(q_in_210), .Y(g945));
CLKBUFX1 gbuf_d_211(.A(n_7562), .Y(d_out_211));
CLKBUFX1 gbuf_q_211(.A(q_in_211), .Y(g948));
CLKBUFX1 gbuf_d_212(.A(n_7565), .Y(d_out_212));
CLKBUFX1 gbuf_q_212(.A(q_in_212), .Y(g951));
MX2X1 g60005(.A (g936), .B (n_7647), .S0 (n_7675), .Y (n_7649));
MX2X1 g60006(.A (g939), .B (n_7647), .S0 (g6518), .Y (n_7648));
MX2X1 g60007(.A (g942), .B (n_7647), .S0 (n_3589), .Y (n_7646));
CLKBUFX1 gbuf_d_213(.A(n_7559), .Y(d_out_213));
CLKBUFX1 gbuf_q_213(.A(q_in_213), .Y(g3060));
CLKBUFX1 gbuf_d_214(.A(n_7560), .Y(d_out_214));
CLKBUFX1 gbuf_q_214(.A(q_in_214), .Y(g3059));
NAND2X1 g60043(.A (n_5937), .B (n_7590), .Y (n_7645));
AND2X1 g60048(.A (n_8542), .B (n_9644), .Y (n_7748));
INVX1 g60059(.A (n_7642), .Y (n_7643));
INVX1 g60061(.A (n_7640), .Y (n_7641));
OAI21X1 g60063(.A0 (n_7530), .A1 (g2580), .B0 (n_6645), .Y (n_7639));
OAI21X1 g60105(.A0 (n_7508), .A1 (n_896), .B0 (n_7634), .Y (n_7638));
INVX1 g60106(.A (n_7594), .Y (n_7637));
OAI21X1 g60108(.A0 (n_7507), .A1 (n_896), .B0 (n_7634), .Y (n_7636));
OAI21X1 g60109(.A0 (n_7506), .A1 (n_896), .B0 (n_7631), .Y (n_7633));
OAI21X1 g60110(.A0 (n_7505), .A1 (n_896), .B0 (n_7631), .Y (n_7632));
INVX1 g60111(.A (n_7593), .Y (n_7630));
AOI21X1 g60113(.A0 (n_6422), .A1 (n_7587), .B0 (n_7992), .Y (n_7957));
NOR2X1 g60119(.A (n_7550), .B (n_7546), .Y (n_7779));
NAND2X1 g60132(.A (n_7555), .B (n_7403), .Y (n_7629));
OAI21X1 g60136(.A0 (n_7397), .A1 (n_7403), .B0 (n_7553), .Y (n_7742));
OAI21X1 g60137(.A0 (n_7491), .A1 (n_7448), .B0 (n_7552), .Y (n_7738));
AOI22X1 g60141(.A0 (n_7607), .A1 (g7014), .B0 (g1686), .B1 (n_3036),.Y (n_7627));
NAND2X1 g60157(.A (n_4324), .B (n_7624), .Y (n_7626));
NAND2X1 g60158(.A (n_4323), .B (n_7624), .Y (n_7625));
NAND2X1 g60159(.A (n_4322), .B (n_7624), .Y (n_7623));
NAND2X1 g60161(.A (n_4320), .B (n_7624), .Y (n_7622));
NAND2X1 g60160(.A (n_4321), .B (n_7624), .Y (n_7621));
AOI21X1 g60193(.A0 (n_7519), .A1 (g1916), .B0 (n_7892), .Y (n_7620));
AOI21X1 g60194(.A0 (n_7519), .A1 (g1917), .B0 (n_7892), .Y (n_7619));
NOR2X1 g60268(.A (n_7380), .B (n_7892), .Y (n_7618));
NAND2X1 g60272(.A (n_7540), .B (n_7499), .Y (n_7617));
NAND2X1 g60313(.A (n_7539), .B (n_9077), .Y (n_7616));
NAND2X1 g60315(.A (n_7568), .B (n_7696), .Y (n_7615));
MX2X1 g59900(.A (g1005), .B (n_7612), .S0 (g5472), .Y (n_7614));
MX2X1 g59901(.A (g1006), .B (n_7612), .S0 (g6712), .Y (n_7613));
MX2X1 g59902(.A (n_7612), .B (g1007), .S0 (n_6420), .Y (n_7611));
INVX2 g60371(.A (n_9562), .Y (n_7726));
NAND3X1 g59934(.A (n_7548), .B (n_7433), .C (n_7566), .Y (n_7609));
MX2X1 g60475(.A (n_4444), .B (n_5947), .S0 (n_7536), .Y (n_7608));
INVX1 g59982(.A (n_7567), .Y (n_7676));
CLKBUFX1 gbuf_d_215(.A(n_7529), .Y(d_out_215));
CLKBUFX1 gbuf_q_215(.A(q_in_215), .Y(g2387));
CLKBUFX1 gbuf_d_216(.A(n_7528), .Y(d_out_216));
CLKBUFX1 gbuf_q_216(.A(q_in_216), .Y(g2388));
CLKBUFX1 gbuf_d_217(.A(n_7526), .Y(d_out_217));
CLKBUFX1 gbuf_q_217(.A(q_in_217), .Y(g2389));
CLKBUFX1 gbuf_d_218(.A(n_7521), .Y(d_out_218));
CLKBUFX1 gbuf_q_218(.A(q_in_218), .Y(g1695));
CLKBUFX1 gbuf_d_219(.A(n_7524), .Y(d_out_219));
CLKBUFX1 gbuf_q_219(.A(q_in_219), .Y(g1694));
CLKBUFX1 gbuf_d_220(.A(n_7607), .Y(d_out_220));
CLKBUFX1 gbuf_q_220(.A(q_in_220), .Y(g992));
NAND2X1 g60060(.A (n_7532), .B (n_9347), .Y (n_7642));
NAND2X1 g60062(.A (n_7531), .B (n_6969), .Y (n_7640));
NAND3X1 g60094(.A (n_7403), .B (n_9147), .C (n_436), .Y (n_9575));
NAND2X1 g60095(.A (n_4534), .B (n_7600), .Y (n_7605));
NAND3X1 g60096(.A (n_7407), .B (n_8635), .C (n_435), .Y (n_9616));
NAND3X1 g60097(.A (n_7403), .B (n_9144), .C (n_8759), .Y (n_9576));
NAND2X1 g60098(.A (n_4780), .B (n_7600), .Y (n_7601));
NAND2X1 g60099(.A (n_5189), .B (n_7595), .Y (n_7599));
NAND3X1 g60100(.A (n_7407), .B (n_8635), .C (n_364), .Y (n_9596));
NAND2X1 g60101(.A (n_4976), .B (n_7595), .Y (n_7596));
AOI21X1 g60107(.A0 (n_7464), .A1 (n_882), .B0 (n_7591), .Y (n_7594));
AOI21X1 g60112(.A0 (n_7465), .A1 (n_882), .B0 (n_7591), .Y (n_7593));
INVX1 g60142(.A (n_7590), .Y (n_7710));
XOR2X1 g60150(.A (n_7187), .B (n_7470), .Y (n_7589));
XOR2X1 g60151(.A (n_7452), .B (n_7454), .Y (n_7588));
OR2X1 g60169(.A (n_7992), .B (n_7587), .Y (n_8004));
AND2X1 g60168(.A (n_6441), .B (n_7587), .Y (n_7586));
NAND2X1 g60185(.A (n_7482), .B (n_9075), .Y (n_7583));
NAND2X1 g60186(.A (n_7478), .B (n_7577), .Y (n_7582));
NAND2X1 g60187(.A (n_7476), .B (n_9075), .Y (n_7581));
NAND2X1 g60188(.A (n_7475), .B (n_9075), .Y (n_7579));
NAND2X1 g60189(.A (n_7472), .B (n_7577), .Y (n_7578));
NAND2X1 g60191(.A (n_7471), .B (n_7577), .Y (n_7576));
NAND2X1 g60221(.A (n_7518), .B (n_7441), .Y (n_7575));
NAND2X2 g59915(.A (n_7533), .B (n_7047), .Y (n_7571));
INVX1 g59925(.A (n_7543), .Y (n_7668));
CLKBUFX1 gbuf_d_221(.A(n_7525), .Y(d_out_221));
CLKBUFX1 gbuf_q_221(.A(q_in_221), .Y(g1693));
MX2X1 g60476(.A (n_5233), .B (n_5051), .S0 (n_7493), .Y (n_7569));
INVX1 g59974(.A (n_7538), .Y (n_7684));
XOR2X1 g60539(.A (n_4676), .B (n_8462), .Y (n_7568));
NAND3X1 g59983(.A (n_7566), .B (n_7389), .C (n_9608), .Y (n_7567));
CLKBUFX1 gbuf_d_222(.A(n_7460), .Y(d_out_222));
CLKBUFX1 gbuf_qn_222(.A(qn_in_222), .Y(g3103));
CLKBUFX1 gbuf_d_223(.A(n_7461), .Y(d_out_223));
CLKBUFX1 gbuf_qn_223(.A(qn_in_223), .Y(g3104));
CLKBUFX1 gbuf_d_224(.A(n_7445), .Y(d_out_224));
CLKBUFX1 gbuf_q_224(.A(q_in_224), .Y(g_16936));
CLKBUFX1 gbuf_d_225(.A(n_7444), .Y(d_out_225));
CLKBUFX1 gbuf_q_225(.A(q_in_225), .Y(g322));
CLKBUFX1 gbuf_d_226(.A(n_7442), .Y(d_out_226));
CLKBUFX1 gbuf_q_226(.A(q_in_226), .Y(g_8008));
MX2X1 g60004(.A (g951), .B (n_7563), .S0 (n_3589), .Y (n_7565));
MX2X1 g60008(.A (g945), .B (n_7563), .S0 (n_7675), .Y (n_7564));
MX2X1 g60009(.A (g948), .B (n_7563), .S0 (g6518), .Y (n_7562));
AOI21X1 g60122(.A0 (n_6065), .A1 (n_7561), .B0 (n_7486), .Y (n_7654));
AOI21X1 g60124(.A0 (n_6978), .A1 (n_7561), .B0 (n_7485), .Y (n_7651));
AOI21X1 g60135(.A0 (n_7251), .A1 (n_7561), .B0 (n_7483), .Y (n_7705));
AOI22X1 g60143(.A0 (n_7420), .A1 (n_5749), .B0 (g2618), .B1 (g2574),.Y (n_7590));
OAI22X1 g60144(.A0 (n_7422), .A1 (n_896), .B0 (n_7456), .B1 (n_7558),.Y (n_7560));
OAI22X1 g60145(.A0 (n_7421), .A1 (n_896), .B0 (n_7455), .B1 (n_7558),.Y (n_7559));
XOR2X1 g60148(.A (n_9021), .B (n_7423), .Y (n_9644));
XOR2X1 g60152(.A (n_7416), .B (n_7419), .Y (n_7556));
NAND2X1 g60166(.A (n_9147), .B (n_2719), .Y (n_7555));
NAND2X1 g60167(.A (n_7474), .B (n_454), .Y (n_7554));
NAND2X2 g60178(.A (n_9144), .B (n_9074), .Y (n_9139));
NAND3X1 g60190(.A (n_7403), .B (n_7344), .C (n_482), .Y (n_7553));
NAND3X1 g60192(.A (n_7448), .B (n_7343), .C (n_473), .Y (n_7552));
AOI22X1 g60218(.A0 (n_7252), .A1 (n_7466), .B0 (n_7406), .B1 (n_471),.Y (n_7550));
INVX2 g60265(.A (n_7694), .Y (n_7624));
CLKBUFX1 gbuf_d_227(.A(n_7458), .Y(d_out_227));
CLKBUFX1 gbuf_qn_227(.A(qn_in_227), .Y(g3105));
NAND3X1 g60285(.A (n_7561), .B (n_7439), .C (n_7399), .Y (n_7548));
INVX1 g60299(.A (n_7577), .Y (n_7546));
NAND2X1 g60305(.A (n_7496), .B (n_7697), .Y (n_7545));
NAND2X1 g59908(.A (n_7489), .B (n_7566), .Y (n_7701));
NAND3X1 g59926(.A (n_8253), .B (n_8254), .C (n_7566), .Y (n_7543));
AND2X1 g60404(.A (n_7495), .B (n_7891), .Y (n_7678));
AOI22X1 g60455(.A0 (n_5486), .A1 (n_7498), .B0 (n_5485), .B1(n_9219), .Y (n_7540));
MX2X1 g60474(.A (n_3991), .B (n_5779), .S0 (n_7438), .Y (n_7539));
NAND3X1 g59975(.A (n_7566), .B (n_7392), .C (n_9598), .Y (n_7538));
MX2X1 g60537(.A (n_5232), .B (n_6697), .S0 (n_7492), .Y (n_7537));
NAND2X1 g60582(.A (n_8462), .B (n_6841), .Y (n_7536));
AND2X1 g60049(.A (n_7431), .B (n_9375), .Y (n_7612));
AOI22X1 g60064(.A0 (n_7386), .A1 (n_3701), .B0 (n_7223), .B1 (g557),.Y (n_7533));
NAND2X1 g60079(.A (n_7429), .B (n_7194), .Y (n_7532));
NAND2X1 g60080(.A (n_7430), .B (n_5477), .Y (n_7531));
NOR2X1 g60103(.A (n_7387), .B (n_7426), .Y (n_7647));
NOR2X1 g60179(.A (n_9077), .B (n_9148), .Y (n_7600));
NOR2X1 g60182(.A (n_7477), .B (n_8636), .Y (n_7595));
AOI22X1 g60201(.A0 (n_7494), .A1 (g7390), .B0 (g16437), .B1 (n_1596),.Y (n_7530));
MX2X1 g60211(.A (g2387), .B (n_7527), .S0 (g5555), .Y (n_7529));
MX2X1 g60212(.A (g2388), .B (n_7527), .S0 (g7264), .Y (n_7528));
MX2X1 g60213(.A (g2389), .B (n_7527), .S0 (n_6611), .Y (n_7526));
MX2X1 g60214(.A (g1693), .B (n_7523), .S0 (g5511), .Y (n_7525));
MX2X1 g60215(.A (g1694), .B (n_7523), .S0 (n_3190), .Y (n_7524));
MX2X1 g60216(.A (g1695), .B (n_7523), .S0 (n_6832), .Y (n_7521));
NAND2X2 g60266(.A (n_7519), .B (n_6461), .Y (n_7694));
OR2X1 g60267(.A (n_7519), .B (n_6440), .Y (n_7587));
NAND3X1 g60271(.A (n_7517), .B (n_7376), .C (n_7258), .Y (n_7518));
NAND2X1 g60292(.A (n_6824), .B (n_9077), .Y (n_8191));
INVX1 g60300(.A (n_8630), .Y (n_7577));
NAND2X1 g60304(.A (n_6967), .B (n_7511), .Y (n_9617));
NAND2X1 g60310(.A (n_6658), .B (n_9077), .Y (n_8189));
NAND2X1 g60318(.A (n_6795), .B (n_7511), .Y (n_9597));
NAND2X1 g60330(.A (n_7415), .B (n_7264), .Y (n_7508));
NAND2X1 g60333(.A (n_7413), .B (n_7263), .Y (n_7507));
NAND2X1 g60334(.A (n_7411), .B (n_7262), .Y (n_7506));
NAND2X1 g60335(.A (n_7410), .B (n_7261), .Y (n_7505));
OAI21X1 g60339(.A0 (n_7375), .A1 (g986), .B0 (n_7003), .Y (n_7607));
INVX1 g60360(.A (n_8876), .Y (n_7504));
INVX1 g60387(.A (n_7380), .Y (n_7856));
NAND4X1 g60430(.A (n_7498), .B (n_5337), .C (n_9219), .D (n_7209), .Y(n_7499));
XOR2X1 g60538(.A (n_4678), .B (n_8395), .Y (n_7496));
XOR2X1 g60540(.A (n_5485), .B (n_7372), .Y (n_7495));
CLKBUFX1 gbuf_d_228(.A(n_7494), .Y(d_out_228));
CLKBUFX1 gbuf_q_228(.A(q_in_228), .Y(g16399));
NAND2X1 g60583(.A (n_7492), .B (n_6772), .Y (n_7493));
XOR2X1 g60619(.A (n_4596), .B (n_8463), .Y (n_7491));
AOI21X1 g60620(.A0 (n_5463), .A1 (n_8483), .B0 (n_7395), .Y (n_7490));
OR2X1 g60052(.A (n_7295), .B (n_7388), .Y (n_7489));
INVX1 g60057(.A (n_9379), .Y (n_7488));
NAND2X1 g60198(.A (n_7353), .B (n_7484), .Y (n_7486));
NAND2X1 g60199(.A (n_7351), .B (n_7484), .Y (n_7485));
NAND2X1 g60200(.A (n_7349), .B (n_7484), .Y (n_7483));
OR2X1 g60291(.A (n_9077), .B (g2165), .Y (n_7482));
OR2X1 g60297(.A (n_7477), .B (g1471), .Y (n_7478));
OR2X1 g60298(.A (n_9077), .B (g2185), .Y (n_7476));
OR2X1 g60303(.A (n_9077), .B (g2195), .Y (n_7475));
INVX1 g60306(.A (n_8636), .Y (n_7474));
OR2X1 g60312(.A (n_7477), .B (n_600), .Y (n_7472));
OR2X1 g60314(.A (n_7477), .B (g1501), .Y (n_7471));
NAND2X1 g60323(.A (n_7377), .B (n_7342), .Y (n_7470));
NAND2X1 g60326(.A (n_6926), .B (n_9077), .Y (n_7469));
AOI22X1 g60331(.A0 (n_1257), .A1 (n_7463), .B0 (n_7451), .B1(n_7462), .Y (n_7465));
AOI22X1 g60332(.A0 (n_1443), .A1 (n_7463), .B0 (n_7453), .B1(n_7462), .Y (n_7464));
MX2X1 g60336(.A (n_1197), .B (n_7459), .S0 (g8030), .Y (n_7461));
MX2X1 g60337(.A (n_911), .B (n_7459), .S0 (g8106), .Y (n_7460));
MX2X1 g60338(.A (n_1170), .B (n_7459), .S0 (g3109), .Y (n_7458));
XOR2X1 g60341(.A (n_7456), .B (n_7455), .Y (n_7457));
XOR2X1 g60342(.A (n_7412), .B (n_7453), .Y (n_7454));
XOR2X1 g60343(.A (n_7414), .B (n_7451), .Y (n_7452));
INVX1 g60399(.A (n_7511), .Y (n_7448));
MX2X1 g60462(.A (g_16936), .B (n_7443), .S0 (n_7362), .Y (n_7445));
MX2X1 g60463(.A (g322), .B (n_7443), .S0 (n_7361), .Y (n_7444));
MX2X1 g60464(.A (g_8008), .B (n_7443), .S0 (n_7359), .Y (n_7442));
CLKBUFX1 gbuf_d_229(.A(n_7366), .Y(d_out_229));
CLKBUFX1 gbuf_qn_229(.A(qn_in_229), .Y(g_18564));
CLKBUFX1 gbuf_d_230(.A(n_7459), .Y(d_out_230));
CLKBUFX1 gbuf_q_230(.A(q_in_230), .Y(g1928));
NAND2X1 g60560(.A (n_9224), .B (n_5099), .Y (n_7498));
NAND2X1 g60564(.A (n_7365), .B (n_5099), .Y (n_7441));
NAND2X1 g60579(.A (n_7370), .B (n_4001), .Y (n_7439));
NAND2X1 g60581(.A (n_8394), .B (n_6700), .Y (n_7438));
AOI21X1 g60714(.A0 (n_6603), .A1 (n_8464), .B0 (n_7358), .Y (n_7435));
OR2X1 g60091(.A (n_4280), .B (n_7432), .Y (n_8253));
OR2X1 g60092(.A (n_4281), .B (n_7432), .Y (n_7433));
OAI21X1 g60138(.A0 (n_7315), .A1 (n_7246), .B0 (n_7354), .Y (n_7563));
XOR2X1 g60149(.A (n_7155), .B (n_7296), .Y (n_7431));
NAND2X2 g60173(.A (n_7385), .B (n_9309), .Y (n_7566));
NAND2X1 g60219(.A (n_7346), .B (n_7278), .Y (n_7430));
NAND2X1 g60220(.A (n_7348), .B (n_7232), .Y (n_7429));
CLKBUFX1 gbuf_d_231(.A(n_7339), .Y(d_out_231));
CLKBUFX1 gbuf_q_231(.A(q_in_231), .Y(g3044));
CLKBUFX1 gbuf_d_232(.A(n_7338), .Y(d_out_232));
CLKBUFX1 gbuf_q_232(.A(q_in_232), .Y(g3045));
CLKBUFX1 gbuf_d_233(.A(n_7331), .Y(d_out_233));
CLKBUFX1 gbuf_q_233(.A(q_in_233), .Y(g3048));
CLKBUFX1 gbuf_d_234(.A(n_7332), .Y(d_out_234));
CLKBUFX1 gbuf_q_234(.A(q_in_234), .Y(g3047));
CLKBUFX1 gbuf_d_235(.A(n_7335), .Y(d_out_235));
CLKBUFX1 gbuf_q_235(.A(q_in_235), .Y(g3043));
CLKBUFX1 gbuf_d_236(.A(n_7334), .Y(d_out_236));
CLKBUFX1 gbuf_q_236(.A(q_in_236), .Y(g3046));
NAND2X1 g60273(.A (n_7373), .B (n_7561), .Y (n_8254));
INVX1 g60277(.A (n_7484), .Y (n_7426));
NAND2X1 g60319(.A (n_7329), .B (n_7292), .Y (n_7423));
AOI21X1 g60324(.A0 (n_7417), .A1 (n_7462), .B0 (n_7319), .Y (n_7422));
AOI21X1 g60325(.A0 (n_7418), .A1 (n_7462), .B0 (n_7318), .Y (n_7421));
OAI21X1 g60340(.A0 (n_7280), .A1 (n_6822), .B0 (n_632), .Y (n_7420));
XOR2X1 g60344(.A (n_7418), .B (n_7417), .Y (n_7419));
XOR2X1 g60345(.A (n_7324), .B (n_7326), .Y (n_7416));
NAND2X1 g60359(.A (n_7414), .B (n_7462), .Y (n_7415));
NAND2X1 g60362(.A (n_7412), .B (n_7462), .Y (n_7413));
NAND2X1 g60363(.A (n_7327), .B (n_7462), .Y (n_7411));
NAND2X1 g60364(.A (n_7325), .B (n_7462), .Y (n_7410));
INVX2 g60391(.A (n_7380), .Y (n_7519));
INVX2 g60395(.A (n_7466), .Y (n_7407));
CLKBUFX3 g60396(.A (n_7466), .Y (n_7696));
CLKBUFX3 g60400(.A (n_7477), .Y (n_7511));
INVX1 g60401(.A (n_7477), .Y (n_7406));
INVX4 g60418(.A (n_9077), .Y (n_7403));
CLKBUFX1 g60419(.A (n_9077), .Y (n_7697));
CLKBUFX1 gbuf_d_237(.A(n_7308), .Y(d_out_237));
CLKBUFX1 gbuf_qn_237(.A(qn_in_237), .Y(g_27975));
CLKBUFX1 gbuf_d_238(.A(n_7301), .Y(d_out_238));
CLKBUFX1 gbuf_q_238(.A(q_in_238), .Y(g1000));
CLKBUFX1 gbuf_d_239(.A(n_7306), .Y(d_out_239));
CLKBUFX1 gbuf_q_239(.A(q_in_239), .Y(g999));
CLKBUFX1 gbuf_d_240(.A(n_7289), .Y(d_out_240));
CLKBUFX1 gbuf_q_240(.A(q_in_240), .Y(g2396));
CLKBUFX1 gbuf_d_241(.A(n_7288), .Y(d_out_241));
CLKBUFX1 gbuf_q_241(.A(q_in_241), .Y(g2397));
CLKBUFX1 gbuf_d_242(.A(n_7286), .Y(d_out_242));
CLKBUFX1 gbuf_q_242(.A(q_in_242), .Y(g2398));
CLKBUFX1 gbuf_d_243(.A(n_7285), .Y(d_out_243));
CLKBUFX1 gbuf_q_243(.A(q_in_243), .Y(g1702));
CLKBUFX1 gbuf_d_244(.A(n_7284), .Y(d_out_244));
CLKBUFX1 gbuf_q_244(.A(q_in_244), .Y(g1703));
CLKBUFX1 gbuf_d_245(.A(n_7282), .Y(d_out_245));
CLKBUFX1 gbuf_q_245(.A(q_in_245), .Y(g1704));
CLKBUFX1 gbuf_d_246(.A(n_7311), .Y(d_out_246));
CLKBUFX1 gbuf_q_246(.A(q_in_246), .Y(g402));
CLKBUFX1 gbuf_d_247(.A(n_7312), .Y(d_out_247));
CLKBUFX1 gbuf_q_247(.A(q_in_247), .Y(g403));
CLKBUFX1 gbuf_d_248(.A(n_7309), .Y(d_out_248));
CLKBUFX1 gbuf_q_248(.A(q_in_248), .Y(g404));
NAND2X1 g60580(.A (n_7369), .B (n_8884), .Y (n_7399));
NAND4X1 g60584(.A (n_7317), .B (n_882), .C (n_461), .D (n_1367), .Y(n_7398));
XOR2X1 g60618(.A (n_4206), .B (n_8397), .Y (n_7397));
NOR2X1 g60673(.A (n_6619), .B (n_8483), .Y (n_7492));
NOR2X1 g60678(.A (n_5463), .B (n_8483), .Y (n_7395));
NAND3X1 g60115(.A (n_7246), .B (n_9309), .C (n_3171), .Y (n_7392));
NAND3X1 g60116(.A (n_7246), .B (n_9309), .C (n_4110), .Y (n_7389));
AOI21X1 g60125(.A0 (n_9309), .A1 (n_525), .B0 (n_7247), .Y (n_7388));
AOI22X1 g60202(.A0 (n_7046), .A1 (n_7561), .B0 (n_7355), .B1 (g805),.Y (n_7387));
XOR2X1 g60204(.A (n_7239), .B (n_7238), .Y (n_7386));
CLKBUFX1 gbuf_d_249(.A(n_7304), .Y(d_out_249));
CLKBUFX1 gbuf_q_249(.A(q_in_249), .Y(g1001));
INVX2 g60278(.A (n_7385), .Y (n_7484));
NAND2X2 g60296(.A (n_9627), .B (n_8541), .Y (n_7384));
NAND2X2 g60392(.A (n_5936), .B (n_7322), .Y (n_7380));
INVX1 g60397(.A (n_7379), .Y (n_7466));
INVX2 g60402(.A (n_7379), .Y (n_7477));
AND2X1 g60428(.A (n_7321), .B (n_8542), .Y (n_7527));
AND2X1 g60429(.A (n_7320), .B (n_8476), .Y (n_7523));
OAI21X1 g60441(.A0 (n_7266), .A1 (g1886), .B0 (n_6571), .Y (n_7494));
AOI22X1 g60458(.A0 (n_7341), .A1 (n_9591), .B0 (n_5064), .B1(n_7187), .Y (n_7377));
NAND3X1 g60512(.A (n_6985), .B (n_7260), .C (n_7082), .Y (n_7376));
AOI22X1 g60531(.A0 (n_7374), .A1 (g6712), .B0 (g992), .B1 (n_2361),.Y (n_7375));
CLKBUFX1 gbuf_d_250(.A(n_7374), .Y(d_out_250));
CLKBUFX1 gbuf_q_250(.A(q_in_250), .Y(g_20059));
AOI21X1 g60585(.A0 (n_7218), .A1 (n_7371), .B0 (n_7214), .Y (n_7443));
MX2X1 g60612(.A (n_3985), .B (n_4223), .S0 (n_7316), .Y (n_7373));
AOI21X1 g60658(.A0 (n_7213), .A1 (n_7371), .B0 (n_8863), .Y (n_7372));
INVX1 g60671(.A (n_7369), .Y (n_7370));
NOR2X1 g60047(.A (n_7307), .B (n_9611), .Y (n_7366));
AOI22X1 g60691(.A0 (n_7212), .A1 (n_9219), .B0 (n_8678), .B1(n_7257), .Y (n_7365));
AOI21X1 g60713(.A0 (n_6414), .A1 (n_8398), .B0 (n_7256), .Y (n_7363));
AND2X1 g60785(.A (n_7360), .B (n_6917), .Y (n_7362));
AND2X1 g60787(.A (n_7360), .B (n_6914), .Y (n_7361));
AND2X1 g60788(.A (n_7360), .B (g6447), .Y (n_7359));
NOR2X1 g60795(.A (n_6603), .B (n_8464), .Y (n_7358));
NAND2X1 g60174(.A (n_9309), .B (n_7355), .Y (n_7432));
NAND3X1 g60175(.A (n_7246), .B (n_7204), .C (n_763), .Y (n_7354));
CLKBUFX1 gbuf_d_251(.A(n_7241), .Y(d_out_251));
CLKBUFX1 gbuf_q_251(.A(q_in_251), .Y(g3050));
CLKBUFX1 gbuf_d_252(.A(n_7242), .Y(d_out_252));
CLKBUFX1 gbuf_q_252(.A(q_in_252), .Y(g3049));
NAND2X1 g60276(.A (n_7246), .B (n_590), .Y (n_7353));
INVX2 g60279(.A (n_7297), .Y (n_7385));
NAND2X1 g60281(.A (n_6735), .B (n_7561), .Y (n_9598));
NAND2X1 g60283(.A (n_7246), .B (n_448), .Y (n_7351));
NAND2X1 g60284(.A (n_6483), .B (n_7561), .Y (n_9608));
NAND2X1 g60316(.A (n_7246), .B (n_762), .Y (n_7349));
NAND3X1 g60317(.A (n_7347), .B (n_7198), .C (n_7049), .Y (n_7348));
NAND3X1 g60322(.A (n_7345), .B (n_7197), .C (n_7048), .Y (n_7346));
INVX1 g60367(.A (n_8541), .Y (n_7344));
INVX1 g60369(.A (n_7381), .Y (n_7343));
NAND2X2 g60403(.A (n_7235), .B (n_7293), .Y (n_7379));
NAND4X1 g60433(.A (n_7341), .B (n_5477), .C (n_7187), .D (n_6988), .Y(n_7342));
OAI21X1 g60434(.A0 (n_7229), .A1 (n_7337), .B0 (n_7336), .Y (n_7339));
OAI21X1 g60435(.A0 (n_7227), .A1 (n_7337), .B0 (n_7336), .Y (n_7338));
OAI21X1 g60437(.A0 (n_7230), .A1 (n_7337), .B0 (n_7333), .Y (n_7335));
OAI21X1 g60438(.A0 (n_7226), .A1 (n_7337), .B0 (n_7333), .Y (n_7334));
OAI21X1 g60439(.A0 (n_7225), .A1 (n_7337), .B0 (n_7330), .Y (n_7332));
OAI21X1 g60440(.A0 (n_7224), .A1 (n_7337), .B0 (n_7330), .Y (n_7331));
AOI22X1 g60456(.A0 (n_5481), .A1 (n_7291), .B0 (n_5480), .B1(n_9021), .Y (n_7329));
AOI21X1 g60500(.A0 (n_3115), .A1 (n_7328), .B0 (n_7276), .Y (n_7414));
AOI21X1 g60501(.A0 (n_3275), .A1 (n_7328), .B0 (n_7275), .Y (n_7451));
AOI21X1 g60502(.A0 (n_3113), .A1 (n_7328), .B0 (n_7274), .Y (n_7453));
AOI21X1 g60503(.A0 (n_3276), .A1 (n_7328), .B0 (n_7272), .Y (n_7412));
INVX1 g60504(.A (n_7326), .Y (n_7327));
INVX1 g60506(.A (n_7324), .Y (n_7325));
AOI21X1 g60508(.A0 (n_3111), .A1 (n_7328), .B0 (n_7270), .Y (n_7456));
AOI21X1 g60510(.A0 (n_3537), .A1 (n_7328), .B0 (n_7269), .Y (n_7455));
NAND2X1 g60519(.A (n_7268), .B (n_896), .Y (n_7634));
INVX1 g60520(.A (n_7322), .Y (n_7459));
XOR2X1 g60541(.A (n_5480), .B (n_7195), .Y (n_7321));
XOR2X1 g60543(.A (n_5064), .B (n_7193), .Y (n_7320));
CLKBUFX1 gbuf_d_253(.A(n_7201), .Y(d_out_253));
CLKBUFX1 gbuf_qn_253(.A(qn_in_253), .Y(g_23734));
AOI21X1 g60589(.A0 (n_7463), .A1 (g1222), .B0 (n_7462), .Y (n_7319));
AOI21X1 g60590(.A0 (n_7463), .A1 (g1223), .B0 (n_7462), .Y (n_7318));
NOR2X1 g60669(.A (n_7007), .B (n_7462), .Y (n_7317));
NOR2X1 g60672(.A (n_8266), .B (n_7316), .Y (n_7369));
XOR2X1 g60712(.A (n_4014), .B (n_7166), .Y (n_7315));
NOR2X1 g60789(.A (n_5963), .B (n_8487), .Y (n_7314));
MX2X1 g60831(.A (g403), .B (n_7310), .S0 (n_2667), .Y (n_7312));
MX2X1 g60832(.A (g402), .B (n_7310), .S0 (n_5526), .Y (n_7311));
MX2X1 g60833(.A (g404), .B (n_7310), .S0 (n_3271), .Y (n_7309));
NOR2X1 g60172(.A (n_7199), .B (n_7307), .Y (n_7308));
MX2X1 g60208(.A (g999), .B (n_7303), .S0 (g5472), .Y (n_7306));
MX2X1 g60209(.A (n_7303), .B (g1001), .S0 (n_6420), .Y (n_7304));
MX2X1 g60210(.A (g1000), .B (n_7303), .S0 (g6712), .Y (n_7301));
OAI21X1 g60222(.A0 (n_7150), .A1 (n_9369), .B0 (n_7145), .Y (n_7299));
NAND2X1 g60280(.A (n_7202), .B (n_9308), .Y (n_7297));
NAND2X1 g60320(.A (n_7200), .B (n_7157), .Y (n_7296));
AOI21X1 g60328(.A0 (n_6680), .A1 (n_6654), .B0 (n_7355), .Y (n_7295));
NOR2X1 g60370(.A (n_7293), .B (n_9425), .Y (n_7381));
NAND4X1 g60431(.A (n_7291), .B (n_4840), .C (n_9021), .D (n_6994), .Y(n_7292));
MX2X1 g60465(.A (g2396), .B (n_7287), .S0 (n_7115), .Y (n_7289));
MX2X1 g60466(.A (g2397), .B (n_7287), .S0 (n_7114), .Y (n_7288));
MX2X1 g60467(.A (g2398), .B (n_7287), .S0 (n_7112), .Y (n_7286));
MX2X1 g60471(.A (g1702), .B (n_7283), .S0 (n_7179), .Y (n_7285));
MX2X1 g60472(.A (g1703), .B (n_7283), .S0 (n_7178), .Y (n_7284));
MX2X1 g60473(.A (g1704), .B (n_7283), .S0 (n_7176), .Y (n_7282));
NAND3X1 g60505(.A (n_4290), .B (n_4511), .C (n_7281), .Y (n_7326));
NAND3X1 g60507(.A (n_4288), .B (n_4510), .C (n_7281), .Y (n_7324));
NAND3X1 g60509(.A (n_4286), .B (n_4509), .C (n_7281), .Y (n_7417));
NAND3X1 g60511(.A (n_4284), .B (n_4508), .C (n_7281), .Y (n_7418));
AOI21X1 g60518(.A0 (n_6164), .A1 (n_7267), .B0 (n_882), .Y (n_7591));
INVX1 g60521(.A (n_7279), .Y (n_7322));
INVX1 g60522(.A (n_7279), .Y (n_7280));
CLKBUFX1 gbuf_d_254(.A(n_7154), .Y(d_out_254));
CLKBUFX1 gbuf_q_254(.A(q_in_254), .Y(g1300));
CLKBUFX1 gbuf_d_255(.A(n_7148), .Y(d_out_255));
CLKBUFX1 gbuf_q_255(.A(q_in_255), .Y(g1009));
CLKBUFX1 gbuf_d_256(.A(n_7185), .Y(d_out_256));
CLKBUFX1 gbuf_q_256(.A(q_in_256), .Y(g417));
CLKBUFX1 gbuf_d_257(.A(n_7184), .Y(d_out_257));
CLKBUFX1 gbuf_q_257(.A(q_in_257), .Y(g420));
CLKBUFX1 gbuf_d_258(.A(n_7182), .Y(d_out_258));
CLKBUFX1 gbuf_q_258(.A(q_in_258), .Y(g423));
CLKBUFX1 gbuf_d_259(.A(n_7174), .Y(d_out_259));
CLKBUFX1 gbuf_q_259(.A(q_in_259), .Y(g408));
CLKBUFX1 gbuf_d_260(.A(n_7173), .Y(d_out_260));
CLKBUFX1 gbuf_q_260(.A(q_in_260), .Y(g411));
CLKBUFX1 gbuf_d_261(.A(n_7171), .Y(d_out_261));
CLKBUFX1 gbuf_q_261(.A(q_in_261), .Y(g414));
NAND2X2 g60563(.A (n_7189), .B (n_7277), .Y (n_7341));
NAND2X1 g60567(.A (n_7188), .B (n_7277), .Y (n_7278));
OAI21X1 g60568(.A0 (n_4046), .A1 (n_7273), .B0 (n_7281), .Y (n_7276));
OAI21X1 g60569(.A0 (n_4045), .A1 (n_7271), .B0 (n_7281), .Y (n_7275));
OAI21X1 g60570(.A0 (n_4043), .A1 (n_7273), .B0 (n_7281), .Y (n_7274));
OAI21X1 g60571(.A0 (n_4042), .A1 (n_7271), .B0 (n_7281), .Y (n_7272));
OAI21X1 g60572(.A0 (n_4297), .A1 (n_7273), .B0 (n_7281), .Y (n_7270));
OAI21X1 g60573(.A0 (n_4296), .A1 (n_7271), .B0 (n_7281), .Y (n_7269));
OAI21X1 g60575(.A0 (n_5906), .A1 (n_7190), .B0 (n_7267), .Y (n_7268));
OR2X1 g60576(.A (n_882), .B (n_7267), .Y (n_7631));
AOI22X1 g60600(.A0 (n_7233), .A1 (g7194), .B0 (g16399), .B1 (n_1689),.Y (n_7266));
NAND2X1 g60664(.A (n_1346), .B (n_7463), .Y (n_7264));
NAND2X1 g60666(.A (n_1256), .B (n_7463), .Y (n_7263));
NAND2X1 g60667(.A (n_1258), .B (n_7463), .Y (n_7262));
NAND2X1 g60668(.A (n_1344), .B (n_7463), .Y (n_7261));
NAND3X1 g60681(.A (n_7215), .B (n_8357), .C (n_9227), .Y (n_7260));
OAI21X1 g60694(.A0 (g_7108), .A1 (g_30261), .B0 (n_6310), .Y(n_7374));
CLKBUFX1 gbuf_d_262(.A(n_7146), .Y(d_out_262));
CLKBUFX1 gbuf_q_262(.A(q_in_262), .Y(g1010));
CLKBUFX1 gbuf_d_263(.A(n_7149), .Y(d_out_263));
CLKBUFX1 gbuf_q_263(.A(q_in_263), .Y(g1008));
NAND3X1 g60784(.A (n_5717), .B (n_7090), .C (n_7257), .Y (n_7258));
NOR2X1 g60792(.A (n_6414), .B (n_8398), .Y (n_7256));
NAND2X1 g60817(.A (g2374), .B (g2373), .Y (n_7253));
OAI21X1 g60818(.A0 (n_5163), .A1 (n_9673), .B0 (n_7160), .Y (n_7252));
CLKBUFX1 gbuf_d_264(.A(n_7153), .Y(d_out_264));
CLKBUFX1 gbuf_q_264(.A(q_in_264), .Y(g1303));
AOI21X1 g60853(.A0 (n_3790), .A1 (n_7032), .B0 (n_7168), .Y (n_7251));
XOR2X1 g60147(.A (n_5741), .B (n_7068), .Y (n_9611));
OAI21X1 g60945(.A0 (n_6072), .A1 (n_9222), .B0 (n_5890), .Y (n_7360));
AOI21X1 g60984(.A0 (n_7162), .A1 (n_5162), .B0 (n_7163), .Y (n_7249));
INVX4 g60405(.A (n_7355), .Y (n_7561));
INVX4 g60409(.A (n_7247), .Y (n_7246));
OAI22X1 g60459(.A0 (n_7144), .A1 (n_7337), .B0 (n_7221), .B1(n_7240), .Y (n_7242));
OAI22X1 g60460(.A0 (n_7143), .A1 (n_7337), .B0 (n_7222), .B1(n_7240), .Y (n_7241));
XOR2X1 g60477(.A (n_7138), .B (n_7141), .Y (n_7239));
XOR2X1 g60478(.A (n_7136), .B (n_7137), .Y (n_7238));
INVX1 g60492(.A (n_9063), .Y (n_7237));
INVX1 g60495(.A (n_9425), .Y (n_7235));
NAND2X1 g60523(.A (n_6080), .B (n_7196), .Y (n_7279));
CLKBUFX1 gbuf_d_265(.A(n_7074), .Y(d_out_265));
CLKBUFX1 gbuf_q_265(.A(q_in_265), .Y(g1994));
CLKBUFX1 gbuf_d_266(.A(n_7073), .Y(d_out_266));
CLKBUFX1 gbuf_q_266(.A(q_in_266), .Y(g1997));
CLKBUFX1 gbuf_d_267(.A(n_7070), .Y(d_out_267));
CLKBUFX1 gbuf_q_267(.A(q_in_267), .Y(g2000));
CLKBUFX1 gbuf_d_268(.A(n_7069), .Y(d_out_268));
CLKBUFX1 gbuf_q_268(.A(q_in_268), .Y(g1306));
CLKBUFX1 gbuf_d_269(.A(n_7064), .Y(d_out_269));
CLKBUFX1 gbuf_q_269(.A(q_in_269), .Y(g1985));
CLKBUFX1 gbuf_d_270(.A(n_7062), .Y(d_out_270));
CLKBUFX1 gbuf_q_270(.A(q_in_270), .Y(g1988));
CLKBUFX1 gbuf_d_271(.A(n_7060), .Y(d_out_271));
CLKBUFX1 gbuf_q_271(.A(q_in_271), .Y(g1991));
CLKBUFX1 gbuf_d_272(.A(n_7127), .Y(d_out_272));
CLKBUFX1 gbuf_q_272(.A(q_in_272), .Y(g3100));
CLKBUFX1 gbuf_d_273(.A(n_7126), .Y(d_out_273));
CLKBUFX1 gbuf_q_273(.A(q_in_273), .Y(g3101));
CLKBUFX1 gbuf_d_274(.A(n_7124), .Y(d_out_274));
CLKBUFX1 gbuf_q_274(.A(q_in_274), .Y(g3102));
CLKBUFX1 gbuf_d_275(.A(n_7119), .Y(d_out_275));
CLKBUFX1 gbuf_q_275(.A(q_in_275), .Y(g1801));
CLKBUFX1 gbuf_d_276(.A(n_7116), .Y(d_out_276));
CLKBUFX1 gbuf_q_276(.A(q_in_276), .Y(g1804));
CLKBUFX1 gbuf_d_277(.A(n_7233), .Y(d_out_277));
CLKBUFX1 gbuf_q_277(.A(q_in_277), .Y(g16355));
CLKBUFX1 gbuf_d_278(.A(n_7120), .Y(d_out_278));
CLKBUFX1 gbuf_q_278(.A(q_in_278), .Y(g1798));
CLKBUFX1 gbuf_d_279(.A(n_7110), .Y(d_out_279));
CLKBUFX1 gbuf_q_279(.A(q_in_279), .Y(g2477));
CLKBUFX1 gbuf_d_280(.A(n_7109), .Y(d_out_280));
CLKBUFX1 gbuf_q_280(.A(q_in_280), .Y(g2478));
CLKBUFX1 gbuf_d_281(.A(n_7107), .Y(d_out_281));
CLKBUFX1 gbuf_q_281(.A(q_in_281), .Y(g2479));
CLKBUFX1 gbuf_d_282(.A(n_7099), .Y(d_out_282));
CLKBUFX1 gbuf_q_282(.A(q_in_282), .Y(g1784));
CLKBUFX1 gbuf_d_283(.A(n_7102), .Y(d_out_283));
CLKBUFX1 gbuf_q_283(.A(q_in_283), .Y(g1783));
CLKBUFX1 gbuf_d_284(.A(n_7101), .Y(d_out_284));
CLKBUFX1 gbuf_q_284(.A(q_in_284), .Y(g1785));
CLKBUFX1 gbuf_d_285(.A(n_7106), .Y(d_out_285));
CLKBUFX1 gbuf_q_285(.A(q_in_285), .Y(g1789));
CLKBUFX1 gbuf_d_286(.A(n_7103), .Y(d_out_286));
CLKBUFX1 gbuf_q_286(.A(q_in_286), .Y(g1792));
CLKBUFX1 gbuf_d_287(.A(n_7105), .Y(d_out_287));
CLKBUFX1 gbuf_q_287(.A(q_in_287), .Y(g1795));
CLKBUFX1 gbuf_d_288(.A(n_7096), .Y(d_out_288));
CLKBUFX1 gbuf_q_288(.A(q_in_288), .Y(g426));
CLKBUFX1 gbuf_d_289(.A(n_7095), .Y(d_out_289));
CLKBUFX1 gbuf_q_289(.A(q_in_289), .Y(g427));
CLKBUFX1 gbuf_d_290(.A(n_7093), .Y(d_out_290));
CLKBUFX1 gbuf_q_290(.A(q_in_290), .Y(g428));
CLKBUFX1 gbuf_d_291(.A(n_7080), .Y(d_out_291));
CLKBUFX1 gbuf_q_291(.A(q_in_291), .Y(g447));
CLKBUFX1 gbuf_d_292(.A(n_7079), .Y(d_out_292));
CLKBUFX1 gbuf_q_292(.A(q_in_292), .Y(g448));
CLKBUFX1 gbuf_d_293(.A(n_7077), .Y(d_out_293));
CLKBUFX1 gbuf_q_293(.A(q_in_293), .Y(g449));
NAND2X1 g60561(.A (n_8571), .B (n_4627), .Y (n_7291));
NAND2X1 g60565(.A (n_7123), .B (n_4627), .Y (n_7232));
OAI21X1 g60593(.A0 (n_1337), .A1 (n_7228), .B0 (n_7135), .Y (n_7230));
OAI21X1 g60594(.A0 (n_1347), .A1 (n_7228), .B0 (n_7134), .Y (n_7229));
OAI21X1 g60595(.A0 (n_1343), .A1 (n_7228), .B0 (n_7132), .Y (n_7227));
OAI21X1 g60596(.A0 (n_1186), .A1 (n_7228), .B0 (n_7131), .Y (n_7226));
OAI21X1 g60597(.A0 (n_1189), .A1 (n_7228), .B0 (n_7130), .Y (n_7225));
OAI21X1 g60598(.A0 (n_1259), .A1 (n_7228), .B0 (n_7129), .Y (n_7224));
XOR2X1 g60621(.A (n_7222), .B (n_7221), .Y (n_7223));
AND2X1 g60786(.A (n_9219), .B (n_8357), .Y (n_7218));
NAND2X1 g60790(.A (n_6592), .B (n_7165), .Y (n_7316));
OAI21X1 g60819(.A0 (n_8685), .A1 (n_8484), .B0 (n_7085), .Y (n_7217));
AOI21X1 g60829(.A0 (n_7215), .A1 (n_7214), .B0 (n_6046), .Y (n_8187));
CLKBUFX1 gbuf_d_294(.A(n_7083), .Y(d_out_294));
CLKBUFX1 gbuf_qn_294(.A(qn_in_294), .Y(g1679));
NAND2X1 g60899(.A (n_5292), .B (n_7208), .Y (n_7213));
AOI21X1 g60900(.A0 (n_8929), .A1 (n_9227), .B0 (n_6972), .Y (n_7212));
NOR2X1 g60902(.A (n_7208), .B (g309), .Y (n_7209));
AOI21X1 g60982(.A0 (n_7087), .A1 (n_9637), .B0 (n_7088), .Y (n_7205));
INVX1 g60365(.A (n_9308), .Y (n_7204));
INVX2 g60407(.A (n_7203), .Y (n_7355));
CLKBUFX3 g60413(.A (n_7203), .Y (n_7247));
INVX1 g60414(.A (n_7203), .Y (n_7202));
AOI21X1 g60436(.A0 (n_7022), .A1 (g_23734), .B0 (n_7065), .Y(n_7201));
AOI22X1 g60457(.A0 (n_7156), .A1 (n_9666), .B0 (n_4670), .B1(n_6448), .Y (n_7200));
AOI21X1 g60461(.A0 (n_45), .A1 (n_7067), .B0 (n_7066), .Y (n_7199));
NAND3X1 g60516(.A (n_6718), .B (n_7054), .C (n_6778), .Y (n_7198));
NAND3X1 g60517(.A (n_6715), .B (n_9257), .C (n_6851), .Y (n_7197));
CLKBUFX1 gbuf_d_295(.A(n_7045), .Y(d_out_295));
CLKBUFX1 gbuf_q_295(.A(q_in_295), .Y(g1807));
CLKBUFX1 gbuf_d_296(.A(n_7044), .Y(d_out_296));
CLKBUFX1 gbuf_q_296(.A(q_in_296), .Y(g1808));
CLKBUFX1 gbuf_d_297(.A(n_7042), .Y(d_out_297));
CLKBUFX1 gbuf_q_297(.A(q_in_297), .Y(g1809));
CLKBUFX1 gbuf_d_298(.A(n_7029), .Y(d_out_298));
CLKBUFX1 gbuf_q_298(.A(q_in_298), .Y(g438));
CLKBUFX1 gbuf_d_299(.A(n_7028), .Y(d_out_299));
CLKBUFX1 gbuf_q_299(.A(q_in_299), .Y(g441));
CLKBUFX1 gbuf_d_300(.A(n_7026), .Y(d_out_300));
CLKBUFX1 gbuf_q_300(.A(q_in_300), .Y(g444));
NAND2X1 g60577(.A (n_7050), .B (g1880), .Y (n_7196));
AOI21X1 g60586(.A0 (n_7005), .A1 (n_7194), .B0 (n_6999), .Y (n_7287));
CLKBUFX1 gbuf_d_301(.A(n_7057), .Y(d_out_301));
CLKBUFX1 gbuf_qn_301(.A(qn_in_301), .Y(g_22538));
AOI21X1 g60588(.A0 (n_7004), .A1 (n_5477), .B0 (n_6996), .Y (n_7283));
AOI21X1 g60660(.A0 (n_6995), .A1 (n_7194), .B0 (n_6413), .Y (n_7195));
AOI21X1 g60661(.A0 (n_6992), .A1 (n_5477), .B0 (n_6602), .Y (n_7193));
AND2X1 g60663(.A (n_7463), .B (n_6219), .Y (n_7281));
OR2X1 g60665(.A (n_7463), .B (n_7190), .Y (n_7267));
AOI22X1 g60686(.A0 (n_6989), .A1 (n_7186), .B0 (n_6850), .B1(n_6713), .Y (n_7189));
AOI22X1 g60695(.A0 (n_6991), .A1 (n_7187), .B0 (n_6691), .B1(n_7186), .Y (n_7188));
MX2X1 g60699(.A (g417), .B (n_7183), .S0 (n_6914), .Y (n_7185));
MX2X1 g60700(.A (g420), .B (n_7183), .S0 (g6447), .Y (n_7184));
MX2X1 g60701(.A (g423), .B (n_7183), .S0 (n_6917), .Y (n_7182));
AND2X1 g60808(.A (n_7177), .B (n_6832), .Y (n_7179));
AND2X1 g60810(.A (n_7177), .B (g5511), .Y (n_7178));
AND2X1 g60811(.A (n_7177), .B (n_3190), .Y (n_7176));
MX2X1 g60834(.A (g408), .B (n_7172), .S0 (n_6914), .Y (n_7174));
MX2X1 g60835(.A (g411), .B (n_7172), .S0 (g6447), .Y (n_7173));
MX2X1 g60836(.A (g414), .B (n_7172), .S0 (n_6917), .Y (n_7171));
CLKBUFX1 gbuf_d_302(.A(n_7031), .Y(d_out_302));
CLKBUFX1 gbuf_qn_302(.A(qn_in_302), .Y(g2373));
NOR2X1 g60910(.A (n_3790), .B (n_7032), .Y (n_7168));
INVX1 g60911(.A (n_7165), .Y (n_7166));
AOI21X1 g60983(.A0 (n_7038), .A1 (n_4756), .B0 (n_7039), .Y (n_7164));
OR2X1 g61013(.A (n_9270), .B (n_7091), .Y (n_7310));
NOR2X1 g61049(.A (n_7162), .B (n_5162), .Y (n_7163));
NAND3X1 g61054(.A (n_7162), .B (n_6531), .C (n_5163), .Y (n_7160));
NOR2X1 g60415(.A (n_9311), .B (n_9304), .Y (n_7203));
AND2X1 g60427(.A (n_7058), .B (n_9375), .Y (n_7303));
NAND4X1 g60432(.A (n_7156), .B (n_8653), .C (n_7155), .D (n_6635), .Y(n_7157));
MX2X1 g60449(.A (g1300), .B (n_7152), .S0 (g6750), .Y (n_7154));
MX2X1 g60450(.A (g1303), .B (n_7152), .S0 (g6944), .Y (n_7153));
NAND2X1 g60454(.A (n_7023), .B (n_6788), .Y (n_7150));
MX2X1 g60468(.A (g1008), .B (n_7147), .S0 (n_6944), .Y (n_7149));
MX2X1 g60469(.A (g1009), .B (n_7147), .S0 (n_6943), .Y (n_7148));
MX2X1 g60470(.A (g1010), .B (n_7147), .S0 (n_6941), .Y (n_7146));
CLKBUFX1 gbuf_d_303(.A(n_6968), .Y(d_out_303));
CLKBUFX1 gbuf_q_303(.A(q_in_303), .Y(g614));
CLKBUFX1 gbuf_d_304(.A(n_6966), .Y(d_out_304));
CLKBUFX1 gbuf_q_304(.A(q_in_304), .Y(g617));
CLKBUFX1 gbuf_d_305(.A(n_6960), .Y(d_out_305));
CLKBUFX1 gbuf_q_305(.A(q_in_305), .Y(g608));
CLKBUFX1 gbuf_d_306(.A(n_6958), .Y(d_out_306));
CLKBUFX1 gbuf_q_306(.A(q_in_306), .Y(g611));
CLKBUFX1 gbuf_d_307(.A(n_7002), .Y(d_out_307));
CLKBUFX1 gbuf_q_307(.A(q_in_307), .Y(g_32037));
NAND2X1 g60566(.A (n_7020), .B (n_9369), .Y (n_7145));
AOI21X1 g60610(.A0 (n_7139), .A1 (n_7142), .B0 (n_6932), .Y (n_7144));
AOI21X1 g60611(.A0 (n_7140), .A1 (n_7142), .B0 (n_6931), .Y (n_7143));
XOR2X1 g60622(.A (n_7140), .B (n_7139), .Y (n_7141));
XOR2X1 g60623(.A (n_7010), .B (n_7008), .Y (n_7138));
XOR2X1 g60624(.A (n_7018), .B (n_7016), .Y (n_7137));
XOR2X1 g60625(.A (n_7012), .B (n_7014), .Y (n_7136));
NAND2X1 g60652(.A (n_7019), .B (n_7142), .Y (n_7135));
NAND2X1 g60653(.A (n_7017), .B (n_7142), .Y (n_7134));
NAND2X1 g60654(.A (n_7015), .B (n_7142), .Y (n_7132));
NAND2X1 g60655(.A (n_7013), .B (n_7142), .Y (n_7131));
NAND2X1 g60656(.A (n_7011), .B (n_7142), .Y (n_7130));
NAND2X1 g60657(.A (n_7009), .B (n_7142), .Y (n_7129));
CLKBUFX1 gbuf_d_308(.A(n_6962), .Y(d_out_308));
CLKBUFX1 gbuf_q_308(.A(q_in_308), .Y(g605));
MX2X1 g60688(.A (g3100), .B (n_7125), .S0 (g8106), .Y (n_7127));
MX2X1 g60689(.A (g3101), .B (n_7125), .S0 (g8030), .Y (n_7126));
MX2X1 g60690(.A (g3102), .B (n_7125), .S0 (g3109), .Y (n_7124));
AOI22X1 g60692(.A0 (n_6929), .A1 (n_9021), .B0 (n_6689), .B1(n_9014), .Y (n_7123));
MX2X1 g60705(.A (g1798), .B (n_7118), .S0 (g5511), .Y (n_7120));
MX2X1 g60706(.A (g1801), .B (n_7118), .S0 (n_3190), .Y (n_7119));
MX2X1 g60707(.A (g1804), .B (n_7118), .S0 (n_6832), .Y (n_7116));
AND2X1 g60799(.A (n_7113), .B (n_6611), .Y (n_7115));
AND2X1 g60801(.A (n_7113), .B (g5555), .Y (n_7114));
AND2X1 g60802(.A (n_7113), .B (n_2180), .Y (n_7112));
NAND2X1 g60815(.A (n_6986), .B (n_7337), .Y (n_7336));
CLKBUFX1 gbuf_d_309(.A(n_6963), .Y(d_out_309));
CLKBUFX1 gbuf_q_309(.A(q_in_309), .Y(g620));
MX2X1 g60825(.A (g1193), .B (n_6925), .S0 (g1192), .Y (n_7233));
MX2X1 g60837(.A (g2477), .B (n_7108), .S0 (n_4970), .Y (n_7110));
MX2X1 g60838(.A (g2478), .B (n_7108), .S0 (n_2561), .Y (n_7109));
MX2X1 g60839(.A (g2479), .B (n_7108), .S0 (n_3233), .Y (n_7107));
MX2X1 g60843(.A (g1789), .B (n_7104), .S0 (g5511), .Y (n_7106));
MX2X1 g60844(.A (g1795), .B (n_7104), .S0 (n_6832), .Y (n_7105));
MX2X1 g60845(.A (g1792), .B (n_7104), .S0 (n_3190), .Y (n_7103));
MX2X1 g60850(.A (g1783), .B (n_7100), .S0 (n_5371), .Y (n_7102));
MX2X1 g60851(.A (g1785), .B (n_7100), .S0 (n_3474), .Y (n_7101));
MX2X1 g60852(.A (g1784), .B (n_7100), .S0 (n_2859), .Y (n_7099));
CLKBUFX1 gbuf_d_310(.A(n_6982), .Y(d_out_310));
CLKBUFX1 gbuf_q_310(.A(q_in_310), .Y(g_30261));
NOR2X1 g60912(.A (n_6516), .B (n_8727), .Y (n_7165));
NAND2X1 g60934(.A (n_6979), .B (n_6473), .Y (n_7293));
MX2X1 g60971(.A (n_7094), .B (g426), .S0 (n_6918), .Y (n_7096));
MX2X1 g60972(.A (n_7094), .B (g427), .S0 (n_6916), .Y (n_7095));
MX2X1 g60973(.A (n_7094), .B (g428), .S0 (n_6913), .Y (n_7093));
INVX1 g61023(.A (n_9226), .Y (n_7208));
NAND2X2 g61031(.A (n_7089), .B (n_7091), .Y (n_7891));
NAND2X1 g61032(.A (n_7089), .B (n_7215), .Y (n_7090));
NOR2X1 g61035(.A (n_7087), .B (n_9637), .Y (n_7088));
NAND3X1 g61059(.A (n_7087), .B (n_6432), .C (n_8685), .Y (n_7085));
NAND2X1 g61065(.A (n_6971), .B (n_6472), .Y (n_7083));
INVX1 g61069(.A (n_9225), .Y (n_7082));
MX2X1 g61111(.A (n_7078), .B (g447), .S0 (n_6903), .Y (n_7080));
MX2X1 g61112(.A (n_7078), .B (g448), .S0 (n_6904), .Y (n_7079));
MX2X1 g61113(.A (n_7078), .B (g449), .S0 (n_6901), .Y (n_7077));
MX2X1 g60442(.A (g1994), .B (n_7072), .S0 (g7052), .Y (n_7074));
MX2X1 g60443(.A (g1997), .B (n_7072), .S0 (g7194), .Y (n_7073));
MX2X1 g60444(.A (g2000), .B (n_7072), .S0 (n_6626), .Y (n_7070));
OAI21X1 g60448(.A0 (n_7021), .A1 (n_3220), .B0 (n_3346), .Y (n_7069));
OR2X1 g60494(.A (g_27975), .B (n_7067), .Y (n_7068));
NOR2X1 g60513(.A (n_45), .B (n_7067), .Y (n_7066));
NAND2X1 g60514(.A (n_7067), .B (n_6865), .Y (n_7065));
MX2X1 g60524(.A (g1985), .B (n_7061), .S0 (g7052), .Y (n_7064));
MX2X1 g60525(.A (g1988), .B (n_7061), .S0 (g7194), .Y (n_7062));
MX2X1 g60526(.A (g1991), .B (n_7061), .S0 (n_6626), .Y (n_7060));
XOR2X1 g60542(.A (n_4670), .B (n_6880), .Y (n_7058));
CLKBUFX1 gbuf_d_311(.A(n_6951), .Y(d_out_311));
CLKBUFX1 gbuf_q_311(.A(q_in_311), .Y(g2492));
CLKBUFX1 gbuf_d_312(.A(n_6897), .Y(d_out_312));
CLKBUFX1 gbuf_q_312(.A(q_in_312), .Y(g1291));
CLKBUFX1 gbuf_d_313(.A(n_6956), .Y(d_out_313));
CLKBUFX1 gbuf_q_313(.A(q_in_313), .Y(g1294));
CLKBUFX1 gbuf_d_314(.A(n_6955), .Y(d_out_314));
CLKBUFX1 gbuf_q_314(.A(q_in_314), .Y(g1297));
CLKBUFX1 gbuf_d_315(.A(n_6950), .Y(d_out_315));
CLKBUFX1 gbuf_q_315(.A(q_in_315), .Y(g2495));
CLKBUFX1 gbuf_d_316(.A(n_6948), .Y(d_out_316));
CLKBUFX1 gbuf_q_316(.A(q_in_316), .Y(g2498));
CLKBUFX1 gbuf_d_317(.A(n_6940), .Y(d_out_317));
CLKBUFX1 gbuf_q_317(.A(q_in_317), .Y(g2483));
CLKBUFX1 gbuf_d_318(.A(n_6909), .Y(d_out_318));
CLKBUFX1 gbuf_q_318(.A(q_in_318), .Y(g429));
CLKBUFX1 gbuf_d_319(.A(n_6908), .Y(d_out_319));
CLKBUFX1 gbuf_q_319(.A(q_in_319), .Y(g432));
CLKBUFX1 gbuf_d_320(.A(n_6906), .Y(d_out_320));
CLKBUFX1 gbuf_q_320(.A(q_in_320), .Y(g435));
NAND2X1 g60562(.A (n_6952), .B (n_9369), .Y (n_7156));
NOR2X1 g60578(.A (n_6936), .B (n_7307), .Y (n_7057));
NAND3X1 g60679(.A (n_8419), .B (n_7000), .C (n_8573), .Y (n_7054));
OAI21X1 g60687(.A0 (n_8794), .A1 (n_864), .B0 (n_599), .Y (n_7050));
AND2X1 g60773(.A (n_5103), .B (n_6934), .Y (n_7221));
AND2X1 g60775(.A (n_5100), .B (n_6933), .Y (n_7222));
INVX1 g60782(.A (n_7007), .Y (n_7463));
NAND3X1 g60798(.A (n_5169), .B (n_6855), .C (n_9014), .Y (n_7049));
NAND3X1 g60807(.A (n_5331), .B (n_6853), .C (n_7186), .Y (n_7048));
NAND4X1 g60935(.A (n_1188), .B (n_6692), .C (n_1368), .D (n_593), .Y(n_7047));
OAI21X1 g60937(.A0 (n_3812), .A1 (n_8437), .B0 (n_6924), .Y (n_7046));
OAI21X1 g60961(.A0 (n_6199), .A1 (n_6836), .B0 (n_6035), .Y (n_7177));
MX2X1 g60977(.A (n_7043), .B (g1807), .S0 (n_6833), .Y (n_7045));
MX2X1 g60978(.A (n_7043), .B (g1808), .S0 (n_6831), .Y (n_7044));
MX2X1 g60979(.A (n_7043), .B (g1809), .S0 (n_6828), .Y (n_7042));
NOR2X1 g61018(.A (n_5543), .B (n_9270), .Y (n_7214));
NOR2X1 g61047(.A (n_7038), .B (n_4756), .Y (n_7039));
NAND3X1 g61050(.A (n_7038), .B (n_6319), .C (n_4757), .Y (n_7036));
INVX1 g61057(.A (n_8727), .Y (n_7032));
NAND2X1 g61064(.A (n_6911), .B (n_6368), .Y (n_7031));
OAI21X1 g61074(.A0 (n_9192), .A1 (n_6974), .B0 (n_6900), .Y (n_7030));
MX2X1 g61093(.A (g438), .B (n_7027), .S0 (n_6914), .Y (n_7029));
MX2X1 g61094(.A (g441), .B (n_7027), .S0 (g6447), .Y (n_7028));
MX2X1 g61095(.A (g444), .B (n_7027), .S0 (n_6917), .Y (n_7026));
INVX1 g61261(.A (n_7025), .Y (n_7162));
CLKBUFX1 gbuf_d_321(.A(n_7125), .Y(d_out_321));
CLKBUFX1 gbuf_q_321(.A(q_in_321), .Y(g1234));
CLKBUFX1 gbuf_d_322(.A(n_6937), .Y(d_out_322));
CLKBUFX1 gbuf_q_322(.A(q_in_322), .Y(g2489));
CLKBUFX1 gbuf_d_323(.A(n_6939), .Y(d_out_323));
CLKBUFX1 gbuf_q_323(.A(q_in_323), .Y(g2486));
NAND3X1 g60515(.A (n_6450), .B (n_6877), .C (n_6625), .Y (n_7023));
CLKBUFX1 gbuf_d_324(.A(n_6868), .Y(d_out_324));
CLKBUFX1 gbuf_q_324(.A(q_in_324), .Y(g1101));
CLKBUFX1 gbuf_d_325(.A(n_6872), .Y(d_out_325));
CLKBUFX1 gbuf_q_325(.A(q_in_325), .Y(g1090));
CLKBUFX1 gbuf_d_326(.A(n_6874), .Y(d_out_326));
CLKBUFX1 gbuf_q_326(.A(q_in_326), .Y(g1091));
CLKBUFX1 gbuf_d_327(.A(n_6823), .Y(d_out_327));
CLKBUFX1 gbuf_q_327(.A(q_in_327), .Y(g2688));
CLKBUFX1 gbuf_d_328(.A(n_6818), .Y(d_out_328));
CLKBUFX1 gbuf_q_328(.A(q_in_328), .Y(g2694));
CLKBUFX1 gbuf_d_329(.A(n_6896), .Y(d_out_329));
CLKBUFX1 gbuf_q_329(.A(q_in_329), .Y(g2679));
CLKBUFX1 gbuf_d_330(.A(n_6894), .Y(d_out_330));
CLKBUFX1 gbuf_q_330(.A(q_in_330), .Y(g2682));
CLKBUFX1 gbuf_d_331(.A(n_6875), .Y(d_out_331));
CLKBUFX1 gbuf_q_331(.A(q_in_331), .Y(g1089));
CLKBUFX1 gbuf_d_332(.A(n_6870), .Y(d_out_332));
CLKBUFX1 gbuf_q_332(.A(q_in_332), .Y(g1098));
CLKBUFX1 gbuf_d_333(.A(n_6871), .Y(d_out_333));
CLKBUFX1 gbuf_q_333(.A(q_in_333), .Y(g1095));
CLKBUFX1 gbuf_d_334(.A(n_6861), .Y(d_out_334));
CLKBUFX1 gbuf_q_334(.A(q_in_334), .Y(g2503));
CLKBUFX1 gbuf_d_335(.A(n_6864), .Y(d_out_335));
CLKBUFX1 gbuf_q_335(.A(q_in_335), .Y(g2501));
CLKBUFX1 gbuf_d_336(.A(n_6846), .Y(d_out_336));
CLKBUFX1 gbuf_q_336(.A(q_in_336), .Y(g1828));
CLKBUFX1 gbuf_d_337(.A(n_6843), .Y(d_out_337));
CLKBUFX1 gbuf_q_337(.A(q_in_337), .Y(g1830));
CLKBUFX1 gbuf_d_338(.A(n_6845), .Y(d_out_338));
CLKBUFX1 gbuf_q_338(.A(q_in_338), .Y(g1829));
CLKBUFX1 gbuf_d_339(.A(n_6814), .Y(d_out_339));
CLKBUFX1 gbuf_q_339(.A(q_in_339), .Y(g343));
CLKBUFX1 gbuf_d_340(.A(n_6813), .Y(d_out_340));
CLKBUFX1 gbuf_q_340(.A(q_in_340), .Y(g346));
CLKBUFX1 gbuf_d_341(.A(n_6811), .Y(d_out_341));
CLKBUFX1 gbuf_q_341(.A(q_in_341), .Y(g354));
CLKBUFX1 gbuf_d_342(.A(n_6810), .Y(d_out_342));
CLKBUFX1 gbuf_q_342(.A(q_in_342), .Y(g373));
CLKBUFX1 gbuf_d_343(.A(n_6805), .Y(d_out_343));
CLKBUFX1 gbuf_q_343(.A(q_in_343), .Y(g384));
CLKBUFX1 gbuf_d_344(.A(n_6808), .Y(d_out_344));
CLKBUFX1 gbuf_q_344(.A(q_in_344), .Y(g376));
CLKBUFX1 gbuf_d_345(.A(n_6895), .Y(d_out_345));
CLKBUFX1 gbuf_q_345(.A(q_in_345), .Y(g1724));
CLKBUFX1 gbuf_d_346(.A(n_6891), .Y(d_out_346));
CLKBUFX1 gbuf_q_346(.A(q_in_346), .Y(g1727));
CLKBUFX1 gbuf_d_347(.A(n_6889), .Y(d_out_347));
CLKBUFX1 gbuf_q_347(.A(q_in_347), .Y(g1735));
CLKBUFX1 gbuf_d_348(.A(n_6888), .Y(d_out_348));
CLKBUFX1 gbuf_q_348(.A(q_in_348), .Y(g1754));
CLKBUFX1 gbuf_d_349(.A(n_6883), .Y(d_out_349));
CLKBUFX1 gbuf_q_349(.A(q_in_349), .Y(g1765));
OR2X1 g60574(.A (n_7022), .B (g_23734), .Y (n_7067));
AOI21X1 g60587(.A0 (n_6787), .A1 (n_8653), .B0 (n_8968), .Y (n_7147));
INVX1 g60615(.A (n_7021), .Y (n_7152));
CLKBUFX1 gbuf_d_350(.A(n_6892), .Y(d_out_350));
CLKBUFX1 gbuf_q_350(.A(q_in_350), .Y(g2685));
AOI22X1 g60693(.A0 (n_6786), .A1 (n_6448), .B0 (n_8533), .B1(n_3959), .Y (n_7020));
INVX1 g60761(.A (n_7018), .Y (n_7019));
INVX1 g60763(.A (n_7016), .Y (n_7017));
INVX1 g60765(.A (n_7014), .Y (n_7015));
INVX1 g60767(.A (n_7012), .Y (n_7013));
INVX1 g60769(.A (n_7010), .Y (n_7011));
INVX1 g60771(.A (n_7008), .Y (n_7009));
CLKBUFX1 gbuf_d_351(.A(n_6863), .Y(d_out_351));
CLKBUFX1 gbuf_q_351(.A(q_in_351), .Y(g2502));
NAND3X1 g60783(.A (n_8794), .B (n_31), .C (n_5186), .Y (n_7007));
AND2X1 g60800(.A (n_9021), .B (n_8419), .Y (n_7005));
AND2X1 g60809(.A (n_7187), .B (n_9254), .Y (n_7004));
NAND2X1 g60820(.A (g986), .B (g985), .Y (n_7003));
OAI21X1 g60821(.A0 (n_6443), .A1 (n_6935), .B0 (n_7337), .Y (n_7333));
AOI21X1 g60822(.A0 (n_6712), .A1 (n_43), .B0 (n_6866), .Y (n_7002));
NAND2X1 g60917(.A (n_5332), .B (n_9654), .Y (n_6995));
NOR2X1 g60922(.A (n_9654), .B (g2384), .Y (n_6994));
NAND2X1 g60926(.A (n_5492), .B (n_6987), .Y (n_6992));
AOI21X1 g60927(.A0 (n_8548), .A1 (n_9255), .B0 (n_6690), .Y (n_6991));
NAND2X1 g60928(.A (n_6859), .B (n_6836), .Y (n_6989));
NOR2X1 g60929(.A (n_6987), .B (n_5531), .Y (n_6988));
NAND2X1 g60936(.A (n_6423), .B (n_6860), .Y (n_6986));
OAI21X1 g60953(.A0 (n_6068), .A1 (n_8567), .B0 (n_5886), .Y (n_7113));
CLKBUFX1 gbuf_d_352(.A(n_6821), .Y(d_out_352));
CLKBUFX1 gbuf_q_352(.A(q_in_352), .Y(g2691));
XOR2X1 g60981(.A (n_6212), .B (n_6769), .Y (n_7183));
AND2X1 g61010(.A (n_8929), .B (n_9219), .Y (n_6985));
NAND2X1 g61062(.A (n_6827), .B (n_6231), .Y (n_6982));
CLKBUFX1 gbuf_d_353(.A(n_6886), .Y(d_out_353));
CLKBUFX1 gbuf_q_353(.A(q_in_353), .Y(g1757));
OAI21X1 g61087(.A0 (n_6970), .A1 (n_6602), .B0 (n_6837), .Y (n_6979));
XOR2X1 g61102(.A (n_4339), .B (n_6759), .Y (n_6978));
XOR2X1 g61123(.A (n_6558), .B (n_6752), .Y (n_7172));
INVX1 g61245(.A (n_6975), .Y (n_7087));
NAND3X1 g61262(.A (n_6974), .B (n_6177), .C (n_6055), .Y (n_7025));
INVX1 g61301(.A (n_9270), .Y (n_7089));
OAI21X1 g61335(.A0 (n_6970), .A1 (n_6969), .B0 (n_6815), .Y (n_6971));
MX2X1 g60445(.A (g614), .B (n_6965), .S0 (g6485), .Y (n_6968));
XOR2X1 g61354(.A (n_4433), .B (n_6899), .Y (n_6967));
MX2X1 g60446(.A (g617), .B (n_6965), .S0 (g6642), .Y (n_6966));
MX2X1 g60447(.A (g620), .B (n_6965), .S0 (n_4601), .Y (n_6963));
MX2X1 g60527(.A (g605), .B (n_6959), .S0 (g6485), .Y (n_6962));
MX2X1 g60528(.A (g608), .B (n_6959), .S0 (g6642), .Y (n_6960));
MX2X1 g60529(.A (g611), .B (n_6959), .S0 (n_4601), .Y (n_6958));
MX2X1 g60532(.A (g1294), .B (n_6954), .S0 (g6944), .Y (n_6956));
MX2X1 g60533(.A (n_6954), .B (g1297), .S0 (n_3220), .Y (n_6955));
CLKBUFX1 gbuf_d_354(.A(n_6793), .Y(d_out_354));
CLKBUFX1 gbuf_q_354(.A(q_in_354), .Y(g1104));
CLKBUFX1 gbuf_d_355(.A(n_6792), .Y(d_out_355));
CLKBUFX1 gbuf_q_355(.A(q_in_355), .Y(g1107));
CLKBUFX1 gbuf_d_356(.A(n_6776), .Y(d_out_356));
CLKBUFX1 gbuf_q_356(.A(q_in_356), .Y(g1819));
CLKBUFX1 gbuf_d_357(.A(n_6775), .Y(d_out_357));
CLKBUFX1 gbuf_q_357(.A(q_in_357), .Y(g1822));
CLKBUFX1 gbuf_d_358(.A(n_6763), .Y(d_out_358));
CLKBUFX1 gbuf_q_358(.A(q_in_358), .Y(g1816));
CLKBUFX1 gbuf_d_359(.A(n_6762), .Y(d_out_359));
CLKBUFX1 gbuf_q_359(.A(q_in_359), .Y(g1810));
CLKBUFX1 gbuf_d_360(.A(n_6802), .Y(d_out_360));
CLKBUFX1 gbuf_q_360(.A(q_in_360), .Y(g391));
CLKBUFX1 gbuf_d_361(.A(n_6803), .Y(d_out_361));
CLKBUFX1 gbuf_q_361(.A(q_in_361), .Y(g388));
CLKBUFX1 gbuf_d_362(.A(n_6800), .Y(d_out_362));
CLKBUFX1 gbuf_q_362(.A(q_in_362), .Y(g398));
CLKBUFX1 gbuf_d_363(.A(n_6798), .Y(d_out_363));
CLKBUFX1 gbuf_q_363(.A(q_in_363), .Y(g1772));
CLKBUFX1 gbuf_d_364(.A(n_6799), .Y(d_out_364));
CLKBUFX1 gbuf_q_364(.A(q_in_364), .Y(g1769));
CLKBUFX1 gbuf_d_365(.A(n_6796), .Y(d_out_365));
CLKBUFX1 gbuf_q_365(.A(q_in_365), .Y(g1779));
CLKBUFX1 gbuf_d_366(.A(n_6790), .Y(d_out_366));
CLKBUFX1 gbuf_q_366(.A(q_in_366), .Y(g1110));
OAI22X1 g60613(.A0 (n_6728), .A1 (n_6947), .B0 (n_6946), .B1(n_5323), .Y (n_7072));
MX2X1 g60616(.A (n_6729), .B (n_7271), .S0 (n_6947), .Y (n_7021));
CLKBUFX1 gbuf_d_367(.A(n_6773), .Y(d_out_367));
CLKBUFX1 gbuf_q_367(.A(q_in_367), .Y(g1825));
AOI22X1 g60685(.A0 (n_6723), .A1 (n_3959), .B0 (n_6624), .B1(n_6448), .Y (n_6952));
MX2X1 g60702(.A (g2492), .B (n_6949), .S0 (g5555), .Y (n_6951));
MX2X1 g60703(.A (g2495), .B (n_6949), .S0 (g7264), .Y (n_6950));
MX2X1 g60704(.A (g2498), .B (n_6949), .S0 (n_6611), .Y (n_6948));
OAI22X1 g60708(.A0 (n_6724), .A1 (n_6947), .B0 (n_6946), .B1(n_4317), .Y (n_7061));
NAND3X1 g60762(.A (n_4696), .B (n_4952), .C (n_6945), .Y (n_7018));
NAND3X1 g60764(.A (n_4694), .B (n_4951), .C (n_6945), .Y (n_7016));
NAND3X1 g60766(.A (n_4692), .B (n_4950), .C (n_6945), .Y (n_7014));
NAND3X1 g60768(.A (n_4690), .B (n_4949), .C (n_6945), .Y (n_7012));
NAND3X1 g60770(.A (n_4688), .B (n_4948), .C (n_6945), .Y (n_7010));
NAND3X1 g60772(.A (n_4686), .B (n_4947), .C (n_6945), .Y (n_7008));
NAND3X1 g60774(.A (n_4684), .B (n_4945), .C (n_6945), .Y (n_7139));
NAND3X1 g60776(.A (n_4682), .B (n_4941), .C (n_6945), .Y (n_7140));
NOR2X1 g60803(.A (n_6942), .B (n_6420), .Y (n_6944));
NOR2X1 g60805(.A (n_6942), .B (n_8305), .Y (n_6943));
NOR2X1 g60806(.A (n_6942), .B (n_2343), .Y (n_6941));
MX2X1 g60840(.A (g2483), .B (n_6938), .S0 (g5555), .Y (n_6940));
MX2X1 g60841(.A (g2486), .B (n_6938), .S0 (g7264), .Y (n_6939));
MX2X1 g60842(.A (g2489), .B (n_6938), .S0 (n_6611), .Y (n_6937));
XOR2X1 g60849(.A (n_297), .B (n_6867), .Y (n_6936));
NAND2X1 g60889(.A (n_7337), .B (n_6935), .Y (n_7330));
NOR2X1 g60890(.A (n_4946), .B (n_6782), .Y (n_6934));
NOR2X1 g60891(.A (n_4944), .B (n_6782), .Y (n_6933));
AOI21X1 g60897(.A0 (n_6692), .A1 (g_17483), .B0 (n_7142), .Y(n_6932));
AOI21X1 g60898(.A0 (n_6692), .A1 (g_17001), .B0 (n_7142), .Y(n_6931));
AOI21X1 g60919(.A0 (n_8420), .A1 (n_8573), .B0 (n_6688), .Y (n_6929));
INVX1 g60938(.A (n_8794), .Y (n_7125));
XOR2X1 g60986(.A (n_6465), .B (n_6693), .Y (n_7118));
OR2X1 g61015(.A (n_6765), .B (n_9060), .Y (n_7108));
OR2X1 g61017(.A (n_9366), .B (n_8472), .Y (n_7100));
OAI21X1 g61071(.A0 (n_5778), .A1 (n_8704), .B0 (n_6756), .Y (n_6926));
MX2X1 g61105(.A (g16355), .B (n_6881), .S0 (g6944), .Y (n_6925));
XOR2X1 g61125(.A (n_6464), .B (n_6678), .Y (n_7104));
NAND3X1 g61246(.A (n_6920), .B (n_6174), .C (n_6058), .Y (n_6975));
NAND3X1 g61253(.A (n_6759), .B (n_8725), .C (n_3812), .Y (n_6924));
INVX1 g61255(.A (n_8706), .Y (n_7038));
OR2X1 g61267(.A (n_5234), .B (n_6920), .Y (n_6921));
INVX1 g61284(.A (n_8678), .Y (n_6972));
NAND2X1 g61311(.A (n_6915), .B (n_6917), .Y (n_6918));
NAND2X1 g61312(.A (n_6915), .B (n_6914), .Y (n_6916));
NAND2X1 g61313(.A (n_6915), .B (g6447), .Y (n_6913));
OAI21X1 g61334(.A0 (n_6847), .A1 (n_9347), .B0 (n_6753), .Y (n_6911));
MX2X1 g61341(.A (g429), .B (n_6907), .S0 (n_6914), .Y (n_6909));
MX2X1 g61342(.A (g432), .B (n_6907), .S0 (g6447), .Y (n_6908));
MX2X1 g61343(.A (g435), .B (n_6907), .S0 (n_6917), .Y (n_6906));
XOR2X1 g61352(.A (n_5049), .B (n_6731), .Y (n_6905));
NAND2X1 g61388(.A (n_6902), .B (n_6914), .Y (n_6904));
NAND2X1 g61394(.A (n_6902), .B (n_6917), .Y (n_6903));
NAND2X1 g61395(.A (n_6902), .B (g6447), .Y (n_6901));
NAND3X1 g61416(.A (n_6899), .B (n_6430), .C (n_9192), .Y (n_6900));
MX2X1 g60530(.A (g1291), .B (n_6954), .S0 (g6750), .Y (n_6897));
OAI21X1 g60534(.A0 (n_6893), .A1 (n_6822), .B0 (n_908), .Y (n_6896));
OAI21X1 g61554(.A0 (n_6890), .A1 (n_6887), .B0 (n_6651), .Y (n_6895));
OAI21X1 g60535(.A0 (n_6893), .A1 (n_1596), .B0 (n_2091), .Y (n_6894));
OAI21X1 g60536(.A0 (n_6893), .A1 (n_3448), .B0 (n_3753), .Y (n_6892));
OAI21X1 g61560(.A0 (n_6890), .A1 (n_6884), .B0 (n_6650), .Y (n_6891));
OAI21X1 g61561(.A0 (n_6890), .A1 (n_6882), .B0 (n_6649), .Y (n_6889));
OAI21X1 g61562(.A0 (n_6885), .A1 (n_6887), .B0 (n_6648), .Y (n_6888));
OAI21X1 g61563(.A0 (n_6885), .A1 (n_6884), .B0 (n_6647), .Y (n_6886));
OAI21X1 g61564(.A0 (n_6885), .A1 (n_6882), .B0 (n_6646), .Y (n_6883));
CLKBUFX1 gbuf_d_368(.A(n_6721), .Y(d_out_368));
CLKBUFX1 gbuf_q_368(.A(q_in_368), .Y(g1115));
CLKBUFX1 gbuf_d_369(.A(n_6719), .Y(d_out_369));
CLKBUFX1 gbuf_q_369(.A(q_in_369), .Y(g1114));
CLKBUFX1 gbuf_d_370(.A(n_6722), .Y(d_out_370));
CLKBUFX1 gbuf_q_370(.A(q_in_370), .Y(g1113));
CLKBUFX1 gbuf_d_371(.A(n_6709), .Y(d_out_371));
CLKBUFX1 gbuf_q_371(.A(q_in_371), .Y(g1134));
CLKBUFX1 gbuf_d_372(.A(n_6708), .Y(d_out_372));
CLKBUFX1 gbuf_q_372(.A(q_in_372), .Y(g1135));
CLKBUFX1 gbuf_d_373(.A(n_6706), .Y(d_out_373));
CLKBUFX1 gbuf_q_373(.A(q_in_373), .Y(g1136));
CLKBUFX1 gbuf_d_374(.A(n_6705), .Y(d_out_374));
CLKBUFX1 gbuf_q_374(.A(q_in_374), .Y(g2522));
CLKBUFX1 gbuf_d_375(.A(n_6704), .Y(d_out_375));
CLKBUFX1 gbuf_q_375(.A(q_in_375), .Y(g2523));
CLKBUFX1 gbuf_d_376(.A(n_6702), .Y(d_out_376));
CLKBUFX1 gbuf_q_376(.A(q_in_376), .Y(g2524));
CLKBUFX1 gbuf_d_377(.A(n_6686), .Y(d_out_377));
CLKBUFX1 gbuf_q_377(.A(q_in_377), .Y(g3097));
CLKBUFX1 gbuf_d_378(.A(n_6685), .Y(d_out_378));
CLKBUFX1 gbuf_q_378(.A(q_in_378), .Y(g3098));
CLKBUFX1 gbuf_d_379(.A(n_6683), .Y(d_out_379));
CLKBUFX1 gbuf_q_379(.A(q_in_379), .Y(g3099));
CLKBUFX1 gbuf_d_380(.A(n_6674), .Y(d_out_380));
CLKBUFX1 gbuf_q_380(.A(q_in_380), .Y(g2418));
CLKBUFX1 gbuf_d_381(.A(n_6671), .Y(d_out_381));
CLKBUFX1 gbuf_q_381(.A(q_in_381), .Y(g2421));
CLKBUFX1 gbuf_d_382(.A(n_6748), .Y(d_out_382));
CLKBUFX1 gbuf_q_382(.A(q_in_382), .Y(g2448));
CLKBUFX1 gbuf_d_383(.A(n_6747), .Y(d_out_383));
CLKBUFX1 gbuf_q_383(.A(q_in_383), .Y(g2451));
CLKBUFX1 gbuf_d_384(.A(n_6745), .Y(d_out_384));
CLKBUFX1 gbuf_q_384(.A(q_in_384), .Y(g2459));
CLKBUFX1 gbuf_d_385(.A(n_6749), .Y(d_out_385));
CLKBUFX1 gbuf_q_385(.A(q_in_385), .Y(g2429));
CLKBUFX1 gbuf_d_386(.A(n_6743), .Y(d_out_386));
CLKBUFX1 gbuf_q_386(.A(q_in_386), .Y(g358));
CLKBUFX1 gbuf_d_387(.A(n_6740), .Y(d_out_387));
CLKBUFX1 gbuf_q_387(.A(q_in_387), .Y(g369));
CLKBUFX1 gbuf_d_388(.A(n_6742), .Y(d_out_388));
CLKBUFX1 gbuf_q_388(.A(q_in_388), .Y(g361));
CLKBUFX1 gbuf_d_389(.A(n_6739), .Y(d_out_389));
CLKBUFX1 gbuf_q_389(.A(q_in_389), .Y(g1739));
CLKBUFX1 gbuf_d_390(.A(n_6738), .Y(d_out_390));
CLKBUFX1 gbuf_q_390(.A(q_in_390), .Y(g1742));
CLKBUFX1 gbuf_d_391(.A(n_6736), .Y(d_out_391));
CLKBUFX1 gbuf_q_391(.A(q_in_391), .Y(g1750));
CLKBUFX1 gbuf_d_392(.A(n_6881), .Y(d_out_392));
CLKBUFX1 gbuf_q_392(.A(q_in_392), .Y(g16297));
XOR2X1 g61622(.A (n_6150), .B (n_6642), .Y (n_7027));
CLKBUFX1 gbuf_d_393(.A(n_6687), .Y(d_out_393));
CLKBUFX1 gbuf_q_393(.A(q_in_393), .Y(g1813));
CLKBUFX1 gbuf_d_394(.A(n_6711), .Y(d_out_394));
CLKBUFX1 gbuf_q_394(.A(q_in_394), .Y(g_14626));
AOI21X1 g60659(.A0 (n_6636), .A1 (n_8653), .B0 (n_9129), .Y (n_6880));
NAND3X1 g60683(.A (n_8281), .B (n_6785), .C (n_6726), .Y (n_6877));
MX2X1 g60826(.A (g1089), .B (n_6873), .S0 (n_5135), .Y (n_6875));
MX2X1 g60827(.A (g1091), .B (n_6873), .S0 (n_2969), .Y (n_6874));
MX2X1 g60828(.A (g1090), .B (n_6873), .S0 (n_2972), .Y (n_6872));
MX2X1 g60846(.A (g1095), .B (n_6869), .S0 (g5472), .Y (n_6871));
MX2X1 g60847(.A (g1098), .B (n_6869), .S0 (g6712), .Y (n_6870));
MX2X1 g60848(.A (n_6869), .B (g1101), .S0 (n_6420), .Y (n_6868));
CLKBUFX1 gbuf_d_395(.A(n_6710), .Y(d_out_395));
CLKBUFX1 gbuf_qn_395(.A(qn_in_395), .Y(g985));
OR2X1 g60892(.A (g_22538), .B (n_6867), .Y (n_7022));
NAND2X1 g60907(.A (n_6867), .B (n_6865), .Y (n_6866));
MX2X1 g60974(.A (n_6862), .B (g2501), .S0 (n_6612), .Y (n_6864));
MX2X1 g60975(.A (n_6862), .B (g2502), .S0 (n_6610), .Y (n_6863));
MX2X1 g60976(.A (n_6862), .B (g2503), .S0 (n_6607), .Y (n_6861));
INVX1 g61026(.A (n_6935), .Y (n_6860));
INVX1 g61039(.A (n_6859), .Y (n_6987));
NAND2X1 g61052(.A (n_8607), .B (n_7000), .Y (n_6855));
NAND2X1 g61060(.A (n_8471), .B (n_9256), .Y (n_6853));
INVX1 g61075(.A (n_6850), .Y (n_6851));
OAI21X1 g61081(.A0 (n_6826), .A1 (n_8863), .B0 (n_6698), .Y (n_6849));
OAI21X1 g61086(.A0 (n_6847), .A1 (n_6413), .B0 (n_6696), .Y (n_6848));
MX2X1 g61107(.A (n_6844), .B (g1828), .S0 (n_6600), .Y (n_6846));
MX2X1 g61108(.A (n_6844), .B (g1829), .S0 (n_6599), .Y (n_6845));
MX2X1 g61109(.A (n_6844), .B (g1830), .S0 (n_6597), .Y (n_6843));
XOR2X1 g62833(.A (n_4676), .B (n_6602), .Y (n_6841));
NAND4X1 g61257(.A (n_4677), .B (n_4610), .C (n_6522), .D (n_5610), .Y(n_6837));
INVX1 g61271(.A (n_9255), .Y (n_6836));
NAND2X1 g61328(.A (n_6830), .B (n_6832), .Y (n_6833));
NAND2X1 g61329(.A (n_6830), .B (g5511), .Y (n_6831));
NAND2X1 g61330(.A (n_6830), .B (g7014), .Y (n_6828));
OAI21X1 g61332(.A0 (n_6826), .A1 (n_5898), .B0 (n_6682), .Y (n_6827));
XOR2X1 g61353(.A (n_4228), .B (n_6755), .Y (n_6824));
OAI21X1 g60451(.A0 (n_6820), .A1 (n_6822), .B0 (n_850), .Y (n_6823));
OAI21X1 g60452(.A0 (n_6820), .A1 (n_1596), .B0 (n_2094), .Y (n_6821));
OAI21X1 g60453(.A0 (n_6820), .A1 (n_3448), .B0 (n_3752), .Y (n_6818));
NOR2X1 g61413(.A (n_6429), .B (n_6794), .Y (n_6974));
NAND3X1 g61417(.A (n_6731), .B (n_6321), .C (n_5234), .Y (n_6816));
NAND4X1 g61419(.A (n_6247), .B (n_6640), .C (n_5318), .D (n_4902), .Y(n_6815));
OAI21X1 g61530(.A0 (n_6812), .A1 (n_6809), .B0 (n_6497), .Y (n_6814));
OAI21X1 g61531(.A0 (n_6812), .A1 (n_6806), .B0 (n_6496), .Y (n_6813));
OAI21X1 g61532(.A0 (n_6812), .A1 (n_6804), .B0 (n_6495), .Y (n_6811));
OAI21X1 g61533(.A0 (n_6807), .A1 (n_6809), .B0 (n_6494), .Y (n_6810));
OAI21X1 g61534(.A0 (n_6807), .A1 (n_6806), .B0 (n_6493), .Y (n_6808));
OAI21X1 g61535(.A0 (n_6807), .A1 (n_6804), .B0 (n_6492), .Y (n_6805));
CLKBUFX1 gbuf_d_396(.A(n_6664), .Y(d_out_396));
CLKBUFX1 gbuf_q_396(.A(q_in_396), .Y(g2436));
CLKBUFX1 gbuf_d_397(.A(n_6634), .Y(d_out_397));
CLKBUFX1 gbuf_q_397(.A(q_in_397), .Y(g1967));
CLKBUFX1 gbuf_d_398(.A(n_6631), .Y(d_out_398));
CLKBUFX1 gbuf_q_398(.A(q_in_398), .Y(g1973));
CLKBUFX1 gbuf_d_399(.A(n_6633), .Y(d_out_399));
CLKBUFX1 gbuf_q_399(.A(q_in_399), .Y(g1970));
CLKBUFX1 gbuf_d_400(.A(n_6630), .Y(d_out_400));
CLKBUFX1 gbuf_q_400(.A(q_in_400), .Y(g1976));
CLKBUFX1 gbuf_d_401(.A(n_6629), .Y(d_out_401));
CLKBUFX1 gbuf_q_401(.A(q_in_401), .Y(g1979));
CLKBUFX1 gbuf_d_402(.A(n_6627), .Y(d_out_402));
CLKBUFX1 gbuf_q_402(.A(q_in_402), .Y(g1982));
CLKBUFX1 gbuf_d_403(.A(n_6622), .Y(d_out_403));
CLKBUFX1 gbuf_q_403(.A(q_in_403), .Y(g2516));
CLKBUFX1 gbuf_d_404(.A(n_6620), .Y(d_out_404));
CLKBUFX1 gbuf_q_404(.A(q_in_404), .Y(g2519));
CLKBUFX1 gbuf_d_405(.A(n_6623), .Y(d_out_405));
CLKBUFX1 gbuf_q_405(.A(q_in_405), .Y(g2513));
CLKBUFX1 gbuf_d_406(.A(n_6669), .Y(d_out_406));
CLKBUFX1 gbuf_q_406(.A(q_in_406), .Y(g1030));
CLKBUFX1 gbuf_d_407(.A(n_6666), .Y(d_out_407));
CLKBUFX1 gbuf_q_407(.A(q_in_407), .Y(g1041));
CLKBUFX1 gbuf_d_408(.A(n_6668), .Y(d_out_408));
CLKBUFX1 gbuf_q_408(.A(q_in_408), .Y(g1033));
CLKBUFX1 gbuf_d_409(.A(n_6665), .Y(d_out_409));
CLKBUFX1 gbuf_q_409(.A(q_in_409), .Y(g2433));
CLKBUFX1 gbuf_d_410(.A(n_6589), .Y(d_out_410));
CLKBUFX1 gbuf_q_410(.A(q_in_410), .Y(g_9172));
CLKBUFX1 gbuf_d_411(.A(n_6595), .Y(d_out_411));
CLKBUFX1 gbuf_q_411(.A(q_in_411), .Y(g_22536));
CLKBUFX1 gbuf_d_412(.A(n_6662), .Y(d_out_412));
CLKBUFX1 gbuf_q_412(.A(q_in_412), .Y(g2463));
CLKBUFX1 gbuf_d_413(.A(n_6661), .Y(d_out_413));
CLKBUFX1 gbuf_q_413(.A(q_in_413), .Y(g2466));
CLKBUFX1 gbuf_d_414(.A(n_6659), .Y(d_out_414));
CLKBUFX1 gbuf_q_414(.A(q_in_414), .Y(g2473));
MX2X1 g61590(.A (n_6801), .B (g388), .S0 (n_6809), .Y (n_6803));
MX2X1 g61591(.A (n_6801), .B (g391), .S0 (n_6806), .Y (n_6802));
MX2X1 g61592(.A (n_6801), .B (g398), .S0 (n_6804), .Y (n_6800));
MX2X1 g61614(.A (n_6797), .B (g1769), .S0 (n_6887), .Y (n_6799));
MX2X1 g61615(.A (n_6797), .B (g1772), .S0 (n_6884), .Y (n_6798));
MX2X1 g61616(.A (n_6797), .B (g1779), .S0 (n_6882), .Y (n_6796));
XOR2X1 g61619(.A (n_4827), .B (n_6730), .Y (n_6795));
NAND3X1 g61685(.A (n_7078), .B (n_6453), .C (n_6308), .Y (n_6902));
OAI22X1 g60614(.A0 (n_6567), .A1 (n_6947), .B0 (n_6946), .B1(n_4737), .Y (n_6965));
INVX1 g61776(.A (n_6794), .Y (n_6899));
MX2X1 g60696(.A (g1104), .B (n_6791), .S0 (g5472), .Y (n_6793));
MX2X1 g60697(.A (g1107), .B (n_6791), .S0 (g6712), .Y (n_6792));
MX2X1 g60698(.A (n_6791), .B (g1110), .S0 (n_6420), .Y (n_6790));
OAI22X1 g60710(.A0 (n_6550), .A1 (n_6947), .B0 (n_6946), .B1(n_5101), .Y (n_6959));
NAND3X1 g60797(.A (n_6543), .B (n_6545), .C (n_3959), .Y (n_6788));
AND2X1 g60804(.A (n_7155), .B (n_8281), .Y (n_6787));
AOI21X1 g60920(.A0 (n_8534), .A1 (n_6785), .B0 (n_6314), .Y (n_6786));
AOI21X1 g60960(.A0 (n_8960), .A1 (n_6785), .B0 (n_4927), .Y (n_6942));
CLKBUFX1 gbuf_d_415(.A(n_6606), .Y(d_out_415));
CLKBUFX1 gbuf_q_415(.A(q_in_415), .Y(g2444));
NOR2X1 g61021(.A (n_9366), .B (n_5712), .Y (n_6996));
NOR2X1 g61022(.A (n_5539), .B (n_9058), .Y (n_6999));
NOR2X1 g61027(.A (n_6692), .B (n_6442), .Y (n_6935));
INVX1 g61028(.A (n_6945), .Y (n_6782));
INVX1 g61040(.A (n_9418), .Y (n_6859));
INVX1 g61072(.A (n_8566), .Y (n_6778));
OAI21X1 g61076(.A0 (n_8667), .A1 (n_5141), .B0 (n_5331), .Y (n_6850));
MX2X1 g61089(.A (g1819), .B (n_6774), .S0 (g5511), .Y (n_6776));
MX2X1 g61090(.A (g1822), .B (n_6774), .S0 (n_3190), .Y (n_6775));
MX2X1 g61091(.A (g1825), .B (n_6774), .S0 (n_6832), .Y (n_6773));
AOI22X1 g62834(.A0 (n_5232), .A1 (n_8863), .B0 (n_6697), .B1(n_8862), .Y (n_6772));
AND2X1 g61244(.A (n_6560), .B (n_6594), .Y (n_6769));
INVX1 g61321(.A (n_8607), .Y (n_6765));
MX2X1 g61337(.A (g1816), .B (n_6761), .S0 (n_6832), .Y (n_6763));
MX2X1 g61347(.A (g1810), .B (n_6761), .S0 (g5511), .Y (n_6762));
NOR2X1 g61397(.A (n_6320), .B (n_6732), .Y (n_6920));
INVX1 g61406(.A (n_8598), .Y (n_6759));
NAND3X1 g61412(.A (n_6755), .B (n_6188), .C (n_5778), .Y (n_6756));
NAND4X1 g61414(.A (n_6120), .B (n_6563), .C (n_5133), .D (n_4901), .Y(n_6753));
AOI21X1 g61428(.A0 (n_6168), .A1 (n_6204), .B0 (n_6644), .Y (n_6752));
NAND2X1 g61502(.A (n_6657), .B (n_7094), .Y (n_6915));
OAI21X1 g61548(.A0 (n_6673), .A1 (n_6744), .B0 (n_6576), .Y (n_6749));
OAI21X1 g61549(.A0 (n_6746), .A1 (n_6672), .B0 (n_6575), .Y (n_6748));
OAI21X1 g61550(.A0 (n_6746), .A1 (n_6670), .B0 (n_6574), .Y (n_6747));
OAI21X1 g61551(.A0 (n_6746), .A1 (n_6744), .B0 (n_6573), .Y (n_6745));
MX2X1 g61567(.A (n_6741), .B (g358), .S0 (n_6809), .Y (n_6743));
MX2X1 g61568(.A (n_6741), .B (g361), .S0 (n_6806), .Y (n_6742));
MX2X1 g61569(.A (n_6741), .B (g369), .S0 (n_6804), .Y (n_6740));
MX2X1 g61573(.A (n_6737), .B (g1739), .S0 (n_6887), .Y (n_6739));
MX2X1 g61574(.A (n_6737), .B (g1742), .S0 (n_6884), .Y (n_6738));
MX2X1 g61575(.A (n_6737), .B (g1750), .S0 (n_6882), .Y (n_6736));
CLKBUFX1 gbuf_d_416(.A(n_6541), .Y(d_out_416));
CLKBUFX1 gbuf_q_416(.A(q_in_416), .Y(g1128));
CLKBUFX1 gbuf_d_417(.A(n_6511), .Y(d_out_417));
CLKBUFX1 gbuf_q_417(.A(q_in_417), .Y(g1063));
CLKBUFX1 gbuf_d_418(.A(n_6508), .Y(d_out_418));
CLKBUFX1 gbuf_q_418(.A(q_in_418), .Y(g1071));
CLKBUFX1 gbuf_d_419(.A(n_6513), .Y(d_out_419));
CLKBUFX1 gbuf_q_419(.A(q_in_419), .Y(g1060));
XOR2X1 g61583(.A (n_8730), .B (n_6475), .Y (n_6735));
CLKBUFX1 gbuf_d_420(.A(n_6519), .Y(d_out_420));
CLKBUFX1 gbuf_q_420(.A(q_in_420), .Y(g2120));
CLKBUFX1 gbuf_d_421(.A(n_6557), .Y(d_out_421));
CLKBUFX1 gbuf_q_421(.A(q_in_421), .Y(g3088));
CLKBUFX1 gbuf_d_422(.A(n_6556), .Y(d_out_422));
CLKBUFX1 gbuf_q_422(.A(q_in_422), .Y(g3155));
CLKBUFX1 gbuf_d_423(.A(n_6551), .Y(d_out_423));
CLKBUFX1 gbuf_q_423(.A(q_in_423), .Y(g3158));
CLKBUFX1 gbuf_d_424(.A(n_6555), .Y(d_out_424));
CLKBUFX1 gbuf_q_424(.A(q_in_424), .Y(g3161));
CLKBUFX1 gbuf_d_425(.A(n_6554), .Y(d_out_425));
CLKBUFX1 gbuf_q_425(.A(q_in_425), .Y(g3182));
CLKBUFX1 gbuf_d_426(.A(n_6552), .Y(d_out_426));
CLKBUFX1 gbuf_q_426(.A(q_in_426), .Y(g3185));
CLKBUFX1 gbuf_d_427(.A(n_6566), .Y(d_out_427));
CLKBUFX1 gbuf_q_427(.A(q_in_427), .Y(g1430));
CLKBUFX1 gbuf_d_428(.A(n_6538), .Y(d_out_428));
CLKBUFX1 gbuf_qn_428(.A(qn_in_428), .Y(g1836));
CLKBUFX1 gbuf_d_429(.A(n_6537), .Y(d_out_429));
CLKBUFX1 gbuf_qn_429(.A(qn_in_429), .Y(g1839));
CLKBUFX1 gbuf_d_430(.A(n_6535), .Y(d_out_430));
CLKBUFX1 gbuf_qn_430(.A(qn_in_430), .Y(g1842));
XOR2X1 g61618(.A (n_6100), .B (n_6656), .Y (n_6734));
CLKBUFX1 gbuf_d_431(.A(n_6539), .Y(d_out_431));
CLKBUFX1 gbuf_q_431(.A(q_in_431), .Y(g1131));
INVX1 g61755(.A (n_6732), .Y (n_6731));
CLKBUFX1 gbuf_d_432(.A(n_6542), .Y(d_out_432));
CLKBUFX1 gbuf_q_432(.A(q_in_432), .Y(g1125));
NAND2X2 g61777(.A (n_6186), .B (n_6730), .Y (n_6794));
XOR2X1 g61848(.A (n_6151), .B (n_6445), .Y (n_6907));
OAI22X1 g60709(.A0 (n_6458), .A1 (n_6947), .B0 (n_6946), .B1(n_7273), .Y (n_6954));
NAND2X1 g60812(.A (n_6547), .B (n_6191), .Y (n_6729));
NAND2X1 g60814(.A (n_6548), .B (n_6532), .Y (n_6728));
NAND2X1 g60903(.A (n_6534), .B (n_6053), .Y (n_6724));
OR2X1 g60923(.A (n_6526), .B (n_8843), .Y (n_6723));
MX2X1 g60968(.A (n_6720), .B (g1113), .S0 (n_6421), .Y (n_6722));
MX2X1 g60969(.A (n_6720), .B (g1115), .S0 (n_6416), .Y (n_6721));
MX2X1 g60970(.A (n_6720), .B (g1114), .S0 (n_6418), .Y (n_6719));
XOR2X1 g60985(.A (n_6106), .B (n_6425), .Y (n_6949));
AND2X1 g61014(.A (n_8420), .B (n_9021), .Y (n_6718));
AND2X1 g61016(.A (n_8548), .B (n_6713), .Y (n_6715));
OR2X1 g61019(.A (n_6712), .B (n_43), .Y (n_6867));
NOR2X1 g61030(.A (n_7228), .B (n_5929), .Y (n_6945));
NOR2X1 g61037(.A (n_6583), .B (n_7307), .Y (n_6711));
NAND2X1 g61063(.A (n_6521), .B (n_5757), .Y (n_6710));
MX2X1 g61114(.A (n_6707), .B (g1134), .S0 (n_6400), .Y (n_6709));
MX2X1 g61115(.A (n_6707), .B (g1135), .S0 (n_6399), .Y (n_6708));
MX2X1 g61116(.A (n_6707), .B (g1136), .S0 (n_6397), .Y (n_6706));
MX2X1 g61117(.A (n_6703), .B (g2522), .S0 (n_6394), .Y (n_6705));
MX2X1 g61118(.A (n_6703), .B (g2523), .S0 (n_6393), .Y (n_6704));
MX2X1 g61119(.A (n_6703), .B (g2524), .S0 (n_6391), .Y (n_6702));
XOR2X1 g61124(.A (n_6105), .B (n_6395), .Y (n_6938));
XOR2X1 g62830(.A (n_4678), .B (n_6413), .Y (n_6700));
NAND3X1 g61233(.A (n_6520), .B (n_5233), .C (n_6697), .Y (n_6698));
NAND4X1 g61254(.A (n_4679), .B (n_4432), .C (n_6311), .D (n_5412), .Y(n_6696));
AND2X1 g61280(.A (n_6466), .B (n_6518), .Y (n_6693));
INVX1 g61294(.A (n_6690), .Y (n_6691));
INVX1 g61297(.A (n_6688), .Y (n_6689));
OAI21X1 g61336(.A0 (n_6568), .A1 (n_3036), .B0 (n_3433), .Y (n_6687));
MX2X1 g61348(.A (g3097), .B (n_6684), .S0 (g8106), .Y (n_6686));
MX2X1 g61349(.A (g3098), .B (n_6684), .S0 (g8030), .Y (n_6685));
MX2X1 g61350(.A (g3099), .B (n_6684), .S0 (g3109), .Y (n_6683));
NAND4X1 g61380(.A (n_6581), .B (n_6470), .C (n_5742), .D (n_5827), .Y(n_6682));
NAND3X1 g61405(.A (n_8734), .B (n_4001), .C (n_3985), .Y (n_8210));
OR2X1 g61409(.A (n_6653), .B (n_8726), .Y (n_6680));
AOI21X1 g61427(.A0 (n_5738), .A1 (n_6189), .B0 (n_6570), .Y (n_6678));
NAND2X1 g61513(.A (n_6582), .B (n_7043), .Y (n_6830));
OAI21X1 g61539(.A0 (g_25348), .A1 (g_8090), .B0 (n_6561), .Y(n_6881));
OAI21X1 g61544(.A0 (n_6673), .A1 (n_6672), .B0 (n_6578), .Y (n_6674));
OAI21X1 g61547(.A0 (n_6673), .A1 (n_6670), .B0 (n_6577), .Y (n_6671));
OAI21X1 g61552(.A0 (n_6667), .A1 (n_6512), .B0 (n_6110), .Y (n_6669));
OAI21X1 g61565(.A0 (n_6667), .A1 (n_6509), .B0 (n_6109), .Y (n_6668));
OAI21X1 g61566(.A0 (n_6667), .A1 (n_6507), .B0 (n_6108), .Y (n_6666));
CLKBUFX1 gbuf_d_433(.A(n_6406), .Y(d_out_433));
CLKBUFX1 gbuf_q_433(.A(q_in_433), .Y(g2504));
MX2X1 g61570(.A (n_6663), .B (g2433), .S0 (n_6672), .Y (n_6665));
MX2X1 g61571(.A (n_6663), .B (g2436), .S0 (n_6670), .Y (n_6664));
CLKBUFX1 gbuf_d_434(.A(n_6407), .Y(d_out_434));
CLKBUFX1 gbuf_q_434(.A(q_in_434), .Y(g1122));
CLKBUFX1 gbuf_d_435(.A(n_6498), .Y(d_out_435));
CLKBUFX1 gbuf_qn_435(.A(qn_in_435), .Y(g2808));
CLKBUFX1 gbuf_d_436(.A(n_6505), .Y(d_out_436));
CLKBUFX1 gbuf_qn_436(.A(qn_in_436), .Y(g2809));
CLKBUFX1 gbuf_d_437(.A(n_6504), .Y(d_out_437));
CLKBUFX1 gbuf_qn_437(.A(qn_in_437), .Y(g2810));
CLKBUFX1 gbuf_d_438(.A(n_6502), .Y(d_out_438));
CLKBUFX1 gbuf_qn_438(.A(qn_in_438), .Y(g734));
CLKBUFX1 gbuf_d_439(.A(n_6501), .Y(d_out_439));
CLKBUFX1 gbuf_qn_439(.A(qn_in_439), .Y(g735));
CLKBUFX1 gbuf_d_440(.A(n_6499), .Y(d_out_440));
CLKBUFX1 gbuf_qn_440(.A(qn_in_440), .Y(g736));
CLKBUFX1 gbuf_d_441(.A(n_6456), .Y(d_out_441));
CLKBUFX1 gbuf_q_441(.A(q_in_441), .Y(g593));
CLKBUFX1 gbuf_d_442(.A(n_6457), .Y(d_out_442));
CLKBUFX1 gbuf_q_442(.A(q_in_442), .Y(g587));
CLKBUFX1 gbuf_d_443(.A(n_6454), .Y(d_out_443));
CLKBUFX1 gbuf_q_443(.A(q_in_443), .Y(g590));
CLKBUFX1 gbuf_d_444(.A(n_6412), .Y(d_out_444));
CLKBUFX1 gbuf_q_444(.A(q_in_444), .Y(g1116));
CLKBUFX1 gbuf_d_445(.A(n_6410), .Y(d_out_445));
CLKBUFX1 gbuf_q_445(.A(q_in_445), .Y(g1119));
CLKBUFX1 gbuf_d_446(.A(n_6405), .Y(d_out_446));
CLKBUFX1 gbuf_q_446(.A(q_in_446), .Y(g2507));
CLKBUFX1 gbuf_d_447(.A(n_6488), .Y(d_out_447));
CLKBUFX1 gbuf_q_447(.A(q_in_447), .Y(g1056));
CLKBUFX1 gbuf_d_448(.A(n_6485), .Y(d_out_448));
CLKBUFX1 gbuf_q_448(.A(q_in_448), .Y(g1048));
CLKBUFX1 gbuf_d_449(.A(n_6487), .Y(d_out_449));
CLKBUFX1 gbuf_q_449(.A(q_in_449), .Y(g1045));
CLKBUFX1 gbuf_d_450(.A(n_6684), .Y(d_out_450));
CLKBUFX1 gbuf_q_450(.A(q_in_450), .Y(g548));
CLKBUFX1 gbuf_d_451(.A(n_6460), .Y(d_out_451));
CLKBUFX1 gbuf_q_451(.A(q_in_451), .Y(g3179));
CLKBUFX1 gbuf_d_452(.A(n_6462), .Y(d_out_452));
CLKBUFX1 gbuf_q_452(.A(q_in_452), .Y(g3176));
CLKBUFX1 gbuf_d_453(.A(n_6463), .Y(d_out_453));
CLKBUFX1 gbuf_q_453(.A(q_in_453), .Y(g3173));
CLKBUFX1 gbuf_d_454(.A(n_6479), .Y(d_out_454));
CLKBUFX1 gbuf_q_454(.A(q_in_454), .Y(g2124));
CLKBUFX1 gbuf_d_455(.A(n_6439), .Y(d_out_455));
CLKBUFX1 gbuf_qn_455(.A(qn_in_455), .Y(g1846));
CLKBUFX1 gbuf_d_456(.A(n_6438), .Y(d_out_456));
CLKBUFX1 gbuf_qn_456(.A(qn_in_456), .Y(g1849));
CLKBUFX1 gbuf_d_457(.A(n_6437), .Y(d_out_457));
CLKBUFX1 gbuf_qn_457(.A(qn_in_457), .Y(g1852));
CLKBUFX1 gbuf_d_458(.A(n_6436), .Y(d_out_458));
CLKBUFX1 gbuf_qn_458(.A(qn_in_458), .Y(g2530));
CLKBUFX1 gbuf_d_459(.A(n_6435), .Y(d_out_459));
CLKBUFX1 gbuf_qn_459(.A(qn_in_459), .Y(g2533));
CLKBUFX1 gbuf_d_460(.A(n_6433), .Y(d_out_460));
CLKBUFX1 gbuf_qn_460(.A(qn_in_460), .Y(g2536));
MX2X1 g61605(.A (n_6660), .B (g2463), .S0 (n_6672), .Y (n_6662));
MX2X1 g61606(.A (n_6660), .B (g2466), .S0 (n_6670), .Y (n_6661));
MX2X1 g61607(.A (n_6660), .B (g2473), .S0 (n_6744), .Y (n_6659));
XOR2X1 g61617(.A (n_4825), .B (n_6579), .Y (n_6658));
NAND2X1 g61703(.A (n_6655), .B (n_6166), .Y (n_6657));
MX2X1 g60617(.A (n_6370), .B (n_4517), .S0 (n_6947), .Y (n_6820));
NAND2X2 g61756(.A (n_6062), .B (n_6656), .Y (n_6732));
NAND3X1 g61764(.A (n_6655), .B (n_6643), .C (n_6593), .Y (n_7094));
NAND3X1 g61770(.A (n_6475), .B (n_6300), .C (n_6653), .Y (n_6654));
INVX1 g61774(.A (n_6652), .Y (n_6755));
NAND2X1 g61789(.A (n_6887), .B (g1724), .Y (n_6651));
NAND2X1 g61790(.A (n_6884), .B (g1727), .Y (n_6650));
NAND2X1 g61791(.A (g1735), .B (n_6882), .Y (n_6649));
NAND2X1 g61792(.A (n_6887), .B (g1754), .Y (n_6648));
NAND2X1 g61793(.A (n_6884), .B (g1757), .Y (n_6647));
NAND2X1 g61794(.A (g1765), .B (n_6882), .Y (n_6646));
NAND2X1 g61799(.A (g2580), .B (g2581), .Y (n_6645));
AOI21X1 g61821(.A0 (n_6336), .A1 (n_6643), .B0 (n_6354), .Y (n_6644));
AOI22X1 g60715(.A0 (n_6361), .A1 (n_6946), .B0 (n_6947), .B1(n_3260), .Y (n_6893));
NAND2X1 g62155(.A (n_5715), .B (n_6641), .Y (n_6642));
NAND3X1 g62157(.A (n_6641), .B (n_5714), .C (n_6451), .Y (n_7078));
NAND4X1 g62213(.A (n_6638), .B (n_6251), .C (n_6243), .D (n_6140), .Y(n_6885));
NAND3X1 g62218(.A (n_6639), .B (n_6245), .C (n_6302), .Y (n_6807));
INVX1 g62244(.A (n_6562), .Y (n_6640));
NAND4X1 g62260(.A (n_6424), .B (n_6639), .C (n_6255), .D (n_6158), .Y(n_6812));
NAND4X1 g62272(.A (n_6402), .B (n_6638), .C (n_6253), .D (n_6270), .Y(n_6890));
NAND2X1 g60918(.A (n_4671), .B (n_8844), .Y (n_6636));
NOR2X1 g60924(.A (g996), .B (n_8844), .Y (n_6635));
MX2X1 g60940(.A (g1967), .B (n_6632), .S0 (g7052), .Y (n_6634));
MX2X1 g60941(.A (g1970), .B (n_6632), .S0 (g7194), .Y (n_6633));
MX2X1 g60942(.A (g1973), .B (n_6632), .S0 (n_6626), .Y (n_6631));
MX2X1 g60943(.A (g1976), .B (n_6628), .S0 (g7052), .Y (n_6630));
MX2X1 g60944(.A (g1979), .B (n_6628), .S0 (g7194), .Y (n_6629));
MX2X1 g60946(.A (g1982), .B (n_6628), .S0 (n_6626), .Y (n_6627));
OR2X1 g61012(.A (n_6427), .B (n_6546), .Y (n_6873));
INVX1 g61077(.A (n_6624), .Y (n_6625));
MX2X1 g61098(.A (g2513), .B (n_6621), .S0 (g5555), .Y (n_6623));
MX2X1 g61099(.A (g2516), .B (n_6621), .S0 (g7264), .Y (n_6622));
MX2X1 g61100(.A (g2519), .B (n_6621), .S0 (n_6611), .Y (n_6620));
XOR2X1 g61122(.A (n_5420), .B (n_6296), .Y (n_6869));
XOR2X1 g62808(.A (n_5463), .B (n_8863), .Y (n_6619));
OR2X1 g62963(.A (n_5163), .B (n_6602), .Y (n_6618));
INVX1 g61291(.A (n_7228), .Y (n_6692));
INVX1 g61295(.A (n_8655), .Y (n_6690));
INVX1 g61298(.A (n_8786), .Y (n_6688));
NAND2X1 g61324(.A (n_6609), .B (n_6611), .Y (n_6612));
NAND2X1 g61325(.A (n_6609), .B (g5555), .Y (n_6610));
NAND2X1 g61326(.A (n_6609), .B (n_2180), .Y (n_6607));
MX2X1 g61572(.A (n_6663), .B (g2444), .S0 (n_6744), .Y (n_6606));
NAND2X1 g61377(.A (n_6598), .B (n_6832), .Y (n_6600));
NAND2X1 g61378(.A (n_6598), .B (g5511), .Y (n_6599));
NAND2X1 g61379(.A (n_6598), .B (g7014), .Y (n_6597));
NOR2X1 g61391(.A (n_6484), .B (n_6565), .Y (n_6595));
NAND4X1 g61393(.A (n_6593), .B (n_6165), .C (n_6167), .D (n_6213), .Y(n_6594));
MX2X1 g63356(.A (n_4014), .B (n_4455), .S0 (n_9303), .Y (n_6592));
OAI22X1 g63363(.A0 (n_3985), .A1 (n_9303), .B0 (n_4223), .B1(n_9129), .Y (n_8266));
CLKBUFX1 gbuf_d_461(.A(n_6403), .Y(d_out_461));
CLKBUFX1 gbuf_q_461(.A(q_in_461), .Y(g2510));
AOI21X1 g61514(.A0 (n_6064), .A1 (n_5825), .B0 (n_6490), .Y (n_6589));
CLKBUFX1 gbuf_d_462(.A(n_6358), .Y(d_out_462));
CLKBUFX1 gbuf_q_462(.A(q_in_462), .Y(g599));
CLKBUFX1 gbuf_d_463(.A(n_6353), .Y(d_out_463));
CLKBUFX1 gbuf_q_463(.A(q_in_463), .Y(g1273));
CLKBUFX1 gbuf_d_464(.A(n_6351), .Y(d_out_464));
CLKBUFX1 gbuf_q_464(.A(q_in_464), .Y(g1276));
CLKBUFX1 gbuf_d_465(.A(n_6349), .Y(d_out_465));
CLKBUFX1 gbuf_q_465(.A(q_in_465), .Y(g1279));
CLKBUFX1 gbuf_d_466(.A(n_6345), .Y(d_out_466));
CLKBUFX1 gbuf_q_466(.A(q_in_466), .Y(g1288));
CLKBUFX1 gbuf_d_467(.A(n_6344), .Y(d_out_467));
CLKBUFX1 gbuf_q_467(.A(q_in_467), .Y(g2670));
CLKBUFX1 gbuf_d_468(.A(n_6341), .Y(d_out_468));
CLKBUFX1 gbuf_q_468(.A(q_in_468), .Y(g2676));
CLKBUFX1 gbuf_d_469(.A(n_6347), .Y(d_out_469));
CLKBUFX1 gbuf_q_469(.A(q_in_469), .Y(g1285));
CLKBUFX1 gbuf_d_470(.A(n_6287), .Y(d_out_470));
CLKBUFX1 gbuf_q_470(.A(q_in_470), .Y(g1956));
CLKBUFX1 gbuf_d_471(.A(n_6288), .Y(d_out_471));
CLKBUFX1 gbuf_q_471(.A(q_in_471), .Y(g1955));
XOR2X1 g61582(.A (g_14626), .B (n_6489), .Y (n_6583));
CLKBUFX1 gbuf_d_472(.A(n_6304), .Y(d_out_472));
CLKBUFX1 gbuf_q_472(.A(q_in_472), .Y(g_21690));
CLKBUFX1 gbuf_d_473(.A(n_6379), .Y(d_out_473));
CLKBUFX1 gbuf_q_473(.A(q_in_473), .Y(g1075));
CLKBUFX1 gbuf_d_474(.A(n_6376), .Y(d_out_474));
CLKBUFX1 gbuf_q_474(.A(q_in_474), .Y(g1085));
CLKBUFX1 gbuf_d_475(.A(n_6378), .Y(d_out_475));
CLKBUFX1 gbuf_q_475(.A(q_in_475), .Y(g1078));
CLKBUFX1 gbuf_d_476(.A(n_6371), .Y(d_out_476));
CLKBUFX1 gbuf_q_476(.A(q_in_476), .Y(g1435));
CLKBUFX1 gbuf_d_477(.A(n_6367), .Y(d_out_477));
CLKBUFX1 gbuf_q_477(.A(q_in_477), .Y(g_29227));
CLKBUFX1 gbuf_d_478(.A(n_6327), .Y(d_out_478));
CLKBUFX1 gbuf_qn_478(.A(qn_in_478), .Y(g465));
CLKBUFX1 gbuf_d_479(.A(n_6326), .Y(d_out_479));
CLKBUFX1 gbuf_qn_479(.A(qn_in_479), .Y(g468));
XOR2X1 g61620(.A (n_5555), .B (n_6234), .Y (n_6774));
NAND2X1 g61704(.A (g_14626), .B (n_6375), .Y (n_6712));
NAND2X1 g61721(.A (n_6572), .B (n_5736), .Y (n_6582));
NOR2X1 g61724(.A (n_6365), .B (n_6282), .Y (n_6581));
CLKBUFX1 gbuf_d_480(.A(n_6325), .Y(d_out_480));
CLKBUFX1 gbuf_qn_480(.A(qn_in_480), .Y(g471));
NAND2X2 g61775(.A (n_6579), .B (n_8236), .Y (n_6652));
NAND2X1 g61779(.A (n_6672), .B (g2418), .Y (n_6578));
NAND2X1 g61780(.A (n_6670), .B (g2421), .Y (n_6577));
NAND2X1 g61781(.A (g2429), .B (n_6744), .Y (n_6576));
NAND2X1 g61782(.A (n_6672), .B (g2448), .Y (n_6575));
NAND2X1 g61783(.A (n_6670), .B (g2451), .Y (n_6574));
NAND2X1 g61784(.A (g2459), .B (n_6744), .Y (n_6573));
NAND3X1 g61795(.A (n_6572), .B (n_6569), .C (n_6517), .Y (n_7043));
NAND2X1 g61796(.A (g1886), .B (g1887), .Y (n_6571));
AOI21X1 g61815(.A0 (n_6206), .A1 (n_6569), .B0 (n_6210), .Y (n_6570));
INVX1 g61851(.A (n_6568), .Y (n_6761));
NAND2X1 g60794(.A (n_6334), .B (n_6323), .Y (n_6567));
NOR2X1 g62145(.A (n_6303), .B (n_6565), .Y (n_6566));
INVX2 g62188(.A (n_6474), .Y (n_6730));
INVX1 g62241(.A (n_6469), .Y (n_6563));
NAND4X1 g62245(.A (n_4898), .B (n_5696), .C (n_6141), .D (n_5683), .Y(n_6562));
OAI21X1 g62264(.A0 (g16297), .A1 (g6642), .B0 (g_25348), .Y (n_6561));
NAND4X1 g62282(.A (n_6482), .B (n_6212), .C (n_6558), .D (n_6036), .Y(n_6560));
MX2X1 g62301(.A (g3088), .B (n_6553), .S0 (g3109), .Y (n_6557));
NAND2X1 g62302(.A (n_570), .B (n_6340), .Y (n_6556));
NAND2X1 g62303(.A (n_6337), .B (n_902), .Y (n_6555));
MX2X1 g62309(.A (g3182), .B (n_6553), .S0 (g8106), .Y (n_6554));
MX2X1 g62311(.A (g3185), .B (n_6553), .S0 (g8030), .Y (n_6552));
NAND2X1 g62319(.A (n_687), .B (n_6338), .Y (n_6551));
NAND2X1 g60905(.A (n_6324), .B (n_5888), .Y (n_6550));
XOR2X1 g60980(.A (n_5414), .B (n_6181), .Y (n_6791));
OAI21X1 g60989(.A0 (n_6332), .A1 (n_6533), .B0 (n_6333), .Y (n_6548));
AOI22X1 g62555(.A0 (n_6149), .A1 (n_5798), .B0 (n_6254), .B1(n_6170), .Y (n_6801));
OAI21X1 g60990(.A0 (n_6330), .A1 (n_6190), .B0 (n_6331), .Y (n_6547));
AOI22X1 g62562(.A0 (n_6145), .A1 (n_5796), .B0 (n_6252), .B1(n_6161), .Y (n_6797));
NAND2X1 g61053(.A (n_6544), .B (n_6726), .Y (n_6545));
OAI21X1 g61078(.A0 (n_9235), .A1 (n_4505), .B0 (n_6543), .Y (n_6624));
MX2X1 g61092(.A (g1125), .B (n_6540), .S0 (g5472), .Y (n_6542));
MX2X1 g61096(.A (g1128), .B (n_6540), .S0 (g6712), .Y (n_6541));
MX2X1 g61097(.A (n_6540), .B (g1131), .S0 (n_6420), .Y (n_6539));
CLKBUFX1 gbuf_d_481(.A(n_6348), .Y(d_out_481));
CLKBUFX1 gbuf_q_481(.A(q_in_481), .Y(g1282));
MX2X1 g62705(.A (n_376), .B (n_6012), .S0 (g8012), .Y (n_6538));
MX2X1 g62706(.A (n_372), .B (n_6012), .S0 (g8082), .Y (n_6537));
MX2X1 g62707(.A (n_6012), .B (n_349), .S0 (g1866), .Y (n_6535));
OAI21X1 g61110(.A0 (n_6533), .A1 (n_6532), .B0 (n_6315), .Y (n_6534));
CLKBUFX1 gbuf_d_482(.A(n_6343), .Y(d_out_482));
CLKBUFX1 gbuf_q_482(.A(q_in_482), .Y(g2673));
CLKBUFX1 gbuf_d_483(.A(n_6359), .Y(d_out_483));
CLKBUFX1 gbuf_q_483(.A(q_in_483), .Y(g596));
INVX1 g62831(.A (n_6530), .Y (n_6531));
OR2X1 g62962(.A (n_3997), .B (n_6144), .Y (n_6527));
INVX1 g61258(.A (n_6525), .Y (n_6785));
INVX1 g61259(.A (n_6525), .Y (n_6526));
CLKBUFX1 gbuf_d_484(.A(n_6356), .Y(d_out_484));
CLKBUFX1 gbuf_q_484(.A(q_in_484), .Y(g602));
NAND4X1 g61292(.A (n_8796), .B (n_30), .C (n_6381), .D (g559), .Y(n_7228));
NOR2X1 g63136(.A (n_9192), .B (n_6144), .Y (n_6522));
OAI21X1 g61333(.A0 (n_8887), .A1 (n_5136), .B0 (n_6305), .Y (n_6521));
NOR2X1 g61385(.A (n_6384), .B (n_5049), .Y (n_6520));
NOR2X1 g61403(.A (n_6380), .B (n_6478), .Y (n_6519));
NAND4X1 g61434(.A (n_6517), .B (n_5879), .C (n_5737), .D (n_6086), .Y(n_6518));
MX2X1 g63357(.A (n_9303), .B (n_9129), .S0 (n_3790), .Y (n_6516));
CLKBUFX1 gbuf_d_485(.A(n_6284), .Y(d_out_485));
CLKBUFX1 gbuf_q_485(.A(q_in_485), .Y(g1957));
OAI21X1 g61524(.A0 (n_6510), .A1 (n_6512), .B0 (n_6115), .Y (n_6513));
OAI21X1 g61525(.A0 (n_6510), .A1 (n_6509), .B0 (n_6114), .Y (n_6511));
OAI21X1 g61526(.A0 (n_6510), .A1 (n_6507), .B0 (n_6113), .Y (n_6508));
CLKBUFX1 gbuf_d_486(.A(n_6264), .Y(d_out_486));
CLKBUFX1 gbuf_qn_486(.A(qn_in_486), .Y(g1421));
CLKBUFX1 gbuf_d_487(.A(n_6263), .Y(d_out_487));
CLKBUFX1 gbuf_qn_487(.A(qn_in_487), .Y(g2114));
CLKBUFX1 gbuf_d_488(.A(n_6280), .Y(d_out_488));
CLKBUFX1 gbuf_q_488(.A(q_in_488), .Y(g1962));
CLKBUFX1 gbuf_d_489(.A(n_6278), .Y(d_out_489));
CLKBUFX1 gbuf_q_489(.A(q_in_489), .Y(g1963));
CLKBUFX1 gbuf_d_490(.A(n_6275), .Y(d_out_490));
CLKBUFX1 gbuf_q_490(.A(q_in_490), .Y(g1958));
CLKBUFX1 gbuf_d_491(.A(n_6273), .Y(d_out_491));
CLKBUFX1 gbuf_q_491(.A(q_in_491), .Y(g1959));
CLKBUFX1 gbuf_d_492(.A(n_6271), .Y(d_out_492));
CLKBUFX1 gbuf_q_492(.A(q_in_492), .Y(g1960));
CLKBUFX1 gbuf_d_493(.A(n_6238), .Y(d_out_493));
CLKBUFX1 gbuf_q_493(.A(q_in_493), .Y(g1874));
CLKBUFX1 gbuf_d_494(.A(n_6236), .Y(d_out_494));
CLKBUFX1 gbuf_q_494(.A(q_in_494), .Y(g1877));
CLKBUFX1 gbuf_d_495(.A(n_6223), .Y(d_out_495));
CLKBUFX1 gbuf_q_495(.A(q_in_495), .Y(g_27924));
CLKBUFX1 gbuf_d_496(.A(n_6222), .Y(d_out_496));
CLKBUFX1 gbuf_q_496(.A(q_in_496), .Y(g3084));
CLKBUFX1 gbuf_d_497(.A(n_6221), .Y(d_out_497));
CLKBUFX1 gbuf_q_497(.A(q_in_497), .Y(g3164));
CLKBUFX1 gbuf_d_498(.A(n_6217), .Y(d_out_498));
CLKBUFX1 gbuf_q_498(.A(q_in_498), .Y(g3210));
CLKBUFX1 gbuf_d_499(.A(n_6229), .Y(d_out_499));
CLKBUFX1 gbuf_q_499(.A(q_in_499), .Y(g1444));
CLKBUFX1 gbuf_d_500(.A(n_6228), .Y(d_out_500));
CLKBUFX1 gbuf_q_500(.A(q_in_500), .Y(g_25523));
CLKBUFX1 gbuf_d_501(.A(n_6226), .Y(d_out_501));
CLKBUFX1 gbuf_q_501(.A(q_in_501), .Y(g2129));
CLKBUFX1 gbuf_d_502(.A(n_6203), .Y(d_out_502));
CLKBUFX1 gbuf_qn_502(.A(qn_in_502), .Y(g2540));
CLKBUFX1 gbuf_d_503(.A(n_6202), .Y(d_out_503));
CLKBUFX1 gbuf_qn_503(.A(qn_in_503), .Y(g2543));
CLKBUFX1 gbuf_d_504(.A(n_6201), .Y(d_out_504));
CLKBUFX1 gbuf_qn_504(.A(qn_in_504), .Y(g2546));
CLKBUFX1 gbuf_d_505(.A(n_6200), .Y(d_out_505));
CLKBUFX1 gbuf_qn_505(.A(qn_in_505), .Y(g1858));
CLKBUFX1 gbuf_d_506(.A(n_6198), .Y(d_out_506));
CLKBUFX1 gbuf_q_506(.A(q_in_506), .Y(g1859));
CLKBUFX1 gbuf_d_507(.A(n_6197), .Y(d_out_507));
CLKBUFX1 gbuf_qn_507(.A(qn_in_507), .Y(g1860));
CLKBUFX1 gbuf_d_508(.A(n_6214), .Y(d_out_508));
CLKBUFX1 gbuf_q_508(.A(q_in_508), .Y(g1439));
CLKBUFX1 gbuf_d_509(.A(n_6196), .Y(d_out_509));
CLKBUFX1 gbuf_qn_509(.A(qn_in_509), .Y(g455));
CLKBUFX1 gbuf_d_510(.A(n_6195), .Y(d_out_510));
CLKBUFX1 gbuf_qn_510(.A(qn_in_510), .Y(g458));
OAI21X1 g60591(.A0 (n_6503), .A1 (n_1785), .B0 (n_1569), .Y (n_6505));
OAI21X1 g60592(.A0 (n_6503), .A1 (n_1979), .B0 (n_1679), .Y (n_6504));
CLKBUFX1 gbuf_d_511(.A(n_6260), .Y(d_out_511));
CLKBUFX1 gbuf_qn_511(.A(qn_in_511), .Y(g2115));
CLKBUFX1 gbuf_d_512(.A(n_6262), .Y(d_out_512));
CLKBUFX1 gbuf_qn_512(.A(qn_in_512), .Y(g2116));
OAI21X1 g60604(.A0 (n_6500), .A1 (n_3307), .B0 (n_2848), .Y (n_6502));
OAI21X1 g60605(.A0 (n_6500), .A1 (n_2201), .B0 (n_1817), .Y (n_6501));
OAI21X1 g60606(.A0 (n_6500), .A1 (n_2207), .B0 (n_1815), .Y (n_6499));
NAND3X1 g61684(.A (n_6844), .B (n_5939), .C (n_5877), .Y (n_6598));
OAI21X1 g60609(.A0 (n_6503), .A1 (n_3151), .B0 (n_2974), .Y (n_6498));
CLKBUFX1 gbuf_d_513(.A(n_6266), .Y(d_out_513));
CLKBUFX1 gbuf_qn_513(.A(qn_in_513), .Y(g1422));
NAND2X1 g61757(.A (n_6809), .B (g343), .Y (n_6497));
NAND2X1 g61758(.A (n_6806), .B (g346), .Y (n_6496));
NAND2X1 g61759(.A (g354), .B (n_6804), .Y (n_6495));
NAND2X1 g61760(.A (n_6809), .B (g373), .Y (n_6494));
NAND2X1 g61761(.A (n_6806), .B (g376), .Y (n_6493));
NAND2X1 g61762(.A (g384), .B (n_6804), .Y (n_6492));
NAND2X1 g61767(.A (n_6489), .B (n_6865), .Y (n_6490));
INVX1 g61772(.A (n_8796), .Y (n_6684));
CLKBUFX1 gbuf_d_514(.A(n_6267), .Y(d_out_514));
CLKBUFX1 gbuf_qn_514(.A(qn_in_514), .Y(g1420));
MX2X1 g61816(.A (n_6486), .B (g1056), .S0 (n_6507), .Y (n_6488));
MX2X1 g61817(.A (n_6486), .B (g1045), .S0 (n_6512), .Y (n_6487));
MX2X1 g61818(.A (n_6486), .B (g1048), .S0 (n_6509), .Y (n_6485));
XOR2X1 g61829(.A (g_22536), .B (n_6026), .Y (n_6484));
CLKBUFX1 gbuf_d_515(.A(n_6216), .Y(d_out_515));
CLKBUFX1 gbuf_q_515(.A(q_in_515), .Y(g3211));
XOR2X1 g61847(.A (n_4240), .B (n_6096), .Y (n_6483));
XOR2X1 g61852(.A (n_5556), .B (n_6074), .Y (n_6568));
CLKBUFX1 gbuf_d_516(.A(n_6220), .Y(d_out_516));
CLKBUFX1 gbuf_q_516(.A(q_in_516), .Y(g3170));
CLKBUFX1 gbuf_d_517(.A(n_6218), .Y(d_out_517));
CLKBUFX1 gbuf_q_517(.A(q_in_517), .Y(g3167));
OAI21X1 g62116(.A0 (n_6482), .A1 (n_6212), .B0 (n_6335), .Y (n_6655));
NAND3X1 g62137(.A (n_6159), .B (n_6033), .C (n_5570), .Y (n_6481));
NAND3X1 g62138(.A (n_8234), .B (n_6047), .C (n_5687), .Y (n_6480));
INVX2 g62142(.A (n_6373), .Y (n_6656));
NOR2X1 g62169(.A (n_6153), .B (n_6478), .Y (n_6479));
INVX1 g62185(.A (n_6476), .Y (n_6475));
NAND3X1 g62189(.A (n_6473), .B (n_6056), .C (n_5901), .Y (n_6474));
NAND3X1 g62197(.A (n_6467), .B (n_5969), .C (n_6027), .Y (n_6746));
NAND2X1 g62208(.A (n_6472), .B (g7014), .Y (n_6887));
NAND2X1 g62211(.A (n_6472), .B (n_6832), .Y (n_6884));
NAND2X1 g62212(.A (n_6472), .B (g5511), .Y (n_6882));
INVX1 g62220(.A (n_6366), .Y (n_6470));
NAND4X1 g62242(.A (n_4715), .B (n_5518), .C (n_6014), .D (n_5685), .Y(n_6469));
NAND4X1 g62269(.A (n_6162), .B (n_6467), .C (n_5980), .D (n_5997), .Y(n_6673));
NAND4X1 g62284(.A (n_6374), .B (n_6465), .C (n_6464), .D (n_5880), .Y(n_6466));
MX2X1 g62306(.A (g3173), .B (n_6461), .S0 (g8106), .Y (n_6463));
MX2X1 g62307(.A (g3176), .B (n_6461), .S0 (g8030), .Y (n_6462));
MX2X1 g62308(.A (g3179), .B (n_6461), .S0 (g3109), .Y (n_6460));
XOR2X1 g62315(.A (n_4244), .B (n_6473), .Y (n_6459));
CLKBUFX1 gbuf_d_518(.A(n_6163), .Y(d_out_518));
CLKBUFX1 gbuf_q_518(.A(q_in_518), .Y(g1961));
NAND2X1 g60925(.A (n_6192), .B (n_6042), .Y (n_6458));
CLKBUFX1 gbuf_d_519(.A(n_6553), .Y(d_out_519));
CLKBUFX1 gbuf_q_519(.A(q_in_519), .Y(g2580));
MX2X1 g60947(.A (g587), .B (n_6455), .S0 (g6485), .Y (n_6457));
MX2X1 g60948(.A (g593), .B (n_6455), .S0 (n_4601), .Y (n_6456));
MX2X1 g60949(.A (g590), .B (n_6455), .S0 (g6642), .Y (n_6454));
NOR2X1 g62442(.A (n_6152), .B (n_6452), .Y (n_6641));
NAND3X1 g62443(.A (n_5444), .B (n_6452), .C (n_6451), .Y (n_6453));
AND2X1 g61011(.A (n_8534), .B (n_6448), .Y (n_6450));
OAI21X1 g62598(.A0 (n_6307), .A1 (n_6452), .B0 (n_6451), .Y (n_6445));
NOR2X1 g61079(.A (n_6183), .B (n_6442), .Y (n_6443));
OR2X1 g61082(.A (n_6180), .B (n_6440), .Y (n_6441));
OAI21X1 g62689(.A0 (g1846), .A1 (g8012), .B0 (n_6173), .Y (n_6439));
OAI21X1 g62690(.A0 (g1849), .A1 (g8082), .B0 (n_6172), .Y (n_6438));
OAI21X1 g62691(.A0 (n_6969), .A1 (g1866), .B0 (n_1007), .Y (n_6437));
MX2X1 g62742(.A (n_370), .B (n_5854), .S0 (g8087), .Y (n_6436));
MX2X1 g62743(.A (n_363), .B (n_5854), .S0 (g8167), .Y (n_6435));
MX2X1 g62744(.A (n_5854), .B (n_339), .S0 (g2560), .Y (n_6433));
INVX1 g62820(.A (n_6431), .Y (n_6432));
INVX1 g62828(.A (n_6429), .Y (n_6430));
OAI22X1 g62832(.A0 (n_4230), .A1 (n_6144), .B0 (n_5162), .B1(n_6602), .Y (n_6530));
CLKBUFX1 gbuf_d_520(.A(n_6193), .Y(d_out_520));
CLKBUFX1 gbuf_qn_520(.A(qn_in_520), .Y(g461));
OR2X1 g62956(.A (n_4757), .B (n_5902), .Y (n_9570));
INVX1 g61248(.A (n_6544), .Y (n_6427));
NAND2X1 g61260(.A (n_9235), .B (n_8839), .Y (n_6525));
AND2X1 g61268(.A (n_6107), .B (n_6155), .Y (n_6425));
AND2X1 g63041(.A (n_6269), .B (n_6424), .Y (n_6741));
OR2X1 g61303(.A (n_6208), .B (n_6182), .Y (n_6423));
OR2X1 g61306(.A (n_6207), .B (n_6179), .Y (n_6422));
OR2X1 g61307(.A (n_6417), .B (n_6420), .Y (n_6421));
NAND3X1 g61308(.A (n_5562), .B (n_6328), .C (n_6553), .Y (n_6419));
OR2X1 g61309(.A (n_6417), .B (n_8305), .Y (n_6418));
OR2X1 g61310(.A (n_6417), .B (n_2343), .Y (n_6416));
OAI21X1 g61338(.A0 (n_6409), .A1 (n_8305), .B0 (n_1402), .Y (n_6412));
OAI21X1 g61339(.A0 (n_6409), .A1 (n_2343), .B0 (n_2705), .Y (n_6410));
OAI21X1 g61340(.A0 (n_6409), .A1 (n_6420), .B0 (n_5198), .Y (n_6407));
MX2X1 g61344(.A (g2504), .B (n_6404), .S0 (g5555), .Y (n_6406));
MX2X1 g61345(.A (g2507), .B (n_6404), .S0 (g7264), .Y (n_6405));
MX2X1 g61346(.A (g2510), .B (n_6404), .S0 (n_6611), .Y (n_6403));
AND2X1 g63189(.A (n_6268), .B (n_6402), .Y (n_6737));
NAND2X1 g61396(.A (n_6398), .B (n_3808), .Y (n_6400));
NAND2X1 g61398(.A (n_6398), .B (g5472), .Y (n_6399));
NAND2X1 g61399(.A (n_6398), .B (g6712), .Y (n_6397));
NOR2X1 g61410(.A (n_8837), .B (n_4501), .Y (n_6396));
NAND4X1 g61415(.A (n_8221), .B (n_5129), .C (n_5567), .D (n_8222), .Y(n_6616));
AOI21X1 g61418(.A0 (n_5356), .A1 (n_5750), .B0 (n_6241), .Y (n_6395));
NAND2X1 g61421(.A (n_6392), .B (n_6611), .Y (n_6394));
NAND2X1 g61422(.A (n_6392), .B (g5555), .Y (n_6393));
NAND2X1 g61423(.A (n_6392), .B (n_2180), .Y (n_6391));
NAND2X1 g61509(.A (n_6256), .B (n_6862), .Y (n_6609));
CLKBUFX1 gbuf_d_521(.A(n_6239), .Y(d_out_521));
CLKBUFX1 gbuf_q_521(.A(q_in_521), .Y(g1871));
CLKBUFX1 gbuf_d_522(.A(n_6093), .Y(d_out_522));
CLKBUFX1 gbuf_q_522(.A(q_in_522), .Y(g2661));
CLKBUFX1 gbuf_d_523(.A(n_6089), .Y(d_out_523));
CLKBUFX1 gbuf_q_523(.A(q_in_523), .Y(g2667));
CLKBUFX1 gbuf_d_524(.A(n_6011), .Y(d_out_524));
CLKBUFX1 gbuf_q_524(.A(q_in_524), .Y(g1262));
CLKBUFX1 gbuf_d_525(.A(n_6009), .Y(d_out_525));
CLKBUFX1 gbuf_q_525(.A(q_in_525), .Y(g1263));
CLKBUFX1 gbuf_d_526(.A(n_6013), .Y(d_out_526));
CLKBUFX1 gbuf_q_526(.A(q_in_526), .Y(g1261));
CLKBUFX1 gbuf_d_527(.A(n_6133), .Y(d_out_527));
CLKBUFX1 gbuf_q_527(.A(q_in_527), .Y(g1966));
CLKBUFX1 gbuf_d_528(.A(n_6104), .Y(d_out_528));
CLKBUFX1 gbuf_q_528(.A(q_in_528), .Y(g3091));
CLKBUFX1 gbuf_d_529(.A(n_6102), .Y(d_out_529));
CLKBUFX1 gbuf_q_529(.A(q_in_529), .Y(g3092));
CLKBUFX1 gbuf_d_530(.A(n_6112), .Y(d_out_530));
CLKBUFX1 gbuf_q_530(.A(q_in_530), .Y(g1453));
CLKBUFX1 gbuf_d_531(.A(n_6111), .Y(d_out_531));
CLKBUFX1 gbuf_q_531(.A(q_in_531), .Y(g2138));
CLKBUFX1 gbuf_d_532(.A(n_6098), .Y(d_out_532));
CLKBUFX1 gbuf_q_532(.A(q_in_532), .Y(g1448));
CLKBUFX1 gbuf_d_533(.A(n_6073), .Y(d_out_533));
CLKBUFX1 gbuf_qn_533(.A(qn_in_533), .Y(g477));
CLKBUFX1 gbuf_d_534(.A(n_6071), .Y(d_out_534));
CLKBUFX1 gbuf_q_534(.A(q_in_534), .Y(g478));
CLKBUFX1 gbuf_d_535(.A(n_6070), .Y(d_out_535));
CLKBUFX1 gbuf_qn_535(.A(qn_in_535), .Y(g479));
CLKBUFX1 gbuf_d_536(.A(n_6097), .Y(d_out_536));
CLKBUFX1 gbuf_q_536(.A(q_in_536), .Y(g2133));
CLKBUFX1 gbuf_d_537(.A(n_6067), .Y(d_out_537));
CLKBUFX1 gbuf_q_537(.A(q_in_537), .Y(g2553));
CLKBUFX1 gbuf_d_538(.A(n_6066), .Y(d_out_538));
CLKBUFX1 gbuf_qn_538(.A(qn_in_538), .Y(g2554));
CLKBUFX1 gbuf_d_539(.A(n_6118), .Y(d_out_539));
CLKBUFX1 gbuf_q_539(.A(q_in_539), .Y(g1867));
CLKBUFX1 gbuf_d_540(.A(n_6123), .Y(d_out_540));
CLKBUFX1 gbuf_q_540(.A(q_in_540), .Y(g1868));
CLKBUFX1 gbuf_d_541(.A(n_6131), .Y(d_out_541));
CLKBUFX1 gbuf_qn_541(.A(qn_in_541), .Y(g1869));
CLKBUFX1 gbuf_d_542(.A(n_6136), .Y(d_out_542));
CLKBUFX1 gbuf_q_542(.A(q_in_542), .Y(g486));
CLKBUFX1 gbuf_d_543(.A(n_6128), .Y(d_out_543));
CLKBUFX1 gbuf_q_543(.A(q_in_543), .Y(g487));
XOR2X1 g61623(.A (n_5154), .B (n_5950), .Y (n_6621));
NAND2X1 g61744(.A (n_6101), .B (n_6045), .Y (n_6384));
CLKBUFX1 gbuf_d_544(.A(n_6116), .Y(d_out_544));
CLKBUFX1 gbuf_q_544(.A(q_in_544), .Y(g1964));
XOR2X1 g61836(.A (g2120), .B (n_5865), .Y (n_6380));
MX2X1 g61844(.A (n_6377), .B (g1075), .S0 (n_6512), .Y (n_6379));
MX2X1 g61845(.A (n_6377), .B (g1078), .S0 (n_6509), .Y (n_6378));
MX2X1 g61846(.A (n_6377), .B (g1085), .S0 (n_6507), .Y (n_6376));
CLKBUFX1 gbuf_d_545(.A(n_6134), .Y(d_out_545));
CLKBUFX1 gbuf_q_545(.A(q_in_545), .Y(g1965));
CLKBUFX1 gbuf_d_546(.A(n_6103), .Y(d_out_546));
CLKBUFX1 gbuf_q_546(.A(q_in_546), .Y(g3093));
INVX1 g62105(.A (n_6489), .Y (n_6375));
OAI21X1 g62114(.A0 (n_6374), .A1 (n_6465), .B0 (n_6205), .Y (n_6572));
NAND3X1 g62143(.A (n_6372), .B (n_5907), .C (n_5748), .Y (n_6373));
NOR2X1 g62146(.A (n_6099), .B (n_6079), .Y (n_6371));
NAND2X1 g60813(.A (n_6078), .B (n_5559), .Y (n_6370));
INVX2 g62182(.A (n_9346), .Y (n_6579));
NAND3X1 g62186(.A (n_6096), .B (n_5726), .C (n_5551), .Y (n_6476));
NAND2X1 g62194(.A (n_6368), .B (g7264), .Y (n_6672));
NAND2X1 g62195(.A (n_6368), .B (n_6611), .Y (n_6670));
NAND2X1 g62196(.A (n_6368), .B (g5555), .Y (n_6744));
NOR2X1 g62206(.A (n_6028), .B (n_7307), .Y (n_6367));
NAND4X1 g62221(.A (n_6124), .B (n_5897), .C (n_5719), .D (n_5686), .Y(n_6366));
CLKBUFX1 gbuf_d_547(.A(n_6069), .Y(d_out_547));
CLKBUFX1 gbuf_qn_547(.A(qn_in_547), .Y(g2552));
NAND4X1 g62222(.A (n_4088), .B (n_6001), .C (n_5824), .D (n_5826), .Y(n_6365));
NAND4X1 g62230(.A (n_6083), .B (n_5051), .C (n_5234), .D (n_5232), .Y(n_6826));
NAND3X1 g62252(.A (n_6048), .B (n_5878), .C (n_5832), .Y (n_6363));
NAND4X1 g62270(.A (n_6034), .B (n_6232), .C (n_5821), .D (n_5843), .Y(n_6667));
XOR2X1 g62293(.A (n_8694), .B (n_6372), .Y (n_6362));
AOI21X1 g60930(.A0 (n_5893), .A1 (n_5891), .B0 (n_6077), .Y (n_6361));
CLKBUFX1 gbuf_d_548(.A(n_6461), .Y(d_out_548));
CLKBUFX1 gbuf_q_548(.A(q_in_548), .Y(g1886));
CLKBUFX1 gbuf_d_549(.A(n_6339), .Y(d_out_549));
CLKBUFX1 gbuf_qn_549(.A(qn_in_549), .Y(g_25348));
MX2X1 g60950(.A (g596), .B (n_6357), .S0 (g6485), .Y (n_6359));
MX2X1 g60951(.A (g599), .B (n_6357), .S0 (g6642), .Y (n_6358));
MX2X1 g60952(.A (g602), .B (n_6357), .S0 (n_4601), .Y (n_6356));
NAND2X1 g62440(.A (n_6052), .B (n_6451), .Y (n_6354));
MX2X1 g60954(.A (g1273), .B (n_6350), .S0 (g6750), .Y (n_6353));
MX2X1 g60955(.A (g1276), .B (n_6350), .S0 (g6944), .Y (n_6351));
MX2X1 g60956(.A (n_6350), .B (g1279), .S0 (n_3220), .Y (n_6349));
MX2X1 g60957(.A (g1282), .B (n_6346), .S0 (g6750), .Y (n_6348));
MX2X1 g60958(.A (g1285), .B (n_6346), .S0 (g6944), .Y (n_6347));
MX2X1 g60959(.A (n_6346), .B (g1288), .S0 (n_3220), .Y (n_6345));
MX2X1 g60965(.A (g2670), .B (n_6342), .S0 (g7302), .Y (n_6344));
MX2X1 g60966(.A (g2673), .B (n_6342), .S0 (g7390), .Y (n_6343));
MX2X1 g60967(.A (n_6342), .B (g2676), .S0 (n_3448), .Y (n_6341));
NAND2X1 g62513(.A (n_6339), .B (g8106), .Y (n_6340));
NAND2X1 g62514(.A (n_6339), .B (g8030), .Y (n_6338));
NAND2X1 g62519(.A (g3109), .B (n_6339), .Y (n_6337));
INVX1 g62520(.A (n_6335), .Y (n_6336));
OAI21X1 g60987(.A0 (n_6075), .A1 (n_6322), .B0 (n_6076), .Y (n_6334));
AOI22X1 g62559(.A0 (n_5863), .A1 (n_5465), .B0 (n_5979), .B1(n_5884), .Y (n_6660));
NAND2X1 g61033(.A (n_6332), .B (n_6054), .Y (n_6333));
NAND2X1 g61061(.A (n_6330), .B (n_6043), .Y (n_6331));
OAI21X1 g61083(.A0 (n_5561), .A1 (n_5749), .B0 (n_6328), .Y (n_6329));
OAI21X1 g62694(.A0 (g465), .A1 (g7909), .B0 (n_6041), .Y (n_6327));
OAI21X1 g62695(.A0 (g468), .A1 (g7956), .B0 (n_6040), .Y (n_6326));
OAI21X1 g62696(.A0 (n_5868), .A1 (g485), .B0 (n_1046), .Y (n_6325));
OAI21X1 g61120(.A0 (n_6323), .A1 (n_6322), .B0 (n_6044), .Y (n_6324));
CLKBUFX1 gbuf_d_550(.A(n_6092), .Y(d_out_550));
CLKBUFX1 gbuf_q_550(.A(q_in_550), .Y(g2664));
INVX1 g62818(.A (n_6320), .Y (n_6321));
OAI22X1 g62821(.A0 (n_9633), .A1 (n_8862), .B0 (n_9637), .B1(n_8861), .Y (n_6431));
INVX1 g62825(.A (n_8708), .Y (n_6319));
OAI22X1 g62829(.A0 (n_4610), .A1 (n_6185), .B0 (n_4433), .B1(n_5713), .Y (n_6429));
AND2X1 g61222(.A (n_6533), .B (n_6947), .Y (n_6632));
NOR2X1 g61223(.A (n_6332), .B (n_6946), .Y (n_6628));
OR2X1 g62957(.A (n_3994), .B (n_5857), .Y (n_6316));
NAND2X1 g61241(.A (n_6332), .B (n_6533), .Y (n_6315));
INVX1 g61249(.A (n_9111), .Y (n_6544));
INVX1 g61286(.A (n_8533), .Y (n_6314));
NOR2X1 g63131(.A (n_5778), .B (n_5857), .Y (n_6311));
NAND2X1 g63171(.A (n_6127), .B (g_20059), .Y (n_6310));
NAND3X1 g63244(.A (n_6307), .B (n_6150), .C (n_6451), .Y (n_6308));
CLKBUFX1 gbuf_d_551(.A(n_6137), .Y(d_out_551));
CLKBUFX1 gbuf_qn_551(.A(qn_in_551), .Y(g488));
NAND4X1 g61382(.A (n_5811), .B (n_5948), .C (n_4537), .D (n_4717), .Y(n_6305));
NOR2X1 g61404(.A (n_6117), .B (n_6227), .Y (n_6304));
XOR2X1 g63344(.A (g1430), .B (n_5965), .Y (n_6303));
AOI22X1 g63350(.A0 (n_5961), .A1 (n_6157), .B0 (n_6156), .B1(n_6148), .Y (n_6302));
INVX1 g63359(.A (n_6299), .Y (n_6300));
AOI21X1 g61456(.A0 (n_5617), .A1 (n_5379), .B0 (n_6119), .Y (n_6296));
NAND3X1 g61507(.A (n_5783), .B (n_5773), .C (n_8985), .Y (n_6289));
OAI21X1 g61527(.A0 (n_6286), .A1 (n_6274), .B0 (n_5983), .Y (n_6288));
OAI21X1 g61528(.A0 (n_6286), .A1 (n_6279), .B0 (n_5982), .Y (n_6287));
OAI21X1 g61529(.A0 (n_6286), .A1 (n_6276), .B0 (n_5981), .Y (n_6284));
INVX1 g63638(.A (n_6413), .Y (n_9627));
NAND2X1 g63768(.A (n_5803), .B (n_5964), .Y (n_6282));
MX2X1 g61577(.A (n_6277), .B (g1962), .S0 (n_6279), .Y (n_6280));
MX2X1 g61578(.A (n_6277), .B (g1963), .S0 (n_6276), .Y (n_6278));
CLKBUFX1 gbuf_d_552(.A(n_5856), .Y(d_out_552));
CLKBUFX1 gbuf_q_552(.A(q_in_552), .Y(g575));
CLKBUFX1 gbuf_d_553(.A(n_5853), .Y(d_out_553));
CLKBUFX1 gbuf_q_553(.A(q_in_553), .Y(g576));
CLKBUFX1 gbuf_d_554(.A(n_6007), .Y(d_out_554));
CLKBUFX1 gbuf_q_554(.A(q_in_554), .Y(g2649));
CLKBUFX1 gbuf_d_555(.A(n_6006), .Y(d_out_555));
CLKBUFX1 gbuf_q_555(.A(q_in_555), .Y(g2650));
CLKBUFX1 gbuf_d_556(.A(n_6004), .Y(d_out_556));
CLKBUFX1 gbuf_q_556(.A(q_in_556), .Y(g2651));
CLKBUFX1 gbuf_d_557(.A(n_5972), .Y(d_out_557));
CLKBUFX1 gbuf_q_557(.A(q_in_557), .Y(g581));
CLKBUFX1 gbuf_d_558(.A(n_5999), .Y(d_out_558));
CLKBUFX1 gbuf_q_558(.A(q_in_558), .Y(g583));
MX2X1 g61584(.A (n_6272), .B (g1958), .S0 (n_6274), .Y (n_6275));
CLKBUFX1 gbuf_d_559(.A(n_5994), .Y(d_out_559));
CLKBUFX1 gbuf_q_559(.A(q_in_559), .Y(g1264));
CLKBUFX1 gbuf_d_560(.A(n_5989), .Y(d_out_560));
CLKBUFX1 gbuf_q_560(.A(q_in_560), .Y(g1266));
MX2X1 g61585(.A (n_6272), .B (g1959), .S0 (n_6279), .Y (n_6273));
MX2X1 g61586(.A (n_6272), .B (g1960), .S0 (n_6276), .Y (n_6271));
CLKBUFX1 gbuf_d_561(.A(n_5943), .Y(d_out_561));
CLKBUFX1 gbuf_q_561(.A(q_in_561), .Y(g3094));
CLKBUFX1 gbuf_d_562(.A(n_5941), .Y(d_out_562));
CLKBUFX1 gbuf_q_562(.A(q_in_562), .Y(g3095));
CLKBUFX1 gbuf_d_563(.A(n_5957), .Y(d_out_563));
CLKBUFX1 gbuf_q_563(.A(q_in_563), .Y(g_21927));
CLKBUFX1 gbuf_d_564(.A(n_5956), .Y(d_out_564));
CLKBUFX1 gbuf_q_564(.A(q_in_564), .Y(g2147));
AOI22X1 g63895(.A0 (n_6250), .A1 (n_6139), .B0 (n_5800), .B1 (g3229),.Y (n_6270));
CLKBUFX1 gbuf_d_565(.A(n_5934), .Y(d_out_565));
CLKBUFX1 gbuf_q_565(.A(q_in_565), .Y(g2142));
AOI22X1 g63904(.A0 (n_5799), .A1 (n_5647), .B0 (n_5967), .B1(n_5798), .Y (n_6269));
CLKBUFX1 gbuf_d_566(.A(n_5874), .Y(d_out_566));
CLKBUFX1 gbuf_qn_566(.A(qn_in_566), .Y(g1152));
CLKBUFX1 gbuf_d_567(.A(n_5875), .Y(d_out_567));
CLKBUFX1 gbuf_qn_567(.A(qn_in_567), .Y(g1155));
CLKBUFX1 gbuf_d_568(.A(n_5872), .Y(d_out_568));
CLKBUFX1 gbuf_qn_568(.A(qn_in_568), .Y(g1158));
AOI22X1 g63913(.A0 (n_5797), .A1 (n_5644), .B0 (n_5966), .B1(n_5796), .Y (n_6268));
XOR2X1 g61621(.A (n_4441), .B (n_5782), .Y (n_6540));
OAI21X1 g60599(.A0 (n_6265), .A1 (n_2889), .B0 (n_2541), .Y (n_6267));
OAI21X1 g60601(.A0 (n_6265), .A1 (n_2160), .B0 (n_1830), .Y (n_6266));
OAI21X1 g60602(.A0 (n_6265), .A1 (n_2203), .B0 (n_1831), .Y (n_6264));
OAI21X1 g60603(.A0 (n_6261), .A1 (n_2840), .B0 (n_2526), .Y (n_6263));
CLKBUFX1 gbuf_d_569(.A(n_5992), .Y(d_out_569));
CLKBUFX1 gbuf_q_569(.A(q_in_569), .Y(g1265));
OAI21X1 g60607(.A0 (n_6261), .A1 (n_1804), .B0 (n_1545), .Y (n_6262));
OAI21X1 g60608(.A0 (n_6261), .A1 (n_1802), .B0 (n_1558), .Y (n_6260));
NAND3X1 g61686(.A (n_6707), .B (n_5761), .C (n_5352), .Y (n_6398));
NAND3X1 g61687(.A (n_6703), .B (n_5606), .C (n_5348), .Y (n_6392));
OR2X1 g61702(.A (n_8887), .B (n_9136), .Y (n_8211));
NAND2X1 g61714(.A (n_6246), .B (n_5354), .Y (n_6256));
NAND2X1 g64252(.A (n_5967), .B (n_6254), .Y (n_6255));
NAND2X1 g64259(.A (n_5966), .B (n_6252), .Y (n_6253));
NAND2X1 g64260(.A (n_5962), .B (n_6250), .Y (n_6251));
NOR2X1 g61785(.A (n_5775), .B (n_6008), .Y (n_6247));
NAND3X1 g61786(.A (n_6246), .B (n_6240), .C (n_6154), .Y (n_6862));
NAND3X1 g64429(.A (n_5647), .B (n_5967), .C (g3229), .Y (n_6245));
NAND3X1 g64442(.A (n_5644), .B (n_5966), .C (g3229), .Y (n_6243));
AOI21X1 g61814(.A0 (n_5756), .A1 (n_6240), .B0 (n_5927), .Y (n_6241));
MX2X1 g61826(.A (g1871), .B (n_6237), .S0 (g7052), .Y (n_6239));
MX2X1 g61827(.A (g1874), .B (n_6237), .S0 (g7194), .Y (n_6238));
MX2X1 g61828(.A (g1877), .B (n_6237), .S0 (n_6626), .Y (n_6236));
NAND2X1 g62106(.A (n_6063), .B (g_9172), .Y (n_6489));
NAND2X1 g62117(.A (n_5723), .B (n_6233), .Y (n_6234));
NAND3X1 g62119(.A (n_6233), .B (n_5722), .C (n_6209), .Y (n_6844));
NAND4X1 g62120(.A (n_6232), .B (n_5681), .C (n_5679), .D (n_5548), .Y(n_6510));
NAND2X1 g62130(.A (n_6231), .B (n_6914), .Y (n_6804));
CLKBUFX1 gbuf_d_570(.A(n_6000), .Y(d_out_570));
CLKBUFX1 gbuf_q_570(.A(q_in_570), .Y(g582));
NOR2X1 g62147(.A (n_5940), .B (n_5876), .Y (n_6229));
NAND2X1 g62151(.A (n_6231), .B (g6447), .Y (n_6809));
NAND2X1 g62153(.A (n_6231), .B (n_6917), .Y (n_6806));
NOR2X1 g62164(.A (n_5870), .B (n_6227), .Y (n_6228));
NOR2X1 g62170(.A (n_5935), .B (n_5917), .Y (n_6226));
AOI21X1 g62285(.A0 (n_5435), .A1 (n_28), .B0 (n_5933), .Y (n_6223));
NAND2X1 g62297(.A (n_5919), .B (n_879), .Y (n_6222));
MX2X1 g62304(.A (g3164), .B (n_6219), .S0 (g8106), .Y (n_6221));
MX2X1 g62305(.A (g3170), .B (n_6219), .S0 (g3109), .Y (n_6220));
MX2X1 g62310(.A (g3167), .B (n_6219), .S0 (g8030), .Y (n_6218));
NAND2X1 g62312(.A (n_602), .B (n_5926), .Y (n_6217));
NAND2X1 g62313(.A (n_713), .B (n_5921), .Y (n_6216));
XOR2X1 g62316(.A (n_4900), .B (n_9345), .Y (n_6215));
NOR2X1 g62435(.A (n_5889), .B (n_6565), .Y (n_6214));
NAND3X1 g62441(.A (n_6212), .B (n_6643), .C (n_5717), .Y (n_6213));
NAND2X1 g62489(.A (n_5900), .B (n_6209), .Y (n_6210));
CLKBUFX1 gbuf_d_571(.A(n_5942), .Y(d_out_571));
CLKBUFX1 gbuf_q_571(.A(q_in_571), .Y(g3096));
OR2X1 g62506(.A (n_6442), .B (n_5913), .Y (n_6208));
OR2X1 g62509(.A (n_6440), .B (g1880), .Y (n_6207));
NAND3X1 g62521(.A (n_6482), .B (n_6212), .C (n_5717), .Y (n_6335));
INVX1 g62539(.A (n_6205), .Y (n_6206));
AOI21X1 g62560(.A0 (n_920), .A1 (n_6037), .B0 (n_6012), .Y (n_6472));
MX2X1 g62692(.A (n_6051), .B (n_5717), .S0 (n_6212), .Y (n_6204));
OAI21X1 g62698(.A0 (g2540), .A1 (g8087), .B0 (n_5883), .Y (n_6203));
OAI21X1 g62699(.A0 (g2543), .A1 (g8167), .B0 (n_5882), .Y (n_6202));
OAI21X1 g62700(.A0 (n_9347), .A1 (g2560), .B0 (n_1043), .Y (n_6201));
MX2X1 g62708(.A (n_4419), .B (n_6199), .S0 (g8012), .Y (n_6200));
MX2X1 g62709(.A (g1859), .B (n_6199), .S0 (g8082), .Y (n_6198));
MX2X1 g62710(.A (n_6199), .B (n_1093), .S0 (g1866), .Y (n_6197));
MX2X1 g62711(.A (n_378), .B (n_5545), .S0 (g7909), .Y (n_6196));
MX2X1 g62712(.A (n_348), .B (n_5545), .S0 (g7956), .Y (n_6195));
MX2X1 g62713(.A (n_5545), .B (n_367), .S0 (g485), .Y (n_6193));
OAI21X1 g61121(.A0 (n_6191), .A1 (n_6190), .B0 (n_5894), .Y (n_6192));
AOI21X1 g62748(.A0 (n_6465), .A1 (n_5138), .B0 (n_5533), .Y (n_6189));
OAI22X1 g62819(.A0 (n_8995), .A1 (n_8862), .B0 (n_5049), .B1(n_8861), .Y (n_6320));
INVX1 g62823(.A (n_6187), .Y (n_6188));
MX2X1 g62827(.A (n_4615), .B (n_4827), .S0 (n_6185), .Y (n_6186));
NOR2X1 g61232(.A (n_6182), .B (n_5929), .Y (n_6183));
AND2X1 g61235(.A (n_5422), .B (n_5871), .Y (n_6181));
NOR2X1 g61236(.A (n_6179), .B (g1880), .Y (n_6180));
OR2X1 g62961(.A (n_9192), .B (n_6602), .Y (n_6177));
OR2X1 g62965(.A (n_5234), .B (n_8863), .Y (n_6174));
NAND2X1 g62980(.A (n_6171), .B (g8012), .Y (n_6173));
NAND2X1 g62981(.A (n_6171), .B (g8082), .Y (n_6172));
NAND3X1 g63040(.A (n_5628), .B (n_6170), .C (g3229), .Y (n_6639));
AND2X1 g63046(.A (n_6167), .B (n_6166), .Y (n_6168));
OAI21X1 g63048(.A0 (n_6482), .A1 (n_6643), .B0 (n_5037), .Y (n_6165));
OR2X1 g61305(.A (n_5925), .B (n_5905), .Y (n_6164));
CLKBUFX1 gbuf_d_572(.A(n_5850), .Y(d_out_572));
CLKBUFX1 gbuf_q_572(.A(q_in_572), .Y(g577));
MX2X1 g61576(.A (n_6277), .B (g1961), .S0 (n_6274), .Y (n_6163));
AND2X1 g63164(.A (n_5984), .B (n_6162), .Y (n_6663));
NAND3X1 g63185(.A (n_5625), .B (n_6161), .C (g3229), .Y (n_6638));
AOI22X1 g63833(.A0 (n_6157), .A1 (n_6156), .B0 (n_5801), .B1 (g3229),.Y (n_6158));
NAND4X1 g61433(.A (n_6154), .B (n_5576), .C (n_5355), .D (n_5609), .Y(n_6155));
XOR2X1 g63346(.A (g2124), .B (n_5805), .Y (n_6153));
MX2X1 g63353(.A (n_6019), .B (n_6151), .S0 (n_6150), .Y (n_6152));
NAND2X1 g63360(.A (n_5725), .B (n_5867), .Y (n_6299));
AND2X1 g63465(.A (n_6148), .B (g3229), .Y (n_6149));
AOI21X1 g61500(.A0 (n_5819), .A1 (n_5615), .B0 (n_5976), .Y (n_6417));
AND2X1 g63492(.A (n_6138), .B (g3229), .Y (n_6145));
INVX2 g63639(.A (n_5857), .Y (n_6413));
NAND2X1 g63721(.A (n_6139), .B (n_6138), .Y (n_6140));
MX2X1 g63835(.A (n_5444), .B (n_1101), .S0 (g485), .Y (n_6137));
MX2X1 g63837(.A (g486), .B (n_5444), .S0 (g7909), .Y (n_6136));
CLKBUFX1 gbuf_d_573(.A(n_5706), .Y(d_out_573));
CLKBUFX1 gbuf_q_573(.A(q_in_573), .Y(g1269));
CLKBUFX1 gbuf_d_574(.A(n_5822), .Y(d_out_574));
CLKBUFX1 gbuf_q_574(.A(q_in_574), .Y(g578));
CLKBUFX1 gbuf_d_575(.A(n_5842), .Y(d_out_575));
CLKBUFX1 gbuf_q_575(.A(q_in_575), .Y(g580));
CLKBUFX1 gbuf_d_576(.A(n_5766), .Y(d_out_576));
CLKBUFX1 gbuf_q_576(.A(q_in_576), .Y(g3085));
CLKBUFX1 gbuf_d_577(.A(n_5765), .Y(d_out_577));
CLKBUFX1 gbuf_q_577(.A(q_in_577), .Y(g3086));
CLKBUFX1 gbuf_d_578(.A(n_5785), .Y(d_out_578));
CLKBUFX1 gbuf_q_578(.A(q_in_578), .Y(g_18173));
MX2X1 g61588(.A (n_6132), .B (g1965), .S0 (n_6279), .Y (n_6134));
MX2X1 g61589(.A (n_6132), .B (g1966), .S0 (n_6276), .Y (n_6133));
CLKBUFX1 gbuf_d_579(.A(n_5760), .Y(d_out_579));
CLKBUFX1 gbuf_q_579(.A(q_in_579), .Y(g_26529));
CLKBUFX1 gbuf_d_580(.A(n_5759), .Y(d_out_580));
CLKBUFX1 gbuf_q_580(.A(q_in_580), .Y(g_15687));
CLKBUFX1 gbuf_d_581(.A(n_5754), .Y(d_out_581));
CLKBUFX1 gbuf_q_581(.A(q_in_581), .Y(g_14677));
CLKBUFX1 gbuf_d_582(.A(n_5753), .Y(d_out_582));
CLKBUFX1 gbuf_q_582(.A(q_in_582), .Y(g_29207));
CLKBUFX1 gbuf_d_583(.A(n_5751), .Y(d_out_583));
CLKBUFX1 gbuf_q_583(.A(q_in_583), .Y(g_24922));
CLKBUFX1 gbuf_d_584(.A(n_5728), .Y(d_out_584));
CLKBUFX1 gbuf_qn_584(.A(qn_in_584), .Y(g1142));
CLKBUFX1 gbuf_d_585(.A(n_5731), .Y(d_out_585));
CLKBUFX1 gbuf_qn_585(.A(qn_in_585), .Y(g1145));
CLKBUFX1 gbuf_d_586(.A(n_5847), .Y(d_out_586));
CLKBUFX1 gbuf_q_586(.A(q_in_586), .Y(g2561));
CLKBUFX1 gbuf_d_587(.A(n_5810), .Y(d_out_587));
CLKBUFX1 gbuf_q_587(.A(q_in_587), .Y(g2562));
CLKBUFX1 gbuf_d_588(.A(n_5846), .Y(d_out_588));
CLKBUFX1 gbuf_qn_588(.A(qn_in_588), .Y(g2563));
CLKBUFX1 gbuf_d_589(.A(n_5837), .Y(d_out_589));
CLKBUFX1 gbuf_qn_589(.A(qn_in_589), .Y(g464));
CLKBUFX1 gbuf_d_590(.A(n_5834), .Y(d_out_590));
CLKBUFX1 gbuf_q_590(.A(q_in_590), .Y(g480));
CLKBUFX1 gbuf_d_591(.A(n_5836), .Y(d_out_591));
CLKBUFX1 gbuf_q_591(.A(q_in_591), .Y(g484));
MX2X1 g63829(.A (n_5445), .B (n_1136), .S0 (g1866), .Y (n_6131));
MX2X1 g63838(.A (g487), .B (n_5444), .S0 (g7956), .Y (n_6128));
AND2X1 g63811(.A (g_7108), .B (n_2874), .Y (n_6127));
XOR2X1 g64082(.A (g_27975), .B (n_6697), .Y (n_6124));
MX2X1 g63828(.A (g1868), .B (n_5445), .S0 (g8082), .Y (n_6123));
NOR2X1 g61778(.A (n_5777), .B (n_5697), .Y (n_6120));
CLKBUFX1 gbuf_d_592(.A(n_5844), .Y(d_out_592));
CLKBUFX1 gbuf_q_592(.A(q_in_592), .Y(g579));
AOI21X1 g61802(.A0 (n_5210), .A1 (n_5818), .B0 (n_5788), .Y (n_6119));
MX2X1 g63827(.A (g1867), .B (n_5445), .S0 (g8012), .Y (n_6118));
NAND3X1 g64461(.A (n_6250), .B (n_5768), .C (g3229), .Y (n_6402));
NAND3X1 g64464(.A (n_6157), .B (n_5770), .C (g3229), .Y (n_6424));
XOR2X1 g61835(.A (g_21690), .B (n_5553), .Y (n_6117));
XOR2X1 g61849(.A (n_4953), .B (n_5595), .Y (n_6409));
XOR2X1 g61850(.A (n_5155), .B (n_5592), .Y (n_6404));
MX2X1 g61587(.A (n_6132), .B (g1964), .S0 (n_6274), .Y (n_6116));
NAND3X1 g60759(.A (n_3108), .B (n_2815), .C (n_5594), .Y (n_6500));
NAND3X1 g60760(.A (n_2956), .B (n_2672), .C (n_5593), .Y (n_6503));
NAND2X1 g62118(.A (n_6512), .B (g1060), .Y (n_6115));
NAND2X1 g62121(.A (n_6509), .B (g1063), .Y (n_6114));
NAND2X1 g62122(.A (g1071), .B (n_6507), .Y (n_6113));
NOR2X1 g62150(.A (n_5762), .B (n_5527), .Y (n_6112));
NOR2X1 g62171(.A (n_5763), .B (n_5732), .Y (n_6111));
NAND2X1 g62205(.A (n_6512), .B (g1030), .Y (n_6110));
NAND2X1 g62215(.A (n_6509), .B (g1033), .Y (n_6109));
NAND2X1 g62216(.A (g1041), .B (n_6507), .Y (n_6108));
NAND4X1 g62283(.A (n_5958), .B (n_6106), .C (n_6105), .D (n_5353), .Y(n_6107));
MX2X1 g62294(.A (g3091), .B (g1939), .S0 (g8106), .Y (n_6104));
MX2X1 g62314(.A (g3093), .B (g1939), .S0 (g3109), .Y (n_6103));
MX2X1 g62317(.A (g3092), .B (g1939), .S0 (g8030), .Y (n_6102));
CLKBUFX1 gbuf_d_593(.A(n_6219), .Y(d_out_593));
CLKBUFX1 gbuf_qn_593(.A(qn_in_593), .Y(g1192));
NOR2X1 g62427(.A (n_8693), .B (n_6100), .Y (n_6101));
OR2X1 g62434(.A (n_6025), .B (n_6565), .Y (n_6099));
NOR2X1 g62436(.A (n_5804), .B (n_6565), .Y (n_6098));
NOR2X1 g62459(.A (n_5848), .B (n_6478), .Y (n_6097));
INVX2 g62464(.A (n_6094), .Y (n_6096));
MX2X1 g60962(.A (g2661), .B (n_6091), .S0 (g7302), .Y (n_6093));
MX2X1 g60963(.A (g2664), .B (n_6091), .S0 (g7390), .Y (n_6092));
MX2X1 g60964(.A (n_6091), .B (g2667), .S0 (n_3448), .Y (n_6089));
NAND3X1 g62493(.A (n_6465), .B (n_6569), .C (n_5331), .Y (n_6086));
NOR2X1 g62498(.A (n_5489), .B (n_8693), .Y (n_6083));
OR2X1 g62510(.A (g1924), .B (g1880), .Y (n_6080));
AOI21X1 g62515(.A0 (n_5651), .A1 (g1439), .B0 (g1435), .Y (n_6079));
NAND3X1 g62540(.A (n_6374), .B (n_6465), .C (n_5331), .Y (n_6205));
MX2X1 g60988(.A (n_5892), .B (n_6077), .S0 (n_5908), .Y (n_6078));
AOI21X1 g62557(.A0 (n_3873), .A1 (n_9347), .B0 (n_5854), .Y (n_6368));
NAND2X1 g61036(.A (n_6075), .B (n_5887), .Y (n_6076));
CLKBUFX1 gbuf_d_594(.A(n_5764), .Y(d_out_594));
CLKBUFX1 gbuf_q_594(.A(q_in_594), .Y(g3087));
AOI21X1 g62688(.A0 (n_5704), .A1 (n_5703), .B0 (n_5531), .Y (n_6074));
MX2X1 g62714(.A (n_3971), .B (n_6072), .S0 (g7909), .Y (n_6073));
MX2X1 g62715(.A (g478), .B (n_6072), .S0 (g7956), .Y (n_6071));
MX2X1 g62716(.A (n_6072), .B (n_1141), .S0 (g485), .Y (n_6070));
MX2X1 g62745(.A (n_3978), .B (n_6068), .S0 (g8087), .Y (n_6069));
MX2X1 g62746(.A (g2553), .B (n_6068), .S0 (g8167), .Y (n_6067));
MX2X1 g62747(.A (n_6068), .B (n_845), .S0 (g2560), .Y (n_6066));
XOR2X1 g62789(.A (n_8411), .B (n_5325), .Y (n_6065));
INVX1 g62813(.A (n_6063), .Y (n_6064));
MX2X1 g62817(.A (n_5307), .B (n_6100), .S0 (n_8862), .Y (n_6062));
OAI22X1 g62824(.A0 (n_4432), .A1 (n_5915), .B0 (n_4228), .B1(n_5902), .Y (n_6187));
AND2X1 g61224(.A (n_6322), .B (n_6947), .Y (n_6455));
OR2X1 g62951(.A (n_5053), .B (n_8862), .Y (n_6058));
NAND2X1 g62958(.A (n_4004), .B (n_5335), .Y (n_6056));
OR2X1 g62960(.A (n_9188), .B (n_6185), .Y (n_6055));
INVX1 g61242(.A (n_6053), .Y (n_6054));
AOI21X1 g62969(.A0 (n_5494), .A1 (n_6051), .B0 (n_6558), .Y (n_6052));
NAND2X1 g63009(.A (n_9116), .B (n_9000), .Y (n_6050));
NAND2X1 g63010(.A (n_9116), .B (n_6002), .Y (n_6049));
NAND2X1 g63013(.A (n_9678), .B (n_5985), .Y (n_6048));
NAND2X1 g63014(.A (n_5985), .B (n_6032), .Y (n_6047));
AND2X1 g63015(.A (n_5337), .B (n_5716), .Y (n_6046));
NOR2X1 g63016(.A (n_5234), .B (n_8862), .Y (n_6045));
CLKBUFX1 gbuf_d_595(.A(n_5709), .Y(d_out_595));
CLKBUFX1 gbuf_q_595(.A(q_in_595), .Y(g1267));
CLKBUFX1 gbuf_d_596(.A(n_5708), .Y(d_out_596));
CLKBUFX1 gbuf_q_596(.A(q_in_596), .Y(g1268));
NAND2X1 g61269(.A (n_6075), .B (n_6322), .Y (n_6044));
INVX1 g61275(.A (n_6042), .Y (n_6043));
NAND2X1 g63038(.A (n_6039), .B (g7909), .Y (n_6041));
NAND2X1 g63052(.A (n_6039), .B (g7956), .Y (n_6040));
CLKBUFX1 gbuf_d_597(.A(n_5730), .Y(d_out_597));
CLKBUFX1 gbuf_qn_597(.A(qn_in_597), .Y(g1148));
NAND2X2 g63098(.A (n_5335), .B (n_6037), .Y (n_6473));
NOR2X1 g63179(.A (n_5717), .B (g309), .Y (n_6036));
NAND2X1 g63180(.A (n_6199), .B (n_6209), .Y (n_6035));
AND2X1 g63206(.A (n_5839), .B (n_6034), .Y (n_6486));
NAND2X1 g63221(.A (n_5987), .B (n_6032), .Y (n_6033));
NAND2X1 g63224(.A (n_9677), .B (n_5987), .Y (n_8234));
XOR2X1 g63347(.A (g_29227), .B (n_5932), .Y (n_6028));
AOI22X1 g63349(.A0 (n_5655), .A1 (n_5996), .B0 (n_5995), .B1(n_5862), .Y (n_6027));
NAND2X1 g63463(.A (n_6025), .B (g1430), .Y (n_6026));
NOR2X1 g63493(.A (n_8879), .B (n_9303), .Y (n_6023));
AND2X1 g63534(.A (n_6019), .B (n_6151), .Y (n_6307));
OAI21X1 g61516(.A0 (n_2493), .A1 (n_1691), .B0 (n_5809), .Y (n_6533));
AND2X1 g61517(.A (n_5808), .B (n_2772), .Y (n_6332));
NOR2X1 g63581(.A (n_6019), .B (n_6151), .Y (n_6452));
INVX2 g63621(.A (n_6602), .Y (n_6144));
OAI21X1 g61540(.A0 (n_6010), .A1 (n_5993), .B0 (n_4714), .Y (n_6013));
INVX1 g63693(.A (n_6012), .Y (n_6141));
OAI21X1 g61541(.A0 (n_6010), .A1 (n_5990), .B0 (n_4713), .Y (n_6011));
OAI21X1 g61542(.A0 (n_6010), .A1 (n_5988), .B0 (n_4712), .Y (n_6009));
NAND2X1 g63809(.A (n_5660), .B (n_5076), .Y (n_6008));
OAI21X1 g61553(.A0 (n_6005), .A1 (n_5528), .B0 (n_5113), .Y (n_6007));
OAI21X1 g61555(.A0 (n_6005), .A1 (n_5701), .B0 (n_5300), .Y (n_6006));
OAI21X1 g61556(.A0 (n_6005), .A1 (n_5698), .B0 (n_5297), .Y (n_6004));
NAND2X1 g63800(.A (n_6032), .B (n_6002), .Y (n_6003));
XOR2X1 g63831(.A (g_14626), .B (n_9637), .Y (n_6001));
MX2X1 g61580(.A (n_5998), .B (g582), .S0 (n_5851), .Y (n_6000));
MX2X1 g61581(.A (n_5998), .B (g583), .S0 (n_5849), .Y (n_5999));
CLKBUFX1 gbuf_d_598(.A(n_5702), .Y(d_out_598));
CLKBUFX1 gbuf_q_598(.A(q_in_598), .Y(g2656));
CLKBUFX1 gbuf_d_599(.A(n_5565), .Y(d_out_599));
CLKBUFX1 gbuf_q_599(.A(q_in_599), .Y(g585));
CLKBUFX1 gbuf_d_600(.A(n_5633), .Y(d_out_600));
CLKBUFX1 gbuf_q_600(.A(q_in_600), .Y(g586));
CLKBUFX1 gbuf_d_601(.A(n_5637), .Y(d_out_601));
CLKBUFX1 gbuf_q_601(.A(q_in_601), .Y(g1462));
CLKBUFX1 gbuf_d_602(.A(n_5634), .Y(d_out_602));
CLKBUFX1 gbuf_q_602(.A(q_in_602), .Y(g_17877));
AOI22X1 g63887(.A0 (n_5996), .A1 (n_5995), .B0 (n_5472), .B1 (g3229),.Y (n_5997));
CLKBUFX1 gbuf_d_603(.A(n_5584), .Y(d_out_603));
CLKBUFX1 gbuf_q_603(.A(q_in_603), .Y(g_19472));
CLKBUFX1 gbuf_d_604(.A(n_5583), .Y(d_out_604));
CLKBUFX1 gbuf_q_604(.A(q_in_604), .Y(g_18364));
CLKBUFX1 gbuf_d_605(.A(n_5604), .Y(d_out_605));
CLKBUFX1 gbuf_q_605(.A(q_in_605), .Y(g1457));
CLKBUFX1 gbuf_d_606(.A(n_5613), .Y(d_out_606));
CLKBUFX1 gbuf_q_606(.A(q_in_606), .Y(g_28142));
CLKBUFX1 gbuf_d_607(.A(n_5589), .Y(d_out_607));
CLKBUFX1 gbuf_q_607(.A(q_in_607), .Y(g_14751));
CLKBUFX1 gbuf_d_608(.A(n_5586), .Y(d_out_608));
CLKBUFX1 gbuf_q_608(.A(q_in_608), .Y(g_23490));
MX2X1 g61599(.A (n_5991), .B (g1264), .S0 (n_5993), .Y (n_5994));
MX2X1 g61600(.A (n_5991), .B (g1265), .S0 (n_5990), .Y (n_5992));
MX2X1 g61601(.A (n_5991), .B (g1266), .S0 (n_5988), .Y (n_5989));
CLKBUFX1 gbuf_d_609(.A(n_5558), .Y(d_out_609));
CLKBUFX1 gbuf_qn_609(.A(qn_in_609), .Y(g1164));
CLKBUFX1 gbuf_d_610(.A(n_5693), .Y(d_out_610));
CLKBUFX1 gbuf_qn_610(.A(qn_in_610), .Y(g1845));
CLKBUFX1 gbuf_d_611(.A(n_5690), .Y(d_out_611));
CLKBUFX1 gbuf_q_611(.A(q_in_611), .Y(g1865));
CLKBUFX1 gbuf_d_612(.A(n_5669), .Y(d_out_612));
CLKBUFX1 gbuf_q_612(.A(q_in_612), .Y(g_25466));
CLKBUFX1 gbuf_d_613(.A(n_5667), .Y(d_out_613));
CLKBUFX1 gbuf_q_613(.A(q_in_613), .Y(g_5159));
CLKBUFX1 gbuf_d_614(.A(n_5665), .Y(d_out_614));
CLKBUFX1 gbuf_q_614(.A(q_in_614), .Y(g_25960));
CLKBUFX1 gbuf_d_615(.A(n_5664), .Y(d_out_615));
CLKBUFX1 gbuf_q_615(.A(q_in_615), .Y(g_29721));
INVX1 g64023(.A (n_5985), .Y (n_6159));
AOI22X1 g63911(.A0 (n_5466), .A1 (n_5237), .B0 (n_5673), .B1(n_5465), .Y (n_5984));
NAND2X1 g61698(.A (n_6274), .B (g1955), .Y (n_5983));
NAND2X1 g61700(.A (n_6279), .B (g1956), .Y (n_5982));
NAND2X1 g61701(.A (n_6276), .B (g1957), .Y (n_5981));
NAND2X1 g64258(.A (n_5673), .B (n_5979), .Y (n_5980));
INVX1 g61752(.A (n_6720), .Y (n_5976));
MX2X1 g61579(.A (n_5998), .B (g581), .S0 (n_5855), .Y (n_5972));
NAND3X1 g64391(.A (n_5237), .B (n_5673), .C (g3229), .Y (n_5969));
CLKBUFX1 gbuf_d_616(.A(n_5694), .Y(d_out_616));
CLKBUFX1 gbuf_q_616(.A(q_in_616), .Y(g584));
NOR2X1 g64421(.A (n_6157), .B (n_5967), .Y (n_6148));
NOR2X1 g64428(.A (n_6250), .B (n_5966), .Y (n_6138));
INVX1 g64444(.A (n_6025), .Y (n_5965));
CLKBUFX1 gbuf_d_617(.A(n_5692), .Y(d_out_617));
CLKBUFX1 gbuf_q_617(.A(q_in_617), .Y(g1861));
AOI22X1 g64566(.A0 (n_5026), .A1 (g_22538), .B0 (n_5963), .B1(n_297), .Y (n_5964));
NOR2X1 g64599(.A (n_5770), .B (g3229), .Y (n_6254));
NOR2X1 g64614(.A (n_5768), .B (g3229), .Y (n_6252));
NOR2X1 g64682(.A (n_5767), .B (g3229), .Y (n_5962));
NOR2X1 g64696(.A (n_5774), .B (g3229), .Y (n_5961));
OAI21X1 g62110(.A0 (n_5958), .A1 (n_6106), .B0 (n_5755), .Y (n_6246));
NOR2X1 g62165(.A (n_5614), .B (n_5600), .Y (n_5957));
NOR2X1 g62172(.A (n_5612), .B (n_5183), .Y (n_5956));
NAND2X1 g62202(.A (n_5327), .B (n_5949), .Y (n_5950));
NAND3X1 g62203(.A (n_5949), .B (n_5326), .C (n_5885), .Y (n_6703));
INVX1 g62236(.A (n_5780), .Y (n_5948));
NAND4X1 g62240(.A (n_5603), .B (n_5947), .C (n_9192), .D (n_4676), .Y(n_6970));
NAND4X1 g62277(.A (n_5522), .B (n_5787), .C (n_4650), .D (n_5312), .Y(n_6286));
MX2X1 g62295(.A (g3094), .B (g2633), .S0 (g8106), .Y (n_5943));
MX2X1 g62296(.A (g3096), .B (g2633), .S0 (g3109), .Y (n_5942));
MX2X1 g62318(.A (g3095), .B (g2633), .S0 (g8030), .Y (n_5941));
OR2X1 g62414(.A (n_5651), .B (n_6565), .Y (n_5940));
NOR2X1 g62417(.A (n_5557), .B (n_5938), .Y (n_6233));
NAND3X1 g62419(.A (n_5445), .B (n_5938), .C (n_6209), .Y (n_5939));
AND2X1 g62421(.A (n_69), .B (n_5580), .Y (n_5937));
CLKBUFX1 gbuf_d_618(.A(n_5624), .Y(d_out_618));
CLKBUFX1 gbuf_q_618(.A(q_in_618), .Y(g692));
NOR2X1 g62430(.A (g1943), .B (g1939), .Y (n_5936));
OR2X1 g62458(.A (n_5864), .B (n_6478), .Y (n_5935));
NOR2X1 g62460(.A (n_5668), .B (n_6478), .Y (n_5934));
NAND3X1 g62466(.A (n_8208), .B (n_5325), .C (n_5149), .Y (n_6094));
NAND2X1 g62467(.A (n_5932), .B (n_6865), .Y (n_5933));
NAND2X1 g62472(.A (n_106), .B (n_5929), .Y (n_5930));
NOR2X1 g62477(.A (n_5577), .B (n_5134), .Y (n_8221));
NAND2X1 g62479(.A (n_5578), .B (n_5885), .Y (n_5927));
CLKBUFX1 gbuf_d_619(.A(n_5591), .Y(d_out_619));
CLKBUFX1 gbuf_q_619(.A(q_in_619), .Y(g_28702));
NAND2X1 g62507(.A (n_5920), .B (g8106), .Y (n_5926));
OR2X1 g62508(.A (n_7190), .B (n_8792), .Y (n_5925));
NAND2X1 g62518(.A (n_5920), .B (g8030), .Y (n_5921));
NAND2X1 g62522(.A (g3109), .B (n_5920), .Y (n_5919));
OR2X1 g62529(.A (n_5581), .B (g544), .Y (n_5918));
AOI21X1 g62531(.A0 (n_5462), .A1 (g2133), .B0 (g2129), .Y (n_5917));
AOI22X1 g62552(.A0 (n_5342), .A1 (n_5838), .B0 (n_5820), .B1(n_5575), .Y (n_6377));
AOI21X1 g62553(.A0 (n_920), .A1 (n_5898), .B0 (n_5545), .Y (n_6231));
CLKBUFX1 gbuf_d_620(.A(n_5700), .Y(d_out_620));
CLKBUFX1 gbuf_q_620(.A(q_in_620), .Y(g2657));
MX2X1 g62822(.A (n_4613), .B (n_4825), .S0 (n_5915), .Y (n_8236));
INVX1 g62905(.A (n_6339), .Y (n_5913));
NOR2X1 g61225(.A (n_6075), .B (n_6946), .Y (n_6357));
AND2X1 g61228(.A (n_6190), .B (n_6947), .Y (n_6350));
NOR2X1 g61229(.A (n_6330), .B (n_6946), .Y (n_6346));
NOR2X1 g61231(.A (n_5908), .B (n_6946), .Y (n_6342));
NAND2X1 g62943(.A (n_8689), .B (n_8862), .Y (n_5907));
NOR2X1 g61234(.A (n_5905), .B (n_8792), .Y (n_5906));
NAND2X1 g62959(.A (n_4244), .B (n_5713), .Y (n_5901));
NOR2X1 g61243(.A (n_5550), .B (n_5263), .Y (n_6053));
AOI21X1 g62971(.A0 (n_5493), .A1 (n_5532), .B0 (n_6464), .Y (n_5900));
NAND2X2 g62989(.A (n_8862), .B (n_5898), .Y (n_6372));
AOI22X1 g63834(.A0 (n_5049), .A1 (g_29227), .B0 (n_5446), .B1(n_5866), .Y (n_5897));
NAND2X1 g61270(.A (n_6330), .B (n_6190), .Y (n_5894));
NOR2X1 g61276(.A (n_5541), .B (n_4879), .Y (n_6042));
NAND2X1 g61277(.A (n_5892), .B (n_5560), .Y (n_5893));
NAND2X1 g61278(.A (n_5908), .B (n_5336), .Y (n_5891));
NAND2X1 g63037(.A (n_6072), .B (n_6451), .Y (n_5890));
XOR2X1 g63842(.A (g1439), .B (n_5806), .Y (n_5889));
INVX1 g61314(.A (n_5887), .Y (n_5888));
NAND2X1 g63160(.A (n_6068), .B (n_5885), .Y (n_5886));
NAND3X1 g63163(.A (n_5215), .B (n_5884), .C (g3229), .Y (n_6467));
NAND2X1 g63172(.A (n_5881), .B (g8087), .Y (n_5883));
NAND2X1 g63173(.A (n_5881), .B (g8167), .Y (n_5882));
NOR2X1 g63203(.A (n_5331), .B (n_5531), .Y (n_5880));
OR2X1 g63204(.A (n_5549), .B (n_6465), .Y (n_5879));
NAND2X1 g63223(.A (n_5569), .B (n_6032), .Y (n_5878));
NAND3X1 g63236(.A (n_5705), .B (n_5555), .C (n_6209), .Y (n_5877));
AOI21X1 g63258(.A0 (n_5223), .A1 (g1448), .B0 (g1444), .Y (n_5876));
MX2X1 g63334(.A (n_360), .B (n_5290), .S0 (g8007), .Y (n_5875));
MX2X1 g63335(.A (n_351), .B (n_5290), .S0 (g7961), .Y (n_5874));
MX2X1 g63336(.A (n_352), .B (n_5290), .S0 (g1172), .Y (n_5872));
NAND4X1 g61431(.A (n_5817), .B (n_5415), .C (n_5616), .D (n_5014), .Y(n_5871));
XOR2X1 g63345(.A (g_25523), .B (n_5475), .Y (n_5870));
INVX1 g63454(.A (n_6039), .Y (n_5868));
NAND2X1 g63468(.A (n_8730), .B (n_9129), .Y (n_5867));
INVX1 g63472(.A (n_6969), .Y (n_6171));
NOR2X1 g63485(.A (n_5866), .B (n_5932), .Y (n_6063));
NAND2X1 g63486(.A (n_5864), .B (g2124), .Y (n_5865));
AND2X1 g63488(.A (n_5862), .B (g3229), .Y (n_5863));
NAND2X1 g63552(.A (n_6051), .B (n_6212), .Y (n_6167));
INVX4 g63622(.A (n_6185), .Y (n_6602));
OAI21X1 g61536(.A0 (n_5852), .A1 (n_5855), .B0 (n_5116), .Y (n_5856));
INVX1 g63676(.A (n_5854), .Y (n_6014));
OAI21X1 g61537(.A0 (n_5852), .A1 (n_5851), .B0 (n_5115), .Y (n_5853));
OAI21X1 g61538(.A0 (n_5852), .A1 (n_5849), .B0 (n_5114), .Y (n_5850));
AND2X1 g63694(.A (n_7186), .B (n_5334), .Y (n_6012));
CLKBUFX1 gbuf_d_621(.A(n_5502), .Y(d_out_621));
CLKBUFX1 gbuf_q_621(.A(q_in_621), .Y(g2660));
CLKBUFX1 gbuf_d_622(.A(n_5381), .Y(d_out_622));
CLKBUFX1 gbuf_q_622(.A(q_in_622), .Y(g_22340));
CLKBUFX1 gbuf_d_623(.A(n_5373), .Y(d_out_623));
CLKBUFX1 gbuf_q_623(.A(q_in_623), .Y(g686));
CLKBUFX1 gbuf_d_624(.A(n_5524), .Y(d_out_624));
CLKBUFX1 gbuf_q_624(.A(q_in_624), .Y(g1270));
CLKBUFX1 gbuf_d_625(.A(n_5514), .Y(d_out_625));
CLKBUFX1 gbuf_q_625(.A(q_in_625), .Y(g1271));
CLKBUFX1 gbuf_d_626(.A(n_5506), .Y(d_out_626));
CLKBUFX1 gbuf_q_626(.A(q_in_626), .Y(g2654));
CLKBUFX1 gbuf_d_627(.A(n_5508), .Y(d_out_627));
CLKBUFX1 gbuf_q_627(.A(q_in_627), .Y(g2652));
CLKBUFX1 gbuf_d_628(.A(n_5503), .Y(d_out_628));
CLKBUFX1 gbuf_q_628(.A(q_in_628), .Y(g2659));
XOR2X1 g63883(.A (g2133), .B (n_5670), .Y (n_5848));
MX2X1 g63892(.A (g2561), .B (n_5036), .S0 (g8087), .Y (n_5847));
CLKBUFX1 gbuf_d_629(.A(n_5387), .Y(d_out_629));
CLKBUFX1 gbuf_q_629(.A(q_in_629), .Y(g_13546));
CLKBUFX1 gbuf_d_630(.A(n_5385), .Y(d_out_630));
CLKBUFX1 gbuf_q_630(.A(q_in_630), .Y(g_5095));
CLKBUFX1 gbuf_d_631(.A(n_5386), .Y(d_out_631));
CLKBUFX1 gbuf_q_631(.A(q_in_631), .Y(g_25878));
MX2X1 g63894(.A (n_5036), .B (n_819), .S0 (g2560), .Y (n_5846));
CLKBUFX1 gbuf_d_632(.A(n_5384), .Y(d_out_632));
CLKBUFX1 gbuf_q_632(.A(q_in_632), .Y(g_12505));
MX2X1 g61594(.A (n_5841), .B (g579), .S0 (n_5851), .Y (n_5844));
AOI22X1 g63896(.A0 (n_5680), .A1 (n_5547), .B0 (n_5251), .B1 (g3229),.Y (n_5843));
MX2X1 g61595(.A (n_5841), .B (g580), .S0 (n_5849), .Y (n_5842));
CLKBUFX1 gbuf_d_633(.A(n_5383), .Y(d_out_633));
CLKBUFX1 gbuf_q_633(.A(q_in_633), .Y(g_27846));
CLKBUFX1 gbuf_d_634(.A(n_5413), .Y(d_out_634));
CLKBUFX1 gbuf_q_634(.A(q_in_634), .Y(g1466));
CLKBUFX1 gbuf_d_635(.A(n_5411), .Y(d_out_635));
CLKBUFX1 gbuf_q_635(.A(q_in_635), .Y(g2151));
CLKBUFX1 gbuf_d_636(.A(n_5346), .Y(d_out_636));
CLKBUFX1 gbuf_q_636(.A(q_in_636), .Y(g1165));
CLKBUFX1 gbuf_d_637(.A(n_5345), .Y(d_out_637));
CLKBUFX1 gbuf_qn_637(.A(qn_in_637), .Y(g1166));
CLKBUFX1 gbuf_d_638(.A(n_5521), .Y(d_out_638));
CLKBUFX1 gbuf_q_638(.A(q_in_638), .Y(g1174));
CLKBUFX1 gbuf_d_639(.A(n_5500), .Y(d_out_639));
CLKBUFX1 gbuf_q_639(.A(q_in_639), .Y(g1173));
CLKBUFX1 gbuf_d_640(.A(n_5511), .Y(d_out_640));
CLKBUFX1 gbuf_qn_640(.A(qn_in_640), .Y(g1151));
CLKBUFX1 gbuf_d_641(.A(n_5510), .Y(d_out_641));
CLKBUFX1 gbuf_q_641(.A(q_in_641), .Y(g1167));
CLKBUFX1 gbuf_d_642(.A(n_5507), .Y(d_out_642));
CLKBUFX1 gbuf_q_642(.A(q_in_642), .Y(g1171));
AOI22X1 g63915(.A0 (n_5245), .A1 (n_4624), .B0 (n_5104), .B1(n_5838), .Y (n_5839));
MX2X1 g63920(.A (n_6212), .B (n_1112), .S0 (g485), .Y (n_5837));
MX2X1 g63921(.A (g484), .B (n_6212), .S0 (g7956), .Y (n_5836));
MX2X1 g63927(.A (g480), .B (n_6212), .S0 (g7909), .Y (n_5834));
CLKBUFX1 gbuf_d_643(.A(n_5433), .Y(d_out_643));
CLKBUFX1 gbuf_q_643(.A(q_in_643), .Y(g2156));
INVX1 g63980(.A (n_5832), .Y (n_5987));
CLKBUFX1 gbuf_d_644(.A(n_5504), .Y(d_out_644));
CLKBUFX1 gbuf_q_644(.A(q_in_644), .Y(g2653));
INVX1 g64024(.A (n_5828), .Y (n_5985));
XOR2X1 g64083(.A (g_32037), .B (n_8685), .Y (n_5827));
XOR2X1 g64084(.A (n_5825), .B (n_5053), .Y (n_5826));
XOR2X1 g64085(.A (g_15687), .B (n_8694), .Y (n_5824));
CLKBUFX1 gbuf_d_645(.A(n_5037), .Y(d_out_645));
CLKBUFX1 gbuf_q_645(.A(q_in_645), .Y(g_7108));
MX2X1 g61593(.A (n_5841), .B (g578), .S0 (n_5855), .Y (n_5822));
NOR2X1 g64238(.A (n_5647), .B (n_5967), .Y (n_6170));
NOR2X1 g64246(.A (n_5644), .B (n_5966), .Y (n_6161));
NAND2X1 g64253(.A (n_5104), .B (n_5820), .Y (n_5821));
NAND3X1 g61753(.A (n_5819), .B (n_5818), .C (n_5817), .Y (n_6720));
NOR2X1 g64306(.A (n_5460), .B (n_5663), .Y (n_6019));
INVX1 g64336(.A (n_6051), .Y (n_6482));
NOR2X1 g61771(.A (n_5431), .B (n_4921), .Y (n_5811));
MX2X1 g63893(.A (g2562), .B (n_5036), .S0 (g8167), .Y (n_5810));
CLKBUFX1 gbuf_d_646(.A(n_5512), .Y(d_out_646));
CLKBUFX1 gbuf_q_646(.A(q_in_646), .Y(g1272));
AOI21X1 g61804(.A0 (g1973), .A1 (n_6626), .B0 (n_5439), .Y (n_5809));
AOI21X1 g61805(.A0 (g1982), .A1 (n_6626), .B0 (n_5438), .Y (n_5808));
NOR2X1 g64445(.A (n_183), .B (n_5806), .Y (n_6025));
INVX1 g64457(.A (n_5864), .Y (n_5805));
NAND3X1 g64459(.A (n_5996), .B (n_5425), .C (g3229), .Y (n_6162));
XOR2X1 g64522(.A (g1448), .B (n_5429), .Y (n_5804));
XOR2X1 g64559(.A (g_23734), .B (n_5463), .Y (n_5803));
NOR2X1 g64600(.A (n_5801), .B (g3229), .Y (n_6156));
NOR2X1 g64613(.A (n_5800), .B (g3229), .Y (n_6139));
NOR2X1 g64662(.A (n_5798), .B (g3229), .Y (n_5799));
NOR2X1 g64702(.A (n_5796), .B (g3229), .Y (n_5797));
NAND3X1 g60757(.A (n_2823), .B (n_2468), .C (n_5193), .Y (n_6265));
NAND3X1 g60758(.A (n_2821), .B (n_2463), .C (n_5192), .Y (n_6261));
NAND2X1 g62136(.A (n_5416), .B (n_5786), .Y (n_5788));
AND2X1 g62144(.A (n_5405), .B (n_5787), .Y (n_6277));
NAND3X1 g62159(.A (n_5781), .B (n_5329), .C (n_5786), .Y (n_6707));
NOR2X1 g62166(.A (n_5417), .B (n_5350), .Y (n_5785));
NAND3X1 g62181(.A (n_5566), .B (n_5176), .C (n_5175), .Y (n_5783));
NAND2X1 g62201(.A (n_5330), .B (n_5781), .Y (n_5782));
NAND4X1 g62237(.A (n_5124), .B (n_4669), .C (n_5275), .D (n_5122), .Y(n_5780));
NAND4X1 g62239(.A (n_5410), .B (n_5779), .C (n_5778), .D (n_4678), .Y(n_6847));
NAND4X1 g62243(.A (n_4088), .B (n_4500), .C (n_4899), .D (n_5120), .Y(n_5777));
NAND4X1 g62246(.A (n_4088), .B (n_4913), .C (n_4897), .D (n_5119), .Y(n_5775));
NAND3X1 g62267(.A (n_9292), .B (n_4767), .C (n_5205), .Y (n_5773));
CLKBUFX1 gbuf_d_647(.A(n_5418), .Y(d_out_647));
CLKBUFX1 gbuf_q_647(.A(q_in_647), .Y(g2766));
NAND2X1 g62298(.A (n_588), .B (n_5406), .Y (n_5766));
NAND2X1 g62299(.A (n_700), .B (n_5408), .Y (n_5765));
NAND2X1 g62300(.A (n_881), .B (n_5407), .Y (n_5764));
OR2X1 g62411(.A (n_5462), .B (n_6478), .Y (n_5763));
OR2X1 g62438(.A (n_5223), .B (n_6565), .Y (n_5762));
NAND3X1 g62445(.A (n_4618), .B (n_4937), .C (n_5786), .Y (n_5761));
NOR2X1 g62453(.A (n_5516), .B (n_6227), .Y (n_5760));
NOR2X1 g62468(.A (n_5419), .B (n_7307), .Y (n_5759));
INVX1 g62470(.A (n_9462), .Y (n_5758));
NAND2X1 g62486(.A (n_5757), .B (g6712), .Y (n_6512));
NAND2X1 g62492(.A (n_5757), .B (n_3808), .Y (n_6509));
NAND2X1 g62495(.A (n_5757), .B (g5472), .Y (n_6507));
OR2X1 g62530(.A (g499), .B (n_1498), .Y (n_6381));
INVX1 g62535(.A (n_5755), .Y (n_5756));
CLKBUFX1 gbuf_d_648(.A(n_5529), .Y(d_out_648));
CLKBUFX1 gbuf_q_648(.A(q_in_648), .Y(g2655));
OAI21X1 g62738(.A0 (n_5974), .A1 (n_5590), .B0 (n_5165), .Y (n_5754));
OAI21X1 g62739(.A0 (n_5974), .A1 (n_5587), .B0 (n_2535), .Y (n_5753));
OAI21X1 g62740(.A0 (n_5974), .A1 (n_5585), .B0 (n_2998), .Y (n_5751));
AOI21X1 g62741(.A0 (n_6106), .A1 (n_4932), .B0 (n_4929), .Y (n_5750));
XOR2X1 g62804(.A (n_3646), .B (n_5324), .Y (n_6237));
INVX1 g62866(.A (g1880), .Y (n_6461));
CLKBUFX1 gbuf_d_649(.A(gbuf163), .Y(d_out_649));
CLKBUFX1 gbuf_qn_649(.A(qn_in_649), .Y(g1924));
INVX1 g62906(.A (n_5929), .Y (n_6339));
INVX1 g62919(.A (n_5749), .Y (n_6553));
NAND2X1 g62944(.A (n_8690), .B (n_8861), .Y (n_5748));
NAND4X1 g61315(.A (n_5338), .B (n_4574), .C (n_4361), .D (n_4354), .Y(n_5887));
NAND2X1 g63108(.A (n_5515), .B (n_4936), .Y (n_5743));
NOR2X1 g63116(.A (n_5523), .B (n_4376), .Y (n_6272));
XOR2X1 g63830(.A (n_5741), .B (n_5051), .Y (n_5742));
CLKBUFX1 gbuf_d_650(.A(n_5349), .Y(d_out_650));
CLKBUFX1 gbuf_qn_650(.A(qn_in_650), .Y(g1175));
AND2X1 g63200(.A (n_5737), .B (n_5736), .Y (n_5738));
NAND2X1 g63216(.A (n_9002), .B (n_6002), .Y (n_5735));
NAND2X1 g63219(.A (n_5573), .B (n_6002), .Y (n_5734));
AOI21X1 g63229(.A0 (n_5024), .A1 (g2142), .B0 (g2138), .Y (n_5732));
NOR2X1 g61430(.A (n_5476), .B (n_5277), .Y (n_6532));
MX2X1 g63338(.A (n_359), .B (n_5086), .S0 (g8007), .Y (n_5731));
MX2X1 g63342(.A (n_338), .B (n_5086), .S0 (g1172), .Y (n_5730));
MX2X1 g63343(.A (n_384), .B (n_5086), .S0 (g7961), .Y (n_5728));
INVX1 g63455(.A (n_5898), .Y (n_6039));
CLKBUFX1 g63473(.A (n_6037), .Y (n_6969));
NAND2X1 g63480(.A (n_4000), .B (n_9137), .Y (n_5726));
NAND2X1 g63484(.A (n_8736), .B (n_9137), .Y (n_5725));
NOR2X1 g63496(.A (n_5722), .B (n_5531), .Y (n_5723));
INVX1 g63545(.A (n_5717), .Y (n_5716));
NAND2X1 g61518(.A (n_5479), .B (n_2774), .Y (n_6322));
NOR2X1 g63582(.A (n_5714), .B (g309), .Y (n_5715));
INVX2 g63623(.A (n_5713), .Y (n_6185));
INVX1 g63643(.A (n_5902), .Y (n_5857));
INVX1 g63661(.A (n_5712), .Y (n_6199));
AND2X1 g63677(.A (n_9014), .B (n_4934), .Y (n_5854));
OAI21X1 g61543(.A0 (n_5707), .A1 (n_5993), .B0 (n_4711), .Y (n_5709));
OAI21X1 g61545(.A0 (n_5707), .A1 (n_5990), .B0 (n_4710), .Y (n_5708));
OAI21X1 g61546(.A0 (n_5707), .A1 (n_5988), .B0 (n_4709), .Y (n_5706));
INVX1 g63760(.A (n_5704), .Y (n_5705));
INVX1 g63763(.A (n_5938), .Y (n_5703));
OAI21X1 g61558(.A0 (n_5699), .A1 (n_5701), .B0 (n_5296), .Y (n_5702));
OAI21X1 g61559(.A0 (n_5699), .A1 (n_5698), .B0 (n_5295), .Y (n_5700));
NAND2X1 g63797(.A (n_5253), .B (n_4652), .Y (n_5697));
CLKBUFX1 gbuf_d_651(.A(n_5316), .Y(d_out_651));
CLKBUFX1 gbuf_q_651(.A(q_in_651), .Y(g2555));
CLKBUFX1 gbuf_d_652(.A(n_5313), .Y(d_out_652));
CLKBUFX1 gbuf_q_652(.A(q_in_652), .Y(g2658));
CLKBUFX1 gbuf_d_653(.A(n_5310), .Y(d_out_653));
CLKBUFX1 gbuf_q_653(.A(q_in_653), .Y(g2110));
CLKBUFX1 gbuf_d_654(.A(n_5182), .Y(d_out_654));
CLKBUFX1 gbuf_q_654(.A(q_in_654), .Y(g2760));
CLKBUFX1 gbuf_d_655(.A(n_5262), .Y(d_out_655));
CLKBUFX1 gbuf_q_655(.A(q_in_655), .Y(g_27699));
CLKBUFX1 gbuf_d_656(.A(n_5259), .Y(d_out_656));
CLKBUFX1 gbuf_q_656(.A(q_in_656), .Y(g_25958));
CLKBUFX1 gbuf_d_657(.A(n_5257), .Y(d_out_657));
CLKBUFX1 gbuf_q_657(.A(q_in_657), .Y(g2568));
CLKBUFX1 gbuf_d_658(.A(n_5258), .Y(d_out_658));
CLKBUFX1 gbuf_q_658(.A(q_in_658), .Y(g2565));
XOR2X1 g63889(.A (g1462), .B (n_4827), .Y (n_5696));
CLKBUFX1 gbuf_d_659(.A(n_5188), .Y(d_out_659));
CLKBUFX1 gbuf_q_659(.A(q_in_659), .Y(g1542));
CLKBUFX1 gbuf_d_660(.A(n_5187), .Y(d_out_660));
CLKBUFX1 gbuf_q_660(.A(q_in_660), .Y(g1543));
MX2X1 g61597(.A (n_5632), .B (g584), .S0 (n_5855), .Y (n_5694));
CLKBUFX1 gbuf_d_661(.A(n_5207), .Y(d_out_661));
CLKBUFX1 gbuf_q_661(.A(q_in_661), .Y(g2160));
CLKBUFX1 gbuf_d_662(.A(n_5309), .Y(d_out_662));
CLKBUFX1 gbuf_q_662(.A(q_in_662), .Y(g2109));
CLKBUFX1 gbuf_d_663(.A(n_5317), .Y(d_out_663));
CLKBUFX1 gbuf_qn_663(.A(qn_in_663), .Y(g2539));
MX2X1 g63916(.A (n_6465), .B (n_1131), .S0 (g1866), .Y (n_5693));
MX2X1 g63917(.A (g1861), .B (n_6465), .S0 (g8012), .Y (n_5692));
MX2X1 g63918(.A (g1865), .B (n_6465), .S0 (g8082), .Y (n_5690));
CLKBUFX1 gbuf_d_664(.A(n_5314), .Y(d_out_664));
CLKBUFX1 gbuf_q_664(.A(q_in_664), .Y(g2559));
NAND2X1 g63982(.A (n_5288), .B (n_5098), .Y (n_5832));
NAND2X1 g64026(.A (n_5294), .B (n_5111), .Y (n_5828));
XOR2X1 g64081(.A (g_27924), .B (n_6100), .Y (n_5686));
XOR2X1 g64092(.A (g2156), .B (n_4825), .Y (n_5685));
XOR2X1 g64097(.A (g1457), .B (n_4433), .Y (n_5683));
CLKBUFX1 gbuf_d_665(.A(n_5229), .Y(d_out_665));
CLKBUFX1 gbuf_qn_665(.A(qn_in_665), .Y(g1680));
NAND2X1 g64250(.A (n_5250), .B (n_5680), .Y (n_5681));
NAND2X2 g64251(.A (n_5434), .B (g_27924), .Y (n_5932));
NAND3X1 g64267(.A (n_4624), .B (n_5104), .C (g3229), .Y (n_5679));
NAND3X1 g64337(.A (n_1055), .B (n_5974), .C (n_8747), .Y (n_6051));
NOR2X1 g64338(.A (n_5996), .B (n_5673), .Y (n_5862));
NOR2X1 g64407(.A (n_5064), .B (n_7345), .Y (n_9591));
NOR2X1 g64458(.A (n_289), .B (n_5670), .Y (n_5864));
NAND3X1 g64462(.A (n_5680), .B (n_5022), .C (g3229), .Y (n_6034));
MX2X1 g64506(.A (g_25466), .B (n_3390), .S0 (n_5666), .Y (n_5669));
XOR2X1 g64523(.A (g2142), .B (n_5220), .Y (n_5668));
CLKBUFX1 gbuf_d_666(.A(n_5638), .Y(d_out_666));
CLKBUFX1 gbuf_q_666(.A(q_in_666), .Y(g1887));
MX2X1 g64548(.A (g_5159), .B (n_5380), .S0 (n_5666), .Y (n_5667));
MX2X1 g64551(.A (g_25960), .B (n_5382), .S0 (n_5666), .Y (n_5665));
MX2X1 g64553(.A (g_29721), .B (n_5663), .S0 (n_5666), .Y (n_5664));
INVX1 g64556(.A (n_5474), .Y (n_6032));
OAI21X1 g64581(.A0 (n_4596), .A1 (g1435), .B0 (n_5246), .Y (n_5660));
NOR2X1 g64609(.A (n_5425), .B (g3229), .Y (n_5979));
OR2X1 g64683(.A (n_5653), .B (n_5382), .Y (n_5658));
NAND2X1 g64686(.A (n_9403), .B (n_5298), .Y (n_5973));
NAND2X1 g64687(.A (n_5656), .B (g125), .Y (n_5970));
NOR2X1 g64694(.A (n_5423), .B (g3229), .Y (n_5655));
NAND2X1 g64701(.A (n_5653), .B (n_5382), .Y (n_5654));
INVX1 g64715(.A (n_5806), .Y (n_5651));
INVX1 g64879(.A (n_5647), .Y (n_6157));
INVX1 g65019(.A (n_5644), .Y (n_6250));
NAND2X1 g62140(.A (n_5638), .B (n_6626), .Y (n_6274));
NAND2X1 g62141(.A (n_5638), .B (g7052), .Y (n_6279));
NOR2X1 g62152(.A (n_5212), .B (n_4883), .Y (n_5637));
NAND2X1 g62156(.A (n_5638), .B (g7194), .Y (n_6276));
NOR2X1 g62167(.A (n_5208), .B (n_4920), .Y (n_5634));
MX2X1 g61598(.A (n_5632), .B (g586), .S0 (n_5849), .Y (n_5633));
INVX1 g65647(.A (n_5967), .Y (n_5774));
INVX1 g65649(.A (n_5801), .Y (n_5628));
NAND4X1 g62279(.A (n_4925), .B (n_5226), .C (n_3521), .D (n_4912), .Y(n_6010));
INVX1 g65764(.A (n_5798), .Y (n_5770));
INVX1 g65776(.A (n_5796), .Y (n_5768));
INVX1 g65786(.A (n_5966), .Y (n_5767));
INVX1 g65788(.A (n_5800), .Y (n_5625));
NOR2X1 g60906(.A (n_5191), .B (n_5372), .Y (n_5624));
NOR2X1 g62413(.A (n_9199), .B (n_9202), .Y (n_8222));
CLKBUFX1 gbuf_d_667(.A(n_5213), .Y(d_out_667));
CLKBUFX1 gbuf_q_667(.A(q_in_667), .Y(g2072));
AND2X1 g62428(.A (n_5616), .B (n_5615), .Y (n_5617));
OR2X1 g62452(.A (n_5552), .B (n_6227), .Y (n_5614));
NOR2X1 g62454(.A (n_5254), .B (n_6227), .Y (n_5613));
OR2X1 g62461(.A (n_5024), .B (n_6478), .Y (n_5612));
NOR2X1 g62474(.A (n_5602), .B (n_4827), .Y (n_5610));
NAND3X1 g62480(.A (n_6106), .B (n_6240), .C (n_5169), .Y (n_5609));
NOR2X1 g62482(.A (n_5156), .B (n_5605), .Y (n_5949));
NAND3X1 g62483(.A (n_5036), .B (n_5605), .C (n_5885), .Y (n_5606));
NOR2X1 g62496(.A (n_5238), .B (n_6565), .Y (n_5604));
NOR2X1 g62502(.A (n_5087), .B (n_5602), .Y (n_5603));
NAND2X1 g66239(.A (g_14632), .B (n_5004), .Y (n_9689));
AOI21X1 g62527(.A0 (n_5067), .A1 (g_26529), .B0 (g_21927), .Y(n_5600));
NAND3X1 g62536(.A (n_5958), .B (n_6106), .C (n_5169), .Y (n_5755));
NAND2X1 g66459(.A (g1698), .B (n_5008), .Y (n_9588));
AOI21X1 g62603(.A0 (n_4938), .A1 (n_5143), .B0 (g996), .Y (n_5595));
AOI21X1 g61085(.A0 (n_2302), .A1 (n_2797), .B0 (n_5179), .Y (n_5594));
AOI21X1 g61088(.A0 (n_2303), .A1 (n_2653), .B0 (n_5168), .Y (n_5593));
OAI21X1 g62684(.A0 (n_5347), .A1 (n_5605), .B0 (n_5885), .Y (n_5592));
CLKBUFX1 gbuf_d_668(.A(n_5214), .Y(d_out_668));
CLKBUFX1 gbuf_q_668(.A(q_in_668), .Y(g1378));
OAI21X1 g62735(.A0 (n_8747), .A1 (n_5590), .B0 (n_5166), .Y (n_5591));
OAI21X1 g62736(.A0 (n_8747), .A1 (n_5587), .B0 (n_2536), .Y (n_5589));
OAI21X1 g62737(.A0 (n_8747), .A1 (n_5585), .B0 (n_2999), .Y (n_5586));
OAI21X1 g62762(.A0 (n_733), .A1 (n_5590), .B0 (n_5180), .Y (n_5584));
OAI21X1 g62791(.A0 (g125), .A1 (n_5590), .B0 (n_5167), .Y (n_5583));
CLKBUFX1 gbuf_d_669(.A(n_5311), .Y(d_out_669));
CLKBUFX1 gbuf_q_669(.A(q_in_669), .Y(g2108));
INVX1 g62859(.A (g559), .Y (n_5920));
CLKBUFX1 gbuf_d_670(.A(gbuf164), .Y(d_out_670));
CLKBUFX1 gbuf_qn_670(.A(qn_in_670), .Y(g1880));
CLKBUFX1 gbuf_d_671(.A(gbuf165), .Y(d_out_671));
CLKBUFX1 gbuf_q_671(.A(q_in_671), .Y(g1939));
INVX1 g62907(.A (g499), .Y (n_5929));
INVX1 g62908(.A (g499), .Y (n_5581));
INVX1 g62920(.A (g2574), .Y (n_5749));
INVX1 g62925(.A (g2633), .Y (n_5580));
NOR2X1 g61230(.A (n_5892), .B (n_6946), .Y (n_6091));
AOI21X1 g62970(.A0 (n_5106), .A1 (n_4930), .B0 (n_6105), .Y (n_5578));
NAND4X1 g61327(.A (n_5145), .B (n_3936), .C (n_3905), .D (n_3734), .Y(n_6077));
NAND2X1 g63156(.A (n_4915), .B (n_5206), .Y (n_5577));
OR2X1 g63169(.A (n_5148), .B (n_6106), .Y (n_5576));
NAND3X1 g63201(.A (n_5020), .B (n_5575), .C (g3229), .Y (n_6232));
NAND2X1 g63218(.A (n_5573), .B (n_9000), .Y (n_5574));
NAND2X1 g63222(.A (n_9678), .B (n_5569), .Y (n_5570));
NAND4X1 g63238(.A (n_5068), .B (n_4856), .C (n_4602), .D (n_4848), .Y(n_5568));
NOR2X1 g63247(.A (n_4924), .B (n_5566), .Y (n_5567));
MX2X1 g61596(.A (n_5632), .B (g585), .S0 (n_5851), .Y (n_5565));
INVX1 g61389(.A (n_5561), .Y (n_5562));
NOR2X1 g61400(.A (n_5265), .B (n_5285), .Y (n_6323));
NOR2X1 g61420(.A (n_5264), .B (n_5279), .Y (n_6191));
INVX1 g61425(.A (n_5559), .Y (n_5560));
OAI21X1 g63339(.A0 (g1164), .A1 (g7961), .B0 (n_5137), .Y (n_5558));
MX2X1 g63352(.A (n_5530), .B (n_5556), .S0 (n_5555), .Y (n_5557));
CLKBUFX1 gbuf_d_672(.A(n_5255), .Y(d_out_672));
CLKBUFX1 gbuf_q_672(.A(q_in_672), .Y(g2571));
CLKBUFX1 gbuf_d_673(.A(n_5261), .Y(d_out_673));
CLKBUFX1 gbuf_q_673(.A(q_in_673), .Y(g_29095));
NAND2X2 g63474(.A (n_5064), .B (n_8710), .Y (n_6037));
INVX1 g63476(.A (n_9347), .Y (n_5881));
NAND2X1 g63479(.A (n_5552), .B (g_25523), .Y (n_5553));
NAND2X1 g63482(.A (n_3805), .B (n_9129), .Y (n_5551));
NAND4X1 g61501(.A (n_5286), .B (n_4550), .C (n_4315), .D (n_4084), .Y(n_5550));
NOR2X1 g63495(.A (n_6374), .B (n_6569), .Y (n_5549));
NAND2X1 g63504(.A (n_5547), .B (n_5341), .Y (n_5548));
INVX1 g63524(.A (n_5545), .Y (n_5719));
INVX1 g63541(.A (n_5543), .Y (n_6072));
NAND4X1 g61511(.A (n_5278), .B (n_4114), .C (n_3869), .D (n_3728), .Y(n_5541));
NAND2X1 g63546(.A (n_9547), .B (g_22408), .Y (n_5717));
AOI21X1 g61515(.A0 (n_2488), .A1 (n_3498), .B0 (n_5274), .Y (n_6075));
OAI21X1 g61519(.A0 (n_2391), .A1 (n_1598), .B0 (n_5272), .Y (n_6190));
AND2X1 g61520(.A (n_5271), .B (n_2618), .Y (n_6330));
CLKBUFX1 gbuf_d_674(.A(n_5190), .Y(d_out_674));
CLKBUFX1 gbuf_q_674(.A(q_in_674), .Y(g1541));
AOI21X1 g61523(.A0 (n_2172), .A1 (n_2925), .B0 (n_5267), .Y (n_5908));
INVX2 g63624(.A (n_5335), .Y (n_5713));
INVX2 g63644(.A (n_5915), .Y (n_5902));
INVX1 g63653(.A (n_5539), .Y (n_6068));
NAND2X1 g63663(.A (n_5491), .B (n_5477), .Y (n_5712));
NOR2X1 g63728(.A (n_6558), .B (g309), .Y (n_6593));
AND2X1 g63735(.A (n_6464), .B (n_6209), .Y (n_5736));
NOR2X1 g63737(.A (n_5532), .B (n_6465), .Y (n_5533));
NOR2X1 g63748(.A (n_6464), .B (n_5531), .Y (n_6517));
NAND2X1 g63761(.A (n_5530), .B (n_5556), .Y (n_5704));
NOR2X1 g63764(.A (n_5530), .B (n_5556), .Y (n_5938));
OAI21X1 g61557(.A0 (n_5699), .A1 (n_5528), .B0 (n_5110), .Y (n_5529));
AOI21X1 g63786(.A0 (n_5211), .A1 (g1457), .B0 (g1453), .Y (n_5527));
AND2X1 g63791(.A (n_6451), .B (n_6917), .Y (n_5526));
CLKBUFX1 gbuf_d_675(.A(n_4974), .Y(d_out_675));
CLKBUFX1 gbuf_q_675(.A(q_in_675), .Y(g1545));
MX2X1 g61602(.A (n_5513), .B (g1270), .S0 (n_5993), .Y (n_5524));
OAI21X1 g63806(.A0 (n_4850), .A1 (n_4096), .B0 (n_5522), .Y (n_5523));
MX2X1 g63840(.A (g1174), .B (n_4618), .S0 (g8007), .Y (n_5521));
XOR2X1 g63884(.A (g2151), .B (n_4228), .Y (n_5518));
XOR2X1 g63888(.A (g_26529), .B (n_5266), .Y (n_5516));
CLKBUFX1 gbuf_d_676(.A(n_4977), .Y(d_out_676));
CLKBUFX1 gbuf_q_676(.A(q_in_676), .Y(g1544));
CLKBUFX1 gbuf_d_677(.A(n_4972), .Y(d_out_677));
CLKBUFX1 gbuf_q_677(.A(q_in_677), .Y(g1546));
CLKBUFX1 gbuf_d_678(.A(n_5012), .Y(d_out_678));
CLKBUFX1 gbuf_q_678(.A(q_in_678), .Y(g771));
AOI22X1 g63908(.A0 (n_5282), .A1 (g1501), .B0 (n_5280), .B1 (n_473),.Y (n_5515));
MX2X1 g61603(.A (n_5513), .B (g1271), .S0 (n_5990), .Y (n_5514));
MX2X1 g61604(.A (n_5513), .B (g1272), .S0 (n_5988), .Y (n_5512));
CLKBUFX1 gbuf_d_679(.A(n_5082), .Y(d_out_679));
CLKBUFX1 gbuf_q_679(.A(q_in_679), .Y(g2244));
CLKBUFX1 gbuf_d_680(.A(n_5078), .Y(d_out_680));
CLKBUFX1 gbuf_q_680(.A(q_in_680), .Y(g2253));
MX2X1 g63919(.A (n_1145), .B (n_5414), .S0 (g1172), .Y (n_5511));
MX2X1 g63922(.A (g1167), .B (n_5414), .S0 (g7961), .Y (n_5510));
MX2X1 g61608(.A (n_5505), .B (g2652), .S0 (n_5528), .Y (n_5508));
MX2X1 g63923(.A (g1171), .B (n_5414), .S0 (g8007), .Y (n_5507));
MX2X1 g61609(.A (n_5505), .B (g2654), .S0 (n_5698), .Y (n_5506));
MX2X1 g61610(.A (n_5505), .B (g2653), .S0 (n_5701), .Y (n_5504));
MX2X1 g61612(.A (n_5501), .B (g2659), .S0 (n_5701), .Y (n_5503));
MX2X1 g61613(.A (n_5501), .B (g2660), .S0 (n_5698), .Y (n_5502));
MX2X1 g63839(.A (g1173), .B (n_4618), .S0 (g7961), .Y (n_5500));
INVX1 g63968(.A (n_9002), .Y (n_5498));
INVX1 g63970(.A (n_5573), .Y (n_5922));
INVX1 g63986(.A (n_5569), .Y (n_5687));
CLKBUFX1 gbuf_d_681(.A(n_4245), .Y(d_out_681));
CLKBUFX1 gbuf_qn_681(.A(qn_in_681), .Y(g986));
AND2X1 g64205(.A (n_5037), .B (n_6643), .Y (n_5494));
AND2X1 g64220(.A (n_5229), .B (n_6569), .Y (n_5493));
INVX1 g64235(.A (n_5491), .Y (n_5492));
NOR2X1 g64239(.A (n_5237), .B (n_5673), .Y (n_5884));
NAND2X1 g64283(.A (n_5049), .B (n_6100), .Y (n_5489));
NOR2X1 g64299(.A (n_5485), .B (n_7517), .Y (n_5486));
CLKBUFX1 gbuf_d_682(.A(n_5033), .Y(d_out_682));
CLKBUFX1 gbuf_q_682(.A(q_in_682), .Y(g776));
NOR2X1 g64384(.A (n_5480), .B (n_4838), .Y (n_5481));
AOI21X1 g61807(.A0 (g593), .A1 (n_4601), .B0 (n_5034), .Y (n_5479));
NAND4X1 g61813(.A (n_4965), .B (n_4377), .C (n_4353), .D (n_4099), .Y(n_5476));
INVX1 g64448(.A (n_5552), .Y (n_5475));
MX2X1 g64557(.A (n_5473), .B (g121), .S0 (n_5026), .Y (n_5474));
MX2X1 g64558(.A (n_467), .B (g125), .S0 (n_5027), .Y (n_6002));
NOR2X1 g64608(.A (n_5472), .B (g3229), .Y (n_5995));
NOR2X1 g64616(.A (n_5022), .B (g3229), .Y (n_5820));
NOR2X1 g64667(.A (n_5465), .B (g3229), .Y (n_5466));
NAND3X1 g64717(.A (n_5223), .B (g1448), .C (g1444), .Y (n_5806));
INVX1 g64730(.A (n_5670), .Y (n_5462));
AOI21X1 g64752(.A0 (n_3353), .A1 (n_5035), .B0 (n_5010), .Y (n_5722));
AOI21X1 g64789(.A0 (n_3066), .A1 (n_9055), .B0 (n_4999), .Y (n_5460));
AOI21X1 g64836(.A0 (n_3352), .A1 (n_5044), .B0 (n_5005), .Y (n_5714));
AOI21X1 g64881(.A0 (n_3235), .A1 (n_5044), .B0 (n_5007), .Y (n_5647));
INVX1 g64917(.A (n_7186), .Y (n_7187));
AOI21X1 g65021(.A0 (n_3061), .A1 (n_5035), .B0 (n_5003), .Y (n_5644));
OAI21X1 g62103(.A0 (n_5015), .A1 (n_5414), .B0 (n_5209), .Y (n_5819));
NOR2X1 g62148(.A (n_5016), .B (n_3856), .Y (n_5439));
NOR2X1 g62149(.A (n_5013), .B (n_3855), .Y (n_5438));
AND2X1 g62161(.A (n_4979), .B (n_5424), .Y (n_5998));
INVX1 g65378(.A (n_5434), .Y (n_5435));
NOR2X1 g62173(.A (n_5018), .B (n_4667), .Y (n_5433));
NAND4X1 g62238(.A (n_4088), .B (n_4553), .C (n_4298), .D (n_4716), .Y(n_5431));
NAND2X1 g65648(.A (n_5001), .B (n_3237), .Y (n_5967));
NAND2X1 g65650(.A (n_5002), .B (n_3354), .Y (n_5801));
NAND4X1 g62278(.A (n_4867), .B (n_5424), .C (n_4021), .D (n_4727), .Y(n_5852));
NAND4X1 g62280(.A (n_4335), .B (n_4826), .C (n_3384), .D (n_4725), .Y(n_6005));
NAND4X1 g62281(.A (n_5015), .B (n_5414), .C (n_5420), .D (n_4529), .Y(n_5422));
AOI21X1 g65766(.A0 (n_2875), .A1 (n_5044), .B0 (n_5000), .Y (n_5798));
AOI21X1 g65778(.A0 (n_3035), .A1 (n_5035), .B0 (n_5009), .Y (n_5796));
NAND2X1 g65787(.A (n_4997), .B (n_3355), .Y (n_5966));
NAND2X1 g65789(.A (n_5006), .B (n_3356), .Y (n_5800));
XOR2X1 g65816(.A (g_15687), .B (n_4792), .Y (n_5419));
NOR2X1 g60931(.A (n_4978), .B (n_5181), .Y (n_5418));
OR2X1 g62409(.A (n_5067), .B (n_6227), .Y (n_5417));
AOI21X1 g62416(.A0 (n_4708), .A1 (n_5378), .B0 (n_5420), .Y (n_5416));
OR2X1 g62431(.A (n_4966), .B (n_5414), .Y (n_5415));
NOR2X1 g62439(.A (n_5019), .B (n_6565), .Y (n_5413));
NOR2X1 g62473(.A (n_5409), .B (n_4825), .Y (n_5412));
NOR2X1 g62476(.A (n_5059), .B (n_6478), .Y (n_5411));
NOR2X1 g62485(.A (n_4954), .B (n_4937), .Y (n_5781));
NOR2X1 g62501(.A (n_5088), .B (n_5409), .Y (n_5410));
NAND2X1 g62511(.A (g1245), .B (g8030), .Y (n_5408));
NAND2X1 g62512(.A (g1245), .B (g3109), .Y (n_5407));
NAND2X1 g62517(.A (g1245), .B (g8106), .Y (n_5406));
AOI21X1 g62601(.A0 (n_4253), .A1 (n_4096), .B0 (n_4957), .Y (n_5405));
INVX1 g66651(.A (n_5008), .Y (n_6832));
MX2X1 g62753(.A (g105), .B (g_13546), .S0 (n_5590), .Y (n_5387));
MX2X1 g62756(.A (n_5247), .B (g_25878), .S0 (n_5590), .Y (n_5386));
MX2X1 g62757(.A (n_3187), .B (g_5095), .S0 (n_5590), .Y (n_5385));
MX2X1 g62765(.A (n_3161), .B (g_12505), .S0 (n_5590), .Y (n_5384));
MX2X1 g62795(.A (n_5382), .B (g_27846), .S0 (n_5590), .Y (n_5383));
MX2X1 g62799(.A (n_5380), .B (g_22340), .S0 (n_5590), .Y (n_5381));
MX2X1 g62805(.A (n_5378), .B (n_6543), .S0 (n_5414), .Y (n_5379));
CLKBUFX1 gbuf_d_683(.A(gbuf67), .Y(d_out_683));
CLKBUFX1 gbuf_qn_683(.A(qn_in_683), .Y(g559));
CLKBUFX1 gbuf_d_684(.A(gbuf66), .Y(d_out_684));
CLKBUFX1 gbuf_q_684(.A(q_in_684), .Y(g499));
CLKBUFX1 gbuf_d_685(.A(gbuf65), .Y(d_out_685));
CLKBUFX1 gbuf_q_685(.A(q_in_685), .Y(g544));
CLKBUFX1 gbuf_d_686(.A(gbuf213), .Y(d_out_686));
CLKBUFX1 gbuf_q_686(.A(q_in_686), .Y(g2574));
CLKBUFX1 gbuf_d_687(.A(gbuf212), .Y(d_out_687));
CLKBUFX1 gbuf_q_687(.A(q_in_687), .Y(g2618));
CLKBUFX1 gbuf_d_688(.A(gbuf214), .Y(d_out_688));
CLKBUFX1 gbuf_q_688(.A(q_in_688), .Y(g2633));
NAND2X1 g62935(.A (n_8551), .B (n_5368), .Y (n_5376));
NAND2X1 g62938(.A (n_9641), .B (n_9085), .Y (n_5374));
NOR2X1 g61251(.A (n_5081), .B (n_5372), .Y (n_5373));
AND2X1 g63821(.A (n_6209), .B (n_6832), .Y (n_5371));
NAND2X1 g63110(.A (n_9072), .B (n_5368), .Y (n_5369));
NAND2X1 g63112(.A (n_9072), .B (n_5319), .Y (n_5367));
NAND2X1 g63115(.A (n_9696), .B (n_5184), .Y (n_5365));
NAND2X1 g63128(.A (n_9085), .B (n_5320), .Y (n_5359));
NAND2X1 g63129(.A (n_8771), .B (n_9641), .Y (n_5358));
AND2X1 g63133(.A (n_5477), .B (n_5138), .Y (n_5357));
NOR2X1 g63157(.A (n_4926), .B (n_4362), .Y (n_5991));
AND2X1 g63167(.A (n_5355), .B (n_5354), .Y (n_5356));
NOR2X1 g63168(.A (n_5169), .B (g2384), .Y (n_5353));
INVX1 g63196(.A (n_6865), .Y (n_7307));
NAND3X1 g63228(.A (n_4939), .B (n_4441), .C (n_5786), .Y (n_5352));
AOI21X1 g63235(.A0 (n_4597), .A1 (g_28142), .B0 (g_18173), .Y(n_5350));
MX2X1 g63841(.A (n_1125), .B (n_4618), .S0 (g1172), .Y (n_5349));
NAND3X1 g63251(.A (n_5347), .B (n_5154), .C (n_5885), .Y (n_5348));
AOI21X1 g63263(.A0 (n_3873), .A1 (n_5136), .B0 (n_5086), .Y (n_5757));
NOR2X1 g61383(.A (n_5118), .B (n_1917), .Y (n_6182));
NOR2X1 g61390(.A (n_5117), .B (n_1949), .Y (n_5561));
NOR2X1 g61426(.A (n_4707), .B (n_5109), .Y (n_5559));
MX2X1 g63340(.A (g1165), .B (n_5344), .S0 (g8007), .Y (n_5346));
MX2X1 g63341(.A (n_1114), .B (n_5344), .S0 (g1172), .Y (n_5345));
INVX1 g61435(.A (n_5159), .Y (n_5343));
CLKBUFX1 gbuf_d_689(.A(n_5083), .Y(d_out_689));
CLKBUFX1 gbuf_q_689(.A(q_in_689), .Y(gbuf163));
CLKBUFX1 gbuf_d_690(.A(n_4968), .Y(d_out_690));
CLKBUFX1 gbuf_q_690(.A(q_in_690), .Y(g2066));
AND2X1 g63453(.A (n_5341), .B (g3229), .Y (n_5342));
NAND2X2 g63457(.A (n_5485), .B (n_9267), .Y (n_5898));
NAND2X1 g63467(.A (n_3643), .B (n_9302), .Y (n_8208));
NOR2X1 g61503(.A (n_4594), .B (n_5097), .Y (n_5338));
AND2X1 g63525(.A (n_7257), .B (n_5146), .Y (n_5545));
NAND2X1 g63543(.A (n_5291), .B (n_5337), .Y (n_5543));
CLKBUFX1 gbuf_d_691(.A(n_4964), .Y(d_out_691));
CLKBUFX1 gbuf_q_691(.A(q_in_691), .Y(g1372));
INVX1 g61521(.A (n_5892), .Y (n_5336));
AND2X1 g63580(.A (n_6558), .B (n_6451), .Y (n_6166));
NAND2X2 g63625(.A (n_5293), .B (n_5334), .Y (n_5335));
INVX1 g63645(.A (n_9340), .Y (n_5915));
OR2X1 g63655(.A (n_5332), .B (n_5480), .Y (n_5539));
NAND2X1 g63684(.A (n_5532), .B (n_6465), .Y (n_5737));
NOR2X1 g63688(.A (n_5329), .B (g996), .Y (n_5330));
NOR2X1 g63698(.A (n_5326), .B (g2384), .Y (n_5327));
AOI21X1 g63778(.A0 (n_5323), .A1 (n_5322), .B0 (n_5201), .Y (n_5324));
CLKBUFX1 gbuf_d_692(.A(n_4796), .Y(d_out_692));
CLKBUFX1 gbuf_q_692(.A(q_in_692), .Y(g780));
NAND2X1 g63812(.A (n_5320), .B (n_5319), .Y (n_5321));
CLKBUFX1 gbuf_d_693(.A(n_4828), .Y(d_out_693));
CLKBUFX1 gbuf_q_693(.A(q_in_693), .Y(n_3203));
CLKBUFX1 gbuf_d_694(.A(n_4787), .Y(d_out_694));
CLKBUFX1 gbuf_q_694(.A(q_in_694), .Y(g1529));
CLKBUFX1 gbuf_d_695(.A(n_4786), .Y(d_out_695));
CLKBUFX1 gbuf_q_695(.A(q_in_695), .Y(g1532));
CLKBUFX1 gbuf_d_696(.A(n_4785), .Y(d_out_696));
CLKBUFX1 gbuf_q_696(.A(q_in_696), .Y(g1535));
CLKBUFX1 gbuf_d_697(.A(n_4784), .Y(d_out_697));
CLKBUFX1 gbuf_q_697(.A(q_in_697), .Y(g1538));
XOR2X1 g63890(.A (g1448), .B (n_5162), .Y (n_5318));
CLKBUFX1 gbuf_d_698(.A(n_4779), .Y(d_out_698));
CLKBUFX1 gbuf_q_698(.A(q_in_698), .Y(g2239));
CLKBUFX1 gbuf_d_699(.A(n_4871), .Y(d_out_699));
CLKBUFX1 gbuf_q_699(.A(q_in_699), .Y(g1550));
CLKBUFX1 gbuf_d_700(.A(n_4878), .Y(d_out_700));
CLKBUFX1 gbuf_q_700(.A(q_in_700), .Y(g1553));
CLKBUFX1 gbuf_d_701(.A(n_4876), .Y(d_out_701));
CLKBUFX1 gbuf_q_701(.A(q_in_701), .Y(g2247));
CLKBUFX1 gbuf_d_702(.A(n_4875), .Y(d_out_702));
CLKBUFX1 gbuf_q_702(.A(q_in_702), .Y(g2250));
CLKBUFX1 gbuf_d_703(.A(n_4882), .Y(d_out_703));
CLKBUFX1 gbuf_q_703(.A(q_in_703), .Y(g1556));
CLKBUFX1 gbuf_d_704(.A(n_4862), .Y(d_out_704));
CLKBUFX1 gbuf_q_704(.A(q_in_704), .Y(g1559));
MX2X1 g63924(.A (n_6106), .B (n_836), .S0 (g2560), .Y (n_5317));
MX2X1 g63925(.A (g2555), .B (n_6106), .S0 (g8087), .Y (n_5316));
MX2X1 g63926(.A (g2559), .B (n_6106), .S0 (g8167), .Y (n_5314));
MX2X1 g61611(.A (n_5501), .B (g2658), .S0 (n_5528), .Y (n_5313));
AOI22X1 g63928(.A0 (n_4096), .A1 (n_4503), .B0 (n_4116), .B1(n_5200), .Y (n_5312));
MX2X1 g63944(.A (n_5323), .B (g2108), .S0 (n_3691), .Y (n_5311));
MX2X1 g63945(.A (g2110), .B (n_5323), .S0 (n_4967), .Y (n_5310));
MX2X1 g63954(.A (n_5323), .B (g2109), .S0 (n_3689), .Y (n_5309));
MX2X1 g63971(.A (n_5380), .B (g101), .S0 (n_5307), .Y (n_5573));
MX2X1 g63987(.A (n_5382), .B (g97), .S0 (n_8688), .Y (n_5569));
INVX1 g64071(.A (n_5126), .Y (n_5566));
CLKBUFX1 gbuf_d_705(.A(n_4822), .Y(d_out_705));
CLKBUFX1 gbuf_qn_705(.A(qn_in_705), .Y(g2374));
NAND2X1 g61716(.A (n_5701), .B (g2650), .Y (n_5300));
NAND2X1 g64190(.A (n_9651), .B (n_5298), .Y (n_5299));
NAND2X1 g61717(.A (n_5698), .B (g2651), .Y (n_5297));
NAND2X1 g61719(.A (n_5701), .B (g2656), .Y (n_5296));
NAND2X1 g61720(.A (n_5698), .B (g2657), .Y (n_5295));
NAND2X1 g64217(.A (n_5047), .B (n_8515), .Y (n_5294));
NOR2X1 g64236(.A (n_5287), .B (n_5293), .Y (n_5491));
INVX1 g64241(.A (n_5291), .Y (n_5292));
NAND2X1 g64279(.A (n_9632), .B (n_5247), .Y (n_5288));
AND2X1 g61763(.A (n_4805), .B (n_3895), .Y (n_5286));
NAND2X1 g61765(.A (n_4595), .B (n_4773), .Y (n_5285));
NAND2X1 g64356(.A (n_4852), .B (n_5282), .Y (n_5283));
NAND2X1 g64357(.A (n_4851), .B (n_5280), .Y (n_5281));
NAND2X1 g61787(.A (n_4593), .B (n_4765), .Y (n_5279));
AND2X1 g61788(.A (n_4804), .B (n_3737), .Y (n_5278));
NAND4X1 g61797(.A (n_4092), .B (n_4341), .C (n_4375), .D (n_4097), .Y(n_5277));
OAI21X1 g61806(.A0 (n_4580), .A1 (n_3549), .B0 (n_3347), .Y (n_5274));
AOI21X1 g61809(.A0 (g1279), .A1 (n_5270), .B0 (n_4817), .Y (n_5272));
AOI21X1 g61810(.A0 (g1288), .A1 (n_5270), .B0 (n_4816), .Y (n_5271));
INVX1 g64436(.A (n_5532), .Y (n_6374));
OAI21X1 g61812(.A0 (n_4579), .A1 (n_3548), .B0 (n_3334), .Y (n_5267));
NOR2X1 g64449(.A (n_216), .B (n_5266), .Y (n_5552));
NAND4X1 g61819(.A (n_4128), .B (n_4382), .C (n_4086), .D (n_4345), .Y(n_5265));
NAND4X1 g61820(.A (n_4363), .B (n_4381), .C (n_4338), .D (n_3886), .Y(n_5264));
NAND4X1 g61822(.A (n_4333), .B (n_4311), .C (n_4117), .D (n_4352), .Y(n_5263));
MX2X1 g61830(.A (g_27699), .B (n_5260), .S0 (g6485), .Y (n_5262));
MX2X1 g61831(.A (g_29095), .B (n_5260), .S0 (g6642), .Y (n_5261));
MX2X1 g61832(.A (g_25958), .B (n_5260), .S0 (n_4601), .Y (n_5259));
MX2X1 g61840(.A (g2565), .B (n_5256), .S0 (g7302), .Y (n_5258));
MX2X1 g61841(.A (g2568), .B (n_5256), .S0 (g7390), .Y (n_5257));
MX2X1 g61842(.A (n_5256), .B (g2571), .S0 (n_3448), .Y (n_5255));
XOR2X1 g64528(.A (g_28142), .B (n_4813), .Y (n_5254));
OAI21X1 g64579(.A0 (n_4206), .A1 (g2129), .B0 (n_4847), .Y (n_5253));
NOR2X1 g64615(.A (n_5251), .B (g3229), .Y (n_5547));
NOR2X1 g64640(.A (n_5023), .B (g3229), .Y (n_5250));
NAND2X1 g64697(.A (n_4596), .B (g1435), .Y (n_5246));
NOR2X1 g64705(.A (n_5838), .B (g3229), .Y (n_5245));
NAND3X1 g64732(.A (n_5024), .B (g2142), .C (g2138), .Y (n_5670));
CLKBUFX1 gbuf_d_706(.A(n_4788), .Y(d_out_706));
CLKBUFX1 gbuf_q_706(.A(q_in_706), .Y(g1511));
INVX1 g64774(.A (n_5485), .Y (n_7371));
INVX1 g64918(.A (n_6713), .Y (n_7186));
INVX1 g64927(.A (n_7277), .Y (n_7345));
INVX1 g64953(.A (n_7347), .Y (n_5239));
XOR2X1 g64963(.A (g1457), .B (n_5025), .Y (n_5238));
INVX1 g64997(.A (n_5237), .Y (n_5996));
INVX1 g65072(.A (n_5049), .Y (n_5446));
INVX1 g65080(.A (n_5232), .Y (n_6697));
INVX1 g65118(.A (n_5231), .Y (n_5230));
INVX1 g65125(.A (n_5555), .Y (n_5445));
INVX1 g65146(.A (n_6150), .Y (n_5444));
INVX1 g65309(.A (n_6465), .Y (n_5229));
NOR2X1 g65421(.A (n_4798), .B (n_1234), .Y (n_5227));
NAND3X1 g62193(.A (n_5226), .B (n_4675), .C (n_4524), .Y (n_5707));
OR2X1 g65514(.A (n_4797), .B (n_1107), .Y (n_5656));
INVX1 g65525(.A (n_5028), .Y (n_5653));
INVX1 g65542(.A (n_5026), .Y (n_5963));
INVX1 g65563(.A (n_5223), .Y (n_5429));
CLKBUFX1 gbuf_d_707(.A(n_4778), .Y(d_out_707));
CLKBUFX1 gbuf_q_707(.A(q_in_707), .Y(g2240));
INVX1 g65692(.A (n_5465), .Y (n_5425));
INVX1 g65747(.A (n_5673), .Y (n_5423));
INVX1 g65749(.A (n_5472), .Y (n_5215));
NOR2X1 g65828(.A (n_4791), .B (n_87), .Y (n_5434));
NOR2X1 g60896(.A (n_4783), .B (n_4963), .Y (n_5214));
NOR2X1 g60904(.A (n_4782), .B (n_4967), .Y (n_5213));
OR2X1 g62406(.A (n_5211), .B (n_6565), .Y (n_5212));
INVX1 g62424(.A (n_5209), .Y (n_5210));
OR2X1 g62455(.A (n_4597), .B (n_6227), .Y (n_5208));
NOR2X1 g62462(.A (n_4801), .B (n_6478), .Y (n_5207));
INVX1 g63864(.A (n_5205), .Y (n_5206));
NAND2X1 g66206(.A (g_16638), .B (n_9314), .Y (n_8257));
NAND2X1 g66325(.A (g1004), .B (n_6420), .Y (n_5202));
OAI21X1 g62544(.A0 (n_4731), .A1 (n_5201), .B0 (n_3529), .Y (n_5638));
AOI22X1 g62554(.A0 (n_3723), .A1 (n_3363), .B0 (n_5200), .B1(n_4355), .Y (n_6132));
NAND2X1 g66401(.A (g_26067), .B (n_9314), .Y (n_5199));
NAND2X1 g66404(.A (g1122), .B (n_6420), .Y (n_5198));
NAND2X1 g66419(.A (g237), .B (n_9314), .Y (n_9621));
NAND2X1 g66425(.A (g2392), .B (n_4576), .Y (n_5196));
NAND2X1 g66495(.A (g273), .B (n_9314), .Y (n_8230));
AOI21X1 g61080(.A0 (n_2168), .A1 (n_2635), .B0 (n_4772), .Y (n_5193));
AOI21X1 g61084(.A0 (n_2167), .A1 (n_2508), .B0 (n_4771), .Y (n_5192));
XOR2X1 g61104(.A (g692), .B (n_4614), .Y (n_5191));
MX2X1 g62717(.A (n_5189), .B (g1541), .S0 (n_4975), .Y (n_5190));
MX2X1 g62718(.A (n_5189), .B (g1542), .S0 (n_4973), .Y (n_5188));
MX2X1 g62719(.A (n_5189), .B (g1543), .S0 (n_4971), .Y (n_5187));
INVX1 g62911(.A (g1245), .Y (n_5186));
NAND2X1 g62942(.A (n_5378), .B (n_5414), .Y (n_5616));
AOI21X1 g63802(.A0 (n_5017), .A1 (g2151), .B0 (g2147), .Y (n_5183));
NOR2X1 g61279(.A (n_4866), .B (n_5181), .Y (n_5182));
NAND2X1 g63050(.A (g_19472), .B (n_5590), .Y (n_5180));
NOR2X1 g61317(.A (n_4752), .B (n_3951), .Y (n_5179));
NAND2X1 g63109(.A (n_4769), .B (n_5319), .Y (n_5178));
NAND2X1 g63122(.A (n_5011), .B (n_4923), .Y (n_5176));
NAND2X1 g63123(.A (n_9289), .B (n_8986), .Y (n_5175));
NAND2X1 g63127(.A (n_5171), .B (n_5320), .Y (n_5172));
NOR2X1 g61331(.A (n_4751), .B (n_3773), .Y (n_5168));
NAND2X1 g63138(.A (g_18364), .B (n_5590), .Y (n_5167));
NAND2X1 g63149(.A (g_28702), .B (n_5590), .Y (n_5166));
NAND2X1 g63162(.A (g_14677), .B (n_5590), .Y (n_5165));
NOR2X1 g63170(.A (n_4869), .B (n_4127), .Y (n_5841));
OR2X1 g63197(.A (n_4088), .B (n_5590), .Y (n_6865));
NAND4X1 g63240(.A (n_4846), .B (n_4244), .C (n_5163), .D (n_5162), .Y(n_5602));
CLKBUFX1 gbuf_d_708(.A(n_4781), .Y(d_out_708));
CLKBUFX1 gbuf_q_708(.A(q_in_708), .Y(g2238));
AOI21X1 g61436(.A0 (n_4894), .A1 (n_2657), .B0 (n_4515), .Y (n_5159));
INVX1 g61437(.A (n_4955), .Y (n_5157));
MX2X1 g63354(.A (n_4928), .B (n_5155), .S0 (n_5154), .Y (n_5156));
CLKBUFX1 gbuf_d_709(.A(n_4873), .Y(d_out_709));
CLKBUFX1 gbuf_q_709(.A(q_in_709), .Y(g1183));
CLKBUFX1 gbuf_d_710(.A(n_4865), .Y(d_out_710));
CLKBUFX1 gbuf_q_710(.A(q_in_710), .Y(gbuf164));
CLKBUFX1 gbuf_d_711(.A(n_4881), .Y(d_out_711));
CLKBUFX1 gbuf_q_711(.A(q_in_711), .Y(gbuf165));
CLKBUFX1 gbuf_d_712(.A(n_4870), .Y(d_out_712));
CLKBUFX1 gbuf_q_712(.A(q_in_712), .Y(g1177));
CLKBUFX1 gbuf_d_713(.A(n_4874), .Y(d_out_713));
CLKBUFX1 gbuf_q_713(.A(q_in_713), .Y(g1180));
NAND2X1 g63481(.A (n_8411), .B (n_9119), .Y (n_5149));
NOR2X1 g63494(.A (n_5958), .B (n_6240), .Y (n_5148));
NOR2X1 g61512(.A (n_4411), .B (n_4885), .Y (n_5145));
AOI21X1 g61522(.A0 (n_2177), .A1 (n_2925), .B0 (n_4884), .Y (n_5892));
INVX1 g63627(.A (n_6529), .Y (n_5141));
INVX1 g63668(.A (n_5138), .Y (n_5331));
NAND2X1 g63685(.A (n_5344), .B (g7961), .Y (n_5137));
NAND2X2 g63709(.A (n_5136), .B (n_9302), .Y (n_5325));
NOR2X1 g63770(.A (g996), .B (n_6420), .Y (n_5135));
CLKBUFX1 gbuf_d_714(.A(n_4547), .Y(d_out_714));
CLKBUFX1 gbuf_q_714(.A(q_in_714), .Y(g848));
CLKBUFX1 gbuf_d_715(.A(n_4542), .Y(d_out_715));
CLKBUFX1 gbuf_q_715(.A(q_in_715), .Y(g851));
CLKBUFX1 gbuf_d_716(.A(n_4598), .Y(d_out_716));
CLKBUFX1 gbuf_q_716(.A(q_in_716), .Y(g2740));
INVX1 g63876(.A (n_9289), .Y (n_5134));
XOR2X1 g63885(.A (g2142), .B (n_4756), .Y (n_5133));
CLKBUFX1 gbuf_d_717(.A(n_4551), .Y(d_out_717));
CLKBUFX1 gbuf_q_717(.A(q_in_717), .Y(g2229));
CLKBUFX1 gbuf_d_718(.A(n_4563), .Y(d_out_718));
CLKBUFX1 gbuf_q_718(.A(q_in_718), .Y(g2232));
CLKBUFX1 gbuf_d_719(.A(n_4559), .Y(d_out_719));
CLKBUFX1 gbuf_q_719(.A(q_in_719), .Y(g1523));
CLKBUFX1 gbuf_d_720(.A(n_4548), .Y(d_out_720));
CLKBUFX1 gbuf_q_720(.A(q_in_720), .Y(g847));
CLKBUFX1 gbuf_d_721(.A(n_4544), .Y(d_out_721));
CLKBUFX1 gbuf_q_721(.A(q_in_721), .Y(g850));
CLKBUFX1 gbuf_d_722(.A(n_4539), .Y(d_out_722));
CLKBUFX1 gbuf_q_722(.A(q_in_722), .Y(g852));
CLKBUFX1 gbuf_d_723(.A(n_4535), .Y(d_out_723));
CLKBUFX1 gbuf_q_723(.A(q_in_723), .Y(g2235));
NAND2X1 g63907(.A (n_4666), .B (n_4665), .Y (n_5132));
INVX1 g64063(.A (n_5129), .Y (n_5303));
INVX2 g64073(.A (n_9290), .Y (n_5126));
XOR2X1 g64087(.A (g_25523), .B (n_4223), .Y (n_5124));
XOR2X1 g64088(.A (g776), .B (n_4240), .Y (n_5122));
XOR2X1 g64095(.A (g2124), .B (n_4678), .Y (n_5120));
XOR2X1 g64099(.A (g1430), .B (n_4676), .Y (n_5119));
OAI21X1 g61695(.A0 (n_2847), .A1 (n_2814), .B0 (n_4693), .Y (n_5118));
OAI21X1 g61699(.A0 (n_2973), .A1 (n_2674), .B0 (n_4894), .Y (n_5117));
NAND2X1 g61705(.A (n_5855), .B (g575), .Y (n_5116));
NAND2X1 g61706(.A (n_5851), .B (g576), .Y (n_5115));
NAND2X1 g61707(.A (n_5849), .B (g577), .Y (n_5114));
NAND2X1 g61715(.A (n_5528), .B (g2649), .Y (n_5113));
NAND2X1 g64191(.A (n_9444), .B (n_9509), .Y (n_5112));
NAND2X1 g64193(.A (n_4831), .B (n_8740), .Y (n_5111));
NAND2X1 g61718(.A (n_5528), .B (g2655), .Y (n_5110));
NAND4X1 g61723(.A (n_3879), .B (n_4342), .C (n_3909), .D (n_3580), .Y(n_5109));
NAND3X1 g61725(.A (n_4894), .B (n_2657), .C (n_4515), .Y (n_5108));
AND2X1 g64218(.A (n_4822), .B (n_6240), .Y (n_5106));
NAND2X1 g64234(.A (n_4838), .B (n_9014), .Y (n_5332));
NOR2X1 g64237(.A (n_4844), .B (n_4842), .Y (n_5334));
NOR2X1 g64242(.A (n_5099), .B (n_9216), .Y (n_5291));
NOR2X1 g64247(.A (n_4624), .B (n_5104), .Y (n_5575));
NAND3X1 g61740(.A (n_4693), .B (n_2646), .C (n_5101), .Y (n_5103));
INVX1 g64256(.A (n_5136), .Y (n_5290));
NAND3X1 g61742(.A (n_4693), .B (n_3313), .C (n_4737), .Y (n_5100));
NOR2X1 g64265(.A (n_5680), .B (n_5104), .Y (n_5341));
CLKBUFX1 gbuf_d_724(.A(n_4612), .Y(d_out_724));
CLKBUFX1 gbuf_q_724(.A(q_in_724), .Y(n_3143));
NAND2X1 g64281(.A (n_9640), .B (g113), .Y (n_5098));
NAND4X1 g61766(.A (n_3741), .B (n_3892), .C (n_4090), .D (n_4095), .Y(n_5097));
NOR2X1 g64358(.A (n_4626), .B (n_4861), .Y (n_5530));
AND2X1 g64361(.A (n_4840), .B (n_7000), .Y (n_8280));
NAND2X1 g64378(.A (n_4228), .B (n_4825), .Y (n_5088));
NAND2X1 g64380(.A (n_4433), .B (n_4827), .Y (n_5087));
INVX1 g64415(.A (n_5086), .Y (n_5275));
NAND3X1 g64437(.A (n_775), .B (n_4477), .C (n_4410), .Y (n_5532));
CLKBUFX1 gbuf_d_725(.A(n_4603), .Y(d_out_725));
CLKBUFX1 gbuf_q_725(.A(q_in_725), .Y(g666));
CLKBUFX1 gbuf_d_726(.A(n_4545), .Y(d_out_726));
CLKBUFX1 gbuf_q_726(.A(q_in_726), .Y(g849));
AOI21X1 g64475(.A0 (n_4420), .A1 (n_4880), .B0 (n_1094), .Y (n_5083));
OAI21X1 g64484(.A0 (n_2952), .A1 (n_5077), .B0 (n_4649), .Y (n_5082));
XOR2X1 g61834(.A (g686), .B (n_4357), .Y (n_5081));
OAI21X1 g64544(.A0 (n_4674), .A1 (n_5077), .B0 (n_4648), .Y (n_5078));
CLKBUFX1 gbuf_d_727(.A(n_4561), .Y(d_out_727));
CLKBUFX1 gbuf_q_727(.A(q_in_727), .Y(g1514));
CLKBUFX1 gbuf_d_728(.A(n_4558), .Y(d_out_728));
CLKBUFX1 gbuf_q_728(.A(q_in_728), .Y(g1526));
XOR2X1 g64582(.A (g1439), .B (n_6603), .Y (n_5076));
OR2X1 g64629(.A (n_5071), .B (n_454), .Y (n_5073));
NAND2X1 g64630(.A (n_5071), .B (n_454), .Y (n_5072));
NAND2X1 g64664(.A (n_5069), .B (n_4410), .Y (n_5482));
NAND2X1 g64676(.A (n_4213), .B (n_293), .Y (n_5068));
INVX1 g64720(.A (n_5266), .Y (n_5067));
AOI21X1 g64767(.A0 (n_2599), .A1 (n_3810), .B0 (n_4572), .Y (n_5329));
INVX1 g64784(.A (n_5099), .Y (n_7517));
INVX1 g64849(.A (n_5064), .Y (n_5477));
CLKBUFX1 gbuf_d_729(.A(n_4663), .Y(d_out_729));
CLKBUFX1 gbuf_q_729(.A(q_in_729), .Y(g856));
INVX1 g64908(.A (n_9219), .Y (n_7257));
CLKBUFX1 g64919(.A (n_5293), .Y (n_6713));
CLKBUFX1 g64929(.A (n_5287), .Y (n_7277));
INVX1 g64947(.A (n_5480), .Y (n_7194));
INVX1 g64954(.A (n_4627), .Y (n_7347));
XOR2X1 g64991(.A (g2151), .B (n_4809), .Y (n_5059));
AOI21X1 g64999(.A0 (n_3063), .A1 (n_4604), .B0 (n_4568), .Y (n_5237));
AOI21X1 g65001(.A0 (n_2901), .A1 (n_5044), .B0 (n_4573), .Y (n_6643));
AOI21X1 g65006(.A0 (n_3232), .A1 (n_4604), .B0 (n_4567), .Y (n_5326));
AOI21X1 g65027(.A0 (n_2751), .A1 (n_5035), .B0 (n_4564), .Y (n_6569));
INVX1 g65051(.A (n_5053), .Y (n_5234));
INVX1 g65057(.A (n_5051), .Y (n_5233));
INVX1 g65081(.A (n_5047), .Y (n_5232));
INVX1 g65119(.A (n_8685), .Y (n_5231));
AOI22X1 g65126(.A0 (n_2913), .A1 (n_5035), .B0 (n_6832), .B1 (g1825),.Y (n_5555));
AOI22X1 g65143(.A0 (n_3073), .A1 (n_5044), .B0 (g435), .B1 (n_6917),.Y (n_6151));
AOI22X1 g65147(.A0 (n_3072), .A1 (n_5044), .B0 (n_6917), .B1 (g444),.Y (n_6150));
AOI22X1 g65165(.A0 (n_3069), .A1 (n_5044), .B0 (g414), .B1 (n_6917),.Y (n_6558));
AOI22X1 g65363(.A0 (n_2903), .A1 (n_5035), .B0 (g1795), .B1 (n_6832),.Y (n_6464));
NOR2X1 g62162(.A (n_4581), .B (n_3547), .Y (n_5034));
NOR2X1 g62168(.A (n_4583), .B (n_4265), .Y (n_5033));
INVX1 g65418(.A (n_4818), .Y (n_5469));
INVX1 g65439(.A (n_5031), .Y (n_5032));
NAND3X1 g65444(.A (n_1121), .B (n_2568), .C (n_4394), .Y (n_5030));
OR2X1 g65463(.A (n_4585), .B (n_1108), .Y (n_5029));
NOR2X1 g65510(.A (n_2915), .B (n_9314), .Y (n_5666));
NAND3X1 g65526(.A (n_1030), .B (n_2572), .C (n_4379), .Y (n_5028));
CLKBUFX1 g65536(.A (n_5027), .Y (n_5463));
NOR2X1 g65564(.A (n_182), .B (n_5025), .Y (n_5223));
INVX1 g65600(.A (n_5024), .Y (n_5220));
INVX1 g65688(.A (n_5838), .Y (n_5022));
AOI21X1 g65694(.A0 (n_2738), .A1 (n_4604), .B0 (n_4570), .Y (n_5465));
CLKBUFX1 g65743(.A (n_5298), .Y (n_5974));
NAND2X1 g65748(.A (n_4577), .B (n_3068), .Y (n_5673));
NAND2X1 g65750(.A (n_4578), .B (n_3236), .Y (n_5472));
INVX1 g65790(.A (n_5251), .Y (n_5020));
XOR2X1 g65813(.A (g1466), .B (n_4393), .Y (n_5019));
OR2X1 g62412(.A (n_5017), .B (n_6478), .Y (n_5018));
NAND2X1 g62423(.A (g1904), .B (g185), .Y (n_5016));
NAND3X1 g62425(.A (n_5015), .B (n_5414), .C (n_6543), .Y (n_5209));
NAND3X1 g62432(.A (n_5414), .B (n_5818), .C (n_6543), .Y (n_5014));
NAND2X1 g62437(.A (g1922), .B (g185), .Y (n_5013));
NOR2X1 g62456(.A (n_4625), .B (n_6227), .Y (n_5012));
INVX1 g63865(.A (n_5011), .Y (n_5205));
NOR2X1 g66202(.A (g1828), .B (n_5008), .Y (n_5010));
NOR2X1 g66204(.A (g1757), .B (n_5008), .Y (n_5009));
NOR2X1 g66205(.A (g346), .B (n_5004), .Y (n_5007));
OR2X1 g66280(.A (g1772), .B (n_5008), .Y (n_5006));
NOR2X1 g66289(.A (g447), .B (n_5004), .Y (n_5005));
NOR2X1 g66293(.A (g1727), .B (n_5008), .Y (n_5003));
OR2X1 g66342(.A (g391), .B (n_5004), .Y (n_5002));
OR2X1 g66360(.A (g361), .B (n_5004), .Y (n_5001));
NOR2X1 g66385(.A (g376), .B (n_5004), .Y (n_5000));
AOI22X1 g62556(.A0 (n_4319), .A1 (n_3684), .B0 (n_4726), .B1(n_3893), .Y (n_5632));
NOR2X1 g66441(.A (g_29721), .B (n_9314), .Y (n_4999));
OR2X1 g66467(.A (g1742), .B (n_5008), .Y (n_4997));
INVX1 g66864(.A (n_4576), .Y (n_4985));
AOI21X1 g62680(.A0 (n_4019), .A1 (n_3685), .B0 (n_4525), .Y (n_4979));
XOR2X1 g61106(.A (g2766), .B (n_4436), .Y (n_4978));
MX2X1 g62720(.A (n_4976), .B (g1544), .S0 (n_4975), .Y (n_4977));
MX2X1 g62721(.A (n_4976), .B (g1545), .S0 (n_4973), .Y (n_4974));
MX2X1 g62722(.A (n_4976), .B (g1546), .S0 (n_4971), .Y (n_4972));
AND2X1 g63803(.A (n_5885), .B (n_6611), .Y (n_4970));
CLKBUFX1 gbuf_d_730(.A(gbuf115), .Y(d_out_730));
CLKBUFX1 gbuf_q_730(.A(q_in_730), .Y(n_6219));
CLKBUFX1 gbuf_d_731(.A(gbuf114), .Y(d_out_731));
CLKBUFX1 gbuf_q_731(.A(q_in_731), .Y(g1230));
CLKBUFX1 gbuf_d_732(.A(gbuf116), .Y(d_out_732));
CLKBUFX1 gbuf_q_732(.A(q_in_732), .Y(g1245));
NOR2X1 g61247(.A (n_4659), .B (n_4967), .Y (n_4968));
NOR2X1 g63023(.A (n_5015), .B (n_5818), .Y (n_4966));
OR4X1 g63039(.A (n_4096), .B (n_4351), .C (n_1750), .D (n_4278), .Y(n_4965));
NOR2X1 g61281(.A (n_4662), .B (n_4963), .Y (n_4964));
CLKBUFX1 gbuf_d_733(.A(n_4531), .Y(d_out_733));
CLKBUFX1 gbuf_q_733(.A(q_in_733), .Y(g2236));
CLKBUFX1 gbuf_d_734(.A(n_4533), .Y(d_out_734));
CLKBUFX1 gbuf_q_734(.A(q_in_734), .Y(g2237));
NAND2X1 g63268(.A (n_4504), .B (n_4471), .Y (n_4957));
AOI21X1 g61438(.A0 (n_4894), .A1 (n_3136), .B0 (n_4517), .Y (n_4955));
MX2X1 g63355(.A (n_4732), .B (n_4953), .S0 (n_4441), .Y (n_4954));
INVX1 g61459(.A (n_4742), .Y (n_4952));
INVX1 g61461(.A (n_4741), .Y (n_4951));
INVX1 g61463(.A (n_4739), .Y (n_4950));
INVX1 g61465(.A (n_4738), .Y (n_4949));
INVX1 g61467(.A (n_4736), .Y (n_4948));
CLKBUFX1 gbuf_d_735(.A(n_4661), .Y(d_out_735));
CLKBUFX1 gbuf_q_735(.A(q_in_735), .Y(gbuf65));
INVX1 g61469(.A (n_4735), .Y (n_4947));
CLKBUFX1 gbuf_d_736(.A(n_4664), .Y(d_out_736));
CLKBUFX1 gbuf_q_736(.A(q_in_736), .Y(gbuf67));
AOI21X1 g61471(.A0 (n_4693), .A1 (n_2646), .B0 (n_5101), .Y (n_4946));
INVX1 g61472(.A (n_4734), .Y (n_4945));
AOI21X1 g61474(.A0 (n_4693), .A1 (n_3313), .B0 (n_4737), .Y (n_4944));
CLKBUFX1 gbuf_d_737(.A(n_4658), .Y(d_out_737));
CLKBUFX1 gbuf_q_737(.A(q_in_737), .Y(gbuf66));
INVX1 g61475(.A (n_4733), .Y (n_4941));
CLKBUFX1 gbuf_d_738(.A(n_4656), .Y(d_out_738));
CLKBUFX1 gbuf_q_738(.A(q_in_738), .Y(gbuf213));
CLKBUFX1 gbuf_d_739(.A(n_4657), .Y(d_out_739));
CLKBUFX1 gbuf_q_739(.A(q_in_739), .Y(gbuf212));
CLKBUFX1 gbuf_d_740(.A(n_4654), .Y(d_out_740));
CLKBUFX1 gbuf_q_740(.A(q_in_740), .Y(gbuf214));
INVX1 g63569(.A (n_4938), .Y (n_4939));
INVX1 g63573(.A (n_4937), .Y (n_5143));
CLKBUFX1 g63628(.A (n_4936), .Y (n_6529));
NOR2X1 g63669(.A (n_4591), .B (n_4055), .Y (n_5138));
NAND2X1 g63689(.A (n_4930), .B (n_6106), .Y (n_5355));
AND2X1 g63690(.A (n_6105), .B (n_5885), .Y (n_5354));
NOR2X1 g63691(.A (n_4930), .B (n_6106), .Y (n_4929));
NOR2X1 g63695(.A (n_6105), .B (g2384), .Y (n_6154));
AND2X1 g63696(.A (n_4928), .B (n_5155), .Y (n_5347));
NOR2X1 g63697(.A (n_4928), .B (n_5155), .Y (n_5605));
NOR2X1 g63699(.A (n_8960), .B (g996), .Y (n_4927));
OAI21X1 g63799(.A0 (n_4449), .A1 (n_3648), .B0 (n_4925), .Y (n_4926));
NAND2X1 g63798(.A (n_4923), .B (n_9538), .Y (n_4924));
NAND2X1 g63793(.A (n_4456), .B (n_4457), .Y (n_4921));
AOI21X1 g63795(.A0 (n_4582), .A1 (g771), .B0 (g_17877), .Y (n_4920));
CLKBUFX1 gbuf_d_741(.A(n_4435), .Y(d_out_741));
CLKBUFX1 gbuf_q_741(.A(q_in_741), .Y(n_2880));
NAND2X1 g63818(.A (g_22408), .B (n_9315), .Y (n_5590));
INVX1 g63873(.A (n_4918), .Y (n_4919));
CLKBUFX1 gbuf_d_742(.A(n_4423), .Y(d_out_742));
CLKBUFX1 gbuf_q_742(.A(q_in_742), .Y(g1352));
INVX1 g63878(.A (n_9288), .Y (n_4917));
INVX1 g63880(.A (n_8984), .Y (n_4915));
CLKBUFX1 gbuf_d_743(.A(n_4366), .Y(d_out_743));
CLKBUFX1 gbuf_q_743(.A(q_in_743), .Y(g2220));
XOR2X1 g63891(.A (g_22536), .B (n_5947), .Y (n_4913));
CLKBUFX1 gbuf_d_744(.A(n_4364), .Y(d_out_744));
CLKBUFX1 gbuf_q_744(.A(q_in_744), .Y(g2226));
CLKBUFX1 gbuf_d_745(.A(n_4397), .Y(d_out_745));
CLKBUFX1 gbuf_q_745(.A(q_in_745), .Y(g2746));
CLKBUFX1 gbuf_d_746(.A(n_4462), .Y(d_out_746));
CLKBUFX1 gbuf_qn_746(.A(qn_in_746), .Y(g1934));
CLKBUFX1 gbuf_d_747(.A(n_4459), .Y(d_out_747));
CLKBUFX1 gbuf_q_747(.A(q_in_747), .Y(g859));
CLKBUFX1 gbuf_d_748(.A(n_4458), .Y(d_out_748));
CLKBUFX1 gbuf_q_748(.A(q_in_748), .Y(g865));
CLKBUFX1 gbuf_d_749(.A(n_4401), .Y(d_out_749));
CLKBUFX1 gbuf_q_749(.A(q_in_749), .Y(g1937));
AOI22X1 g63931(.A0 (n_3648), .A1 (n_4523), .B0 (n_3515), .B1(n_4789), .Y (n_4912));
INVX1 g63972(.A (n_9448), .Y (n_4910));
INVX2 g64064(.A (n_8990), .Y (n_5129));
XOR2X1 g64086(.A (g1466), .B (n_4244), .Y (n_4902));
XOR2X1 g64094(.A (g2160), .B (n_4900), .Y (n_4901));
XOR2X1 g64096(.A (g2138), .B (n_4757), .Y (n_4899));
XOR2X1 g64098(.A (g1453), .B (n_9192), .Y (n_4898));
XOR2X1 g64100(.A (g1444), .B (n_5163), .Y (n_4897));
NOR2X1 g64202(.A (n_2651), .B (n_4037), .Y (n_4896));
NAND3X1 g61728(.A (n_4894), .B (n_2942), .C (n_4515), .Y (n_4895));
CLKBUFX1 gbuf_d_750(.A(n_4461), .Y(d_out_750));
CLKBUFX1 gbuf_q_750(.A(q_in_750), .Y(g862));
NOR2X1 g64240(.A (n_4631), .B (n_4630), .Y (n_5146));
NAND2X2 g64257(.A (n_4670), .B (n_8894), .Y (n_5136));
NOR2X1 g64359(.A (n_4627), .B (n_9024), .Y (n_5150));
INVX1 g64395(.A (n_4930), .Y (n_5958));
OAI21X1 g61800(.A0 (n_3412), .A1 (n_1962), .B0 (n_4409), .Y (n_4885));
INVX1 g64400(.A (n_8960), .Y (n_5344));
AND2X1 g64416(.A (n_3959), .B (n_8652), .Y (n_5086));
CLKBUFX1 gbuf_d_751(.A(n_4439), .Y(d_out_751));
CLKBUFX1 gbuf_q_751(.A(q_in_751), .Y(n_2834));
OAI21X1 g61811(.A0 (n_4183), .A1 (n_3290), .B0 (n_3056), .Y (n_4884));
AOI21X1 g64446(.A0 (n_4584), .A1 (g1466), .B0 (g1462), .Y (n_4883));
NAND3X1 g64460(.A (n_4096), .B (n_3628), .C (g3229), .Y (n_5522));
MX2X1 g64472(.A (g1556), .B (n_365), .S0 (n_4877), .Y (n_4882));
AOI21X1 g64473(.A0 (n_4205), .A1 (n_4880), .B0 (n_1137), .Y (n_4881));
NAND4X1 g61824(.A (n_4083), .B (n_4054), .C (n_3907), .D (n_3880), .Y(n_4879));
MX2X1 g64477(.A (g1553), .B (n_364), .S0 (n_4877), .Y (n_4878));
MX2X1 g64487(.A (n_2809), .B (g2247), .S0 (n_5077), .Y (n_4876));
MX2X1 g64490(.A (n_4368), .B (g2250), .S0 (n_5077), .Y (n_4875));
MX2X1 g61837(.A (g1180), .B (n_4872), .S0 (g6944), .Y (n_4874));
MX2X1 g61838(.A (g1183), .B (n_4872), .S0 (n_5270), .Y (n_4873));
CLKBUFX1 gbuf_d_752(.A(n_4428), .Y(d_out_752));
CLKBUFX1 gbuf_q_752(.A(q_in_752), .Y(g2046));
MX2X1 g64502(.A (g1550), .B (n_2946), .S0 (n_4877), .Y (n_4871));
MX2X1 g61839(.A (g1177), .B (n_4872), .S0 (g6750), .Y (n_4870));
OAI21X1 g63808(.A0 (n_4018), .A1 (n_3685), .B0 (n_4867), .Y (n_4869));
XOR2X1 g61843(.A (g2760), .B (n_4101), .Y (n_4866));
AOI21X1 g64511(.A0 (n_4201), .A1 (n_4880), .B0 (n_1132), .Y (n_4865));
XOR2X1 g64527(.A (g2195), .B (n_4210), .Y (n_4863));
CLKBUFX1 gbuf_d_753(.A(n_4815), .Y(d_out_753));
CLKBUFX1 gbuf_q_753(.A(q_in_753), .Y(g2581));
MX2X1 g64547(.A (g1559), .B (n_4861), .S0 (n_4877), .Y (n_4862));
CLKBUFX1 gbuf_d_754(.A(n_4378), .Y(d_out_754));
CLKBUFX1 gbuf_q_754(.A(q_in_754), .Y(g2208));
INVX1 g64567(.A (n_4859), .Y (n_5319));
INVX1 g64573(.A (n_4857), .Y (n_5320));
MX2X1 g64586(.A (n_365), .B (g1471), .S0 (n_4208), .Y (n_4856));
XOR2X1 g64589(.A (n_482), .B (n_4216), .Y (n_4853));
NAND2X1 g64633(.A (n_4852), .B (g1501), .Y (n_5282));
NAND2X1 g64634(.A (n_4851), .B (n_473), .Y (n_5280));
OR2X1 g64657(.A (n_3363), .B (g3229), .Y (n_4850));
CLKBUFX1 gbuf_d_755(.A(n_4367), .Y(d_out_755));
CLKBUFX1 gbuf_q_755(.A(q_in_755), .Y(g2217));
OR2X1 g64671(.A (n_4426), .B (n_435), .Y (n_4849));
NAND2X1 g64677(.A (n_4599), .B (n_600), .Y (n_4848));
NAND2X1 g64698(.A (n_4206), .B (g2129), .Y (n_4847));
NAND3X1 g64722(.A (n_4597), .B (g_18173), .C (g_28142), .Y (n_5266));
NOR2X1 g64729(.A (n_4653), .B (n_4202), .Y (n_4846));
INVX1 g64776(.A (n_5485), .Y (n_5337));
INVX1 g64850(.A (n_4844), .Y (n_5064));
CLKBUFX1 gbuf_d_756(.A(n_4365), .Y(d_out_756));
CLKBUFX1 gbuf_q_756(.A(q_in_756), .Y(g2223));
INVX2 g64920(.A (n_4843), .Y (n_5293));
INVX1 g64930(.A (n_4842), .Y (n_5287));
INVX1 g65039(.A (n_5307), .Y (n_6100));
CLKBUFX1 g65053(.A (n_4836), .Y (n_5053));
INVX1 g65058(.A (n_9509), .Y (n_5051));
INVX1 g65059(.A (n_9509), .Y (n_9651));
INVX1 g65075(.A (n_8995), .Y (n_5049));
INVX1 g65082(.A (n_4831), .Y (n_5047));
CLKBUFX1 gbuf_d_757(.A(n_4359), .Y(d_out_757));
CLKBUFX1 gbuf_q_757(.A(q_in_757), .Y(g838));
NOR2X1 g62108(.A (n_4330), .B (n_5372), .Y (n_4828));
NAND3X1 g62111(.A (n_4826), .B (n_3862), .C (n_4079), .Y (n_5699));
INVX1 g65285(.A (n_6106), .Y (n_4822));
INVX1 g65296(.A (n_6212), .Y (n_5037));
INVX1 g65318(.A (n_5154), .Y (n_5036));
NAND3X1 g65419(.A (n_1109), .B (n_2418), .C (n_4164), .Y (n_4818));
NAND3X1 g65440(.A (n_8206), .B (n_4175), .C (n_8207), .Y (n_5031));
NOR2X1 g62198(.A (n_4399), .B (n_3398), .Y (n_4817));
NOR2X1 g62199(.A (n_4398), .B (n_3397), .Y (n_4816));
NAND2X1 g62209(.A (n_4815), .B (g7302), .Y (n_5701));
NAND2X1 g62210(.A (n_4815), .B (g7390), .Y (n_5698));
NAND3X1 g65537(.A (n_1138), .B (n_2253), .C (n_4160), .Y (n_5027));
NAND3X1 g65545(.A (n_1117), .B (n_2250), .C (n_4176), .Y (n_5026));
NOR2X1 g65601(.A (n_131), .B (n_4809), .Y (n_5024));
INVX1 g65616(.A (n_5104), .Y (n_5023));
AOI21X1 g65690(.A0 (n_2362), .A1 (n_3810), .B0 (n_4392), .Y (n_5838));
AOI21X1 g62274(.A0 (n_4374), .A1 (n_4098), .B0 (n_4389), .Y (n_4805));
AOI21X1 g62275(.A0 (n_4592), .A1 (n_4380), .B0 (n_4387), .Y (n_4804));
INVX1 g65744(.A (n_9444), .Y (n_5298));
OAI21X1 g65791(.A0 (g1078), .A1 (n_3336), .B0 (n_2907), .Y (n_5251));
CLKBUFX1 gbuf_d_758(.A(n_4358), .Y(d_out_758));
CLKBUFX1 gbuf_q_758(.A(q_in_758), .Y(g844));
XOR2X1 g65815(.A (g2160), .B (n_4152), .Y (n_4801));
NAND3X1 g65837(.A (n_4395), .B (n_2569), .C (n_1134), .Y (n_4800));
INVX2 g63866(.A (n_9285), .Y (n_5011));
CLKBUFX1 gbuf_d_759(.A(n_4400), .Y(d_out_759));
CLKBUFX1 gbuf_q_759(.A(q_in_759), .Y(n_5322));
OAI22X1 g66031(.A0 (g_12505), .A1 (n_9314), .B0 (g_19162), .B1(n_2579), .Y (n_4798));
INVX1 g66032(.A (n_5025), .Y (n_5211));
OAI21X1 g66075(.A0 (g_18364), .A1 (n_9314), .B0 (n_2436), .Y(n_4797));
CLKBUFX1 gbuf_d_760(.A(n_4369), .Y(d_out_760));
CLKBUFX1 gbuf_q_760(.A(q_in_760), .Y(g2205));
NOR2X1 g62457(.A (n_4403), .B (n_6227), .Y (n_4796));
INVX1 g66297(.A (n_4790), .Y (n_4792));
INVX1 g66298(.A (n_4790), .Y (n_4791));
NOR2X1 g62537(.A (n_4337), .B (n_3559), .Y (n_5505));
AOI22X1 g62558(.A0 (n_3722), .A1 (n_3524), .B0 (n_4789), .B1(n_4081), .Y (n_5513));
OAI21X1 g62607(.A0 (n_4975), .A1 (g1471), .B0 (n_4350), .Y (n_4788));
OAI21X1 g62619(.A0 (n_4975), .A1 (n_600), .B0 (n_4349), .Y (n_4787));
OAI21X1 g62622(.A0 (n_4975), .A1 (n_471), .B0 (n_4346), .Y (n_4786));
OAI21X1 g62626(.A0 (n_4975), .A1 (g1501), .B0 (n_4348), .Y (n_4785));
OAI21X1 g62629(.A0 (n_4975), .A1 (n_473), .B0 (n_4347), .Y (n_4784));
XOR2X1 g61101(.A (g1378), .B (n_4239), .Y (n_4783));
XOR2X1 g61103(.A (g2072), .B (n_4234), .Y (n_4782));
MX2X1 g62732(.A (n_4780), .B (g2238), .S0 (n_4562), .Y (n_4781));
MX2X1 g62733(.A (g2239), .B (n_4780), .S0 (n_4530), .Y (n_4779));
MX2X1 g62734(.A (g2240), .B (n_4780), .S0 (n_4532), .Y (n_4778));
NAND2X1 g62991(.A (n_4718), .B (n_8609), .Y (n_4777));
NAND4X1 g63063(.A (n_3822), .B (n_3863), .C (n_2039), .D (n_4029), .Y(n_4773));
NOR2X1 g61304(.A (n_4334), .B (n_3766), .Y (n_4772));
NOR2X1 g61316(.A (n_4331), .B (n_3765), .Y (n_4771));
NAND2X1 g63111(.A (n_9296), .B (n_9538), .Y (n_4770));
NAND2X1 g63124(.A (n_8986), .B (n_4923), .Y (n_4767));
NAND4X1 g63182(.A (n_4053), .B (n_3735), .C (n_1754), .D (n_4028), .Y(n_4765));
NAND4X1 g63239(.A (n_4448), .B (n_4900), .C (n_4757), .D (n_4756), .Y(n_5409));
NAND2X1 g63249(.A (n_8909), .B (n_4729), .Y (n_4755));
NAND2X1 g63254(.A (n_8609), .B (n_9229), .Y (n_8255));
NOR2X1 g61386(.A (n_4480), .B (n_1603), .Y (n_5905));
NOR2X1 g61387(.A (n_4479), .B (n_1730), .Y (n_6179));
NAND4X1 g61402(.A (n_3120), .B (n_4207), .C (n_2961), .D (n_3293), .Y(n_4752));
NAND4X1 g61429(.A (n_3301), .B (n_4203), .C (n_3130), .D (n_3131), .Y(n_4751));
INVX1 g61439(.A (n_4522), .Y (n_4750));
INVX1 g61441(.A (n_4521), .Y (n_4749));
INVX1 g61443(.A (n_4519), .Y (n_4748));
INVX1 g61445(.A (n_4518), .Y (n_4747));
INVX1 g61447(.A (n_4516), .Y (n_4746));
INVX1 g61449(.A (n_4514), .Y (n_4745));
INVX1 g61451(.A (n_4513), .Y (n_4744));
INVX1 g61453(.A (n_4512), .Y (n_4743));
AOI21X1 g61460(.A0 (n_4740), .A1 (n_4695), .B0 (n_5101), .Y (n_4742));
AOI21X1 g61462(.A0 (n_4740), .A1 (n_2786), .B0 (n_4737), .Y (n_4741));
AOI21X1 g61464(.A0 (n_4740), .A1 (n_4691), .B0 (n_5101), .Y (n_4739));
AOI21X1 g61466(.A0 (n_4740), .A1 (n_4689), .B0 (n_4737), .Y (n_4738));
AOI21X1 g61468(.A0 (n_4740), .A1 (n_4687), .B0 (n_5101), .Y (n_4736));
AOI21X1 g61470(.A0 (n_4740), .A1 (n_4685), .B0 (n_4737), .Y (n_4735));
AOI21X1 g61473(.A0 (n_4740), .A1 (n_4683), .B0 (n_5101), .Y (n_4734));
AOI21X1 g61476(.A0 (n_4740), .A1 (n_4681), .B0 (n_4737), .Y (n_4733));
INVX1 g63461(.A (n_5015), .Y (n_5378));
NAND2X1 g63570(.A (n_4732), .B (n_4953), .Y (n_4938));
NOR2X1 g63574(.A (n_4732), .B (n_4953), .Y (n_4937));
NOR2X1 g63629(.A (n_4590), .B (n_4055), .Y (n_4936));
INVX1 g63659(.A (n_5169), .Y (n_4932));
AOI21X1 g63780(.A0 (n_4037), .A1 (n_5322), .B0 (n_4151), .Y (n_4731));
INVX1 g63874(.A (n_5171), .Y (n_4918));
INVX1 g63845(.A (n_4769), .Y (n_4728));
CLKBUFX1 gbuf_d_761(.A(n_4113), .Y(d_out_761));
CLKBUFX1 gbuf_q_761(.A(q_in_761), .Y(g817));
CLKBUFX1 gbuf_d_762(.A(n_4187), .Y(d_out_762));
CLKBUFX1 gbuf_q_762(.A(q_in_762), .Y(g2052));
CLKBUFX1 gbuf_d_763(.A(n_4181), .Y(d_out_763));
CLKBUFX1 gbuf_q_763(.A(q_in_763), .Y(g1358));
CLKBUFX1 gbuf_d_764(.A(n_4308), .Y(d_out_764));
CLKBUFX1 gbuf_q_764(.A(q_in_764), .Y(g2802));
CLKBUFX1 gbuf_d_765(.A(n_4305), .Y(d_out_765));
CLKBUFX1 gbuf_q_765(.A(q_in_765), .Y(g2804));
CLKBUFX1 gbuf_d_766(.A(n_4301), .Y(d_out_766));
CLKBUFX1 gbuf_q_766(.A(q_in_766), .Y(g2806));
AOI22X1 g63933(.A0 (n_3685), .A1 (n_3834), .B0 (n_3359), .B1(n_4726), .Y (n_4727));
AOI22X1 g63934(.A0 (n_4078), .A1 (n_4569), .B0 (n_3534), .B1(n_4077), .Y (n_4725));
OAI22X1 g63994(.A0 (n_4011), .A1 (n_496), .B0 (n_4010), .B1 (g805),.Y (n_4722));
INVX2 g64039(.A (n_4718), .Y (n_4958));
CLKBUFX1 gbuf_d_767(.A(n_4309), .Y(d_out_767));
CLKBUFX1 gbuf_q_767(.A(q_in_767), .Y(g2807));
XOR2X1 g64089(.A (g_18173), .B (n_3812), .Y (n_4717));
XOR2X1 g64090(.A (g_17877), .B (n_6653), .Y (n_4716));
XOR2X1 g64093(.A (g2147), .B (n_5778), .Y (n_4715));
NAND2X1 g61708(.A (n_5993), .B (g1261), .Y (n_4714));
NAND2X1 g61709(.A (n_5990), .B (g1262), .Y (n_4713));
NAND2X1 g61710(.A (n_5988), .B (g1263), .Y (n_4712));
NAND2X1 g61711(.A (n_5993), .B (g1267), .Y (n_4711));
NAND2X1 g61712(.A (n_5990), .B (g1268), .Y (n_4710));
NAND2X1 g61713(.A (n_5988), .B (g1269), .Y (n_4709));
AND2X1 g64189(.A (n_4245), .B (n_5818), .Y (n_4708));
NAND4X1 g61722(.A (n_3726), .B (n_3931), .C (n_3428), .D (n_3414), .Y(n_4707));
OR2X1 g61726(.A (n_3289), .B (n_4698), .Y (n_4706));
OR2X1 g61727(.A (n_3287), .B (n_4698), .Y (n_4704));
OR2X1 g61729(.A (n_3285), .B (n_4698), .Y (n_4703));
OR2X1 g61730(.A (n_3283), .B (n_4698), .Y (n_4701));
OR2X1 g61731(.A (n_3282), .B (n_4698), .Y (n_4700));
OR2X1 g61732(.A (n_3280), .B (n_4698), .Y (n_4699));
OR2X1 g61733(.A (n_3278), .B (n_4698), .Y (n_4697));
NAND3X1 g61734(.A (n_4693), .B (n_4695), .C (n_5101), .Y (n_4696));
NOR2X1 g64233(.A (n_4446), .B (n_9437), .Y (n_4934));
NAND3X1 g61735(.A (n_4693), .B (n_2786), .C (n_4737), .Y (n_4694));
NAND3X1 g61736(.A (n_4693), .B (n_4691), .C (n_5101), .Y (n_4692));
NAND3X1 g61737(.A (n_4693), .B (n_4689), .C (n_4737), .Y (n_4690));
NAND3X1 g61738(.A (n_4693), .B (n_4687), .C (n_5101), .Y (n_4688));
NAND3X1 g61739(.A (n_4693), .B (n_4685), .C (n_4737), .Y (n_4686));
NAND3X1 g61741(.A (n_4693), .B (n_4683), .C (n_5101), .Y (n_4684));
NAND3X1 g61743(.A (n_4693), .B (n_4681), .C (n_4737), .Y (n_4682));
NOR2X1 g64379(.A (n_5779), .B (n_4678), .Y (n_4679));
NOR2X1 g64381(.A (n_5947), .B (n_4676), .Y (n_4677));
NAND3X1 g64385(.A (n_4053), .B (n_3515), .C (g3229), .Y (n_4675));
NAND3X1 g64396(.A (n_4674), .B (n_9463), .C (n_4672), .Y (n_4930));
AND2X1 g64398(.A (n_4246), .B (n_4674), .Y (n_4928));
XOR2X1 g63836(.A (g771), .B (n_8730), .Y (n_4669));
AOI21X1 g64451(.A0 (n_4402), .A1 (g2160), .B0 (g2156), .Y (n_4667));
NOR2X1 g64452(.A (n_3981), .B (n_4221), .Y (n_4666));
NOR2X1 g64453(.A (n_4220), .B (n_4219), .Y (n_4665));
AOI21X1 g64474(.A0 (n_3974), .A1 (n_4660), .B0 (n_1102), .Y (n_4664));
OAI21X1 g64479(.A0 (n_2811), .A1 (n_4460), .B0 (n_4254), .Y (n_4663));
XOR2X1 g61825(.A (g1372), .B (n_3901), .Y (n_4662));
AOI21X1 g64483(.A0 (n_3972), .A1 (n_4660), .B0 (n_1142), .Y (n_4661));
XOR2X1 g61833(.A (g2066), .B (n_3903), .Y (n_4659));
AOI21X1 g64494(.A0 (n_3977), .A1 (n_4660), .B0 (n_1113), .Y (n_4658));
AOI21X1 g64507(.A0 (n_3979), .A1 (n_4655), .B0 (n_846), .Y (n_4657));
AOI21X1 g64508(.A0 (n_3968), .A1 (n_4655), .B0 (n_837), .Y (n_4656));
AOI21X1 g64510(.A0 (n_3966), .A1 (n_4655), .B0 (n_820), .Y (n_4654));
CLKBUFX1 gbuf_d_768(.A(n_4605), .Y(d_out_768));
CLKBUFX1 gbuf_qn_768(.A(qn_in_768), .Y(g_8090));
MX2X1 g64569(.A (n_473), .B (n_337), .S0 (n_4202), .Y (n_4859));
MX2X1 g64575(.A (g1501), .B (n_343), .S0 (n_4653), .Y (n_4857));
XOR2X1 g64580(.A (g2133), .B (n_6414), .Y (n_4652));
NOR2X1 g64596(.A (n_3628), .B (g3229), .Y (n_5200));
NAND2X1 g64597(.A (n_3625), .B (g3229), .Y (n_4650));
NAND2X1 g64625(.A (n_5077), .B (g2244), .Y (n_4649));
NAND2X1 g64628(.A (n_5077), .B (g2253), .Y (n_4648));
OR2X1 g64672(.A (n_4425), .B (g1481), .Y (n_4644));
NAND2X1 g64674(.A (n_4640), .B (n_4639), .Y (n_4642));
OR2X1 g64675(.A (n_4640), .B (n_4639), .Y (n_4641));
NAND2X1 g64678(.A (n_8939), .B (n_4672), .Y (n_5089));
NAND2X1 g64679(.A (n_4635), .B (n_436), .Y (n_4637));
OR2X1 g64680(.A (n_4635), .B (n_436), .Y (n_4636));
NOR2X1 g64695(.A (n_4670), .B (n_4192), .Y (n_9666));
INVX1 g64777(.A (n_4631), .Y (n_5485));
INVX1 g64787(.A (n_4630), .Y (n_5099));
OR2X1 g64818(.A (n_4161), .B (n_2920), .Y (n_7091));
OAI21X1 g64851(.A0 (n_2480), .A1 (n_2336), .B0 (n_4145), .Y (n_4844));
NAND2X1 g64921(.A (n_4153), .B (n_2765), .Y (n_4843));
CLKBUFX1 gbuf_d_769(.A(n_4182), .Y(d_out_769));
CLKBUFX1 gbuf_q_769(.A(q_in_769), .Y(g2734));
AOI21X1 g64931(.A0 (n_2602), .A1 (n_2046), .B0 (n_4062), .Y (n_4842));
INVX1 g64950(.A (n_5480), .Y (n_4840));
INVX1 g64957(.A (n_4627), .Y (n_4838));
AOI21X1 g64960(.A0 (n_2589), .A1 (n_4412), .B0 (n_4155), .Y (n_4626));
XOR2X1 g64967(.A (g771), .B (n_4418), .Y (n_4625));
AOI21X1 g65002(.A0 (n_2752), .A1 (n_4604), .B0 (n_4140), .Y (n_6240));
NAND2X1 g65022(.A (n_4137), .B (n_2917), .Y (n_7215));
INVX1 g65023(.A (n_5680), .Y (n_4624));
NAND2X2 g65040(.A (n_4171), .B (n_8810), .Y (n_5307));
OAI21X1 g65054(.A0 (n_2613), .A1 (n_2346), .B0 (n_4170), .Y (n_4836));
AOI21X1 g65083(.A0 (n_2492), .A1 (n_2921), .B0 (n_4139), .Y (n_4831));
AOI22X1 g65177(.A0 (n_2902), .A1 (n_5035), .B0 (g1816), .B1 (n_6832),.Y (n_5556));
NAND2X1 g62109(.A (n_4356), .B (g686), .Y (n_4614));
NOR2X1 g62112(.A (n_4080), .B (n_5181), .Y (n_4612));
AOI22X1 g65298(.A0 (n_2761), .A1 (n_5044), .B0 (g423), .B1 (n_6917),.Y (n_6212));
AOI22X1 g65307(.A0 (n_2909), .A1 (n_4604), .B0 (g2489), .B1 (n_6611),.Y (n_6105));
AOI22X1 g65314(.A0 (n_2608), .A1 (n_5035), .B0 (g1804), .B1 (n_6832),.Y (n_6465));
NAND2X1 g62139(.A (n_4605), .B (g6485), .Y (n_5851));
AOI22X1 g65319(.A0 (n_2904), .A1 (n_4604), .B0 (g2476), .B1 (g2519),.Y (n_5154));
NOR2X1 g62163(.A (n_4063), .B (n_3940), .Y (n_4603));
MX2X1 g65379(.A (n_79), .B (g1476), .S0 (n_3954), .Y (n_4602));
NAND2X1 g62191(.A (n_4605), .B (n_4601), .Y (n_5855));
NAND3X1 g65446(.A (n_1028), .B (n_2322), .C (n_3929), .Y (n_5069));
NAND2X1 g62204(.A (n_4605), .B (g6642), .Y (n_5849));
OR2X1 g62207(.A (n_4388), .B (n_3448), .Y (n_5528));
NOR2X1 g62214(.A (n_4060), .B (n_4159), .Y (n_4598));
INVX1 g65480(.A (n_4424), .Y (n_5071));
INVX1 g65576(.A (n_4597), .Y (n_4813));
OAI21X1 g65617(.A0 (g1048), .A1 (n_3336), .B0 (n_2910), .Y (n_5104));
AOI21X1 g62262(.A0 (n_3891), .A1 (n_4360), .B0 (n_4105), .Y (n_4595));
NAND4X1 g62263(.A (n_3420), .B (n_3743), .C (n_3709), .D (n_3731), .Y(n_4594));
AOI21X1 g62271(.A0 (n_4592), .A1 (n_3906), .B0 (n_4103), .Y (n_4593));
INVX1 g65704(.A (n_4590), .Y (n_4591));
INVX1 g65709(.A (n_4410), .Y (n_5189));
INVX1 g65754(.A (n_3959), .Y (n_7155));
NAND2X1 g65983(.A (n_2441), .B (n_4179), .Y (n_4585));
NAND3X1 g66033(.A (n_4584), .B (g1462), .C (g1466), .Y (n_5025));
OR2X1 g62410(.A (n_4582), .B (n_6227), .Y (n_4583));
INVX1 g66050(.A (n_4809), .Y (n_5017));
CLKBUFX1 gbuf_d_770(.A(n_4185), .Y(d_out_770));
CLKBUFX1 gbuf_q_770(.A(q_in_770), .Y(g672));
NAND2X1 g62447(.A (g524), .B (g185), .Y (n_4581));
NAND2X1 g62448(.A (g542), .B (g185), .Y (n_4580));
CLKBUFX1 gbuf_d_771(.A(n_4106), .Y(d_out_771));
CLKBUFX1 gbuf_q_771(.A(q_in_771), .Y(g841));
NAND2X1 g62488(.A (g2616), .B (g185), .Y (n_4579));
CLKBUFX1 gbuf_d_772(.A(n_4188), .Y(d_out_772));
CLKBUFX1 gbuf_q_772(.A(q_in_772), .Y(g660));
NOR2X1 g66299(.A (n_3873), .B (n_9314), .Y (n_4790));
OR2X1 g66327(.A (g2466), .B (n_4576), .Y (n_4578));
OR2X1 g66329(.A (g2436), .B (n_4576), .Y (n_4577));
AOI21X1 g62542(.A0 (n_3844), .A1 (n_1756), .B0 (n_4089), .Y (n_4574));
NOR2X1 g66421(.A (g426), .B (n_5004), .Y (n_4573));
NOR2X1 g66426(.A (g1134), .B (n_3336), .Y (n_4572));
NOR2X1 g66434(.A (g2451), .B (n_4576), .Y (n_4570));
AOI22X1 g62561(.A0 (n_3423), .A1 (n_3533), .B0 (n_4569), .B1(n_3430), .Y (n_5501));
NOR2X1 g66436(.A (g2421), .B (n_4576), .Y (n_4568));
NOR2X1 g66450(.A (g2522), .B (n_4576), .Y (n_4567));
NOR2X1 g66491(.A (g1807), .B (n_5008), .Y (n_4564));
OAI21X1 g62602(.A0 (n_4562), .A1 (n_482), .B0 (n_4087), .Y (n_4563));
MX2X1 g62610(.A (n_364), .B (g1514), .S0 (n_4975), .Y (n_4561));
MX2X1 g62613(.A (n_435), .B (g1523), .S0 (n_4975), .Y (n_4559));
MX2X1 g62616(.A (n_454), .B (g1526), .S0 (n_4975), .Y (n_4558));
INVX1 g66925(.A (n_3808), .Y (n_6420));
XOR2X1 g63844(.A (g_28142), .B (n_4339), .Y (n_4553));
CLKBUFX1 gbuf_d_773(.A(n_4306), .Y(d_out_773));
CLKBUFX1 gbuf_q_773(.A(q_in_773), .Y(g2803));
OAI21X1 g62674(.A0 (n_4562), .A1 (g2195), .B0 (n_4093), .Y (n_4551));
AOI21X1 g62703(.A0 (n_3872), .A1 (n_4096), .B0 (n_3871), .Y (n_4550));
OAI21X1 g62723(.A0 (n_4280), .A1 (n_4543), .B0 (n_3876), .Y (n_4548));
OAI21X1 g62724(.A0 (n_4280), .A1 (n_4540), .B0 (n_3006), .Y (n_4547));
OAI21X1 g62725(.A0 (n_4280), .A1 (n_4538), .B0 (n_3005), .Y (n_4545));
OAI21X1 g62726(.A0 (n_4281), .A1 (n_4543), .B0 (n_3889), .Y (n_4544));
OAI21X1 g62727(.A0 (n_4281), .A1 (n_4540), .B0 (n_3004), .Y (n_4542));
OAI21X1 g62728(.A0 (n_4281), .A1 (n_4538), .B0 (n_3000), .Y (n_4539));
XOR2X1 g63843(.A (g_21690), .B (n_8884), .Y (n_4537));
MX2X1 g62729(.A (n_4534), .B (g2235), .S0 (n_4562), .Y (n_4535));
MX2X1 g62730(.A (g2237), .B (n_4534), .S0 (n_4532), .Y (n_4533));
MX2X1 g62731(.A (g2236), .B (n_4534), .S0 (n_4530), .Y (n_4531));
CLKBUFX1 gbuf_d_774(.A(n_4304), .Y(d_out_774));
CLKBUFX1 gbuf_q_774(.A(q_in_774), .Y(g2805));
XOR2X1 g62806(.A (n_3499), .B (n_4058), .Y (n_5260));
XOR2X1 g62811(.A (n_3636), .B (n_4051), .Y (n_5256));
CLKBUFX1 gbuf_d_775(.A(n_4107), .Y(d_out_775));
CLKBUFX1 gbuf_q_775(.A(q_in_775), .Y(g835));
CLKBUFX1 gbuf_d_776(.A(gbuf152), .Y(d_out_776));
CLKBUFX1 gbuf_q_776(.A(q_in_776), .Y(g1904));
CLKBUFX1 gbuf_d_777(.A(gbuf162), .Y(d_out_777));
CLKBUFX1 gbuf_q_777(.A(q_in_777), .Y(g1922));
CLKBUFX1 gbuf_d_778(.A(n_4108), .Y(d_out_778));
CLKBUFX1 gbuf_q_778(.A(q_in_778), .Y(g832));
CLKBUFX1 gbuf_d_779(.A(n_4109), .Y(d_out_779));
CLKBUFX1 gbuf_q_779(.A(q_in_779), .Y(g829));
NOR2X1 g63020(.A (g996), .B (n_6543), .Y (n_4529));
NOR2X1 g63097(.A (n_4670), .B (n_6543), .Y (n_4528));
NAND2X1 g63212(.A (n_9229), .B (n_4729), .Y (n_4527));
OAI21X1 g63279(.A0 (n_3833), .A1 (n_3677), .B0 (n_4270), .Y (n_4525));
AOI22X1 g63348(.A0 (n_4017), .A1 (n_3648), .B0 (n_4523), .B1(n_3721), .Y (n_4524));
AOI21X1 g61440(.A0 (n_4520), .A1 (n_3288), .B0 (n_4515), .Y (n_4522));
AOI21X1 g61442(.A0 (n_4520), .A1 (n_3286), .B0 (n_4517), .Y (n_4521));
AOI21X1 g61444(.A0 (n_4520), .A1 (n_2942), .B0 (n_4515), .Y (n_4519));
AOI21X1 g61446(.A0 (n_4520), .A1 (n_3284), .B0 (n_4517), .Y (n_4518));
AOI21X1 g61448(.A0 (n_4520), .A1 (n_3311), .B0 (n_4515), .Y (n_4516));
AOI21X1 g61450(.A0 (n_4520), .A1 (n_3281), .B0 (n_4517), .Y (n_4514));
AOI21X1 g61452(.A0 (n_4520), .A1 (n_3279), .B0 (n_4515), .Y (n_4513));
AOI21X1 g61454(.A0 (n_4520), .A1 (n_3277), .B0 (n_4517), .Y (n_4512));
CLKBUFX1 gbuf_d_780(.A(n_4111), .Y(d_out_780));
CLKBUFX1 gbuf_q_780(.A(q_in_780), .Y(g820));
INVX1 g61477(.A (n_4329), .Y (n_4511));
CLKBUFX1 gbuf_d_781(.A(n_4264), .Y(d_out_781));
CLKBUFX1 gbuf_q_781(.A(q_in_781), .Y(gbuf114));
CLKBUFX1 gbuf_d_782(.A(n_4261), .Y(d_out_782));
CLKBUFX1 gbuf_q_782(.A(q_in_782), .Y(gbuf116));
CLKBUFX1 gbuf_d_783(.A(n_4263), .Y(d_out_783));
CLKBUFX1 gbuf_q_783(.A(q_in_783), .Y(gbuf115));
INVX1 g61479(.A (n_4328), .Y (n_4510));
INVX1 g61481(.A (n_4326), .Y (n_4509));
INVX1 g61483(.A (n_4325), .Y (n_4508));
NOR2X1 g63462(.A (n_4282), .B (n_4464), .Y (n_5015));
AOI21X1 g61498(.A0 (n_7732), .A1 (n_2799), .B0 (n_5323), .Y (n_4507));
INVX1 g63529(.A (n_8839), .Y (n_4505));
NAND2X1 g63568(.A (n_4503), .B (n_3897), .Y (n_4504));
INVX1 g63648(.A (n_6528), .Y (n_4502));
INVX1 g63649(.A (n_6528), .Y (n_4501));
NAND2X1 g63660(.A (n_4195), .B (g2257), .Y (n_5169));
XOR2X1 g63886(.A (g2120), .B (n_5779), .Y (n_4500));
CLKBUFX1 gbuf_d_784(.A(n_3899), .Y(d_out_784));
CLKBUFX1 gbuf_q_784(.A(q_in_784), .Y(g646));
CLKBUFX1 gbuf_d_785(.A(n_3877), .Y(d_out_785));
CLKBUFX1 gbuf_q_785(.A(q_in_785), .Y(g2727));
CLKBUFX1 gbuf_d_786(.A(n_4025), .Y(d_out_786));
CLKBUFX1 gbuf_qn_786(.A(qn_in_786), .Y(g554));
CLKBUFX1 gbuf_d_787(.A(n_3950), .Y(d_out_787));
CLKBUFX1 gbuf_q_787(.A(q_in_787), .Y(g557));
CLKBUFX1 gbuf_d_788(.A(n_3945), .Y(d_out_788));
CLKBUFX1 gbuf_q_788(.A(q_in_788), .Y(n_3701));
CLKBUFX1 gbuf_d_789(.A(n_3943), .Y(d_out_789));
CLKBUFX1 gbuf_q_789(.A(q_in_789), .Y(g2584));
INVX2 g63961(.A (n_4497), .Y (n_4763));
INVX1 g63962(.A (n_4497), .Y (n_4498));
INVX1 g63991(.A (n_8825), .Y (n_9661));
INVX1 g64036(.A (n_9431), .Y (n_4486));
INVX2 g64040(.A (n_4483), .Y (n_4718));
INVX1 g64041(.A (n_4483), .Y (n_4484));
CLKBUFX1 gbuf_d_790(.A(n_4023), .Y(d_out_790));
CLKBUFX1 gbuf_qn_790(.A(qn_in_790), .Y(g2628));
OAI21X1 g61696(.A0 (n_2540), .A1 (n_2410), .B0 (n_7328), .Y (n_4480));
OAI21X1 g61697(.A0 (n_2525), .A1 (n_2292), .B0 (n_7732), .Y (n_4479));
MX2X1 g63875(.A (n_365), .B (g1471), .S0 (n_4004), .Y (n_5171));
NAND2X2 g64208(.A (n_4477), .B (n_4242), .Y (n_4478));
NAND2X1 g64213(.A (n_4227), .B (n_4193), .Y (n_4476));
NAND2X1 g64214(.A (n_4226), .B (n_3804), .Y (n_4475));
NAND3X1 g61751(.A (n_7732), .B (n_4064), .C (n_5323), .Y (n_4474));
NAND3X1 g64298(.A (n_3651), .B (n_4116), .C (g3229), .Y (n_4471));
NAND2X1 g64364(.A (n_4233), .B (n_79), .Y (n_4469));
NAND2X2 g64368(.A (n_4231), .B (n_8759), .Y (n_4468));
NAND2X1 g64370(.A (n_4230), .B (n_293), .Y (n_4466));
NAND2X1 g64375(.A (n_4229), .B (n_78), .Y (n_4465));
NOR2X1 g64392(.A (n_4009), .B (n_4464), .Y (n_4732));
NAND3X1 g64443(.A (n_3685), .B (n_3361), .C (g3229), .Y (n_4867));
NAND3X1 g64454(.A (n_3648), .B (n_3415), .C (g3229), .Y (n_4925));
MX2X1 g63851(.A (n_454), .B (g1486), .S0 (n_4463), .Y (n_5368));
MX2X1 g64515(.A (n_26), .B (n_6947), .S0 (n_6626), .Y (n_4462));
MX2X1 g64532(.A (n_4112), .B (g862), .S0 (n_4460), .Y (n_4461));
MX2X1 g64534(.A (n_4110), .B (g859), .S0 (n_4460), .Y (n_4459));
MX2X1 g64540(.A (n_4464), .B (g865), .S0 (n_4460), .Y (n_4458));
XOR2X1 g64564(.A (g_26529), .B (n_3790), .Y (n_4457));
XOR2X1 g64565(.A (g_21927), .B (n_4455), .Y (n_4456));
INVX1 g64571(.A (n_9535), .Y (n_4454));
INVX1 g64576(.A (n_4451), .Y (n_4923));
OR2X1 g64690(.A (n_3524), .B (g3229), .Y (n_4449));
NOR2X1 g64728(.A (n_8641), .B (n_4206), .Y (n_4448));
OAI21X1 g64778(.A0 (n_2474), .A1 (n_2378), .B0 (n_3938), .Y (n_4631));
AOI21X1 g64788(.A0 (n_2604), .A1 (n_2061), .B0 (n_3928), .Y (n_4630));
INVX1 g64951(.A (n_4446), .Y (n_5480));
INVX1 g64958(.A (n_9437), .Y (n_4627));
OAI21X1 g65026(.A0 (g1033), .A1 (n_3336), .B0 (n_2763), .Y (n_5680));
INVX1 g65107(.A (n_5947), .Y (n_4444));
CLKBUFX1 gbuf_d_791(.A(n_3952), .Y(d_out_791));
CLKBUFX1 gbuf_q_791(.A(q_in_791), .Y(g2040));
INVX1 g65175(.A (n_4441), .Y (n_4618));
NOR2X1 g62104(.A (n_3875), .B (n_4967), .Y (n_4439));
INVX1 g65205(.A (n_4827), .Y (n_4615));
INVX1 g65221(.A (n_4825), .Y (n_4613));
NAND2X1 g62113(.A (n_4100), .B (g2760), .Y (n_4436));
NOR2X1 g62115(.A (n_3874), .B (n_4963), .Y (n_4435));
INVX1 g65242(.A (n_4433), .Y (n_4610));
INVX2 g62125(.A (n_4698), .Y (n_4894));
NOR2X1 g62158(.A (n_3710), .B (n_3941), .Y (n_4428));
INVX1 g65471(.A (n_4425), .Y (n_4426));
INVX1 g65476(.A (n_4213), .Y (n_4599));
NAND3X1 g65481(.A (n_2195), .B (n_1034), .C (n_3760), .Y (n_4424));
NAND3X1 g65482(.A (n_1031), .B (n_2083), .C (n_3759), .Y (n_4852));
NAND3X1 g65483(.A (n_8277), .B (n_8278), .C (n_3756), .Y (n_4851));
NOR2X1 g62217(.A (n_3867), .B (n_3937), .Y (n_4423));
AOI22X1 g65559(.A0 (n_3763), .A1 (n_4419), .B0 (g1859), .B1 (n_1689),.Y (n_4420));
NOR2X1 g65577(.A (n_275), .B (n_4418), .Y (n_4597));
INVX1 g65582(.A (n_4416), .Y (n_4596));
INVX1 g65684(.A (n_4477), .Y (n_4976));
AOI21X1 g65705(.A0 (n_2267), .A1 (n_4412), .B0 (n_3935), .Y (n_4590));
NAND4X1 g62273(.A (n_2987), .B (n_3578), .C (n_3573), .D (n_3571), .Y(n_4411));
AOI21X1 g62276(.A0 (n_3908), .A1 (n_3930), .B0 (n_3933), .Y (n_4409));
XOR2X1 g65814(.A (g780), .B (n_3761), .Y (n_4403));
MX2X1 g63846(.A (n_4639), .B (n_471), .S0 (n_3997), .Y (n_4769));
NAND3X1 g66051(.A (n_4402), .B (g2156), .C (g2160), .Y (n_4809));
MX2X1 g66105(.A (g1937), .B (g1934), .S0 (n_6626), .Y (n_4401));
MX2X1 g66118(.A (n_5322), .B (g1937), .S0 (n_6626), .Y (n_4400));
NAND2X1 g62478(.A (g1210), .B (g185), .Y (n_4399));
NAND2X1 g62481(.A (g1228), .B (g185), .Y (n_4398));
NOR2X1 g62491(.A (n_4052), .B (n_5181), .Y (n_4397));
INVX1 g66221(.A (n_4174), .Y (n_4395));
INVX1 g66224(.A (n_4173), .Y (n_4394));
INVX1 g66269(.A (n_4584), .Y (n_4393));
NOR2X1 g66303(.A (g1063), .B (n_3336), .Y (n_4392));
NAND2X1 g66347(.A (g1627), .B (n_7800), .Y (n_4390));
OAI21X1 g62545(.A0 (n_3713), .A1 (n_4351), .B0 (n_3898), .Y (n_4389));
INVX1 g62548(.A (n_4388), .Y (n_4815));
OAI21X1 g62550(.A0 (n_3563), .A1 (n_3882), .B0 (n_3883), .Y (n_4387));
NAND2X1 g66391(.A (g1618), .B (n_7800), .Y (n_9625));
NAND2X1 g66408(.A (g1582), .B (n_7800), .Y (n_4385));
NAND2X1 g66423(.A (g1609), .B (n_7800), .Y (n_4384));
NAND2X1 g66443(.A (g1654), .B (n_7800), .Y (n_8216));
AOI22X1 g62563(.A0 (n_3708), .A1 (n_3684), .B0 (n_4104), .B1(n_3890), .Y (n_4382));
AOI22X1 g62564(.A0 (n_3704), .A1 (n_3524), .B0 (n_4102), .B1(n_4380), .Y (n_4381));
INVX1 g66473(.A (n_4138), .Y (n_4379));
MX2X1 g62599(.A (n_2809), .B (g2208), .S0 (n_4562), .Y (n_4378));
AOI22X1 g62604(.A0 (n_3720), .A1 (n_3651), .B0 (n_4376), .B1(n_4332), .Y (n_4377));
AOI22X1 g62606(.A0 (n_3715), .A1 (n_3848), .B0 (n_4374), .B1(n_4115), .Y (n_4375));
MX2X1 g62663(.A (n_4368), .B (g2205), .S0 (n_4562), .Y (n_4369));
MX2X1 g62666(.A (n_436), .B (g2217), .S0 (n_4562), .Y (n_4367));
MX2X1 g62667(.A (n_2719), .B (g2220), .S0 (n_4562), .Y (n_4366));
MX2X1 g62675(.A (n_2716), .B (g2223), .S0 (n_4562), .Y (n_4365));
MX2X1 g62679(.A (n_385), .B (g2226), .S0 (n_4562), .Y (n_4364));
CLKBUFX1 gbuf_d_792(.A(n_4049), .Y(d_out_792));
CLKBUFX1 gbuf_q_792(.A(q_in_792), .Y(g728));
AOI22X1 g62685(.A0 (n_3707), .A1 (n_4053), .B0 (n_4362), .B1(n_4082), .Y (n_4363));
AOI22X1 g62697(.A0 (n_2212), .A1 (n_3359), .B0 (n_4343), .B1(n_4360), .Y (n_4361));
OAI21X1 g62754(.A0 (n_4543), .A1 (g805), .B0 (n_3887), .Y (n_4359));
OAI21X1 g62785(.A0 (n_4543), .A1 (n_763), .B0 (n_3888), .Y (n_4358));
CLKBUFX1 gbuf_d_793(.A(n_4048), .Y(d_out_793));
CLKBUFX1 gbuf_q_793(.A(q_in_793), .Y(g729));
INVX1 g62815(.A (n_4356), .Y (n_4357));
CLKBUFX1 gbuf_d_794(.A(n_4047), .Y(d_out_794));
CLKBUFX1 gbuf_q_794(.A(q_in_794), .Y(g730));
NAND3X1 g63032(.A (n_3848), .B (n_4355), .C (g3229), .Y (n_5787));
NOR2X1 g63034(.A (n_4088), .B (n_4975), .Y (n_6565));
NAND3X1 g63036(.A (n_1662), .B (n_2211), .C (n_3830), .Y (n_4354));
NAND3X1 g63042(.A (n_3363), .B (n_1532), .C (n_4355), .Y (n_4353));
NAND3X1 g63047(.A (n_4351), .B (n_1766), .C (n_4277), .Y (n_4352));
NAND2X1 g63051(.A (n_4975), .B (g1511), .Y (n_4350));
NAND2X1 g63057(.A (n_4975), .B (g1529), .Y (n_4349));
NAND2X1 g63061(.A (n_4975), .B (g1535), .Y (n_4348));
NAND2X1 g63065(.A (n_4975), .B (g1538), .Y (n_4347));
NAND2X1 g63152(.A (n_4975), .B (g1532), .Y (n_4346));
NAND3X1 g63161(.A (n_1662), .B (n_4343), .C (n_4094), .Y (n_4345));
CLKBUFX1 gbuf_d_795(.A(n_3948), .Y(d_out_795));
CLKBUFX1 gbuf_q_795(.A(q_in_795), .Y(n_655));
OR4X1 g63191(.A (n_3534), .B (n_1536), .C (n_1370), .D (n_3663), .Y(n_4342));
NAND4X1 g63231(.A (n_4020), .B (n_4096), .C (n_3896), .D (n_4351), .Y(n_4341));
CLKBUFX1 gbuf_d_796(.A(n_3942), .Y(d_out_796));
CLKBUFX1 gbuf_q_796(.A(q_in_796), .Y(g1346));
NAND4X1 g63253(.A (n_3828), .B (n_3648), .C (n_3881), .D (n_3882), .Y(n_4338));
OAI21X1 g63264(.A0 (n_3536), .A1 (n_3533), .B0 (n_4335), .Y (n_4337));
NAND4X1 g61384(.A (n_2964), .B (n_3794), .C (n_2960), .D (n_3127), .Y(n_4334));
AOI22X1 g63267(.A0 (n_3849), .A1 (n_1728), .B0 (n_4332), .B1(n_4355), .Y (n_4333));
NAND4X1 g61401(.A (n_3117), .B (n_3792), .C (n_3298), .D (n_3121), .Y(n_4331));
XOR2X1 g63291(.A (n_3203), .B (n_4073), .Y (n_4330));
AOI21X1 g61478(.A0 (n_4044), .A1 (n_4289), .B0 (n_7273), .Y (n_4329));
AOI21X1 g61480(.A0 (n_4044), .A1 (n_4287), .B0 (n_7271), .Y (n_4328));
AOI21X1 g61482(.A0 (n_4044), .A1 (n_4285), .B0 (n_7273), .Y (n_4326));
AOI21X1 g61484(.A0 (n_4044), .A1 (n_4283), .B0 (n_7271), .Y (n_4325));
INVX1 g61485(.A (n_4076), .Y (n_4324));
INVX1 g61487(.A (n_4075), .Y (n_4323));
INVX1 g61489(.A (n_4072), .Y (n_4322));
INVX1 g61492(.A (n_4069), .Y (n_4321));
INVX1 g61494(.A (n_4068), .Y (n_4320));
AND2X1 g63469(.A (g3229), .B (n_3845), .Y (n_4319));
AOI21X1 g61496(.A0 (n_7732), .A1 (n_2626), .B0 (n_4317), .Y (n_4318));
NAND3X1 g63576(.A (n_3651), .B (n_3628), .C (n_1532), .Y (n_4315));
AND2X1 g63650(.A (n_4194), .B (g2257), .Y (n_6528));
MX2X1 g63863(.A (n_2719), .B (g2180), .S0 (n_4312), .Y (n_5184));
NAND4X1 g63905(.A (n_3651), .B (n_3848), .C (n_1532), .D (n_1665), .Y(n_4311));
CLKBUFX1 gbuf_d_797(.A(n_3732), .Y(d_out_797));
CLKBUFX1 gbuf_q_797(.A(q_in_797), .Y(g1339));
MX2X1 g63937(.A (g2807), .B (n_4515), .S0 (n_5181), .Y (n_4309));
MX2X1 g63956(.A (n_4517), .B (g2802), .S0 (n_4302), .Y (n_4308));
MX2X1 g63957(.A (n_4517), .B (g2803), .S0 (n_4300), .Y (n_4306));
MX2X1 g63958(.A (g2804), .B (n_4517), .S0 (n_5181), .Y (n_4305));
MX2X1 g63959(.A (n_4515), .B (g2805), .S0 (n_4302), .Y (n_4304));
MX2X1 g63960(.A (n_4515), .B (g2806), .S0 (n_4300), .Y (n_4301));
NAND2X2 g63963(.A (n_3846), .B (n_3682), .Y (n_4497));
NAND2X2 g64042(.A (n_3853), .B (n_3854), .Y (n_4483));
XOR2X1 g64091(.A (g780), .B (n_8411), .Y (n_4298));
AND2X1 g61692(.A (n_7328), .B (n_3110), .Y (n_4297));
AND2X1 g61693(.A (n_7328), .B (n_2512), .Y (n_4296));
CLKBUFX1 gbuf_d_798(.A(n_3739), .Y(d_out_798));
CLKBUFX1 gbuf_q_798(.A(q_in_798), .Y(g653));
NAND2X1 g64209(.A (n_9676), .B (n_4003), .Y (n_4295));
NAND2X1 g64215(.A (n_3986), .B (n_3620), .Y (n_4292));
NAND2X1 g64216(.A (n_3987), .B (n_3960), .Y (n_4291));
NAND3X1 g61745(.A (n_7328), .B (n_4289), .C (n_7273), .Y (n_4290));
NAND3X1 g61746(.A (n_7328), .B (n_4287), .C (n_7271), .Y (n_4288));
NAND3X1 g61747(.A (n_7328), .B (n_4285), .C (n_7273), .Y (n_4286));
NAND3X1 g61748(.A (n_7328), .B (n_4283), .C (n_7271), .Y (n_4284));
NAND2X1 g64280(.A (n_4281), .B (n_4280), .Y (n_4282));
NAND3X1 g61750(.A (n_7732), .B (n_4066), .C (n_4317), .Y (n_4279));
NAND2X1 g64301(.A (n_1521), .B (n_4277), .Y (n_4278));
NAND2X1 g64365(.A (n_3996), .B (g1476), .Y (n_4275));
NAND2X1 g64371(.A (n_3993), .B (g2170), .Y (n_4274));
NAND2X1 g64372(.A (n_3992), .B (n_600), .Y (n_4273));
NAND3X1 g64382(.A (n_3822), .B (n_3359), .C (g3229), .Y (n_4270));
NAND2X1 g64383(.A (n_3824), .B (g813), .Y (n_4267));
NAND2X1 g64390(.A (n_3989), .B (g1481), .Y (n_4266));
AOI21X1 g64450(.A0 (n_3953), .A1 (g780), .B0 (g776), .Y (n_4265));
CLKBUFX1 gbuf_d_799(.A(n_3744), .Y(d_out_799));
CLKBUFX1 gbuf_q_799(.A(q_in_799), .Y(g2720));
AOI21X1 g64493(.A0 (n_3633), .A1 (n_4262), .B0 (n_1115), .Y (n_4264));
AOI21X1 g64495(.A0 (n_3629), .A1 (n_4262), .B0 (n_1146), .Y (n_4263));
AOI21X1 g64496(.A0 (n_3632), .A1 (n_4262), .B0 (n_1126), .Y (n_4261));
CLKBUFX1 gbuf_d_800(.A(n_4218), .Y(d_out_800));
CLKBUFX1 gbuf_q_800(.A(q_in_800), .Y(g1193));
INVX1 g64560(.A (n_4259), .Y (n_4760));
INVX1 g64561(.A (n_4259), .Y (n_9662));
MX2X1 g64578(.A (g2195), .B (n_447), .S0 (n_8641), .Y (n_4451));
INVX2 g64583(.A (n_4256), .Y (n_4729));
NOR2X1 g64598(.A (n_3625), .B (g3229), .Y (n_4503));
NOR2X1 g64602(.A (n_3415), .B (g3229), .Y (n_4789));
NAND2X1 g64621(.A (n_9370), .B (n_3959), .Y (n_4671));
NAND2X1 g64637(.A (n_4460), .B (g856), .Y (n_4254));
NOR2X1 g64660(.A (n_3485), .B (g3229), .Y (n_4253));
AOI21X1 g64815(.A0 (n_2483), .A1 (n_3810), .B0 (n_3762), .Y (n_5818));
NAND2X1 g64925(.A (n_3711), .B (n_2770), .Y (n_7000));
OAI21X1 g64952(.A0 (n_2476), .A1 (n_9438), .B0 (n_3725), .Y (n_4446));
OAI21X1 g65005(.A0 (g2253), .A1 (n_7809), .B0 (n_2916), .Y (n_4246));
CLKBUFX1 g65108(.A (n_4242), .Y (n_5947));
AOI22X1 g65176(.A0 (n_2610), .A1 (n_3810), .B0 (g1131), .B1 (n_3808),.Y (n_4441));
NAND2X1 g62101(.A (n_3900), .B (g1372), .Y (n_4239));
CLKBUFX1 g65192(.A (n_4237), .Y (n_4900));
INVX1 g65193(.A (n_4237), .Y (n_4236));
NAND2X1 g62107(.A (n_3902), .B (g2066), .Y (n_4234));
INVX1 g65206(.A (n_4233), .Y (n_4827));
INVX1 g65222(.A (n_4231), .Y (n_4825));
INVX1 g65227(.A (n_4230), .Y (n_5162));
INVX1 g65235(.A (n_4756), .Y (n_4434));
INVX1 g65243(.A (n_4229), .Y (n_4433));
INVX1 g65249(.A (n_4228), .Y (n_4432));
INVX1 g65254(.A (n_4227), .Y (n_4676));
INVX1 g65258(.A (n_4226), .Y (n_4678));
INVX2 g62126(.A (n_4520), .Y (n_4698));
AOI22X1 g65290(.A0 (n_2609), .A1 (n_4604), .B0 (g2498), .B1 (g2476),.Y (n_6106));
AOI22X1 g65315(.A0 (n_2908), .A1 (n_4604), .B0 (g2510), .B1 (g2476),.Y (n_5155));
XOR2X1 g65375(.A (g797), .B (n_3616), .Y (n_4221));
XOR2X1 g65376(.A (g789), .B (n_3615), .Y (n_4220));
XOR2X1 g65377(.A (g785), .B (n_3614), .Y (n_4219));
NAND2X1 g62187(.A (n_4218), .B (n_5270), .Y (n_5993));
NAND2X1 g62190(.A (n_4218), .B (g6750), .Y (n_5990));
NAND2X1 g62192(.A (n_4218), .B (g6944), .Y (n_5988));
NOR2X1 g65441(.A (n_3767), .B (n_1157), .Y (n_4216));
OAI21X1 g65452(.A0 (g2225), .A1 (n_3770), .B0 (n_3772), .Y (n_4645));
NAND3X1 g65454(.A (n_9692), .B (n_9693), .C (n_3606), .Y (n_4214));
NAND3X1 g65458(.A (n_923), .B (n_2092), .C (n_3605), .Y (n_4635));
NOR2X1 g65459(.A (n_2915), .B (n_7800), .Y (n_4877));
NOR2X1 g65472(.A (n_3774), .B (n_1023), .Y (n_4425));
NAND3X1 g65474(.A (n_1022), .B (n_2067), .C (n_3603), .Y (n_4640));
NAND3X1 g65477(.A (n_1021), .B (n_3592), .C (n_2242), .Y (n_4213));
NAND2X1 g65478(.A (n_3793), .B (n_3588), .Y (n_5077));
NOR2X1 g65491(.A (n_3771), .B (n_1092), .Y (n_4211));
NOR2X1 g65492(.A (n_3769), .B (n_1129), .Y (n_4210));
CLKBUFX1 g62225(.A (n_4209), .Y (n_4693));
CLKBUFX1 g62226(.A (n_4209), .Y (n_4740));
NAND3X1 g65523(.A (n_2231), .B (n_1016), .C (n_3602), .Y (n_4208));
INVX1 g62233(.A (n_3980), .Y (n_4207));
AOI22X1 g65560(.A0 (n_3607), .A1 (g1867), .B0 (g1868), .B1 (n_1689),.Y (n_4205));
INVX1 g62247(.A (n_3970), .Y (n_4203));
INVX1 g65584(.A (n_4202), .Y (n_4416));
INVX1 g65588(.A (n_4653), .Y (n_6603));
AOI22X1 g65603(.A0 (n_3595), .A1 (g1861), .B0 (g1865), .B1 (n_1689),.Y (n_4201));
INVX1 g65706(.A (n_4194), .Y (n_4195));
INVX2 g65711(.A (n_4193), .Y (n_4410));
INVX1 g65733(.A (n_9369), .Y (n_4192));
INVX1 g66043(.A (n_4418), .Y (n_4582));
NOR2X1 g62426(.A (n_3676), .B (n_3729), .Y (n_4188));
NOR2X1 g62446(.A (n_3861), .B (n_4967), .Y (n_4187));
NOR2X1 g62449(.A (n_3860), .B (n_5372), .Y (n_4185));
NAND2X1 g62487(.A (g2598), .B (g185), .Y (n_4183));
NOR2X1 g62490(.A (n_3837), .B (n_3572), .Y (n_4182));
NOR2X1 g62497(.A (n_3859), .B (n_4963), .Y (n_4181));
OR2X1 g66214(.A (g_19472), .B (n_9314), .Y (n_4179));
OR2X1 g66216(.A (g_28702), .B (n_9314), .Y (n_4178));
OR2X1 g66219(.A (n_0), .B (n_4172), .Y (n_4176));
OR2X1 g66220(.A (g_25878), .B (n_4172), .Y (n_4175));
NOR2X1 g66222(.A (g_5095), .B (n_9314), .Y (n_4174));
NOR2X1 g66225(.A (g_22340), .B (n_4172), .Y (n_4173));
OR2X1 g66230(.A (n_14), .B (n_4172), .Y (n_4171));
OR2X1 g66232(.A (n_9316), .B (n_4172), .Y (n_4170));
NOR2X1 g66237(.A (n_222), .B (n_4172), .Y (n_4169));
NAND2X1 g66241(.A (g933), .B (n_4162), .Y (n_4168));
NOR2X1 g66270(.A (n_3873), .B (n_7800), .Y (n_4584));
NAND2X1 g66272(.A (g2276), .B (n_7809), .Y (n_9603));
OR2X1 g66275(.A (g_13546), .B (n_9314), .Y (n_4164));
NAND2X1 g66291(.A (g915), .B (n_4162), .Y (n_4163));
NOR2X1 g66302(.A (g402), .B (n_5004), .Y (n_4161));
OR2X1 g66316(.A (n_98), .B (n_4172), .Y (n_4160));
AOI21X1 g62538(.A0 (n_3508), .A1 (g2746), .B0 (g2740), .Y (n_4159));
NOR2X1 g66341(.A (g1559), .B (n_7800), .Y (n_4155));
OAI21X1 g62546(.A0 (n_3702), .A1 (n_4056), .B0 (n_3396), .Y (n_4605));
OR2X1 g66353(.A (g1701), .B (n_5008), .Y (n_4153));
INVX1 g66354(.A (n_4402), .Y (n_4152));
AOI22X1 g62549(.A0 (n_3696), .A1 (n_3636), .B0 (n_4151), .B1(n_4515), .Y (n_4388));
OR2X1 g66397(.A (g1783), .B (n_5008), .Y (n_4149));
OR2X1 g66406(.A (n_96), .B (n_4172), .Y (n_4147));
NAND2X1 g66407(.A (g2312), .B (n_7809), .Y (n_9605));
OR2X1 g66411(.A (g1695), .B (n_5008), .Y (n_4145));
NAND2X1 g66412(.A (g2321), .B (n_7809), .Y (n_8248));
NAND2X1 g66414(.A (g888), .B (n_4162), .Y (n_4143));
NAND2X1 g66416(.A (g2348), .B (n_7809), .Y (n_8263));
NAND2X1 g66422(.A (g924), .B (n_4162), .Y (n_4141));
NOR2X1 g66446(.A (g2501), .B (n_4576), .Y (n_4140));
NOR2X1 g66458(.A (n_319), .B (n_4172), .Y (n_4139));
NOR2X1 g66474(.A (g_27846), .B (n_9314), .Y (n_4138));
OR2X1 g66476(.A (g_16936), .B (n_5004), .Y (n_4137));
NAND2X1 g66478(.A (g2303), .B (n_7809), .Y (n_4135));
NAND2X1 g66480(.A (g960), .B (n_4162), .Y (n_8272));
OR2X1 g66488(.A (g1702), .B (n_5008), .Y (n_4133));
AOI22X1 g62625(.A0 (n_3565), .A1 (n_3822), .B0 (n_4127), .B1(n_3716), .Y (n_4128));
AOI22X1 g62693(.A0 (n_1767), .A1 (n_4116), .B0 (n_4091), .B1(n_4115), .Y (n_4117));
AOI21X1 g62704(.A0 (n_4102), .A1 (n_2032), .B0 (n_3738), .Y (n_4114));
MX2X1 g62767(.A (n_4112), .B (g817), .S0 (n_4543), .Y (n_4113));
MX2X1 g62770(.A (n_4110), .B (g820), .S0 (n_4543), .Y (n_4111));
MX2X1 g62773(.A (n_3171), .B (g829), .S0 (n_4543), .Y (n_4109));
MX2X1 g62775(.A (n_3169), .B (g832), .S0 (n_4543), .Y (n_4108));
MX2X1 g62777(.A (n_3167), .B (g835), .S0 (n_4543), .Y (n_4107));
MX2X1 g62782(.A (n_3164), .B (g841), .S0 (n_4543), .Y (n_4106));
OAI33X1 g62802(.A0 (n_3531), .A1 (n_3530), .A2 (n_3419), .B0(n_4104), .B1 (n_3677), .B2 (n_1954), .Y (n_4105));
OAI33X1 g62803(.A0 (n_4053), .A1 (n_3382), .A2 (n_2031), .B0(n_4102), .B1 (n_3527), .B2 (n_2036), .Y (n_4103));
XOR2X1 g62807(.A (n_3263), .B (n_3700), .Y (n_4872));
INVX1 g62816(.A (n_4100), .Y (n_4101));
CLKBUFX1 gbuf_d_801(.A(gbuf54), .Y(d_out_801));
CLKBUFX1 gbuf_q_801(.A(q_in_801), .Y(g524));
CLKBUFX1 gbuf_d_802(.A(gbuf64), .Y(d_out_802));
CLKBUFX1 gbuf_q_802(.A(q_in_802), .Y(g542));
CLKBUFX1 gbuf_d_803(.A(gbuf211), .Y(d_out_803));
CLKBUFX1 gbuf_q_803(.A(q_in_803), .Y(g2616));
NAND2X1 g62941(.A (n_3625), .B (n_4098), .Y (n_4099));
NAND3X1 g62945(.A (n_4096), .B (n_4116), .C (n_3870), .Y (n_4097));
NAND3X1 g63017(.A (n_3863), .B (n_4094), .C (n_4127), .Y (n_4095));
NAND2X1 g63030(.A (n_4562), .B (g2229), .Y (n_4093));
NAND3X1 g63043(.A (n_4351), .B (n_4091), .C (n_3712), .Y (n_4092));
NAND3X1 g63067(.A (n_1662), .B (n_3845), .C (n_4085), .Y (n_4090));
NAND2X1 g63069(.A (n_3717), .B (n_3865), .Y (n_4089));
NOR2X1 g63088(.A (n_4088), .B (n_4562), .Y (n_6478));
NAND2X1 g63106(.A (n_4562), .B (g2232), .Y (n_4087));
NAND4X1 g63234(.A (n_3827), .B (n_3685), .C (n_4085), .D (n_1662), .Y(n_4086));
NAND3X1 g63250(.A (n_4116), .B (n_3363), .C (n_3714), .Y (n_4084));
AOI22X1 g63300(.A0 (n_3669), .A1 (n_2035), .B0 (n_4082), .B1(n_4081), .Y (n_4083));
XOR2X1 g63301(.A (n_3143), .B (n_4059), .Y (n_4080));
AOI22X1 g63351(.A0 (n_3671), .A1 (n_4078), .B0 (n_4077), .B1(n_3576), .Y (n_4079));
CLKBUFX1 gbuf_d_804(.A(n_3742), .Y(d_out_804));
CLKBUFX1 gbuf_q_804(.A(q_in_804), .Y(g2033));
CLKBUFX1 gbuf_d_805(.A(gbuf151), .Y(d_out_805));
CLKBUFX1 gbuf_q_805(.A(q_in_805), .Y(gbuf152));
CLKBUFX1 gbuf_d_806(.A(gbuf161), .Y(d_out_806));
CLKBUFX1 gbuf_q_806(.A(q_in_806), .Y(gbuf162));
AOI21X1 g61486(.A0 (n_9630), .A1 (n_3544), .B0 (n_4317), .Y (n_4076));
AOI21X1 g61488(.A0 (n_9630), .A1 (n_2990), .B0 (n_5323), .Y (n_4075));
NOR2X1 g63451(.A (n_4073), .B (n_163), .Y (n_4356));
AOI21X1 g61490(.A0 (n_9630), .A1 (n_3542), .B0 (n_4317), .Y (n_4072));
AOI21X1 g61491(.A0 (n_9630), .A1 (n_2625), .B0 (n_5323), .Y (n_4071));
AOI21X1 g61493(.A0 (n_9630), .A1 (n_3540), .B0 (n_4317), .Y (n_4069));
AOI21X1 g61495(.A0 (n_9631), .A1 (n_2816), .B0 (n_5323), .Y (n_4068));
AOI21X1 g61497(.A0 (n_9631), .A1 (n_4066), .B0 (n_4317), .Y (n_4067));
AOI21X1 g61499(.A0 (n_9631), .A1 (n_4064), .B0 (n_5323), .Y (n_4065));
AND2X1 g63551(.A (n_5420), .B (n_5786), .Y (n_5615));
NOR2X1 g63561(.A (n_5420), .B (g996), .Y (n_5817));
NAND2X1 g63601(.A (n_4073), .B (n_3674), .Y (n_4063));
NOR2X1 g66349(.A (g1698), .B (n_5008), .Y (n_4062));
NAND2X1 g63681(.A (n_4061), .B (n_2416), .Y (n_6543));
NAND2X1 g63732(.A (n_4059), .B (n_3835), .Y (n_4060));
AOI21X1 g63779(.A0 (n_4737), .A1 (n_3701), .B0 (n_4056), .Y (n_4058));
OR2X1 g63785(.A (n_4055), .B (n_7800), .Y (n_4975));
CLKBUFX1 gbuf_d_807(.A(n_3581), .Y(d_out_807));
CLKBUFX1 gbuf_q_807(.A(q_in_807), .Y(g2026));
NAND4X1 g63912(.A (n_4053), .B (n_3736), .C (n_4027), .D (n_3735), .Y(n_4054));
CLKBUFX1 gbuf_d_808(.A(n_3692), .Y(d_out_808));
CLKBUFX1 gbuf_q_808(.A(q_in_808), .Y(g2111));
CLKBUFX1 gbuf_d_809(.A(n_3703), .Y(d_out_809));
CLKBUFX1 gbuf_q_809(.A(q_in_809), .Y(g2707));
CLKBUFX1 gbuf_d_810(.A(n_3655), .Y(d_out_810));
CLKBUFX1 gbuf_q_810(.A(q_in_810), .Y(g640));
NAND3X1 g63816(.A (n_3239), .B (n_3534), .C (g3229), .Y (n_4335));
XOR2X1 g63935(.A (g2746), .B (n_3836), .Y (n_4052));
AOI21X1 g63813(.A0 (n_4517), .A1 (n_4050), .B0 (n_3795), .Y (n_4051));
MX2X1 g63949(.A (n_4737), .B (g728), .S0 (n_3554), .Y (n_4049));
MX2X1 g63950(.A (n_4737), .B (g729), .S0 (n_3552), .Y (n_4048));
MX2X1 g63951(.A (g730), .B (n_4737), .S0 (n_5372), .Y (n_4047));
AND2X1 g61688(.A (n_4044), .B (n_3114), .Y (n_4046));
AND2X1 g61689(.A (n_4044), .B (n_2993), .Y (n_4045));
AND2X1 g61690(.A (n_4044), .B (n_3112), .Y (n_4043));
AND2X1 g61691(.A (n_4044), .B (n_2938), .Y (n_4042));
CLKBUFX1 gbuf_d_811(.A(n_3694), .Y(d_out_811));
CLKBUFX1 gbuf_q_811(.A(q_in_811), .Y(g1415));
NOR2X1 g64200(.A (n_2652), .B (n_4037), .Y (n_4039));
NOR2X1 g64207(.A (n_2623), .B (n_4037), .Y (n_4038));
AND2X1 g61749(.A (n_3686), .B (n_9631), .Y (n_4035));
NAND2X1 g64307(.A (n_3823), .B (n_763), .Y (n_4034));
CLKBUFX1 gbuf_d_812(.A(n_3695), .Y(d_out_812));
CLKBUFX1 gbuf_q_812(.A(q_in_812), .Y(g1414));
NAND2X1 g64341(.A (n_3820), .B (n_656), .Y (n_4031));
NOR2X1 g64402(.A (n_3864), .B (n_3829), .Y (n_4029));
NOR2X1 g64412(.A (n_4027), .B (n_3657), .Y (n_4028));
CLKBUFX1 gbuf_d_813(.A(n_3579), .Y(d_out_813));
CLKBUFX1 gbuf_q_813(.A(q_in_813), .Y(g1332));
MX2X1 g64516(.A (n_23), .B (n_6947), .S0 (n_4601), .Y (n_4025));
MX2X1 g64517(.A (n_6947), .B (n_103), .S0 (n_3448), .Y (n_4023));
MX2X1 g64562(.A (n_763), .B (g813), .S0 (n_3630), .Y (n_4259));
MX2X1 g64585(.A (n_656), .B (g809), .S0 (n_4015), .Y (n_4256));
NOR2X1 g64601(.A (n_3239), .B (g3229), .Y (n_4569));
NAND2X1 g64605(.A (n_4104), .B (g3229), .Y (n_4021));
NOR2X1 g64663(.A (n_4116), .B (n_3625), .Y (n_4020));
NOR2X1 g64685(.A (n_3530), .B (g3229), .Y (n_4019));
OR2X1 g64689(.A (n_3684), .B (g3229), .Y (n_4018));
NOR2X1 g64693(.A (n_3382), .B (g3229), .Y (n_4017));
NOR2X1 g64723(.A (n_4015), .B (n_4014), .Y (n_4016));
INVX1 g64988(.A (n_4010), .Y (n_4011));
AOI21X1 g64990(.A0 (n_2482), .A1 (n_3816), .B0 (n_3596), .Y (n_4009));
INVX1 g65101(.A (n_5414), .Y (n_4245));
INVX1 g65105(.A (n_4004), .Y (n_4244));
INVX1 g65109(.A (n_4003), .Y (n_4242));
INVX1 g65154(.A (n_4000), .Y (n_4240));
INVX1 g65194(.A (n_8982), .Y (n_4237));
INVX1 g65199(.A (n_3997), .Y (n_5163));
INVX1 g65207(.A (n_3996), .Y (n_4233));
INVX1 g65215(.A (n_3994), .Y (n_4757));
INVX2 g65223(.A (n_3993), .Y (n_4231));
INVX1 g65228(.A (n_3992), .Y (n_4230));
INVX1 g65230(.A (n_5779), .Y (n_3991));
INVX1 g65236(.A (n_9284), .Y (n_4756));
INVX1 g65244(.A (n_3989), .Y (n_4229));
INVX1 g65250(.A (n_3988), .Y (n_4228));
INVX1 g65255(.A (n_3987), .Y (n_4227));
INVX1 g65259(.A (n_3986), .Y (n_4226));
NAND2X2 g62129(.A (n_3608), .B (n_3139), .Y (n_4520));
XOR2X1 g65374(.A (g801), .B (n_3480), .Y (n_3981));
OR2X1 g65490(.A (n_3613), .B (n_1144), .Y (n_4450));
NAND3X1 g62227(.A (n_3609), .B (n_3109), .C (n_4687), .Y (n_4209));
NAND4X1 g62234(.A (n_2962), .B (n_3556), .C (n_3294), .D (n_3295), .Y(n_3980));
AOI22X1 g65538(.A0 (n_3449), .A1 (n_3978), .B0 (g2553), .B1 (n_1596),.Y (n_3979));
AOI22X1 g65547(.A0 (n_3445), .A1 (g480), .B0 (g484), .B1 (n_1911), .Y(n_3977));
INVX1 g65552(.A (n_3975), .Y (n_4206));
AOI22X1 g65565(.A0 (n_3459), .A1 (g486), .B0 (g487), .B1 (n_1911), .Y(n_3974));
AOI22X1 g65573(.A0 (n_3442), .A1 (n_3971), .B0 (g478), .B1 (n_1911),.Y (n_3972));
NAND4X1 g62248(.A (n_3403), .B (n_3156), .C (n_3399), .D (n_3116), .Y(n_3970));
NAND3X1 g65585(.A (n_949), .B (n_2075), .C (n_3461), .Y (n_4202));
NAND3X1 g65589(.A (n_940), .B (n_2076), .C (n_3451), .Y (n_4653));
AOI22X1 g65605(.A0 (n_3438), .A1 (g2555), .B0 (g2559), .B1 (n_1596),.Y (n_3968));
AOI22X1 g65606(.A0 (n_3465), .A1 (g2561), .B0 (g2562), .B1 (n_1596),.Y (n_3966));
INVX2 g65686(.A (n_9675), .Y (n_4477));
INVX1 g65696(.A (n_4672), .Y (n_4534));
OAI21X1 g65707(.A0 (n_2363), .A1 (n_2407), .B0 (n_3610), .Y (n_4194));
INVX2 g65712(.A (n_3960), .Y (n_4193));
INVX1 g65759(.A (n_3959), .Y (n_6448));
INVX1 g65899(.A (n_3955), .Y (n_3956));
NAND3X1 g65941(.A (n_8241), .B (n_953), .C (n_8242), .Y (n_3954));
NAND3X1 g66044(.A (n_3953), .B (g776), .C (g780), .Y (n_4418));
NOR2X1 g62444(.A (n_3666), .B (n_3429), .Y (n_3952));
NAND3X1 g62451(.A (n_3291), .B (n_3550), .C (n_3292), .Y (n_3951));
MX2X1 g66109(.A (g557), .B (g554), .S0 (n_4601), .Y (n_3950));
OAI22X1 g66110(.A0 (n_103), .A1 (n_3448), .B0 (n_2863), .B1 (n_300),.Y (n_3948));
MX2X1 g66117(.A (n_3701), .B (g557), .S0 (n_4601), .Y (n_3945));
MX2X1 g66122(.A (n_655), .B (n_4050), .S0 (n_3448), .Y (n_3943));
NOR2X1 g62494(.A (n_3680), .B (n_3425), .Y (n_3942));
AOI21X1 g62523(.A0 (n_3381), .A1 (g2052), .B0 (g2046), .Y (n_3941));
AOI21X1 g62526(.A0 (n_3509), .A1 (g672), .B0 (g666), .Y (n_3940));
OR2X1 g66292(.A (g_24632), .B (n_5004), .Y (n_3939));
OR2X1 g66312(.A (g_18093), .B (n_5004), .Y (n_3938));
AOI21X1 g62541(.A0 (n_3380), .A1 (g1358), .B0 (g1352), .Y (n_3937));
AOI21X1 g62543(.A0 (n_3395), .A1 (n_1951), .B0 (n_3574), .Y (n_3936));
NOR2X1 g66372(.A (g1550), .B (n_7800), .Y (n_3935));
OAI21X1 g62551(.A0 (n_3561), .A1 (n_1536), .B0 (n_3577), .Y (n_3933));
AOI22X1 g62565(.A0 (n_3310), .A1 (n_3533), .B0 (n_2986), .B1(n_3930), .Y (n_3931));
OR2X1 g66477(.A (g1541), .B (n_3467), .Y (n_3929));
NOR2X1 g66481(.A (g_14632), .B (n_5004), .Y (n_3928));
INVX1 g66737(.A (n_4162), .Y (n_3919));
INVX1 g66759(.A (n_7809), .Y (n_3914));
INVX1 g66795(.A (n_5004), .Y (n_6917));
INVX1 g66873(.A (n_4576), .Y (n_6611));
AOI22X1 g62687(.A0 (n_3411), .A1 (n_3393), .B0 (n_3908), .B1(n_3904), .Y (n_3909));
AOI22X1 g62701(.A0 (n_1964), .A1 (n_3515), .B0 (n_3884), .B1(n_3906), .Y (n_3907));
AOI22X1 g62702(.A0 (n_1960), .A1 (n_4078), .B0 (n_3878), .B1(n_3904), .Y (n_3905));
INVX1 g62812(.A (n_3902), .Y (n_3903));
INVX1 g62814(.A (n_3900), .Y (n_3901));
CLKBUFX1 gbuf_d_814(.A(gbuf103), .Y(d_out_814));
CLKBUFX1 gbuf_q_814(.A(q_in_814), .Y(g1210));
CLKBUFX1 gbuf_d_815(.A(gbuf113), .Y(d_out_815));
CLKBUFX1 gbuf_q_815(.A(q_in_815), .Y(g1228));
CLKBUFX1 gbuf_d_816(.A(n_3693), .Y(d_out_816));
CLKBUFX1 gbuf_q_816(.A(q_in_816), .Y(g1416));
NOR2X1 g62947(.A (n_3660), .B (n_5372), .Y (n_3899));
CLKBUFX1 gbuf_d_817(.A(n_3612), .Y(d_out_817));
CLKBUFX1 gbuf_q_817(.A(q_in_817), .Y(g1243));
NAND3X1 g63044(.A (n_4351), .B (n_3897), .C (n_3896), .Y (n_3898));
NAND4X1 g63045(.A (n_4096), .B (n_3848), .C (n_3718), .D (n_1665), .Y(n_3895));
NAND3X1 g63056(.A (n_3842), .B (g3229), .C (n_3893), .Y (n_5424));
NAND2X1 g63066(.A (n_3891), .B (n_3890), .Y (n_3892));
NAND2X1 g63094(.A (n_4543), .B (g850), .Y (n_3889));
CLKBUFX1 gbuf_d_818(.A(n_3690), .Y(d_out_818));
CLKBUFX1 gbuf_q_818(.A(q_in_818), .Y(g2112));
NOR2X1 g63135(.A (n_4088), .B (n_4543), .Y (n_6227));
NAND3X1 g63143(.A (n_3736), .B (n_4081), .C (g3229), .Y (n_5226));
NAND2X1 g63151(.A (n_4543), .B (g844), .Y (n_3888));
NAND2X1 g63177(.A (n_4543), .B (g838), .Y (n_3887));
NAND3X1 g63178(.A (n_3882), .B (n_3884), .C (n_3562), .Y (n_3886));
NAND3X1 g63186(.A (n_3882), .B (n_3721), .C (n_3881), .Y (n_3883));
NAND3X1 g63188(.A (n_3882), .B (n_1963), .C (n_3656), .Y (n_3880));
NAND3X1 g63190(.A (n_1536), .B (n_3878), .C (n_3560), .Y (n_3879));
NOR2X1 g63199(.A (n_3658), .B (n_3476), .Y (n_3877));
NAND2X1 g63205(.A (n_4543), .B (g847), .Y (n_3876));
XOR2X1 g63270(.A (n_2834), .B (n_3724), .Y (n_3875));
XOR2X1 g63332(.A (n_2880), .B (n_3866), .Y (n_3874));
CLKBUFX1 gbuf_d_819(.A(n_3659), .Y(d_out_819));
CLKBUFX1 gbuf_qn_819(.A(qn_in_819), .Y(g1240));
NOR2X1 g63452(.A (n_4059), .B (n_213), .Y (n_4100));
NOR2X1 g66355(.A (n_3873), .B (n_3344), .Y (n_4402));
NOR2X1 g63575(.A (n_3363), .B (n_1755), .Y (n_3872));
CLKBUFX1 gbuf_d_820(.A(n_3688), .Y(d_out_820));
CLKBUFX1 gbuf_q_820(.A(q_in_820), .Y(g2113));
AND2X1 g63704(.A (n_3625), .B (n_3870), .Y (n_3871));
NAND3X1 g63714(.A (n_4053), .B (n_3415), .C (n_4027), .Y (n_3869));
NAND2X1 g63758(.A (n_3866), .B (n_3678), .Y (n_3867));
NAND2X1 g63771(.A (g2257), .B (n_3588), .Y (n_4562));
NAND4X1 g63903(.A (n_3531), .B (n_3842), .C (n_3864), .D (n_3863), .Y(n_3865));
NAND3X1 g63817(.A (n_4078), .B (n_3394), .C (g3229), .Y (n_3862));
CLKBUFX1 gbuf_d_821(.A(n_3551), .Y(d_out_821));
CLKBUFX1 gbuf_q_821(.A(q_in_821), .Y(g733));
XOR2X1 g63929(.A (g2052), .B (n_3665), .Y (n_3861));
XOR2X1 g63932(.A (g672), .B (n_3675), .Y (n_3860));
XOR2X1 g63936(.A (g1358), .B (n_3679), .Y (n_3859));
CLKBUFX1 gbuf_d_822(.A(n_3513), .Y(d_out_822));
CLKBUFX1 gbuf_q_822(.A(q_in_822), .Y(g2714));
CLKBUFX1 gbuf_d_823(.A(n_3856), .Y(d_out_823));
CLKBUFX1 gbuf_q_823(.A(q_in_823), .Y(gbuf151));
CLKBUFX1 gbuf_d_824(.A(n_3855), .Y(d_out_824));
CLKBUFX1 gbuf_q_824(.A(q_in_824), .Y(gbuf161));
CLKBUFX1 gbuf_d_825(.A(n_3553), .Y(d_out_825));
CLKBUFX1 gbuf_q_825(.A(q_in_825), .Y(g732));
NAND2X1 g64180(.A (n_8880), .B (n_8499), .Y (n_3854));
NAND2X1 g64192(.A (n_8881), .B (n_8498), .Y (n_3853));
NOR2X1 g64223(.A (n_4096), .B (n_3363), .Y (n_4374));
NOR2X1 g64229(.A (n_3651), .B (n_4116), .Y (n_4355));
NOR2X1 g64285(.A (n_3651), .B (n_3848), .Y (n_3849));
NAND2X1 g64287(.A (n_3642), .B (g789), .Y (n_3847));
NAND2X1 g64293(.A (n_8878), .B (g797), .Y (n_3846));
NOR2X1 g64340(.A (n_3531), .B (n_3684), .Y (n_4343));
NOR2X1 g64360(.A (n_3531), .B (n_3842), .Y (n_3844));
NAND2X1 g64399(.A (n_3638), .B (n_448), .Y (n_3841));
NAND2X1 g64424(.A (n_8736), .B (n_3171), .Y (n_3840));
NAND2X1 g64432(.A (n_3836), .B (n_3835), .Y (n_3837));
NAND3X1 g64455(.A (n_3509), .B (g672), .C (g666), .Y (n_4073));
INVX1 g64606(.A (n_3833), .Y (n_3834));
NOR2X1 g64610(.A (n_3361), .B (g3229), .Y (n_4726));
INVX1 g64658(.A (n_3829), .Y (n_3830));
NOR2X1 g64661(.A (n_4116), .B (n_3628), .Y (n_4277));
NOR2X1 g64669(.A (n_3515), .B (n_4102), .Y (n_3828));
NOR2X1 g64670(.A (n_3359), .B (n_4104), .Y (n_3827));
INVX1 g64757(.A (n_8492), .Y (n_4280));
INVX1 g64873(.A (n_3825), .Y (n_4281));
INVX1 g64887(.A (n_3823), .Y (n_3824));
INVX1 g64913(.A (n_3820), .Y (n_3821));
AOI21X1 g64989(.A0 (n_2485), .A1 (n_3816), .B0 (n_3450), .Y (n_4010));
AOI21X1 g65000(.A0 (n_2600), .A1 (n_3816), .B0 (n_3447), .Y (n_4061));
INVX1 g65003(.A (n_3814), .Y (n_3815));
INVX1 g65031(.A (n_4312), .Y (n_5778));
AOI22X1 g65084(.A0 (n_2398), .A1 (n_3810), .B0 (g1101), .B1 (n_3808),.Y (n_5420));
INVX1 g65088(.A (n_3646), .Y (n_5201));
AOI22X1 g65102(.A0 (n_2405), .A1 (n_3810), .B0 (g1110), .B1 (n_3808),.Y (n_5414));
NAND2X2 g65106(.A (n_3472), .B (n_2617), .Y (n_4004));
OAI21X1 g65110(.A0 (n_2397), .A1 (n_3781), .B0 (n_3458), .Y (n_4003));
INVX1 g65129(.A (n_8884), .Y (n_4001));
INVX1 g65155(.A (n_3805), .Y (n_4000));
AOI22X1 g65164(.A0 (n_2404), .A1 (n_3810), .B0 (g1122), .B1 (n_3808),.Y (n_4953));
INVX2 g65697(.A (n_3804), .Y (n_4672));
NAND2X2 g65200(.A (n_3460), .B (n_2505), .Y (n_3997));
AOI21X1 g65208(.A0 (n_2311), .A1 (n_8945), .B0 (n_3464), .Y (n_3996));
NAND2X2 g65212(.A (n_3468), .B (n_2507), .Y (n_4463));
NAND2X2 g65216(.A (n_3454), .B (n_2504), .Y (n_3994));
AOI21X1 g65224(.A0 (n_2310), .A1 (n_3799), .B0 (n_3452), .Y (n_3993));
AOI21X1 g65229(.A0 (n_2309), .A1 (n_8945), .B0 (n_3439), .Y (n_3992));
CLKBUFX1 g65231(.A (n_8988), .Y (n_5779));
AOI21X1 g65245(.A0 (n_2307), .A1 (n_8945), .B0 (n_3471), .Y (n_3989));
INVX2 g65251(.A (n_3800), .Y (n_3988));
AOI21X1 g65256(.A0 (n_2312), .A1 (n_8945), .B0 (n_3457), .Y (n_3987));
AOI21X1 g65260(.A0 (n_2304), .A1 (n_3799), .B0 (n_3473), .Y (n_3986));
CLKBUFX1 gbuf_d_826(.A(n_3475), .Y(d_out_826));
CLKBUFX1 gbuf_q_826(.A(q_in_826), .Y(n_3698));
INVX1 g65303(.A (n_4223), .Y (n_3985));
INVX1 g65321(.A (n_4339), .Y (n_3984));
INVX1 g62228(.A (n_3635), .Y (n_3794));
NAND2X1 g65511(.A (n_3793), .B (n_3589), .Y (n_4460));
INVX1 g62231(.A (n_3634), .Y (n_3792));
INVX1 g65554(.A (n_9531), .Y (n_3975));
INVX1 g65591(.A (n_8641), .Y (n_6414));
INVX1 g65595(.A (n_4014), .Y (n_4455));
CLKBUFX3 g62254(.A (n_4044), .Y (n_7328));
CLKBUFX3 g62258(.A (n_9631), .Y (n_7732));
INVX2 g65659(.A (n_8653), .Y (n_4670));
OAI21X1 g65713(.A0 (n_2266), .A1 (n_3781), .B0 (n_3466), .Y (n_3960));
INVX1 g65760(.A (n_8644), .Y (n_3959));
NAND3X1 g65900(.A (n_9667), .B (n_9668), .C (n_2206), .Y (n_3955));
OAI21X1 g66052(.A0 (g1523), .A1 (n_3467), .B0 (n_2087), .Y (n_3774));
NAND3X1 g62418(.A (n_3128), .B (n_3402), .C (n_3300), .Y (n_3773));
NOR2X1 g66058(.A (n_941), .B (n_3455), .Y (n_3772));
OAI22X1 g66060(.A0 (g2226), .A1 (n_3768), .B0 (g2228), .B1 (n_3770),.Y (n_3771));
OAI21X1 g66061(.A0 (g2229), .A1 (n_3768), .B0 (n_2056), .Y (n_3769));
OAI21X1 g66062(.A0 (g2232), .A1 (n_3768), .B0 (n_2106), .Y (n_3767));
NAND3X1 g62429(.A (n_2963), .B (n_3401), .C (n_3296), .Y (n_3766));
NAND3X1 g62450(.A (n_3123), .B (n_3400), .C (n_3299), .Y (n_3765));
NAND2X1 g66253(.A (n_56), .B (n_6626), .Y (n_3763));
NOR2X1 g66265(.A (g1113), .B (n_3336), .Y (n_3762));
INVX1 g66330(.A (n_3953), .Y (n_3761));
OAI21X1 g62547(.A0 (n_3405), .A1 (n_3697), .B0 (n_3106), .Y (n_4218));
INVX1 g66365(.A (n_3568), .Y (n_3760));
INVX1 g66367(.A (n_3601), .Y (n_3759));
OR2X1 g66369(.A (g2395), .B (n_4576), .Y (n_9670));
INVX1 g66370(.A (n_3569), .Y (n_3756));
OR2X1 g66396(.A (g2477), .B (n_4576), .Y (n_3755));
OR2X1 g66466(.A (g_25960), .B (n_4172), .Y (n_3754));
NAND2X1 g66486(.A (g2685), .B (n_3448), .Y (n_3753));
NAND2X1 g66487(.A (n_3448), .B (g2694), .Y (n_3752));
INVX2 g66660(.A (g1782), .Y (n_5008));
CLKBUFX1 gbuf_d_827(.A(n_3555), .Y(d_out_827));
CLKBUFX1 gbuf_q_827(.A(q_in_827), .Y(g731));
CLKBUFX1 gbuf_d_828(.A(n_3558), .Y(d_out_828));
CLKBUFX1 gbuf_q_828(.A(q_in_828), .Y(g1319));
CLKBUFX1 gbuf_d_829(.A(n_3417), .Y(d_out_829));
CLKBUFX1 gbuf_q_829(.A(q_in_829), .Y(g633));
CLKBUFX1 gbuf_d_830(.A(gbuf201), .Y(d_out_830));
CLKBUFX1 gbuf_q_830(.A(q_in_830), .Y(g2598));
NOR2X1 g62967(.A (n_3523), .B (n_5181), .Y (n_3744));
NAND2X1 g63019(.A (n_3422), .B (n_3685), .Y (n_3743));
NOR2X1 g63053(.A (n_3518), .B (n_3407), .Y (n_3742));
NAND4X1 g63068(.A (n_3685), .B (n_3842), .C (n_2197), .D (n_3863), .Y(n_3741));
NOR2X1 g63072(.A (n_3517), .B (n_3406), .Y (n_3739));
NOR2X1 g63183(.A (n_3416), .B (n_3525), .Y (n_3738));
NAND4X1 g63187(.A (n_3648), .B (n_3736), .C (n_3705), .D (n_3735), .Y(n_3737));
NAND3X1 g63195(.A (n_1536), .B (n_1959), .C (n_3662), .Y (n_3734));
NOR2X1 g63202(.A (n_3514), .B (n_3374), .Y (n_3732));
NAND3X1 g63241(.A (n_3359), .B (n_3684), .C (n_1955), .Y (n_3731));
AOI21X1 g63242(.A0 (n_3249), .A1 (g646), .B0 (g660), .Y (n_3729));
NAND3X1 g63255(.A (n_3515), .B (n_3524), .C (n_2037), .Y (n_3728));
CLKBUFX1 gbuf_d_831(.A(n_3418), .Y(d_out_831));
CLKBUFX1 gbuf_q_831(.A(q_in_831), .Y(g2013));
NAND3X1 g63337(.A (n_3413), .B (n_1536), .C (n_3575), .Y (n_3726));
OR2X1 g66373(.A (g2389), .B (n_3546), .Y (n_3725));
CLKBUFX1 gbuf_d_832(.A(gbuf53), .Y(d_out_832));
CLKBUFX1 gbuf_q_832(.A(q_in_832), .Y(gbuf54));
CLKBUFX1 gbuf_d_833(.A(gbuf210), .Y(d_out_833));
CLKBUFX1 gbuf_q_833(.A(q_in_833), .Y(gbuf211));
CLKBUFX1 gbuf_d_834(.A(gbuf63), .Y(d_out_834));
CLKBUFX1 gbuf_q_834(.A(q_in_834), .Y(gbuf64));
NOR2X1 g63449(.A (n_3866), .B (n_2959), .Y (n_3900));
NOR2X1 g63450(.A (n_3724), .B (n_245), .Y (n_3902));
AND2X1 g63483(.A (n_3897), .B (g3229), .Y (n_3723));
AND2X1 g63487(.A (n_3721), .B (g3229), .Y (n_3722));
AND2X1 g63547(.A (n_4116), .B (n_3718), .Y (n_3720));
NAND2X1 g63559(.A (n_3716), .B (n_3893), .Y (n_3717));
AND2X1 g63571(.A (n_3897), .B (n_3714), .Y (n_3715));
NAND2X1 g63579(.A (n_3712), .B (n_4376), .Y (n_3713));
OR2X1 g66350(.A (g2396), .B (n_4576), .Y (n_3711));
NAND2X1 g63599(.A (n_3724), .B (n_3664), .Y (n_3710));
NAND3X1 g63682(.A (n_3531), .B (n_3361), .C (n_3864), .Y (n_3709));
AND2X1 g63702(.A (n_3864), .B (n_3893), .Y (n_3708));
AND2X1 g63703(.A (n_3515), .B (n_3705), .Y (n_3707));
AND2X1 g63706(.A (n_4027), .B (n_4081), .Y (n_3704));
NOR2X1 g63730(.A (n_3368), .B (n_5181), .Y (n_3703));
AOI21X1 g63767(.A0 (n_3372), .A1 (n_3701), .B0 (n_4151), .Y (n_3702));
OR2X1 g63781(.A (g869), .B (n_4162), .Y (n_4543));
AOI21X1 g63787(.A0 (n_7271), .A1 (n_3698), .B0 (n_3697), .Y (n_3700));
CLKBUFX1 gbuf_d_835(.A(n_3335), .Y(d_out_835));
CLKBUFX1 gbuf_q_835(.A(q_in_835), .Y(g2811));
INVX1 g63814(.A (n_3557), .Y (n_3696));
CLKBUFX1 gbuf_d_836(.A(n_3357), .Y(d_out_836));
CLKBUFX1 gbuf_q_836(.A(q_in_836), .Y(g737));
CLKBUFX1 gbuf_d_837(.A(n_3377), .Y(d_out_837));
CLKBUFX1 gbuf_q_837(.A(q_in_837), .Y(g1326));
MX2X1 g63938(.A (n_7271), .B (g1414), .S0 (n_3305), .Y (n_3695));
MX2X1 g63939(.A (n_7271), .B (g1415), .S0 (n_3303), .Y (n_3694));
MX2X1 g63940(.A (g1416), .B (n_7271), .S0 (n_4963), .Y (n_3693));
MX2X1 g63946(.A (n_4317), .B (g2111), .S0 (n_3691), .Y (n_3692));
MX2X1 g63947(.A (n_4317), .B (g2112), .S0 (n_3689), .Y (n_3690));
MX2X1 g63948(.A (g2113), .B (n_4317), .S0 (n_4967), .Y (n_3688));
NOR2X1 g64181(.A (n_3129), .B (n_3256), .Y (n_3687));
NOR2X1 g64206(.A (n_2783), .B (n_4037), .Y (n_3686));
NOR2X1 g64231(.A (n_3685), .B (n_3684), .Y (n_3891));
NOR2X1 g64244(.A (n_3648), .B (n_3524), .Y (n_4592));
NAND2X1 g64289(.A (n_8877), .B (n_465), .Y (n_3682));
NAND2X1 g64292(.A (n_9672), .B (n_468), .Y (n_3681));
NAND2X1 g64308(.A (n_3679), .B (n_3678), .Y (n_3680));
INVX1 g64332(.A (n_3677), .Y (n_3845));
NAND2X1 g64342(.A (n_3675), .B (n_3674), .Y (n_3676));
CLKBUFX1 gbuf_d_838(.A(n_3317), .Y(d_out_838));
CLKBUFX1 gbuf_q_838(.A(q_in_838), .Y(g846));
NOR2X1 g64397(.A (n_3651), .B (n_3363), .Y (n_4091));
NOR2X1 g64418(.A (n_3394), .B (g3229), .Y (n_3671));
NOR2X1 g64419(.A (n_3525), .B (n_3736), .Y (n_3669));
NAND2X1 g64420(.A (n_3489), .B (g801), .Y (n_3667));
NAND2X1 g64422(.A (n_3665), .B (n_3664), .Y (n_3666));
NAND2X1 g64427(.A (n_1359), .B (n_3662), .Y (n_3663));
NAND2X1 g64433(.A (n_8778), .B (g793), .Y (n_3661));
CLKBUFX1 gbuf_d_839(.A(n_3386), .Y(d_out_839));
CLKBUFX1 gbuf_q_839(.A(q_in_839), .Y(g_17170));
NAND3X1 g64465(.A (n_3508), .B (g2746), .C (g2740), .Y (n_4059));
CLKBUFX1 gbuf_d_840(.A(n_3316), .Y(d_out_840));
CLKBUFX1 gbuf_q_840(.A(q_in_840), .Y(g_23514));
XOR2X1 g64512(.A (g646), .B (n_3516), .Y (n_3660));
MX2X1 g64518(.A (n_3611), .B (n_6947), .S0 (n_5270), .Y (n_3659));
OR2X1 g64607(.A (n_4104), .B (g3229), .Y (n_3833));
NOR2X1 g64619(.A (n_3530), .B (n_3361), .Y (n_4127));
NAND2X1 g64659(.A (n_3530), .B (n_3684), .Y (n_3829));
NAND2X1 g64668(.A (n_3378), .B (n_3835), .Y (n_3658));
INVX1 g64699(.A (n_3656), .Y (n_3657));
NOR2X1 g64719(.A (n_3367), .B (n_2759), .Y (n_3655));
AOI21X1 g64870(.A0 (n_2594), .A1 (n_3816), .B0 (n_3338), .Y (n_3650));
INVX1 g64874(.A (n_9043), .Y (n_3825));
AOI21X1 g64888(.A0 (n_2603), .A1 (n_3816), .B0 (n_3339), .Y (n_3823));
INVX1 g64895(.A (n_3685), .Y (n_3822));
AOI21X1 g64914(.A0 (n_2595), .A1 (n_3816), .B0 (n_3350), .Y (n_3820));
CLKBUFX1 gbuf_d_841(.A(n_3322), .Y(d_out_841));
CLKBUFX1 gbuf_q_841(.A(q_in_841), .Y(g839));
INVX1 g64977(.A (n_3648), .Y (n_4053));
OAI21X1 g64986(.A0 (g1008), .A1 (n_3336), .B0 (n_2501), .Y (n_6726));
AOI21X1 g65004(.A0 (n_2598), .A1 (n_3816), .B0 (n_3349), .Y (n_3814));
NAND2X1 g65033(.A (n_3345), .B (n_2502), .Y (n_4312));
INVX1 g65044(.A (n_9449), .Y (n_3812));
AOI22X1 g65089(.A0 (n_2486), .A1 (n_3264), .B0 (g1877), .B1 (n_6626),.Y (n_3646));
INVX1 g65092(.A (n_3499), .Y (n_4056));
INVX1 g65156(.A (n_3642), .Y (n_3805));
AOI21X1 g65252(.A0 (n_2306), .A1 (n_3799), .B0 (n_3370), .Y (n_3800));
INVX1 g65322(.A (n_3638), .Y (n_4339));
INVX1 g65344(.A (n_3636), .Y (n_3795));
CLKBUFX1 gbuf_d_842(.A(n_3391), .Y(d_out_842));
CLKBUFX1 gbuf_q_842(.A(q_in_842), .Y(g_14013));
NAND4X1 g62229(.A (n_3124), .B (n_2954), .C (n_3125), .D (n_3126), .Y(n_3635));
NAND4X1 g62232(.A (n_3119), .B (n_3216), .C (n_3118), .D (n_3122), .Y(n_3634));
AOI22X1 g65586(.A0 (n_3153), .A1 (n_313), .B0 (g1165), .B1 (n_1660),.Y (n_3633));
AOI22X1 g65593(.A0 (n_3221), .A1 (g1173), .B0 (g1174), .B1 (n_1660),.Y (n_3632));
CLKBUFX1 g65596(.A (n_3630), .Y (n_4014));
AOI22X1 g65604(.A0 (n_3222), .A1 (g1167), .B0 (g1171), .B1 (n_1660),.Y (n_3629));
NAND4X1 g62256(.A (n_2994), .B (n_3155), .C (n_3110), .D (n_2958), .Y(n_4044));
INVX1 g65608(.A (n_4015), .Y (n_3790));
INVX1 g65644(.A (n_3848), .Y (n_3625));
INVX1 g65698(.A (n_3620), .Y (n_3804));
OAI21X1 g65708(.A0 (g1089), .A1 (n_3336), .B0 (n_2395), .Y (n_6546));
INVX1 g65897(.A (n_3479), .Y (n_3616));
INVX1 g65903(.A (n_3478), .Y (n_3615));
INVX1 g65905(.A (n_3477), .Y (n_3614));
OAI22X1 g66059(.A0 (g2238), .A1 (n_3224), .B0 (g2240), .B1 (n_3770),.Y (n_3613));
CLKBUFX1 gbuf_d_843(.A(n_3320), .Y(d_out_843));
CLKBUFX1 gbuf_q_843(.A(q_in_843), .Y(g840));
OAI21X1 g66107(.A0 (n_3611), .A1 (n_3220), .B0 (n_3342), .Y (n_3612));
OR2X1 g66215(.A (g2244), .B (n_3344), .Y (n_3610));
NOR2X1 g62503(.A (n_3138), .B (n_3314), .Y (n_3609));
NOR2X1 g62505(.A (n_3137), .B (n_3312), .Y (n_3608));
OR2X1 g66296(.A (g1868), .B (g1930), .Y (n_3607));
INVX1 g66306(.A (n_3463), .Y (n_3606));
OR2X1 g66313(.A (g2217), .B (n_3768), .Y (n_3605));
NOR2X1 g66331(.A (n_3873), .B (n_4162), .Y (n_3953));
OR2X1 g66358(.A (g1532), .B (n_3467), .Y (n_3603));
INVX1 g66361(.A (n_3424), .Y (n_3602));
NOR2X1 g66368(.A (g1535), .B (n_3467), .Y (n_3601));
INVX1 g66378(.A (n_3426), .Y (n_3597));
NOR2X1 g66381(.A (g865), .B (n_4162), .Y (n_3596));
OR2X1 g66429(.A (g1865), .B (g1930), .Y (n_3595));
INVX1 g66470(.A (n_3441), .Y (n_8242));
INVX1 g66482(.A (n_3440), .Y (n_3592));
NAND2X1 g66605(.A (g1930), .B (n_1689), .Y (n_4880));
CLKBUFX1 gbuf_d_844(.A(g7014), .Y(d_out_844));
CLKBUFX1 gbuf_q_844(.A(q_in_844), .Y(g1782));
INVX1 g66765(.A (n_3588), .Y (n_7809));
INVX2 g66797(.A (g401), .Y (n_5004));
INVX4 g66852(.A (n_4125), .Y (n_7800));
CLKBUFX1 gbuf_d_845(.A(n_3351), .Y(d_out_845));
CLKBUFX1 gbuf_q_845(.A(q_in_845), .Y(g2733));
NOR2X1 g62946(.A (n_3389), .B (n_4967), .Y (n_3581));
NAND3X1 g62966(.A (n_4078), .B (n_3534), .C (n_2985), .Y (n_3580));
NOR2X1 g62968(.A (n_3392), .B (n_4963), .Y (n_3579));
CLKBUFX1 gbuf_d_846(.A(n_3319), .Y(d_out_846));
CLKBUFX1 gbuf_q_846(.A(q_in_846), .Y(g845));
NAND3X1 g63192(.A (n_3239), .B (n_3534), .C (n_3427), .Y (n_3578));
NAND3X1 g63193(.A (n_1536), .B (n_3576), .C (n_3575), .Y (n_3577));
NAND2X1 g63194(.A (n_3409), .B (n_3325), .Y (n_3574));
CLKBUFX1 gbuf_d_847(.A(n_3404), .Y(d_out_847));
CLKBUFX1 gbuf_q_847(.A(q_in_847), .Y(g659));
NAND3X1 g63257(.A (n_4078), .B (n_3533), .C (n_3410), .Y (n_3573));
AOI21X1 g63259(.A0 (n_3364), .A1 (g2720), .B0 (g2734), .Y (n_3572));
CLKBUFX1 gbuf_d_848(.A(n_3379), .Y(d_out_848));
CLKBUFX1 gbuf_q_848(.A(q_in_848), .Y(g2020));
NAND3X1 g63819(.A (n_3239), .B (n_2929), .C (n_1264), .Y (n_3571));
NOR2X1 g66371(.A (g1538), .B (n_3467), .Y (n_3569));
NOR2X1 g66366(.A (g1526), .B (n_3467), .Y (n_3568));
CLKBUFX1 gbuf_d_849(.A(n_3388), .Y(d_out_849));
CLKBUFX1 gbuf_q_849(.A(q_in_849), .Y(g_26381));
CLKBUFX1 gbuf_d_850(.A(gbuf102), .Y(d_out_850));
CLKBUFX1 gbuf_q_850(.A(q_in_850), .Y(gbuf103));
CLKBUFX1 gbuf_d_851(.A(gbuf112), .Y(d_out_851));
CLKBUFX1 gbuf_q_851(.A(q_in_851), .Y(gbuf113));
CLKBUFX1 gbuf_d_852(.A(n_3324), .Y(d_out_852));
CLKBUFX1 gbuf_q_852(.A(q_in_852), .Y(g_30039));
OR2X1 g66357(.A (g1544), .B (n_3467), .Y (n_3567));
CLKBUFX1 gbuf_d_853(.A(n_3385), .Y(d_out_853));
CLKBUFX1 gbuf_q_853(.A(q_in_853), .Y(g_30213));
NOR2X1 g63680(.A (n_3530), .B (n_3421), .Y (n_3565));
NAND2X1 g63715(.A (n_3562), .B (n_4362), .Y (n_3563));
NAND2X1 g63724(.A (n_3560), .B (n_3559), .Y (n_3561));
NOR2X1 g63729(.A (n_3253), .B (n_4963), .Y (n_3558));
CLKBUFX1 gbuf_d_854(.A(n_3178), .Y(d_out_854));
CLKBUFX1 gbuf_q_854(.A(q_in_854), .Y(g_19132));
CLKBUFX1 gbuf_d_855(.A(n_3205), .Y(d_out_855));
CLKBUFX1 gbuf_q_855(.A(q_in_855), .Y(g716));
AOI21X1 g63815(.A0 (n_3256), .A1 (g2584), .B0 (n_4151), .Y (n_3557));
CLKBUFX1 gbuf_d_856(.A(n_3207), .Y(d_out_856));
CLKBUFX1 gbuf_q_856(.A(q_in_856), .Y(g707));
CLKBUFX1 gbuf_d_857(.A(n_3308), .Y(d_out_857));
CLKBUFX1 gbuf_q_857(.A(q_in_857), .Y(g713));
CLKBUFX1 gbuf_d_858(.A(n_3168), .Y(d_out_858));
CLKBUFX1 gbuf_q_858(.A(q_in_858), .Y(g836));
AOI22X1 g63898(.A0 (n_2941), .A1 (n_3203), .B0 (n_4695), .B1 (n_163),.Y (n_3556));
CLKBUFX1 gbuf_d_859(.A(n_3152), .Y(d_out_859));
CLKBUFX1 gbuf_q_859(.A(q_in_859), .Y(g2772));
CLKBUFX1 gbuf_d_860(.A(n_3149), .Y(d_out_860));
CLKBUFX1 gbuf_q_860(.A(q_in_860), .Y(g2778));
CLKBUFX1 gbuf_d_861(.A(n_3148), .Y(d_out_861));
CLKBUFX1 gbuf_q_861(.A(q_in_861), .Y(g2781));
CLKBUFX1 gbuf_d_862(.A(n_3142), .Y(d_out_862));
CLKBUFX1 gbuf_q_862(.A(q_in_862), .Y(g2796));
CLKBUFX1 gbuf_d_863(.A(n_3302), .Y(d_out_863));
CLKBUFX1 gbuf_q_863(.A(q_in_863), .Y(g1419));
CLKBUFX1 gbuf_d_864(.A(n_3212), .Y(d_out_864));
CLKBUFX1 gbuf_q_864(.A(q_in_864), .Y(g701));
MX2X1 g63952(.A (n_5101), .B (g731), .S0 (n_3554), .Y (n_3555));
MX2X1 g63953(.A (n_5101), .B (g732), .S0 (n_3552), .Y (n_3553));
MX2X1 g63955(.A (g733), .B (n_5101), .S0 (n_5372), .Y (n_3551));
CLKBUFX1 gbuf_d_865(.A(n_3180), .Y(d_out_865));
CLKBUFX1 gbuf_q_865(.A(q_in_865), .Y(g_24593));
XOR2X1 g64052(.A (g640), .B (n_2940), .Y (n_3550));
CLKBUFX1 gbuf_d_866(.A(n_3213), .Y(d_out_866));
CLKBUFX1 gbuf_q_866(.A(q_in_866), .Y(g698));
CLKBUFX1 gbuf_d_867(.A(n_3549), .Y(d_out_867));
CLKBUFX1 gbuf_q_867(.A(q_in_867), .Y(gbuf63));
CLKBUFX1 gbuf_d_868(.A(n_3548), .Y(d_out_868));
CLKBUFX1 gbuf_q_868(.A(q_in_868), .Y(gbuf210));
CLKBUFX1 gbuf_d_869(.A(n_3547), .Y(d_out_869));
CLKBUFX1 gbuf_q_869(.A(q_in_869), .Y(gbuf53));
INVX1 g66878(.A (g2476), .Y (n_3546));
AND2X1 g64197(.A (n_3544), .B (n_4317), .Y (n_3545));
AND2X1 g64198(.A (n_3542), .B (n_4317), .Y (n_3543));
AND2X1 g64199(.A (n_3540), .B (n_4317), .Y (n_3541));
AND2X1 g64201(.A (n_2626), .B (n_4317), .Y (n_3539));
NOR2X1 g64219(.A (n_2637), .B (n_2927), .Y (n_3537));
OR2X1 g64221(.A (n_3534), .B (g3229), .Y (n_3536));
NOR2X1 g64225(.A (n_3525), .B (n_3515), .Y (n_4081));
NOR2X1 g64232(.A (n_3531), .B (n_3359), .Y (n_3893));
NOR2X1 g64249(.A (n_3533), .B (n_3534), .Y (n_3908));
CLKBUFX1 gbuf_d_870(.A(n_3150), .Y(d_out_870));
CLKBUFX1 gbuf_q_870(.A(q_in_870), .Y(g2775));
INVX2 g66854(.A (n_3467), .Y (n_4125));
NOR2X1 g64273(.A (n_3533), .B (n_2929), .Y (n_3878));
CLKBUFX1 gbuf_d_871(.A(n_3157), .Y(d_out_871));
CLKBUFX1 gbuf_q_871(.A(q_in_871), .Y(g_20947));
NOR2X1 g64297(.A (n_4096), .B (n_4116), .Y (n_3897));
CLKBUFX1 gbuf_d_872(.A(n_3274), .Y(d_out_872));
CLKBUFX1 gbuf_q_872(.A(q_in_872), .Y(g704));
NAND2X1 g64333(.A (n_3531), .B (n_3530), .Y (n_3677));
NAND2X1 g64369(.A (n_4151), .B (n_4317), .Y (n_3529));
INVX1 g64386(.A (n_3527), .Y (n_3721));
NOR2X1 g64409(.A (n_3525), .B (n_3524), .Y (n_3884));
NAND3X1 g64447(.A (n_3381), .B (g2046), .C (g2052), .Y (n_3724));
NAND3X1 g64463(.A (n_3380), .B (g1358), .C (g1352), .Y (n_3866));
XOR2X1 g64513(.A (g2720), .B (n_3378), .Y (n_3523));
CLKBUFX1 gbuf_d_873(.A(n_3188), .Y(d_out_873));
CLKBUFX1 gbuf_q_873(.A(q_in_873), .Y(g_16484));
CLKBUFX1 gbuf_d_874(.A(n_3141), .Y(d_out_874));
CLKBUFX1 gbuf_q_874(.A(q_in_874), .Y(g2799));
NAND2X1 g64603(.A (n_4102), .B (g3229), .Y (n_3521));
NOR2X1 g64604(.A (n_4102), .B (g3229), .Y (n_4523));
AND2X1 g64618(.A (n_4116), .B (n_3363), .Y (n_4376));
NAND2X1 g64666(.A (n_3270), .B (n_3664), .Y (n_3518));
NAND2X1 g64684(.A (n_3516), .B (n_3674), .Y (n_3517));
CLKBUFX1 gbuf_d_875(.A(n_3162), .Y(d_out_875));
CLKBUFX1 gbuf_q_875(.A(q_in_875), .Y(g_19162));
NOR2X1 g64700(.A (n_3515), .B (n_3415), .Y (n_3656));
NAND2X1 g64704(.A (n_3269), .B (n_3678), .Y (n_3514));
NOR2X1 g64708(.A (n_3252), .B (n_2756), .Y (n_3513));
INVX1 g66767(.A (n_3344), .Y (n_3588));
INVX1 g64726(.A (n_3675), .Y (n_3509));
INVX1 g64735(.A (n_3508), .Y (n_3836));
CLKBUFX1 gbuf_d_876(.A(n_3147), .Y(d_out_876));
CLKBUFX1 gbuf_q_876(.A(q_in_876), .Y(g2784));
CLKBUFX1 gbuf_d_877(.A(n_3144), .Y(d_out_877));
CLKBUFX1 gbuf_q_877(.A(q_in_877), .Y(g2793));
INVX1 g64978(.A (n_3525), .Y (n_3648));
AOI22X1 g65093(.A0 (n_2403), .A1 (n_3498), .B0 (g_25958), .B1(n_4601), .Y (n_3499));
CLKBUFX1 gbuf_d_878(.A(n_3165), .Y(d_out_878));
CLKBUFX1 gbuf_q_878(.A(q_in_878), .Y(g842));
INVX1 g65149(.A (n_8411), .Y (n_3643));
INVX1 g65157(.A (n_9671), .Y (n_3642));
AOI22X1 g65163(.A0 (n_2169), .A1 (n_3264), .B0 (g1953), .B1 (n_6626),.Y (n_3856));
AOI22X1 g65182(.A0 (n_2506), .A1 (n_3264), .B0 (g1870), .B1 (n_6626),.Y (n_3855));
INVX2 g65189(.A (n_4037), .Y (n_5323));
INVX1 g65323(.A (n_3489), .Y (n_3638));
AOI22X1 g65345(.A0 (n_2174), .A1 (n_2925), .B0 (g2571), .B1 (n_2863),.Y (n_3636));
CLKBUFX1 gbuf_d_879(.A(n_3163), .Y(d_out_879));
CLKBUFX1 gbuf_q_879(.A(q_in_879), .Y(g843));
NAND3X1 g65597(.A (n_9698), .B (n_9699), .C (n_3053), .Y (n_3630));
NAND3X1 g65609(.A (n_1140), .B (n_2246), .C (n_2988), .Y (n_4015));
INVX1 g65628(.A (n_3363), .Y (n_3628));
AOI21X1 g65645(.A0 (n_2008), .A1 (n_3264), .B0 (n_3218), .Y (n_3848));
OAI21X1 g65699(.A0 (n_2269), .A1 (n_3482), .B0 (n_3217), .Y (n_3620));
NAND3X1 g65896(.A (n_3140), .B (n_1015), .C (n_2069), .Y (n_3480));
NAND3X1 g65898(.A (n_8365), .B (n_1105), .C (n_8366), .Y (n_3479));
NAND3X1 g65904(.A (n_3227), .B (n_1127), .C (n_2254), .Y (n_3478));
NAND3X1 g65906(.A (n_8367), .B (n_1083), .C (n_8368), .Y (n_3477));
CLKBUFX1 gbuf_d_880(.A(n_3229), .Y(d_out_880));
CLKBUFX1 gbuf_q_880(.A(q_in_880), .Y(g2704));
CLKBUFX1 gbuf_d_881(.A(n_3231), .Y(d_out_881));
CLKBUFX1 gbuf_q_881(.A(q_in_881), .Y(g630));
AOI21X1 g63824(.A0 (n_2905), .A1 (g2707), .B0 (g2727), .Y (n_3476));
MX2X1 g66120(.A (g1243), .B (n_3698), .S0 (n_3220), .Y (n_3475));
NOR2X1 g63823(.A (n_5531), .B (n_3036), .Y (n_3474));
NOR2X1 g66212(.A (n_112), .B (n_3224), .Y (n_3473));
OR2X1 g66217(.A (n_334), .B (n_3467), .Y (n_3472));
NOR2X1 g66218(.A (n_207), .B (n_3467), .Y (n_3471));
OR2X1 g66285(.A (n_143), .B (n_3467), .Y (n_3468));
OR2X1 g66288(.A (g1556), .B (n_3467), .Y (n_3466));
OR2X1 g66294(.A (g2562), .B (n_3448), .Y (n_3465));
NOR2X1 g66304(.A (n_4), .B (n_3467), .Y (n_3464));
NOR2X1 g66307(.A (g2205), .B (n_3224), .Y (n_3463));
OR2X1 g66308(.A (n_44), .B (n_3467), .Y (n_3461));
OR2X1 g66328(.A (n_125), .B (n_3467), .Y (n_3460));
OR2X1 g66332(.A (g487), .B (n_2748), .Y (n_3459));
OR2X1 g66337(.A (n_209), .B (n_3467), .Y (n_3458));
NOR2X1 g66346(.A (n_54), .B (n_3467), .Y (n_3457));
OR2X1 g66377(.A (g2220), .B (n_3224), .Y (n_9668));
NOR2X1 g66380(.A (g2223), .B (n_3224), .Y (n_3455));
OR2X1 g66383(.A (n_75), .B (n_3224), .Y (n_3454));
NOR2X1 g66386(.A (n_113), .B (n_3224), .Y (n_3452));
OR2X1 g66390(.A (n_38), .B (n_3467), .Y (n_3451));
NOR2X1 g66399(.A (g838), .B (n_4162), .Y (n_3450));
OR2X1 g66413(.A (g2553), .B (n_3448), .Y (n_3449));
NOR2X1 g66418(.A (g856), .B (n_4162), .Y (n_3447));
OR2X1 g66430(.A (g484), .B (n_2748), .Y (n_3445));
OR2X1 g66437(.A (n_239), .B (n_3224), .Y (n_3443));
OR2X1 g66452(.A (g478), .B (n_2748), .Y (n_3442));
NOR2X1 g66471(.A (g1514), .B (n_3467), .Y (n_3441));
NOR2X1 g66483(.A (g1529), .B (n_3467), .Y (n_3440));
NOR2X1 g66492(.A (n_76), .B (n_3467), .Y (n_3439));
OR2X1 g66494(.A (g2559), .B (n_3448), .Y (n_3438));
NAND2X1 g66567(.A (n_2748), .B (n_1911), .Y (n_4660));
NAND2X1 g66598(.A (n_3448), .B (n_1596), .Y (n_4655));
CLKBUFX1 gbuf_d_882(.A(g6447), .Y(d_out_882));
CLKBUFX1 gbuf_q_882(.A(q_in_882), .Y(g401));
INVX4 g66877(.A (g2476), .Y (n_4576));
NAND2X1 g66943(.A (g1813), .B (n_3036), .Y (n_3433));
NAND2X1 g66960(.A (g1697), .B (n_3036), .Y (n_3431));
CLKBUFX1 gbuf_d_883(.A(n_3173), .Y(d_out_883));
CLKBUFX1 gbuf_q_883(.A(q_in_883), .Y(g822));
CLKBUFX1 gbuf_d_884(.A(n_3160), .Y(d_out_884));
CLKBUFX1 gbuf_q_884(.A(q_in_884), .Y(g834));
CLKBUFX1 gbuf_d_885(.A(n_3170), .Y(d_out_885));
CLKBUFX1 gbuf_q_885(.A(q_in_885), .Y(g833));
CLKBUFX1 gbuf_d_886(.A(n_3145), .Y(d_out_886));
CLKBUFX1 gbuf_q_886(.A(q_in_886), .Y(g2790));
CLKBUFX1 gbuf_d_887(.A(n_3172), .Y(d_out_887));
CLKBUFX1 gbuf_q_887(.A(q_in_887), .Y(g831));
CLKBUFX1 gbuf_d_888(.A(n_3202), .Y(d_out_888));
CLKBUFX1 gbuf_q_888(.A(q_in_888), .Y(g722));
CLKBUFX1 gbuf_d_889(.A(n_3159), .Y(d_out_889));
CLKBUFX1 gbuf_q_889(.A(q_in_889), .Y(g830));
NAND3X1 g63184(.A (n_3393), .B (n_3430), .C (g3229), .Y (n_4826));
CLKBUFX1 gbuf_d_890(.A(n_3158), .Y(d_out_890));
CLKBUFX1 gbuf_q_890(.A(q_in_890), .Y(g_14855));
CLKBUFX1 gbuf_d_891(.A(n_3146), .Y(d_out_891));
CLKBUFX1 gbuf_q_891(.A(q_in_891), .Y(g2787));
AOI21X1 g63233(.A0 (n_3247), .A1 (g2026), .B0 (g2040), .Y (n_3429));
CLKBUFX1 gbuf_d_892(.A(n_3166), .Y(d_out_892));
CLKBUFX1 gbuf_q_892(.A(q_in_892), .Y(g837));
NAND3X1 g63256(.A (n_4078), .B (n_3394), .C (n_3427), .Y (n_3428));
NOR2X1 g66379(.A (g2208), .B (n_3224), .Y (n_3426));
AOI21X1 g63260(.A0 (n_3245), .A1 (g1332), .B0 (g1346), .Y (n_3425));
CLKBUFX1 gbuf_d_893(.A(n_3306), .Y(d_out_893));
CLKBUFX1 gbuf_q_893(.A(q_in_893), .Y(g1417));
CLKBUFX1 gbuf_d_894(.A(n_3174), .Y(d_out_894));
CLKBUFX1 gbuf_q_894(.A(q_in_894), .Y(g821));
CLKBUFX1 gbuf_d_895(.A(n_3175), .Y(d_out_895));
CLKBUFX1 gbuf_q_895(.A(q_in_895), .Y(g819));
CLKBUFX1 gbuf_d_896(.A(n_3204), .Y(d_out_896));
CLKBUFX1 gbuf_q_896(.A(q_in_896), .Y(g719));
NOR2X1 g66362(.A (g1511), .B (n_3467), .Y (n_3424));
CLKBUFX1 gbuf_d_897(.A(gbuf200), .Y(d_out_897));
CLKBUFX1 gbuf_q_897(.A(q_in_897), .Y(gbuf201));
CLKBUFX1 gbuf_d_898(.A(n_3304), .Y(d_out_898));
CLKBUFX1 gbuf_q_898(.A(q_in_898), .Y(g1418));
CLKBUFX1 gbuf_d_899(.A(n_3206), .Y(d_out_899));
CLKBUFX1 gbuf_q_899(.A(q_in_899), .Y(g710));
AND2X1 g63490(.A (n_3576), .B (g3229), .Y (n_3423));
CLKBUFX1 gbuf_d_900(.A(n_3201), .Y(d_out_900));
CLKBUFX1 gbuf_q_900(.A(q_in_900), .Y(g725));
NOR2X1 g63556(.A (n_3684), .B (n_3421), .Y (n_3422));
OR2X1 g63557(.A (n_3842), .B (n_3419), .Y (n_3420));
NOR2X1 g63583(.A (n_3255), .B (n_4967), .Y (n_3418));
NOR2X1 g63600(.A (n_3254), .B (n_5372), .Y (n_3417));
CLKBUFX1 gbuf_d_901(.A(n_3176), .Y(d_out_901));
CLKBUFX1 gbuf_q_901(.A(q_in_901), .Y(g818));
NAND2X1 g63712(.A (n_3415), .B (n_3705), .Y (n_3416));
NAND2X1 g63718(.A (n_3559), .B (n_3408), .Y (n_3414));
NOR2X1 g63720(.A (n_3412), .B (n_4078), .Y (n_3413));
AND2X1 g63722(.A (n_3576), .B (n_3410), .Y (n_3411));
NAND2X1 g63726(.A (n_3408), .B (n_3430), .Y (n_3409));
AOI21X1 g63788(.A0 (n_2760), .A1 (g2013), .B0 (g2033), .Y (n_3407));
AOI21X1 g63790(.A0 (n_3070), .A1 (g633), .B0 (g653), .Y (n_3406));
AOI21X1 g63794(.A0 (n_2927), .A1 (n_3698), .B0 (n_4151), .Y (n_3405));
CLKBUFX1 gbuf_d_902(.A(n_3022), .Y(d_out_902));
CLKBUFX1 gbuf_q_902(.A(q_in_902), .Y(g2117));
CLKBUFX1 gbuf_d_903(.A(n_3058), .Y(d_out_903));
CLKBUFX1 gbuf_q_903(.A(q_in_903), .Y(g2039));
OAI21X1 g66104(.A0 (n_4151), .A1 (n_2814), .B0 (n_2989), .Y (n_3404));
XOR2X1 g64008(.A (g2746), .B (n_2805), .Y (n_3403));
XOR2X1 g64012(.A (g2707), .B (n_2779), .Y (n_3402));
XOR2X1 g64029(.A (g1346), .B (n_2788), .Y (n_3401));
CLKBUFX1 gbuf_d_904(.A(n_3023), .Y(d_out_904));
CLKBUFX1 gbuf_q_904(.A(q_in_904), .Y(g1540));
XOR2X1 g64075(.A (g2040), .B (n_2783), .Y (n_3400));
XOR2X1 g64080(.A (n_3143), .B (n_2785), .Y (n_3399));
CLKBUFX1 gbuf_d_905(.A(n_3089), .Y(d_out_905));
CLKBUFX1 gbuf_q_905(.A(q_in_905), .Y(g1534));
CLKBUFX1 gbuf_d_906(.A(n_3398), .Y(d_out_906));
CLKBUFX1 gbuf_q_906(.A(q_in_906), .Y(gbuf102));
CLKBUFX1 gbuf_d_907(.A(n_3397), .Y(d_out_907));
CLKBUFX1 gbuf_q_907(.A(q_in_907), .Y(gbuf112));
NAND2X1 g64286(.A (n_4151), .B (n_5101), .Y (n_3396));
CLKBUFX1 gbuf_d_908(.A(n_3094), .Y(d_out_908));
CLKBUFX1 gbuf_q_908(.A(q_in_908), .Y(g1537));
CLKBUFX1 gbuf_d_909(.A(n_3096), .Y(d_out_909));
CLKBUFX1 gbuf_q_909(.A(q_in_909), .Y(g1536));
CLKBUFX1 gbuf_d_910(.A(n_3034), .Y(d_out_910));
CLKBUFX1 gbuf_q_910(.A(q_in_910), .Y(g1512));
NAND2X1 g64388(.A (n_3525), .B (n_3382), .Y (n_3527));
CLKBUFX1 gbuf_d_911(.A(n_3078), .Y(d_out_911));
CLKBUFX1 gbuf_q_911(.A(q_in_911), .Y(g1531));
NOR2X1 g64430(.A (n_3394), .B (n_3393), .Y (n_3395));
XOR2X1 g64476(.A (g1332), .B (n_3269), .Y (n_3392));
CLKBUFX1 gbuf_d_912(.A(n_3029), .Y(d_out_912));
CLKBUFX1 gbuf_q_912(.A(q_in_912), .Y(g1533));
CLKBUFX1 gbuf_d_913(.A(n_3027), .Y(d_out_913));
CLKBUFX1 gbuf_q_913(.A(q_in_913), .Y(g1539));
MX2X1 g64509(.A (g_14013), .B (n_3390), .S0 (n_3387), .Y (n_3391));
CLKBUFX1 gbuf_d_914(.A(n_3032), .Y(d_out_914));
CLKBUFX1 gbuf_q_914(.A(q_in_914), .Y(g1513));
XOR2X1 g64514(.A (g2026), .B (n_3270), .Y (n_3389));
MX2X1 g64531(.A (g_26381), .B (n_5663), .S0 (n_3387), .Y (n_3388));
MX2X1 g64533(.A (g_17170), .B (n_5382), .S0 (n_3387), .Y (n_3386));
MX2X1 g64550(.A (g_30213), .B (n_5380), .S0 (n_3387), .Y (n_3385));
NOR2X1 g64611(.A (n_2986), .B (g3229), .Y (n_4077));
NAND2X1 g64612(.A (n_2986), .B (g3229), .Y (n_3384));
NOR2X1 g64620(.A (n_3382), .B (n_3075), .Y (n_4362));
NOR2X1 g64643(.A (n_4078), .B (n_3239), .Y (n_3662));
INVX1 g64710(.A (n_3381), .Y (n_3665));
INVX1 g64713(.A (n_3380), .Y (n_3679));
NOR2X1 g64718(.A (n_3083), .B (n_2612), .Y (n_3379));
CLKBUFX1 gbuf_d_915(.A(n_3031), .Y(d_out_915));
CLKBUFX1 gbuf_q_915(.A(q_in_915), .Y(g1530));
NAND3X1 g64727(.A (n_3249), .B (g646), .C (g660), .Y (n_3675));
NOR2X1 g64736(.A (n_234), .B (n_3378), .Y (n_3508));
NOR2X1 g64737(.A (n_3081), .B (n_2607), .Y (n_3377));
INVX1 g64868(.A (n_4096), .Y (n_3651));
INVX1 g64899(.A (n_3531), .Y (n_3685));
AOI21X1 g63826(.A0 (n_2757), .A1 (g1319), .B0 (g1339), .Y (n_3374));
INVX1 g65180(.A (n_3263), .Y (n_3697));
OAI21X1 g65190(.A0 (n_2176), .A1 (n_1691), .B0 (n_3045), .Y (n_4037));
NOR2X1 g66484(.A (n_48), .B (n_3344), .Y (n_3370));
AOI21X1 g65324(.A0 (n_2390), .A1 (n_8408), .B0 (n_3039), .Y (n_3489));
XOR2X1 g65370(.A (g2707), .B (n_3251), .Y (n_3368));
NAND2X1 g65461(.A (n_3079), .B (n_3674), .Y (n_3367));
INVX1 g65636(.A (n_4116), .Y (n_3485));
INVX1 g65666(.A (n_3684), .Y (n_3361));
OAI21X1 g62290(.A0 (n_3064), .A1 (g630), .B0 (n_3065), .Y (n_3357));
NAND2X1 g65878(.A (n_3037), .B (n_5035), .Y (n_3356));
NAND2X1 g65888(.A (n_2732), .B (n_5035), .Y (n_3355));
NAND2X1 g65958(.A (n_3038), .B (n_5044), .Y (n_3354));
AOI22X1 g66080(.A0 (n_2862), .A1 (g1829), .B0 (g1830), .B1 (n_1235),.Y (n_3353));
AOI22X1 g66092(.A0 (n_2861), .A1 (g448), .B0 (g449), .B1 (n_1237), .Y(n_3352));
OAI21X1 g66106(.A0 (n_4151), .A1 (n_2674), .B0 (n_3047), .Y (n_3351));
NOR2X1 g66242(.A (g841), .B (n_4162), .Y (n_3350));
NOR2X1 g66277(.A (g850), .B (n_4162), .Y (n_3349));
NAND2X1 g66290(.A (g602), .B (n_4601), .Y (n_3347));
NAND2X1 g66317(.A (g1306), .B (n_3220), .Y (n_3346));
OR2X1 g66388(.A (n_176), .B (n_3344), .Y (n_3345));
NOR2X1 g66392(.A (n_51), .B (n_3344), .Y (n_3343));
NAND2X1 g66398(.A (n_3220), .B (g1243), .Y (n_3342));
OR2X1 g66402(.A (g1001), .B (n_3336), .Y (n_3340));
NOR2X1 g66409(.A (g844), .B (n_4162), .Y (n_3339));
NOR2X1 g66420(.A (g829), .B (n_4162), .Y (n_3338));
NOR2X1 g66439(.A (g1007), .B (n_3336), .Y (n_3337));
OAI21X1 g62568(.A0 (n_3010), .A1 (g2704), .B0 (n_3011), .Y (n_3335));
NAND2X1 g66479(.A (g2676), .B (n_2863), .Y (n_3334));
NOR2X1 g66493(.A (g2247), .B (n_3344), .Y (n_3333));
OR2X1 g66497(.A (g847), .B (n_4162), .Y (n_3332));
OR2X1 g66424(.A (g1004), .B (n_3336), .Y (n_3331));
CLKBUFX1 gbuf_d_916(.A(g6313), .Y(d_out_916));
CLKBUFX1 gbuf_q_916(.A(q_in_916), .Y(g_5550));
CLKBUFX1 g66754(.A (n_3224), .Y (n_3768));
CLKBUFX1 gbuf_d_917(.A(g7264), .Y(d_out_917));
CLKBUFX1 gbuf_q_917(.A(q_in_917), .Y(g2476));
INVX1 g66932(.A (n_3336), .Y (n_3808));
NAND2X1 g67147(.A (g_10841), .B (n_2874), .Y (n_9691));
CLKBUFX1 gbuf_d_918(.A(n_3074), .Y(d_out_918));
CLKBUFX1 gbuf_q_918(.A(q_in_918), .Y(g1423));
NAND4X1 g63914(.A (n_3394), .B (n_3393), .C (n_1264), .D (n_1518), .Y(n_3325));
OAI21X1 g62764(.A0 (n_5585), .A1 (n_733), .B0 (n_3003), .Y (n_3324));
OAI21X1 g62780(.A0 (n_4540), .A1 (g805), .B0 (n_3009), .Y (n_3322));
OAI21X1 g62781(.A0 (n_4538), .A1 (g805), .B0 (n_3002), .Y (n_3320));
OAI21X1 g62786(.A0 (n_4540), .A1 (n_763), .B0 (n_3008), .Y (n_3319));
OAI21X1 g62787(.A0 (n_4538), .A1 (n_763), .B0 (n_3007), .Y (n_3317));
OAI21X1 g62794(.A0 (n_5585), .A1 (g125), .B0 (n_3001), .Y (n_3316));
NAND4X1 g63209(.A (n_3313), .B (n_9569), .C (n_2646), .D (n_4685), .Y(n_3314));
NAND4X1 g63215(.A (n_2996), .B (n_2805), .C (n_2657), .D (n_3311), .Y(n_3312));
CLKBUFX1 gbuf_d_919(.A(n_3059), .Y(d_out_919));
CLKBUFX1 gbuf_q_919(.A(q_in_919), .Y(g1345));
AND2X1 g63719(.A (n_1264), .B (n_3430), .Y (n_3310));
CLKBUFX1 gbuf_d_920(.A(g26104), .Y(d_out_920));
CLKBUFX1 gbuf_qn_920(.A(qn_in_920), .Y(g3136));
CLKBUFX1 gbuf_d_921(.A(n_2890), .Y(d_out_921));
CLKBUFX1 gbuf_q_921(.A(q_in_921), .Y(g1384));
CLKBUFX1 gbuf_d_922(.A(n_2881), .Y(d_out_922));
CLKBUFX1 gbuf_q_922(.A(q_in_922), .Y(g1405));
CLKBUFX1 gbuf_d_923(.A(n_2879), .Y(d_out_923));
CLKBUFX1 gbuf_q_923(.A(q_in_923), .Y(g1408));
CLKBUFX1 gbuf_d_924(.A(n_2838), .Y(d_out_924));
CLKBUFX1 gbuf_q_924(.A(q_in_924), .Y(g2084));
CLKBUFX1 gbuf_d_925(.A(n_2837), .Y(d_out_925));
CLKBUFX1 gbuf_q_925(.A(q_in_925), .Y(g2087));
CLKBUFX1 gbuf_d_926(.A(n_2833), .Y(d_out_926));
CLKBUFX1 gbuf_q_926(.A(q_in_926), .Y(g2102));
OAI21X1 g62646(.A0 (n_3307), .A1 (g672), .B0 (n_2850), .Y (n_3308));
CLKBUFX1 gbuf_d_927(.A(n_2949), .Y(d_out_927));
CLKBUFX1 gbuf_q_927(.A(q_in_927), .Y(g1555));
CLKBUFX1 gbuf_d_928(.A(n_2944), .Y(d_out_928));
CLKBUFX1 gbuf_q_928(.A(q_in_928), .Y(g2255));
CLKBUFX1 gbuf_d_929(.A(n_2951), .Y(d_out_929));
CLKBUFX1 gbuf_q_929(.A(q_in_929), .Y(g1558));
MX2X1 g63941(.A (n_7273), .B (g1417), .S0 (n_3305), .Y (n_3306));
MX2X1 g63942(.A (n_7273), .B (g1418), .S0 (n_3303), .Y (n_3304));
MX2X1 g63943(.A (g1419), .B (n_7273), .S0 (n_4963), .Y (n_3302));
XOR2X1 g64011(.A (g2734), .B (n_2656), .Y (n_3301));
XOR2X1 g64013(.A (g2714), .B (n_2655), .Y (n_3300));
XOR2X1 g64030(.A (g2020), .B (n_2650), .Y (n_3299));
XOR2X1 g64031(.A (g2066), .B (n_2651), .Y (n_3298));
XOR2X1 g64032(.A (g1326), .B (n_2634), .Y (n_3296));
XOR2X1 g64046(.A (g666), .B (n_2633), .Y (n_3295));
XOR2X1 g64047(.A (g646), .B (n_2794), .Y (n_3294));
XOR2X1 g64049(.A (g672), .B (n_2648), .Y (n_3293));
XOR2X1 g64053(.A (g660), .B (n_2795), .Y (n_3292));
XOR2X1 g64054(.A (g633), .B (n_2638), .Y (n_3291));
CLKBUFX1 gbuf_d_930(.A(n_3290), .Y(d_out_930));
CLKBUFX1 gbuf_q_930(.A(q_in_930), .Y(gbuf200));
NAND2X1 g64182(.A (n_3288), .B (n_4515), .Y (n_3289));
NAND2X1 g64183(.A (n_3286), .B (n_4517), .Y (n_3287));
NAND2X1 g64184(.A (n_3284), .B (n_4517), .Y (n_3285));
NAND2X1 g64185(.A (n_3311), .B (n_4515), .Y (n_3283));
NAND2X1 g64186(.A (n_3281), .B (n_4517), .Y (n_3282));
NAND2X1 g64187(.A (n_3279), .B (n_4515), .Y (n_3280));
NAND2X1 g64188(.A (n_3277), .B (n_4517), .Y (n_3278));
NOR2X1 g64195(.A (n_2788), .B (n_2927), .Y (n_3276));
NOR2X1 g64210(.A (n_2629), .B (n_2927), .Y (n_3275));
NAND2X1 g64248(.A (n_3534), .B (n_3393), .Y (n_3412));
OAI21X1 g62637(.A0 (n_3307), .A1 (g653), .B0 (n_2844), .Y (n_3274));
CLKBUFX1 gbuf_d_931(.A(n_2835), .Y(d_out_931));
CLKBUFX1 gbuf_q_931(.A(q_in_931), .Y(g2099));
CLKBUFX1 gbuf_d_932(.A(g26104), .Y(d_out_932));
CLKBUFX1 gbuf_qn_932(.A(qn_in_932), .Y(g3142));
CLKBUFX1 gbuf_d_933(.A(g26104), .Y(d_out_933));
CLKBUFX1 gbuf_q_933(.A(q_in_933), .Y(g3207));
CLKBUFX1 gbuf_d_934(.A(g26104), .Y(d_out_934));
CLKBUFX1 gbuf_qn_934(.A(qn_in_934), .Y(g3132));
NOR2X1 g64417(.A (n_4078), .B (n_3534), .Y (n_3576));
CLKBUFX1 gbuf_d_935(.A(g26104), .Y(d_out_935));
CLKBUFX1 gbuf_q_935(.A(q_in_935), .Y(g3120));
CLKBUFX1 gbuf_d_936(.A(n_2945), .Y(d_out_936));
CLKBUFX1 gbuf_q_936(.A(q_in_936), .Y(g1561));
CLKBUFX1 gbuf_d_937(.A(n_2867), .Y(d_out_937));
CLKBUFX1 gbuf_q_937(.A(q_in_937), .Y(g1527));
CLKBUFX1 gbuf_d_938(.A(n_2865), .Y(d_out_938));
CLKBUFX1 gbuf_q_938(.A(q_in_938), .Y(g1528));
CLKBUFX1 gbuf_d_939(.A(n_2868), .Y(d_out_939));
CLKBUFX1 gbuf_q_939(.A(q_in_939), .Y(g1525));
CLKBUFX1 gbuf_d_940(.A(n_2873), .Y(d_out_940));
CLKBUFX1 gbuf_q_940(.A(q_in_940), .Y(g1515));
CLKBUFX1 gbuf_d_941(.A(n_2870), .Y(d_out_941));
CLKBUFX1 gbuf_q_941(.A(q_in_941), .Y(g1524));
AND2X1 g64622(.A (n_4078), .B (n_3533), .Y (n_3559));
CLKBUFX1 gbuf_d_942(.A(n_2872), .Y(d_out_942));
CLKBUFX1 gbuf_q_942(.A(q_in_942), .Y(g1516));
CLKBUFX1 gbuf_d_943(.A(n_2898), .Y(d_out_943));
CLKBUFX1 gbuf_q_943(.A(q_in_943), .Y(g1316));
AND2X1 g63807(.A (n_6451), .B (g6447), .Y (n_3271));
NOR2X1 g64711(.A (n_187), .B (n_3270), .Y (n_3381));
NOR2X1 g64714(.A (n_282), .B (n_3269), .Y (n_3380));
CLKBUFX1 gbuf_d_944(.A(n_2854), .Y(d_out_944));
CLKBUFX1 gbuf_q_944(.A(q_in_944), .Y(g_27738));
NAND2X2 g64869(.A (n_2895), .B (n_2316), .Y (n_4096));
AOI21X1 g64900(.A0 (n_2171), .A1 (n_3498), .B0 (n_2892), .Y (n_3531));
CLKBUFX1 gbuf_d_945(.A(n_2878), .Y(d_out_945));
CLKBUFX1 gbuf_q_945(.A(q_in_945), .Y(g1411));
AOI22X1 g65066(.A0 (n_2012), .A1 (n_3498), .B0 (g573), .B1 (n_4601),.Y (n_3547));
INVX1 g65069(.A (n_4737), .Y (n_3372));
AOI22X1 g65090(.A0 (n_2013), .A1 (n_3264), .B0 (g1991), .B1 (n_6626),.Y (n_4317));
AOI21X1 g65178(.A0 (n_2166), .A1 (n_2925), .B0 (n_2882), .Y (n_3548));
AOI22X1 g65181(.A0 (n_2393), .A1 (n_3093), .B0 (g1183), .B1 (n_5270),.Y (n_3263));
AOI22X1 g65335(.A0 (n_2379), .A1 (n_3498), .B0 (g489), .B1 (n_4601),.Y (n_3549));
XOR2X1 g65366(.A (g2013), .B (n_3082), .Y (n_3255));
XOR2X1 g65367(.A (g633), .B (n_3079), .Y (n_3254));
XOR2X1 g65369(.A (g1319), .B (n_3080), .Y (n_3253));
NAND2X1 g65435(.A (n_3251), .B (n_3835), .Y (n_3252));
AOI21X1 g65667(.A0 (n_1912), .A1 (n_3498), .B0 (n_2896), .Y (n_3684));
INVX1 g65557(.A (n_3249), .Y (n_3516));
INVX1 g65611(.A (n_3378), .Y (n_3364));
AOI21X1 g65630(.A0 (n_1731), .A1 (n_3264), .B0 (n_2893), .Y (n_3363));
CLKBUFX1 gbuf_d_946(.A(n_2830), .Y(d_out_946));
CLKBUFX1 gbuf_q_946(.A(q_in_946), .Y(g2096));
INVX1 g65674(.A (n_3530), .Y (n_3359));
INVX1 g65680(.A (n_4104), .Y (n_3842));
INVX1 g65720(.A (n_3382), .Y (n_3515));
INVX1 g65725(.A (n_3736), .Y (n_4102));
NAND2X2 g65637(.A (n_2894), .B (n_2016), .Y (n_4116));
INVX1 g65798(.A (n_3524), .Y (n_3415));
CLKBUFX1 gbuf_d_947(.A(n_2836), .Y(d_out_947));
CLKBUFX1 gbuf_q_947(.A(q_in_947), .Y(g2093));
NAND2X1 g65919(.A (n_2877), .B (n_5044), .Y (n_3237));
NAND2X1 g65925(.A (n_2876), .B (n_4604), .Y (n_3236));
CLKBUFX1 gbuf_d_948(.A(n_2831), .Y(d_out_948));
CLKBUFX1 gbuf_q_948(.A(q_in_948), .Y(g2105));
AOI22X1 g65982(.A0 (n_2704), .A1 (g354), .B0 (g343), .B1 (n_1237), .Y(n_3235));
AND2X1 g63805(.A (n_5885), .B (n_2180), .Y (n_3233));
CLKBUFX1 gbuf_d_949(.A(n_2953), .Y(d_out_949));
CLKBUFX1 gbuf_q_949(.A(q_in_949), .Y(g2246));
AOI22X1 g66079(.A0 (n_2709), .A1 (g2523), .B0 (g2524), .B1 (n_9512),.Y (n_3232));
MX2X1 g66119(.A (n_3701), .B (g630), .S0 (n_2814), .Y (n_3231));
MX2X1 g66124(.A (n_4050), .B (g2704), .S0 (n_2674), .Y (n_3229));
CLKBUFX1 gbuf_d_950(.A(n_2832), .Y(d_out_950));
CLKBUFX1 gbuf_q_950(.A(q_in_950), .Y(g2090));
CLKBUFX1 gbuf_d_951(.A(n_2947), .Y(d_out_951));
CLKBUFX1 gbuf_q_951(.A(q_in_951), .Y(g1552));
INVX1 g66300(.A (n_3107), .Y (n_3227));
CLKBUFX1 gbuf_d_952(.A(n_2900), .Y(d_out_952));
CLKBUFX1 gbuf_q_952(.A(q_in_952), .Y(g2010));
OR2X1 g66389(.A (n_255), .B (n_3224), .Y (n_3225));
OR2X1 g66394(.A (g1171), .B (n_3220), .Y (n_3222));
OR2X1 g66400(.A (g1174), .B (n_3220), .Y (n_3221));
INVX1 g66448(.A (n_3040), .Y (n_8368));
NOR2X1 g66472(.A (g1964), .B (g1930), .Y (n_3218));
OR2X1 g66496(.A (g2250), .B (n_3224), .Y (n_3217));
AOI22X1 g63899(.A0 (n_2624), .A1 (n_2834), .B0 (n_3544), .B1 (n_245),.Y (n_3216));
NAND2X1 g66562(.A (n_3220), .B (n_1660), .Y (n_4262));
OAI21X1 g62631(.A0 (n_3307), .A1 (g640), .B0 (n_2849), .Y (n_3213));
OAI21X1 g62634(.A0 (n_3307), .A1 (g633), .B0 (n_2842), .Y (n_3212));
INVX4 g66840(.A (g1547), .Y (n_3467));
OAI21X1 g62640(.A0 (n_3307), .A1 (g646), .B0 (n_2846), .Y (n_3207));
OAI21X1 g62643(.A0 (n_3307), .A1 (g660), .B0 (n_2852), .Y (n_3206));
OAI21X1 g62649(.A0 (n_3307), .A1 (g666), .B0 (n_2853), .Y (n_3205));
OAI21X1 g62652(.A0 (n_3307), .A1 (n_3203), .B0 (n_2851), .Y (n_3204));
OAI21X1 g62655(.A0 (n_3307), .A1 (g686), .B0 (n_2845), .Y (n_3202));
OAI21X1 g62658(.A0 (n_3307), .A1 (g692), .B0 (n_2843), .Y (n_3201));
NAND2X1 g67001(.A (g243), .B (n_3195), .Y (n_3200));
NAND2X1 g67022(.A (g2391), .B (n_2736), .Y (n_3199));
NAND2X1 g67074(.A (g270), .B (n_3195), .Y (n_8228));
NAND2X1 g67161(.A (g_26724), .B (n_3195), .Y (n_8260));
NAND2X1 g67186(.A (g_30665), .B (n_3195), .Y (n_3194));
NAND2X1 g67213(.A (g234), .B (n_3195), .Y (n_9595));
MX2X1 g62758(.A (n_3187), .B (g_16484), .S0 (n_5585), .Y (n_3188));
MX2X1 g62760(.A (g105), .B (g_24593), .S0 (n_5585), .Y (n_3180));
MX2X1 g62761(.A (n_5247), .B (g_19132), .S0 (n_5585), .Y (n_3178));
MX2X1 g62768(.A (n_4112), .B (g818), .S0 (n_4540), .Y (n_3176));
MX2X1 g62769(.A (n_4112), .B (g819), .S0 (n_4538), .Y (n_3175));
MX2X1 g62771(.A (n_4110), .B (g821), .S0 (n_4540), .Y (n_3174));
MX2X1 g62772(.A (n_4110), .B (g822), .S0 (n_4538), .Y (n_3173));
MX2X1 g62774(.A (n_3171), .B (g831), .S0 (n_4538), .Y (n_3172));
MX2X1 g62776(.A (n_3169), .B (g833), .S0 (n_4540), .Y (n_3170));
MX2X1 g62778(.A (n_3167), .B (g836), .S0 (n_4540), .Y (n_3168));
MX2X1 g62779(.A (n_3167), .B (g837), .S0 (n_4538), .Y (n_3166));
MX2X1 g62783(.A (n_3164), .B (g842), .S0 (n_4540), .Y (n_3165));
MX2X1 g62784(.A (n_3164), .B (g843), .S0 (n_4538), .Y (n_3163));
MX2X1 g62788(.A (n_3161), .B (g_19162), .S0 (n_5585), .Y (n_3162));
MX2X1 g62790(.A (n_3169), .B (g834), .S0 (n_4538), .Y (n_3160));
MX2X1 g62793(.A (n_3171), .B (g830), .S0 (n_4540), .Y (n_3159));
MX2X1 g62798(.A (n_5382), .B (g_14855), .S0 (n_5585), .Y (n_3158));
MX2X1 g62801(.A (n_5380), .B (g_20947), .S0 (n_5585), .Y (n_3157));
CLKBUFX1 gbuf_d_953(.A(n_2883), .Y(d_out_953));
CLKBUFX1 gbuf_q_953(.A(q_in_953), .Y(g1402));
CLKBUFX1 gbuf_d_954(.A(n_2841), .Y(d_out_954));
CLKBUFX1 gbuf_q_954(.A(q_in_954), .Y(g2078));
XOR2X1 g63900(.A (g2740), .B (n_2658), .Y (n_3156));
NOR2X1 g63227(.A (n_2967), .B (n_2828), .Y (n_3155));
INVX1 g66375(.A (n_3042), .Y (n_8366));
OR2X1 g66382(.A (g1165), .B (n_3220), .Y (n_3153));
OAI21X1 g63302(.A0 (n_3151), .A1 (g2714), .B0 (n_2984), .Y (n_3152));
OAI21X1 g63305(.A0 (n_3151), .A1 (g2707), .B0 (n_2983), .Y (n_3150));
OAI21X1 g63308(.A0 (n_3151), .A1 (g2727), .B0 (n_2982), .Y (n_3149));
OAI21X1 g63311(.A0 (n_3151), .A1 (g2720), .B0 (n_2981), .Y (n_3148));
OAI21X1 g63314(.A0 (n_3151), .A1 (g2734), .B0 (n_2980), .Y (n_3147));
OAI21X1 g63317(.A0 (n_3151), .A1 (g2746), .B0 (n_2979), .Y (n_3146));
OAI21X1 g63319(.A0 (n_3151), .A1 (g2740), .B0 (n_2978), .Y (n_3145));
OAI21X1 g63322(.A0 (n_3151), .A1 (n_3143), .B0 (n_2977), .Y (n_3144));
CLKBUFX1 gbuf_d_955(.A(n_2884), .Y(d_out_955));
CLKBUFX1 gbuf_q_955(.A(q_in_955), .Y(g1399));
OAI21X1 g63326(.A0 (n_3151), .A1 (g2760), .B0 (n_2976), .Y (n_3142));
OAI21X1 g63329(.A0 (n_3151), .A1 (g2766), .B0 (n_2975), .Y (n_3141));
CLKBUFX1 gbuf_d_956(.A(n_2888), .Y(d_out_956));
CLKBUFX1 gbuf_q_956(.A(q_in_956), .Y(g1387));
CLKBUFX1 gbuf_d_957(.A(n_2885), .Y(d_out_957));
CLKBUFX1 gbuf_q_957(.A(q_in_957), .Y(g1396));
INVX1 g66363(.A (n_3044), .Y (n_3140));
AND2X1 g63458(.A (n_2957), .B (n_3281), .Y (n_3139));
CLKBUFX1 gbuf_d_958(.A(n_2857), .Y(d_out_958));
CLKBUFX1 gbuf_q_958(.A(q_in_958), .Y(g_15404));
CLKBUFX1 gbuf_d_959(.A(n_2886), .Y(d_out_959));
CLKBUFX1 gbuf_q_959(.A(q_in_959), .Y(g1393));
NAND3X1 g63578(.A (n_2940), .B (n_2649), .C (n_2941), .Y (n_3138));
CLKBUFX1 gbuf_d_960(.A(n_2887), .Y(d_out_960));
CLKBUFX1 gbuf_q_960(.A(q_in_960), .Y(g1390));
CLKBUFX1 gbuf_d_961(.A(n_2839), .Y(d_out_961));
CLKBUFX1 gbuf_q_961(.A(q_in_961), .Y(g2081));
NAND3X1 g63769(.A (n_3136), .B (n_2615), .C (n_2785), .Y (n_3137));
NOR2X1 g63775(.A (n_2818), .B (n_2638), .Y (n_9569));
NOR2X1 g63782(.A (n_2820), .B (n_2651), .Y (n_3134));
AND2X1 g63783(.A (n_2822), .B (n_2626), .Y (n_3133));
CLKBUFX1 gbuf_d_962(.A(n_2689), .Y(d_out_962));
CLKBUFX1 gbuf_q_962(.A(q_in_962), .Y(g_24187));
CLKBUFX1 gbuf_d_963(.A(n_2813), .Y(d_out_963));
CLKBUFX1 gbuf_q_963(.A(q_in_963), .Y(g1425));
CLKBUFX1 gbuf_d_964(.A(n_2723), .Y(d_out_964));
CLKBUFX1 gbuf_q_964(.A(q_in_964), .Y(g2207));
CLKBUFX1 gbuf_d_965(.A(n_2693), .Y(d_out_965));
CLKBUFX1 gbuf_q_965(.A(q_in_965), .Y(g_5844));
CLKBUFX1 gbuf_d_966(.A(n_2808), .Y(d_out_966));
CLKBUFX1 gbuf_q_966(.A(q_in_966), .Y(g2252));
CLKBUFX1 gbuf_d_967(.A(n_2692), .Y(d_out_967));
CLKBUFX1 gbuf_q_967(.A(q_in_967), .Y(g_29016));
XOR2X1 g64009(.A (g2766), .B (n_2803), .Y (n_3131));
XOR2X1 g64010(.A (g2760), .B (n_3129), .Y (n_3130));
XOR2X1 g64014(.A (g2727), .B (n_2654), .Y (n_3128));
XOR2X1 g64015(.A (g1332), .B (n_2636), .Y (n_3127));
XOR2X1 g64021(.A (g1358), .B (n_2639), .Y (n_3126));
XOR2X1 g64022(.A (g1378), .B (n_2790), .Y (n_3125));
XOR2X1 g64027(.A (g1352), .B (n_2629), .Y (n_3124));
XOR2X1 g64038(.A (g2013), .B (n_2631), .Y (n_3123));
XOR2X1 g64044(.A (g2026), .B (n_2627), .Y (n_3122));
XOR2X1 g64045(.A (g2052), .B (n_2632), .Y (n_3121));
XOR2X1 g64050(.A (g653), .B (n_2647), .Y (n_3120));
XOR2X1 g64056(.A (g2072), .B (n_2784), .Y (n_3119));
XOR2X1 g64076(.A (g2046), .B (n_2623), .Y (n_3118));
XOR2X1 g64078(.A (g2033), .B (n_2652), .Y (n_3117));
XOR2X1 g64079(.A (g2720), .B (n_2621), .Y (n_3116));
AND2X1 g64194(.A (n_3114), .B (n_7273), .Y (n_3115));
AND2X1 g64203(.A (n_3112), .B (n_7273), .Y (n_3113));
AND2X1 g64222(.A (n_3110), .B (n_7273), .Y (n_3111));
CLKBUFX1 gbuf_d_968(.A(n_2688), .Y(d_out_968));
CLKBUFX1 gbuf_q_968(.A(q_in_968), .Y(g_26130));
NOR2X1 g64224(.A (n_3108), .B (n_4689), .Y (n_3109));
NOR2X1 g66301(.A (g820), .B (n_4162), .Y (n_3107));
NOR2X1 g64245(.A (n_4078), .B (n_2929), .Y (n_3430));
NAND2X1 g64272(.A (n_4151), .B (n_7273), .Y (n_3106));
CLKBUFX1 gbuf_d_969(.A(n_2722), .Y(d_out_969));
CLKBUFX1 gbuf_q_969(.A(q_in_969), .Y(g2210));
CLKBUFX1 gbuf_d_970(.A(n_2690), .Y(d_out_970));
CLKBUFX1 gbuf_q_970(.A(q_in_970), .Y(g_20789));
AOI21X1 g65726(.A0 (n_1909), .A1 (n_3093), .B0 (n_2744), .Y (n_3736));
CLKBUFX1 gbuf_d_971(.A(n_2707), .Y(d_out_971));
CLKBUFX1 gbuf_q_971(.A(q_in_971), .Y(g2234));
NOR2X1 g66223(.A (n_89), .B (n_4162), .Y (n_3103));
CLKBUFX1 gbuf_d_972(.A(n_2712), .Y(d_out_972));
CLKBUFX1 gbuf_q_972(.A(q_in_972), .Y(g2228));
CLKBUFX1 gbuf_d_973(.A(n_2703), .Y(d_out_973));
CLKBUFX1 gbuf_q_973(.A(q_in_973), .Y(g2209));
CLKBUFX1 gbuf_d_974(.A(n_2714), .Y(d_out_974));
CLKBUFX1 gbuf_q_974(.A(q_in_974), .Y(g2227));
CLKBUFX1 gbuf_d_975(.A(n_2710), .Y(d_out_975));
CLKBUFX1 gbuf_q_975(.A(q_in_975), .Y(g2233));
CLKBUFX1 gbuf_d_976(.A(n_2702), .Y(d_out_976));
CLKBUFX1 gbuf_q_976(.A(q_in_976), .Y(g2230));
CLKBUFX1 gbuf_d_977(.A(n_2711), .Y(d_out_977));
CLKBUFX1 gbuf_q_977(.A(q_in_977), .Y(g2231));
CLKBUFX1 gbuf_d_978(.A(n_2715), .Y(d_out_978));
CLKBUFX1 gbuf_q_978(.A(q_in_978), .Y(g2225));
CLKBUFX1 gbuf_d_979(.A(n_2735), .Y(d_out_979));
CLKBUFX1 gbuf_q_979(.A(q_in_979), .Y(g2219));
OAI21X1 g62627(.A0 (n_4973), .A1 (g1501), .B0 (n_2680), .Y (n_3096));
OAI21X1 g62628(.A0 (n_4971), .A1 (g1501), .B0 (n_2679), .Y (n_3094));
CLKBUFX1 gbuf_d_980(.A(n_2717), .Y(d_out_980));
CLKBUFX1 gbuf_q_980(.A(q_in_980), .Y(g2224));
AOI21X1 g64982(.A0 (n_1920), .A1 (n_3093), .B0 (n_2826), .Y (n_3525));
INVX1 g65011(.A (n_3534), .Y (n_3394));
CLKBUFX1 gbuf_d_981(.A(n_2733), .Y(d_out_981));
CLKBUFX1 gbuf_q_981(.A(q_in_981), .Y(g2218));
CLKBUFX1 gbuf_d_982(.A(n_2720), .Y(d_out_982));
CLKBUFX1 gbuf_q_982(.A(q_in_982), .Y(g2221));
AOI22X1 g65070(.A0 (n_2313), .A1 (n_3498), .B0 (g620), .B1 (g550), .Y(n_4737));
CLKBUFX1 gbuf_d_983(.A(n_2718), .Y(d_out_983));
CLKBUFX1 gbuf_q_983(.A(q_in_983), .Y(g2222));
CLKBUFX1 gbuf_d_984(.A(n_2724), .Y(d_out_984));
CLKBUFX1 gbuf_q_984(.A(q_in_984), .Y(g2206));
AOI22X1 g65191(.A0 (n_2040), .A1 (n_3093), .B0 (g1259), .B1 (n_5270),.Y (n_3398));
AOI22X1 g65196(.A0 (n_2382), .A1 (n_3093), .B0 (g1176), .B1 (n_5270),.Y (n_3397));
INVX1 g65267(.A (n_4515), .Y (n_3260));
AOI21X1 g65292(.A0 (n_2018), .A1 (n_3498), .B0 (n_2750), .Y (n_5101));
OAI21X1 g62624(.A0 (n_4971), .A1 (n_471), .B0 (n_2681), .Y (n_3089));
INVX1 g65341(.A (n_4517), .Y (n_3256));
INVX1 g67726(.A (n_2736), .Y (n_3085));
NAND2X1 g65683(.A (n_2746), .B (n_2175), .Y (n_4104));
NAND2X1 g65451(.A (n_3082), .B (n_3664), .Y (n_3083));
CLKBUFX1 gbuf_d_985(.A(n_2810), .Y(d_out_985));
CLKBUFX1 gbuf_q_985(.A(q_in_985), .Y(g2249));
NAND2X1 g65529(.A (n_3080), .B (n_3678), .Y (n_3081));
NOR2X1 g65558(.A (n_269), .B (n_3079), .Y (n_3249));
INVX1 g65570(.A (n_3269), .Y (n_3245));
CLKBUFX1 gbuf_d_986(.A(n_2812), .Y(d_out_986));
CLKBUFX1 gbuf_q_986(.A(q_in_986), .Y(g858));
OAI21X1 g62620(.A0 (n_4971), .A1 (n_600), .B0 (n_2682), .Y (n_3078));
AOI21X1 g65676(.A0 (n_1914), .A1 (n_3498), .B0 (n_2749), .Y (n_3530));
AOI21X1 g65721(.A0 (n_1605), .A1 (n_3093), .B0 (n_2745), .Y (n_3382));
INVX2 g65773(.A (n_3533), .Y (n_3239));
INVX1 g65799(.A (n_3075), .Y (n_3524));
OAI21X1 g62288(.A0 (n_2753), .A1 (g1316), .B0 (n_2754), .Y (n_3074));
NOR2X1 g65872(.A (n_1118), .B (n_2739), .Y (n_3073));
NOR2X1 g65874(.A (n_1104), .B (n_2741), .Y (n_3072));
NOR2X1 g65914(.A (n_1135), .B (n_2742), .Y (n_3069));
NAND2X1 g65924(.A (n_2737), .B (n_4604), .Y (n_3068));
AOI22X1 g66022(.A0 (n_2570), .A1 (g_24794), .B0 (g_26381), .B1(n_1382), .Y (n_3066));
NAND2X1 g62407(.A (n_3064), .B (g737), .Y (n_3065));
AOI22X1 g66074(.A0 (n_2571), .A1 (g2429), .B0 (g2418), .B1 (n_9512),.Y (n_3063));
AOI22X1 g66087(.A0 (n_2593), .A1 (g1735), .B0 (g1724), .B1 (n_1235),.Y (n_3061));
OAI21X1 g66102(.A0 (n_4151), .A1 (n_2410), .B0 (n_2743), .Y (n_3059));
OAI21X1 g66108(.A0 (n_4151), .A1 (n_2292), .B0 (n_2747), .Y (n_3058));
NOR2X1 g66209(.A (n_118), .B (n_4162), .Y (n_3057));
NAND2X1 g66213(.A (g2667), .B (n_2863), .Y (n_3056));
NOR2X1 g66236(.A (n_68), .B (n_4162), .Y (n_3055));
OR2X1 g66263(.A (n_52), .B (n_4162), .Y (n_3053));
NOR2X1 g66282(.A (n_107), .B (n_4162), .Y (n_3052));
NOR2X1 g66283(.A (g862), .B (n_4162), .Y (n_3051));
NAND3X1 g65612(.A (n_2905), .B (g2707), .C (g2727), .Y (n_3378));
NAND2X1 g66319(.A (g2733), .B (n_2674), .Y (n_3047));
NOR2X1 g66333(.A (n_27), .B (n_4162), .Y (n_3046));
NAND2X1 g66343(.A (n_6626), .B (g2000), .Y (n_3045));
NOR2X1 g66364(.A (g835), .B (n_4162), .Y (n_3044));
NOR2X1 g66376(.A (g832), .B (n_4162), .Y (n_3042));
NOR2X1 g66445(.A (g859), .B (n_4162), .Y (n_3041));
NOR2X1 g66449(.A (g817), .B (n_4162), .Y (n_3040));
NOR2X1 g66454(.A (n_4162), .B (n_81), .Y (n_3039));
AOI22X1 g66523(.A0 (n_1315), .A1 (g388), .B0 (g398), .B1 (n_2874), .Y(n_3038));
AOI22X1 g66533(.A0 (n_1314), .A1 (g1769), .B0 (g1779), .B1 (n_3036),.Y (n_3037));
AOI22X1 g66601(.A0 (n_1288), .A1 (g1754), .B0 (g1765), .B1 (n_3036),.Y (n_3035));
OAI21X1 g62608(.A0 (n_4973), .A1 (g1471), .B0 (n_2675), .Y (n_3034));
OAI21X1 g62609(.A0 (n_4971), .A1 (g1471), .B0 (n_2684), .Y (n_3032));
OAI21X1 g62621(.A0 (n_4973), .A1 (n_600), .B0 (n_2683), .Y (n_3031));
OAI21X1 g62623(.A0 (n_4973), .A1 (n_471), .B0 (n_2676), .Y (n_3029));
CLKBUFX3 g66753(.A (n_3224), .Y (n_3344));
OAI21X1 g62630(.A0 (n_4973), .A1 (n_473), .B0 (n_2678), .Y (n_3027));
INVX2 g66934(.A (g1088), .Y (n_3336));
OAI21X1 g62682(.A0 (n_4971), .A1 (n_473), .B0 (n_2677), .Y (n_3023));
OAI21X1 g62683(.A0 (n_2685), .A1 (g2010), .B0 (n_2686), .Y (n_3022));
CLKBUFX1 gbuf_d_987(.A(n_2762), .Y(d_out_987));
CLKBUFX1 gbuf_q_987(.A(q_in_987), .Y(g1424));
INVX1 g67756(.A (n_3195), .Y (n_8028));
INVX1 g65567(.A (n_3270), .Y (n_3247));
NAND2X1 g62939(.A (n_3010), .B (g2811), .Y (n_3011));
NAND2X1 g63089(.A (n_4540), .B (g839), .Y (n_3009));
NAND2X1 g63090(.A (n_4540), .B (g845), .Y (n_3008));
NAND2X1 g63091(.A (n_4538), .B (g846), .Y (n_3007));
NAND2X1 g63092(.A (n_4540), .B (g848), .Y (n_3006));
NAND2X1 g63093(.A (n_4538), .B (g849), .Y (n_3005));
NAND2X1 g63095(.A (n_4540), .B (g851), .Y (n_3004));
NAND2X1 g63102(.A (n_5585), .B (g_30039), .Y (n_3003));
NAND2X1 g63137(.A (n_4538), .B (g840), .Y (n_3002));
NAND2X1 g63145(.A (n_5585), .B (g_23514), .Y (n_3001));
NAND2X1 g63148(.A (n_4538), .B (g852), .Y (n_3000));
NAND2X1 g63159(.A (n_5585), .B (g_23490), .Y (n_2999));
NAND2X1 g63166(.A (n_5585), .B (g_24922), .Y (n_2998));
INVX1 g67504(.A (n_3036), .Y (n_3190));
INVX1 g63532(.A (n_2829), .Y (n_2996));
NOR2X1 g63549(.A (n_2824), .B (n_2993), .Y (n_2994));
NOR2X1 g63554(.A (n_2817), .B (n_2625), .Y (n_2992));
NOR2X1 g63558(.A (n_2819), .B (n_2990), .Y (n_2991));
NAND2X1 g66351(.A (n_2814), .B (g659), .Y (n_2989));
CLKBUFX1 gbuf_d_988(.A(n_2691), .Y(d_out_988));
CLKBUFX1 gbuf_q_988(.A(q_in_988), .Y(g_7184));
OR2X1 g66345(.A (n_18), .B (n_4162), .Y (n_2988));
NAND2X1 g63723(.A (n_2986), .B (n_2985), .Y (n_2987));
NAND2X1 g63733(.A (n_3151), .B (g2772), .Y (n_2984));
NAND2X1 g63736(.A (n_3151), .B (g2775), .Y (n_2983));
NAND2X1 g63740(.A (n_3151), .B (g2778), .Y (n_2982));
NAND2X1 g63742(.A (n_3151), .B (g2781), .Y (n_2981));
NAND2X1 g63744(.A (n_3151), .B (g2784), .Y (n_2980));
NAND2X1 g63746(.A (n_3151), .B (g2787), .Y (n_2979));
NAND2X1 g63750(.A (n_3151), .B (g2790), .Y (n_2978));
NAND2X1 g63752(.A (n_3151), .B (g2793), .Y (n_2977));
NAND2X1 g63755(.A (n_3151), .B (g2796), .Y (n_2976));
NAND2X1 g63757(.A (n_3151), .B (g2799), .Y (n_2975));
NAND2X1 g63762(.A (n_3151), .B (n_2973), .Y (n_2974));
NOR2X1 g63772(.A (g996), .B (n_8305), .Y (n_2972));
NOR2X1 g63774(.A (g996), .B (n_2343), .Y (n_2969));
NAND3X1 g63777(.A (n_4285), .B (n_2512), .C (n_2634), .Y (n_2967));
CLKBUFX1 gbuf_d_989(.A(g6712), .Y(d_out_989));
CLKBUFX1 gbuf_q_989(.A(q_in_989), .Y(g1088));
CLKBUFX1 gbuf_d_990(.A(n_2665), .Y(d_out_990));
CLKBUFX1 gbuf_q_990(.A(q_in_990), .Y(g861));
XOR2X1 g64028(.A (g1339), .B (n_2511), .Y (n_2964));
XOR2X1 g64033(.A (g1319), .B (n_2509), .Y (n_2963));
XOR2X1 g64048(.A (g692), .B (n_2645), .Y (n_2962));
XOR2X1 g64051(.A (g686), .B (n_2641), .Y (n_2961));
XOR2X1 g64077(.A (n_2959), .B (n_3114), .Y (n_2960));
NOR2X1 g64226(.A (n_2614), .B (n_3114), .Y (n_2958));
NOR2X1 g64271(.A (n_2956), .B (n_2779), .Y (n_2957));
XOR2X1 g63897(.A (g1372), .B (n_2637), .Y (n_2954));
OAI21X1 g64486(.A0 (n_2952), .A1 (n_2943), .B0 (n_2660), .Y (n_2953));
MX2X1 g64497(.A (g1558), .B (n_365), .S0 (n_2948), .Y (n_2951));
MX2X1 g64503(.A (g1555), .B (n_364), .S0 (n_2948), .Y (n_2949));
MX2X1 g64504(.A (g1552), .B (n_2946), .S0 (n_2948), .Y (n_2947));
MX2X1 g64537(.A (g1561), .B (n_4861), .S0 (n_2948), .Y (n_2945));
OAI21X1 g64546(.A0 (n_4674), .A1 (n_2943), .B0 (n_2659), .Y (n_2944));
INVX4 g66771(.A (g2241), .Y (n_3224));
CLKBUFX1 gbuf_d_991(.A(n_2662), .Y(d_out_991));
CLKBUFX1 gbuf_q_991(.A(q_in_991), .Y(g867));
INVX1 g64795(.A (n_2941), .Y (n_4695));
INVX1 g64798(.A (n_2940), .Y (n_4681));
INVX1 g66745(.A (n_4162), .Y (n_3589));
INVX2 g65014(.A (n_2929), .Y (n_3534));
AOI21X1 g65268(.A0 (n_1926), .A1 (n_2925), .B0 (n_2586), .Y (n_4515));
INVX1 g65269(.A (n_7271), .Y (n_2927));
AOI21X1 g65342(.A0 (n_1631), .A1 (n_2925), .B0 (n_2588), .Y (n_4517));
AOI22X1 g65348(.A0 (n_1753), .A1 (n_2925), .B0 (g2647), .B1 (n_2863),.Y (n_3290));
NAND3X1 g65424(.A (n_9647), .B (n_937), .C (n_2921), .Y (n_2922));
AND2X1 g65432(.A (n_2601), .B (n_5044), .Y (n_2920));
NAND2X1 g65496(.A (n_2591), .B (n_5044), .Y (n_2917));
NAND2X1 g65517(.A (n_2605), .B (n_2408), .Y (n_2916));
NOR2X1 g65521(.A (n_2915), .B (n_3195), .Y (n_3387));
NAND3X1 g65568(.A (n_2760), .B (g2013), .C (g2033), .Y (n_3270));
NAND3X1 g65571(.A (n_2757), .B (g1319), .C (g1339), .Y (n_3269));
AOI21X1 g65774(.A0 (n_1506), .A1 (n_2925), .B0 (n_2585), .Y (n_3533));
INVX1 g65783(.A (n_2986), .Y (n_3393));
OAI21X1 g65800(.A0 (g1267), .A1 (n_2499), .B0 (n_1922), .Y (n_3075));
NOR2X1 g65830(.A (n_1100), .B (n_2576), .Y (n_2913));
INVX1 g65886(.A (n_3079), .Y (n_3070));
NAND2X1 g65895(.A (n_2360), .B (n_3810), .Y (n_2910));
NOR2X1 g65928(.A (n_1120), .B (n_2581), .Y (n_2909));
NOR2X1 g65933(.A (n_1143), .B (n_2584), .Y (n_2908));
NAND2X1 g65945(.A (n_2356), .B (n_3810), .Y (n_2907));
INVX1 g65950(.A (n_2905), .Y (n_3251));
NOR2X1 g65952(.A (n_1211), .B (n_2578), .Y (n_2904));
NOR2X1 g65956(.A (n_1099), .B (n_2582), .Y (n_2903));
NOR2X1 g65959(.A (n_1116), .B (n_2583), .Y (n_2902));
AOI22X1 g66034(.A0 (n_2439), .A1 (g427), .B0 (g428), .B1 (n_1237), .Y(n_2901));
MX2X1 g66121(.A (n_5322), .B (g2010), .S0 (n_2292), .Y (n_2900));
MX2X1 g66123(.A (n_3698), .B (g1316), .S0 (n_2410), .Y (n_2898));
NOR2X1 g66247(.A (g581), .B (n_2748), .Y (n_2896));
OR2X1 g66261(.A (g1955), .B (g1930), .Y (n_2895));
OR2X1 g66262(.A (g1958), .B (g1930), .Y (n_2894));
NOR2X1 g66438(.A (g1961), .B (g1930), .Y (n_2893));
NOR2X1 g66315(.A (g575), .B (n_2748), .Y (n_2892));
NAND2X1 g66326(.A (n_2264), .B (g630), .Y (n_3554));
NAND2X1 g66451(.A (g2704), .B (n_2451), .Y (n_4302));
OAI21X1 g62566(.A0 (n_2889), .A1 (g1326), .B0 (n_2551), .Y (n_2890));
OAI21X1 g62571(.A0 (n_2889), .A1 (g1319), .B0 (n_2550), .Y (n_2888));
OAI21X1 g62574(.A0 (n_2889), .A1 (g1339), .B0 (n_2549), .Y (n_2887));
OAI21X1 g62577(.A0 (n_2889), .A1 (g1332), .B0 (n_2548), .Y (n_2886));
OAI21X1 g62580(.A0 (n_2889), .A1 (g1346), .B0 (n_2547), .Y (n_2885));
OAI21X1 g62583(.A0 (n_2889), .A1 (g1358), .B0 (n_2546), .Y (n_2884));
OAI21X1 g62586(.A0 (n_2889), .A1 (g1352), .B0 (n_2545), .Y (n_2883));
NOR2X1 g66546(.A (g2564), .B (n_3448), .Y (n_2882));
OAI21X1 g62589(.A0 (n_2889), .A1 (n_2880), .B0 (n_2544), .Y (n_2881));
OAI21X1 g62592(.A0 (n_2889), .A1 (g1372), .B0 (n_2543), .Y (n_2879));
OAI21X1 g62595(.A0 (n_2889), .A1 (g1378), .B0 (n_2542), .Y (n_2878));
AOI22X1 g66575(.A0 (n_1238), .A1 (g358), .B0 (g369), .B1 (n_2874), .Y(n_2877));
AOI22X1 g66578(.A0 (n_1313), .A1 (g2463), .B0 (g2473), .B1 (n_2736),.Y (n_2876));
AOI22X1 g66588(.A0 (n_1253), .A1 (g373), .B0 (g384), .B1 (n_2874), .Y(n_2875));
MX2X1 g62611(.A (n_364), .B (g1515), .S0 (n_4973), .Y (n_2873));
MX2X1 g62612(.A (n_364), .B (g1516), .S0 (n_4971), .Y (n_2872));
MX2X1 g62614(.A (n_435), .B (g1524), .S0 (n_4973), .Y (n_2870));
MX2X1 g62615(.A (n_435), .B (g1525), .S0 (n_4971), .Y (n_2868));
MX2X1 g62617(.A (n_454), .B (g1527), .S0 (n_4973), .Y (n_2867));
MX2X1 g62618(.A (n_454), .B (g1528), .S0 (n_4971), .Y (n_2865));
CLKBUFX1 gbuf_d_992(.A(n_2663), .Y(d_out_992));
CLKBUFX1 gbuf_q_992(.A(q_in_992), .Y(g864));
CLKBUFX1 gbuf_d_993(.A(g6782), .Y(d_out_993));
CLKBUFX1 gbuf_q_993(.A(q_in_993), .Y(g1547));
NAND3X1 g61068(.A (n_2539), .B (n_1090), .C (n_1169), .Y (g26104));
OR2X1 g67107(.A (g1830), .B (n_3036), .Y (n_2862));
OR2X1 g67122(.A (g449), .B (n_2874), .Y (n_2861));
AND2X1 g63822(.A (n_6209), .B (g5511), .Y (n_2859));
OAI21X1 g62763(.A0 (n_5587), .A1 (n_733), .B0 (n_2538), .Y (n_2857));
OAI21X1 g62792(.A0 (n_5587), .A1 (g125), .B0 (n_2537), .Y (n_2854));
NAND2X1 g63018(.A (n_3307), .B (g716), .Y (n_2853));
NAND2X1 g63022(.A (n_3307), .B (g710), .Y (n_2852));
NAND2X1 g63024(.A (n_3307), .B (g719), .Y (n_2851));
NAND2X1 g63027(.A (n_3307), .B (g713), .Y (n_2850));
NAND2X1 g63073(.A (n_3307), .B (g698), .Y (n_2849));
NAND2X1 g63084(.A (n_3307), .B (n_2847), .Y (n_2848));
NAND2X1 g63099(.A (n_3307), .B (g707), .Y (n_2846));
NAND2X1 g63132(.A (n_3307), .B (g722), .Y (n_2845));
NAND2X1 g63134(.A (n_3307), .B (g704), .Y (n_2844));
NAND2X1 g63142(.A (n_3307), .B (g725), .Y (n_2843));
NAND2X1 g63147(.A (n_3307), .B (g701), .Y (n_2842));
OAI21X1 g63271(.A0 (n_2840), .A1 (g2020), .B0 (n_2534), .Y (n_2841));
OAI21X1 g63273(.A0 (n_2840), .A1 (g2013), .B0 (n_2533), .Y (n_2839));
OAI21X1 g63276(.A0 (n_2840), .A1 (g2033), .B0 (n_2532), .Y (n_2838));
OAI21X1 g63278(.A0 (n_2840), .A1 (g2026), .B0 (n_2524), .Y (n_2837));
OAI21X1 g63281(.A0 (n_2840), .A1 (g2052), .B0 (n_2531), .Y (n_2836));
OAI21X1 g63284(.A0 (n_2840), .A1 (n_2834), .B0 (n_2530), .Y (n_2835));
OAI21X1 g63287(.A0 (n_2840), .A1 (g2066), .B0 (n_2529), .Y (n_2833));
OAI21X1 g63293(.A0 (n_2840), .A1 (g2040), .B0 (n_2527), .Y (n_2832));
OAI21X1 g63296(.A0 (n_2840), .A1 (g2072), .B0 (n_2528), .Y (n_2831));
OAI21X1 g63323(.A0 (n_2840), .A1 (g2046), .B0 (n_2668), .Y (n_2830));
NAND3X1 g63533(.A (n_2655), .B (n_2656), .C (n_2658), .Y (n_2829));
NAND3X1 g63548(.A (n_4287), .B (n_2788), .C (n_4289), .Y (n_2828));
NAND2X1 g63773(.A (n_2416), .B (g6518), .Y (n_4538));
NAND2X1 g63784(.A (n_2416), .B (g6368), .Y (n_4540));
AOI21X1 g65016(.A0 (n_1511), .A1 (n_2925), .B0 (n_2497), .Y (n_2929));
NAND2X1 g63825(.A (g_22408), .B (g6313), .Y (n_5585));
CLKBUFX1 gbuf_d_994(.A(n_2444), .Y(d_out_994));
CLKBUFX1 gbuf_q_994(.A(q_in_994), .Y(g2118));
NOR2X1 g66335(.A (g1261), .B (n_2499), .Y (n_2826));
OAI21X1 g65784(.A0 (g2658), .A1 (n_2587), .B0 (n_1718), .Y (n_2986));
OR2X1 g64227(.A (n_2823), .B (n_3112), .Y (n_2824));
NOR2X1 g64228(.A (n_2821), .B (n_3542), .Y (n_2822));
NAND2X1 g64230(.A (n_4066), .B (n_2650), .Y (n_2820));
NAND2X1 g64243(.A (n_2409), .B (n_2624), .Y (n_2819));
NAND2X1 g64291(.A (n_2633), .B (n_2648), .Y (n_2818));
NAND2X1 g64339(.A (n_2816), .B (n_3540), .Y (n_2817));
OR2X1 g66287(.A (g728), .B (n_2814), .Y (n_2815));
OAI21X1 g61803(.A0 (n_2381), .A1 (n_4963), .B0 (n_2340), .Y (n_2813));
OAI21X1 g64481(.A0 (n_2811), .A1 (n_2664), .B0 (n_2517), .Y (n_2812));
MX2X1 g64489(.A (n_2809), .B (g2249), .S0 (n_2943), .Y (n_2810));
MX2X1 g64492(.A (n_4368), .B (g2252), .S0 (n_2943), .Y (n_2808));
CLKBUFX1 gbuf_d_995(.A(n_2518), .Y(d_out_995));
CLKBUFX1 gbuf_q_995(.A(q_in_995), .Y(g739));
INVX1 g64744(.A (n_2805), .Y (n_2942));
AOI21X1 g64796(.A0 (n_1628), .A1 (n_2020), .B0 (n_2466), .Y (n_2941));
AOI21X1 g64799(.A0 (n_1615), .A1 (n_2797), .B0 (n_2469), .Y (n_2940));
AOI21X1 g64812(.A0 (n_1711), .A1 (n_2797), .B0 (n_2465), .Y (n_3108));
INVX1 g64813(.A (n_4689), .Y (n_2795));
INVX1 g64816(.A (n_4687), .Y (n_2794));
INVX1 g64830(.A (n_2790), .Y (n_3110));
INVX1 g64839(.A (n_2788), .Y (n_2938));
INVX1 g64885(.A (n_2785), .Y (n_3288));
INVX8 g66746(.A (n_2780), .Y (n_4162));
INVX1 g64993(.A (n_2779), .Y (n_3279));
AOI22X1 g65275(.A0 (n_2015), .A1 (n_3093), .B0 (g1306), .B1 (n_5270),.Y (n_7271));
AOI22X1 g65291(.A0 (n_2017), .A1 (n_3093), .B0 (n_5270), .B1 (g1297),.Y (n_7273));
NAND3X1 g65415(.A (n_2061), .B (n_754), .C (n_2374), .Y (n_2776));
INVX1 g66684(.A (n_2748), .Y (n_4601));
NAND2X1 g65450(.A (n_2489), .B (n_3498), .Y (n_2774));
NAND2X1 g65457(.A (n_2477), .B (n_5035), .Y (n_2773));
NAND2X1 g65464(.A (n_2490), .B (n_3264), .Y (n_2772));
NAND3X1 g65485(.A (n_2769), .B (n_818), .C (n_2376), .Y (n_9669));
NAND2X1 g65487(.A (n_2475), .B (n_2769), .Y (n_2770));
NAND2X1 g65498(.A (n_2484), .B (n_2769), .Y (n_2768));
NAND2X1 g65508(.A (n_2473), .B (n_5035), .Y (n_2767));
NAND3X1 g65509(.A (n_2046), .B (n_839), .C (n_2377), .Y (n_2765));
NAND3X1 g65513(.A (n_3816), .B (n_1059), .C (n_2375), .Y (n_2764));
NAND2X1 g65524(.A (n_2472), .B (n_3810), .Y (n_2763));
OAI21X1 g62289(.A0 (n_2478), .A1 (g1316), .B0 (n_2479), .Y (n_2762));
NOR2X1 g65839(.A (n_951), .B (n_2458), .Y (n_2761));
INVX1 g65883(.A (n_2760), .Y (n_3082));
NAND2X1 g65887(.A (n_2758), .B (g640), .Y (n_3079));
NOR2X1 g65894(.A (n_2758), .B (g640), .Y (n_2759));
INVX1 g65947(.A (n_2757), .Y (n_3080));
AND2X1 g65951(.A (n_2755), .B (g2714), .Y (n_2905));
NOR2X1 g65953(.A (n_2755), .B (g2714), .Y (n_2756));
NAND2X1 g62404(.A (n_2753), .B (g1423), .Y (n_2754));
AOI22X1 g66076(.A0 (n_2354), .A1 (g2502), .B0 (g2503), .B1 (n_9512),.Y (n_2752));
AOI22X1 g66095(.A0 (n_2353), .A1 (g1808), .B0 (g1809), .B1 (n_1235),.Y (n_2751));
NOR2X1 g66440(.A (n_2748), .B (n_84), .Y (n_2750));
NOR2X1 g66248(.A (g578), .B (n_2748), .Y (n_2749));
NAND2X1 g66267(.A (g2039), .B (n_2292), .Y (n_2747));
OR2X1 g66403(.A (g584), .B (n_2748), .Y (n_2746));
NOR2X1 g66415(.A (g1264), .B (n_2499), .Y (n_2745));
NOR2X1 g66417(.A (g1270), .B (n_3220), .Y (n_2744));
NAND2X1 g66444(.A (g1345), .B (n_2410), .Y (n_2743));
AOI21X1 g66527(.A0 (g411), .A1 (g6447), .B0 (g408), .Y (n_2742));
AOI21X1 g66558(.A0 (g441), .A1 (g6447), .B0 (g438), .Y (n_2741));
AOI21X1 g66563(.A0 (g432), .A1 (g6447), .B0 (g429), .Y (n_2739));
AOI22X1 g66564(.A0 (n_1241), .A1 (g2448), .B0 (g2459), .B1 (n_2736),.Y (n_2738));
CLKBUFX1 gbuf_d_996(.A(n_2496), .Y(d_out_996));
CLKBUFX1 gbuf_q_996(.A(q_in_996), .Y(g2813));
AOI22X1 g66577(.A0 (n_1240), .A1 (g2433), .B0 (g2444), .B1 (n_2736),.Y (n_2737));
MX2X1 g62600(.A (g2219), .B (n_436), .S0 (n_4532), .Y (n_2735));
MX2X1 g62605(.A (g2218), .B (n_436), .S0 (n_4530), .Y (n_2733));
AOI22X1 g66603(.A0 (n_1236), .A1 (g1739), .B0 (g1750), .B1 (n_3036),.Y (n_2732));
CLKBUFX1 gbuf_d_997(.A(g7084), .Y(d_out_997));
CLKBUFX1 gbuf_q_997(.A(q_in_997), .Y(g2241));
INVX2 g66822(.A (g1930), .Y (n_6626));
MX2X1 g62662(.A (g2206), .B (n_4368), .S0 (n_4530), .Y (n_2724));
MX2X1 g62664(.A (g2207), .B (n_4368), .S0 (n_4532), .Y (n_2723));
MX2X1 g62665(.A (g2210), .B (n_2809), .S0 (n_4532), .Y (n_2722));
MX2X1 g62668(.A (g2221), .B (n_2719), .S0 (n_4530), .Y (n_2720));
MX2X1 g62669(.A (g2222), .B (n_2719), .S0 (n_4532), .Y (n_2718));
MX2X1 g62670(.A (g2224), .B (n_2716), .S0 (n_4530), .Y (n_2717));
MX2X1 g62671(.A (g2225), .B (n_2716), .S0 (n_4532), .Y (n_2715));
MX2X1 g62672(.A (g2227), .B (n_385), .S0 (n_4530), .Y (n_2714));
MX2X1 g62673(.A (g2228), .B (n_385), .S0 (n_4532), .Y (n_2712));
MX2X1 g62676(.A (g2231), .B (n_447), .S0 (n_4532), .Y (n_2711));
MX2X1 g62677(.A (g2233), .B (n_2706), .S0 (n_4530), .Y (n_2710));
OR2X1 g67110(.A (g2524), .B (n_2736), .Y (n_2709));
MX2X1 g62678(.A (g2234), .B (n_2706), .S0 (n_4532), .Y (n_2707));
NAND2X1 g67117(.A (g1119), .B (n_2343), .Y (n_2705));
OR2X1 g67128(.A (g343), .B (n_2874), .Y (n_2704));
MX2X1 g62681(.A (g2209), .B (n_2809), .S0 (n_4530), .Y (n_2703));
CLKBUFX1 gbuf_d_998(.A(n_2495), .Y(d_out_998));
CLKBUFX1 gbuf_q_998(.A(q_in_998), .Y(g2119));
MX2X1 g62686(.A (g2230), .B (n_447), .S0 (n_4530), .Y (n_2702));
NAND2X1 g67170(.A (g1615), .B (n_2433), .Y (n_9613));
NAND2X1 g67173(.A (g1624), .B (n_2433), .Y (n_9574));
NAND2X1 g67183(.A (g1651), .B (n_2433), .Y (n_8220));
NAND2X1 g67199(.A (g1579), .B (n_2433), .Y (n_9649));
CLKBUFX1 gbuf_d_999(.A(n_2494), .Y(d_out_999));
CLKBUFX1 gbuf_q_999(.A(q_in_999), .Y(g738));
MX2X1 g62755(.A (g105), .B (g_5844), .S0 (n_5587), .Y (n_2693));
MX2X1 g62759(.A (n_5247), .B (g_29016), .S0 (n_5587), .Y (n_2692));
MX2X1 g62766(.A (n_3161), .B (g_7184), .S0 (n_5587), .Y (n_2691));
MX2X1 g62796(.A (n_5382), .B (g_20789), .S0 (n_5587), .Y (n_2690));
MX2X1 g62797(.A (n_3187), .B (g_24187), .S0 (n_5587), .Y (n_2689));
MX2X1 g62800(.A (n_5380), .B (g_26130), .S0 (n_5587), .Y (n_2688));
NAND2X1 g67025(.A (g1606), .B (n_2433), .Y (n_2687));
NAND2X1 g62948(.A (n_2685), .B (g2117), .Y (n_2686));
NAND2X1 g63054(.A (n_4971), .B (g1513), .Y (n_2684));
NAND2X1 g63058(.A (n_4973), .B (g1530), .Y (n_2683));
NAND2X1 g63059(.A (n_4971), .B (g1531), .Y (n_2682));
NAND2X1 g63060(.A (n_4971), .B (g1534), .Y (n_2681));
NAND2X1 g63062(.A (n_4973), .B (g1536), .Y (n_2680));
NAND2X1 g63064(.A (n_4971), .B (g1537), .Y (n_2679));
NAND2X1 g63070(.A (n_4973), .B (g1539), .Y (n_2678));
NAND2X1 g63071(.A (n_4971), .B (g1540), .Y (n_2677));
OR2X1 g63087(.A (n_2814), .B (n_1678), .Y (n_3064));
NAND2X1 g63158(.A (n_4973), .B (g1533), .Y (n_2676));
NAND2X1 g63198(.A (n_4973), .B (g1512), .Y (n_2675));
OR2X1 g63501(.A (n_1531), .B (n_2674), .Y (n_3010));
OR2X1 g66352(.A (g2802), .B (n_2674), .Y (n_2672));
NAND2X1 g66954(.A (g1003), .B (n_2343), .Y (n_2670));
NAND2X1 g63754(.A (n_2840), .B (g2096), .Y (n_2668));
AND2X1 g63810(.A (n_6451), .B (n_6914), .Y (n_2667));
AND2X1 g65948(.A (n_2606), .B (g1326), .Y (n_2757));
CLKBUFX1 gbuf_d_1000(.A(g7194), .Y(d_out_1000));
CLKBUFX1 gbuf_qn_1000(.A(qn_in_1000), .Y(g1930));
NAND2X1 g64439(.A (n_1530), .B (n_2451), .Y (n_3151));
MX2X1 g64536(.A (n_4110), .B (g861), .S0 (n_2664), .Y (n_2665));
MX2X1 g64539(.A (n_4112), .B (g864), .S0 (n_2664), .Y (n_2663));
MX2X1 g64542(.A (n_4464), .B (g867), .S0 (n_2664), .Y (n_2662));
NAND2X1 g67148(.A (g2318), .B (n_7811), .Y (n_8246));
NAND2X1 g64627(.A (n_2943), .B (g2246), .Y (n_2660));
NAND2X1 g64632(.A (n_2943), .B (g2255), .Y (n_2659));
INVX1 g64740(.A (n_2658), .Y (n_3286));
AOI21X1 g64745(.A0 (n_1717), .A1 (n_2653), .B0 (n_2373), .Y (n_2805));
INVX1 g64748(.A (n_2657), .Y (n_2803));
INVX1 g64750(.A (n_3136), .Y (n_3129));
INVX1 g64754(.A (n_2656), .Y (n_3284));
INVX1 g64762(.A (n_2655), .Y (n_3277));
INVX1 g64764(.A (n_3281), .Y (n_2654));
AOI21X1 g64766(.A0 (n_1715), .A1 (n_2653), .B0 (n_2372), .Y (n_2956));
INVX1 g64768(.A (n_2816), .Y (n_2652));
INVX1 g64780(.A (n_2651), .Y (n_2799));
INVX1 g64791(.A (n_2650), .Y (n_4064));
OAI21X1 g64793(.A0 (n_2814), .A1 (g737), .B0 (n_1938), .Y (n_2649));
INVX1 g64801(.A (n_2648), .Y (n_4691));
INVX1 g64803(.A (n_4685), .Y (n_2647));
INVX1 g64805(.A (n_2645), .Y (n_2646));
OAI21X1 g64814(.A0 (g710), .A1 (g629), .B0 (n_2021), .Y (n_4689));
OAI21X1 g64817(.A0 (g707), .A1 (n_2814), .B0 (n_2022), .Y (n_4687));
INVX1 g64819(.A (n_3112), .Y (n_2639));
INVX1 g64822(.A (n_2638), .Y (n_4683));
INVX1 g64828(.A (n_4289), .Y (n_2636));
AOI21X1 g64832(.A0 (n_1629), .A1 (n_2635), .B0 (n_2368), .Y (n_2790));
AOI21X1 g64840(.A0 (n_1435), .A1 (n_2635), .B0 (n_2369), .Y (n_2788));
INVX1 g64842(.A (n_2634), .Y (n_4283));
INVX1 g64855(.A (n_2633), .Y (n_2786));
INVX1 g64857(.A (n_3542), .Y (n_2632));
INVX1 g64882(.A (n_4066), .Y (n_2631));
AOI21X1 g64886(.A0 (n_1705), .A1 (n_2653), .B0 (n_2338), .Y (n_2785));
INVX1 g64889(.A (n_2993), .Y (n_2629));
INVX1 g64903(.A (n_3540), .Y (n_2627));
INVX1 g64923(.A (n_2626), .Y (n_2784));
INVX1 g64934(.A (n_2625), .Y (n_2783));
INVX1 g64965(.A (n_2624), .Y (n_3544));
INVX1 g64983(.A (n_2990), .Y (n_2623));
AOI21X1 g64994(.A0 (n_1707), .A1 (n_2653), .B0 (n_2370), .Y (n_2779));
INVX1 g65028(.A (n_3311), .Y (n_2621));
INVX1 g67729(.A (n_2736), .Y (g7264));
NAND3X1 g65484(.A (n_2503), .B (n_943), .C (n_2268), .Y (n_2619));
NAND2X1 g65516(.A (n_2406), .B (n_3093), .Y (n_2618));
NAND3X1 g65518(.A (n_4412), .B (n_831), .C (n_2276), .Y (n_2617));
OAI21X1 g65618(.A0 (g2811), .A1 (n_2419), .B0 (n_1719), .Y (n_2615));
AOI21X1 g65651(.A0 (n_1429), .A1 (n_2635), .B0 (n_2413), .Y (n_2614));
OAI21X1 g65732(.A0 (g2652), .A1 (n_2587), .B0 (n_1517), .Y (n_4078));
OAI21X1 g65843(.A0 (n_2238), .A1 (g240), .B0 (n_934), .Y (n_2613));
NOR2X1 g65875(.A (n_2611), .B (g2020), .Y (n_2612));
AND2X1 g65884(.A (n_2611), .B (g2020), .Y (n_2760));
AOI21X1 g65917(.A0 (n_301), .A1 (n_8305), .B0 (n_2357), .Y (n_2610));
NOR2X1 g65921(.A (n_910), .B (n_2358), .Y (n_2609));
NOR2X1 g65934(.A (n_978), .B (n_2365), .Y (n_2608));
NOR2X1 g65955(.A (n_2606), .B (g1326), .Y (n_2607));
AOI22X1 g65976(.A0 (n_2259), .A1 (g2254), .B0 (g2255), .B1 (n_1305),.Y (n_2605));
AOI21X1 g65978(.A0 (n_2257), .A1 (g_12763), .B0 (n_751), .Y (n_2604));
AOI22X1 g65979(.A0 (n_2318), .A1 (g845), .B0 (g846), .B1 (n_2597), .Y(n_2603));
AOI21X1 g65981(.A0 (n_2215), .A1 (g1696), .B0 (n_729), .Y (n_2602));
AOI22X1 g65996(.A0 (n_2237), .A1 (g403), .B0 (g404), .B1 (n_753), .Y(n_2601));
AOI22X1 g66003(.A0 (n_2256), .A1 (g857), .B0 (g858), .B1 (n_1032), .Y(n_2600));
AOI22X1 g66007(.A0 (n_2320), .A1 (g1135), .B0 (g1136), .B1 (n_8305),.Y (n_2599));
AOI22X1 g66029(.A0 (n_2258), .A1 (g851), .B0 (g852), .B1 (n_2597), .Y(n_2598));
AOI22X1 g66072(.A0 (n_2228), .A1 (g842), .B0 (g843), .B1 (n_2597), .Y(n_2595));
AOI22X1 g66073(.A0 (n_2252), .A1 (g830), .B0 (g831), .B1 (n_2597), .Y(n_2594));
OR2X1 g67072(.A (g1724), .B (n_3036), .Y (n_2593));
AOI22X1 g66077(.A0 (n_2235), .A1 (g322), .B0 (g_8008), .B1 (n_753),.Y (n_2591));
AOI22X1 g66097(.A0 (n_2245), .A1 (g1560), .B0 (g1561), .B1 (n_853),.Y (n_2589));
NAND2X1 g66228(.A (g1316), .B (n_2450), .Y (n_3305));
NOR2X1 g66234(.A (n_2587), .B (n_91), .Y (n_2588));
NAND2X1 g66427(.A (g2010), .B (g2009), .Y (n_3691));
NOR2X1 g66460(.A (n_36), .B (n_2587), .Y (n_2586));
NOR2X1 g66465(.A (g2655), .B (n_2587), .Y (n_2585));
AOI21X1 g66499(.A0 (g2507), .A1 (n_2180), .B0 (g2504), .Y (n_2584));
AOI21X1 g66510(.A0 (g1813), .A1 (g7014), .B0 (g1810), .Y (n_2583));
AOI21X1 g66539(.A0 (g1792), .A1 (g7014), .B0 (g1789), .Y (n_2582));
AOI21X1 g66584(.A0 (g2486), .A1 (n_2180), .B0 (g2483), .Y (n_2581));
AOI21X1 g66609(.A0 (g2516), .A1 (n_2180), .B0 (g2513), .Y (n_2578));
AOI21X1 g66611(.A0 (g1822), .A1 (g7014), .B0 (g1819), .Y (n_2576));
INVX1 g66893(.A (n_2863), .Y (n_3448));
INVX1 g67063(.A (n_2470), .Y (n_2572));
OR2X1 g67080(.A (g2418), .B (n_2736), .Y (n_2571));
OR2X1 g67087(.A (g_26381), .B (n_9398), .Y (n_2570));
INVX1 g67114(.A (n_2437), .Y (n_2569));
INVX1 g67137(.A (n_2516), .Y (n_2568));
NAND2X1 g67143(.A (g2273), .B (n_7811), .Y (n_9601));
NAND2X1 g67144(.A (g2300), .B (n_7811), .Y (n_2566));
NAND2X1 g67175(.A (g2309), .B (n_7811), .Y (n_2563));
NAND2X1 g67221(.A (g2345), .B (n_7811), .Y (n_8276));
AND2X1 g63804(.A (n_5885), .B (g5555), .Y (n_2561));
INVX1 g67340(.A (n_2378), .Y (n_5044));
INVX1 g67767(.A (g6313), .Y (n_3195));
NAND2X1 g62972(.A (n_2889), .B (g1384), .Y (n_2551));
NAND2X1 g62976(.A (n_2889), .B (g1387), .Y (n_2550));
NAND2X1 g62979(.A (n_2889), .B (g1390), .Y (n_2549));
NAND2X1 g62984(.A (n_2889), .B (g1393), .Y (n_2548));
NAND2X1 g62987(.A (n_2889), .B (g1396), .Y (n_2547));
NAND2X1 g62992(.A (n_2889), .B (g1399), .Y (n_2546));
NAND2X1 g62996(.A (n_2889), .B (g1402), .Y (n_2545));
NAND2X1 g62999(.A (n_2889), .B (g1405), .Y (n_2544));
NAND2X1 g63002(.A (n_2889), .B (g1408), .Y (n_2543));
NAND2X1 g63006(.A (n_2889), .B (g1411), .Y (n_2542));
NAND2X1 g63011(.A (n_2889), .B (n_2540), .Y (n_2541));
NOR2X1 g61293(.A (n_1386), .B (n_2337), .Y (n_2539));
NAND2X1 g63055(.A (n_5587), .B (g_15404), .Y (n_2538));
NAND2X1 g63141(.A (n_5587), .B (g_27738), .Y (n_2537));
NAND2X1 g63155(.A (n_5587), .B (g_14751), .Y (n_2536));
NAND2X1 g63165(.A (n_5587), .B (g_29207), .Y (n_2535));
NAND2X1 g63584(.A (n_2840), .B (g2078), .Y (n_2534));
NAND2X1 g63586(.A (n_2840), .B (g2081), .Y (n_2533));
NAND2X1 g63589(.A (n_2840), .B (g2084), .Y (n_2532));
NAND2X1 g63591(.A (n_2840), .B (g2093), .Y (n_2531));
NAND2X1 g63593(.A (n_2840), .B (g2099), .Y (n_2530));
NAND2X1 g63596(.A (n_2840), .B (g2102), .Y (n_2529));
NAND2X1 g63597(.A (n_2840), .B (g2105), .Y (n_2528));
NAND2X1 g63626(.A (n_2840), .B (g2090), .Y (n_2527));
NAND2X1 g63672(.A (n_2840), .B (n_2525), .Y (n_2526));
NAND2X1 g63679(.A (n_2840), .B (g2087), .Y (n_2524));
NAND2X1 g63686(.A (n_1566), .B (n_2264), .Y (n_3307));
OR2X1 g63776(.A (n_4055), .B (n_1285), .Y (n_4973));
OR2X1 g63789(.A (n_4055), .B (n_2194), .Y (n_4971));
INVX1 g66894(.A (n_2587), .Y (n_2863));
INVX1 g67810(.A (n_7811), .Y (n_2520));
OAI21X1 g61808(.A0 (n_2163), .A1 (n_5372), .B0 (n_2051), .Y (n_2518));
INVX1 g67768(.A (n_9398), .Y (g6313));
NAND2X1 g64624(.A (n_2664), .B (g858), .Y (n_2517));
NOR2X1 g67138(.A (g_20947), .B (n_2446), .Y (n_2516));
AOI21X1 g64741(.A0 (n_1516), .A1 (n_2653), .B0 (n_2286), .Y (n_2658));
OAI21X1 g64749(.A0 (g2799), .A1 (n_2419), .B0 (n_2025), .Y (n_2657));
OAI21X1 g64751(.A0 (g2796), .A1 (n_2419), .B0 (n_2023), .Y (n_3136));
AOI21X1 g64755(.A0 (n_1462), .A1 (n_2653), .B0 (n_2315), .Y (n_2656));
AOI21X1 g64763(.A0 (n_1515), .A1 (n_2653), .B0 (n_2298), .Y (n_2655));
OAI21X1 g64765(.A0 (g2778), .A1 (n_2419), .B0 (n_2024), .Y (n_3281));
NAND2X1 g64770(.A (n_2280), .B (n_1932), .Y (n_2816));
AOI21X1 g64781(.A0 (n_1622), .A1 (n_2508), .B0 (n_2283), .Y (n_2651));
AOI21X1 g64792(.A0 (n_1616), .A1 (n_2508), .B0 (n_2287), .Y (n_2650));
AOI21X1 g64802(.A0 (n_1514), .A1 (n_9211), .B0 (n_2297), .Y (n_2648));
NAND2X2 g64804(.A (n_9583), .B (n_9584), .Y (n_4685));
AOI21X1 g64808(.A0 (n_1513), .A1 (n_9211), .B0 (n_2296), .Y (n_2645));
INVX1 g64810(.A (n_3313), .Y (n_2641));
NAND2X1 g64820(.A (n_2295), .B (n_1642), .Y (n_3112));
AOI21X1 g64823(.A0 (n_2020), .A1 (n_9590), .B0 (n_2294), .Y (n_2638));
INVX1 g64826(.A (n_2512), .Y (n_2637));
NAND2X1 g64829(.A (n_2334), .B (n_1641), .Y (n_4289));
OAI21X1 g64833(.A0 (g1405), .A1 (n_2410), .B0 (n_1638), .Y (n_3114));
INVX1 g64834(.A (n_4287), .Y (n_2511));
AOI21X1 g64843(.A0 (n_1437), .A1 (n_8623), .B0 (n_2279), .Y (n_2634));
AOI21X1 g64852(.A0 (n_1436), .A1 (n_2635), .B0 (n_2291), .Y (n_2823));
AOI21X1 g64856(.A0 (n_1627), .A1 (n_9211), .B0 (n_2289), .Y (n_2633));
NAND2X1 g64858(.A (n_2288), .B (n_2019), .Y (n_3542));
NAND2X1 g64883(.A (n_2284), .B (n_1933), .Y (n_4066));
OAI21X1 g64891(.A0 (g1402), .A1 (n_2410), .B0 (n_1935), .Y (n_2993));
INVX1 g64901(.A (n_4285), .Y (n_2509));
NAND2X1 g64904(.A (n_9609), .B (n_9610), .Y (n_3540));
CLKBUFX1 gbuf_d_1001(.A(g6518), .Y(d_out_1001));
CLKBUFX1 gbuf_q_1001(.A(q_in_1001), .Y(n_2780));
NAND2X1 g64924(.A (n_2293), .B (n_1934), .Y (n_2626));
OAI21X1 g64935(.A0 (g2090), .A1 (n_2292), .B0 (n_1930), .Y (n_2625));
AOI21X1 g64966(.A0 (n_1611), .A1 (n_2508), .B0 (n_2290), .Y (n_2624));
NAND2X1 g64985(.A (n_2282), .B (n_1929), .Y (n_2990));
AOI21X1 g64987(.A0 (n_1612), .A1 (n_2508), .B0 (n_2281), .Y (n_2821));
NAND3X1 g65448(.A (n_8945), .B (n_842), .C (n_2200), .Y (n_2507));
AOI21X1 g66035(.A0 (g1947), .A1 (n_864), .B0 (n_2261), .Y (n_2506));
NAND3X1 g65486(.A (n_8948), .B (n_844), .C (n_2134), .Y (n_2505));
NAND3X1 g65493(.A (n_2503), .B (n_807), .C (n_2156), .Y (n_2504));
NAND3X1 g65494(.A (n_3799), .B (n_812), .C (n_2130), .Y (n_2502));
NOR2X1 g65512(.A (n_2915), .B (n_2433), .Y (n_2948));
NAND2X1 g65522(.A (n_2299), .B (n_3810), .Y (n_2501));
INVX1 g66674(.A (n_5270), .Y (n_3220));
INVX1 g66666(.A (n_5270), .Y (n_2499));
NOR2X1 g66462(.A (g2649), .B (n_2587), .Y (n_2497));
OAI21X1 g62287(.A0 (n_2058), .A1 (n_5181), .B0 (n_1772), .Y (n_2496));
OAI21X1 g62291(.A0 (n_2055), .A1 (n_4967), .B0 (n_2043), .Y (n_2495));
OAI21X1 g62292(.A0 (n_2300), .A1 (g630), .B0 (n_2301), .Y (n_2494));
OR2X1 g65841(.A (n_956), .B (n_2273), .Y (n_2493));
AOI21X1 g65849(.A0 (n_2103), .A1 (n_94), .B0 (n_727), .Y (n_2492));
AOI21X1 g65867(.A0 (n_2090), .A1 (n_97), .B0 (n_750), .Y (n_9685));
AOI21X1 g65870(.A0 (n_174), .A1 (n_864), .B0 (n_2277), .Y (n_2490));
AOI21X1 g65880(.A0 (n_147), .A1 (n_2170), .B0 (n_2272), .Y (n_2489));
AOI21X1 g65881(.A0 (n_298), .A1 (n_2170), .B0 (n_2270), .Y (n_2488));
AOI21X1 g65915(.A0 (n_59), .A1 (n_864), .B0 (n_2275), .Y (n_2486));
AOI22X1 g66008(.A0 (n_2065), .A1 (g839), .B0 (g840), .B1 (n_2597), .Y(n_2485));
AOI21X1 g66011(.A0 (n_2074), .A1 (g2478), .B0 (n_852), .Y (n_2484));
AOI22X1 g66013(.A0 (n_2093), .A1 (g1114), .B0 (g1115), .B1 (n_8305),.Y (n_2483));
AOI22X1 g66015(.A0 (n_2080), .A1 (g866), .B0 (g867), .B1 (n_1032), .Y(n_2482));
OAI21X1 g66016(.A0 (n_2099), .A1 (n_276), .B0 (n_756), .Y (n_2480));
NAND2X1 g62405(.A (n_2478), .B (g1424), .Y (n_2479));
AOI21X1 g66046(.A0 (n_2110), .A1 (g1703), .B0 (n_856), .Y (n_2477));
OAI21X1 g66055(.A0 (n_2073), .A1 (n_129), .B0 (n_792), .Y (n_2476));
AOI21X1 g66057(.A0 (n_2096), .A1 (g2397), .B0 (n_904), .Y (n_2475));
OAI21X1 g66063(.A0 (n_2179), .A1 (n_149), .B0 (n_798), .Y (n_2474));
AOI21X1 g66064(.A0 (n_2095), .A1 (g1784), .B0 (n_821), .Y (n_2473));
AOI22X1 g66088(.A0 (n_2084), .A1 (g1041), .B0 (g1030), .B1 (n_8305),.Y (n_2472));
NOR2X1 g67064(.A (g_14855), .B (n_9398), .Y (n_2470));
NOR2X1 g66207(.A (n_2814), .B (g659), .Y (n_2758));
NOR2X1 g66227(.A (g698), .B (n_2814), .Y (n_2469));
OR2X1 g66238(.A (g1414), .B (n_2410), .Y (n_2468));
NOR2X1 g66268(.A (g719), .B (n_2814), .Y (n_2466));
NOR2X1 g66279(.A (g731), .B (n_2814), .Y (n_2465));
OR2X1 g66318(.A (g2108), .B (n_2292), .Y (n_2463));
NOR2X1 g66455(.A (g2733), .B (n_2419), .Y (n_2755));
AOI21X1 g66519(.A0 (g420), .A1 (g6447), .B0 (g417), .Y (n_2458));
NAND2X1 g66525(.A (n_2218), .B (n_220), .Y (n_2457));
NAND2X1 g66541(.A (n_2243), .B (n_237), .Y (n_2456));
NAND2X1 g66550(.A (n_2210), .B (n_326), .Y (n_9647));
OAI21X1 g66572(.A0 (n_909), .A1 (n_228), .B0 (n_2233), .Y (n_2454));
CLKBUFX1 gbuf_d_1002(.A(n_2278), .Y(d_out_1002));
CLKBUFX1 gbuf_q_1002(.A(q_in_1002), .Y(g2812));
INVX1 g66687(.A (g550), .Y (n_2748));
INVX1 g66900(.A (n_2451), .Y (n_2674));
NAND2X1 g66966(.A (g912), .B (n_8339), .Y (n_2449));
OR2X1 g66969(.A (g_19132), .B (n_2446), .Y (n_8207));
NAND2X1 g66978(.A (g921), .B (n_8339), .Y (n_2445));
OAI21X1 g62661(.A0 (n_2220), .A1 (g2010), .B0 (n_2221), .Y (n_2444));
OR2X1 g67035(.A (g_23490), .B (n_2579), .Y (n_2443));
NAND2X1 g67046(.A (g885), .B (n_8339), .Y (n_2442));
OR2X1 g67079(.A (g_30039), .B (n_9398), .Y (n_2441));
OR2X1 g67100(.A (g428), .B (n_2874), .Y (n_2439));
NOR2X1 g67115(.A (g_16484), .B (n_2446), .Y (n_2437));
OR2X1 g67172(.A (g_23514), .B (n_2579), .Y (n_2436));
NAND2X1 g67229(.A (g957), .B (n_8339), .Y (n_8270));
CLKBUFX1 g67313(.A (n_2769), .Y (n_4604));
INVX1 g67809(.A (n_7811), .Y (g7084));
INVX1 g67561(.A (n_2433), .Y (n_2422));
OR2X1 g63029(.A (n_1968), .B (n_2410), .Y (n_2753));
OAI21X1 g65029(.A0 (g2781), .A1 (n_2419), .B0 (n_1721), .Y (n_3311));
OR2X1 g66968(.A (g_24593), .B (n_9398), .Y (n_2418));
CLKBUFX1 g67249(.A (n_2046), .Y (n_5035));
OR2X1 g63603(.A (n_1749), .B (n_2292), .Y (n_2685));
AND2X1 g63792(.A (g2257), .B (g6837), .Y (n_4530));
CLKBUFX1 gbuf_d_1003(.A(n_2199), .Y(d_out_1003));
CLKBUFX1 gbuf_q_1003(.A(q_in_1003), .Y(g708));
CLKBUFX1 gbuf_d_1004(.A(n_2202), .Y(d_out_1004));
CLKBUFX1 gbuf_q_1004(.A(q_in_1004), .Y(g711));
CLKBUFX1 gbuf_d_1005(.A(n_2120), .Y(d_out_1005));
CLKBUFX1 gbuf_q_1005(.A(q_in_1005), .Y(g715));
CLKBUFX1 gbuf_d_1006(.A(n_2124), .Y(d_out_1006));
CLKBUFX1 gbuf_q_1006(.A(q_in_1006), .Y(g700));
CLKBUFX1 gbuf_d_1007(.A(n_2191), .Y(d_out_1007));
CLKBUFX1 gbuf_q_1007(.A(q_in_1007), .Y(g702));
CLKBUFX1 gbuf_d_1008(.A(n_2121), .Y(d_out_1008));
CLKBUFX1 gbuf_q_1008(.A(q_in_1008), .Y(g714));
INVX1 g66916(.A (n_2410), .Y (n_2450));
INVX1 g66901(.A (n_2419), .Y (n_2451));
CLKBUFX1 gbuf_d_1009(.A(n_2122), .Y(d_out_1009));
CLKBUFX1 gbuf_q_1009(.A(q_in_1009), .Y(g709));
CLKBUFX1 gbuf_d_1010(.A(n_2208), .Y(d_out_1010));
CLKBUFX1 gbuf_q_1010(.A(q_in_1010), .Y(g712));
NOR2X1 g66295(.A (g1423), .B (n_2410), .Y (n_2413));
INVX1 g67813(.A (n_2339), .Y (n_7811));
OR2X1 g64327(.A (n_1449), .B (n_2292), .Y (n_2840));
CLKBUFX1 gbuf_d_1011(.A(n_2204), .Y(d_out_1011));
CLKBUFX1 gbuf_q_1011(.A(q_in_1011), .Y(g1409));
CLKBUFX1 gbuf_d_1012(.A(n_2135), .Y(d_out_1012));
CLKBUFX1 gbuf_q_1012(.A(q_in_1012), .Y(g1407));
CLKBUFX1 gbuf_d_1013(.A(n_2105), .Y(d_out_1013));
CLKBUFX1 gbuf_q_1013(.A(q_in_1013), .Y(g726));
CLKBUFX1 gbuf_d_1014(.A(n_2131), .Y(d_out_1014));
CLKBUFX1 gbuf_q_1014(.A(q_in_1014), .Y(g1413));
CLKBUFX1 gbuf_d_1015(.A(n_2133), .Y(d_out_1015));
CLKBUFX1 gbuf_q_1015(.A(q_in_1015), .Y(g1410));
OAI21X1 g64811(.A0 (g722), .A1 (g629), .B0 (n_1936), .Y (n_3313));
OAI21X1 g64827(.A0 (g1408), .A1 (n_2410), .B0 (n_1606), .Y (n_2512));
OAI21X1 g64835(.A0 (g1390), .A1 (n_2410), .B0 (n_1639), .Y (n_4287));
OAI21X1 g64902(.A0 (g1387), .A1 (n_2410), .B0 (n_1634), .Y (n_4285));
CLKBUFX1 gbuf_d_1016(.A(n_2132), .Y(d_out_1016));
CLKBUFX1 gbuf_q_1016(.A(q_in_1016), .Y(g1412));
CLKBUFX1 gbuf_d_1017(.A(n_2137), .Y(d_out_1017));
CLKBUFX1 gbuf_q_1017(.A(q_in_1017), .Y(g1406));
CLKBUFX1 gbuf_d_1018(.A(n_2192), .Y(d_out_1018));
CLKBUFX1 gbuf_q_1018(.A(q_in_1018), .Y(g703));
CLKBUFX1 gbuf_d_1019(.A(n_2193), .Y(d_out_1019));
CLKBUFX1 gbuf_q_1019(.A(q_in_1019), .Y(g705));
CLKBUFX1 gbuf_d_1020(.A(n_2142), .Y(d_out_1020));
CLKBUFX1 gbuf_q_1020(.A(q_in_1020), .Y(g1400));
CLKBUFX1 gbuf_d_1021(.A(g6642), .Y(d_out_1021));
CLKBUFX1 gbuf_q_1021(.A(q_in_1021), .Y(g550));
CLKBUFX1 gbuf_d_1022(.A(g6944), .Y(d_out_1022));
CLKBUFX1 gbuf_q_1022(.A(q_in_1022), .Y(n_5270));
CLKBUFX1 gbuf_d_1023(.A(n_2138), .Y(d_out_1023));
CLKBUFX1 gbuf_q_1023(.A(q_in_1023), .Y(g1404));
NAND2X1 g65527(.A (n_3793), .B (n_2339), .Y (n_2943));
OAI21X1 g65762(.A0 (g2117), .A1 (n_2292), .B0 (n_1632), .Y (n_2409));
INVX1 g67372(.A (n_2407), .Y (n_2408));
AOI21X1 g65838(.A0 (n_231), .A1 (n_2014), .B0 (n_2157), .Y (n_2406));
AOI21X1 g65842(.A0 (n_198), .A1 (n_8305), .B0 (n_2128), .Y (n_2405));
AOI21X1 g65846(.A0 (n_67), .A1 (n_8305), .B0 (n_2190), .Y (n_2404));
AOI21X1 g65854(.A0 (n_42), .A1 (n_2170), .B0 (n_2145), .Y (n_2403));
AOI22X1 g65862(.A0 (n_1967), .A1 (n_317), .B0 (n_1768), .B1 (n_8400),.Y (n_9650));
AOI22X1 g65869(.A0 (n_2005), .A1 (n_315), .B0 (n_1841), .B1 (n_8400),.Y (n_9660));
AOI22X1 g65876(.A0 (n_2034), .A1 (n_137), .B0 (n_1884), .B1 (n_2389),.Y (n_2399));
AOI21X1 g65879(.A0 (n_37), .A1 (n_8305), .B0 (n_2153), .Y (n_2398));
OAI21X1 g65902(.A0 (n_2003), .A1 (g1648), .B0 (n_835), .Y (n_2397));
OAI21X1 g65909(.A0 (n_2001), .A1 (g2342), .B0 (n_797), .Y (n_2396));
NAND2X1 g65911(.A (n_2007), .B (n_3810), .Y (n_2395));
AOI21X1 g65920(.A0 (n_108), .A1 (n_2014), .B0 (n_2147), .Y (n_2393));
OR2X1 g65927(.A (n_922), .B (n_2129), .Y (n_2391));
AOI22X1 g65935(.A0 (n_1998), .A1 (n_155), .B0 (n_1875), .B1 (n_2389),.Y (n_2390));
AOI22X1 g65937(.A0 (n_2004), .A1 (n_157), .B0 (n_1895), .B1 (n_8400),.Y (n_2388));
AOI22X1 g65943(.A0 (n_1999), .A1 (n_322), .B0 (n_1878), .B1 (n_8400),.Y (n_2386));
AOI22X1 g65969(.A0 (n_2006), .A1 (g863), .B0 (g864), .B1 (n_2389), .Y(n_2384));
AOI22X1 g65998(.A0 (n_1989), .A1 (g860), .B0 (g861), .B1 (n_8400), .Y(n_2383));
AOI21X1 g66054(.A0 (g1253), .A1 (n_2014), .B0 (n_2126), .Y (n_2382));
AOI21X1 g62433(.A0 (n_2217), .A1 (g7161), .B0 (g1425), .Y (n_2381));
AOI21X1 g66091(.A0 (g567), .A1 (n_2170), .B0 (n_2127), .Y (n_2379));
CLKBUFX1 gbuf_d_1024(.A(n_2178), .Y(d_out_1024));
CLKBUFX1 gbuf_q_1024(.A(q_in_1024), .Y(g1385));
CLKBUFX1 gbuf_d_1025(.A(n_2125), .Y(d_out_1025));
CLKBUFX1 gbuf_q_1025(.A(q_in_1025), .Y(g699));
NAND2X1 g66188(.A (n_2123), .B (g1699), .Y (n_2377));
NAND2X1 g66189(.A (n_2072), .B (g2393), .Y (n_2376));
NAND2X1 g66193(.A (n_2101), .B (g848), .Y (n_2375));
NAND2X1 g66195(.A (n_2068), .B (g_5496), .Y (n_2374));
NOR2X1 g66201(.A (g2787), .B (n_2419), .Y (n_2373));
NOR2X1 g66203(.A (g2805), .B (n_2419), .Y (n_2372));
NOR2X1 g66211(.A (g1345), .B (n_2410), .Y (n_2606));
NOR2X1 g66246(.A (g2775), .B (n_2419), .Y (n_2370));
NOR2X1 g66249(.A (g1396), .B (n_2410), .Y (n_2369));
NOR2X1 g66251(.A (g1411), .B (n_2410), .Y (n_2368));
NOR2X1 g66260(.A (g2039), .B (n_2292), .Y (n_2611));
INVX1 g67351(.A (n_9505), .Y (n_9686));
AOI21X1 g66506(.A0 (g1801), .A1 (g7014), .B0 (g1798), .Y (n_2365));
NAND2X1 g66522(.A (n_2097), .B (n_1039), .Y (n_2363));
AOI22X1 g66534(.A0 (n_955), .A1 (g1060), .B0 (g1071), .B1 (n_2361),.Y (n_2362));
AOI22X1 g66540(.A0 (n_939), .A1 (g1045), .B0 (g1056), .B1 (n_2361),.Y (n_2360));
CLKBUFX1 gbuf_d_1026(.A(n_2140), .Y(d_out_1026));
CLKBUFX1 gbuf_q_1026(.A(q_in_1026), .Y(g1403));
AOI21X1 g66574(.A0 (g2495), .A1 (n_2180), .B0 (g2492), .Y (n_2358));
CLKBUFX1 gbuf_d_1027(.A(n_2048), .Y(d_out_1027));
CLKBUFX1 gbuf_q_1027(.A(q_in_1027), .Y(g2920));
AOI21X1 g66590(.A0 (g1128), .A1 (n_1983), .B0 (g1125), .Y (n_2357));
AOI22X1 g66610(.A0 (n_1073), .A1 (g1075), .B0 (g1085), .B1 (n_2361),.Y (n_2356));
CLKBUFX1 gbuf_d_1028(.A(n_2119), .Y(d_out_1028));
CLKBUFX1 gbuf_q_1028(.A(q_in_1028), .Y(g717));
NAND2X1 g67011(.A (g930), .B (n_8339), .Y (n_2355));
OR2X1 g67185(.A (g2503), .B (n_2736), .Y (n_2354));
OR2X1 g67226(.A (g1809), .B (n_3036), .Y (n_2353));
INVX2 g67314(.A (n_9438), .Y (n_2769));
CLKBUFX1 gbuf_d_1029(.A(n_2196), .Y(d_out_1029));
CLKBUFX1 gbuf_q_1029(.A(q_in_1029), .Y(g706));
INVX2 g67347(.A (n_2921), .Y (n_2346));
CLKBUFX1 gbuf_d_1030(.A(n_2141), .Y(d_out_1030));
CLKBUFX1 gbuf_q_1030(.A(q_in_1030), .Y(g1401));
CLKBUFX1 gbuf_d_1031(.A(n_2104), .Y(d_out_1031));
CLKBUFX1 gbuf_q_1031(.A(q_in_1031), .Y(g727));
NAND2X1 g63033(.A (n_1968), .B (g1425), .Y (n_2340));
NAND2X1 g63820(.A (g_22408), .B (g6231), .Y (n_5587));
AND2X1 g63801(.A (g2257), .B (n_2339), .Y (n_4532));
NOR2X1 g66387(.A (g2793), .B (n_2419), .Y (n_2338));
CLKBUFX1 gbuf_d_1032(.A(n_2044), .Y(d_out_1032));
CLKBUFX1 gbuf_q_1032(.A(q_in_1032), .Y(g718));
CLKBUFX1 gbuf_d_1033(.A(n_2161), .Y(d_out_1033));
CLKBUFX1 gbuf_q_1033(.A(q_in_1033), .Y(g1386));
CLKBUFX1 gbuf_d_1034(.A(n_2149), .Y(d_out_1034));
CLKBUFX1 gbuf_q_1034(.A(q_in_1034), .Y(g1395));
NAND4X1 g61432(.A (n_2189), .B (n_1052), .C (n_983), .D (n_1533), .Y(n_2337));
CLKBUFX1 gbuf_d_1035(.A(n_2143), .Y(d_out_1035));
CLKBUFX1 gbuf_q_1035(.A(q_in_1035), .Y(g1398));
CLKBUFX1 gbuf_d_1036(.A(n_2148), .Y(d_out_1036));
CLKBUFX1 gbuf_q_1036(.A(q_in_1036), .Y(g1397));
CLKBUFX1 gbuf_d_1037(.A(n_2114), .Y(d_out_1037));
CLKBUFX1 gbuf_q_1037(.A(q_in_1037), .Y(g720));
OR2X1 g63497(.A (n_1663), .B (n_2410), .Y (n_2889));
CLKBUFX1 gbuf_d_1038(.A(n_2154), .Y(d_out_1038));
CLKBUFX1 gbuf_q_1038(.A(q_in_1038), .Y(g1392));
CLKBUFX1 gbuf_d_1039(.A(n_2159), .Y(d_out_1039));
CLKBUFX1 gbuf_q_1039(.A(q_in_1039), .Y(g1388));
CLKBUFX1 gbuf_d_1040(.A(n_2151), .Y(d_out_1040));
CLKBUFX1 gbuf_q_1040(.A(q_in_1040), .Y(g1394));
CLKBUFX1 gbuf_d_1041(.A(n_2158), .Y(d_out_1041));
CLKBUFX1 gbuf_q_1041(.A(q_in_1041), .Y(g1389));
CLKBUFX1 gbuf_d_1042(.A(n_2111), .Y(d_out_1042));
CLKBUFX1 gbuf_q_1042(.A(q_in_1042), .Y(g723));
CLKBUFX1 gbuf_d_1043(.A(n_2155), .Y(d_out_1043));
CLKBUFX1 gbuf_q_1043(.A(q_in_1043), .Y(g1391));
CLKBUFX1 gbuf_d_1044(.A(n_2112), .Y(d_out_1044));
CLKBUFX1 gbuf_q_1044(.A(q_in_1044), .Y(g721));
CLKBUFX1 gbuf_d_1045(.A(n_2109), .Y(d_out_1045));
CLKBUFX1 gbuf_q_1045(.A(q_in_1045), .Y(g724));
OR2X1 g66340(.A (g1393), .B (n_2410), .Y (n_2334));
CLKBUFX1 gbuf_d_1046(.A(n_1978), .Y(d_out_1046));
CLKBUFX1 gbuf_q_1046(.A(q_in_1046), .Y(g2777));
CLKBUFX1 gbuf_d_1047(.A(n_1970), .Y(d_out_1047));
CLKBUFX1 gbuf_q_1047(.A(q_in_1047), .Y(g2801));
INVX1 g64117(.A (g869), .Y (n_2416));
INVX1 g64127(.A (g309), .Y (n_6451));
INVX1 g64136(.A (g2384), .Y (n_5885));
INVX1 g64141(.A (g996), .Y (n_5786));
INVX1 g64148(.A (n_6209), .Y (n_5531));
NOR2X1 g64161(.A (n_1662), .B (n_2039), .Y (n_4360));
CLKBUFX1 gbuf_d_1048(.A(n_2041), .Y(d_out_1048));
CLKBUFX1 gbuf_q_1048(.A(q_in_1048), .Y(g2917));
NOR2X1 g64282(.A (n_3863), .B (n_2039), .Y (n_3716));
CLKBUFX1 gbuf_d_1049(.A(n_1975), .Y(d_out_1049));
CLKBUFX1 gbuf_q_1049(.A(q_in_1049), .Y(g2786));
INVX1 g67345(.A (n_2061), .Y (n_2378));
INVX4 g66834(.A (n_2264), .Y (n_2814));
AOI21X1 g61798(.A0 (n_1918), .A1 (g3151), .B0 (n_296), .Y (n_2326));
CLKBUFX1 gbuf_d_1050(.A(n_1971), .Y(d_out_1050));
CLKBUFX1 gbuf_q_1050(.A(q_in_1050), .Y(g2798));
CLKBUFX1 gbuf_d_1051(.A(n_1972), .Y(d_out_1051));
CLKBUFX1 gbuf_q_1051(.A(q_in_1051), .Y(g2795));
CLKBUFX1 gbuf_d_1052(.A(n_1976), .Y(d_out_1052));
CLKBUFX1 gbuf_q_1052(.A(q_in_1052), .Y(g2783));
CLKBUFX1 gbuf_d_1053(.A(n_1973), .Y(d_out_1053));
CLKBUFX1 gbuf_q_1053(.A(q_in_1053), .Y(g2792));
CLKBUFX1 gbuf_d_1054(.A(n_1977), .Y(d_out_1054));
CLKBUFX1 gbuf_q_1054(.A(q_in_1054), .Y(g2780));
OR2X1 g67119(.A (g1543), .B (n_2194), .Y (n_2322));
INVX1 g67112(.A (n_2181), .Y (n_8241));
CLKBUFX1 gbuf_d_1055(.A(n_1980), .Y(d_out_1055));
CLKBUFX1 gbuf_q_1055(.A(q_in_1055), .Y(g2774));
OR2X1 g67106(.A (g1136), .B (n_2361), .Y (n_2320));
NAND2X1 g65469(.A (n_3793), .B (g6518), .Y (n_2664));
INVX1 g67101(.A (n_2089), .Y (n_2318));
NAND2X1 g65443(.A (n_2011), .B (n_3264), .Y (n_2316));
NOR2X1 g66453(.A (g2784), .B (n_2419), .Y (n_2315));
INVX1 g67373(.A (n_2503), .Y (n_2407));
AOI22X1 g65831(.A0 (n_1901), .A1 (n_200), .B0 (n_1900), .B1 (n_810),.Y (n_2314));
AOI21X1 g65868(.A0 (n_33), .A1 (n_2170), .B0 (n_2009), .Y (n_2313));
AOI22X1 g65890(.A0 (n_1943), .A1 (n_286), .B0 (n_1942), .B1 (n_2308),.Y (n_2312));
AOI21X1 g65901(.A0 (n_1864), .A1 (n_17), .B0 (n_759), .Y (n_2311));
AOI21X1 g65907(.A0 (n_1907), .A1 (n_86), .B0 (n_800), .Y (n_2310));
AOI22X1 g65908(.A0 (n_1894), .A1 (n_328), .B0 (n_1893), .B1 (n_2308),.Y (n_2309));
AOI22X1 g65910(.A0 (n_1957), .A1 (n_330), .B0 (n_1956), .B1 (n_2308),.Y (n_2307));
AOI22X1 g65912(.A0 (n_9382), .A1 (n_271), .B0 (n_9383), .B1 (n_810),.Y (n_2306));
AOI22X1 g65913(.A0 (n_1883), .A1 (n_283), .B0 (n_1882), .B1 (n_810),.Y (n_2304));
AOI22X1 g65965(.A0 (n_1898), .A1 (g2803), .B0 (g2804), .B1 (n_1245),.Y (n_2303));
AOI22X1 g65995(.A0 (n_1897), .A1 (g729), .B0 (g730), .B1 (n_1916), .Y(n_2302));
NAND2X1 g62408(.A (n_2300), .B (g738), .Y (n_2301));
AOI22X1 g66085(.A0 (n_1886), .A1 (g1009), .B0 (g1010), .B1 (n_8305),.Y (n_2299));
NOR2X1 g66226(.A (g2772), .B (n_2419), .Y (n_2298));
NOR2X1 g66229(.A (g713), .B (g629), .Y (n_2297));
NOR2X1 g66231(.A (g725), .B (g629), .Y (n_2296));
OR2X1 g66240(.A (g1399), .B (n_2410), .Y (n_2295));
NOR2X1 g66243(.A (g701), .B (g629), .Y (n_2294));
OR2X1 g66252(.A (g2105), .B (n_2292), .Y (n_2293));
NOR2X1 g66255(.A (g1417), .B (n_2410), .Y (n_2291));
NOR2X1 g66257(.A (g2099), .B (n_2292), .Y (n_2290));
NOR2X1 g66258(.A (g716), .B (g629), .Y (n_2289));
OR2X1 g66259(.A (g2093), .B (n_2292), .Y (n_2288));
NOR2X1 g66271(.A (g2078), .B (n_2292), .Y (n_2287));
NOR2X1 g66276(.A (g2790), .B (n_2419), .Y (n_2286));
OR2X1 g66320(.A (g704), .B (g629), .Y (n_9584));
OR2X1 g66321(.A (g2081), .B (n_2292), .Y (n_2284));
NOR2X1 g66356(.A (g2102), .B (n_2292), .Y (n_2283));
OR2X1 g66405(.A (g2096), .B (n_2292), .Y (n_2282));
NOR2X1 g66428(.A (g2111), .B (n_2292), .Y (n_2281));
OR2X1 g66447(.A (g2084), .B (n_2292), .Y (n_2280));
NOR2X1 g66485(.A (g1384), .B (n_2410), .Y (n_2279));
OAI21X1 g62570(.A0 (n_1984), .A1 (g2704), .B0 (n_1985), .Y (n_2278));
AOI21X1 g66500(.A0 (g1979), .A1 (g7194), .B0 (g1976), .Y (n_2277));
NAND2X1 g66502(.A (n_2000), .B (n_306), .Y (n_2276));
AOI21X1 g66511(.A0 (g1874), .A1 (g7194), .B0 (g1871), .Y (n_2275));
AOI21X1 g66518(.A0 (g1970), .A1 (g7194), .B0 (g1967), .Y (n_2273));
AOI21X1 g66542(.A0 (g590), .A1 (g6642), .B0 (g587), .Y (n_2272));
AOI21X1 g66551(.A0 (g599), .A1 (g6642), .B0 (g596), .Y (n_2270));
OAI21X1 g66553(.A0 (n_814), .A1 (n_332), .B0 (n_8892), .Y (n_2269));
NAND2X1 g66557(.A (n_2030), .B (n_303), .Y (n_2268));
AOI22X1 g66559(.A0 (n_1020), .A1 (g1552), .B0 (g1551), .B1 (n_2194),.Y (n_2267));
OAI21X1 g66569(.A0 (n_730), .A1 (n_189), .B0 (n_1986), .Y (n_2266));
NOR2X1 g66622(.A (n_1992), .B (g1945), .Y (n_2261));
CLKBUFX1 gbuf_d_1056(.A(g7390), .Y(d_out_1056));
CLKBUFX1 gbuf_qn_1056(.A(qn_in_1056), .Y(n_2587));
OR2X1 g66959(.A (g2255), .B (n_3770), .Y (n_2259));
INVX1 g66961(.A (n_2118), .Y (n_2258));
INVX1 g66963(.A (n_2116), .Y (n_2257));
INVX1 g66971(.A (n_2113), .Y (n_2256));
INVX1 g66993(.A (n_2108), .Y (n_9698));
INVX1 g66995(.A (n_2107), .Y (n_2254));
OR2X1 g67000(.A (n_83), .B (n_9397), .Y (n_2253));
INVX1 g67023(.A (n_2100), .Y (n_2252));
INVX1 g67056(.A (n_2164), .Y (n_2251));
OR2X1 g67066(.A (n_7), .B (n_9397), .Y (n_2250));
INVX1 g67075(.A (n_2182), .Y (n_2246));
OR2X1 g67077(.A (g1561), .B (n_2194), .Y (n_2245));
OR2X1 g67098(.A (n_971), .B (n_2232), .Y (n_2243));
INVX1 g67108(.A (n_2086), .Y (n_2242));
INVX1 g67123(.A (n_2081), .Y (n_8365));
INVX1 g67131(.A (n_2183), .Y (n_8367));
NOR2X1 g67177(.A (n_933), .B (n_9397), .Y (n_2238));
OR2X1 g67178(.A (g404), .B (n_2874), .Y (n_2237));
CLKBUFX1 gbuf_d_1057(.A(g26149), .Y(d_out_1057));
CLKBUFX1 gbuf_qn_1057(.A(qn_in_1057), .Y(g3113));
OR2X1 g67181(.A (g_8008), .B (n_2874), .Y (n_2235));
NAND2X1 g67189(.A (g_19787), .B (n_2232), .Y (n_2233));
INVX1 g67201(.A (n_2070), .Y (n_2231));
INVX1 g67233(.A (n_2042), .Y (n_2228));
CLKBUFX3 g67348(.A (n_9049), .Y (n_2921));
CLKBUFX3 g67365(.A (n_8408), .Y (n_3816));
OR2X1 g66410(.A (g2087), .B (n_2292), .Y (n_9610));
INVX2 g67771(.A (n_8756), .Y (n_2446));
INVX1 g67773(.A (n_8756), .Y (n_2579));
NAND2X1 g62949(.A (n_2220), .B (g2118), .Y (n_2221));
INVX1 g67568(.A (g6782), .Y (n_2433));
OR2X1 g67021(.A (n_917), .B (n_2232), .Y (n_2218));
NAND2X1 g63031(.A (n_2217), .B (g6979), .Y (n_2478));
CLKBUFX1 gbuf_d_1058(.A(g26149), .Y(d_out_1058));
CLKBUFX1 gbuf_q_1058(.A(q_in_1058), .Y(g3201));
INVX1 g66997(.A (n_2053), .Y (n_2215));
INVX1 g67538(.A (g6712), .Y (n_2343));
CLKBUFX1 gbuf_d_1059(.A(n_1974), .Y(d_out_1059));
CLKBUFX1 gbuf_q_1059(.A(q_in_1059), .Y(g2789));
CLKBUFX1 gbuf_d_1060(.A(g26149), .Y(d_out_1060));
CLKBUFX1 gbuf_qn_1060(.A(qn_in_1060), .Y(g3127));
CLKBUFX1 gbuf_d_1061(.A(g26149), .Y(d_out_1061));
CLKBUFX1 gbuf_qn_1061(.A(qn_in_1061), .Y(g3135));
CLKBUFX1 gbuf_d_1062(.A(n_2033), .Y(d_out_1062));
CLKBUFX1 gbuf_q_1062(.A(q_in_1062), .Y(g3028));
INVX1 g67252(.A (n_2046), .Y (n_2336));
AND2X1 g63553(.A (n_3863), .B (n_2211), .Y (n_2212));
OR2X1 g67096(.A (n_936), .B (n_2232), .Y (n_2210));
OR2X1 g67058(.A (g2207), .B (n_2205), .Y (n_9693));
OAI21X1 g62645(.A0 (g660), .A1 (n_2207), .B0 (n_1823), .Y (n_2208));
CLKBUFX1 gbuf_d_1063(.A(n_1784), .Y(d_out_1063));
CLKBUFX1 gbuf_q_1063(.A(q_in_1063), .Y(g2088));
OR2X1 g67214(.A (g2222), .B (n_2205), .Y (n_2206));
OAI21X1 g62593(.A0 (n_2203), .A1 (g1372), .B0 (n_1836), .Y (n_2204));
OAI21X1 g62644(.A0 (n_2201), .A1 (g660), .B0 (n_1829), .Y (n_2202));
NAND2X1 g66561(.A (n_1902), .B (n_202), .Y (n_2200));
OAI21X1 g62641(.A0 (n_2201), .A1 (g646), .B0 (n_1824), .Y (n_2199));
OAI21X1 g66552(.A0 (n_737), .A1 (n_308), .B0 (n_1888), .Y (n_2198));
CLKBUFX1 gbuf_d_1064(.A(g5595), .Y(d_out_1064));
CLKBUFX1 gbuf_qn_1064(.A(qn_in_1064), .Y(g869));
CLKBUFX1 gbuf_d_1065(.A(g5612), .Y(d_out_1065));
CLKBUFX1 gbuf_qn_1065(.A(qn_in_1065), .Y(n_4055));
CLKBUFX1 gbuf_d_1066(.A(g5549), .Y(d_out_1066));
CLKBUFX1 gbuf_qn_1066(.A(qn_in_1066), .Y(g309));
CLKBUFX1 gbuf_d_1067(.A(g5637), .Y(d_out_1067));
CLKBUFX1 gbuf_qn_1067(.A(qn_in_1067), .Y(g2384));
CLKBUFX1 gbuf_d_1068(.A(g5595), .Y(d_out_1068));
CLKBUFX1 gbuf_qn_1068(.A(qn_in_1068), .Y(g996));
CLKBUFX1 gbuf_d_1069(.A(g5612), .Y(d_out_1069));
CLKBUFX1 gbuf_q_1069(.A(q_in_1069), .Y(n_6209));
CLKBUFX1 gbuf_d_1070(.A(g5637), .Y(d_out_1070));
CLKBUFX1 gbuf_q_1070(.A(q_in_1070), .Y(g2257));
CLKBUFX1 gbuf_d_1071(.A(g5549), .Y(d_out_1071));
CLKBUFX1 gbuf_q_1071(.A(q_in_1071), .Y(g_22408));
CLKBUFX1 gbuf_d_1072(.A(n_1803), .Y(d_out_1072));
CLKBUFX1 gbuf_q_1072(.A(q_in_1072), .Y(g2103));
INVX1 g64162(.A (n_3421), .Y (n_2197));
OAI21X1 g62639(.A0 (g653), .A1 (n_2207), .B0 (n_1813), .Y (n_2196));
CLKBUFX1 gbuf_d_1073(.A(n_1793), .Y(d_out_1073));
CLKBUFX1 gbuf_q_1073(.A(q_in_1073), .Y(g2100));
OR2X1 g67190(.A (g1528), .B (n_2194), .Y (n_2195));
OAI21X1 g62638(.A0 (n_2201), .A1 (g653), .B0 (n_1812), .Y (n_2193));
CLKBUFX1 gbuf_d_1074(.A(n_1797), .Y(d_out_1074));
CLKBUFX1 gbuf_q_1074(.A(q_in_1074), .Y(g2085));
INVX1 g67815(.A (n_3770), .Y (n_2339));
NOR2X1 g64290(.A (n_1727), .B (n_3864), .Y (n_4094));
OAI21X1 g62636(.A0 (g633), .A1 (n_2207), .B0 (n_1825), .Y (n_2192));
OAI21X1 g62635(.A0 (n_2201), .A1 (g633), .B0 (n_1809), .Y (n_2191));
AOI21X1 g66521(.A0 (g1119), .A1 (g6712), .B0 (g1116), .Y (n_2190));
AOI22X1 g61823(.A0 (n_2188), .A1 (g3095), .B0 (n_2187), .B1 (n_2186),.Y (n_2189));
AOI21X1 g66524(.A0 (n_832), .A1 (g1006), .B0 (n_1887), .Y (n_8265));
CLKBUFX1 gbuf_d_1075(.A(n_1773), .Y(d_out_1075));
CLKBUFX1 gbuf_q_1075(.A(q_in_1075), .Y(g2800));
CLKBUFX1 gbuf_d_1076(.A(n_1776), .Y(d_out_1076));
CLKBUFX1 gbuf_q_1076(.A(q_in_1076), .Y(g2791));
CLKBUFX1 gbuf_d_1077(.A(n_1777), .Y(d_out_1077));
CLKBUFX1 gbuf_q_1077(.A(q_in_1077), .Y(g2785));
CLKBUFX1 gbuf_d_1078(.A(n_1774), .Y(d_out_1078));
CLKBUFX1 gbuf_q_1078(.A(q_in_1078), .Y(g2797));
CLKBUFX1 gbuf_d_1079(.A(n_1780), .Y(d_out_1079));
CLKBUFX1 gbuf_q_1079(.A(q_in_1079), .Y(g2776));
CLKBUFX1 gbuf_d_1080(.A(n_1778), .Y(d_out_1080));
CLKBUFX1 gbuf_q_1080(.A(q_in_1080), .Y(g2782));
NOR2X1 g67132(.A (g819), .B (n_8346), .Y (n_2183));
CLKBUFX1 gbuf_d_1081(.A(n_1775), .Y(d_out_1081));
CLKBUFX1 gbuf_q_1081(.A(q_in_1081), .Y(g2794));
CLKBUFX1 gbuf_d_1082(.A(n_1779), .Y(d_out_1082));
CLKBUFX1 gbuf_q_1082(.A(q_in_1082), .Y(g2779));
CLKBUFX1 gbuf_d_1083(.A(n_1789), .Y(d_out_1083));
CLKBUFX1 gbuf_q_1083(.A(q_in_1083), .Y(g2107));
NOR2X1 g67076(.A (n_99), .B (n_8326), .Y (n_2182));
CLKBUFX1 gbuf_d_1084(.A(n_1788), .Y(d_out_1084));
CLKBUFX1 gbuf_q_1084(.A(q_in_1084), .Y(g2091));
NOR2X1 g67113(.A (g1516), .B (n_2194), .Y (n_2181));
INVX1 g67734(.A (n_2180), .Y (n_2736));
CLKBUFX1 gbuf_d_1085(.A(n_1795), .Y(d_out_1085));
CLKBUFX1 gbuf_q_1085(.A(q_in_1085), .Y(g2095));
CLKBUFX1 gbuf_d_1086(.A(n_1781), .Y(d_out_1086));
CLKBUFX1 gbuf_q_1086(.A(q_in_1086), .Y(g2773));
CLKBUFX1 gbuf_d_1087(.A(n_1794), .Y(d_out_1087));
CLKBUFX1 gbuf_q_1087(.A(q_in_1087), .Y(g2097));
NOR2X1 g67089(.A (g313), .B (n_2115), .Y (n_2179));
CLKBUFX1 gbuf_d_1088(.A(n_1791), .Y(d_out_1088));
CLKBUFX1 gbuf_q_1088(.A(q_in_1088), .Y(g2104));
OAI21X1 g62567(.A0 (n_2203), .A1 (g1326), .B0 (n_1854), .Y (n_2178));
CLKBUFX1 gbuf_d_1089(.A(n_1801), .Y(d_out_1089));
CLKBUFX1 gbuf_q_1089(.A(q_in_1089), .Y(g2092));
CLKBUFX1 gbuf_d_1090(.A(n_1783), .Y(d_out_1090));
CLKBUFX1 gbuf_q_1090(.A(q_in_1090), .Y(g2098));
AOI21X1 g65833(.A0 (n_170), .A1 (n_6822), .B0 (n_1856), .Y (n_2177));
CLKBUFX1 gbuf_d_1091(.A(n_1782), .Y(d_out_1091));
CLKBUFX1 gbuf_q_1091(.A(q_in_1091), .Y(g2094));
OR2X1 g65852(.A (n_745), .B (n_1915), .Y (n_2176));
NAND2X1 g65877(.A (n_1913), .B (n_3498), .Y (n_2175));
AOI21X1 g65891(.A0 (n_167), .A1 (n_6822), .B0 (n_1806), .Y (n_2174));
AOI21X1 g65940(.A0 (n_294), .A1 (n_6822), .B0 (n_1910), .Y (n_2172));
AOI22X1 g65967(.A0 (n_1697), .A1 (g576), .B0 (g577), .B1 (n_2170), .Y(n_2171));
CLKBUFX1 gbuf_d_1092(.A(n_1787), .Y(d_out_1092));
CLKBUFX1 gbuf_q_1092(.A(q_in_1092), .Y(g2086));
AOI21X1 g66002(.A0 (g1949), .A1 (n_1689), .B0 (n_1040), .Y (n_2169));
AOI22X1 g66005(.A0 (n_1696), .A1 (g1415), .B0 (g1416), .B1 (n_8625),.Y (n_2168));
AOI22X1 g66038(.A0 (n_1693), .A1 (g2109), .B0 (g2110), .B1 (n_562),.Y (n_2167));
AOI21X1 g66045(.A0 (g2641), .A1 (n_6822), .B0 (n_1908), .Y (n_2166));
CLKBUFX1 gbuf_d_1093(.A(n_1790), .Y(d_out_1093));
CLKBUFX1 gbuf_q_1093(.A(q_in_1093), .Y(g2106));
NOR2X1 g67057(.A (g2210), .B (n_2205), .Y (n_2164));
AOI21X1 g62475(.A0 (n_1982), .A1 (g6911), .B0 (g739), .Y (n_2163));
OAI21X1 g62569(.A0 (g1326), .A1 (n_2160), .B0 (n_1853), .Y (n_2161));
OAI21X1 g62572(.A0 (n_2203), .A1 (g1319), .B0 (n_1852), .Y (n_2159));
OAI21X1 g62573(.A0 (g1319), .A1 (n_2160), .B0 (n_1851), .Y (n_2158));
AOI21X1 g66503(.A0 (g1285), .A1 (g6944), .B0 (g1282), .Y (n_2157));
NAND2X1 g66507(.A (n_1904), .B (n_204), .Y (n_2156));
OAI21X1 g62575(.A0 (n_2203), .A1 (g1339), .B0 (n_1850), .Y (n_2155));
OAI21X1 g62576(.A0 (g1339), .A1 (n_2160), .B0 (n_1849), .Y (n_2154));
AOI21X1 g66517(.A0 (g1098), .A1 (g6712), .B0 (g1095), .Y (n_2153));
OAI21X1 g62578(.A0 (n_2203), .A1 (g1332), .B0 (n_1848), .Y (n_2151));
OAI21X1 g66520(.A0 (n_752), .A1 (n_141), .B0 (n_1906), .Y (n_8362));
OAI21X1 g62579(.A0 (g1332), .A1 (n_2160), .B0 (n_1847), .Y (n_2149));
OAI21X1 g62581(.A0 (n_2203), .A1 (g1346), .B0 (n_1846), .Y (n_2148));
AOI21X1 g66528(.A0 (g1180), .A1 (g6944), .B0 (g1177), .Y (n_2147));
AOI21X1 g66529(.A0 (g_29095), .A1 (g6642), .B0 (g_27699), .Y(n_2145));
OAI21X1 g62582(.A0 (g1346), .A1 (n_2160), .B0 (n_1845), .Y (n_2143));
OAI21X1 g62584(.A0 (n_2203), .A1 (g1358), .B0 (n_1844), .Y (n_2142));
OAI21X1 g62585(.A0 (g1358), .A1 (n_2160), .B0 (n_1843), .Y (n_2141));
OAI21X1 g62587(.A0 (n_2203), .A1 (g1352), .B0 (n_1840), .Y (n_2140));
OAI21X1 g62588(.A0 (g1352), .A1 (n_2160), .B0 (n_1839), .Y (n_2138));
OAI21X1 g62590(.A0 (n_2203), .A1 (n_2880), .B0 (n_1838), .Y (n_2137));
AOI22X1 g66555(.A0 (n_894), .A1 (g2249), .B0 (g2248), .B1 (n_8891),.Y (n_2136));
OAI21X1 g62591(.A0 (n_2880), .A1 (n_2160), .B0 (n_1837), .Y (n_2135));
NAND2X1 g66560(.A (n_1919), .B (n_249), .Y (n_2134));
OAI21X1 g62594(.A0 (g1372), .A1 (n_2160), .B0 (n_1835), .Y (n_2133));
OAI21X1 g62596(.A0 (n_2203), .A1 (g1378), .B0 (n_1834), .Y (n_2132));
OAI21X1 g62597(.A0 (g1378), .A1 (n_2160), .B0 (n_1833), .Y (n_2131));
NAND2X1 g66579(.A (n_1868), .B (n_193), .Y (n_2130));
AOI21X1 g66583(.A0 (g1276), .A1 (g6944), .B0 (g1273), .Y (n_2129));
AOI21X1 g66585(.A0 (g1107), .A1 (g6712), .B0 (g1104), .Y (n_2128));
NOR2X1 g66625(.A (n_1924), .B (g565), .Y (n_2127));
NOR2X1 g66628(.A (n_1866), .B (g1251), .Y (n_2126));
OAI21X1 g62632(.A0 (n_2201), .A1 (g640), .B0 (n_1827), .Y (n_2125));
OAI21X1 g62633(.A0 (g640), .A1 (n_2207), .B0 (n_1826), .Y (n_2124));
INVX1 g66837(.A (g629), .Y (n_2264));
OR2X1 g67047(.A (g1700), .B (n_2052), .Y (n_2123));
OAI21X1 g62642(.A0 (g646), .A1 (n_2207), .B0 (n_1828), .Y (n_2122));
OAI21X1 g62647(.A0 (n_2201), .A1 (g672), .B0 (n_1832), .Y (n_2121));
OAI21X1 g62648(.A0 (g672), .A1 (n_2207), .B0 (n_1822), .Y (n_2120));
OAI21X1 g62650(.A0 (n_2201), .A1 (g666), .B0 (n_1808), .Y (n_2119));
NOR2X1 g66962(.A (g852), .B (n_8346), .Y (n_2118));
NOR2X1 g66964(.A (g_10841), .B (n_2115), .Y (n_2116));
OAI21X1 g62653(.A0 (n_2201), .A1 (n_3203), .B0 (n_1807), .Y (n_2114));
NOR2X1 g66972(.A (g858), .B (n_8326), .Y (n_2113));
OAI21X1 g62654(.A0 (n_3203), .A1 (n_2207), .B0 (n_1820), .Y (n_2112));
OAI21X1 g62656(.A0 (n_2201), .A1 (g686), .B0 (n_1814), .Y (n_2111));
OR2X1 g66988(.A (g1704), .B (n_2098), .Y (n_2110));
OAI21X1 g62657(.A0 (g686), .A1 (n_2207), .B0 (n_1819), .Y (n_2109));
NOR2X1 g66994(.A (n_60), .B (n_8346), .Y (n_2108));
NOR2X1 g66996(.A (g822), .B (n_8326), .Y (n_2107));
OR2X1 g66999(.A (g2234), .B (n_3770), .Y (n_2106));
OAI21X1 g62659(.A0 (n_2201), .A1 (g692), .B0 (n_1810), .Y (n_2105));
OAI21X1 g62660(.A0 (g692), .A1 (n_2207), .B0 (n_1818), .Y (n_2104));
OR2X1 g67012(.A (n_726), .B (n_2102), .Y (n_2103));
OR2X1 g67017(.A (g849), .B (n_8346), .Y (n_2101));
NOR2X1 g67024(.A (g831), .B (n_8326), .Y (n_2100));
NOR2X1 g67029(.A (g1694), .B (n_2098), .Y (n_2099));
NAND2X1 g67037(.A (g2245), .B (n_3770), .Y (n_2097));
OR2X1 g67048(.A (g2398), .B (n_2078), .Y (n_2096));
OR2X1 g67041(.A (g1785), .B (n_2098), .Y (n_2095));
NAND2X1 g67042(.A (g2691), .B (n_1596), .Y (n_2094));
OR2X1 g67044(.A (g1115), .B (n_2343), .Y (n_2093));
OR2X1 g67069(.A (g2219), .B (n_3770), .Y (n_2092));
NAND2X1 g67078(.A (g2682), .B (n_1596), .Y (n_2091));
OR2X1 g67086(.A (n_749), .B (n_2102), .Y (n_2090));
CLKBUFX1 gbuf_d_1094(.A(n_1796), .Y(d_out_1094));
CLKBUFX1 gbuf_q_1094(.A(q_in_1094), .Y(g2089));
NOR2X1 g67102(.A (g846), .B (n_8346), .Y (n_2089));
OR2X1 g67103(.A (g1525), .B (n_2194), .Y (n_2087));
NOR2X1 g67109(.A (g1531), .B (n_2194), .Y (n_2086));
OR2X1 g67116(.A (g1030), .B (n_2361), .Y (n_2084));
OR2X1 g67118(.A (g1537), .B (n_2194), .Y (n_2083));
OR2X1 g67121(.A (g1540), .B (n_2194), .Y (n_8277));
NOR2X1 g67124(.A (g834), .B (n_8346), .Y (n_2081));
OR2X1 g67125(.A (g867), .B (n_8339), .Y (n_2080));
OR2X1 g67135(.A (n_72), .B (n_8949), .Y (n_2076));
OR2X1 g67140(.A (n_39), .B (n_8949), .Y (n_2075));
OR2X1 g67141(.A (g2479), .B (n_2078), .Y (n_2074));
NOR2X1 g67142(.A (g2388), .B (n_2078), .Y (n_2073));
OR2X1 g67146(.A (g2394), .B (n_2078), .Y (n_2072));
OR2X1 g67149(.A (n_848), .B (n_2102), .Y (n_2071));
NOR2X1 g67202(.A (g1513), .B (n_2194), .Y (n_2070));
OR2X1 g67208(.A (g837), .B (n_8346), .Y (n_2069));
OR2X1 g67220(.A (g_10959), .B (n_2115), .Y (n_2068));
OR2X1 g67222(.A (g1534), .B (n_2194), .Y (n_2067));
OR2X1 g67223(.A (g1546), .B (n_2194), .Y (n_2066));
OR2X1 g67230(.A (g840), .B (n_8326), .Y (n_2065));
INVX1 g67331(.A (n_2063), .Y (n_3810));
INVX1 g67332(.A (n_2063), .Y (n_8264));
NAND2X2 g67346(.A (n_2115), .B (n_666), .Y (n_2061));
INVX1 g67374(.A (n_3482), .Y (n_2503));
INVX1 g67516(.A (g7014), .Y (n_3036));
INVX4 g67610(.A (n_2874), .Y (g6447));
INVX1 g67570(.A (n_2194), .Y (g6782));
AOI21X1 g62975(.A0 (n_1675), .A1 (g7487), .B0 (g2813), .Y (n_2058));
OR2X1 g67013(.A (g2231), .B (n_3770), .Y (n_2056));
CLKBUFX1 gbuf_d_1095(.A(n_1792), .Y(d_out_1095));
CLKBUFX1 gbuf_q_1095(.A(q_in_1095), .Y(g2101));
AOI21X1 g63101(.A0 (n_1966), .A1 (g7357), .B0 (g2119), .Y (n_2055));
NOR2X1 g66998(.A (g1697), .B (n_2052), .Y (n_2053));
CLKBUFX1 gbuf_d_1096(.A(n_1798), .Y(d_out_1096));
CLKBUFX1 gbuf_q_1096(.A(q_in_1096), .Y(g2083));
NAND2X1 g63175(.A (n_1678), .B (g739), .Y (n_2051));
CLKBUFX1 gbuf_d_1097(.A(n_1786), .Y(d_out_1097));
CLKBUFX1 gbuf_q_1097(.A(q_in_1097), .Y(g2788));
INVX2 g67254(.A (n_3781), .Y (n_4412));
CLKBUFX1 gbuf_d_1098(.A(n_1799), .Y(d_out_1098));
CLKBUFX1 gbuf_q_1098(.A(q_in_1098), .Y(g2082));
CLKBUFX1 gbuf_d_1099(.A(n_1800), .Y(d_out_1099));
CLKBUFX1 gbuf_q_1099(.A(q_in_1099), .Y(g2079));
AND2X1 g63466(.A (n_3863), .B (n_4085), .Y (n_3890));
AOI21X1 g62286(.A0 (n_1181), .A1 (n_32), .B0 (n_1921), .Y (n_2048));
CLKBUFX1 gbuf_d_1100(.A(n_1805), .Y(d_out_1100));
CLKBUFX1 gbuf_q_1100(.A(q_in_1100), .Y(g2080));
NAND2X2 g67253(.A (n_2052), .B (n_755), .Y (n_2046));
OAI21X1 g62651(.A0 (g666), .A1 (n_2207), .B0 (n_1821), .Y (n_2044));
NAND2X1 g63604(.A (n_1749), .B (g2119), .Y (n_2043));
NOR2X1 g67234(.A (g843), .B (n_8346), .Y (n_2042));
NOR2X1 g63766(.A (n_1747), .B (n_1355), .Y (n_2041));
CLKBUFX1 gbuf_d_1101(.A(n_1722), .Y(d_out_1101));
CLKBUFX1 gbuf_q_1101(.A(q_in_1101), .Y(g3018));
BUFX3 g66920(.A (g1315), .Y (n_2410));
INVX1 g67333(.A (n_8720), .Y (n_2063));
CLKBUFX1 gbuf_d_1102(.A(g7487), .Y(d_out_1102));
CLKBUFX1 gbuf_qn_1102(.A(qn_in_1102), .Y(n_2419));
CLKBUFX1 gbuf_d_1103(.A(n_1734), .Y(d_out_1103));
CLKBUFX1 gbuf_q_1103(.A(q_in_1103), .Y(g_24786));
AOI21X1 g66096(.A0 (g1255), .A1 (n_1660), .B0 (n_963), .Y (n_2040));
OR2X1 g64163(.A (n_2039), .B (n_2038), .Y (n_3421));
AND2X1 g64168(.A (n_2039), .B (n_2038), .Y (n_2211));
INVX1 g64170(.A (n_2036), .Y (n_2037));
NOR2X1 g64172(.A (n_3735), .B (n_4027), .Y (n_2035));
INVX1 g67191(.A (n_1885), .Y (n_2034));
CLKBUFX1 gbuf_d_1104(.A(n_1676), .Y(d_out_1104));
CLKBUFX1 gbuf_q_1104(.A(q_in_1104), .Y(g2924));
CLKBUFX1 gbuf_d_1105(.A(g6911), .Y(d_out_1105));
CLKBUFX1 gbuf_qn_1105(.A(qn_in_1105), .Y(g629));
AOI21X1 g61801(.A0 (n_1219), .A1 (n_116), .B0 (n_1703), .Y (n_2033));
INVX1 g64410(.A (n_2031), .Y (n_2032));
CLKBUFX1 gbuf_d_1106(.A(n_1737), .Y(d_out_1106));
CLKBUFX1 gbuf_q_1106(.A(q_in_1106), .Y(g1560));
CLKBUFX1 gbuf_d_1107(.A(n_1724), .Y(d_out_1107));
CLKBUFX1 gbuf_q_1107(.A(q_in_1107), .Y(g3032));
OR2X1 g67168(.A (n_942), .B (n_8891), .Y (n_2030));
CLKBUFX1 gbuf_d_1108(.A(n_1736), .Y(d_out_1108));
CLKBUFX1 gbuf_q_1108(.A(q_in_1108), .Y(g2254));
CLKBUFX1 gbuf_d_1109(.A(n_1733), .Y(d_out_1109));
CLKBUFX1 gbuf_q_1109(.A(q_in_1109), .Y(g_19787));
INVX2 g66723(.A (g2009), .Y (n_2292));
CLKBUFX1 gbuf_d_1110(.A(n_1742), .Y(d_out_1110));
CLKBUFX1 gbuf_q_1110(.A(q_in_1110), .Y(g1557));
CLKBUFX1 gbuf_d_1111(.A(n_1739), .Y(d_out_1111));
CLKBUFX1 gbuf_q_1111(.A(q_in_1111), .Y(g_24794));
CLKBUFX1 gbuf_d_1112(.A(n_1752), .Y(d_out_1112));
CLKBUFX1 gbuf_q_1112(.A(q_in_1112), .Y(g2912));
NAND3X1 g62504(.A (n_1682), .B (n_1196), .C (n_1165), .Y (g26149));
CLKBUFX1 gbuf_d_1113(.A(n_1743), .Y(d_out_1113));
CLKBUFX1 gbuf_q_1113(.A(q_in_1113), .Y(g2245));
CLKBUFX1 gbuf_d_1114(.A(n_1746), .Y(d_out_1114));
CLKBUFX1 gbuf_q_1114(.A(q_in_1114), .Y(g1554));
NAND2X1 g65411(.A (n_1716), .B (n_2653), .Y (n_2025));
NAND2X1 g65412(.A (n_1681), .B (n_2653), .Y (n_2024));
NAND2X1 g65413(.A (n_1714), .B (n_2653), .Y (n_2023));
NAND2X1 g65427(.A (n_1712), .B (n_2797), .Y (n_2022));
NAND2X1 g65428(.A (n_1710), .B (n_2020), .Y (n_2021));
NAND2X1 g65497(.A (n_1708), .B (n_2508), .Y (n_2019));
INVX1 g67375(.A (n_1990), .Y (n_3482));
CLKBUFX1 gbuf_d_1115(.A(n_1745), .Y(d_out_1115));
CLKBUFX1 gbuf_q_1115(.A(q_in_1115), .Y(g857));
AOI21X1 g65864(.A0 (n_1501), .A1 (n_2170), .B0 (n_1748), .Y (n_2018));
AOI21X1 g65873(.A0 (n_1466), .A1 (n_2014), .B0 (n_1702), .Y (n_2017));
NAND2X1 g65922(.A (n_1700), .B (n_3264), .Y (n_2016));
AOI21X1 g65926(.A0 (n_66), .A1 (n_2014), .B0 (n_1701), .Y (n_2015));
AOI21X1 g65957(.A0 (n_1469), .A1 (n_864), .B0 (n_1732), .Y (n_2013));
CLKBUFX1 gbuf_d_1116(.A(n_1744), .Y(d_out_1116));
CLKBUFX1 gbuf_q_1116(.A(q_in_1116), .Y(g_25781));
AOI21X1 g66028(.A0 (g569), .A1 (n_1911), .B0 (n_966), .Y (n_2012));
AOI22X1 g66037(.A0 (n_1573), .A1 (g1956), .B0 (g1957), .B1 (n_864),.Y (n_2011));
CLKBUFX1 gbuf_d_1117(.A(n_1740), .Y(d_out_1117));
CLKBUFX1 gbuf_q_1117(.A(q_in_1117), .Y(g1551));
AOI21X1 g66513(.A0 (g617), .A1 (n_1494), .B0 (g614), .Y (n_2009));
AOI22X1 g66531(.A0 (n_709), .A1 (g1966), .B0 (g1965), .B1 (n_1689),.Y (n_2008));
AOI22X1 g66565(.A0 (n_809), .A1 (g1091), .B0 (g1090), .B1 (n_8719),.Y (n_2007));
INVX1 g66957(.A (n_1770), .Y (n_2006));
CLKBUFX1 gbuf_d_1118(.A(n_1725), .Y(d_out_1118));
CLKBUFX1 gbuf_q_1118(.A(q_in_1118), .Y(g3036));
INVX1 g67015(.A (n_1842), .Y (n_2005));
INVX1 g67061(.A (n_1896), .Y (n_2004));
NOR2X1 g67129(.A (n_834), .B (n_8941), .Y (n_2003));
NOR2X1 g67134(.A (n_796), .B (n_8891), .Y (n_2001));
OR2X1 g67159(.A (n_830), .B (n_8941), .Y (n_2000));
CLKBUFX2 g67611(.A (n_2115), .Y (n_2874));
INVX1 g67206(.A (n_1879), .Y (n_1999));
INVX1 g67211(.A (n_1876), .Y (n_1998));
INVX1 g67216(.A (n_1874), .Y (n_1997));
INVX2 g67256(.A (n_8948), .Y (n_3781));
NOR2X1 g67363(.A (g1947), .B (n_1689), .Y (n_1992));
CLKBUFX3 g67376(.A (n_1990), .Y (n_3799));
INVX1 g67038(.A (n_1899), .Y (n_1989));
INVX1 g67517(.A (n_2098), .Y (g7014));
INVX1 g67735(.A (n_2078), .Y (n_2180));
INVX2 g67754(.A (n_9439), .Y (n_2232));
NAND2X1 g67030(.A (g1557), .B (n_8941), .Y (n_1986));
NAND2X1 g62940(.A (n_1984), .B (g2812), .Y (n_1985));
INVX1 g67542(.A (n_2361), .Y (n_1983));
NAND2X1 g63150(.A (n_1982), .B (g6677), .Y (n_2300));
OAI21X1 g63304(.A0 (g2714), .A1 (n_1979), .B0 (n_1677), .Y (n_1980));
OAI21X1 g63307(.A0 (g2707), .A1 (n_1979), .B0 (n_1764), .Y (n_1978));
OAI21X1 g63310(.A0 (g2727), .A1 (n_1979), .B0 (n_1763), .Y (n_1977));
OAI21X1 g63313(.A0 (g2720), .A1 (n_1979), .B0 (n_1765), .Y (n_1976));
OAI21X1 g63316(.A0 (g2734), .A1 (n_1979), .B0 (n_1762), .Y (n_1975));
OAI21X1 g63318(.A0 (g2746), .A1 (n_1979), .B0 (n_1761), .Y (n_1974));
OAI21X1 g63321(.A0 (g2740), .A1 (n_1979), .B0 (n_1760), .Y (n_1973));
OAI21X1 g63325(.A0 (n_3143), .A1 (n_1979), .B0 (n_1673), .Y (n_1972));
OAI21X1 g63328(.A0 (g2760), .A1 (n_1979), .B0 (n_1759), .Y (n_1971));
OAI21X1 g63331(.A0 (g2766), .A1 (n_1979), .B0 (n_1758), .Y (n_1970));
INVX1 g63564(.A (n_1968), .Y (n_2217));
INVX1 g66955(.A (n_1769), .Y (n_1967));
NAND2X1 g63674(.A (n_1966), .B (g7229), .Y (n_2220));
AND2X1 g63717(.A (n_1952), .B (n_1963), .Y (n_1964));
NAND2X1 g63725(.A (n_1518), .B (n_3427), .Y (n_1962));
AND2X1 g63727(.A (n_1518), .B (n_1959), .Y (n_1960));
CLKBUFX1 gbuf_d_1119(.A(n_1577), .Y(d_out_1119));
CLKBUFX1 gbuf_qn_1119(.A(qn_in_1119), .Y(g2877));
CLKBUFX1 gbuf_d_1120(.A(g25442), .Y(d_out_1120));
CLKBUFX1 gbuf_qn_1120(.A(qn_in_1120), .Y(g3111));
OR2X1 g67215(.A (n_1956), .B (n_8949), .Y (n_1957));
CLKBUFX1 gbuf_d_1121(.A(g7161), .Y(d_out_1121));
CLKBUFX1 gbuf_qn_1121(.A(qn_in_1121), .Y(g1315));
CLKBUFX1 gbuf_d_1122(.A(n_1593), .Y(d_out_1122));
CLKBUFX1 gbuf_q_1122(.A(q_in_1122), .Y(g8096));
INVX1 g64158(.A (n_1954), .Y (n_1955));
NOR2X1 g64169(.A (n_3882), .B (n_1754), .Y (n_3906));
NAND2X1 g64171(.A (n_1952), .B (n_1944), .Y (n_2036));
NOR2X1 g64178(.A (n_1518), .B (n_1264), .Y (n_1951));
CLKBUFX1 gbuf_d_1123(.A(n_1594), .Y(d_out_1123));
CLKBUFX1 gbuf_q_1123(.A(q_in_1123), .Y(g7519));
CLKBUFX1 gbuf_d_1124(.A(n_1651), .Y(d_out_1124));
CLKBUFX1 gbuf_q_1124(.A(q_in_1124), .Y(g863));
CLKBUFX1 gbuf_d_1125(.A(gbuf73), .Y(d_out_1125));
CLKBUFX1 gbuf_q_1125(.A(q_in_1125), .Y(g5595));
OAI21X1 g66544(.A0 (n_1568), .A1 (n_1245), .B0 (n_1601), .Y (n_1949));
CLKBUFX1 gbuf_d_1126(.A(g25442), .Y(d_out_1126));
CLKBUFX1 gbuf_q_1126(.A(q_in_1126), .Y(g3124));
INVX1 g67803(.A (n_1945), .Y (n_2205));
CLKBUFX1 gbuf_d_1127(.A(n_1650), .Y(d_out_1127));
CLKBUFX1 gbuf_q_1127(.A(q_in_1127), .Y(g866));
INVX1 g67802(.A (n_1945), .Y (n_1946));
NOR2X1 g64403(.A (n_1952), .B (n_1754), .Y (n_4082));
NOR2X1 g64405(.A (n_1727), .B (n_2038), .Y (n_4085));
NAND2X1 g64411(.A (n_3882), .B (n_1944), .Y (n_2031));
CLKBUFX1 gbuf_d_1128(.A(gbuf24), .Y(d_out_1128));
CLKBUFX1 gbuf_q_1128(.A(q_in_1128), .Y(g5549));
CLKBUFX1 gbuf_d_1129(.A(gbuf122), .Y(d_out_1129));
CLKBUFX1 gbuf_q_1129(.A(q_in_1129), .Y(g5612));
CLKBUFX1 gbuf_d_1130(.A(gbuf171), .Y(d_out_1130));
CLKBUFX1 gbuf_q_1130(.A(q_in_1130), .Y(g5637));
CLKBUFX1 gbuf_d_1131(.A(n_1653), .Y(d_out_1131));
CLKBUFX1 gbuf_q_1131(.A(q_in_1131), .Y(g860));
CLKBUFX1 gbuf_d_1132(.A(g25442), .Y(d_out_1132));
CLKBUFX1 gbuf_q_1132(.A(q_in_1132), .Y(g3194));
OR2X1 g67139(.A (n_1942), .B (n_8949), .Y (n_1943));
CLKBUFX1 gbuf_d_1133(.A(g25420), .Y(d_out_1133));
CLKBUFX1 gbuf_q_1133(.A(q_in_1133), .Y(g3126));
NAND2X1 g65423(.A (n_1619), .B (n_2020), .Y (n_1938));
NAND2X1 g65425(.A (n_1626), .B (n_9211), .Y (n_9583));
NAND2X1 g65426(.A (n_1624), .B (n_9211), .Y (n_1936));
CLKBUFX1 gbuf_d_1134(.A(g25420), .Y(d_out_1134));
CLKBUFX1 gbuf_q_1134(.A(q_in_1134), .Y(g3198));
NAND2X1 g65434(.A (n_1618), .B (n_2635), .Y (n_1935));
NAND2X1 g65437(.A (n_1621), .B (n_2508), .Y (n_1934));
NAND2X1 g65460(.A (n_1608), .B (n_2508), .Y (n_1933));
NAND2X1 g65466(.A (n_1649), .B (n_2508), .Y (n_1932));
NAND2X1 g65467(.A (n_1613), .B (n_2508), .Y (n_1930));
NAND2X1 g65470(.A (n_1610), .B (n_2508), .Y (n_1929));
NAND2X1 g65515(.A (n_1609), .B (n_2508), .Y (n_9609));
NAND2X1 g67377(.A (n_9592), .B (n_9593), .Y (n_1990));
INVX1 g67083(.A (n_3835), .Y (n_5181));
AOI21X1 g65832(.A0 (n_132), .A1 (n_6822), .B0 (n_1572), .Y (n_1926));
CLKBUFX1 gbuf_d_1135(.A(n_1656), .Y(d_out_1135));
CLKBUFX1 gbuf_q_1135(.A(q_in_1135), .Y(g2251));
NOR2X1 g67371(.A (g567), .B (n_1911), .Y (n_1924));
NAND2X1 g65916(.A (n_1667), .B (n_3093), .Y (n_1922));
CLKBUFX1 gbuf_d_1136(.A(n_1657), .Y(d_out_1136));
CLKBUFX1 gbuf_q_1136(.A(q_in_1136), .Y(g2248));
OR2X1 g62420(.A (n_1751), .B (n_1571), .Y (n_1921));
AOI22X1 g66066(.A0 (n_1500), .A1 (g1262), .B0 (g1263), .B1 (n_2014),.Y (n_1920));
OR2X1 g67071(.A (n_843), .B (n_8949), .Y (n_1919));
CLKBUFX1 gbuf_d_1137(.A(g25420), .Y(d_out_1137));
CLKBUFX1 gbuf_qn_1137(.A(qn_in_1137), .Y(g3112));
INVX1 g62524(.A (n_2186), .Y (n_1918));
OAI21X1 g66505(.A0 (n_1816), .A1 (n_1916), .B0 (n_1636), .Y (n_1917));
AOI21X1 g66509(.A0 (g1997), .A1 (g7194), .B0 (g1994), .Y (n_1915));
AOI22X1 g66532(.A0 (n_718), .A1 (g580), .B0 (g579), .B1 (n_1911), .Y(n_1914));
AOI22X1 g66581(.A0 (n_721), .A1 (g586), .B0 (g585), .B1 (n_1499), .Y(n_1913));
AOI22X1 g66591(.A0 (n_686), .A1 (g583), .B0 (g582), .B1 (n_1911), .Y(n_1912));
AOI21X1 g66607(.A0 (g2673), .A1 (g7390), .B0 (g2670), .Y (n_1910));
AOI22X1 g66608(.A0 (n_719), .A1 (g1272), .B0 (g1271), .B1 (n_1660),.Y (n_1909));
NOR2X1 g66635(.A (n_1597), .B (g2639), .Y (n_1908));
CLKBUFX1 gbuf_d_1138(.A(g7357), .Y(d_out_1138));
CLKBUFX1 gbuf_q_1138(.A(q_in_1138), .Y(g2009));
OR2X1 g66951(.A (n_799), .B (n_9380), .Y (n_1907));
NAND2X1 g66981(.A (g999), .B (n_8719), .Y (n_1906));
OR2X1 g66989(.A (n_806), .B (n_9380), .Y (n_1904));
OR2X1 g67002(.A (n_841), .B (n_8949), .Y (n_1902));
OR2X1 g67032(.A (n_1900), .B (n_9380), .Y (n_1901));
NOR2X1 g67039(.A (g861), .B (n_8351), .Y (n_1899));
OR2X1 g67045(.A (g2804), .B (n_1265), .Y (n_1898));
OR2X1 g67050(.A (g730), .B (n_1497), .Y (n_1897));
NOR2X1 g67062(.A (n_1895), .B (n_8355), .Y (n_1896));
OR2X1 g67073(.A (n_1893), .B (n_8949), .Y (n_1894));
INVX1 g67093(.A (n_3674), .Y (n_5372));
NAND2X1 g67174(.A (g1002), .B (n_8719), .Y (n_1888));
AND2X1 g67184(.A (g1005), .B (n_8719), .Y (n_1887));
OR2X1 g67187(.A (g1010), .B (n_8719), .Y (n_1886));
NOR2X1 g67192(.A (n_1884), .B (n_8353), .Y (n_1885));
OR2X1 g67193(.A (n_1882), .B (n_9380), .Y (n_1883));
NOR2X1 g67207(.A (n_1878), .B (n_8355), .Y (n_1879));
NOR2X1 g67212(.A (n_1875), .B (n_8355), .Y (n_1876));
NOR2X1 g67217(.A (n_1873), .B (n_8353), .Y (n_1874));
OR2X1 g67227(.A (n_811), .B (n_9380), .Y (n_1868));
NOR2X1 g67307(.A (g1253), .B (n_1660), .Y (n_1866));
OR2X1 g67040(.A (n_758), .B (n_8949), .Y (n_1864));
INVX1 g67518(.A (g_8670), .Y (n_2098));
INVX1 g67543(.A (g6712), .Y (n_2361));
INVX2 g67612(.A (g_19017), .Y (n_2115));
INVX2 g67736(.A (g_10341), .Y (n_2078));
INVX2 g67753(.A (g_20948), .Y (n_2102));
INVX2 g67817(.A (n_1945), .Y (n_3770));
AOI21X1 g66606(.A0 (g2664), .A1 (g7390), .B0 (g2661), .Y (n_1856));
INVX4 g67572(.A (n_1861), .Y (n_2194));
NAND2X1 g62973(.A (n_2203), .B (g1385), .Y (n_1854));
NAND2X1 g62974(.A (n_2160), .B (g1386), .Y (n_1853));
NAND2X1 g62977(.A (n_2203), .B (g1388), .Y (n_1852));
NAND2X1 g62978(.A (n_2160), .B (g1389), .Y (n_1851));
NAND2X1 g62982(.A (n_2203), .B (g1391), .Y (n_1850));
NAND2X1 g62983(.A (n_2160), .B (g1392), .Y (n_1849));
NAND2X1 g62985(.A (n_2203), .B (g1394), .Y (n_1848));
NAND2X1 g62986(.A (n_2160), .B (g1395), .Y (n_1847));
NAND2X1 g62988(.A (n_2203), .B (g1397), .Y (n_1846));
NAND2X1 g62990(.A (n_2160), .B (g1398), .Y (n_1845));
NAND2X1 g62994(.A (n_2203), .B (g1400), .Y (n_1844));
NAND2X1 g62995(.A (n_2160), .B (g1401), .Y (n_1843));
NOR2X1 g67016(.A (n_1841), .B (n_8353), .Y (n_1842));
NAND2X1 g62997(.A (n_2203), .B (g1403), .Y (n_1840));
NAND2X1 g62998(.A (n_2160), .B (g1404), .Y (n_1839));
NAND2X1 g63000(.A (n_2203), .B (g1406), .Y (n_1838));
NAND2X1 g63001(.A (n_2160), .B (g1407), .Y (n_1837));
NAND2X1 g63003(.A (n_2203), .B (g1409), .Y (n_1836));
NAND2X1 g63004(.A (n_2160), .B (g1410), .Y (n_1835));
NAND2X1 g63007(.A (n_2203), .B (g1412), .Y (n_1834));
NAND2X1 g63008(.A (n_2160), .B (g1413), .Y (n_1833));
NAND2X1 g63021(.A (n_2201), .B (g714), .Y (n_1832));
NAND2X1 g63025(.A (n_2203), .B (n_21), .Y (n_1831));
NAND2X1 g63026(.A (n_2160), .B (n_25), .Y (n_1830));
NAND2X1 g63028(.A (n_2201), .B (g711), .Y (n_1829));
NAND2X1 g63035(.A (g709), .B (n_2207), .Y (n_1828));
NAND2X1 g63074(.A (n_2201), .B (g699), .Y (n_1827));
NAND2X1 g63075(.A (g700), .B (n_2207), .Y (n_1826));
NAND2X1 g63076(.A (g703), .B (n_2207), .Y (n_1825));
NAND2X1 g63077(.A (n_2201), .B (g708), .Y (n_1824));
NAND2X1 g63078(.A (g712), .B (n_2207), .Y (n_1823));
NAND2X1 g63079(.A (g715), .B (n_2207), .Y (n_1822));
NAND2X1 g63080(.A (g718), .B (n_2207), .Y (n_1821));
NAND2X1 g63081(.A (g721), .B (n_2207), .Y (n_1820));
NAND2X1 g63082(.A (g724), .B (n_2207), .Y (n_1819));
NAND2X1 g63083(.A (g727), .B (n_2207), .Y (n_1818));
NAND2X1 g63085(.A (n_2201), .B (n_1816), .Y (n_1817));
NAND2X1 g63086(.A (n_2207), .B (n_1635), .Y (n_1815));
NAND2X1 g63096(.A (n_2201), .B (g723), .Y (n_1814));
NAND2X1 g63100(.A (g706), .B (n_2207), .Y (n_1813));
NAND2X1 g63105(.A (n_2201), .B (g705), .Y (n_1812));
NAND2X1 g63144(.A (n_2201), .B (g726), .Y (n_1810));
NAND2X1 g63146(.A (n_2201), .B (g702), .Y (n_1809));
NAND2X1 g63174(.A (n_2201), .B (g717), .Y (n_1808));
NAND2X1 g63181(.A (n_2201), .B (g720), .Y (n_1807));
AOI21X1 g66593(.A0 (g2568), .A1 (g7390), .B0 (g2565), .Y (n_1806));
CLKBUFX1 gbuf_d_1139(.A(n_1575), .Y(d_out_1139));
CLKBUFX1 gbuf_qn_1139(.A(qn_in_1139), .Y(g2878));
OAI21X1 g63265(.A0 (g2020), .A1 (n_1804), .B0 (n_1564), .Y (n_1805));
OAI21X1 g63266(.A0 (n_1802), .A1 (g2066), .B0 (n_1561), .Y (n_1803));
OAI21X1 g63269(.A0 (g2040), .A1 (n_1804), .B0 (n_1551), .Y (n_1801));
OAI21X1 g63272(.A0 (n_1802), .A1 (g2020), .B0 (n_1554), .Y (n_1800));
OAI21X1 g63274(.A0 (n_1802), .A1 (g2013), .B0 (n_1553), .Y (n_1799));
OAI21X1 g63275(.A0 (g2013), .A1 (n_1804), .B0 (n_1552), .Y (n_1798));
OAI21X1 g63277(.A0 (n_1802), .A1 (g2033), .B0 (n_1543), .Y (n_1797));
INVX2 g67519(.A (g_8670), .Y (n_2052));
OAI21X1 g63280(.A0 (g2026), .A1 (n_1804), .B0 (n_1546), .Y (n_1796));
OAI21X1 g63282(.A0 (g2052), .A1 (n_1804), .B0 (n_1556), .Y (n_1795));
OAI21X1 g63283(.A0 (n_1802), .A1 (g2046), .B0 (n_1563), .Y (n_1794));
OAI21X1 g63285(.A0 (n_1802), .A1 (n_2834), .B0 (n_1550), .Y (n_1793));
OAI21X1 g63286(.A0 (n_2834), .A1 (n_1804), .B0 (n_1549), .Y (n_1792));
OAI21X1 g63288(.A0 (g2066), .A1 (n_1804), .B0 (n_1559), .Y (n_1791));
OAI21X1 g63289(.A0 (n_1802), .A1 (g2072), .B0 (n_1560), .Y (n_1790));
OAI21X1 g63290(.A0 (g2072), .A1 (n_1804), .B0 (n_1548), .Y (n_1789));
OAI21X1 g63292(.A0 (n_1802), .A1 (g2040), .B0 (n_1547), .Y (n_1788));
OAI21X1 g63294(.A0 (g2033), .A1 (n_1804), .B0 (n_1542), .Y (n_1787));
OAI21X1 g63295(.A0 (n_1785), .A1 (g2746), .B0 (n_1669), .Y (n_1786));
OAI21X1 g63297(.A0 (n_1802), .A1 (g2026), .B0 (n_1544), .Y (n_1784));
OAI21X1 g63298(.A0 (g2046), .A1 (n_1804), .B0 (n_1541), .Y (n_1783));
OAI21X1 g63299(.A0 (n_1802), .A1 (g2052), .B0 (n_1540), .Y (n_1782));
OAI21X1 g63303(.A0 (n_1785), .A1 (g2714), .B0 (n_1672), .Y (n_1781));
OAI21X1 g63306(.A0 (n_1785), .A1 (g2707), .B0 (n_1671), .Y (n_1780));
OAI21X1 g63309(.A0 (n_1785), .A1 (g2727), .B0 (n_1562), .Y (n_1779));
OAI21X1 g63312(.A0 (n_1785), .A1 (g2720), .B0 (n_1670), .Y (n_1778));
OAI21X1 g63315(.A0 (n_1785), .A1 (g2734), .B0 (n_1539), .Y (n_1777));
OAI21X1 g63320(.A0 (n_1785), .A1 (g2740), .B0 (n_1555), .Y (n_1776));
OAI21X1 g63324(.A0 (n_1785), .A1 (n_3143), .B0 (n_1668), .Y (n_1775));
OAI21X1 g63327(.A0 (n_1785), .A1 (g2760), .B0 (n_1565), .Y (n_1774));
OAI21X1 g63330(.A0 (n_1785), .A1 (g2766), .B0 (n_1538), .Y (n_1773));
AND2X1 g63489(.A (n_1952), .B (n_3881), .Y (n_4380));
NAND2X1 g63503(.A (n_1531), .B (g2813), .Y (n_1772));
NOR2X1 g63565(.A (n_1567), .B (g1316), .Y (n_1968));
NOR2X1 g66958(.A (g864), .B (n_8355), .Y (n_1770));
NOR2X1 g66956(.A (n_1768), .B (n_8353), .Y (n_1769));
AND2X1 g63711(.A (n_1665), .B (n_1766), .Y (n_1767));
NAND2X1 g63731(.A (n_1979), .B (g2783), .Y (n_1765));
NAND2X1 g63739(.A (n_1979), .B (g2777), .Y (n_1764));
NAND2X1 g63741(.A (n_1979), .B (g2780), .Y (n_1763));
NAND2X1 g63745(.A (n_1979), .B (g2786), .Y (n_1762));
NAND2X1 g63749(.A (n_1979), .B (g2789), .Y (n_1761));
NAND2X1 g63751(.A (n_1979), .B (g2792), .Y (n_1760));
NAND2X1 g63756(.A (n_1979), .B (g2798), .Y (n_1759));
NAND2X1 g63759(.A (n_1979), .B (g2801), .Y (n_1758));
CLKBUFX1 gbuf_d_1140(.A(n_1529), .Y(d_out_1140));
CLKBUFX1 gbuf_qn_1140(.A(qn_in_1140), .Y(g3125));
NAND2X1 g64159(.A (n_3863), .B (n_2038), .Y (n_1954));
NOR2X1 g64160(.A (n_4351), .B (n_1666), .Y (n_3714));
NOR2X1 g64164(.A (n_3863), .B (n_3864), .Y (n_1756));
INVX1 g64165(.A (n_1755), .Y (n_3718));
NOR2X1 g64167(.A (n_1754), .B (n_1944), .Y (n_3705));
AND2X1 g64173(.A (n_1754), .B (n_1944), .Y (n_1963));
AOI21X1 g66086(.A0 (g2643), .A1 (n_1596), .B0 (n_871), .Y (n_1753));
OR2X1 g64266(.A (n_1348), .B (n_1751), .Y (n_1752));
AND2X1 g64294(.A (n_4351), .B (n_1750), .Y (n_4332));
INVX1 g64346(.A (n_1749), .Y (n_1966));
NOR2X1 g66530(.A (n_1502), .B (g605), .Y (n_1748));
OR2X1 g64466(.A (n_1260), .B (n_1751), .Y (n_1747));
MX2X1 g64478(.A (g1554), .B (n_364), .S0 (n_1741), .Y (n_1746));
OAI21X1 g64480(.A0 (n_2811), .A1 (n_1652), .B0 (n_1528), .Y (n_1745));
MX2X1 g64482(.A (g_25781), .B (n_3390), .S0 (n_1738), .Y (n_1744));
OAI21X1 g64485(.A0 (n_2952), .A1 (n_1735), .B0 (n_1527), .Y (n_1743));
MX2X1 g64498(.A (g1557), .B (n_365), .S0 (n_1741), .Y (n_1742));
MX2X1 g64501(.A (g1551), .B (n_2946), .S0 (n_1741), .Y (n_1740));
MX2X1 g64530(.A (g_24794), .B (n_5663), .S0 (n_1738), .Y (n_1739));
MX2X1 g64543(.A (g1560), .B (n_4861), .S0 (n_1741), .Y (n_1737));
OAI21X1 g64545(.A0 (n_4674), .A1 (n_1735), .B0 (n_1526), .Y (n_1736));
MX2X1 g64549(.A (g_24786), .B (n_5380), .S0 (n_1738), .Y (n_1734));
MX2X1 g64552(.A (g_19787), .B (n_5382), .S0 (n_1738), .Y (n_1733));
NOR2X1 g66514(.A (n_1470), .B (g1985), .Y (n_1732));
AOI22X1 g66498(.A0 (n_678), .A1 (g1963), .B0 (g1962), .B1 (n_1689),.Y (n_1731));
NAND2X1 g67085(.A (g2704), .B (g7487), .Y (n_3835));
OAI21X1 g66501(.A0 (n_1557), .A1 (n_562), .B0 (n_1504), .Y (n_1730));
NOR2X1 g64156(.A (n_1665), .B (n_1532), .Y (n_1728));
INVX1 g65161(.A (n_1727), .Y (n_2039));
AND2X1 g62097(.A (n_1454), .B (n_1723), .Y (n_1725));
AND2X1 g62102(.A (n_1723), .B (n_1496), .Y (n_1724));
NAND2X1 g62131(.A (n_1263), .B (n_1723), .Y (n_1722));
INVX1 g65328(.A (n_3882), .Y (n_3735));
NAND2X1 g65530(.A (n_1510), .B (n_2653), .Y (n_1721));
NAND2X1 g67095(.A (g630), .B (g6911), .Y (n_3674));
NAND2X1 g65836(.A (n_1507), .B (n_2653), .Y (n_1719));
NAND2X1 g65939(.A (n_1505), .B (n_2925), .Y (n_1718));
AOI22X1 g65962(.A0 (n_1426), .A1 (g2788), .B0 (g2789), .B1 (n_1245),.Y (n_1717));
AOI22X1 g65963(.A0 (n_1384), .A1 (g2800), .B0 (g2801), .B1 (n_1245),.Y (n_1716));
AOI22X1 g65966(.A0 (n_1420), .A1 (g2806), .B0 (g2807), .B1 (n_1245),.Y (n_1715));
AOI22X1 g65968(.A0 (n_1421), .A1 (g2797), .B0 (g2798), .B1 (n_1245),.Y (n_1714));
AOI22X1 g65989(.A0 (n_1425), .A1 (g708), .B0 (g709), .B1 (n_9208), .Y(n_1712));
AOI22X1 g65992(.A0 (n_1418), .A1 (g732), .B0 (g733), .B1 (n_9208), .Y(n_1711));
AOI22X1 g65993(.A0 (n_1424), .A1 (g711), .B0 (g712), .B1 (n_9208), .Y(n_1710));
NOR2X1 g66021(.A (n_664), .B (n_1508), .Y (n_1708));
AOI22X1 g66026(.A0 (n_1422), .A1 (g2776), .B0 (g2777), .B1 (n_1245),.Y (n_1707));
AOI22X1 g66098(.A0 (n_1410), .A1 (g2794), .B0 (g2795), .B1 (n_1245),.Y (n_1705));
INVX1 g67655(.A (n_1911), .Y (g6642));
NAND2X1 g62133(.A (n_1723), .B (n_1453), .Y (n_1703));
NAND2X1 g62525(.A (g2985), .B (g2984), .Y (n_2186));
CLKBUFX1 gbuf_d_1141(.A(g5437), .Y(d_out_1141));
CLKBUFX1 gbuf_q_1141(.A(q_in_1141), .Y(g_19017));
NOR2X1 g66556(.A (n_1467), .B (g1291), .Y (n_1702));
AOI21X1 g66566(.A0 (g1303), .A1 (n_1492), .B0 (g1300), .Y (n_1701));
AOI22X1 g66604(.A0 (n_535), .A1 (g1960), .B0 (g1959), .B1 (n_1689),.Y (n_1700));
OR2X1 g66992(.A (g577), .B (n_1911), .Y (n_1697));
OR2X1 g67068(.A (g1416), .B (n_8626), .Y (n_1696));
INVX1 g67164(.A (n_3664), .Y (n_4967));
OR2X1 g67197(.A (g2110), .B (n_1327), .Y (n_1693));
CLKBUFX1 gbuf_d_1142(.A(g5511), .Y(d_out_1142));
CLKBUFX1 gbuf_q_1142(.A(q_in_1142), .Y(g_8670));
INVX1 g67545(.A (n_8719), .Y (g6712));
INVX2 g67574(.A (n_8949), .Y (n_1861));
CLKBUFX1 gbuf_d_1143(.A(g5555), .Y(d_out_1143));
CLKBUFX1 gbuf_q_1143(.A(q_in_1143), .Y(g_10341));
CLKBUFX1 gbuf_d_1144(.A(g6231), .Y(d_out_1144));
CLKBUFX1 gbuf_q_1144(.A(q_in_1144), .Y(g_20948));
INVX1 g67786(.A (n_1660), .Y (g6944));
INVX1 g67818(.A (n_9380), .Y (n_1945));
CLKBUFX1 gbuf_d_1145(.A(n_1525), .Y(d_out_1145));
CLKBUFX1 gbuf_q_1145(.A(q_in_1145), .Y(g2883));
CLKBUFX1 gbuf_d_1146(.A(n_1524), .Y(d_out_1146));
CLKBUFX1 gbuf_q_1146(.A(q_in_1146), .Y(n_517));
CLKBUFX1 gbuf_d_1147(.A(n_1523), .Y(d_out_1147));
CLKBUFX1 gbuf_q_1147(.A(q_in_1147), .Y(g2888));
NOR2X1 g63210(.A (n_1372), .B (n_1537), .Y (n_1682));
AOI22X1 g65980(.A0 (n_1461), .A1 (g2779), .B0 (g2780), .B1 (n_1245),.Y (n_1681));
AND2X1 g63464(.A (n_1665), .B (n_3896), .Y (n_4098));
INVX1 g66948(.A (n_3678), .Y (n_4963));
NAND2X1 g63500(.A (n_1979), .B (n_1600), .Y (n_1679));
INVX1 g63527(.A (n_1678), .Y (n_1982));
NAND2X1 g63590(.A (n_1979), .B (g2774), .Y (n_1677));
NOR2X1 g63602(.A (n_1364), .B (n_1751), .Y (n_1676));
NAND2X1 g63605(.A (n_1675), .B (g7425), .Y (n_1984));
NAND2X1 g63652(.A (n_1979), .B (g2795), .Y (n_1673));
NAND2X1 g63734(.A (n_1785), .B (g2773), .Y (n_1672));
NAND2X1 g63738(.A (n_1785), .B (g2776), .Y (n_1671));
NAND2X1 g63743(.A (n_1785), .B (g2782), .Y (n_1670));
NAND2X1 g63747(.A (n_1785), .B (g2788), .Y (n_1669));
NAND2X1 g63753(.A (n_1785), .B (g2794), .Y (n_1668));
AOI22X1 g66570(.A0 (n_669), .A1 (g1269), .B0 (g1268), .B1 (n_1604),.Y (n_1667));
NOR2X1 g64157(.A (n_1750), .B (n_1666), .Y (n_1766));
NAND2X1 g64166(.A (n_1750), .B (n_1666), .Y (n_1755));
AND2X1 g64174(.A (n_1665), .B (n_1750), .Y (n_4115));
NOR2X1 g64300(.A (n_1665), .B (n_1666), .Y (n_3870));
NAND2X1 g64305(.A (n_1662), .B (n_2038), .Y (n_3419));
NOR2X1 g64347(.A (n_1457), .B (g2010), .Y (n_1749));
NOR2X1 g64406(.A (n_1658), .B (n_1944), .Y (n_3881));
NOR2X1 g64408(.A (n_1658), .B (n_4027), .Y (n_3562));
NOR2X1 g64423(.A (n_1518), .B (n_1535), .Y (n_3408));
NAND2X1 g67166(.A (g2010), .B (g7357), .Y (n_3664));
CLKBUFX1 gbuf_d_1148(.A(n_1387), .Y(d_out_1148));
CLKBUFX1 gbuf_q_1148(.A(q_in_1148), .Y(g2908));
MX2X1 g64488(.A (n_2809), .B (g2248), .S0 (n_1735), .Y (n_1657));
MX2X1 g64491(.A (n_4368), .B (g2251), .S0 (n_1735), .Y (n_1656));
OAI21X1 g64499(.A0 (n_1352), .A1 (n_1655), .B0 (n_1385), .Y (g25420));
OAI21X1 g64500(.A0 (n_1295), .A1 (n_1655), .B0 (n_1385), .Y (g25442));
MX2X1 g64535(.A (n_4110), .B (g860), .S0 (n_1652), .Y (n_1653));
MX2X1 g64538(.A (n_4112), .B (g863), .S0 (n_1652), .Y (n_1651));
MX2X1 g64541(.A (n_4464), .B (g866), .S0 (n_1652), .Y (n_1650));
NOR2X1 g66047(.A (n_662), .B (n_1430), .Y (n_1649));
AOI22X1 g65162(.A0 (n_1340), .A1 (n_1447), .B0 (g_27149), .B1(g_28034), .Y (n_1727));
INVX1 g65133(.A (n_1665), .Y (n_4351));
INVX2 g65329(.A (n_1952), .Y (n_3882));
CLKBUFX1 gbuf_d_1149(.A(n_3793), .Y(d_out_1149));
CLKBUFX1 gbuf_q_1149(.A(q_in_1149), .Y(gbuf122));
CLKBUFX1 gbuf_d_1150(.A(n_3793), .Y(d_out_1150));
CLKBUFX1 gbuf_q_1150(.A(q_in_1150), .Y(gbuf171));
CLKBUFX1 gbuf_d_1151(.A(n_3793), .Y(d_out_1151));
CLKBUFX1 gbuf_q_1151(.A(q_in_1151), .Y(gbuf24));
CLKBUFX1 gbuf_d_1152(.A(n_3793), .Y(d_out_1152));
CLKBUFX1 gbuf_q_1152(.A(q_in_1152), .Y(gbuf73));
NAND2X1 g65430(.A (n_1432), .B (n_8623), .Y (n_1642));
NAND2X1 g65436(.A (n_1439), .B (n_8623), .Y (n_1641));
NAND2X1 g65438(.A (n_1442), .B (n_8623), .Y (n_1639));
NAND2X1 g65462(.A (n_1438), .B (n_8623), .Y (n_1638));
OR2X1 g67088(.A (n_1635), .B (n_1497), .Y (n_1636));
NAND2X1 g65449(.A (n_1433), .B (n_8623), .Y (n_1634));
NAND2X1 g65923(.A (n_1428), .B (n_2508), .Y (n_1632));
AOI21X1 g65936(.A0 (n_151), .A1 (n_6822), .B0 (n_1427), .Y (n_1631));
AOI22X1 g65984(.A0 (n_1336), .A1 (g1412), .B0 (g1413), .B1 (n_8625),.Y (n_1629));
AOI22X1 g65985(.A0 (n_1329), .A1 (g720), .B0 (g721), .B1 (n_9208), .Y(n_1628));
AOI22X1 g65986(.A0 (n_1326), .A1 (g717), .B0 (g718), .B1 (n_9208), .Y(n_1627));
AOI22X1 g65988(.A0 (n_1334), .A1 (g705), .B0 (g706), .B1 (n_9208), .Y(n_1626));
AOI22X1 g65991(.A0 (n_1369), .A1 (g723), .B0 (g724), .B1 (n_9208), .Y(n_1624));
AOI22X1 g65994(.A0 (n_1375), .A1 (g702), .B0 (g703), .B1 (n_9208), .Y(n_9590));
AOI22X1 g66000(.A0 (n_1371), .A1 (g2103), .B0 (g2104), .B1 (n_562),.Y (n_1622));
AOI22X1 g66009(.A0 (n_1323), .A1 (g2106), .B0 (g2107), .B1 (n_562),.Y (n_1621));
AOI22X1 g66012(.A0 (n_1332), .A1 (g738), .B0 (g739), .B1 (n_9208), .Y(n_1619));
AOI22X1 g66020(.A0 (n_1304), .A1 (g1403), .B0 (g1404), .B1 (n_8625),.Y (n_1618));
AOI22X1 g66024(.A0 (n_1330), .A1 (g2079), .B0 (g2080), .B1 (n_562),.Y (n_1616));
AOI22X1 g66027(.A0 (n_1302), .A1 (g699), .B0 (g700), .B1 (n_9208), .Y(n_1615));
AOI22X1 g66041(.A0 (n_1328), .A1 (g2091), .B0 (g2092), .B1 (n_562),.Y (n_1613));
AOI22X1 g66042(.A0 (n_1321), .A1 (g2112), .B0 (g2113), .B1 (n_562),.Y (n_1612));
AOI22X1 g66049(.A0 (n_1325), .A1 (g2100), .B0 (g2101), .B1 (n_562),.Y (n_1611));
AOI22X1 g66067(.A0 (n_1322), .A1 (g2097), .B0 (g2098), .B1 (n_562),.Y (n_1610));
NOR2X1 g66068(.A (n_660), .B (n_1431), .Y (n_1609));
NOR2X1 g66071(.A (n_563), .B (n_1445), .Y (n_1608));
CLKBUFX1 gbuf_d_1153(.A(g25435), .Y(d_out_1153));
CLKBUFX1 gbuf_q_1153(.A(q_in_1153), .Y(g3197));
NAND2X1 g65433(.A (n_1441), .B (n_8623), .Y (n_1606));
AOI22X1 g66571(.A0 (n_633), .A1 (g1266), .B0 (g1265), .B1 (n_1604),.Y (n_1605));
OAI22X1 g66587(.A0 (n_21), .A1 (n_8625), .B0 (n_25), .B1 (n_8626), .Y(n_1603));
CLKBUFX1 gbuf_d_1154(.A(g25435), .Y(d_out_1154));
CLKBUFX1 gbuf_q_1154(.A(q_in_1154), .Y(g3110));
OR2X1 g66986(.A (n_1600), .B (n_1265), .Y (n_1601));
INVX1 g67285(.A (n_3264), .Y (n_1691));
NOR2X1 g67305(.A (g2641), .B (n_1596), .Y (n_1597));
MX2X1 g62749(.A (n_1574), .B (g7519), .S0 (g2879), .Y (n_1594));
MX2X1 g62750(.A (n_1576), .B (g8096), .S0 (g2879), .Y (n_1593));
NAND2X1 g67832(.A (g1696), .B (n_1235), .Y (n_1587));
NAND2X1 g67871(.A (g_20070), .B (n_1382), .Y (n_1586));
NAND2X1 g67954(.A (g231), .B (n_1382), .Y (n_9619));
NAND2X1 g67957(.A (g267), .B (n_1382), .Y (n_8226));
NAND2X1 g67958(.A (g_24437), .B (n_1382), .Y (n_1581));
NAND2X1 g67965(.A (g240), .B (n_1382), .Y (n_1580));
NAND2X1 g67972(.A (g_12763), .B (n_1237), .Y (n_9659));
MX2X1 g62835(.A (n_350), .B (n_1576), .S0 (g2879), .Y (n_1577));
MX2X1 g62836(.A (n_374), .B (n_1574), .S0 (g2879), .Y (n_1575));
OR2X1 g67014(.A (g1957), .B (n_1689), .Y (n_1573));
AOI21X1 g66595(.A0 (g2682), .A1 (g7390), .B0 (g2679), .Y (n_1572));
AOI21X1 g63213(.A0 (n_1357), .A1 (g2920), .B0 (n_476), .Y (n_1571));
NOR2X1 g63491(.A (n_1536), .B (n_1456), .Y (n_3930));
NAND2X1 g63498(.A (n_1567), .B (g6979), .Y (n_2203));
NAND2X1 g63499(.A (n_1785), .B (n_1568), .Y (n_1569));
NAND2X1 g63502(.A (n_1567), .B (g7161), .Y (n_2160));
NOR2X1 g63528(.A (n_1566), .B (g630), .Y (n_1678));
NAND2X1 g63538(.A (n_1785), .B (g2797), .Y (n_1565));
NAND2X1 g63539(.A (n_1804), .B (g2080), .Y (n_1564));
NAND2X1 g63540(.A (n_1802), .B (g2097), .Y (n_1563));
NAND2X1 g63550(.A (n_1785), .B (g2779), .Y (n_1562));
NAND2X1 g63555(.A (n_1802), .B (g2103), .Y (n_1561));
NAND2X1 g63560(.A (n_1802), .B (g2106), .Y (n_1560));
NAND2X1 g63562(.A (n_1804), .B (g2104), .Y (n_1559));
NAND2X1 g63566(.A (n_1802), .B (n_1557), .Y (n_1558));
NAND2X1 g63567(.A (n_1804), .B (g2095), .Y (n_1556));
NAND2X1 g63577(.A (n_1785), .B (g2791), .Y (n_1555));
NAND2X1 g63585(.A (n_1802), .B (g2079), .Y (n_1554));
NAND2X1 g63587(.A (n_1802), .B (g2082), .Y (n_1553));
NAND2X1 g63588(.A (n_1804), .B (g2083), .Y (n_1552));
NAND2X1 g63592(.A (n_1804), .B (g2092), .Y (n_1551));
NAND2X1 g63594(.A (n_1802), .B (g2100), .Y (n_1550));
NAND2X1 g63595(.A (n_1804), .B (g2101), .Y (n_1549));
NAND2X1 g63598(.A (n_1804), .B (g2107), .Y (n_1548));
NAND2X1 g63606(.A (n_1802), .B (g2091), .Y (n_1547));
NAND2X1 g63670(.A (n_1804), .B (g2089), .Y (n_1546));
NAND2X1 g63671(.A (n_1804), .B (n_1503), .Y (n_1545));
NAND2X1 g63673(.A (n_1802), .B (g2088), .Y (n_1544));
NAND2X1 g66950(.A (g1316), .B (g7161), .Y (n_3678));
NAND2X1 g63683(.A (n_1802), .B (g2085), .Y (n_1543));
NAND2X1 g63687(.A (n_1566), .B (g6911), .Y (n_2207));
NAND2X1 g63700(.A (n_1804), .B (g2086), .Y (n_1542));
NAND2X1 g63701(.A (n_1804), .B (g2098), .Y (n_1541));
NAND2X1 g63705(.A (n_1566), .B (g6677), .Y (n_2201));
NAND2X1 g63710(.A (n_1802), .B (g2094), .Y (n_1540));
NAND2X1 g63713(.A (n_1785), .B (g2785), .Y (n_1539));
NAND2X1 g63716(.A (n_1785), .B (g2800), .Y (n_1538));
NAND4X1 g63765(.A (n_1054), .B (n_1065), .C (n_1060), .D (n_1194), .Y(n_1537));
CLKBUFX1 gbuf_d_1155(.A(n_1353), .Y(d_out_1155));
CLKBUFX1 gbuf_q_1155(.A(q_in_1155), .Y(g2896));
CLKBUFX1 gbuf_d_1156(.A(n_1373), .Y(d_out_1156));
CLKBUFX1 gbuf_q_1156(.A(q_in_1156), .Y(g3002));
CLKBUFX1 gbuf_d_1157(.A(n_1292), .Y(d_out_1157));
CLKBUFX1 gbuf_q_1157(.A(q_in_1157), .Y(g2900));
NOR2X1 g64176(.A (n_1536), .B (n_1535), .Y (n_3904));
CLKBUFX1 gbuf_d_1158(.A(n_1339), .Y(d_out_1158));
CLKBUFX1 gbuf_q_1158(.A(q_in_1158), .Y(g3024));
INVX1 g68356(.A (n_1237), .Y (g5437));
INVX1 g64263(.A (n_1567), .Y (n_1663));
AOI22X1 g63910(.A0 (n_1271), .A1 (n_1464), .B0 (n_1463), .B1 (g3086),.Y (n_1533));
NOR2X1 g64288(.A (n_1750), .B (n_1532), .Y (n_3712));
NOR2X1 g64303(.A (n_1750), .B (n_1448), .Y (n_3896));
INVX1 g64351(.A (n_1531), .Y (n_1675));
AND2X1 g64438(.A (n_1536), .B (n_1459), .Y (n_2985));
NAND2X1 g64441(.A (n_1530), .B (g7487), .Y (n_1979));
INVX1 g64467(.A (g25435), .Y (n_1529));
NAND2X1 g64623(.A (n_1652), .B (g857), .Y (n_1528));
NAND2X1 g64626(.A (n_1735), .B (g2245), .Y (n_1527));
NAND2X1 g64631(.A (n_1735), .B (g2254), .Y (n_1526));
NAND2X1 g64641(.A (n_1349), .B (n_676), .Y (n_1525));
NOR2X1 g64642(.A (n_1354), .B (n_794), .Y (n_1524));
NAND2X1 g64644(.A (n_1299), .B (g2814), .Y (n_1751));
AOI21X1 g64738(.A0 (n_442), .A1 (n_100), .B0 (n_1320), .Y (n_1523));
INVX1 g65170(.A (n_1662), .Y (n_3863));
OAI21X1 g65331(.A0 (g1040), .A1 (g1024), .B0 (n_1300), .Y (n_1952));
INVX1 g65333(.A (n_1658), .Y (n_1754));
NAND2X1 g65938(.A (n_1338), .B (n_2925), .Y (n_1517));
AOI22X1 g65961(.A0 (n_1250), .A1 (g2791), .B0 (g2792), .B1 (n_1245),.Y (n_1516));
AOI22X1 g65971(.A0 (n_1252), .A1 (g2773), .B0 (g2774), .B1 (n_1245),.Y (n_1515));
AOI22X1 g65987(.A0 (n_1223), .A1 (g714), .B0 (g715), .B1 (n_9208), .Y(n_1514));
AOI22X1 g65990(.A0 (n_1251), .A1 (g726), .B0 (g727), .B1 (n_9208), .Y(n_1513));
AOI22X1 g66023(.A0 (n_1248), .A1 (g2650), .B0 (g2651), .B1 (n_6822),.Y (n_1511));
AOI21X1 g62403(.A0 (n_1220), .A1 (n_386), .B0 (g3234), .Y (n_1723));
AOI22X1 g66039(.A0 (n_1266), .A1 (g2782), .B0 (g2783), .B1 (n_1245),.Y (n_1510));
NOR2X1 g66187(.A (n_1335), .B (n_22), .Y (n_1508));
AOI22X1 g66580(.A0 (n_715), .A1 (g2813), .B0 (g2812), .B1 (n_1265),.Y (n_1507));
AOI22X1 g66589(.A0 (n_565), .A1 (g2657), .B0 (g2656), .B1 (n_1596),.Y (n_1506));
AOI22X1 g66602(.A0 (n_587), .A1 (g2660), .B0 (g2659), .B1 (n_1247),.Y (n_1505));
OR2X1 g66975(.A (n_1503), .B (n_1327), .Y (n_1504));
NOR2X1 g67052(.A (n_1501), .B (n_1499), .Y (n_1502));
OR2X1 g67154(.A (g1263), .B (n_1604), .Y (n_1500));
NAND2X1 g67262(.A (n_1499), .B (n_1498), .Y (n_3498));
NAND2X2 g67286(.A (n_1689), .B (n_864), .Y (n_3264));
INVX2 g67482(.A (n_1689), .Y (g7194));
XOR2X1 g62752(.A (g3032), .B (n_1275), .Y (n_1496));
CLKBUFX1 gbuf_d_1159(.A(g5472), .Y(d_out_1159));
CLKBUFX1 gbuf_q_1159(.A(q_in_1159), .Y(g_20180));
INVX2 g67658(.A (n_1494), .Y (n_1911));
INVX1 g67788(.A (n_1492), .Y (n_1660));
CLKBUFX1 gbuf_d_1160(.A(g6837), .Y(d_out_1160));
CLKBUFX1 gbuf_q_1160(.A(q_in_1160), .Y(g_9470));
CLKBUFX1 gbuf_d_1161(.A(n_1376), .Y(d_out_1161));
CLKBUFX1 gbuf_qn_1161(.A(qn_in_1161), .Y(g3123));
INVX1 g68164(.A (n_1235), .Y (n_1483));
CLKBUFX1 gbuf_d_1162(.A(n_1378), .Y(d_out_1162));
CLKBUFX1 gbuf_qn_1162(.A(qn_in_1162), .Y(g2985));
CLKBUFX1 gbuf_d_1163(.A(n_1380), .Y(d_out_1163));
CLKBUFX1 gbuf_qn_1163(.A(qn_in_1163), .Y(g2984));
CLKBUFX1 gbuf_d_1164(.A(g6573), .Y(d_out_1164));
CLKBUFX1 gbuf_q_1164(.A(q_in_1164), .Y(g_21829));
INVX2 g68440(.A (n_9512), .Y (g5555));
INVX1 g67277(.A (n_3093), .Y (n_1598));
NOR2X1 g66987(.A (n_1469), .B (n_1689), .Y (n_1470));
CLKBUFX1 gbuf_d_1165(.A(n_1366), .Y(d_out_1165));
CLKBUFX1 gbuf_q_1165(.A(q_in_1165), .Y(n_782));
NOR2X1 g66965(.A (n_1466), .B (n_1604), .Y (n_1467));
AOI22X1 g63902(.A0 (n_1273), .A1 (n_1464), .B0 (g3101), .B1 (n_1463),.Y (n_1465));
AOI22X1 g65964(.A0 (n_1268), .A1 (g2785), .B0 (g2786), .B1 (n_1245),.Y (n_1462));
OR2X1 g66945(.A (g2780), .B (n_1265), .Y (n_1461));
CLKBUFX1 gbuf_d_1166(.A(n_1278), .Y(d_out_1166));
CLKBUFX1 gbuf_q_1166(.A(q_in_1166), .Y(n_458));
AND2X1 g64177(.A (n_1518), .B (n_1459), .Y (n_3410));
AND2X1 g64179(.A (n_1535), .B (n_1459), .Y (n_1959));
CLKBUFX1 gbuf_d_1167(.A(n_1280), .Y(d_out_1167));
CLKBUFX1 gbuf_q_1167(.A(q_in_1167), .Y(g2998));
NAND3X1 g64261(.A (n_1064), .B (n_1087), .C (n_1385), .Y (n_1458));
NOR2X1 g64264(.A (n_1270), .B (g1345), .Y (n_1567));
NAND2X1 g64328(.A (n_1457), .B (g7229), .Y (n_1802));
NAND2X1 g64329(.A (n_1457), .B (g7357), .Y (n_1804));
NOR2X1 g64343(.A (n_1269), .B (g659), .Y (n_1566));
NOR2X1 g64352(.A (n_1530), .B (g2704), .Y (n_1531));
INVX1 g64425(.A (n_3575), .Y (n_1456));
NAND2X1 g64440(.A (n_1530), .B (g7425), .Y (n_1785));
INVX1 g67789(.A (n_1604), .Y (n_1492));
AOI21X1 g64456(.A0 (n_985), .A1 (n_1202), .B0 (n_969), .Y (n_1455));
OAI21X1 g64468(.A0 (n_1201), .A1 (n_1655), .B0 (n_1385), .Y (g25435));
OAI21X1 g64471(.A0 (n_1453), .A1 (g3036), .B0 (n_1274), .Y (n_1454));
NAND2X1 g67947(.A (g909), .B (n_1032), .Y (n_1452));
NOR2X1 g64175(.A (n_1535), .B (n_1459), .Y (n_3427));
INVX1 g65085(.A (n_1448), .Y (n_1666));
NAND2X1 g65139(.A (n_913), .B (n_1262), .Y (n_1665));
INVX1 g65141(.A (n_1532), .Y (n_1521));
AOI22X1 g65171(.A0 (n_1180), .A1 (n_1447), .B0 (g_13227), .B1(g_28034), .Y (n_1662));
AOI21X1 g65334(.A0 (n_1176), .A1 (n_1446), .B0 (n_1004), .Y (n_1658));
AOI21X1 g65336(.A0 (n_1174), .A1 (n_1446), .B0 (n_1003), .Y (n_1944));
AOI21X1 g65346(.A0 (n_1173), .A1 (n_1446), .B0 (n_1041), .Y (n_4027));
AOI22X1 g65347(.A0 (n_1208), .A1 (n_1447), .B0 (g_28035), .B1(g_28034), .Y (n_3864));
NOR2X1 g65416(.A (n_2915), .B (n_1285), .Y (n_1741));
CLKBUFX1 gbuf_d_1168(.A(g6368), .Y(d_out_1168));
CLKBUFX1 gbuf_q_1168(.A(q_in_1168), .Y(g_14662));
NOR2X1 g66194(.A (n_1287), .B (n_95), .Y (n_1445));
NOR2X1 g65866(.A (n_7462), .B (g1217), .Y (n_1443));
AOI22X1 g65276(.A0 (n_1179), .A1 (n_1447), .B0 (g_7905), .B1(g_28034), .Y (n_2038));
AOI22X1 g65977(.A0 (n_1218), .A1 (g1391), .B0 (g1392), .B1 (n_8625),.Y (n_1442));
AOI22X1 g65997(.A0 (n_1203), .A1 (g1409), .B0 (g1410), .B1 (n_8625),.Y (n_1441));
AOI22X1 g65999(.A0 (n_1164), .A1 (g1394), .B0 (g1395), .B1 (n_8625),.Y (n_1439));
AOI22X1 g66001(.A0 (n_1095), .A1 (g1406), .B0 (g1407), .B1 (n_8625),.Y (n_1438));
AOI22X1 g66004(.A0 (n_1155), .A1 (g1385), .B0 (g1386), .B1 (n_8625),.Y (n_1437));
AOI22X1 g66006(.A0 (n_1085), .A1 (g1418), .B0 (g1419), .B1 (n_8625),.Y (n_1436));
AOI22X1 g66014(.A0 (n_1154), .A1 (g1397), .B0 (g1398), .B1 (n_8625),.Y (n_1435));
AOI22X1 g66030(.A0 (n_1217), .A1 (g1388), .B0 (g1389), .B1 (n_8625),.Y (n_1433));
AOI22X1 g66065(.A0 (n_1088), .A1 (g1400), .B0 (g1401), .B1 (n_8625),.Y (n_1432));
NOR2X1 g66190(.A (n_1249), .B (n_70), .Y (n_1431));
NOR2X1 g66191(.A (n_1277), .B (n_53), .Y (n_1430));
AOI22X1 g66508(.A0 (n_614), .A1 (g1425), .B0 (g1424), .B1 (n_8626),.Y (n_1429));
AOI22X1 g66516(.A0 (n_624), .A1 (g2119), .B0 (g2118), .B1 (n_1327),.Y (n_1428));
AOI21X1 g66592(.A0 (g2691), .A1 (g7390), .B0 (g2688), .Y (n_1427));
OR2X1 g66944(.A (g2789), .B (n_1265), .Y (n_1426));
OR2X1 g66979(.A (g709), .B (n_1333), .Y (n_1425));
OR2X1 g66983(.A (g712), .B (n_1333), .Y (n_1424));
OR2X1 g67053(.A (g2777), .B (n_1265), .Y (n_1422));
OR2X1 g67120(.A (g2798), .B (n_1265), .Y (n_1421));
OR2X1 g67160(.A (g2807), .B (n_1265), .Y (n_1420));
OR2X1 g67198(.A (g733), .B (n_1333), .Y (n_1418));
CLKBUFX1 gbuf_d_1169(.A(g24734), .Y(d_out_1169));
CLKBUFX1 gbuf_q_1169(.A(q_in_1169), .Y(g3191));
INVX1 g67268(.A (n_1416), .Y (n_2797));
INVX2 g67269(.A (n_1416), .Y (n_2020));
NAND2X2 g67278(.A (n_1604), .B (n_2014), .Y (n_3093));
INVX1 g67464(.A (g6911), .Y (n_1497));
OR2X1 g67036(.A (g2795), .B (n_1265), .Y (n_1410));
INVX1 g67660(.A (n_1499), .Y (n_1494));
NAND2X1 g67856(.A (g2315), .B (n_1305), .Y (n_8244));
NAND2X1 g67861(.A (g1612), .B (n_1285), .Y (n_9623));
NAND2X1 g67881(.A (g2306), .B (n_1305), .Y (n_1403));
NAND2X1 g67894(.A (g1116), .B (n_8305), .Y (n_1402));
NAND2X1 g67936(.A (g1576), .B (n_1285), .Y (n_1401));
NAND2X1 g67948(.A (g882), .B (n_1032), .Y (n_1399));
NAND2X1 g67955(.A (g954), .B (n_1032), .Y (n_8268));
CLKBUFX1 gbuf_d_1170(.A(n_1225), .Y(d_out_1170));
CLKBUFX1 gbuf_q_1170(.A(q_in_1170), .Y(g3010));
NAND2X1 g68015(.A (g2342), .B (n_1305), .Y (n_8274));
NAND2X1 g68017(.A (g1002), .B (n_8305), .Y (n_1396));
NAND2X1 g68020(.A (g2270), .B (n_1305), .Y (n_9607));
NAND2X1 g68023(.A (g1621), .B (n_1392), .Y (n_9615));
NAND2X1 g68027(.A (g918), .B (n_1032), .Y (n_1391));
NAND2X1 g68035(.A (g1648), .B (n_1392), .Y (n_8218));
NAND2X1 g68048(.A (g2297), .B (n_1305), .Y (n_1389));
NAND2X1 g68050(.A (g1603), .B (n_1285), .Y (n_1388));
AOI21X1 g63207(.A0 (n_1214), .A1 (n_539), .B0 (n_1365), .Y (n_1387));
NAND3X1 g64404(.A (n_1062), .B (n_1200), .C (n_1385), .Y (n_1386));
OR2X1 g66967(.A (g2801), .B (n_1265), .Y (n_1384));
NOR2X1 g65520(.A (n_2915), .B (n_1382), .Y (n_1738));
INVX1 g68387(.A (n_1382), .Y (n_8024));
INVX2 g68391(.A (n_1382), .Y (g6231));
CLKBUFX1 gbuf_d_1171(.A(n_1190), .Y(d_out_1171));
CLKBUFX1 gbuf_q_1171(.A(q_in_1171), .Y(n_379));
XOR2X1 g63964(.A (n_1381), .B (n_1377), .Y (n_1574));
XOR2X1 g63965(.A (n_1381), .B (n_1379), .Y (n_1576));
XOR2X1 g63966(.A (g2934), .B (n_1379), .Y (n_1380));
XOR2X1 g63967(.A (g2962), .B (n_1377), .Y (n_1378));
INVX1 g66099(.A (g24734), .Y (n_1376));
OR2X1 g67059(.A (g703), .B (n_1331), .Y (n_1375));
NAND2X1 g64274(.A (n_501), .B (n_1206), .Y (n_1374));
NOR2X1 g64275(.A (n_1210), .B (n_793), .Y (n_1373));
NAND3X1 g64302(.A (n_1166), .B (n_984), .C (n_1385), .Y (n_1372));
OR2X1 g67179(.A (g2104), .B (n_1327), .Y (n_1371));
NOR2X1 g64373(.A (n_1370), .B (n_1264), .Y (n_3560));
NOR2X1 g64426(.A (n_1370), .B (n_1459), .Y (n_3575));
OR2X1 g67157(.A (g724), .B (n_1333), .Y (n_1369));
MX2X1 g64520(.A (g_16317), .B (g_22696), .S0 (g3229), .Y (n_1368));
MX2X1 g64521(.A (g1227), .B (g1224), .S0 (g3229), .Y (n_1367));
NOR2X1 g64645(.A (n_976), .B (n_1365), .Y (n_1366));
INVX1 g64654(.A (n_1457), .Y (n_1449));
XOR2X1 g64782(.A (g2924), .B (n_1181), .Y (n_1364));
CLKBUFX1 gbuf_d_1172(.A(n_1187), .Y(d_out_1172));
CLKBUFX1 gbuf_q_1172(.A(q_in_1172), .Y(g3080));
AOI22X1 g65086(.A0 (n_1057), .A1 (n_1363), .B0 (g1764), .B1 (g1718),.Y (n_1448));
AOI22X1 g65142(.A0 (n_1056), .A1 (n_1363), .B0 (g1705), .B1 (g1718),.Y (n_1532));
INVX1 g65283(.A (n_1518), .Y (n_1536));
AOI22X1 g65308(.A0 (n_1079), .A1 (n_1363), .B0 (g1749), .B1 (g1718),.Y (n_1750));
NAND2X1 g65406(.A (n_1182), .B (g2924), .Y (n_1357));
OR2X1 g65407(.A (n_1182), .B (n_986), .Y (n_1355));
OR2X1 g65410(.A (n_783), .B (n_1365), .Y (n_1354));
NOR2X1 g65422(.A (n_680), .B (n_1365), .Y (n_1353));
NAND2X1 g65431(.A (n_7337), .B (n_1192), .Y (n_7240));
OR2X1 g65445(.A (n_878), .B (n_1184), .Y (n_1352));
NAND2X1 g65465(.A (n_3793), .B (g6368), .Y (n_1652));
NAND2X1 g65479(.A (n_3793), .B (g6837), .Y (n_1735));
AOI21X1 g65614(.A0 (g2883), .A1 (n_233), .B0 (n_1365), .Y (n_1349));
XOR2X1 g65817(.A (g2912), .B (n_1001), .Y (n_1348));
NAND2X1 g65845(.A (n_1342), .B (g_11640), .Y (n_1347));
NOR2X1 g65851(.A (n_7462), .B (g1215), .Y (n_1346));
NOR2X1 g65865(.A (n_7462), .B (g1220), .Y (n_1344));
NAND2X1 g65889(.A (n_1342), .B (g_19993), .Y (n_1343));
AOI21X1 g66048(.A0 (g_9473), .A1 (g_24889), .B0 (n_1156), .Y(n_1340));
NOR2X1 g62132(.A (n_1150), .B (n_1279), .Y (n_1339));
AOI22X1 g66600(.A0 (n_494), .A1 (g2654), .B0 (g2653), .B1 (n_1247),.Y (n_1338));
NAND2X1 g65844(.A (n_1342), .B (g_9014), .Y (n_1337));
OR2X1 g66985(.A (g1413), .B (n_8626), .Y (n_1336));
NOR2X1 g67019(.A (g2095), .B (n_1327), .Y (n_1335));
OR2X1 g67020(.A (g706), .B (n_1333), .Y (n_1334));
OR2X1 g67028(.A (g739), .B (n_1331), .Y (n_1332));
INVX1 g67033(.A (n_1244), .Y (n_1330));
OR2X1 g67065(.A (g721), .B (n_1331), .Y (n_1329));
OR2X1 g67090(.A (g2092), .B (n_1327), .Y (n_1328));
OR2X1 g67097(.A (g718), .B (n_9209), .Y (n_1326));
OR2X1 g67105(.A (g2101), .B (n_1327), .Y (n_1325));
OR2X1 g67169(.A (g2107), .B (n_1327), .Y (n_1323));
OR2X1 g67176(.A (g2098), .B (n_1327), .Y (n_1322));
OR2X1 g67210(.A (g2113), .B (n_1327), .Y (n_1321));
OR2X1 g65414(.A (n_478), .B (n_1365), .Y (n_1320));
INVX1 g67271(.A (n_9211), .Y (n_1416));
CLKBUFX1 gbuf_d_1173(.A(n_1212), .Y(d_out_1173));
CLKBUFX1 gbuf_q_1173(.A(q_in_1173), .Y(g3013));
INVX1 g67465(.A (n_1333), .Y (g6911));
INVX2 g67484(.A (g_10301), .Y (n_1689));
INVX1 g67661(.A (g_15095), .Y (n_1499));
INVX1 g67744(.A (n_1265), .Y (g7487));
OR2X1 g67896(.A (g398), .B (n_1237), .Y (n_1315));
OR2X1 g67916(.A (g1779), .B (n_1235), .Y (n_1314));
OR2X1 g68009(.A (g2473), .B (n_9512), .Y (n_1313));
NAND2X1 g68019(.A (g927), .B (n_1032), .Y (n_1312));
CLKBUFX1 gbuf_d_1174(.A(n_1213), .Y(d_out_1174));
CLKBUFX1 gbuf_q_1174(.A(q_in_1174), .Y(g3006));
OR2X1 g66990(.A (g1404), .B (n_8626), .Y (n_1304));
OR2X1 g66991(.A (g700), .B (n_1331), .Y (n_1302));
INVX1 g68462(.A (n_1305), .Y (n_1301));
NAND2X1 g65519(.A (n_1177), .B (n_1446), .Y (n_1300));
NAND4X1 g65531(.A (n_1191), .B (g2912), .C (n_358), .D (g2920), .Y(n_1299));
OR2X1 g65528(.A (n_875), .B (n_1178), .Y (n_1295));
NOR2X1 g63505(.A (n_1076), .B (n_1365), .Y (n_1292));
INVX1 g67237(.A (n_1290), .Y (n_2635));
OR2X1 g67837(.A (g1765), .B (n_1235), .Y (n_1288));
NOR2X1 g67204(.A (g2083), .B (n_1327), .Y (n_1287));
INVX1 g68255(.A (n_1032), .Y (n_7675));
CLKBUFX1 gbuf_d_1175(.A(g6750), .Y(d_out_1175));
CLKBUFX1 gbuf_qn_1175(.A(qn_in_1175), .Y(n_1604));
MX2X1 g64470(.A (n_714), .B (g3234), .S0 (n_1279), .Y (n_1280));
MX2X1 g64505(.A (n_470), .B (n_310), .S0 (n_1279), .Y (n_1278));
NOR2X1 g67155(.A (g2086), .B (n_1327), .Y (n_1277));
NOR2X1 g64595(.A (n_1453), .B (n_9), .Y (n_1275));
NAND2X1 g64651(.A (n_1453), .B (g3036), .Y (n_1274));
AOI21X1 g64652(.A0 (n_117), .A1 (n_893), .B0 (n_1008), .Y (n_1273));
NOR2X1 g64655(.A (n_1068), .B (g2039), .Y (n_1457));
NOR2X1 g64665(.A (n_1066), .B (g2733), .Y (n_1530));
CLKBUFX1 gbuf_d_1176(.A(g16496), .Y(d_out_1176));
CLKBUFX1 gbuf_q_1176(.A(q_in_1176), .Y(g2987));
AOI21X1 g64688(.A0 (n_892), .A1 (n_122), .B0 (n_1067), .Y (n_1271));
NAND2X1 g64706(.A (g1211), .B (g1224), .Y (n_1270));
NAND2X1 g64733(.A (g_18792), .B (g_22696), .Y (n_1269));
OR2X1 g67133(.A (g2786), .B (n_1265), .Y (n_1268));
NAND2X1 g65284(.A (n_777), .B (n_1070), .Y (n_1518));
OR2X1 g67060(.A (g2783), .B (n_1265), .Y (n_1266));
INVX1 g65350(.A (n_1370), .Y (n_1535));
INVX1 g65355(.A (n_1264), .Y (n_1359));
XOR2X1 g65365(.A (g3018), .B (n_891), .Y (n_1263));
NAND2X1 g65447(.A (n_1058), .B (n_1363), .Y (n_1262));
NOR2X1 g65829(.A (n_1001), .B (g2917), .Y (n_1260));
NAND2X1 g65848(.A (n_1342), .B (g_11807), .Y (n_1259));
INVX1 g65859(.A (n_3793), .Y (n_2915));
NOR2X1 g65871(.A (n_7462), .B (g1219), .Y (n_1258));
OR2X1 g65892(.A (n_8103), .B (n_970), .Y (n_8111));
NOR2X1 g65893(.A (n_7462), .B (g1216), .Y (n_1257));
NOR2X1 g65918(.A (n_7462), .B (g1218), .Y (n_1256));
OAI21X1 g66100(.A0 (n_801), .A1 (n_12), .B0 (n_1385), .Y (g24734));
CLKBUFX1 gbuf_d_1177(.A(g966), .Y(d_out_1177));
CLKBUFX1 gbuf_q_1177(.A(q_in_1177), .Y(g1217));
OR2X1 g67952(.A (g384), .B (n_1237), .Y (n_1253));
OR2X1 g67049(.A (g2774), .B (n_1265), .Y (n_1252));
OR2X1 g66982(.A (g727), .B (n_9210), .Y (n_1251));
OR2X1 g67031(.A (g2792), .B (n_1265), .Y (n_1250));
NOR2X1 g67043(.A (g2089), .B (n_1327), .Y (n_1249));
OR2X1 g67205(.A (g2651), .B (n_1247), .Y (n_1248));
NAND2X2 g67294(.A (n_1265), .B (n_1245), .Y (n_2653));
NAND2X2 g67359(.A (n_1247), .B (g_14726), .Y (n_2925));
NOR2X1 g67034(.A (g2080), .B (n_1327), .Y (n_1244));
INVX2 g67627(.A (g7390), .Y (n_1596));
CLKBUFX1 gbuf_d_1178(.A(g6485), .Y(d_out_1178));
CLKBUFX1 gbuf_q_1178(.A(q_in_1178), .Y(g_15095));
OR2X1 g67833(.A (g2459), .B (n_9512), .Y (n_1241));
OR2X1 g67860(.A (g2444), .B (n_9512), .Y (n_1240));
OR2X1 g67906(.A (g369), .B (n_1237), .Y (n_1238));
OR2X1 g67910(.A (g1750), .B (n_1235), .Y (n_1236));
NOR2X1 g67935(.A (g_7184), .B (n_1382), .Y (n_1234));
INVX1 g67582(.A (n_8626), .Y (g7161));
INVX1 g68253(.A (n_1032), .Y (n_7686));
INVX1 g68334(.A (g6573), .Y (n_1392));
NOR2X1 g63005(.A (n_1074), .B (n_1279), .Y (n_1225));
OR2X1 g66980(.A (g715), .B (n_9210), .Y (n_1223));
CLKBUFX1 gbuf_d_1179(.A(g7052), .Y(d_out_1179));
CLKBUFX1 gbuf_q_1179(.A(q_in_1179), .Y(g_10301));
INVX1 g67238(.A (n_8623), .Y (n_1290));
NOR2X1 g63678(.A (n_1219), .B (g3036), .Y (n_1220));
OR2X1 g67218(.A (g1392), .B (n_8626), .Y (n_1218));
OR2X1 g67188(.A (g1389), .B (n_8626), .Y (n_1217));
AOI21X1 g64469(.A0 (n_1075), .A1 (n_420), .B0 (n_999), .Y (n_1214));
NOR2X1 g64639(.A (n_705), .B (n_1279), .Y (n_1213));
NOR2X1 g64650(.A (n_886), .B (n_1279), .Y (n_1212));
NOR2X1 g67932(.A (g2516), .B (g5555), .Y (n_1211));
OR2X1 g64703(.A (n_706), .B (n_1279), .Y (n_1210));
AOI22X1 g65351(.A0 (n_887), .A1 (n_1209), .B0 (g2443), .B1 (g2412),.Y (n_1370));
AOI22X1 g65122(.A0 (n_889), .A1 (n_1209), .B0 (g2458), .B1 (g2412),.Y (n_1459));
AOI21X1 g66040(.A0 (n_866), .A1 (g394), .B0 (n_688), .Y (n_1208));
AOI22X1 g65356(.A0 (n_890), .A1 (n_1209), .B0 (g2399), .B1 (g2412),.Y (n_1264));
MX2X1 g65364(.A (g2615), .B (g2612), .S0 (g3229), .Y (n_1206));
MX2X1 g65368(.A (g1921), .B (g1918), .S0 (g3229), .Y (n_1205));
NOR2X1 g66475(.A (n_8084), .B (g2607), .Y (n_1204));
OR2X1 g67099(.A (g1410), .B (n_8626), .Y (n_1203));
AOI21X1 g65578(.A0 (n_111), .A1 (g3133), .B0 (n_977), .Y (n_1202));
OAI22X1 g65751(.A0 (n_880), .A1 (g3125), .B0 (g3110), .B1 (n_1051),.Y (n_1201));
AOI22X1 g65803(.A0 (n_1195), .A1 (g3085), .B0 (n_1086), .B1 (n_185),.Y (n_1200));
AOI22X1 g65806(.A0 (n_1089), .A1 (n_1198), .B0 (n_1197), .B1(n_1193), .Y (n_1199));
AOI22X1 g65807(.A0 (g3164), .A1 (n_1195), .B0 (g3161), .B1 (n_779),.Y (n_1196));
AOI22X1 g65811(.A0 (g3176), .A1 (n_1193), .B0 (g3173), .B1 (n_982),.Y (n_1194));
INVX1 g65826(.A (n_6442), .Y (n_1192));
NOR2X1 g65834(.A (n_1185), .B (g2917), .Y (n_1191));
OR2X1 g65835(.A (g2933), .B (g51), .Y (n_1190));
NAND2X1 g65847(.A (n_1342), .B (g_8187), .Y (n_1189));
NOR2X1 g65850(.A (n_7142), .B (n_7337), .Y (n_1188));
NAND2X1 g65863(.A (n_310), .B (g3079), .Y (n_1187));
NAND2X1 g65944(.A (n_1342), .B (g_17474), .Y (n_1186));
NAND2X1 g65960(.A (n_1185), .B (g2814), .Y (n_1365));
AOI21X1 g65970(.A0 (g3126), .A1 (n_1051), .B0 (n_120), .Y (n_1184));
INVX1 g65974(.A (n_1181), .Y (n_1182));
AOI21X1 g66018(.A0 (n_862), .A1 (g_19985), .B0 (n_642), .Y (n_1180));
AOI21X1 g66036(.A0 (n_867), .A1 (g_16164), .B0 (n_646), .Y (n_1179));
AOI21X1 g66070(.A0 (g3124), .A1 (n_1051), .B0 (n_63), .Y (n_1178));
AOI21X1 g66081(.A0 (g1038), .A1 (n_404), .B0 (n_975), .Y (n_1177));
AOI21X1 g66082(.A0 (g1053), .A1 (n_404), .B0 (n_967), .Y (n_1176));
AOI21X1 g66083(.A0 (g1068), .A1 (n_404), .B0 (n_964), .Y (n_1174));
AOI21X1 g66084(.A0 (g1083), .A1 (n_404), .B0 (n_965), .Y (n_1173));
AOI22X1 g66111(.A0 (n_1171), .A1 (n_1168), .B0 (n_1170), .B1(n_1167), .Y (n_1172));
AOI22X1 g66112(.A0 (n_1168), .A1 (g3094), .B0 (n_1167), .B1 (g3093),.Y (n_1169));
AOI22X1 g66113(.A0 (g3182), .A1 (n_1168), .B0 (g3179), .B1 (n_1167),.Y (n_1166));
AOI22X1 g66115(.A0 (n_2), .A1 (n_1086), .B0 (g3167), .B1 (n_1463), .Y(n_1165));
OR2X1 g67051(.A (g1395), .B (n_8626), .Y (n_1164));
CLKBUFX1 gbuf_d_1180(.A(g_23988), .Y(d_out_1180));
CLKBUFX1 gbuf_qn_1180(.A(qn_in_1180), .Y(g_17001));
CLKBUFX1 gbuf_d_1181(.A(g451), .Y(d_out_1181));
CLKBUFX1 gbuf_qn_1181(.A(qn_in_1181), .Y(g_9014));
CLKBUFX1 gbuf_d_1182(.A(g1138), .Y(d_out_1182));
CLKBUFX1 gbuf_q_1182(.A(q_in_1182), .Y(g1215));
CLKBUFX1 gbuf_d_1183(.A(g972), .Y(d_out_1183));
CLKBUFX1 gbuf_q_1183(.A(q_in_1183), .Y(g1220));
CLKBUFX1 gbuf_d_1184(.A(g_26059), .Y(d_out_1184));
CLKBUFX1 gbuf_qn_1184(.A(qn_in_1184), .Y(g_19993));
CLKBUFX1 gbuf_d_1185(.A(g453), .Y(d_out_1185));
CLKBUFX1 gbuf_qn_1185(.A(qn_in_1185), .Y(g_11640));
NOR2X1 g66244(.A (n_8084), .B (g2604), .Y (n_1163));
NOR2X1 g66245(.A (n_7892), .B (g1914), .Y (n_1162));
NOR2X1 g66254(.A (n_7892), .B (g1913), .Y (n_1161));
NOR2X1 g66256(.A (n_7892), .B (g1911), .Y (n_1160));
NOR2X1 g66264(.A (n_8084), .B (g2608), .Y (n_1159));
AND2X1 g65860(.A (n_987), .B (n_608), .Y (n_3793));
NOR2X1 g66464(.A (n_8084), .B (g2603), .Y (n_1158));
NOR2X1 g67862(.A (g2233), .B (n_1305), .Y (n_1157));
NOR2X1 g66632(.A (n_960), .B (g_19959), .Y (n_1156));
OR2X1 g66984(.A (g1386), .B (n_8626), .Y (n_1155));
OR2X1 g67209(.A (g1398), .B (n_8626), .Y (n_1154));
NAND2X2 g67303(.A (n_1327), .B (n_562), .Y (n_2508));
INVX1 g67460(.A (n_1152), .Y (n_1331));
INVX1 g67467(.A (n_1152), .Y (n_1333));
XOR2X1 g62751(.A (g3024), .B (n_899), .Y (n_1150));
INVX4 g67629(.A (n_1247), .Y (g7390));
NOR2X1 g67834(.A (n_1145), .B (n_2014), .Y (n_1146));
NOR2X1 g67835(.A (g2239), .B (n_1305), .Y (n_1144));
NOR2X1 g67841(.A (g2507), .B (g5555), .Y (n_1143));
NOR2X1 g67848(.A (n_1141), .B (n_2170), .Y (n_1142));
INVX1 g67853(.A (n_1084), .Y (n_1140));
INVX1 g67866(.A (n_1036), .Y (n_1138));
NOR2X1 g67868(.A (n_1136), .B (n_864), .Y (n_1137));
NOR2X1 g67869(.A (g411), .B (n_6914), .Y (n_1135));
INVX1 g67879(.A (n_1006), .Y (n_1134));
OR2X1 g67883(.A (g_25781), .B (n_1122), .Y (n_1133));
NOR2X1 g67889(.A (n_1131), .B (n_864), .Y (n_1132));
NOR2X1 g67895(.A (g2230), .B (n_1305), .Y (n_1129));
INVX1 g67898(.A (n_1033), .Y (n_1127));
NOR2X1 g67902(.A (n_1125), .B (n_2014), .Y (n_1126));
OR2X1 g67913(.A (g_14751), .B (n_1122), .Y (n_1123));
INVX1 g67920(.A (n_1026), .Y (n_1121));
NOR2X1 g67923(.A (g2486), .B (g5555), .Y (n_1120));
NOR2X1 g67925(.A (g432), .B (n_6914), .Y (n_1118));
INVX1 g67929(.A (n_1025), .Y (n_1117));
NOR2X1 g67931(.A (g1813), .B (g5511), .Y (n_1116));
NOR2X1 g67944(.A (n_1114), .B (n_2014), .Y (n_1115));
NOR2X1 g67973(.A (n_1112), .B (n_2170), .Y (n_1113));
OR2X1 g67979(.A (g_5844), .B (n_1122), .Y (n_1109));
NOR2X1 g67981(.A (g_15404), .B (n_1122), .Y (n_1108));
NOR2X1 g67983(.A (g_27738), .B (n_9395), .Y (n_1107));
INVX1 g67989(.A (n_1019), .Y (n_1105));
NOR2X1 g68002(.A (g441), .B (n_6914), .Y (n_1104));
NOR2X1 g68005(.A (n_1101), .B (n_2170), .Y (n_1102));
NOR2X1 g68018(.A (g1822), .B (g5511), .Y (n_1100));
NOR2X1 g68021(.A (g1792), .B (g5511), .Y (n_1099));
INVX1 g68056(.A (n_1014), .Y (n_9699));
OR2X1 g67018(.A (g1407), .B (n_8626), .Y (n_1095));
INVX1 g68337(.A (n_1285), .Y (g6573));
NOR2X1 g67914(.A (n_1093), .B (n_864), .Y (n_1094));
NOR2X1 g67905(.A (g2227), .B (n_1305), .Y (n_1092));
AOI22X1 g65812(.A0 (n_1089), .A1 (g3096), .B0 (n_1193), .B1 (g3092),.Y (n_1090));
OR2X1 g66970(.A (g1401), .B (n_8626), .Y (n_1088));
AOI22X1 g65801(.A0 (g3100), .A1 (n_1195), .B0 (n_88), .B1 (n_1086),.Y (n_1087));
OR2X1 g66952(.A (g1419), .B (n_8626), .Y (n_1085));
NOR2X1 g67854(.A (n_104), .B (n_901), .Y (n_1084));
OR2X1 g67842(.A (g818), .B (n_1032), .Y (n_1083));
CLKBUFX1 gbuf_d_1186(.A(g970), .Y(d_out_1186));
CLKBUFX1 gbuf_q_1186(.A(q_in_1186), .Y(g1219));
XOR2X1 g65373(.A (n_785), .B (n_786), .Y (n_1379));
AOI21X1 g66103(.A0 (g3114), .A1 (n_1053), .B0 (n_883), .Y (n_1082));
INVX1 g68338(.A (n_1077), .Y (n_1285));
AOI21X1 g66078(.A0 (g1747), .A1 (g_32166), .B0 (n_872), .Y (n_1079));
CLKBUFX1 gbuf_d_1187(.A(gbuf79), .Y(d_out_1187));
CLKBUFX1 gbuf_qn_1187(.A(qn_in_1187), .Y(g966));
XOR2X1 g64519(.A (n_268), .B (n_1075), .Y (n_1076));
XOR2X1 g64529(.A (g3010), .B (n_732), .Y (n_1074));
OR2X1 g67922(.A (g1085), .B (n_8305), .Y (n_1073));
XOR2X1 g65371(.A (n_787), .B (n_788), .Y (n_1377));
CLKBUFX1 gbuf_d_1188(.A(n_885), .Y(d_out_1188));
CLKBUFX1 gbuf_q_1188(.A(q_in_1188), .Y(g_22696));
CLKBUFX1 gbuf_d_1189(.A(n_884), .Y(d_out_1189));
CLKBUFX1 gbuf_q_1189(.A(q_in_1189), .Y(g1224));
NAND2X1 g65408(.A (n_1069), .B (g3018), .Y (n_1219));
NAND2X1 g65495(.A (n_888), .B (n_1209), .Y (n_1070));
NAND3X1 g65534(.A (n_1069), .B (g3018), .C (g3028), .Y (n_1453));
NAND2X1 g65572(.A (g1905), .B (g1918), .Y (n_1068));
AOI21X1 g65602(.A0 (n_781), .A1 (g3211), .B0 (g3084), .Y (n_1067));
NAND2X1 g65613(.A (g2612), .B (g2599), .Y (n_1066));
AOI22X1 g65804(.A0 (g3158), .A1 (n_781), .B0 (g3155), .B1 (n_1063),.Y (n_1065));
AOI22X1 g65808(.A0 (n_1061), .A1 (g3147), .B0 (n_1063), .B1 (g3097),.Y (n_1064));
AOI22X1 g65809(.A0 (n_1061), .A1 (n_296), .B0 (n_1063), .B1 (g3210),.Y (n_1062));
NAND2X1 g65825(.A (n_1089), .B (g3088), .Y (n_1060));
NAND2X1 g65827(.A (n_1342), .B (n_7337), .Y (n_6442));
OR2X1 g65853(.A (n_882), .B (n_7190), .Y (n_7558));
OR2X1 g65861(.A (n_7992), .B (n_6440), .Y (n_8054));
NAND3X1 g65975(.A (n_1001), .B (g2917), .C (g2912), .Y (n_1181));
CLKBUFX1 gbuf_d_1190(.A(g_11049), .Y(d_out_1190));
CLKBUFX1 gbuf_qn_1190(.A(qn_in_1190), .Y(g_11807));
NAND2X1 g67870(.A (g849), .B (n_2597), .Y (n_1059));
AOI21X1 g66019(.A0 (g1732), .A1 (g_32166), .B0 (n_874), .Y (n_1058));
AOI21X1 g66025(.A0 (g1762), .A1 (g_32166), .B0 (n_873), .Y (n_1057));
AOI21X1 g66069(.A0 (g1777), .A1 (g_32166), .B0 (n_870), .Y (n_1056));
INVX1 g66093(.A (n_1055), .Y (n_5663));
CLKBUFX1 gbuf_d_1191(.A(g974), .Y(d_out_1191));
CLKBUFX1 gbuf_qn_1191(.A(qn_in_1191), .Y(g1222));
AOI22X1 g66114(.A0 (n_24), .A1 (n_1051), .B0 (n_35), .B1 (n_1053), .Y(n_1054));
AOI22X1 g66116(.A0 (n_62), .A1 (n_1051), .B0 (g3120), .B1 (n_1053),.Y (n_1052));
CLKBUFX1 gbuf_d_1192(.A(g968), .Y(d_out_1192));
CLKBUFX1 gbuf_q_1192(.A(q_in_1192), .Y(g1218));
CLKBUFX1 gbuf_d_1193(.A(g1140), .Y(d_out_1193));
CLKBUFX1 gbuf_q_1193(.A(q_in_1193), .Y(g1216));
CLKBUFX1 gbuf_d_1194(.A(g976), .Y(d_out_1194));
CLKBUFX1 gbuf_qn_1194(.A(qn_in_1194), .Y(g1223));
NOR2X1 g66250(.A (n_8084), .B (g2605), .Y (n_1049));
NOR2X1 g66309(.A (n_7892), .B (g1910), .Y (n_1048));
NOR2X1 g66310(.A (n_7892), .B (g1912), .Y (n_1047));
NOR2X1 g66311(.A (n_1053), .B (n_1051), .Y (n_1655));
NAND2X1 g66314(.A (g485), .B (n_336), .Y (n_1046));
NOR2X1 g66435(.A (n_8084), .B (g2606), .Y (n_1044));
NAND2X1 g66456(.A (g2560), .B (n_342), .Y (n_1043));
NAND2X1 g66568(.A (n_863), .B (g2987), .Y (g16496));
NOR2X1 g66594(.A (g1011), .B (g1024), .Y (n_1041));
NOR2X1 g66624(.A (n_865), .B (g1951), .Y (n_1040));
OAI21X1 g66942(.A0 (g2245), .A1 (n_8934), .B0 (g2246), .Y (n_1039));
INVX1 g67937(.A (n_950), .Y (n_9692));
INVX2 g67630(.A (g_17921), .Y (n_1247));
INVX1 g67677(.A (n_1327), .Y (g7357));
INVX2 g67748(.A (g_5793), .Y (n_1265));
NOR2X1 g67867(.A (n_247), .B (n_1024), .Y (n_1036));
OR2X1 g67878(.A (g_29016), .B (n_9395), .Y (n_8206));
INVX1 g67891(.A (n_952), .Y (n_1034));
NOR2X1 g67899(.A (g821), .B (n_1032), .Y (n_1033));
OR2X1 g67903(.A (g1536), .B (n_853), .Y (n_1031));
OR2X1 g67904(.A (g_20789), .B (n_9395), .Y (n_1030));
OR2X1 g67917(.A (g1542), .B (n_853), .Y (n_1028));
NOR2X1 g67921(.A (g_26130), .B (n_9395), .Y (n_1026));
NOR2X1 g67930(.A (n_251), .B (n_1024), .Y (n_1025));
NOR2X1 g67959(.A (g1524), .B (n_853), .Y (n_1023));
OR2X1 g67960(.A (g1533), .B (n_853), .Y (n_1022));
INVX1 g67961(.A (n_946), .Y (n_1021));
INVX1 g67986(.A (n_944), .Y (n_1020));
NOR2X1 g67990(.A (g833), .B (n_1032), .Y (n_1019));
OR2X1 g68003(.A (g1539), .B (n_853), .Y (n_8278));
OR2X1 g68008(.A (g1545), .B (n_853), .Y (n_1017));
INVX1 g68029(.A (n_938), .Y (n_1016));
OR2X1 g68039(.A (g836), .B (n_2597), .Y (n_1015));
NOR2X1 g68057(.A (n_278), .B (n_901), .Y (n_1014));
INVX1 g68060(.A (n_930), .Y (n_1013));
INVX1 g68257(.A (n_1032), .Y (g6368));
BUFX3 g68394(.A (n_9395), .Y (n_1382));
AOI21X1 g65546(.A0 (g3099), .A1 (n_779), .B0 (g3098), .Y (n_1008));
INVX1 g68471(.A (n_1305), .Y (g6837));
NAND2X1 g66359(.A (g1866), .B (n_389), .Y (n_1007));
NOR2X1 g67880(.A (g_24187), .B (n_1024), .Y (n_1006));
INVX1 g67469(.A (n_9209), .Y (n_1152));
NOR2X1 g66576(.A (g1055), .B (g1024), .Y (n_1004));
NOR2X1 g66573(.A (g1070), .B (g1024), .Y (n_1003));
CLKBUFX1 gbuf_d_1195(.A(g1660), .Y(d_out_1195));
CLKBUFX1 gbuf_q_1195(.A(q_in_1195), .Y(g1911));
CLKBUFX1 gbuf_d_1196(.A(gbuf30), .Y(d_out_1196));
CLKBUFX1 gbuf_qn_1196(.A(qn_in_1196), .Y(g_26059));
CLKBUFX1 gbuf_d_1197(.A(g1664), .Y(d_out_1197));
CLKBUFX1 gbuf_q_1197(.A(q_in_1197), .Y(g1913));
CLKBUFX1 gbuf_d_1198(.A(g2360), .Y(d_out_1198));
CLKBUFX1 gbuf_q_1198(.A(q_in_1198), .Y(g2608));
CLKBUFX1 gbuf_d_1199(.A(g1670), .Y(d_out_1199));
CLKBUFX1 gbuf_qn_1199(.A(qn_in_1199), .Y(g1917));
INVX1 g66537(.A (n_1001), .Y (n_1185));
CLKBUFX1 gbuf_d_1200(.A(gbuf82), .Y(d_out_1200));
CLKBUFX1 gbuf_qn_1200(.A(qn_in_1200), .Y(g972));
CLKBUFX1 gbuf_d_1201(.A(gbuf29), .Y(d_out_1201));
CLKBUFX1 gbuf_qn_1201(.A(qn_in_1201), .Y(g453));
CLKBUFX1 gbuf_d_1202(.A(gbuf28), .Y(d_out_1202));
CLKBUFX1 gbuf_qn_1202(.A(qn_in_1202), .Y(g451));
CLKBUFX1 gbuf_d_1203(.A(g2358), .Y(d_out_1203));
CLKBUFX1 gbuf_q_1203(.A(q_in_1203), .Y(g2607));
CLKBUFX1 gbuf_d_1204(.A(n_816), .Y(d_out_1204));
CLKBUFX1 gbuf_qn_1204(.A(qn_in_1204), .Y(g3079));
CLKBUFX1 gbuf_d_1205(.A(gbuf35), .Y(d_out_1205));
CLKBUFX1 gbuf_qn_1205(.A(qn_in_1205), .Y(g_23988));
NOR2X1 g64707(.A (n_419), .B (n_1075), .Y (n_999));
NOR2X1 g66233(.A (n_8084), .B (n_905), .Y (n_998));
CLKBUFX1 gbuf_d_1206(.A(g2528), .Y(d_out_1206));
CLKBUFX1 gbuf_q_1206(.A(q_in_1206), .Y(g2604));
CLKBUFX1 gbuf_d_1207(.A(g7425), .Y(d_out_1207));
CLKBUFX1 gbuf_q_1207(.A(q_in_1207), .Y(g_5793));
NAND2X1 g65409(.A (n_891), .B (n_310), .Y (n_1279));
OR2X1 g67901(.A (g2221), .B (n_8934), .Y (n_9667));
CLKBUFX1 gbuf_d_1208(.A(gbuf77), .Y(d_out_1208));
CLKBUFX1 gbuf_qn_1208(.A(qn_in_1208), .Y(g1138));
NAND4X1 g65548(.A (n_776), .B (n_465), .C (g793), .D (n_763), .Y(n_4464));
AND2X1 g66192(.A (n_3873), .B (n_986), .Y (n_987));
NAND2X1 g66185(.A (g3133), .B (n_868), .Y (n_985));
AOI22X1 g65805(.A0 (g3170), .A1 (n_981), .B0 (g3185), .B1 (n_2188),.Y (n_984));
AOI22X1 g65810(.A0 (n_982), .A1 (g3091), .B0 (n_981), .B1 (g3087), .Y(n_983));
INVX4 g67678(.A (g_21556), .Y (n_1327));
NAND2X1 g65824(.A (n_1061), .B (g3151), .Y (n_980));
CLKBUFX1 gbuf_d_1209(.A(n_805), .Y(d_out_1209));
CLKBUFX1 gbuf_q_1209(.A(q_in_1209), .Y(g2879));
NOR2X1 g67975(.A (g1801), .B (g5511), .Y (n_978));
AOI21X1 g66053(.A0 (g3139), .A1 (n_1086), .B0 (n_1051), .Y (n_977));
NOR2X1 g66094(.A (n_735), .B (n_647), .Y (n_1055));
XOR2X1 g66101(.A (n_782), .B (n_518), .Y (n_976));
NOR2X1 g66633(.A (n_772), .B (g1036), .Y (n_975));
CLKBUFX1 gbuf_d_1210(.A(n_774), .Y(d_out_1210));
CLKBUFX1 gbuf_q_1210(.A(q_in_1210), .Y(g2933));
CLKBUFX1 gbuf_d_1211(.A(g_25350), .Y(d_out_1211));
CLKBUFX1 gbuf_qn_1211(.A(qn_in_1211), .Y(g_17474));
CLKBUFX1 gbuf_d_1212(.A(g_22901), .Y(d_out_1212));
CLKBUFX1 gbuf_qn_1212(.A(qn_in_1212), .Y(g_17483));
CLKBUFX1 gbuf_d_1213(.A(g_25247), .Y(d_out_1213));
CLKBUFX1 gbuf_qn_1213(.A(qn_in_1213), .Y(g_8187));
NOR2X1 g66281(.A (n_7892), .B (g1909), .Y (n_973));
NAND2X1 g67956(.A (n_971), .B (n_935), .Y (n_972));
INVX1 g66198(.A (n_970), .Y (n_6328));
AOI21X1 g66554(.A0 (n_903), .A1 (n_802), .B0 (n_699), .Y (n_969));
NOR2X1 g66619(.A (n_773), .B (g1051), .Y (n_967));
NOR2X1 g66626(.A (n_769), .B (g571), .Y (n_966));
NOR2X1 g66627(.A (n_771), .B (g1081), .Y (n_965));
NOR2X1 g66634(.A (n_770), .B (g1066), .Y (n_964));
NOR2X1 g66636(.A (n_766), .B (g1257), .Y (n_963));
CLKBUFX1 gbuf_d_1214(.A(g2364), .Y(d_out_1214));
CLKBUFX1 gbuf_qn_1214(.A(qn_in_1214), .Y(g2611));
CLKBUFX1 gbuf_d_1215(.A(g2526), .Y(d_out_1215));
CLKBUFX1 gbuf_q_1215(.A(q_in_1215), .Y(g2603));
CLKBUFX1 gbuf_d_1216(.A(g1666), .Y(d_out_1216));
CLKBUFX1 gbuf_q_1216(.A(q_in_1216), .Y(g1914));
NOR2X1 g67291(.A (g_9473), .B (n_761), .Y (n_960));
NAND2X1 g67292(.A (n_761), .B (g_24889), .Y (n_1447));
CLKBUFX1 gbuf_d_1217(.A(g7302), .Y(d_out_1217));
CLKBUFX1 gbuf_q_1217(.A(q_in_1217), .Y(g_17921));
NOR2X1 g67838(.A (g1970), .B (g7052), .Y (n_956));
OR2X1 g67851(.A (g1071), .B (n_8305), .Y (n_955));
INVX1 g67874(.A (n_854), .Y (n_953));
NOR2X1 g67892(.A (g1527), .B (n_840), .Y (n_952));
NOR2X1 g67897(.A (g420), .B (n_6914), .Y (n_951));
NOR2X1 g67938(.A (g2206), .B (n_8934), .Y (n_950));
INVX1 g67939(.A (n_857), .Y (n_949));
NOR2X1 g67962(.A (g1530), .B (n_840), .Y (n_946));
NOR2X1 g67987(.A (g1551), .B (n_840), .Y (n_944));
NAND2X1 g67998(.A (n_942), .B (n_8643), .Y (n_943));
NOR2X1 g68014(.A (g2224), .B (n_8934), .Y (n_941));
INVX1 g68024(.A (n_833), .Y (n_940));
OR2X1 g68028(.A (g1056), .B (n_8305), .Y (n_939));
NOR2X1 g68030(.A (g1512), .B (n_840), .Y (n_938));
NAND2X1 g68032(.A (n_936), .B (n_935), .Y (n_937));
NAND2X1 g68033(.A (n_933), .B (n_748), .Y (n_934));
NAND2X1 g68058(.A (g2704), .B (g7425), .Y (n_4300));
NOR2X1 g68061(.A (g2209), .B (n_8934), .Y (n_930));
INVX1 g68340(.A (n_853), .Y (n_1077));
CLKBUFX3 g68397(.A (n_1024), .Y (n_1122));
OR2X1 g68034(.A (g2218), .B (n_8934), .Y (n_923));
NOR2X1 g67915(.A (g1276), .B (g6750), .Y (n_922));
INVX1 g67006(.A (n_4088), .Y (n_920));
INVX4 g68472(.A (n_8935), .Y (n_1305));
NAND2X1 g67863(.A (n_917), .B (n_935), .Y (n_918));
NAND2X1 g66586(.A (g1734), .B (g1718), .Y (n_913));
AOI22X1 g65802(.A0 (n_911), .A1 (n_982), .B0 (g3102), .B1 (n_981), .Y(n_912));
NOR2X1 g67864(.A (g2495), .B (g5555), .Y (n_910));
CLKBUFX1 gbuf_d_1218(.A(gbuf83), .Y(d_out_1218));
CLKBUFX1 gbuf_qn_1218(.A(qn_in_1218), .Y(g974));
NOR2X1 g67839(.A (g_19787), .B (n_9393), .Y (n_909));
NAND2X1 g67836(.A (g2679), .B (n_6822), .Y (n_908));
CLKBUFX1 gbuf_d_1219(.A(g1662), .Y(d_out_1219));
CLKBUFX1 gbuf_q_1219(.A(q_in_1219), .Y(g1912));
CLKBUFX1 gbuf_d_1220(.A(gbuf80), .Y(d_out_1220));
CLKBUFX1 gbuf_qn_1220(.A(qn_in_1220), .Y(g968));
CLKBUFX1 gbuf_d_1221(.A(g2362), .Y(d_out_1221));
CLKBUFX1 gbuf_qn_1221(.A(qn_in_1221), .Y(g2610));
CLKBUFX1 gbuf_d_1222(.A(g2354), .Y(d_out_1222));
CLKBUFX1 gbuf_q_1222(.A(q_in_1222), .Y(g2605));
INVX1 g65506(.A (n_6947), .Y (n_6946));
CLKBUFX1 gbuf_d_1223(.A(g1834), .Y(d_out_1223));
CLKBUFX1 gbuf_q_1223(.A(q_in_1223), .Y(g1910));
CLKBUFX1 gbuf_d_1224(.A(g5686), .Y(d_out_1224));
CLKBUFX1 gbuf_qn_1224(.A(qn_in_1224), .Y(g1024));
AND2X1 g67968(.A (g2398), .B (n_9510), .Y (n_904));
NOR2X1 g67182(.A (n_803), .B (n_903), .Y (n_1168));
NOR2X1 g66538(.A (n_677), .B (n_487), .Y (n_1001));
NAND2X1 g66284(.A (n_701), .B (g3161), .Y (n_902));
CLKBUFX1 gbuf_d_1225(.A(g8082), .Y(d_out_1225));
CLKBUFX1 gbuf_qn_1225(.A(qn_in_1225), .Y(g1866));
CLKBUFX1 gbuf_d_1226(.A(g2356), .Y(d_out_1226));
CLKBUFX1 gbuf_q_1226(.A(q_in_1226), .Y(g2606));
INVX2 g68262(.A (n_900), .Y (n_2597));
CLKBUFX1 gbuf_d_1227(.A(gbuf78), .Y(d_out_1227));
CLKBUFX1 gbuf_qn_1227(.A(qn_in_1227), .Y(g1140));
INVX1 g68261(.A (n_900), .Y (n_901));
CLKBUFX1 gbuf_d_1228(.A(g8007), .Y(d_out_1228));
CLKBUFX1 gbuf_q_1228(.A(q_in_1228), .Y(g1172));
NAND2X1 g64638(.A (n_731), .B (g3010), .Y (n_899));
OR2X1 g66199(.A (n_8084), .B (n_8103), .Y (n_970));
CLKBUFX1 gbuf_d_1229(.A(g8167), .Y(d_out_1229));
CLKBUFX1 gbuf_qn_1229(.A(qn_in_1229), .Y(g2560));
AND2X1 g66489(.A (n_877), .B (n_710), .Y (n_1193));
CLKBUFX1 gbuf_d_1230(.A(n_496), .Y(d_out_1230));
CLKBUFX1 gbuf_q_1230(.A(q_in_1230), .Y(gbuf79));
CLKBUFX1 gbuf_d_1231(.A(gbuf84), .Y(d_out_1231));
CLKBUFX1 gbuf_qn_1231(.A(qn_in_1231), .Y(g976));
INVX1 g68172(.A (g5511), .Y (n_1235));
CLKBUFX1 gbuf_d_1232(.A(n_723), .Y(d_out_1232));
CLKBUFX1 gbuf_q_1232(.A(q_in_1232), .Y(g1918));
CLKBUFX1 gbuf_d_1233(.A(n_703), .Y(d_out_1233));
CLKBUFX1 gbuf_q_1233(.A(q_in_1233), .Y(g2612));
INVX1 g67876(.A (n_790), .Y (n_894));
CLKBUFX1 gbuf_d_1234(.A(gbuf33), .Y(d_out_1234));
CLKBUFX1 gbuf_qn_1234(.A(qn_in_1234), .Y(g_11049));
NAND2X1 g65929(.A (n_893), .B (n_892), .Y (n_1464));
INVX1 g65931(.A (n_891), .Y (n_1069));
AOI21X1 g66010(.A0 (n_651), .A1 (g2469), .B0 (n_667), .Y (n_890));
AOI21X1 g66017(.A0 (n_650), .A1 (g2454), .B0 (n_649), .Y (n_889));
INVX4 g68259(.A (n_900), .Y (n_1032));
AOI21X1 g66089(.A0 (n_648), .A1 (g2424), .B0 (n_609), .Y (n_888));
AOI21X1 g66090(.A0 (n_665), .A1 (g2439), .B0 (n_617), .Y (n_887));
XOR2X1 g66129(.A (g3013), .B (n_652), .Y (n_886));
MX2X1 g66130(.A (g_20059), .B (g_31512), .S0 (g3229), .Y (n_885));
MX2X1 g66131(.A (g992), .B (g978), .S0 (g3229), .Y (n_884));
NOR2X1 g66186(.A (n_34), .B (n_801), .Y (n_883));
OR2X1 g66196(.A (n_7892), .B (n_7992), .Y (n_6440));
OR2X1 g66200(.A (n_7462), .B (n_882), .Y (n_7190));
NAND2X1 g66208(.A (n_701), .B (g3087), .Y (n_881));
AND2X1 g66235(.A (g3110), .B (n_1053), .Y (n_880));
NAND2X1 g66266(.A (n_701), .B (g3084), .Y (n_879));
NOR2X1 g66278(.A (n_1053), .B (g3126), .Y (n_878));
AND2X1 g66336(.A (n_619), .B (n_877), .Y (n_1089));
NOR2X1 g66348(.A (n_2187), .B (n_479), .Y (n_876));
AND2X1 g66463(.A (n_877), .B (n_712), .Y (n_1195));
NOR2X1 g66490(.A (g3124), .B (n_1053), .Y (n_875));
INVX1 g66616(.A (n_7142), .Y (n_1342));
NOR2X1 g66620(.A (n_690), .B (g1730), .Y (n_874));
NOR2X1 g66623(.A (n_693), .B (g1760), .Y (n_873));
NOR2X1 g66631(.A (n_692), .B (g1745), .Y (n_872));
NOR2X1 g66637(.A (n_689), .B (g2645), .Y (n_871));
NOR2X1 g66638(.A (n_691), .B (g1775), .Y (n_870));
CLKBUFX1 gbuf_d_1235(.A(g7956), .Y(d_out_1235));
CLKBUFX1 gbuf_qn_1235(.A(qn_in_1235), .Y(g485));
CLKBUFX1 gbuf_d_1236(.A(g5648), .Y(d_out_1236));
CLKBUFX1 gbuf_q_1236(.A(q_in_1236), .Y(g_28034));
CLKBUFX1 gbuf_d_1237(.A(gbuf81), .Y(d_out_1237));
CLKBUFX1 gbuf_qn_1237(.A(qn_in_1237), .Y(g970));
NAND2X1 g67240(.A (g_18059), .B (g5648), .Y (n_867));
OR2X1 g67265(.A (g5686), .B (g5657), .Y (n_1446));
NAND2X1 g67304(.A (g396), .B (g5648), .Y (n_866));
NOR2X1 g67306(.A (g1949), .B (n_864), .Y (n_865));
NAND2X1 g67319(.A (g2986), .B (g5388), .Y (n_863));
NAND2X1 g67320(.A (g_27919), .B (g5648), .Y (n_862));
NOR2X1 g67940(.A (n_61), .B (n_853), .Y (n_857));
CLKBUFX1 gbuf_d_1238(.A(g6677), .Y(d_out_1238));
CLKBUFX1 gbuf_q_1238(.A(q_in_1238), .Y(g_21387));
CLKBUFX1 gbuf_d_1239(.A(g7229), .Y(d_out_1239));
CLKBUFX1 gbuf_q_1239(.A(q_in_1239), .Y(g_21556));
AND2X1 g67840(.A (g1704), .B (n_755), .Y (n_856));
NOR2X1 g67875(.A (g1515), .B (n_853), .Y (n_854));
AND2X1 g67884(.A (g2479), .B (n_9510), .Y (n_852));
NAND2X1 g67885(.A (g2688), .B (n_6822), .Y (n_850));
NAND2X1 g67888(.A (g2010), .B (g7229), .Y (n_3689));
NAND2X1 g67909(.A (g1316), .B (g6979), .Y (n_3303));
NOR2X1 g67912(.A (n_845), .B (n_6822), .Y (n_846));
NAND2X1 g67969(.A (n_843), .B (n_840), .Y (n_844));
NAND2X1 g67970(.A (n_841), .B (n_840), .Y (n_842));
NAND2X1 g67995(.A (g1700), .B (n_755), .Y (n_839));
NOR2X1 g68000(.A (n_836), .B (n_6822), .Y (n_837));
NAND2X1 g68010(.A (n_834), .B (n_2308), .Y (n_835));
NAND2X1 g68016(.A (g630), .B (g6677), .Y (n_3552));
NOR2X1 g68025(.A (n_211), .B (n_853), .Y (n_833));
CLKBUFX1 gbuf_d_1240(.A(g6979), .Y(d_out_1240));
CLKBUFX1 gbuf_q_1240(.A(q_in_1240), .Y(g_9980));
INVX1 g68042(.A (n_747), .Y (n_832));
NAND2X1 g68046(.A (n_830), .B (n_840), .Y (n_831));
INVX1 g68363(.A (n_6914), .Y (n_1237));
INVX2 g68398(.A (n_9394), .Y (n_1024));
INVX1 g67008(.A (n_3873), .Y (n_4088));
AND2X1 g67911(.A (g1785), .B (n_755), .Y (n_821));
NOR2X1 g67893(.A (n_819), .B (n_6822), .Y (n_820));
NAND2X1 g67872(.A (g2394), .B (n_9510), .Y (n_818));
CLKBUFX1 gbuf_d_1241(.A(n_639), .Y(d_out_1241));
CLKBUFX1 gbuf_q_1241(.A(q_in_1241), .Y(g1471));
CLKBUFX1 gbuf_d_1242(.A(n_638), .Y(d_out_1242));
CLKBUFX1 gbuf_q_1242(.A(q_in_1242), .Y(g2195));
NOR2X1 g67219(.A (g3054), .B (g3234), .Y (n_816));
CLKBUFX1 gbuf_d_1243(.A(n_671), .Y(d_out_1243));
CLKBUFX1 gbuf_q_1243(.A(q_in_1243), .Y(g2165));
NOR2X1 g68052(.A (g2251), .B (n_810), .Y (n_814));
CLKBUFX1 gbuf_d_1244(.A(gbuf179), .Y(d_out_1244));
CLKBUFX1 gbuf_qn_1244(.A(qn_in_1244), .Y(g2358));
CLKBUFX1 gbuf_d_1245(.A(g5738), .Y(d_out_1245));
CLKBUFX1 gbuf_q_1245(.A(q_in_1245), .Y(g1718));
NAND2X1 g67980(.A (n_811), .B (n_810), .Y (n_812));
OR2X1 g67971(.A (g1090), .B (n_8305), .Y (n_809));
CLKBUFX1 gbuf_d_1246(.A(g1668), .Y(d_out_1246));
CLKBUFX1 gbuf_qn_1246(.A(qn_in_1246), .Y(g1916));
INVX1 g67195(.A (n_1086), .Y (n_868));
CLKBUFX1 gbuf_d_1247(.A(n_466), .Y(d_out_1247));
CLKBUFX1 gbuf_q_1247(.A(q_in_1247), .Y(gbuf30));
NAND2X1 g67882(.A (n_806), .B (n_810), .Y (n_807));
NAND2X1 g66543(.A (n_613), .B (g2879), .Y (n_805));
CLKBUFX1 gbuf_d_1248(.A(gbuf180), .Y(d_out_1248));
CLKBUFX1 gbuf_qn_1248(.A(qn_in_1248), .Y(g2360));
CLKBUFX1 gbuf_d_1249(.A(gbuf32), .Y(d_out_1249));
CLKBUFX1 gbuf_qn_1249(.A(qn_in_1249), .Y(g_25247));
CLKBUFX1 gbuf_d_1250(.A(gbuf34), .Y(d_out_1250));
CLKBUFX1 gbuf_qn_1250(.A(qn_in_1250), .Y(g_22901));
CLKBUFX1 gbuf_d_1251(.A(gbuf133), .Y(d_out_1251));
CLKBUFX1 gbuf_qn_1251(.A(qn_in_1251), .Y(g1670));
CLKBUFX1 gbuf_d_1252(.A(n_672), .Y(d_out_1252));
CLKBUFX1 gbuf_q_1252(.A(q_in_1252), .Y(g1486));
NOR2X1 g67156(.A (n_803), .B (n_802), .Y (n_1167));
INVX1 g67152(.A (n_801), .Y (n_1051));
CLKBUFX1 gbuf_d_1253(.A(gbuf31), .Y(d_out_1253));
CLKBUFX1 gbuf_qn_1253(.A(qn_in_1253), .Y(g_25350));
AND2X1 g67924(.A (n_799), .B (n_810), .Y (n_800));
CLKBUFX1 gbuf_d_1254(.A(n_467), .Y(d_out_1254));
CLKBUFX1 gbuf_q_1254(.A(q_in_1254), .Y(gbuf28));
CLKBUFX1 gbuf_d_1255(.A(gbuf175), .Y(d_out_1255));
CLKBUFX1 gbuf_qn_1255(.A(qn_in_1255), .Y(g2526));
CLKBUFX1 gbuf_d_1256(.A(n_634), .Y(d_out_1256));
CLKBUFX1 gbuf_q_1256(.A(q_in_1256), .Y(n_482));
CLKBUFX3 g68263(.A (n_742), .Y (n_900));
NAND2X1 g67974(.A (g313), .B (n_753), .Y (n_798));
NAND2X1 g68001(.A (n_796), .B (n_810), .Y (n_797));
CLKBUFX1 gbuf_d_1257(.A(n_3161), .Y(d_out_1257));
CLKBUFX1 gbuf_q_1257(.A(q_in_1257), .Y(gbuf29));
NAND4X1 g65507(.A (n_789), .B (g3018), .C (n_9), .D (n_375), .Y(n_6947));
AOI21X1 g65532(.A0 (n_478), .A1 (n_679), .B0 (n_517), .Y (n_794));
AOI21X1 g65533(.A0 (n_542), .A1 (g3006), .B0 (g3002), .Y (n_793));
NAND2X1 g67988(.A (g2388), .B (n_9510), .Y (n_792));
NOR2X1 g67877(.A (g2248), .B (n_810), .Y (n_790));
NAND2X1 g65932(.A (n_789), .B (g3080), .Y (n_891));
XOR2X1 g66125(.A (n_553), .B (n_584), .Y (n_788));
XOR2X1 g66126(.A (n_552), .B (n_549), .Y (n_787));
XOR2X1 g66127(.A (n_585), .B (n_551), .Y (n_786));
XOR2X1 g66128(.A (n_550), .B (n_548), .Y (n_785));
CLKBUFX1 gbuf_d_1258(.A(g978), .Y(d_out_1258));
CLKBUFX1 gbuf_q_1258(.A(q_in_1258), .Y(g1227));
CLKBUFX1 gbuf_d_1259(.A(g_31512), .Y(d_out_1259));
CLKBUFX1 gbuf_q_1259(.A(q_in_1259), .Y(g_16317));
NAND2X1 g66184(.A (n_783), .B (n_782), .Y (n_1075));
CLKBUFX1 gbuf_d_1260(.A(n_3171), .Y(d_out_1260));
CLKBUFX1 gbuf_q_1260(.A(q_in_1260), .Y(gbuf82));
INVX1 g66322(.A (n_893), .Y (n_781));
INVX1 g66431(.A (n_892), .Y (n_779));
NAND2X1 g66504(.A (g2428), .B (g2412), .Y (n_777));
NOR2X1 g66526(.A (n_630), .B (n_657), .Y (n_776));
INVX1 g66548(.A (n_775), .Y (n_4861));
CLKBUFX1 gbuf_d_1261(.A(n_661), .Y(d_out_1261));
CLKBUFX1 gbuf_q_1261(.A(q_in_1261), .Y(g1481));
INVX1 g66629(.A (n_704), .Y (n_1061));
INVX1 g67393(.A (n_882), .Y (n_896));
CLKBUFX1 gbuf_d_1262(.A(g1832), .Y(d_out_1262));
CLKBUFX1 gbuf_q_1262(.A(q_in_1262), .Y(g1909));
AOI21X1 g66618(.A0 (g557), .A1 (n_321), .B0 (n_767), .Y (n_7142));
NOR2X1 g67111(.A (g2817), .B (g51), .Y (n_774));
AND2X1 g67263(.A (n_734), .B (n_636), .Y (n_3390));
NOR2X1 g67266(.A (g1053), .B (g_25914), .Y (n_773));
NOR2X1 g67288(.A (g1038), .B (g_25914), .Y (n_772));
NOR2X1 g67290(.A (g1083), .B (g_25914), .Y (n_771));
NOR2X1 g67296(.A (g1068), .B (g_25914), .Y (n_770));
NOR2X1 g67297(.A (g569), .B (n_2170), .Y (n_769));
AOI21X1 g66612(.A0 (n_77), .A1 (n_3701), .B0 (n_767), .Y (n_7337));
NOR2X1 g67370(.A (g1255), .B (n_2014), .Y (n_766));
INVX1 g67382(.A (n_8103), .Y (n_905));
NAND4X1 g67396(.A (n_763), .B (n_496), .C (g801), .D (n_762), .Y(n_2811));
CLKBUFX1 gbuf_d_1263(.A(gbuf128), .Y(d_out_1263));
CLKBUFX1 gbuf_qn_1263(.A(qn_in_1263), .Y(g1660));
CLKBUFX1 gbuf_d_1264(.A(gbuf182), .Y(d_out_1264));
CLKBUFX1 gbuf_qn_1264(.A(qn_in_1264), .Y(g2364));
INVX1 g67488(.A (g5648), .Y (n_761));
CLKBUFX1 gbuf_d_1265(.A(n_5382), .Y(d_out_1265));
CLKBUFX1 gbuf_q_1265(.A(q_in_1265), .Y(gbuf35));
CLKBUFX1 gbuf_d_1266(.A(gbuf176), .Y(d_out_1266));
CLKBUFX1 gbuf_qn_1266(.A(qn_in_1266), .Y(g2528));
CLKBUFX1 gbuf_d_1267(.A(gbuf130), .Y(d_out_1267));
CLKBUFX1 gbuf_qn_1267(.A(qn_in_1267), .Y(g1664));
CLKBUFX1 gbuf_d_1268(.A(gbuf131), .Y(d_out_1268));
CLKBUFX1 gbuf_qn_1268(.A(qn_in_1268), .Y(g1666));
AND2X1 g67850(.A (n_758), .B (n_757), .Y (n_759));
NAND2X1 g67907(.A (g1694), .B (n_755), .Y (n_756));
NAND2X1 g67919(.A (g_10959), .B (n_753), .Y (n_754));
NOR2X1 g67942(.A (g999), .B (n_8718), .Y (n_752));
AND2X1 g67985(.A (g_10841), .B (n_753), .Y (n_751));
AND2X1 g67997(.A (n_749), .B (n_748), .Y (n_750));
NOR2X1 g68043(.A (g1005), .B (n_8718), .Y (n_747));
NOR2X1 g68041(.A (g1997), .B (g7052), .Y (n_745));
AND2X1 g68064(.A (n_616), .B (n_569), .Y (n_744));
INVX1 g68173(.A (n_755), .Y (g5511));
INVX1 g68243(.A (n_2014), .Y (g6750));
INVX1 g68265(.A (n_742), .Y (n_2389));
INVX1 g68364(.A (n_753), .Y (n_6914));
INVX1 g68383(.A (n_739), .Y (n_935));
INVX1 g68421(.A (n_6822), .Y (g7302));
NOR2X1 g67926(.A (g1002), .B (n_8718), .Y (n_737));
CLKBUFX1 gbuf_d_1269(.A(n_670), .Y(d_out_1269));
CLKBUFX1 gbuf_q_1269(.A(q_in_1269), .Y(g2180));
NAND4X1 g66599(.A (g101), .B (n_734), .C (n_733), .D (n_5473), .Y(n_735));
INVX1 g65818(.A (n_731), .Y (n_732));
NOR2X1 g66596(.A (n_654), .B (n_483), .Y (n_4674));
NOR2X1 g67933(.A (g1557), .B (n_757), .Y (n_730));
AND2X1 g67900(.A (g1697), .B (n_755), .Y (n_729));
CLKBUFX1 gbuf_d_1270(.A(g813), .Y(d_out_1270));
CLKBUFX1 gbuf_q_1270(.A(q_in_1270), .Y(gbuf77));
AND2X1 g67934(.A (n_726), .B (n_748), .Y (n_727));
CLKBUFX1 gbuf_d_1271(.A(n_640), .Y(d_out_1271));
CLKBUFX1 gbuf_q_1271(.A(q_in_1271), .Y(g2175));
CLKBUFX1 gbuf_d_1272(.A(n_643), .Y(d_out_1272));
CLKBUFX1 gbuf_q_1272(.A(q_in_1272), .Y(n_471));
CLKBUFX3 g68346(.A (n_757), .Y (n_853));
CLKBUFX1 gbuf_d_1273(.A(n_591), .Y(d_out_1273));
CLKBUFX1 gbuf_q_1273(.A(q_in_1273), .Y(g2170));
CLKBUFX1 gbuf_d_1274(.A(n_568), .Y(d_out_1274));
CLKBUFX1 gbuf_q_1274(.A(q_in_1274), .Y(g2190));
CLKBUFX1 gbuf_d_1275(.A(n_578), .Y(d_out_1275));
CLKBUFX1 gbuf_q_1275(.A(q_in_1275), .Y(g8249));
CLKBUFX1 gbuf_d_1276(.A(n_594), .Y(d_out_1276));
CLKBUFX1 gbuf_q_1276(.A(q_in_1276), .Y(g1476));
CLKBUFX1 gbuf_d_1277(.A(n_580), .Y(d_out_1277));
CLKBUFX1 gbuf_q_1277(.A(q_in_1277), .Y(g3993));
CLKBUFX1 gbuf_d_1278(.A(n_589), .Y(d_out_1278));
CLKBUFX1 gbuf_q_1278(.A(q_in_1278), .Y(g2185));
MX2X1 g66640(.A (g1686), .B (g1672), .S0 (g3229), .Y (n_723));
CLKBUFX1 gbuf_d_1279(.A(n_581), .Y(d_out_1279));
CLKBUFX1 gbuf_q_1279(.A(q_in_1279), .Y(g6442));
CLKBUFX1 gbuf_d_1280(.A(n_4110), .Y(d_out_1280));
CLKBUFX1 gbuf_q_1280(.A(q_in_1280), .Y(gbuf83));
CLKBUFX1 gbuf_d_1281(.A(g7961), .Y(d_out_1281));
CLKBUFX1 gbuf_q_1281(.A(q_in_1281), .Y(g8007));
NOR2X1 g66549(.A (n_601), .B (n_474), .Y (n_775));
NOR2X1 g67196(.A (n_695), .B (n_699), .Y (n_1086));
CLKBUFX1 gbuf_d_1282(.A(n_605), .Y(d_out_1282));
CLKBUFX1 gbuf_q_1282(.A(q_in_1282), .Y(g8251));
CLKBUFX1 gbuf_d_1283(.A(n_579), .Y(d_out_1283));
CLKBUFX1 gbuf_q_1283(.A(q_in_1283), .Y(g4200));
INVX1 g68308(.A (n_2170), .Y (g6485));
OR2X1 g68036(.A (g585), .B (n_2170), .Y (n_721));
INVX1 g68266(.A (n_8413), .Y (n_742));
OR2X1 g68026(.A (g1271), .B (n_2014), .Y (n_719));
OR2X1 g67943(.A (g579), .B (n_2170), .Y (n_718));
CLKBUFX1 gbuf_d_1284(.A(n_556), .Y(d_out_1284));
CLKBUFX1 gbuf_q_1284(.A(q_in_1284), .Y(g7334));
CLKBUFX1 gbuf_d_1285(.A(n_555), .Y(d_out_1285));
CLKBUFX1 gbuf_q_1285(.A(q_in_1285), .Y(g6895));
CLKBUFX1 gbuf_d_1286(.A(n_554), .Y(d_out_1286));
CLKBUFX1 gbuf_q_1286(.A(q_in_1286), .Y(g6225));
CLKBUFX1 gbuf_d_1287(.A(g5629), .Y(d_out_1287));
CLKBUFX1 gbuf_q_1287(.A(q_in_1287), .Y(g5648));
OR2X1 g67999(.A (g2812), .B (n_1245), .Y (n_715));
CLKBUFX1 gbuf_d_1288(.A(g5388), .Y(d_out_1288));
CLKBUFX1 gbuf_qn_1288(.A(qn_in_1288), .Y(g2986));
CLKBUFX1 gbuf_d_1289(.A(n_4112), .Y(d_out_1289));
CLKBUFX1 gbuf_q_1289(.A(q_in_1289), .Y(gbuf84));
CLKBUFX1 gbuf_d_1290(.A(g8012), .Y(d_out_1290));
CLKBUFX1 gbuf_q_1290(.A(q_in_1290), .Y(g8082));
CLKBUFX1 gbuf_d_1291(.A(g105), .Y(d_out_1291));
CLKBUFX1 gbuf_q_1291(.A(q_in_1291), .Y(gbuf33));
CLKBUFX1 gbuf_d_1292(.A(gbuf178), .Y(d_out_1292));
CLKBUFX1 gbuf_qn_1292(.A(qn_in_1292), .Y(g2356));
CLKBUFX1 gbuf_d_1293(.A(n_571), .Y(d_out_1293));
CLKBUFX1 gbuf_q_1293(.A(q_in_1293), .Y(n_600));
OAI21X1 g67383(.A0 (n_655), .A1 (n_377), .B0 (n_528), .Y (n_8103));
CLKBUFX1 gbuf_d_1294(.A(n_583), .Y(d_out_1294));
CLKBUFX1 gbuf_q_1294(.A(q_in_1294), .Y(g4321));
NOR2X1 g65823(.A (n_459), .B (n_542), .Y (n_714));
NAND2X1 g67067(.A (g3211), .B (n_545), .Y (n_713));
NAND2X1 g66324(.A (n_711), .B (n_712), .Y (n_893));
NAND2X1 g66433(.A (n_707), .B (n_712), .Y (n_892));
AND2X1 g66457(.A (n_711), .B (n_710), .Y (n_981));
OR2X1 g67949(.A (g1965), .B (n_864), .Y (n_709));
AND2X1 g66461(.A (n_707), .B (n_710), .Y (n_982));
AND2X1 g66468(.A (n_706), .B (g3013), .Y (n_731));
XOR2X1 g66621(.A (g3006), .B (n_456), .Y (n_705));
NAND4X1 g66630(.A (n_597), .B (n_417), .C (g3201), .D (n_344), .Y(n_704));
MX2X1 g66641(.A (n_101), .B (g2366), .S0 (g3229), .Y (n_703));
INVX1 g66778(.A (g3109), .Y (n_701));
NOR2X1 g66953(.A (n_803), .B (n_698), .Y (n_2188));
NAND2X1 g67027(.A (g3086), .B (n_545), .Y (n_700));
NOR2X1 g67054(.A (n_803), .B (n_694), .Y (n_1063));
NOR2X1 g67055(.A (n_699), .B (n_697), .Y (n_1053));
NOR2X1 g67104(.A (n_564), .B (n_803), .Y (n_877));
OR2X1 g67153(.A (n_699), .B (n_698), .Y (n_801));
NOR2X1 g67158(.A (n_803), .B (n_697), .Y (n_1463));
NOR2X1 g67200(.A (n_803), .B (n_695), .Y (n_696));
NOR2X1 g67231(.A (n_699), .B (n_694), .Y (n_2187));
NOR2X1 g67281(.A (g1762), .B (g_29316), .Y (n_693));
NOR2X1 g67287(.A (g1747), .B (g_29316), .Y (n_692));
NOR2X1 g67309(.A (g1777), .B (g_29316), .Y (n_691));
NAND2X1 g67318(.A (g_29316), .B (g_32166), .Y (n_1363));
NOR2X1 g67336(.A (g1732), .B (g_29316), .Y (n_690));
NOR2X1 g67360(.A (g2643), .B (n_6822), .Y (n_689));
OAI21X1 g67394(.A0 (g1243), .A1 (n_645), .B0 (n_538), .Y (n_882));
NOR2X1 g67321(.A (g396), .B (g5629), .Y (n_688));
CLKBUFX1 gbuf_d_1295(.A(gbuf181), .Y(d_out_1295));
CLKBUFX1 gbuf_qn_1295(.A(qn_in_1295), .Y(g2362));
CLKBUFX1 gbuf_d_1296(.A(n_3169), .Y(d_out_1296));
CLKBUFX1 gbuf_q_1296(.A(q_in_1296), .Y(gbuf81));
CLKBUFX1 gbuf_d_1297(.A(gbuf129), .Y(d_out_1297));
CLKBUFX1 gbuf_qn_1297(.A(qn_in_1297), .Y(g1662));
NAND2X1 g67026(.A (g3158), .B (n_545), .Y (n_687));
CLKBUFX1 gbuf_d_1298(.A(gbuf177), .Y(d_out_1298));
CLKBUFX1 gbuf_qn_1298(.A(qn_in_1298), .Y(g2354));
CLKBUFX1 gbuf_d_1299(.A(n_3167), .Y(d_out_1299));
CLKBUFX1 gbuf_q_1299(.A(q_in_1299), .Y(gbuf80));
CLKBUFX1 gbuf_d_1300(.A(g7909), .Y(d_out_1300));
CLKBUFX1 gbuf_q_1300(.A(q_in_1300), .Y(g7956));
OR2X1 g68040(.A (g582), .B (n_2170), .Y (n_686));
NAND3X1 g68062(.A (n_631), .B (n_357), .C (n_411), .Y (n_903));
CLKBUFX1 gbuf_d_1301(.A(n_561), .Y(d_out_1301));
CLKBUFX1 gbuf_q_1301(.A(q_in_1301), .Y(g4090));
INVX2 g68321(.A (n_682), .Y (n_840));
INVX2 g68322(.A (n_682), .Y (n_2308));
INVX1 g68385(.A (n_748), .Y (n_739));
CLKBUFX1 gbuf_d_1302(.A(n_558), .Y(d_out_1302));
CLKBUFX1 gbuf_q_1302(.A(q_in_1302), .Y(g4450));
XOR2X1 g66639(.A (n_679), .B (n_603), .Y (n_680));
OR2X1 g67953(.A (g1962), .B (n_864), .Y (n_678));
NOR2X1 g67010(.A (n_369), .B (n_595), .Y (n_3873));
CLKBUFX1 gbuf_d_1303(.A(g8087), .Y(d_out_1303));
CLKBUFX1 gbuf_q_1303(.A(q_in_1303), .Y(g8167));
OR2X1 g67289(.A (n_540), .B (n_676), .Y (n_677));
OAI21X1 g67385(.A0 (g1937), .A1 (n_659), .B0 (n_522), .Y (n_7992));
INVX1 g67522(.A (g_25914), .Y (g5686));
CLKBUFX1 gbuf_d_1304(.A(n_560), .Y(d_out_1304));
CLKBUFX1 gbuf_q_1304(.A(q_in_1304), .Y(g8023));
CLKBUFX1 gbuf_d_1305(.A(n_557), .Y(d_out_1305));
CLKBUFX1 gbuf_q_1305(.A(q_in_1305), .Y(g4088));
CLKBUFX1 gbuf_d_1306(.A(n_3164), .Y(d_out_1306));
CLKBUFX1 gbuf_q_1306(.A(q_in_1306), .Y(gbuf78));
CLKBUFX1 gbuf_d_1307(.A(n_576), .Y(d_out_1307));
CLKBUFX1 gbuf_q_1307(.A(q_in_1307), .Y(g8175));
CLKBUFX1 gbuf_d_1308(.A(gbuf127), .Y(d_out_1308));
CLKBUFX1 gbuf_qn_1308(.A(qn_in_1308), .Y(g1834));
CLKBUFX1 gbuf_d_1309(.A(n_559), .Y(d_out_1309));
CLKBUFX1 gbuf_q_1309(.A(q_in_1309), .Y(g4323));
CLKBUFX1 gbuf_d_1310(.A(n_546), .Y(d_out_1310));
CLKBUFX1 gbuf_q_1310(.A(q_in_1310), .Y(g1501));
CLKBUFX1 gbuf_d_1311(.A(n_592), .Y(d_out_1311));
CLKBUFX1 gbuf_q_1311(.A(q_in_1311), .Y(g4590));
CLKBUFX1 gbuf_d_1312(.A(n_547), .Y(d_out_1312));
CLKBUFX1 gbuf_q_1312(.A(q_in_1312), .Y(n_473));
CLKBUFX1 gbuf_d_1313(.A(n_365), .Y(d_out_1313));
CLKBUFX1 gbuf_q_1313(.A(q_in_1313), .Y(gbuf133));
NOR2X1 g66941(.A (n_475), .B (g557), .Y (n_767));
CLKBUFX1 gbuf_d_1314(.A(n_447), .Y(d_out_1314));
CLKBUFX1 gbuf_q_1314(.A(q_in_1314), .Y(gbuf176));
CLKBUFX1 gbuf_d_1315(.A(n_454), .Y(d_out_1315));
CLKBUFX1 gbuf_q_1315(.A(q_in_1315), .Y(gbuf130));
INVX1 g68386(.A (g_4886), .Y (n_748));
MX2X1 g67432(.A (g1486), .B (g2944), .S0 (g2879), .Y (n_672));
MX2X1 g67430(.A (g2165), .B (g2963), .S0 (g2879), .Y (n_671));
CLKBUFX1 gbuf_d_1316(.A(gbuf36), .Y(d_out_1316));
CLKBUFX1 gbuf_qn_1316(.A(qn_in_1316), .Y(g_31512));
MX2X1 g67428(.A (g2180), .B (g2972), .S0 (g2879), .Y (n_670));
CLKBUFX1 gbuf_d_1317(.A(g1672), .Y(d_out_1317));
CLKBUFX1 gbuf_q_1317(.A(q_in_1317), .Y(g1921));
CLKBUFX1 gbuf_d_1318(.A(gbuf85), .Y(d_out_1318));
CLKBUFX1 gbuf_qn_1318(.A(qn_in_1318), .Y(g978));
OR2X1 g67976(.A (g1268), .B (n_2014), .Y (n_669));
NOR2X1 g67322(.A (g2471), .B (g5747), .Y (n_667));
INVX1 g68351(.A (g_9649), .Y (n_666));
CLKBUFX2 g68324(.A (g_12670), .Y (n_682));
NAND2X1 g67282(.A (g2441), .B (g5796), .Y (n_665));
AND2X1 g67946(.A (g2095), .B (n_562), .Y (n_664));
CLKBUFX1 gbuf_d_1319(.A(g5796), .Y(d_out_1319));
CLKBUFX1 gbuf_q_1319(.A(q_in_1319), .Y(g2412));
CLKBUFX1 gbuf_d_1320(.A(g8030), .Y(d_out_1320));
CLKBUFX1 gbuf_q_1320(.A(q_in_1320), .Y(g3109));
AND2X1 g67886(.A (g2086), .B (n_562), .Y (n_662));
MX2X1 g67424(.A (g1481), .B (g2941), .S0 (g2879), .Y (n_661));
CLKBUFX1 gbuf_d_1321(.A(n_505), .Y(d_out_1321));
CLKBUFX1 gbuf_qn_1321(.A(qn_in_1321), .Y(g2817));
INVX1 g68207(.A (n_864), .Y (g7052));
AND2X1 g67887(.A (g2089), .B (n_562), .Y (n_660));
AOI21X1 g67395(.A0 (g1937), .A1 (n_659), .B0 (n_521), .Y (n_7892));
CLKBUFX1 gbuf_d_1322(.A(n_3187), .Y(d_out_1322));
CLKBUFX1 gbuf_q_1322(.A(q_in_1322), .Y(gbuf32));
INVX2 g68175(.A (g_15833), .Y (n_755));
CLKBUFX1 gbuf_d_1323(.A(g2366), .Y(d_out_1323));
CLKBUFX1 gbuf_q_1323(.A(q_in_1323), .Y(g2615));
NAND3X1 g67369(.A (n_504), .B (n_656), .C (g801), .Y (n_657));
AOI21X1 g67384(.A0 (n_655), .A1 (n_377), .B0 (n_527), .Y (n_8084));
NOR2X1 g66395(.A (n_455), .B (n_254), .Y (n_789));
CLKBUFX1 gbuf_d_1324(.A(n_2706), .Y(d_out_1324));
CLKBUFX1 gbuf_q_1324(.A(q_in_1324), .Y(gbuf175));
CLKBUFX1 gbuf_d_1325(.A(n_2719), .Y(d_out_1325));
CLKBUFX1 gbuf_q_1325(.A(q_in_1325), .Y(gbuf179));
NAND4X1 g66940(.A (g2185), .B (n_415), .C (g2180), .D (g2175), .Y(n_654));
CLKBUFX1 gbuf_d_1326(.A(n_4639), .Y(d_out_1326));
CLKBUFX1 gbuf_q_1326(.A(q_in_1326), .Y(gbuf128));
INVX1 g66973(.A (n_706), .Y (n_652));
CLKBUFX1 gbuf_d_1327(.A(n_4368), .Y(d_out_1327));
CLKBUFX1 gbuf_q_1327(.A(q_in_1327), .Y(gbuf182));
INVX1 g67260(.A (n_518), .Y (n_783));
NAND2X1 g67273(.A (g2471), .B (g5796), .Y (n_651));
NAND2X1 g67279(.A (g2456), .B (g5796), .Y (n_650));
NOR2X1 g67280(.A (g2456), .B (g5747), .Y (n_649));
NAND2X1 g67295(.A (g2426), .B (g5796), .Y (n_648));
OR2X1 g67308(.A (g5796), .B (g5747), .Y (n_1209));
NAND3X1 g67323(.A (g97), .B (n_9490), .C (g109), .Y (n_647));
NOR2X1 g67362(.A (g_18059), .B (g5629), .Y (n_646));
AOI21X1 g67386(.A0 (g1243), .A1 (n_645), .B0 (n_537), .Y (n_7462));
MX2X1 g67421(.A (n_471), .B (g2953), .S0 (g2879), .Y (n_643));
NOR2X1 g67317(.A (g_27919), .B (g5629), .Y (n_642));
MX2X1 g67433(.A (g2175), .B (g2969), .S0 (g2879), .Y (n_640));
MX2X1 g67434(.A (g1471), .B (g2935), .S0 (g2879), .Y (n_639));
MX2X1 g67435(.A (g2195), .B (g2981), .S0 (g2879), .Y (n_638));
CLKBUFX1 gbuf_d_1328(.A(gbuf132), .Y(d_out_1328));
CLKBUFX1 gbuf_qn_1328(.A(qn_in_1328), .Y(g1668));
NOR2X1 g68065(.A (n_5473), .B (n_733), .Y (n_636));
INVX2 g68347(.A (g_12670), .Y (n_757));
CLKBUFX1 gbuf_d_1329(.A(n_5247), .Y(d_out_1329));
CLKBUFX1 gbuf_q_1329(.A(q_in_1329), .Y(gbuf31));
INVX1 g67644(.A (g_29316), .Y (g5738));
MX2X1 g67431(.A (n_482), .B (g2874), .S0 (g2879), .Y (n_634));
CLKBUFX1 gbuf_d_1330(.A(n_5380), .Y(d_out_1330));
CLKBUFX1 gbuf_q_1330(.A(q_in_1330), .Y(gbuf34));
OR2X1 g67852(.A (g1265), .B (n_2014), .Y (n_633));
NAND2X1 g67928(.A (g2622), .B (n_6822), .Y (n_632));
NAND2X1 g67984(.A (n_631), .B (n_536), .Y (n_802));
NOR2X1 g68049(.A (n_413), .B (n_460), .Y (n_2946));
NAND2X1 g68063(.A (n_468), .B (g805), .Y (n_630));
CLKBUFX1 gbuf_d_1331(.A(n_435), .Y(d_out_1331));
CLKBUFX1 gbuf_q_1331(.A(q_in_1331), .Y(gbuf131));
INVX1 g68096(.A (g6677), .Y (n_1916));
INVX1 g68127(.A (n_1245), .Y (g7425));
OR2X1 g67927(.A (g2118), .B (n_562), .Y (n_624));
INVX2 g68366(.A (g_9649), .Y (n_753));
NOR2X1 g68558(.A (n_344), .B (n_264), .Y (n_619));
NOR2X1 g67361(.A (g2441), .B (g5747), .Y (n_617));
NOR2X1 g68575(.A (n_355), .B (n_264), .Y (n_616));
OR2X1 g67918(.A (g1424), .B (n_8625), .Y (n_614));
NAND2X1 g67267(.A (g2929), .B (g8021), .Y (n_613));
CLKBUFX1 gbuf_d_1332(.A(g5657), .Y(d_out_1332));
CLKBUFX1 gbuf_qn_1332(.A(qn_in_1332), .Y(g_25914));
CLKBUFX1 g68489(.A (g121), .Y (n_3161));
INVX1 g68481(.A (g_19064), .Y (n_9593));
NOR2X1 g67264(.A (g2426), .B (g5747), .Y (n_609));
CLKBUFX1 gbuf_d_1333(.A(n_484), .Y(d_out_1333));
CLKBUFX1 gbuf_qn_1333(.A(qn_in_1333), .Y(g3054));
NOR2X1 g66976(.A (n_477), .B (g2888), .Y (n_608));
INVX2 g68459(.A (g_19064), .Y (n_810));
NAND4X1 g67873(.A (g2185), .B (n_482), .C (n_385), .D (n_447), .Y(n_2952));
CLKBUFX1 gbuf_d_1334(.A(gbuf126), .Y(d_out_1334));
CLKBUFX1 gbuf_qn_1334(.A(qn_in_1334), .Y(g1832));
CLKBUFX1 gbuf_d_1335(.A(n_436), .Y(d_out_1335));
CLKBUFX1 gbuf_q_1335(.A(q_in_1335), .Y(gbuf180));
MX2X1 g67403(.A (g2874), .B (g8251), .S0 (g2879), .Y (n_605));
NAND2X1 g67857(.A (g3210), .B (n_422), .Y (n_602));
CLKBUFX1 gbuf_d_1336(.A(n_379), .Y(d_out_1336));
CLKBUFX1 gbuf_q_1336(.A(q_in_1336), .Y(g_9649));
CLKBUFX1 gbuf_d_1337(.A(n_379), .Y(d_out_1337));
CLKBUFX1 gbuf_q_1337(.A(q_in_1337), .Y(g_4886));
NAND4X1 g66939(.A (n_600), .B (n_366), .C (g1486), .D (g1481), .Y(n_601));
NAND2X1 g68059(.A (g1928), .B (n_864), .Y (n_599));
CLKBUFX1 gbuf_d_1338(.A(n_2809), .Y(d_out_1338));
CLKBUFX1 gbuf_q_1338(.A(q_in_1338), .Y(gbuf181));
NAND2X1 g67826(.A (n_431), .B (n_180), .Y (n_595));
MX2X1 g67426(.A (g1476), .B (g2938), .S0 (g2879), .Y (n_594));
NOR2X1 g68593(.A (g557), .B (n_3701), .Y (n_593));
MX2X1 g67401(.A (g2975), .B (g4590), .S0 (g2879), .Y (n_592));
CLKBUFX1 gbuf_d_1339(.A(g3234), .Y(d_out_1339));
CLKBUFX1 gbuf_q_1339(.A(q_in_1339), .Y(g5388));
MX2X1 g67423(.A (g2170), .B (g2966), .S0 (g2879), .Y (n_591));
CLKBUFX1 g68316(.A (n_590), .Y (n_4112));
MX2X1 g67422(.A (g2185), .B (g2975), .S0 (g2879), .Y (n_589));
NAND2X1 g67963(.A (g3085), .B (n_422), .Y (n_588));
OR2X1 g68031(.A (g2659), .B (n_6822), .Y (n_587));
XOR2X1 g67417(.A (g2944), .B (g2941), .Y (n_585));
CLKBUFX1 gbuf_d_1340(.A(n_379), .Y(d_out_1340));
CLKBUFX1 gbuf_q_1340(.A(q_in_1340), .Y(g_13515));
XOR2X1 g67413(.A (g2978), .B (g2975), .Y (n_584));
MX2X1 g67412(.A (g2953), .B (g4321), .S0 (g2879), .Y (n_583));
CLKBUFX1 gbuf_d_1341(.A(g5695), .Y(d_out_1341));
CLKBUFX1 gbuf_qn_1341(.A(qn_in_1341), .Y(g_29316));
MX2X1 g67408(.A (g2969), .B (g6442), .S0 (g2879), .Y (n_581));
MX2X1 g67407(.A (g2941), .B (g3993), .S0 (g2879), .Y (n_580));
MX2X1 g67405(.A (g2938), .B (g4200), .S0 (g2879), .Y (n_579));
MX2X1 g67402(.A (g2959), .B (g8249), .S0 (g2879), .Y (n_578));
MX2X1 g67397(.A (g2944), .B (g8175), .S0 (g2879), .Y (n_576));
CLKBUFX1 gbuf_d_1342(.A(n_379), .Y(d_out_1342));
CLKBUFX1 gbuf_q_1342(.A(q_in_1342), .Y(g_8360));
MX2X1 g67436(.A (n_600), .B (g2947), .S0 (g2879), .Y (n_571));
NAND2X1 g67982(.A (g3155), .B (n_422), .Y (n_570));
NAND2X1 g67977(.A (n_425), .B (n_569), .Y (n_697));
MX2X1 g67425(.A (g2190), .B (g2978), .S0 (g2879), .Y (n_568));
OR2X1 g68038(.A (g2656), .B (n_6822), .Y (n_565));
NAND2X1 g68563(.A (n_411), .B (g3207), .Y (n_564));
CLKBUFX1 gbuf_d_1343(.A(n_2716), .Y(d_out_1343));
CLKBUFX1 gbuf_q_1343(.A(q_in_1343), .Y(gbuf178));
CLKBUFX1 gbuf_d_1344(.A(n_293), .Y(d_out_1344));
CLKBUFX1 gbuf_q_1344(.A(q_in_1344), .Y(gbuf129));
NOR2X1 g68066(.A (n_5247), .B (n_467), .Y (n_734));
AND2X1 g67945(.A (g2083), .B (n_562), .Y (n_563));
NOR2X1 g67171(.A (n_803), .B (n_416), .Y (n_707));
NOR2X1 g67180(.A (n_356), .B (n_803), .Y (n_711));
MX2X1 g67398(.A (g2981), .B (g4090), .S0 (g2879), .Y (n_561));
MX2X1 g67399(.A (g2947), .B (g8023), .S0 (g2879), .Y (n_560));
MX2X1 g67400(.A (g2978), .B (g4323), .S0 (g2879), .Y (n_559));
MX2X1 g67404(.A (g2935), .B (g4450), .S0 (g2879), .Y (n_558));
MX2X1 g67406(.A (g2956), .B (g4088), .S0 (g2879), .Y (n_557));
MX2X1 g67409(.A (g2963), .B (g7334), .S0 (g2879), .Y (n_556));
MX2X1 g67410(.A (g2966), .B (g6895), .S0 (g2879), .Y (n_555));
MX2X1 g67411(.A (g2972), .B (g6225), .S0 (g2879), .Y (n_554));
XOR2X1 g67414(.A (g2874), .B (g2981), .Y (n_553));
XOR2X1 g67415(.A (g2972), .B (g2969), .Y (n_552));
XOR2X1 g67416(.A (g2938), .B (g2935), .Y (n_551));
XOR2X1 g67418(.A (g2953), .B (g2947), .Y (n_550));
XOR2X1 g67419(.A (g2966), .B (g2963), .Y (n_549));
XOR2X1 g67420(.A (g2959), .B (g2956), .Y (n_548));
MX2X1 g67427(.A (n_473), .B (g2959), .S0 (g2879), .Y (n_547));
MX2X1 g67429(.A (g1501), .B (g2956), .S0 (g2879), .Y (n_546));
INVX1 g67438(.A (g8030), .Y (n_545));
INVX1 g67991(.A (n_456), .Y (n_542));
OR2X1 g67996(.A (n_539), .B (n_100), .Y (n_540));
INVX1 g68006(.A (n_537), .Y (n_538));
NAND3X1 g68013(.A (n_536), .B (g3201), .C (g3207), .Y (n_698));
OR2X1 g68022(.A (g1959), .B (n_864), .Y (n_535));
NAND3X1 g68067(.A (n_569), .B (n_355), .C (g3201), .Y (n_695));
CLKBUFX1 gbuf_d_1345(.A(n_385), .Y(d_out_1345));
CLKBUFX1 gbuf_q_1345(.A(q_in_1345), .Y(gbuf177));
CLKBUFX1 gbuf_d_1346(.A(n_343), .Y(d_out_1346));
CLKBUFX1 gbuf_q_1346(.A(q_in_1346), .Y(gbuf127));
INVX1 g68097(.A (n_9208), .Y (g6677));
CLKBUFX1 g68141(.A (n_762), .Y (n_3164));
CLKBUFX1 gbuf_d_1347(.A(n_379), .Y(d_out_1347));
CLKBUFX1 gbuf_q_1347(.A(q_in_1347), .Y(g7909));
INVX2 g68310(.A (n_529), .Y (n_2170));
INVX1 g68044(.A (n_527), .Y (n_528));
CLKBUFX1 gbuf_d_1348(.A(n_379), .Y(d_out_1348));
CLKBUFX1 gbuf_q_1348(.A(q_in_1348), .Y(g_12670));
CLKBUFX1 gbuf_d_1349(.A(n_379), .Y(d_out_1349));
CLKBUFX1 gbuf_q_1349(.A(q_in_1349), .Y(g8012));
CLKBUFX1 g68503(.A (n_525), .Y (n_3169));
INVX1 g68526(.A (n_8625), .Y (g6979));
CLKBUFX1 gbuf_d_1350(.A(n_379), .Y(d_out_1350));
CLKBUFX1 gbuf_q_1350(.A(q_in_1350), .Y(g_19064));
INVX1 g67966(.A (n_521), .Y (n_522));
NOR2X1 g67145(.A (n_803), .B (g185), .Y (n_519));
NAND2X1 g67890(.A (n_410), .B (n_536), .Y (n_694));
OR4X1 g66977(.A (g3002), .B (g3006), .C (g3013), .D (n_288), .Y(n_4151));
NOR2X1 g66974(.A (n_225), .B (n_456), .Y (n_706));
NAND3X1 g67261(.A (n_478), .B (n_517), .C (n_679), .Y (n_518));
CLKBUFX1 gbuf_d_1351(.A(n_379), .Y(d_out_1351));
CLKBUFX1 gbuf_q_1351(.A(q_in_1351), .Y(g_17130));
CLKBUFX1 gbuf_d_1352(.A(n_379), .Y(d_out_1352));
CLKBUFX1 gbuf_q_1352(.A(q_in_1352), .Y(g_15833));
CLKBUFX1 gbuf_d_1353(.A(n_379), .Y(d_out_1353));
CLKBUFX1 gbuf_q_1353(.A(q_in_1353), .Y(g7961));
INVX1 g68414(.A (g801), .Y (n_3167));
INVX1 g68406(.A (n_562), .Y (g7229));
CLKBUFX1 gbuf_d_1354(.A(n_379), .Y(d_out_1354));
CLKBUFX1 gbuf_q_1354(.A(q_in_1354), .Y(g8087));
CLKBUFX1 gbuf_d_1355(.A(gbuf97), .Y(d_out_1355));
CLKBUFX1 gbuf_qn_1355(.A(qn_in_1355), .Y(g1011));
CLKBUFX1 gbuf_d_1356(.A(g8106), .Y(d_out_1356));
CLKBUFX1 gbuf_q_1356(.A(q_in_1356), .Y(g8030));
NOR2X1 g68554(.A (g51), .B (n_233), .Y (n_505));
CLKBUFX1 gbuf_d_1357(.A(gbuf106), .Y(d_out_1357));
CLKBUFX1 gbuf_q_1357(.A(q_in_1357), .Y(g1259));
CLKBUFX1 gbuf_d_1358(.A(gbuf44), .Y(d_out_1358));
CLKBUFX1 gbuf_q_1358(.A(q_in_1358), .Y(g_18059));
CLKBUFX1 gbuf_d_1359(.A(gbuf135), .Y(d_out_1359));
CLKBUFX1 gbuf_q_1359(.A(q_in_1359), .Y(g1730));
CLKBUFX1 gbuf_d_1360(.A(g5747), .Y(d_out_1360));
CLKBUFX1 gbuf_q_1360(.A(q_in_1360), .Y(g5796));
CLKBUFX1 gbuf_d_1361(.A(gbuf144), .Y(d_out_1361));
CLKBUFX1 gbuf_q_1361(.A(q_in_1361), .Y(g1775));
CLKBUFX1 gbuf_d_1362(.A(gbuf107), .Y(d_out_1362));
CLKBUFX1 gbuf_q_1362(.A(q_in_1362), .Y(g1251));
INVX1 g68317(.A (n_504), .Y (n_590));
CLKBUFX1 gbuf_d_1363(.A(gbuf189), .Y(d_out_1363));
CLKBUFX1 gbuf_q_1363(.A(q_in_1363), .Y(g2443));
CLKBUFX1 gbuf_d_1364(.A(gbuf92), .Y(d_out_1364));
CLKBUFX1 gbuf_q_1364(.A(q_in_1364), .Y(g1066));
CLKBUFX1 gbuf_d_1365(.A(gbuf45), .Y(d_out_1365));
CLKBUFX1 gbuf_q_1365(.A(q_in_1365), .Y(g_7905));
CLKBUFX1 gbuf_d_1366(.A(gbuf89), .Y(d_out_1366));
CLKBUFX1 gbuf_q_1366(.A(q_in_1366), .Y(g1051));
CLKBUFX1 gbuf_d_1367(.A(gbuf56), .Y(d_out_1367));
CLKBUFX1 gbuf_q_1367(.A(q_in_1367), .Y(g571));
CLKBUFX1 gbuf_d_1368(.A(gbuf194), .Y(d_out_1368));
CLKBUFX1 gbuf_q_1368(.A(q_in_1368), .Y(g2471));
CLKBUFX1 gbuf_d_1369(.A(gbuf157), .Y(d_out_1369));
CLKBUFX1 gbuf_qn_1369(.A(qn_in_1369), .Y(g1947));
AND2X1 g68045(.A (n_501), .B (g2599), .Y (n_527));
CLKBUFX1 gbuf_d_1370(.A(gbuf37), .Y(d_out_1370));
CLKBUFX1 gbuf_qn_1370(.A(qn_in_1370), .Y(g_19985));
INVX1 g68312(.A (n_1498), .Y (n_529));
CLKBUFX1 gbuf_d_1371(.A(gbuf155), .Y(d_out_1371));
CLKBUFX1 gbuf_q_1371(.A(q_in_1371), .Y(g1953));
CLKBUFX1 gbuf_d_1372(.A(gbuf207), .Y(d_out_1372));
CLKBUFX1 gbuf_qn_1372(.A(qn_in_1372), .Y(g2564));
CLKBUFX1 gbuf_d_1373(.A(gbuf88), .Y(d_out_1373));
CLKBUFX1 gbuf_qn_1373(.A(qn_in_1373), .Y(g1040));
CLKBUFX1 gbuf_d_1374(.A(gbuf203), .Y(d_out_1374));
CLKBUFX1 gbuf_q_1374(.A(q_in_1374), .Y(g2645));
CLKBUFX1 gbuf_d_1375(.A(gbuf183), .Y(d_out_1375));
CLKBUFX1 gbuf_qn_1375(.A(qn_in_1375), .Y(g2366));
CLKBUFX1 gbuf_d_1376(.A(gbuf146), .Y(d_out_1376));
CLKBUFX1 gbuf_q_1376(.A(q_in_1376), .Y(g1705));
CLKBUFX1 gbuf_d_1377(.A(gbuf95), .Y(d_out_1377));
CLKBUFX1 gbuf_q_1377(.A(q_in_1377), .Y(g1081));
NAND3X1 g68011(.A (n_296), .B (g3151), .C (g3097), .Y (n_495));
CLKBUFX1 gbuf_d_1378(.A(gbuf204), .Y(d_out_1378));
CLKBUFX1 gbuf_q_1378(.A(q_in_1378), .Y(g2647));
OR2X1 g68047(.A (g2653), .B (g_14726), .Y (n_494));
CLKBUFX1 gbuf_d_1379(.A(gbuf91), .Y(d_out_1379));
CLKBUFX1 gbuf_qn_1379(.A(qn_in_1379), .Y(g1055));
CLKBUFX1 gbuf_d_1380(.A(gbuf134), .Y(d_out_1380));
CLKBUFX1 gbuf_qn_1380(.A(qn_in_1380), .Y(g1672));
CLKBUFX1 gbuf_d_1381(.A(g2857), .Y(d_out_1381));
CLKBUFX1 gbuf_q_1381(.A(q_in_1381), .Y(gbuf36));
CLKBUFX1 gbuf_d_1382(.A(gbuf143), .Y(d_out_1382));
CLKBUFX1 gbuf_q_1382(.A(q_in_1382), .Y(g1764));
CLKBUFX1 gbuf_d_1383(.A(gbuf141), .Y(d_out_1383));
CLKBUFX1 gbuf_q_1383(.A(q_in_1383), .Y(g1760));
CLKBUFX1 gbuf_d_1384(.A(gbuf40), .Y(d_out_1384));
CLKBUFX1 gbuf_q_1384(.A(q_in_1384), .Y(g_19959));
CLKBUFX1 gbuf_d_1385(.A(gbuf138), .Y(d_out_1385));
CLKBUFX1 gbuf_q_1385(.A(q_in_1385), .Y(g1745));
CLKBUFX1 gbuf_d_1386(.A(gbuf158), .Y(d_out_1386));
CLKBUFX1 gbuf_q_1386(.A(q_in_1386), .Y(g1870));
CLKBUFX1 gbuf_d_1387(.A(gbuf39), .Y(d_out_1387));
CLKBUFX1 gbuf_q_1387(.A(q_in_1387), .Y(g_13227));
CLKBUFX1 gbuf_d_1388(.A(g8021), .Y(d_out_1388));
CLKBUFX1 gbuf_qn_1388(.A(qn_in_1388), .Y(g2929));
CLKBUFX1 gbuf_d_1389(.A(gbuf137), .Y(d_out_1389));
CLKBUFX1 gbuf_q_1389(.A(q_in_1389), .Y(g1734));
CLKBUFX1 gbuf_d_1390(.A(gbuf90), .Y(d_out_1390));
CLKBUFX1 gbuf_qn_1390(.A(qn_in_1390), .Y(g1053));
CLKBUFX1 gbuf_d_1391(.A(gbuf94), .Y(d_out_1391));
CLKBUFX1 gbuf_qn_1391(.A(qn_in_1391), .Y(g1070));
CLKBUFX1 gbuf_d_1392(.A(gbuf191), .Y(d_out_1392));
CLKBUFX1 gbuf_q_1392(.A(q_in_1392), .Y(g2456));
CLKBUFX1 gbuf_d_1393(.A(gbuf188), .Y(d_out_1393));
CLKBUFX1 gbuf_q_1393(.A(q_in_1393), .Y(g2441));
CLKBUFX1 gbuf_d_1394(.A(gbuf190), .Y(d_out_1394));
CLKBUFX1 gbuf_qn_1394(.A(qn_in_1394), .Y(g2454));
CLKBUFX1 gbuf_d_1395(.A(gbuf42), .Y(d_out_1395));
CLKBUFX1 gbuf_q_1395(.A(q_in_1395), .Y(g_27149));
CLKBUFX1 gbuf_d_1396(.A(gbuf48), .Y(d_out_1396));
CLKBUFX1 gbuf_q_1396(.A(q_in_1396), .Y(g_28035));
CLKBUFX1 gbuf_d_1397(.A(gbuf58), .Y(d_out_1397));
CLKBUFX1 gbuf_q_1397(.A(q_in_1397), .Y(g565));
NOR2X1 g68539(.A (n_357), .B (g3201), .Y (n_710));
CLKBUFX1 gbuf_d_1398(.A(gbuf57), .Y(d_out_1398));
CLKBUFX1 gbuf_q_1398(.A(q_in_1398), .Y(g573));
INVX1 g69050(.A (g2180), .Y (n_2719));
CLKBUFX1 gbuf_d_1399(.A(gbuf105), .Y(d_out_1399));
CLKBUFX1 gbuf_q_1399(.A(q_in_1399), .Y(g1257));
NAND3X1 g67865(.A (n_517), .B (n_368), .C (n_782), .Y (n_487));
CLKBUFX1 gbuf_d_1400(.A(gbuf184), .Y(d_out_1400));
CLKBUFX1 gbuf_qn_1400(.A(qn_in_1400), .Y(g2424));
CLKBUFX1 gbuf_d_1401(.A(gbuf154), .Y(d_out_1401));
CLKBUFX1 gbuf_q_1401(.A(q_in_1401), .Y(g1951));
CLKBUFX1 gbuf_d_1402(.A(gbuf87), .Y(d_out_1402));
CLKBUFX1 gbuf_qn_1402(.A(qn_in_1402), .Y(g1038));
AND2X1 g67967(.A (n_485), .B (g1905), .Y (n_521));
AND2X1 g68559(.A (n_310), .B (g3080), .Y (n_484));
NAND3X1 g67849(.A (n_482), .B (g2195), .C (g2190), .Y (n_483));
CLKBUFX1 gbuf_d_1403(.A(gbuf108), .Y(d_out_1403));
CLKBUFX1 gbuf_qn_1403(.A(qn_in_1403), .Y(g1253));
CLKBUFX1 gbuf_d_1404(.A(gbuf206), .Y(d_out_1404));
CLKBUFX1 gbuf_qn_1404(.A(qn_in_1404), .Y(g2641));
INVX1 g67844(.A (n_699), .Y (n_597));
CLKBUFX1 gbuf_d_1405(.A(n_337), .Y(d_out_1405));
CLKBUFX1 gbuf_q_1405(.A(q_in_1405), .Y(gbuf126));
CLKBUFX1 gbuf_d_1406(.A(gbuf185), .Y(d_out_1406));
CLKBUFX1 gbuf_q_1406(.A(q_in_1406), .Y(g2426));
INVX1 g67829(.A (n_478), .Y (n_603));
CLKBUFX1 gbuf_d_1407(.A(gbuf142), .Y(d_out_1407));
CLKBUFX1 gbuf_qn_1407(.A(qn_in_1407), .Y(g1762));
CLKBUFX1 gbuf_d_1408(.A(n_364), .Y(d_out_1408));
CLKBUFX1 gbuf_q_1408(.A(q_in_1408), .Y(gbuf132));
CLKBUFX1 gbuf_d_1409(.A(gbuf86), .Y(d_out_1409));
CLKBUFX1 gbuf_q_1409(.A(q_in_1409), .Y(g1036));
CLKBUFX1 gbuf_d_1410(.A(gbuf59), .Y(d_out_1410));
CLKBUFX1 gbuf_qn_1410(.A(qn_in_1410), .Y(g567));
CLKBUFX1 gbuf_d_1411(.A(gbuf153), .Y(d_out_1411));
CLKBUFX1 gbuf_qn_1411(.A(qn_in_1411), .Y(g1949));
CLKBUFX1 gbuf_d_1412(.A(gbuf47), .Y(d_out_1412));
CLKBUFX1 gbuf_q_1412(.A(q_in_1412), .Y(g396));
CLKBUFX1 gbuf_d_1413(.A(gbuf186), .Y(d_out_1413));
CLKBUFX1 gbuf_q_1413(.A(q_in_1413), .Y(g2428));
CLKBUFX1 gbuf_d_1414(.A(gbuf38), .Y(d_out_1414));
CLKBUFX1 gbuf_q_1414(.A(q_in_1414), .Y(g_27919));
CLKBUFX1 gbuf_d_1415(.A(gbuf93), .Y(d_out_1415));
CLKBUFX1 gbuf_qn_1415(.A(qn_in_1415), .Y(g1068));
CLKBUFX1 gbuf_d_1416(.A(gbuf55), .Y(d_out_1416));
CLKBUFX1 gbuf_qn_1416(.A(qn_in_1416), .Y(g569));
CLKBUFX1 gbuf_d_1417(.A(gbuf195), .Y(d_out_1417));
CLKBUFX1 gbuf_q_1417(.A(q_in_1417), .Y(g2399));
CLKBUFX1 gbuf_d_1418(.A(gbuf104), .Y(d_out_1418));
CLKBUFX1 gbuf_qn_1418(.A(qn_in_1418), .Y(g1255));
CLKBUFX1 gbuf_d_1419(.A(gbuf202), .Y(d_out_1419));
CLKBUFX1 gbuf_qn_1419(.A(qn_in_1419), .Y(g2643));
CLKBUFX1 gbuf_d_1420(.A(gbuf156), .Y(d_out_1420));
CLKBUFX1 gbuf_q_1420(.A(q_in_1420), .Y(g1945));
NAND2X1 g67941(.A (n_476), .B (g2883), .Y (n_477));
NAND2X1 g68012(.A (n_321), .B (g_18792), .Y (n_475));
NAND3X1 g68055(.A (n_473), .B (g1501), .C (n_471), .Y (n_474));
XOR2X1 g68068(.A (n_458), .B (g3080), .Y (n_470));
INVX1 g68142(.A (n_656), .Y (n_762));
INVX1 g68295(.A (n_468), .Y (n_4110));
CLKBUFX1 gbuf_d_1421(.A(gbuf192), .Y(d_out_1421));
CLKBUFX1 gbuf_q_1421(.A(q_in_1421), .Y(g2458));
INVX1 g68455(.A (n_466), .Y (n_733));
NOR2X1 g68544(.A (n_264), .B (g3207), .Y (n_631));
CLKBUFX1 gbuf_d_1422(.A(gbuf43), .Y(d_out_1422));
CLKBUFX1 gbuf_qn_1422(.A(qn_in_1422), .Y(g_16164));
INVX1 g68504(.A (n_465), .Y (n_525));
CLKBUFX1 gbuf_d_1423(.A(gbuf96), .Y(d_out_1423));
CLKBUFX1 gbuf_qn_1423(.A(qn_in_1423), .Y(g1083));
CLKBUFX1 gbuf_d_1424(.A(g2873), .Y(d_out_1424));
CLKBUFX1 gbuf_q_1424(.A(q_in_1424), .Y(gbuf85));
CLKBUFX1 gbuf_d_1425(.A(gbuf60), .Y(d_out_1425));
CLKBUFX1 gbuf_q_1425(.A(q_in_1425), .Y(g489));
CLKBUFX1 gbuf_d_1426(.A(gbuf145), .Y(d_out_1426));
CLKBUFX1 gbuf_qn_1426(.A(qn_in_1426), .Y(g1777));
CLKBUFX1 gbuf_d_1427(.A(gbuf187), .Y(d_out_1427));
CLKBUFX1 gbuf_qn_1427(.A(qn_in_1427), .Y(g2439));
CLKBUFX1 gbuf_d_1428(.A(gbuf193), .Y(d_out_1428));
CLKBUFX1 gbuf_qn_1428(.A(qn_in_1428), .Y(g2469));
AND2X1 g68007(.A (n_461), .B (g1211), .Y (n_537));
CLKBUFX1 gbuf_d_1429(.A(gbuf109), .Y(d_out_1429));
CLKBUFX1 gbuf_q_1429(.A(q_in_1429), .Y(g1176));
CLKBUFX1 gbuf_d_1430(.A(gbuf46), .Y(d_out_1430));
CLKBUFX1 gbuf_qn_1430(.A(qn_in_1430), .Y(g394));
NAND2X1 g68566(.A (n_343), .B (n_4639), .Y (n_460));
CLKBUFX1 gbuf_d_1431(.A(gbuf140), .Y(d_out_1431));
CLKBUFX1 gbuf_q_1431(.A(q_in_1431), .Y(g1749));
AOI21X1 g66582(.A0 (n_458), .A1 (g3080), .B0 (g2998), .Y (n_459));
CLKBUFX1 gbuf_d_1432(.A(gbuf41), .Y(d_out_1432));
CLKBUFX1 gbuf_qn_1432(.A(qn_in_1432), .Y(g_9473));
CLKBUFX1 gbuf_d_1433(.A(gbuf136), .Y(d_out_1433));
CLKBUFX1 gbuf_qn_1433(.A(qn_in_1433), .Y(g1732));
CLKBUFX1 gbuf_d_1434(.A(gbuf139), .Y(d_out_1434));
CLKBUFX1 gbuf_qn_1434(.A(qn_in_1434), .Y(g1747));
CLKBUFX1 gbuf_d_1435(.A(gbuf205), .Y(d_out_1435));
CLKBUFX1 gbuf_q_1435(.A(q_in_1435), .Y(g2639));
NAND4X1 g67235(.A (g3002), .B (n_206), .C (g2998), .D (n_215), .Y(n_455));
INVX1 g68413(.A (g801), .Y (n_448));
INVX4 g68408(.A (g_18628), .Y (n_562));
NAND2X1 g67845(.A (n_236), .B (n_433), .Y (n_699));
NOR2X1 g67830(.A (n_442), .B (n_100), .Y (n_478));
INVX1 g68371(.A (g113), .Y (n_5247));
INVX1 g68282(.A (g_24889), .Y (g5629));
INVX1 g68313(.A (g_20137), .Y (n_1498));
INVX1 g68220(.A (g805), .Y (n_496));
NAND3X1 g68004(.A (n_433), .B (n_47), .C (g3197), .Y (n_803));
INVX1 g68590(.A (n_373), .Y (n_431));
NOR2X1 g68555(.A (g3231), .B (g3136), .Y (n_8163));
INVX1 g68143(.A (g809), .Y (n_656));
NOR2X1 g68560(.A (n_411), .B (g3201), .Y (n_425));
INVX1 g68109(.A (g101), .Y (n_5380));
INVX1 g68284(.A (g8106), .Y (n_422));
INVX1 g68296(.A (g789), .Y (n_468));
INVX1 g68318(.A (g785), .Y (n_504));
BUFX3 g68430(.A (g_14726), .Y (n_6822));
INVX1 g68542(.A (n_1385), .Y (n_479));
NAND2X1 g68547(.A (n_418), .B (n_420), .Y (n_539));
OR2X1 g68550(.A (n_418), .B (n_420), .Y (n_419));
INVX1 g68551(.A (n_416), .Y (n_417));
NOR2X1 g68565(.A (n_4368), .B (n_8759), .Y (n_415));
NAND2X1 g68568(.A (n_600), .B (n_473), .Y (n_413));
OR2X1 g68577(.A (g3151), .B (g3147), .Y (n_412));
NOR2X1 g68581(.A (n_344), .B (n_411), .Y (n_536));
NOR2X1 g68588(.A (g3201), .B (g3207), .Y (n_410));
INVX4 g68211(.A (g_21144), .Y (n_864));
INVX1 g68511(.A (g97), .Y (n_5382));
NAND3X1 g67994(.A (n_458), .B (g2998), .C (g3080), .Y (n_456));
INVX1 g68505(.A (g797), .Y (n_465));
INVX1 g68121(.A (g813), .Y (n_763));
INVX1 g68138(.A (g5657), .Y (n_404));
INVX1 g68492(.A (g121), .Y (n_5473));
INVX4 g68132(.A (g_24459), .Y (n_1245));
INVX1 g68973(.A (g2170), .Y (n_2809));
INVX1 g68536(.A (g793), .Y (n_3171));
INVX1 g68456(.A (g117), .Y (n_466));
INVX1 g68418(.A (g_32166), .Y (g5695));
INVX1 g68380(.A (g125), .Y (n_467));
CLKBUFX1 gbuf_d_1436(.A(g1075), .Y(d_out_1436));
CLKBUFX1 gbuf_q_1436(.A(q_in_1436), .Y(gbuf96));
CLKBUFX1 gbuf_d_1437(.A(g4590), .Y(d_out_1437));
CLKBUFX1 gbuf_q_1437(.A(q_in_1437), .Y(g801));
CLKBUFX1 gbuf_d_1438(.A(n_389), .Y(d_out_1438));
CLKBUFX1 gbuf_q_1438(.A(q_in_1438), .Y(gbuf158));
CLKBUFX1 gbuf_d_1439(.A(g2429), .Y(d_out_1439));
CLKBUFX1 gbuf_q_1439(.A(q_in_1439), .Y(gbuf184));
CLKBUFX1 gbuf_d_1440(.A(g1030), .Y(d_out_1440));
CLKBUFX1 gbuf_q_1440(.A(q_in_1440), .Y(gbuf87));
CLKBUFX1 gbuf_d_1441(.A(g1060), .Y(d_out_1441));
CLKBUFX1 gbuf_q_1441(.A(q_in_1441), .Y(gbuf93));
CLKBUFX1 gbuf_d_1442(.A(g16437), .Y(d_out_1442));
CLKBUFX1 gbuf_q_1442(.A(q_in_1442), .Y(g2599));
CLKBUFX1 gbuf_d_1443(.A(g8249), .Y(d_out_1443));
CLKBUFX1 gbuf_q_1443(.A(q_in_1443), .Y(g125));
AND2X1 g68579(.A (n_357), .B (n_264), .Y (n_712));
AND2X1 g68548(.A (g3032), .B (n_116), .Y (n_386));
CLKBUFX1 gbuf_d_1444(.A(g3080), .Y(d_out_1444));
CLKBUFX1 gbuf_q_1444(.A(q_in_1444), .Y(g8106));
CLKBUFX1 gbuf_d_1445(.A(g3226), .Y(d_out_1445));
CLKBUFX1 gbuf_q_1445(.A(q_in_1445), .Y(g2941));
CLKBUFX1 gbuf_d_1446(.A(g7334), .Y(d_out_1446));
CLKBUFX1 gbuf_qn_1446(.A(qn_in_1446), .Y(g785));
CLKBUFX1 gbuf_d_1447(.A(n_3), .Y(d_out_1447));
CLKBUFX1 gbuf_q_1447(.A(q_in_1447), .Y(gbuf156));
CLKBUFX1 gbuf_d_1448(.A(g3221), .Y(d_out_1448));
CLKBUFX1 gbuf_q_1448(.A(q_in_1448), .Y(g2959));
CLKBUFX1 gbuf_d_1449(.A(g3080), .Y(d_out_1449));
CLKBUFX1 gbuf_q_1449(.A(q_in_1449), .Y(g_20137));
CLKBUFX1 gbuf_d_1450(.A(g16297), .Y(d_out_1450));
CLKBUFX1 gbuf_q_1450(.A(q_in_1450), .Y(g_18792));
CLKBUFX1 gbuf_d_1451(.A(g1085), .Y(d_out_1451));
CLKBUFX1 gbuf_q_1451(.A(q_in_1451), .Y(gbuf95));
CLKBUFX1 gbuf_d_1452(.A(g3214), .Y(d_out_1452));
CLKBUFX1 gbuf_q_1452(.A(q_in_1452), .Y(g2981));
CLKBUFX1 gbuf_d_1453(.A(g1739), .Y(d_out_1453));
CLKBUFX1 gbuf_q_1453(.A(q_in_1453), .Y(gbuf139));
CLKBUFX1 gbuf_d_1454(.A(g2436), .Y(d_out_1454));
CLKBUFX1 gbuf_q_1454(.A(q_in_1454), .Y(gbuf189));
CLKBUFX1 gbuf_d_1455(.A(g1071), .Y(d_out_1455));
CLKBUFX1 gbuf_q_1455(.A(q_in_1455), .Y(gbuf92));
CLKBUFX1 gbuf_d_1456(.A(n_384), .Y(d_out_1456));
CLKBUFX1 gbuf_q_1456(.A(q_in_1456), .Y(gbuf104));
CLKBUFX1 gbuf_d_1457(.A(g1041), .Y(d_out_1457));
CLKBUFX1 gbuf_q_1457(.A(q_in_1457), .Y(gbuf86));
CLKBUFX1 gbuf_d_1458(.A(g1048), .Y(d_out_1458));
CLKBUFX1 gbuf_q_1458(.A(q_in_1458), .Y(gbuf91));
CLKBUFX1 gbuf_d_1459(.A(g3080), .Y(d_out_1459));
CLKBUFX1 gbuf_qn_1459(.A(qn_in_1459), .Y(g_24889));
CLKBUFX1 gbuf_d_1460(.A(g3213), .Y(d_out_1460));
CLKBUFX1 gbuf_q_1460(.A(q_in_1460), .Y(g2874));
CLKBUFX1 gbuf_d_1461(.A(g1742), .Y(d_out_1461));
CLKBUFX1 gbuf_q_1461(.A(q_in_1461), .Y(gbuf140));
CLKBUFX1 gbuf_d_1462(.A(g3080), .Y(d_out_1462));
CLKBUFX1 gbuf_q_1462(.A(q_in_1462), .Y(g5747));
CLKBUFX1 gbuf_d_1463(.A(g3216), .Y(d_out_1463));
CLKBUFX1 gbuf_q_1463(.A(q_in_1463), .Y(g2975));
CLKBUFX1 gbuf_d_1464(.A(g2451), .Y(d_out_1464));
CLKBUFX1 gbuf_q_1464(.A(q_in_1464), .Y(gbuf192));
NOR2X1 g68543(.A (g3230), .B (n_55), .Y (n_1385));
CLKBUFX1 gbuf_d_1465(.A(g1772), .Y(d_out_1465));
CLKBUFX1 gbuf_q_1465(.A(q_in_1465), .Y(gbuf146));
INVX1 g68647(.A (n_482), .Y (n_2706));
CLKBUFX1 gbuf_d_1466(.A(g1754), .Y(d_out_1466));
CLKBUFX1 gbuf_q_1466(.A(q_in_1466), .Y(gbuf142));
CLKBUFX1 gbuf_d_1467(.A(g346), .Y(d_out_1467));
CLKBUFX1 gbuf_q_1467(.A(q_in_1467), .Y(gbuf39));
CLKBUFX1 gbuf_d_1468(.A(n_378), .Y(d_out_1468));
CLKBUFX1 gbuf_q_1468(.A(q_in_1468), .Y(gbuf55));
OR2X1 g68546(.A (g3231), .B (n_111), .Y (n_1381));
AND2X1 g68564(.A (n_300), .B (n_377), .Y (n_501));
CLKBUFX1 gbuf_d_1469(.A(n_376), .Y(d_out_1469));
CLKBUFX1 gbuf_q_1469(.A(q_in_1469), .Y(gbuf153));
CLKBUFX1 gbuf_d_1470(.A(g3225), .Y(d_out_1470));
CLKBUFX1 gbuf_q_1470(.A(q_in_1470), .Y(g2944));
CLKBUFX1 gbuf_d_1471(.A(g51), .Y(d_out_1471));
CLKBUFX1 gbuf_q_1471(.A(q_in_1471), .Y(g8021));
CLKBUFX1 gbuf_d_1472(.A(g8175), .Y(d_out_1472));
CLKBUFX1 gbuf_q_1472(.A(q_in_1472), .Y(g109));
NOR2X1 g68556(.A (g3032), .B (n_116), .Y (n_375));
CLKBUFX1 gbuf_d_1473(.A(n_121), .Y(d_out_1473));
CLKBUFX1 gbuf_q_1473(.A(q_in_1473), .Y(gbuf205));
CLKBUFX1 gbuf_d_1474(.A(g16399), .Y(d_out_1474));
CLKBUFX1 gbuf_q_1474(.A(q_in_1474), .Y(g1905));
CLKBUFX1 gbuf_d_1475(.A(g2421), .Y(d_out_1475));
CLKBUFX1 gbuf_q_1475(.A(q_in_1475), .Y(gbuf186));
CLKBUFX1 gbuf_d_1476(.A(g2473), .Y(d_out_1476));
CLKBUFX1 gbuf_q_1476(.A(q_in_1476), .Y(gbuf193));
CLKBUFX1 gbuf_d_1477(.A(g3993), .Y(d_out_1477));
CLKBUFX1 gbuf_qn_1477(.A(qn_in_1477), .Y(g105));
CLKBUFX1 gbuf_d_1478(.A(g3080), .Y(d_out_1478));
CLKBUFX1 gbuf_q_1478(.A(q_in_1478), .Y(g_21144));
CLKBUFX1 gbuf_d_1479(.A(g391), .Y(d_out_1479));
CLKBUFX1 gbuf_q_1479(.A(q_in_1479), .Y(gbuf48));
CLKBUFX1 gbuf_d_1480(.A(g376), .Y(d_out_1480));
CLKBUFX1 gbuf_q_1480(.A(q_in_1480), .Y(gbuf45));
CLKBUFX1 gbuf_d_1481(.A(n_374), .Y(d_out_1481));
CLKBUFX1 gbuf_q_1481(.A(q_in_1481), .Y(gbuf183));
CLKBUFX1 gbuf_d_1482(.A(g3228), .Y(d_out_1482));
CLKBUFX1 gbuf_q_1482(.A(q_in_1482), .Y(g2935));
NAND2X1 g68591(.A (n_418), .B (n_260), .Y (n_373));
CLKBUFX1 gbuf_d_1483(.A(g2466), .Y(d_out_1483));
CLKBUFX1 gbuf_q_1483(.A(q_in_1483), .Y(gbuf195));
CLKBUFX1 gbuf_d_1484(.A(n_372), .Y(d_out_1484));
CLKBUFX1 gbuf_q_1484(.A(q_in_1484), .Y(gbuf154));
CLKBUFX1 gbuf_d_1485(.A(g1727), .Y(d_out_1485));
CLKBUFX1 gbuf_q_1485(.A(q_in_1485), .Y(gbuf137));
CLKBUFX1 gbuf_d_1486(.A(g1056), .Y(d_out_1486));
CLKBUFX1 gbuf_q_1486(.A(q_in_1486), .Y(gbuf89));
CLKBUFX1 gbuf_d_1487(.A(g1063), .Y(d_out_1487));
CLKBUFX1 gbuf_q_1487(.A(q_in_1487), .Y(gbuf94));
CLKBUFX1 gbuf_d_1488(.A(n_370), .Y(d_out_1488));
CLKBUFX1 gbuf_q_1488(.A(q_in_1488), .Y(gbuf202));
CLKBUFX1 gbuf_d_1489(.A(g1045), .Y(d_out_1489));
CLKBUFX1 gbuf_q_1489(.A(q_in_1489), .Y(gbuf90));
CLKBUFX1 gbuf_d_1490(.A(g3220), .Y(d_out_1490));
CLKBUFX1 gbuf_q_1490(.A(q_in_1490), .Y(g2963));
CLKBUFX1 gbuf_d_1491(.A(g373), .Y(d_out_1491));
CLKBUFX1 gbuf_q_1491(.A(q_in_1491), .Y(gbuf44));
CLKBUFX1 gbuf_d_1492(.A(g1769), .Y(d_out_1492));
CLKBUFX1 gbuf_q_1492(.A(q_in_1492), .Y(gbuf145));
CLKBUFX1 gbuf_d_1493(.A(g3080), .Y(d_out_1493));
CLKBUFX1 gbuf_q_1493(.A(q_in_1493), .Y(g5657));
CLKBUFX1 gbuf_d_1494(.A(g2433), .Y(d_out_1494));
CLKBUFX1 gbuf_q_1494(.A(q_in_1494), .Y(gbuf188));
CLKBUFX1 gbuf_d_1495(.A(g8096), .Y(d_out_1495));
CLKBUFX1 gbuf_q_1495(.A(q_in_1495), .Y(g2857));
CLKBUFX1 gbuf_d_1496(.A(g3215), .Y(d_out_1496));
CLKBUFX1 gbuf_q_1496(.A(q_in_1496), .Y(g2978));
CLKBUFX1 gbuf_d_1497(.A(g3232), .Y(d_out_1497));
CLKBUFX1 gbuf_q_1497(.A(q_in_1497), .Y(g2962));
CLKBUFX1 gbuf_d_1498(.A(n_10), .Y(d_out_1498));
CLKBUFX1 gbuf_q_1498(.A(q_in_1498), .Y(gbuf206));
CLKBUFX1 gbuf_d_1499(.A(g3080), .Y(d_out_1499));
CLKBUFX1 gbuf_q_1499(.A(q_in_1499), .Y(g_18412));
CLKBUFX1 gbuf_d_1500(.A(g8251), .Y(d_out_1500));
CLKBUFX1 gbuf_qn_1500(.A(qn_in_1500), .Y(g813));
NAND2X1 g68562(.A (n_166), .B (n_368), .Y (n_369));
CLKBUFX1 gbuf_d_1501(.A(g384), .Y(d_out_1501));
CLKBUFX1 gbuf_q_1501(.A(q_in_1501), .Y(gbuf43));
CLKBUFX1 gbuf_d_1502(.A(g2448), .Y(d_out_1502));
CLKBUFX1 gbuf_q_1502(.A(q_in_1502), .Y(gbuf191));
CLKBUFX1 gbuf_d_1503(.A(n_6), .Y(d_out_1503));
CLKBUFX1 gbuf_q_1503(.A(q_in_1503), .Y(gbuf59));
CLKBUFX1 gbuf_d_1504(.A(n_367), .Y(d_out_1504));
CLKBUFX1 gbuf_q_1504(.A(q_in_1504), .Y(gbuf57));
CLKBUFX1 gbuf_d_1505(.A(g1735), .Y(d_out_1505));
CLKBUFX1 gbuf_q_1505(.A(q_in_1505), .Y(gbuf135));
NOR2X1 g68582(.A (n_365), .B (n_364), .Y (n_366));
CLKBUFX1 gbuf_d_1506(.A(g358), .Y(d_out_1506));
CLKBUFX1 gbuf_q_1506(.A(q_in_1506), .Y(gbuf41));
CLKBUFX1 gbuf_d_1507(.A(g361), .Y(d_out_1507));
CLKBUFX1 gbuf_q_1507(.A(q_in_1507), .Y(gbuf42));
CLKBUFX1 gbuf_d_1508(.A(n_363), .Y(d_out_1508));
CLKBUFX1 gbuf_q_1508(.A(q_in_1508), .Y(gbuf203));
CLKBUFX1 gbuf_d_1509(.A(g3217), .Y(d_out_1509));
CLKBUFX1 gbuf_q_1509(.A(q_in_1509), .Y(g2972));
CLKBUFX1 gbuf_d_1510(.A(g1033), .Y(d_out_1510));
CLKBUFX1 gbuf_q_1510(.A(q_in_1510), .Y(gbuf88));
NAND2X1 g68552(.A (n_355), .B (g3207), .Y (n_416));
CLKBUFX1 gbuf_d_1511(.A(g4200), .Y(d_out_1511));
CLKBUFX1 gbuf_q_1511(.A(q_in_1511), .Y(g101));
CLKBUFX1 gbuf_d_1512(.A(g1078), .Y(d_out_1512));
CLKBUFX1 gbuf_q_1512(.A(q_in_1512), .Y(gbuf97));
CLKBUFX1 gbuf_d_1513(.A(g4090), .Y(d_out_1513));
CLKBUFX1 gbuf_qn_1513(.A(qn_in_1513), .Y(g809));
CLKBUFX1 gbuf_d_1514(.A(g4323), .Y(d_out_1514));
CLKBUFX1 gbuf_q_1514(.A(q_in_1514), .Y(g805));
CLKBUFX1 gbuf_d_1515(.A(n_360), .Y(d_out_1515));
CLKBUFX1 gbuf_q_1515(.A(q_in_1515), .Y(gbuf108));
CLKBUFX1 gbuf_d_1516(.A(g3080), .Y(d_out_1516));
CLKBUFX1 gbuf_q_1516(.A(q_in_1516), .Y(g_8082));
CLKBUFX1 gbuf_d_1517(.A(n_359), .Y(d_out_1517));
CLKBUFX1 gbuf_q_1517(.A(q_in_1517), .Y(gbuf105));
CLKBUFX1 gbuf_d_1518(.A(g369), .Y(d_out_1518));
CLKBUFX1 gbuf_q_1518(.A(q_in_1518), .Y(gbuf40));
CLKBUFX1 gbuf_d_1519(.A(g6895), .Y(d_out_1519));
CLKBUFX1 gbuf_qn_1519(.A(qn_in_1519), .Y(g789));
CLKBUFX1 gbuf_d_1520(.A(g7519), .Y(d_out_1520));
CLKBUFX1 gbuf_q_1520(.A(q_in_1520), .Y(g2873));
NOR2X1 g68549(.A (g2920), .B (n_358), .Y (n_476));
NOR2X1 g68553(.A (n_357), .B (g3207), .Y (n_569));
OR2X1 g68557(.A (n_355), .B (g3207), .Y (n_356));
CLKBUFX1 gbuf_d_1521(.A(g2463), .Y(d_out_1521));
CLKBUFX1 gbuf_q_1521(.A(q_in_1521), .Y(gbuf194));
CLKBUFX1 gbuf_d_1522(.A(g3222), .Y(d_out_1522));
CLKBUFX1 gbuf_q_1522(.A(q_in_1522), .Y(g2956));
CLKBUFX1 gbuf_d_1523(.A(g3218), .Y(d_out_1523));
CLKBUFX1 gbuf_q_1523(.A(q_in_1523), .Y(g2969));
CLKBUFX1 gbuf_d_1524(.A(g2444), .Y(d_out_1524));
CLKBUFX1 gbuf_q_1524(.A(q_in_1524), .Y(gbuf187));
CLKBUFX1 gbuf_d_1525(.A(n_352), .Y(d_out_1525));
CLKBUFX1 gbuf_q_1525(.A(q_in_1525), .Y(gbuf109));
CLKBUFX1 gbuf_d_1526(.A(g3224), .Y(d_out_1526));
CLKBUFX1 gbuf_q_1526(.A(q_in_1526), .Y(g2947));
CLKBUFX1 gbuf_d_1527(.A(g1779), .Y(d_out_1527));
CLKBUFX1 gbuf_q_1527(.A(q_in_1527), .Y(gbuf144));
CLKBUFX1 gbuf_d_1528(.A(g1724), .Y(d_out_1528));
CLKBUFX1 gbuf_q_1528(.A(q_in_1528), .Y(gbuf136));
CLKBUFX1 gbuf_d_1529(.A(g3227), .Y(d_out_1529));
CLKBUFX1 gbuf_q_1529(.A(q_in_1529), .Y(g2938));
CLKBUFX1 gbuf_d_1530(.A(g4450), .Y(d_out_1530));
CLKBUFX1 gbuf_q_1530(.A(q_in_1530), .Y(g97));
CLKBUFX1 gbuf_d_1531(.A(g6225), .Y(d_out_1531));
CLKBUFX1 gbuf_qn_1531(.A(qn_in_1531), .Y(g797));
CLKBUFX1 gbuf_d_1532(.A(g1750), .Y(d_out_1532));
CLKBUFX1 gbuf_q_1532(.A(q_in_1532), .Y(gbuf138));
CLKBUFX1 gbuf_d_1533(.A(g51), .Y(d_out_1533));
CLKBUFX1 gbuf_qn_1533(.A(qn_in_1533), .Y(g2814));
CLKBUFX1 gbuf_d_1534(.A(n_351), .Y(d_out_1534));
CLKBUFX1 gbuf_q_1534(.A(q_in_1534), .Y(gbuf107));
CLKBUFX1 gbuf_d_1535(.A(g3223), .Y(d_out_1535));
CLKBUFX1 gbuf_q_1535(.A(q_in_1535), .Y(g2953));
CLKBUFX1 gbuf_d_1536(.A(g8023), .Y(d_out_1536));
CLKBUFX1 gbuf_q_1536(.A(q_in_1536), .Y(g113));
CLKBUFX1 gbuf_d_1537(.A(g1757), .Y(d_out_1537));
CLKBUFX1 gbuf_q_1537(.A(q_in_1537), .Y(gbuf143));
CLKBUFX1 gbuf_d_1538(.A(n_350), .Y(d_out_1538));
CLKBUFX1 gbuf_q_1538(.A(q_in_1538), .Y(gbuf134));
CLKBUFX1 gbuf_d_1539(.A(n_349), .Y(d_out_1539));
CLKBUFX1 gbuf_q_1539(.A(q_in_1539), .Y(gbuf155));
CLKBUFX1 gbuf_d_1540(.A(g388), .Y(d_out_1540));
CLKBUFX1 gbuf_q_1540(.A(q_in_1540), .Y(gbuf47));
CLKBUFX1 gbuf_d_1541(.A(g3080), .Y(d_out_1541));
CLKBUFX1 gbuf_q_1541(.A(q_in_1541), .Y(g_24459));
CLKBUFX1 gbuf_d_1542(.A(g3080), .Y(d_out_1542));
CLKBUFX1 gbuf_q_1542(.A(q_in_1542), .Y(g_17832));
CLKBUFX1 gbuf_d_1543(.A(g4088), .Y(d_out_1543));
CLKBUFX1 gbuf_qn_1543(.A(qn_in_1543), .Y(g121));
CLKBUFX1 gbuf_d_1544(.A(n_348), .Y(d_out_1544));
CLKBUFX1 gbuf_q_1544(.A(q_in_1544), .Y(gbuf56));
CLKBUFX1 gbuf_d_1545(.A(n_80), .Y(d_out_1545));
CLKBUFX1 gbuf_q_1545(.A(q_in_1545), .Y(gbuf58));
CLKBUFX1 gbuf_d_1546(.A(g3212), .Y(d_out_1546));
CLKBUFX1 gbuf_q_1546(.A(q_in_1546), .Y(g2934));
INVX2 g69143(.A (n_377), .Y (n_4050));
CLKBUFX1 gbuf_d_1547(.A(g16355), .Y(d_out_1547));
CLKBUFX1 gbuf_q_1547(.A(q_in_1547), .Y(g1211));
CLKBUFX1 gbuf_d_1548(.A(g343), .Y(d_out_1548));
CLKBUFX1 gbuf_q_1548(.A(q_in_1548), .Y(gbuf38));
CLKBUFX1 gbuf_d_1549(.A(g2418), .Y(d_out_1549));
CLKBUFX1 gbuf_q_1549(.A(q_in_1549), .Y(gbuf185));
CLKBUFX1 gbuf_d_1550(.A(n_342), .Y(d_out_1550));
CLKBUFX1 gbuf_q_1550(.A(q_in_1550), .Y(gbuf207));
CLKBUFX1 gbuf_d_1551(.A(g398), .Y(d_out_1551));
CLKBUFX1 gbuf_q_1551(.A(q_in_1551), .Y(gbuf46));
CLKBUFX1 gbuf_d_1552(.A(g354), .Y(d_out_1552));
CLKBUFX1 gbuf_q_1552(.A(q_in_1552), .Y(gbuf37));
CLKBUFX1 gbuf_d_1553(.A(g6442), .Y(d_out_1553));
CLKBUFX1 gbuf_q_1553(.A(q_in_1553), .Y(g793));
CLKBUFX1 gbuf_d_1554(.A(n_58), .Y(d_out_1554));
CLKBUFX1 gbuf_q_1554(.A(q_in_1554), .Y(gbuf157));
CLKBUFX1 gbuf_d_1555(.A(g3219), .Y(d_out_1555));
CLKBUFX1 gbuf_q_1555(.A(q_in_1555), .Y(g2966));
CLKBUFX1 gbuf_d_1556(.A(n_339), .Y(d_out_1556));
CLKBUFX1 gbuf_q_1556(.A(q_in_1556), .Y(gbuf204));
CLKBUFX1 gbuf_d_1557(.A(g4321), .Y(d_out_1557));
CLKBUFX1 gbuf_q_1557(.A(q_in_1557), .Y(g117));
OR2X1 g68545(.A (g2883), .B (n_233), .Y (n_676));
CLKBUFX1 gbuf_d_1558(.A(g3080), .Y(d_out_1558));
CLKBUFX1 gbuf_qn_1558(.A(qn_in_1558), .Y(g_14726));
CLKBUFX1 gbuf_d_1559(.A(g3080), .Y(d_out_1559));
CLKBUFX1 gbuf_qn_1559(.A(qn_in_1559), .Y(g_32166));
CLKBUFX1 gbuf_d_1560(.A(g1765), .Y(d_out_1560));
CLKBUFX1 gbuf_q_1560(.A(q_in_1560), .Y(gbuf141));
CLKBUFX1 gbuf_d_1561(.A(n_338), .Y(d_out_1561));
CLKBUFX1 gbuf_q_1561(.A(q_in_1561), .Y(gbuf106));
INVX1 g68813(.A (n_473), .Y (n_337));
CLKBUFX1 gbuf_d_1562(.A(g2459), .Y(d_out_1562));
CLKBUFX1 gbuf_q_1562(.A(q_in_1562), .Y(gbuf190));
CLKBUFX1 gbuf_d_1563(.A(g3080), .Y(d_out_1563));
CLKBUFX1 gbuf_q_1563(.A(q_in_1563), .Y(g_18628));
CLKBUFX1 gbuf_d_1564(.A(n_336), .Y(d_out_1564));
CLKBUFX1 gbuf_q_1564(.A(q_in_1564), .Y(gbuf60));
INVX1 g69149(.A (n_368), .Y (n_679));
NAND2X1 g68574(.A (g2883), .B (n_379), .Y (n_442));
NAND2X1 g68567(.A (g2129), .B (g2133), .Y (n_289));
OR2X1 g68572(.A (g3010), .B (g3024), .Y (n_288));
NAND2X1 g68586(.A (g1332), .B (g1346), .Y (n_282));
NAND2X1 g68595(.A (g771), .B (g_17877), .Y (n_275));
NAND2X1 g68594(.A (g633), .B (g653), .Y (n_269));
INVX1 g69044(.A (n_418), .Y (n_268));
INVX1 g68636(.A (n_260), .Y (n_420));
NAND2X1 g68573(.A (g3013), .B (g3024), .Y (n_254));
NOR2X1 g68578(.A (g1243), .B (n_3698), .Y (n_461));
NOR2X1 g68592(.A (g1937), .B (n_5322), .Y (n_485));
NOR2X1 g68589(.A (g3198), .B (g3197), .Y (n_236));
NOR2X1 g68587(.A (g3191), .B (g3194), .Y (n_433));
NAND2X1 g68584(.A (g2720), .B (g2734), .Y (n_234));
NAND2X1 g68576(.A (g3002), .B (g3006), .Y (n_225));
NAND2X1 g68580(.A (g_21927), .B (g_26529), .Y (n_216));
NOR2X1 g68561(.A (g3006), .B (g3010), .Y (n_206));
INVX1 g68985(.A (g2190), .Y (n_385));
NAND2X1 g68571(.A (g2026), .B (g2040), .Y (n_187));
NAND2X1 g68570(.A (g1435), .B (g1439), .Y (n_183));
NOR2X1 g68569(.A (g2917), .B (g2912), .Y (n_986));
INVX1 g68863(.A (g1501), .Y (n_343));
NAND2X1 g68583(.A (g1457), .B (g1453), .Y (n_182));
INVX1 g68918(.A (g2185), .Y (n_2716));
NAND2X1 g68585(.A (g2151), .B (g2147), .Y (n_131));
INVX1 g69085(.A (g479), .Y (n_1141));
INVX1 g69058(.A (g267), .Y (n_139));
INVX1 g68633(.A (g2165), .Y (n_126));
INVX1 g68664(.A (g1636), .Y (n_125));
INVX1 g68734(.A (g936), .Y (n_157));
INVX1 g68754(.A (g927), .Y (n_317));
INVX1 g68823(.A (g2387), .Y (n_129));
INVX1 g69084(.A (g1158), .Y (n_352));
INVX1 g68662(.A (g2294), .Y (n_123));
INVX1 g68905(.A (g_18003), .Y (n_251));
INVX1 g68875(.A (n_344), .Y (n_357));
INVX1 g68857(.A (g_26724), .Y (n_917));
INVX1 g68949(.A (g3211), .Y (n_122));
INVX1 g69146(.A (g2584), .Y (n_377));
INVX1 g68752(.A (g3106), .Y (n_1171));
INVX1 g68921(.A (n_782), .Y (n_180));
INVX1 g68621(.A (g1633), .Y (n_843));
INVX1 g68981(.A (g1869), .Y (n_1136));
INVX1 g68691(.A (g2540), .Y (n_121));
INVX1 g68884(.A (g2552), .Y (n_3978));
INVX1 g68948(.A (g3112), .Y (n_120));
INVX1 g69091(.A (g2546), .Y (n_342));
INVX1 g68896(.A (g_30665), .Y (n_726));
INVX1 g69001(.A (g960), .Y (n_118));
INVX1 g68721(.A (g3099), .Y (n_117));
INVX1 g68870(.A (g2115), .Y (n_1557));
INVX1 g68712(.A (g2568), .Y (n_167));
INVX1 g68800(.A (g3028), .Y (n_116));
INVX1 g69078(.A (g_25929), .Y (n_971));
INVX1 g69080(.A (n_3143), .Y (n_213));
INVX1 g69022(.A (g1860), .Y (n_1093));
INVX1 g69137(.A (g2261), .Y (n_303));
INVX1 g68638(.A (g2539), .Y (n_836));
INVX1 g69116(.A (g2267), .Y (n_239));
INVX1 g68898(.A (g2312), .Y (n_113));
INVX1 g68824(.A (g2303), .Y (n_112));
INVX1 g68654(.A (g2554), .Y (n_845));
INVX1 g68616(.A (n_379), .Y (n_233));
INVX1 g68997(.A (g3139), .Y (n_111));
INVX1 g68968(.A (g2682), .Y (n_132));
INVX1 g69027(.A (g2321), .Y (n_176));
INVX1 g68902(.A (n_600), .Y (n_293));
INVX1 g68977(.A (g1180), .Y (n_108));
INVX1 g68907(.A (g_9172), .Y (n_5825));
INVX1 g69090(.A (g942), .Y (n_107));
INVX1 g68781(.A (g918), .Y (n_322));
INVX1 g69004(.A (g548), .Y (n_106));
INVX1 g68808(.A (g1145), .Y (n_359));
INVX1 g69038(.A (g1627), .Y (n_143));
INVX1 g68751(.A (g879), .Y (n_105));
INVX1 g68619(.A (g2348), .Y (n_255));
INVX1 g68643(.A (g1294), .Y (n_1466));
INVX1 g68655(.A (g900), .Y (n_104));
INVX1 g68777(.A (g2628), .Y (n_103));
INVX1 g69107(.A (g2270), .Y (n_271));
INVX1 g68858(.A (g2380), .Y (n_101));
INVX1 g68970(.A (g2664), .Y (n_170));
INVX1 g69141(.A (g_19110), .Y (n_222));
INVX1 g68706(.A (g930), .Y (n_1768));
INVX1 g68853(.A (g2888), .Y (n_100));
INVX1 g68676(.A (g1579), .Y (n_1956));
INVX1 g68894(.A (g1615), .Y (n_758));
INVX1 g68656(.A (g903), .Y (n_99));
INVX1 g68877(.A (g1000), .Y (n_141));
INVX1 g68598(.A (g264), .Y (n_98));
INVX1 g68624(.A (g2309), .Y (n_799));
INVX1 g69100(.A (g945), .Y (n_278));
INVX1 g68833(.A (g3105), .Y (n_1170));
INVX1 g68844(.A (g_28592), .Y (n_97));
INVX1 g68663(.A (g2877), .Y (n_350));
INVX1 g69109(.A (n_517), .Y (n_166));
INVX1 g68809(.A (g255), .Y (n_96));
INVX1 g68821(.A (g2533), .Y (n_363));
INVX1 g68774(.A (g1285), .Y (n_231));
INVX1 g68831(.A (g2082), .Y (n_95));
INVX1 g68789(.A (g_24437), .Y (n_94));
INVX1 g68693(.A (g2333), .Y (n_93));
INVX1 g68740(.A (g1845), .Y (n_1131));
INVX1 g68739(.A (g2878), .Y (n_374));
INVX1 g68741(.A (g3103), .Y (n_911));
INVX1 g68779(.A (g2694), .Y (n_91));
INVX1 g69032(.A (g234), .Y (n_931));
INVX1 g69121(.A (g1693), .Y (n_276));
INVX1 g69069(.A (g933), .Y (n_89));
INVX1 g68709(.A (g3134), .Y (n_88));
INVX1 g69110(.A (g_15687), .Y (n_87));
INVX1 g69128(.A (g3201), .Y (n_264));
INVX1 g69071(.A (g2306), .Y (n_86));
INVX1 g68661(.A (g611), .Y (n_84));
INVX1 g68669(.A (g261), .Y (n_83));
INVX1 g69048(.A (g921), .Y (n_1878));
INVX1 g68657(.A (g897), .Y (n_81));
INVX1 g68681(.A (g465), .Y (n_80));
INVX1 g68846(.A (g1476), .Y (n_79));
INVX1 g68732(.A (g_26067), .Y (n_319));
INVX1 g69019(.A (g1481), .Y (n_78));
INVX1 g68883(.A (g608), .Y (n_1501));
INVX1 g68938(.A (g557), .Y (n_77));
INVX1 g69060(.A (g1988), .Y (n_1469));
INVX1 g68866(.A (g3107), .Y (n_7712));
INVX1 g69135(.A (n_3698), .Y (n_645));
INVX1 g68690(.A (g1591), .Y (n_76));
INVX1 g68820(.A (g2536), .Y (n_339));
INVX1 g69034(.A (g1594), .Y (n_211));
INVX1 g68737(.A (g2330), .Y (n_75));
INVX1 g68786(.A (g1585), .Y (n_328));
INVX1 g68811(.A (g1654), .Y (n_209));
INVX1 g68689(.A (g599), .Y (n_298));
INVX1 g68735(.A (g458), .Y (n_348));
INVX1 g68819(.A (g882), .Y (n_153));
INVX1 g68697(.A (g1128), .Y (n_301));
INVX1 g68680(.A (g1651), .Y (n_834));
INVX1 g69029(.A (g_30245), .Y (n_237));
INVX1 g69156(.A (g243), .Y (n_933));
INVX1 g68926(.A (g258), .Y (n_247));
INVX1 g69112(.A (g954), .Y (n_137));
INVX1 g68666(.A (blif_reset_net), .Y (n_8183));
INVX1 g68635(.A (g2327), .Y (n_806));
INVX1 g68806(.A (g3142), .Y (n_296));
INVX1 g68719(.A (g3234), .Y (n_310));
INVX1 g69081(.A (g1597), .Y (n_72));
INVX1 g68798(.A (g1486), .Y (n_454));
INVX1 g69089(.A (n_3203), .Y (n_163));
INVX1 g68695(.A (g_20070), .Y (n_220));
INVX1 g68993(.A (g1836), .Y (n_376));
INVX1 g69148(.A (g957), .Y (n_1884));
INVX1 g68745(.A (g2088), .Y (n_70));
INVX1 g68597(.A (g2637), .Y (n_69));
INVX1 g69117(.A (g924), .Y (n_68));
INVX1 g68759(.A (n_471), .Y (n_4639));
INVX1 g68890(.A (g455), .Y (n_378));
INVX1 g68839(.A (g1852), .Y (n_389));
INVX1 g68641(.A (g1603), .Y (n_286));
INVX1 g68660(.A (g_22538), .Y (n_297));
INVX1 g68828(.A (g1119), .Y (n_67));
INVX1 g68750(.A (g1303), .Y (n_66));
INVX1 g68951(.A (g2114), .Y (n_2525));
INVX1 g68784(.A (g3151), .Y (n_324));
INVX1 g69132(.A (g2339), .Y (n_64));
INVX1 g69043(.A (g3104), .Y (n_1197));
INVX1 g68678(.A (g2282), .Y (n_1900));
INVX1 g68892(.A (g2924), .Y (n_358));
INVX1 g68701(.A (n_655), .Y (n_300));
INVX1 g69068(.A (g1582), .Y (n_207));
INVX1 g68738(.A (g3111), .Y (n_63));
INVX1 g69119(.A (g888), .Y (n_266));
INVX1 g69041(.A (g3132), .Y (n_62));
INVX1 g68653(.A (n_5322), .Y (n_659));
INVX1 g68765(.A (g461), .Y (n_367));
INVX2 g69045(.A (g2900), .Y (n_418));
INVX1 g68692(.A (g1639), .Y (n_61));
INVX1 g69075(.A (g3136), .Y (n_185));
INVX1 g69142(.A (g1240), .Y (n_3611));
INVX1 g68906(.A (g_18564), .Y (n_5741));
INVX1 g69009(.A (g948), .Y (n_60));
INVX1 g68888(.A (g894), .Y (n_1875));
INVX1 g68889(.A (g1874), .Y (n_59));
INVX1 g68743(.A (g1849), .Y (n_58));
INVX1 g69040(.A (g2264), .Y (n_942));
INVX1 g68746(.A (g1859), .Y (n_56));
INVX1 g69011(.A (g_13736), .Y (n_749));
INVX1 g68923(.A (g1630), .Y (n_249));
INVX1 g68928(.A (g1164), .Y (n_313));
INVX1 g68879(.A (g1624), .Y (n_841));
INVX1 g69021(.A (g2297), .Y (n_283));
INVX1 g69097(.A (g2175), .Y (n_436));
INVX1 g68639(.A (g3233), .Y (n_55));
INVX1 g69139(.A (g1107), .Y (n_198));
INVX1 g68807(.A (g464), .Y (n_1112));
INVX1 g68601(.A (g1609), .Y (n_54));
INVX1 g68775(.A (g2085), .Y (n_53));
INVX1 g68776(.A (g951), .Y (n_52));
INVX1 g69113(.A (g1858), .Y (n_4419));
INVX1 g68687(.A (n_411), .Y (n_355));
INVX1 g68604(.A (g2252), .Y (n_332));
INVX1 g68673(.A (g885), .Y (n_1873));
INVX1 g69152(.A (g_29227), .Y (n_5866));
INVX1 g69023(.A (g2285), .Y (n_51));
INVX1 g69105(.A (g939), .Y (n_1895));
INVX1 g68924(.A (g2276), .Y (n_48));
INVX1 g68914(.A (g1979), .Y (n_174));
INVX1 g68843(.A (g3108), .Y (n_1198));
INVX1 g68827(.A (g3198), .Y (n_47));
INVX1 g68637(.A (g2908), .Y (n_260));
INVX1 g68909(.A (g_27975), .Y (n_45));
INVX1 g68851(.A (g1476), .Y (n_364));
INVX1 g68908(.A (g1645), .Y (n_44));
INVX1 g68764(.A (g891), .Y (n_155));
INVX1 g68978(.A (g_32037), .Y (n_43));
INVX1 g68885(.A (g_29095), .Y (n_42));
INVX1 g68958(.A (g1642), .Y (n_39));
INVX1 g68940(.A (g590), .Y (n_147));
INVX1 g68600(.A (g1600), .Y (n_38));
INVX1 g68838(.A (g2691), .Y (n_151));
INVX1 g69036(.A (g1098), .Y (n_37));
INVX1 g69066(.A (g1573), .Y (n_334));
INVX1 g68868(.A (g2685), .Y (n_36));
INVX1 g68744(.A (g1839), .Y (n_372));
INVX1 g68865(.A (g3113), .Y (n_35));
INVX1 g68599(.A (g3128), .Y (n_34));
INVX1 g68955(.A (g617), .Y (n_33));
INVX1 g69042(.A (g2920), .Y (n_32));
INVX1 g68632(.A (g2165), .Y (n_4368));
INVX1 g68766(.A (g2563), .Y (n_819));
INVX1 g68842(.A (g1249), .Y (n_31));
INVX1 g68886(.A (g1151), .Y (n_1145));
INVX1 g69150(.A (g2896), .Y (n_368));
INVX1 g68966(.A (g1471), .Y (n_365));
INVX1 g69025(.A (g1570), .Y (n_830));
INVX1 g69000(.A (g_16638), .Y (n_172));
INVX1 g69008(.A (g1621), .Y (n_202));
INVX1 g68859(.A (g563), .Y (n_30));
INVX1 g68788(.A (g2315), .Y (n_193));
INVX1 g68714(.A (g2300), .Y (n_1882));
INVX1 g69073(.A (g_27924), .Y (n_28));
INVX1 g68957(.A (g1588), .Y (n_1893));
INVX1 g68950(.A (g915), .Y (n_27));
INVX1 g69103(.A (g270), .Y (n_848));
INVX1 g68702(.A (g1934), .Y (n_26));
INVX1 g68762(.A (g1422), .Y (n_25));
INVX1 g68897(.A (g3127), .Y (n_24));
INVX1 g68742(.A (g554), .Y (n_23));
INVX1 g69101(.A (g2116), .Y (n_1503));
INVX1 g68792(.A (g1576), .Y (n_330));
INVX1 g69006(.A (g735), .Y (n_1816));
INVX1 g68622(.A (g736), .Y (n_1635));
INVX1 g68832(.A (g734), .Y (n_2847));
INVX1 g68736(.A (g2094), .Y (n_22));
INVX1 g68804(.A (g1421), .Y (n_21));
INVX1 g68710(.A (g1420), .Y (n_2540));
INVX1 g69005(.A (g2810), .Y (n_1600));
INVX1 g68959(.A (g2808), .Y (n_2973));
INVX1 g69076(.A (g1842), .Y (n_349));
INVX1 g68602(.A (g906), .Y (n_18));
INVX1 g69056(.A (g1612), .Y (n_17));
INVX1 g68708(.A (g1003), .Y (n_308));
INVX1 g68826(.A (g_17170), .Y (n_228));
INVX1 g68912(.A (g471), .Y (n_336));
INVX1 g69070(.A (g488), .Y (n_1101));
INVX1 g68932(.A (n_2834), .Y (n_245));
INVX1 g68995(.A (g_19223), .Y (n_241));
INVX1 g68980(.A (g2809), .Y (n_1568));
INVX1 g68596(.A (g237), .Y (n_14));
INVX1 g69035(.A (g1175), .Y (n_1125));
INVX1 g68771(.A (n_3701), .Y (n_321));
INVX1 g69083(.A (n_458), .Y (n_215));
INVX1 g68674(.A (g3123), .Y (n_12));
INVX1 g68704(.A (g252), .Y (n_936));
INVX1 g68626(.A (g2279), .Y (n_200));
INVX1 g68668(.A (g2345), .Y (n_796));
INVX1 g69072(.A (g2530), .Y (n_370));
INVX1 g69098(.A (g2175), .Y (n_11));
INVX1 g68852(.A (g1142), .Y (n_384));
INVX1 g68722(.A (g1166), .Y (n_1114));
INVX1 g68817(.A (g912), .Y (n_1841));
INVX1 g68952(.A (g2543), .Y (n_10));
INVX1 g68841(.A (g1606), .Y (n_1942));
INVX1 g68992(.A (g3036), .Y (n_9));
INVX1 g68867(.A (g2336), .Y (n_8));
INVX1 g68936(.A (g2673), .Y (n_294));
INVX1 g68998(.A (g1152), .Y (n_351));
INVX1 g68911(.A (g_18819), .Y (n_7));
INVX1 g68835(.A (g273), .Y (n_226));
INVX1 g68988(.A (g477), .Y (n_3971));
INVX1 g69114(.A (g468), .Y (n_6));
INVX1 g68665(.A (g2291), .Y (n_5));
INVX1 g68749(.A (g1618), .Y (n_4));
INVX1 g68934(.A (g312), .Y (n_149));
INVX1 g68748(.A (g909), .Y (n_315));
INVX1 g69018(.A (g1481), .Y (n_435));
INVX1 g68790(.A (g1846), .Y (n_3));
INVX1 g68729(.A (g2195), .Y (n_447));
INVX1 g68954(.A (g1558), .Y (n_189));
INVX1 g69154(.A (g1567), .Y (n_306));
INVX1 g68836(.A (g1148), .Y (n_338));
INVX1 g68881(.A (g2318), .Y (n_811));
INVX1 g68947(.A (g249), .Y (n_326));
INVX1 g69030(.A (g3135), .Y (n_2));
INVX1 g68830(.A (n_2880), .Y (n_2959));
INVX1 g68945(.A (g_22281), .Y (n_0));
INVX1 g68869(.A (g1155), .Y (n_360));
INVX1 g68942(.A (g2324), .Y (n_204));
CLKBUFX1 g70721(.A (n_9113), .Y (n_8281));
INVX1 g70734(.A (n_8305), .Y (g5472));
CLKBUFX1 g70755(.A (n_8718), .Y (n_8305));
INVX2 g70762(.A (n_8339), .Y (g6518));
CLKBUFX1 g70770(.A (n_8326), .Y (n_8339));
CLKBUFX3 g70771(.A (n_8351), .Y (n_8326));
CLKBUFX3 g70772(.A (n_8351), .Y (n_8346));
INVX1 g70774(.A (g_14662), .Y (n_8351));
INVX1 g70775(.A (g_14662), .Y (n_8353));
INVX1 g70776(.A (g_14662), .Y (n_8355));
CLKBUFX1 g70778(.A (n_9272), .Y (n_8357));
MX2X1 g54(.A (n_3171), .B (g793), .S0 (n_3650), .Y (n_8376));
INVX1 g61(.A (n_4267), .Y (n_8377));
NOR2X1 g57(.A (n_3825), .B (n_3815), .Y (n_8379));
NAND2X1 g55(.A (n_4031), .B (n_4034), .Y (n_8380));
NOR2X1 g56(.A (n_8492), .B (n_8497), .Y (n_8383));
NOR2X1 g31(.A (n_8387), .B (n_8393), .Y (n_8394));
OAI21X1 g38(.A0 (n_6413), .A1 (n_6414), .B0 (n_8386), .Y (n_8387));
NAND2X1 g41(.A (n_6413), .B (n_6414), .Y (n_8386));
NAND2X1 g33(.A (n_8389), .B (n_8392), .Y (n_8393));
INVX1 g43(.A (n_8388), .Y (n_8389));
NAND3X1 g37(.A (n_8703), .B (n_6316), .C (n_9570), .Y (n_8388));
OAI21X1 g39(.A0 (n_6413), .A1 (n_4206), .B0 (n_8391), .Y (n_8392));
NAND2X1 g40(.A (n_6413), .B (n_4206), .Y (n_8391));
CLKBUFX1 g1(.A (n_8394), .Y (n_8395));
OR2X1 g32(.A (n_8387), .B (n_8396), .Y (n_8397));
CLKBUFX1 g45(.A (n_8388), .Y (n_8396));
INVX1 g44(.A (n_8396), .Y (n_8398));
AOI21X1 g70781(.A0 (n_8404), .A1 (n_8408), .B0 (n_8409), .Y (n_8410));
AOI21X1 g70782(.A0 (n_8400), .A1 (n_8401), .B0 (n_8403), .Y (n_8404));
INVX2 g47(.A (n_8774), .Y (n_8400));
INVX1 g70783(.A (g876), .Y (n_8401));
AOI21X1 g70784(.A0 (n_8402), .A1 (g876), .B0 (g873), .Y (n_8403));
INVX1 g70785(.A (n_8351), .Y (n_8402));
INVX4 g70786(.A (n_8775), .Y (n_8408));
NOR2X1 g70789(.A (n_105), .B (n_4162), .Y (n_8409));
CLKBUFX1 g70790(.A (n_8410), .Y (n_8411));
INVX1 g70792(.A (g_13515), .Y (n_8413));
CLKBUFX1 g70793(.A (n_8784), .Y (n_8419));
CLKBUFX1 g20(.A (n_8785), .Y (n_8420));
NAND3X1 g70796(.A (n_1017), .B (n_2066), .C (n_3567), .Y (n_8421));
INVX1 g70797(.A (n_8422), .Y (n_8423));
CLKBUFX2 g70798(.A (n_4477), .Y (n_8422));
NAND2X1 g70799(.A (n_4641), .B (n_4642), .Y (n_8424));
NAND2X1 g70802(.A (n_8421), .B (n_8422), .Y (n_8427));
OR2X1 g35(.A (n_9136), .B (n_4339), .Y (n_8432));
NOR2X1 g70805(.A (n_8597), .B (n_8598), .Y (n_8437));
NAND2X1 g70816(.A (n_2443), .B (n_4178), .Y (n_8445));
INVX1 g70817(.A (n_1123), .Y (n_8446));
INVX2 g70822(.A (n_8461), .Y (n_8462));
NAND3X1 g70823(.A (n_8455), .B (n_8457), .C (n_8460), .Y (n_8461));
INVX2 g70824(.A (n_8454), .Y (n_8455));
NAND3X1 g70825(.A (n_9674), .B (n_6527), .C (n_6618), .Y (n_8454));
AOI21X1 g70826(.A0 (n_6602), .A1 (n_6603), .B0 (n_8456), .Y (n_8457));
NOR2X1 g70827(.A (n_6603), .B (n_6602), .Y (n_8456));
OAI21X1 g70828(.A0 (n_6602), .A1 (n_4596), .B0 (n_8459), .Y (n_8460));
NAND2X1 g70829(.A (n_6602), .B (n_4596), .Y (n_8459));
NAND2X1 g70831(.A (n_8457), .B (n_8455), .Y (n_8463));
CLKBUFX1 g70832(.A (n_8455), .Y (n_8464));
INVX2 g70838(.A (n_9366), .Y (n_8471));
NAND2X1 g70843(.A (n_2767), .B (n_4149), .Y (n_8472));
INVX1 g70844(.A (n_9426), .Y (n_8476));
NAND3X1 g70846(.A (n_9577), .B (n_9578), .C (n_8482), .Y (n_8483));
AOI21X1 g70847(.A0 (n_8861), .A1 (n_5963), .B0 (n_8478), .Y (n_9578));
AOI21X1 g70848(.A0 (n_5230), .A1 (n_5963), .B0 (n_8863), .Y (n_8478));
INVX1 g70849(.A (n_6975), .Y (n_9577));
NOR2X1 g70850(.A (n_8481), .B (n_6431), .Y (n_8482));
NOR2X1 g70851(.A (n_8862), .B (n_5231), .Y (n_8481));
AND2X1 g70852(.A (n_8484), .B (n_8486), .Y (n_8487));
NOR2X1 g70853(.A (n_6431), .B (n_6975), .Y (n_8484));
NOR2X1 g70854(.A (n_8481), .B (n_8485), .Y (n_8486));
NOR2X1 g70855(.A (n_5230), .B (n_8863), .Y (n_8485));
NOR2X1 g67(.A (n_8376), .B (n_8377), .Y (n_8488));
AOI21X1 g66(.A0 (n_3821), .A1 (g809), .B0 (n_8380), .Y (n_8489));
AOI21X1 g70857(.A0 (n_3815), .A1 (n_3825), .B0 (n_8493), .Y (n_8494));
AND2X1 g70858(.A (n_8490), .B (n_8492), .Y (n_8493));
NAND2X1 g68_dup(.A (n_3332), .B (n_2764), .Y (n_8490));
AOI21X1 g65_dup(.A0 (n_2384), .A1 (n_8408), .B0 (n_3051), .Y(n_8492));
NOR2X1 g69(.A (n_8383), .B (n_8379), .Y (n_8495));
NAND2X1 g68(.A (n_3332), .B (n_2764), .Y (n_8497));
INVX1 g62(.A (n_8498), .Y (n_8499));
AOI21X1 g65(.A0 (n_2384), .A1 (n_8408), .B0 (n_3051), .Y (n_8498));
AND2X1 g70861(.A (n_9560), .B (n_8876), .Y (n_9198));
INVX1 g70866(.A (n_8740), .Y (n_8515));
AOI21X1 g70870(.A0 (n_8968), .A1 (n_6726), .B0 (n_4528), .Y (n_8517));
NOR2X1 g70879(.A (n_9041), .B (n_9101), .Y (n_8527));
CLKBUFX1 g70883(.A (n_8842), .Y (n_8533));
CLKBUFX1 g70884(.A (n_8841), .Y (n_8534));
NOR2X1 g70885(.A (n_8540), .B (n_9063), .Y (n_8541));
NAND2X1 g70891(.A (n_6848), .B (n_9345), .Y (n_8540));
CLKBUFX1 g70892(.A (n_9061), .Y (n_8542));
CLKBUFX1 g23(.A (n_8656), .Y (n_8548));
INVX1 g59(.A (n_8551), .Y (n_8552));
INVX2 g70898(.A (n_8550), .Y (n_8551));
NAND2X2 g70899(.A (n_4478), .B (n_4295), .Y (n_8550));
NAND2X2 g70903(.A (n_4465), .B (n_4266), .Y (n_8557));
AOI22X1 g70904(.A0 (n_9021), .A1 (n_8566), .B0 (n_8570), .B1(n_9014), .Y (n_8571));
NAND2X1 g70907(.A (n_9670), .B (n_9669), .Y (n_8563));
OAI21X1 g70908(.A0 (n_6616), .A1 (n_4502), .B0 (n_5169), .Y (n_8566));
NAND2X1 g70909(.A (n_9655), .B (n_8567), .Y (n_8570));
NAND2X2 g70910(.A (n_6616), .B (n_6528), .Y (n_8567));
INVX1 g70914(.A (n_8567), .Y (n_8573));
NOR2X1 g70915(.A (n_8574), .B (n_8584), .Y (n_8585));
INVX1 g70916(.A (n_7751), .Y (n_8574));
NAND2X1 g70917(.A (n_8583), .B (n_9195), .Y (n_8584));
NAND2X1 g70918(.A (n_8575), .B (n_8582), .Y (n_8583));
AOI21X1 g70919(.A0 (n_8487), .A1 (n_5963), .B0 (n_7314), .Y (n_8575));
INVX2 g70920(.A (n_8874), .Y (n_8582));
NAND2X1 g70925(.A (n_6849), .B (n_6372), .Y (n_8576));
NAND3X1 g70926(.A (n_8187), .B (n_9273), .C (n_7891), .Y (n_8578));
NOR2X1 g70935(.A (n_3984), .B (n_9303), .Y (n_8590));
INVX1 g70936(.A (n_8432), .Y (n_8591));
INVX1 g70938(.A (n_8725), .Y (n_8597));
NAND2X1 g70939(.A (n_8726), .B (n_8722), .Y (n_8598));
CLKBUFX1 g70948(.A (n_9059), .Y (n_8607));
INVX2 g70953(.A (n_8608), .Y (n_8609));
NAND2X2 g70954(.A (n_3840), .B (n_3661), .Y (n_8608));
NAND2X2 g8(.A (n_8621), .B (n_8622), .Y (n_8623));
INVX1 g12(.A (g_17832), .Y (n_8621));
INVX1 g13(.A (g_9980), .Y (n_8622));
INVX2 g11(.A (g_17832), .Y (n_8625));
INVX2 g14(.A (g_9980), .Y (n_8626));
AOI21X1 g70963(.A0 (n_8628), .A1 (n_8629), .B0 (n_8633), .Y (n_8634));
NAND2X1 g70964(.A (n_7554), .B (n_7407), .Y (n_8628));
NAND2X1 g70965(.A (n_7030), .B (n_7466), .Y (n_8629));
INVX1 g30(.A (n_8632), .Y (n_8633));
NAND2X1 g70966(.A (n_8630), .B (n_8631), .Y (n_8632));
AND2X1 g70967(.A (n_7379), .B (n_7381), .Y (n_8630));
NAND2X2 g36(.A (n_6144), .B (n_7381), .Y (n_8631));
CLKBUFX1 g70968(.A (n_8631), .Y (n_8635));
INVX2 g34(.A (n_8631), .Y (n_8636));
OAI21X1 g70969(.A0 (n_1946), .A1 (n_5), .B0 (n_8640), .Y (n_8641));
AOI21X1 g70970(.A0 (n_8933), .A1 (g2288), .B0 (n_8639), .Y (n_8640));
NOR2X1 g25(.A (n_3224), .B (n_123), .Y (n_8639));
INVX1 g70974(.A (n_8933), .Y (n_8643));
AOI21X1 g70976(.A0 (n_8264), .A1 (n_8265), .B0 (n_3337), .Y (n_8644));
NAND2X1 g70978(.A (n_8720), .B (n_8646), .Y (n_8647));
INVX1 g70980(.A (n_2198), .Y (n_8646));
INVX1 g70981(.A (n_8649), .Y (n_8650));
OAI21X1 g70982(.A0 (n_8362), .A1 (n_2063), .B0 (n_3340), .Y (n_8649));
AND2X1 g70983(.A (n_8650), .B (n_9369), .Y (n_8652));
INVX4 g70984(.A (n_8650), .Y (n_8653));
NAND2X2 g70988(.A (n_9090), .B (n_6529), .Y (n_8655));
NAND2X2 g70989(.A (n_9071), .B (n_6529), .Y (n_8656));
NOR2X1 g70996(.A (n_9067), .B (n_5321), .Y (n_8663));
CLKBUFX1 g70998(.A (n_8770), .Y (n_8667));
NAND2X1 g71005(.A (n_9502), .B (n_8924), .Y (n_8678));
NAND4X1 g49(.A (n_8682), .B (n_8685), .C (n_8690), .D (n_9637), .Y(n_8693));
NOR2X1 g71007(.A (n_5463), .B (n_5026), .Y (n_8682));
INVX1 g71008(.A (n_8998), .Y (n_8685));
INVX1 g50(.A (n_8689), .Y (n_8690));
CLKBUFX1 g71011(.A (n_8688), .Y (n_8689));
NAND2X2 g71012(.A (n_8686), .B (n_8687), .Y (n_8688));
NAND3X1 g71013(.A (n_9055), .B (n_972), .C (n_2456), .Y (n_8686));
OR2X1 g71014(.A (n_241), .B (n_9314), .Y (n_8687));
AOI21X1 g71016(.A0 (n_9685), .A1 (n_9686), .B0 (n_4169), .Y (n_9640));
INVX1 g52(.A (n_8689), .Y (n_8694));
AND2X1 g71018(.A (n_8700), .B (n_8702), .Y (n_8703));
NOR2X1 g71019(.A (n_8699), .B (n_6187), .Y (n_8700));
OAI21X1 g71020(.A0 (n_5902), .A1 (n_8697), .B0 (n_8698), .Y (n_8699));
AND2X1 g71022(.A (n_5778), .B (n_4756), .Y (n_8697));
OR2X1 g71023(.A (n_5915), .B (n_4312), .Y (n_8698));
NOR2X1 g71024(.A (n_8701), .B (n_6652), .Y (n_8702));
NOR2X1 g71025(.A (n_4434), .B (n_5857), .Y (n_8701));
NAND3X1 g71026(.A (n_8704), .B (n_8705), .C (n_8698), .Y (n_8706));
NOR2X1 g71027(.A (n_6652), .B (n_6187), .Y (n_8704));
OR2X1 g71028(.A (n_5778), .B (n_5902), .Y (n_8705));
OR2X1 g71029(.A (n_8707), .B (n_8701), .Y (n_8708));
NOR2X1 g71030(.A (n_4756), .B (n_5902), .Y (n_8707));
NOR2X1 g71035(.A (n_4843), .B (n_5287), .Y (n_8710));
NAND2X1 g71040(.A (n_8718), .B (n_8719), .Y (n_8720));
INVX2 g9(.A (g_8360), .Y (n_8718));
INVX2 g10(.A (g_20180), .Y (n_8719));
NAND3X1 g71042(.A (n_8724), .B (n_8725), .C (n_8726), .Y (n_8727));
NOR2X1 g71043(.A (n_8721), .B (n_8723), .Y (n_8724));
NOR2X1 g71044(.A (n_9449), .B (n_9303), .Y (n_8721));
OAI21X1 g71045(.A0 (n_9136), .A1 (n_3812), .B0 (n_8722), .Y (n_8723));
AOI21X1 g71046(.A0 (n_9137), .A1 (n_8879), .B0 (n_6023), .Y (n_8722));
NOR2X1 g71047(.A (n_8591), .B (n_8590), .Y (n_8725));
NOR2X1 g71048(.A (n_6299), .B (n_6476), .Y (n_8726));
AND2X1 g71049(.A (n_8732), .B (n_8733), .Y (n_8734));
NOR2X1 g71050(.A (n_8731), .B (n_8886), .Y (n_8732));
OR2X1 g71051(.A (n_8730), .B (n_4240), .Y (n_8731));
CLKBUFX1 g71052(.A (n_8778), .Y (n_8730));
NOR2X1 g71054(.A (n_6653), .B (n_9137), .Y (n_8733));
INVX1 g71056(.A (n_8778), .Y (n_8736));
INVX1 g71063(.A (n_8740), .Y (n_8741));
OAI21X1 g71064(.A0 (n_2454), .A1 (n_9505), .B0 (n_3754), .Y (n_8740));
NOR2X1 g71065(.A (n_8445), .B (n_8446), .Y (n_8743));
CLKBUFX1 g71067(.A (n_9541), .Y (n_8747));
INVX2 g71076(.A (n_9397), .Y (n_8756));
AOI21X1 g71078(.A0 (n_2719), .A1 (n_3955), .B0 (n_8757), .Y (n_8758));
NOR2X1 g71079(.A (n_126), .B (n_4214), .Y (n_8757));
MX2X1 g71080(.A (n_8759), .B (g2170), .S0 (n_8760), .Y (n_8761));
INVX1 g71081(.A (g2170), .Y (n_8759));
NAND3X1 g71082(.A (n_1013), .B (n_3597), .C (n_2251), .Y (n_8760));
NAND2X1 g71083(.A (n_3956), .B (g2180), .Y (n_8762));
NAND2X1 g71084(.A (n_4214), .B (n_126), .Y (n_8764));
NAND4X1 g71085(.A (n_8768), .B (n_4919), .C (n_8663), .D (n_8769), .Y(n_8770));
NOR2X1 g71086(.A (n_8552), .B (n_8767), .Y (n_8768));
OR2X1 g71087(.A (n_8766), .B (n_9066), .Y (n_8767));
NAND2X2 g71088(.A (n_4466), .B (n_4273), .Y (n_8766));
NOR2X1 g71089(.A (n_8557), .B (n_9091), .Y (n_8769));
INVX1 g71091(.A (n_8766), .Y (n_8771));
AOI21X1 g71092(.A0 (n_9585), .A1 (n_9586), .B0 (n_8777), .Y (n_8778));
NAND2X1 g71093(.A (n_1997), .B (n_153), .Y (n_9586));
AOI21X1 g71094(.A0 (n_8413), .A1 (n_1873), .B0 (n_8775), .Y (n_9585));
NOR2X1 g71095(.A (g_14662), .B (n_8774), .Y (n_8775));
CLKBUFX2 g71096(.A (g_13515), .Y (n_8774));
NOR2X1 g71097(.A (n_266), .B (n_4162), .Y (n_8777));
NOR2X1 g71099(.A (n_9058), .B (n_8783), .Y (n_8784));
NOR2X1 g71101(.A (n_8781), .B (n_8782), .Y (n_8783));
INVX1 g71102(.A (n_6528), .Y (n_8781));
NOR2X1 g71103(.A (n_6289), .B (n_9301), .Y (n_8782));
NAND2X1 g71104(.A (n_8785), .B (n_8786), .Y (n_9656));
NAND2X1 g71105(.A (n_9301), .B (n_6528), .Y (n_8785));
NAND2X1 g71106(.A (n_6289), .B (n_6528), .Y (n_8786));
NAND2X1 g71108(.A (n_8791), .B (n_8793), .Y (n_8794));
OAI21X1 g71109(.A0 (n_8788), .A1 (n_8789), .B0 (n_8790), .Y (n_8791));
NAND2X1 g71110(.A (n_5930), .B (n_5918), .Y (n_8788));
NAND2X1 g71111(.A (n_6381), .B (g_8082), .Y (n_8789));
AOI21X1 g71112(.A0 (n_2014), .A1 (g1234), .B0 (n_6219), .Y (n_8790));
OR2X1 g71113(.A (g1230), .B (n_8792), .Y (n_8793));
INVX1 g71114(.A (n_6219), .Y (n_8792));
NAND3X1 g71115(.A (n_5930), .B (n_5918), .C (n_6381), .Y (n_8796));
INVX4 g71116(.A (g_8082), .Y (n_2014));
NAND2X1 g71124(.A (n_8806), .B (n_8809), .Y (n_8810));
OAI21X1 g71125(.A0 (n_935), .A1 (n_8805), .B0 (n_931), .Y (n_8806));
INVX1 g71126(.A (g231), .Y (n_8805));
AOI21X1 g71127(.A0 (n_2232), .A1 (n_8805), .B0 (n_9050), .Y (n_8809));
NAND2X1 g71143(.A (n_4760), .B (n_9432), .Y (n_8823));
NAND2X1 g71144(.A (n_4763), .B (n_4910), .Y (n_8824));
NAND2X2 g71145(.A (n_3847), .B (n_3681), .Y (n_8825));
INVX1 g71147(.A (n_8829), .Y (n_8830));
INVX1 g71148(.A (n_8825), .Y (n_8829));
NAND3X1 g46(.A (n_8833), .B (n_8834), .C (n_8836), .Y (n_8837));
AOI21X1 g71149(.A0 (n_8831), .A1 (n_5089), .B0 (n_8832), .Y (n_8833));
OR2X1 g71150(.A (n_4672), .B (n_8939), .Y (n_8831));
NAND4X1 g71151(.A (n_8758), .B (n_8761), .C (n_8762), .D (n_8764), .Y(n_8832));
AND2X1 g71152(.A (n_4636), .B (n_4637), .Y (n_8834));
OAI21X1 g48(.A0 (n_4645), .A1 (g2185), .B0 (n_8835), .Y (n_8836));
NAND2X1 g71153(.A (n_4645), .B (g2185), .Y (n_8835));
NAND2X1 g71154(.A (n_8841), .B (n_8842), .Y (n_8843));
NAND2X1 g71155(.A (n_8839), .B (n_9041), .Y (n_8841));
INVX1 g71156(.A (n_8838), .Y (n_8839));
OR2X1 g71157(.A (g869), .B (n_4061), .Y (n_8838));
NAND2X1 g71158(.A (n_9101), .B (n_8839), .Y (n_8842));
CLKBUFX1 g71159(.A (n_8843), .Y (n_8844));
AOI21X1 g71174(.A0 (n_8865), .A1 (n_9680), .B0 (n_8867), .Y (n_8868));
OR2X1 g71175(.A (n_8863), .B (n_9679), .Y (n_8865));
INVX1 g71176(.A (n_8862), .Y (n_8863));
INVX4 g71177(.A (n_8861), .Y (n_8862));
AND2X1 g71178(.A (n_9216), .B (n_5146), .Y (n_8861));
INVX1 g71180(.A (n_8866), .Y (n_8867));
INVX1 g71181(.A (n_8578), .Y (n_8866));
NAND2X1 g42_dup(.A (n_9679), .B (n_8873), .Y (n_8874));
INVX2 g71186(.A (n_8578), .Y (n_8873));
NOR2X1 g71188(.A (n_9679), .B (n_8578), .Y (n_8876));
OR2X1 g71189(.A (n_8885), .B (n_8886), .Y (n_8887));
NAND4X1 g71190(.A (n_4240), .B (n_8730), .C (n_8882), .D (n_8884), .Y(n_8885));
NOR2X1 g71191(.A (n_8879), .B (n_8881), .Y (n_8882));
CLKBUFX1 g73(.A (n_8878), .Y (n_8879));
INVX1 g74(.A (n_8877), .Y (n_8878));
AOI21X1 g75(.A0 (n_8408), .A1 (n_9650), .B0 (n_3103), .Y (n_8877));
INVX2 g71192(.A (n_8880), .Y (n_8881));
AOI21X1 g70(.A0 (n_8408), .A1 (n_9660), .B0 (n_3046), .Y (n_8880));
CLKBUFX1 g71193(.A (n_9044), .Y (n_8884));
NAND4X1 g63(.A (n_8411), .B (n_4016), .C (n_3812), .D (n_4339), .Y(n_8886));
INVX1 g71195(.A (n_9044), .Y (n_8888));
INVX1 g71(.A (n_8879), .Y (n_6653));
INVX1 g71196(.A (n_8881), .Y (n_4223));
NAND2X1 g6(.A (n_8891), .B (g2251), .Y (n_8892));
INVX1 g71197(.A (g_9470), .Y (n_8891));
INVX1 g7(.A (g_9470), .Y (n_9592));
AND2X1 g71201(.A (n_9370), .B (n_8644), .Y (n_8894));
NAND2X2 g71208(.A (n_3841), .B (n_3667), .Y (n_8901));
NAND2X1 g71211(.A (n_4910), .B (n_4763), .Y (n_8905));
INVX2 g71214(.A (n_8901), .Y (n_8909));
NAND3X1 g71217(.A (n_8911), .B (n_8912), .C (n_4644), .Y (n_8913));
NAND2X1 g71218(.A (n_5073), .B (n_5072), .Y (n_8911));
INVX1 g71219(.A (n_8424), .Y (n_8912));
NAND2X1 g71227(.A (n_8924), .B (n_9501), .Y (n_8929));
INVX1 g71228(.A (n_9556), .Y (n_8924));
NAND2X1 g71235(.A (n_8931), .B (n_8938), .Y (n_8939));
OR2X1 g71236(.A (g2237), .B (n_3770), .Y (n_8931));
AOI21X1 g71237(.A0 (n_8935), .A1 (n_8936), .B0 (n_8937), .Y (n_8938));
INVX2 g71238(.A (n_8934), .Y (n_8935));
INVX2 g71239(.A (n_8933), .Y (n_8934));
INVX2 g71240(.A (n_810), .Y (n_8933));
INVX1 g71242(.A (g2236), .Y (n_8936));
NOR2X1 g71243(.A (g2235), .B (n_3344), .Y (n_8937));
AOI22X1 g71245(.A0 (g1554), .A1 (n_8941), .B0 (n_8942), .B1 (g1555),.Y (n_8943));
CLKBUFX3 g71246(.A (n_8940), .Y (n_8941));
INVX1 g71247(.A (g_21829), .Y (n_8940));
OR2X1 g71248(.A (g1554), .B (n_757), .Y (n_8942));
CLKBUFX3 g71249(.A (n_8944), .Y (n_8945));
NAND2X1 g35_dup(.A (n_8940), .B (n_757), .Y (n_8944));
NOR2X1 g71250(.A (g1553), .B (n_3467), .Y (n_8946));
NAND2X1 g71251(.A (n_8940), .B (n_757), .Y (n_8948));
INVX2 g71252(.A (g_21829), .Y (n_8949));
NAND4X1 g71253(.A (n_8951), .B (n_8953), .C (n_8956), .D (n_8957), .Y(n_8958));
NOR2X1 g71254(.A (n_6159), .B (n_5687), .Y (n_8951));
AND2X1 g71256(.A (n_5987), .B (n_9677), .Y (n_8953));
NOR2X1 g71258(.A (n_8954), .B (n_9001), .Y (n_8956));
NAND2X2 g71260(.A (n_5299), .B (n_5112), .Y (n_8954));
NOR2X1 g71261(.A (n_5922), .B (n_6003), .Y (n_8957));
NOR2X1 g71263(.A (n_8960), .B (n_8967), .Y (n_8968));
OR2X1 g71264(.A (n_4670), .B (n_4671), .Y (n_8960));
NAND3X1 g36_dup(.A (n_8963), .B (n_9682), .C (n_8961), .Y (n_8967));
AND2X1 g71265(.A (n_8494), .B (n_8489), .Y (n_8961));
NOR2X1 g71266(.A (n_5132), .B (n_8962), .Y (n_8963));
INVX1 g71267(.A (n_8488), .Y (n_8962));
NAND2X1 g71269(.A (n_8964), .B (n_8495), .Y (n_8965));
INVX1 g71270(.A (n_8838), .Y (n_8964));
NAND3X1 g71280(.A (n_8979), .B (n_8980), .C (n_8984), .Y (n_8985));
NAND2X1 g71281(.A (n_5126), .B (n_4923), .Y (n_8979));
NAND2X1 g71282(.A (n_5011), .B (n_4917), .Y (n_8980));
INVX1 g26(.A (n_8983), .Y (n_8984));
MX2X1 g27_dup(.A (n_126), .B (g2165), .S0 (n_8982), .Y (n_8983));
NAND2X2 g71284(.A (n_3443), .B (n_2619), .Y (n_8982));
MX2X1 g71285(.A (n_126), .B (g2165), .S0 (n_8982), .Y (n_8986));
MX2X1 g71286(.A (n_8988), .B (n_8987), .S0 (n_9458), .Y (n_8990));
INVX1 g71287(.A (n_8987), .Y (n_8988));
OAI21X1 g71288(.A0 (n_2396), .A1 (n_3482), .B0 (n_3225), .Y (n_8987));
NAND2X2 g71293(.A (n_8993), .B (n_8994), .Y (n_8995));
NAND3X1 g71294(.A (n_2457), .B (n_918), .C (n_2921), .Y (n_8993));
OR2X1 g71295(.A (n_172), .B (n_4172), .Y (n_8994));
NAND2X1 g71296(.A (n_8999), .B (n_9000), .Y (n_9001));
MX2X1 g24_dup(.A (n_466), .B (g117), .S0 (n_8998), .Y (n_8999));
NAND2X2 g71298(.A (n_4147), .B (n_2922), .Y (n_8998));
MX2X1 g71299(.A (n_3187), .B (g109), .S0 (n_4836), .Y (n_9000));
MX2X1 g71300(.A (n_466), .B (g117), .S0 (n_8998), .Y (n_9002));
AOI21X1 g71301(.A0 (n_9003), .A1 (n_5970), .B0 (n_9005), .Y (n_9006));
OR2X1 g71302(.A (n_5656), .B (g125), .Y (n_9003));
XOR2X1 g71303(.A (g121), .B (n_5227), .Y (n_9005));
NAND3X1 g71308(.A (n_7545), .B (n_7605), .C (n_9139), .Y (n_9010));
NAND3X1 g59931_dup(.A (n_7545), .B (n_7605), .C (n_9140), .Y(n_9011));
INVX1 g71317(.A (n_9014), .Y (n_9021));
CLKBUFX1 g71319(.A (n_9024), .Y (n_9014));
INVX1 g71320(.A (n_9025), .Y (n_9024));
INVX1 g71321(.A (n_8563), .Y (n_9025));
NAND3X1 g71331(.A (n_9434), .B (n_9036), .C (n_9040), .Y (n_9041));
NAND3X1 g71333(.A (n_8823), .B (n_8824), .C (n_8825), .Y (n_9036));
NAND3X1 g71334(.A (n_9037), .B (n_9038), .C (n_9448), .Y (n_9040));
NAND2X1 g71335(.A (n_4486), .B (n_4498), .Y (n_9037));
NAND2X1 g71336(.A (n_9661), .B (n_9662), .Y (n_9038));
INVX1 g71340(.A (n_9042), .Y (n_9043));
AOI21X1 g71341(.A0 (n_8408), .A1 (n_2383), .B0 (n_3041), .Y (n_9042));
AOI21X1 g71342(.A0 (n_2399), .A1 (n_8408), .B0 (n_3057), .Y (n_9044));
NAND2X1 g24(.A (n_9052), .B (n_9053), .Y (n_9054));
NAND2X1 g71344(.A (n_9048), .B (n_9051), .Y (n_9052));
NAND2X1 g71345(.A (n_1133), .B (g_14013), .Y (n_9048));
AOI21X1 g71346(.A0 (n_2579), .A1 (g_25781), .B0 (n_9050), .Y(n_9051));
INVX1 g71347(.A (n_9049), .Y (n_9050));
NAND2X1 g71348(.A (n_2102), .B (n_9404), .Y (n_9049));
OR2X1 g71349(.A (g_25466), .B (n_9314), .Y (n_9053));
INVX1 g71350(.A (n_9050), .Y (n_9055));
NAND4X1 g71351(.A (n_9056), .B (n_9057), .C (n_9061), .D (n_9062), .Y(n_9063));
NAND3X1 g71352(.A (n_8784), .B (n_8280), .C (n_5150), .Y (n_9056));
NAND2X1 g71353(.A (n_6999), .B (n_7000), .Y (n_9057));
NAND2X1 g71354(.A (n_9059), .B (n_9060), .Y (n_9061));
INVX1 g71355(.A (n_9058), .Y (n_9059));
NAND2X2 g71356(.A (n_5758), .B (n_6396), .Y (n_9058));
NAND2X1 g71357(.A (n_2768), .B (n_3755), .Y (n_9060));
OR2X1 g71358(.A (n_5480), .B (n_5169), .Y (n_9062));
NAND3X1 g71359(.A (n_9571), .B (n_9572), .C (n_9070), .Y (n_9071));
NAND3X1 g71360(.A (n_5376), .B (n_5367), .C (n_4728), .Y (n_9572));
NAND3X1 g71361(.A (n_9065), .B (n_9066), .C (n_9067), .Y (n_9571));
NAND2X1 g71362(.A (n_8551), .B (n_5319), .Y (n_9065));
NAND2X1 g71363(.A (n_5368), .B (n_4769), .Y (n_9066));
NAND2X2 g71365(.A (n_4469), .B (n_4275), .Y (n_9067));
NAND3X1 g71366(.A (n_8550), .B (n_5369), .C (n_5178), .Y (n_9070));
INVX2 g71367(.A (n_9067), .Y (n_9072));
NOR2X1 g71368(.A (n_9076), .B (n_9080), .Y (n_9081));
INVX1 g71369(.A (n_9075), .Y (n_9076));
INVX2 g71370(.A (n_9074), .Y (n_9075));
AND2X1 g71371(.A (n_9073), .B (n_8541), .Y (n_9074));
NAND2X2 g71372(.A (n_7237), .B (n_8540), .Y (n_9073));
AOI22X1 g71373(.A0 (g2190), .A1 (n_7403), .B0 (n_9077), .B1 (n_9079),.Y (n_9080));
INVX4 g71375(.A (n_9073), .Y (n_9077));
OAI21X1 g71376(.A0 (n_8703), .A1 (n_4757), .B0 (n_7036), .Y (n_9079));
NAND3X1 g71378(.A (n_9087), .B (n_9088), .C (n_9089), .Y (n_9090));
NAND2X1 g71379(.A (n_9083), .B (n_9086), .Y (n_9087));
NAND2X1 g71380(.A (n_8771), .B (n_5320), .Y (n_9083));
AOI21X1 g71381(.A0 (n_5171), .A1 (n_9641), .B0 (n_9085), .Y (n_9086));
INVX2 g71382(.A (n_9084), .Y (n_9085));
NAND2X2 g71383(.A (n_4476), .B (n_4291), .Y (n_9084));
NAND3X1 g71384(.A (n_5358), .B (n_5359), .C (n_4918), .Y (n_9088));
NAND3X1 g71385(.A (n_5374), .B (n_8766), .C (n_5172), .Y (n_9089));
INVX1 g71386(.A (n_9085), .Y (n_9091));
NAND3X1 g71387(.A (n_9663), .B (n_9093), .C (n_9664), .Y (n_9101));
NAND3X1 g71388(.A (n_4777), .B (n_4527), .C (n_8901), .Y (n_9664));
NAND3X1 g71389(.A (n_4755), .B (n_8255), .C (n_4958), .Y (n_9093));
NAND3X1 g71390(.A (n_9683), .B (n_9684), .C (n_9236), .Y (n_9663));
NAND2X1 g71391(.A (n_4484), .B (n_4729), .Y (n_9684));
NAND2X1 g71392(.A (n_8909), .B (n_8609), .Y (n_9683));
NAND2X1 g71401(.A (n_5281), .B (n_5283), .Y (n_9104));
AND2X1 g71403(.A (n_5482), .B (n_5069), .Y (n_9106));
NAND2X1 g71404(.A (n_9110), .B (n_9113), .Y (n_9114));
INVX1 g71405(.A (n_9109), .Y (n_9110));
NAND3X1 g71406(.A (n_8653), .B (n_8894), .C (n_6726), .Y (n_9109));
NOR2X1 g71407(.A (n_9111), .B (n_9112), .Y (n_9113));
NAND3X1 g71408(.A (n_9629), .B (n_8961), .C (n_8963), .Y (n_9111));
NOR2X1 g71409(.A (n_4505), .B (n_8527), .Y (n_9112));
INVX1 g71412(.A (n_8954), .Y (n_9116));
INVX1 g71413(.A (n_9302), .Y (n_9119));
INVX2 g71420(.A (n_9303), .Y (n_9129));
INVX1 g71426(.A (n_9137), .Y (n_9136));
CLKBUFX1 g71427(.A (n_9302), .Y (n_9137));
INVX1 g71429(.A (n_9141), .Y (n_9140));
INVX2 g71430(.A (n_9139), .Y (n_9141));
INVX2 g71432(.A (n_9148), .Y (n_9144));
INVX2 g71434(.A (n_9148), .Y (n_9147));
INVX2 g71435(.A (n_7384), .Y (n_9148));
INVX1 g71471(.A (n_9188), .Y (n_9192));
CLKBUFX1 g71472(.A (n_4463), .Y (n_9188));
INVX1 g71473(.A (n_9195), .Y (n_9196));
INVX1 g71474(.A (n_9198), .Y (n_9195));
NAND2X1 g71477(.A (n_9296), .B (n_5184), .Y (n_9199));
NAND2X1 g71478(.A (n_5129), .B (n_4454), .Y (n_9200));
CLKBUFX1 g71479(.A (n_9529), .Y (n_9202));
NAND2X2 g71484(.A (n_9208), .B (n_9210), .Y (n_9211));
INVX4 g71485(.A (g_18412), .Y (n_9208));
CLKBUFX2 g71486(.A (n_9209), .Y (n_9210));
INVX1 g71487(.A (g_21387), .Y (n_9209));
NAND2X1 g71488(.A (n_9220), .B (n_9223), .Y (n_9224));
NAND3X1 g71489(.A (n_9214), .B (n_5717), .C (n_9219), .Y (n_9220));
NAND2X1 g71490(.A (n_9212), .B (n_8924), .Y (n_9214));
INVX1 g71491(.A (n_8958), .Y (n_9212));
INVX1 g71493(.A (n_9217), .Y (n_9219));
INVX1 g71495(.A (n_9216), .Y (n_9217));
INVX1 g71496(.A (n_9215), .Y (n_9216));
NAND2X1 g71497(.A (n_2776), .B (n_3939), .Y (n_9215));
NAND4X1 g71498(.A (n_9222), .B (n_8678), .C (n_8929), .D (n_9217), .Y(n_9223));
NAND2X1 g71499(.A (n_8924), .B (n_8958), .Y (n_9222));
NAND2X1 g71501(.A (n_9214), .B (n_5717), .Y (n_9225));
AND2X1 g71502(.A (n_8678), .B (n_8929), .Y (n_9226));
INVX1 g71503(.A (n_9222), .Y (n_9227));
NAND4X1 g71504(.A (n_9231), .B (n_9232), .C (n_9233), .D (n_9234), .Y(n_9235));
INVX1 g71505(.A (n_9230), .Y (n_9231));
NAND4X1 g71506(.A (n_4760), .B (n_8909), .C (n_9229), .D (n_4729), .Y(n_9230));
MX2X1 g71508(.A (n_504), .B (g785), .S0 (n_8410), .Y (n_9229));
NOR2X1 g71509(.A (n_8830), .B (n_4958), .Y (n_9232));
INVX1 g71510(.A (n_8905), .Y (n_9233));
NOR2X1 g71511(.A (n_8608), .B (n_9433), .Y (n_9234));
INVX1 g71512(.A (n_9229), .Y (n_9236));
MX2X1 g71516(.A (n_5380), .B (g101), .S0 (n_5030), .Y (n_9237));
NAND2X1 g71517(.A (n_5031), .B (n_5247), .Y (n_9238));
NAND2X1 g71518(.A (n_4800), .B (n_3187), .Y (n_9240));
NAND2X1 g78(.A (n_5032), .B (g113), .Y (n_9242));
OR2X1 g77(.A (n_3187), .B (n_4800), .Y (n_9243));
NAND3X1 g71521(.A (n_9254), .B (n_9255), .C (n_9256), .Y (n_9257));
NOR2X1 g71522(.A (n_9418), .B (n_9687), .Y (n_9254));
INVX1 g71523(.A (n_8471), .Y (n_9687));
AND2X1 g71527(.A (n_8770), .B (n_6529), .Y (n_9255));
NAND2X1 g71528(.A (n_2773), .B (n_4133), .Y (n_9256));
NAND2X1 g71538(.A (n_9272), .B (n_9657), .Y (n_9273));
AND2X1 g71539(.A (n_9267), .B (n_9268), .Y (n_9657));
NOR2X1 g71540(.A (n_5099), .B (n_9217), .Y (n_9267));
AND2X1 g71541(.A (n_7215), .B (n_5337), .Y (n_9268));
NOR2X1 g71542(.A (n_9270), .B (n_9271), .Y (n_9272));
NAND2X2 g71543(.A (n_9555), .B (n_9006), .Y (n_9270));
NOR2X1 g71544(.A (n_9556), .B (n_9503), .Y (n_9271));
XOR2X1 g71554(.A (g2185), .B (n_9284), .Y (n_9285));
INVX1 g21(.A (n_9283), .Y (n_9284));
AOI21X1 g22(.A0 (n_2314), .A1 (n_3799), .B0 (n_3343), .Y (n_9283));
NAND2X1 g71555(.A (n_9289), .B (n_5126), .Y (n_9292));
INVX2 g71556(.A (n_9288), .Y (n_9289));
NAND2X2 g71557(.A (n_9286), .B (n_9287), .Y (n_9288));
NAND2X2 g71558(.A (n_3988), .B (n_11), .Y (n_9286));
NAND2X1 g71559(.A (g2175), .B (n_3800), .Y (n_9287));
NAND2X1 g71561(.A (n_4475), .B (n_4292), .Y (n_9290));
NAND3X1 g71563(.A (n_9294), .B (n_9295), .C (n_9300), .Y (n_9301));
NAND3X1 g71564(.A (n_9199), .B (n_9200), .C (n_9202), .Y (n_9294));
NAND3X1 g71565(.A (n_4770), .B (n_5365), .C (n_5303), .Y (n_9295));
NAND3X1 g71566(.A (n_9297), .B (n_9298), .C (n_9537), .Y (n_9300));
INVX1 g71567(.A (n_9296), .Y (n_9297));
MX2X1 g71568(.A (n_385), .B (g2190), .S0 (n_3994), .Y (n_9296));
NAND2X1 g71569(.A (n_5129), .B (n_5184), .Y (n_9298));
NAND2X2 g71571(.A (n_9303), .B (n_9308), .Y (n_9309));
CLKBUFX3 g71572(.A (n_9302), .Y (n_9303));
NAND3X1 g71573(.A (n_8650), .B (n_8644), .C (n_9369), .Y (n_9302));
NOR2X1 g71574(.A (n_9307), .B (n_9304), .Y (n_9308));
NAND3X1 g71575(.A (n_9114), .B (n_8517), .C (n_9374), .Y (n_9304));
NAND2X1 g71576(.A (n_9305), .B (n_5325), .Y (n_9307));
NAND2X1 g71577(.A (n_8210), .B (n_8211), .Y (n_9305));
INVX1 g71580(.A (n_9307), .Y (n_9311));
OAI21X1 g71581(.A0 (n_9315), .A1 (n_9316), .B0 (n_9320), .Y (n_9321));
INVX1 g71582(.A (n_9314), .Y (n_9315));
INVX4 g71584(.A (n_9312), .Y (n_9314));
CLKBUFX3 g71585(.A (g_5550), .Y (n_9312));
INVX1 g71586(.A (g246), .Y (n_9316));
NAND3X1 g71587(.A (n_9315), .B (n_9318), .C (n_9566), .Y (n_9320));
CLKBUFX1 g71588(.A (n_9486), .Y (n_9318));
NAND2X2 g71591(.A (n_9318), .B (n_9566), .Y (n_9322));
INVX2 g71592(.A (g_5550), .Y (n_4172));
NAND2X2 g71607(.A (n_9343), .B (n_9345), .Y (n_9346));
AOI22X1 g71608(.A0 (n_4237), .A1 (n_9342), .B0 (n_9341), .B1(n_4236), .Y (n_9343));
INVX1 g71609(.A (n_9341), .Y (n_9342));
INVX1 g71610(.A (n_9340), .Y (n_9341));
AND2X1 g71611(.A (n_9025), .B (n_4934), .Y (n_9340));
NAND2X2 g29(.A (n_9344), .B (n_9341), .Y (n_9345));
NAND2X2 g71612(.A (n_5150), .B (n_5480), .Y (n_9344));
CLKBUFX1 g71613(.A (n_9344), .Y (n_9347));
NAND4X1 g71625(.A (n_9579), .B (n_9580), .C (n_9364), .D (n_9365), .Y(n_9366));
AOI21X1 g71626(.A0 (n_4410), .A1 (n_5482), .B0 (n_5568), .Y (n_9580));
AOI21X1 g71628(.A0 (n_8427), .A1 (n_4477), .B0 (n_9362), .Y (n_9579));
NAND2X1 g71629(.A (n_9361), .B (n_4849), .Y (n_9362));
NAND2X1 g71630(.A (n_8423), .B (n_8421), .Y (n_9361));
NOR2X1 g71631(.A (n_8913), .B (n_9106), .Y (n_9364));
NOR2X1 g71632(.A (n_9104), .B (n_5743), .Y (n_9365));
NAND2X2 g71633(.A (n_9367), .B (n_9377), .Y (n_9378));
NAND2X1 g71634(.A (n_7488), .B (n_9370), .Y (n_9367));
AOI21X1 g71635(.A0 (n_9368), .A1 (n_9373), .B0 (n_9376), .Y (n_9377));
NAND2X1 g71636(.A (n_8653), .B (n_7299), .Y (n_9368));
NOR2X1 g71637(.A (n_4192), .B (n_5290), .Y (n_9373));
INVX2 g71640(.A (n_9369), .Y (n_9370));
NAND2X2 g71641(.A (n_8647), .B (n_3331), .Y (n_9369));
INVX1 g71642(.A (n_9375), .Y (n_9376));
CLKBUFX1 g71643(.A (n_9374), .Y (n_9375));
NAND2X1 g71644(.A (n_6544), .B (n_6546), .Y (n_9374));
AOI21X1 g71645(.A0 (n_7299), .A1 (n_8653), .B0 (n_5290), .Y (n_9379));
NAND2X1 g71646(.A (n_9381), .B (g2273), .Y (n_9382));
INVX1 g71647(.A (n_9380), .Y (n_9381));
INVX2 g71648(.A (g_9470), .Y (n_9380));
INVX1 g71649(.A (g2273), .Y (n_9383));
INVX1 g71658(.A (n_9515), .Y (n_9392));
OAI21X1 g71659(.A0 (n_9395), .A1 (g_29207), .B0 (n_9402), .Y(n_9403));
INVX1 g71660(.A (n_9394), .Y (n_9395));
INVX2 g71661(.A (n_9393), .Y (n_9394));
INVX1 g71662(.A (g_4886), .Y (n_9393));
AOI21X1 g71663(.A0 (n_9399), .A1 (n_9400), .B0 (n_9401), .Y (n_9402));
INVX1 g71664(.A (n_9398), .Y (n_9399));
CLKBUFX3 g71665(.A (n_9397), .Y (n_9398));
INVX2 g71666(.A (n_9439), .Y (n_9397));
INVX1 g71668(.A (g_24922), .Y (n_9400));
NOR2X1 g71669(.A (g_14677), .B (n_9314), .Y (n_9401));
INVX1 g71670(.A (g_4886), .Y (n_9404));
NAND3X1 g71677(.A (n_9422), .B (n_9423), .C (n_9424), .Y (n_9425));
NAND3X1 g71678(.A (n_9419), .B (n_8471), .C (n_9421), .Y (n_9422));
INVX1 g71679(.A (n_9418), .Y (n_9419));
NAND2X2 g71680(.A (n_8655), .B (n_8656), .Y (n_9418));
INVX1 g71681(.A (n_9420), .Y (n_9421));
NAND3X1 g71682(.A (n_9256), .B (n_8710), .C (n_5477), .Y (n_9420));
NAND2X1 g71683(.A (n_6996), .B (n_9256), .Y (n_9423));
AOI21X1 g71684(.A0 (n_8471), .A1 (n_8472), .B0 (n_5357), .Y (n_9424));
AND2X1 g71685(.A (n_8471), .B (n_8472), .Y (n_9426));
NAND3X1 g71686(.A (n_9427), .B (n_9428), .C (n_9433), .Y (n_9434));
NAND2X1 g71687(.A (n_4910), .B (n_4760), .Y (n_9427));
NAND2X1 g71688(.A (n_8829), .B (n_4763), .Y (n_9428));
INVX1 g71689(.A (n_9432), .Y (n_9433));
INVX2 g71690(.A (n_9431), .Y (n_9432));
NAND2X2 g71691(.A (n_9429), .B (n_9430), .Y (n_9431));
NAND2X1 g71692(.A (n_9043), .B (n_9044), .Y (n_9429));
NAND2X1 g71693(.A (n_8888), .B (n_9042), .Y (n_9430));
NOR2X1 g71694(.A (n_9695), .B (n_9694), .Y (n_9437));
NOR2X1 g71695(.A (g2392), .B (n_4576), .Y (n_9694));
OAI22X1 g71696(.A0 (n_9510), .A1 (g2390), .B0 (g2391), .B1 (n_2078),.Y (n_9695));
AND2X1 g71697(.A (n_9510), .B (n_2078), .Y (n_9438));
AOI21X1 g71698(.A0 (n_9441), .A1 (n_9442), .B0 (n_9443), .Y (n_9444));
AOI22X1 g71699(.A0 (g_24786), .A1 (n_9440), .B0 (n_9404), .B1(n_2102), .Y (n_9441));
INVX1 g71700(.A (n_9439), .Y (n_9440));
BUFX1 g71701(.A (g_20948), .Y (n_9439));
OAI21X1 g71702(.A0 (n_748), .A1 (g_24786), .B0 (g_30213), .Y(n_9442));
NOR2X1 g71703(.A (g_5159), .B (n_4172), .Y (n_9443));
MX2X1 g71705(.A (n_496), .B (g805), .S0 (n_9447), .Y (n_9448));
AOI21X1 g71707(.A0 (n_2388), .A1 (n_8408), .B0 (n_3052), .Y (n_9447));
INVX1 g71708(.A (n_9447), .Y (n_9449));
OAI21X1 g71714(.A0 (n_5469), .A1 (n_9490), .B0 (n_9243), .Y (n_9453));
NAND4X1 g71717(.A (n_9460), .B (n_4853), .C (n_4863), .D (n_9461), .Y(n_9462));
XOR2X1 g71718(.A (n_4780), .B (n_4450), .Y (n_9460));
CLKBUFX1 g71719(.A (n_9458), .Y (n_4780));
AOI21X1 g71720(.A0 (n_2136), .A1 (n_3799), .B0 (n_3333), .Y (n_9458));
XOR2X1 g71721(.A (g2190), .B (n_4211), .Y (n_9461));
INVX1 g71722(.A (n_4780), .Y (n_9463));
OR2X1 g71736(.A (n_8), .B (n_1946), .Y (n_9475));
OR2X1 g71737(.A (n_93), .B (n_8643), .Y (n_9476));
OR2X1 g71738(.A (n_3224), .B (n_64), .Y (n_9477));
NAND3X1 g71739(.A (n_9485), .B (n_9486), .C (n_9487), .Y (n_9488));
NAND3X1 g71740(.A (n_9557), .B (n_9484), .C (g105), .Y (n_9485));
INVX1 g71742(.A (n_9483), .Y (n_9484));
CLKBUFX3 g71743(.A (n_9561), .Y (n_9483));
NAND2X2 g71746(.A (n_9198), .B (n_9557), .Y (n_9486));
NAND2X1 g71747(.A (n_7726), .B (n_6905), .Y (n_9487));
INVX1 g71748(.A (n_9483), .Y (n_9489));
INVX1 g71749(.A (g105), .Y (n_9490));
NOR2X1 g71755(.A (n_9501), .B (n_9502), .Y (n_9503));
NAND3X1 g71756(.A (n_9498), .B (n_9499), .C (n_9500), .Y (n_9501));
NAND3X1 g71757(.A (n_6049), .B (n_9001), .C (n_5922), .Y (n_9498));
NAND3X1 g71758(.A (n_6050), .B (n_5734), .C (n_5498), .Y (n_9499));
NAND3X1 g71759(.A (n_5735), .B (n_5574), .C (n_8954), .Y (n_9500));
NAND3X1 g71760(.A (n_6481), .B (n_6480), .C (n_6363), .Y (n_9502));
NAND2X2 g71761(.A (n_9507), .B (n_9508), .Y (n_9509));
NAND2X1 g71762(.A (n_9581), .B (n_9582), .Y (n_9507));
NAND2X1 g71763(.A (n_2071), .B (n_139), .Y (n_9582));
AOI21X1 g71764(.A0 (n_848), .A1 (n_9393), .B0 (n_9505), .Y (n_9581));
AND2X1 g71765(.A (n_9404), .B (n_2102), .Y (n_9505));
OR2X1 g27(.A (n_226), .B (n_4172), .Y (n_9508));
OAI21X1 g18(.A0 (g5555), .A1 (n_9514), .B0 (n_9517), .Y (n_9518));
BUFX3 g71767(.A (n_9510), .Y (n_9512));
INVX2 g71768(.A (g_17130), .Y (n_9510));
INVX1 g71769(.A (g2390), .Y (n_9514));
INVX1 g19(.A (n_9516), .Y (n_9517));
NOR2X1 g71770(.A (n_9515), .B (n_9512), .Y (n_9516));
NAND3X1 g71771(.A (n_7723), .B (n_7660), .C (n_8542), .Y (n_9515));
NAND2X1 g71782(.A (n_9696), .B (n_9697), .Y (n_9537));
INVX2 g71783(.A (n_9529), .Y (n_9696));
NAND2X2 g71784(.A (n_4468), .B (n_4274), .Y (n_9529));
INVX1 g71785(.A (n_9535), .Y (n_9697));
OAI21X1 g71786(.A0 (n_9531), .A1 (n_2706), .B0 (n_9534), .Y (n_9535));
NAND3X1 g71787(.A (n_9475), .B (n_9476), .C (n_9477), .Y (n_9531));
NAND2X1 g71789(.A (n_9533), .B (n_2706), .Y (n_9534));
NAND3X1 g29_dup(.A (n_9475), .B (n_9476), .C (n_9477), .Y (n_9533));
INVX1 g71790(.A (n_9535), .Y (n_9538));
NOR2X1 g76(.A (n_9545), .B (n_9554), .Y (n_9555));
NAND4X1 g71791(.A (n_9540), .B (n_9542), .C (n_9543), .D (n_9544), .Y(n_9545));
INVX1 g81(.A (n_9539), .Y (n_9540));
NAND4X1 g82(.A (n_9237), .B (n_9242), .C (n_9238), .D (n_9240), .Y(n_9539));
AOI22X1 g80(.A0 (n_9541), .A1 (n_8743), .B0 (n_5469), .B1 (n_9490),.Y (n_9542));
INVX1 g91(.A (n_8741), .Y (n_9541));
NAND2X1 g88(.A (n_5658), .B (n_5654), .Y (n_9543));
MX2X1 g83(.A (n_466), .B (g117), .S0 (n_5029), .Y (n_9544));
NAND4X1 g71792(.A (n_9589), .B (n_9549), .C (n_9548), .D (n_9553), .Y(n_9554));
NOR2X1 g86(.A (n_9546), .B (n_9547), .Y (n_9548));
INVX1 g89(.A (g_22408), .Y (n_9546));
INVX1 g92(.A (n_9054), .Y (n_9547));
NAND2X1 g87(.A (n_5973), .B (n_9403), .Y (n_9549));
AOI21X1 g71793(.A0 (n_9550), .A1 (n_8741), .B0 (n_9453), .Y (n_9589));
INVX1 g93(.A (n_8743), .Y (n_9550));
NAND2X1 g84(.A (n_5973), .B (n_5974), .Y (n_9553));
INVX1 g85(.A (n_9548), .Y (n_9556));
OAI21X1 g71794(.A0 (n_9559), .A1 (n_7726), .B0 (n_9565), .Y (n_9566));
AND2X1 g71795(.A (n_9557), .B (n_3187), .Y (n_9559));
NAND3X1 g71796(.A (n_8866), .B (n_9680), .C (n_8862), .Y (n_9557));
INVX1 g71797(.A (g109), .Y (n_3187));
INVX2 g71799(.A (n_9561), .Y (n_9562));
INVX2 g71800(.A (n_9560), .Y (n_9561));
NAND2X2 g71801(.A (n_8873), .B (n_9679), .Y (n_9560));
INVX1 g71802(.A (n_9564), .Y (n_9565));
AOI21X1 g71803(.A0 (n_6921), .A1 (n_6816), .B0 (n_9562), .Y (n_9564));
NOR2X1 g71804(.A (n_4722), .B (n_8965), .Y (n_9682));
NOR2X1 g71268_dup(.A (n_4722), .B (n_8965), .Y (n_9629));
NAND4X1 g71805(.A (n_3133), .B (n_2991), .C (n_2992), .D (n_3134), .Y(n_9630));
NAND4X1 g62259_dup(.A (n_3133), .B (n_2991), .C (n_2992), .D(n_3134), .Y (n_9631));
INVX1 g71806(.A (n_9640), .Y (n_9632));
INVX1 g71807(.A (n_9637), .Y (n_9633));
CLKBUFX1 g71813(.A (n_9640), .Y (n_9637));
INVX2 g71815(.A (n_8557), .Y (n_9641));
CLKBUFX1 g71817(.A (n_9656), .Y (n_9654));
INVX1 g71818(.A (n_9656), .Y (n_9655));
AOI21X1 g71819(.A0 (n_2386), .A1 (n_8408), .B0 (n_3055), .Y (n_9671));
AOI21X1 g65158_dup(.A0 (n_2386), .A1 (n_8408), .B0 (n_3055), .Y(n_9672));
NOR2X1 g71820(.A (n_6530), .B (n_7025), .Y (n_9673));
NOR2X1 g61051_dup(.A (n_6530), .B (n_7025), .Y (n_9674));
AOI21X1 g71821(.A0 (n_8943), .A1 (n_8945), .B0 (n_8946), .Y (n_9675));
AOI21X1 g71244_dup(.A0 (n_8943), .A1 (n_8945), .B0 (n_8946), .Y(n_9676));
MX2X1 g71822(.A (g105), .B (n_9490), .S0 (n_8995), .Y (n_9677));
MX2X1 g71291_dup(.A (g105), .B (n_9490), .S0 (n_8995), .Y (n_9678));
INVX1 g71823(.A (n_9679), .Y (n_9680));
CLKBUFX3 g71824(.A (n_8576), .Y (n_9679));
endmodule
