module gcm_aes_v0(clk, rst, dii_data, dii_data_vld, dii_data_type, dii_data_not_ready, dii_last_word, dii_data_size, cii_ctl_vld, cii_IV_vld, cii_K, Out_data, Out_vld, Out_data_size, Out_last_word, Tag_vld, ddout__1, qq_in1, qnn_in_1, ddout__2, qq_in2, qnn_in_2, ddout__3, qq_in3, qnn_in_3, ddout__4, qq_in4, qnn_in_4, ddout__5, qq_in5, qnn_in_5, ddout__6, qq_in6, qnn_in_6, ddout__7, qq_in7, qnn_in_7, ddout__8, qq_in8, qnn_in_8, ddout__9, qq_in9, qnn_in_9, ddout__10, qq_in10, qnn_in_10, ddout__11, qq_in11, qnn_in_11, ddout__12, qq_in12, qnn_in_12, ddout__13, qq_in13, qnn_in_13, ddout__14, qq_in14, qnn_in_14, ddout__15, qq_in15, qnn_in_15, ddout__16, qq_in16, qnn_in_16, ddout__17, qq_in17, qnn_in_17, ddout__18, qq_in18, qnn_in_18, ddout__19, qq_in19, qnn_in_19, ddout__20, qq_in20, qnn_in_20, ddout__21, qq_in21, qnn_in_21, ddout__22, qq_in22, qnn_in_22, ddout__23, qq_in23, qnn_in_23, ddout__24, qq_in24, qnn_in_24, ddout__25, qq_in25, qnn_in_25, ddout__26, qq_in26, qnn_in_26, ddout__27, qq_in27, qnn_in_27, ddout__28, qq_in28, qnn_in_28, ddout__29, qq_in29, qnn_in_29, ddout__30, qq_in30, qnn_in_30, ddout__31, qq_in31, qnn_in_31, ddout__32, qq_in32, qnn_in_32, ddout__33, qq_in33, qnn_in_33, ddout__34, qq_in34, qnn_in_34, ddout__35, qq_in35, qnn_in_35, ddout__36, qq_in36, qnn_in_36, ddout__37, qq_in37, qnn_in_37, ddout__38, qq_in38, qnn_in_38, ddout__39, qq_in39, qnn_in_39, ddout__40, qq_in40, qnn_in_40, ddout__41, qq_in41, qnn_in_41, ddout__42, qq_in42, qnn_in_42, ddout__43, qq_in43, qnn_in_43, ddout__44, qq_in44, qnn_in_44, ddout__45, qq_in45, qnn_in_45, ddout__46, qq_in46, qnn_in_46, ddout__47, qq_in47, qnn_in_47, ddout__48, qq_in48, qnn_in_48, ddout__49, qq_in49, qnn_in_49, ddout__50, qq_in50, qnn_in_50, ddout__51, qq_in51, qnn_in_51, ddout__52, qq_in52, qnn_in_52, ddout__53, qq_in53, qnn_in_53, ddout__54, qq_in54, qnn_in_54, ddout__55, qq_in55, qnn_in_55, ddout__56, qq_in56, qnn_in_56, ddout__57, qq_in57, qnn_in_57, ddout__58, qq_in58, qnn_in_58, ddout__59, qq_in59, qnn_in_59, ddout__60, qq_in60, qnn_in_60, ddout__61, qq_in61, qnn_in_61, ddout__62, qq_in62, qnn_in_62, ddout__63, qq_in63, qnn_in_63, ddout__64, qq_in64, qnn_in_64, ddout__65, qq_in65, qnn_in_65, ddout__66, qq_in66, qnn_in_66, ddout__67, qq_in67, qnn_in_67, ddout__68, qq_in68, qnn_in_68, ddout__69, qq_in69, qnn_in_69, ddout__70, qq_in70, qnn_in_70, ddout__71, qq_in71, qnn_in_71, ddout__72, qq_in72, qnn_in_72, ddout__73, qq_in73, qnn_in_73, ddout__74, qq_in74, qnn_in_74, ddout__75, qq_in75, qnn_in_75, ddout__76, qq_in76, qnn_in_76, ddout__77, qq_in77, qnn_in_77, ddout__78, qq_in78, qnn_in_78, ddout__79, qq_in79, qnn_in_79, ddout__80, qq_in80, qnn_in_80, ddout__81, qq_in81, qnn_in_81, ddout__82, qq_in82, qnn_in_82, ddout__83, qq_in83, qnn_in_83, ddout__84, qq_in84, qnn_in_84, ddout__85, qq_in85, qnn_in_85, ddout__86, qq_in86, qnn_in_86, ddout__87, qq_in87, qnn_in_87, ddout__88, qq_in88, qnn_in_88, ddout__89, qq_in89, qnn_in_89, ddout__90, qq_in90, qnn_in_90, ddout__91, qq_in91, qnn_in_91, ddout__92, qq_in92, qnn_in_92, ddout__93, qq_in93, qnn_in_93, ddout__94, qq_in94, qnn_in_94, ddout__95, qq_in95, qnn_in_95, ddout__96, qq_in96, qnn_in_96, ddout__97, qq_in97, qnn_in_97, ddout__98, qq_in98, qnn_in_98, ddout__99, qq_in99, qnn_in_99, ddout__100, qq_in100, qnn_in_100, ddout__101, qq_in101, qnn_in_101, ddout__102, qq_in102, qnn_in_102, ddout__103, qq_in103, qnn_in_103, ddout__104, qq_in104, qnn_in_104, ddout__105, qq_in105, qnn_in_105, ddout__106, qq_in106, qnn_in_106, ddout__107, qq_in107, qnn_in_107, ddout__108, qq_in108, qnn_in_108, ddout__109, qq_in109, qnn_in_109, ddout__110, qq_in110, qnn_in_110, ddout__111, qq_in111, qnn_in_111, ddout__112, qq_in112, qnn_in_112, ddout__113, qq_in113, qnn_in_113, ddout__114, qq_in114, qnn_in_114, ddout__115, qq_in115, qnn_in_115, ddout__116, qq_in116, qnn_in_116, ddout__117, qq_in117, qnn_in_117, ddout__118, qq_in118, qnn_in_118, ddout__119, qq_in119, qnn_in_119, ddout__120, qq_in120, qnn_in_120, ddout__121, qq_in121, qnn_in_121, ddout__122, qq_in122, qnn_in_122, ddout__123, qq_in123, qnn_in_123, ddout__124, qq_in124, qnn_in_124, ddout__125, qq_in125, qnn_in_125, ddout__126, qq_in126, qnn_in_126, ddout__127, qq_in127, qnn_in_127, ddout__128, qq_in128, qnn_in_128, ddout__129, qq_in129, ddout__130, qq_in130, ddout__131, qq_in131, ddout__132, qq_in132, ddout__133, qq_in133, ddout__134, qq_in134, ddout__135, qq_in135, ddout__136, qq_in136, ddout__137, qq_in137, ddout__138, qq_in138, ddout__139, qq_in139, ddout__140, qq_in140, ddout__141, qq_in141, ddout__142, qq_in142, ddout__143, qq_in143, ddout__144, qq_in144, ddout__145, qq_in145, ddout__146, qq_in146, ddout__147, qq_in147, ddout__148, qq_in148, ddout__149, qq_in149, ddout__150, qq_in150, ddout__151, qq_in151, ddout__152, qq_in152, ddout__153, qq_in153, ddout__154, qq_in154, ddout__155, qq_in155, ddout__156, qq_in156, ddout__157, qq_in157, ddout__158, qq_in158, ddout__159, qq_in159, ddout__160, qq_in160, ddout__161, qq_in161, ddout__162, qq_in162, ddout__163, qq_in163, ddout__164, qq_in164, ddout__165, qq_in165, ddout__166, qq_in166, ddout__167, qq_in167, ddout__168, qq_in168, ddout__169, qq_in169, ddout__170, qq_in170, ddout__171, qq_in171, ddout__172, qq_in172, ddout__173, qq_in173, ddout__174, qq_in174, ddout__175, qq_in175, ddout__176, qq_in176, ddout__177, qq_in177, ddout__178, qq_in178, ddout__179, qq_in179, ddout__180, qq_in180, ddout__181, qq_in181, ddout__182, qq_in182, ddout__183, qq_in183, ddout__184, qq_in184, ddout__185, qq_in185, ddout__186, qq_in186, ddout__187, qq_in187, ddout__188, qq_in188, ddout__189, qq_in189, ddout__190, qq_in190, ddout__191, qq_in191, ddout__192, qq_in192, ddout__193, qq_in193, ddout__194, qq_in194, ddout__195, qq_in195, ddout__196, qq_in196, ddout__197, qq_in197, ddout__198, qq_in198, ddout__199, qq_in199, ddout__200, qq_in200, ddout__201, qq_in201, ddout__202, qq_in202, ddout__203, qq_in203, ddout__204, qq_in204, ddout__205, qq_in205, ddout__206, qq_in206, ddout__207, qq_in207, ddout__208, qq_in208, ddout__209, qq_in209, ddout__210, qq_in210, ddout__211, qq_in211, ddout__212, qq_in212, ddout__213, qq_in213, ddout__214, qq_in214, ddout__215, qq_in215, ddout__216, qq_in216, ddout__217, qq_in217, ddout__218, qq_in218, ddout__219, qq_in219, ddout__220, qq_in220, ddout__221, qq_in221, ddout__222, qq_in222, ddout__223, qq_in223, ddout__224, qq_in224, ddout__225, qq_in225, ddout__226, qq_in226, ddout__227, qq_in227, ddout__228, qq_in228, ddout__229, qq_in229, ddout__230, qq_in230, ddout__231, qq_in231, ddout__232, qq_in232, ddout__233, qq_in233, ddout__234, qq_in234, ddout__235, qq_in235, ddout__236, qq_in236, ddout__237, qq_in237, ddout__238, qq_in238, ddout__239, qq_in239, ddout__240, qq_in240, ddout__241, qq_in241, ddout__242, qq_in242, ddout__243, qq_in243, ddout__244, qq_in244, ddout__245, qq_in245, ddout__246, qq_in246, ddout__247, qq_in247, ddout__248, qq_in248, ddout__249, qq_in249, ddout__250, qq_in250, ddout__251, qq_in251, ddout__252, qq_in252, ddout__253, qq_in253, ddout__254, qq_in254, ddout__255, qq_in255, ddout__256, qq_in256, ddout__257, qq_in257, ddout__258, qq_in258, ddout__259, qq_in259, ddout__260, qq_in260, ddout__261, qq_in261, ddout__262, qq_in262, ddout__263, qq_in263, ddout__264, qq_in264, ddout__265, qq_in265, ddout__266, qq_in266, ddout__267, qq_in267, ddout__268, qq_in268, ddout__269, qq_in269, ddout__270, qq_in270, ddout__271, qq_in271, ddout__272, qq_in272, ddout__273, qq_in273, ddout__274, qq_in274, ddout__275, qq_in275, ddout__276, qq_in276, ddout__277, qq_in277, ddout__278, qq_in278, ddout__279, qq_in279, ddout__280, qq_in280, ddout__281, qq_in281, ddout__282, qq_in282, ddout__283, qq_in283, ddout__284, qq_in284, ddout__285, qq_in285, ddout__286, qq_in286, ddout__287, qq_in287, ddout__288, qq_in288, ddout__289, qq_in289, ddout__290, qq_in290, ddout__291, qq_in291, ddout__292, qq_in292, ddout__293, qq_in293, ddout__294, qq_in294, ddout__295, qq_in295, ddout__296, qq_in296, ddout__297, qq_in297, ddout__298, qq_in298, ddout__299, qq_in299, ddout__300, qq_in300, ddout__301, qq_in301, ddout__302, qq_in302, ddout__303, qq_in303, ddout__304, qq_in304, ddout__305, qq_in305, ddout__306, qq_in306, ddout__307, qq_in307, ddout__308, qq_in308, ddout__309, qq_in309, ddout__310, qq_in310, ddout__311, qq_in311, ddout__312, qq_in312, ddout__313, qq_in313, ddout__314, qq_in314, ddout__315, qq_in315, ddout__316, qq_in316, ddout__317, qq_in317, ddout__318, qq_in318, ddout__319, qq_in319, ddout__320, qq_in320, ddout__321, qq_in321, ddout__322, qq_in322, ddout__323, qq_in323, ddout__324, qq_in324, ddout__325, qq_in325, ddout__326, qq_in326, ddout__327, qq_in327, ddout__328, qq_in328, ddout__329, qq_in329, ddout__330, qq_in330, ddout__331, qq_in331, ddout__332, qq_in332, ddout__333, qq_in333, ddout__334, qq_in334, ddout__335, qq_in335, ddout__336, qq_in336, ddout__337, qq_in337, ddout__338, qq_in338, ddout__339, qq_in339, ddout__340, qq_in340, ddout__341, qq_in341, ddout__342, qq_in342, ddout__343, qq_in343, ddout__344, qq_in344, ddout__345, qq_in345, ddout__346, qq_in346, ddout__347, qq_in347, ddout__348, qq_in348, ddout__349, qq_in349, ddout__350, qq_in350, ddout__351, qq_in351, ddout__352, qq_in352, ddout__353, qq_in353, ddout__354, qq_in354, ddout__355, qq_in355, ddout__356, qq_in356, ddout__357, qq_in357, ddout__358, qq_in358, ddout__359, qq_in359, ddout__360, qq_in360, ddout__361, qq_in361, ddout__362, qq_in362, ddout__363, qq_in363, ddout__364, qq_in364, ddout__365, qq_in365, ddout__366, qq_in366, ddout__367, qq_in367, ddout__368, qq_in368, ddout__369, qq_in369, ddout__370, qq_in370, ddout__371, qq_in371, ddout__372, qq_in372, ddout__373, qq_in373, ddout__374, qq_in374, ddout__375, qq_in375, ddout__376, qq_in376, ddout__377, qq_in377, ddout__378, qq_in378, ddout__379, qq_in379, ddout__380, qq_in380, ddout__381, qq_in381, ddout__382, qq_in382, ddout__383, qq_in383, ddout__384, qq_in384, ddout__385, qq_in385, ddout__386, qq_in386, ddout__387, qq_in387, ddout__388, qq_in388, ddout__389, qq_in389, ddout__390, qq_in390, ddout__391, qq_in391, ddout__392, qq_in392, ddout__393, qq_in393, ddout__394, qq_in394, ddout__395, qq_in395, ddout__396, qq_in396, ddout__397, qq_in397, ddout__398, qq_in398, ddout__399, qq_in399, ddout__400, qq_in400, ddout__401, qq_in401, ddout__402, qq_in402, ddout__403, qq_in403, ddout__404, qq_in404, ddout__405, qq_in405, ddout__406, qq_in406, ddout__407, qq_in407, ddout__408, qq_in408, ddout__409, qq_in409, ddout__410, qq_in410, ddout__411, qq_in411, ddout__412, qq_in412, ddout__413, qq_in413, ddout__414, qq_in414, ddout__415, qq_in415, ddout__416, qq_in416, ddout__417, qq_in417, ddout__418, qq_in418, ddout__419, qq_in419, ddout__420, qq_in420, ddout__421, qq_in421, ddout__422, qq_in422, ddout__423, qq_in423, ddout__424, qq_in424, ddout__425, qq_in425, ddout__426, qq_in426, ddout__427, qq_in427, ddout__428, qq_in428, ddout__429, qq_in429, ddout__430, qq_in430, ddout__431, qq_in431, ddout__432, qq_in432, ddout__433, qq_in433, ddout__434, qq_in434, ddout__435, qq_in435, ddout__436, qq_in436, ddout__437, qq_in437, ddout__438, qq_in438, ddout__439, qq_in439, ddout__440, qq_in440, ddout__441, qq_in441, ddout__442, qq_in442, ddout__443, qq_in443, ddout__444, qq_in444, ddout__445, qq_in445, ddout__446, qq_in446, ddout__447, qq_in447, ddout__448, qq_in448, ddout__449, qq_in449, ddout__450, qq_in450, ddout__451, qq_in451, ddout__452, qq_in452, ddout__453, qq_in453, ddout__454, qq_in454, ddout__455, qq_in455, ddout__456, qq_in456, ddout__457, qq_in457, ddout__458, qq_in458, ddout__459, qq_in459, ddout__460, qq_in460, ddout__461, qq_in461, ddout__462, qq_in462, ddout__463, qq_in463, ddout__464, qq_in464, ddout__465, qq_in465, ddout__466, qq_in466, ddout__467, qq_in467, ddout__468, qq_in468, ddout__469, qq_in469, ddout__470, qq_in470, ddout__471, qq_in471, ddout__472, qq_in472, ddout__473, qq_in473, ddout__474, qq_in474, ddout__475, qq_in475, ddout__476, qq_in476, ddout__477, qq_in477, ddout__478, qq_in478, ddout__479, qq_in479, ddout__480, qq_in480, ddout__481, qq_in481, ddout__482, qq_in482, ddout__483, qq_in483, ddout__484, qq_in484, ddout__485, qq_in485, ddout__486, qq_in486, ddout__487, qq_in487, ddout__488, qq_in488, ddout__489, qq_in489, ddout__490, qq_in490, ddout__491, qq_in491, ddout__492, qq_in492, ddout__493, qq_in493, ddout__494, qq_in494, ddout__495, qq_in495, ddout__496, qq_in496, ddout__497, qq_in497, ddout__498, qq_in498, ddout__499, qq_in499, ddout__500, qq_in500, ddout__501, qq_in501, ddout__502, qq_in502, ddout__503, qq_in503, ddout__504, qq_in504, ddout__505, qq_in505, ddout__506, qq_in506, ddout__507, qq_in507, ddout__508, qq_in508, ddout__509, qq_in509, ddout__510, qq_in510, ddout__511, qq_in511, ddout__512, qq_in512, ddout__513, qq_in513, ddout__514, qq_in514, ddout__515, qq_in515, ddout__516, qq_in516, ddout__517, qq_in517, ddout__518, qq_in518, ddout__519, qq_in519, ddout__520, qq_in520, ddout__521, qq_in521, ddout__522, qq_in522, ddout__523, qq_in523, ddout__524, qq_in524, ddout__525, qq_in525, ddout__526, qq_in526, ddout__527, qq_in527, ddout__528, qq_in528, ddout__529, qq_in529, ddout__530, qq_in530, ddout__531, qq_in531, ddout__532, qq_in532, ddout__533, qq_in533, ddout__534, qq_in534, ddout__535, qq_in535, ddout__536, qq_in536, ddout__537, qq_in537, ddout__538, qq_in538, ddout__539, qq_in539, ddout__540, qq_in540, ddout__541, qq_in541, ddout__542, qq_in542, ddout__543, qq_in543, ddout__544, qq_in544, ddout__545, qq_in545, ddout__546, qq_in546, ddout__547, qq_in547, ddout__548, qq_in548, ddout__549, qq_in549, ddout__550, qq_in550, ddout__551, qq_in551, ddout__552, qq_in552, ddout__553, qq_in553, ddout__554, qq_in554, ddout__555, qq_in555, ddout__556, qq_in556, ddout__557, qq_in557, ddout__558, qq_in558, ddout__559, qq_in559, ddout__560, qq_in560, ddout__561, qq_in561, ddout__562, qq_in562, ddout__563, qq_in563, ddout__564, qq_in564, ddout__565, qq_in565, ddout__566, qq_in566, ddout__567, qq_in567, ddout__568, qq_in568, ddout__569, qq_in569, ddout__570, qq_in570, ddout__571, qq_in571, ddout__572, qq_in572, ddout__573, qq_in573, ddout__574, qq_in574, ddout__575, qq_in575, ddout__576, qq_in576, ddout__577, qq_in577, ddout__578, qq_in578, ddout__579, qq_in579, ddout__580, qq_in580, ddout__581, qq_in581, ddout__582, qq_in582, ddout__583, qq_in583, ddout__584, qq_in584, ddout__585, qq_in585, ddout__586, qq_in586, ddout__587, qq_in587, ddout__588, qq_in588, ddout__589, qq_in589, ddout__590, qq_in590, ddout__591, qq_in591, ddout__592, qq_in592, ddout__593, qq_in593, ddout__594, qq_in594, ddout__595, qq_in595, ddout__596, qq_in596, ddout__597, qq_in597, ddout__598, qq_in598, ddout__599, qq_in599, ddout__600, qq_in600, ddout__601, qq_in601, ddout__602, qq_in602, ddout__603, qq_in603, ddout__604, qq_in604, ddout__605, qq_in605, ddout__606, qq_in606, ddout__607, qq_in607, ddout__608, qq_in608, ddout__609, qq_in609, ddout__610, qq_in610, ddout__611, qq_in611, ddout__612, qq_in612, ddout__613, qq_in613, ddout__614, qq_in614, ddout__615, qq_in615, ddout__616, qq_in616, ddout__617, qq_in617, ddout__618, qq_in618, ddout__619, qq_in619, ddout__620, qq_in620, ddout__621, qq_in621, ddout__622, qq_in622, ddout__623, qq_in623, ddout__624, qq_in624, ddout__625, qq_in625, ddout__626, qq_in626, ddout__627, qq_in627, ddout__628, qq_in628, ddout__629, qq_in629, ddout__630, qq_in630, ddout__631, qq_in631, ddout__632, qq_in632, ddout__633, qq_in633, ddout__634, qq_in634, ddout__635, qq_in635, ddout__636, qq_in636, ddout__637, qq_in637, ddout__638, qq_in638, ddout__639, qq_in639, ddout__640, qq_in640, ddout__641, qq_in641, ddout__642, qq_in642, ddout__643, qq_in643, ddout__644, qq_in644, ddout__645, qq_in645, ddout__646, qq_in646, ddout__647, qq_in647, ddout__648, qq_in648, ddout__649, qq_in649, qnn_in_649, ddout__650, qq_in650, qnn_in_650, ddout__651, qq_in651, qnn_in_651, ddout__652, qq_in652, ddout__653, qq_in653, ddout__654, qq_in654, qnn_in_654, ddout__655, qq_in655, ddout__656, qq_in656, ddout__657, qq_in657, ddout__658, qq_in658, ddout__659, qq_in659, ddout__660, qq_in660, ddout__661, qq_in661, ddout__662, qq_in662, ddout__663, qq_in663, ddout__664, qq_in664, ddout__665, qq_in665, ddout__666, qq_in666, ddout__667, qq_in667, qnn_in_667, ddout__668, qq_in668, qnn_in_668, ddout__669, qq_in669, qnn_in_669, ddout__670, qq_in670, qnn_in_670, ddout__671, qq_in671, ddout__672, qq_in672, ddout__673, qq_in673, ddout__674, qq_in674, ddout__675, qq_in675, ddout__676, qq_in676, ddout__677, qq_in677, ddout__678, qq_in678, ddout__679, qq_in679, ddout__680, qq_in680, ddout__681, qq_in681, ddout__682, qq_in682, ddout__683, qq_in683, ddout__684, qq_in684, ddout__685, qq_in685, ddout__686, qq_in686, ddout__687, qq_in687, ddout__688, qq_in688, ddout__689, qq_in689, ddout__690, qq_in690, ddout__691, qq_in691, ddout__692, qq_in692, ddout__693, qq_in693, ddout__694, qq_in694, ddout__695, qq_in695, ddout__696, qq_in696, ddout__697, qq_in697, ddout__698, qq_in698, ddout__699, qq_in699, ddout__700, qq_in700, ddout__701, qq_in701, ddout__702, qq_in702, ddout__703, qq_in703, ddout__704, qq_in704, ddout__705, qq_in705, ddout__706, qq_in706, ddout__707, qq_in707, ddout__708, qq_in708, ddout__709, qq_in709, ddout__710, qq_in710, ddout__711, qq_in711, ddout__712, qq_in712, ddout__713, qq_in713, ddout__714, qq_in714, ddout__715, qq_in715, ddout__716, qq_in716, ddout__717, qq_in717, ddout__718, qq_in718, ddout__719, qq_in719, ddout__720, qq_in720, ddout__721, qq_in721, ddout__722, qq_in722, ddout__723, qq_in723, ddout__724, qq_in724, ddout__725, qq_in725, ddout__726, qq_in726, ddout__727, qq_in727, ddout__728, qq_in728, ddout__729, qq_in729, ddout__730, qq_in730, ddout__731, qq_in731, ddout__732, qq_in732, ddout__733, qq_in733, ddout__734, qq_in734, ddout__735, qq_in735, ddout__736, qq_in736, ddout__737, qq_in737, ddout__738, qq_in738, ddout__739, qq_in739, ddout__740, qq_in740, ddout__741, qq_in741, ddout__742, qq_in742, ddout__743, qq_in743, ddout__744, qq_in744, ddout__745, qq_in745, ddout__746, qq_in746, ddout__747, qq_in747, ddout__748, qq_in748, ddout__749, qq_in749, ddout__750, qq_in750, ddout__751, qq_in751, ddout__752, qq_in752, ddout__753, qq_in753, ddout__754, qq_in754, ddout__755, qq_in755, ddout__756, qq_in756, ddout__757, qq_in757, ddout__758, qq_in758, ddout__759, qq_in759, ddout__760, qq_in760, qnn_in_760, ddout__761, qq_in761, qnn_in_761, ddout__762, qq_in762, qnn_in_762, ddout__763, qq_in763, qnn_in_763, ddout__764, qq_in764, qnn_in_764, ddout__765, qq_in765, ddout__766, qq_in766, qnn_in_766, ddout__767, qq_in767, qnn_in_767, ddout__768, qq_in768, qnn_in_768, ddout__769, qq_in769, ddout__770, qq_in770, ddout__771, qq_in771, ddout__772, qq_in772, ddout__773, qq_in773, ddout__774, qq_in774, ddout__775, qq_in775, ddout__776, qq_in776, ddout__777, qq_in777, qnn_in_777, ddout__778, qq_in778, qnn_in_778, ddout__779, qq_in779, qnn_in_779, ddout__780, qq_in780, qnn_in_780, ddout__781, qq_in781, ddout__782, qq_in782, ddout__783, qq_in783, ddout__784, qq_in784, ddout__785, qq_in785, ddout__786, qq_in786, ddout__787, qq_in787, ddout__788, qq_in788, ddout__789, qq_in789, ddout__790, qq_in790, ddout__791, qq_in791, ddout__792, qq_in792, ddout__793, qq_in793, ddout__794, qq_in794, ddout__795, qq_in795, ddout__796, qq_in796, ddout__797, qq_in797, ddout__798, qq_in798, ddout__799, qq_in799, ddout__800, qq_in800, ddout__801, qq_in801, ddout__802, qq_in802, ddout__803, qq_in803, ddout__804, qq_in804, ddout__805, qq_in805, ddout__806, qq_in806, ddout__807, qq_in807, ddout__808, qq_in808, ddout__809, qq_in809, ddout__810, qq_in810, ddout__811, qq_in811, ddout__812, qq_in812, ddout__813, qq_in813, ddout__814, qq_in814, ddout__815, qq_in815, ddout__816, qq_in816, ddout__817, qq_in817, ddout__818, qq_in818, ddout__819, qq_in819, ddout__820, qq_in820, ddout__821, qq_in821, ddout__822, qq_in822, ddout__823, qq_in823, ddout__824, qq_in824, ddout__825, qq_in825, ddout__826, qq_in826, ddout__827, qq_in827, ddout__828, qq_in828, ddout__829, qq_in829, ddout__830, qq_in830, ddout__831, qq_in831, ddout__832, qq_in832, ddout__833, qq_in833, ddout__834, qq_in834, ddout__835, qq_in835, ddout__836, qq_in836, ddout__837, qq_in837, ddout__838, qq_in838, ddout__839, qq_in839, ddout__840, qq_in840, ddout__841, qq_in841, ddout__842, qq_in842, ddout__843, qq_in843, ddout__844, qq_in844, ddout__845, qq_in845, ddout__846, qq_in846, ddout__847, qq_in847, ddout__848, qq_in848, ddout__849, qq_in849, ddout__850, qq_in850, ddout__851, qq_in851, ddout__852, qq_in852, ddout__853, qq_in853, ddout__854, qq_in854, ddout__855, qq_in855, ddout__856, qq_in856, ddout__857, qq_in857, ddout__858, qq_in858, ddout__859, qq_in859, ddout__860, qq_in860, ddout__861, qq_in861, ddout__862, qq_in862, ddout__863, qq_in863, ddout__864, qq_in864, ddout__865, qq_in865, ddout__866, qq_in866, ddout__867, qq_in867, ddout__868, qq_in868, ddout__869, qq_in869, ddout__870, qq_in870, ddout__871, qq_in871, ddout__872, qq_in872, ddout__873, qq_in873, ddout__874, qq_in874, ddout__875, qq_in875, ddout__876, qq_in876, ddout__877, qq_in877, ddout__878, qq_in878, ddout__879, qq_in879, ddout__880, qq_in880, ddout__881, qq_in881, ddout__882, qq_in882, ddout__883, qq_in883, ddout__884, qq_in884, ddout__885, qq_in885, ddout__886, qq_in886, ddout__887, qq_in887, ddout__888, qq_in888, ddout__889, qq_in889, ddout__890, qq_in890, ddout__891, qq_in891, ddout__892, qq_in892, ddout__893, qq_in893, ddout__894, qq_in894, ddout__895, qq_in895, ddout__896, qq_in896, ddout__897, qq_in897, ddout__898, qq_in898, ddout__899, qq_in899, ddout__900, qq_in900, ddout__901, qq_in901, ddout__902, qq_in902, ddout__903, qq_in903, ddout__904, qq_in904, ddout__905, qq_in905, ddout__906, qq_in906, ddout__907, qq_in907, ddout__908, qq_in908, ddout__909, qq_in909, ddout__910, qq_in910, ddout__911, qq_in911, ddout__912, qq_in912, ddout__913, qq_in913, ddout__914, qq_in914, ddout__915, qq_in915, ddout__916, qq_in916, ddout__917, qq_in917, ddout__918, qq_in918, ddout__919, qq_in919, ddout__920, qq_in920, ddout__921, qq_in921, ddout__922, qq_in922, ddout__923, qq_in923, ddout__924, qq_in924, ddout__925, qq_in925, ddout__926, qq_in926, ddout__927, qq_in927, ddout__928, qq_in928, ddout__929, qq_in929, ddout__930, qq_in930, ddout__931, qq_in931, ddout__932, qq_in932, ddout__933, qq_in933, ddout__934, qq_in934, ddout__935, qq_in935, ddout__936, qq_in936, ddout__937, qq_in937, ddout__938, qq_in938, ddout__939, qq_in939, ddout__940, qq_in940, ddout__941, qq_in941, ddout__942, qq_in942, ddout__943, qq_in943, ddout__944, qq_in944, ddout__945, qq_in945, ddout__946, qq_in946, ddout__947, qq_in947, ddout__948, qq_in948, ddout__949, qq_in949, ddout__950, qq_in950, ddout__951, qq_in951, ddout__952, qq_in952, ddout__953, qq_in953, ddout__954, qq_in954, ddout__955, qq_in955, ddout__956, qq_in956, ddout__957, qq_in957, ddout__958, qq_in958, ddout__959, qq_in959, ddout__960, qq_in960, ddout__961, qq_in961, ddout__962, qq_in962, ddout__963, qq_in963, ddout__964, qq_in964, ddout__965, qq_in965, ddout__966, qq_in966, ddout__967, qq_in967, ddout__968, qq_in968, ddout__969, qq_in969, ddout__970, qq_in970, ddout__971, qq_in971, ddout__972, qq_in972, ddout__973, qq_in973, ddout__974, qq_in974, ddout__975, qq_in975, ddout__976, qq_in976, ddout__977, qq_in977, ddout__978, qq_in978, ddout__979, qq_in979, ddout__980, qq_in980, ddout__981, qq_in981, ddout__982, qq_in982, ddout__983, qq_in983, ddout__984, qq_in984, ddout__985, qq_in985, ddout__986, qq_in986, ddout__987, qq_in987, ddout__988, qq_in988, ddout__989, qq_in989, ddout__990, qq_in990, ddout__991, qq_in991, ddout__992, qq_in992, ddout__993, qq_in993, ddout__994, qq_in994, ddout__995, qq_in995, ddout__996, qq_in996, ddout__997, qq_in997, ddout__998, qq_in998, ddout__999, qq_in999, ddout__1000, qq_in1000, ddout__1001, qq_in1001, ddout__1002, qq_in1002, ddout__1003, qq_in1003, ddout__1004, qq_in1004, ddout__1005, qq_in1005, ddout__1006, qq_in1006, ddout__1007, qq_in1007, ddout__1008, qq_in1008, ddout__1009, qq_in1009, ddout__1010, qq_in1010, ddout__1011, qq_in1011, ddout__1012, qq_in1012, ddout__1013, qq_in1013, ddout__1014, qq_in1014, ddout__1015, qq_in1015, ddout__1016, qq_in1016, ddout__1017, qq_in1017, ddout__1018, qq_in1018, ddout__1019, qq_in1019, ddout__1020, qq_in1020, ddout__1021, qq_in1021, ddout__1022, qq_in1022, ddout__1023, qq_in1023, ddout__1024, qq_in1024, ddout__1025, qq_in1025, ddout__1026, qq_in1026, ddout__1027, qq_in1027, ddout__1028, qq_in1028, ddout__1029, qq_in1029, ddout__1030, qq_in1030, ddout__1031, qq_in1031, ddout__1032, qq_in1032, ddout__1033, qq_in1033, ddout__1034, qq_in1034, ddout__1035, qq_in1035, ddout__1036, qq_in1036, ddout__1037, qq_in1037, ddout__1038, qq_in1038, ddout__1039, qq_in1039, ddout__1040, qq_in1040, ddout__1041, qq_in1041, ddout__1042, qq_in1042, ddout__1043, qq_in1043, ddout__1044, qq_in1044, ddout__1045, qq_in1045, ddout__1046, qq_in1046, ddout__1047, qq_in1047, ddout__1048, qq_in1048, ddout__1049, qq_in1049, ddout__1050, qq_in1050, ddout__1051, qq_in1051, ddout__1052, qq_in1052, ddout__1053, qq_in1053, ddout__1054, qq_in1054, ddout__1055, qq_in1055, ddout__1056, qq_in1056, ddout__1057, qq_in1057, ddout__1058, qq_in1058, ddout__1059, qq_in1059, ddout__1060, qq_in1060, ddout__1061, qq_in1061, ddout__1062, qq_in1062, ddout__1063, qq_in1063, ddout__1064, qq_in1064, ddout__1065, qq_in1065, ddout__1066, qq_in1066, ddout__1067, qq_in1067, ddout__1068, qq_in1068, ddout__1069, qq_in1069, ddout__1070, qq_in1070, ddout__1071, qq_in1071, ddout__1072, qq_in1072, ddout__1073, qq_in1073, ddout__1074, qq_in1074, ddout__1075, qq_in1075, ddout__1076, qq_in1076, ddout__1077, qq_in1077, ddout__1078, qq_in1078, ddout__1079, qq_in1079, ddout__1080, qq_in1080, ddout__1081, qq_in1081, ddout__1082, qq_in1082, ddout__1083, qq_in1083, ddout__1084, qq_in1084, ddout__1085, qq_in1085, ddout__1086, qq_in1086, ddout__1087, qq_in1087, ddout__1088, qq_in1088, ddout__1089, qq_in1089, ddout__1090, qq_in1090, ddout__1091, qq_in1091, ddout__1092, qq_in1092, ddout__1093, qq_in1093, ddout__1094, qq_in1094, ddout__1095, qq_in1095, ddout__1096, qq_in1096, ddout__1097, qq_in1097, ddout__1098, qq_in1098, ddout__1099, qq_in1099, ddout__1100, qq_in1100, ddout__1101, qq_in1101, ddout__1102, qq_in1102, ddout__1103, qq_in1103, ddout__1104, qq_in1104, ddout__1105, qq_in1105, ddout__1106, qq_in1106, ddout__1107, qq_in1107, ddout__1108, qq_in1108, ddout__1109, qq_in1109, ddout__1110, qq_in1110, ddout__1111, qq_in1111, ddout__1112, qq_in1112, ddout__1113, qq_in1113, ddout__1114, qq_in1114, ddout__1115, qq_in1115, ddout__1116, qq_in1116, ddout__1117, qq_in1117, ddout__1118, qq_in1118, ddout__1119, qq_in1119, ddout__1120, qq_in1120, ddout__1121, qq_in1121, ddout__1122, qq_in1122, ddout__1123, qq_in1123, ddout__1124, qq_in1124, ddout__1125, qq_in1125, ddout__1126, qq_in1126, ddout__1127, qq_in1127, ddout__1128, qq_in1128, ddout__1129, qq_in1129, ddout__1130, qq_in1130, ddout__1131, qq_in1131, ddout__1132, qq_in1132, ddout__1133, qq_in1133, ddout__1134, qq_in1134, ddout__1135, qq_in1135, ddout__1136, qq_in1136, ddout__1137, qq_in1137, ddout__1138, qq_in1138, ddout__1139, qq_in1139, ddout__1140, qq_in1140, ddout__1141, qq_in1141, ddout__1142, qq_in1142, ddout__1143, qq_in1143, ddout__1144, qq_in1144, ddout__1145, qq_in1145, ddout__1146, qq_in1146, ddout__1147, qq_in1147, ddout__1148, qq_in1148, ddout__1149, qq_in1149, ddout__1150, qq_in1150, ddout__1151, qq_in1151, ddout__1152, qq_in1152, ddout__1153, qq_in1153, ddout__1154, qq_in1154, ddout__1155, qq_in1155, ddout__1156, qq_in1156, ddout__1157, qq_in1157, ddout__1158, qq_in1158, ddout__1159, qq_in1159, ddout__1160, qq_in1160, ddout__1161, qq_in1161, ddout__1162, qq_in1162, ddout__1163, qq_in1163, ddout__1164, qq_in1164, ddout__1165, qq_in1165, ddout__1166, qq_in1166, ddout__1167, qq_in1167, ddout__1168, qq_in1168, ddout__1169, qq_in1169, ddout__1170, qq_in1170, ddout__1171, qq_in1171, ddout__1172, qq_in1172, ddout__1173, qq_in1173, ddout__1174, qq_in1174, ddout__1175, qq_in1175, ddout__1176, qq_in1176, ddout__1177, qq_in1177, ddout__1178, qq_in1178, ddout__1179, qq_in1179, ddout__1180, qq_in1180, ddout__1181, qq_in1181, ddout__1182, qq_in1182, ddout__1183, qq_in1183, ddout__1184, qq_in1184, ddout__1185, qq_in1185, ddout__1186, qq_in1186, ddout__1187, qq_in1187, ddout__1188, qq_in1188, ddout__1189, qq_in1189, ddout__1190, qq_in1190, ddout__1191, qq_in1191, ddout__1192, qq_in1192, ddout__1193, qq_in1193, ddout__1194, qq_in1194, ddout__1195, qq_in1195, ddout__1196, qq_in1196, ddout__1197, qq_in1197, ddout__1198, qq_in1198, ddout__1199, qq_in1199, ddout__1200, qq_in1200, ddout__1201, qq_in1201, ddout__1202, qq_in1202, ddout__1203, qq_in1203, ddout__1204, qq_in1204, ddout__1205, qq_in1205, ddout__1206, qq_in1206, ddout__1207, qq_in1207, ddout__1208, qq_in1208, ddout__1209, qq_in1209, ddout__1210, qq_in1210, ddout__1211, qq_in1211, ddout__1212, qq_in1212, ddout__1213, qq_in1213, ddout__1214, qq_in1214, ddout__1215, qq_in1215, ddout__1216, qq_in1216, ddout__1217, qq_in1217, ddout__1218, qq_in1218, ddout__1219, qq_in1219, ddout__1220, qq_in1220, ddout__1221, qq_in1221, ddout__1222, qq_in1222, ddout__1223, qq_in1223, ddout__1224, qq_in1224, ddout__1225, qq_in1225, ddout__1226, qq_in1226, ddout__1227, qq_in1227, ddout__1228, qq_in1228, ddout__1229, qq_in1229, ddout__1230, qq_in1230, ddout__1231, qq_in1231, ddout__1232, qq_in1232, ddout__1233, qq_in1233, ddout__1234, qq_in1234, ddout__1235, qq_in1235, ddout__1236, qq_in1236, ddout__1237, qq_in1237, ddout__1238, qq_in1238, ddout__1239, qq_in1239, ddout__1240, qq_in1240, ddout__1241, qq_in1241, ddout__1242, qq_in1242, ddout__1243, qq_in1243, ddout__1244, qq_in1244, ddout__1245, qq_in1245, ddout__1246, qq_in1246, ddout__1247, qq_in1247, ddout__1248, qq_in1248, ddout__1249, qq_in1249, ddout__1250, qq_in1250, ddout__1251, qq_in1251, ddout__1252, qq_in1252, ddout__1253, qq_in1253, ddout__1254, qq_in1254, ddout__1255, qq_in1255, ddout__1256, qq_in1256, ddout__1257, qq_in1257, ddout__1258, qq_in1258, ddout__1259, qq_in1259, ddout__1260, qq_in1260, ddout__1261, qq_in1261, ddout__1262, qq_in1262, ddout__1263, qq_in1263, ddout__1264, qq_in1264, ddout__1265, qq_in1265, ddout__1266, qq_in1266, ddout__1267, qq_in1267, ddout__1268, qq_in1268, ddout__1269, qq_in1269, ddout__1270, qq_in1270, ddout__1271, qq_in1271, ddout__1272, qq_in1272, ddout__1273, qq_in1273, ddout__1274, qq_in1274, ddout__1275, qq_in1275, ddout__1276, qq_in1276, ddout__1277, qq_in1277, ddout__1278, qq_in1278, ddout__1279, qq_in1279, ddout__1280, qq_in1280, ddout__1281, qq_in1281, ddout__1282, qq_in1282, ddout__1283, qq_in1283, ddout__1284, qq_in1284, ddout__1285, qq_in1285, ddout__1286, qq_in1286, ddout__1287, qq_in1287, ddout__1288, qq_in1288, ddout__1289, qq_in1289, ddout__1290, qq_in1290, ddout__1291, qq_in1291, ddout__1292, qq_in1292, ddout__1293, qq_in1293, ddout__1294, qq_in1294, ddout__1295, qq_in1295, ddout__1296, qq_in1296, ddout__1297, qq_in1297, ddout__1298, qq_in1298, ddout__1299, qq_in1299, ddout__1300, qq_in1300, ddout__1301, qnn_in_1301, ddout__1302, qq_in1302, ddout__1303, qq_in1303, qnn_in_1303, ddout__1304, qq_in1304, ddout__1305, qq_in1305, d_out_1, q_in_1, d_out_2, q_in_2, d_out_3, q_in_3, d_out_4, q_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, q_in_7, d_out_8, q_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, d_out_12, q_in_12, d_out_13, q_in_13, d_out_14, q_in_14, d_out_15, q_in_15, d_out_16, q_in_16, d_out_17, q_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, q_in_20, d_out_21, q_in_21, d_out_22, q_in_22, d_out_23, q_in_23, d_out_24, q_in_24, d_out_25, q_in_25, d_out_26, q_in_26, d_out_27, q_in_27, d_out_28, q_in_28, d_out_29, q_in_29, d_out_30, q_in_30, d_out_31, q_in_31, d_out_32, q_in_32, d_out_33, q_in_33, d_out_34, q_in_34, d_out_35, q_in_35, d_out_36, q_in_36, d_out_37, q_in_37, d_out_38, q_in_38, d_out_39, q_in_39, d_out_40, q_in_40, d_out_41, q_in_41, d_out_42, q_in_42, d_out_43, q_in_43, d_out_44, q_in_44, d_out_45, q_in_45, d_out_46, q_in_46, d_out_47, q_in_47, d_out_48, q_in_48, d_out_49, q_in_49, d_out_50, q_in_50, d_out_51, q_in_51, d_out_52, q_in_52, d_out_53, q_in_53, d_out_54, q_in_54, d_out_55, q_in_55, d_out_56, q_in_56, d_out_57, q_in_57, d_out_58, q_in_58, d_out_59, q_in_59, d_out_60, q_in_60, d_out_61, q_in_61, d_out_62, q_in_62, d_out_63, q_in_63, d_out_64, q_in_64, d_out_65, q_in_65, d_out_66, q_in_66, d_out_67, q_in_67, d_out_68, q_in_68, d_out_69, q_in_69, d_out_70, q_in_70, d_out_71, q_in_71, d_out_72, q_in_72, d_out_73, q_in_73, d_out_74, q_in_74, d_out_75, q_in_75, d_out_76, q_in_76, d_out_77, q_in_77, d_out_78, q_in_78, d_out_79, q_in_79, d_out_80, q_in_80, d_out_81, q_in_81, d_out_82, q_in_82, d_out_83, q_in_83, d_out_84, qn_in_84, d_out_85, qn_in_85, d_out_86, qn_in_86, d_out_87, qn_in_87, d_out_88, qn_in_88, d_out_89, qn_in_89, d_out_90, qn_in_90, d_out_91, qn_in_91, d_out_92, qn_in_92, d_out_93, qn_in_93, d_out_94, qn_in_94, d_out_95, qn_in_95, d_out_96, qn_in_96, d_out_97, qn_in_97, d_out_98, qn_in_98, d_out_99, qn_in_99, d_out_100, qn_in_100, d_out_101, qn_in_101, d_out_102, qn_in_102, d_out_103, qn_in_103, d_out_104, qn_in_104, d_out_105, qn_in_105, d_out_106, qn_in_106, d_out_107, qn_in_107, d_out_108, qn_in_108, d_out_109, qn_in_109, d_out_110, qn_in_110, d_out_111, qn_in_111, d_out_112, qn_in_112, d_out_113, qn_in_113, d_out_114, qn_in_114, d_out_115, qn_in_115, d_out_116, qn_in_116, d_out_117, qn_in_117, d_out_118, qn_in_118, d_out_119, qn_in_119, d_out_120, qn_in_120, d_out_121, qn_in_121, d_out_122, qn_in_122, d_out_123, qn_in_123, d_out_124, qn_in_124, d_out_125, qn_in_125, d_out_126, qn_in_126, d_out_127, qn_in_127, d_out_128, qn_in_128, d_out_129, qn_in_129, d_out_130, qn_in_130, d_out_131, qn_in_131, d_out_132, qn_in_132, d_out_133, qn_in_133, d_out_134, qn_in_134, d_out_135, qn_in_135, d_out_136, qn_in_136, d_out_137, qn_in_137, d_out_138, qn_in_138, d_out_139, qn_in_139, d_out_140, qn_in_140, d_out_141, qn_in_141, d_out_142, qn_in_142, d_out_143, qn_in_143, d_out_144, qn_in_144, d_out_145, qn_in_145, d_out_146, qn_in_146, d_out_147, qn_in_147, d_out_148, qn_in_148, d_out_149, qn_in_149, d_out_150, qn_in_150, d_out_151, qn_in_151, d_out_152, qn_in_152, d_out_153, qn_in_153, d_out_154, qn_in_154, d_out_155, qn_in_155, d_out_156, qn_in_156, d_out_157, qn_in_157, d_out_158, qn_in_158, d_out_159, qn_in_159, d_out_160, qn_in_160, d_out_161, qn_in_161, d_out_162, qn_in_162, d_out_163, qn_in_163, d_out_164, qn_in_164, d_out_165, qn_in_165, d_out_166, qn_in_166, d_out_167, qn_in_167, d_out_168, qn_in_168, d_out_169, qn_in_169, d_out_170, qn_in_170, d_out_171, qn_in_171, d_out_172, qn_in_172, d_out_173, qn_in_173, d_out_174, qn_in_174, d_out_175, qn_in_175, d_out_176, qn_in_176, d_out_177, qn_in_177, d_out_178, qn_in_178, d_out_179, qn_in_179, d_out_180, qn_in_180, d_out_181, qn_in_181, d_out_182, qn_in_182, d_out_183, qn_in_183, d_out_184, qn_in_184, d_out_185, qn_in_185, d_out_186, qn_in_186, d_out_187, qn_in_187, d_out_188, qn_in_188, d_out_189, qn_in_189, d_out_190, qn_in_190, d_out_191, qn_in_191, d_out_192, q_in_192, qn_in_192, d_out_193, q_in_193, qn_in_193, d_out_194, q_in_194, qn_in_194, d_out_195, q_in_195, qn_in_195, d_out_196, q_in_196, d_out_197, q_in_197, qn_in_197, d_out_198, q_in_198, qn_in_198, d_out_199, q_in_199, d_out_200, q_in_200, d_out_201, q_in_201, d_out_202, q_in_202, d_out_203, q_in_203, d_out_204, q_in_204, d_out_205, q_in_205, d_out_206, q_in_206, qn_in_206, d_out_207, q_in_207, qn_in_207, d_out_208, q_in_208, qn_in_208, d_out_209, q_in_209, d_out_210, q_in_210, qn_in_210, d_out_211, q_in_211, d_out_212, q_in_212, d_out_213, q_in_213, d_out_214, q_in_214, d_out_215, q_in_215, d_out_216, q_in_216, d_out_217, q_in_217, d_out_218, q_in_218, d_out_219, q_in_219, d_out_220, q_in_220, d_out_221, q_in_221, d_out_222, q_in_222, d_out_223, q_in_223, qn_in_223, d_out_224, q_in_224, d_out_225, q_in_225, d_out_226, q_in_226, d_out_227, q_in_227, d_out_228, q_in_228, d_out_229, q_in_229, d_out_230, q_in_230, d_out_231, q_in_231, d_out_232, q_in_232, d_out_233, q_in_233, d_out_234, q_in_234, d_out_235, q_in_235, d_out_236, q_in_236, d_out_237, q_in_237, d_out_238, q_in_238, qn_in_238, d_out_239, q_in_239, d_out_240, q_in_240, qn_in_240, d_out_241, q_in_241, d_out_242, q_in_242, d_out_243, q_in_243, d_out_244, q_in_244, d_out_245, q_in_245, qn_in_245, d_out_246, q_in_246, d_out_247, q_in_247, d_out_248, q_in_248, d_out_249, q_in_249, qn_in_249, d_out_250, q_in_250, qn_in_250, d_out_251, q_in_251, d_out_252, q_in_252, d_out_253, q_in_253, d_out_254, q_in_254, d_out_255, q_in_255, d_out_256, q_in_256, d_out_257, q_in_257, d_out_258, q_in_258, qn_in_258, d_out_259, q_in_259, qn_in_259, d_out_260, q_in_260, qn_in_260, d_out_261, q_in_261, d_out_262, q_in_262, d_out_263, q_in_263, d_out_264, q_in_264, d_out_265, q_in_265, d_out_266, q_in_266, d_out_267, q_in_267, d_out_268, q_in_268, d_out_269, q_in_269, d_out_270, q_in_270, d_out_271, q_in_271, d_out_272, q_in_272, d_out_273, q_in_273, d_out_274, q_in_274, qn_in_274, d_out_275, q_in_275, d_out_276, q_in_276, d_out_277, q_in_277, d_out_278, q_in_278, qn_in_278, d_out_279, q_in_279, qn_in_279, d_out_280, q_in_280, d_out_281, q_in_281, d_out_282, q_in_282, d_out_283, q_in_283, d_out_284, q_in_284, d_out_285, q_in_285, d_out_286, q_in_286, qn_in_286, d_out_287, q_in_287, qn_in_287, d_out_288, q_in_288, d_out_289, q_in_289, qn_in_289, d_out_290, q_in_290, d_out_291, q_in_291, d_out_292, q_in_292, d_out_293, q_in_293, d_out_294, q_in_294, d_out_295, q_in_295, qn_in_295, d_out_296, q_in_296, d_out_297, q_in_297, qn_in_297, d_out_298, q_in_298, qn_in_298, d_out_299, q_in_299, d_out_300, q_in_300, d_out_301, q_in_301, d_out_302, q_in_302, d_out_303, q_in_303, d_out_304, q_in_304, d_out_305, q_in_305, d_out_306, q_in_306, d_out_307, q_in_307, d_out_308, q_in_308, d_out_309, q_in_309, d_out_310, q_in_310, d_out_311, q_in_311, d_out_312, q_in_312, d_out_313, q_in_313, qn_in_313, d_out_314, q_in_314, qn_in_314, d_out_315, q_in_315, qn_in_315, d_out_316, q_in_316, d_out_317, q_in_317, d_out_318, q_in_318, d_out_319, q_in_319, d_out_320, q_in_320, d_out_321, q_in_321, d_out_322, q_in_322, qn_in_322, d_out_323, q_in_323, qn_in_323, d_out_324, q_in_324, qn_in_324, d_out_325, q_in_325, qn_in_325, d_out_326, q_in_326, qn_in_326, d_out_327, q_in_327, qn_in_327, d_out_328, q_in_328, qn_in_328, d_out_329, q_in_329, qn_in_329, d_out_330, q_in_330, d_out_331, q_in_331, d_out_332, q_in_332, d_out_333, q_in_333, d_out_334, q_in_334, d_out_335, q_in_335, d_out_336, q_in_336, d_out_337, q_in_337, d_out_338, q_in_338, d_out_339, q_in_339, d_out_340, q_in_340, d_out_341, q_in_341, d_out_342, q_in_342, d_out_343, q_in_343, d_out_344, q_in_344, d_out_345, q_in_345, d_out_346, q_in_346, d_out_347, q_in_347, d_out_348, q_in_348, d_out_349, q_in_349, d_out_350, q_in_350, d_out_351, q_in_351, d_out_352, q_in_352, d_out_353, q_in_353, d_out_354, q_in_354, d_out_355, q_in_355, d_out_356, q_in_356, d_out_357, q_in_357, d_out_358, q_in_358, d_out_359, q_in_359, d_out_360, q_in_360, d_out_361, q_in_361, d_out_362, q_in_362, d_out_363, q_in_363, d_out_364, q_in_364, d_out_365, q_in_365, d_out_366, q_in_366, d_out_367, q_in_367, d_out_368, q_in_368, d_out_369, q_in_369, d_out_370, q_in_370, d_out_371, q_in_371, d_out_372, q_in_372, d_out_373, q_in_373, d_out_374, q_in_374, d_out_375, qn_in_375, d_out_376, qn_in_376, d_out_377, qn_in_377, d_out_378, qn_in_378, d_out_379, qn_in_379, d_out_380, qn_in_380, d_out_381, qn_in_381, d_out_382, qn_in_382, d_out_383, qn_in_383, d_out_384, qn_in_384, d_out_385, qn_in_385, d_out_386, qn_in_386, d_out_387, qn_in_387, d_out_388, qn_in_388, d_out_389, qn_in_389, d_out_390, qn_in_390, d_out_391, qn_in_391, d_out_392, qn_in_392, d_out_393, qn_in_393, d_out_394, qn_in_394, d_out_395, q_in_395, d_out_396, q_in_396, qn_in_396, d_out_397, q_in_397, qn_in_397, d_out_398, q_in_398, qn_in_398);
input qn_in_210;
input qn_in_208;
input qn_in_207;
input qn_in_206;
input qn_in_198;
input qn_in_197;
input qn_in_195;
input qn_in_194;
input qn_in_193;
input qn_in_192;
input qn_in_191;
input qn_in_190;
input qn_in_189;
input qn_in_188;
input qn_in_187;
input qn_in_186;
input qn_in_185;
input qn_in_184;
input qn_in_183;
input qn_in_182;
input qn_in_181;
input qn_in_180;
input qn_in_179;
input qn_in_178;
input qn_in_177;
input qn_in_176;
input qn_in_175;
input qn_in_174;
input qn_in_173;
input qn_in_172;
input qn_in_171;
input qn_in_170;
input qn_in_169;
input qn_in_168;
input qn_in_167;
input qn_in_166;
input qn_in_165;
input qn_in_164;
input qn_in_163;
input qn_in_162;
input qn_in_161;
input qn_in_160;
input qn_in_159;
input qn_in_158;
input qn_in_157;
input qn_in_156;
input qn_in_155;
input qn_in_154;
input qn_in_153;
input qn_in_152;
input qn_in_151;
input qn_in_150;
input qn_in_149;
input qn_in_148;
input qn_in_147;
input qn_in_146;
input qn_in_145;
input qn_in_144;
input qn_in_143;
input qn_in_142;
input qn_in_141;
input qn_in_140;
input qn_in_139;
input qn_in_138;
input qn_in_137;
input qn_in_136;
input qn_in_135;
input qn_in_134;
input qn_in_133;
input qn_in_132;
input qn_in_131;
input qn_in_130;
input qn_in_129;
input qn_in_128;
input qn_in_127;
input qn_in_126;
input qn_in_125;
input qn_in_124;
input qn_in_123;
input qn_in_122;
input qn_in_121;
input qn_in_120;
input qn_in_119;
input qn_in_118;
input qn_in_117;
input qn_in_116;
input qn_in_115;
input qn_in_114;
input qn_in_113;
input qn_in_112;
input qn_in_111;
input qn_in_110;
input qn_in_109;
input qn_in_108;
input qn_in_107;
input qn_in_106;
input qn_in_105;
input qn_in_104;
input qn_in_103;
input qn_in_102;
input qn_in_101;
input qn_in_100;
input qn_in_99;
input qn_in_98;
input qn_in_97;
input qn_in_96;
input qn_in_95;
input qn_in_94;
input qn_in_93;
input qn_in_92;
input qn_in_91;
input qn_in_90;
input qn_in_89;
input qn_in_88;
input qn_in_87;
input qn_in_86;
input qn_in_85;
input qn_in_84;
input qn_in_394;
input qn_in_393;
input qn_in_392;
input qn_in_391;
input qn_in_390;
input qn_in_389;
input qn_in_388;
input qn_in_387;
input qn_in_386;
input qn_in_385;
input qn_in_384;
input qn_in_383;
input qn_in_382;
input qn_in_381;
input qn_in_380;
input qn_in_379;
input qn_in_378;
input qn_in_377;
input qn_in_376;
input qn_in_375;
input qn_in_329;
input qn_in_328;
input qn_in_327;
input qn_in_326;
input qn_in_325;
input qn_in_324;
input qn_in_323;
input qn_in_322;
input qn_in_315;
input qn_in_314;
input qn_in_313;
input qn_in_298;
input qn_in_297;
input qn_in_295;
input qn_in_289;
input qn_in_287;
input qn_in_286;
input qn_in_279;
input qn_in_278;
input qn_in_274;
input qn_in_260;
input qn_in_259;
input qn_in_258;
input qn_in_250;
input qn_in_249;
input qn_in_245;
input qn_in_240;
input qn_in_238;
input qn_in_398;
input qn_in_397;
input qn_in_396;
input qn_in_223;
input q_in_211;
input q_in_210;
input q_in_209;
input q_in_208;
input q_in_207;
input q_in_206;
input q_in_205;
input q_in_204;
input q_in_203;
input q_in_202;
input q_in_201;
input q_in_200;
input q_in_199;
input q_in_198;
input q_in_197;
input q_in_196;
input q_in_195;
input q_in_194;
input q_in_193;
input q_in_192;
input q_in_83;
input q_in_82;
input q_in_81;
input q_in_80;
input q_in_79;
input q_in_78;
input q_in_77;
input q_in_76;
input q_in_75;
input q_in_74;
input q_in_73;
input q_in_72;
input q_in_71;
input q_in_70;
input q_in_69;
input q_in_68;
input q_in_67;
input q_in_66;
input q_in_65;
input q_in_64;
input q_in_63;
input q_in_62;
input q_in_61;
input q_in_60;
input q_in_59;
input q_in_58;
input q_in_57;
input q_in_56;
input q_in_55;
input q_in_54;
input q_in_53;
input q_in_52;
input q_in_51;
input q_in_50;
input q_in_49;
input q_in_48;
input q_in_47;
input q_in_46;
input q_in_45;
input q_in_44;
input q_in_43;
input q_in_42;
input q_in_41;
input q_in_40;
input q_in_39;
input q_in_38;
input q_in_37;
input q_in_36;
input q_in_35;
input q_in_34;
input q_in_33;
input q_in_32;
input q_in_31;
input q_in_30;
input q_in_29;
input q_in_28;
input q_in_27;
input q_in_26;
input q_in_25;
input q_in_24;
input q_in_23;
input q_in_22;
input q_in_21;
input q_in_20;
input q_in_19;
input q_in_18;
input q_in_17;
input q_in_16;
input q_in_15;
input q_in_14;
input q_in_13;
input q_in_12;
input q_in_11;
input q_in_10;
input q_in_9;
input q_in_8;
input q_in_7;
input q_in_6;
input q_in_5;
input q_in_4;
input q_in_3;
input q_in_2;
input q_in_1;
input q_in_398;
input q_in_395;
input q_in_397;
input q_in_396;
input q_in_374;
input q_in_373;
input q_in_372;
input q_in_371;
input q_in_370;
input q_in_369;
input q_in_368;
input q_in_367;
input q_in_366;
input q_in_365;
input q_in_364;
input q_in_363;
input q_in_362;
input q_in_361;
input q_in_360;
input q_in_359;
input q_in_358;
input q_in_357;
input q_in_356;
input q_in_355;
input q_in_354;
input q_in_353;
input q_in_352;
input q_in_351;
input q_in_350;
input q_in_349;
input q_in_348;
input q_in_347;
input q_in_346;
input q_in_345;
input q_in_344;
input q_in_343;
input q_in_342;
input q_in_341;
input q_in_340;
input q_in_339;
input q_in_338;
input q_in_337;
input q_in_336;
input q_in_335;
input q_in_334;
input q_in_333;
input q_in_332;
input q_in_331;
input q_in_330;
input q_in_329;
input q_in_328;
input q_in_327;
input q_in_326;
input q_in_325;
input q_in_324;
input q_in_323;
input q_in_322;
input q_in_321;
input q_in_320;
input q_in_319;
input q_in_318;
input q_in_317;
input q_in_316;
input q_in_315;
input q_in_314;
input q_in_313;
input q_in_312;
input q_in_311;
input q_in_310;
input q_in_309;
input q_in_308;
input q_in_307;
input q_in_306;
input q_in_305;
input q_in_304;
input q_in_303;
input q_in_302;
input q_in_301;
input q_in_300;
input q_in_299;
input q_in_298;
input q_in_297;
input q_in_296;
input q_in_295;
input q_in_294;
input q_in_293;
input q_in_292;
input q_in_291;
input q_in_290;
input q_in_289;
input q_in_288;
input q_in_287;
input q_in_286;
input q_in_285;
input q_in_284;
input q_in_283;
input q_in_282;
input q_in_281;
input q_in_280;
input q_in_279;
input q_in_278;
input q_in_277;
input q_in_276;
input q_in_275;
input q_in_274;
input q_in_273;
input q_in_272;
input q_in_271;
input q_in_270;
input q_in_269;
input q_in_268;
input q_in_267;
input q_in_266;
input q_in_265;
input q_in_264;
input q_in_263;
input q_in_262;
input q_in_261;
input q_in_260;
input q_in_259;
input q_in_258;
input q_in_257;
input q_in_256;
input q_in_255;
input q_in_254;
input q_in_253;
input q_in_252;
input q_in_251;
input q_in_250;
input q_in_249;
input q_in_248;
input q_in_247;
input q_in_246;
input q_in_245;
input q_in_244;
input q_in_243;
input q_in_242;
input q_in_241;
input q_in_240;
input q_in_239;
input q_in_238;
input q_in_237;
input q_in_236;
input q_in_235;
input q_in_234;
input q_in_233;
input q_in_232;
input q_in_231;
input q_in_230;
input q_in_229;
input q_in_228;
input q_in_227;
input q_in_226;
input q_in_225;
input q_in_224;
input q_in_223;
input q_in_222;
input q_in_221;
input q_in_220;
input q_in_219;
input q_in_218;
input q_in_217;
input q_in_216;
input q_in_215;
input q_in_214;
input q_in_213;
input q_in_212;
input [127:0] dii_data;
input [3:0] dii_data_size;
input [127:0] cii_K;
input clk, rst, dii_data_vld, dii_data_type, dii_last_word, cii_ctl_vld, cii_IV_vld;
input qq_in1;
input qq_in2;
input qq_in3;
input qq_in4;
input qq_in5;
input qq_in6;
input qq_in7;
input qq_in8;
input qq_in9;
input qq_in10;
input qq_in11;
input qq_in12;
input qq_in13;
input qq_in14;
input qq_in15;
input qq_in16;
input qq_in17;
input qq_in18;
input qq_in19;
input qq_in20;
input qq_in21;
input qq_in22;
input qq_in23;
input qq_in24;
input qq_in25;
input qq_in26;
input qq_in27;
input qq_in28;
input qq_in29;
input qq_in30;
input qq_in31;
input qq_in32;
input qq_in33;
input qq_in34;
input qq_in35;
input qq_in36;
input qq_in37;
input qq_in38;
input qq_in39;
input qq_in40;
input qq_in41;
input qq_in42;
input qq_in43;
input qq_in44;
input qq_in45;
input qq_in46;
input qq_in47;
input qq_in48;
input qq_in49;
input qq_in50;
input qq_in51;
input qq_in52;
input qq_in53;
input qq_in54;
input qq_in55;
input qq_in56;
input qq_in57;
input qq_in58;
input qq_in59;
input qq_in60;
input qq_in61;
input qq_in62;
input qq_in63;
input qq_in64;
input qq_in65;
input qq_in66;
input qq_in67;
input qq_in68;
input qq_in69;
input qq_in70;
input qq_in71;
input qq_in72;
input qq_in73;
input qq_in74;
input qq_in75;
input qq_in76;
input qq_in77;
input qq_in78;
input qq_in79;
input qq_in80;
input qq_in81;
input qq_in82;
input qq_in83;
input qq_in84;
input qq_in85;
input qq_in86;
input qq_in87;
input qq_in88;
input qq_in89;
input qq_in90;
input qq_in91;
input qq_in92;
input qq_in93;
input qq_in94;
input qq_in95;
input qq_in96;
input qq_in97;
input qq_in98;
input qq_in99;
input qq_in100;
input qq_in101;
input qq_in102;
input qq_in103;
input qq_in104;
input qq_in105;
input qq_in106;
input qq_in107;
input qq_in108;
input qq_in109;
input qq_in110;
input qq_in111;
input qq_in112;
input qq_in113;
input qq_in114;
input qq_in115;
input qq_in116;
input qq_in117;
input qq_in118;
input qq_in119;
input qq_in120;
input qq_in121;
input qq_in122;
input qq_in123;
input qq_in124;
input qq_in125;
input qq_in126;
input qq_in127;
input qq_in128;
input qq_in129;
input qq_in130;
input qq_in131;
input qq_in132;
input qq_in133;
input qq_in134;
input qq_in135;
input qq_in136;
input qq_in137;
input qq_in138;
input qq_in139;
input qq_in140;
input qq_in141;
input qq_in142;
input qq_in143;
input qq_in144;
input qq_in145;
input qq_in146;
input qq_in147;
input qq_in148;
input qq_in149;
input qq_in150;
input qq_in151;
input qq_in152;
input qq_in153;
input qq_in154;
input qq_in155;
input qq_in156;
input qq_in157;
input qq_in158;
input qq_in159;
input qq_in160;
input qq_in161;
input qq_in162;
input qq_in163;
input qq_in164;
input qq_in165;
input qq_in166;
input qq_in167;
input qq_in168;
input qq_in169;
input qq_in170;
input qq_in171;
input qq_in172;
input qq_in173;
input qq_in174;
input qq_in175;
input qq_in176;
input qq_in177;
input qq_in178;
input qq_in179;
input qq_in180;
input qq_in181;
input qq_in182;
input qq_in183;
input qq_in184;
input qq_in185;
input qq_in186;
input qq_in187;
input qq_in188;
input qq_in189;
input qq_in190;
input qq_in191;
input qq_in192;
input qq_in193;
input qq_in194;
input qq_in195;
input qq_in196;
input qq_in197;
input qq_in198;
input qq_in199;
input qq_in200;
input qq_in201;
input qq_in202;
input qq_in203;
input qq_in204;
input qq_in205;
input qq_in206;
input qq_in207;
input qq_in208;
input qq_in209;
input qq_in210;
input qq_in211;
input qq_in212;
input qq_in213;
input qq_in214;
input qq_in215;
input qq_in216;
input qq_in217;
input qq_in218;
input qq_in219;
input qq_in220;
input qq_in221;
input qq_in222;
input qq_in223;
input qq_in224;
input qq_in225;
input qq_in226;
input qq_in227;
input qq_in228;
input qq_in229;
input qq_in230;
input qq_in231;
input qq_in232;
input qq_in233;
input qq_in234;
input qq_in235;
input qq_in236;
input qq_in237;
input qq_in238;
input qq_in239;
input qq_in240;
input qq_in241;
input qq_in242;
input qq_in243;
input qq_in244;
input qq_in245;
input qq_in246;
input qq_in247;
input qq_in248;
input qq_in249;
input qq_in250;
input qq_in251;
input qq_in252;
input qq_in253;
input qq_in254;
input qq_in255;
input qq_in256;
input qq_in257;
input qq_in258;
input qq_in259;
input qq_in260;
input qq_in261;
input qq_in262;
input qq_in263;
input qq_in264;
input qq_in265;
input qq_in266;
input qq_in267;
input qq_in268;
input qq_in269;
input qq_in270;
input qq_in271;
input qq_in272;
input qq_in273;
input qq_in274;
input qq_in275;
input qq_in276;
input qq_in277;
input qq_in278;
input qq_in279;
input qq_in280;
input qq_in281;
input qq_in282;
input qq_in283;
input qq_in284;
input qq_in285;
input qq_in286;
input qq_in287;
input qq_in288;
input qq_in289;
input qq_in290;
input qq_in291;
input qq_in292;
input qq_in293;
input qq_in294;
input qq_in295;
input qq_in296;
input qq_in297;
input qq_in298;
input qq_in299;
input qq_in300;
input qq_in301;
input qq_in302;
input qq_in303;
input qq_in304;
input qq_in305;
input qq_in306;
input qq_in307;
input qq_in308;
input qq_in309;
input qq_in310;
input qq_in311;
input qq_in312;
input qq_in313;
input qq_in314;
input qq_in315;
input qq_in316;
input qq_in317;
input qq_in318;
input qq_in319;
input qq_in320;
input qq_in321;
input qq_in322;
input qq_in323;
input qq_in324;
input qq_in325;
input qq_in326;
input qq_in327;
input qq_in328;
input qq_in329;
input qq_in330;
input qq_in331;
input qq_in332;
input qq_in333;
input qq_in334;
input qq_in335;
input qq_in336;
input qq_in337;
input qq_in338;
input qq_in339;
input qq_in340;
input qq_in341;
input qq_in342;
input qq_in343;
input qq_in344;
input qq_in345;
input qq_in346;
input qq_in347;
input qq_in348;
input qq_in349;
input qq_in350;
input qq_in351;
input qq_in352;
input qq_in353;
input qq_in354;
input qq_in355;
input qq_in356;
input qq_in357;
input qq_in358;
input qq_in359;
input qq_in360;
input qq_in361;
input qq_in362;
input qq_in363;
input qq_in364;
input qq_in365;
input qq_in366;
input qq_in367;
input qq_in368;
input qq_in369;
input qq_in370;
input qq_in371;
input qq_in372;
input qq_in373;
input qq_in374;
input qq_in375;
input qq_in376;
input qq_in377;
input qq_in378;
input qq_in379;
input qq_in380;
input qq_in381;
input qq_in382;
input qq_in383;
input qq_in384;
input qq_in385;
input qq_in386;
input qq_in387;
input qq_in388;
input qq_in389;
input qq_in390;
input qq_in391;
input qq_in392;
input qq_in393;
input qq_in394;
input qq_in395;
input qq_in396;
input qq_in397;
input qq_in398;
input qq_in399;
input qq_in400;
input qq_in401;
input qq_in402;
input qq_in403;
input qq_in404;
input qq_in405;
input qq_in406;
input qq_in407;
input qq_in408;
input qq_in409;
input qq_in410;
input qq_in411;
input qq_in412;
input qq_in413;
input qq_in414;
input qq_in415;
input qq_in416;
input qq_in417;
input qq_in418;
input qq_in419;
input qq_in420;
input qq_in421;
input qq_in422;
input qq_in423;
input qq_in424;
input qq_in425;
input qq_in426;
input qq_in427;
input qq_in428;
input qq_in429;
input qq_in430;
input qq_in431;
input qq_in432;
input qq_in433;
input qq_in434;
input qq_in435;
input qq_in436;
input qq_in437;
input qq_in438;
input qq_in439;
input qq_in440;
input qq_in441;
input qq_in442;
input qq_in443;
input qq_in444;
input qq_in445;
input qq_in446;
input qq_in447;
input qq_in448;
input qq_in449;
input qq_in450;
input qq_in451;
input qq_in452;
input qq_in453;
input qq_in454;
input qq_in455;
input qq_in456;
input qq_in457;
input qq_in458;
input qq_in459;
input qq_in460;
input qq_in461;
input qq_in462;
input qq_in463;
input qq_in464;
input qq_in465;
input qq_in466;
input qq_in467;
input qq_in468;
input qq_in469;
input qq_in470;
input qq_in471;
input qq_in472;
input qq_in473;
input qq_in474;
input qq_in475;
input qq_in476;
input qq_in477;
input qq_in478;
input qq_in479;
input qq_in480;
input qq_in481;
input qq_in482;
input qq_in483;
input qq_in484;
input qq_in485;
input qq_in486;
input qq_in487;
input qq_in488;
input qq_in489;
input qq_in490;
input qq_in491;
input qq_in492;
input qq_in493;
input qq_in494;
input qq_in495;
input qq_in496;
input qq_in497;
input qq_in498;
input qq_in499;
input qq_in500;
input qq_in501;
input qq_in502;
input qq_in503;
input qq_in504;
input qq_in505;
input qq_in506;
input qq_in507;
input qq_in508;
input qq_in509;
input qq_in510;
input qq_in511;
input qq_in512;
input qq_in513;
input qq_in514;
input qq_in515;
input qq_in516;
input qq_in517;
input qq_in518;
input qq_in519;
input qq_in520;
input qq_in521;
input qq_in522;
input qq_in523;
input qq_in524;
input qq_in525;
input qq_in526;
input qq_in527;
input qq_in528;
input qq_in529;
input qq_in530;
input qq_in531;
input qq_in532;
input qq_in533;
input qq_in534;
input qq_in535;
input qq_in536;
input qq_in537;
input qq_in538;
input qq_in539;
input qq_in540;
input qq_in541;
input qq_in542;
input qq_in543;
input qq_in544;
input qq_in545;
input qq_in546;
input qq_in547;
input qq_in548;
input qq_in549;
input qq_in550;
input qq_in551;
input qq_in552;
input qq_in553;
input qq_in554;
input qq_in555;
input qq_in556;
input qq_in557;
input qq_in558;
input qq_in559;
input qq_in560;
input qq_in561;
input qq_in562;
input qq_in563;
input qq_in564;
input qq_in565;
input qq_in566;
input qq_in567;
input qq_in568;
input qq_in569;
input qq_in570;
input qq_in571;
input qq_in572;
input qq_in573;
input qq_in574;
input qq_in575;
input qq_in576;
input qq_in577;
input qq_in578;
input qq_in579;
input qq_in580;
input qq_in581;
input qq_in582;
input qq_in583;
input qq_in584;
input qq_in585;
input qq_in586;
input qq_in587;
input qq_in588;
input qq_in589;
input qq_in590;
input qq_in591;
input qq_in592;
input qq_in593;
input qq_in594;
input qq_in595;
input qq_in596;
input qq_in597;
input qq_in598;
input qq_in599;
input qq_in600;
input qq_in601;
input qq_in602;
input qq_in603;
input qq_in604;
input qq_in605;
input qq_in606;
input qq_in607;
input qq_in608;
input qq_in609;
input qq_in610;
input qq_in611;
input qq_in612;
input qq_in613;
input qq_in614;
input qq_in615;
input qq_in616;
input qq_in617;
input qq_in618;
input qq_in619;
input qq_in620;
input qq_in621;
input qq_in622;
input qq_in623;
input qq_in624;
input qq_in625;
input qq_in626;
input qq_in627;
input qq_in628;
input qq_in629;
input qq_in630;
input qq_in631;
input qq_in632;
input qq_in633;
input qq_in634;
input qq_in635;
input qq_in636;
input qq_in637;
input qq_in638;
input qq_in639;
input qq_in640;
input qq_in641;
input qq_in642;
input qq_in643;
input qq_in644;
input qq_in645;
input qq_in646;
input qq_in647;
input qq_in648;
input qq_in1166;
input qq_in1167;
input qq_in1168;
input qq_in1169;
input qq_in1170;
input qq_in1171;
input qq_in1172;
input qq_in1173;
input qq_in1174;
input qq_in1175;
input qq_in1176;
input qq_in1177;
input qq_in1178;
input qq_in1179;
input qq_in1180;
input qq_in1181;
input qq_in1182;
input qq_in1183;
input qq_in1184;
input qq_in1185;
input qq_in1186;
input qq_in1187;
input qq_in1188;
input qq_in1189;
input qq_in1190;
input qq_in1191;
input qq_in1192;
input qq_in1193;
input qq_in1194;
input qq_in1195;
input qq_in1196;
input qq_in1197;
input qq_in1198;
input qq_in1199;
input qq_in1200;
input qq_in1201;
input qq_in1202;
input qq_in1203;
input qq_in1204;
input qq_in1205;
input qq_in1206;
input qq_in1207;
input qq_in1208;
input qq_in1209;
input qq_in1210;
input qq_in1211;
input qq_in1212;
input qq_in1213;
input qq_in1214;
input qq_in1215;
input qq_in1216;
input qq_in1217;
input qq_in1218;
input qq_in1219;
input qq_in1220;
input qq_in1221;
input qq_in1222;
input qq_in1223;
input qq_in1224;
input qq_in1225;
input qq_in1226;
input qq_in1227;
input qq_in1228;
input qq_in1229;
input qq_in1230;
input qq_in1231;
input qq_in1232;
input qq_in1233;
input qq_in1234;
input qq_in1235;
input qq_in1236;
input qq_in1237;
input qq_in1238;
input qq_in1239;
input qq_in1240;
input qq_in1241;
input qq_in1242;
input qq_in1243;
input qq_in1244;
input qq_in1245;
input qq_in1246;
input qq_in1247;
input qq_in1248;
input qq_in1249;
input qq_in1250;
input qq_in1251;
input qq_in1252;
input qq_in1253;
input qq_in1254;
input qq_in1255;
input qq_in1256;
input qq_in1257;
input qq_in1258;
input qq_in1259;
input qq_in1260;
input qq_in1261;
input qq_in1262;
input qq_in1263;
input qq_in1264;
input qq_in1265;
input qq_in1266;
input qq_in1267;
input qq_in1268;
input qq_in1269;
input qq_in1270;
input qq_in1271;
input qq_in1272;
input qq_in1273;
input qq_in1274;
input qq_in1275;
input qq_in1276;
input qq_in1277;
input qq_in1278;
input qq_in1279;
input qq_in1280;
input qq_in1281;
input qq_in1282;
input qq_in1283;
input qq_in1284;
input qq_in1285;
input qq_in1286;
input qq_in1287;
input qq_in1288;
input qq_in1289;
input qq_in1290;
input qq_in1291;
input qq_in1292;
input qq_in1293;
input qq_in649;
input qq_in650;
input qq_in651;
input qq_in652;
input qq_in653;
input qq_in654;
input qq_in655;
input qq_in656;
input qq_in657;
input qq_in658;
input qq_in659;
input qq_in660;
input qq_in661;
input qq_in662;
input qq_in663;
input qq_in664;
input qq_in665;
input qq_in666;
input qq_in667;
input qq_in668;
input qq_in669;
input qq_in670;
input qq_in671;
input qq_in672;
input qq_in673;
input qq_in674;
input qq_in675;
input qq_in676;
input qq_in677;
input qq_in678;
input qq_in679;
input qq_in680;
input qq_in681;
input qq_in682;
input qq_in683;
input qq_in684;
input qq_in685;
input qq_in686;
input qq_in687;
input qq_in688;
input qq_in689;
input qq_in690;
input qq_in691;
input qq_in692;
input qq_in693;
input qq_in694;
input qq_in695;
input qq_in696;
input qq_in697;
input qq_in698;
input qq_in699;
input qq_in700;
input qq_in701;
input qq_in702;
input qq_in703;
input qq_in704;
input qq_in705;
input qq_in706;
input qq_in707;
input qq_in708;
input qq_in709;
input qq_in710;
input qq_in711;
input qq_in712;
input qq_in713;
input qq_in714;
input qq_in715;
input qq_in716;
input qq_in717;
input qq_in718;
input qq_in719;
input qq_in720;
input qq_in721;
input qq_in722;
input qq_in723;
input qq_in724;
input qq_in725;
input qq_in726;
input qq_in727;
input qq_in728;
input qq_in729;
input qq_in730;
input qq_in731;
input qq_in732;
input qq_in733;
input qq_in734;
input qq_in735;
input qq_in736;
input qq_in737;
input qq_in738;
input qq_in739;
input qq_in740;
input qq_in741;
input qq_in742;
input qq_in743;
input qq_in744;
input qq_in745;
input qq_in746;
input qq_in747;
input qq_in748;
input qq_in749;
input qq_in750;
input qq_in751;
input qq_in752;
input qq_in753;
input qq_in754;
input qq_in755;
input qq_in756;
input qq_in757;
input qq_in758;
input qq_in759;
input qq_in760;
input qq_in761;
input qq_in762;
input qq_in763;
input qq_in764;
input qq_in765;
input qq_in766;
input qq_in767;
input qq_in768;
input qq_in769;
input qq_in770;
input qq_in771;
input qq_in772;
input qq_in773;
input qq_in774;
input qq_in775;
input qq_in776;
input qq_in777;
input qq_in778;
input qq_in779;
input qq_in934;
input qq_in1294;
input qq_in1295;
input qq_in1296;
input qq_in1297;
input qq_in1298;
input qq_in1299;
input qq_in1300;
input qq_in1302;
input qq_in1303;
input qq_in1304;
input qq_in1305;
input qq_in781;
input qq_in782;
input qq_in783;
input qq_in784;
input qq_in785;
input qq_in786;
input qq_in787;
input qq_in788;
input qq_in789;
input qq_in780;
input qq_in791;
input qq_in792;
input qq_in793;
input qq_in794;
input qq_in795;
input qq_in796;
input qq_in797;
input qq_in798;
input qq_in799;
input qq_in800;
input qq_in801;
input qq_in802;
input qq_in803;
input qq_in804;
input qq_in805;
input qq_in806;
input qq_in807;
input qq_in808;
input qq_in809;
input qq_in810;
input qq_in811;
input qq_in812;
input qq_in813;
input qq_in814;
input qq_in815;
input qq_in816;
input qq_in817;
input qq_in818;
input qq_in819;
input qq_in820;
input qq_in821;
input qq_in822;
input qq_in823;
input qq_in824;
input qq_in825;
input qq_in826;
input qq_in827;
input qq_in828;
input qq_in829;
input qq_in830;
input qq_in831;
input qq_in832;
input qq_in833;
input qq_in834;
input qq_in835;
input qq_in836;
input qq_in837;
input qq_in838;
input qq_in839;
input qq_in840;
input qq_in841;
input qq_in842;
input qq_in843;
input qq_in844;
input qq_in845;
input qq_in846;
input qq_in847;
input qq_in848;
input qq_in849;
input qq_in850;
input qq_in851;
input qq_in852;
input qq_in853;
input qq_in854;
input qq_in855;
input qq_in856;
input qq_in857;
input qq_in858;
input qq_in859;
input qq_in860;
input qq_in861;
input qq_in862;
input qq_in863;
input qq_in864;
input qq_in865;
input qq_in866;
input qq_in867;
input qq_in868;
input qq_in869;
input qq_in870;
input qq_in871;
input qq_in872;
input qq_in873;
input qq_in874;
input qq_in875;
input qq_in876;
input qq_in877;
input qq_in878;
input qq_in879;
input qq_in880;
input qq_in881;
input qq_in882;
input qq_in883;
input qq_in884;
input qq_in885;
input qq_in886;
input qq_in887;
input qq_in888;
input qq_in889;
input qq_in890;
input qq_in891;
input qq_in892;
input qq_in893;
input qq_in894;
input qq_in895;
input qq_in896;
input qq_in897;
input qq_in898;
input qq_in899;
input qq_in900;
input qq_in901;
input qq_in902;
input qq_in903;
input qq_in904;
input qq_in905;
input qq_in906;
input qq_in907;
input qq_in908;
input qq_in909;
input qq_in910;
input qq_in911;
input qq_in912;
input qq_in913;
input qq_in914;
input qq_in915;
input qq_in916;
input qq_in917;
input qq_in918;
input qq_in919;
input qq_in920;
input qq_in921;
input qq_in922;
input qq_in923;
input qq_in924;
input qq_in925;
input qq_in926;
input qq_in927;
input qq_in928;
input qq_in929;
input qq_in930;
input qq_in931;
input qq_in932;
input qq_in933;
input qq_in790;
input qq_in935;
input qq_in936;
input qq_in937;
input qq_in938;
input qq_in939;
input qq_in940;
input qq_in941;
input qq_in942;
input qq_in943;
input qq_in944;
input qq_in945;
input qq_in946;
input qq_in947;
input qq_in948;
input qq_in949;
input qq_in950;
input qq_in951;
input qq_in952;
input qq_in953;
input qq_in954;
input qq_in955;
input qq_in956;
input qq_in957;
input qq_in958;
input qq_in959;
input qq_in960;
input qq_in961;
input qq_in962;
input qq_in963;
input qq_in964;
input qq_in965;
input qq_in966;
input qq_in967;
input qq_in968;
input qq_in969;
input qq_in970;
input qq_in971;
input qq_in972;
input qq_in973;
input qq_in974;
input qq_in975;
input qq_in976;
input qq_in977;
input qq_in978;
input qq_in979;
input qq_in980;
input qq_in981;
input qq_in982;
input qq_in983;
input qq_in984;
input qq_in985;
input qq_in986;
input qq_in987;
input qq_in988;
input qq_in989;
input qq_in990;
input qq_in991;
input qq_in992;
input qq_in993;
input qq_in994;
input qq_in995;
input qq_in996;
input qq_in997;
input qq_in998;
input qq_in999;
input qq_in1000;
input qq_in1001;
input qq_in1002;
input qq_in1003;
input qq_in1004;
input qq_in1005;
input qq_in1006;
input qq_in1007;
input qq_in1008;
input qq_in1009;
input qq_in1010;
input qq_in1011;
input qq_in1012;
input qq_in1013;
input qq_in1014;
input qq_in1015;
input qq_in1016;
input qq_in1017;
input qq_in1018;
input qq_in1019;
input qq_in1020;
input qq_in1021;
input qq_in1022;
input qq_in1023;
input qq_in1024;
input qq_in1025;
input qq_in1026;
input qq_in1027;
input qq_in1028;
input qq_in1029;
input qq_in1030;
input qq_in1031;
input qq_in1032;
input qq_in1033;
input qq_in1034;
input qq_in1035;
input qq_in1036;
input qq_in1037;
input qq_in1038;
input qq_in1039;
input qq_in1040;
input qq_in1041;
input qq_in1042;
input qq_in1043;
input qq_in1044;
input qq_in1045;
input qq_in1046;
input qq_in1047;
input qq_in1048;
input qq_in1049;
input qq_in1050;
input qq_in1051;
input qq_in1052;
input qq_in1053;
input qq_in1054;
input qq_in1055;
input qq_in1056;
input qq_in1057;
input qq_in1058;
input qq_in1059;
input qq_in1060;
input qq_in1061;
input qq_in1062;
input qq_in1063;
input qq_in1064;
input qq_in1065;
input qq_in1066;
input qq_in1067;
input qq_in1068;
input qq_in1069;
input qq_in1070;
input qq_in1071;
input qq_in1072;
input qq_in1073;
input qq_in1074;
input qq_in1075;
input qq_in1076;
input qq_in1077;
input qq_in1078;
input qq_in1079;
input qq_in1080;
input qq_in1081;
input qq_in1082;
input qq_in1083;
input qq_in1084;
input qq_in1085;
input qq_in1086;
input qq_in1087;
input qq_in1088;
input qq_in1089;
input qq_in1090;
input qq_in1091;
input qq_in1092;
input qq_in1093;
input qq_in1094;
input qq_in1095;
input qq_in1096;
input qq_in1097;
input qq_in1098;
input qq_in1099;
input qq_in1100;
input qq_in1101;
input qq_in1102;
input qq_in1103;
input qq_in1104;
input qq_in1105;
input qq_in1106;
input qq_in1107;
input qq_in1108;
input qq_in1109;
input qq_in1110;
input qq_in1111;
input qq_in1112;
input qq_in1113;
input qq_in1114;
input qq_in1115;
input qq_in1116;
input qq_in1117;
input qq_in1118;
input qq_in1119;
input qq_in1120;
input qq_in1121;
input qq_in1122;
input qq_in1123;
input qq_in1124;
input qq_in1125;
input qq_in1126;
input qq_in1127;
input qq_in1128;
input qq_in1129;
input qq_in1130;
input qq_in1131;
input qq_in1132;
input qq_in1133;
input qq_in1134;
input qq_in1135;
input qq_in1136;
input qq_in1137;
input qq_in1138;
input qq_in1139;
input qq_in1140;
input qq_in1141;
input qq_in1142;
input qq_in1143;
input qq_in1144;
input qq_in1145;
input qq_in1146;
input qq_in1147;
input qq_in1148;
input qq_in1149;
input qq_in1150;
input qq_in1151;
input qq_in1152;
input qq_in1153;
input qq_in1154;
input qq_in1155;
input qq_in1156;
input qq_in1157;
input qq_in1158;
input qq_in1159;
input qq_in1160;
input qq_in1161;
input qq_in1162;
input qq_in1163;
input qq_in1164;
input qq_in1165;
input qnn_in_1301;
input qnn_in_1303;
input qnn_in_760;
input qnn_in_761;
input qnn_in_762;
input qnn_in_763;
input qnn_in_764;
input qnn_in_766;
input qnn_in_767;
input qnn_in_768;
input qnn_in_780;
input qnn_in_777;
input qnn_in_778;
input qnn_in_779;
input qnn_in_649;
input qnn_in_650;
input qnn_in_651;
input qnn_in_654;
input qnn_in_1;
input qnn_in_2;
input qnn_in_3;
input qnn_in_4;
input qnn_in_5;
input qnn_in_6;
input qnn_in_7;
input qnn_in_8;
input qnn_in_9;
input qnn_in_10;
input qnn_in_11;
input qnn_in_12;
input qnn_in_13;
input qnn_in_14;
input qnn_in_15;
input qnn_in_16;
input qnn_in_17;
input qnn_in_18;
input qnn_in_19;
input qnn_in_20;
input qnn_in_21;
input qnn_in_22;
input qnn_in_23;
input qnn_in_24;
input qnn_in_25;
input qnn_in_26;
input qnn_in_27;
input qnn_in_28;
input qnn_in_29;
input qnn_in_30;
input qnn_in_31;
input qnn_in_32;
input qnn_in_33;
input qnn_in_34;
input qnn_in_35;
input qnn_in_36;
input qnn_in_37;
input qnn_in_38;
input qnn_in_39;
input qnn_in_40;
input qnn_in_41;
input qnn_in_42;
input qnn_in_43;
input qnn_in_44;
input qnn_in_45;
input qnn_in_46;
input qnn_in_47;
input qnn_in_48;
input qnn_in_49;
input qnn_in_50;
input qnn_in_51;
input qnn_in_52;
input qnn_in_53;
input qnn_in_54;
input qnn_in_55;
input qnn_in_56;
input qnn_in_57;
input qnn_in_58;
input qnn_in_59;
input qnn_in_60;
input qnn_in_61;
input qnn_in_62;
input qnn_in_63;
input qnn_in_64;
input qnn_in_65;
input qnn_in_66;
input qnn_in_67;
input qnn_in_68;
input qnn_in_69;
input qnn_in_70;
input qnn_in_71;
input qnn_in_72;
input qnn_in_73;
input qnn_in_74;
input qnn_in_75;
input qnn_in_76;
input qnn_in_77;
input qnn_in_78;
input qnn_in_79;
input qnn_in_80;
input qnn_in_81;
input qnn_in_82;
input qnn_in_83;
input qnn_in_84;
input qnn_in_85;
input qnn_in_86;
input qnn_in_87;
input qnn_in_88;
input qnn_in_89;
input qnn_in_90;
input qnn_in_91;
input qnn_in_92;
input qnn_in_93;
input qnn_in_94;
input qnn_in_95;
input qnn_in_96;
input qnn_in_97;
input qnn_in_98;
input qnn_in_99;
input qnn_in_100;
input qnn_in_101;
input qnn_in_102;
input qnn_in_103;
input qnn_in_104;
input qnn_in_105;
input qnn_in_106;
input qnn_in_107;
input qnn_in_108;
input qnn_in_109;
input qnn_in_110;
input qnn_in_111;
input qnn_in_112;
input qnn_in_113;
input qnn_in_114;
input qnn_in_115;
input qnn_in_116;
input qnn_in_117;
input qnn_in_118;
input qnn_in_119;
input qnn_in_120;
input qnn_in_121;
input qnn_in_122;
input qnn_in_123;
input qnn_in_124;
input qnn_in_125;
input qnn_in_126;
input qnn_in_127;
input qnn_in_128;
input qnn_in_667;
input qnn_in_668;
input qnn_in_669;
input qnn_in_670;
output d_out_398;
output d_out_397;
output d_out_396;
output d_out_395;
output d_out_191;
output d_out_190;
output d_out_189;
output d_out_188;
output d_out_187;
output d_out_186;
output d_out_185;
output d_out_184;
output d_out_183;
output d_out_182;
output d_out_181;
output d_out_180;
output d_out_179;
output d_out_178;
output d_out_177;
output d_out_176;
output d_out_175;
output d_out_174;
output d_out_173;
output d_out_172;
output d_out_171;
output d_out_170;
output d_out_169;
output d_out_168;
output d_out_167;
output d_out_166;
output d_out_165;
output d_out_164;
output d_out_163;
output d_out_162;
output d_out_161;
output d_out_160;
output d_out_159;
output d_out_158;
output d_out_157;
output d_out_156;
output d_out_155;
output d_out_154;
output d_out_153;
output d_out_152;
output d_out_151;
output d_out_150;
output d_out_149;
output d_out_148;
output d_out_147;
output d_out_146;
output d_out_145;
output d_out_144;
output d_out_143;
output d_out_142;
output d_out_141;
output d_out_140;
output d_out_139;
output d_out_138;
output d_out_137;
output d_out_136;
output d_out_135;
output d_out_134;
output d_out_133;
output d_out_132;
output d_out_131;
output d_out_130;
output d_out_129;
output d_out_128;
output d_out_127;
output d_out_126;
output d_out_125;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_121;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_116;
output d_out_115;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_111;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_83;
output d_out_82;
output d_out_81;
output d_out_80;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_76;
output d_out_75;
output d_out_74;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_64;
output d_out_63;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_50;
output d_out_49;
output d_out_48;
output d_out_47;
output d_out_46;
output d_out_45;
output d_out_44;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_30;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_5;
output d_out_4;
output d_out_3;
output d_out_2;
output d_out_1;
output [127:0] Out_data;
output [3:0] Out_data_size;
output dii_data_not_ready, Out_vld, Out_last_word, Tag_vld;
output ddout__1;
output ddout__2;
output ddout__3;
output ddout__4;
output ddout__5;
output ddout__6;
output ddout__7;
output ddout__8;
output ddout__9;
output ddout__10;
output ddout__11;
output ddout__12;
output ddout__13;
output ddout__14;
output ddout__15;
output ddout__16;
output ddout__17;
output ddout__18;
output ddout__19;
output ddout__20;
output ddout__21;
output ddout__22;
output ddout__23;
output ddout__24;
output ddout__25;
output ddout__26;
output ddout__27;
output ddout__28;
output ddout__29;
output ddout__30;
output ddout__31;
output ddout__32;
output ddout__33;
output ddout__34;
output ddout__35;
output ddout__36;
output ddout__37;
output ddout__38;
output ddout__39;
output ddout__40;
output ddout__41;
output ddout__42;
output ddout__43;
output ddout__44;
output ddout__45;
output ddout__46;
output ddout__47;
output ddout__48;
output ddout__49;
output ddout__50;
output ddout__51;
output ddout__52;
output ddout__53;
output ddout__54;
output ddout__55;
output ddout__56;
output ddout__57;
output ddout__58;
output ddout__59;
output ddout__60;
output ddout__61;
output ddout__62;
output ddout__63;
output ddout__64;
output ddout__65;
output ddout__66;
output ddout__67;
output ddout__68;
output ddout__69;
output ddout__70;
output ddout__71;
output ddout__72;
output ddout__73;
output ddout__74;
output ddout__75;
output ddout__76;
output ddout__77;
output ddout__78;
output ddout__79;
output ddout__80;
output ddout__81;
output ddout__82;
output ddout__83;
output ddout__84;
output ddout__85;
output ddout__86;
output ddout__87;
output ddout__88;
output ddout__89;
output ddout__90;
output ddout__91;
output ddout__92;
output ddout__93;
output ddout__94;
output ddout__95;
output ddout__96;
output ddout__97;
output ddout__98;
output ddout__99;
output ddout__100;
output ddout__101;
output ddout__102;
output ddout__103;
output ddout__104;
output ddout__105;
output ddout__106;
output ddout__107;
output ddout__108;
output ddout__109;
output ddout__110;
output ddout__111;
output ddout__112;
output ddout__113;
output ddout__114;
output ddout__115;
output ddout__116;
output ddout__117;
output ddout__118;
output ddout__119;
output ddout__120;
output ddout__121;
output ddout__122;
output ddout__123;
output ddout__124;
output ddout__125;
output ddout__126;
output ddout__127;
output ddout__128;
output ddout__129;
output ddout__130;
output ddout__131;
output ddout__132;
output ddout__133;
output ddout__134;
output ddout__135;
output ddout__136;
output ddout__137;
output ddout__138;
output ddout__139;
output ddout__140;
output ddout__141;
output ddout__142;
output ddout__143;
output ddout__144;
output ddout__145;
output ddout__146;
output ddout__147;
output ddout__148;
output ddout__149;
output ddout__150;
output ddout__151;
output ddout__152;
output ddout__153;
output ddout__154;
output ddout__155;
output ddout__156;
output ddout__157;
output ddout__158;
output ddout__159;
output ddout__160;
output ddout__161;
output ddout__162;
output ddout__163;
output ddout__164;
output ddout__165;
output ddout__166;
output ddout__167;
output ddout__168;
output ddout__169;
output ddout__170;
output ddout__171;
output ddout__172;
output ddout__173;
output ddout__174;
output ddout__175;
output ddout__176;
output ddout__177;
output ddout__178;
output ddout__179;
output ddout__180;
output ddout__181;
output ddout__182;
output ddout__183;
output ddout__184;
output ddout__185;
output ddout__186;
output ddout__187;
output ddout__188;
output ddout__189;
output ddout__190;
output ddout__191;
output ddout__192;
output ddout__193;
output ddout__194;
output ddout__195;
output ddout__196;
output ddout__197;
output ddout__198;
output ddout__199;
output ddout__200;
output ddout__201;
output ddout__202;
output ddout__203;
output ddout__204;
output ddout__205;
output ddout__206;
output ddout__207;
output ddout__208;
output ddout__209;
output ddout__210;
output ddout__211;
output ddout__212;
output ddout__213;
output ddout__214;
output ddout__215;
output ddout__216;
output ddout__217;
output ddout__218;
output ddout__219;
output ddout__220;
output ddout__221;
output ddout__222;
output ddout__223;
output ddout__224;
output ddout__225;
output ddout__226;
output ddout__227;
output ddout__228;
output ddout__229;
output ddout__230;
output ddout__231;
output ddout__232;
output ddout__233;
output ddout__234;
output ddout__235;
output ddout__236;
output ddout__237;
output ddout__238;
output ddout__239;
output ddout__240;
output ddout__241;
output ddout__242;
output ddout__243;
output ddout__244;
output ddout__245;
output ddout__246;
output ddout__247;
output ddout__248;
output ddout__249;
output ddout__250;
output ddout__251;
output ddout__252;
output ddout__253;
output ddout__254;
output ddout__255;
output ddout__256;
output ddout__257;
output ddout__258;
output ddout__259;
output ddout__260;
output ddout__261;
output ddout__262;
output ddout__263;
output ddout__264;
output ddout__265;
output ddout__266;
output ddout__267;
output ddout__268;
output ddout__269;
output ddout__270;
output ddout__271;
output ddout__272;
output ddout__273;
output ddout__274;
output ddout__275;
output ddout__276;
output ddout__277;
output ddout__278;
output ddout__279;
output ddout__280;
output ddout__281;
output ddout__282;
output ddout__283;
output ddout__284;
output ddout__285;
output ddout__286;
output ddout__287;
output ddout__288;
output ddout__289;
output ddout__290;
output ddout__291;
output ddout__292;
output ddout__293;
output ddout__294;
output ddout__295;
output ddout__296;
output ddout__297;
output ddout__298;
output ddout__299;
output ddout__300;
output ddout__301;
output ddout__302;
output ddout__303;
output ddout__304;
output ddout__305;
output ddout__306;
output ddout__307;
output ddout__308;
output ddout__309;
output ddout__310;
output ddout__311;
output ddout__312;
output ddout__313;
output ddout__314;
output ddout__315;
output ddout__316;
output ddout__317;
output ddout__318;
output ddout__319;
output ddout__320;
output ddout__321;
output ddout__322;
output ddout__323;
output ddout__324;
output ddout__325;
output ddout__326;
output ddout__327;
output ddout__328;
output ddout__329;
output ddout__330;
output ddout__331;
output ddout__332;
output ddout__333;
output ddout__334;
output ddout__335;
output ddout__336;
output ddout__337;
output ddout__338;
output ddout__339;
output ddout__340;
output ddout__341;
output ddout__342;
output ddout__343;
output ddout__344;
output ddout__345;
output ddout__346;
output ddout__347;
output ddout__348;
output ddout__349;
output ddout__350;
output ddout__351;
output ddout__352;
output ddout__353;
output ddout__354;
output ddout__355;
output ddout__356;
output ddout__357;
output ddout__358;
output ddout__359;
output ddout__360;
output ddout__361;
output ddout__362;
output ddout__363;
output ddout__364;
output ddout__365;
output ddout__366;
output ddout__367;
output ddout__368;
output ddout__369;
output ddout__370;
output ddout__371;
output ddout__372;
output ddout__373;
output ddout__374;
output ddout__375;
output ddout__376;
output ddout__377;
output ddout__378;
output ddout__379;
output ddout__380;
output ddout__381;
output ddout__382;
output ddout__383;
output ddout__384;
output ddout__385;
output ddout__386;
output ddout__387;
output ddout__388;
output ddout__389;
output ddout__390;
output ddout__391;
output ddout__392;
output ddout__393;
output ddout__394;
output ddout__395;
output ddout__396;
output ddout__397;
output ddout__398;
output ddout__399;
output ddout__400;
output ddout__401;
output ddout__402;
output ddout__403;
output ddout__404;
output ddout__405;
output ddout__406;
output ddout__407;
output ddout__408;
output ddout__409;
output ddout__410;
output ddout__411;
output ddout__412;
output ddout__413;
output ddout__414;
output ddout__415;
output ddout__416;
output ddout__417;
output ddout__418;
output ddout__419;
output ddout__420;
output ddout__421;
output ddout__422;
output ddout__423;
output ddout__424;
output ddout__425;
output ddout__426;
output ddout__427;
output ddout__428;
output ddout__429;
output ddout__430;
output ddout__431;
output ddout__432;
output ddout__433;
output ddout__434;
output ddout__435;
output ddout__436;
output ddout__437;
output ddout__438;
output ddout__439;
output ddout__440;
output ddout__441;
output ddout__442;
output ddout__443;
output ddout__444;
output ddout__445;
output ddout__446;
output ddout__447;
output ddout__448;
output ddout__449;
output ddout__450;
output ddout__451;
output ddout__452;
output ddout__453;
output ddout__454;
output ddout__455;
output ddout__456;
output ddout__457;
output ddout__458;
output ddout__459;
output ddout__460;
output ddout__461;
output ddout__462;
output ddout__463;
output ddout__464;
output ddout__465;
output ddout__466;
output ddout__467;
output ddout__468;
output ddout__469;
output ddout__470;
output ddout__471;
output ddout__472;
output ddout__473;
output ddout__474;
output ddout__475;
output ddout__476;
output ddout__477;
output ddout__478;
output ddout__479;
output ddout__480;
output ddout__481;
output ddout__482;
output ddout__483;
output ddout__484;
output ddout__485;
output ddout__486;
output ddout__487;
output ddout__488;
output ddout__489;
output ddout__490;
output ddout__491;
output ddout__492;
output ddout__493;
output ddout__494;
output ddout__495;
output ddout__496;
output ddout__497;
output ddout__498;
output ddout__499;
output ddout__500;
output ddout__501;
output ddout__502;
output ddout__503;
output ddout__504;
output ddout__505;
output ddout__506;
output ddout__507;
output ddout__508;
output ddout__509;
output ddout__510;
output ddout__511;
output ddout__512;
output ddout__513;
output ddout__514;
output ddout__515;
output ddout__516;
output ddout__517;
output ddout__518;
output ddout__519;
output ddout__520;
output ddout__521;
output ddout__522;
output ddout__523;
output ddout__524;
output ddout__525;
output ddout__526;
output ddout__527;
output ddout__528;
output ddout__529;
output ddout__530;
output ddout__531;
output ddout__532;
output ddout__533;
output ddout__534;
output ddout__535;
output ddout__536;
output ddout__537;
output ddout__538;
output ddout__539;
output ddout__540;
output ddout__541;
output ddout__542;
output ddout__543;
output ddout__544;
output ddout__545;
output ddout__546;
output ddout__547;
output ddout__548;
output ddout__549;
output ddout__550;
output ddout__551;
output ddout__552;
output ddout__553;
output ddout__554;
output ddout__555;
output ddout__556;
output ddout__557;
output ddout__558;
output ddout__559;
output ddout__560;
output ddout__561;
output ddout__562;
output ddout__563;
output ddout__564;
output ddout__565;
output ddout__566;
output ddout__567;
output ddout__568;
output ddout__569;
output ddout__570;
output ddout__571;
output ddout__572;
output ddout__573;
output ddout__574;
output ddout__575;
output ddout__576;
output ddout__577;
output ddout__578;
output ddout__579;
output ddout__580;
output ddout__581;
output ddout__582;
output ddout__583;
output ddout__584;
output ddout__585;
output ddout__586;
output ddout__587;
output ddout__588;
output ddout__589;
output ddout__590;
output ddout__591;
output ddout__592;
output ddout__593;
output ddout__594;
output ddout__595;
output ddout__596;
output ddout__597;
output ddout__598;
output ddout__599;
output ddout__600;
output ddout__601;
output ddout__602;
output ddout__603;
output ddout__604;
output ddout__605;
output ddout__606;
output ddout__607;
output ddout__608;
output ddout__609;
output ddout__610;
output ddout__611;
output ddout__612;
output ddout__613;
output ddout__614;
output ddout__615;
output ddout__616;
output ddout__617;
output ddout__618;
output ddout__619;
output ddout__620;
output ddout__621;
output ddout__622;
output ddout__623;
output ddout__624;
output ddout__625;
output ddout__626;
output ddout__627;
output ddout__628;
output ddout__629;
output ddout__630;
output ddout__631;
output ddout__632;
output ddout__633;
output ddout__634;
output ddout__635;
output ddout__636;
output ddout__637;
output ddout__638;
output ddout__639;
output ddout__640;
output ddout__641;
output ddout__642;
output ddout__643;
output ddout__644;
output ddout__645;
output ddout__646;
output ddout__647;
output ddout__648;
output ddout__1166;
output ddout__1167;
output ddout__1168;
output ddout__1169;
output ddout__1170;
output ddout__1171;
output ddout__1172;
output ddout__1173;
output ddout__1174;
output ddout__1175;
output ddout__1176;
output ddout__1177;
output ddout__1178;
output ddout__1179;
output ddout__1180;
output ddout__1181;
output ddout__1182;
output ddout__1183;
output ddout__1184;
output ddout__1185;
output ddout__1186;
output ddout__1187;
output ddout__1188;
output ddout__1189;
output ddout__1190;
output ddout__1191;
output ddout__1192;
output ddout__1193;
output ddout__1194;
output ddout__1195;
output ddout__1196;
output ddout__1197;
output ddout__1198;
output ddout__1199;
output ddout__1200;
output ddout__1201;
output ddout__1202;
output ddout__1203;
output ddout__1204;
output ddout__1205;
output ddout__1206;
output ddout__1207;
output ddout__1208;
output ddout__1209;
output ddout__1210;
output ddout__1211;
output ddout__1212;
output ddout__1213;
output ddout__1214;
output ddout__1215;
output ddout__1216;
output ddout__1217;
output ddout__1218;
output ddout__1219;
output ddout__1220;
output ddout__1221;
output ddout__1222;
output ddout__1223;
output ddout__1224;
output ddout__1225;
output ddout__1226;
output ddout__1227;
output ddout__1228;
output ddout__1229;
output ddout__1230;
output ddout__1231;
output ddout__1232;
output ddout__1233;
output ddout__1234;
output ddout__1235;
output ddout__1236;
output ddout__1237;
output ddout__1238;
output ddout__1239;
output ddout__1240;
output ddout__1241;
output ddout__1242;
output ddout__1243;
output ddout__1244;
output ddout__1245;
output ddout__1246;
output ddout__1247;
output ddout__1248;
output ddout__1249;
output ddout__1250;
output ddout__1251;
output ddout__1252;
output ddout__1253;
output ddout__1254;
output ddout__1255;
output ddout__1256;
output ddout__1257;
output ddout__1258;
output ddout__1259;
output ddout__1260;
output ddout__1261;
output ddout__1262;
output ddout__1263;
output ddout__1264;
output ddout__1265;
output ddout__1266;
output ddout__1267;
output ddout__1268;
output ddout__1269;
output ddout__1270;
output ddout__1271;
output ddout__1272;
output ddout__1273;
output ddout__1274;
output ddout__1275;
output ddout__1276;
output ddout__1277;
output ddout__1278;
output ddout__1279;
output ddout__1280;
output ddout__1281;
output ddout__1282;
output ddout__1283;
output ddout__1284;
output ddout__1285;
output ddout__1286;
output ddout__1287;
output ddout__1288;
output ddout__1289;
output ddout__1290;
output ddout__1291;
output ddout__1292;
output ddout__1293;
output ddout__649;
output ddout__650;
output ddout__651;
output ddout__652;
output ddout__653;
output ddout__654;
output ddout__655;
output ddout__656;
output ddout__657;
output ddout__658;
output ddout__659;
output ddout__660;
output ddout__661;
output ddout__662;
output ddout__663;
output ddout__664;
output ddout__665;
output ddout__666;
output ddout__667;
output ddout__668;
output ddout__669;
output ddout__670;
output ddout__671;
output ddout__672;
output ddout__673;
output ddout__674;
output ddout__675;
output ddout__676;
output ddout__677;
output ddout__678;
output ddout__679;
output ddout__680;
output ddout__681;
output ddout__682;
output ddout__683;
output ddout__684;
output ddout__685;
output ddout__686;
output ddout__687;
output ddout__688;
output ddout__689;
output ddout__690;
output ddout__691;
output ddout__692;
output ddout__693;
output ddout__694;
output ddout__695;
output ddout__696;
output ddout__697;
output ddout__698;
output ddout__699;
output ddout__700;
output ddout__701;
output ddout__702;
output ddout__703;
output ddout__704;
output ddout__705;
output ddout__706;
output ddout__707;
output ddout__708;
output ddout__709;
output ddout__710;
output ddout__711;
output ddout__712;
output ddout__713;
output ddout__714;
output ddout__715;
output ddout__716;
output ddout__717;
output ddout__718;
output ddout__719;
output ddout__720;
output ddout__721;
output ddout__722;
output ddout__723;
output ddout__724;
output ddout__725;
output ddout__726;
output ddout__727;
output ddout__728;
output ddout__729;
output ddout__730;
output ddout__731;
output ddout__732;
output ddout__733;
output ddout__734;
output ddout__735;
output ddout__736;
output ddout__737;
output ddout__738;
output ddout__739;
output ddout__740;
output ddout__741;
output ddout__742;
output ddout__743;
output ddout__744;
output ddout__745;
output ddout__746;
output ddout__747;
output ddout__748;
output ddout__749;
output ddout__750;
output ddout__751;
output ddout__752;
output ddout__753;
output ddout__754;
output ddout__755;
output ddout__756;
output ddout__757;
output ddout__758;
output ddout__759;
output ddout__760;
output ddout__761;
output ddout__762;
output ddout__763;
output ddout__764;
output ddout__765;
output ddout__766;
output ddout__767;
output ddout__768;
output ddout__769;
output ddout__770;
output ddout__771;
output ddout__772;
output ddout__773;
output ddout__774;
output ddout__775;
output ddout__776;
output ddout__777;
output ddout__778;
output ddout__779;
output ddout__934;
output ddout__1294;
output ddout__1295;
output ddout__1296;
output ddout__1297;
output ddout__1298;
output ddout__1299;
output ddout__1300;
output ddout__1301;
output ddout__1302;
output ddout__1303;
output ddout__1304;
output ddout__1305;
output ddout__781;
output ddout__782;
output ddout__783;
output ddout__784;
output ddout__785;
output ddout__786;
output ddout__787;
output ddout__788;
output ddout__789;
output ddout__780;
output ddout__791;
output ddout__792;
output ddout__793;
output ddout__794;
output ddout__795;
output ddout__796;
output ddout__797;
output ddout__798;
output ddout__799;
output ddout__800;
output ddout__801;
output ddout__802;
output ddout__803;
output ddout__804;
output ddout__805;
output ddout__806;
output ddout__807;
output ddout__808;
output ddout__809;
output ddout__810;
output ddout__811;
output ddout__812;
output ddout__813;
output ddout__814;
output ddout__815;
output ddout__816;
output ddout__817;
output ddout__818;
output ddout__819;
output ddout__820;
output ddout__821;
output ddout__822;
output ddout__823;
output ddout__824;
output ddout__825;
output ddout__826;
output ddout__827;
output ddout__828;
output ddout__829;
output ddout__830;
output ddout__831;
output ddout__832;
output ddout__833;
output ddout__834;
output ddout__835;
output ddout__836;
output ddout__837;
output ddout__838;
output ddout__839;
output ddout__840;
output ddout__841;
output ddout__842;
output ddout__843;
output ddout__844;
output ddout__845;
output ddout__846;
output ddout__847;
output ddout__848;
output ddout__849;
output ddout__850;
output ddout__851;
output ddout__852;
output ddout__853;
output ddout__854;
output ddout__855;
output ddout__856;
output ddout__857;
output ddout__858;
output ddout__859;
output ddout__860;
output ddout__861;
output ddout__862;
output ddout__863;
output ddout__864;
output ddout__865;
output ddout__866;
output ddout__867;
output ddout__868;
output ddout__869;
output ddout__870;
output ddout__871;
output ddout__872;
output ddout__873;
output ddout__874;
output ddout__875;
output ddout__876;
output ddout__877;
output ddout__878;
output ddout__879;
output ddout__880;
output ddout__881;
output ddout__882;
output ddout__883;
output ddout__884;
output ddout__885;
output ddout__886;
output ddout__887;
output ddout__888;
output ddout__889;
output ddout__890;
output ddout__891;
output ddout__892;
output ddout__893;
output ddout__894;
output ddout__895;
output ddout__896;
output ddout__897;
output ddout__898;
output ddout__899;
output ddout__900;
output ddout__901;
output ddout__902;
output ddout__903;
output ddout__904;
output ddout__905;
output ddout__906;
output ddout__907;
output ddout__908;
output ddout__909;
output ddout__910;
output ddout__911;
output ddout__912;
output ddout__913;
output ddout__914;
output ddout__915;
output ddout__916;
output ddout__917;
output ddout__918;
output ddout__919;
output ddout__920;
output ddout__921;
output ddout__922;
output ddout__923;
output ddout__924;
output ddout__925;
output ddout__926;
output ddout__927;
output ddout__928;
output ddout__929;
output ddout__930;
output ddout__931;
output ddout__932;
output ddout__933;
output ddout__790;
output ddout__935;
output ddout__936;
output ddout__937;
output ddout__938;
output ddout__939;
output ddout__940;
output ddout__941;
output ddout__942;
output ddout__943;
output ddout__944;
output ddout__945;
output ddout__946;
output ddout__947;
output ddout__948;
output ddout__949;
output ddout__950;
output ddout__951;
output ddout__952;
output ddout__953;
output ddout__954;
output ddout__955;
output ddout__956;
output ddout__957;
output ddout__958;
output ddout__959;
output ddout__960;
output ddout__961;
output ddout__962;
output ddout__963;
output ddout__964;
output ddout__965;
output ddout__966;
output ddout__967;
output ddout__968;
output ddout__969;
output ddout__970;
output ddout__971;
output ddout__972;
output ddout__973;
output ddout__974;
output ddout__975;
output ddout__976;
output ddout__977;
output ddout__978;
output ddout__979;
output ddout__980;
output ddout__981;
output ddout__982;
output ddout__983;
output ddout__984;
output ddout__985;
output ddout__986;
output ddout__987;
output ddout__988;
output ddout__989;
output ddout__990;
output ddout__991;
output ddout__992;
output ddout__993;
output ddout__994;
output ddout__995;
output ddout__996;
output ddout__997;
output ddout__998;
output ddout__999;
output ddout__1000;
output ddout__1001;
output ddout__1002;
output ddout__1003;
output ddout__1004;
output ddout__1005;
output ddout__1006;
output ddout__1007;
output ddout__1008;
output ddout__1009;
output ddout__1010;
output ddout__1011;
output ddout__1012;
output ddout__1013;
output ddout__1014;
output ddout__1015;
output ddout__1016;
output ddout__1017;
output ddout__1018;
output ddout__1019;
output ddout__1020;
output ddout__1021;
output ddout__1022;
output ddout__1023;
output ddout__1024;
output ddout__1025;
output ddout__1026;
output ddout__1027;
output ddout__1028;
output ddout__1029;
output ddout__1030;
output ddout__1031;
output ddout__1032;
output ddout__1033;
output ddout__1034;
output ddout__1035;
output ddout__1036;
output ddout__1037;
output ddout__1038;
output ddout__1039;
output ddout__1040;
output ddout__1041;
output ddout__1042;
output ddout__1043;
output ddout__1044;
output ddout__1045;
output ddout__1046;
output ddout__1047;
output ddout__1048;
output ddout__1049;
output ddout__1050;
output ddout__1051;
output ddout__1052;
output ddout__1053;
output ddout__1054;
output ddout__1055;
output ddout__1056;
output ddout__1057;
output ddout__1058;
output ddout__1059;
output ddout__1060;
output ddout__1061;
output ddout__1062;
output ddout__1063;
output ddout__1064;
output ddout__1065;
output ddout__1066;
output ddout__1067;
output ddout__1068;
output ddout__1069;
output ddout__1070;
output ddout__1071;
output ddout__1072;
output ddout__1073;
output ddout__1074;
output ddout__1075;
output ddout__1076;
output ddout__1077;
output ddout__1078;
output ddout__1079;
output ddout__1080;
output ddout__1081;
output ddout__1082;
output ddout__1083;
output ddout__1084;
output ddout__1085;
output ddout__1086;
output ddout__1087;
output ddout__1088;
output ddout__1089;
output ddout__1090;
output ddout__1091;
output ddout__1092;
output ddout__1093;
output ddout__1094;
output ddout__1095;
output ddout__1096;
output ddout__1097;
output ddout__1098;
output ddout__1099;
output ddout__1100;
output ddout__1101;
output ddout__1102;
output ddout__1103;
output ddout__1104;
output ddout__1105;
output ddout__1106;
output ddout__1107;
output ddout__1108;
output ddout__1109;
output ddout__1110;
output ddout__1111;
output ddout__1112;
output ddout__1113;
output ddout__1114;
output ddout__1115;
output ddout__1116;
output ddout__1117;
output ddout__1118;
output ddout__1119;
output ddout__1120;
output ddout__1121;
output ddout__1122;
output ddout__1123;
output ddout__1124;
output ddout__1125;
output ddout__1126;
output ddout__1127;
output ddout__1128;
output ddout__1129;
output ddout__1130;
output ddout__1131;
output ddout__1132;
output ddout__1133;
output ddout__1134;
output ddout__1135;
output ddout__1136;
output ddout__1137;
output ddout__1138;
output ddout__1139;
output ddout__1140;
output ddout__1141;
output ddout__1142;
output ddout__1143;
output ddout__1144;
output ddout__1145;
output ddout__1146;
output ddout__1147;
output ddout__1148;
output ddout__1149;
output ddout__1150;
output ddout__1151;
output ddout__1152;
output ddout__1153;
output ddout__1154;
output ddout__1155;
output ddout__1156;
output ddout__1157;
output ddout__1158;
output ddout__1159;
output ddout__1160;
output ddout__1161;
output ddout__1162;
output ddout__1163;
output ddout__1164;
output ddout__1165;
output d_out_394;
output d_out_393;
output d_out_392;
output d_out_391;
output d_out_390;
output d_out_389;
output d_out_388;
output d_out_387;
output d_out_386;
output d_out_385;
output d_out_384;
output d_out_383;
output d_out_382;
output d_out_381;
output d_out_380;
output d_out_379;
output d_out_378;
output d_out_377;
output d_out_376;
output d_out_375;
output d_out_374;
output d_out_373;
output d_out_372;
output d_out_371;
output d_out_370;
output d_out_369;
output d_out_368;
output d_out_367;
output d_out_366;
output d_out_365;
output d_out_364;
output d_out_363;
output d_out_362;
output d_out_361;
output d_out_360;
output d_out_359;
output d_out_358;
output d_out_357;
output d_out_356;
output d_out_355;
output d_out_354;
output d_out_353;
output d_out_352;
output d_out_351;
output d_out_350;
output d_out_349;
output d_out_348;
output d_out_347;
output d_out_346;
output d_out_345;
output d_out_344;
output d_out_343;
output d_out_342;
output d_out_341;
output d_out_340;
output d_out_339;
output d_out_338;
output d_out_337;
output d_out_336;
output d_out_335;
output d_out_334;
output d_out_333;
output d_out_332;
output d_out_331;
output d_out_330;
output d_out_329;
output d_out_328;
output d_out_327;
output d_out_326;
output d_out_325;
output d_out_324;
output d_out_323;
output d_out_322;
output d_out_321;
output d_out_320;
output d_out_319;
output d_out_318;
output d_out_317;
output d_out_316;
output d_out_315;
output d_out_314;
output d_out_313;
output d_out_312;
output d_out_311;
output d_out_310;
output d_out_309;
output d_out_308;
output d_out_307;
output d_out_306;
output d_out_305;
output d_out_304;
output d_out_303;
output d_out_302;
output d_out_301;
output d_out_300;
output d_out_299;
output d_out_298;
output d_out_297;
output d_out_296;
output d_out_295;
output d_out_294;
output d_out_293;
output d_out_292;
output d_out_291;
output d_out_290;
output d_out_289;
output d_out_288;
output d_out_287;
output d_out_286;
output d_out_285;
output d_out_284;
output d_out_283;
output d_out_282;
output d_out_281;
output d_out_280;
output d_out_279;
output d_out_278;
output d_out_277;
output d_out_276;
output d_out_275;
output d_out_274;
output d_out_273;
output d_out_272;
output d_out_271;
output d_out_270;
output d_out_269;
output d_out_268;
output d_out_267;
output d_out_266;
output d_out_265;
output d_out_264;
output d_out_263;
output d_out_262;
output d_out_261;
output d_out_260;
output d_out_259;
output d_out_258;
output d_out_257;
output d_out_256;
output d_out_255;
output d_out_254;
output d_out_253;
output d_out_252;
output d_out_251;
output d_out_250;
output d_out_249;
output d_out_248;
output d_out_247;
output d_out_246;
output d_out_245;
output d_out_244;
output d_out_243;
output d_out_242;
output d_out_241;
output d_out_240;
output d_out_239;
output d_out_238;
output d_out_237;
output d_out_236;
output d_out_235;
output d_out_234;
output d_out_233;
output d_out_232;
output d_out_231;
output d_out_230;
output d_out_229;
output d_out_228;
output d_out_227;
output d_out_226;
output d_out_225;
output d_out_224;
output d_out_223;
output d_out_222;
output d_out_221;
output d_out_220;
output d_out_219;
output d_out_218;
output d_out_217;
output d_out_216;
output d_out_215;
output d_out_214;
output d_out_213;
output d_out_212;
output d_out_211;
output d_out_210;
output d_out_209;
output d_out_208;
output d_out_207;
output d_out_206;
output d_out_205;
output d_out_204;
output d_out_203;
output d_out_202;
output d_out_201;
output d_out_200;
output d_out_199;
output d_out_198;
output d_out_197;
output d_out_196;
output d_out_195;
output d_out_194;
output d_out_193;
output d_out_192;
wire aes_done, aes_kld, N2027, N2028, N2029, N2030, N2031, N2032, N2033, N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2075, 
  N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083, N2084, N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114, N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2123, N2124, N2125, 
  N2126, N2127, N2128, N2129, N2130, N2131, N2132, N2133, N2134, N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153, N2154, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369, 
  N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407, N2408, N2409, N2410, N2411, N2412, N2479, N2480, N2481, N2482, N2483, N2484, N2485, 
  N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, 
  N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, 
  N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, 
  N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, 
  N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, 
  N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055, N3056, N3057, 
  N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, 
  N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135, N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, N3156, N3157, 
  N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3198, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5342, 
  n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, 
  n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
  n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
  n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, 
  n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
  n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
  n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
  n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
  n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
  n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
  n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
  n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
  n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
  n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
  n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
  n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
  n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
  n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
  n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6850, n6859, n11921, n11922, n11923, n11924, n11926, n11927, n11928, n11929, n11930, n11931, n11935, n11936, n11937, n11939, 
  n11940, n11941, n11942, n11943, n11944, n11946, n11947, n11948, n11949, n11950, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11970, n11971, n11973, n11976, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, 
  n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, 
  n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, 
  n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, 
  n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, 
  n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, 
  n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, 
  n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, 
  n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, 
  n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, 
  n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, 
  n12499, n12500, n12501, n12502, n13019, n13020, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, 
  n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, 
  n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, 
  n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, 
  n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, 
  n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, 
  n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, 
  n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, 
  n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, 
  n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, 
  n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, 
  n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, 
  n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, 
  n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, 
  n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, 
  n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, 
  n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, 
  n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, 
  n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, 
  n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, 
  n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14155, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, 
  n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, 
  n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, 
  n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, 
  n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14391, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, 
  n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, 
  n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, 
  n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, 
  n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, 
  n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, 
  n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, 
  n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, 
  n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, 
  n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, 
  n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, 
  n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14949, n14950, n14951, n14952, n14953, 
  n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, 
  n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, 
  n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, 
  n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, 
  n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, 
  n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, 
  n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, 
  n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, 
  n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, 
  n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, 
  n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15504, n15505, 
  n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15553, n15554, n15555, n15556, n15557, 
  n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, 
  n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, 
  n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, 
  n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, 
  n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, 
  n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, 
  n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, 
  n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, 
  n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, 
  n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, 
  n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, 
  n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, 
  n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, 
  n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, 
  n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, 
  n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, 
  n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, 
  n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16458, n16459, n16460, n16461, n16462, n16463, 
  n16464, n16465, n16466, n16467, n16468, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16523, 
  n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16553, n16554, n16555, n16556, n16558, n16559, n16560, n16561, n16563, n16564, n16565, n16566, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, 
  n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, 
  n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, 
  n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, 
  n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, 
  n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, 
  n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17041, n17043, n17045, n17047, n17049, n17051, n17053, n17055, n17057, n17059, n17061, n17063, n17065, n17067, n17069, n17071, n17073, n17075, n17077, n17079, n17081, n17083, n17085, n17087, 
  n17089, n17091, n17093, n17095, n17097, n17099, n17101, n17103, n17105, n17107, n17109, n17111, n17113, n17115, n17117, n17119, n17121, n17123, n17125, n17127, n17129, n17131, n17133, n17135, n17137, n17139, n17141, n17143, n17145, n17147, n17149, n17151, n17153, n17155, n17157, n17159, n17161, n17163, n17165, n17167, n17169, n17171, n17173, n17175, n17177, n17179, n17181, n17183, n17185, n17187, 
  n17189, n17191, n17193, n17195, n17197, n17199, n17201, n17203, n17205, n17207, n17209, n17211, n17213, n17215, n17217, n17219, n17221, n17223, n17225, n17227, n17229, n17231, n17233, n17235, n17237, n17239, n17241, n17243, n17245, n17247, n17249, n17251, n17253, n17255, n17257, n17259, n17261, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, 
  n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, 
  n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, 
  n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, 
  n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, 
  n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, 
  n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, 
  n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, 
  n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, 
  n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, 
  n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, 
  n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, 
  n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, 
  n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, 
  n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, 
  n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, 
  n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, 
  n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, 
  n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, 
  n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, 
  n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, 
  n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, 
  n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, 
  n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, 
  n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, 
  n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, 
  n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, 
  n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, 
  n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, 
  n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, 
  n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, 
  n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, 
  n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, 
  n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, 
  n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, 
  n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, 
  n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, 
  n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, 
  n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, 
  n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, _GFM_n2699, _GFM_n26980, _GFM_n2697, _GFM_n2696, _GFM_n2695, _GFM_n26940, _GFM_n26930, _GFM_n26921, _GFM_n26910, _GFM_n26900, _GFM_n2689, _GFM_n2688, _GFM_n26870, _GFM_n26860, _GFM_n2685, _GFM_n26840, _GFM_n2683, _GFM_n26820, _GFM_n26810, 
  _GFM_n26801, _GFM_n2679, _GFM_n2678, _GFM_n26770, _GFM_n26760, _GFM_n2675, _GFM_n26740, _GFM_n26730, _GFM_n2672, _GFM_n2671, _GFM_n26700, _GFM_n26690, _GFM_n2668, _GFM_n26670, _GFM_n2666, _GFM_n2665, _GFM_n2664, _GFM_n26630, _GFM_n26620, _GFM_n26611, _GFM_n26600, _GFM_n26590, _GFM_n2658, _GFM_n2657, _GFM_n26560, _GFM_n26550, _GFM_n2654, _GFM_n26530, _GFM_n2652, _GFM_n26510, _GFM_n26500, _GFM_n2649, _GFM_n2648, _GFM_n2647, _GFM_n26460, _GFM_n26450, _GFM_n2644, _GFM_n26430, _GFM_n26420, _GFM_n2641, _GFM_n26401, _GFM_n26390, _GFM_n26380, _GFM_n2637, _GFM_n26360, _GFM_n2635, _GFM_n2634, _GFM_n2633, _GFM_n26320, _GFM_n26310, 
  _GFM_n26301, _GFM_n26290, _GFM_n26280, _GFM_n2627, _GFM_n2626, _GFM_n26250, _GFM_n26240, _GFM_n2623, _GFM_n26220, _GFM_n2621, _GFM_n26200, _GFM_n26190, _GFM_n2618, _GFM_n2617, _GFM_n2616, _GFM_n26150, _GFM_n26140, _GFM_n2613, _GFM_n26120, _GFM_n26110, _GFM_n2610, _GFM_n2609, _GFM_n26080, _GFM_n26070, _GFM_n2606, _GFM_n26050, _GFM_n2604, _GFM_n2603, _GFM_n2602, _GFM_n26010, _GFM_n26000, _GFM_n2599, _GFM_n25980, _GFM_n25970, _GFM_n2596, _GFM_n2595, _GFM_n25940, _GFM_n25930, _GFM_n2592, _GFM_n25910, _GFM_n25901, _GFM_n25890, _GFM_n25880, _GFM_n2587, _GFM_n2586, _GFM_n2585, _GFM_n25840, _GFM_n25830, _GFM_n25821, _GFM_n25810, 
  _GFM_n25800, _GFM_n2579, _GFM_n2578, _GFM_n25770, _GFM_n25760, _GFM_n2575, _GFM_n25740, _GFM_n2573, _GFM_n2572, _GFM_n2571, _GFM_n25700, _GFM_n25690, _GFM_n2568, _GFM_n25670, _GFM_n25660, _GFM_n2565, _GFM_n2564, _GFM_n25630, _GFM_n25620, _GFM_n25611, _GFM_n25600, _GFM_n2559, _GFM_n25580, _GFM_n25570, _GFM_n2556, _GFM_n2555, _GFM_n2554, _GFM_n25530, _GFM_n25520, _GFM_n25511, _GFM_n25500, _GFM_n25490, _GFM_n2548, _GFM_n2547, _GFM_n25460, _GFM_n25450, _GFM_n2544, _GFM_n25430, _GFM_n2542, _GFM_n2541, _GFM_n2540, _GFM_n25390, _GFM_n25380, _GFM_n2537, _GFM_n25360, _GFM_n25350, _GFM_n2534, _GFM_n2533, _GFM_n25320, _GFM_n25310, 
  _GFM_n2530, _GFM_n25290, _GFM_n2528, _GFM_n25270, _GFM_n25260, _GFM_n2525, _GFM_n2524, _GFM_n2523, _GFM_n25220, _GFM_n25210, _GFM_n25201, _GFM_n25190, _GFM_n25180, _GFM_n2517, _GFM_n2516, _GFM_n25150, _GFM_n25140, _GFM_n2513, _GFM_n25120, _GFM_n2511, _GFM_n25101, _GFM_n2509, _GFM_n25080, _GFM_n25070, _GFM_n2506, _GFM_n25050, _GFM_n25040, _GFM_n2503, _GFM_n2502, _GFM_n25010, _GFM_n25000, _GFM_n2499, _GFM_n24980, _GFM_n2497, _GFM_n24960, _GFM_n24950, _GFM_n2494, _GFM_n2493, _GFM_n24921, _GFM_n24910, _GFM_n24900, _GFM_n2489, _GFM_n24880, _GFM_n24870, _GFM_n2486, _GFM_n2485, _GFM_n24840, _GFM_n24830, _GFM_n2482, _GFM_n24810, 
  _GFM_n2480, _GFM_n2479, _GFM_n2478, _GFM_n24770, _GFM_n24760, _GFM_n2475, _GFM_n24740, _GFM_n24730, _GFM_n2472, _GFM_n2471, _GFM_n24700, _GFM_n24690, _GFM_n2468, _GFM_n24670, _GFM_n2466, _GFM_n24650, _GFM_n24640, _GFM_n2463, _GFM_n2462, _GFM_n2461, _GFM_n24600, _GFM_n24590, _GFM_n2458, _GFM_n24570, _GFM_n24560, _GFM_n2455, _GFM_n2454, _GFM_n24530, _GFM_n24520, _GFM_n24511, _GFM_n24500, _GFM_n2449, _GFM_n2448, _GFM_n2447, _GFM_n24460, _GFM_n24450, _GFM_n2444, _GFM_n24430, _GFM_n24420, _GFM_n2441, _GFM_n24401, _GFM_n24390, _GFM_n24380, _GFM_n2437, _GFM_n24360, _GFM_n2435, _GFM_n24340, _GFM_n24330, _GFM_n2432, _GFM_n2431, 
  _GFM_n2430, _GFM_n24290, _GFM_n24280, _GFM_n2427, _GFM_n24260, _GFM_n24250, _GFM_n2424, _GFM_n2423, _GFM_n24220, _GFM_n24210, _GFM_n24201, _GFM_n24190, _GFM_n2418, _GFM_n2417, _GFM_n2416, _GFM_n24150, _GFM_n24140, _GFM_n2413, _GFM_n24120, _GFM_n24110, _GFM_n24101, _GFM_n2409, _GFM_n24080, _GFM_n24070, _GFM_n2406, _GFM_n24050, _GFM_n2404, _GFM_n24030, _GFM_n24020, _GFM_n2401, _GFM_n2400, _GFM_n2399, _GFM_n23980, _GFM_n23970, _GFM_n2396, _GFM_n23950, _GFM_n23940, _GFM_n2393, _GFM_n2392, _GFM_n23910, _GFM_n23900, _GFM_n2389, _GFM_n23880, _GFM_n2387, _GFM_n21360, _GFM_n21350, _GFM_n2134, _GFM_n21330, _GFM_n21320, _GFM_n2131, 
  _GFM_n21301, _GFM_n21290, _GFM_n21280, _GFM_n2127, _GFM_n21260, _GFM_n2125, _GFM_n21240, _GFM_n21230, _GFM_n2122, _GFM_n2121, _GFM_n184, _GFM_n18310, _GFM_n18210, _GFM_n181, _GFM_n18011, _GFM_n17911, _GFM_n178, _GFM_n177, _GFM_n17611, _GFM_n17511, _GFM_n174, _GFM_n17310, _GFM_n172, _GFM_n17110, _GFM_n17011, _GFM_n2120, _GFM_n21190, _GFM_n21180, _GFM_n2117, _GFM_n21160, _GFM_n21150, _GFM_n2114, _GFM_n2113, _GFM_n21120, _GFM_n21110, _GFM_n21101, _GFM_n21090, _GFM_n2108, _GFM_n2107, _GFM_n2106, _GFM_n21050, _GFM_n21040, _GFM_n2103, _GFM_n21020, _GFM_n21010, _GFM_n21001, _GFM_n2099, _GFM_n20980, _GFM_n20970, _GFM_n2096, 
  _GFM_n20950, _GFM_n2094, _GFM_n20930, _GFM_n20920, _GFM_n2091, _GFM_n2090, _GFM_n2089, _GFM_n20880, _GFM_n20870, _GFM_n2086, _GFM_n20850, _GFM_n20840, _GFM_n2083, _GFM_n2082, _GFM_n20810, _GFM_n20800, _GFM_n2079, _GFM_n20780, _GFM_n2077, _GFM_n2076, _GFM_n2075, _GFM_n20740, _GFM_n20730, _GFM_n20721, _GFM_n20710, _GFM_n20700, _GFM_n2069, _GFM_n2068, _GFM_n20670, _GFM_n20660, _GFM_n2065, _GFM_n20640, _GFM_n2063, _GFM_n20620, _GFM_n20610, _GFM_n20601, _GFM_n2059, _GFM_n2058, _GFM_n20570, _GFM_n20560, _GFM_n2055, _GFM_n20540, _GFM_n20530, _GFM_n2052, _GFM_n2051, _GFM_n20500, _GFM_n20490, _GFM_n2048, _GFM_n20470, _GFM_n2046, 
  _GFM_n2045, _GFM_n2044, _GFM_n20430, _GFM_n20420, _GFM_n20411, _GFM_n20400, _GFM_n20390, _GFM_n2038, _GFM_n2037, _GFM_n20360, _GFM_n20350, _GFM_n2034, _GFM_n20330, _GFM_n2032, _GFM_n20310, _GFM_n20300, _GFM_n2029, _GFM_n2028, _GFM_n2027, _GFM_n20260, _GFM_n20250, _GFM_n2024, _GFM_n20230, _GFM_n20220, _GFM_n2021, _GFM_n20201, _GFM_n20190, _GFM_n20180, _GFM_n2017, _GFM_n20160, _GFM_n2015, _GFM_n2014, _GFM_n2013, _GFM_n20120, _GFM_n20110, _GFM_n20101, _GFM_n20090, _GFM_n20080, _GFM_n2007, _GFM_n2006, _GFM_n20050, _GFM_n20040, _GFM_n2003, _GFM_n20020, _GFM_n2001, _GFM_n20000, _GFM_n19990, _GFM_n1998, _GFM_n1997, _GFM_n1996, 
  _GFM_n19950, _GFM_n19940, _GFM_n1993, _GFM_n19920, _GFM_n19910, _GFM_n1990, _GFM_n1989, _GFM_n19880, _GFM_n19870, _GFM_n1986, _GFM_n19850, _GFM_n1984, _GFM_n1983, _GFM_n1982, _GFM_n19810, _GFM_n19800, _GFM_n1979, _GFM_n19780, _GFM_n19770, _GFM_n1976, _GFM_n1975, _GFM_n19740, _GFM_n19730, _GFM_n1972, _GFM_n19710, _GFM_n19701, _GFM_n19690, _GFM_n19680, _GFM_n1967, _GFM_n1966, _GFM_n1965, _GFM_n19640, _GFM_n19630, _GFM_n19621, _GFM_n19610, _GFM_n19600, _GFM_n1959, _GFM_n1958, _GFM_n19570, _GFM_n19560, _GFM_n1955, _GFM_n19540, _GFM_n1953, _GFM_n1952, _GFM_n1951, _GFM_n19500, _GFM_n19490, _GFM_n1948, _GFM_n19470, _GFM_n19460, 
  _GFM_n1945, _GFM_n1944, _GFM_n19430, _GFM_n19420, _GFM_n19411, _GFM_n19400, _GFM_n1939, _GFM_n19380, _GFM_n19370, _GFM_n1936, _GFM_n1935, _GFM_n1934, _GFM_n19330, _GFM_n19320, _GFM_n19311, _GFM_n19300, _GFM_n19290, _GFM_n1928, _GFM_n1927, _GFM_n19260, _GFM_n19250, _GFM_n1924, _GFM_n19230, _GFM_n1922, _GFM_n1921, _GFM_n1920, _GFM_n19190, _GFM_n19180, _GFM_n1917, _GFM_n19160, _GFM_n19150, _GFM_n1914, _GFM_n1913, _GFM_n19120, _GFM_n19110, _GFM_n1910, _GFM_n19090, _GFM_n1908, _GFM_n19070, _GFM_n19060, _GFM_n1905, _GFM_n1904, _GFM_n1903, _GFM_n19020, _GFM_n19010, _GFM_n19001, _GFM_n18990, _GFM_n18980, _GFM_n1897, _GFM_n1896, 
  _GFM_n18950, _GFM_n18940, _GFM_n1893, _GFM_n18920, _GFM_n1891, _GFM_n18901, _GFM_n1889, _GFM_n18880, _GFM_n18870, _GFM_n1886, _GFM_n18850, _GFM_n18840, _GFM_n1883, _GFM_n1882, _GFM_n18810, _GFM_n18800, _GFM_n1879, _GFM_n18780, _GFM_n1877, _GFM_n18760, _GFM_n18750, _GFM_n1874, _GFM_n1873, _GFM_n18721, _GFM_n18710, _GFM_n18700, _GFM_n1869, _GFM_n18680, _GFM_n18670, _GFM_n1866, _GFM_n1865, _GFM_n18640, _GFM_n18630, _GFM_n1862, _GFM_n18610, _GFM_n1860, _GFM_n1859, _GFM_n1858, _GFM_n18570, _GFM_n18560, _GFM_n1855, _GFM_n18540, _GFM_n18530, _GFM_n1852, _GFM_n1851, _GFM_n18500, _GFM_n18490, _GFM_n1848, _GFM_n18470, _GFM_n1846, 
  _GFM_n18450, _GFM_n18440, _GFM_n1843, _GFM_n1842, _GFM_n1841, _GFM_n18400, _GFM_n18390, _GFM_n1838, _GFM_n18370, _GFM_n18360, _GFM_n1835, _GFM_n1834, _GFM_n18330, _GFM_n18320, _GFM_n1831, _GFM_n18300, _GFM_n1829, _GFM_n1828, _GFM_n1827, _GFM_n18260, _GFM_n18250, _GFM_n1824, _GFM_n18230, _GFM_n18220, _GFM_n1821, _GFM_n1820, _GFM_n18190, _GFM_n18180, _GFM_n1817, _GFM_n18160, _GFM_n1815, _GFM_n18140, _GFM_n18130, _GFM_n1812, _GFM_n1811, _GFM_n1810, _GFM_n18090, _GFM_n18080, _GFM_n1807, _GFM_n18060, _GFM_n18050, _GFM_n1804, _GFM_n1803, _GFM_n18020, _GFM_n18010, _GFM_n1800, _GFM_n17990, _GFM_n1798, _GFM_n1797, _GFM_n1796, 
  _GFM_n17950, _GFM_n17940, _GFM_n1793, _GFM_n17920, _GFM_n17910, _GFM_n1790, _GFM_n1789, _GFM_n17880, _GFM_n17870, _GFM_n1786, _GFM_n17850, _GFM_n1784, _GFM_n17830, _GFM_n17820, _GFM_n1781, _GFM_n1780, _GFM_n1779, _GFM_n17780, _GFM_n17770, _GFM_n1776, _GFM_n17750, _GFM_n17740, _GFM_n1773, _GFM_n1772, _GFM_n17710, _GFM_n17700, _GFM_n1769, _GFM_n17680, _GFM_n1767, _GFM_n1766, _GFM_n1765, _GFM_n17640, _GFM_n17630, _GFM_n1762, _GFM_n17610, _GFM_n17600, _GFM_n1759, _GFM_n1758, _GFM_n17570, _GFM_n17560, _GFM_n1755, _GFM_n17540, _GFM_n1753, _GFM_n17520, _GFM_n17510, _GFM_n1750, _GFM_n1749, _GFM_n1748, _GFM_n17470, _GFM_n17460, 
  _GFM_n1745, _GFM_n17440, _GFM_n17430, _GFM_n1742, _GFM_n1741, _GFM_n17400, _GFM_n17390, _GFM_n1738, _GFM_n17370, _GFM_n1736, _GFM_n1735, _GFM_n1734, _GFM_n17330, _GFM_n17320, _GFM_n1731, _GFM_n17300, _GFM_n17290, _GFM_n1728, _GFM_n1727, _GFM_n17260, _GFM_n17250, _GFM_n1724, _GFM_n17230, _GFM_n1722, _GFM_n17210, _GFM_n17200, _GFM_n1719, _GFM_n1718, _GFM_n1717, _GFM_n17160, _GFM_n17150, _GFM_n1714, _GFM_n17130, _GFM_n17120, _GFM_n1711, _GFM_n1710, _GFM_n17090, _GFM_n17080, _GFM_n1707, _GFM_n17060, _GFM_n1705, _GFM_n1704, _GFM_n1703, _GFM_n17020, _GFM_n17010, _GFM_n1700, _GFM_n16990, _GFM_n16980, _GFM_n1697, _GFM_n1696, 
  _GFM_n16950, _GFM_n16940, _GFM_n1693, _GFM_n16920, _GFM_n1691, _GFM_n16900, _GFM_n16890, _GFM_n1688, _GFM_n1687, _GFM_n1686, _GFM_n16850, _GFM_n16840, _GFM_n1683, _GFM_n16820, _GFM_n16810, _GFM_n1680, _GFM_n1679, _GFM_n16780, _GFM_n16770, _GFM_n1676, _GFM_n16750, _GFM_n1674, _GFM_n1673, _GFM_n1672, _GFM_n16710, _GFM_n16700, _GFM_n1669, _GFM_n16680, _GFM_n16670, _GFM_n1666, _GFM_n1665, _GFM_n16640, _GFM_n16630, _GFM_n1662, _GFM_n16610, _GFM_n1660, _GFM_n16590, _GFM_n16580, _GFM_n1657, _GFM_n1656, _GFM_n1655, _GFM_n16540, _GFM_n16530, _GFM_n1652, _GFM_n16510, _GFM_n16500, _GFM_n1649, _GFM_n1648, _GFM_n16470, _GFM_n16460, 
  _GFM_n1645, _GFM_n16440, _GFM_n1643, _GFM_n1642, _GFM_n1641, _GFM_n16400, _GFM_n16390, _GFM_n1638, _GFM_n16370, _GFM_n16360, _GFM_n1635, _GFM_n1634, _GFM_n16330, _GFM_n16320, _GFM_n1631, _GFM_n16300, _GFM_n1629, _GFM_n16280, _GFM_n16270, _GFM_n1626, _GFM_n1625, _GFM_n1624, _GFM_n16230, _GFM_n16220, _GFM_n1621, _GFM_n16200, _GFM_n16190, _GFM_n1618, _GFM_n1617, _GFM_n16160, _GFM_n16150, _GFM_n1614, _GFM_n16130, _GFM_n1612, _GFM_n1611, _GFM_n1610, _GFM_n16090, _GFM_n16080, _GFM_n1607, _GFM_n16060, _GFM_n16050, _GFM_n1604, _GFM_n1603, _GFM_n16020, _GFM_n16010, _GFM_n1600, _GFM_n15990, _GFM_n1598, _GFM_n15970, _GFM_n15960, 
  _GFM_n1595, _GFM_n1594, _GFM_n1593, _GFM_n15920, _GFM_n15910, _GFM_n1590, _GFM_n15890, _GFM_n15880, _GFM_n1587, _GFM_n1586, _GFM_n15850, _GFM_n15840, _GFM_n1583, _GFM_n15820, _GFM_n1581, _GFM_n1580, _GFM_n1579, _GFM_n15780, _GFM_n15770, _GFM_n1576, _GFM_n15750, _GFM_n15740, _GFM_n1573, _GFM_n1572, _GFM_n15710, _GFM_n15700, _GFM_n1569, _GFM_n15680, _GFM_n1567, _GFM_n15660, _GFM_n15650, _GFM_n1564, _GFM_n1563, _GFM_n1562, _GFM_n15610, _GFM_n15600, _GFM_n1559, _GFM_n15580, _GFM_n15570, _GFM_n1556, _GFM_n1555, _GFM_n15540, _GFM_n15530, _GFM_n1552, _GFM_n15510, _GFM_n1550, _GFM_n1549, _GFM_n1548, _GFM_n15470, _GFM_n15460, 
  _GFM_n1545, _GFM_n15440, _GFM_n15430, _GFM_n1542, _GFM_n1541, _GFM_n15400, _GFM_n15390, _GFM_n1538, _GFM_n15370, _GFM_n1536, _GFM_n15350, _GFM_n15340, _GFM_n1533, _GFM_n1532, _GFM_n1531, _GFM_n15300, _GFM_n15290, _GFM_n1528, _GFM_n15270, _GFM_n15260, _GFM_n1525, _GFM_n1524, _GFM_n15230, _GFM_n15220, _GFM_n1521, _GFM_n15200, _GFM_n1519, _GFM_n1518, _GFM_n1517, _GFM_n15160, _GFM_n15150, _GFM_n1514, _GFM_n15130, _GFM_n15120, _GFM_n1511, _GFM_n1510, _GFM_n15090, _GFM_n15080, _GFM_n1507, _GFM_n15060, _GFM_n1505, _GFM_n15040, _GFM_n15030, _GFM_n1502, _GFM_n1501, _GFM_n1500, _GFM_n14990, _GFM_n14980, _GFM_n1497, _GFM_n14960, 
  _GFM_n14950, _GFM_n1494, _GFM_n1493, _GFM_n14920, _GFM_n14910, _GFM_n1490, _GFM_n14890, _GFM_n1488, _GFM_n1487, _GFM_n1486, _GFM_n14850, _GFM_n14840, _GFM_n1483, _GFM_n14820, _GFM_n14810, _GFM_n1480, _GFM_n1479, _GFM_n14780, _GFM_n14770, _GFM_n1476, _GFM_n14750, _GFM_n1474, _GFM_n14730, _GFM_n14720, _GFM_n1471, _GFM_n1470, _GFM_n1469, _GFM_n14680, _GFM_n14670, _GFM_n1466, _GFM_n14650, _GFM_n14640, _GFM_n1463, _GFM_n1462, _GFM_n14610, _GFM_n14600, _GFM_n1459, _GFM_n14580, _GFM_n1457, _GFM_n1456, _GFM_n1455, _GFM_n14540, _GFM_n14530, _GFM_n1452, _GFM_n14510, _GFM_n14500, _GFM_n1449, _GFM_n1448, _GFM_n14470, _GFM_n14460, 
  _GFM_n1445, _GFM_n14440, _GFM_n1443, _GFM_n14420, _GFM_n14410, _GFM_n1440, _GFM_n1439, _GFM_n1438, _GFM_n14370, _GFM_n14360, _GFM_n1435, _GFM_n14340, _GFM_n14330, _GFM_n1432, _GFM_n1431, _GFM_n14300, _GFM_n14290, _GFM_n1428, _GFM_n14270, _GFM_n1426, _GFM_n1425, _GFM_n1424, _GFM_n14230, _GFM_n14220, _GFM_n1421, _GFM_n14200, _GFM_n14190, _GFM_n1418, _GFM_n1417, _GFM_n14160, _GFM_n14150, _GFM_n1414, _GFM_n14130, _GFM_n1412, _GFM_n14110, _GFM_n14100, _GFM_n1409, _GFM_n1408, _GFM_n1407, _GFM_n14060, _GFM_n14050, _GFM_n1404, _GFM_n14030, _GFM_n14020, _GFM_n1401, _GFM_n1400, _GFM_n13990, _GFM_n13980, _GFM_n1397, _GFM_n13960, 
  _GFM_n1395, _GFM_n1394, _GFM_n1393, _GFM_n13920, _GFM_n13910, _GFM_n1390, _GFM_n13890, _GFM_n13880, _GFM_n1387, _GFM_n1386, _GFM_n13850, _GFM_n13840, _GFM_n1383, _GFM_n13820, _GFM_n1381, _GFM_n13800, _GFM_n13790, _GFM_n1378, _GFM_n1377, _GFM_n1376, _GFM_n13750, _GFM_n13740, _GFM_n1373, _GFM_n13720, _GFM_n13710, _GFM_n1370, _GFM_n1369, _GFM_n13680, _GFM_n13670, _GFM_n1366, _GFM_n13650, _GFM_n1364, _GFM_n1363, _GFM_n1362, _GFM_n13610, _GFM_n13600, _GFM_n1359, _GFM_n13580, _GFM_n13570, _GFM_n1356, _GFM_n1355, _GFM_n13540, _GFM_n13530, _GFM_n1352, _GFM_n13510, _GFM_n1350, _GFM_n13490, _GFM_n13480, _GFM_n1347, _GFM_n1346, 
  _GFM_n1345, _GFM_n13440, _GFM_n13430, _GFM_n1342, _GFM_n13410, _GFM_n13400, _GFM_n1339, _GFM_n1338, _GFM_n13370, _GFM_n13360, _GFM_n1335, _GFM_n13340, _GFM_n1333, _GFM_n1332, _GFM_n1331, _GFM_n13300, _GFM_n13290, _GFM_n1328, _GFM_n13270, _GFM_n13260, _GFM_n1325, _GFM_n1324, _GFM_n13230, _GFM_n13220, _GFM_n1321, _GFM_n13200, _GFM_n1319, _GFM_n13180, _GFM_n13170, _GFM_n1316, _GFM_n1315, _GFM_n1314, _GFM_n13130, _GFM_n13120, _GFM_n1311, _GFM_n13100, _GFM_n13090, _GFM_n1308, _GFM_n1307, _GFM_n13060, _GFM_n13050, _GFM_n1304, _GFM_n13030, _GFM_n1302, _GFM_n1301, _GFM_n1300, _GFM_n12990, _GFM_n12980, _GFM_n1297, _GFM_n12960, 
  _GFM_n12950, _GFM_n1294, _GFM_n1293, _GFM_n12920, _GFM_n12910, _GFM_n1290, _GFM_n12890, _GFM_n1288, _GFM_n12870, _GFM_n12860, _GFM_n1285, _GFM_n1284, _GFM_n1283, _GFM_n12820, _GFM_n12810, _GFM_n1280, _GFM_n12790, _GFM_n12780, _GFM_n1277, _GFM_n1276, _GFM_n12750, _GFM_n12740, _GFM_n1273, _GFM_n12720, _GFM_n1271, _GFM_n1270, _GFM_n1269, _GFM_n12680, _GFM_n12670, _GFM_n1266, _GFM_n12650, _GFM_n12640, _GFM_n1263, _GFM_n1262, _GFM_n12610, _GFM_n12600, _GFM_n1259, _GFM_n12580, _GFM_n1257, _GFM_n12560, _GFM_n12550, _GFM_n1254, _GFM_n1253, _GFM_n1252, _GFM_n12510, _GFM_n12500, _GFM_n1249, _GFM_n12480, _GFM_n12470, _GFM_n1246, 
  _GFM_n1245, _GFM_n12440, _GFM_n12430, _GFM_n1242, _GFM_n12410, _GFM_n1240, _GFM_n1239, _GFM_n1238, _GFM_n12370, _GFM_n12360, _GFM_n1235, _GFM_n12340, _GFM_n12330, _GFM_n1232, _GFM_n1231, _GFM_n12300, _GFM_n12290, _GFM_n1228, _GFM_n12270, _GFM_n1226, _GFM_n12250, _GFM_n12240, _GFM_n1223, _GFM_n1222, _GFM_n1221, _GFM_n12200, _GFM_n12190, _GFM_n1218, _GFM_n12170, _GFM_n12160, _GFM_n1215, _GFM_n1214, _GFM_n12130, _GFM_n12120, _GFM_n1211, _GFM_n12100, _GFM_n1209, _GFM_n1208, _GFM_n1207, _GFM_n12060, _GFM_n12050, _GFM_n1204, _GFM_n12030, _GFM_n12020, _GFM_n1201, _GFM_n1200, _GFM_n11990, _GFM_n11980, _GFM_n1197, _GFM_n11960, 
  _GFM_n1195, _GFM_n11940, _GFM_n11930, _GFM_n1192, _GFM_n1191, _GFM_n1190, _GFM_n11890, _GFM_n11880, _GFM_n1187, _GFM_n11860, _GFM_n11850, _GFM_n1184, _GFM_n1183, _GFM_n11820, _GFM_n11810, _GFM_n1180, _GFM_n11790, _GFM_n1178, _GFM_n1177, _GFM_n1176, _GFM_n11750, _GFM_n11740, _GFM_n1173, _GFM_n11720, _GFM_n11710, _GFM_n1170, _GFM_n1169, _GFM_n11680, _GFM_n11670, _GFM_n1166, _GFM_n11650, _GFM_n1164, _GFM_n11630, _GFM_n11620, _GFM_n1161, _GFM_n1160, _GFM_n1159, _GFM_n11580, _GFM_n11570, _GFM_n1156, _GFM_n11550, _GFM_n11540, _GFM_n1153, _GFM_n1152, _GFM_n11510, _GFM_n11500, _GFM_n1149, _GFM_n11480, _GFM_n1147, _GFM_n1146, 
  _GFM_n1145, _GFM_n11440, _GFM_n11430, _GFM_n1142, _GFM_n11410, _GFM_n11400, _GFM_n1139, _GFM_n1138, _GFM_n11370, _GFM_n11360, _GFM_n1135, _GFM_n11340, _GFM_n1133, _GFM_n11320, _GFM_n11310, _GFM_n1130, _GFM_n1129, _GFM_n1128, _GFM_n11270, _GFM_n11260, _GFM_n1125, _GFM_n11240, _GFM_n11230, _GFM_n1122, _GFM_n1121, _GFM_n11200, _GFM_n11190, _GFM_n1118, _GFM_n11170, _GFM_n1116, _GFM_n1115, _GFM_n1114, _GFM_n11130, _GFM_n11120, _GFM_n1111, _GFM_n11100, _GFM_n11090, _GFM_n1108, _GFM_n1107, _GFM_n11060, _GFM_n11050, _GFM_n1104, _GFM_n11030, _GFM_n1102, _GFM_n11010, _GFM_n11000, _GFM_n1099, _GFM_n1098, _GFM_n1097, _GFM_n10960, 
  _GFM_n10950, _GFM_n1094, _GFM_n10930, _GFM_n10920, _GFM_n1091, _GFM_n1090, _GFM_n10890, _GFM_n10880, _GFM_n1087, _GFM_n10860, _GFM_n1085, _GFM_n1084, _GFM_n1083, _GFM_n10820, _GFM_n10810, _GFM_n1080, _GFM_n10790, _GFM_n10780, _GFM_n1077, _GFM_n1076, _GFM_n10750, _GFM_n10740, _GFM_n1073, _GFM_n10720, _GFM_n1071, _GFM_n10700, _GFM_n10690, _GFM_n1068, _GFM_n1067, _GFM_n1066, _GFM_n10650, _GFM_n10640, _GFM_n1063, _GFM_n10620, _GFM_n10610, _GFM_n1060, _GFM_n1059, _GFM_n10580, _GFM_n10570, _GFM_n1056, _GFM_n10550, _GFM_n1054, _GFM_n1053, _GFM_n1052, _GFM_n10510, _GFM_n10500, _GFM_n1049, _GFM_n10480, _GFM_n10470, _GFM_n1046, 
  _GFM_n1045, _GFM_n10440, _GFM_n10430, _GFM_n1042, _GFM_n10410, _GFM_n1040, _GFM_n10390, _GFM_n10380, _GFM_n1037, _GFM_n1036, _GFM_n1035, _GFM_n10340, _GFM_n10330, _GFM_n1032, _GFM_n10310, _GFM_n10300, _GFM_n1029, _GFM_n1028, _GFM_n10270, _GFM_n10260, _GFM_n1025, _GFM_n10240, _GFM_n1023, _GFM_n1022, _GFM_n1021, _GFM_n10200, _GFM_n10190, _GFM_n1018, _GFM_n10170, _GFM_n10160, _GFM_n1015, _GFM_n1014, _GFM_n10130, _GFM_n10120, _GFM_n1011, _GFM_n10100, _GFM_n1009, _GFM_n10080, _GFM_n10070, _GFM_n1006, _GFM_n1005, _GFM_n1004, _GFM_n10030, _GFM_n10020, _GFM_n1001, _GFM_n10000, _GFM_n9990, _GFM_n998, _GFM_n997, _GFM_n9960, 
  _GFM_n9950, _GFM_n994, _GFM_n9930, _GFM_n992, _GFM_n991, _GFM_n990, _GFM_n9890, _GFM_n9880, _GFM_n987, _GFM_n9860, _GFM_n9850, _GFM_n984, _GFM_n983, _GFM_n9820, _GFM_n9810, _GFM_n980, _GFM_n9790, _GFM_n978, _GFM_n9770, _GFM_n9760, _GFM_n975, _GFM_n974, _GFM_n973, _GFM_n9720, _GFM_n9710, _GFM_n970, _GFM_n9690, _GFM_n9680, _GFM_n967, _GFM_n966, _GFM_n9650, _GFM_n9640, _GFM_n963, _GFM_n9620, _GFM_n961, _GFM_n960, _GFM_n959, _GFM_n9580, _GFM_n9570, _GFM_n956, _GFM_n9550, _GFM_n9540, _GFM_n953, _GFM_n952, _GFM_n9510, _GFM_n9500, _GFM_n949, _GFM_n9480, _GFM_n947, _GFM_n9460, 
  _GFM_n9450, _GFM_n944, _GFM_n943, _GFM_n942, _GFM_n9410, _GFM_n9400, _GFM_n939, _GFM_n9380, _GFM_n9370, _GFM_n936, _GFM_n935, _GFM_n9340, _GFM_n9330, _GFM_n932, _GFM_n9310, _GFM_n930, _GFM_n929, _GFM_n928, _GFM_n9270, _GFM_n9260, _GFM_n925, _GFM_n9240, _GFM_n9230, _GFM_n922, _GFM_n921, _GFM_n9200, _GFM_n9190, _GFM_n918, _GFM_n9170, _GFM_n916, _GFM_n9150, _GFM_n9140, _GFM_n913, _GFM_n912, _GFM_n911, _GFM_n9100, _GFM_n9090, _GFM_n908, _GFM_n9070, _GFM_n9060, _GFM_n905, _GFM_n904, _GFM_n9030, _GFM_n9020, _GFM_n901, _GFM_n9000, _GFM_n899, _GFM_n898, _GFM_n897, _GFM_n8960, 
  _GFM_n8950, _GFM_n894, _GFM_n8930, _GFM_n8920, _GFM_n891, _GFM_n890, _GFM_n8890, _GFM_n8880, _GFM_n887, _GFM_n8860, _GFM_n885, _GFM_n8840, _GFM_n8830, _GFM_n882, _GFM_n881, _GFM_n880, _GFM_n8790, _GFM_n8780, _GFM_n877, _GFM_n8760, _GFM_n8750, _GFM_n874, _GFM_n873, _GFM_n8720, _GFM_n8710, _GFM_n870, _GFM_n8690, _GFM_n868, _GFM_n867, _GFM_n866, _GFM_n8650, _GFM_n8640, _GFM_n863, _GFM_n8620, _GFM_n8610, _GFM_n860, _GFM_n859, _GFM_n8580, _GFM_n8570, _GFM_n856, _GFM_n8550, _GFM_n854, _GFM_n8530, _GFM_n8520, _GFM_n851, _GFM_n850, _GFM_n849, _GFM_n8480, _GFM_n8470, _GFM_n846, 
  _GFM_n8450, _GFM_n8440, _GFM_n843, _GFM_n842, _GFM_n8410, _GFM_n8400, _GFM_n839, _GFM_n8380, _GFM_n837, _GFM_n836, _GFM_n835, _GFM_n8340, _GFM_n8330, _GFM_n832, _GFM_n8310, _GFM_n8300, _GFM_n829, _GFM_n828, _GFM_n8270, _GFM_n8260, _GFM_n825, _GFM_n8240, _GFM_n823, _GFM_n8220, _GFM_n8210, _GFM_n820, _GFM_n819, _GFM_n818, _GFM_n8170, _GFM_n8160, _GFM_n815, _GFM_n8140, _GFM_n8130, _GFM_n812, _GFM_n811, _GFM_n8100, _GFM_n8090, _GFM_n808, _GFM_n8070, _GFM_n806, _GFM_n805, _GFM_n804, _GFM_n8030, _GFM_n8020, _GFM_n801, _GFM_n8000, _GFM_n7990, _GFM_n798, _GFM_n797, _GFM_n7960, 
  _GFM_n7950, _GFM_n794, _GFM_n7930, _GFM_n792, _GFM_n7910, _GFM_n7900, _GFM_n789, _GFM_n788, _GFM_n787, _GFM_n7860, _GFM_n7850, _GFM_n784, _GFM_n7830, _GFM_n7820, _GFM_n781, _GFM_n780, _GFM_n7790, _GFM_n7780, _GFM_n777, _GFM_n7760, _GFM_n775, _GFM_n774, _GFM_n773, _GFM_n7720, _GFM_n7710, _GFM_n770, _GFM_n7690, _GFM_n7680, _GFM_n767, _GFM_n766, _GFM_n7650, _GFM_n7640, _GFM_n763, _GFM_n7620, _GFM_n761, _GFM_n7600, _GFM_n7590, _GFM_n758, _GFM_n757, _GFM_n756, _GFM_n7550, _GFM_n7540, _GFM_n753, _GFM_n7520, _GFM_n7510, _GFM_n750, _GFM_n749, _GFM_n7480, _GFM_n7470, _GFM_n746, 
  _GFM_n7450, _GFM_n744, _GFM_n743, _GFM_n742, _GFM_n7410, _GFM_n7400, _GFM_n739, _GFM_n7380, _GFM_n7370, _GFM_n736, _GFM_n735, _GFM_n7340, _GFM_n7330, _GFM_n732, _GFM_n7310, _GFM_n730, _GFM_n7290, _GFM_n7280, _GFM_n727, _GFM_n726, _GFM_n725, _GFM_n7240, _GFM_n7230, _GFM_n722, _GFM_n7210, _GFM_n7200, _GFM_n719, _GFM_n718, _GFM_n7170, _GFM_n7160, _GFM_n715, _GFM_n7140, _GFM_n713, _GFM_n712, _GFM_n711, _GFM_n7100, _GFM_n7090, _GFM_n708, _GFM_n7070, _GFM_n7060, _GFM_n705, _GFM_n704, _GFM_n7030, _GFM_n7020, _GFM_n701, _GFM_n7000, _GFM_n699, _GFM_n6980, _GFM_n6970, _GFM_n696, 
  _GFM_n695, _GFM_n694, _GFM_n6930, _GFM_n6920, _GFM_n691, _GFM_n6900, _GFM_n6890, _GFM_n688, _GFM_n687, _GFM_n6860, _GFM_n6850, _GFM_n684, _GFM_n6830, _GFM_n682, _GFM_n681, _GFM_n680, _GFM_n6790, _GFM_n6780, _GFM_n677, _GFM_n6760, _GFM_n6750, _GFM_n674, _GFM_n673, _GFM_n6720, _GFM_n6710, _GFM_n670, _GFM_n6690, _GFM_n668, _GFM_n6670, _GFM_n6660, _GFM_n665, _GFM_n664, _GFM_n663, _GFM_n6620, _GFM_n6610, _GFM_n660, _GFM_n6590, _GFM_n6580, _GFM_n657, _GFM_n656, _GFM_n6550, _GFM_n6540, _GFM_n653, _GFM_n6520, _GFM_n651, _GFM_n650, _GFM_n649, _GFM_n6480, _GFM_n6470, _GFM_n646, 
  _GFM_n6450, _GFM_n6440, _GFM_n643, _GFM_n642, _GFM_n6410, _GFM_n6400, _GFM_n639, _GFM_n6380, _GFM_n637, _GFM_n6360, _GFM_n6350, _GFM_n634, _GFM_n633, _GFM_n632, _GFM_n6310, _GFM_n6300, _GFM_n629, _GFM_n6280, _GFM_n6270, _GFM_n626, _GFM_n625, _GFM_n6240, _GFM_n6230, _GFM_n622, _GFM_n6210, _GFM_n620, _GFM_n619, _GFM_n618, _GFM_n6170, _GFM_n6160, _GFM_n615, _GFM_n6140, _GFM_n6130, _GFM_n612, _GFM_n611, _GFM_n6100, _GFM_n6090, _GFM_n608, _GFM_n6070, _GFM_n606, _GFM_n6050, _GFM_n6040, _GFM_n603, _GFM_n602, _GFM_n601, _GFM_n6000, _GFM_n5990, _GFM_n598, _GFM_n5970, _GFM_n5960, 
  _GFM_n595, _GFM_n594, _GFM_n5930, _GFM_n5920, _GFM_n591, _GFM_n5900, _GFM_n589, _GFM_n588, _GFM_n587, _GFM_n5860, _GFM_n5850, _GFM_n584, _GFM_n5830, _GFM_n5820, _GFM_n581, _GFM_n580, _GFM_n5790, _GFM_n5780, _GFM_n577, _GFM_n5760, _GFM_n575, _GFM_n5740, _GFM_n5730, _GFM_n572, _GFM_n571, _GFM_n570, _GFM_n5690, _GFM_n5680, _GFM_n567, _GFM_n5660, _GFM_n5650, _GFM_n564, _GFM_n563, _GFM_n5620, _GFM_n5610, _GFM_n560, _GFM_n5590, _GFM_n558, _GFM_n557, _GFM_n556, _GFM_n5550, _GFM_n5540, _GFM_n553, _GFM_n5520, _GFM_n5510, _GFM_n550, _GFM_n549, _GFM_n5480, _GFM_n5470, _GFM_n546, 
  _GFM_n5450, _GFM_n544, _GFM_n5430, _GFM_n5420, _GFM_n541, _GFM_n540, _GFM_n539, _GFM_n5380, _GFM_n5370, _GFM_n536, _GFM_n5350, _GFM_n5340, _GFM_n533, _GFM_n532, _GFM_n5310, _GFM_n5300, _GFM_n529, _GFM_n5280, _GFM_n527, _GFM_n526, _GFM_n525, _GFM_n5240, _GFM_n5230, _GFM_n522, _GFM_n5210, _GFM_n5200, _GFM_n519, _GFM_n518, _GFM_n5170, _GFM_n5160, _GFM_n515, _GFM_n5140, _GFM_n513, _GFM_n5120, _GFM_n5110, _GFM_n510, _GFM_n509, _GFM_n508, _GFM_n5070, _GFM_n5060, _GFM_n505, _GFM_n5040, _GFM_n5030, _GFM_n502, _GFM_n501, _GFM_n5000, _GFM_n4990, _GFM_n498, _GFM_n4970, _GFM_n496, 
  _GFM_n495, _GFM_n494, _GFM_n4930, _GFM_n4920, _GFM_n491, _GFM_n4900, _GFM_n4890, _GFM_n488, _GFM_n487, _GFM_n4860, _GFM_n4850, _GFM_n484, _GFM_n4830, _GFM_n482, _GFM_n4810, _GFM_n4800, _GFM_n479, _GFM_n478, _GFM_n477, _GFM_n4760, _GFM_n4750, _GFM_n474, _GFM_n4730, _GFM_n4720, _GFM_n471, _GFM_n470, _GFM_n4690, _GFM_n4680, _GFM_n467, _GFM_n4660, _GFM_n465, _GFM_n464, _GFM_n463, _GFM_n4620, _GFM_n4610, _GFM_n460, _GFM_n4590, _GFM_n4580, _GFM_n457, _GFM_n456, _GFM_n4550, _GFM_n4540, _GFM_n453, _GFM_n4520, _GFM_n451, _GFM_n4500, _GFM_n4490, _GFM_n448, _GFM_n447, _GFM_n446, 
  _GFM_n4450, _GFM_n4440, _GFM_n443, _GFM_n4420, _GFM_n4410, _GFM_n440, _GFM_n439, _GFM_n4380, _GFM_n4370, _GFM_n436, _GFM_n4350, _GFM_n434, _GFM_n433, _GFM_n432, _GFM_n4310, _GFM_n4301, _GFM_n429, _GFM_n4280, _GFM_n4270, _GFM_n426, _GFM_n425, _GFM_n4241, _GFM_n4230, _GFM_n422, _GFM_n4211, _GFM_n420, _GFM_n4190, _GFM_n4180, _GFM_n417, _GFM_n416, _GFM_n415, _GFM_n4140, _GFM_n4130, _GFM_n412, _GFM_n4110, _GFM_n4100, _GFM_n409, _GFM_n408, _GFM_n4070, _GFM_n4060, _GFM_n405, _GFM_n4040, _GFM_n403, _GFM_n402, _GFM_n401, _GFM_n4000, _GFM_n3991, _GFM_n398, _GFM_n3970, _GFM_n3960, 
  _GFM_n395, _GFM_n394, _GFM_n3930, _GFM_n3920, _GFM_n391, _GFM_n3900, _GFM_n389, _GFM_n3880, _GFM_n3870, _GFM_n386, _GFM_n385, _GFM_n384, _GFM_n3830, _GFM_n3820, _GFM_n381, _GFM_n3800, _GFM_n3790, _GFM_n378, _GFM_n377, _GFM_n3760, _GFM_n3751, _GFM_n374, _GFM_n3730, _GFM_n372, _GFM_n371, _GFM_n370, _GFM_n3691, _GFM_n3680, _GFM_n367, _GFM_n3660, _GFM_n3650, _GFM_n364, _GFM_n363, _GFM_n3621, _GFM_n3610, _GFM_n360, _GFM_n3590, _GFM_n358, _GFM_n3570, _GFM_n3560, _GFM_n355, _GFM_n354, _GFM_n353, _GFM_n3520, _GFM_n3510, _GFM_n350, _GFM_n3490, _GFM_n3480, _GFM_n347, _GFM_n346, 
  _GFM_n3451, _GFM_n3440, _GFM_n343, _GFM_n3420, _GFM_n341, _GFM_n340, _GFM_n339, _GFM_n3381, _GFM_n3370, _GFM_n336, _GFM_n3350, _GFM_n3342, _GFM_n333, _GFM_n332, _GFM_n3310, _GFM_n3300, _GFM_n329, _GFM_n3281, _GFM_n327, _GFM_n3260, _GFM_n3250, _GFM_n324, _GFM_n323, _GFM_n322, _GFM_n3210, _GFM_n3202, _GFM_n319, _GFM_n3181, _GFM_n3171, _GFM_n316, _GFM_n315, _GFM_n3140, _GFM_n3130, _GFM_n312, _GFM_n3112, _GFM_n310, _GFM_n309, _GFM_n308, _GFM_n3071, _GFM_n3060, _GFM_n305, _GFM_n3040, _GFM_n3030, _GFM_n302, _GFM_n301, _GFM_n3002, _GFM_n2990, _GFM_n298, _GFM_n2971, _GFM_n296, 
  _GFM_n2950, _GFM_n2940, _GFM_n293, _GFM_n292, _GFM_n291, _GFM_n2900, _GFM_n2892, _GFM_n288, _GFM_n2871, _GFM_n2861, _GFM_n285, _GFM_n284, _GFM_n2830, _GFM_n2820, _GFM_n281, _GFM_n2802, _GFM_n279, _GFM_n278, _GFM_n277, _GFM_n2761, _GFM_n2750, _GFM_n274, _GFM_n2730, _GFM_n2720, _GFM_n271, _GFM_n270, _GFM_n26920, _GFM_n26800, _GFM_n267, _GFM_n26610, _GFM_n265, _GFM_n26400, _GFM_n26300, _GFM_n262, _GFM_n261, _GFM_n260, _GFM_n25900, _GFM_n25820, _GFM_n257, _GFM_n25610, _GFM_n25510, _GFM_n254, _GFM_n253, _GFM_n25200, _GFM_n25100, _GFM_n250, _GFM_n24920, _GFM_n248, _GFM_n247, _GFM_n246, 
  _GFM_n24510, _GFM_n24400, _GFM_n243, _GFM_n24200, _GFM_n24100, _GFM_n240, _GFM_n239, _GFM_n2382, _GFM_n2370, _GFM_n236, _GFM_n2351, _GFM_n234, _GFM_n2330, _GFM_n2320, _GFM_n231, _GFM_n230, _GFM_n229, _GFM_n2280, _GFM_n2272, _GFM_n226, _GFM_n2251, _GFM_n2241, _GFM_n223, _GFM_n222, _GFM_n2210, _GFM_n2200, _GFM_n219, _GFM_n2182, _GFM_n217, _GFM_n216, _GFM_n215, _GFM_n2141, _GFM_n21300, _GFM_n212, _GFM_n21100, _GFM_n21000, _GFM_n209, _GFM_n208, _GFM_n20720, _GFM_n20600, _GFM_n205, _GFM_n20410, _GFM_n203, _GFM_n20200, _GFM_n20100, _GFM_n200, _GFM_n199, _GFM_n198, _GFM_n19700, _GFM_n19620, 
  _GFM_n195, _GFM_n19410, _GFM_n19310, _GFM_n192, _GFM_n191, _GFM_n19000, _GFM_n18900, _GFM_n188, _GFM_n18720, _GFM_n186, _GFM_n185, _GFM_N4349, _GFM_N4348, _GFM_N4346, _GFM_N4345, _GFM_N4342, _GFM_N4341, _GFM_N4339, _GFM_N4337, _GFM_N4336, _GFM_N4332, _GFM_N4331, _GFM_N4329, _GFM_N4328, _GFM_N4325, _GFM_N4324, _GFM_N4322, _GFM_N4318, _GFM_N4316, _GFM_N4313, _GFM_N4311, _GFM_N4307, _GFM_N4305, _GFM_N4302, _GFM_N4300, _GFM_N4295, _GFM_N4293, _GFM_N4290, _GFM_N4288, _GFM_N4284, _GFM_N4282, _GFM_N4279, _GFM_N4276, _GFM_N4272, _GFM_N4269, _GFM_N4265, _GFM_N4263, _GFM_N4258, _GFM_N4257, _GFM_N4255, 
  _GFM_N4254, _GFM_N4251, _GFM_N4250, _GFM_N4249, _GFM_N4248, _GFM_N4243, _GFM_N4242, _GFM_N4240, _GFM_N4239, _GFM_N4236, _GFM_N4235, _GFM_N4233, _GFM_N4232, _GFM_N4228, _GFM_N4227, _GFM_N4225, _GFM_N4224, _GFM_N4221, _GFM_N4218, _GFM_N4213, _GFM_N4210, _GFM_N4206, _GFM_N4203, _GFM_N4198, _GFM_N4195, _GFM_N4191, _GFM_N4188, _GFM_N4182, _GFM_N4179, _GFM_N4175, _GFM_N4172, _GFM_N4167, _GFM_N4164, _GFM_N4160, _GFM_N4159, _GFM_N4154, _GFM_N4151, _GFM_N4147, _GFM_N4144, _GFM_N4139, _GFM_N4136, _GFM_N4132, _GFM_N4129, _GFM_N4123, _GFM_N4120, _GFM_N4116, _GFM_N4113, _GFM_N4108, _GFM_N4106, _GFM_N4103, 
  _GFM_N4102, _GFM_N4097, _GFM_N4094, _GFM_N4090, _GFM_N4087, _GFM_N4082, _GFM_N4079, _GFM_N4075, _GFM_N4072, _GFM_N4066, _GFM_N4063, _GFM_N4059, _GFM_N4057, _GFM_N4052, _GFM_N4050, _GFM_N4049, _GFM_N4047, _GFM_N4042, _GFM_N4039, _GFM_N4035, _GFM_N4032, _GFM_N4027, _GFM_N4024, _GFM_N4020, _GFM_N4017, _GFM_N4012, _GFM_N4007, _GFM_N4006, _GFM_N4004, _GFM_N3999, _GFM_N3997, _GFM_N3996, _GFM_N3994, _GFM_N3990, _GFM_N3985, _GFM_N3981, _GFM_N3975, _GFM_N3971, _GFM_N3966, _GFM_N3962, _GFM_N3955, _GFM_N3951, _GFM_N3946, _GFM_N3944, _GFM_N3939, _GFM_N3936, _GFM_N3934, _GFM_N3931, _GFM_N3928, _GFM_N3923, 
  _GFM_N3918, _GFM_N3914, _GFM_N3908, _GFM_N3904, _GFM_N3899, _GFM_N3895, _GFM_N3889, _GFM_N3883, _GFM_N3881, _GFM_N3879, _GFM_N3874, _GFM_N3871, _GFM_N3869, _GFM_N3865, _GFM_N3864, _GFM_N3859, _GFM_N3854, _GFM_N3850, _GFM_N3844, _GFM_N3840, _GFM_N3835, _GFM_N3831, _GFM_N3825, _GFM_N3821, _GFM_N3818, _GFM_N3816, _GFM_N3812, _GFM_N3809, _GFM_N3808, _GFM_N3804, _GFM_N3803, _GFM_N3798, _GFM_N3793, _GFM_N3789, _GFM_N3783, _GFM_N3780, _GFM_N3775, _GFM_N3771, _GFM_N3764, _GFM_N3762, _GFM_N3759, _GFM_N3756, _GFM_N3754, _GFM_N3750, _GFM_N3748, _GFM_N3747, _GFM_N3745, _GFM_N3740, _GFM_N3735, _GFM_N3731, 
  _GFM_N3725, _GFM_N3723, _GFM_N3719, _GFM_N3715, _GFM_N3708, _GFM_N3706, _GFM_N3703, _GFM_N3701, _GFM_N3699, _GFM_N3695, _GFM_N3693, _GFM_N3692, _GFM_N3690, _GFM_N3685, _GFM_N3681, _GFM_N3674, _GFM_N3672, _GFM_N3670, _GFM_N3666, _GFM_N3662, _GFM_N3655, _GFM_N3653, _GFM_N3649, _GFM_N3648, _GFM_N3647, _GFM_N3643, _GFM_N3641, _GFM_N3640, _GFM_N3638, _GFM_N3633, _GFM_N3629, _GFM_N3623, _GFM_N3620, _GFM_N3618, _GFM_N3615, _GFM_N3611, _GFM_N3605, _GFM_N3603, _GFM_N3600, _GFM_N3598, _GFM_N3597, _GFM_N3594, _GFM_N3592, _GFM_N3591, _GFM_N3589, _GFM_N3584, _GFM_N3580, _GFM_N3574, _GFM_N3571, _GFM_N3569, 
  _GFM_N3566, _GFM_N3563, _GFM_N3558, _GFM_N3556, _GFM_N3554, _GFM_N3552, _GFM_N3551, _GFM_N3548, _GFM_N3546, _GFM_N3545, _GFM_N3543, _GFM_N3538, _GFM_N3534, _GFM_N3529, _GFM_N3527, _GFM_N3524, _GFM_N3521, _GFM_N3519, _GFM_N3514, _GFM_N3513, _GFM_N3511, _GFM_N3509, _GFM_N3508, _GFM_N3505, _GFM_N3503, _GFM_N3502, _GFM_N3500, _GFM_N3495, _GFM_N3491, _GFM_N3489, _GFM_N3484, _GFM_N3483, _GFM_N3482, _GFM_N3479, _GFM_N3477, _GFM_N3472, _GFM_N3471, _GFM_N3469, _GFM_N3467, _GFM_N3466, _GFM_N3463, _GFM_N3462, _GFM_N3460, _GFM_N3455, _GFM_N3452, _GFM_N3450, _GFM_N3446, _GFM_N3444, _GFM_N3443, _GFM_N3441, 
  _GFM_N3439, _GFM_N3434, _GFM_N3433, _GFM_N3431, _GFM_N3429, _GFM_N3428, _GFM_N3425, _GFM_N3424, _GFM_N3422, _GFM_N3418, _GFM_N3415, _GFM_N3413, _GFM_N3409, _GFM_N3407, _GFM_N3406, _GFM_N3404, _GFM_N3402, _GFM_N3398, _GFM_N3397, _GFM_N3395, _GFM_N3393, _GFM_N3392, _GFM_N3389, _GFM_N3388, _GFM_N3386, _GFM_N3383, _GFM_N3380, _GFM_N3378, _GFM_N3374, _GFM_N3373, _GFM_N3371, _GFM_N3369, _GFM_N3368, _GFM_N3364, _GFM_N3363, _GFM_N3361, _GFM_N3359, _GFM_N3358, _GFM_N3355, _GFM_N3354, _GFM_N3352, _GFM_N3349, _GFM_N3346, _GFM_N3345, _GFM_N3341, _GFM_N3340, _GFM_N3338, _GFM_N3336, _GFM_N3335, _GFM_N3331, 
  _GFM_N3330, _GFM_N3328, _GFM_N3326, _GFM_N3325, _GFM_N3322, _GFM_N3321, _GFM_N3319, _GFM_N3316, _GFM_N3313, _GFM_N3312, _GFM_N3309, _GFM_N3308, _GFM_N3306, _GFM_N3304, _GFM_N3303, _GFM_N3299, _GFM_N3298, _GFM_N3296, _GFM_N3294, _GFM_N3293, _GFM_N3290, _GFM_N3289, _GFM_N3287, _GFM_N3283, _GFM_N3282, _GFM_N3280, _GFM_N3279, _GFM_N3276, _GFM_N3275, _GFM_N3273, _GFM_N3271, _GFM_N3270, _GFM_N3266, _GFM_N3265, _GFM_N3263, _GFM_N3262, _GFM_N3259, _GFM_N3258, _GFM_N3256, _GFM_N3252, _GFM_N3251, _GFM_N3249, _GFM_N3248, _GFM_N3245, _GFM_N3244, _GFM_N3242, _GFM_N3240, _GFM_N3239, _GFM_N3235, _GFM_N3234, 
  _GFM_N3232, _GFM_N3231, _GFM_N3228, _GFM_N3227, _GFM_N3225, _GFM_N3221, _GFM_N3220, _GFM_N3218, _GFM_N3217, _GFM_N3214, _GFM_N3213, _GFM_N3211, _GFM_N3209, _GFM_N3208, _GFM_N3204, _GFM_N3203, _GFM_N3201, _GFM_N3200, _GFM_N3197, _GFM_N3196, _GFM_N3194, _GFM_N3190, _GFM_N3189, _GFM_N3187, _GFM_N3186, _GFM_N3183, _GFM_N3182, _GFM_N3180, _GFM_N3178, _GFM_N3177, _GFM_N3173, _GFM_N3172, _GFM_N3170, _GFM_N3169, _GFM_N3166, _GFM_N3165, _GFM_N3163, _GFM_N3159, _GFM_N3158, _GFM_N3156, _GFM_N3155, _GFM_N3152, _GFM_N3151, _GFM_N3149, _GFM_N3147, _GFM_N3146, _GFM_N3142, _GFM_N3141, _GFM_N3139, _GFM_N3138, 
  _GFM_N3135, _GFM_N3134, _GFM_N3132, _GFM_N3128, _GFM_N3127, _GFM_N3125, _GFM_N3124, _GFM_N3121, _GFM_N3120, _GFM_N3118, _GFM_N3116, _GFM_N3115, _GFM_N3111, _GFM_N3110, _GFM_N3108, _GFM_N3107, _GFM_N3104, _GFM_N3103, _GFM_N3101, _GFM_N3097, _GFM_N3096, _GFM_N3094, _GFM_N3093, _GFM_N3090, _GFM_N3089, _GFM_N3087, _GFM_N3085, _GFM_N3084, _GFM_N3080, _GFM_N3079, _GFM_N3077, _GFM_N3076, _GFM_N3073, _GFM_N3072, _GFM_N3070, _GFM_N3066, _GFM_N3065, _GFM_N3063, _GFM_N3062, _GFM_N3059, _GFM_N3058, _GFM_N3056, _GFM_N3054, _GFM_N3053, _GFM_N3049, _GFM_N3048, _GFM_N3046, _GFM_N3045, _GFM_N3042, _GFM_N3041, 
  _GFM_N3039, _GFM_N3035, _GFM_N3034, _GFM_N3032, _GFM_N3031, _GFM_N3028, _GFM_N3027, _GFM_N3025, _GFM_N3023, _GFM_N3022, _GFM_N3018, _GFM_N3017, _GFM_N3015, _GFM_N3014, _GFM_N3011, _GFM_N3010, _GFM_N3008, _GFM_N3004, _GFM_N3003, _GFM_N3001, _GFM_N3000, _GFM_N2997, _GFM_N2996, _GFM_N2994, _GFM_N2992, _GFM_N2991, _GFM_N2987, _GFM_N2986, _GFM_N2984, _GFM_N2983, _GFM_N2980, _GFM_N2979, _GFM_N2977, _GFM_N2973, _GFM_N2972, _GFM_N2970, _GFM_N2969, _GFM_N2966, _GFM_N2965, _GFM_N2963, _GFM_N2961, _GFM_N2960, _GFM_N2956, _GFM_N2955, _GFM_N2953, _GFM_N2952, _GFM_N2949, _GFM_N2948, _GFM_N2946, _GFM_N2942, 
  _GFM_N2941, _GFM_N2939, _GFM_N2938, _GFM_N2935, _GFM_N2934, _GFM_N2932, _GFM_N2930, _GFM_N2929, _GFM_N2925, _GFM_N2924, _GFM_N2922, _GFM_N2921, _GFM_N2918, _GFM_N2917, _GFM_N2915, _GFM_N2911, _GFM_N2910, _GFM_N2908, _GFM_N2907, _GFM_N2904, _GFM_N2903, _GFM_N2901, _GFM_N2899, _GFM_N2898, _GFM_N2894, _GFM_N2893, _GFM_N2891, _GFM_N2890, _GFM_N2887, _GFM_N2886, _GFM_N2884, _GFM_N2880, _GFM_N2879, _GFM_N2877, _GFM_N2876, _GFM_N2873, _GFM_N2872, _GFM_N2870, _GFM_N2868, _GFM_N2867, _GFM_N2863, _GFM_N2862, _GFM_N2860, _GFM_N2859, _GFM_N2856, _GFM_N2855, _GFM_N2853, _GFM_N2849, _GFM_N2848, _GFM_N2846, 
  _GFM_N2845, _GFM_N2842, _GFM_N2841, _GFM_N2839, _GFM_N2837, _GFM_N2836, _GFM_N2832, _GFM_N2831, _GFM_N2829, _GFM_N2828, _GFM_N2825, _GFM_N2824, _GFM_N2822, _GFM_N2818, _GFM_N2817, _GFM_N2815, _GFM_N2814, _GFM_N2811, _GFM_N2810, _GFM_N2808, _GFM_N2806, _GFM_N2805, _GFM_N2801, _GFM_N2800, _GFM_N2798, _GFM_N2797, _GFM_N2794, _GFM_N2793, _GFM_N2791, _GFM_N2787, _GFM_N2786, _GFM_N2784, _GFM_N2783, _GFM_N2780, _GFM_N2779, _GFM_N2777, _GFM_N2775, _GFM_N2774, _GFM_N2770, _GFM_N2769, _GFM_N2767, _GFM_N2766, _GFM_N2763, _GFM_N2762, _GFM_N2760, _GFM_N2756, _GFM_N2755, _GFM_N2753, _GFM_N2752, _GFM_N2749, 
  _GFM_N2748, _GFM_N2746, _GFM_N2744, _GFM_N2743, _GFM_N2739, _GFM_N2738, _GFM_N2736, _GFM_N2735, _GFM_N2732, _GFM_N2731, _GFM_N2729, _GFM_N2725, _GFM_N2724, _GFM_N2722, _GFM_N2721, _GFM_N2718, _GFM_N2717, _GFM_N2715, _GFM_N2713, _GFM_N2712, _GFM_N2708, _GFM_N2707, _GFM_N2705, _GFM_N2704, _GFM_N2701, _GFM_N2700, _GFM_N2698, _GFM_N2694, _GFM_N2693, _GFM_N2691, _GFM_N2690, _GFM_N2687, _GFM_N2686, _GFM_N2684, _GFM_N2682, _GFM_N2681, _GFM_N2677, _GFM_N2676, _GFM_N2674, _GFM_N2673, _GFM_N2670, _GFM_N2669, _GFM_N2667, _GFM_N2663, _GFM_N2662, _GFM_N2660, _GFM_N2659, _GFM_N2656, _GFM_N2655, _GFM_N2653, 
  _GFM_N2651, _GFM_N2650, _GFM_N2646, _GFM_N2645, _GFM_N2643, _GFM_N2642, _GFM_N2639, _GFM_N2638, _GFM_N2636, _GFM_N2632, _GFM_N2631, _GFM_N2629, _GFM_N2628, _GFM_N2625, _GFM_N2624, _GFM_N2622, _GFM_N2620, _GFM_N2619, _GFM_N2615, _GFM_N2614, _GFM_N2612, _GFM_N2611, _GFM_N2608, _GFM_N2607, _GFM_N2605, _GFM_N2601, _GFM_N2600, _GFM_N2598, _GFM_N2597, _GFM_N2594, _GFM_N2593, _GFM_N2591, _GFM_N2589, _GFM_N2588, _GFM_N2584, _GFM_N2583, _GFM_N2581, _GFM_N2580, _GFM_N2577, _GFM_N2576, _GFM_N2574, _GFM_N2570, _GFM_N2569, _GFM_N2567, _GFM_N2566, _GFM_N2563, _GFM_N2562, _GFM_N2560, _GFM_N2558, _GFM_N2557, 
  _GFM_N2553, _GFM_N2552, _GFM_N2550, _GFM_N2549, _GFM_N2546, _GFM_N2545, _GFM_N2543, _GFM_N2539, _GFM_N2538, _GFM_N2536, _GFM_N2535, _GFM_N2532, _GFM_N2531, _GFM_N2529, _GFM_N2527, _GFM_N2526, _GFM_N2522, _GFM_N2521, _GFM_N2519, _GFM_N2518, _GFM_N2515, _GFM_N2514, _GFM_N2512, _GFM_N2508, _GFM_N2507, _GFM_N2505, _GFM_N2504, _GFM_N2501, _GFM_N2500, _GFM_N2498, _GFM_N2496, _GFM_N2495, _GFM_N2491, _GFM_N2490, _GFM_N2488, _GFM_N2487, _GFM_N2484, _GFM_N2483, _GFM_N2481, _GFM_N2477, _GFM_N2476, _GFM_N2474, _GFM_N2473, _GFM_N2470, _GFM_N2469, _GFM_N2467, _GFM_N2465, _GFM_N2464, _GFM_N2460, _GFM_N2459, 
  _GFM_N2457, _GFM_N2456, _GFM_N2453, _GFM_N2452, _GFM_N2450, _GFM_N2446, _GFM_N2445, _GFM_N2443, _GFM_N2442, _GFM_N2439, _GFM_N2438, _GFM_N2436, _GFM_N2434, _GFM_N2433, _GFM_N2429, _GFM_N2428, _GFM_N2426, _GFM_N2425, _GFM_N2422, _GFM_N2421, _GFM_N2419, _GFM_N2415, _GFM_N2414, _GFM_N2412, _GFM_N2411, _GFM_N2408, _GFM_N2407, _GFM_N2405, _GFM_N2403, _GFM_N2402, _GFM_N2398, _GFM_N2397, _GFM_N2395, _GFM_N2394, _GFM_N2391, _GFM_N2390, _GFM_N2388, _GFM_N2384, _GFM_N2383, _GFM_N2381, _GFM_N2380, _GFM_N2377, _GFM_N2376, _GFM_N2374, _GFM_N2372, _GFM_N2371, _GFM_N2367, _GFM_N2366, _GFM_N2364, _GFM_N2363, 
  _GFM_N2360, _GFM_N2359, _GFM_N2357, _GFM_N2353, _GFM_N2352, _GFM_N2350, _GFM_N2349, _GFM_N2346, _GFM_N2345, _GFM_N2343, _GFM_N2341, _GFM_N2340, _GFM_N2336, _GFM_N2335, _GFM_N2333, _GFM_N2332, _GFM_N2329, _GFM_N2328, _GFM_N2326, _GFM_N2322, _GFM_N2321, _GFM_N2319, _GFM_N2318, _GFM_N2315, _GFM_N2314, _GFM_N2312, _GFM_N2310, _GFM_N2309, _GFM_N2305, _GFM_N2304, _GFM_N2302, _GFM_N2301, _GFM_N2298, _GFM_N2297, _GFM_N2295, _GFM_N2291, _GFM_N2290, _GFM_N2288, _GFM_N2287, _GFM_N2284, _GFM_N2283, _GFM_N2281, _GFM_N2279, _GFM_N2278, _GFM_N2274, _GFM_N2273, _GFM_N2271, _GFM_N2270, _GFM_N2267, _GFM_N2266, 
  _GFM_N2264, _GFM_N2260, _GFM_N2259, _GFM_N2257, _GFM_N2256, _GFM_N2253, _GFM_N2252, _GFM_N2250, _GFM_N2248, _GFM_N2247, _GFM_N2243, _GFM_N2242, _GFM_N2240, _GFM_N2239, _GFM_N2236, _GFM_N2235, _GFM_N2233, _GFM_N2229, _GFM_N2228, _GFM_N2226, _GFM_N2225, _GFM_N2222, _GFM_N2221, _GFM_N2219, _GFM_N2217, _GFM_N2216, _GFM_N2212, _GFM_N2211, _GFM_N2209, _GFM_N2208, _GFM_N2205, _GFM_N2204, _GFM_N2202, _GFM_N2198, _GFM_N2197, _GFM_N2195, _GFM_N2194, _GFM_N2191, _GFM_N2190, _GFM_N2188, _GFM_N2186, _GFM_N2185, _GFM_N2181, _GFM_N2180, _GFM_N2178, _GFM_N2177, _GFM_N2174, _GFM_N2173, _GFM_N2171, _GFM_N2167, 
  _GFM_N2166, _GFM_N2164, _GFM_N2163, _GFM_N2160, _GFM_N2159, _GFM_N2157, _GFM_N2155, _GFM_N2154, _GFM_N2150, _GFM_N2149, _GFM_N2147, _GFM_N2146, _GFM_N2143, _GFM_N2142, _GFM_N2140, _GFM_N2136, _GFM_N2135, _GFM_N2133, _GFM_N2132, _GFM_N2129, _GFM_N2128, _GFM_N2126, _GFM_N2124, _GFM_N2123, _GFM_N2119, _GFM_N2118, _GFM_N2116, _GFM_N2115, _GFM_N2112, _GFM_N2111, _GFM_N2109, _GFM_N2105, _GFM_N2104, _GFM_N2102, _GFM_N2101, _GFM_N2098, _GFM_N2097, _GFM_N2095, _GFM_N2093, _GFM_N2092, _GFM_N2088, _GFM_N2087, _GFM_N2085, _GFM_N2084, _GFM_N2081, _GFM_N2080, _GFM_N2078, _GFM_N2074, _GFM_N2073, _GFM_N2071, 
  _GFM_N2070, _GFM_N2067, _GFM_N2066, _GFM_N2064, _GFM_N2062, _GFM_N2061, _GFM_N2057, _GFM_N2056, _GFM_N2054, _GFM_N2053, _GFM_N2050, _GFM_N2049, _GFM_N2047, _GFM_N2043, _GFM_N2042, _GFM_N2040, _GFM_N2039, _GFM_N2036, _GFM_N2035, _GFM_N2033, _GFM_N2031, _GFM_N2030, _GFM_N2026, _GFM_N2025, _GFM_N2023, _GFM_N2022, _GFM_N2019, _GFM_N2018, _GFM_N2016, _GFM_N2012, _GFM_N2011, _GFM_N2009, _GFM_N2008, _GFM_N2005, _GFM_N2004, _GFM_N2002, _GFM_N2000, _GFM_N1999, _GFM_N1995, _GFM_N1994, _GFM_N1992, _GFM_N1991, _GFM_N1988, _GFM_N1987, _GFM_N1985, _GFM_N1981, _GFM_N1980, _GFM_N1978, _GFM_N1977, _GFM_N1974, 
  _GFM_N1973, _GFM_N1971, _GFM_N1969, _GFM_N1968, _GFM_N1964, _GFM_N1963, _GFM_N1961, _GFM_N1960, _GFM_N1957, _GFM_N1956, _GFM_N1954, _GFM_N1950, _GFM_N1949, _GFM_N1947, _GFM_N1946, _GFM_N1943, _GFM_N1942, _GFM_N1940, _GFM_N1938, _GFM_N1937, _GFM_N1933, _GFM_N1932, _GFM_N1930, _GFM_N1929, _GFM_N1926, _GFM_N1925, _GFM_N1923, _GFM_N1919, _GFM_N1918, _GFM_N1916, _GFM_N1915, _GFM_N1912, _GFM_N1911, _GFM_N1909, _GFM_N1907, _GFM_N1906, _GFM_N1902, _GFM_N1901, _GFM_N1899, _GFM_N1898, _GFM_N1895, _GFM_N1894, _GFM_N1892, _GFM_N1888, _GFM_N1887, _GFM_N1885, _GFM_N1884, _GFM_N1881, _GFM_N1880, _GFM_N1878, 
  _GFM_N1876, _GFM_N1875, _GFM_N1871, _GFM_N1870, _GFM_N1868, _GFM_N1867, _GFM_N1864, _GFM_N1863, _GFM_N1861, _GFM_N1857, _GFM_N1856, _GFM_N1854, _GFM_N1853, _GFM_N1850, _GFM_N1849, _GFM_N1847, _GFM_N1845, _GFM_N1844, _GFM_N1840, _GFM_N1839, _GFM_N1837, _GFM_N1836, _GFM_N1833, _GFM_N1832, _GFM_N1830, _GFM_N1826, _GFM_N1825, _GFM_N1823, _GFM_N1822, _GFM_N1819, _GFM_N1818, _GFM_N1816, _GFM_N1814, _GFM_N1813, _GFM_N1809, _GFM_N1808, _GFM_N1806, _GFM_N1805, _GFM_N1802, _GFM_N1801, _GFM_N1799, _GFM_N1795, _GFM_N1794, _GFM_N1792, _GFM_N1791, _GFM_N1788, _GFM_N1787, _GFM_N1785, _GFM_N1783, _GFM_N1782, 
  _GFM_N1778, _GFM_N1777, _GFM_N1775, _GFM_N1774, _GFM_N1771, _GFM_N1770, _GFM_N1768, _GFM_N1764, _GFM_N1763, _GFM_N1761, _GFM_N1760, _GFM_N1757, _GFM_N1756, _GFM_N1754, _GFM_N1752, _GFM_N1751, _GFM_N1747, _GFM_N1746, _GFM_N1744, _GFM_N1743, _GFM_N1740, _GFM_N1739, _GFM_N1737, _GFM_N1733, _GFM_N1732, _GFM_N1730, _GFM_N1729, _GFM_N1726, _GFM_N1725, _GFM_N1723, _GFM_N1721, _GFM_N1720, _GFM_N1716, _GFM_N1715, _GFM_N1713, _GFM_N1712, _GFM_N1709, _GFM_N1708, _GFM_N1706, _GFM_N1702, _GFM_N1701, _GFM_N1699, _GFM_N1698, _GFM_N1695, _GFM_N1694, _GFM_N1692, _GFM_N1690, _GFM_N1689, _GFM_N1685, _GFM_N1684, 
  _GFM_N1682, _GFM_N1681, _GFM_N1678, _GFM_N1677, _GFM_N1675, _GFM_N1671, _GFM_N1670, _GFM_N1668, _GFM_N1667, _GFM_N1664, _GFM_N1663, _GFM_N1661, _GFM_N1659, _GFM_N1658, _GFM_N1654, _GFM_N1653, _GFM_N1651, _GFM_N1650, _GFM_N1647, _GFM_N1646, _GFM_N1644, _GFM_N1640, _GFM_N1639, _GFM_N1637, _GFM_N1636, _GFM_N1633, _GFM_N1632, _GFM_N1630, _GFM_N1628, _GFM_N1627, _GFM_N1623, _GFM_N1622, _GFM_N1620, _GFM_N1619, _GFM_N1616, _GFM_N1615, _GFM_N1613, _GFM_N1609, _GFM_N1608, _GFM_N1606, _GFM_N1605, _GFM_N1602, _GFM_N1601, _GFM_N1599, _GFM_N1597, _GFM_N1596, _GFM_N1592, _GFM_N1591, _GFM_N1589, _GFM_N1588, 
  _GFM_N1585, _GFM_N1584, _GFM_N1582, _GFM_N1578, _GFM_N1577, _GFM_N1575, _GFM_N1574, _GFM_N1571, _GFM_N1570, _GFM_N1568, _GFM_N1566, _GFM_N1565, _GFM_N1561, _GFM_N1560, _GFM_N1558, _GFM_N1557, _GFM_N1554, _GFM_N1553, _GFM_N1551, _GFM_N1547, _GFM_N1546, _GFM_N1544, _GFM_N1543, _GFM_N1540, _GFM_N1539, _GFM_N1537, _GFM_N1535, _GFM_N1534, _GFM_N1530, _GFM_N1529, _GFM_N1527, _GFM_N1526, _GFM_N1523, _GFM_N1522, _GFM_N1520, _GFM_N1516, _GFM_N1515, _GFM_N1513, _GFM_N1512, _GFM_N1509, _GFM_N1508, _GFM_N1506, _GFM_N1504, _GFM_N1503, _GFM_N1499, _GFM_N1498, _GFM_N1496, _GFM_N1495, _GFM_N1492, _GFM_N1491, 
  _GFM_N1489, _GFM_N1485, _GFM_N1484, _GFM_N1482, _GFM_N1481, _GFM_N1478, _GFM_N1477, _GFM_N1475, _GFM_N1473, _GFM_N1472, _GFM_N1468, _GFM_N1467, _GFM_N1465, _GFM_N1464, _GFM_N1461, _GFM_N1460, _GFM_N1458, _GFM_N1454, _GFM_N1453, _GFM_N1451, _GFM_N1450, _GFM_N1447, _GFM_N1446, _GFM_N1444, _GFM_N1442, _GFM_N1441, _GFM_N1437, _GFM_N1436, _GFM_N1434, _GFM_N1433, _GFM_N1430, _GFM_N1429, _GFM_N1427, _GFM_N1423, _GFM_N1422, _GFM_N1420, _GFM_N1419, _GFM_N1416, _GFM_N1415, _GFM_N1413, _GFM_N1411, _GFM_N1410, _GFM_N1406, _GFM_N1405, _GFM_N1403, _GFM_N1402, _GFM_N1399, _GFM_N1398, _GFM_N1396, _GFM_N1392, 
  _GFM_N1391, _GFM_N1389, _GFM_N1388, _GFM_N1385, _GFM_N1384, _GFM_N1382, _GFM_N1380, _GFM_N1379, _GFM_N1375, _GFM_N1374, _GFM_N1372, _GFM_N1371, _GFM_N1368, _GFM_N1367, _GFM_N1365, _GFM_N1361, _GFM_N1360, _GFM_N1358, _GFM_N1357, _GFM_N1354, _GFM_N1353, _GFM_N1351, _GFM_N1349, _GFM_N1348, _GFM_N1344, _GFM_N1343, _GFM_N1341, _GFM_N1340, _GFM_N1337, _GFM_N1336, _GFM_N1334, _GFM_N1330, _GFM_N1329, _GFM_N1327, _GFM_N1326, _GFM_N1323, _GFM_N1322, _GFM_N1320, _GFM_N1318, _GFM_N1317, _GFM_N1313, _GFM_N1312, _GFM_N1310, _GFM_N1309, _GFM_N1306, _GFM_N1305, _GFM_N1303, _GFM_N1299, _GFM_N1298, _GFM_N1296, 
  _GFM_N1295, _GFM_N1292, _GFM_N1291, _GFM_N1289, _GFM_N1287, _GFM_N1286, _GFM_N1282, _GFM_N1281, _GFM_N1279, _GFM_N1278, _GFM_N1275, _GFM_N1274, _GFM_N1272, _GFM_N1268, _GFM_N1267, _GFM_N1265, _GFM_N1264, _GFM_N1261, _GFM_N1260, _GFM_N1258, _GFM_N1256, _GFM_N1255, _GFM_N1251, _GFM_N1250, _GFM_N1248, _GFM_N1247, _GFM_N1244, _GFM_N1243, _GFM_N1241, _GFM_N1237, _GFM_N1236, _GFM_N1234, _GFM_N1233, _GFM_N1230, _GFM_N1229, _GFM_N1227, _GFM_N1225, _GFM_N1224, _GFM_N1220, _GFM_N1219, _GFM_N1217, _GFM_N1216, _GFM_N1213, _GFM_N1212, _GFM_N1210, _GFM_N1206, _GFM_N1205, _GFM_N1203, _GFM_N1202, _GFM_N1199, 
  _GFM_N1198, _GFM_N1196, _GFM_N1194, _GFM_N1193, _GFM_N1189, _GFM_N1188, _GFM_N1186, _GFM_N1185, _GFM_N1182, _GFM_N1181, _GFM_N1179, _GFM_N1175, _GFM_N1174, _GFM_N1172, _GFM_N1171, _GFM_N1168, _GFM_N1167, _GFM_N1165, _GFM_N1163, _GFM_N1162, _GFM_N1158, _GFM_N1157, _GFM_N1155, _GFM_N1154, _GFM_N1151, _GFM_N1150, _GFM_N1148, _GFM_N1144, _GFM_N1143, _GFM_N1141, _GFM_N1140, _GFM_N1137, _GFM_N1136, _GFM_N1134, _GFM_N1132, _GFM_N1131, _GFM_N1127, _GFM_N1126, _GFM_N1124, _GFM_N1123, _GFM_N1120, _GFM_N1119, _GFM_N1117, _GFM_N1113, _GFM_N1112, _GFM_N1110, _GFM_N1109, _GFM_N1106, _GFM_N1105, _GFM_N1103, 
  _GFM_N1101, _GFM_N1100, _GFM_N1096, _GFM_N1095, _GFM_N1093, _GFM_N1092, _GFM_N1089, _GFM_N1088, _GFM_N1086, _GFM_N1082, _GFM_N1081, _GFM_N1079, _GFM_N1078, _GFM_N1075, _GFM_N1074, _GFM_N1072, _GFM_N1070, _GFM_N1069, _GFM_N1065, _GFM_N1064, _GFM_N1062, _GFM_N1061, _GFM_N1058, _GFM_N1057, _GFM_N1055, _GFM_N1051, _GFM_N1050, _GFM_N1048, _GFM_N1047, _GFM_N1044, _GFM_N1043, _GFM_N1041, _GFM_N1039, _GFM_N1038, _GFM_N1034, _GFM_N1033, _GFM_N1031, _GFM_N1030, _GFM_N1027, _GFM_N1026, _GFM_N1024, _GFM_N1020, _GFM_N1019, _GFM_N1017, _GFM_N1016, _GFM_N1013, _GFM_N1012, _GFM_N1010, _GFM_N1008, _GFM_N1007, 
  _GFM_N1003, _GFM_N1002, _GFM_N1000, _GFM_N999, _GFM_N996, _GFM_N995, _GFM_N993, _GFM_N989, _GFM_N988, _GFM_N986, _GFM_N985, _GFM_N982, _GFM_N981, _GFM_N979, _GFM_N977, _GFM_N976, _GFM_N972, _GFM_N971, _GFM_N969, _GFM_N968, _GFM_N965, _GFM_N964, _GFM_N962, _GFM_N958, _GFM_N957, _GFM_N955, _GFM_N954, _GFM_N951, _GFM_N950, _GFM_N948, _GFM_N946, _GFM_N945, _GFM_N941, _GFM_N940, _GFM_N938, _GFM_N937, _GFM_N934, _GFM_N933, _GFM_N931, _GFM_N927, _GFM_N926, _GFM_N924, _GFM_N923, _GFM_N920, _GFM_N919, _GFM_N917, _GFM_N915, _GFM_N914, _GFM_N910, _GFM_N909, 
  _GFM_N907, _GFM_N906, _GFM_N903, _GFM_N902, _GFM_N900, _GFM_N896, _GFM_N895, _GFM_N893, _GFM_N892, _GFM_N889, _GFM_N888, _GFM_N886, _GFM_N884, _GFM_N883, _GFM_N879, _GFM_N878, _GFM_N876, _GFM_N875, _GFM_N872, _GFM_N871, _GFM_N869, _GFM_N865, _GFM_N864, _GFM_N862, _GFM_N861, _GFM_N858, _GFM_N857, _GFM_N855, _GFM_N853, _GFM_N852, _GFM_N848, _GFM_N847, _GFM_N845, _GFM_N844, _GFM_N841, _GFM_N840, _GFM_N838, _GFM_N834, _GFM_N833, _GFM_N831, _GFM_N830, _GFM_N827, _GFM_N826, _GFM_N824, _GFM_N822, _GFM_N821, _GFM_N817, _GFM_N816, _GFM_N814, _GFM_N813, 
  _GFM_N810, _GFM_N809, _GFM_N807, _GFM_N803, _GFM_N802, _GFM_N800, _GFM_N799, _GFM_N796, _GFM_N795, _GFM_N793, _GFM_N791, _GFM_N790, _GFM_N786, _GFM_N785, _GFM_N783, _GFM_N782, _GFM_N779, _GFM_N778, _GFM_N776, _GFM_N772, _GFM_N771, _GFM_N769, _GFM_N768, _GFM_N765, _GFM_N764, _GFM_N762, _GFM_N760, _GFM_N759, _GFM_N755, _GFM_N754, _GFM_N752, _GFM_N751, _GFM_N748, _GFM_N747, _GFM_N745, _GFM_N741, _GFM_N740, _GFM_N738, _GFM_N737, _GFM_N734, _GFM_N733, _GFM_N731, _GFM_N729, _GFM_N728, _GFM_N724, _GFM_N723, _GFM_N721, _GFM_N720, _GFM_N717, _GFM_N716, 
  _GFM_N714, _GFM_N710, _GFM_N709, _GFM_N707, _GFM_N706, _GFM_N703, _GFM_N702, _GFM_N700, _GFM_N698, _GFM_N697, _GFM_N693, _GFM_N692, _GFM_N690, _GFM_N689, _GFM_N686, _GFM_N685, _GFM_N683, _GFM_N679, _GFM_N678, _GFM_N676, _GFM_N675, _GFM_N672, _GFM_N671, _GFM_N669, _GFM_N667, _GFM_N666, _GFM_N662, _GFM_N661, _GFM_N659, _GFM_N658, _GFM_N655, _GFM_N654, _GFM_N652, _GFM_N648, _GFM_N647, _GFM_N645, _GFM_N644, _GFM_N641, _GFM_N640, _GFM_N638, _GFM_N636, _GFM_N635, _GFM_N631, _GFM_N630, _GFM_N628, _GFM_N627, _GFM_N624, _GFM_N623, _GFM_N621, _GFM_N617, 
  _GFM_N616, _GFM_N614, _GFM_N613, _GFM_N610, _GFM_N609, _GFM_N607, _GFM_N605, _GFM_N604, _GFM_N600, _GFM_N599, _GFM_N597, _GFM_N596, _GFM_N593, _GFM_N592, _GFM_N590, _GFM_N586, _GFM_N585, _GFM_N583, _GFM_N582, _GFM_N579, _GFM_N578, _GFM_N576, _GFM_N574, _GFM_N573, _GFM_N569, _GFM_N568, _GFM_N566, _GFM_N565, _GFM_N562, _GFM_N561, _GFM_N559, _GFM_N555, _GFM_N554, _GFM_N552, _GFM_N551, _GFM_N548, _GFM_N547, _GFM_N545, _GFM_N543, _GFM_N542, _GFM_N538, _GFM_N537, _GFM_N535, _GFM_N534, _GFM_N531, _GFM_N530, _GFM_N528, _GFM_N524, _GFM_N523, _GFM_N521, 
  _GFM_N520, _GFM_N517, _GFM_N516, _GFM_N514, _GFM_N512, _GFM_N511, _GFM_N507, _GFM_N506, _GFM_N504, _GFM_N503, _GFM_N500, _GFM_N499, _GFM_N497, _GFM_N493, _GFM_N492, _GFM_N490, _GFM_N489, _GFM_N486, _GFM_N485, _GFM_N483, _GFM_N481, _GFM_N480, _GFM_N476, _GFM_N475, _GFM_N473, _GFM_N472, _GFM_N469, _GFM_N468, _GFM_N466, _GFM_N462, _GFM_N461, _GFM_N459, _GFM_N458, _GFM_N455, _GFM_N454, _GFM_N452, _GFM_N450, _GFM_N449, _GFM_N445, _GFM_N444, _GFM_N442, _GFM_N441, _GFM_N438, _GFM_N437, _GFM_N435, _GFM_N431, _GFM_N430, _GFM_N428, _GFM_N427, _GFM_N424, 
  _GFM_N423, _GFM_N421, _GFM_N419, _GFM_N418, _GFM_N414, _GFM_N413, _GFM_N411, _GFM_N410, _GFM_N407, _GFM_N406, _GFM_N404, _GFM_N400, _GFM_N399, _GFM_N397, _GFM_N396, _GFM_N393, _GFM_N392, _GFM_N390, _GFM_N388, _GFM_N387, _GFM_N383, _GFM_N382, _GFM_N380, _GFM_N379, _GFM_N376, _GFM_N375, _GFM_N373, _GFM_N369, _GFM_N368, _GFM_N366, _GFM_N365, _GFM_N362, _GFM_N361, _GFM_N359, _GFM_N357, _GFM_N356, _GFM_N352, _GFM_N351, _GFM_N349, _GFM_N348, _GFM_N345, _GFM_N344, _GFM_N342, _GFM_N338, _GFM_N337, _GFM_N335, _GFM_N334, _GFM_N331, _GFM_N330, _GFM_N328, 
  _GFM_N326, _GFM_N325, _GFM_N321, _GFM_N320, _GFM_N318, _GFM_N317, _GFM_N314, _GFM_N313, _GFM_N311, _GFM_N307, _GFM_N306, _GFM_N304, _GFM_N303, _GFM_N300, _GFM_N299, _GFM_N297, _GFM_N295, _GFM_N294, _GFM_N290, _GFM_N289, _GFM_N287, _GFM_N286, _GFM_N283, _GFM_N282, _GFM_N280, _GFM_N276, _GFM_N275, _GFM_N273, _GFM_N272, _GFM_N269, _GFM_N268, _GFM_N266, _GFM_N264, _GFM_N263, _GFM_N259, _GFM_N258, _GFM_N256, _GFM_N255, _GFM_N252, _GFM_N251, _GFM_N249, _GFM_N245, _GFM_N244, _GFM_N242, _GFM_N241, _GFM_N238, _GFM_N237, _GFM_N235, _GFM_N233, _GFM_N232, 
  _GFM_N228, _GFM_N227, _GFM_N225, _GFM_N224, _GFM_N221, _GFM_N220, _GFM_N218, _GFM_N214, _GFM_N213, _GFM_N211, _GFM_N210, _GFM_N207, _GFM_N206, _GFM_N204, _GFM_N202, _GFM_N201, _GFM_N197, _GFM_N196, _GFM_N194, _GFM_N193, _GFM_N190, _GFM_N189, _GFM_N187, _GFM_N183, _GFM_N182, _GFM_N180, _GFM_N179, _GFM_N176, _GFM_N175, _GFM_N173, _GFM_N171, _GFM_N170, _GFM_N166, _GFM_N165, _GFM_N163, _GFM_N162, _GFM_N159, _GFM_N158, _GFM_N156, _GFM_N152, _GFM_N151, _GFM_N149, _GFM_N148, _GFM_N145, _GFM_N144, _GFM_N142, _GFM_N140, _GFM_N139, _GFM_N135, _GFM_N134, 
  _GFM_N132, _GFM_N131, _GFM_N128, _GFM_N127, _GFM_N125, _GFM_N121, _GFM_N120, _GFM_N118, _GFM_N117, _GFM_N114, _GFM_N113, _GFM_N111, _GFM_N109, _GFM_N108, _GFM_N104, _GFM_N103, _GFM_N101, _GFM_N100, _GFM_N97, _GFM_N96, _GFM_N94, _GFM_N90, _GFM_N89, _GFM_N87, _GFM_N86, _GFM_N83, _GFM_N82, _GFM_N80, _GFM_N78, _GFM_N77, _GFM_N73, _GFM_N72, _GFM_N70, _GFM_N69, _GFM_N66, _GFM_N65, _GFM_N63, _GFM_N59, _GFM_N58, _GFM_N56, _GFM_N55, _GFM_N52, _GFM_N51, _GFM_N49, _GFM_N47, _GFM_N46, _GFM_N42, _GFM_N41, _GFM_N39, _GFM_N38, 
  _GFM_N35, _GFM_N34, _GFM_N32, _GFM_N28, _GFM_N27, _GFM_N25, _GFM_N24, _GFM_N21, _GFM_N20, _GFM_N18, _GFM_N16, _GFM_N15, _GFM_N11, _GFM_N10, _GFM_N8, _GFM_N7, _GFM_N4, _GFM_N3, _GFM_N1, _AES_ENC_n1267, _AES_ENC_n1266, _AES_ENC_n1265, _AES_ENC_n1264, _AES_ENC_n1263, _AES_ENC_n1262, _AES_ENC_n1261, _AES_ENC_n12601, _AES_ENC_n1259, _AES_ENC_n1258, _AES_ENC_n1257, _AES_ENC_n1256, _AES_ENC_n1255, _AES_ENC_n1254, _AES_ENC_n1253, _AES_ENC_n1252, _AES_ENC_n1251, _AES_ENC_n1250, _AES_ENC_n1249, _AES_ENC_n1248, _AES_ENC_n1247, _AES_ENC_n1246, _AES_ENC_n1245, _AES_ENC_n1244, _AES_ENC_n1243, _AES_ENC_n1242, _AES_ENC_n1241, _AES_ENC_n1240, _AES_ENC_n1239, _AES_ENC_n1238, _AES_ENC_n1237, 
  _AES_ENC_n1236, _AES_ENC_n1235, _AES_ENC_n1234, _AES_ENC_n1233, _AES_ENC_n1232, _AES_ENC_n1231, _AES_ENC_n793, _AES_ENC_n794, _AES_ENC_n792, _AES_ENC_n791, _AES_ENC_n7901, _AES_ENC_n7891, _AES_ENC_n6601, _AES_ENC_n659, _AES_ENC_n658, _AES_ENC_n657, _AES_ENC_n656, _AES_ENC_n655, _AES_ENC_n654, _AES_ENC_n653, _AES_ENC_n652, _AES_ENC_n651, _AES_ENC_n6501, _AES_ENC_n649, _AES_ENC_n648, _AES_ENC_n647, _AES_ENC_n646, _AES_ENC_n645, _AES_ENC_n644, _AES_ENC_n643, _AES_ENC_n642, _AES_ENC_n641, _AES_ENC_n6401, _AES_ENC_n639, _AES_ENC_n638, _AES_ENC_n637, _AES_ENC_n636, _AES_ENC_n635, _AES_ENC_n634, _AES_ENC_n633, _AES_ENC_n632, _AES_ENC_n631, _AES_ENC_n6301, _AES_ENC_n629, _AES_ENC_n628, _AES_ENC_n627, _AES_ENC_n626, _AES_ENC_n625, _AES_ENC_n624, _AES_ENC_n623, 
  _AES_ENC_n622, _AES_ENC_n621, _AES_ENC_n6201, _AES_ENC_n619, _AES_ENC_n618, _AES_ENC_n617, _AES_ENC_n616, _AES_ENC_n615, _AES_ENC_n614, _AES_ENC_n613, _AES_ENC_n612, _AES_ENC_n611, _AES_ENC_n610, _AES_ENC_n609, _AES_ENC_n608, _AES_ENC_n607, _AES_ENC_n606, _AES_ENC_n605, _AES_ENC_n604, _AES_ENC_n603, _AES_ENC_n602, _AES_ENC_n601, _AES_ENC_n600, _AES_ENC_n599, _AES_ENC_n598, _AES_ENC_n597, _AES_ENC_n596, _AES_ENC_n595, _AES_ENC_n594, _AES_ENC_n593, _AES_ENC_n592, _AES_ENC_n591, _AES_ENC_n590, _AES_ENC_n589, _AES_ENC_n588, _AES_ENC_n587, _AES_ENC_n586, _AES_ENC_n585, _AES_ENC_n584, _AES_ENC_n583, _AES_ENC_n582, _AES_ENC_n581, _AES_ENC_n580, _AES_ENC_n579, _AES_ENC_n578, _AES_ENC_n577, _AES_ENC_n576, _AES_ENC_n575, _AES_ENC_n574, _AES_ENC_n573, 
  _AES_ENC_n572, _AES_ENC_n571, _AES_ENC_n570, _AES_ENC_n569, _AES_ENC_n568, _AES_ENC_n567, _AES_ENC_n566, _AES_ENC_n565, _AES_ENC_n564, _AES_ENC_n563, _AES_ENC_n562, _AES_ENC_n561, _AES_ENC_n560, _AES_ENC_n559, _AES_ENC_n558, _AES_ENC_n557, _AES_ENC_n556, _AES_ENC_n555, _AES_ENC_n554, _AES_ENC_n553, _AES_ENC_n552, _AES_ENC_n551, _AES_ENC_n550, _AES_ENC_n549, _AES_ENC_n548, _AES_ENC_n547, _AES_ENC_n546, _AES_ENC_n545, _AES_ENC_n544, _AES_ENC_n543, _AES_ENC_n542, _AES_ENC_n541, _AES_ENC_n540, _AES_ENC_n539, _AES_ENC_n538, _AES_ENC_n537, _AES_ENC_n536, _AES_ENC_n535, _AES_ENC_n534, _AES_ENC_n533, _AES_ENC_n532, _AES_ENC_n531, _AES_ENC_n5301, _AES_ENC_n529, _AES_ENC_n528, _AES_ENC_n527, _AES_ENC_n526, _AES_ENC_n525, _AES_ENC_n524, _AES_ENC_n523, 
  _AES_ENC_n522, _AES_ENC_n521, _AES_ENC_n5201, _AES_ENC_n519, _AES_ENC_n518, _AES_ENC_n517, _AES_ENC_n516, _AES_ENC_n515, _AES_ENC_n514, _AES_ENC_n513, _AES_ENC_n512, _AES_ENC_n511, _AES_ENC_n5101, _AES_ENC_n509, _AES_ENC_n508, _AES_ENC_n507, _AES_ENC_n506, _AES_ENC_n505, _AES_ENC_n504, _AES_ENC_n503, _AES_ENC_n5021, _AES_ENC_n5010, _AES_ENC_n5000, _AES_ENC_n4990, _AES_ENC_n4980, _AES_ENC_n4970, _AES_ENC_n4960, _AES_ENC_n4950, _AES_ENC_n4940, _AES_ENC_n4930, _AES_ENC_n4920, _AES_ENC_n4911, _AES_ENC_n4900, _AES_ENC_n4890, _AES_ENC_n4880, _AES_ENC_n4870, _AES_ENC_n4860, _AES_ENC_n4850, _AES_ENC_n4840, _AES_ENC_n4830, _AES_ENC_n4820, _AES_ENC_n4811, _AES_ENC_n4800, _AES_ENC_n4790, _AES_ENC_n4780, _AES_ENC_n4770, _AES_ENC_n4760, _AES_ENC_n4750, _AES_ENC_n4740, _AES_ENC_n4730, 
  _AES_ENC_n4720, _AES_ENC_n4711, _AES_ENC_n4700, _AES_ENC_n4690, _AES_ENC_n4680, _AES_ENC_n4670, _AES_ENC_n4660, _AES_ENC_n4650, _AES_ENC_n4640, _AES_ENC_n4630, _AES_ENC_n4620, _AES_ENC_n4611, _AES_ENC_n4600, _AES_ENC_n4590, _AES_ENC_n4580, _AES_ENC_n4570, _AES_ENC_n4560, _AES_ENC_n4550, _AES_ENC_n4540, _AES_ENC_n4530, _AES_ENC_n4520, _AES_ENC_n4510, _AES_ENC_n4500, _AES_ENC_n4490, _AES_ENC_n4480, _AES_ENC_n4470, _AES_ENC_n4460, _AES_ENC_n4450, _AES_ENC_n4440, _AES_ENC_n4430, _AES_ENC_n4420, _AES_ENC_n4410, _AES_ENC_n4400, _AES_ENC_n4390, _AES_ENC_n4380, _AES_ENC_n4370, _AES_ENC_n4360, _AES_ENC_n4350, _AES_ENC_n4340, _AES_ENC_n4330, _AES_ENC_n4320, _AES_ENC_n4310, _AES_ENC_n4300, _AES_ENC_n4290, _AES_ENC_n4280, _AES_ENC_n4270, _AES_ENC_n4260, _AES_ENC_n4250, _AES_ENC_n4240, _AES_ENC_n4230, 
  _AES_ENC_n4220, _AES_ENC_n4210, _AES_ENC_n4200, _AES_ENC_n4190, _AES_ENC_n4180, _AES_ENC_n4170, _AES_ENC_n4160, _AES_ENC_n4150, _AES_ENC_n4140, _AES_ENC_n4130, _AES_ENC_n4120, _AES_ENC_n4110, _AES_ENC_n4100, _AES_ENC_n4090, _AES_ENC_n4080, _AES_ENC_n4070, _AES_ENC_n4060, _AES_ENC_n4050, _AES_ENC_n4040, _AES_ENC_n4030, _AES_ENC_n4020, _AES_ENC_n4010, _AES_ENC_n4000, _AES_ENC_n3990, _AES_ENC_n3980, _AES_ENC_n3970, _AES_ENC_n3960, _AES_ENC_n3950, _AES_ENC_n3940, _AES_ENC_n3930, _AES_ENC_n3920, _AES_ENC_n3910, _AES_ENC_n3900, _AES_ENC_n3890, _AES_ENC_n3880, _AES_ENC_n3870, _AES_ENC_n3860, _AES_ENC_n3850, _AES_ENC_n3840, _AES_ENC_n3830, _AES_ENC_n3820, _AES_ENC_n3810, _AES_ENC_n3800, _AES_ENC_n3790, _AES_ENC_n3780, _AES_ENC_n3770, _AES_ENC_n3760, _AES_ENC_n3750, _AES_ENC_n3740, _AES_ENC_n373, 
  _AES_ENC_n372, _AES_ENC_n371, _AES_ENC_n3701, _AES_ENC_n369, _AES_ENC_n368, _AES_ENC_n367, _AES_ENC_n366, _AES_ENC_n365, _AES_ENC_n364, _AES_ENC_n363, _AES_ENC_n362, _AES_ENC_n361, _AES_ENC_n3601, _AES_ENC_n359, _AES_ENC_n358, _AES_ENC_n357, _AES_ENC_n356, _AES_ENC_n355, _AES_ENC_n354, _AES_ENC_n353, _AES_ENC_n352, _AES_ENC_n351, _AES_ENC_n3501, _AES_ENC_n349, _AES_ENC_n348, _AES_ENC_n347, _AES_ENC_n346, _AES_ENC_n345, _AES_ENC_n344, _AES_ENC_n343, _AES_ENC_n342, _AES_ENC_n341, _AES_ENC_n3401, _AES_ENC_n339, _AES_ENC_n338, _AES_ENC_n337, _AES_ENC_n336, _AES_ENC_n335, _AES_ENC_n334, _AES_ENC_n333, _AES_ENC_n332, _AES_ENC_n331, _AES_ENC_n3301, _AES_ENC_n329, _AES_ENC_n328, _AES_ENC_n327, _AES_ENC_n326, _AES_ENC_n325, _AES_ENC_n324, _AES_ENC_n323, 
  _AES_ENC_n322, _AES_ENC_n321, _AES_ENC_n3201, _AES_ENC_n319, _AES_ENC_n318, _AES_ENC_n317, _AES_ENC_n316, _AES_ENC_n315, _AES_ENC_n314, _AES_ENC_n313, _AES_ENC_n312, _AES_ENC_n311, _AES_ENC_n3101, _AES_ENC_n309, _AES_ENC_n308, _AES_ENC_n307, _AES_ENC_n306, _AES_ENC_n305, _AES_ENC_n304, _AES_ENC_n303, _AES_ENC_n302, _AES_ENC_n301, _AES_ENC_n3001, _AES_ENC_n299, _AES_ENC_n298, _AES_ENC_n297, _AES_ENC_n296, _AES_ENC_n295, _AES_ENC_n294, _AES_ENC_n293, _AES_ENC_n292, _AES_ENC_n291, _AES_ENC_n290, _AES_ENC_n289, _AES_ENC_n288, _AES_ENC_n287, _AES_ENC_n286, _AES_ENC_n285, _AES_ENC_n284, _AES_ENC_n283, _AES_ENC_n282, _AES_ENC_n281, _AES_ENC_n280, _AES_ENC_n279, _AES_ENC_n278, _AES_ENC_n2770, _AES_ENC_n2760, _AES_ENC_n2750, _AES_ENC_n2740, _AES_ENC_n2730, 
  _AES_ENC_n2720, _AES_ENC_n2710, _AES_ENC_n2700, _AES_ENC_n269, _AES_ENC_n268, _AES_ENC_n267, _AES_ENC_n266, _AES_ENC_n265, _AES_ENC_n264, _AES_ENC_n263, _AES_ENC_n262, _AES_ENC_n2610, _AES_ENC_n2600, _AES_ENC_n2590, _AES_ENC_n2580, _AES_ENC_n2570, _AES_ENC_n2560, _AES_ENC_n2550, _AES_ENC_n2540, _AES_ENC_n253, _AES_ENC_n252, _AES_ENC_n251, _AES_ENC_n250, _AES_ENC_n249, _AES_ENC_n248, _AES_ENC_n247, _AES_ENC_n246, _AES_ENC_n2450, _AES_ENC_n2440, _AES_ENC_n2430, _AES_ENC_n2420, _AES_ENC_n2410, _AES_ENC_n2400, _AES_ENC_n2390, _AES_ENC_n2380, _AES_ENC_n237, _AES_ENC_n236, _AES_ENC_n235, _AES_ENC_n234, _AES_ENC_n233, _AES_ENC_n232, _AES_ENC_n231, _AES_ENC_n230, _AES_ENC_n2290, _AES_ENC_n2280, _AES_ENC_n2270, _AES_ENC_n2260, _AES_ENC_n2250, _AES_ENC_n2240, _AES_ENC_n2230, 
  _AES_ENC_n2220, _AES_ENC_n221, _AES_ENC_n220, _AES_ENC_n219, _AES_ENC_n218, _AES_ENC_n217, _AES_ENC_n216, _AES_ENC_n215, _AES_ENC_n214, _AES_ENC_n2130, _AES_ENC_n2120, _AES_ENC_n2110, _AES_ENC_n2100, _AES_ENC_n2090, _AES_ENC_n2080, _AES_ENC_n2070, _AES_ENC_n2060, _AES_ENC_n205, _AES_ENC_n204, _AES_ENC_n203, _AES_ENC_n202, _AES_ENC_n201, _AES_ENC_n200, _AES_ENC_n199, _AES_ENC_n1981, _AES_ENC_n1970, _AES_ENC_n1960, _AES_ENC_n1950, _AES_ENC_n1940, _AES_ENC_n1930, _AES_ENC_n1920, _AES_ENC_n1910, _AES_ENC_n1900, _AES_ENC_n189, _AES_ENC_n188, _AES_ENC_n187, _AES_ENC_n186, _AES_ENC_n185, _AES_ENC_n184, _AES_ENC_n183, _AES_ENC_n182, _AES_ENC_n1810, _AES_ENC_n1800, _AES_ENC_n1790, _AES_ENC_n1780, _AES_ENC_n1770, _AES_ENC_n1760, _AES_ENC_n1750, _AES_ENC_n1740, _AES_ENC_n173, 
  _AES_ENC_n172, _AES_ENC_n171, _AES_ENC_n170, _AES_ENC_n169, _AES_ENC_n168, _AES_ENC_n167, _AES_ENC_n166, _AES_ENC_n1650, _AES_ENC_n1640, _AES_ENC_n1630, _AES_ENC_n1620, _AES_ENC_n1610, _AES_ENC_n1600, _AES_ENC_n1590, _AES_ENC_n1580, _AES_ENC_n157, _AES_ENC_n156, _AES_ENC_n155, _AES_ENC_n154, _AES_ENC_n153, _AES_ENC_n152, _AES_ENC_n151, _AES_ENC_n150, _AES_ENC_n1490, _AES_ENC_n1480, _AES_ENC_n1470, _AES_ENC_n1460, _AES_ENC_n1450, _AES_ENC_n1440, _AES_ENC_n1430, _AES_ENC_n1420, _AES_ENC_n141, _AES_ENC_n140, _AES_ENC_n139, _AES_ENC_n138, _AES_ENC_n137, _AES_ENC_n136, _AES_ENC_n135, _AES_ENC_n134, _AES_ENC_n1330, _AES_ENC_n1320, _AES_ENC_n1310, _AES_ENC_n1300, _AES_ENC_n1290, _AES_ENC_n1280, _AES_ENC_n1270, _AES_ENC_n12600, _AES_ENC_n125, _AES_ENC_n124, _AES_ENC_n123, 
  _AES_ENC_n122, _AES_ENC_n121, _AES_ENC_n120, _AES_ENC_n119, _AES_ENC_n118, _AES_ENC_n11710, _AES_ENC_n11610, _AES_ENC_n11510, _AES_ENC_n11410, _AES_ENC_n11310, _AES_ENC_n11210, _AES_ENC_n11110, _AES_ENC_n11010, _AES_ENC_n109, _AES_ENC_n108, _AES_ENC_n107, _AES_ENC_n106, _AES_ENC_n105, _AES_ENC_n104, _AES_ENC_n103, _AES_ENC_n102, _AES_ENC_n10110, _AES_ENC_n10010, _AES_ENC_n9910, _AES_ENC_n9810, _AES_ENC_n9710, _AES_ENC_n9610, _AES_ENC_n9510, _AES_ENC_n9410, _AES_ENC_n93, _AES_ENC_n92, _AES_ENC_n91, _AES_ENC_n90, _AES_ENC_n89, _AES_ENC_n88, _AES_ENC_n87, _AES_ENC_n86, _AES_ENC_n8510, _AES_ENC_n8410, _AES_ENC_n8310, _AES_ENC_n8210, _AES_ENC_n8110, _AES_ENC_n8010, _AES_ENC_n7900, _AES_ENC_n7890, _AES_ENC_n77, _AES_ENC_n76, _AES_ENC_n75, _AES_ENC_n74, _AES_ENC_n73, 
  _AES_ENC_n72, _AES_ENC_n71, _AES_ENC_n70, _AES_ENC_n6910, _AES_ENC_n6810, _AES_ENC_n6710, _AES_ENC_n6600, _AES_ENC_n6500, _AES_ENC_n6400, _AES_ENC_n6300, _AES_ENC_n6200, _AES_ENC_n61, _AES_ENC_n60, _AES_ENC_n59, _AES_ENC_n58, _AES_ENC_n57, _AES_ENC_n56, _AES_ENC_n55, _AES_ENC_n54, _AES_ENC_n5300, _AES_ENC_n5200, _AES_ENC_n5100, _AES_ENC_n5020, _AES_ENC_n4910, _AES_ENC_n4810, _AES_ENC_n4710, _AES_ENC_n4610, _AES_ENC_n45, _AES_ENC_n44, _AES_ENC_n43, _AES_ENC_n42, _AES_ENC_n41, _AES_ENC_n40, _AES_ENC_n39, _AES_ENC_n38, _AES_ENC_n3700, _AES_ENC_n3600, _AES_ENC_n3500, _AES_ENC_n3400, _AES_ENC_n3300, _AES_ENC_n3200, _AES_ENC_n3100, _AES_ENC_n3000, _AES_ENC_n29, _AES_ENC_n28, _AES_ENC_n27, _AES_ENC_n26, _AES_ENC_n25, _AES_ENC_n24, _AES_ENC_n23, 
  _AES_ENC_n22, _AES_ENC_n21, _AES_ENC_n20, _AES_ENC_n1980, _AES_ENC_n18, _AES_ENC_n17, _AES_ENC_n16, _AES_ENC_n15, _AES_ENC_n14, _AES_ENC_n13, _AES_ENC_n12, _AES_ENC_n11, _AES_ENC_n2, _AES_ENC_n1230, _AES_ENC_n1229, _AES_ENC_n1228, _AES_ENC_n1227, _AES_ENC_n1226, _AES_ENC_n1225, _AES_ENC_n1224, _AES_ENC_n1223, _AES_ENC_n1222, _AES_ENC_n1221, _AES_ENC_n1220, _AES_ENC_n1219, _AES_ENC_n1218, _AES_ENC_n1217, _AES_ENC_n1216, _AES_ENC_n1215, _AES_ENC_n1214, _AES_ENC_n1213, _AES_ENC_n1212, _AES_ENC_n1211, _AES_ENC_n1210, _AES_ENC_n1209, _AES_ENC_n1208, _AES_ENC_n1207, _AES_ENC_n1206, _AES_ENC_n1205, _AES_ENC_n1204, _AES_ENC_n1203, _AES_ENC_n1202, _AES_ENC_n1201, _AES_ENC_n1200, _AES_ENC_n1199, _AES_ENC_n1198, _AES_ENC_n1197, _AES_ENC_n1196, _AES_ENC_n1195, _AES_ENC_n1194, 
  _AES_ENC_n1193, _AES_ENC_n1192, _AES_ENC_n1191, _AES_ENC_n1190, _AES_ENC_n1189, _AES_ENC_n1188, _AES_ENC_n1187, _AES_ENC_n1186, _AES_ENC_n1185, _AES_ENC_n1184, _AES_ENC_n1183, _AES_ENC_n1182, _AES_ENC_n1181, _AES_ENC_n1180, _AES_ENC_n1179, _AES_ENC_n1178, _AES_ENC_n1177, _AES_ENC_n1176, _AES_ENC_n1175, _AES_ENC_n1174, _AES_ENC_n1173, _AES_ENC_n1172, _AES_ENC_n1171, _AES_ENC_n1170, _AES_ENC_n1169, _AES_ENC_n1168, _AES_ENC_n1167, _AES_ENC_n1166, _AES_ENC_n1165, _AES_ENC_n1164, _AES_ENC_n1163, _AES_ENC_n1162, _AES_ENC_n1161, _AES_ENC_n1160, _AES_ENC_n1159, _AES_ENC_n1158, _AES_ENC_n1157, _AES_ENC_n1156, _AES_ENC_n1155, _AES_ENC_n1154, _AES_ENC_n1153, _AES_ENC_n1152, _AES_ENC_n1151, _AES_ENC_n1150, _AES_ENC_n1149, _AES_ENC_n1148, _AES_ENC_n1147, _AES_ENC_n1146, _AES_ENC_n1145, _AES_ENC_n1144, 
  _AES_ENC_n1143, _AES_ENC_n1142, _AES_ENC_n1141, _AES_ENC_n1140, _AES_ENC_n1139, _AES_ENC_n1138, _AES_ENC_n1137, _AES_ENC_n1136, _AES_ENC_n1135, _AES_ENC_n1134, _AES_ENC_n1133, _AES_ENC_n1132, _AES_ENC_n1131, _AES_ENC_n1130, _AES_ENC_n1129, _AES_ENC_n1128, _AES_ENC_n1127, _AES_ENC_n1126, _AES_ENC_n1125, _AES_ENC_n1124, _AES_ENC_n1123, _AES_ENC_n1122, _AES_ENC_n1121, _AES_ENC_n1120, _AES_ENC_n1119, _AES_ENC_n1118, _AES_ENC_n1117, _AES_ENC_n1116, _AES_ENC_n1115, _AES_ENC_n1114, _AES_ENC_n1113, _AES_ENC_n1112, _AES_ENC_n1111, _AES_ENC_n1110, _AES_ENC_n1109, _AES_ENC_n1108, _AES_ENC_n1107, _AES_ENC_n1106, _AES_ENC_n1105, _AES_ENC_n1104, _AES_ENC_n1103, _AES_ENC_n1102, _AES_ENC_n1101, _AES_ENC_n1100, _AES_ENC_n1099, _AES_ENC_n1098, _AES_ENC_n1097, _AES_ENC_n1096, _AES_ENC_n1095, _AES_ENC_n1094, 
  _AES_ENC_n1093, _AES_ENC_n1092, _AES_ENC_n1091, _AES_ENC_n1090, _AES_ENC_n1089, _AES_ENC_n1088, _AES_ENC_n1087, _AES_ENC_n1086, _AES_ENC_n1085, _AES_ENC_n1084, _AES_ENC_n1083, _AES_ENC_n1082, _AES_ENC_n1081, _AES_ENC_n1080, _AES_ENC_n1079, _AES_ENC_n1078, _AES_ENC_n1077, _AES_ENC_n1076, _AES_ENC_n1075, _AES_ENC_n1074, _AES_ENC_n1073, _AES_ENC_n1072, _AES_ENC_n1071, _AES_ENC_n1070, _AES_ENC_n1069, _AES_ENC_n1068, _AES_ENC_n1067, _AES_ENC_n1066, _AES_ENC_n1065, _AES_ENC_n1064, _AES_ENC_n1063, _AES_ENC_n1062, _AES_ENC_n1061, _AES_ENC_n1060, _AES_ENC_n1059, _AES_ENC_n1058, _AES_ENC_n1057, _AES_ENC_n1056, _AES_ENC_n1055, _AES_ENC_n1054, _AES_ENC_n1053, _AES_ENC_n1052, _AES_ENC_n1051, _AES_ENC_n1050, _AES_ENC_n1049, _AES_ENC_n1048, _AES_ENC_n1047, _AES_ENC_n1046, _AES_ENC_n1045, _AES_ENC_n1044, 
  _AES_ENC_n1043, _AES_ENC_n1042, _AES_ENC_n1041, _AES_ENC_n1040, _AES_ENC_n1039, _AES_ENC_n1038, _AES_ENC_n1037, _AES_ENC_n1036, _AES_ENC_n1035, _AES_ENC_n1034, _AES_ENC_n1033, _AES_ENC_n1032, _AES_ENC_n1031, _AES_ENC_n1030, _AES_ENC_n1029, _AES_ENC_n1028, _AES_ENC_n1027, _AES_ENC_n1026, _AES_ENC_n1025, _AES_ENC_n1024, _AES_ENC_n1023, _AES_ENC_n1022, _AES_ENC_n1021, _AES_ENC_n1020, _AES_ENC_n1019, _AES_ENC_n1018, _AES_ENC_n1017, _AES_ENC_n1016, _AES_ENC_n1015, _AES_ENC_n1014, _AES_ENC_n1013, _AES_ENC_n1012, _AES_ENC_n1011, _AES_ENC_n1010, _AES_ENC_n1009, _AES_ENC_n1008, _AES_ENC_n1007, _AES_ENC_n1006, _AES_ENC_n1005, _AES_ENC_n1004, _AES_ENC_n1003, _AES_ENC_n1002, _AES_ENC_n1001, _AES_ENC_n1000, _AES_ENC_n999, _AES_ENC_n998, _AES_ENC_n997, _AES_ENC_n996, _AES_ENC_n995, _AES_ENC_n994, 
  _AES_ENC_n993, _AES_ENC_n992, _AES_ENC_n991, _AES_ENC_n990, _AES_ENC_n989, _AES_ENC_n988, _AES_ENC_n987, _AES_ENC_n986, _AES_ENC_n985, _AES_ENC_n984, _AES_ENC_n983, _AES_ENC_n982, _AES_ENC_n981, _AES_ENC_n980, _AES_ENC_n979, _AES_ENC_n978, _AES_ENC_n977, _AES_ENC_n976, _AES_ENC_n975, _AES_ENC_n974, _AES_ENC_n973, _AES_ENC_n972, _AES_ENC_n971, _AES_ENC_n970, _AES_ENC_n969, _AES_ENC_n968, _AES_ENC_n967, _AES_ENC_n966, _AES_ENC_n965, _AES_ENC_n964, _AES_ENC_n963, _AES_ENC_n962, _AES_ENC_n961, _AES_ENC_n960, _AES_ENC_n959, _AES_ENC_n958, _AES_ENC_n957, _AES_ENC_n956, _AES_ENC_n955, _AES_ENC_n954, _AES_ENC_n953, _AES_ENC_n952, _AES_ENC_n951, _AES_ENC_n950, _AES_ENC_n949, _AES_ENC_n948, _AES_ENC_n947, _AES_ENC_n946, _AES_ENC_n945, _AES_ENC_n944, 
  _AES_ENC_n943, _AES_ENC_n942, _AES_ENC_n941, _AES_ENC_n940, _AES_ENC_n939, _AES_ENC_n938, _AES_ENC_n937, _AES_ENC_n936, _AES_ENC_n935, _AES_ENC_n934, _AES_ENC_n933, _AES_ENC_n932, _AES_ENC_n931, _AES_ENC_n930, _AES_ENC_n929, _AES_ENC_n928, _AES_ENC_n927, _AES_ENC_n926, _AES_ENC_n925, _AES_ENC_n924, _AES_ENC_n923, _AES_ENC_n922, _AES_ENC_n921, _AES_ENC_n920, _AES_ENC_n919, _AES_ENC_n918, _AES_ENC_n917, _AES_ENC_n916, _AES_ENC_n915, _AES_ENC_n914, _AES_ENC_n913, _AES_ENC_n912, _AES_ENC_n911, _AES_ENC_n910, _AES_ENC_n909, _AES_ENC_n908, _AES_ENC_n907, _AES_ENC_n906, _AES_ENC_n905, _AES_ENC_n904, _AES_ENC_n903, _AES_ENC_n902, _AES_ENC_n901, _AES_ENC_n900, _AES_ENC_n899, _AES_ENC_n898, _AES_ENC_n897, _AES_ENC_n896, _AES_ENC_n895, _AES_ENC_n894, 
  _AES_ENC_n893, _AES_ENC_n892, _AES_ENC_n891, _AES_ENC_n890, _AES_ENC_n889, _AES_ENC_n888, _AES_ENC_n887, _AES_ENC_n886, _AES_ENC_n885, _AES_ENC_n884, _AES_ENC_n883, _AES_ENC_n882, _AES_ENC_n881, _AES_ENC_n880, _AES_ENC_n879, _AES_ENC_n878, _AES_ENC_n877, _AES_ENC_n876, _AES_ENC_n875, _AES_ENC_n874, _AES_ENC_n873, _AES_ENC_n872, _AES_ENC_n871, _AES_ENC_n870, _AES_ENC_n869, _AES_ENC_n868, _AES_ENC_n867, _AES_ENC_n866, _AES_ENC_n865, _AES_ENC_n864, _AES_ENC_n863, _AES_ENC_n862, _AES_ENC_n861, _AES_ENC_n860, _AES_ENC_n859, _AES_ENC_n858, _AES_ENC_n857, _AES_ENC_n856, _AES_ENC_n855, _AES_ENC_n854, _AES_ENC_n853, _AES_ENC_n852, _AES_ENC_n851, _AES_ENC_n850, _AES_ENC_n849, _AES_ENC_n848, _AES_ENC_n847, _AES_ENC_n846, _AES_ENC_n845, _AES_ENC_n844, 
  _AES_ENC_n843, _AES_ENC_n842, _AES_ENC_n841, _AES_ENC_n840, _AES_ENC_n839, _AES_ENC_n838, _AES_ENC_n837, _AES_ENC_n836, _AES_ENC_n835, _AES_ENC_n834, _AES_ENC_n833, _AES_ENC_n832, _AES_ENC_n831, _AES_ENC_n830, _AES_ENC_n829, _AES_ENC_n828, _AES_ENC_n827, _AES_ENC_n826, _AES_ENC_n825, _AES_ENC_n824, _AES_ENC_n823, _AES_ENC_n822, _AES_ENC_n821, _AES_ENC_n820, _AES_ENC_n819, _AES_ENC_n818, _AES_ENC_n817, _AES_ENC_n816, _AES_ENC_n815, _AES_ENC_n814, _AES_ENC_n813, _AES_ENC_n812, _AES_ENC_n811, _AES_ENC_n810, _AES_ENC_n809, _AES_ENC_n808, _AES_ENC_n807, _AES_ENC_n806, _AES_ENC_n805, _AES_ENC_n804, _AES_ENC_n803, _AES_ENC_n802, _AES_ENC_n801, _AES_ENC_n800, _AES_ENC_n799, _AES_ENC_n798, _AES_ENC_n797, _AES_ENC_n796, _AES_ENC_n795, _AES_ENC_n788, 
  _AES_ENC_n787, _AES_ENC_n786, _AES_ENC_n785, _AES_ENC_n784, _AES_ENC_n783, _AES_ENC_n782, _AES_ENC_n781, _AES_ENC_n780, _AES_ENC_n779, _AES_ENC_n778, _AES_ENC_n777, _AES_ENC_n776, _AES_ENC_n775, _AES_ENC_n774, _AES_ENC_n773, _AES_ENC_n772, _AES_ENC_n771, _AES_ENC_n770, _AES_ENC_n769, _AES_ENC_n768, _AES_ENC_n767, _AES_ENC_n766, _AES_ENC_n765, _AES_ENC_n764, _AES_ENC_n763, _AES_ENC_n762, _AES_ENC_n761, _AES_ENC_n760, _AES_ENC_n759, _AES_ENC_n758, _AES_ENC_n757, _AES_ENC_n756, _AES_ENC_n755, _AES_ENC_n754, _AES_ENC_n753, _AES_ENC_n752, _AES_ENC_n751, _AES_ENC_n750, _AES_ENC_n749, _AES_ENC_n748, _AES_ENC_n747, _AES_ENC_n746, _AES_ENC_n745, _AES_ENC_n744, _AES_ENC_n743, _AES_ENC_n742, _AES_ENC_n741, _AES_ENC_n740, _AES_ENC_n739, _AES_ENC_n738, 
  _AES_ENC_n737, _AES_ENC_n736, _AES_ENC_n735, _AES_ENC_n734, _AES_ENC_n733, _AES_ENC_n732, _AES_ENC_n731, _AES_ENC_n730, _AES_ENC_n729, _AES_ENC_n728, _AES_ENC_n727, _AES_ENC_n726, _AES_ENC_n725, _AES_ENC_n724, _AES_ENC_n723, _AES_ENC_n722, _AES_ENC_n721, _AES_ENC_n720, _AES_ENC_n719, _AES_ENC_n718, _AES_ENC_n717, _AES_ENC_n716, _AES_ENC_n715, _AES_ENC_n714, _AES_ENC_n713, _AES_ENC_n712, _AES_ENC_n711, _AES_ENC_n710, _AES_ENC_n709, _AES_ENC_n708, _AES_ENC_n707, _AES_ENC_n706, _AES_ENC_n705, _AES_ENC_n704, _AES_ENC_n703, _AES_ENC_n702, _AES_ENC_n701, _AES_ENC_n700, _AES_ENC_n699, _AES_ENC_n698, _AES_ENC_n697, _AES_ENC_n696, _AES_ENC_n695, _AES_ENC_n694, _AES_ENC_n693, _AES_ENC_n692, _AES_ENC_n691, _AES_ENC_n690, _AES_ENC_n689, _AES_ENC_n688, 
  _AES_ENC_n687, _AES_ENC_n686, _AES_ENC_n685, _AES_ENC_n684, _AES_ENC_n683, _AES_ENC_n682, _AES_ENC_n681, _AES_ENC_n680, _AES_ENC_n679, _AES_ENC_n678, _AES_ENC_n677, _AES_ENC_n676, _AES_ENC_n675, _AES_ENC_n674, _AES_ENC_n673, _AES_ENC_n672, _AES_ENC_n671, _AES_ENC_n670, _AES_ENC_n669, _AES_ENC_n668, _AES_ENC_n667, _AES_ENC_n666, _AES_ENC_n665, _AES_ENC_n664, _AES_ENC_n663, _AES_ENC_n662, _AES_ENC_n661, _AES_ENC_N501, _AES_ENC_N500, _AES_ENC_N499, _AES_ENC_N498, _AES_ENC_N497, _AES_ENC_N496, _AES_ENC_N495, _AES_ENC_N494, _AES_ENC_N493, _AES_ENC_N492, _AES_ENC_N491, _AES_ENC_N490, _AES_ENC_N489, _AES_ENC_N488, _AES_ENC_N487, _AES_ENC_N486, _AES_ENC_N485, _AES_ENC_N484, _AES_ENC_N483, _AES_ENC_N482, _AES_ENC_N481, _AES_ENC_N480, _AES_ENC_N479, 
  _AES_ENC_N478, _AES_ENC_N477, _AES_ENC_N476, _AES_ENC_N475, _AES_ENC_N474, _AES_ENC_N473, _AES_ENC_N472, _AES_ENC_N471, _AES_ENC_N470, _AES_ENC_N469, _AES_ENC_N468, _AES_ENC_N467, _AES_ENC_N466, _AES_ENC_N465, _AES_ENC_N464, _AES_ENC_N463, _AES_ENC_N462, _AES_ENC_N461, _AES_ENC_N460, _AES_ENC_N459, _AES_ENC_N458, _AES_ENC_N457, _AES_ENC_N456, _AES_ENC_N455, _AES_ENC_N454, _AES_ENC_N453, _AES_ENC_N452, _AES_ENC_N451, _AES_ENC_N450, _AES_ENC_N449, _AES_ENC_N448, _AES_ENC_N447, _AES_ENC_N446, _AES_ENC_N445, _AES_ENC_N444, _AES_ENC_N443, _AES_ENC_N442, _AES_ENC_N441, _AES_ENC_N440, _AES_ENC_N439, _AES_ENC_N438, _AES_ENC_N437, _AES_ENC_N436, _AES_ENC_N435, _AES_ENC_N434, _AES_ENC_N433, _AES_ENC_N432, _AES_ENC_N431, _AES_ENC_N430, _AES_ENC_N429, 
  _AES_ENC_N428, _AES_ENC_N427, _AES_ENC_N426, _AES_ENC_N425, _AES_ENC_N424, _AES_ENC_N423, _AES_ENC_N422, _AES_ENC_N421, _AES_ENC_N420, _AES_ENC_N419, _AES_ENC_N418, _AES_ENC_N417, _AES_ENC_N416, _AES_ENC_N415, _AES_ENC_N414, _AES_ENC_N413, _AES_ENC_N412, _AES_ENC_N411, _AES_ENC_N410, _AES_ENC_N409, _AES_ENC_N408, _AES_ENC_N407, _AES_ENC_N406, _AES_ENC_N405, _AES_ENC_N404, _AES_ENC_N403, _AES_ENC_N402, _AES_ENC_N401, _AES_ENC_N400, _AES_ENC_N399, _AES_ENC_N398, _AES_ENC_N397, _AES_ENC_N396, _AES_ENC_N395, _AES_ENC_N394, _AES_ENC_N393, _AES_ENC_N392, _AES_ENC_N391, _AES_ENC_N390, _AES_ENC_N389, _AES_ENC_N388, _AES_ENC_N387, _AES_ENC_N386, _AES_ENC_N385, _AES_ENC_N384, _AES_ENC_N383, _AES_ENC_N382, _AES_ENC_N381, _AES_ENC_N380, _AES_ENC_N379, 
  _AES_ENC_N378, _AES_ENC_N377, _AES_ENC_N376, _AES_ENC_N375, _AES_ENC_N374, _AES_ENC_sa33_sub[0], _AES_ENC_sa33_sub[1], _AES_ENC_sa33_sub[2], _AES_ENC_sa33_sub[3], _AES_ENC_sa33_sub[4], _AES_ENC_sa33_sub[5], _AES_ENC_sa33_sub[6], _AES_ENC_sa33_sub[7], _AES_ENC_sa32_sub[0], _AES_ENC_sa32_sub[1], _AES_ENC_sa32_sub[2], _AES_ENC_sa32_sub[3], _AES_ENC_sa32_sub[4], _AES_ENC_sa32_sub[5], _AES_ENC_sa32_sub[6], _AES_ENC_sa32_sub[7], _AES_ENC_sa31_sub[0], _AES_ENC_sa31_sub[1], _AES_ENC_sa31_sub[2], _AES_ENC_sa31_sub[3], _AES_ENC_sa31_sub[4], _AES_ENC_sa31_sub[5], _AES_ENC_sa31_sub[6], _AES_ENC_sa31_sub[7], _AES_ENC_sa30_sub[0], _AES_ENC_sa30_sub[1], _AES_ENC_sa30_sub[2], _AES_ENC_sa30_sub[3], _AES_ENC_sa30_sub[4], _AES_ENC_sa30_sub[5], _AES_ENC_sa30_sub[6], _AES_ENC_sa30_sub[7], _AES_ENC_sa23_sub[0], _AES_ENC_sa23_sub[1], _AES_ENC_sa23_sub[2], _AES_ENC_sa23_sub[3], _AES_ENC_sa23_sub[4], _AES_ENC_sa23_sub[5], _AES_ENC_sa23_sub[6], _AES_ENC_sa23_sub[7], _AES_ENC_sa22_sub[0], _AES_ENC_sa22_sub[1], _AES_ENC_sa22_sub[2], _AES_ENC_sa22_sub[3], _AES_ENC_sa22_sub[4], 
  _AES_ENC_sa22_sub[5], _AES_ENC_sa22_sub[6], _AES_ENC_sa22_sub[7], _AES_ENC_sa21_sub[0], _AES_ENC_sa21_sub[1], _AES_ENC_sa21_sub[2], _AES_ENC_sa21_sub[3], _AES_ENC_sa21_sub[4], _AES_ENC_sa21_sub[5], _AES_ENC_sa21_sub[6], _AES_ENC_sa21_sub[7], _AES_ENC_sa20_sub[0], _AES_ENC_sa20_sub[1], _AES_ENC_sa20_sub[2], _AES_ENC_sa20_sub[3], _AES_ENC_sa20_sub[4], _AES_ENC_sa20_sub[5], _AES_ENC_sa20_sub[6], _AES_ENC_sa20_sub[7], _AES_ENC_sa13_sub[0], _AES_ENC_sa13_sub[1], _AES_ENC_sa13_sub[2], _AES_ENC_sa13_sub[3], _AES_ENC_sa13_sub[4], _AES_ENC_sa13_sub[5], _AES_ENC_sa13_sub[6], _AES_ENC_sa13_sub[7], _AES_ENC_sa12_sub[0], _AES_ENC_sa12_sub[1], _AES_ENC_sa12_sub[2], _AES_ENC_sa12_sub[3], _AES_ENC_sa12_sub[4], _AES_ENC_sa12_sub[5], _AES_ENC_sa12_sub[6], _AES_ENC_sa12_sub[7], _AES_ENC_sa11_sub[0], _AES_ENC_sa11_sub[1], _AES_ENC_sa11_sub[2], _AES_ENC_sa11_sub[3], _AES_ENC_sa11_sub[4], _AES_ENC_sa11_sub[5], _AES_ENC_sa11_sub[6], _AES_ENC_sa11_sub[7], _AES_ENC_sa10_sub[0], _AES_ENC_sa10_sub[1], _AES_ENC_sa10_sub[2], _AES_ENC_sa10_sub[3], _AES_ENC_sa10_sub[4], _AES_ENC_sa10_sub[5], _AES_ENC_sa10_sub[6], 
  _AES_ENC_sa10_sub[7], _AES_ENC_sa03_sub[0], _AES_ENC_sa03_sub[1], _AES_ENC_sa03_sub[2], _AES_ENC_sa03_sub[3], _AES_ENC_sa03_sub[4], _AES_ENC_sa03_sub[5], _AES_ENC_sa03_sub[6], _AES_ENC_sa03_sub[7], _AES_ENC_sa02_sub[0], _AES_ENC_sa02_sub[1], _AES_ENC_sa02_sub[2], _AES_ENC_sa02_sub[3], _AES_ENC_sa02_sub[4], _AES_ENC_sa02_sub[5], _AES_ENC_sa02_sub[6], _AES_ENC_sa02_sub[7], _AES_ENC_sa01_sub[0], _AES_ENC_sa01_sub[1], _AES_ENC_sa01_sub[2], _AES_ENC_sa01_sub[3], _AES_ENC_sa01_sub[4], _AES_ENC_sa01_sub[5], _AES_ENC_sa01_sub[6], _AES_ENC_sa01_sub[7], _AES_ENC_sa00_sub[0], _AES_ENC_sa00_sub[1], _AES_ENC_sa00_sub[2], _AES_ENC_sa00_sub[3], _AES_ENC_sa00_sub[4], _AES_ENC_sa00_sub[5], _AES_ENC_sa00_sub[6], _AES_ENC_sa00_sub[7], _AES_ENC_N277, _AES_ENC_N276, _AES_ENC_N275, _AES_ENC_N274, _AES_ENC_N273, _AES_ENC_N272, _AES_ENC_N271, _AES_ENC_N270, _AES_ENC_N261, _AES_ENC_N260, _AES_ENC_N259, _AES_ENC_N258, _AES_ENC_N257, _AES_ENC_N256, _AES_ENC_N255, _AES_ENC_N254, _AES_ENC_N245, 
  _AES_ENC_N244, _AES_ENC_N243, _AES_ENC_N242, _AES_ENC_N241, _AES_ENC_N240, _AES_ENC_N239, _AES_ENC_N238, _AES_ENC_N229, _AES_ENC_N228, _AES_ENC_N227, _AES_ENC_N226, _AES_ENC_N225, _AES_ENC_N224, _AES_ENC_N223, _AES_ENC_N222, _AES_ENC_w0[0], _AES_ENC_w0[1], _AES_ENC_w0[2], _AES_ENC_w0[3], _AES_ENC_w0[4], _AES_ENC_w0[5], _AES_ENC_w0[6], _AES_ENC_w0[7], _AES_ENC_w0[8], _AES_ENC_w0[9], _AES_ENC_w0[10], _AES_ENC_w0[11], _AES_ENC_w0[12], _AES_ENC_w0[13], _AES_ENC_w0[14], _AES_ENC_w0[15], _AES_ENC_w0[16], _AES_ENC_w0[17], _AES_ENC_w0[18], _AES_ENC_w0[19], _AES_ENC_w0[20], _AES_ENC_w0[21], _AES_ENC_w0[22], _AES_ENC_w0[23], _AES_ENC_w0[24], _AES_ENC_w0[25], _AES_ENC_w0[26], _AES_ENC_w0[27], _AES_ENC_w0[28], _AES_ENC_w0[29], _AES_ENC_w0[30], _AES_ENC_w0[31], _AES_ENC_N213, _AES_ENC_N212, _AES_ENC_N211, 
  _AES_ENC_N210, _AES_ENC_N209, _AES_ENC_N208, _AES_ENC_N207, _AES_ENC_N206, _AES_ENC_N197, _AES_ENC_N196, _AES_ENC_N195, _AES_ENC_N194, _AES_ENC_N193, _AES_ENC_N192, _AES_ENC_N191, _AES_ENC_N190, _AES_ENC_N181, _AES_ENC_N180, _AES_ENC_N179, _AES_ENC_N178, _AES_ENC_N177, _AES_ENC_N176, _AES_ENC_N175, _AES_ENC_N174, _AES_ENC_N165, _AES_ENC_N164, _AES_ENC_N163, _AES_ENC_N162, _AES_ENC_N161, _AES_ENC_N160, _AES_ENC_N159, _AES_ENC_N158, _AES_ENC_w1[0], _AES_ENC_w1[1], _AES_ENC_w1[2], _AES_ENC_w1[3], _AES_ENC_w1[4], _AES_ENC_w1[5], _AES_ENC_w1[6], _AES_ENC_w1[7], _AES_ENC_w1[8], _AES_ENC_w1[9], _AES_ENC_w1[10], _AES_ENC_w1[11], _AES_ENC_w1[12], _AES_ENC_w1[13], _AES_ENC_w1[14], _AES_ENC_w1[15], _AES_ENC_w1[16], _AES_ENC_w1[17], _AES_ENC_w1[18], _AES_ENC_w1[19], _AES_ENC_w1[20], 
  _AES_ENC_w1[21], _AES_ENC_w1[22], _AES_ENC_w1[23], _AES_ENC_w1[24], _AES_ENC_w1[25], _AES_ENC_w1[26], _AES_ENC_w1[27], _AES_ENC_w1[28], _AES_ENC_w1[29], _AES_ENC_w1[30], _AES_ENC_w1[31], _AES_ENC_N149, _AES_ENC_N148, _AES_ENC_N147, _AES_ENC_N146, _AES_ENC_N145, _AES_ENC_N144, _AES_ENC_N143, _AES_ENC_N142, _AES_ENC_N133, _AES_ENC_N132, _AES_ENC_N131, _AES_ENC_N130, _AES_ENC_N129, _AES_ENC_N128, _AES_ENC_N127, _AES_ENC_N126, _AES_ENC_N117, _AES_ENC_N116, _AES_ENC_N115, _AES_ENC_N114, _AES_ENC_N113, _AES_ENC_N112, _AES_ENC_N111, _AES_ENC_N110, _AES_ENC_N101, _AES_ENC_N100, _AES_ENC_N99, _AES_ENC_N98, _AES_ENC_N97, _AES_ENC_N96, _AES_ENC_N95, _AES_ENC_N94, _AES_ENC_w2[0], _AES_ENC_w2[1], _AES_ENC_w2[2], _AES_ENC_w2[3], _AES_ENC_w2[4], _AES_ENC_w2[5], _AES_ENC_w2[6], 
  _AES_ENC_w2[7], _AES_ENC_w2[8], _AES_ENC_w2[9], _AES_ENC_w2[10], _AES_ENC_w2[11], _AES_ENC_w2[12], _AES_ENC_w2[13], _AES_ENC_w2[14], _AES_ENC_w2[15], _AES_ENC_w2[16], _AES_ENC_w2[17], _AES_ENC_w2[18], _AES_ENC_w2[19], _AES_ENC_w2[20], _AES_ENC_w2[21], _AES_ENC_w2[22], _AES_ENC_w2[23], _AES_ENC_w2[24], _AES_ENC_w2[25], _AES_ENC_w2[26], _AES_ENC_w2[27], _AES_ENC_w2[28], _AES_ENC_w2[29], _AES_ENC_w2[30], _AES_ENC_w2[31], _AES_ENC_N85, _AES_ENC_N84, _AES_ENC_N83, _AES_ENC_N82, _AES_ENC_N81, _AES_ENC_N80, _AES_ENC_N79, _AES_ENC_N78, _AES_ENC_N69, _AES_ENC_N68, _AES_ENC_N67, _AES_ENC_N66, _AES_ENC_N65, _AES_ENC_N64, _AES_ENC_N63, _AES_ENC_N62, _AES_ENC_N53, _AES_ENC_N52, _AES_ENC_N51, _AES_ENC_N50, _AES_ENC_N49, _AES_ENC_N48, _AES_ENC_N47, _AES_ENC_N46, _AES_ENC_N37, 
  _AES_ENC_N36, _AES_ENC_N35, _AES_ENC_N34, _AES_ENC_N33, _AES_ENC_N32, _AES_ENC_N31, _AES_ENC_N30, _AES_ENC_w3[0], _AES_ENC_w3[1], _AES_ENC_w3[2], _AES_ENC_w3[3], _AES_ENC_w3[4], _AES_ENC_w3[5], _AES_ENC_w3[6], _AES_ENC_w3[7], _AES_ENC_w3[8], _AES_ENC_w3[9], _AES_ENC_w3[10], _AES_ENC_w3[11], _AES_ENC_w3[12], _AES_ENC_w3[13], _AES_ENC_w3[14], _AES_ENC_w3[15], _AES_ENC_w3[16], _AES_ENC_w3[17], _AES_ENC_w3[18], _AES_ENC_w3[19], _AES_ENC_w3[20], _AES_ENC_w3[21], _AES_ENC_w3[22], _AES_ENC_w3[23], _AES_ENC_w3[24], _AES_ENC_w3[25], _AES_ENC_w3[26], _AES_ENC_w3[27], _AES_ENC_w3[28], _AES_ENC_w3[29], _AES_ENC_w3[30], _AES_ENC_w3[31], _AES_ENC_text_in_r[0], _AES_ENC_text_in_r[1], _AES_ENC_text_in_r[2], _AES_ENC_text_in_r[3], _AES_ENC_text_in_r[4], _AES_ENC_text_in_r[5], _AES_ENC_text_in_r[6], _AES_ENC_text_in_r[7], _AES_ENC_text_in_r[8], _AES_ENC_text_in_r[9], _AES_ENC_text_in_r[10], 
  _AES_ENC_text_in_r[11], _AES_ENC_text_in_r[12], _AES_ENC_text_in_r[13], _AES_ENC_text_in_r[14], _AES_ENC_text_in_r[15], _AES_ENC_text_in_r[16], _AES_ENC_text_in_r[17], _AES_ENC_text_in_r[18], _AES_ENC_text_in_r[19], _AES_ENC_text_in_r[20], _AES_ENC_text_in_r[21], _AES_ENC_text_in_r[22], _AES_ENC_text_in_r[23], _AES_ENC_text_in_r[24], _AES_ENC_text_in_r[25], _AES_ENC_text_in_r[26], _AES_ENC_text_in_r[27], _AES_ENC_text_in_r[28], _AES_ENC_text_in_r[29], _AES_ENC_text_in_r[30], _AES_ENC_text_in_r[31], _AES_ENC_text_in_r[32], _AES_ENC_text_in_r[33], _AES_ENC_text_in_r[34], _AES_ENC_text_in_r[35], _AES_ENC_text_in_r[36], _AES_ENC_text_in_r[37], _AES_ENC_text_in_r[38], _AES_ENC_text_in_r[39], _AES_ENC_text_in_r[40], _AES_ENC_text_in_r[41], _AES_ENC_text_in_r[42], _AES_ENC_text_in_r[43], _AES_ENC_text_in_r[44], _AES_ENC_text_in_r[45], _AES_ENC_text_in_r[46], _AES_ENC_text_in_r[47], _AES_ENC_text_in_r[48], _AES_ENC_text_in_r[49], _AES_ENC_text_in_r[50], _AES_ENC_text_in_r[51], _AES_ENC_text_in_r[52], _AES_ENC_text_in_r[53], _AES_ENC_text_in_r[54], _AES_ENC_text_in_r[55], _AES_ENC_text_in_r[56], _AES_ENC_text_in_r[57], _AES_ENC_text_in_r[58], _AES_ENC_text_in_r[59], _AES_ENC_text_in_r[60], 
  _AES_ENC_text_in_r[61], _AES_ENC_text_in_r[62], _AES_ENC_text_in_r[63], _AES_ENC_text_in_r[64], _AES_ENC_text_in_r[65], _AES_ENC_text_in_r[66], _AES_ENC_text_in_r[67], _AES_ENC_text_in_r[68], _AES_ENC_text_in_r[69], _AES_ENC_text_in_r[70], _AES_ENC_text_in_r[71], _AES_ENC_text_in_r[72], _AES_ENC_text_in_r[73], _AES_ENC_text_in_r[74], _AES_ENC_text_in_r[75], _AES_ENC_text_in_r[76], _AES_ENC_text_in_r[77], _AES_ENC_text_in_r[78], _AES_ENC_text_in_r[79], _AES_ENC_text_in_r[80], _AES_ENC_text_in_r[81], _AES_ENC_text_in_r[82], _AES_ENC_text_in_r[83], _AES_ENC_text_in_r[84], _AES_ENC_text_in_r[85], _AES_ENC_text_in_r[86], _AES_ENC_text_in_r[87], _AES_ENC_text_in_r[88], _AES_ENC_text_in_r[89], _AES_ENC_text_in_r[90], _AES_ENC_text_in_r[91], _AES_ENC_text_in_r[92], _AES_ENC_text_in_r[93], _AES_ENC_text_in_r[94], _AES_ENC_text_in_r[95], _AES_ENC_text_in_r[96], _AES_ENC_text_in_r[97], _AES_ENC_text_in_r[98], _AES_ENC_text_in_r[99], _AES_ENC_text_in_r[100], _AES_ENC_text_in_r[101], _AES_ENC_text_in_r[102], _AES_ENC_text_in_r[103], _AES_ENC_text_in_r[104], _AES_ENC_text_in_r[105], _AES_ENC_text_in_r[106], _AES_ENC_text_in_r[107], _AES_ENC_text_in_r[108], _AES_ENC_text_in_r[109], _AES_ENC_text_in_r[110], 
  _AES_ENC_text_in_r[111], _AES_ENC_text_in_r[112], _AES_ENC_text_in_r[113], _AES_ENC_text_in_r[114], _AES_ENC_text_in_r[115], _AES_ENC_text_in_r[116], _AES_ENC_text_in_r[117], _AES_ENC_text_in_r[118], _AES_ENC_text_in_r[119], _AES_ENC_text_in_r[120], _AES_ENC_text_in_r[121], _AES_ENC_text_in_r[122], _AES_ENC_text_in_r[123], _AES_ENC_text_in_r[124], _AES_ENC_text_in_r[125], _AES_ENC_text_in_r[126], _AES_ENC_text_in_r[127], _AES_ENC_N19, _AES_ENC_u0_n325, _AES_ENC_u0_n324, _AES_ENC_u0_n323, _AES_ENC_u0_n322, _AES_ENC_u0_n321, _AES_ENC_u0_n320, _AES_ENC_u0_n319, _AES_ENC_u0_n318, _AES_ENC_u0_n317, _AES_ENC_u0_n316, _AES_ENC_u0_n315, _AES_ENC_u0_n314, _AES_ENC_u0_n281, _AES_ENC_u0_n280, _AES_ENC_u0_n279, _AES_ENC_u0_n278, _AES_ENC_u0_n277, _AES_ENC_u0_n276, _AES_ENC_u0_n275, _AES_ENC_u0_n274, _AES_ENC_u0_n273, _AES_ENC_u0_n272, _AES_ENC_u0_n2710, _AES_ENC_u0_n2700, _AES_ENC_u0_n2690, _AES_ENC_u0_n2680, _AES_ENC_u0_n2670, _AES_ENC_u0_n2660, _AES_ENC_u0_n2650, _AES_ENC_u0_n2640, _AES_ENC_u0_n2630, _AES_ENC_u0_n2620, 
  _AES_ENC_u0_n2610, _AES_ENC_u0_n2600, _AES_ENC_u0_n2590, _AES_ENC_u0_n2580, _AES_ENC_u0_n2570, _AES_ENC_u0_n2560, _AES_ENC_u0_n2550, _AES_ENC_u0_n2540, _AES_ENC_u0_n2530, _AES_ENC_u0_n2520, _AES_ENC_u0_n2510, _AES_ENC_u0_n2500, _AES_ENC_u0_n2490, _AES_ENC_u0_n2480, _AES_ENC_u0_n2470, _AES_ENC_u0_n2460, _AES_ENC_u0_n2450, _AES_ENC_u0_n2440, _AES_ENC_u0_n2430, _AES_ENC_u0_n2420, _AES_ENC_u0_n2410, _AES_ENC_u0_n2400, _AES_ENC_u0_n2390, _AES_ENC_u0_n2380, _AES_ENC_u0_n2370, _AES_ENC_u0_n2360, _AES_ENC_u0_n2350, _AES_ENC_u0_n2340, _AES_ENC_u0_n2330, _AES_ENC_u0_n2320, _AES_ENC_u0_n2310, _AES_ENC_u0_n2300, _AES_ENC_u0_n2290, _AES_ENC_u0_n2280, _AES_ENC_u0_n2270, _AES_ENC_u0_n2260, _AES_ENC_u0_n2250, _AES_ENC_u0_n2240, _AES_ENC_u0_n2230, _AES_ENC_u0_n2220, _AES_ENC_u0_n2210, _AES_ENC_u0_n2200, _AES_ENC_u0_n2190, _AES_ENC_u0_n2180, _AES_ENC_u0_n2170, _AES_ENC_u0_n2160, _AES_ENC_u0_n2150, _AES_ENC_u0_n2140, _AES_ENC_u0_n2130, _AES_ENC_u0_n2120, 
  _AES_ENC_u0_n2110, _AES_ENC_u0_n2100, _AES_ENC_u0_n2090, _AES_ENC_u0_n2080, _AES_ENC_u0_n207, _AES_ENC_u0_n206, _AES_ENC_u0_n2050, _AES_ENC_u0_n2040, _AES_ENC_u0_n2030, _AES_ENC_u0_n2020, _AES_ENC_u0_n2010, _AES_ENC_u0_n2000, _AES_ENC_u0_n1990, _AES_ENC_u0_n1980, _AES_ENC_u0_n1970, _AES_ENC_u0_n1960, _AES_ENC_u0_n1950, _AES_ENC_u0_n1940, _AES_ENC_u0_n1930, _AES_ENC_u0_n1920, _AES_ENC_u0_n1910, _AES_ENC_u0_n1900, _AES_ENC_u0_n1890, _AES_ENC_u0_n1880, _AES_ENC_u0_n1870, _AES_ENC_u0_n1860, _AES_ENC_u0_n1850, _AES_ENC_u0_n1840, _AES_ENC_u0_n1830, _AES_ENC_u0_n1820, _AES_ENC_u0_n1810, _AES_ENC_u0_n1800, _AES_ENC_u0_n1790, _AES_ENC_u0_n1780, _AES_ENC_u0_n1770, _AES_ENC_u0_n1760, _AES_ENC_u0_n1750, _AES_ENC_u0_n1740, _AES_ENC_u0_n1730, _AES_ENC_u0_n1720, _AES_ENC_u0_n1711, _AES_ENC_u0_n1700, _AES_ENC_u0_n1690, _AES_ENC_u0_n1680, _AES_ENC_u0_n1670, _AES_ENC_u0_n1660, _AES_ENC_u0_n1650, _AES_ENC_u0_n1640, _AES_ENC_u0_n1630, _AES_ENC_u0_n1620, 
  _AES_ENC_u0_n1611, _AES_ENC_u0_n1600, _AES_ENC_u0_n1590, _AES_ENC_u0_n1580, _AES_ENC_u0_n1570, _AES_ENC_u0_n1560, _AES_ENC_u0_n1550, _AES_ENC_u0_n1540, _AES_ENC_u0_n1530, _AES_ENC_u0_n1520, _AES_ENC_u0_n1511, _AES_ENC_u0_n1500, _AES_ENC_u0_n1490, _AES_ENC_u0_n1480, _AES_ENC_u0_n1470, _AES_ENC_u0_n1460, _AES_ENC_u0_n1450, _AES_ENC_u0_n1440, _AES_ENC_u0_n1430, _AES_ENC_u0_n1420, _AES_ENC_u0_n141, _AES_ENC_u0_n1401, _AES_ENC_u0_n1390, _AES_ENC_u0_n1380, _AES_ENC_u0_n1370, _AES_ENC_u0_n1360, _AES_ENC_u0_n1350, _AES_ENC_u0_n1340, _AES_ENC_u0_n1330, _AES_ENC_u0_n1320, _AES_ENC_u0_n1311, _AES_ENC_u0_n1300, _AES_ENC_u0_n1290, _AES_ENC_u0_n1280, _AES_ENC_u0_n1270, _AES_ENC_u0_n1260, _AES_ENC_u0_n1250, _AES_ENC_u0_n1240, _AES_ENC_u0_n1230, _AES_ENC_u0_n1220, _AES_ENC_u0_n1211, _AES_ENC_u0_n1200, _AES_ENC_u0_n1190, _AES_ENC_u0_n1180, _AES_ENC_u0_n1170, _AES_ENC_u0_n1160, _AES_ENC_u0_n1150, _AES_ENC_u0_n1140, _AES_ENC_u0_n1130, _AES_ENC_u0_n1120, 
  _AES_ENC_u0_n1111, _AES_ENC_u0_n1100, _AES_ENC_u0_n1090, _AES_ENC_u0_n1080, _AES_ENC_u0_n1070, _AES_ENC_u0_n1060, _AES_ENC_u0_n1050, _AES_ENC_u0_n1040, _AES_ENC_u0_n1030, _AES_ENC_u0_n1020, _AES_ENC_u0_n1011, _AES_ENC_u0_n1000, _AES_ENC_u0_n990, _AES_ENC_u0_n980, _AES_ENC_u0_n970, _AES_ENC_u0_n960, _AES_ENC_u0_n950, _AES_ENC_u0_n940, _AES_ENC_u0_n930, _AES_ENC_u0_n920, _AES_ENC_u0_n910, _AES_ENC_u0_n900, _AES_ENC_u0_n890, _AES_ENC_u0_n880, _AES_ENC_u0_n870, _AES_ENC_u0_n860, _AES_ENC_u0_n850, _AES_ENC_u0_n840, _AES_ENC_u0_n830, _AES_ENC_u0_n820, _AES_ENC_u0_n810, _AES_ENC_u0_n800, _AES_ENC_u0_n790, _AES_ENC_u0_n780, _AES_ENC_u0_n770, _AES_ENC_u0_n760, _AES_ENC_u0_n75, _AES_ENC_u0_n74, _AES_ENC_u0_n730, _AES_ENC_u0_n720, _AES_ENC_u0_n710, _AES_ENC_u0_n700, _AES_ENC_u0_n690, _AES_ENC_u0_n680, _AES_ENC_u0_n670, _AES_ENC_u0_n660, _AES_ENC_u0_n650, _AES_ENC_u0_n640, _AES_ENC_u0_n630, _AES_ENC_u0_n620, 
  _AES_ENC_u0_n610, _AES_ENC_u0_n600, _AES_ENC_u0_n590, _AES_ENC_u0_n580, _AES_ENC_u0_n570, _AES_ENC_u0_n560, _AES_ENC_u0_n550, _AES_ENC_u0_n540, _AES_ENC_u0_n530, _AES_ENC_u0_n520, _AES_ENC_u0_n510, _AES_ENC_u0_n500, _AES_ENC_u0_n490, _AES_ENC_u0_n480, _AES_ENC_u0_n470, _AES_ENC_u0_n460, _AES_ENC_u0_n450, _AES_ENC_u0_n440, _AES_ENC_u0_n430, _AES_ENC_u0_n420, _AES_ENC_u0_n41, _AES_ENC_u0_n40, _AES_ENC_u0_n39, _AES_ENC_u0_n38, _AES_ENC_u0_n37, _AES_ENC_u0_n36, _AES_ENC_u0_n35, _AES_ENC_u0_n34, _AES_ENC_u0_n33, _AES_ENC_u0_n32, _AES_ENC_u0_n31, _AES_ENC_u0_n30, _AES_ENC_u0_n29, _AES_ENC_u0_n28, _AES_ENC_u0_n27, _AES_ENC_u0_n26, _AES_ENC_u0_n25, _AES_ENC_u0_n24, _AES_ENC_u0_n23, _AES_ENC_u0_n22, _AES_ENC_u0_n21, _AES_ENC_u0_n20, _AES_ENC_u0_n19, _AES_ENC_u0_n18, _AES_ENC_u0_n1710, _AES_ENC_u0_n1610, _AES_ENC_u0_n1510, _AES_ENC_u0_n1400, _AES_ENC_u0_n1310, _AES_ENC_u0_n1210, 
  _AES_ENC_u0_n1110, _AES_ENC_u0_n1010, _AES_ENC_u0_n9, _AES_ENC_u0_n8, _AES_ENC_u0_n7, _AES_ENC_u0_n6, _AES_ENC_u0_n5, _AES_ENC_u0_n4, _AES_ENC_u0_n3, _AES_ENC_u0_n2, _AES_ENC_u0_n313, _AES_ENC_u0_n312, _AES_ENC_u0_n311, _AES_ENC_u0_n310, _AES_ENC_u0_n309, _AES_ENC_u0_n308, _AES_ENC_u0_n307, _AES_ENC_u0_n306, _AES_ENC_u0_n305, _AES_ENC_u0_n304, _AES_ENC_u0_n303, _AES_ENC_u0_n302, _AES_ENC_u0_n301, _AES_ENC_u0_n300, _AES_ENC_u0_n299, _AES_ENC_u0_n298, _AES_ENC_u0_n297, _AES_ENC_u0_n296, _AES_ENC_u0_n295, _AES_ENC_u0_n294, _AES_ENC_u0_n293, _AES_ENC_u0_n292, _AES_ENC_u0_n291, _AES_ENC_u0_n290, _AES_ENC_u0_n289, _AES_ENC_u0_n288, _AES_ENC_u0_n287, _AES_ENC_u0_n286, _AES_ENC_u0_n285, _AES_ENC_u0_n284, _AES_ENC_u0_n283, _AES_ENC_u0_n282, _AES_ENC_u0_N271, _AES_ENC_u0_N270, _AES_ENC_u0_N269, _AES_ENC_u0_N268, _AES_ENC_u0_N267, _AES_ENC_u0_N266, _AES_ENC_u0_N265, _AES_ENC_u0_N264, 
  _AES_ENC_u0_N263, _AES_ENC_u0_N262, _AES_ENC_u0_N261, _AES_ENC_u0_N260, _AES_ENC_u0_N259, _AES_ENC_u0_N258, _AES_ENC_u0_N257, _AES_ENC_u0_N256, _AES_ENC_u0_N255, _AES_ENC_u0_N254, _AES_ENC_u0_N253, _AES_ENC_u0_N252, _AES_ENC_u0_N251, _AES_ENC_u0_N250, _AES_ENC_u0_N249, _AES_ENC_u0_N248, _AES_ENC_u0_N247, _AES_ENC_u0_N246, _AES_ENC_u0_N245, _AES_ENC_u0_N244, _AES_ENC_u0_N243, _AES_ENC_u0_N242, _AES_ENC_u0_N241, _AES_ENC_u0_N240, _AES_ENC_u0_N239, _AES_ENC_u0_N238, _AES_ENC_u0_N237, _AES_ENC_u0_N236, _AES_ENC_u0_N235, _AES_ENC_u0_N234, _AES_ENC_u0_N233, _AES_ENC_u0_N232, _AES_ENC_u0_N231, _AES_ENC_u0_N230, _AES_ENC_u0_N229, _AES_ENC_u0_N228, _AES_ENC_u0_N227, _AES_ENC_u0_N226, _AES_ENC_u0_N225, _AES_ENC_u0_N224, _AES_ENC_u0_N223, _AES_ENC_u0_N222, _AES_ENC_u0_N221, _AES_ENC_u0_N220, _AES_ENC_u0_N219, _AES_ENC_u0_N218, _AES_ENC_u0_N217, _AES_ENC_u0_N216, _AES_ENC_u0_N215, _AES_ENC_u0_N214, 
  _AES_ENC_u0_N213, _AES_ENC_u0_N212, _AES_ENC_u0_N211, _AES_ENC_u0_N210, _AES_ENC_u0_N209, _AES_ENC_u0_N208, _AES_ENC_u0_N205, _AES_ENC_u0_N204, _AES_ENC_u0_N203, _AES_ENC_u0_N202, _AES_ENC_u0_N201, _AES_ENC_u0_N200, _AES_ENC_u0_N199, _AES_ENC_u0_N198, _AES_ENC_u0_N197, _AES_ENC_u0_N196, _AES_ENC_u0_N195, _AES_ENC_u0_N194, _AES_ENC_u0_N193, _AES_ENC_u0_N192, _AES_ENC_u0_N191, _AES_ENC_u0_N190, _AES_ENC_u0_N189, _AES_ENC_u0_N188, _AES_ENC_u0_N187, _AES_ENC_u0_N186, _AES_ENC_u0_N185, _AES_ENC_u0_N184, _AES_ENC_u0_N183, _AES_ENC_u0_N182, _AES_ENC_u0_N181, _AES_ENC_u0_N180, _AES_ENC_u0_N179, _AES_ENC_u0_N178, _AES_ENC_u0_N177, _AES_ENC_u0_N176, _AES_ENC_u0_N175, _AES_ENC_u0_N174, _AES_ENC_u0_N173, _AES_ENC_u0_N172, _AES_ENC_u0_N171, _AES_ENC_u0_N170, _AES_ENC_u0_N169, _AES_ENC_u0_N168, _AES_ENC_u0_N167, _AES_ENC_u0_N166, _AES_ENC_u0_N165, _AES_ENC_u0_N164, _AES_ENC_u0_N163, _AES_ENC_u0_N162, 
  _AES_ENC_u0_N161, _AES_ENC_u0_N160, _AES_ENC_u0_N159, _AES_ENC_u0_N158, _AES_ENC_u0_N157, _AES_ENC_u0_N156, _AES_ENC_u0_N155, _AES_ENC_u0_N154, _AES_ENC_u0_N153, _AES_ENC_u0_N152, _AES_ENC_u0_N151, _AES_ENC_u0_N150, _AES_ENC_u0_N149, _AES_ENC_u0_N148, _AES_ENC_u0_N147, _AES_ENC_u0_N146, _AES_ENC_u0_N145, _AES_ENC_u0_N144, _AES_ENC_u0_N143, _AES_ENC_u0_N142, _AES_ENC_u0_N139, _AES_ENC_u0_N138, _AES_ENC_u0_N137, _AES_ENC_u0_N136, _AES_ENC_u0_N135, _AES_ENC_u0_N134, _AES_ENC_u0_N133, _AES_ENC_u0_N132, _AES_ENC_u0_N131, _AES_ENC_u0_N130, _AES_ENC_u0_N129, _AES_ENC_u0_N128, _AES_ENC_u0_N127, _AES_ENC_u0_N126, _AES_ENC_u0_N125, _AES_ENC_u0_N124, _AES_ENC_u0_N123, _AES_ENC_u0_N122, _AES_ENC_u0_N121, _AES_ENC_u0_N120, _AES_ENC_u0_N119, _AES_ENC_u0_N118, _AES_ENC_u0_N117, _AES_ENC_u0_N116, _AES_ENC_u0_N115, _AES_ENC_u0_N114, _AES_ENC_u0_N113, _AES_ENC_u0_N112, _AES_ENC_u0_N111, _AES_ENC_u0_N110, 
  _AES_ENC_u0_N109, _AES_ENC_u0_N108, _AES_ENC_u0_N107, _AES_ENC_u0_N106, _AES_ENC_u0_N105, _AES_ENC_u0_N104, _AES_ENC_u0_N103, _AES_ENC_u0_N102, _AES_ENC_u0_N101, _AES_ENC_u0_N100, _AES_ENC_u0_N99, _AES_ENC_u0_N98, _AES_ENC_u0_N97, _AES_ENC_u0_N96, _AES_ENC_u0_N95, _AES_ENC_u0_N94, _AES_ENC_u0_N93, _AES_ENC_u0_N92, _AES_ENC_u0_N91, _AES_ENC_u0_N90, _AES_ENC_u0_N89, _AES_ENC_u0_N88, _AES_ENC_u0_N87, _AES_ENC_u0_N86, _AES_ENC_u0_N85, _AES_ENC_u0_N84, _AES_ENC_u0_N83, _AES_ENC_u0_N82, _AES_ENC_u0_N81, _AES_ENC_u0_N80, _AES_ENC_u0_N79, _AES_ENC_u0_N78, _AES_ENC_u0_N77, _AES_ENC_u0_N76, _AES_ENC_u0_N73, _AES_ENC_u0_N72, _AES_ENC_u0_N71, _AES_ENC_u0_N70, _AES_ENC_u0_N69, _AES_ENC_u0_N68, _AES_ENC_u0_N67, _AES_ENC_u0_N66, _AES_ENC_u0_N65, _AES_ENC_u0_N64, _AES_ENC_u0_N63, _AES_ENC_u0_N62, _AES_ENC_u0_N61, _AES_ENC_u0_N60, _AES_ENC_u0_N59, _AES_ENC_u0_N58, 
  _AES_ENC_u0_N57, _AES_ENC_u0_N56, _AES_ENC_u0_N55, _AES_ENC_u0_N54, _AES_ENC_u0_N53, _AES_ENC_u0_N52, _AES_ENC_u0_N51, _AES_ENC_u0_N50, _AES_ENC_u0_N49, _AES_ENC_u0_N48, _AES_ENC_u0_N47, _AES_ENC_u0_N46, _AES_ENC_u0_N45, _AES_ENC_u0_N44, _AES_ENC_u0_N43, _AES_ENC_u0_N42, _AES_ENC_u0_N17, _AES_ENC_u0_N16, _AES_ENC_u0_N15, _AES_ENC_u0_N14, _AES_ENC_u0_N13, _AES_ENC_u0_N12, _AES_ENC_u0_N11, _AES_ENC_u0_N10, _AES_ENC_u0_subword[0], _AES_ENC_u0_subword[1], _AES_ENC_u0_subword[2], _AES_ENC_u0_subword[3], _AES_ENC_u0_subword[4], _AES_ENC_u0_subword[5], _AES_ENC_u0_subword[6], _AES_ENC_u0_subword[7], _AES_ENC_u0_subword[8], _AES_ENC_u0_subword[9], _AES_ENC_u0_subword[10], _AES_ENC_u0_subword[11], _AES_ENC_u0_subword[12], _AES_ENC_u0_subword[13], _AES_ENC_u0_subword[14], _AES_ENC_u0_subword[15], _AES_ENC_u0_subword[16], _AES_ENC_u0_subword[17], _AES_ENC_u0_subword[18], _AES_ENC_u0_subword[19], _AES_ENC_u0_subword[20], _AES_ENC_u0_subword[21], _AES_ENC_u0_subword[22], _AES_ENC_u0_subword[23], _AES_ENC_u0_subword[24], _AES_ENC_u0_subword[25], 
  _AES_ENC_u0_subword[26], _AES_ENC_u0_subword[27], _AES_ENC_u0_subword[28], _AES_ENC_u0_subword[29], _AES_ENC_u0_subword[30], _AES_ENC_u0_subword[31], _AES_ENC_u0_u0_n1135, _AES_ENC_u0_u0_n1134, _AES_ENC_u0_u0_n1133, _AES_ENC_u0_u0_n1132, _AES_ENC_u0_u0_n1131, _AES_ENC_u0_u0_n1130, _AES_ENC_u0_u0_n1129, _AES_ENC_u0_u0_n1128, _AES_ENC_u0_u0_n1127, _AES_ENC_u0_u0_n1126, _AES_ENC_u0_u0_n1125, _AES_ENC_u0_u0_n1124, _AES_ENC_u0_u0_n1123, _AES_ENC_u0_u0_n1122, _AES_ENC_u0_u0_n1121, _AES_ENC_u0_u0_n1120, _AES_ENC_u0_u0_n1119, _AES_ENC_u0_u0_n1118, _AES_ENC_u0_u0_n1117, _AES_ENC_u0_u0_n1116, _AES_ENC_u0_u0_n1115, _AES_ENC_u0_u0_n1114, _AES_ENC_u0_u0_n1113, _AES_ENC_u0_u0_n1112, _AES_ENC_u0_u0_n1111, _AES_ENC_u0_u0_n1110, _AES_ENC_u0_u0_n1109, _AES_ENC_u0_u0_n1108, _AES_ENC_u0_u0_n1107, _AES_ENC_u0_u0_n1106, _AES_ENC_u0_u0_n1105, _AES_ENC_u0_u0_n1104, _AES_ENC_u0_u0_n1103, _AES_ENC_u0_u0_n1102, _AES_ENC_u0_u0_n1101, _AES_ENC_u0_u0_n1100, _AES_ENC_u0_u0_n1099, _AES_ENC_u0_u0_n1098, _AES_ENC_u0_u0_n1097, _AES_ENC_u0_u0_n1096, _AES_ENC_u0_u0_n1095, _AES_ENC_u0_u0_n1094, _AES_ENC_u0_u0_n1093, _AES_ENC_u0_u0_n1092, 
  _AES_ENC_u0_u0_n1091, _AES_ENC_u0_u0_n1090, _AES_ENC_u0_u0_n1089, _AES_ENC_u0_u0_n1088, _AES_ENC_u0_u0_n1087, _AES_ENC_u0_u0_n1086, _AES_ENC_u0_u0_n1085, _AES_ENC_u0_u0_n1084, _AES_ENC_u0_u0_n1083, _AES_ENC_u0_u0_n1082, _AES_ENC_u0_u0_n1081, _AES_ENC_u0_u0_n1080, _AES_ENC_u0_u0_n1079, _AES_ENC_u0_u0_n1078, _AES_ENC_u0_u0_n1077, _AES_ENC_u0_u0_n1076, _AES_ENC_u0_u0_n1075, _AES_ENC_u0_u0_n1074, _AES_ENC_u0_u0_n1073, _AES_ENC_u0_u0_n1072, _AES_ENC_u0_u0_n1071, _AES_ENC_u0_u0_n1070, _AES_ENC_u0_u0_n1069, _AES_ENC_u0_u0_n1068, _AES_ENC_u0_u0_n1067, _AES_ENC_u0_u0_n1066, _AES_ENC_u0_u0_n1065, _AES_ENC_u0_u0_n1064, _AES_ENC_u0_u0_n1063, _AES_ENC_u0_u0_n1062, _AES_ENC_u0_u0_n1061, _AES_ENC_u0_u0_n1060, _AES_ENC_u0_u0_n1059, _AES_ENC_u0_u0_n1058, _AES_ENC_u0_u0_n1057, _AES_ENC_u0_u0_n1056, _AES_ENC_u0_u0_n1055, _AES_ENC_u0_u0_n1054, _AES_ENC_u0_u0_n1053, _AES_ENC_u0_u0_n1052, _AES_ENC_u0_u0_n1051, _AES_ENC_u0_u0_n1050, _AES_ENC_u0_u0_n1049, _AES_ENC_u0_u0_n1048, _AES_ENC_u0_u0_n1047, _AES_ENC_u0_u0_n1046, _AES_ENC_u0_u0_n1045, _AES_ENC_u0_u0_n1044, _AES_ENC_u0_u0_n1043, _AES_ENC_u0_u0_n1042, 
  _AES_ENC_u0_u0_n1041, _AES_ENC_u0_u0_n1040, _AES_ENC_u0_u0_n1039, _AES_ENC_u0_u0_n1038, _AES_ENC_u0_u0_n1037, _AES_ENC_u0_u0_n1036, _AES_ENC_u0_u0_n1035, _AES_ENC_u0_u0_n1034, _AES_ENC_u0_u0_n1033, _AES_ENC_u0_u0_n1032, _AES_ENC_u0_u0_n1031, _AES_ENC_u0_u0_n1030, _AES_ENC_u0_u0_n1029, _AES_ENC_u0_u0_n1028, _AES_ENC_u0_u0_n1027, _AES_ENC_u0_u0_n1026, _AES_ENC_u0_u0_n1025, _AES_ENC_u0_u0_n1024, _AES_ENC_u0_u0_n1023, _AES_ENC_u0_u0_n1022, _AES_ENC_u0_u0_n1021, _AES_ENC_u0_u0_n1020, _AES_ENC_u0_u0_n1019, _AES_ENC_u0_u0_n1018, _AES_ENC_u0_u0_n1017, _AES_ENC_u0_u0_n1016, _AES_ENC_u0_u0_n1015, _AES_ENC_u0_u0_n1014, _AES_ENC_u0_u0_n1013, _AES_ENC_u0_u0_n1012, _AES_ENC_u0_u0_n1011, _AES_ENC_u0_u0_n1010, _AES_ENC_u0_u0_n1009, _AES_ENC_u0_u0_n1008, _AES_ENC_u0_u0_n1007, _AES_ENC_u0_u0_n1006, _AES_ENC_u0_u0_n1005, _AES_ENC_u0_u0_n1004, _AES_ENC_u0_u0_n1003, _AES_ENC_u0_u0_n1002, _AES_ENC_u0_u0_n1001, _AES_ENC_u0_u0_n1000, _AES_ENC_u0_u0_n999, _AES_ENC_u0_u0_n998, _AES_ENC_u0_u0_n997, _AES_ENC_u0_u0_n996, _AES_ENC_u0_u0_n995, _AES_ENC_u0_u0_n994, _AES_ENC_u0_u0_n993, _AES_ENC_u0_u0_n992, 
  _AES_ENC_u0_u0_n991, _AES_ENC_u0_u0_n990, _AES_ENC_u0_u0_n989, _AES_ENC_u0_u0_n988, _AES_ENC_u0_u0_n987, _AES_ENC_u0_u0_n986, _AES_ENC_u0_u0_n985, _AES_ENC_u0_u0_n984, _AES_ENC_u0_u0_n983, _AES_ENC_u0_u0_n982, _AES_ENC_u0_u0_n981, _AES_ENC_u0_u0_n980, _AES_ENC_u0_u0_n979, _AES_ENC_u0_u0_n978, _AES_ENC_u0_u0_n977, _AES_ENC_u0_u0_n976, _AES_ENC_u0_u0_n975, _AES_ENC_u0_u0_n974, _AES_ENC_u0_u0_n973, _AES_ENC_u0_u0_n972, _AES_ENC_u0_u0_n971, _AES_ENC_u0_u0_n970, _AES_ENC_u0_u0_n969, _AES_ENC_u0_u0_n968, _AES_ENC_u0_u0_n967, _AES_ENC_u0_u0_n966, _AES_ENC_u0_u0_n965, _AES_ENC_u0_u0_n964, _AES_ENC_u0_u0_n963, _AES_ENC_u0_u0_n962, _AES_ENC_u0_u0_n961, _AES_ENC_u0_u0_n960, _AES_ENC_u0_u0_n959, _AES_ENC_u0_u0_n958, _AES_ENC_u0_u0_n957, _AES_ENC_u0_u0_n956, _AES_ENC_u0_u0_n955, _AES_ENC_u0_u0_n954, _AES_ENC_u0_u0_n953, _AES_ENC_u0_u0_n952, _AES_ENC_u0_u0_n951, _AES_ENC_u0_u0_n950, _AES_ENC_u0_u0_n949, _AES_ENC_u0_u0_n948, _AES_ENC_u0_u0_n947, _AES_ENC_u0_u0_n946, _AES_ENC_u0_u0_n945, _AES_ENC_u0_u0_n944, _AES_ENC_u0_u0_n943, _AES_ENC_u0_u0_n942, 
  _AES_ENC_u0_u0_n941, _AES_ENC_u0_u0_n940, _AES_ENC_u0_u0_n939, _AES_ENC_u0_u0_n938, _AES_ENC_u0_u0_n937, _AES_ENC_u0_u0_n936, _AES_ENC_u0_u0_n935, _AES_ENC_u0_u0_n934, _AES_ENC_u0_u0_n933, _AES_ENC_u0_u0_n932, _AES_ENC_u0_u0_n931, _AES_ENC_u0_u0_n930, _AES_ENC_u0_u0_n929, _AES_ENC_u0_u0_n928, _AES_ENC_u0_u0_n927, _AES_ENC_u0_u0_n926, _AES_ENC_u0_u0_n925, _AES_ENC_u0_u0_n924, _AES_ENC_u0_u0_n923, _AES_ENC_u0_u0_n922, _AES_ENC_u0_u0_n921, _AES_ENC_u0_u0_n920, _AES_ENC_u0_u0_n919, _AES_ENC_u0_u0_n918, _AES_ENC_u0_u0_n917, _AES_ENC_u0_u0_n916, _AES_ENC_u0_u0_n915, _AES_ENC_u0_u0_n914, _AES_ENC_u0_u0_n913, _AES_ENC_u0_u0_n912, _AES_ENC_u0_u0_n911, _AES_ENC_u0_u0_n910, _AES_ENC_u0_u0_n909, _AES_ENC_u0_u0_n908, _AES_ENC_u0_u0_n907, _AES_ENC_u0_u0_n906, _AES_ENC_u0_u0_n905, _AES_ENC_u0_u0_n904, _AES_ENC_u0_u0_n903, _AES_ENC_u0_u0_n902, _AES_ENC_u0_u0_n901, _AES_ENC_u0_u0_n900, _AES_ENC_u0_u0_n899, _AES_ENC_u0_u0_n898, _AES_ENC_u0_u0_n897, _AES_ENC_u0_u0_n896, _AES_ENC_u0_u0_n895, _AES_ENC_u0_u0_n894, _AES_ENC_u0_u0_n893, _AES_ENC_u0_u0_n892, 
  _AES_ENC_u0_u0_n891, _AES_ENC_u0_u0_n890, _AES_ENC_u0_u0_n889, _AES_ENC_u0_u0_n888, _AES_ENC_u0_u0_n887, _AES_ENC_u0_u0_n886, _AES_ENC_u0_u0_n885, _AES_ENC_u0_u0_n884, _AES_ENC_u0_u0_n883, _AES_ENC_u0_u0_n882, _AES_ENC_u0_u0_n881, _AES_ENC_u0_u0_n880, _AES_ENC_u0_u0_n879, _AES_ENC_u0_u0_n878, _AES_ENC_u0_u0_n877, _AES_ENC_u0_u0_n876, _AES_ENC_u0_u0_n875, _AES_ENC_u0_u0_n874, _AES_ENC_u0_u0_n873, _AES_ENC_u0_u0_n872, _AES_ENC_u0_u0_n871, _AES_ENC_u0_u0_n870, _AES_ENC_u0_u0_n869, _AES_ENC_u0_u0_n868, _AES_ENC_u0_u0_n867, _AES_ENC_u0_u0_n866, _AES_ENC_u0_u0_n865, _AES_ENC_u0_u0_n864, _AES_ENC_u0_u0_n863, _AES_ENC_u0_u0_n862, _AES_ENC_u0_u0_n861, _AES_ENC_u0_u0_n860, _AES_ENC_u0_u0_n859, _AES_ENC_u0_u0_n858, _AES_ENC_u0_u0_n857, _AES_ENC_u0_u0_n856, _AES_ENC_u0_u0_n855, _AES_ENC_u0_u0_n854, _AES_ENC_u0_u0_n853, _AES_ENC_u0_u0_n852, _AES_ENC_u0_u0_n851, _AES_ENC_u0_u0_n850, _AES_ENC_u0_u0_n849, _AES_ENC_u0_u0_n848, _AES_ENC_u0_u0_n847, _AES_ENC_u0_u0_n846, _AES_ENC_u0_u0_n845, _AES_ENC_u0_u0_n844, _AES_ENC_u0_u0_n843, _AES_ENC_u0_u0_n842, 
  _AES_ENC_u0_u0_n841, _AES_ENC_u0_u0_n840, _AES_ENC_u0_u0_n839, _AES_ENC_u0_u0_n838, _AES_ENC_u0_u0_n837, _AES_ENC_u0_u0_n836, _AES_ENC_u0_u0_n835, _AES_ENC_u0_u0_n834, _AES_ENC_u0_u0_n833, _AES_ENC_u0_u0_n832, _AES_ENC_u0_u0_n831, _AES_ENC_u0_u0_n830, _AES_ENC_u0_u0_n829, _AES_ENC_u0_u0_n828, _AES_ENC_u0_u0_n827, _AES_ENC_u0_u0_n826, _AES_ENC_u0_u0_n825, _AES_ENC_u0_u0_n824, _AES_ENC_u0_u0_n823, _AES_ENC_u0_u0_n822, _AES_ENC_u0_u0_n821, _AES_ENC_u0_u0_n820, _AES_ENC_u0_u0_n819, _AES_ENC_u0_u0_n818, _AES_ENC_u0_u0_n817, _AES_ENC_u0_u0_n816, _AES_ENC_u0_u0_n815, _AES_ENC_u0_u0_n814, _AES_ENC_u0_u0_n813, _AES_ENC_u0_u0_n812, _AES_ENC_u0_u0_n811, _AES_ENC_u0_u0_n810, _AES_ENC_u0_u0_n809, _AES_ENC_u0_u0_n808, _AES_ENC_u0_u0_n807, _AES_ENC_u0_u0_n806, _AES_ENC_u0_u0_n805, _AES_ENC_u0_u0_n804, _AES_ENC_u0_u0_n803, _AES_ENC_u0_u0_n802, _AES_ENC_u0_u0_n801, _AES_ENC_u0_u0_n800, _AES_ENC_u0_u0_n799, _AES_ENC_u0_u0_n798, _AES_ENC_u0_u0_n797, _AES_ENC_u0_u0_n796, _AES_ENC_u0_u0_n795, _AES_ENC_u0_u0_n794, _AES_ENC_u0_u0_n793, _AES_ENC_u0_u0_n792, 
  _AES_ENC_u0_u0_n791, _AES_ENC_u0_u0_n790, _AES_ENC_u0_u0_n789, _AES_ENC_u0_u0_n788, _AES_ENC_u0_u0_n787, _AES_ENC_u0_u0_n786, _AES_ENC_u0_u0_n785, _AES_ENC_u0_u0_n784, _AES_ENC_u0_u0_n783, _AES_ENC_u0_u0_n782, _AES_ENC_u0_u0_n781, _AES_ENC_u0_u0_n780, _AES_ENC_u0_u0_n779, _AES_ENC_u0_u0_n778, _AES_ENC_u0_u0_n777, _AES_ENC_u0_u0_n776, _AES_ENC_u0_u0_n775, _AES_ENC_u0_u0_n774, _AES_ENC_u0_u0_n773, _AES_ENC_u0_u0_n772, _AES_ENC_u0_u0_n771, _AES_ENC_u0_u0_n770, _AES_ENC_u0_u0_n769, _AES_ENC_u0_u0_n768, _AES_ENC_u0_u0_n767, _AES_ENC_u0_u0_n766, _AES_ENC_u0_u0_n765, _AES_ENC_u0_u0_n764, _AES_ENC_u0_u0_n763, _AES_ENC_u0_u0_n762, _AES_ENC_u0_u0_n761, _AES_ENC_u0_u0_n760, _AES_ENC_u0_u0_n759, _AES_ENC_u0_u0_n758, _AES_ENC_u0_u0_n757, _AES_ENC_u0_u0_n756, _AES_ENC_u0_u0_n755, _AES_ENC_u0_u0_n754, _AES_ENC_u0_u0_n753, _AES_ENC_u0_u0_n752, _AES_ENC_u0_u0_n751, _AES_ENC_u0_u0_n750, _AES_ENC_u0_u0_n749, _AES_ENC_u0_u0_n748, _AES_ENC_u0_u0_n747, _AES_ENC_u0_u0_n746, _AES_ENC_u0_u0_n745, _AES_ENC_u0_u0_n744, _AES_ENC_u0_u0_n743, _AES_ENC_u0_u0_n742, 
  _AES_ENC_u0_u0_n741, _AES_ENC_u0_u0_n740, _AES_ENC_u0_u0_n739, _AES_ENC_u0_u0_n738, _AES_ENC_u0_u0_n737, _AES_ENC_u0_u0_n736, _AES_ENC_u0_u0_n735, _AES_ENC_u0_u0_n734, _AES_ENC_u0_u0_n733, _AES_ENC_u0_u0_n732, _AES_ENC_u0_u0_n731, _AES_ENC_u0_u0_n730, _AES_ENC_u0_u0_n729, _AES_ENC_u0_u0_n728, _AES_ENC_u0_u0_n727, _AES_ENC_u0_u0_n726, _AES_ENC_u0_u0_n725, _AES_ENC_u0_u0_n724, _AES_ENC_u0_u0_n723, _AES_ENC_u0_u0_n722, _AES_ENC_u0_u0_n721, _AES_ENC_u0_u0_n720, _AES_ENC_u0_u0_n719, _AES_ENC_u0_u0_n718, _AES_ENC_u0_u0_n717, _AES_ENC_u0_u0_n716, _AES_ENC_u0_u0_n715, _AES_ENC_u0_u0_n714, _AES_ENC_u0_u0_n713, _AES_ENC_u0_u0_n712, _AES_ENC_u0_u0_n711, _AES_ENC_u0_u0_n710, _AES_ENC_u0_u0_n709, _AES_ENC_u0_u0_n708, _AES_ENC_u0_u0_n707, _AES_ENC_u0_u0_n706, _AES_ENC_u0_u0_n705, _AES_ENC_u0_u0_n704, _AES_ENC_u0_u0_n703, _AES_ENC_u0_u0_n702, _AES_ENC_u0_u0_n701, _AES_ENC_u0_u0_n700, _AES_ENC_u0_u0_n699, _AES_ENC_u0_u0_n698, _AES_ENC_u0_u0_n697, _AES_ENC_u0_u0_n696, _AES_ENC_u0_u0_n695, _AES_ENC_u0_u0_n694, _AES_ENC_u0_u0_n693, _AES_ENC_u0_u0_n692, 
  _AES_ENC_u0_u0_n691, _AES_ENC_u0_u0_n690, _AES_ENC_u0_u0_n689, _AES_ENC_u0_u0_n688, _AES_ENC_u0_u0_n687, _AES_ENC_u0_u0_n686, _AES_ENC_u0_u0_n685, _AES_ENC_u0_u0_n684, _AES_ENC_u0_u0_n683, _AES_ENC_u0_u0_n682, _AES_ENC_u0_u0_n681, _AES_ENC_u0_u0_n680, _AES_ENC_u0_u0_n679, _AES_ENC_u0_u0_n678, _AES_ENC_u0_u0_n677, _AES_ENC_u0_u0_n676, _AES_ENC_u0_u0_n675, _AES_ENC_u0_u0_n674, _AES_ENC_u0_u0_n673, _AES_ENC_u0_u0_n672, _AES_ENC_u0_u0_n671, _AES_ENC_u0_u0_n670, _AES_ENC_u0_u0_n669, _AES_ENC_u0_u0_n668, _AES_ENC_u0_u0_n667, _AES_ENC_u0_u0_n666, _AES_ENC_u0_u0_n665, _AES_ENC_u0_u0_n664, _AES_ENC_u0_u0_n663, _AES_ENC_u0_u0_n662, _AES_ENC_u0_u0_n661, _AES_ENC_u0_u0_n660, _AES_ENC_u0_u0_n659, _AES_ENC_u0_u0_n658, _AES_ENC_u0_u0_n657, _AES_ENC_u0_u0_n656, _AES_ENC_u0_u0_n655, _AES_ENC_u0_u0_n654, _AES_ENC_u0_u0_n653, _AES_ENC_u0_u0_n652, _AES_ENC_u0_u0_n651, _AES_ENC_u0_u0_n650, _AES_ENC_u0_u0_n649, _AES_ENC_u0_u0_n648, _AES_ENC_u0_u0_n647, _AES_ENC_u0_u0_n646, _AES_ENC_u0_u0_n645, _AES_ENC_u0_u0_n644, _AES_ENC_u0_u0_n643, _AES_ENC_u0_u0_n642, 
  _AES_ENC_u0_u0_n641, _AES_ENC_u0_u0_n640, _AES_ENC_u0_u0_n639, _AES_ENC_u0_u0_n638, _AES_ENC_u0_u0_n637, _AES_ENC_u0_u0_n636, _AES_ENC_u0_u0_n635, _AES_ENC_u0_u0_n634, _AES_ENC_u0_u0_n633, _AES_ENC_u0_u0_n632, _AES_ENC_u0_u0_n631, _AES_ENC_u0_u0_n630, _AES_ENC_u0_u0_n629, _AES_ENC_u0_u0_n628, _AES_ENC_u0_u0_n627, _AES_ENC_u0_u0_n626, _AES_ENC_u0_u0_n625, _AES_ENC_u0_u0_n624, _AES_ENC_u0_u0_n623, _AES_ENC_u0_u0_n622, _AES_ENC_u0_u0_n621, _AES_ENC_u0_u0_n620, _AES_ENC_u0_u0_n619, _AES_ENC_u0_u0_n618, _AES_ENC_u0_u0_n617, _AES_ENC_u0_u0_n616, _AES_ENC_u0_u0_n615, _AES_ENC_u0_u0_n614, _AES_ENC_u0_u0_n613, _AES_ENC_u0_u0_n612, _AES_ENC_u0_u0_n611, _AES_ENC_u0_u0_n610, _AES_ENC_u0_u0_n609, _AES_ENC_u0_u0_n608, _AES_ENC_u0_u0_n607, _AES_ENC_u0_u0_n606, _AES_ENC_u0_u0_n605, _AES_ENC_u0_u0_n604, _AES_ENC_u0_u0_n603, _AES_ENC_u0_u0_n602, _AES_ENC_u0_u0_n601, _AES_ENC_u0_u0_n600, _AES_ENC_u0_u0_n599, _AES_ENC_u0_u0_n598, _AES_ENC_u0_u0_n597, _AES_ENC_u0_u0_n596, _AES_ENC_u0_u0_n595, _AES_ENC_u0_u0_n594, _AES_ENC_u0_u0_n593, _AES_ENC_u0_u0_n592, 
  _AES_ENC_u0_u0_n591, _AES_ENC_u0_u0_n590, _AES_ENC_u0_u0_n589, _AES_ENC_u0_u0_n588, _AES_ENC_u0_u0_n587, _AES_ENC_u0_u0_n586, _AES_ENC_u0_u0_n585, _AES_ENC_u0_u0_n584, _AES_ENC_u0_u0_n583, _AES_ENC_u0_u0_n582, _AES_ENC_u0_u0_n581, _AES_ENC_u0_u0_n580, _AES_ENC_u0_u0_n579, _AES_ENC_u0_u0_n578, _AES_ENC_u0_u0_n577, _AES_ENC_u0_u0_n576, _AES_ENC_u0_u0_n575, _AES_ENC_u0_u0_n574, _AES_ENC_u0_u0_n573, _AES_ENC_u0_u0_n572, _AES_ENC_u0_u0_n571, _AES_ENC_u0_u0_n570, _AES_ENC_u0_u0_n569, _AES_ENC_u0_u1_n1135, _AES_ENC_u0_u1_n1134, _AES_ENC_u0_u1_n1133, _AES_ENC_u0_u1_n1132, _AES_ENC_u0_u1_n1131, _AES_ENC_u0_u1_n1130, _AES_ENC_u0_u1_n1129, _AES_ENC_u0_u1_n1128, _AES_ENC_u0_u1_n1127, _AES_ENC_u0_u1_n1126, _AES_ENC_u0_u1_n1125, _AES_ENC_u0_u1_n1124, _AES_ENC_u0_u1_n1123, _AES_ENC_u0_u1_n1122, _AES_ENC_u0_u1_n1121, _AES_ENC_u0_u1_n1120, _AES_ENC_u0_u1_n1119, _AES_ENC_u0_u1_n1118, _AES_ENC_u0_u1_n1117, _AES_ENC_u0_u1_n1116, _AES_ENC_u0_u1_n1115, _AES_ENC_u0_u1_n1114, _AES_ENC_u0_u1_n1113, _AES_ENC_u0_u1_n1112, _AES_ENC_u0_u1_n1111, _AES_ENC_u0_u1_n1110, _AES_ENC_u0_u1_n1109, 
  _AES_ENC_u0_u1_n1108, _AES_ENC_u0_u1_n1107, _AES_ENC_u0_u1_n1106, _AES_ENC_u0_u1_n1105, _AES_ENC_u0_u1_n1104, _AES_ENC_u0_u1_n1103, _AES_ENC_u0_u1_n1102, _AES_ENC_u0_u1_n1101, _AES_ENC_u0_u1_n1100, _AES_ENC_u0_u1_n1099, _AES_ENC_u0_u1_n1098, _AES_ENC_u0_u1_n1097, _AES_ENC_u0_u1_n1096, _AES_ENC_u0_u1_n1095, _AES_ENC_u0_u1_n1094, _AES_ENC_u0_u1_n1093, _AES_ENC_u0_u1_n1092, _AES_ENC_u0_u1_n1091, _AES_ENC_u0_u1_n1090, _AES_ENC_u0_u1_n1089, _AES_ENC_u0_u1_n1088, _AES_ENC_u0_u1_n1087, _AES_ENC_u0_u1_n1086, _AES_ENC_u0_u1_n1085, _AES_ENC_u0_u1_n1084, _AES_ENC_u0_u1_n1083, _AES_ENC_u0_u1_n1082, _AES_ENC_u0_u1_n1081, _AES_ENC_u0_u1_n1080, _AES_ENC_u0_u1_n1079, _AES_ENC_u0_u1_n1078, _AES_ENC_u0_u1_n1077, _AES_ENC_u0_u1_n1076, _AES_ENC_u0_u1_n1075, _AES_ENC_u0_u1_n1074, _AES_ENC_u0_u1_n1073, _AES_ENC_u0_u1_n1072, _AES_ENC_u0_u1_n1071, _AES_ENC_u0_u1_n1070, _AES_ENC_u0_u1_n1069, _AES_ENC_u0_u1_n1068, _AES_ENC_u0_u1_n1067, _AES_ENC_u0_u1_n1066, _AES_ENC_u0_u1_n1065, _AES_ENC_u0_u1_n1064, _AES_ENC_u0_u1_n1063, _AES_ENC_u0_u1_n1062, _AES_ENC_u0_u1_n1061, _AES_ENC_u0_u1_n1060, _AES_ENC_u0_u1_n1059, 
  _AES_ENC_u0_u1_n1058, _AES_ENC_u0_u1_n1057, _AES_ENC_u0_u1_n1056, _AES_ENC_u0_u1_n1055, _AES_ENC_u0_u1_n1054, _AES_ENC_u0_u1_n1053, _AES_ENC_u0_u1_n1052, _AES_ENC_u0_u1_n1051, _AES_ENC_u0_u1_n1050, _AES_ENC_u0_u1_n1049, _AES_ENC_u0_u1_n1048, _AES_ENC_u0_u1_n1047, _AES_ENC_u0_u1_n1046, _AES_ENC_u0_u1_n1045, _AES_ENC_u0_u1_n1044, _AES_ENC_u0_u1_n1043, _AES_ENC_u0_u1_n1042, _AES_ENC_u0_u1_n1041, _AES_ENC_u0_u1_n1040, _AES_ENC_u0_u1_n1039, _AES_ENC_u0_u1_n1038, _AES_ENC_u0_u1_n1037, _AES_ENC_u0_u1_n1036, _AES_ENC_u0_u1_n1035, _AES_ENC_u0_u1_n1034, _AES_ENC_u0_u1_n1033, _AES_ENC_u0_u1_n1032, _AES_ENC_u0_u1_n1031, _AES_ENC_u0_u1_n1030, _AES_ENC_u0_u1_n1029, _AES_ENC_u0_u1_n1028, _AES_ENC_u0_u1_n1027, _AES_ENC_u0_u1_n1026, _AES_ENC_u0_u1_n1025, _AES_ENC_u0_u1_n1024, _AES_ENC_u0_u1_n1023, _AES_ENC_u0_u1_n1022, _AES_ENC_u0_u1_n1021, _AES_ENC_u0_u1_n1020, _AES_ENC_u0_u1_n1019, _AES_ENC_u0_u1_n1018, _AES_ENC_u0_u1_n1017, _AES_ENC_u0_u1_n1016, _AES_ENC_u0_u1_n1015, _AES_ENC_u0_u1_n1014, _AES_ENC_u0_u1_n1013, _AES_ENC_u0_u1_n1012, _AES_ENC_u0_u1_n1011, _AES_ENC_u0_u1_n1010, _AES_ENC_u0_u1_n1009, 
  _AES_ENC_u0_u1_n1008, _AES_ENC_u0_u1_n1007, _AES_ENC_u0_u1_n1006, _AES_ENC_u0_u1_n1005, _AES_ENC_u0_u1_n1004, _AES_ENC_u0_u1_n1003, _AES_ENC_u0_u1_n1002, _AES_ENC_u0_u1_n1001, _AES_ENC_u0_u1_n1000, _AES_ENC_u0_u1_n999, _AES_ENC_u0_u1_n998, _AES_ENC_u0_u1_n997, _AES_ENC_u0_u1_n996, _AES_ENC_u0_u1_n995, _AES_ENC_u0_u1_n994, _AES_ENC_u0_u1_n993, _AES_ENC_u0_u1_n992, _AES_ENC_u0_u1_n991, _AES_ENC_u0_u1_n990, _AES_ENC_u0_u1_n989, _AES_ENC_u0_u1_n988, _AES_ENC_u0_u1_n987, _AES_ENC_u0_u1_n986, _AES_ENC_u0_u1_n985, _AES_ENC_u0_u1_n984, _AES_ENC_u0_u1_n983, _AES_ENC_u0_u1_n982, _AES_ENC_u0_u1_n981, _AES_ENC_u0_u1_n980, _AES_ENC_u0_u1_n979, _AES_ENC_u0_u1_n978, _AES_ENC_u0_u1_n977, _AES_ENC_u0_u1_n976, _AES_ENC_u0_u1_n975, _AES_ENC_u0_u1_n974, _AES_ENC_u0_u1_n973, _AES_ENC_u0_u1_n972, _AES_ENC_u0_u1_n971, _AES_ENC_u0_u1_n970, _AES_ENC_u0_u1_n969, _AES_ENC_u0_u1_n968, _AES_ENC_u0_u1_n967, _AES_ENC_u0_u1_n966, _AES_ENC_u0_u1_n965, _AES_ENC_u0_u1_n964, _AES_ENC_u0_u1_n963, _AES_ENC_u0_u1_n962, _AES_ENC_u0_u1_n961, _AES_ENC_u0_u1_n960, _AES_ENC_u0_u1_n959, 
  _AES_ENC_u0_u1_n958, _AES_ENC_u0_u1_n957, _AES_ENC_u0_u1_n956, _AES_ENC_u0_u1_n955, _AES_ENC_u0_u1_n954, _AES_ENC_u0_u1_n953, _AES_ENC_u0_u1_n952, _AES_ENC_u0_u1_n951, _AES_ENC_u0_u1_n950, _AES_ENC_u0_u1_n949, _AES_ENC_u0_u1_n948, _AES_ENC_u0_u1_n947, _AES_ENC_u0_u1_n946, _AES_ENC_u0_u1_n945, _AES_ENC_u0_u1_n944, _AES_ENC_u0_u1_n943, _AES_ENC_u0_u1_n942, _AES_ENC_u0_u1_n941, _AES_ENC_u0_u1_n940, _AES_ENC_u0_u1_n939, _AES_ENC_u0_u1_n938, _AES_ENC_u0_u1_n937, _AES_ENC_u0_u1_n936, _AES_ENC_u0_u1_n935, _AES_ENC_u0_u1_n934, _AES_ENC_u0_u1_n933, _AES_ENC_u0_u1_n932, _AES_ENC_u0_u1_n931, _AES_ENC_u0_u1_n930, _AES_ENC_u0_u1_n929, _AES_ENC_u0_u1_n928, _AES_ENC_u0_u1_n927, _AES_ENC_u0_u1_n926, _AES_ENC_u0_u1_n925, _AES_ENC_u0_u1_n924, _AES_ENC_u0_u1_n923, _AES_ENC_u0_u1_n922, _AES_ENC_u0_u1_n921, _AES_ENC_u0_u1_n920, _AES_ENC_u0_u1_n919, _AES_ENC_u0_u1_n918, _AES_ENC_u0_u1_n917, _AES_ENC_u0_u1_n916, _AES_ENC_u0_u1_n915, _AES_ENC_u0_u1_n914, _AES_ENC_u0_u1_n913, _AES_ENC_u0_u1_n912, _AES_ENC_u0_u1_n911, _AES_ENC_u0_u1_n910, _AES_ENC_u0_u1_n909, 
  _AES_ENC_u0_u1_n908, _AES_ENC_u0_u1_n907, _AES_ENC_u0_u1_n906, _AES_ENC_u0_u1_n905, _AES_ENC_u0_u1_n904, _AES_ENC_u0_u1_n903, _AES_ENC_u0_u1_n902, _AES_ENC_u0_u1_n901, _AES_ENC_u0_u1_n900, _AES_ENC_u0_u1_n899, _AES_ENC_u0_u1_n898, _AES_ENC_u0_u1_n897, _AES_ENC_u0_u1_n896, _AES_ENC_u0_u1_n895, _AES_ENC_u0_u1_n894, _AES_ENC_u0_u1_n893, _AES_ENC_u0_u1_n892, _AES_ENC_u0_u1_n891, _AES_ENC_u0_u1_n890, _AES_ENC_u0_u1_n889, _AES_ENC_u0_u1_n888, _AES_ENC_u0_u1_n887, _AES_ENC_u0_u1_n886, _AES_ENC_u0_u1_n885, _AES_ENC_u0_u1_n884, _AES_ENC_u0_u1_n883, _AES_ENC_u0_u1_n882, _AES_ENC_u0_u1_n881, _AES_ENC_u0_u1_n880, _AES_ENC_u0_u1_n879, _AES_ENC_u0_u1_n878, _AES_ENC_u0_u1_n877, _AES_ENC_u0_u1_n876, _AES_ENC_u0_u1_n875, _AES_ENC_u0_u1_n874, _AES_ENC_u0_u1_n873, _AES_ENC_u0_u1_n872, _AES_ENC_u0_u1_n871, _AES_ENC_u0_u1_n870, _AES_ENC_u0_u1_n869, _AES_ENC_u0_u1_n868, _AES_ENC_u0_u1_n867, _AES_ENC_u0_u1_n866, _AES_ENC_u0_u1_n865, _AES_ENC_u0_u1_n864, _AES_ENC_u0_u1_n863, _AES_ENC_u0_u1_n862, _AES_ENC_u0_u1_n861, _AES_ENC_u0_u1_n860, _AES_ENC_u0_u1_n859, 
  _AES_ENC_u0_u1_n858, _AES_ENC_u0_u1_n857, _AES_ENC_u0_u1_n856, _AES_ENC_u0_u1_n855, _AES_ENC_u0_u1_n854, _AES_ENC_u0_u1_n853, _AES_ENC_u0_u1_n852, _AES_ENC_u0_u1_n851, _AES_ENC_u0_u1_n850, _AES_ENC_u0_u1_n849, _AES_ENC_u0_u1_n848, _AES_ENC_u0_u1_n847, _AES_ENC_u0_u1_n846, _AES_ENC_u0_u1_n845, _AES_ENC_u0_u1_n844, _AES_ENC_u0_u1_n843, _AES_ENC_u0_u1_n842, _AES_ENC_u0_u1_n841, _AES_ENC_u0_u1_n840, _AES_ENC_u0_u1_n839, _AES_ENC_u0_u1_n838, _AES_ENC_u0_u1_n837, _AES_ENC_u0_u1_n836, _AES_ENC_u0_u1_n835, _AES_ENC_u0_u1_n834, _AES_ENC_u0_u1_n833, _AES_ENC_u0_u1_n832, _AES_ENC_u0_u1_n831, _AES_ENC_u0_u1_n830, _AES_ENC_u0_u1_n829, _AES_ENC_u0_u1_n828, _AES_ENC_u0_u1_n827, _AES_ENC_u0_u1_n826, _AES_ENC_u0_u1_n825, _AES_ENC_u0_u1_n824, _AES_ENC_u0_u1_n823, _AES_ENC_u0_u1_n822, _AES_ENC_u0_u1_n821, _AES_ENC_u0_u1_n820, _AES_ENC_u0_u1_n819, _AES_ENC_u0_u1_n818, _AES_ENC_u0_u1_n817, _AES_ENC_u0_u1_n816, _AES_ENC_u0_u1_n815, _AES_ENC_u0_u1_n814, _AES_ENC_u0_u1_n813, _AES_ENC_u0_u1_n812, _AES_ENC_u0_u1_n811, _AES_ENC_u0_u1_n810, _AES_ENC_u0_u1_n809, 
  _AES_ENC_u0_u1_n808, _AES_ENC_u0_u1_n807, _AES_ENC_u0_u1_n806, _AES_ENC_u0_u1_n805, _AES_ENC_u0_u1_n804, _AES_ENC_u0_u1_n803, _AES_ENC_u0_u1_n802, _AES_ENC_u0_u1_n801, _AES_ENC_u0_u1_n800, _AES_ENC_u0_u1_n799, _AES_ENC_u0_u1_n798, _AES_ENC_u0_u1_n797, _AES_ENC_u0_u1_n796, _AES_ENC_u0_u1_n795, _AES_ENC_u0_u1_n794, _AES_ENC_u0_u1_n793, _AES_ENC_u0_u1_n792, _AES_ENC_u0_u1_n791, _AES_ENC_u0_u1_n790, _AES_ENC_u0_u1_n789, _AES_ENC_u0_u1_n788, _AES_ENC_u0_u1_n787, _AES_ENC_u0_u1_n786, _AES_ENC_u0_u1_n785, _AES_ENC_u0_u1_n784, _AES_ENC_u0_u1_n783, _AES_ENC_u0_u1_n782, _AES_ENC_u0_u1_n781, _AES_ENC_u0_u1_n780, _AES_ENC_u0_u1_n779, _AES_ENC_u0_u1_n778, _AES_ENC_u0_u1_n777, _AES_ENC_u0_u1_n776, _AES_ENC_u0_u1_n775, _AES_ENC_u0_u1_n774, _AES_ENC_u0_u1_n773, _AES_ENC_u0_u1_n772, _AES_ENC_u0_u1_n771, _AES_ENC_u0_u1_n770, _AES_ENC_u0_u1_n769, _AES_ENC_u0_u1_n768, _AES_ENC_u0_u1_n767, _AES_ENC_u0_u1_n766, _AES_ENC_u0_u1_n765, _AES_ENC_u0_u1_n764, _AES_ENC_u0_u1_n763, _AES_ENC_u0_u1_n762, _AES_ENC_u0_u1_n761, _AES_ENC_u0_u1_n760, _AES_ENC_u0_u1_n759, 
  _AES_ENC_u0_u1_n758, _AES_ENC_u0_u1_n757, _AES_ENC_u0_u1_n756, _AES_ENC_u0_u1_n755, _AES_ENC_u0_u1_n754, _AES_ENC_u0_u1_n753, _AES_ENC_u0_u1_n752, _AES_ENC_u0_u1_n751, _AES_ENC_u0_u1_n750, _AES_ENC_u0_u1_n749, _AES_ENC_u0_u1_n748, _AES_ENC_u0_u1_n747, _AES_ENC_u0_u1_n746, _AES_ENC_u0_u1_n745, _AES_ENC_u0_u1_n744, _AES_ENC_u0_u1_n743, _AES_ENC_u0_u1_n742, _AES_ENC_u0_u1_n741, _AES_ENC_u0_u1_n740, _AES_ENC_u0_u1_n739, _AES_ENC_u0_u1_n738, _AES_ENC_u0_u1_n737, _AES_ENC_u0_u1_n736, _AES_ENC_u0_u1_n735, _AES_ENC_u0_u1_n734, _AES_ENC_u0_u1_n733, _AES_ENC_u0_u1_n732, _AES_ENC_u0_u1_n731, _AES_ENC_u0_u1_n730, _AES_ENC_u0_u1_n729, _AES_ENC_u0_u1_n728, _AES_ENC_u0_u1_n727, _AES_ENC_u0_u1_n726, _AES_ENC_u0_u1_n725, _AES_ENC_u0_u1_n724, _AES_ENC_u0_u1_n723, _AES_ENC_u0_u1_n722, _AES_ENC_u0_u1_n721, _AES_ENC_u0_u1_n720, _AES_ENC_u0_u1_n719, _AES_ENC_u0_u1_n718, _AES_ENC_u0_u1_n717, _AES_ENC_u0_u1_n716, _AES_ENC_u0_u1_n715, _AES_ENC_u0_u1_n714, _AES_ENC_u0_u1_n713, _AES_ENC_u0_u1_n712, _AES_ENC_u0_u1_n711, _AES_ENC_u0_u1_n710, _AES_ENC_u0_u1_n709, 
  _AES_ENC_u0_u1_n708, _AES_ENC_u0_u1_n707, _AES_ENC_u0_u1_n706, _AES_ENC_u0_u1_n705, _AES_ENC_u0_u1_n704, _AES_ENC_u0_u1_n703, _AES_ENC_u0_u1_n702, _AES_ENC_u0_u1_n701, _AES_ENC_u0_u1_n700, _AES_ENC_u0_u1_n699, _AES_ENC_u0_u1_n698, _AES_ENC_u0_u1_n697, _AES_ENC_u0_u1_n696, _AES_ENC_u0_u1_n695, _AES_ENC_u0_u1_n694, _AES_ENC_u0_u1_n693, _AES_ENC_u0_u1_n692, _AES_ENC_u0_u1_n691, _AES_ENC_u0_u1_n690, _AES_ENC_u0_u1_n689, _AES_ENC_u0_u1_n688, _AES_ENC_u0_u1_n687, _AES_ENC_u0_u1_n686, _AES_ENC_u0_u1_n685, _AES_ENC_u0_u1_n684, _AES_ENC_u0_u1_n683, _AES_ENC_u0_u1_n682, _AES_ENC_u0_u1_n681, _AES_ENC_u0_u1_n680, _AES_ENC_u0_u1_n679, _AES_ENC_u0_u1_n678, _AES_ENC_u0_u1_n677, _AES_ENC_u0_u1_n676, _AES_ENC_u0_u1_n675, _AES_ENC_u0_u1_n674, _AES_ENC_u0_u1_n673, _AES_ENC_u0_u1_n672, _AES_ENC_u0_u1_n671, _AES_ENC_u0_u1_n670, _AES_ENC_u0_u1_n669, _AES_ENC_u0_u1_n668, _AES_ENC_u0_u1_n667, _AES_ENC_u0_u1_n666, _AES_ENC_u0_u1_n665, _AES_ENC_u0_u1_n664, _AES_ENC_u0_u1_n663, _AES_ENC_u0_u1_n662, _AES_ENC_u0_u1_n661, _AES_ENC_u0_u1_n660, _AES_ENC_u0_u1_n659, 
  _AES_ENC_u0_u1_n658, _AES_ENC_u0_u1_n657, _AES_ENC_u0_u1_n656, _AES_ENC_u0_u1_n655, _AES_ENC_u0_u1_n654, _AES_ENC_u0_u1_n653, _AES_ENC_u0_u1_n652, _AES_ENC_u0_u1_n651, _AES_ENC_u0_u1_n650, _AES_ENC_u0_u1_n649, _AES_ENC_u0_u1_n648, _AES_ENC_u0_u1_n647, _AES_ENC_u0_u1_n646, _AES_ENC_u0_u1_n645, _AES_ENC_u0_u1_n644, _AES_ENC_u0_u1_n643, _AES_ENC_u0_u1_n642, _AES_ENC_u0_u1_n641, _AES_ENC_u0_u1_n640, _AES_ENC_u0_u1_n639, _AES_ENC_u0_u1_n638, _AES_ENC_u0_u1_n637, _AES_ENC_u0_u1_n636, _AES_ENC_u0_u1_n635, _AES_ENC_u0_u1_n634, _AES_ENC_u0_u1_n633, _AES_ENC_u0_u1_n632, _AES_ENC_u0_u1_n631, _AES_ENC_u0_u1_n630, _AES_ENC_u0_u1_n629, _AES_ENC_u0_u1_n628, _AES_ENC_u0_u1_n627, _AES_ENC_u0_u1_n626, _AES_ENC_u0_u1_n625, _AES_ENC_u0_u1_n624, _AES_ENC_u0_u1_n623, _AES_ENC_u0_u1_n622, _AES_ENC_u0_u1_n621, _AES_ENC_u0_u1_n620, _AES_ENC_u0_u1_n619, _AES_ENC_u0_u1_n618, _AES_ENC_u0_u1_n617, _AES_ENC_u0_u1_n616, _AES_ENC_u0_u1_n615, _AES_ENC_u0_u1_n614, _AES_ENC_u0_u1_n613, _AES_ENC_u0_u1_n612, _AES_ENC_u0_u1_n611, _AES_ENC_u0_u1_n610, _AES_ENC_u0_u1_n609, 
  _AES_ENC_u0_u1_n608, _AES_ENC_u0_u1_n607, _AES_ENC_u0_u1_n606, _AES_ENC_u0_u1_n605, _AES_ENC_u0_u1_n604, _AES_ENC_u0_u1_n603, _AES_ENC_u0_u1_n602, _AES_ENC_u0_u1_n601, _AES_ENC_u0_u1_n600, _AES_ENC_u0_u1_n599, _AES_ENC_u0_u1_n598, _AES_ENC_u0_u1_n597, _AES_ENC_u0_u1_n596, _AES_ENC_u0_u1_n595, _AES_ENC_u0_u1_n594, _AES_ENC_u0_u1_n593, _AES_ENC_u0_u1_n592, _AES_ENC_u0_u1_n591, _AES_ENC_u0_u1_n590, _AES_ENC_u0_u1_n589, _AES_ENC_u0_u1_n588, _AES_ENC_u0_u1_n587, _AES_ENC_u0_u1_n586, _AES_ENC_u0_u1_n585, _AES_ENC_u0_u1_n584, _AES_ENC_u0_u1_n583, _AES_ENC_u0_u1_n582, _AES_ENC_u0_u1_n581, _AES_ENC_u0_u1_n580, _AES_ENC_u0_u1_n579, _AES_ENC_u0_u1_n578, _AES_ENC_u0_u1_n577, _AES_ENC_u0_u1_n576, _AES_ENC_u0_u1_n575, _AES_ENC_u0_u1_n574, _AES_ENC_u0_u1_n573, _AES_ENC_u0_u1_n572, _AES_ENC_u0_u1_n571, _AES_ENC_u0_u1_n570, _AES_ENC_u0_u1_n569, _AES_ENC_u0_u2_n1135, _AES_ENC_u0_u2_n1134, _AES_ENC_u0_u2_n1133, _AES_ENC_u0_u2_n1132, _AES_ENC_u0_u2_n1131, _AES_ENC_u0_u2_n1130, _AES_ENC_u0_u2_n1129, _AES_ENC_u0_u2_n1128, _AES_ENC_u0_u2_n1127, _AES_ENC_u0_u2_n1126, 
  _AES_ENC_u0_u2_n1125, _AES_ENC_u0_u2_n1124, _AES_ENC_u0_u2_n1123, _AES_ENC_u0_u2_n1122, _AES_ENC_u0_u2_n1121, _AES_ENC_u0_u2_n1120, _AES_ENC_u0_u2_n1119, _AES_ENC_u0_u2_n1118, _AES_ENC_u0_u2_n1117, _AES_ENC_u0_u2_n1116, _AES_ENC_u0_u2_n1115, _AES_ENC_u0_u2_n1114, _AES_ENC_u0_u2_n1113, _AES_ENC_u0_u2_n1112, _AES_ENC_u0_u2_n1111, _AES_ENC_u0_u2_n1110, _AES_ENC_u0_u2_n1109, _AES_ENC_u0_u2_n1108, _AES_ENC_u0_u2_n1107, _AES_ENC_u0_u2_n1106, _AES_ENC_u0_u2_n1105, _AES_ENC_u0_u2_n1104, _AES_ENC_u0_u2_n1103, _AES_ENC_u0_u2_n1102, _AES_ENC_u0_u2_n1101, _AES_ENC_u0_u2_n1100, _AES_ENC_u0_u2_n1099, _AES_ENC_u0_u2_n1098, _AES_ENC_u0_u2_n1097, _AES_ENC_u0_u2_n1096, _AES_ENC_u0_u2_n1095, _AES_ENC_u0_u2_n1094, _AES_ENC_u0_u2_n1093, _AES_ENC_u0_u2_n1092, _AES_ENC_u0_u2_n1091, _AES_ENC_u0_u2_n1090, _AES_ENC_u0_u2_n1089, _AES_ENC_u0_u2_n1088, _AES_ENC_u0_u2_n1087, _AES_ENC_u0_u2_n1086, _AES_ENC_u0_u2_n1085, _AES_ENC_u0_u2_n1084, _AES_ENC_u0_u2_n1083, _AES_ENC_u0_u2_n1082, _AES_ENC_u0_u2_n1081, _AES_ENC_u0_u2_n1080, _AES_ENC_u0_u2_n1079, _AES_ENC_u0_u2_n1078, _AES_ENC_u0_u2_n1077, _AES_ENC_u0_u2_n1076, 
  _AES_ENC_u0_u2_n1075, _AES_ENC_u0_u2_n1074, _AES_ENC_u0_u2_n1073, _AES_ENC_u0_u2_n1072, _AES_ENC_u0_u2_n1071, _AES_ENC_u0_u2_n1070, _AES_ENC_u0_u2_n1069, _AES_ENC_u0_u2_n1068, _AES_ENC_u0_u2_n1067, _AES_ENC_u0_u2_n1066, _AES_ENC_u0_u2_n1065, _AES_ENC_u0_u2_n1064, _AES_ENC_u0_u2_n1063, _AES_ENC_u0_u2_n1062, _AES_ENC_u0_u2_n1061, _AES_ENC_u0_u2_n1060, _AES_ENC_u0_u2_n1059, _AES_ENC_u0_u2_n1058, _AES_ENC_u0_u2_n1057, _AES_ENC_u0_u2_n1056, _AES_ENC_u0_u2_n1055, _AES_ENC_u0_u2_n1054, _AES_ENC_u0_u2_n1053, _AES_ENC_u0_u2_n1052, _AES_ENC_u0_u2_n1051, _AES_ENC_u0_u2_n1050, _AES_ENC_u0_u2_n1049, _AES_ENC_u0_u2_n1048, _AES_ENC_u0_u2_n1047, _AES_ENC_u0_u2_n1046, _AES_ENC_u0_u2_n1045, _AES_ENC_u0_u2_n1044, _AES_ENC_u0_u2_n1043, _AES_ENC_u0_u2_n1042, _AES_ENC_u0_u2_n1041, _AES_ENC_u0_u2_n1040, _AES_ENC_u0_u2_n1039, _AES_ENC_u0_u2_n1038, _AES_ENC_u0_u2_n1037, _AES_ENC_u0_u2_n1036, _AES_ENC_u0_u2_n1035, _AES_ENC_u0_u2_n1034, _AES_ENC_u0_u2_n1033, _AES_ENC_u0_u2_n1032, _AES_ENC_u0_u2_n1031, _AES_ENC_u0_u2_n1030, _AES_ENC_u0_u2_n1029, _AES_ENC_u0_u2_n1028, _AES_ENC_u0_u2_n1027, _AES_ENC_u0_u2_n1026, 
  _AES_ENC_u0_u2_n1025, _AES_ENC_u0_u2_n1024, _AES_ENC_u0_u2_n1023, _AES_ENC_u0_u2_n1022, _AES_ENC_u0_u2_n1021, _AES_ENC_u0_u2_n1020, _AES_ENC_u0_u2_n1019, _AES_ENC_u0_u2_n1018, _AES_ENC_u0_u2_n1017, _AES_ENC_u0_u2_n1016, _AES_ENC_u0_u2_n1015, _AES_ENC_u0_u2_n1014, _AES_ENC_u0_u2_n1013, _AES_ENC_u0_u2_n1012, _AES_ENC_u0_u2_n1011, _AES_ENC_u0_u2_n1010, _AES_ENC_u0_u2_n1009, _AES_ENC_u0_u2_n1008, _AES_ENC_u0_u2_n1007, _AES_ENC_u0_u2_n1006, _AES_ENC_u0_u2_n1005, _AES_ENC_u0_u2_n1004, _AES_ENC_u0_u2_n1003, _AES_ENC_u0_u2_n1002, _AES_ENC_u0_u2_n1001, _AES_ENC_u0_u2_n1000, _AES_ENC_u0_u2_n999, _AES_ENC_u0_u2_n998, _AES_ENC_u0_u2_n997, _AES_ENC_u0_u2_n996, _AES_ENC_u0_u2_n995, _AES_ENC_u0_u2_n994, _AES_ENC_u0_u2_n993, _AES_ENC_u0_u2_n992, _AES_ENC_u0_u2_n991, _AES_ENC_u0_u2_n990, _AES_ENC_u0_u2_n989, _AES_ENC_u0_u2_n988, _AES_ENC_u0_u2_n987, _AES_ENC_u0_u2_n986, _AES_ENC_u0_u2_n985, _AES_ENC_u0_u2_n984, _AES_ENC_u0_u2_n983, _AES_ENC_u0_u2_n982, _AES_ENC_u0_u2_n981, _AES_ENC_u0_u2_n980, _AES_ENC_u0_u2_n979, _AES_ENC_u0_u2_n978, _AES_ENC_u0_u2_n977, _AES_ENC_u0_u2_n976, 
  _AES_ENC_u0_u2_n975, _AES_ENC_u0_u2_n974, _AES_ENC_u0_u2_n973, _AES_ENC_u0_u2_n972, _AES_ENC_u0_u2_n971, _AES_ENC_u0_u2_n970, _AES_ENC_u0_u2_n969, _AES_ENC_u0_u2_n968, _AES_ENC_u0_u2_n967, _AES_ENC_u0_u2_n966, _AES_ENC_u0_u2_n965, _AES_ENC_u0_u2_n964, _AES_ENC_u0_u2_n963, _AES_ENC_u0_u2_n962, _AES_ENC_u0_u2_n961, _AES_ENC_u0_u2_n960, _AES_ENC_u0_u2_n959, _AES_ENC_u0_u2_n958, _AES_ENC_u0_u2_n957, _AES_ENC_u0_u2_n956, _AES_ENC_u0_u2_n955, _AES_ENC_u0_u2_n954, _AES_ENC_u0_u2_n953, _AES_ENC_u0_u2_n952, _AES_ENC_u0_u2_n951, _AES_ENC_u0_u2_n950, _AES_ENC_u0_u2_n949, _AES_ENC_u0_u2_n948, _AES_ENC_u0_u2_n947, _AES_ENC_u0_u2_n946, _AES_ENC_u0_u2_n945, _AES_ENC_u0_u2_n944, _AES_ENC_u0_u2_n943, _AES_ENC_u0_u2_n942, _AES_ENC_u0_u2_n941, _AES_ENC_u0_u2_n940, _AES_ENC_u0_u2_n939, _AES_ENC_u0_u2_n938, _AES_ENC_u0_u2_n937, _AES_ENC_u0_u2_n936, _AES_ENC_u0_u2_n935, _AES_ENC_u0_u2_n934, _AES_ENC_u0_u2_n933, _AES_ENC_u0_u2_n932, _AES_ENC_u0_u2_n931, _AES_ENC_u0_u2_n930, _AES_ENC_u0_u2_n929, _AES_ENC_u0_u2_n928, _AES_ENC_u0_u2_n927, _AES_ENC_u0_u2_n926, 
  _AES_ENC_u0_u2_n925, _AES_ENC_u0_u2_n924, _AES_ENC_u0_u2_n923, _AES_ENC_u0_u2_n922, _AES_ENC_u0_u2_n921, _AES_ENC_u0_u2_n920, _AES_ENC_u0_u2_n919, _AES_ENC_u0_u2_n918, _AES_ENC_u0_u2_n917, _AES_ENC_u0_u2_n916, _AES_ENC_u0_u2_n915, _AES_ENC_u0_u2_n914, _AES_ENC_u0_u2_n913, _AES_ENC_u0_u2_n912, _AES_ENC_u0_u2_n911, _AES_ENC_u0_u2_n910, _AES_ENC_u0_u2_n909, _AES_ENC_u0_u2_n908, _AES_ENC_u0_u2_n907, _AES_ENC_u0_u2_n906, _AES_ENC_u0_u2_n905, _AES_ENC_u0_u2_n904, _AES_ENC_u0_u2_n903, _AES_ENC_u0_u2_n902, _AES_ENC_u0_u2_n901, _AES_ENC_u0_u2_n900, _AES_ENC_u0_u2_n899, _AES_ENC_u0_u2_n898, _AES_ENC_u0_u2_n897, _AES_ENC_u0_u2_n896, _AES_ENC_u0_u2_n895, _AES_ENC_u0_u2_n894, _AES_ENC_u0_u2_n893, _AES_ENC_u0_u2_n892, _AES_ENC_u0_u2_n891, _AES_ENC_u0_u2_n890, _AES_ENC_u0_u2_n889, _AES_ENC_u0_u2_n888, _AES_ENC_u0_u2_n887, _AES_ENC_u0_u2_n886, _AES_ENC_u0_u2_n885, _AES_ENC_u0_u2_n884, _AES_ENC_u0_u2_n883, _AES_ENC_u0_u2_n882, _AES_ENC_u0_u2_n881, _AES_ENC_u0_u2_n880, _AES_ENC_u0_u2_n879, _AES_ENC_u0_u2_n878, _AES_ENC_u0_u2_n877, _AES_ENC_u0_u2_n876, 
  _AES_ENC_u0_u2_n875, _AES_ENC_u0_u2_n874, _AES_ENC_u0_u2_n873, _AES_ENC_u0_u2_n872, _AES_ENC_u0_u2_n871, _AES_ENC_u0_u2_n870, _AES_ENC_u0_u2_n869, _AES_ENC_u0_u2_n868, _AES_ENC_u0_u2_n867, _AES_ENC_u0_u2_n866, _AES_ENC_u0_u2_n865, _AES_ENC_u0_u2_n864, _AES_ENC_u0_u2_n863, _AES_ENC_u0_u2_n862, _AES_ENC_u0_u2_n861, _AES_ENC_u0_u2_n860, _AES_ENC_u0_u2_n859, _AES_ENC_u0_u2_n858, _AES_ENC_u0_u2_n857, _AES_ENC_u0_u2_n856, _AES_ENC_u0_u2_n855, _AES_ENC_u0_u2_n854, _AES_ENC_u0_u2_n853, _AES_ENC_u0_u2_n852, _AES_ENC_u0_u2_n851, _AES_ENC_u0_u2_n850, _AES_ENC_u0_u2_n849, _AES_ENC_u0_u2_n848, _AES_ENC_u0_u2_n847, _AES_ENC_u0_u2_n846, _AES_ENC_u0_u2_n845, _AES_ENC_u0_u2_n844, _AES_ENC_u0_u2_n843, _AES_ENC_u0_u2_n842, _AES_ENC_u0_u2_n841, _AES_ENC_u0_u2_n840, _AES_ENC_u0_u2_n839, _AES_ENC_u0_u2_n838, _AES_ENC_u0_u2_n837, _AES_ENC_u0_u2_n836, _AES_ENC_u0_u2_n835, _AES_ENC_u0_u2_n834, _AES_ENC_u0_u2_n833, _AES_ENC_u0_u2_n832, _AES_ENC_u0_u2_n831, _AES_ENC_u0_u2_n830, _AES_ENC_u0_u2_n829, _AES_ENC_u0_u2_n828, _AES_ENC_u0_u2_n827, _AES_ENC_u0_u2_n826, 
  _AES_ENC_u0_u2_n825, _AES_ENC_u0_u2_n824, _AES_ENC_u0_u2_n823, _AES_ENC_u0_u2_n822, _AES_ENC_u0_u2_n821, _AES_ENC_u0_u2_n820, _AES_ENC_u0_u2_n819, _AES_ENC_u0_u2_n818, _AES_ENC_u0_u2_n817, _AES_ENC_u0_u2_n816, _AES_ENC_u0_u2_n815, _AES_ENC_u0_u2_n814, _AES_ENC_u0_u2_n813, _AES_ENC_u0_u2_n812, _AES_ENC_u0_u2_n811, _AES_ENC_u0_u2_n810, _AES_ENC_u0_u2_n809, _AES_ENC_u0_u2_n808, _AES_ENC_u0_u2_n807, _AES_ENC_u0_u2_n806, _AES_ENC_u0_u2_n805, _AES_ENC_u0_u2_n804, _AES_ENC_u0_u2_n803, _AES_ENC_u0_u2_n802, _AES_ENC_u0_u2_n801, _AES_ENC_u0_u2_n800, _AES_ENC_u0_u2_n799, _AES_ENC_u0_u2_n798, _AES_ENC_u0_u2_n797, _AES_ENC_u0_u2_n796, _AES_ENC_u0_u2_n795, _AES_ENC_u0_u2_n794, _AES_ENC_u0_u2_n793, _AES_ENC_u0_u2_n792, _AES_ENC_u0_u2_n791, _AES_ENC_u0_u2_n790, _AES_ENC_u0_u2_n789, _AES_ENC_u0_u2_n788, _AES_ENC_u0_u2_n787, _AES_ENC_u0_u2_n786, _AES_ENC_u0_u2_n785, _AES_ENC_u0_u2_n784, _AES_ENC_u0_u2_n783, _AES_ENC_u0_u2_n782, _AES_ENC_u0_u2_n781, _AES_ENC_u0_u2_n780, _AES_ENC_u0_u2_n779, _AES_ENC_u0_u2_n778, _AES_ENC_u0_u2_n777, _AES_ENC_u0_u2_n776, 
  _AES_ENC_u0_u2_n775, _AES_ENC_u0_u2_n774, _AES_ENC_u0_u2_n773, _AES_ENC_u0_u2_n772, _AES_ENC_u0_u2_n771, _AES_ENC_u0_u2_n770, _AES_ENC_u0_u2_n769, _AES_ENC_u0_u2_n768, _AES_ENC_u0_u2_n767, _AES_ENC_u0_u2_n766, _AES_ENC_u0_u2_n765, _AES_ENC_u0_u2_n764, _AES_ENC_u0_u2_n763, _AES_ENC_u0_u2_n762, _AES_ENC_u0_u2_n761, _AES_ENC_u0_u2_n760, _AES_ENC_u0_u2_n759, _AES_ENC_u0_u2_n758, _AES_ENC_u0_u2_n757, _AES_ENC_u0_u2_n756, _AES_ENC_u0_u2_n755, _AES_ENC_u0_u2_n754, _AES_ENC_u0_u2_n753, _AES_ENC_u0_u2_n752, _AES_ENC_u0_u2_n751, _AES_ENC_u0_u2_n750, _AES_ENC_u0_u2_n749, _AES_ENC_u0_u2_n748, _AES_ENC_u0_u2_n747, _AES_ENC_u0_u2_n746, _AES_ENC_u0_u2_n745, _AES_ENC_u0_u2_n744, _AES_ENC_u0_u2_n743, _AES_ENC_u0_u2_n742, _AES_ENC_u0_u2_n741, _AES_ENC_u0_u2_n740, _AES_ENC_u0_u2_n739, _AES_ENC_u0_u2_n738, _AES_ENC_u0_u2_n737, _AES_ENC_u0_u2_n736, _AES_ENC_u0_u2_n735, _AES_ENC_u0_u2_n734, _AES_ENC_u0_u2_n733, _AES_ENC_u0_u2_n732, _AES_ENC_u0_u2_n731, _AES_ENC_u0_u2_n730, _AES_ENC_u0_u2_n729, _AES_ENC_u0_u2_n728, _AES_ENC_u0_u2_n727, _AES_ENC_u0_u2_n726, 
  _AES_ENC_u0_u2_n725, _AES_ENC_u0_u2_n724, _AES_ENC_u0_u2_n723, _AES_ENC_u0_u2_n722, _AES_ENC_u0_u2_n721, _AES_ENC_u0_u2_n720, _AES_ENC_u0_u2_n719, _AES_ENC_u0_u2_n718, _AES_ENC_u0_u2_n717, _AES_ENC_u0_u2_n716, _AES_ENC_u0_u2_n715, _AES_ENC_u0_u2_n714, _AES_ENC_u0_u2_n713, _AES_ENC_u0_u2_n712, _AES_ENC_u0_u2_n711, _AES_ENC_u0_u2_n710, _AES_ENC_u0_u2_n709, _AES_ENC_u0_u2_n708, _AES_ENC_u0_u2_n707, _AES_ENC_u0_u2_n706, _AES_ENC_u0_u2_n705, _AES_ENC_u0_u2_n704, _AES_ENC_u0_u2_n703, _AES_ENC_u0_u2_n702, _AES_ENC_u0_u2_n701, _AES_ENC_u0_u2_n700, _AES_ENC_u0_u2_n699, _AES_ENC_u0_u2_n698, _AES_ENC_u0_u2_n697, _AES_ENC_u0_u2_n696, _AES_ENC_u0_u2_n695, _AES_ENC_u0_u2_n694, _AES_ENC_u0_u2_n693, _AES_ENC_u0_u2_n692, _AES_ENC_u0_u2_n691, _AES_ENC_u0_u2_n690, _AES_ENC_u0_u2_n689, _AES_ENC_u0_u2_n688, _AES_ENC_u0_u2_n687, _AES_ENC_u0_u2_n686, _AES_ENC_u0_u2_n685, _AES_ENC_u0_u2_n684, _AES_ENC_u0_u2_n683, _AES_ENC_u0_u2_n682, _AES_ENC_u0_u2_n681, _AES_ENC_u0_u2_n680, _AES_ENC_u0_u2_n679, _AES_ENC_u0_u2_n678, _AES_ENC_u0_u2_n677, _AES_ENC_u0_u2_n676, 
  _AES_ENC_u0_u2_n675, _AES_ENC_u0_u2_n674, _AES_ENC_u0_u2_n673, _AES_ENC_u0_u2_n672, _AES_ENC_u0_u2_n671, _AES_ENC_u0_u2_n670, _AES_ENC_u0_u2_n669, _AES_ENC_u0_u2_n668, _AES_ENC_u0_u2_n667, _AES_ENC_u0_u2_n666, _AES_ENC_u0_u2_n665, _AES_ENC_u0_u2_n664, _AES_ENC_u0_u2_n663, _AES_ENC_u0_u2_n662, _AES_ENC_u0_u2_n661, _AES_ENC_u0_u2_n660, _AES_ENC_u0_u2_n659, _AES_ENC_u0_u2_n658, _AES_ENC_u0_u2_n657, _AES_ENC_u0_u2_n656, _AES_ENC_u0_u2_n655, _AES_ENC_u0_u2_n654, _AES_ENC_u0_u2_n653, _AES_ENC_u0_u2_n652, _AES_ENC_u0_u2_n651, _AES_ENC_u0_u2_n650, _AES_ENC_u0_u2_n649, _AES_ENC_u0_u2_n648, _AES_ENC_u0_u2_n647, _AES_ENC_u0_u2_n646, _AES_ENC_u0_u2_n645, _AES_ENC_u0_u2_n644, _AES_ENC_u0_u2_n643, _AES_ENC_u0_u2_n642, _AES_ENC_u0_u2_n641, _AES_ENC_u0_u2_n640, _AES_ENC_u0_u2_n639, _AES_ENC_u0_u2_n638, _AES_ENC_u0_u2_n637, _AES_ENC_u0_u2_n636, _AES_ENC_u0_u2_n635, _AES_ENC_u0_u2_n634, _AES_ENC_u0_u2_n633, _AES_ENC_u0_u2_n632, _AES_ENC_u0_u2_n631, _AES_ENC_u0_u2_n630, _AES_ENC_u0_u2_n629, _AES_ENC_u0_u2_n628, _AES_ENC_u0_u2_n627, _AES_ENC_u0_u2_n626, 
  _AES_ENC_u0_u2_n625, _AES_ENC_u0_u2_n624, _AES_ENC_u0_u2_n623, _AES_ENC_u0_u2_n622, _AES_ENC_u0_u2_n621, _AES_ENC_u0_u2_n620, _AES_ENC_u0_u2_n619, _AES_ENC_u0_u2_n618, _AES_ENC_u0_u2_n617, _AES_ENC_u0_u2_n616, _AES_ENC_u0_u2_n615, _AES_ENC_u0_u2_n614, _AES_ENC_u0_u2_n613, _AES_ENC_u0_u2_n612, _AES_ENC_u0_u2_n611, _AES_ENC_u0_u2_n610, _AES_ENC_u0_u2_n609, _AES_ENC_u0_u2_n608, _AES_ENC_u0_u2_n607, _AES_ENC_u0_u2_n606, _AES_ENC_u0_u2_n605, _AES_ENC_u0_u2_n604, _AES_ENC_u0_u2_n603, _AES_ENC_u0_u2_n602, _AES_ENC_u0_u2_n601, _AES_ENC_u0_u2_n600, _AES_ENC_u0_u2_n599, _AES_ENC_u0_u2_n598, _AES_ENC_u0_u2_n597, _AES_ENC_u0_u2_n596, _AES_ENC_u0_u2_n595, _AES_ENC_u0_u2_n594, _AES_ENC_u0_u2_n593, _AES_ENC_u0_u2_n592, _AES_ENC_u0_u2_n591, _AES_ENC_u0_u2_n590, _AES_ENC_u0_u2_n589, _AES_ENC_u0_u2_n588, _AES_ENC_u0_u2_n587, _AES_ENC_u0_u2_n586, _AES_ENC_u0_u2_n585, _AES_ENC_u0_u2_n584, _AES_ENC_u0_u2_n583, _AES_ENC_u0_u2_n582, _AES_ENC_u0_u2_n581, _AES_ENC_u0_u2_n580, _AES_ENC_u0_u2_n579, _AES_ENC_u0_u2_n578, _AES_ENC_u0_u2_n577, _AES_ENC_u0_u2_n576, 
  _AES_ENC_u0_u2_n575, _AES_ENC_u0_u2_n574, _AES_ENC_u0_u2_n573, _AES_ENC_u0_u2_n572, _AES_ENC_u0_u2_n571, _AES_ENC_u0_u2_n570, _AES_ENC_u0_u2_n569, _AES_ENC_u0_u3_n1135, _AES_ENC_u0_u3_n1134, _AES_ENC_u0_u3_n1133, _AES_ENC_u0_u3_n1132, _AES_ENC_u0_u3_n1131, _AES_ENC_u0_u3_n1130, _AES_ENC_u0_u3_n1129, _AES_ENC_u0_u3_n1128, _AES_ENC_u0_u3_n1127, _AES_ENC_u0_u3_n1126, _AES_ENC_u0_u3_n1125, _AES_ENC_u0_u3_n1124, _AES_ENC_u0_u3_n1123, _AES_ENC_u0_u3_n1122, _AES_ENC_u0_u3_n1121, _AES_ENC_u0_u3_n1120, _AES_ENC_u0_u3_n1119, _AES_ENC_u0_u3_n1118, _AES_ENC_u0_u3_n1117, _AES_ENC_u0_u3_n1116, _AES_ENC_u0_u3_n1115, _AES_ENC_u0_u3_n1114, _AES_ENC_u0_u3_n1113, _AES_ENC_u0_u3_n1112, _AES_ENC_u0_u3_n1111, _AES_ENC_u0_u3_n1110, _AES_ENC_u0_u3_n1109, _AES_ENC_u0_u3_n1108, _AES_ENC_u0_u3_n1107, _AES_ENC_u0_u3_n1106, _AES_ENC_u0_u3_n1105, _AES_ENC_u0_u3_n1104, _AES_ENC_u0_u3_n1103, _AES_ENC_u0_u3_n1102, _AES_ENC_u0_u3_n1101, _AES_ENC_u0_u3_n1100, _AES_ENC_u0_u3_n1099, _AES_ENC_u0_u3_n1098, _AES_ENC_u0_u3_n1097, _AES_ENC_u0_u3_n1096, _AES_ENC_u0_u3_n1095, _AES_ENC_u0_u3_n1094, _AES_ENC_u0_u3_n1093, 
  _AES_ENC_u0_u3_n1092, _AES_ENC_u0_u3_n1091, _AES_ENC_u0_u3_n1090, _AES_ENC_u0_u3_n1089, _AES_ENC_u0_u3_n1088, _AES_ENC_u0_u3_n1087, _AES_ENC_u0_u3_n1086, _AES_ENC_u0_u3_n1085, _AES_ENC_u0_u3_n1084, _AES_ENC_u0_u3_n1083, _AES_ENC_u0_u3_n1082, _AES_ENC_u0_u3_n1081, _AES_ENC_u0_u3_n1080, _AES_ENC_u0_u3_n1079, _AES_ENC_u0_u3_n1078, _AES_ENC_u0_u3_n1077, _AES_ENC_u0_u3_n1076, _AES_ENC_u0_u3_n1075, _AES_ENC_u0_u3_n1074, _AES_ENC_u0_u3_n1073, _AES_ENC_u0_u3_n1072, _AES_ENC_u0_u3_n1071, _AES_ENC_u0_u3_n1070, _AES_ENC_u0_u3_n1069, _AES_ENC_u0_u3_n1068, _AES_ENC_u0_u3_n1067, _AES_ENC_u0_u3_n1066, _AES_ENC_u0_u3_n1065, _AES_ENC_u0_u3_n1064, _AES_ENC_u0_u3_n1063, _AES_ENC_u0_u3_n1062, _AES_ENC_u0_u3_n1061, _AES_ENC_u0_u3_n1060, _AES_ENC_u0_u3_n1059, _AES_ENC_u0_u3_n1058, _AES_ENC_u0_u3_n1057, _AES_ENC_u0_u3_n1056, _AES_ENC_u0_u3_n1055, _AES_ENC_u0_u3_n1054, _AES_ENC_u0_u3_n1053, _AES_ENC_u0_u3_n1052, _AES_ENC_u0_u3_n1051, _AES_ENC_u0_u3_n1050, _AES_ENC_u0_u3_n1049, _AES_ENC_u0_u3_n1048, _AES_ENC_u0_u3_n1047, _AES_ENC_u0_u3_n1046, _AES_ENC_u0_u3_n1045, _AES_ENC_u0_u3_n1044, _AES_ENC_u0_u3_n1043, 
  _AES_ENC_u0_u3_n1042, _AES_ENC_u0_u3_n1041, _AES_ENC_u0_u3_n1040, _AES_ENC_u0_u3_n1039, _AES_ENC_u0_u3_n1038, _AES_ENC_u0_u3_n1037, _AES_ENC_u0_u3_n1036, _AES_ENC_u0_u3_n1035, _AES_ENC_u0_u3_n1034, _AES_ENC_u0_u3_n1033, _AES_ENC_u0_u3_n1032, _AES_ENC_u0_u3_n1031, _AES_ENC_u0_u3_n1030, _AES_ENC_u0_u3_n1029, _AES_ENC_u0_u3_n1028, _AES_ENC_u0_u3_n1027, _AES_ENC_u0_u3_n1026, _AES_ENC_u0_u3_n1025, _AES_ENC_u0_u3_n1024, _AES_ENC_u0_u3_n1023, _AES_ENC_u0_u3_n1022, _AES_ENC_u0_u3_n1021, _AES_ENC_u0_u3_n1020, _AES_ENC_u0_u3_n1019, _AES_ENC_u0_u3_n1018, _AES_ENC_u0_u3_n1017, _AES_ENC_u0_u3_n1016, _AES_ENC_u0_u3_n1015, _AES_ENC_u0_u3_n1014, _AES_ENC_u0_u3_n1013, _AES_ENC_u0_u3_n1012, _AES_ENC_u0_u3_n1011, _AES_ENC_u0_u3_n1010, _AES_ENC_u0_u3_n1009, _AES_ENC_u0_u3_n1008, _AES_ENC_u0_u3_n1007, _AES_ENC_u0_u3_n1006, _AES_ENC_u0_u3_n1005, _AES_ENC_u0_u3_n1004, _AES_ENC_u0_u3_n1003, _AES_ENC_u0_u3_n1002, _AES_ENC_u0_u3_n1001, _AES_ENC_u0_u3_n1000, _AES_ENC_u0_u3_n999, _AES_ENC_u0_u3_n998, _AES_ENC_u0_u3_n997, _AES_ENC_u0_u3_n996, _AES_ENC_u0_u3_n995, _AES_ENC_u0_u3_n994, _AES_ENC_u0_u3_n993, 
  _AES_ENC_u0_u3_n992, _AES_ENC_u0_u3_n991, _AES_ENC_u0_u3_n990, _AES_ENC_u0_u3_n989, _AES_ENC_u0_u3_n988, _AES_ENC_u0_u3_n987, _AES_ENC_u0_u3_n986, _AES_ENC_u0_u3_n985, _AES_ENC_u0_u3_n984, _AES_ENC_u0_u3_n983, _AES_ENC_u0_u3_n982, _AES_ENC_u0_u3_n981, _AES_ENC_u0_u3_n980, _AES_ENC_u0_u3_n979, _AES_ENC_u0_u3_n978, _AES_ENC_u0_u3_n977, _AES_ENC_u0_u3_n976, _AES_ENC_u0_u3_n975, _AES_ENC_u0_u3_n974, _AES_ENC_u0_u3_n973, _AES_ENC_u0_u3_n972, _AES_ENC_u0_u3_n971, _AES_ENC_u0_u3_n970, _AES_ENC_u0_u3_n969, _AES_ENC_u0_u3_n968, _AES_ENC_u0_u3_n967, _AES_ENC_u0_u3_n966, _AES_ENC_u0_u3_n965, _AES_ENC_u0_u3_n964, _AES_ENC_u0_u3_n963, _AES_ENC_u0_u3_n962, _AES_ENC_u0_u3_n961, _AES_ENC_u0_u3_n960, _AES_ENC_u0_u3_n959, _AES_ENC_u0_u3_n958, _AES_ENC_u0_u3_n957, _AES_ENC_u0_u3_n956, _AES_ENC_u0_u3_n955, _AES_ENC_u0_u3_n954, _AES_ENC_u0_u3_n953, _AES_ENC_u0_u3_n952, _AES_ENC_u0_u3_n951, _AES_ENC_u0_u3_n950, _AES_ENC_u0_u3_n949, _AES_ENC_u0_u3_n948, _AES_ENC_u0_u3_n947, _AES_ENC_u0_u3_n946, _AES_ENC_u0_u3_n945, _AES_ENC_u0_u3_n944, _AES_ENC_u0_u3_n943, 
  _AES_ENC_u0_u3_n942, _AES_ENC_u0_u3_n941, _AES_ENC_u0_u3_n940, _AES_ENC_u0_u3_n939, _AES_ENC_u0_u3_n938, _AES_ENC_u0_u3_n937, _AES_ENC_u0_u3_n936, _AES_ENC_u0_u3_n935, _AES_ENC_u0_u3_n934, _AES_ENC_u0_u3_n933, _AES_ENC_u0_u3_n932, _AES_ENC_u0_u3_n931, _AES_ENC_u0_u3_n930, _AES_ENC_u0_u3_n929, _AES_ENC_u0_u3_n928, _AES_ENC_u0_u3_n927, _AES_ENC_u0_u3_n926, _AES_ENC_u0_u3_n925, _AES_ENC_u0_u3_n924, _AES_ENC_u0_u3_n923, _AES_ENC_u0_u3_n922, _AES_ENC_u0_u3_n921, _AES_ENC_u0_u3_n920, _AES_ENC_u0_u3_n919, _AES_ENC_u0_u3_n918, _AES_ENC_u0_u3_n917, _AES_ENC_u0_u3_n916, _AES_ENC_u0_u3_n915, _AES_ENC_u0_u3_n914, _AES_ENC_u0_u3_n913, _AES_ENC_u0_u3_n912, _AES_ENC_u0_u3_n911, _AES_ENC_u0_u3_n910, _AES_ENC_u0_u3_n909, _AES_ENC_u0_u3_n908, _AES_ENC_u0_u3_n907, _AES_ENC_u0_u3_n906, _AES_ENC_u0_u3_n905, _AES_ENC_u0_u3_n904, _AES_ENC_u0_u3_n903, _AES_ENC_u0_u3_n902, _AES_ENC_u0_u3_n901, _AES_ENC_u0_u3_n900, _AES_ENC_u0_u3_n899, _AES_ENC_u0_u3_n898, _AES_ENC_u0_u3_n897, _AES_ENC_u0_u3_n896, _AES_ENC_u0_u3_n895, _AES_ENC_u0_u3_n894, _AES_ENC_u0_u3_n893, 
  _AES_ENC_u0_u3_n892, _AES_ENC_u0_u3_n891, _AES_ENC_u0_u3_n890, _AES_ENC_u0_u3_n889, _AES_ENC_u0_u3_n888, _AES_ENC_u0_u3_n887, _AES_ENC_u0_u3_n886, _AES_ENC_u0_u3_n885, _AES_ENC_u0_u3_n884, _AES_ENC_u0_u3_n883, _AES_ENC_u0_u3_n882, _AES_ENC_u0_u3_n881, _AES_ENC_u0_u3_n880, _AES_ENC_u0_u3_n879, _AES_ENC_u0_u3_n878, _AES_ENC_u0_u3_n877, _AES_ENC_u0_u3_n876, _AES_ENC_u0_u3_n875, _AES_ENC_u0_u3_n874, _AES_ENC_u0_u3_n873, _AES_ENC_u0_u3_n872, _AES_ENC_u0_u3_n871, _AES_ENC_u0_u3_n870, _AES_ENC_u0_u3_n869, _AES_ENC_u0_u3_n868, _AES_ENC_u0_u3_n867, _AES_ENC_u0_u3_n866, _AES_ENC_u0_u3_n865, _AES_ENC_u0_u3_n864, _AES_ENC_u0_u3_n863, _AES_ENC_u0_u3_n862, _AES_ENC_u0_u3_n861, _AES_ENC_u0_u3_n860, _AES_ENC_u0_u3_n859, _AES_ENC_u0_u3_n858, _AES_ENC_u0_u3_n857, _AES_ENC_u0_u3_n856, _AES_ENC_u0_u3_n855, _AES_ENC_u0_u3_n854, _AES_ENC_u0_u3_n853, _AES_ENC_u0_u3_n852, _AES_ENC_u0_u3_n851, _AES_ENC_u0_u3_n850, _AES_ENC_u0_u3_n849, _AES_ENC_u0_u3_n848, _AES_ENC_u0_u3_n847, _AES_ENC_u0_u3_n846, _AES_ENC_u0_u3_n845, _AES_ENC_u0_u3_n844, _AES_ENC_u0_u3_n843, 
  _AES_ENC_u0_u3_n842, _AES_ENC_u0_u3_n841, _AES_ENC_u0_u3_n840, _AES_ENC_u0_u3_n839, _AES_ENC_u0_u3_n838, _AES_ENC_u0_u3_n837, _AES_ENC_u0_u3_n836, _AES_ENC_u0_u3_n835, _AES_ENC_u0_u3_n834, _AES_ENC_u0_u3_n833, _AES_ENC_u0_u3_n832, _AES_ENC_u0_u3_n831, _AES_ENC_u0_u3_n830, _AES_ENC_u0_u3_n829, _AES_ENC_u0_u3_n828, _AES_ENC_u0_u3_n827, _AES_ENC_u0_u3_n826, _AES_ENC_u0_u3_n825, _AES_ENC_u0_u3_n824, _AES_ENC_u0_u3_n823, _AES_ENC_u0_u3_n822, _AES_ENC_u0_u3_n821, _AES_ENC_u0_u3_n820, _AES_ENC_u0_u3_n819, _AES_ENC_u0_u3_n818, _AES_ENC_u0_u3_n817, _AES_ENC_u0_u3_n816, _AES_ENC_u0_u3_n815, _AES_ENC_u0_u3_n814, _AES_ENC_u0_u3_n813, _AES_ENC_u0_u3_n812, _AES_ENC_u0_u3_n811, _AES_ENC_u0_u3_n810, _AES_ENC_u0_u3_n809, _AES_ENC_u0_u3_n808, _AES_ENC_u0_u3_n807, _AES_ENC_u0_u3_n806, _AES_ENC_u0_u3_n805, _AES_ENC_u0_u3_n804, _AES_ENC_u0_u3_n803, _AES_ENC_u0_u3_n802, _AES_ENC_u0_u3_n801, _AES_ENC_u0_u3_n800, _AES_ENC_u0_u3_n799, _AES_ENC_u0_u3_n798, _AES_ENC_u0_u3_n797, _AES_ENC_u0_u3_n796, _AES_ENC_u0_u3_n795, _AES_ENC_u0_u3_n794, _AES_ENC_u0_u3_n793, 
  _AES_ENC_u0_u3_n792, _AES_ENC_u0_u3_n791, _AES_ENC_u0_u3_n790, _AES_ENC_u0_u3_n789, _AES_ENC_u0_u3_n788, _AES_ENC_u0_u3_n787, _AES_ENC_u0_u3_n786, _AES_ENC_u0_u3_n785, _AES_ENC_u0_u3_n784, _AES_ENC_u0_u3_n783, _AES_ENC_u0_u3_n782, _AES_ENC_u0_u3_n781, _AES_ENC_u0_u3_n780, _AES_ENC_u0_u3_n779, _AES_ENC_u0_u3_n778, _AES_ENC_u0_u3_n777, _AES_ENC_u0_u3_n776, _AES_ENC_u0_u3_n775, _AES_ENC_u0_u3_n774, _AES_ENC_u0_u3_n773, _AES_ENC_u0_u3_n772, _AES_ENC_u0_u3_n771, _AES_ENC_u0_u3_n770, _AES_ENC_u0_u3_n769, _AES_ENC_u0_u3_n768, _AES_ENC_u0_u3_n767, _AES_ENC_u0_u3_n766, _AES_ENC_u0_u3_n765, _AES_ENC_u0_u3_n764, _AES_ENC_u0_u3_n763, _AES_ENC_u0_u3_n762, _AES_ENC_u0_u3_n761, _AES_ENC_u0_u3_n760, _AES_ENC_u0_u3_n759, _AES_ENC_u0_u3_n758, _AES_ENC_u0_u3_n757, _AES_ENC_u0_u3_n756, _AES_ENC_u0_u3_n755, _AES_ENC_u0_u3_n754, _AES_ENC_u0_u3_n753, _AES_ENC_u0_u3_n752, _AES_ENC_u0_u3_n751, _AES_ENC_u0_u3_n750, _AES_ENC_u0_u3_n749, _AES_ENC_u0_u3_n748, _AES_ENC_u0_u3_n747, _AES_ENC_u0_u3_n746, _AES_ENC_u0_u3_n745, _AES_ENC_u0_u3_n744, _AES_ENC_u0_u3_n743, 
  _AES_ENC_u0_u3_n742, _AES_ENC_u0_u3_n741, _AES_ENC_u0_u3_n740, _AES_ENC_u0_u3_n739, _AES_ENC_u0_u3_n738, _AES_ENC_u0_u3_n737, _AES_ENC_u0_u3_n736, _AES_ENC_u0_u3_n735, _AES_ENC_u0_u3_n734, _AES_ENC_u0_u3_n733, _AES_ENC_u0_u3_n732, _AES_ENC_u0_u3_n731, _AES_ENC_u0_u3_n730, _AES_ENC_u0_u3_n729, _AES_ENC_u0_u3_n728, _AES_ENC_u0_u3_n727, _AES_ENC_u0_u3_n726, _AES_ENC_u0_u3_n725, _AES_ENC_u0_u3_n724, _AES_ENC_u0_u3_n723, _AES_ENC_u0_u3_n722, _AES_ENC_u0_u3_n721, _AES_ENC_u0_u3_n720, _AES_ENC_u0_u3_n719, _AES_ENC_u0_u3_n718, _AES_ENC_u0_u3_n717, _AES_ENC_u0_u3_n716, _AES_ENC_u0_u3_n715, _AES_ENC_u0_u3_n714, _AES_ENC_u0_u3_n713, _AES_ENC_u0_u3_n712, _AES_ENC_u0_u3_n711, _AES_ENC_u0_u3_n710, _AES_ENC_u0_u3_n709, _AES_ENC_u0_u3_n708, _AES_ENC_u0_u3_n707, _AES_ENC_u0_u3_n706, _AES_ENC_u0_u3_n705, _AES_ENC_u0_u3_n704, _AES_ENC_u0_u3_n703, _AES_ENC_u0_u3_n702, _AES_ENC_u0_u3_n701, _AES_ENC_u0_u3_n700, _AES_ENC_u0_u3_n699, _AES_ENC_u0_u3_n698, _AES_ENC_u0_u3_n697, _AES_ENC_u0_u3_n696, _AES_ENC_u0_u3_n695, _AES_ENC_u0_u3_n694, _AES_ENC_u0_u3_n693, 
  _AES_ENC_u0_u3_n692, _AES_ENC_u0_u3_n691, _AES_ENC_u0_u3_n690, _AES_ENC_u0_u3_n689, _AES_ENC_u0_u3_n688, _AES_ENC_u0_u3_n687, _AES_ENC_u0_u3_n686, _AES_ENC_u0_u3_n685, _AES_ENC_u0_u3_n684, _AES_ENC_u0_u3_n683, _AES_ENC_u0_u3_n682, _AES_ENC_u0_u3_n681, _AES_ENC_u0_u3_n680, _AES_ENC_u0_u3_n679, _AES_ENC_u0_u3_n678, _AES_ENC_u0_u3_n677, _AES_ENC_u0_u3_n676, _AES_ENC_u0_u3_n675, _AES_ENC_u0_u3_n674, _AES_ENC_u0_u3_n673, _AES_ENC_u0_u3_n672, _AES_ENC_u0_u3_n671, _AES_ENC_u0_u3_n670, _AES_ENC_u0_u3_n669, _AES_ENC_u0_u3_n668, _AES_ENC_u0_u3_n667, _AES_ENC_u0_u3_n666, _AES_ENC_u0_u3_n665, _AES_ENC_u0_u3_n664, _AES_ENC_u0_u3_n663, _AES_ENC_u0_u3_n662, _AES_ENC_u0_u3_n661, _AES_ENC_u0_u3_n660, _AES_ENC_u0_u3_n659, _AES_ENC_u0_u3_n658, _AES_ENC_u0_u3_n657, _AES_ENC_u0_u3_n656, _AES_ENC_u0_u3_n655, _AES_ENC_u0_u3_n654, _AES_ENC_u0_u3_n653, _AES_ENC_u0_u3_n652, _AES_ENC_u0_u3_n651, _AES_ENC_u0_u3_n650, _AES_ENC_u0_u3_n649, _AES_ENC_u0_u3_n648, _AES_ENC_u0_u3_n647, _AES_ENC_u0_u3_n646, _AES_ENC_u0_u3_n645, _AES_ENC_u0_u3_n644, _AES_ENC_u0_u3_n643, 
  _AES_ENC_u0_u3_n642, _AES_ENC_u0_u3_n641, _AES_ENC_u0_u3_n640, _AES_ENC_u0_u3_n639, _AES_ENC_u0_u3_n638, _AES_ENC_u0_u3_n637, _AES_ENC_u0_u3_n636, _AES_ENC_u0_u3_n635, _AES_ENC_u0_u3_n634, _AES_ENC_u0_u3_n633, _AES_ENC_u0_u3_n632, _AES_ENC_u0_u3_n631, _AES_ENC_u0_u3_n630, _AES_ENC_u0_u3_n629, _AES_ENC_u0_u3_n628, _AES_ENC_u0_u3_n627, _AES_ENC_u0_u3_n626, _AES_ENC_u0_u3_n625, _AES_ENC_u0_u3_n624, _AES_ENC_u0_u3_n623, _AES_ENC_u0_u3_n622, _AES_ENC_u0_u3_n621, _AES_ENC_u0_u3_n620, _AES_ENC_u0_u3_n619, _AES_ENC_u0_u3_n618, _AES_ENC_u0_u3_n617, _AES_ENC_u0_u3_n616, _AES_ENC_u0_u3_n615, _AES_ENC_u0_u3_n614, _AES_ENC_u0_u3_n613, _AES_ENC_u0_u3_n612, _AES_ENC_u0_u3_n611, _AES_ENC_u0_u3_n610, _AES_ENC_u0_u3_n609, _AES_ENC_u0_u3_n608, _AES_ENC_u0_u3_n607, _AES_ENC_u0_u3_n606, _AES_ENC_u0_u3_n605, _AES_ENC_u0_u3_n604, _AES_ENC_u0_u3_n603, _AES_ENC_u0_u3_n602, _AES_ENC_u0_u3_n601, _AES_ENC_u0_u3_n600, _AES_ENC_u0_u3_n599, _AES_ENC_u0_u3_n598, _AES_ENC_u0_u3_n597, _AES_ENC_u0_u3_n596, _AES_ENC_u0_u3_n595, _AES_ENC_u0_u3_n594, _AES_ENC_u0_u3_n593, 
  _AES_ENC_u0_u3_n592, _AES_ENC_u0_u3_n591, _AES_ENC_u0_u3_n590, _AES_ENC_u0_u3_n589, _AES_ENC_u0_u3_n588, _AES_ENC_u0_u3_n587, _AES_ENC_u0_u3_n586, _AES_ENC_u0_u3_n585, _AES_ENC_u0_u3_n584, _AES_ENC_u0_u3_n583, _AES_ENC_u0_u3_n582, _AES_ENC_u0_u3_n581, _AES_ENC_u0_u3_n580, _AES_ENC_u0_u3_n579, _AES_ENC_u0_u3_n578, _AES_ENC_u0_u3_n577, _AES_ENC_u0_u3_n576, _AES_ENC_u0_u3_n575, _AES_ENC_u0_u3_n574, _AES_ENC_u0_u3_n573, _AES_ENC_u0_u3_n572, _AES_ENC_u0_u3_n571, _AES_ENC_u0_u3_n570, _AES_ENC_u0_u3_n569, _AES_ENC_u0_r0_n38, _AES_ENC_u0_r0_n37, _AES_ENC_u0_r0_n36, _AES_ENC_u0_r0_n35, _AES_ENC_u0_r0_n34, _AES_ENC_u0_r0_n33, _AES_ENC_u0_r0_n29, _AES_ENC_u0_r0_n28, _AES_ENC_u0_r0_n27, _AES_ENC_u0_r0_n26, _AES_ENC_u0_r0_n25, _AES_ENC_u0_r0_n24, _AES_ENC_u0_r0_n23, _AES_ENC_u0_r0_n22, _AES_ENC_u0_r0_n21, _AES_ENC_u0_r0_n20, _AES_ENC_u0_r0_n19, _AES_ENC_u0_r0_n18, _AES_ENC_u0_r0_n17, _AES_ENC_u0_r0_n16, _AES_ENC_u0_r0_n15, _AES_ENC_u0_r0_n14, _AES_ENC_u0_r0_n13, _AES_ENC_u0_r0_n12, _AES_ENC_u0_r0_n11, _AES_ENC_u0_r0_n10, 
  _AES_ENC_u0_r0_n9, _AES_ENC_u0_r0_n8, _AES_ENC_u0_r0_n7, _AES_ENC_u0_r0_n32, _AES_ENC_u0_r0_N55, _AES_ENC_u0_r0_N54, _AES_ENC_u0_r0_N53, _AES_ENC_u0_r0_rcnt[0], _AES_ENC_u0_r0_rcnt[1], _AES_ENC_u0_r0_rcnt[2], _AES_ENC_u0_r0_N51, _AES_ENC_u0_r0_N50, _AES_ENC_u0_r0_N49, _AES_ENC_u0_r0_N48, _AES_ENC_u0_r0_N47, _AES_ENC_u0_r0_N46, _AES_ENC_u0_r0_N45, _AES_ENC_u0_r0_N44, _AES_ENC_us00_n627, _AES_ENC_us00_n626, _AES_ENC_us00_n625, _AES_ENC_us00_n624, _AES_ENC_us00_n623, _AES_ENC_us00_n622, _AES_ENC_us00_n621, _AES_ENC_us00_n620, _AES_ENC_us00_n619, _AES_ENC_us00_n618, _AES_ENC_us00_n617, _AES_ENC_us00_n616, _AES_ENC_us00_n615, _AES_ENC_us00_n614, _AES_ENC_us00_n613, _AES_ENC_us00_n612, _AES_ENC_us00_n611, _AES_ENC_us00_n610, _AES_ENC_us00_n609, _AES_ENC_us00_n608, _AES_ENC_us00_n607, _AES_ENC_us00_n606, _AES_ENC_us00_n605, _AES_ENC_us00_n604, _AES_ENC_us00_n603, _AES_ENC_us00_n602, _AES_ENC_us00_n601, _AES_ENC_us00_n600, _AES_ENC_us00_n599, _AES_ENC_us00_n598, _AES_ENC_us00_n597, _AES_ENC_us00_n596, 
  _AES_ENC_us00_n595, _AES_ENC_us00_n594, _AES_ENC_us00_n593, _AES_ENC_us00_n592, _AES_ENC_us00_n591, _AES_ENC_us00_n590, _AES_ENC_us00_n589, _AES_ENC_us00_n588, _AES_ENC_us00_n587, _AES_ENC_us00_n586, _AES_ENC_us00_n585, _AES_ENC_us00_n584, _AES_ENC_us00_n583, _AES_ENC_us00_n582, _AES_ENC_us00_n581, _AES_ENC_us00_n580, _AES_ENC_us00_n579, _AES_ENC_us00_n578, _AES_ENC_us00_n577, _AES_ENC_us00_n576, _AES_ENC_us00_n575, _AES_ENC_us00_n574, _AES_ENC_us00_n573, _AES_ENC_us00_n572, _AES_ENC_us00_n571, _AES_ENC_us00_n570, _AES_ENC_us00_n569, _AES_ENC_us00_n568, _AES_ENC_us00_n567, _AES_ENC_us00_n566, _AES_ENC_us00_n565, _AES_ENC_us00_n564, _AES_ENC_us00_n563, _AES_ENC_us00_n562, _AES_ENC_us00_n561, _AES_ENC_us00_n560, _AES_ENC_us00_n559, _AES_ENC_us00_n558, _AES_ENC_us00_n557, _AES_ENC_us00_n556, _AES_ENC_us00_n555, _AES_ENC_us00_n554, _AES_ENC_us00_n553, _AES_ENC_us00_n552, _AES_ENC_us00_n551, _AES_ENC_us00_n550, _AES_ENC_us00_n549, _AES_ENC_us00_n548, _AES_ENC_us00_n547, _AES_ENC_us00_n546, 
  _AES_ENC_us00_n545, _AES_ENC_us00_n544, _AES_ENC_us00_n543, _AES_ENC_us00_n542, _AES_ENC_us00_n541, _AES_ENC_us00_n540, _AES_ENC_us00_n539, _AES_ENC_us00_n538, _AES_ENC_us00_n537, _AES_ENC_us00_n536, _AES_ENC_us00_n535, _AES_ENC_us00_n534, _AES_ENC_us00_n533, _AES_ENC_us00_n532, _AES_ENC_us00_n531, _AES_ENC_us00_n530, _AES_ENC_us00_n529, _AES_ENC_us00_n528, _AES_ENC_us00_n527, _AES_ENC_us00_n526, _AES_ENC_us00_n525, _AES_ENC_us00_n524, _AES_ENC_us00_n523, _AES_ENC_us00_n522, _AES_ENC_us00_n521, _AES_ENC_us00_n520, _AES_ENC_us00_n519, _AES_ENC_us00_n518, _AES_ENC_us00_n517, _AES_ENC_us00_n516, _AES_ENC_us00_n515, _AES_ENC_us00_n514, _AES_ENC_us00_n513, _AES_ENC_us00_n512, _AES_ENC_us00_n511, _AES_ENC_us00_n510, _AES_ENC_us00_n509, _AES_ENC_us00_n508, _AES_ENC_us00_n507, _AES_ENC_us00_n506, _AES_ENC_us00_n505, _AES_ENC_us00_n504, _AES_ENC_us00_n503, _AES_ENC_us00_n502, _AES_ENC_us00_n501, _AES_ENC_us00_n500, _AES_ENC_us00_n499, _AES_ENC_us00_n498, _AES_ENC_us00_n497, _AES_ENC_us00_n496, 
  _AES_ENC_us00_n495, _AES_ENC_us00_n494, _AES_ENC_us00_n493, _AES_ENC_us00_n492, _AES_ENC_us00_n491, _AES_ENC_us00_n490, _AES_ENC_us00_n489, _AES_ENC_us00_n488, _AES_ENC_us00_n487, _AES_ENC_us00_n486, _AES_ENC_us00_n485, _AES_ENC_us00_n484, _AES_ENC_us00_n483, _AES_ENC_us00_n482, _AES_ENC_us00_n481, _AES_ENC_us00_n480, _AES_ENC_us00_n479, _AES_ENC_us00_n478, _AES_ENC_us00_n477, _AES_ENC_us00_n476, _AES_ENC_us00_n475, _AES_ENC_us00_n474, _AES_ENC_us00_n473, _AES_ENC_us00_n472, _AES_ENC_us00_n471, _AES_ENC_us00_n470, _AES_ENC_us00_n469, _AES_ENC_us00_n468, _AES_ENC_us00_n467, _AES_ENC_us00_n466, _AES_ENC_us00_n465, _AES_ENC_us00_n464, _AES_ENC_us00_n463, _AES_ENC_us00_n462, _AES_ENC_us00_n461, _AES_ENC_us00_n460, _AES_ENC_us00_n459, _AES_ENC_us00_n458, _AES_ENC_us00_n457, _AES_ENC_us00_n456, _AES_ENC_us00_n455, _AES_ENC_us00_n454, _AES_ENC_us00_n453, _AES_ENC_us00_n452, _AES_ENC_us00_n451, _AES_ENC_us00_n450, _AES_ENC_us00_n449, _AES_ENC_us00_n448, _AES_ENC_us00_n447, _AES_ENC_us00_n446, 
  _AES_ENC_us00_n445, _AES_ENC_us00_n444, _AES_ENC_us00_n443, _AES_ENC_us00_n442, _AES_ENC_us00_n441, _AES_ENC_us00_n440, _AES_ENC_us00_n439, _AES_ENC_us00_n438, _AES_ENC_us00_n437, _AES_ENC_us00_n436, _AES_ENC_us00_n435, _AES_ENC_us00_n434, _AES_ENC_us00_n433, _AES_ENC_us00_n432, _AES_ENC_us00_n431, _AES_ENC_us00_n430, _AES_ENC_us00_n429, _AES_ENC_us00_n428, _AES_ENC_us00_n427, _AES_ENC_us00_n426, _AES_ENC_us00_n425, _AES_ENC_us00_n424, _AES_ENC_us00_n423, _AES_ENC_us00_n422, _AES_ENC_us00_n421, _AES_ENC_us00_n420, _AES_ENC_us00_n419, _AES_ENC_us00_n418, _AES_ENC_us00_n417, _AES_ENC_us00_n416, _AES_ENC_us00_n415, _AES_ENC_us00_n414, _AES_ENC_us00_n413, _AES_ENC_us00_n412, _AES_ENC_us00_n411, _AES_ENC_us00_n410, _AES_ENC_us00_n409, _AES_ENC_us00_n408, _AES_ENC_us00_n407, _AES_ENC_us00_n406, _AES_ENC_us00_n405, _AES_ENC_us00_n404, _AES_ENC_us00_n403, _AES_ENC_us00_n402, _AES_ENC_us00_n401, _AES_ENC_us00_n400, _AES_ENC_us00_n399, _AES_ENC_us00_n398, _AES_ENC_us00_n397, _AES_ENC_us00_n396, 
  _AES_ENC_us00_n395, _AES_ENC_us00_n394, _AES_ENC_us00_n393, _AES_ENC_us00_n392, _AES_ENC_us00_n391, _AES_ENC_us00_n390, _AES_ENC_us00_n389, _AES_ENC_us00_n388, _AES_ENC_us00_n387, _AES_ENC_us00_n386, _AES_ENC_us00_n385, _AES_ENC_us00_n384, _AES_ENC_us00_n383, _AES_ENC_us00_n382, _AES_ENC_us00_n381, _AES_ENC_us00_n380, _AES_ENC_us00_n379, _AES_ENC_us00_n378, _AES_ENC_us00_n377, _AES_ENC_us00_n376, _AES_ENC_us00_n375, _AES_ENC_us00_n374, _AES_ENC_us00_n373, _AES_ENC_us00_n372, _AES_ENC_us00_n371, _AES_ENC_us00_n370, _AES_ENC_us00_n369, _AES_ENC_us00_n368, _AES_ENC_us00_n367, _AES_ENC_us00_n366, _AES_ENC_us00_n365, _AES_ENC_us00_n364, _AES_ENC_us00_n363, _AES_ENC_us00_n362, _AES_ENC_us00_n361, _AES_ENC_us00_n360, _AES_ENC_us00_n359, _AES_ENC_us00_n358, _AES_ENC_us00_n357, _AES_ENC_us00_n356, _AES_ENC_us00_n355, _AES_ENC_us00_n354, _AES_ENC_us00_n353, _AES_ENC_us00_n352, _AES_ENC_us00_n351, _AES_ENC_us00_n350, _AES_ENC_us00_n349, _AES_ENC_us00_n348, _AES_ENC_us00_n347, _AES_ENC_us00_n346, 
  _AES_ENC_us00_n345, _AES_ENC_us00_n344, _AES_ENC_us00_n343, _AES_ENC_us00_n342, _AES_ENC_us00_n341, _AES_ENC_us00_n340, _AES_ENC_us00_n339, _AES_ENC_us00_n338, _AES_ENC_us00_n337, _AES_ENC_us00_n336, _AES_ENC_us00_n335, _AES_ENC_us00_n334, _AES_ENC_us00_n333, _AES_ENC_us00_n332, _AES_ENC_us00_n331, _AES_ENC_us00_n330, _AES_ENC_us00_n329, _AES_ENC_us00_n328, _AES_ENC_us00_n327, _AES_ENC_us00_n326, _AES_ENC_us00_n325, _AES_ENC_us00_n324, _AES_ENC_us00_n323, _AES_ENC_us00_n322, _AES_ENC_us00_n321, _AES_ENC_us00_n320, _AES_ENC_us00_n319, _AES_ENC_us00_n318, _AES_ENC_us00_n317, _AES_ENC_us00_n316, _AES_ENC_us00_n315, _AES_ENC_us00_n314, _AES_ENC_us00_n313, _AES_ENC_us00_n312, _AES_ENC_us00_n311, _AES_ENC_us00_n310, _AES_ENC_us00_n309, _AES_ENC_us00_n308, _AES_ENC_us00_n307, _AES_ENC_us00_n306, _AES_ENC_us00_n305, _AES_ENC_us00_n304, _AES_ENC_us00_n303, _AES_ENC_us00_n302, _AES_ENC_us00_n301, _AES_ENC_us00_n300, _AES_ENC_us00_n299, _AES_ENC_us00_n298, _AES_ENC_us00_n297, _AES_ENC_us00_n296, 
  _AES_ENC_us00_n295, _AES_ENC_us00_n294, _AES_ENC_us00_n293, _AES_ENC_us00_n292, _AES_ENC_us00_n291, _AES_ENC_us00_n290, _AES_ENC_us00_n289, _AES_ENC_us00_n288, _AES_ENC_us00_n287, _AES_ENC_us00_n286, _AES_ENC_us00_n285, _AES_ENC_us00_n284, _AES_ENC_us00_n283, _AES_ENC_us00_n282, _AES_ENC_us00_n281, _AES_ENC_us00_n280, _AES_ENC_us00_n279, _AES_ENC_us00_n278, _AES_ENC_us00_n277, _AES_ENC_us00_n276, _AES_ENC_us00_n275, _AES_ENC_us00_n274, _AES_ENC_us00_n273, _AES_ENC_us00_n272, _AES_ENC_us00_n271, _AES_ENC_us00_n270, _AES_ENC_us00_n269, _AES_ENC_us00_n268, _AES_ENC_us00_n267, _AES_ENC_us00_n266, _AES_ENC_us00_n265, _AES_ENC_us00_n264, _AES_ENC_us00_n263, _AES_ENC_us00_n262, _AES_ENC_us00_n261, _AES_ENC_us00_n260, _AES_ENC_us00_n259, _AES_ENC_us00_n258, _AES_ENC_us00_n257, _AES_ENC_us00_n256, _AES_ENC_us00_n255, _AES_ENC_us00_n254, _AES_ENC_us00_n253, _AES_ENC_us00_n252, _AES_ENC_us00_n251, _AES_ENC_us00_n250, _AES_ENC_us00_n249, _AES_ENC_us00_n248, _AES_ENC_us00_n247, _AES_ENC_us00_n246, 
  _AES_ENC_us00_n245, _AES_ENC_us00_n244, _AES_ENC_us00_n243, _AES_ENC_us00_n242, _AES_ENC_us00_n241, _AES_ENC_us00_n240, _AES_ENC_us00_n239, _AES_ENC_us00_n238, _AES_ENC_us00_n237, _AES_ENC_us00_n235, _AES_ENC_us00_n234, _AES_ENC_us00_n233, _AES_ENC_us00_n232, _AES_ENC_us00_n231, _AES_ENC_us00_n230, _AES_ENC_us00_n229, _AES_ENC_us00_n228, _AES_ENC_us00_n227, _AES_ENC_us00_n226, _AES_ENC_us00_n225, _AES_ENC_us00_n224, _AES_ENC_us00_n223, _AES_ENC_us00_n222, _AES_ENC_us00_n221, _AES_ENC_us00_n220, _AES_ENC_us00_n219, _AES_ENC_us00_n218, _AES_ENC_us00_n217, _AES_ENC_us00_n216, _AES_ENC_us00_n215, _AES_ENC_us00_n214, _AES_ENC_us00_n213, _AES_ENC_us00_n212, _AES_ENC_us00_n211, _AES_ENC_us00_n210, _AES_ENC_us00_n209, _AES_ENC_us00_n208, _AES_ENC_us00_n207, _AES_ENC_us00_n206, _AES_ENC_us00_n205, _AES_ENC_us00_n204, _AES_ENC_us00_n203, _AES_ENC_us00_n202, _AES_ENC_us00_n201, _AES_ENC_us00_n200, _AES_ENC_us00_n199, _AES_ENC_us00_n198, _AES_ENC_us00_n197, _AES_ENC_us00_n196, _AES_ENC_us00_n195, 
  _AES_ENC_us00_n194, _AES_ENC_us00_n193, _AES_ENC_us00_n192, _AES_ENC_us00_n191, _AES_ENC_us00_n190, _AES_ENC_us00_n189, _AES_ENC_us00_n188, _AES_ENC_us00_n187, _AES_ENC_us00_n186, _AES_ENC_us00_n185, _AES_ENC_us00_n184, _AES_ENC_us00_n183, _AES_ENC_us00_n182, _AES_ENC_us00_n181, _AES_ENC_us00_n180, _AES_ENC_us00_n179, _AES_ENC_us00_n178, _AES_ENC_us00_n177, _AES_ENC_us00_n176, _AES_ENC_us00_n175, _AES_ENC_us00_n174, _AES_ENC_us00_n173, _AES_ENC_us00_n172, _AES_ENC_us00_n171, _AES_ENC_us00_n170, _AES_ENC_us00_n168, _AES_ENC_us00_n167, _AES_ENC_us00_n166, _AES_ENC_us00_n165, _AES_ENC_us00_n164, _AES_ENC_us00_n163, _AES_ENC_us00_n162, _AES_ENC_us00_n161, _AES_ENC_us00_n160, _AES_ENC_us00_n159, _AES_ENC_us00_n158, _AES_ENC_us00_n157, _AES_ENC_us00_n156, _AES_ENC_us00_n155, _AES_ENC_us00_n154, _AES_ENC_us00_n153, _AES_ENC_us00_n152, _AES_ENC_us00_n151, _AES_ENC_us00_n150, _AES_ENC_us00_n149, _AES_ENC_us00_n148, _AES_ENC_us00_n147, _AES_ENC_us00_n146, _AES_ENC_us00_n145, _AES_ENC_us00_n144, 
  _AES_ENC_us00_n143, _AES_ENC_us00_n142, _AES_ENC_us00_n141, _AES_ENC_us00_n140, _AES_ENC_us00_n139, _AES_ENC_us00_n138, _AES_ENC_us00_n137, _AES_ENC_us00_n136, _AES_ENC_us00_n135, _AES_ENC_us00_n134, _AES_ENC_us00_n133, _AES_ENC_us00_n132, _AES_ENC_us00_n131, _AES_ENC_us00_n130, _AES_ENC_us00_n129, _AES_ENC_us00_n128, _AES_ENC_us00_n127, _AES_ENC_us00_n126, _AES_ENC_us00_n125, _AES_ENC_us00_n124, _AES_ENC_us00_n123, _AES_ENC_us00_n122, _AES_ENC_us00_n121, _AES_ENC_us00_n120, _AES_ENC_us00_n119, _AES_ENC_us00_n118, _AES_ENC_us00_n117, _AES_ENC_us00_n116, _AES_ENC_us00_n115, _AES_ENC_us00_n114, _AES_ENC_us00_n113, _AES_ENC_us00_n112, _AES_ENC_us00_n111, _AES_ENC_us00_n110, _AES_ENC_us00_n109, _AES_ENC_us00_n108, _AES_ENC_us00_n107, _AES_ENC_us00_n106, _AES_ENC_us00_n105, _AES_ENC_us00_n104, _AES_ENC_us00_n103, _AES_ENC_us00_n102, _AES_ENC_us00_n101, _AES_ENC_us00_n100, _AES_ENC_us00_n99, _AES_ENC_us00_n97, _AES_ENC_us00_n96, _AES_ENC_us00_n95, _AES_ENC_us00_n94, _AES_ENC_us00_n93, 
  _AES_ENC_us00_n92, _AES_ENC_us00_n91, _AES_ENC_us00_n90, _AES_ENC_us00_n89, _AES_ENC_us00_n88, _AES_ENC_us00_n87, _AES_ENC_us00_n86, _AES_ENC_us00_n85, _AES_ENC_us00_n84, _AES_ENC_us00_n83, _AES_ENC_us00_n82, _AES_ENC_us00_n81, _AES_ENC_us00_n80, _AES_ENC_us00_n79, _AES_ENC_us00_n78, _AES_ENC_us00_n77, _AES_ENC_us00_n76, _AES_ENC_us00_n75, _AES_ENC_us00_n74, _AES_ENC_us00_n73, _AES_ENC_us00_n72, _AES_ENC_us00_n71, _AES_ENC_us00_n70, _AES_ENC_us00_n69, _AES_ENC_us00_n68, _AES_ENC_us00_n67, _AES_ENC_us00_n66, _AES_ENC_us00_n65, _AES_ENC_us00_n64, _AES_ENC_us00_n63, _AES_ENC_us00_n62, _AES_ENC_us00_n61, _AES_ENC_us00_n60, _AES_ENC_us00_n59, _AES_ENC_us00_n58, _AES_ENC_us01_n1135, _AES_ENC_us01_n1134, _AES_ENC_us01_n1133, _AES_ENC_us01_n1132, _AES_ENC_us01_n1131, _AES_ENC_us01_n1130, _AES_ENC_us01_n1129, _AES_ENC_us01_n1128, _AES_ENC_us01_n1127, _AES_ENC_us01_n1126, _AES_ENC_us01_n1125, _AES_ENC_us01_n1124, _AES_ENC_us01_n1123, _AES_ENC_us01_n1122, _AES_ENC_us01_n1121, 
  _AES_ENC_us01_n1120, _AES_ENC_us01_n1119, _AES_ENC_us01_n1118, _AES_ENC_us01_n1117, _AES_ENC_us01_n1116, _AES_ENC_us01_n1115, _AES_ENC_us01_n1114, _AES_ENC_us01_n1113, _AES_ENC_us01_n1112, _AES_ENC_us01_n1111, _AES_ENC_us01_n1110, _AES_ENC_us01_n1109, _AES_ENC_us01_n1108, _AES_ENC_us01_n1107, _AES_ENC_us01_n1106, _AES_ENC_us01_n1105, _AES_ENC_us01_n1104, _AES_ENC_us01_n1103, _AES_ENC_us01_n1102, _AES_ENC_us01_n1101, _AES_ENC_us01_n1100, _AES_ENC_us01_n1099, _AES_ENC_us01_n1098, _AES_ENC_us01_n1097, _AES_ENC_us01_n1096, _AES_ENC_us01_n1095, _AES_ENC_us01_n1094, _AES_ENC_us01_n1093, _AES_ENC_us01_n1092, _AES_ENC_us01_n1091, _AES_ENC_us01_n1090, _AES_ENC_us01_n1089, _AES_ENC_us01_n1088, _AES_ENC_us01_n1087, _AES_ENC_us01_n1086, _AES_ENC_us01_n1085, _AES_ENC_us01_n1084, _AES_ENC_us01_n1083, _AES_ENC_us01_n1082, _AES_ENC_us01_n1081, _AES_ENC_us01_n1080, _AES_ENC_us01_n1079, _AES_ENC_us01_n1078, _AES_ENC_us01_n1077, _AES_ENC_us01_n1076, _AES_ENC_us01_n1075, _AES_ENC_us01_n1074, _AES_ENC_us01_n1073, _AES_ENC_us01_n1072, _AES_ENC_us01_n1071, 
  _AES_ENC_us01_n1070, _AES_ENC_us01_n1069, _AES_ENC_us01_n1068, _AES_ENC_us01_n1067, _AES_ENC_us01_n1066, _AES_ENC_us01_n1065, _AES_ENC_us01_n1064, _AES_ENC_us01_n1063, _AES_ENC_us01_n1062, _AES_ENC_us01_n1061, _AES_ENC_us01_n1060, _AES_ENC_us01_n1059, _AES_ENC_us01_n1058, _AES_ENC_us01_n1057, _AES_ENC_us01_n1056, _AES_ENC_us01_n1055, _AES_ENC_us01_n1054, _AES_ENC_us01_n1053, _AES_ENC_us01_n1052, _AES_ENC_us01_n1051, _AES_ENC_us01_n1050, _AES_ENC_us01_n1049, _AES_ENC_us01_n1048, _AES_ENC_us01_n1047, _AES_ENC_us01_n1046, _AES_ENC_us01_n1045, _AES_ENC_us01_n1044, _AES_ENC_us01_n1043, _AES_ENC_us01_n1042, _AES_ENC_us01_n1041, _AES_ENC_us01_n1040, _AES_ENC_us01_n1039, _AES_ENC_us01_n1038, _AES_ENC_us01_n1037, _AES_ENC_us01_n1036, _AES_ENC_us01_n1035, _AES_ENC_us01_n1034, _AES_ENC_us01_n1033, _AES_ENC_us01_n1032, _AES_ENC_us01_n1031, _AES_ENC_us01_n1030, _AES_ENC_us01_n1029, _AES_ENC_us01_n1028, _AES_ENC_us01_n1027, _AES_ENC_us01_n1026, _AES_ENC_us01_n1025, _AES_ENC_us01_n1024, _AES_ENC_us01_n1023, _AES_ENC_us01_n1022, _AES_ENC_us01_n1021, 
  _AES_ENC_us01_n1020, _AES_ENC_us01_n1019, _AES_ENC_us01_n1018, _AES_ENC_us01_n1017, _AES_ENC_us01_n1016, _AES_ENC_us01_n1015, _AES_ENC_us01_n1014, _AES_ENC_us01_n1013, _AES_ENC_us01_n1012, _AES_ENC_us01_n1011, _AES_ENC_us01_n1010, _AES_ENC_us01_n1009, _AES_ENC_us01_n1008, _AES_ENC_us01_n1007, _AES_ENC_us01_n1006, _AES_ENC_us01_n1005, _AES_ENC_us01_n1004, _AES_ENC_us01_n1003, _AES_ENC_us01_n1002, _AES_ENC_us01_n1001, _AES_ENC_us01_n1000, _AES_ENC_us01_n999, _AES_ENC_us01_n998, _AES_ENC_us01_n997, _AES_ENC_us01_n996, _AES_ENC_us01_n995, _AES_ENC_us01_n994, _AES_ENC_us01_n993, _AES_ENC_us01_n992, _AES_ENC_us01_n991, _AES_ENC_us01_n990, _AES_ENC_us01_n989, _AES_ENC_us01_n988, _AES_ENC_us01_n987, _AES_ENC_us01_n986, _AES_ENC_us01_n985, _AES_ENC_us01_n984, _AES_ENC_us01_n983, _AES_ENC_us01_n982, _AES_ENC_us01_n981, _AES_ENC_us01_n980, _AES_ENC_us01_n979, _AES_ENC_us01_n978, _AES_ENC_us01_n977, _AES_ENC_us01_n976, _AES_ENC_us01_n975, _AES_ENC_us01_n974, _AES_ENC_us01_n973, _AES_ENC_us01_n972, _AES_ENC_us01_n971, 
  _AES_ENC_us01_n970, _AES_ENC_us01_n969, _AES_ENC_us01_n968, _AES_ENC_us01_n967, _AES_ENC_us01_n966, _AES_ENC_us01_n965, _AES_ENC_us01_n964, _AES_ENC_us01_n963, _AES_ENC_us01_n962, _AES_ENC_us01_n961, _AES_ENC_us01_n960, _AES_ENC_us01_n959, _AES_ENC_us01_n958, _AES_ENC_us01_n957, _AES_ENC_us01_n956, _AES_ENC_us01_n955, _AES_ENC_us01_n954, _AES_ENC_us01_n953, _AES_ENC_us01_n952, _AES_ENC_us01_n951, _AES_ENC_us01_n950, _AES_ENC_us01_n949, _AES_ENC_us01_n948, _AES_ENC_us01_n947, _AES_ENC_us01_n946, _AES_ENC_us01_n945, _AES_ENC_us01_n944, _AES_ENC_us01_n943, _AES_ENC_us01_n942, _AES_ENC_us01_n941, _AES_ENC_us01_n940, _AES_ENC_us01_n939, _AES_ENC_us01_n938, _AES_ENC_us01_n937, _AES_ENC_us01_n936, _AES_ENC_us01_n935, _AES_ENC_us01_n934, _AES_ENC_us01_n933, _AES_ENC_us01_n932, _AES_ENC_us01_n931, _AES_ENC_us01_n930, _AES_ENC_us01_n929, _AES_ENC_us01_n928, _AES_ENC_us01_n927, _AES_ENC_us01_n926, _AES_ENC_us01_n925, _AES_ENC_us01_n924, _AES_ENC_us01_n923, _AES_ENC_us01_n922, _AES_ENC_us01_n921, 
  _AES_ENC_us01_n920, _AES_ENC_us01_n919, _AES_ENC_us01_n918, _AES_ENC_us01_n917, _AES_ENC_us01_n916, _AES_ENC_us01_n915, _AES_ENC_us01_n914, _AES_ENC_us01_n913, _AES_ENC_us01_n912, _AES_ENC_us01_n911, _AES_ENC_us01_n910, _AES_ENC_us01_n909, _AES_ENC_us01_n908, _AES_ENC_us01_n907, _AES_ENC_us01_n906, _AES_ENC_us01_n905, _AES_ENC_us01_n904, _AES_ENC_us01_n903, _AES_ENC_us01_n902, _AES_ENC_us01_n901, _AES_ENC_us01_n900, _AES_ENC_us01_n899, _AES_ENC_us01_n898, _AES_ENC_us01_n897, _AES_ENC_us01_n896, _AES_ENC_us01_n895, _AES_ENC_us01_n894, _AES_ENC_us01_n893, _AES_ENC_us01_n892, _AES_ENC_us01_n891, _AES_ENC_us01_n890, _AES_ENC_us01_n889, _AES_ENC_us01_n888, _AES_ENC_us01_n887, _AES_ENC_us01_n886, _AES_ENC_us01_n885, _AES_ENC_us01_n884, _AES_ENC_us01_n883, _AES_ENC_us01_n882, _AES_ENC_us01_n881, _AES_ENC_us01_n880, _AES_ENC_us01_n879, _AES_ENC_us01_n878, _AES_ENC_us01_n877, _AES_ENC_us01_n876, _AES_ENC_us01_n875, _AES_ENC_us01_n874, _AES_ENC_us01_n873, _AES_ENC_us01_n872, _AES_ENC_us01_n871, 
  _AES_ENC_us01_n870, _AES_ENC_us01_n869, _AES_ENC_us01_n868, _AES_ENC_us01_n867, _AES_ENC_us01_n866, _AES_ENC_us01_n865, _AES_ENC_us01_n864, _AES_ENC_us01_n863, _AES_ENC_us01_n862, _AES_ENC_us01_n861, _AES_ENC_us01_n860, _AES_ENC_us01_n859, _AES_ENC_us01_n858, _AES_ENC_us01_n857, _AES_ENC_us01_n856, _AES_ENC_us01_n855, _AES_ENC_us01_n854, _AES_ENC_us01_n853, _AES_ENC_us01_n852, _AES_ENC_us01_n851, _AES_ENC_us01_n850, _AES_ENC_us01_n849, _AES_ENC_us01_n848, _AES_ENC_us01_n847, _AES_ENC_us01_n846, _AES_ENC_us01_n845, _AES_ENC_us01_n844, _AES_ENC_us01_n843, _AES_ENC_us01_n842, _AES_ENC_us01_n841, _AES_ENC_us01_n840, _AES_ENC_us01_n839, _AES_ENC_us01_n838, _AES_ENC_us01_n837, _AES_ENC_us01_n836, _AES_ENC_us01_n835, _AES_ENC_us01_n834, _AES_ENC_us01_n833, _AES_ENC_us01_n832, _AES_ENC_us01_n831, _AES_ENC_us01_n830, _AES_ENC_us01_n829, _AES_ENC_us01_n828, _AES_ENC_us01_n827, _AES_ENC_us01_n826, _AES_ENC_us01_n825, _AES_ENC_us01_n824, _AES_ENC_us01_n823, _AES_ENC_us01_n822, _AES_ENC_us01_n821, 
  _AES_ENC_us01_n820, _AES_ENC_us01_n819, _AES_ENC_us01_n818, _AES_ENC_us01_n817, _AES_ENC_us01_n816, _AES_ENC_us01_n815, _AES_ENC_us01_n814, _AES_ENC_us01_n813, _AES_ENC_us01_n812, _AES_ENC_us01_n811, _AES_ENC_us01_n810, _AES_ENC_us01_n809, _AES_ENC_us01_n808, _AES_ENC_us01_n807, _AES_ENC_us01_n806, _AES_ENC_us01_n805, _AES_ENC_us01_n804, _AES_ENC_us01_n803, _AES_ENC_us01_n802, _AES_ENC_us01_n801, _AES_ENC_us01_n800, _AES_ENC_us01_n799, _AES_ENC_us01_n798, _AES_ENC_us01_n797, _AES_ENC_us01_n796, _AES_ENC_us01_n795, _AES_ENC_us01_n794, _AES_ENC_us01_n793, _AES_ENC_us01_n792, _AES_ENC_us01_n791, _AES_ENC_us01_n790, _AES_ENC_us01_n789, _AES_ENC_us01_n788, _AES_ENC_us01_n787, _AES_ENC_us01_n786, _AES_ENC_us01_n785, _AES_ENC_us01_n784, _AES_ENC_us01_n783, _AES_ENC_us01_n782, _AES_ENC_us01_n781, _AES_ENC_us01_n780, _AES_ENC_us01_n779, _AES_ENC_us01_n778, _AES_ENC_us01_n777, _AES_ENC_us01_n776, _AES_ENC_us01_n775, _AES_ENC_us01_n774, _AES_ENC_us01_n773, _AES_ENC_us01_n772, _AES_ENC_us01_n771, 
  _AES_ENC_us01_n770, _AES_ENC_us01_n769, _AES_ENC_us01_n768, _AES_ENC_us01_n767, _AES_ENC_us01_n766, _AES_ENC_us01_n765, _AES_ENC_us01_n764, _AES_ENC_us01_n763, _AES_ENC_us01_n762, _AES_ENC_us01_n761, _AES_ENC_us01_n760, _AES_ENC_us01_n759, _AES_ENC_us01_n758, _AES_ENC_us01_n757, _AES_ENC_us01_n756, _AES_ENC_us01_n755, _AES_ENC_us01_n754, _AES_ENC_us01_n753, _AES_ENC_us01_n752, _AES_ENC_us01_n751, _AES_ENC_us01_n750, _AES_ENC_us01_n749, _AES_ENC_us01_n748, _AES_ENC_us01_n747, _AES_ENC_us01_n746, _AES_ENC_us01_n745, _AES_ENC_us01_n744, _AES_ENC_us01_n743, _AES_ENC_us01_n742, _AES_ENC_us01_n741, _AES_ENC_us01_n740, _AES_ENC_us01_n739, _AES_ENC_us01_n738, _AES_ENC_us01_n737, _AES_ENC_us01_n736, _AES_ENC_us01_n735, _AES_ENC_us01_n734, _AES_ENC_us01_n733, _AES_ENC_us01_n732, _AES_ENC_us01_n731, _AES_ENC_us01_n730, _AES_ENC_us01_n729, _AES_ENC_us01_n728, _AES_ENC_us01_n727, _AES_ENC_us01_n726, _AES_ENC_us01_n725, _AES_ENC_us01_n724, _AES_ENC_us01_n723, _AES_ENC_us01_n722, _AES_ENC_us01_n721, 
  _AES_ENC_us01_n720, _AES_ENC_us01_n719, _AES_ENC_us01_n718, _AES_ENC_us01_n717, _AES_ENC_us01_n716, _AES_ENC_us01_n715, _AES_ENC_us01_n714, _AES_ENC_us01_n713, _AES_ENC_us01_n712, _AES_ENC_us01_n711, _AES_ENC_us01_n710, _AES_ENC_us01_n709, _AES_ENC_us01_n708, _AES_ENC_us01_n707, _AES_ENC_us01_n706, _AES_ENC_us01_n705, _AES_ENC_us01_n704, _AES_ENC_us01_n703, _AES_ENC_us01_n702, _AES_ENC_us01_n701, _AES_ENC_us01_n700, _AES_ENC_us01_n699, _AES_ENC_us01_n698, _AES_ENC_us01_n697, _AES_ENC_us01_n696, _AES_ENC_us01_n695, _AES_ENC_us01_n694, _AES_ENC_us01_n693, _AES_ENC_us01_n692, _AES_ENC_us01_n691, _AES_ENC_us01_n690, _AES_ENC_us01_n689, _AES_ENC_us01_n688, _AES_ENC_us01_n687, _AES_ENC_us01_n686, _AES_ENC_us01_n685, _AES_ENC_us01_n684, _AES_ENC_us01_n683, _AES_ENC_us01_n682, _AES_ENC_us01_n681, _AES_ENC_us01_n680, _AES_ENC_us01_n679, _AES_ENC_us01_n678, _AES_ENC_us01_n677, _AES_ENC_us01_n676, _AES_ENC_us01_n675, _AES_ENC_us01_n674, _AES_ENC_us01_n673, _AES_ENC_us01_n672, _AES_ENC_us01_n671, 
  _AES_ENC_us01_n670, _AES_ENC_us01_n669, _AES_ENC_us01_n668, _AES_ENC_us01_n667, _AES_ENC_us01_n666, _AES_ENC_us01_n665, _AES_ENC_us01_n664, _AES_ENC_us01_n663, _AES_ENC_us01_n662, _AES_ENC_us01_n661, _AES_ENC_us01_n660, _AES_ENC_us01_n659, _AES_ENC_us01_n658, _AES_ENC_us01_n657, _AES_ENC_us01_n656, _AES_ENC_us01_n655, _AES_ENC_us01_n654, _AES_ENC_us01_n653, _AES_ENC_us01_n652, _AES_ENC_us01_n651, _AES_ENC_us01_n650, _AES_ENC_us01_n649, _AES_ENC_us01_n648, _AES_ENC_us01_n647, _AES_ENC_us01_n646, _AES_ENC_us01_n645, _AES_ENC_us01_n644, _AES_ENC_us01_n643, _AES_ENC_us01_n642, _AES_ENC_us01_n641, _AES_ENC_us01_n640, _AES_ENC_us01_n639, _AES_ENC_us01_n638, _AES_ENC_us01_n637, _AES_ENC_us01_n636, _AES_ENC_us01_n635, _AES_ENC_us01_n634, _AES_ENC_us01_n633, _AES_ENC_us01_n632, _AES_ENC_us01_n631, _AES_ENC_us01_n630, _AES_ENC_us01_n629, _AES_ENC_us01_n628, _AES_ENC_us01_n627, _AES_ENC_us01_n626, _AES_ENC_us01_n625, _AES_ENC_us01_n624, _AES_ENC_us01_n623, _AES_ENC_us01_n622, _AES_ENC_us01_n621, 
  _AES_ENC_us01_n620, _AES_ENC_us01_n619, _AES_ENC_us01_n618, _AES_ENC_us01_n617, _AES_ENC_us01_n616, _AES_ENC_us01_n615, _AES_ENC_us01_n614, _AES_ENC_us01_n613, _AES_ENC_us01_n612, _AES_ENC_us01_n611, _AES_ENC_us01_n610, _AES_ENC_us01_n609, _AES_ENC_us01_n608, _AES_ENC_us01_n607, _AES_ENC_us01_n606, _AES_ENC_us01_n605, _AES_ENC_us01_n604, _AES_ENC_us01_n603, _AES_ENC_us01_n602, _AES_ENC_us01_n601, _AES_ENC_us01_n600, _AES_ENC_us01_n599, _AES_ENC_us01_n598, _AES_ENC_us01_n597, _AES_ENC_us01_n596, _AES_ENC_us01_n595, _AES_ENC_us01_n594, _AES_ENC_us01_n593, _AES_ENC_us01_n592, _AES_ENC_us01_n591, _AES_ENC_us01_n590, _AES_ENC_us01_n589, _AES_ENC_us01_n588, _AES_ENC_us01_n587, _AES_ENC_us01_n586, _AES_ENC_us01_n585, _AES_ENC_us01_n584, _AES_ENC_us01_n583, _AES_ENC_us01_n582, _AES_ENC_us01_n581, _AES_ENC_us01_n580, _AES_ENC_us01_n579, _AES_ENC_us01_n578, _AES_ENC_us01_n577, _AES_ENC_us01_n576, _AES_ENC_us01_n575, _AES_ENC_us01_n574, _AES_ENC_us01_n573, _AES_ENC_us01_n572, _AES_ENC_us01_n571, 
  _AES_ENC_us01_n570, _AES_ENC_us01_n569, _AES_ENC_us02_n1135, _AES_ENC_us02_n1134, _AES_ENC_us02_n1133, _AES_ENC_us02_n1132, _AES_ENC_us02_n1131, _AES_ENC_us02_n1130, _AES_ENC_us02_n1129, _AES_ENC_us02_n1128, _AES_ENC_us02_n1127, _AES_ENC_us02_n1126, _AES_ENC_us02_n1125, _AES_ENC_us02_n1124, _AES_ENC_us02_n1123, _AES_ENC_us02_n1122, _AES_ENC_us02_n1121, _AES_ENC_us02_n1120, _AES_ENC_us02_n1119, _AES_ENC_us02_n1118, _AES_ENC_us02_n1117, _AES_ENC_us02_n1116, _AES_ENC_us02_n1115, _AES_ENC_us02_n1114, _AES_ENC_us02_n1113, _AES_ENC_us02_n1112, _AES_ENC_us02_n1111, _AES_ENC_us02_n1110, _AES_ENC_us02_n1109, _AES_ENC_us02_n1108, _AES_ENC_us02_n1107, _AES_ENC_us02_n1106, _AES_ENC_us02_n1105, _AES_ENC_us02_n1104, _AES_ENC_us02_n1103, _AES_ENC_us02_n1102, _AES_ENC_us02_n1101, _AES_ENC_us02_n1100, _AES_ENC_us02_n1099, _AES_ENC_us02_n1098, _AES_ENC_us02_n1097, _AES_ENC_us02_n1096, _AES_ENC_us02_n1095, _AES_ENC_us02_n1094, _AES_ENC_us02_n1093, _AES_ENC_us02_n1092, _AES_ENC_us02_n1091, _AES_ENC_us02_n1090, _AES_ENC_us02_n1089, _AES_ENC_us02_n1088, 
  _AES_ENC_us02_n1087, _AES_ENC_us02_n1086, _AES_ENC_us02_n1085, _AES_ENC_us02_n1084, _AES_ENC_us02_n1083, _AES_ENC_us02_n1082, _AES_ENC_us02_n1081, _AES_ENC_us02_n1080, _AES_ENC_us02_n1079, _AES_ENC_us02_n1078, _AES_ENC_us02_n1077, _AES_ENC_us02_n1076, _AES_ENC_us02_n1075, _AES_ENC_us02_n1074, _AES_ENC_us02_n1073, _AES_ENC_us02_n1072, _AES_ENC_us02_n1071, _AES_ENC_us02_n1070, _AES_ENC_us02_n1069, _AES_ENC_us02_n1068, _AES_ENC_us02_n1067, _AES_ENC_us02_n1066, _AES_ENC_us02_n1065, _AES_ENC_us02_n1064, _AES_ENC_us02_n1063, _AES_ENC_us02_n1062, _AES_ENC_us02_n1061, _AES_ENC_us02_n1060, _AES_ENC_us02_n1059, _AES_ENC_us02_n1058, _AES_ENC_us02_n1057, _AES_ENC_us02_n1056, _AES_ENC_us02_n1055, _AES_ENC_us02_n1054, _AES_ENC_us02_n1053, _AES_ENC_us02_n1052, _AES_ENC_us02_n1051, _AES_ENC_us02_n1050, _AES_ENC_us02_n1049, _AES_ENC_us02_n1048, _AES_ENC_us02_n1047, _AES_ENC_us02_n1046, _AES_ENC_us02_n1045, _AES_ENC_us02_n1044, _AES_ENC_us02_n1043, _AES_ENC_us02_n1042, _AES_ENC_us02_n1041, _AES_ENC_us02_n1040, _AES_ENC_us02_n1039, _AES_ENC_us02_n1038, 
  _AES_ENC_us02_n1037, _AES_ENC_us02_n1036, _AES_ENC_us02_n1035, _AES_ENC_us02_n1034, _AES_ENC_us02_n1033, _AES_ENC_us02_n1032, _AES_ENC_us02_n1031, _AES_ENC_us02_n1030, _AES_ENC_us02_n1029, _AES_ENC_us02_n1028, _AES_ENC_us02_n1027, _AES_ENC_us02_n1026, _AES_ENC_us02_n1025, _AES_ENC_us02_n1024, _AES_ENC_us02_n1023, _AES_ENC_us02_n1022, _AES_ENC_us02_n1021, _AES_ENC_us02_n1020, _AES_ENC_us02_n1019, _AES_ENC_us02_n1018, _AES_ENC_us02_n1017, _AES_ENC_us02_n1016, _AES_ENC_us02_n1015, _AES_ENC_us02_n1014, _AES_ENC_us02_n1013, _AES_ENC_us02_n1012, _AES_ENC_us02_n1011, _AES_ENC_us02_n1010, _AES_ENC_us02_n1009, _AES_ENC_us02_n1008, _AES_ENC_us02_n1007, _AES_ENC_us02_n1006, _AES_ENC_us02_n1005, _AES_ENC_us02_n1004, _AES_ENC_us02_n1003, _AES_ENC_us02_n1002, _AES_ENC_us02_n1001, _AES_ENC_us02_n1000, _AES_ENC_us02_n999, _AES_ENC_us02_n998, _AES_ENC_us02_n997, _AES_ENC_us02_n996, _AES_ENC_us02_n995, _AES_ENC_us02_n994, _AES_ENC_us02_n993, _AES_ENC_us02_n992, _AES_ENC_us02_n991, _AES_ENC_us02_n990, _AES_ENC_us02_n989, _AES_ENC_us02_n988, 
  _AES_ENC_us02_n987, _AES_ENC_us02_n986, _AES_ENC_us02_n985, _AES_ENC_us02_n984, _AES_ENC_us02_n983, _AES_ENC_us02_n982, _AES_ENC_us02_n981, _AES_ENC_us02_n980, _AES_ENC_us02_n979, _AES_ENC_us02_n978, _AES_ENC_us02_n977, _AES_ENC_us02_n976, _AES_ENC_us02_n975, _AES_ENC_us02_n974, _AES_ENC_us02_n973, _AES_ENC_us02_n972, _AES_ENC_us02_n971, _AES_ENC_us02_n970, _AES_ENC_us02_n969, _AES_ENC_us02_n968, _AES_ENC_us02_n967, _AES_ENC_us02_n966, _AES_ENC_us02_n965, _AES_ENC_us02_n964, _AES_ENC_us02_n963, _AES_ENC_us02_n962, _AES_ENC_us02_n961, _AES_ENC_us02_n960, _AES_ENC_us02_n959, _AES_ENC_us02_n958, _AES_ENC_us02_n957, _AES_ENC_us02_n956, _AES_ENC_us02_n955, _AES_ENC_us02_n954, _AES_ENC_us02_n953, _AES_ENC_us02_n952, _AES_ENC_us02_n951, _AES_ENC_us02_n950, _AES_ENC_us02_n949, _AES_ENC_us02_n948, _AES_ENC_us02_n947, _AES_ENC_us02_n946, _AES_ENC_us02_n945, _AES_ENC_us02_n944, _AES_ENC_us02_n943, _AES_ENC_us02_n942, _AES_ENC_us02_n941, _AES_ENC_us02_n940, _AES_ENC_us02_n939, _AES_ENC_us02_n938, 
  _AES_ENC_us02_n937, _AES_ENC_us02_n936, _AES_ENC_us02_n935, _AES_ENC_us02_n934, _AES_ENC_us02_n933, _AES_ENC_us02_n932, _AES_ENC_us02_n931, _AES_ENC_us02_n930, _AES_ENC_us02_n929, _AES_ENC_us02_n928, _AES_ENC_us02_n927, _AES_ENC_us02_n926, _AES_ENC_us02_n925, _AES_ENC_us02_n924, _AES_ENC_us02_n923, _AES_ENC_us02_n922, _AES_ENC_us02_n921, _AES_ENC_us02_n920, _AES_ENC_us02_n919, _AES_ENC_us02_n918, _AES_ENC_us02_n917, _AES_ENC_us02_n916, _AES_ENC_us02_n915, _AES_ENC_us02_n914, _AES_ENC_us02_n913, _AES_ENC_us02_n912, _AES_ENC_us02_n911, _AES_ENC_us02_n910, _AES_ENC_us02_n909, _AES_ENC_us02_n908, _AES_ENC_us02_n907, _AES_ENC_us02_n906, _AES_ENC_us02_n905, _AES_ENC_us02_n904, _AES_ENC_us02_n903, _AES_ENC_us02_n902, _AES_ENC_us02_n901, _AES_ENC_us02_n900, _AES_ENC_us02_n899, _AES_ENC_us02_n898, _AES_ENC_us02_n897, _AES_ENC_us02_n896, _AES_ENC_us02_n895, _AES_ENC_us02_n894, _AES_ENC_us02_n893, _AES_ENC_us02_n892, _AES_ENC_us02_n891, _AES_ENC_us02_n890, _AES_ENC_us02_n889, _AES_ENC_us02_n888, 
  _AES_ENC_us02_n887, _AES_ENC_us02_n886, _AES_ENC_us02_n885, _AES_ENC_us02_n884, _AES_ENC_us02_n883, _AES_ENC_us02_n882, _AES_ENC_us02_n881, _AES_ENC_us02_n880, _AES_ENC_us02_n879, _AES_ENC_us02_n878, _AES_ENC_us02_n877, _AES_ENC_us02_n876, _AES_ENC_us02_n875, _AES_ENC_us02_n874, _AES_ENC_us02_n873, _AES_ENC_us02_n872, _AES_ENC_us02_n871, _AES_ENC_us02_n870, _AES_ENC_us02_n869, _AES_ENC_us02_n868, _AES_ENC_us02_n867, _AES_ENC_us02_n866, _AES_ENC_us02_n865, _AES_ENC_us02_n864, _AES_ENC_us02_n863, _AES_ENC_us02_n862, _AES_ENC_us02_n861, _AES_ENC_us02_n860, _AES_ENC_us02_n859, _AES_ENC_us02_n858, _AES_ENC_us02_n857, _AES_ENC_us02_n856, _AES_ENC_us02_n855, _AES_ENC_us02_n854, _AES_ENC_us02_n853, _AES_ENC_us02_n852, _AES_ENC_us02_n851, _AES_ENC_us02_n850, _AES_ENC_us02_n849, _AES_ENC_us02_n848, _AES_ENC_us02_n847, _AES_ENC_us02_n846, _AES_ENC_us02_n845, _AES_ENC_us02_n844, _AES_ENC_us02_n843, _AES_ENC_us02_n842, _AES_ENC_us02_n841, _AES_ENC_us02_n840, _AES_ENC_us02_n839, _AES_ENC_us02_n838, 
  _AES_ENC_us02_n837, _AES_ENC_us02_n836, _AES_ENC_us02_n835, _AES_ENC_us02_n834, _AES_ENC_us02_n833, _AES_ENC_us02_n832, _AES_ENC_us02_n831, _AES_ENC_us02_n830, _AES_ENC_us02_n829, _AES_ENC_us02_n828, _AES_ENC_us02_n827, _AES_ENC_us02_n826, _AES_ENC_us02_n825, _AES_ENC_us02_n824, _AES_ENC_us02_n823, _AES_ENC_us02_n822, _AES_ENC_us02_n821, _AES_ENC_us02_n820, _AES_ENC_us02_n819, _AES_ENC_us02_n818, _AES_ENC_us02_n817, _AES_ENC_us02_n816, _AES_ENC_us02_n815, _AES_ENC_us02_n814, _AES_ENC_us02_n813, _AES_ENC_us02_n812, _AES_ENC_us02_n811, _AES_ENC_us02_n810, _AES_ENC_us02_n809, _AES_ENC_us02_n808, _AES_ENC_us02_n807, _AES_ENC_us02_n806, _AES_ENC_us02_n805, _AES_ENC_us02_n804, _AES_ENC_us02_n803, _AES_ENC_us02_n802, _AES_ENC_us02_n801, _AES_ENC_us02_n800, _AES_ENC_us02_n799, _AES_ENC_us02_n798, _AES_ENC_us02_n797, _AES_ENC_us02_n796, _AES_ENC_us02_n795, _AES_ENC_us02_n794, _AES_ENC_us02_n793, _AES_ENC_us02_n792, _AES_ENC_us02_n791, _AES_ENC_us02_n790, _AES_ENC_us02_n789, _AES_ENC_us02_n788, 
  _AES_ENC_us02_n787, _AES_ENC_us02_n786, _AES_ENC_us02_n785, _AES_ENC_us02_n784, _AES_ENC_us02_n783, _AES_ENC_us02_n782, _AES_ENC_us02_n781, _AES_ENC_us02_n780, _AES_ENC_us02_n779, _AES_ENC_us02_n778, _AES_ENC_us02_n777, _AES_ENC_us02_n776, _AES_ENC_us02_n775, _AES_ENC_us02_n774, _AES_ENC_us02_n773, _AES_ENC_us02_n772, _AES_ENC_us02_n771, _AES_ENC_us02_n770, _AES_ENC_us02_n769, _AES_ENC_us02_n768, _AES_ENC_us02_n767, _AES_ENC_us02_n766, _AES_ENC_us02_n765, _AES_ENC_us02_n764, _AES_ENC_us02_n763, _AES_ENC_us02_n762, _AES_ENC_us02_n761, _AES_ENC_us02_n760, _AES_ENC_us02_n759, _AES_ENC_us02_n758, _AES_ENC_us02_n757, _AES_ENC_us02_n756, _AES_ENC_us02_n755, _AES_ENC_us02_n754, _AES_ENC_us02_n753, _AES_ENC_us02_n752, _AES_ENC_us02_n751, _AES_ENC_us02_n750, _AES_ENC_us02_n749, _AES_ENC_us02_n748, _AES_ENC_us02_n747, _AES_ENC_us02_n746, _AES_ENC_us02_n745, _AES_ENC_us02_n744, _AES_ENC_us02_n743, _AES_ENC_us02_n742, _AES_ENC_us02_n741, _AES_ENC_us02_n740, _AES_ENC_us02_n739, _AES_ENC_us02_n738, 
  _AES_ENC_us02_n737, _AES_ENC_us02_n736, _AES_ENC_us02_n735, _AES_ENC_us02_n734, _AES_ENC_us02_n733, _AES_ENC_us02_n732, _AES_ENC_us02_n731, _AES_ENC_us02_n730, _AES_ENC_us02_n729, _AES_ENC_us02_n728, _AES_ENC_us02_n727, _AES_ENC_us02_n726, _AES_ENC_us02_n725, _AES_ENC_us02_n724, _AES_ENC_us02_n723, _AES_ENC_us02_n722, _AES_ENC_us02_n721, _AES_ENC_us02_n720, _AES_ENC_us02_n719, _AES_ENC_us02_n718, _AES_ENC_us02_n717, _AES_ENC_us02_n716, _AES_ENC_us02_n715, _AES_ENC_us02_n714, _AES_ENC_us02_n713, _AES_ENC_us02_n712, _AES_ENC_us02_n711, _AES_ENC_us02_n710, _AES_ENC_us02_n709, _AES_ENC_us02_n708, _AES_ENC_us02_n707, _AES_ENC_us02_n706, _AES_ENC_us02_n705, _AES_ENC_us02_n704, _AES_ENC_us02_n703, _AES_ENC_us02_n702, _AES_ENC_us02_n701, _AES_ENC_us02_n700, _AES_ENC_us02_n699, _AES_ENC_us02_n698, _AES_ENC_us02_n697, _AES_ENC_us02_n696, _AES_ENC_us02_n695, _AES_ENC_us02_n694, _AES_ENC_us02_n693, _AES_ENC_us02_n692, _AES_ENC_us02_n691, _AES_ENC_us02_n690, _AES_ENC_us02_n689, _AES_ENC_us02_n688, 
  _AES_ENC_us02_n687, _AES_ENC_us02_n686, _AES_ENC_us02_n685, _AES_ENC_us02_n684, _AES_ENC_us02_n683, _AES_ENC_us02_n682, _AES_ENC_us02_n681, _AES_ENC_us02_n680, _AES_ENC_us02_n679, _AES_ENC_us02_n678, _AES_ENC_us02_n677, _AES_ENC_us02_n676, _AES_ENC_us02_n675, _AES_ENC_us02_n674, _AES_ENC_us02_n673, _AES_ENC_us02_n672, _AES_ENC_us02_n671, _AES_ENC_us02_n670, _AES_ENC_us02_n669, _AES_ENC_us02_n668, _AES_ENC_us02_n667, _AES_ENC_us02_n666, _AES_ENC_us02_n665, _AES_ENC_us02_n664, _AES_ENC_us02_n663, _AES_ENC_us02_n662, _AES_ENC_us02_n661, _AES_ENC_us02_n660, _AES_ENC_us02_n659, _AES_ENC_us02_n658, _AES_ENC_us02_n657, _AES_ENC_us02_n656, _AES_ENC_us02_n655, _AES_ENC_us02_n654, _AES_ENC_us02_n653, _AES_ENC_us02_n652, _AES_ENC_us02_n651, _AES_ENC_us02_n650, _AES_ENC_us02_n649, _AES_ENC_us02_n648, _AES_ENC_us02_n647, _AES_ENC_us02_n646, _AES_ENC_us02_n645, _AES_ENC_us02_n644, _AES_ENC_us02_n643, _AES_ENC_us02_n642, _AES_ENC_us02_n641, _AES_ENC_us02_n640, _AES_ENC_us02_n639, _AES_ENC_us02_n638, 
  _AES_ENC_us02_n637, _AES_ENC_us02_n636, _AES_ENC_us02_n635, _AES_ENC_us02_n634, _AES_ENC_us02_n633, _AES_ENC_us02_n632, _AES_ENC_us02_n631, _AES_ENC_us02_n630, _AES_ENC_us02_n629, _AES_ENC_us02_n628, _AES_ENC_us02_n627, _AES_ENC_us02_n626, _AES_ENC_us02_n625, _AES_ENC_us02_n624, _AES_ENC_us02_n623, _AES_ENC_us02_n622, _AES_ENC_us02_n621, _AES_ENC_us02_n620, _AES_ENC_us02_n619, _AES_ENC_us02_n618, _AES_ENC_us02_n617, _AES_ENC_us02_n616, _AES_ENC_us02_n615, _AES_ENC_us02_n614, _AES_ENC_us02_n613, _AES_ENC_us02_n612, _AES_ENC_us02_n611, _AES_ENC_us02_n610, _AES_ENC_us02_n609, _AES_ENC_us02_n608, _AES_ENC_us02_n607, _AES_ENC_us02_n606, _AES_ENC_us02_n605, _AES_ENC_us02_n604, _AES_ENC_us02_n603, _AES_ENC_us02_n602, _AES_ENC_us02_n601, _AES_ENC_us02_n600, _AES_ENC_us02_n599, _AES_ENC_us02_n598, _AES_ENC_us02_n597, _AES_ENC_us02_n596, _AES_ENC_us02_n595, _AES_ENC_us02_n594, _AES_ENC_us02_n593, _AES_ENC_us02_n592, _AES_ENC_us02_n591, _AES_ENC_us02_n590, _AES_ENC_us02_n589, _AES_ENC_us02_n588, 
  _AES_ENC_us02_n587, _AES_ENC_us02_n586, _AES_ENC_us02_n585, _AES_ENC_us02_n584, _AES_ENC_us02_n583, _AES_ENC_us02_n582, _AES_ENC_us02_n581, _AES_ENC_us02_n580, _AES_ENC_us02_n579, _AES_ENC_us02_n578, _AES_ENC_us02_n577, _AES_ENC_us02_n576, _AES_ENC_us02_n575, _AES_ENC_us02_n574, _AES_ENC_us02_n573, _AES_ENC_us02_n572, _AES_ENC_us02_n571, _AES_ENC_us02_n570, _AES_ENC_us02_n569, _AES_ENC_us03_n1135, _AES_ENC_us03_n1134, _AES_ENC_us03_n1133, _AES_ENC_us03_n1132, _AES_ENC_us03_n1131, _AES_ENC_us03_n1130, _AES_ENC_us03_n1129, _AES_ENC_us03_n1128, _AES_ENC_us03_n1127, _AES_ENC_us03_n1126, _AES_ENC_us03_n1125, _AES_ENC_us03_n1124, _AES_ENC_us03_n1123, _AES_ENC_us03_n1122, _AES_ENC_us03_n1121, _AES_ENC_us03_n1120, _AES_ENC_us03_n1119, _AES_ENC_us03_n1118, _AES_ENC_us03_n1117, _AES_ENC_us03_n1116, _AES_ENC_us03_n1115, _AES_ENC_us03_n1114, _AES_ENC_us03_n1113, _AES_ENC_us03_n1112, _AES_ENC_us03_n1111, _AES_ENC_us03_n1110, _AES_ENC_us03_n1109, _AES_ENC_us03_n1108, _AES_ENC_us03_n1107, _AES_ENC_us03_n1106, _AES_ENC_us03_n1105, 
  _AES_ENC_us03_n1104, _AES_ENC_us03_n1103, _AES_ENC_us03_n1102, _AES_ENC_us03_n1101, _AES_ENC_us03_n1100, _AES_ENC_us03_n1099, _AES_ENC_us03_n1098, _AES_ENC_us03_n1097, _AES_ENC_us03_n1096, _AES_ENC_us03_n1095, _AES_ENC_us03_n1094, _AES_ENC_us03_n1093, _AES_ENC_us03_n1092, _AES_ENC_us03_n1091, _AES_ENC_us03_n1090, _AES_ENC_us03_n1089, _AES_ENC_us03_n1088, _AES_ENC_us03_n1087, _AES_ENC_us03_n1086, _AES_ENC_us03_n1085, _AES_ENC_us03_n1084, _AES_ENC_us03_n1083, _AES_ENC_us03_n1082, _AES_ENC_us03_n1081, _AES_ENC_us03_n1080, _AES_ENC_us03_n1079, _AES_ENC_us03_n1078, _AES_ENC_us03_n1077, _AES_ENC_us03_n1076, _AES_ENC_us03_n1075, _AES_ENC_us03_n1074, _AES_ENC_us03_n1073, _AES_ENC_us03_n1072, _AES_ENC_us03_n1071, _AES_ENC_us03_n1070, _AES_ENC_us03_n1069, _AES_ENC_us03_n1068, _AES_ENC_us03_n1067, _AES_ENC_us03_n1066, _AES_ENC_us03_n1065, _AES_ENC_us03_n1064, _AES_ENC_us03_n1063, _AES_ENC_us03_n1062, _AES_ENC_us03_n1061, _AES_ENC_us03_n1060, _AES_ENC_us03_n1059, _AES_ENC_us03_n1058, _AES_ENC_us03_n1057, _AES_ENC_us03_n1056, _AES_ENC_us03_n1055, 
  _AES_ENC_us03_n1054, _AES_ENC_us03_n1053, _AES_ENC_us03_n1052, _AES_ENC_us03_n1051, _AES_ENC_us03_n1050, _AES_ENC_us03_n1049, _AES_ENC_us03_n1048, _AES_ENC_us03_n1047, _AES_ENC_us03_n1046, _AES_ENC_us03_n1045, _AES_ENC_us03_n1044, _AES_ENC_us03_n1043, _AES_ENC_us03_n1042, _AES_ENC_us03_n1041, _AES_ENC_us03_n1040, _AES_ENC_us03_n1039, _AES_ENC_us03_n1038, _AES_ENC_us03_n1037, _AES_ENC_us03_n1036, _AES_ENC_us03_n1035, _AES_ENC_us03_n1034, _AES_ENC_us03_n1033, _AES_ENC_us03_n1032, _AES_ENC_us03_n1031, _AES_ENC_us03_n1030, _AES_ENC_us03_n1029, _AES_ENC_us03_n1028, _AES_ENC_us03_n1027, _AES_ENC_us03_n1026, _AES_ENC_us03_n1025, _AES_ENC_us03_n1024, _AES_ENC_us03_n1023, _AES_ENC_us03_n1022, _AES_ENC_us03_n1021, _AES_ENC_us03_n1020, _AES_ENC_us03_n1019, _AES_ENC_us03_n1018, _AES_ENC_us03_n1017, _AES_ENC_us03_n1016, _AES_ENC_us03_n1015, _AES_ENC_us03_n1014, _AES_ENC_us03_n1013, _AES_ENC_us03_n1012, _AES_ENC_us03_n1011, _AES_ENC_us03_n1010, _AES_ENC_us03_n1009, _AES_ENC_us03_n1008, _AES_ENC_us03_n1007, _AES_ENC_us03_n1006, _AES_ENC_us03_n1005, 
  _AES_ENC_us03_n1004, _AES_ENC_us03_n1003, _AES_ENC_us03_n1002, _AES_ENC_us03_n1001, _AES_ENC_us03_n1000, _AES_ENC_us03_n999, _AES_ENC_us03_n998, _AES_ENC_us03_n997, _AES_ENC_us03_n996, _AES_ENC_us03_n995, _AES_ENC_us03_n994, _AES_ENC_us03_n993, _AES_ENC_us03_n992, _AES_ENC_us03_n991, _AES_ENC_us03_n990, _AES_ENC_us03_n989, _AES_ENC_us03_n988, _AES_ENC_us03_n987, _AES_ENC_us03_n986, _AES_ENC_us03_n985, _AES_ENC_us03_n984, _AES_ENC_us03_n983, _AES_ENC_us03_n982, _AES_ENC_us03_n981, _AES_ENC_us03_n980, _AES_ENC_us03_n979, _AES_ENC_us03_n978, _AES_ENC_us03_n977, _AES_ENC_us03_n976, _AES_ENC_us03_n975, _AES_ENC_us03_n974, _AES_ENC_us03_n973, _AES_ENC_us03_n972, _AES_ENC_us03_n971, _AES_ENC_us03_n970, _AES_ENC_us03_n969, _AES_ENC_us03_n968, _AES_ENC_us03_n967, _AES_ENC_us03_n966, _AES_ENC_us03_n965, _AES_ENC_us03_n964, _AES_ENC_us03_n963, _AES_ENC_us03_n962, _AES_ENC_us03_n961, _AES_ENC_us03_n960, _AES_ENC_us03_n959, _AES_ENC_us03_n958, _AES_ENC_us03_n957, _AES_ENC_us03_n956, _AES_ENC_us03_n955, 
  _AES_ENC_us03_n954, _AES_ENC_us03_n953, _AES_ENC_us03_n952, _AES_ENC_us03_n951, _AES_ENC_us03_n950, _AES_ENC_us03_n949, _AES_ENC_us03_n948, _AES_ENC_us03_n947, _AES_ENC_us03_n946, _AES_ENC_us03_n945, _AES_ENC_us03_n944, _AES_ENC_us03_n943, _AES_ENC_us03_n942, _AES_ENC_us03_n941, _AES_ENC_us03_n940, _AES_ENC_us03_n939, _AES_ENC_us03_n938, _AES_ENC_us03_n937, _AES_ENC_us03_n936, _AES_ENC_us03_n935, _AES_ENC_us03_n934, _AES_ENC_us03_n933, _AES_ENC_us03_n932, _AES_ENC_us03_n931, _AES_ENC_us03_n930, _AES_ENC_us03_n929, _AES_ENC_us03_n928, _AES_ENC_us03_n927, _AES_ENC_us03_n926, _AES_ENC_us03_n925, _AES_ENC_us03_n924, _AES_ENC_us03_n923, _AES_ENC_us03_n922, _AES_ENC_us03_n921, _AES_ENC_us03_n920, _AES_ENC_us03_n919, _AES_ENC_us03_n918, _AES_ENC_us03_n917, _AES_ENC_us03_n916, _AES_ENC_us03_n915, _AES_ENC_us03_n914, _AES_ENC_us03_n913, _AES_ENC_us03_n912, _AES_ENC_us03_n911, _AES_ENC_us03_n910, _AES_ENC_us03_n909, _AES_ENC_us03_n908, _AES_ENC_us03_n907, _AES_ENC_us03_n906, _AES_ENC_us03_n905, 
  _AES_ENC_us03_n904, _AES_ENC_us03_n903, _AES_ENC_us03_n902, _AES_ENC_us03_n901, _AES_ENC_us03_n900, _AES_ENC_us03_n899, _AES_ENC_us03_n898, _AES_ENC_us03_n897, _AES_ENC_us03_n896, _AES_ENC_us03_n895, _AES_ENC_us03_n894, _AES_ENC_us03_n893, _AES_ENC_us03_n892, _AES_ENC_us03_n891, _AES_ENC_us03_n890, _AES_ENC_us03_n889, _AES_ENC_us03_n888, _AES_ENC_us03_n887, _AES_ENC_us03_n886, _AES_ENC_us03_n885, _AES_ENC_us03_n884, _AES_ENC_us03_n883, _AES_ENC_us03_n882, _AES_ENC_us03_n881, _AES_ENC_us03_n880, _AES_ENC_us03_n879, _AES_ENC_us03_n878, _AES_ENC_us03_n877, _AES_ENC_us03_n876, _AES_ENC_us03_n875, _AES_ENC_us03_n874, _AES_ENC_us03_n873, _AES_ENC_us03_n872, _AES_ENC_us03_n871, _AES_ENC_us03_n870, _AES_ENC_us03_n869, _AES_ENC_us03_n868, _AES_ENC_us03_n867, _AES_ENC_us03_n866, _AES_ENC_us03_n865, _AES_ENC_us03_n864, _AES_ENC_us03_n863, _AES_ENC_us03_n862, _AES_ENC_us03_n861, _AES_ENC_us03_n860, _AES_ENC_us03_n859, _AES_ENC_us03_n858, _AES_ENC_us03_n857, _AES_ENC_us03_n856, _AES_ENC_us03_n855, 
  _AES_ENC_us03_n854, _AES_ENC_us03_n853, _AES_ENC_us03_n852, _AES_ENC_us03_n851, _AES_ENC_us03_n850, _AES_ENC_us03_n849, _AES_ENC_us03_n848, _AES_ENC_us03_n847, _AES_ENC_us03_n846, _AES_ENC_us03_n845, _AES_ENC_us03_n844, _AES_ENC_us03_n843, _AES_ENC_us03_n842, _AES_ENC_us03_n841, _AES_ENC_us03_n840, _AES_ENC_us03_n839, _AES_ENC_us03_n838, _AES_ENC_us03_n837, _AES_ENC_us03_n836, _AES_ENC_us03_n835, _AES_ENC_us03_n834, _AES_ENC_us03_n833, _AES_ENC_us03_n832, _AES_ENC_us03_n831, _AES_ENC_us03_n830, _AES_ENC_us03_n829, _AES_ENC_us03_n828, _AES_ENC_us03_n827, _AES_ENC_us03_n826, _AES_ENC_us03_n825, _AES_ENC_us03_n824, _AES_ENC_us03_n823, _AES_ENC_us03_n822, _AES_ENC_us03_n821, _AES_ENC_us03_n820, _AES_ENC_us03_n819, _AES_ENC_us03_n818, _AES_ENC_us03_n817, _AES_ENC_us03_n816, _AES_ENC_us03_n815, _AES_ENC_us03_n814, _AES_ENC_us03_n813, _AES_ENC_us03_n812, _AES_ENC_us03_n811, _AES_ENC_us03_n810, _AES_ENC_us03_n809, _AES_ENC_us03_n808, _AES_ENC_us03_n807, _AES_ENC_us03_n806, _AES_ENC_us03_n805, 
  _AES_ENC_us03_n804, _AES_ENC_us03_n803, _AES_ENC_us03_n802, _AES_ENC_us03_n801, _AES_ENC_us03_n800, _AES_ENC_us03_n799, _AES_ENC_us03_n798, _AES_ENC_us03_n797, _AES_ENC_us03_n796, _AES_ENC_us03_n795, _AES_ENC_us03_n794, _AES_ENC_us03_n793, _AES_ENC_us03_n792, _AES_ENC_us03_n791, _AES_ENC_us03_n790, _AES_ENC_us03_n789, _AES_ENC_us03_n788, _AES_ENC_us03_n787, _AES_ENC_us03_n786, _AES_ENC_us03_n785, _AES_ENC_us03_n784, _AES_ENC_us03_n783, _AES_ENC_us03_n782, _AES_ENC_us03_n781, _AES_ENC_us03_n780, _AES_ENC_us03_n779, _AES_ENC_us03_n778, _AES_ENC_us03_n777, _AES_ENC_us03_n776, _AES_ENC_us03_n775, _AES_ENC_us03_n774, _AES_ENC_us03_n773, _AES_ENC_us03_n772, _AES_ENC_us03_n771, _AES_ENC_us03_n770, _AES_ENC_us03_n769, _AES_ENC_us03_n768, _AES_ENC_us03_n767, _AES_ENC_us03_n766, _AES_ENC_us03_n765, _AES_ENC_us03_n764, _AES_ENC_us03_n763, _AES_ENC_us03_n762, _AES_ENC_us03_n761, _AES_ENC_us03_n760, _AES_ENC_us03_n759, _AES_ENC_us03_n758, _AES_ENC_us03_n757, _AES_ENC_us03_n756, _AES_ENC_us03_n755, 
  _AES_ENC_us03_n754, _AES_ENC_us03_n753, _AES_ENC_us03_n752, _AES_ENC_us03_n751, _AES_ENC_us03_n750, _AES_ENC_us03_n749, _AES_ENC_us03_n748, _AES_ENC_us03_n747, _AES_ENC_us03_n746, _AES_ENC_us03_n745, _AES_ENC_us03_n744, _AES_ENC_us03_n743, _AES_ENC_us03_n742, _AES_ENC_us03_n741, _AES_ENC_us03_n740, _AES_ENC_us03_n739, _AES_ENC_us03_n738, _AES_ENC_us03_n737, _AES_ENC_us03_n736, _AES_ENC_us03_n735, _AES_ENC_us03_n734, _AES_ENC_us03_n733, _AES_ENC_us03_n732, _AES_ENC_us03_n731, _AES_ENC_us03_n730, _AES_ENC_us03_n729, _AES_ENC_us03_n728, _AES_ENC_us03_n727, _AES_ENC_us03_n726, _AES_ENC_us03_n725, _AES_ENC_us03_n724, _AES_ENC_us03_n723, _AES_ENC_us03_n722, _AES_ENC_us03_n721, _AES_ENC_us03_n720, _AES_ENC_us03_n719, _AES_ENC_us03_n718, _AES_ENC_us03_n717, _AES_ENC_us03_n716, _AES_ENC_us03_n715, _AES_ENC_us03_n714, _AES_ENC_us03_n713, _AES_ENC_us03_n712, _AES_ENC_us03_n711, _AES_ENC_us03_n710, _AES_ENC_us03_n709, _AES_ENC_us03_n708, _AES_ENC_us03_n707, _AES_ENC_us03_n706, _AES_ENC_us03_n705, 
  _AES_ENC_us03_n704, _AES_ENC_us03_n703, _AES_ENC_us03_n702, _AES_ENC_us03_n701, _AES_ENC_us03_n700, _AES_ENC_us03_n699, _AES_ENC_us03_n698, _AES_ENC_us03_n697, _AES_ENC_us03_n696, _AES_ENC_us03_n695, _AES_ENC_us03_n694, _AES_ENC_us03_n693, _AES_ENC_us03_n692, _AES_ENC_us03_n691, _AES_ENC_us03_n690, _AES_ENC_us03_n689, _AES_ENC_us03_n688, _AES_ENC_us03_n687, _AES_ENC_us03_n686, _AES_ENC_us03_n685, _AES_ENC_us03_n684, _AES_ENC_us03_n683, _AES_ENC_us03_n682, _AES_ENC_us03_n681, _AES_ENC_us03_n680, _AES_ENC_us03_n679, _AES_ENC_us03_n678, _AES_ENC_us03_n677, _AES_ENC_us03_n676, _AES_ENC_us03_n675, _AES_ENC_us03_n674, _AES_ENC_us03_n673, _AES_ENC_us03_n672, _AES_ENC_us03_n671, _AES_ENC_us03_n670, _AES_ENC_us03_n669, _AES_ENC_us03_n668, _AES_ENC_us03_n667, _AES_ENC_us03_n666, _AES_ENC_us03_n665, _AES_ENC_us03_n664, _AES_ENC_us03_n663, _AES_ENC_us03_n662, _AES_ENC_us03_n661, _AES_ENC_us03_n660, _AES_ENC_us03_n659, _AES_ENC_us03_n658, _AES_ENC_us03_n657, _AES_ENC_us03_n656, _AES_ENC_us03_n655, 
  _AES_ENC_us03_n654, _AES_ENC_us03_n653, _AES_ENC_us03_n652, _AES_ENC_us03_n651, _AES_ENC_us03_n650, _AES_ENC_us03_n649, _AES_ENC_us03_n648, _AES_ENC_us03_n647, _AES_ENC_us03_n646, _AES_ENC_us03_n645, _AES_ENC_us03_n644, _AES_ENC_us03_n643, _AES_ENC_us03_n642, _AES_ENC_us03_n641, _AES_ENC_us03_n640, _AES_ENC_us03_n639, _AES_ENC_us03_n638, _AES_ENC_us03_n637, _AES_ENC_us03_n636, _AES_ENC_us03_n635, _AES_ENC_us03_n634, _AES_ENC_us03_n633, _AES_ENC_us03_n632, _AES_ENC_us03_n631, _AES_ENC_us03_n630, _AES_ENC_us03_n629, _AES_ENC_us03_n628, _AES_ENC_us03_n627, _AES_ENC_us03_n626, _AES_ENC_us03_n625, _AES_ENC_us03_n624, _AES_ENC_us03_n623, _AES_ENC_us03_n622, _AES_ENC_us03_n621, _AES_ENC_us03_n620, _AES_ENC_us03_n619, _AES_ENC_us03_n618, _AES_ENC_us03_n617, _AES_ENC_us03_n616, _AES_ENC_us03_n615, _AES_ENC_us03_n614, _AES_ENC_us03_n613, _AES_ENC_us03_n612, _AES_ENC_us03_n611, _AES_ENC_us03_n610, _AES_ENC_us03_n609, _AES_ENC_us03_n608, _AES_ENC_us03_n607, _AES_ENC_us03_n606, _AES_ENC_us03_n605, 
  _AES_ENC_us03_n604, _AES_ENC_us03_n603, _AES_ENC_us03_n602, _AES_ENC_us03_n601, _AES_ENC_us03_n600, _AES_ENC_us03_n599, _AES_ENC_us03_n598, _AES_ENC_us03_n597, _AES_ENC_us03_n596, _AES_ENC_us03_n595, _AES_ENC_us03_n594, _AES_ENC_us03_n593, _AES_ENC_us03_n592, _AES_ENC_us03_n591, _AES_ENC_us03_n590, _AES_ENC_us03_n589, _AES_ENC_us03_n588, _AES_ENC_us03_n587, _AES_ENC_us03_n586, _AES_ENC_us03_n585, _AES_ENC_us03_n584, _AES_ENC_us03_n583, _AES_ENC_us03_n582, _AES_ENC_us03_n581, _AES_ENC_us03_n580, _AES_ENC_us03_n579, _AES_ENC_us03_n578, _AES_ENC_us03_n577, _AES_ENC_us03_n576, _AES_ENC_us03_n575, _AES_ENC_us03_n574, _AES_ENC_us03_n573, _AES_ENC_us03_n572, _AES_ENC_us03_n571, _AES_ENC_us03_n570, _AES_ENC_us03_n569, _AES_ENC_us10_n1135, _AES_ENC_us10_n1134, _AES_ENC_us10_n1133, _AES_ENC_us10_n1132, _AES_ENC_us10_n1131, _AES_ENC_us10_n1130, _AES_ENC_us10_n1129, _AES_ENC_us10_n1128, _AES_ENC_us10_n1127, _AES_ENC_us10_n1126, _AES_ENC_us10_n1125, _AES_ENC_us10_n1124, _AES_ENC_us10_n1123, _AES_ENC_us10_n1122, 
  _AES_ENC_us10_n1121, _AES_ENC_us10_n1120, _AES_ENC_us10_n1119, _AES_ENC_us10_n1118, _AES_ENC_us10_n1117, _AES_ENC_us10_n1116, _AES_ENC_us10_n1115, _AES_ENC_us10_n1114, _AES_ENC_us10_n1113, _AES_ENC_us10_n1112, _AES_ENC_us10_n1111, _AES_ENC_us10_n1110, _AES_ENC_us10_n1109, _AES_ENC_us10_n1108, _AES_ENC_us10_n1107, _AES_ENC_us10_n1106, _AES_ENC_us10_n1105, _AES_ENC_us10_n1104, _AES_ENC_us10_n1103, _AES_ENC_us10_n1102, _AES_ENC_us10_n1101, _AES_ENC_us10_n1100, _AES_ENC_us10_n1099, _AES_ENC_us10_n1098, _AES_ENC_us10_n1097, _AES_ENC_us10_n1096, _AES_ENC_us10_n1095, _AES_ENC_us10_n1094, _AES_ENC_us10_n1093, _AES_ENC_us10_n1092, _AES_ENC_us10_n1091, _AES_ENC_us10_n1090, _AES_ENC_us10_n1089, _AES_ENC_us10_n1088, _AES_ENC_us10_n1087, _AES_ENC_us10_n1086, _AES_ENC_us10_n1085, _AES_ENC_us10_n1084, _AES_ENC_us10_n1083, _AES_ENC_us10_n1082, _AES_ENC_us10_n1081, _AES_ENC_us10_n1080, _AES_ENC_us10_n1079, _AES_ENC_us10_n1078, _AES_ENC_us10_n1077, _AES_ENC_us10_n1076, _AES_ENC_us10_n1075, _AES_ENC_us10_n1074, _AES_ENC_us10_n1073, _AES_ENC_us10_n1072, 
  _AES_ENC_us10_n1071, _AES_ENC_us10_n1070, _AES_ENC_us10_n1069, _AES_ENC_us10_n1068, _AES_ENC_us10_n1067, _AES_ENC_us10_n1066, _AES_ENC_us10_n1065, _AES_ENC_us10_n1064, _AES_ENC_us10_n1063, _AES_ENC_us10_n1062, _AES_ENC_us10_n1061, _AES_ENC_us10_n1060, _AES_ENC_us10_n1059, _AES_ENC_us10_n1058, _AES_ENC_us10_n1057, _AES_ENC_us10_n1056, _AES_ENC_us10_n1055, _AES_ENC_us10_n1054, _AES_ENC_us10_n1053, _AES_ENC_us10_n1052, _AES_ENC_us10_n1051, _AES_ENC_us10_n1050, _AES_ENC_us10_n1049, _AES_ENC_us10_n1048, _AES_ENC_us10_n1047, _AES_ENC_us10_n1046, _AES_ENC_us10_n1045, _AES_ENC_us10_n1044, _AES_ENC_us10_n1043, _AES_ENC_us10_n1042, _AES_ENC_us10_n1041, _AES_ENC_us10_n1040, _AES_ENC_us10_n1039, _AES_ENC_us10_n1038, _AES_ENC_us10_n1037, _AES_ENC_us10_n1036, _AES_ENC_us10_n1035, _AES_ENC_us10_n1034, _AES_ENC_us10_n1033, _AES_ENC_us10_n1032, _AES_ENC_us10_n1031, _AES_ENC_us10_n1030, _AES_ENC_us10_n1029, _AES_ENC_us10_n1028, _AES_ENC_us10_n1027, _AES_ENC_us10_n1026, _AES_ENC_us10_n1025, _AES_ENC_us10_n1024, _AES_ENC_us10_n1023, _AES_ENC_us10_n1022, 
  _AES_ENC_us10_n1021, _AES_ENC_us10_n1020, _AES_ENC_us10_n1019, _AES_ENC_us10_n1018, _AES_ENC_us10_n1017, _AES_ENC_us10_n1016, _AES_ENC_us10_n1015, _AES_ENC_us10_n1014, _AES_ENC_us10_n1013, _AES_ENC_us10_n1012, _AES_ENC_us10_n1011, _AES_ENC_us10_n1010, _AES_ENC_us10_n1009, _AES_ENC_us10_n1008, _AES_ENC_us10_n1007, _AES_ENC_us10_n1006, _AES_ENC_us10_n1005, _AES_ENC_us10_n1004, _AES_ENC_us10_n1003, _AES_ENC_us10_n1002, _AES_ENC_us10_n1001, _AES_ENC_us10_n1000, _AES_ENC_us10_n999, _AES_ENC_us10_n998, _AES_ENC_us10_n997, _AES_ENC_us10_n996, _AES_ENC_us10_n995, _AES_ENC_us10_n994, _AES_ENC_us10_n993, _AES_ENC_us10_n992, _AES_ENC_us10_n991, _AES_ENC_us10_n990, _AES_ENC_us10_n989, _AES_ENC_us10_n988, _AES_ENC_us10_n987, _AES_ENC_us10_n986, _AES_ENC_us10_n985, _AES_ENC_us10_n984, _AES_ENC_us10_n983, _AES_ENC_us10_n982, _AES_ENC_us10_n981, _AES_ENC_us10_n980, _AES_ENC_us10_n979, _AES_ENC_us10_n978, _AES_ENC_us10_n977, _AES_ENC_us10_n976, _AES_ENC_us10_n975, _AES_ENC_us10_n974, _AES_ENC_us10_n973, _AES_ENC_us10_n972, 
  _AES_ENC_us10_n971, _AES_ENC_us10_n970, _AES_ENC_us10_n969, _AES_ENC_us10_n968, _AES_ENC_us10_n967, _AES_ENC_us10_n966, _AES_ENC_us10_n965, _AES_ENC_us10_n964, _AES_ENC_us10_n963, _AES_ENC_us10_n962, _AES_ENC_us10_n961, _AES_ENC_us10_n960, _AES_ENC_us10_n959, _AES_ENC_us10_n958, _AES_ENC_us10_n957, _AES_ENC_us10_n956, _AES_ENC_us10_n955, _AES_ENC_us10_n954, _AES_ENC_us10_n953, _AES_ENC_us10_n952, _AES_ENC_us10_n951, _AES_ENC_us10_n950, _AES_ENC_us10_n949, _AES_ENC_us10_n948, _AES_ENC_us10_n947, _AES_ENC_us10_n946, _AES_ENC_us10_n945, _AES_ENC_us10_n944, _AES_ENC_us10_n943, _AES_ENC_us10_n942, _AES_ENC_us10_n941, _AES_ENC_us10_n940, _AES_ENC_us10_n939, _AES_ENC_us10_n938, _AES_ENC_us10_n937, _AES_ENC_us10_n936, _AES_ENC_us10_n935, _AES_ENC_us10_n934, _AES_ENC_us10_n933, _AES_ENC_us10_n932, _AES_ENC_us10_n931, _AES_ENC_us10_n930, _AES_ENC_us10_n929, _AES_ENC_us10_n928, _AES_ENC_us10_n927, _AES_ENC_us10_n926, _AES_ENC_us10_n925, _AES_ENC_us10_n924, _AES_ENC_us10_n923, _AES_ENC_us10_n922, 
  _AES_ENC_us10_n921, _AES_ENC_us10_n920, _AES_ENC_us10_n919, _AES_ENC_us10_n918, _AES_ENC_us10_n917, _AES_ENC_us10_n916, _AES_ENC_us10_n915, _AES_ENC_us10_n914, _AES_ENC_us10_n913, _AES_ENC_us10_n912, _AES_ENC_us10_n911, _AES_ENC_us10_n910, _AES_ENC_us10_n909, _AES_ENC_us10_n908, _AES_ENC_us10_n907, _AES_ENC_us10_n906, _AES_ENC_us10_n905, _AES_ENC_us10_n904, _AES_ENC_us10_n903, _AES_ENC_us10_n902, _AES_ENC_us10_n901, _AES_ENC_us10_n900, _AES_ENC_us10_n899, _AES_ENC_us10_n898, _AES_ENC_us10_n897, _AES_ENC_us10_n896, _AES_ENC_us10_n895, _AES_ENC_us10_n894, _AES_ENC_us10_n893, _AES_ENC_us10_n892, _AES_ENC_us10_n891, _AES_ENC_us10_n890, _AES_ENC_us10_n889, _AES_ENC_us10_n888, _AES_ENC_us10_n887, _AES_ENC_us10_n886, _AES_ENC_us10_n885, _AES_ENC_us10_n884, _AES_ENC_us10_n883, _AES_ENC_us10_n882, _AES_ENC_us10_n881, _AES_ENC_us10_n880, _AES_ENC_us10_n879, _AES_ENC_us10_n878, _AES_ENC_us10_n877, _AES_ENC_us10_n876, _AES_ENC_us10_n875, _AES_ENC_us10_n874, _AES_ENC_us10_n873, _AES_ENC_us10_n872, 
  _AES_ENC_us10_n871, _AES_ENC_us10_n870, _AES_ENC_us10_n869, _AES_ENC_us10_n868, _AES_ENC_us10_n867, _AES_ENC_us10_n866, _AES_ENC_us10_n865, _AES_ENC_us10_n864, _AES_ENC_us10_n863, _AES_ENC_us10_n862, _AES_ENC_us10_n861, _AES_ENC_us10_n860, _AES_ENC_us10_n859, _AES_ENC_us10_n858, _AES_ENC_us10_n857, _AES_ENC_us10_n856, _AES_ENC_us10_n855, _AES_ENC_us10_n854, _AES_ENC_us10_n853, _AES_ENC_us10_n852, _AES_ENC_us10_n851, _AES_ENC_us10_n850, _AES_ENC_us10_n849, _AES_ENC_us10_n848, _AES_ENC_us10_n847, _AES_ENC_us10_n846, _AES_ENC_us10_n845, _AES_ENC_us10_n844, _AES_ENC_us10_n843, _AES_ENC_us10_n842, _AES_ENC_us10_n841, _AES_ENC_us10_n840, _AES_ENC_us10_n839, _AES_ENC_us10_n838, _AES_ENC_us10_n837, _AES_ENC_us10_n836, _AES_ENC_us10_n835, _AES_ENC_us10_n834, _AES_ENC_us10_n833, _AES_ENC_us10_n832, _AES_ENC_us10_n831, _AES_ENC_us10_n830, _AES_ENC_us10_n829, _AES_ENC_us10_n828, _AES_ENC_us10_n827, _AES_ENC_us10_n826, _AES_ENC_us10_n825, _AES_ENC_us10_n824, _AES_ENC_us10_n823, _AES_ENC_us10_n822, 
  _AES_ENC_us10_n821, _AES_ENC_us10_n820, _AES_ENC_us10_n819, _AES_ENC_us10_n818, _AES_ENC_us10_n817, _AES_ENC_us10_n816, _AES_ENC_us10_n815, _AES_ENC_us10_n814, _AES_ENC_us10_n813, _AES_ENC_us10_n812, _AES_ENC_us10_n811, _AES_ENC_us10_n810, _AES_ENC_us10_n809, _AES_ENC_us10_n808, _AES_ENC_us10_n807, _AES_ENC_us10_n806, _AES_ENC_us10_n805, _AES_ENC_us10_n804, _AES_ENC_us10_n803, _AES_ENC_us10_n802, _AES_ENC_us10_n801, _AES_ENC_us10_n800, _AES_ENC_us10_n799, _AES_ENC_us10_n798, _AES_ENC_us10_n797, _AES_ENC_us10_n796, _AES_ENC_us10_n795, _AES_ENC_us10_n794, _AES_ENC_us10_n793, _AES_ENC_us10_n792, _AES_ENC_us10_n791, _AES_ENC_us10_n790, _AES_ENC_us10_n789, _AES_ENC_us10_n788, _AES_ENC_us10_n787, _AES_ENC_us10_n786, _AES_ENC_us10_n785, _AES_ENC_us10_n784, _AES_ENC_us10_n783, _AES_ENC_us10_n782, _AES_ENC_us10_n781, _AES_ENC_us10_n780, _AES_ENC_us10_n779, _AES_ENC_us10_n778, _AES_ENC_us10_n777, _AES_ENC_us10_n776, _AES_ENC_us10_n775, _AES_ENC_us10_n774, _AES_ENC_us10_n773, _AES_ENC_us10_n772, 
  _AES_ENC_us10_n771, _AES_ENC_us10_n770, _AES_ENC_us10_n769, _AES_ENC_us10_n768, _AES_ENC_us10_n767, _AES_ENC_us10_n766, _AES_ENC_us10_n765, _AES_ENC_us10_n764, _AES_ENC_us10_n763, _AES_ENC_us10_n762, _AES_ENC_us10_n761, _AES_ENC_us10_n760, _AES_ENC_us10_n759, _AES_ENC_us10_n758, _AES_ENC_us10_n757, _AES_ENC_us10_n756, _AES_ENC_us10_n755, _AES_ENC_us10_n754, _AES_ENC_us10_n753, _AES_ENC_us10_n752, _AES_ENC_us10_n751, _AES_ENC_us10_n750, _AES_ENC_us10_n749, _AES_ENC_us10_n748, _AES_ENC_us10_n747, _AES_ENC_us10_n746, _AES_ENC_us10_n745, _AES_ENC_us10_n744, _AES_ENC_us10_n743, _AES_ENC_us10_n742, _AES_ENC_us10_n741, _AES_ENC_us10_n740, _AES_ENC_us10_n739, _AES_ENC_us10_n738, _AES_ENC_us10_n737, _AES_ENC_us10_n736, _AES_ENC_us10_n735, _AES_ENC_us10_n734, _AES_ENC_us10_n733, _AES_ENC_us10_n732, _AES_ENC_us10_n731, _AES_ENC_us10_n730, _AES_ENC_us10_n729, _AES_ENC_us10_n728, _AES_ENC_us10_n727, _AES_ENC_us10_n726, _AES_ENC_us10_n725, _AES_ENC_us10_n724, _AES_ENC_us10_n723, _AES_ENC_us10_n722, 
  _AES_ENC_us10_n721, _AES_ENC_us10_n720, _AES_ENC_us10_n719, _AES_ENC_us10_n718, _AES_ENC_us10_n717, _AES_ENC_us10_n716, _AES_ENC_us10_n715, _AES_ENC_us10_n714, _AES_ENC_us10_n713, _AES_ENC_us10_n712, _AES_ENC_us10_n711, _AES_ENC_us10_n710, _AES_ENC_us10_n709, _AES_ENC_us10_n708, _AES_ENC_us10_n707, _AES_ENC_us10_n706, _AES_ENC_us10_n705, _AES_ENC_us10_n704, _AES_ENC_us10_n703, _AES_ENC_us10_n702, _AES_ENC_us10_n701, _AES_ENC_us10_n700, _AES_ENC_us10_n699, _AES_ENC_us10_n698, _AES_ENC_us10_n697, _AES_ENC_us10_n696, _AES_ENC_us10_n695, _AES_ENC_us10_n694, _AES_ENC_us10_n693, _AES_ENC_us10_n692, _AES_ENC_us10_n691, _AES_ENC_us10_n690, _AES_ENC_us10_n689, _AES_ENC_us10_n688, _AES_ENC_us10_n687, _AES_ENC_us10_n686, _AES_ENC_us10_n685, _AES_ENC_us10_n684, _AES_ENC_us10_n683, _AES_ENC_us10_n682, _AES_ENC_us10_n681, _AES_ENC_us10_n680, _AES_ENC_us10_n679, _AES_ENC_us10_n678, _AES_ENC_us10_n677, _AES_ENC_us10_n676, _AES_ENC_us10_n675, _AES_ENC_us10_n674, _AES_ENC_us10_n673, _AES_ENC_us10_n672, 
  _AES_ENC_us10_n671, _AES_ENC_us10_n670, _AES_ENC_us10_n669, _AES_ENC_us10_n668, _AES_ENC_us10_n667, _AES_ENC_us10_n666, _AES_ENC_us10_n665, _AES_ENC_us10_n664, _AES_ENC_us10_n663, _AES_ENC_us10_n662, _AES_ENC_us10_n661, _AES_ENC_us10_n660, _AES_ENC_us10_n659, _AES_ENC_us10_n658, _AES_ENC_us10_n657, _AES_ENC_us10_n656, _AES_ENC_us10_n655, _AES_ENC_us10_n654, _AES_ENC_us10_n653, _AES_ENC_us10_n652, _AES_ENC_us10_n651, _AES_ENC_us10_n650, _AES_ENC_us10_n649, _AES_ENC_us10_n648, _AES_ENC_us10_n647, _AES_ENC_us10_n646, _AES_ENC_us10_n645, _AES_ENC_us10_n644, _AES_ENC_us10_n643, _AES_ENC_us10_n642, _AES_ENC_us10_n641, _AES_ENC_us10_n640, _AES_ENC_us10_n639, _AES_ENC_us10_n638, _AES_ENC_us10_n637, _AES_ENC_us10_n636, _AES_ENC_us10_n635, _AES_ENC_us10_n634, _AES_ENC_us10_n633, _AES_ENC_us10_n632, _AES_ENC_us10_n631, _AES_ENC_us10_n630, _AES_ENC_us10_n629, _AES_ENC_us10_n628, _AES_ENC_us10_n627, _AES_ENC_us10_n626, _AES_ENC_us10_n625, _AES_ENC_us10_n624, _AES_ENC_us10_n623, _AES_ENC_us10_n622, 
  _AES_ENC_us10_n621, _AES_ENC_us10_n620, _AES_ENC_us10_n619, _AES_ENC_us10_n618, _AES_ENC_us10_n617, _AES_ENC_us10_n616, _AES_ENC_us10_n615, _AES_ENC_us10_n614, _AES_ENC_us10_n613, _AES_ENC_us10_n612, _AES_ENC_us10_n611, _AES_ENC_us10_n610, _AES_ENC_us10_n609, _AES_ENC_us10_n608, _AES_ENC_us10_n607, _AES_ENC_us10_n606, _AES_ENC_us10_n605, _AES_ENC_us10_n604, _AES_ENC_us10_n603, _AES_ENC_us10_n602, _AES_ENC_us10_n601, _AES_ENC_us10_n600, _AES_ENC_us10_n599, _AES_ENC_us10_n598, _AES_ENC_us10_n597, _AES_ENC_us10_n596, _AES_ENC_us10_n595, _AES_ENC_us10_n594, _AES_ENC_us10_n593, _AES_ENC_us10_n592, _AES_ENC_us10_n591, _AES_ENC_us10_n590, _AES_ENC_us10_n589, _AES_ENC_us10_n588, _AES_ENC_us10_n587, _AES_ENC_us10_n586, _AES_ENC_us10_n585, _AES_ENC_us10_n584, _AES_ENC_us10_n583, _AES_ENC_us10_n582, _AES_ENC_us10_n581, _AES_ENC_us10_n580, _AES_ENC_us10_n579, _AES_ENC_us10_n578, _AES_ENC_us10_n577, _AES_ENC_us10_n576, _AES_ENC_us10_n575, _AES_ENC_us10_n574, _AES_ENC_us10_n573, _AES_ENC_us10_n572, 
  _AES_ENC_us10_n571, _AES_ENC_us10_n570, _AES_ENC_us10_n569, _AES_ENC_us11_n1135, _AES_ENC_us11_n1134, _AES_ENC_us11_n1133, _AES_ENC_us11_n1132, _AES_ENC_us11_n1131, _AES_ENC_us11_n1130, _AES_ENC_us11_n1129, _AES_ENC_us11_n1128, _AES_ENC_us11_n1127, _AES_ENC_us11_n1126, _AES_ENC_us11_n1125, _AES_ENC_us11_n1124, _AES_ENC_us11_n1123, _AES_ENC_us11_n1122, _AES_ENC_us11_n1121, _AES_ENC_us11_n1120, _AES_ENC_us11_n1119, _AES_ENC_us11_n1118, _AES_ENC_us11_n1117, _AES_ENC_us11_n1116, _AES_ENC_us11_n1115, _AES_ENC_us11_n1114, _AES_ENC_us11_n1113, _AES_ENC_us11_n1112, _AES_ENC_us11_n1111, _AES_ENC_us11_n1110, _AES_ENC_us11_n1109, _AES_ENC_us11_n1108, _AES_ENC_us11_n1107, _AES_ENC_us11_n1106, _AES_ENC_us11_n1105, _AES_ENC_us11_n1104, _AES_ENC_us11_n1103, _AES_ENC_us11_n1102, _AES_ENC_us11_n1101, _AES_ENC_us11_n1100, _AES_ENC_us11_n1099, _AES_ENC_us11_n1098, _AES_ENC_us11_n1097, _AES_ENC_us11_n1096, _AES_ENC_us11_n1095, _AES_ENC_us11_n1094, _AES_ENC_us11_n1093, _AES_ENC_us11_n1092, _AES_ENC_us11_n1091, _AES_ENC_us11_n1090, _AES_ENC_us11_n1089, 
  _AES_ENC_us11_n1088, _AES_ENC_us11_n1087, _AES_ENC_us11_n1086, _AES_ENC_us11_n1085, _AES_ENC_us11_n1084, _AES_ENC_us11_n1083, _AES_ENC_us11_n1082, _AES_ENC_us11_n1081, _AES_ENC_us11_n1080, _AES_ENC_us11_n1079, _AES_ENC_us11_n1078, _AES_ENC_us11_n1077, _AES_ENC_us11_n1076, _AES_ENC_us11_n1075, _AES_ENC_us11_n1074, _AES_ENC_us11_n1073, _AES_ENC_us11_n1072, _AES_ENC_us11_n1071, _AES_ENC_us11_n1070, _AES_ENC_us11_n1069, _AES_ENC_us11_n1068, _AES_ENC_us11_n1067, _AES_ENC_us11_n1066, _AES_ENC_us11_n1065, _AES_ENC_us11_n1064, _AES_ENC_us11_n1063, _AES_ENC_us11_n1062, _AES_ENC_us11_n1061, _AES_ENC_us11_n1060, _AES_ENC_us11_n1059, _AES_ENC_us11_n1058, _AES_ENC_us11_n1057, _AES_ENC_us11_n1056, _AES_ENC_us11_n1055, _AES_ENC_us11_n1054, _AES_ENC_us11_n1053, _AES_ENC_us11_n1052, _AES_ENC_us11_n1051, _AES_ENC_us11_n1050, _AES_ENC_us11_n1049, _AES_ENC_us11_n1048, _AES_ENC_us11_n1047, _AES_ENC_us11_n1046, _AES_ENC_us11_n1045, _AES_ENC_us11_n1044, _AES_ENC_us11_n1043, _AES_ENC_us11_n1042, _AES_ENC_us11_n1041, _AES_ENC_us11_n1040, _AES_ENC_us11_n1039, 
  _AES_ENC_us11_n1038, _AES_ENC_us11_n1037, _AES_ENC_us11_n1036, _AES_ENC_us11_n1035, _AES_ENC_us11_n1034, _AES_ENC_us11_n1033, _AES_ENC_us11_n1032, _AES_ENC_us11_n1031, _AES_ENC_us11_n1030, _AES_ENC_us11_n1029, _AES_ENC_us11_n1028, _AES_ENC_us11_n1027, _AES_ENC_us11_n1026, _AES_ENC_us11_n1025, _AES_ENC_us11_n1024, _AES_ENC_us11_n1023, _AES_ENC_us11_n1022, _AES_ENC_us11_n1021, _AES_ENC_us11_n1020, _AES_ENC_us11_n1019, _AES_ENC_us11_n1018, _AES_ENC_us11_n1017, _AES_ENC_us11_n1016, _AES_ENC_us11_n1015, _AES_ENC_us11_n1014, _AES_ENC_us11_n1013, _AES_ENC_us11_n1012, _AES_ENC_us11_n1011, _AES_ENC_us11_n1010, _AES_ENC_us11_n1009, _AES_ENC_us11_n1008, _AES_ENC_us11_n1007, _AES_ENC_us11_n1006, _AES_ENC_us11_n1005, _AES_ENC_us11_n1004, _AES_ENC_us11_n1003, _AES_ENC_us11_n1002, _AES_ENC_us11_n1001, _AES_ENC_us11_n1000, _AES_ENC_us11_n999, _AES_ENC_us11_n998, _AES_ENC_us11_n997, _AES_ENC_us11_n996, _AES_ENC_us11_n995, _AES_ENC_us11_n994, _AES_ENC_us11_n993, _AES_ENC_us11_n992, _AES_ENC_us11_n991, _AES_ENC_us11_n990, _AES_ENC_us11_n989, 
  _AES_ENC_us11_n988, _AES_ENC_us11_n987, _AES_ENC_us11_n986, _AES_ENC_us11_n985, _AES_ENC_us11_n984, _AES_ENC_us11_n983, _AES_ENC_us11_n982, _AES_ENC_us11_n981, _AES_ENC_us11_n980, _AES_ENC_us11_n979, _AES_ENC_us11_n978, _AES_ENC_us11_n977, _AES_ENC_us11_n976, _AES_ENC_us11_n975, _AES_ENC_us11_n974, _AES_ENC_us11_n973, _AES_ENC_us11_n972, _AES_ENC_us11_n971, _AES_ENC_us11_n970, _AES_ENC_us11_n969, _AES_ENC_us11_n968, _AES_ENC_us11_n967, _AES_ENC_us11_n966, _AES_ENC_us11_n965, _AES_ENC_us11_n964, _AES_ENC_us11_n963, _AES_ENC_us11_n962, _AES_ENC_us11_n961, _AES_ENC_us11_n960, _AES_ENC_us11_n959, _AES_ENC_us11_n958, _AES_ENC_us11_n957, _AES_ENC_us11_n956, _AES_ENC_us11_n955, _AES_ENC_us11_n954, _AES_ENC_us11_n953, _AES_ENC_us11_n952, _AES_ENC_us11_n951, _AES_ENC_us11_n950, _AES_ENC_us11_n949, _AES_ENC_us11_n948, _AES_ENC_us11_n947, _AES_ENC_us11_n946, _AES_ENC_us11_n945, _AES_ENC_us11_n944, _AES_ENC_us11_n943, _AES_ENC_us11_n942, _AES_ENC_us11_n941, _AES_ENC_us11_n940, _AES_ENC_us11_n939, 
  _AES_ENC_us11_n938, _AES_ENC_us11_n937, _AES_ENC_us11_n936, _AES_ENC_us11_n935, _AES_ENC_us11_n934, _AES_ENC_us11_n933, _AES_ENC_us11_n932, _AES_ENC_us11_n931, _AES_ENC_us11_n930, _AES_ENC_us11_n929, _AES_ENC_us11_n928, _AES_ENC_us11_n927, _AES_ENC_us11_n926, _AES_ENC_us11_n925, _AES_ENC_us11_n924, _AES_ENC_us11_n923, _AES_ENC_us11_n922, _AES_ENC_us11_n921, _AES_ENC_us11_n920, _AES_ENC_us11_n919, _AES_ENC_us11_n918, _AES_ENC_us11_n917, _AES_ENC_us11_n916, _AES_ENC_us11_n915, _AES_ENC_us11_n914, _AES_ENC_us11_n913, _AES_ENC_us11_n912, _AES_ENC_us11_n911, _AES_ENC_us11_n910, _AES_ENC_us11_n909, _AES_ENC_us11_n908, _AES_ENC_us11_n907, _AES_ENC_us11_n906, _AES_ENC_us11_n905, _AES_ENC_us11_n904, _AES_ENC_us11_n903, _AES_ENC_us11_n902, _AES_ENC_us11_n901, _AES_ENC_us11_n900, _AES_ENC_us11_n899, _AES_ENC_us11_n898, _AES_ENC_us11_n897, _AES_ENC_us11_n896, _AES_ENC_us11_n895, _AES_ENC_us11_n894, _AES_ENC_us11_n893, _AES_ENC_us11_n892, _AES_ENC_us11_n891, _AES_ENC_us11_n890, _AES_ENC_us11_n889, 
  _AES_ENC_us11_n888, _AES_ENC_us11_n887, _AES_ENC_us11_n886, _AES_ENC_us11_n885, _AES_ENC_us11_n884, _AES_ENC_us11_n883, _AES_ENC_us11_n882, _AES_ENC_us11_n881, _AES_ENC_us11_n880, _AES_ENC_us11_n879, _AES_ENC_us11_n878, _AES_ENC_us11_n877, _AES_ENC_us11_n876, _AES_ENC_us11_n875, _AES_ENC_us11_n874, _AES_ENC_us11_n873, _AES_ENC_us11_n872, _AES_ENC_us11_n871, _AES_ENC_us11_n870, _AES_ENC_us11_n869, _AES_ENC_us11_n868, _AES_ENC_us11_n867, _AES_ENC_us11_n866, _AES_ENC_us11_n865, _AES_ENC_us11_n864, _AES_ENC_us11_n863, _AES_ENC_us11_n862, _AES_ENC_us11_n861, _AES_ENC_us11_n860, _AES_ENC_us11_n859, _AES_ENC_us11_n858, _AES_ENC_us11_n857, _AES_ENC_us11_n856, _AES_ENC_us11_n855, _AES_ENC_us11_n854, _AES_ENC_us11_n853, _AES_ENC_us11_n852, _AES_ENC_us11_n851, _AES_ENC_us11_n850, _AES_ENC_us11_n849, _AES_ENC_us11_n848, _AES_ENC_us11_n847, _AES_ENC_us11_n846, _AES_ENC_us11_n845, _AES_ENC_us11_n844, _AES_ENC_us11_n843, _AES_ENC_us11_n842, _AES_ENC_us11_n841, _AES_ENC_us11_n840, _AES_ENC_us11_n839, 
  _AES_ENC_us11_n838, _AES_ENC_us11_n837, _AES_ENC_us11_n836, _AES_ENC_us11_n835, _AES_ENC_us11_n834, _AES_ENC_us11_n833, _AES_ENC_us11_n832, _AES_ENC_us11_n831, _AES_ENC_us11_n830, _AES_ENC_us11_n829, _AES_ENC_us11_n828, _AES_ENC_us11_n827, _AES_ENC_us11_n826, _AES_ENC_us11_n825, _AES_ENC_us11_n824, _AES_ENC_us11_n823, _AES_ENC_us11_n822, _AES_ENC_us11_n821, _AES_ENC_us11_n820, _AES_ENC_us11_n819, _AES_ENC_us11_n818, _AES_ENC_us11_n817, _AES_ENC_us11_n816, _AES_ENC_us11_n815, _AES_ENC_us11_n814, _AES_ENC_us11_n813, _AES_ENC_us11_n812, _AES_ENC_us11_n811, _AES_ENC_us11_n810, _AES_ENC_us11_n809, _AES_ENC_us11_n808, _AES_ENC_us11_n807, _AES_ENC_us11_n806, _AES_ENC_us11_n805, _AES_ENC_us11_n804, _AES_ENC_us11_n803, _AES_ENC_us11_n802, _AES_ENC_us11_n801, _AES_ENC_us11_n800, _AES_ENC_us11_n799, _AES_ENC_us11_n798, _AES_ENC_us11_n797, _AES_ENC_us11_n796, _AES_ENC_us11_n795, _AES_ENC_us11_n794, _AES_ENC_us11_n793, _AES_ENC_us11_n792, _AES_ENC_us11_n791, _AES_ENC_us11_n790, _AES_ENC_us11_n789, 
  _AES_ENC_us11_n788, _AES_ENC_us11_n787, _AES_ENC_us11_n786, _AES_ENC_us11_n785, _AES_ENC_us11_n784, _AES_ENC_us11_n783, _AES_ENC_us11_n782, _AES_ENC_us11_n781, _AES_ENC_us11_n780, _AES_ENC_us11_n779, _AES_ENC_us11_n778, _AES_ENC_us11_n777, _AES_ENC_us11_n776, _AES_ENC_us11_n775, _AES_ENC_us11_n774, _AES_ENC_us11_n773, _AES_ENC_us11_n772, _AES_ENC_us11_n771, _AES_ENC_us11_n770, _AES_ENC_us11_n769, _AES_ENC_us11_n768, _AES_ENC_us11_n767, _AES_ENC_us11_n766, _AES_ENC_us11_n765, _AES_ENC_us11_n764, _AES_ENC_us11_n763, _AES_ENC_us11_n762, _AES_ENC_us11_n761, _AES_ENC_us11_n760, _AES_ENC_us11_n759, _AES_ENC_us11_n758, _AES_ENC_us11_n757, _AES_ENC_us11_n756, _AES_ENC_us11_n755, _AES_ENC_us11_n754, _AES_ENC_us11_n753, _AES_ENC_us11_n752, _AES_ENC_us11_n751, _AES_ENC_us11_n750, _AES_ENC_us11_n749, _AES_ENC_us11_n748, _AES_ENC_us11_n747, _AES_ENC_us11_n746, _AES_ENC_us11_n745, _AES_ENC_us11_n744, _AES_ENC_us11_n743, _AES_ENC_us11_n742, _AES_ENC_us11_n741, _AES_ENC_us11_n740, _AES_ENC_us11_n739, 
  _AES_ENC_us11_n738, _AES_ENC_us11_n737, _AES_ENC_us11_n736, _AES_ENC_us11_n735, _AES_ENC_us11_n734, _AES_ENC_us11_n733, _AES_ENC_us11_n732, _AES_ENC_us11_n731, _AES_ENC_us11_n730, _AES_ENC_us11_n729, _AES_ENC_us11_n728, _AES_ENC_us11_n727, _AES_ENC_us11_n726, _AES_ENC_us11_n725, _AES_ENC_us11_n724, _AES_ENC_us11_n723, _AES_ENC_us11_n722, _AES_ENC_us11_n721, _AES_ENC_us11_n720, _AES_ENC_us11_n719, _AES_ENC_us11_n718, _AES_ENC_us11_n717, _AES_ENC_us11_n716, _AES_ENC_us11_n715, _AES_ENC_us11_n714, _AES_ENC_us11_n713, _AES_ENC_us11_n712, _AES_ENC_us11_n711, _AES_ENC_us11_n710, _AES_ENC_us11_n709, _AES_ENC_us11_n708, _AES_ENC_us11_n707, _AES_ENC_us11_n706, _AES_ENC_us11_n705, _AES_ENC_us11_n704, _AES_ENC_us11_n703, _AES_ENC_us11_n702, _AES_ENC_us11_n701, _AES_ENC_us11_n700, _AES_ENC_us11_n699, _AES_ENC_us11_n698, _AES_ENC_us11_n697, _AES_ENC_us11_n696, _AES_ENC_us11_n695, _AES_ENC_us11_n694, _AES_ENC_us11_n693, _AES_ENC_us11_n692, _AES_ENC_us11_n691, _AES_ENC_us11_n690, _AES_ENC_us11_n689, 
  _AES_ENC_us11_n688, _AES_ENC_us11_n687, _AES_ENC_us11_n686, _AES_ENC_us11_n685, _AES_ENC_us11_n684, _AES_ENC_us11_n683, _AES_ENC_us11_n682, _AES_ENC_us11_n681, _AES_ENC_us11_n680, _AES_ENC_us11_n679, _AES_ENC_us11_n678, _AES_ENC_us11_n677, _AES_ENC_us11_n676, _AES_ENC_us11_n675, _AES_ENC_us11_n674, _AES_ENC_us11_n673, _AES_ENC_us11_n672, _AES_ENC_us11_n671, _AES_ENC_us11_n670, _AES_ENC_us11_n669, _AES_ENC_us11_n668, _AES_ENC_us11_n667, _AES_ENC_us11_n666, _AES_ENC_us11_n665, _AES_ENC_us11_n664, _AES_ENC_us11_n663, _AES_ENC_us11_n662, _AES_ENC_us11_n661, _AES_ENC_us11_n660, _AES_ENC_us11_n659, _AES_ENC_us11_n658, _AES_ENC_us11_n657, _AES_ENC_us11_n656, _AES_ENC_us11_n655, _AES_ENC_us11_n654, _AES_ENC_us11_n653, _AES_ENC_us11_n652, _AES_ENC_us11_n651, _AES_ENC_us11_n650, _AES_ENC_us11_n649, _AES_ENC_us11_n648, _AES_ENC_us11_n647, _AES_ENC_us11_n646, _AES_ENC_us11_n645, _AES_ENC_us11_n644, _AES_ENC_us11_n643, _AES_ENC_us11_n642, _AES_ENC_us11_n641, _AES_ENC_us11_n640, _AES_ENC_us11_n639, 
  _AES_ENC_us11_n638, _AES_ENC_us11_n637, _AES_ENC_us11_n636, _AES_ENC_us11_n635, _AES_ENC_us11_n634, _AES_ENC_us11_n633, _AES_ENC_us11_n632, _AES_ENC_us11_n631, _AES_ENC_us11_n630, _AES_ENC_us11_n629, _AES_ENC_us11_n628, _AES_ENC_us11_n627, _AES_ENC_us11_n626, _AES_ENC_us11_n625, _AES_ENC_us11_n624, _AES_ENC_us11_n623, _AES_ENC_us11_n622, _AES_ENC_us11_n621, _AES_ENC_us11_n620, _AES_ENC_us11_n619, _AES_ENC_us11_n618, _AES_ENC_us11_n617, _AES_ENC_us11_n616, _AES_ENC_us11_n615, _AES_ENC_us11_n614, _AES_ENC_us11_n613, _AES_ENC_us11_n612, _AES_ENC_us11_n611, _AES_ENC_us11_n610, _AES_ENC_us11_n609, _AES_ENC_us11_n608, _AES_ENC_us11_n607, _AES_ENC_us11_n606, _AES_ENC_us11_n605, _AES_ENC_us11_n604, _AES_ENC_us11_n603, _AES_ENC_us11_n602, _AES_ENC_us11_n601, _AES_ENC_us11_n600, _AES_ENC_us11_n599, _AES_ENC_us11_n598, _AES_ENC_us11_n597, _AES_ENC_us11_n596, _AES_ENC_us11_n595, _AES_ENC_us11_n594, _AES_ENC_us11_n593, _AES_ENC_us11_n592, _AES_ENC_us11_n591, _AES_ENC_us11_n590, _AES_ENC_us11_n589, 
  _AES_ENC_us11_n588, _AES_ENC_us11_n587, _AES_ENC_us11_n586, _AES_ENC_us11_n585, _AES_ENC_us11_n584, _AES_ENC_us11_n583, _AES_ENC_us11_n582, _AES_ENC_us11_n581, _AES_ENC_us11_n580, _AES_ENC_us11_n579, _AES_ENC_us11_n578, _AES_ENC_us11_n577, _AES_ENC_us11_n576, _AES_ENC_us11_n575, _AES_ENC_us11_n574, _AES_ENC_us11_n573, _AES_ENC_us11_n572, _AES_ENC_us11_n571, _AES_ENC_us11_n570, _AES_ENC_us11_n569, _AES_ENC_us12_n1135, _AES_ENC_us12_n1134, _AES_ENC_us12_n1133, _AES_ENC_us12_n1132, _AES_ENC_us12_n1131, _AES_ENC_us12_n1130, _AES_ENC_us12_n1129, _AES_ENC_us12_n1128, _AES_ENC_us12_n1127, _AES_ENC_us12_n1126, _AES_ENC_us12_n1125, _AES_ENC_us12_n1124, _AES_ENC_us12_n1123, _AES_ENC_us12_n1122, _AES_ENC_us12_n1121, _AES_ENC_us12_n1120, _AES_ENC_us12_n1119, _AES_ENC_us12_n1118, _AES_ENC_us12_n1117, _AES_ENC_us12_n1116, _AES_ENC_us12_n1115, _AES_ENC_us12_n1114, _AES_ENC_us12_n1113, _AES_ENC_us12_n1112, _AES_ENC_us12_n1111, _AES_ENC_us12_n1110, _AES_ENC_us12_n1109, _AES_ENC_us12_n1108, _AES_ENC_us12_n1107, _AES_ENC_us12_n1106, 
  _AES_ENC_us12_n1105, _AES_ENC_us12_n1104, _AES_ENC_us12_n1103, _AES_ENC_us12_n1102, _AES_ENC_us12_n1101, _AES_ENC_us12_n1100, _AES_ENC_us12_n1099, _AES_ENC_us12_n1098, _AES_ENC_us12_n1097, _AES_ENC_us12_n1096, _AES_ENC_us12_n1095, _AES_ENC_us12_n1094, _AES_ENC_us12_n1093, _AES_ENC_us12_n1092, _AES_ENC_us12_n1091, _AES_ENC_us12_n1090, _AES_ENC_us12_n1089, _AES_ENC_us12_n1088, _AES_ENC_us12_n1087, _AES_ENC_us12_n1086, _AES_ENC_us12_n1085, _AES_ENC_us12_n1084, _AES_ENC_us12_n1083, _AES_ENC_us12_n1082, _AES_ENC_us12_n1081, _AES_ENC_us12_n1080, _AES_ENC_us12_n1079, _AES_ENC_us12_n1078, _AES_ENC_us12_n1077, _AES_ENC_us12_n1076, _AES_ENC_us12_n1075, _AES_ENC_us12_n1074, _AES_ENC_us12_n1073, _AES_ENC_us12_n1072, _AES_ENC_us12_n1071, _AES_ENC_us12_n1070, _AES_ENC_us12_n1069, _AES_ENC_us12_n1068, _AES_ENC_us12_n1067, _AES_ENC_us12_n1066, _AES_ENC_us12_n1065, _AES_ENC_us12_n1064, _AES_ENC_us12_n1063, _AES_ENC_us12_n1062, _AES_ENC_us12_n1061, _AES_ENC_us12_n1060, _AES_ENC_us12_n1059, _AES_ENC_us12_n1058, _AES_ENC_us12_n1057, _AES_ENC_us12_n1056, 
  _AES_ENC_us12_n1055, _AES_ENC_us12_n1054, _AES_ENC_us12_n1053, _AES_ENC_us12_n1052, _AES_ENC_us12_n1051, _AES_ENC_us12_n1050, _AES_ENC_us12_n1049, _AES_ENC_us12_n1048, _AES_ENC_us12_n1047, _AES_ENC_us12_n1046, _AES_ENC_us12_n1045, _AES_ENC_us12_n1044, _AES_ENC_us12_n1043, _AES_ENC_us12_n1042, _AES_ENC_us12_n1041, _AES_ENC_us12_n1040, _AES_ENC_us12_n1039, _AES_ENC_us12_n1038, _AES_ENC_us12_n1037, _AES_ENC_us12_n1036, _AES_ENC_us12_n1035, _AES_ENC_us12_n1034, _AES_ENC_us12_n1033, _AES_ENC_us12_n1032, _AES_ENC_us12_n1031, _AES_ENC_us12_n1030, _AES_ENC_us12_n1029, _AES_ENC_us12_n1028, _AES_ENC_us12_n1027, _AES_ENC_us12_n1026, _AES_ENC_us12_n1025, _AES_ENC_us12_n1024, _AES_ENC_us12_n1023, _AES_ENC_us12_n1022, _AES_ENC_us12_n1021, _AES_ENC_us12_n1020, _AES_ENC_us12_n1019, _AES_ENC_us12_n1018, _AES_ENC_us12_n1017, _AES_ENC_us12_n1016, _AES_ENC_us12_n1015, _AES_ENC_us12_n1014, _AES_ENC_us12_n1013, _AES_ENC_us12_n1012, _AES_ENC_us12_n1011, _AES_ENC_us12_n1010, _AES_ENC_us12_n1009, _AES_ENC_us12_n1008, _AES_ENC_us12_n1007, _AES_ENC_us12_n1006, 
  _AES_ENC_us12_n1005, _AES_ENC_us12_n1004, _AES_ENC_us12_n1003, _AES_ENC_us12_n1002, _AES_ENC_us12_n1001, _AES_ENC_us12_n1000, _AES_ENC_us12_n999, _AES_ENC_us12_n998, _AES_ENC_us12_n997, _AES_ENC_us12_n996, _AES_ENC_us12_n995, _AES_ENC_us12_n994, _AES_ENC_us12_n993, _AES_ENC_us12_n992, _AES_ENC_us12_n991, _AES_ENC_us12_n990, _AES_ENC_us12_n989, _AES_ENC_us12_n988, _AES_ENC_us12_n987, _AES_ENC_us12_n986, _AES_ENC_us12_n985, _AES_ENC_us12_n984, _AES_ENC_us12_n983, _AES_ENC_us12_n982, _AES_ENC_us12_n981, _AES_ENC_us12_n980, _AES_ENC_us12_n979, _AES_ENC_us12_n978, _AES_ENC_us12_n977, _AES_ENC_us12_n976, _AES_ENC_us12_n975, _AES_ENC_us12_n974, _AES_ENC_us12_n973, _AES_ENC_us12_n972, _AES_ENC_us12_n971, _AES_ENC_us12_n970, _AES_ENC_us12_n969, _AES_ENC_us12_n968, _AES_ENC_us12_n967, _AES_ENC_us12_n966, _AES_ENC_us12_n965, _AES_ENC_us12_n964, _AES_ENC_us12_n963, _AES_ENC_us12_n962, _AES_ENC_us12_n961, _AES_ENC_us12_n960, _AES_ENC_us12_n959, _AES_ENC_us12_n958, _AES_ENC_us12_n957, _AES_ENC_us12_n956, 
  _AES_ENC_us12_n955, _AES_ENC_us12_n954, _AES_ENC_us12_n953, _AES_ENC_us12_n952, _AES_ENC_us12_n951, _AES_ENC_us12_n950, _AES_ENC_us12_n949, _AES_ENC_us12_n948, _AES_ENC_us12_n947, _AES_ENC_us12_n946, _AES_ENC_us12_n945, _AES_ENC_us12_n944, _AES_ENC_us12_n943, _AES_ENC_us12_n942, _AES_ENC_us12_n941, _AES_ENC_us12_n940, _AES_ENC_us12_n939, _AES_ENC_us12_n938, _AES_ENC_us12_n937, _AES_ENC_us12_n936, _AES_ENC_us12_n935, _AES_ENC_us12_n934, _AES_ENC_us12_n933, _AES_ENC_us12_n932, _AES_ENC_us12_n931, _AES_ENC_us12_n930, _AES_ENC_us12_n929, _AES_ENC_us12_n928, _AES_ENC_us12_n927, _AES_ENC_us12_n926, _AES_ENC_us12_n925, _AES_ENC_us12_n924, _AES_ENC_us12_n923, _AES_ENC_us12_n922, _AES_ENC_us12_n921, _AES_ENC_us12_n920, _AES_ENC_us12_n919, _AES_ENC_us12_n918, _AES_ENC_us12_n917, _AES_ENC_us12_n916, _AES_ENC_us12_n915, _AES_ENC_us12_n914, _AES_ENC_us12_n913, _AES_ENC_us12_n912, _AES_ENC_us12_n911, _AES_ENC_us12_n910, _AES_ENC_us12_n909, _AES_ENC_us12_n908, _AES_ENC_us12_n907, _AES_ENC_us12_n906, 
  _AES_ENC_us12_n905, _AES_ENC_us12_n904, _AES_ENC_us12_n903, _AES_ENC_us12_n902, _AES_ENC_us12_n901, _AES_ENC_us12_n900, _AES_ENC_us12_n899, _AES_ENC_us12_n898, _AES_ENC_us12_n897, _AES_ENC_us12_n896, _AES_ENC_us12_n895, _AES_ENC_us12_n894, _AES_ENC_us12_n893, _AES_ENC_us12_n892, _AES_ENC_us12_n891, _AES_ENC_us12_n890, _AES_ENC_us12_n889, _AES_ENC_us12_n888, _AES_ENC_us12_n887, _AES_ENC_us12_n886, _AES_ENC_us12_n885, _AES_ENC_us12_n884, _AES_ENC_us12_n883, _AES_ENC_us12_n882, _AES_ENC_us12_n881, _AES_ENC_us12_n880, _AES_ENC_us12_n879, _AES_ENC_us12_n878, _AES_ENC_us12_n877, _AES_ENC_us12_n876, _AES_ENC_us12_n875, _AES_ENC_us12_n874, _AES_ENC_us12_n873, _AES_ENC_us12_n872, _AES_ENC_us12_n871, _AES_ENC_us12_n870, _AES_ENC_us12_n869, _AES_ENC_us12_n868, _AES_ENC_us12_n867, _AES_ENC_us12_n866, _AES_ENC_us12_n865, _AES_ENC_us12_n864, _AES_ENC_us12_n863, _AES_ENC_us12_n862, _AES_ENC_us12_n861, _AES_ENC_us12_n860, _AES_ENC_us12_n859, _AES_ENC_us12_n858, _AES_ENC_us12_n857, _AES_ENC_us12_n856, 
  _AES_ENC_us12_n855, _AES_ENC_us12_n854, _AES_ENC_us12_n853, _AES_ENC_us12_n852, _AES_ENC_us12_n851, _AES_ENC_us12_n850, _AES_ENC_us12_n849, _AES_ENC_us12_n848, _AES_ENC_us12_n847, _AES_ENC_us12_n846, _AES_ENC_us12_n845, _AES_ENC_us12_n844, _AES_ENC_us12_n843, _AES_ENC_us12_n842, _AES_ENC_us12_n841, _AES_ENC_us12_n840, _AES_ENC_us12_n839, _AES_ENC_us12_n838, _AES_ENC_us12_n837, _AES_ENC_us12_n836, _AES_ENC_us12_n835, _AES_ENC_us12_n834, _AES_ENC_us12_n833, _AES_ENC_us12_n832, _AES_ENC_us12_n831, _AES_ENC_us12_n830, _AES_ENC_us12_n829, _AES_ENC_us12_n828, _AES_ENC_us12_n827, _AES_ENC_us12_n826, _AES_ENC_us12_n825, _AES_ENC_us12_n824, _AES_ENC_us12_n823, _AES_ENC_us12_n822, _AES_ENC_us12_n821, _AES_ENC_us12_n820, _AES_ENC_us12_n819, _AES_ENC_us12_n818, _AES_ENC_us12_n817, _AES_ENC_us12_n816, _AES_ENC_us12_n815, _AES_ENC_us12_n814, _AES_ENC_us12_n813, _AES_ENC_us12_n812, _AES_ENC_us12_n811, _AES_ENC_us12_n810, _AES_ENC_us12_n809, _AES_ENC_us12_n808, _AES_ENC_us12_n807, _AES_ENC_us12_n806, 
  _AES_ENC_us12_n805, _AES_ENC_us12_n804, _AES_ENC_us12_n803, _AES_ENC_us12_n802, _AES_ENC_us12_n801, _AES_ENC_us12_n800, _AES_ENC_us12_n799, _AES_ENC_us12_n798, _AES_ENC_us12_n797, _AES_ENC_us12_n796, _AES_ENC_us12_n795, _AES_ENC_us12_n794, _AES_ENC_us12_n793, _AES_ENC_us12_n792, _AES_ENC_us12_n791, _AES_ENC_us12_n790, _AES_ENC_us12_n789, _AES_ENC_us12_n788, _AES_ENC_us12_n787, _AES_ENC_us12_n786, _AES_ENC_us12_n785, _AES_ENC_us12_n784, _AES_ENC_us12_n783, _AES_ENC_us12_n782, _AES_ENC_us12_n781, _AES_ENC_us12_n780, _AES_ENC_us12_n779, _AES_ENC_us12_n778, _AES_ENC_us12_n777, _AES_ENC_us12_n776, _AES_ENC_us12_n775, _AES_ENC_us12_n774, _AES_ENC_us12_n773, _AES_ENC_us12_n772, _AES_ENC_us12_n771, _AES_ENC_us12_n770, _AES_ENC_us12_n769, _AES_ENC_us12_n768, _AES_ENC_us12_n767, _AES_ENC_us12_n766, _AES_ENC_us12_n765, _AES_ENC_us12_n764, _AES_ENC_us12_n763, _AES_ENC_us12_n762, _AES_ENC_us12_n761, _AES_ENC_us12_n760, _AES_ENC_us12_n759, _AES_ENC_us12_n758, _AES_ENC_us12_n757, _AES_ENC_us12_n756, 
  _AES_ENC_us12_n755, _AES_ENC_us12_n754, _AES_ENC_us12_n753, _AES_ENC_us12_n752, _AES_ENC_us12_n751, _AES_ENC_us12_n750, _AES_ENC_us12_n749, _AES_ENC_us12_n748, _AES_ENC_us12_n747, _AES_ENC_us12_n746, _AES_ENC_us12_n745, _AES_ENC_us12_n744, _AES_ENC_us12_n743, _AES_ENC_us12_n742, _AES_ENC_us12_n741, _AES_ENC_us12_n740, _AES_ENC_us12_n739, _AES_ENC_us12_n738, _AES_ENC_us12_n737, _AES_ENC_us12_n736, _AES_ENC_us12_n735, _AES_ENC_us12_n734, _AES_ENC_us12_n733, _AES_ENC_us12_n732, _AES_ENC_us12_n731, _AES_ENC_us12_n730, _AES_ENC_us12_n729, _AES_ENC_us12_n728, _AES_ENC_us12_n727, _AES_ENC_us12_n726, _AES_ENC_us12_n725, _AES_ENC_us12_n724, _AES_ENC_us12_n723, _AES_ENC_us12_n722, _AES_ENC_us12_n721, _AES_ENC_us12_n720, _AES_ENC_us12_n719, _AES_ENC_us12_n718, _AES_ENC_us12_n717, _AES_ENC_us12_n716, _AES_ENC_us12_n715, _AES_ENC_us12_n714, _AES_ENC_us12_n713, _AES_ENC_us12_n712, _AES_ENC_us12_n711, _AES_ENC_us12_n710, _AES_ENC_us12_n709, _AES_ENC_us12_n708, _AES_ENC_us12_n707, _AES_ENC_us12_n706, 
  _AES_ENC_us12_n705, _AES_ENC_us12_n704, _AES_ENC_us12_n703, _AES_ENC_us12_n702, _AES_ENC_us12_n701, _AES_ENC_us12_n700, _AES_ENC_us12_n699, _AES_ENC_us12_n698, _AES_ENC_us12_n697, _AES_ENC_us12_n696, _AES_ENC_us12_n695, _AES_ENC_us12_n694, _AES_ENC_us12_n693, _AES_ENC_us12_n692, _AES_ENC_us12_n691, _AES_ENC_us12_n690, _AES_ENC_us12_n689, _AES_ENC_us12_n688, _AES_ENC_us12_n687, _AES_ENC_us12_n686, _AES_ENC_us12_n685, _AES_ENC_us12_n684, _AES_ENC_us12_n683, _AES_ENC_us12_n682, _AES_ENC_us12_n681, _AES_ENC_us12_n680, _AES_ENC_us12_n679, _AES_ENC_us12_n678, _AES_ENC_us12_n677, _AES_ENC_us12_n676, _AES_ENC_us12_n675, _AES_ENC_us12_n674, _AES_ENC_us12_n673, _AES_ENC_us12_n672, _AES_ENC_us12_n671, _AES_ENC_us12_n670, _AES_ENC_us12_n669, _AES_ENC_us12_n668, _AES_ENC_us12_n667, _AES_ENC_us12_n666, _AES_ENC_us12_n665, _AES_ENC_us12_n664, _AES_ENC_us12_n663, _AES_ENC_us12_n662, _AES_ENC_us12_n661, _AES_ENC_us12_n660, _AES_ENC_us12_n659, _AES_ENC_us12_n658, _AES_ENC_us12_n657, _AES_ENC_us12_n656, 
  _AES_ENC_us12_n655, _AES_ENC_us12_n654, _AES_ENC_us12_n653, _AES_ENC_us12_n652, _AES_ENC_us12_n651, _AES_ENC_us12_n650, _AES_ENC_us12_n649, _AES_ENC_us12_n648, _AES_ENC_us12_n647, _AES_ENC_us12_n646, _AES_ENC_us12_n645, _AES_ENC_us12_n644, _AES_ENC_us12_n643, _AES_ENC_us12_n642, _AES_ENC_us12_n641, _AES_ENC_us12_n640, _AES_ENC_us12_n639, _AES_ENC_us12_n638, _AES_ENC_us12_n637, _AES_ENC_us12_n636, _AES_ENC_us12_n635, _AES_ENC_us12_n634, _AES_ENC_us12_n633, _AES_ENC_us12_n632, _AES_ENC_us12_n631, _AES_ENC_us12_n630, _AES_ENC_us12_n629, _AES_ENC_us12_n628, _AES_ENC_us12_n627, _AES_ENC_us12_n626, _AES_ENC_us12_n625, _AES_ENC_us12_n624, _AES_ENC_us12_n623, _AES_ENC_us12_n622, _AES_ENC_us12_n621, _AES_ENC_us12_n620, _AES_ENC_us12_n619, _AES_ENC_us12_n618, _AES_ENC_us12_n617, _AES_ENC_us12_n616, _AES_ENC_us12_n615, _AES_ENC_us12_n614, _AES_ENC_us12_n613, _AES_ENC_us12_n612, _AES_ENC_us12_n611, _AES_ENC_us12_n610, _AES_ENC_us12_n609, _AES_ENC_us12_n608, _AES_ENC_us12_n607, _AES_ENC_us12_n606, 
  _AES_ENC_us12_n605, _AES_ENC_us12_n604, _AES_ENC_us12_n603, _AES_ENC_us12_n602, _AES_ENC_us12_n601, _AES_ENC_us12_n600, _AES_ENC_us12_n599, _AES_ENC_us12_n598, _AES_ENC_us12_n597, _AES_ENC_us12_n596, _AES_ENC_us12_n595, _AES_ENC_us12_n594, _AES_ENC_us12_n593, _AES_ENC_us12_n592, _AES_ENC_us12_n591, _AES_ENC_us12_n590, _AES_ENC_us12_n589, _AES_ENC_us12_n588, _AES_ENC_us12_n587, _AES_ENC_us12_n586, _AES_ENC_us12_n585, _AES_ENC_us12_n584, _AES_ENC_us12_n583, _AES_ENC_us12_n582, _AES_ENC_us12_n581, _AES_ENC_us12_n580, _AES_ENC_us12_n579, _AES_ENC_us12_n578, _AES_ENC_us12_n577, _AES_ENC_us12_n576, _AES_ENC_us12_n575, _AES_ENC_us12_n574, _AES_ENC_us12_n573, _AES_ENC_us12_n572, _AES_ENC_us12_n571, _AES_ENC_us12_n570, _AES_ENC_us12_n569, _AES_ENC_us13_n1135, _AES_ENC_us13_n1134, _AES_ENC_us13_n1133, _AES_ENC_us13_n1132, _AES_ENC_us13_n1131, _AES_ENC_us13_n1130, _AES_ENC_us13_n1129, _AES_ENC_us13_n1128, _AES_ENC_us13_n1127, _AES_ENC_us13_n1126, _AES_ENC_us13_n1125, _AES_ENC_us13_n1124, _AES_ENC_us13_n1123, 
  _AES_ENC_us13_n1122, _AES_ENC_us13_n1121, _AES_ENC_us13_n1120, _AES_ENC_us13_n1119, _AES_ENC_us13_n1118, _AES_ENC_us13_n1117, _AES_ENC_us13_n1116, _AES_ENC_us13_n1115, _AES_ENC_us13_n1114, _AES_ENC_us13_n1113, _AES_ENC_us13_n1112, _AES_ENC_us13_n1111, _AES_ENC_us13_n1110, _AES_ENC_us13_n1109, _AES_ENC_us13_n1108, _AES_ENC_us13_n1107, _AES_ENC_us13_n1106, _AES_ENC_us13_n1105, _AES_ENC_us13_n1104, _AES_ENC_us13_n1103, _AES_ENC_us13_n1102, _AES_ENC_us13_n1101, _AES_ENC_us13_n1100, _AES_ENC_us13_n1099, _AES_ENC_us13_n1098, _AES_ENC_us13_n1097, _AES_ENC_us13_n1096, _AES_ENC_us13_n1095, _AES_ENC_us13_n1094, _AES_ENC_us13_n1093, _AES_ENC_us13_n1092, _AES_ENC_us13_n1091, _AES_ENC_us13_n1090, _AES_ENC_us13_n1089, _AES_ENC_us13_n1088, _AES_ENC_us13_n1087, _AES_ENC_us13_n1086, _AES_ENC_us13_n1085, _AES_ENC_us13_n1084, _AES_ENC_us13_n1083, _AES_ENC_us13_n1082, _AES_ENC_us13_n1081, _AES_ENC_us13_n1080, _AES_ENC_us13_n1079, _AES_ENC_us13_n1078, _AES_ENC_us13_n1077, _AES_ENC_us13_n1076, _AES_ENC_us13_n1075, _AES_ENC_us13_n1074, _AES_ENC_us13_n1073, 
  _AES_ENC_us13_n1072, _AES_ENC_us13_n1071, _AES_ENC_us13_n1070, _AES_ENC_us13_n1069, _AES_ENC_us13_n1068, _AES_ENC_us13_n1067, _AES_ENC_us13_n1066, _AES_ENC_us13_n1065, _AES_ENC_us13_n1064, _AES_ENC_us13_n1063, _AES_ENC_us13_n1062, _AES_ENC_us13_n1061, _AES_ENC_us13_n1060, _AES_ENC_us13_n1059, _AES_ENC_us13_n1058, _AES_ENC_us13_n1057, _AES_ENC_us13_n1056, _AES_ENC_us13_n1055, _AES_ENC_us13_n1054, _AES_ENC_us13_n1053, _AES_ENC_us13_n1052, _AES_ENC_us13_n1051, _AES_ENC_us13_n1050, _AES_ENC_us13_n1049, _AES_ENC_us13_n1048, _AES_ENC_us13_n1047, _AES_ENC_us13_n1046, _AES_ENC_us13_n1045, _AES_ENC_us13_n1044, _AES_ENC_us13_n1043, _AES_ENC_us13_n1042, _AES_ENC_us13_n1041, _AES_ENC_us13_n1040, _AES_ENC_us13_n1039, _AES_ENC_us13_n1038, _AES_ENC_us13_n1037, _AES_ENC_us13_n1036, _AES_ENC_us13_n1035, _AES_ENC_us13_n1034, _AES_ENC_us13_n1033, _AES_ENC_us13_n1032, _AES_ENC_us13_n1031, _AES_ENC_us13_n1030, _AES_ENC_us13_n1029, _AES_ENC_us13_n1028, _AES_ENC_us13_n1027, _AES_ENC_us13_n1026, _AES_ENC_us13_n1025, _AES_ENC_us13_n1024, _AES_ENC_us13_n1023, 
  _AES_ENC_us13_n1022, _AES_ENC_us13_n1021, _AES_ENC_us13_n1020, _AES_ENC_us13_n1019, _AES_ENC_us13_n1018, _AES_ENC_us13_n1017, _AES_ENC_us13_n1016, _AES_ENC_us13_n1015, _AES_ENC_us13_n1014, _AES_ENC_us13_n1013, _AES_ENC_us13_n1012, _AES_ENC_us13_n1011, _AES_ENC_us13_n1010, _AES_ENC_us13_n1009, _AES_ENC_us13_n1008, _AES_ENC_us13_n1007, _AES_ENC_us13_n1006, _AES_ENC_us13_n1005, _AES_ENC_us13_n1004, _AES_ENC_us13_n1003, _AES_ENC_us13_n1002, _AES_ENC_us13_n1001, _AES_ENC_us13_n1000, _AES_ENC_us13_n999, _AES_ENC_us13_n998, _AES_ENC_us13_n997, _AES_ENC_us13_n996, _AES_ENC_us13_n995, _AES_ENC_us13_n994, _AES_ENC_us13_n993, _AES_ENC_us13_n992, _AES_ENC_us13_n991, _AES_ENC_us13_n990, _AES_ENC_us13_n989, _AES_ENC_us13_n988, _AES_ENC_us13_n987, _AES_ENC_us13_n986, _AES_ENC_us13_n985, _AES_ENC_us13_n984, _AES_ENC_us13_n983, _AES_ENC_us13_n982, _AES_ENC_us13_n981, _AES_ENC_us13_n980, _AES_ENC_us13_n979, _AES_ENC_us13_n978, _AES_ENC_us13_n977, _AES_ENC_us13_n976, _AES_ENC_us13_n975, _AES_ENC_us13_n974, _AES_ENC_us13_n973, 
  _AES_ENC_us13_n972, _AES_ENC_us13_n971, _AES_ENC_us13_n970, _AES_ENC_us13_n969, _AES_ENC_us13_n968, _AES_ENC_us13_n967, _AES_ENC_us13_n966, _AES_ENC_us13_n965, _AES_ENC_us13_n964, _AES_ENC_us13_n963, _AES_ENC_us13_n962, _AES_ENC_us13_n961, _AES_ENC_us13_n960, _AES_ENC_us13_n959, _AES_ENC_us13_n958, _AES_ENC_us13_n957, _AES_ENC_us13_n956, _AES_ENC_us13_n955, _AES_ENC_us13_n954, _AES_ENC_us13_n953, _AES_ENC_us13_n952, _AES_ENC_us13_n951, _AES_ENC_us13_n950, _AES_ENC_us13_n949, _AES_ENC_us13_n948, _AES_ENC_us13_n947, _AES_ENC_us13_n946, _AES_ENC_us13_n945, _AES_ENC_us13_n944, _AES_ENC_us13_n943, _AES_ENC_us13_n942, _AES_ENC_us13_n941, _AES_ENC_us13_n940, _AES_ENC_us13_n939, _AES_ENC_us13_n938, _AES_ENC_us13_n937, _AES_ENC_us13_n936, _AES_ENC_us13_n935, _AES_ENC_us13_n934, _AES_ENC_us13_n933, _AES_ENC_us13_n932, _AES_ENC_us13_n931, _AES_ENC_us13_n930, _AES_ENC_us13_n929, _AES_ENC_us13_n928, _AES_ENC_us13_n927, _AES_ENC_us13_n926, _AES_ENC_us13_n925, _AES_ENC_us13_n924, _AES_ENC_us13_n923, 
  _AES_ENC_us13_n922, _AES_ENC_us13_n921, _AES_ENC_us13_n920, _AES_ENC_us13_n919, _AES_ENC_us13_n918, _AES_ENC_us13_n917, _AES_ENC_us13_n916, _AES_ENC_us13_n915, _AES_ENC_us13_n914, _AES_ENC_us13_n913, _AES_ENC_us13_n912, _AES_ENC_us13_n911, _AES_ENC_us13_n910, _AES_ENC_us13_n909, _AES_ENC_us13_n908, _AES_ENC_us13_n907, _AES_ENC_us13_n906, _AES_ENC_us13_n905, _AES_ENC_us13_n904, _AES_ENC_us13_n903, _AES_ENC_us13_n902, _AES_ENC_us13_n901, _AES_ENC_us13_n900, _AES_ENC_us13_n899, _AES_ENC_us13_n898, _AES_ENC_us13_n897, _AES_ENC_us13_n896, _AES_ENC_us13_n895, _AES_ENC_us13_n894, _AES_ENC_us13_n893, _AES_ENC_us13_n892, _AES_ENC_us13_n891, _AES_ENC_us13_n890, _AES_ENC_us13_n889, _AES_ENC_us13_n888, _AES_ENC_us13_n887, _AES_ENC_us13_n886, _AES_ENC_us13_n885, _AES_ENC_us13_n884, _AES_ENC_us13_n883, _AES_ENC_us13_n882, _AES_ENC_us13_n881, _AES_ENC_us13_n880, _AES_ENC_us13_n879, _AES_ENC_us13_n878, _AES_ENC_us13_n877, _AES_ENC_us13_n876, _AES_ENC_us13_n875, _AES_ENC_us13_n874, _AES_ENC_us13_n873, 
  _AES_ENC_us13_n872, _AES_ENC_us13_n871, _AES_ENC_us13_n870, _AES_ENC_us13_n869, _AES_ENC_us13_n868, _AES_ENC_us13_n867, _AES_ENC_us13_n866, _AES_ENC_us13_n865, _AES_ENC_us13_n864, _AES_ENC_us13_n863, _AES_ENC_us13_n862, _AES_ENC_us13_n861, _AES_ENC_us13_n860, _AES_ENC_us13_n859, _AES_ENC_us13_n858, _AES_ENC_us13_n857, _AES_ENC_us13_n856, _AES_ENC_us13_n855, _AES_ENC_us13_n854, _AES_ENC_us13_n853, _AES_ENC_us13_n852, _AES_ENC_us13_n851, _AES_ENC_us13_n850, _AES_ENC_us13_n849, _AES_ENC_us13_n848, _AES_ENC_us13_n847, _AES_ENC_us13_n846, _AES_ENC_us13_n845, _AES_ENC_us13_n844, _AES_ENC_us13_n843, _AES_ENC_us13_n842, _AES_ENC_us13_n841, _AES_ENC_us13_n840, _AES_ENC_us13_n839, _AES_ENC_us13_n838, _AES_ENC_us13_n837, _AES_ENC_us13_n836, _AES_ENC_us13_n835, _AES_ENC_us13_n834, _AES_ENC_us13_n833, _AES_ENC_us13_n832, _AES_ENC_us13_n831, _AES_ENC_us13_n830, _AES_ENC_us13_n829, _AES_ENC_us13_n828, _AES_ENC_us13_n827, _AES_ENC_us13_n826, _AES_ENC_us13_n825, _AES_ENC_us13_n824, _AES_ENC_us13_n823, 
  _AES_ENC_us13_n822, _AES_ENC_us13_n821, _AES_ENC_us13_n820, _AES_ENC_us13_n819, _AES_ENC_us13_n818, _AES_ENC_us13_n817, _AES_ENC_us13_n816, _AES_ENC_us13_n815, _AES_ENC_us13_n814, _AES_ENC_us13_n813, _AES_ENC_us13_n812, _AES_ENC_us13_n811, _AES_ENC_us13_n810, _AES_ENC_us13_n809, _AES_ENC_us13_n808, _AES_ENC_us13_n807, _AES_ENC_us13_n806, _AES_ENC_us13_n805, _AES_ENC_us13_n804, _AES_ENC_us13_n803, _AES_ENC_us13_n802, _AES_ENC_us13_n801, _AES_ENC_us13_n800, _AES_ENC_us13_n799, _AES_ENC_us13_n798, _AES_ENC_us13_n797, _AES_ENC_us13_n796, _AES_ENC_us13_n795, _AES_ENC_us13_n794, _AES_ENC_us13_n793, _AES_ENC_us13_n792, _AES_ENC_us13_n791, _AES_ENC_us13_n790, _AES_ENC_us13_n789, _AES_ENC_us13_n788, _AES_ENC_us13_n787, _AES_ENC_us13_n786, _AES_ENC_us13_n785, _AES_ENC_us13_n784, _AES_ENC_us13_n783, _AES_ENC_us13_n782, _AES_ENC_us13_n781, _AES_ENC_us13_n780, _AES_ENC_us13_n779, _AES_ENC_us13_n778, _AES_ENC_us13_n777, _AES_ENC_us13_n776, _AES_ENC_us13_n775, _AES_ENC_us13_n774, _AES_ENC_us13_n773, 
  _AES_ENC_us13_n772, _AES_ENC_us13_n771, _AES_ENC_us13_n770, _AES_ENC_us13_n769, _AES_ENC_us13_n768, _AES_ENC_us13_n767, _AES_ENC_us13_n766, _AES_ENC_us13_n765, _AES_ENC_us13_n764, _AES_ENC_us13_n763, _AES_ENC_us13_n762, _AES_ENC_us13_n761, _AES_ENC_us13_n760, _AES_ENC_us13_n759, _AES_ENC_us13_n758, _AES_ENC_us13_n757, _AES_ENC_us13_n756, _AES_ENC_us13_n755, _AES_ENC_us13_n754, _AES_ENC_us13_n753, _AES_ENC_us13_n752, _AES_ENC_us13_n751, _AES_ENC_us13_n750, _AES_ENC_us13_n749, _AES_ENC_us13_n748, _AES_ENC_us13_n747, _AES_ENC_us13_n746, _AES_ENC_us13_n745, _AES_ENC_us13_n744, _AES_ENC_us13_n743, _AES_ENC_us13_n742, _AES_ENC_us13_n741, _AES_ENC_us13_n740, _AES_ENC_us13_n739, _AES_ENC_us13_n738, _AES_ENC_us13_n737, _AES_ENC_us13_n736, _AES_ENC_us13_n735, _AES_ENC_us13_n734, _AES_ENC_us13_n733, _AES_ENC_us13_n732, _AES_ENC_us13_n731, _AES_ENC_us13_n730, _AES_ENC_us13_n729, _AES_ENC_us13_n728, _AES_ENC_us13_n727, _AES_ENC_us13_n726, _AES_ENC_us13_n725, _AES_ENC_us13_n724, _AES_ENC_us13_n723, 
  _AES_ENC_us13_n722, _AES_ENC_us13_n721, _AES_ENC_us13_n720, _AES_ENC_us13_n719, _AES_ENC_us13_n718, _AES_ENC_us13_n717, _AES_ENC_us13_n716, _AES_ENC_us13_n715, _AES_ENC_us13_n714, _AES_ENC_us13_n713, _AES_ENC_us13_n712, _AES_ENC_us13_n711, _AES_ENC_us13_n710, _AES_ENC_us13_n709, _AES_ENC_us13_n708, _AES_ENC_us13_n707, _AES_ENC_us13_n706, _AES_ENC_us13_n705, _AES_ENC_us13_n704, _AES_ENC_us13_n703, _AES_ENC_us13_n702, _AES_ENC_us13_n701, _AES_ENC_us13_n700, _AES_ENC_us13_n699, _AES_ENC_us13_n698, _AES_ENC_us13_n697, _AES_ENC_us13_n696, _AES_ENC_us13_n695, _AES_ENC_us13_n694, _AES_ENC_us13_n693, _AES_ENC_us13_n692, _AES_ENC_us13_n691, _AES_ENC_us13_n690, _AES_ENC_us13_n689, _AES_ENC_us13_n688, _AES_ENC_us13_n687, _AES_ENC_us13_n686, _AES_ENC_us13_n685, _AES_ENC_us13_n684, _AES_ENC_us13_n683, _AES_ENC_us13_n682, _AES_ENC_us13_n681, _AES_ENC_us13_n680, _AES_ENC_us13_n679, _AES_ENC_us13_n678, _AES_ENC_us13_n677, _AES_ENC_us13_n676, _AES_ENC_us13_n675, _AES_ENC_us13_n674, _AES_ENC_us13_n673, 
  _AES_ENC_us13_n672, _AES_ENC_us13_n671, _AES_ENC_us13_n670, _AES_ENC_us13_n669, _AES_ENC_us13_n668, _AES_ENC_us13_n667, _AES_ENC_us13_n666, _AES_ENC_us13_n665, _AES_ENC_us13_n664, _AES_ENC_us13_n663, _AES_ENC_us13_n662, _AES_ENC_us13_n661, _AES_ENC_us13_n660, _AES_ENC_us13_n659, _AES_ENC_us13_n658, _AES_ENC_us13_n657, _AES_ENC_us13_n656, _AES_ENC_us13_n655, _AES_ENC_us13_n654, _AES_ENC_us13_n653, _AES_ENC_us13_n652, _AES_ENC_us13_n651, _AES_ENC_us13_n650, _AES_ENC_us13_n649, _AES_ENC_us13_n648, _AES_ENC_us13_n647, _AES_ENC_us13_n646, _AES_ENC_us13_n645, _AES_ENC_us13_n644, _AES_ENC_us13_n643, _AES_ENC_us13_n642, _AES_ENC_us13_n641, _AES_ENC_us13_n640, _AES_ENC_us13_n639, _AES_ENC_us13_n638, _AES_ENC_us13_n637, _AES_ENC_us13_n636, _AES_ENC_us13_n635, _AES_ENC_us13_n634, _AES_ENC_us13_n633, _AES_ENC_us13_n632, _AES_ENC_us13_n631, _AES_ENC_us13_n630, _AES_ENC_us13_n629, _AES_ENC_us13_n628, _AES_ENC_us13_n627, _AES_ENC_us13_n626, _AES_ENC_us13_n625, _AES_ENC_us13_n624, _AES_ENC_us13_n623, 
  _AES_ENC_us13_n622, _AES_ENC_us13_n621, _AES_ENC_us13_n620, _AES_ENC_us13_n619, _AES_ENC_us13_n618, _AES_ENC_us13_n617, _AES_ENC_us13_n616, _AES_ENC_us13_n615, _AES_ENC_us13_n614, _AES_ENC_us13_n613, _AES_ENC_us13_n612, _AES_ENC_us13_n611, _AES_ENC_us13_n610, _AES_ENC_us13_n609, _AES_ENC_us13_n608, _AES_ENC_us13_n607, _AES_ENC_us13_n606, _AES_ENC_us13_n605, _AES_ENC_us13_n604, _AES_ENC_us13_n603, _AES_ENC_us13_n602, _AES_ENC_us13_n601, _AES_ENC_us13_n600, _AES_ENC_us13_n599, _AES_ENC_us13_n598, _AES_ENC_us13_n597, _AES_ENC_us13_n596, _AES_ENC_us13_n595, _AES_ENC_us13_n594, _AES_ENC_us13_n593, _AES_ENC_us13_n592, _AES_ENC_us13_n591, _AES_ENC_us13_n590, _AES_ENC_us13_n589, _AES_ENC_us13_n588, _AES_ENC_us13_n587, _AES_ENC_us13_n586, _AES_ENC_us13_n585, _AES_ENC_us13_n584, _AES_ENC_us13_n583, _AES_ENC_us13_n582, _AES_ENC_us13_n581, _AES_ENC_us13_n580, _AES_ENC_us13_n579, _AES_ENC_us13_n578, _AES_ENC_us13_n577, _AES_ENC_us13_n576, _AES_ENC_us13_n575, _AES_ENC_us13_n574, _AES_ENC_us13_n573, 
  _AES_ENC_us13_n572, _AES_ENC_us13_n571, _AES_ENC_us13_n570, _AES_ENC_us13_n569, _AES_ENC_us20_n1135, _AES_ENC_us20_n1134, _AES_ENC_us20_n1133, _AES_ENC_us20_n1132, _AES_ENC_us20_n1131, _AES_ENC_us20_n1130, _AES_ENC_us20_n1129, _AES_ENC_us20_n1128, _AES_ENC_us20_n1127, _AES_ENC_us20_n1126, _AES_ENC_us20_n1125, _AES_ENC_us20_n1124, _AES_ENC_us20_n1123, _AES_ENC_us20_n1122, _AES_ENC_us20_n1121, _AES_ENC_us20_n1120, _AES_ENC_us20_n1119, _AES_ENC_us20_n1118, _AES_ENC_us20_n1117, _AES_ENC_us20_n1116, _AES_ENC_us20_n1115, _AES_ENC_us20_n1114, _AES_ENC_us20_n1113, _AES_ENC_us20_n1112, _AES_ENC_us20_n1111, _AES_ENC_us20_n1110, _AES_ENC_us20_n1109, _AES_ENC_us20_n1108, _AES_ENC_us20_n1107, _AES_ENC_us20_n1106, _AES_ENC_us20_n1105, _AES_ENC_us20_n1104, _AES_ENC_us20_n1103, _AES_ENC_us20_n1102, _AES_ENC_us20_n1101, _AES_ENC_us20_n1100, _AES_ENC_us20_n1099, _AES_ENC_us20_n1098, _AES_ENC_us20_n1097, _AES_ENC_us20_n1096, _AES_ENC_us20_n1095, _AES_ENC_us20_n1094, _AES_ENC_us20_n1093, _AES_ENC_us20_n1092, _AES_ENC_us20_n1091, _AES_ENC_us20_n1090, 
  _AES_ENC_us20_n1089, _AES_ENC_us20_n1088, _AES_ENC_us20_n1087, _AES_ENC_us20_n1086, _AES_ENC_us20_n1085, _AES_ENC_us20_n1084, _AES_ENC_us20_n1083, _AES_ENC_us20_n1082, _AES_ENC_us20_n1081, _AES_ENC_us20_n1080, _AES_ENC_us20_n1079, _AES_ENC_us20_n1078, _AES_ENC_us20_n1077, _AES_ENC_us20_n1076, _AES_ENC_us20_n1075, _AES_ENC_us20_n1074, _AES_ENC_us20_n1073, _AES_ENC_us20_n1072, _AES_ENC_us20_n1071, _AES_ENC_us20_n1070, _AES_ENC_us20_n1069, _AES_ENC_us20_n1068, _AES_ENC_us20_n1067, _AES_ENC_us20_n1066, _AES_ENC_us20_n1065, _AES_ENC_us20_n1064, _AES_ENC_us20_n1063, _AES_ENC_us20_n1062, _AES_ENC_us20_n1061, _AES_ENC_us20_n1060, _AES_ENC_us20_n1059, _AES_ENC_us20_n1058, _AES_ENC_us20_n1057, _AES_ENC_us20_n1056, _AES_ENC_us20_n1055, _AES_ENC_us20_n1054, _AES_ENC_us20_n1053, _AES_ENC_us20_n1052, _AES_ENC_us20_n1051, _AES_ENC_us20_n1050, _AES_ENC_us20_n1049, _AES_ENC_us20_n1048, _AES_ENC_us20_n1047, _AES_ENC_us20_n1046, _AES_ENC_us20_n1045, _AES_ENC_us20_n1044, _AES_ENC_us20_n1043, _AES_ENC_us20_n1042, _AES_ENC_us20_n1041, _AES_ENC_us20_n1040, 
  _AES_ENC_us20_n1039, _AES_ENC_us20_n1038, _AES_ENC_us20_n1037, _AES_ENC_us20_n1036, _AES_ENC_us20_n1035, _AES_ENC_us20_n1034, _AES_ENC_us20_n1033, _AES_ENC_us20_n1032, _AES_ENC_us20_n1031, _AES_ENC_us20_n1030, _AES_ENC_us20_n1029, _AES_ENC_us20_n1028, _AES_ENC_us20_n1027, _AES_ENC_us20_n1026, _AES_ENC_us20_n1025, _AES_ENC_us20_n1024, _AES_ENC_us20_n1023, _AES_ENC_us20_n1022, _AES_ENC_us20_n1021, _AES_ENC_us20_n1020, _AES_ENC_us20_n1019, _AES_ENC_us20_n1018, _AES_ENC_us20_n1017, _AES_ENC_us20_n1016, _AES_ENC_us20_n1015, _AES_ENC_us20_n1014, _AES_ENC_us20_n1013, _AES_ENC_us20_n1012, _AES_ENC_us20_n1011, _AES_ENC_us20_n1010, _AES_ENC_us20_n1009, _AES_ENC_us20_n1008, _AES_ENC_us20_n1007, _AES_ENC_us20_n1006, _AES_ENC_us20_n1005, _AES_ENC_us20_n1004, _AES_ENC_us20_n1003, _AES_ENC_us20_n1002, _AES_ENC_us20_n1001, _AES_ENC_us20_n1000, _AES_ENC_us20_n999, _AES_ENC_us20_n998, _AES_ENC_us20_n997, _AES_ENC_us20_n996, _AES_ENC_us20_n995, _AES_ENC_us20_n994, _AES_ENC_us20_n993, _AES_ENC_us20_n992, _AES_ENC_us20_n991, _AES_ENC_us20_n990, 
  _AES_ENC_us20_n989, _AES_ENC_us20_n988, _AES_ENC_us20_n987, _AES_ENC_us20_n986, _AES_ENC_us20_n985, _AES_ENC_us20_n984, _AES_ENC_us20_n983, _AES_ENC_us20_n982, _AES_ENC_us20_n981, _AES_ENC_us20_n980, _AES_ENC_us20_n979, _AES_ENC_us20_n978, _AES_ENC_us20_n977, _AES_ENC_us20_n976, _AES_ENC_us20_n975, _AES_ENC_us20_n974, _AES_ENC_us20_n973, _AES_ENC_us20_n972, _AES_ENC_us20_n971, _AES_ENC_us20_n970, _AES_ENC_us20_n969, _AES_ENC_us20_n968, _AES_ENC_us20_n967, _AES_ENC_us20_n966, _AES_ENC_us20_n965, _AES_ENC_us20_n964, _AES_ENC_us20_n963, _AES_ENC_us20_n962, _AES_ENC_us20_n961, _AES_ENC_us20_n960, _AES_ENC_us20_n959, _AES_ENC_us20_n958, _AES_ENC_us20_n957, _AES_ENC_us20_n956, _AES_ENC_us20_n955, _AES_ENC_us20_n954, _AES_ENC_us20_n953, _AES_ENC_us20_n952, _AES_ENC_us20_n951, _AES_ENC_us20_n950, _AES_ENC_us20_n949, _AES_ENC_us20_n948, _AES_ENC_us20_n947, _AES_ENC_us20_n946, _AES_ENC_us20_n945, _AES_ENC_us20_n944, _AES_ENC_us20_n943, _AES_ENC_us20_n942, _AES_ENC_us20_n941, _AES_ENC_us20_n940, 
  _AES_ENC_us20_n939, _AES_ENC_us20_n938, _AES_ENC_us20_n937, _AES_ENC_us20_n936, _AES_ENC_us20_n935, _AES_ENC_us20_n934, _AES_ENC_us20_n933, _AES_ENC_us20_n932, _AES_ENC_us20_n931, _AES_ENC_us20_n930, _AES_ENC_us20_n929, _AES_ENC_us20_n928, _AES_ENC_us20_n927, _AES_ENC_us20_n926, _AES_ENC_us20_n925, _AES_ENC_us20_n924, _AES_ENC_us20_n923, _AES_ENC_us20_n922, _AES_ENC_us20_n921, _AES_ENC_us20_n920, _AES_ENC_us20_n919, _AES_ENC_us20_n918, _AES_ENC_us20_n917, _AES_ENC_us20_n916, _AES_ENC_us20_n915, _AES_ENC_us20_n914, _AES_ENC_us20_n913, _AES_ENC_us20_n912, _AES_ENC_us20_n911, _AES_ENC_us20_n910, _AES_ENC_us20_n909, _AES_ENC_us20_n908, _AES_ENC_us20_n907, _AES_ENC_us20_n906, _AES_ENC_us20_n905, _AES_ENC_us20_n904, _AES_ENC_us20_n903, _AES_ENC_us20_n902, _AES_ENC_us20_n901, _AES_ENC_us20_n900, _AES_ENC_us20_n899, _AES_ENC_us20_n898, _AES_ENC_us20_n897, _AES_ENC_us20_n896, _AES_ENC_us20_n895, _AES_ENC_us20_n894, _AES_ENC_us20_n893, _AES_ENC_us20_n892, _AES_ENC_us20_n891, _AES_ENC_us20_n890, 
  _AES_ENC_us20_n889, _AES_ENC_us20_n888, _AES_ENC_us20_n887, _AES_ENC_us20_n886, _AES_ENC_us20_n885, _AES_ENC_us20_n884, _AES_ENC_us20_n883, _AES_ENC_us20_n882, _AES_ENC_us20_n881, _AES_ENC_us20_n880, _AES_ENC_us20_n879, _AES_ENC_us20_n878, _AES_ENC_us20_n877, _AES_ENC_us20_n876, _AES_ENC_us20_n875, _AES_ENC_us20_n874, _AES_ENC_us20_n873, _AES_ENC_us20_n872, _AES_ENC_us20_n871, _AES_ENC_us20_n870, _AES_ENC_us20_n869, _AES_ENC_us20_n868, _AES_ENC_us20_n867, _AES_ENC_us20_n866, _AES_ENC_us20_n865, _AES_ENC_us20_n864, _AES_ENC_us20_n863, _AES_ENC_us20_n862, _AES_ENC_us20_n861, _AES_ENC_us20_n860, _AES_ENC_us20_n859, _AES_ENC_us20_n858, _AES_ENC_us20_n857, _AES_ENC_us20_n856, _AES_ENC_us20_n855, _AES_ENC_us20_n854, _AES_ENC_us20_n853, _AES_ENC_us20_n852, _AES_ENC_us20_n851, _AES_ENC_us20_n850, _AES_ENC_us20_n849, _AES_ENC_us20_n848, _AES_ENC_us20_n847, _AES_ENC_us20_n846, _AES_ENC_us20_n845, _AES_ENC_us20_n844, _AES_ENC_us20_n843, _AES_ENC_us20_n842, _AES_ENC_us20_n841, _AES_ENC_us20_n840, 
  _AES_ENC_us20_n839, _AES_ENC_us20_n838, _AES_ENC_us20_n837, _AES_ENC_us20_n836, _AES_ENC_us20_n835, _AES_ENC_us20_n834, _AES_ENC_us20_n833, _AES_ENC_us20_n832, _AES_ENC_us20_n831, _AES_ENC_us20_n830, _AES_ENC_us20_n829, _AES_ENC_us20_n828, _AES_ENC_us20_n827, _AES_ENC_us20_n826, _AES_ENC_us20_n825, _AES_ENC_us20_n824, _AES_ENC_us20_n823, _AES_ENC_us20_n822, _AES_ENC_us20_n821, _AES_ENC_us20_n820, _AES_ENC_us20_n819, _AES_ENC_us20_n818, _AES_ENC_us20_n817, _AES_ENC_us20_n816, _AES_ENC_us20_n815, _AES_ENC_us20_n814, _AES_ENC_us20_n813, _AES_ENC_us20_n812, _AES_ENC_us20_n811, _AES_ENC_us20_n810, _AES_ENC_us20_n809, _AES_ENC_us20_n808, _AES_ENC_us20_n807, _AES_ENC_us20_n806, _AES_ENC_us20_n805, _AES_ENC_us20_n804, _AES_ENC_us20_n803, _AES_ENC_us20_n802, _AES_ENC_us20_n801, _AES_ENC_us20_n800, _AES_ENC_us20_n799, _AES_ENC_us20_n798, _AES_ENC_us20_n797, _AES_ENC_us20_n796, _AES_ENC_us20_n795, _AES_ENC_us20_n794, _AES_ENC_us20_n793, _AES_ENC_us20_n792, _AES_ENC_us20_n791, _AES_ENC_us20_n790, 
  _AES_ENC_us20_n789, _AES_ENC_us20_n788, _AES_ENC_us20_n787, _AES_ENC_us20_n786, _AES_ENC_us20_n785, _AES_ENC_us20_n784, _AES_ENC_us20_n783, _AES_ENC_us20_n782, _AES_ENC_us20_n781, _AES_ENC_us20_n780, _AES_ENC_us20_n779, _AES_ENC_us20_n778, _AES_ENC_us20_n777, _AES_ENC_us20_n776, _AES_ENC_us20_n775, _AES_ENC_us20_n774, _AES_ENC_us20_n773, _AES_ENC_us20_n772, _AES_ENC_us20_n771, _AES_ENC_us20_n770, _AES_ENC_us20_n769, _AES_ENC_us20_n768, _AES_ENC_us20_n767, _AES_ENC_us20_n766, _AES_ENC_us20_n765, _AES_ENC_us20_n764, _AES_ENC_us20_n763, _AES_ENC_us20_n762, _AES_ENC_us20_n761, _AES_ENC_us20_n760, _AES_ENC_us20_n759, _AES_ENC_us20_n758, _AES_ENC_us20_n757, _AES_ENC_us20_n756, _AES_ENC_us20_n755, _AES_ENC_us20_n754, _AES_ENC_us20_n753, _AES_ENC_us20_n752, _AES_ENC_us20_n751, _AES_ENC_us20_n750, _AES_ENC_us20_n749, _AES_ENC_us20_n748, _AES_ENC_us20_n747, _AES_ENC_us20_n746, _AES_ENC_us20_n745, _AES_ENC_us20_n744, _AES_ENC_us20_n743, _AES_ENC_us20_n742, _AES_ENC_us20_n741, _AES_ENC_us20_n740, 
  _AES_ENC_us20_n739, _AES_ENC_us20_n738, _AES_ENC_us20_n737, _AES_ENC_us20_n736, _AES_ENC_us20_n735, _AES_ENC_us20_n734, _AES_ENC_us20_n733, _AES_ENC_us20_n732, _AES_ENC_us20_n731, _AES_ENC_us20_n730, _AES_ENC_us20_n729, _AES_ENC_us20_n728, _AES_ENC_us20_n727, _AES_ENC_us20_n726, _AES_ENC_us20_n725, _AES_ENC_us20_n724, _AES_ENC_us20_n723, _AES_ENC_us20_n722, _AES_ENC_us20_n721, _AES_ENC_us20_n720, _AES_ENC_us20_n719, _AES_ENC_us20_n718, _AES_ENC_us20_n717, _AES_ENC_us20_n716, _AES_ENC_us20_n715, _AES_ENC_us20_n714, _AES_ENC_us20_n713, _AES_ENC_us20_n712, _AES_ENC_us20_n711, _AES_ENC_us20_n710, _AES_ENC_us20_n709, _AES_ENC_us20_n708, _AES_ENC_us20_n707, _AES_ENC_us20_n706, _AES_ENC_us20_n705, _AES_ENC_us20_n704, _AES_ENC_us20_n703, _AES_ENC_us20_n702, _AES_ENC_us20_n701, _AES_ENC_us20_n700, _AES_ENC_us20_n699, _AES_ENC_us20_n698, _AES_ENC_us20_n697, _AES_ENC_us20_n696, _AES_ENC_us20_n695, _AES_ENC_us20_n694, _AES_ENC_us20_n693, _AES_ENC_us20_n692, _AES_ENC_us20_n691, _AES_ENC_us20_n690, 
  _AES_ENC_us20_n689, _AES_ENC_us20_n688, _AES_ENC_us20_n687, _AES_ENC_us20_n686, _AES_ENC_us20_n685, _AES_ENC_us20_n684, _AES_ENC_us20_n683, _AES_ENC_us20_n682, _AES_ENC_us20_n681, _AES_ENC_us20_n680, _AES_ENC_us20_n679, _AES_ENC_us20_n678, _AES_ENC_us20_n677, _AES_ENC_us20_n676, _AES_ENC_us20_n675, _AES_ENC_us20_n674, _AES_ENC_us20_n673, _AES_ENC_us20_n672, _AES_ENC_us20_n671, _AES_ENC_us20_n670, _AES_ENC_us20_n669, _AES_ENC_us20_n668, _AES_ENC_us20_n667, _AES_ENC_us20_n666, _AES_ENC_us20_n665, _AES_ENC_us20_n664, _AES_ENC_us20_n663, _AES_ENC_us20_n662, _AES_ENC_us20_n661, _AES_ENC_us20_n660, _AES_ENC_us20_n659, _AES_ENC_us20_n658, _AES_ENC_us20_n657, _AES_ENC_us20_n656, _AES_ENC_us20_n655, _AES_ENC_us20_n654, _AES_ENC_us20_n653, _AES_ENC_us20_n652, _AES_ENC_us20_n651, _AES_ENC_us20_n650, _AES_ENC_us20_n649, _AES_ENC_us20_n648, _AES_ENC_us20_n647, _AES_ENC_us20_n646, _AES_ENC_us20_n645, _AES_ENC_us20_n644, _AES_ENC_us20_n643, _AES_ENC_us20_n642, _AES_ENC_us20_n641, _AES_ENC_us20_n640, 
  _AES_ENC_us20_n639, _AES_ENC_us20_n638, _AES_ENC_us20_n637, _AES_ENC_us20_n636, _AES_ENC_us20_n635, _AES_ENC_us20_n634, _AES_ENC_us20_n633, _AES_ENC_us20_n632, _AES_ENC_us20_n631, _AES_ENC_us20_n630, _AES_ENC_us20_n629, _AES_ENC_us20_n628, _AES_ENC_us20_n627, _AES_ENC_us20_n626, _AES_ENC_us20_n625, _AES_ENC_us20_n624, _AES_ENC_us20_n623, _AES_ENC_us20_n622, _AES_ENC_us20_n621, _AES_ENC_us20_n620, _AES_ENC_us20_n619, _AES_ENC_us20_n618, _AES_ENC_us20_n617, _AES_ENC_us20_n616, _AES_ENC_us20_n615, _AES_ENC_us20_n614, _AES_ENC_us20_n613, _AES_ENC_us20_n612, _AES_ENC_us20_n611, _AES_ENC_us20_n610, _AES_ENC_us20_n609, _AES_ENC_us20_n608, _AES_ENC_us20_n607, _AES_ENC_us20_n606, _AES_ENC_us20_n605, _AES_ENC_us20_n604, _AES_ENC_us20_n603, _AES_ENC_us20_n602, _AES_ENC_us20_n601, _AES_ENC_us20_n600, _AES_ENC_us20_n599, _AES_ENC_us20_n598, _AES_ENC_us20_n597, _AES_ENC_us20_n596, _AES_ENC_us20_n595, _AES_ENC_us20_n594, _AES_ENC_us20_n593, _AES_ENC_us20_n592, _AES_ENC_us20_n591, _AES_ENC_us20_n590, 
  _AES_ENC_us20_n589, _AES_ENC_us20_n588, _AES_ENC_us20_n587, _AES_ENC_us20_n586, _AES_ENC_us20_n585, _AES_ENC_us20_n584, _AES_ENC_us20_n583, _AES_ENC_us20_n582, _AES_ENC_us20_n581, _AES_ENC_us20_n580, _AES_ENC_us20_n579, _AES_ENC_us20_n578, _AES_ENC_us20_n577, _AES_ENC_us20_n576, _AES_ENC_us20_n575, _AES_ENC_us20_n574, _AES_ENC_us20_n573, _AES_ENC_us20_n572, _AES_ENC_us20_n571, _AES_ENC_us20_n570, _AES_ENC_us20_n569, _AES_ENC_us21_n1135, _AES_ENC_us21_n1134, _AES_ENC_us21_n1133, _AES_ENC_us21_n1132, _AES_ENC_us21_n1131, _AES_ENC_us21_n1130, _AES_ENC_us21_n1129, _AES_ENC_us21_n1128, _AES_ENC_us21_n1127, _AES_ENC_us21_n1126, _AES_ENC_us21_n1125, _AES_ENC_us21_n1124, _AES_ENC_us21_n1123, _AES_ENC_us21_n1122, _AES_ENC_us21_n1121, _AES_ENC_us21_n1120, _AES_ENC_us21_n1119, _AES_ENC_us21_n1118, _AES_ENC_us21_n1117, _AES_ENC_us21_n1116, _AES_ENC_us21_n1115, _AES_ENC_us21_n1114, _AES_ENC_us21_n1113, _AES_ENC_us21_n1112, _AES_ENC_us21_n1111, _AES_ENC_us21_n1110, _AES_ENC_us21_n1109, _AES_ENC_us21_n1108, _AES_ENC_us21_n1107, 
  _AES_ENC_us21_n1106, _AES_ENC_us21_n1105, _AES_ENC_us21_n1104, _AES_ENC_us21_n1103, _AES_ENC_us21_n1102, _AES_ENC_us21_n1101, _AES_ENC_us21_n1100, _AES_ENC_us21_n1099, _AES_ENC_us21_n1098, _AES_ENC_us21_n1097, _AES_ENC_us21_n1096, _AES_ENC_us21_n1095, _AES_ENC_us21_n1094, _AES_ENC_us21_n1093, _AES_ENC_us21_n1092, _AES_ENC_us21_n1091, _AES_ENC_us21_n1090, _AES_ENC_us21_n1089, _AES_ENC_us21_n1088, _AES_ENC_us21_n1087, _AES_ENC_us21_n1086, _AES_ENC_us21_n1085, _AES_ENC_us21_n1084, _AES_ENC_us21_n1083, _AES_ENC_us21_n1082, _AES_ENC_us21_n1081, _AES_ENC_us21_n1080, _AES_ENC_us21_n1079, _AES_ENC_us21_n1078, _AES_ENC_us21_n1077, _AES_ENC_us21_n1076, _AES_ENC_us21_n1075, _AES_ENC_us21_n1074, _AES_ENC_us21_n1073, _AES_ENC_us21_n1072, _AES_ENC_us21_n1071, _AES_ENC_us21_n1070, _AES_ENC_us21_n1069, _AES_ENC_us21_n1068, _AES_ENC_us21_n1067, _AES_ENC_us21_n1066, _AES_ENC_us21_n1065, _AES_ENC_us21_n1064, _AES_ENC_us21_n1063, _AES_ENC_us21_n1062, _AES_ENC_us21_n1061, _AES_ENC_us21_n1060, _AES_ENC_us21_n1059, _AES_ENC_us21_n1058, _AES_ENC_us21_n1057, 
  _AES_ENC_us21_n1056, _AES_ENC_us21_n1055, _AES_ENC_us21_n1054, _AES_ENC_us21_n1053, _AES_ENC_us21_n1052, _AES_ENC_us21_n1051, _AES_ENC_us21_n1050, _AES_ENC_us21_n1049, _AES_ENC_us21_n1048, _AES_ENC_us21_n1047, _AES_ENC_us21_n1046, _AES_ENC_us21_n1045, _AES_ENC_us21_n1044, _AES_ENC_us21_n1043, _AES_ENC_us21_n1042, _AES_ENC_us21_n1041, _AES_ENC_us21_n1040, _AES_ENC_us21_n1039, _AES_ENC_us21_n1038, _AES_ENC_us21_n1037, _AES_ENC_us21_n1036, _AES_ENC_us21_n1035, _AES_ENC_us21_n1034, _AES_ENC_us21_n1033, _AES_ENC_us21_n1032, _AES_ENC_us21_n1031, _AES_ENC_us21_n1030, _AES_ENC_us21_n1029, _AES_ENC_us21_n1028, _AES_ENC_us21_n1027, _AES_ENC_us21_n1026, _AES_ENC_us21_n1025, _AES_ENC_us21_n1024, _AES_ENC_us21_n1023, _AES_ENC_us21_n1022, _AES_ENC_us21_n1021, _AES_ENC_us21_n1020, _AES_ENC_us21_n1019, _AES_ENC_us21_n1018, _AES_ENC_us21_n1017, _AES_ENC_us21_n1016, _AES_ENC_us21_n1015, _AES_ENC_us21_n1014, _AES_ENC_us21_n1013, _AES_ENC_us21_n1012, _AES_ENC_us21_n1011, _AES_ENC_us21_n1010, _AES_ENC_us21_n1009, _AES_ENC_us21_n1008, _AES_ENC_us21_n1007, 
  _AES_ENC_us21_n1006, _AES_ENC_us21_n1005, _AES_ENC_us21_n1004, _AES_ENC_us21_n1003, _AES_ENC_us21_n1002, _AES_ENC_us21_n1001, _AES_ENC_us21_n1000, _AES_ENC_us21_n999, _AES_ENC_us21_n998, _AES_ENC_us21_n997, _AES_ENC_us21_n996, _AES_ENC_us21_n995, _AES_ENC_us21_n994, _AES_ENC_us21_n993, _AES_ENC_us21_n992, _AES_ENC_us21_n991, _AES_ENC_us21_n990, _AES_ENC_us21_n989, _AES_ENC_us21_n988, _AES_ENC_us21_n987, _AES_ENC_us21_n986, _AES_ENC_us21_n985, _AES_ENC_us21_n984, _AES_ENC_us21_n983, _AES_ENC_us21_n982, _AES_ENC_us21_n981, _AES_ENC_us21_n980, _AES_ENC_us21_n979, _AES_ENC_us21_n978, _AES_ENC_us21_n977, _AES_ENC_us21_n976, _AES_ENC_us21_n975, _AES_ENC_us21_n974, _AES_ENC_us21_n973, _AES_ENC_us21_n972, _AES_ENC_us21_n971, _AES_ENC_us21_n970, _AES_ENC_us21_n969, _AES_ENC_us21_n968, _AES_ENC_us21_n967, _AES_ENC_us21_n966, _AES_ENC_us21_n965, _AES_ENC_us21_n964, _AES_ENC_us21_n963, _AES_ENC_us21_n962, _AES_ENC_us21_n961, _AES_ENC_us21_n960, _AES_ENC_us21_n959, _AES_ENC_us21_n958, _AES_ENC_us21_n957, 
  _AES_ENC_us21_n956, _AES_ENC_us21_n955, _AES_ENC_us21_n954, _AES_ENC_us21_n953, _AES_ENC_us21_n952, _AES_ENC_us21_n951, _AES_ENC_us21_n950, _AES_ENC_us21_n949, _AES_ENC_us21_n948, _AES_ENC_us21_n947, _AES_ENC_us21_n946, _AES_ENC_us21_n945, _AES_ENC_us21_n944, _AES_ENC_us21_n943, _AES_ENC_us21_n942, _AES_ENC_us21_n941, _AES_ENC_us21_n940, _AES_ENC_us21_n939, _AES_ENC_us21_n938, _AES_ENC_us21_n937, _AES_ENC_us21_n936, _AES_ENC_us21_n935, _AES_ENC_us21_n934, _AES_ENC_us21_n933, _AES_ENC_us21_n932, _AES_ENC_us21_n931, _AES_ENC_us21_n930, _AES_ENC_us21_n929, _AES_ENC_us21_n928, _AES_ENC_us21_n927, _AES_ENC_us21_n926, _AES_ENC_us21_n925, _AES_ENC_us21_n924, _AES_ENC_us21_n923, _AES_ENC_us21_n922, _AES_ENC_us21_n921, _AES_ENC_us21_n920, _AES_ENC_us21_n919, _AES_ENC_us21_n918, _AES_ENC_us21_n917, _AES_ENC_us21_n916, _AES_ENC_us21_n915, _AES_ENC_us21_n914, _AES_ENC_us21_n913, _AES_ENC_us21_n912, _AES_ENC_us21_n911, _AES_ENC_us21_n910, _AES_ENC_us21_n909, _AES_ENC_us21_n908, _AES_ENC_us21_n907, 
  _AES_ENC_us21_n906, _AES_ENC_us21_n905, _AES_ENC_us21_n904, _AES_ENC_us21_n903, _AES_ENC_us21_n902, _AES_ENC_us21_n901, _AES_ENC_us21_n900, _AES_ENC_us21_n899, _AES_ENC_us21_n898, _AES_ENC_us21_n897, _AES_ENC_us21_n896, _AES_ENC_us21_n895, _AES_ENC_us21_n894, _AES_ENC_us21_n893, _AES_ENC_us21_n892, _AES_ENC_us21_n891, _AES_ENC_us21_n890, _AES_ENC_us21_n889, _AES_ENC_us21_n888, _AES_ENC_us21_n887, _AES_ENC_us21_n886, _AES_ENC_us21_n885, _AES_ENC_us21_n884, _AES_ENC_us21_n883, _AES_ENC_us21_n882, _AES_ENC_us21_n881, _AES_ENC_us21_n880, _AES_ENC_us21_n879, _AES_ENC_us21_n878, _AES_ENC_us21_n877, _AES_ENC_us21_n876, _AES_ENC_us21_n875, _AES_ENC_us21_n874, _AES_ENC_us21_n873, _AES_ENC_us21_n872, _AES_ENC_us21_n871, _AES_ENC_us21_n870, _AES_ENC_us21_n869, _AES_ENC_us21_n868, _AES_ENC_us21_n867, _AES_ENC_us21_n866, _AES_ENC_us21_n865, _AES_ENC_us21_n864, _AES_ENC_us21_n863, _AES_ENC_us21_n862, _AES_ENC_us21_n861, _AES_ENC_us21_n860, _AES_ENC_us21_n859, _AES_ENC_us21_n858, _AES_ENC_us21_n857, 
  _AES_ENC_us21_n856, _AES_ENC_us21_n855, _AES_ENC_us21_n854, _AES_ENC_us21_n853, _AES_ENC_us21_n852, _AES_ENC_us21_n851, _AES_ENC_us21_n850, _AES_ENC_us21_n849, _AES_ENC_us21_n848, _AES_ENC_us21_n847, _AES_ENC_us21_n846, _AES_ENC_us21_n845, _AES_ENC_us21_n844, _AES_ENC_us21_n843, _AES_ENC_us21_n842, _AES_ENC_us21_n841, _AES_ENC_us21_n840, _AES_ENC_us21_n839, _AES_ENC_us21_n838, _AES_ENC_us21_n837, _AES_ENC_us21_n836, _AES_ENC_us21_n835, _AES_ENC_us21_n834, _AES_ENC_us21_n833, _AES_ENC_us21_n832, _AES_ENC_us21_n831, _AES_ENC_us21_n830, _AES_ENC_us21_n829, _AES_ENC_us21_n828, _AES_ENC_us21_n827, _AES_ENC_us21_n826, _AES_ENC_us21_n825, _AES_ENC_us21_n824, _AES_ENC_us21_n823, _AES_ENC_us21_n822, _AES_ENC_us21_n821, _AES_ENC_us21_n820, _AES_ENC_us21_n819, _AES_ENC_us21_n818, _AES_ENC_us21_n817, _AES_ENC_us21_n816, _AES_ENC_us21_n815, _AES_ENC_us21_n814, _AES_ENC_us21_n813, _AES_ENC_us21_n812, _AES_ENC_us21_n811, _AES_ENC_us21_n810, _AES_ENC_us21_n809, _AES_ENC_us21_n808, _AES_ENC_us21_n807, 
  _AES_ENC_us21_n806, _AES_ENC_us21_n805, _AES_ENC_us21_n804, _AES_ENC_us21_n803, _AES_ENC_us21_n802, _AES_ENC_us21_n801, _AES_ENC_us21_n800, _AES_ENC_us21_n799, _AES_ENC_us21_n798, _AES_ENC_us21_n797, _AES_ENC_us21_n796, _AES_ENC_us21_n795, _AES_ENC_us21_n794, _AES_ENC_us21_n793, _AES_ENC_us21_n792, _AES_ENC_us21_n791, _AES_ENC_us21_n790, _AES_ENC_us21_n789, _AES_ENC_us21_n788, _AES_ENC_us21_n787, _AES_ENC_us21_n786, _AES_ENC_us21_n785, _AES_ENC_us21_n784, _AES_ENC_us21_n783, _AES_ENC_us21_n782, _AES_ENC_us21_n781, _AES_ENC_us21_n780, _AES_ENC_us21_n779, _AES_ENC_us21_n778, _AES_ENC_us21_n777, _AES_ENC_us21_n776, _AES_ENC_us21_n775, _AES_ENC_us21_n774, _AES_ENC_us21_n773, _AES_ENC_us21_n772, _AES_ENC_us21_n771, _AES_ENC_us21_n770, _AES_ENC_us21_n769, _AES_ENC_us21_n768, _AES_ENC_us21_n767, _AES_ENC_us21_n766, _AES_ENC_us21_n765, _AES_ENC_us21_n764, _AES_ENC_us21_n763, _AES_ENC_us21_n762, _AES_ENC_us21_n761, _AES_ENC_us21_n760, _AES_ENC_us21_n759, _AES_ENC_us21_n758, _AES_ENC_us21_n757, 
  _AES_ENC_us21_n756, _AES_ENC_us21_n755, _AES_ENC_us21_n754, _AES_ENC_us21_n753, _AES_ENC_us21_n752, _AES_ENC_us21_n751, _AES_ENC_us21_n750, _AES_ENC_us21_n749, _AES_ENC_us21_n748, _AES_ENC_us21_n747, _AES_ENC_us21_n746, _AES_ENC_us21_n745, _AES_ENC_us21_n744, _AES_ENC_us21_n743, _AES_ENC_us21_n742, _AES_ENC_us21_n741, _AES_ENC_us21_n740, _AES_ENC_us21_n739, _AES_ENC_us21_n738, _AES_ENC_us21_n737, _AES_ENC_us21_n736, _AES_ENC_us21_n735, _AES_ENC_us21_n734, _AES_ENC_us21_n733, _AES_ENC_us21_n732, _AES_ENC_us21_n731, _AES_ENC_us21_n730, _AES_ENC_us21_n729, _AES_ENC_us21_n728, _AES_ENC_us21_n727, _AES_ENC_us21_n726, _AES_ENC_us21_n725, _AES_ENC_us21_n724, _AES_ENC_us21_n723, _AES_ENC_us21_n722, _AES_ENC_us21_n721, _AES_ENC_us21_n720, _AES_ENC_us21_n719, _AES_ENC_us21_n718, _AES_ENC_us21_n717, _AES_ENC_us21_n716, _AES_ENC_us21_n715, _AES_ENC_us21_n714, _AES_ENC_us21_n713, _AES_ENC_us21_n712, _AES_ENC_us21_n711, _AES_ENC_us21_n710, _AES_ENC_us21_n709, _AES_ENC_us21_n708, _AES_ENC_us21_n707, 
  _AES_ENC_us21_n706, _AES_ENC_us21_n705, _AES_ENC_us21_n704, _AES_ENC_us21_n703, _AES_ENC_us21_n702, _AES_ENC_us21_n701, _AES_ENC_us21_n700, _AES_ENC_us21_n699, _AES_ENC_us21_n698, _AES_ENC_us21_n697, _AES_ENC_us21_n696, _AES_ENC_us21_n695, _AES_ENC_us21_n694, _AES_ENC_us21_n693, _AES_ENC_us21_n692, _AES_ENC_us21_n691, _AES_ENC_us21_n690, _AES_ENC_us21_n689, _AES_ENC_us21_n688, _AES_ENC_us21_n687, _AES_ENC_us21_n686, _AES_ENC_us21_n685, _AES_ENC_us21_n684, _AES_ENC_us21_n683, _AES_ENC_us21_n682, _AES_ENC_us21_n681, _AES_ENC_us21_n680, _AES_ENC_us21_n679, _AES_ENC_us21_n678, _AES_ENC_us21_n677, _AES_ENC_us21_n676, _AES_ENC_us21_n675, _AES_ENC_us21_n674, _AES_ENC_us21_n673, _AES_ENC_us21_n672, _AES_ENC_us21_n671, _AES_ENC_us21_n670, _AES_ENC_us21_n669, _AES_ENC_us21_n668, _AES_ENC_us21_n667, _AES_ENC_us21_n666, _AES_ENC_us21_n665, _AES_ENC_us21_n664, _AES_ENC_us21_n663, _AES_ENC_us21_n662, _AES_ENC_us21_n661, _AES_ENC_us21_n660, _AES_ENC_us21_n659, _AES_ENC_us21_n658, _AES_ENC_us21_n657, 
  _AES_ENC_us21_n656, _AES_ENC_us21_n655, _AES_ENC_us21_n654, _AES_ENC_us21_n653, _AES_ENC_us21_n652, _AES_ENC_us21_n651, _AES_ENC_us21_n650, _AES_ENC_us21_n649, _AES_ENC_us21_n648, _AES_ENC_us21_n647, _AES_ENC_us21_n646, _AES_ENC_us21_n645, _AES_ENC_us21_n644, _AES_ENC_us21_n643, _AES_ENC_us21_n642, _AES_ENC_us21_n641, _AES_ENC_us21_n640, _AES_ENC_us21_n639, _AES_ENC_us21_n638, _AES_ENC_us21_n637, _AES_ENC_us21_n636, _AES_ENC_us21_n635, _AES_ENC_us21_n634, _AES_ENC_us21_n633, _AES_ENC_us21_n632, _AES_ENC_us21_n631, _AES_ENC_us21_n630, _AES_ENC_us21_n629, _AES_ENC_us21_n628, _AES_ENC_us21_n627, _AES_ENC_us21_n626, _AES_ENC_us21_n625, _AES_ENC_us21_n624, _AES_ENC_us21_n623, _AES_ENC_us21_n622, _AES_ENC_us21_n621, _AES_ENC_us21_n620, _AES_ENC_us21_n619, _AES_ENC_us21_n618, _AES_ENC_us21_n617, _AES_ENC_us21_n616, _AES_ENC_us21_n615, _AES_ENC_us21_n614, _AES_ENC_us21_n613, _AES_ENC_us21_n612, _AES_ENC_us21_n611, _AES_ENC_us21_n610, _AES_ENC_us21_n609, _AES_ENC_us21_n608, _AES_ENC_us21_n607, 
  _AES_ENC_us21_n606, _AES_ENC_us21_n605, _AES_ENC_us21_n604, _AES_ENC_us21_n603, _AES_ENC_us21_n602, _AES_ENC_us21_n601, _AES_ENC_us21_n600, _AES_ENC_us21_n599, _AES_ENC_us21_n598, _AES_ENC_us21_n597, _AES_ENC_us21_n596, _AES_ENC_us21_n595, _AES_ENC_us21_n594, _AES_ENC_us21_n593, _AES_ENC_us21_n592, _AES_ENC_us21_n591, _AES_ENC_us21_n590, _AES_ENC_us21_n589, _AES_ENC_us21_n588, _AES_ENC_us21_n587, _AES_ENC_us21_n586, _AES_ENC_us21_n585, _AES_ENC_us21_n584, _AES_ENC_us21_n583, _AES_ENC_us21_n582, _AES_ENC_us21_n581, _AES_ENC_us21_n580, _AES_ENC_us21_n579, _AES_ENC_us21_n578, _AES_ENC_us21_n577, _AES_ENC_us21_n576, _AES_ENC_us21_n575, _AES_ENC_us21_n574, _AES_ENC_us21_n573, _AES_ENC_us21_n572, _AES_ENC_us21_n571, _AES_ENC_us21_n570, _AES_ENC_us21_n569, _AES_ENC_us22_n1135, _AES_ENC_us22_n1134, _AES_ENC_us22_n1133, _AES_ENC_us22_n1132, _AES_ENC_us22_n1131, _AES_ENC_us22_n1130, _AES_ENC_us22_n1129, _AES_ENC_us22_n1128, _AES_ENC_us22_n1127, _AES_ENC_us22_n1126, _AES_ENC_us22_n1125, _AES_ENC_us22_n1124, 
  _AES_ENC_us22_n1123, _AES_ENC_us22_n1122, _AES_ENC_us22_n1121, _AES_ENC_us22_n1120, _AES_ENC_us22_n1119, _AES_ENC_us22_n1118, _AES_ENC_us22_n1117, _AES_ENC_us22_n1116, _AES_ENC_us22_n1115, _AES_ENC_us22_n1114, _AES_ENC_us22_n1113, _AES_ENC_us22_n1112, _AES_ENC_us22_n1111, _AES_ENC_us22_n1110, _AES_ENC_us22_n1109, _AES_ENC_us22_n1108, _AES_ENC_us22_n1107, _AES_ENC_us22_n1106, _AES_ENC_us22_n1105, _AES_ENC_us22_n1104, _AES_ENC_us22_n1103, _AES_ENC_us22_n1102, _AES_ENC_us22_n1101, _AES_ENC_us22_n1100, _AES_ENC_us22_n1099, _AES_ENC_us22_n1098, _AES_ENC_us22_n1097, _AES_ENC_us22_n1096, _AES_ENC_us22_n1095, _AES_ENC_us22_n1094, _AES_ENC_us22_n1093, _AES_ENC_us22_n1092, _AES_ENC_us22_n1091, _AES_ENC_us22_n1090, _AES_ENC_us22_n1089, _AES_ENC_us22_n1088, _AES_ENC_us22_n1087, _AES_ENC_us22_n1086, _AES_ENC_us22_n1085, _AES_ENC_us22_n1084, _AES_ENC_us22_n1083, _AES_ENC_us22_n1082, _AES_ENC_us22_n1081, _AES_ENC_us22_n1080, _AES_ENC_us22_n1079, _AES_ENC_us22_n1078, _AES_ENC_us22_n1077, _AES_ENC_us22_n1076, _AES_ENC_us22_n1075, _AES_ENC_us22_n1074, 
  _AES_ENC_us22_n1073, _AES_ENC_us22_n1072, _AES_ENC_us22_n1071, _AES_ENC_us22_n1070, _AES_ENC_us22_n1069, _AES_ENC_us22_n1068, _AES_ENC_us22_n1067, _AES_ENC_us22_n1066, _AES_ENC_us22_n1065, _AES_ENC_us22_n1064, _AES_ENC_us22_n1063, _AES_ENC_us22_n1062, _AES_ENC_us22_n1061, _AES_ENC_us22_n1060, _AES_ENC_us22_n1059, _AES_ENC_us22_n1058, _AES_ENC_us22_n1057, _AES_ENC_us22_n1056, _AES_ENC_us22_n1055, _AES_ENC_us22_n1054, _AES_ENC_us22_n1053, _AES_ENC_us22_n1052, _AES_ENC_us22_n1051, _AES_ENC_us22_n1050, _AES_ENC_us22_n1049, _AES_ENC_us22_n1048, _AES_ENC_us22_n1047, _AES_ENC_us22_n1046, _AES_ENC_us22_n1045, _AES_ENC_us22_n1044, _AES_ENC_us22_n1043, _AES_ENC_us22_n1042, _AES_ENC_us22_n1041, _AES_ENC_us22_n1040, _AES_ENC_us22_n1039, _AES_ENC_us22_n1038, _AES_ENC_us22_n1037, _AES_ENC_us22_n1036, _AES_ENC_us22_n1035, _AES_ENC_us22_n1034, _AES_ENC_us22_n1033, _AES_ENC_us22_n1032, _AES_ENC_us22_n1031, _AES_ENC_us22_n1030, _AES_ENC_us22_n1029, _AES_ENC_us22_n1028, _AES_ENC_us22_n1027, _AES_ENC_us22_n1026, _AES_ENC_us22_n1025, _AES_ENC_us22_n1024, 
  _AES_ENC_us22_n1023, _AES_ENC_us22_n1022, _AES_ENC_us22_n1021, _AES_ENC_us22_n1020, _AES_ENC_us22_n1019, _AES_ENC_us22_n1018, _AES_ENC_us22_n1017, _AES_ENC_us22_n1016, _AES_ENC_us22_n1015, _AES_ENC_us22_n1014, _AES_ENC_us22_n1013, _AES_ENC_us22_n1012, _AES_ENC_us22_n1011, _AES_ENC_us22_n1010, _AES_ENC_us22_n1009, _AES_ENC_us22_n1008, _AES_ENC_us22_n1007, _AES_ENC_us22_n1006, _AES_ENC_us22_n1005, _AES_ENC_us22_n1004, _AES_ENC_us22_n1003, _AES_ENC_us22_n1002, _AES_ENC_us22_n1001, _AES_ENC_us22_n1000, _AES_ENC_us22_n999, _AES_ENC_us22_n998, _AES_ENC_us22_n997, _AES_ENC_us22_n996, _AES_ENC_us22_n995, _AES_ENC_us22_n994, _AES_ENC_us22_n993, _AES_ENC_us22_n992, _AES_ENC_us22_n991, _AES_ENC_us22_n990, _AES_ENC_us22_n989, _AES_ENC_us22_n988, _AES_ENC_us22_n987, _AES_ENC_us22_n986, _AES_ENC_us22_n985, _AES_ENC_us22_n984, _AES_ENC_us22_n983, _AES_ENC_us22_n982, _AES_ENC_us22_n981, _AES_ENC_us22_n980, _AES_ENC_us22_n979, _AES_ENC_us22_n978, _AES_ENC_us22_n977, _AES_ENC_us22_n976, _AES_ENC_us22_n975, _AES_ENC_us22_n974, 
  _AES_ENC_us22_n973, _AES_ENC_us22_n972, _AES_ENC_us22_n971, _AES_ENC_us22_n970, _AES_ENC_us22_n969, _AES_ENC_us22_n968, _AES_ENC_us22_n967, _AES_ENC_us22_n966, _AES_ENC_us22_n965, _AES_ENC_us22_n964, _AES_ENC_us22_n963, _AES_ENC_us22_n962, _AES_ENC_us22_n961, _AES_ENC_us22_n960, _AES_ENC_us22_n959, _AES_ENC_us22_n958, _AES_ENC_us22_n957, _AES_ENC_us22_n956, _AES_ENC_us22_n955, _AES_ENC_us22_n954, _AES_ENC_us22_n953, _AES_ENC_us22_n952, _AES_ENC_us22_n951, _AES_ENC_us22_n950, _AES_ENC_us22_n949, _AES_ENC_us22_n948, _AES_ENC_us22_n947, _AES_ENC_us22_n946, _AES_ENC_us22_n945, _AES_ENC_us22_n944, _AES_ENC_us22_n943, _AES_ENC_us22_n942, _AES_ENC_us22_n941, _AES_ENC_us22_n940, _AES_ENC_us22_n939, _AES_ENC_us22_n938, _AES_ENC_us22_n937, _AES_ENC_us22_n936, _AES_ENC_us22_n935, _AES_ENC_us22_n934, _AES_ENC_us22_n933, _AES_ENC_us22_n932, _AES_ENC_us22_n931, _AES_ENC_us22_n930, _AES_ENC_us22_n929, _AES_ENC_us22_n928, _AES_ENC_us22_n927, _AES_ENC_us22_n926, _AES_ENC_us22_n925, _AES_ENC_us22_n924, 
  _AES_ENC_us22_n923, _AES_ENC_us22_n922, _AES_ENC_us22_n921, _AES_ENC_us22_n920, _AES_ENC_us22_n919, _AES_ENC_us22_n918, _AES_ENC_us22_n917, _AES_ENC_us22_n916, _AES_ENC_us22_n915, _AES_ENC_us22_n914, _AES_ENC_us22_n913, _AES_ENC_us22_n912, _AES_ENC_us22_n911, _AES_ENC_us22_n910, _AES_ENC_us22_n909, _AES_ENC_us22_n908, _AES_ENC_us22_n907, _AES_ENC_us22_n906, _AES_ENC_us22_n905, _AES_ENC_us22_n904, _AES_ENC_us22_n903, _AES_ENC_us22_n902, _AES_ENC_us22_n901, _AES_ENC_us22_n900, _AES_ENC_us22_n899, _AES_ENC_us22_n898, _AES_ENC_us22_n897, _AES_ENC_us22_n896, _AES_ENC_us22_n895, _AES_ENC_us22_n894, _AES_ENC_us22_n893, _AES_ENC_us22_n892, _AES_ENC_us22_n891, _AES_ENC_us22_n890, _AES_ENC_us22_n889, _AES_ENC_us22_n888, _AES_ENC_us22_n887, _AES_ENC_us22_n886, _AES_ENC_us22_n885, _AES_ENC_us22_n884, _AES_ENC_us22_n883, _AES_ENC_us22_n882, _AES_ENC_us22_n881, _AES_ENC_us22_n880, _AES_ENC_us22_n879, _AES_ENC_us22_n878, _AES_ENC_us22_n877, _AES_ENC_us22_n876, _AES_ENC_us22_n875, _AES_ENC_us22_n874, 
  _AES_ENC_us22_n873, _AES_ENC_us22_n872, _AES_ENC_us22_n871, _AES_ENC_us22_n870, _AES_ENC_us22_n869, _AES_ENC_us22_n868, _AES_ENC_us22_n867, _AES_ENC_us22_n866, _AES_ENC_us22_n865, _AES_ENC_us22_n864, _AES_ENC_us22_n863, _AES_ENC_us22_n862, _AES_ENC_us22_n861, _AES_ENC_us22_n860, _AES_ENC_us22_n859, _AES_ENC_us22_n858, _AES_ENC_us22_n857, _AES_ENC_us22_n856, _AES_ENC_us22_n855, _AES_ENC_us22_n854, _AES_ENC_us22_n853, _AES_ENC_us22_n852, _AES_ENC_us22_n851, _AES_ENC_us22_n850, _AES_ENC_us22_n849, _AES_ENC_us22_n848, _AES_ENC_us22_n847, _AES_ENC_us22_n846, _AES_ENC_us22_n845, _AES_ENC_us22_n844, _AES_ENC_us22_n843, _AES_ENC_us22_n842, _AES_ENC_us22_n841, _AES_ENC_us22_n840, _AES_ENC_us22_n839, _AES_ENC_us22_n838, _AES_ENC_us22_n837, _AES_ENC_us22_n836, _AES_ENC_us22_n835, _AES_ENC_us22_n834, _AES_ENC_us22_n833, _AES_ENC_us22_n832, _AES_ENC_us22_n831, _AES_ENC_us22_n830, _AES_ENC_us22_n829, _AES_ENC_us22_n828, _AES_ENC_us22_n827, _AES_ENC_us22_n826, _AES_ENC_us22_n825, _AES_ENC_us22_n824, 
  _AES_ENC_us22_n823, _AES_ENC_us22_n822, _AES_ENC_us22_n821, _AES_ENC_us22_n820, _AES_ENC_us22_n819, _AES_ENC_us22_n818, _AES_ENC_us22_n817, _AES_ENC_us22_n816, _AES_ENC_us22_n815, _AES_ENC_us22_n814, _AES_ENC_us22_n813, _AES_ENC_us22_n812, _AES_ENC_us22_n811, _AES_ENC_us22_n810, _AES_ENC_us22_n809, _AES_ENC_us22_n808, _AES_ENC_us22_n807, _AES_ENC_us22_n806, _AES_ENC_us22_n805, _AES_ENC_us22_n804, _AES_ENC_us22_n803, _AES_ENC_us22_n802, _AES_ENC_us22_n801, _AES_ENC_us22_n800, _AES_ENC_us22_n799, _AES_ENC_us22_n798, _AES_ENC_us22_n797, _AES_ENC_us22_n796, _AES_ENC_us22_n795, _AES_ENC_us22_n794, _AES_ENC_us22_n793, _AES_ENC_us22_n792, _AES_ENC_us22_n791, _AES_ENC_us22_n790, _AES_ENC_us22_n789, _AES_ENC_us22_n788, _AES_ENC_us22_n787, _AES_ENC_us22_n786, _AES_ENC_us22_n785, _AES_ENC_us22_n784, _AES_ENC_us22_n783, _AES_ENC_us22_n782, _AES_ENC_us22_n781, _AES_ENC_us22_n780, _AES_ENC_us22_n779, _AES_ENC_us22_n778, _AES_ENC_us22_n777, _AES_ENC_us22_n776, _AES_ENC_us22_n775, _AES_ENC_us22_n774, 
  _AES_ENC_us22_n773, _AES_ENC_us22_n772, _AES_ENC_us22_n771, _AES_ENC_us22_n770, _AES_ENC_us22_n769, _AES_ENC_us22_n768, _AES_ENC_us22_n767, _AES_ENC_us22_n766, _AES_ENC_us22_n765, _AES_ENC_us22_n764, _AES_ENC_us22_n763, _AES_ENC_us22_n762, _AES_ENC_us22_n761, _AES_ENC_us22_n760, _AES_ENC_us22_n759, _AES_ENC_us22_n758, _AES_ENC_us22_n757, _AES_ENC_us22_n756, _AES_ENC_us22_n755, _AES_ENC_us22_n754, _AES_ENC_us22_n753, _AES_ENC_us22_n752, _AES_ENC_us22_n751, _AES_ENC_us22_n750, _AES_ENC_us22_n749, _AES_ENC_us22_n748, _AES_ENC_us22_n747, _AES_ENC_us22_n746, _AES_ENC_us22_n745, _AES_ENC_us22_n744, _AES_ENC_us22_n743, _AES_ENC_us22_n742, _AES_ENC_us22_n741, _AES_ENC_us22_n740, _AES_ENC_us22_n739, _AES_ENC_us22_n738, _AES_ENC_us22_n737, _AES_ENC_us22_n736, _AES_ENC_us22_n735, _AES_ENC_us22_n734, _AES_ENC_us22_n733, _AES_ENC_us22_n732, _AES_ENC_us22_n731, _AES_ENC_us22_n730, _AES_ENC_us22_n729, _AES_ENC_us22_n728, _AES_ENC_us22_n727, _AES_ENC_us22_n726, _AES_ENC_us22_n725, _AES_ENC_us22_n724, 
  _AES_ENC_us22_n723, _AES_ENC_us22_n722, _AES_ENC_us22_n721, _AES_ENC_us22_n720, _AES_ENC_us22_n719, _AES_ENC_us22_n718, _AES_ENC_us22_n717, _AES_ENC_us22_n716, _AES_ENC_us22_n715, _AES_ENC_us22_n714, _AES_ENC_us22_n713, _AES_ENC_us22_n712, _AES_ENC_us22_n711, _AES_ENC_us22_n710, _AES_ENC_us22_n709, _AES_ENC_us22_n708, _AES_ENC_us22_n707, _AES_ENC_us22_n706, _AES_ENC_us22_n705, _AES_ENC_us22_n704, _AES_ENC_us22_n703, _AES_ENC_us22_n702, _AES_ENC_us22_n701, _AES_ENC_us22_n700, _AES_ENC_us22_n699, _AES_ENC_us22_n698, _AES_ENC_us22_n697, _AES_ENC_us22_n696, _AES_ENC_us22_n695, _AES_ENC_us22_n694, _AES_ENC_us22_n693, _AES_ENC_us22_n692, _AES_ENC_us22_n691, _AES_ENC_us22_n690, _AES_ENC_us22_n689, _AES_ENC_us22_n688, _AES_ENC_us22_n687, _AES_ENC_us22_n686, _AES_ENC_us22_n685, _AES_ENC_us22_n684, _AES_ENC_us22_n683, _AES_ENC_us22_n682, _AES_ENC_us22_n681, _AES_ENC_us22_n680, _AES_ENC_us22_n679, _AES_ENC_us22_n678, _AES_ENC_us22_n677, _AES_ENC_us22_n676, _AES_ENC_us22_n675, _AES_ENC_us22_n674, 
  _AES_ENC_us22_n673, _AES_ENC_us22_n672, _AES_ENC_us22_n671, _AES_ENC_us22_n670, _AES_ENC_us22_n669, _AES_ENC_us22_n668, _AES_ENC_us22_n667, _AES_ENC_us22_n666, _AES_ENC_us22_n665, _AES_ENC_us22_n664, _AES_ENC_us22_n663, _AES_ENC_us22_n662, _AES_ENC_us22_n661, _AES_ENC_us22_n660, _AES_ENC_us22_n659, _AES_ENC_us22_n658, _AES_ENC_us22_n657, _AES_ENC_us22_n656, _AES_ENC_us22_n655, _AES_ENC_us22_n654, _AES_ENC_us22_n653, _AES_ENC_us22_n652, _AES_ENC_us22_n651, _AES_ENC_us22_n650, _AES_ENC_us22_n649, _AES_ENC_us22_n648, _AES_ENC_us22_n647, _AES_ENC_us22_n646, _AES_ENC_us22_n645, _AES_ENC_us22_n644, _AES_ENC_us22_n643, _AES_ENC_us22_n642, _AES_ENC_us22_n641, _AES_ENC_us22_n640, _AES_ENC_us22_n639, _AES_ENC_us22_n638, _AES_ENC_us22_n637, _AES_ENC_us22_n636, _AES_ENC_us22_n635, _AES_ENC_us22_n634, _AES_ENC_us22_n633, _AES_ENC_us22_n632, _AES_ENC_us22_n631, _AES_ENC_us22_n630, _AES_ENC_us22_n629, _AES_ENC_us22_n628, _AES_ENC_us22_n627, _AES_ENC_us22_n626, _AES_ENC_us22_n625, _AES_ENC_us22_n624, 
  _AES_ENC_us22_n623, _AES_ENC_us22_n622, _AES_ENC_us22_n621, _AES_ENC_us22_n620, _AES_ENC_us22_n619, _AES_ENC_us22_n618, _AES_ENC_us22_n617, _AES_ENC_us22_n616, _AES_ENC_us22_n615, _AES_ENC_us22_n614, _AES_ENC_us22_n613, _AES_ENC_us22_n612, _AES_ENC_us22_n611, _AES_ENC_us22_n610, _AES_ENC_us22_n609, _AES_ENC_us22_n608, _AES_ENC_us22_n607, _AES_ENC_us22_n606, _AES_ENC_us22_n605, _AES_ENC_us22_n604, _AES_ENC_us22_n603, _AES_ENC_us22_n602, _AES_ENC_us22_n601, _AES_ENC_us22_n600, _AES_ENC_us22_n599, _AES_ENC_us22_n598, _AES_ENC_us22_n597, _AES_ENC_us22_n596, _AES_ENC_us22_n595, _AES_ENC_us22_n594, _AES_ENC_us22_n593, _AES_ENC_us22_n592, _AES_ENC_us22_n591, _AES_ENC_us22_n590, _AES_ENC_us22_n589, _AES_ENC_us22_n588, _AES_ENC_us22_n587, _AES_ENC_us22_n586, _AES_ENC_us22_n585, _AES_ENC_us22_n584, _AES_ENC_us22_n583, _AES_ENC_us22_n582, _AES_ENC_us22_n581, _AES_ENC_us22_n580, _AES_ENC_us22_n579, _AES_ENC_us22_n578, _AES_ENC_us22_n577, _AES_ENC_us22_n576, _AES_ENC_us22_n575, _AES_ENC_us22_n574, 
  _AES_ENC_us22_n573, _AES_ENC_us22_n572, _AES_ENC_us22_n571, _AES_ENC_us22_n570, _AES_ENC_us22_n569, _AES_ENC_us23_n1135, _AES_ENC_us23_n1134, _AES_ENC_us23_n1133, _AES_ENC_us23_n1132, _AES_ENC_us23_n1131, _AES_ENC_us23_n1130, _AES_ENC_us23_n1129, _AES_ENC_us23_n1128, _AES_ENC_us23_n1127, _AES_ENC_us23_n1126, _AES_ENC_us23_n1125, _AES_ENC_us23_n1124, _AES_ENC_us23_n1123, _AES_ENC_us23_n1122, _AES_ENC_us23_n1121, _AES_ENC_us23_n1120, _AES_ENC_us23_n1119, _AES_ENC_us23_n1118, _AES_ENC_us23_n1117, _AES_ENC_us23_n1116, _AES_ENC_us23_n1115, _AES_ENC_us23_n1114, _AES_ENC_us23_n1113, _AES_ENC_us23_n1112, _AES_ENC_us23_n1111, _AES_ENC_us23_n1110, _AES_ENC_us23_n1109, _AES_ENC_us23_n1108, _AES_ENC_us23_n1107, _AES_ENC_us23_n1106, _AES_ENC_us23_n1105, _AES_ENC_us23_n1104, _AES_ENC_us23_n1103, _AES_ENC_us23_n1102, _AES_ENC_us23_n1101, _AES_ENC_us23_n1100, _AES_ENC_us23_n1099, _AES_ENC_us23_n1098, _AES_ENC_us23_n1097, _AES_ENC_us23_n1096, _AES_ENC_us23_n1095, _AES_ENC_us23_n1094, _AES_ENC_us23_n1093, _AES_ENC_us23_n1092, _AES_ENC_us23_n1091, 
  _AES_ENC_us23_n1090, _AES_ENC_us23_n1089, _AES_ENC_us23_n1088, _AES_ENC_us23_n1087, _AES_ENC_us23_n1086, _AES_ENC_us23_n1085, _AES_ENC_us23_n1084, _AES_ENC_us23_n1083, _AES_ENC_us23_n1082, _AES_ENC_us23_n1081, _AES_ENC_us23_n1080, _AES_ENC_us23_n1079, _AES_ENC_us23_n1078, _AES_ENC_us23_n1077, _AES_ENC_us23_n1076, _AES_ENC_us23_n1075, _AES_ENC_us23_n1074, _AES_ENC_us23_n1073, _AES_ENC_us23_n1072, _AES_ENC_us23_n1071, _AES_ENC_us23_n1070, _AES_ENC_us23_n1069, _AES_ENC_us23_n1068, _AES_ENC_us23_n1067, _AES_ENC_us23_n1066, _AES_ENC_us23_n1065, _AES_ENC_us23_n1064, _AES_ENC_us23_n1063, _AES_ENC_us23_n1062, _AES_ENC_us23_n1061, _AES_ENC_us23_n1060, _AES_ENC_us23_n1059, _AES_ENC_us23_n1058, _AES_ENC_us23_n1057, _AES_ENC_us23_n1056, _AES_ENC_us23_n1055, _AES_ENC_us23_n1054, _AES_ENC_us23_n1053, _AES_ENC_us23_n1052, _AES_ENC_us23_n1051, _AES_ENC_us23_n1050, _AES_ENC_us23_n1049, _AES_ENC_us23_n1048, _AES_ENC_us23_n1047, _AES_ENC_us23_n1046, _AES_ENC_us23_n1045, _AES_ENC_us23_n1044, _AES_ENC_us23_n1043, _AES_ENC_us23_n1042, _AES_ENC_us23_n1041, 
  _AES_ENC_us23_n1040, _AES_ENC_us23_n1039, _AES_ENC_us23_n1038, _AES_ENC_us23_n1037, _AES_ENC_us23_n1036, _AES_ENC_us23_n1035, _AES_ENC_us23_n1034, _AES_ENC_us23_n1033, _AES_ENC_us23_n1032, _AES_ENC_us23_n1031, _AES_ENC_us23_n1030, _AES_ENC_us23_n1029, _AES_ENC_us23_n1028, _AES_ENC_us23_n1027, _AES_ENC_us23_n1026, _AES_ENC_us23_n1025, _AES_ENC_us23_n1024, _AES_ENC_us23_n1023, _AES_ENC_us23_n1022, _AES_ENC_us23_n1021, _AES_ENC_us23_n1020, _AES_ENC_us23_n1019, _AES_ENC_us23_n1018, _AES_ENC_us23_n1017, _AES_ENC_us23_n1016, _AES_ENC_us23_n1015, _AES_ENC_us23_n1014, _AES_ENC_us23_n1013, _AES_ENC_us23_n1012, _AES_ENC_us23_n1011, _AES_ENC_us23_n1010, _AES_ENC_us23_n1009, _AES_ENC_us23_n1008, _AES_ENC_us23_n1007, _AES_ENC_us23_n1006, _AES_ENC_us23_n1005, _AES_ENC_us23_n1004, _AES_ENC_us23_n1003, _AES_ENC_us23_n1002, _AES_ENC_us23_n1001, _AES_ENC_us23_n1000, _AES_ENC_us23_n999, _AES_ENC_us23_n998, _AES_ENC_us23_n997, _AES_ENC_us23_n996, _AES_ENC_us23_n995, _AES_ENC_us23_n994, _AES_ENC_us23_n993, _AES_ENC_us23_n992, _AES_ENC_us23_n991, 
  _AES_ENC_us23_n990, _AES_ENC_us23_n989, _AES_ENC_us23_n988, _AES_ENC_us23_n987, _AES_ENC_us23_n986, _AES_ENC_us23_n985, _AES_ENC_us23_n984, _AES_ENC_us23_n983, _AES_ENC_us23_n982, _AES_ENC_us23_n981, _AES_ENC_us23_n980, _AES_ENC_us23_n979, _AES_ENC_us23_n978, _AES_ENC_us23_n977, _AES_ENC_us23_n976, _AES_ENC_us23_n975, _AES_ENC_us23_n974, _AES_ENC_us23_n973, _AES_ENC_us23_n972, _AES_ENC_us23_n971, _AES_ENC_us23_n970, _AES_ENC_us23_n969, _AES_ENC_us23_n968, _AES_ENC_us23_n967, _AES_ENC_us23_n966, _AES_ENC_us23_n965, _AES_ENC_us23_n964, _AES_ENC_us23_n963, _AES_ENC_us23_n962, _AES_ENC_us23_n961, _AES_ENC_us23_n960, _AES_ENC_us23_n959, _AES_ENC_us23_n958, _AES_ENC_us23_n957, _AES_ENC_us23_n956, _AES_ENC_us23_n955, _AES_ENC_us23_n954, _AES_ENC_us23_n953, _AES_ENC_us23_n952, _AES_ENC_us23_n951, _AES_ENC_us23_n950, _AES_ENC_us23_n949, _AES_ENC_us23_n948, _AES_ENC_us23_n947, _AES_ENC_us23_n946, _AES_ENC_us23_n945, _AES_ENC_us23_n944, _AES_ENC_us23_n943, _AES_ENC_us23_n942, _AES_ENC_us23_n941, 
  _AES_ENC_us23_n940, _AES_ENC_us23_n939, _AES_ENC_us23_n938, _AES_ENC_us23_n937, _AES_ENC_us23_n936, _AES_ENC_us23_n935, _AES_ENC_us23_n934, _AES_ENC_us23_n933, _AES_ENC_us23_n932, _AES_ENC_us23_n931, _AES_ENC_us23_n930, _AES_ENC_us23_n929, _AES_ENC_us23_n928, _AES_ENC_us23_n927, _AES_ENC_us23_n926, _AES_ENC_us23_n925, _AES_ENC_us23_n924, _AES_ENC_us23_n923, _AES_ENC_us23_n922, _AES_ENC_us23_n921, _AES_ENC_us23_n920, _AES_ENC_us23_n919, _AES_ENC_us23_n918, _AES_ENC_us23_n917, _AES_ENC_us23_n916, _AES_ENC_us23_n915, _AES_ENC_us23_n914, _AES_ENC_us23_n913, _AES_ENC_us23_n912, _AES_ENC_us23_n911, _AES_ENC_us23_n910, _AES_ENC_us23_n909, _AES_ENC_us23_n908, _AES_ENC_us23_n907, _AES_ENC_us23_n906, _AES_ENC_us23_n905, _AES_ENC_us23_n904, _AES_ENC_us23_n903, _AES_ENC_us23_n902, _AES_ENC_us23_n901, _AES_ENC_us23_n900, _AES_ENC_us23_n899, _AES_ENC_us23_n898, _AES_ENC_us23_n897, _AES_ENC_us23_n896, _AES_ENC_us23_n895, _AES_ENC_us23_n894, _AES_ENC_us23_n893, _AES_ENC_us23_n892, _AES_ENC_us23_n891, 
  _AES_ENC_us23_n890, _AES_ENC_us23_n889, _AES_ENC_us23_n888, _AES_ENC_us23_n887, _AES_ENC_us23_n886, _AES_ENC_us23_n885, _AES_ENC_us23_n884, _AES_ENC_us23_n883, _AES_ENC_us23_n882, _AES_ENC_us23_n881, _AES_ENC_us23_n880, _AES_ENC_us23_n879, _AES_ENC_us23_n878, _AES_ENC_us23_n877, _AES_ENC_us23_n876, _AES_ENC_us23_n875, _AES_ENC_us23_n874, _AES_ENC_us23_n873, _AES_ENC_us23_n872, _AES_ENC_us23_n871, _AES_ENC_us23_n870, _AES_ENC_us23_n869, _AES_ENC_us23_n868, _AES_ENC_us23_n867, _AES_ENC_us23_n866, _AES_ENC_us23_n865, _AES_ENC_us23_n864, _AES_ENC_us23_n863, _AES_ENC_us23_n862, _AES_ENC_us23_n861, _AES_ENC_us23_n860, _AES_ENC_us23_n859, _AES_ENC_us23_n858, _AES_ENC_us23_n857, _AES_ENC_us23_n856, _AES_ENC_us23_n855, _AES_ENC_us23_n854, _AES_ENC_us23_n853, _AES_ENC_us23_n852, _AES_ENC_us23_n851, _AES_ENC_us23_n850, _AES_ENC_us23_n849, _AES_ENC_us23_n848, _AES_ENC_us23_n847, _AES_ENC_us23_n846, _AES_ENC_us23_n845, _AES_ENC_us23_n844, _AES_ENC_us23_n843, _AES_ENC_us23_n842, _AES_ENC_us23_n841, 
  _AES_ENC_us23_n840, _AES_ENC_us23_n839, _AES_ENC_us23_n838, _AES_ENC_us23_n837, _AES_ENC_us23_n836, _AES_ENC_us23_n835, _AES_ENC_us23_n834, _AES_ENC_us23_n833, _AES_ENC_us23_n832, _AES_ENC_us23_n831, _AES_ENC_us23_n830, _AES_ENC_us23_n829, _AES_ENC_us23_n828, _AES_ENC_us23_n827, _AES_ENC_us23_n826, _AES_ENC_us23_n825, _AES_ENC_us23_n824, _AES_ENC_us23_n823, _AES_ENC_us23_n822, _AES_ENC_us23_n821, _AES_ENC_us23_n820, _AES_ENC_us23_n819, _AES_ENC_us23_n818, _AES_ENC_us23_n817, _AES_ENC_us23_n816, _AES_ENC_us23_n815, _AES_ENC_us23_n814, _AES_ENC_us23_n813, _AES_ENC_us23_n812, _AES_ENC_us23_n811, _AES_ENC_us23_n810, _AES_ENC_us23_n809, _AES_ENC_us23_n808, _AES_ENC_us23_n807, _AES_ENC_us23_n806, _AES_ENC_us23_n805, _AES_ENC_us23_n804, _AES_ENC_us23_n803, _AES_ENC_us23_n802, _AES_ENC_us23_n801, _AES_ENC_us23_n800, _AES_ENC_us23_n799, _AES_ENC_us23_n798, _AES_ENC_us23_n797, _AES_ENC_us23_n796, _AES_ENC_us23_n795, _AES_ENC_us23_n794, _AES_ENC_us23_n793, _AES_ENC_us23_n792, _AES_ENC_us23_n791, 
  _AES_ENC_us23_n790, _AES_ENC_us23_n789, _AES_ENC_us23_n788, _AES_ENC_us23_n787, _AES_ENC_us23_n786, _AES_ENC_us23_n785, _AES_ENC_us23_n784, _AES_ENC_us23_n783, _AES_ENC_us23_n782, _AES_ENC_us23_n781, _AES_ENC_us23_n780, _AES_ENC_us23_n779, _AES_ENC_us23_n778, _AES_ENC_us23_n777, _AES_ENC_us23_n776, _AES_ENC_us23_n775, _AES_ENC_us23_n774, _AES_ENC_us23_n773, _AES_ENC_us23_n772, _AES_ENC_us23_n771, _AES_ENC_us23_n770, _AES_ENC_us23_n769, _AES_ENC_us23_n768, _AES_ENC_us23_n767, _AES_ENC_us23_n766, _AES_ENC_us23_n765, _AES_ENC_us23_n764, _AES_ENC_us23_n763, _AES_ENC_us23_n762, _AES_ENC_us23_n761, _AES_ENC_us23_n760, _AES_ENC_us23_n759, _AES_ENC_us23_n758, _AES_ENC_us23_n757, _AES_ENC_us23_n756, _AES_ENC_us23_n755, _AES_ENC_us23_n754, _AES_ENC_us23_n753, _AES_ENC_us23_n752, _AES_ENC_us23_n751, _AES_ENC_us23_n750, _AES_ENC_us23_n749, _AES_ENC_us23_n748, _AES_ENC_us23_n747, _AES_ENC_us23_n746, _AES_ENC_us23_n745, _AES_ENC_us23_n744, _AES_ENC_us23_n743, _AES_ENC_us23_n742, _AES_ENC_us23_n741, 
  _AES_ENC_us23_n740, _AES_ENC_us23_n739, _AES_ENC_us23_n738, _AES_ENC_us23_n737, _AES_ENC_us23_n736, _AES_ENC_us23_n735, _AES_ENC_us23_n734, _AES_ENC_us23_n733, _AES_ENC_us23_n732, _AES_ENC_us23_n731, _AES_ENC_us23_n730, _AES_ENC_us23_n729, _AES_ENC_us23_n728, _AES_ENC_us23_n727, _AES_ENC_us23_n726, _AES_ENC_us23_n725, _AES_ENC_us23_n724, _AES_ENC_us23_n723, _AES_ENC_us23_n722, _AES_ENC_us23_n721, _AES_ENC_us23_n720, _AES_ENC_us23_n719, _AES_ENC_us23_n718, _AES_ENC_us23_n717, _AES_ENC_us23_n716, _AES_ENC_us23_n715, _AES_ENC_us23_n714, _AES_ENC_us23_n713, _AES_ENC_us23_n712, _AES_ENC_us23_n711, _AES_ENC_us23_n710, _AES_ENC_us23_n709, _AES_ENC_us23_n708, _AES_ENC_us23_n707, _AES_ENC_us23_n706, _AES_ENC_us23_n705, _AES_ENC_us23_n704, _AES_ENC_us23_n703, _AES_ENC_us23_n702, _AES_ENC_us23_n701, _AES_ENC_us23_n700, _AES_ENC_us23_n699, _AES_ENC_us23_n698, _AES_ENC_us23_n697, _AES_ENC_us23_n696, _AES_ENC_us23_n695, _AES_ENC_us23_n694, _AES_ENC_us23_n693, _AES_ENC_us23_n692, _AES_ENC_us23_n691, 
  _AES_ENC_us23_n690, _AES_ENC_us23_n689, _AES_ENC_us23_n688, _AES_ENC_us23_n687, _AES_ENC_us23_n686, _AES_ENC_us23_n685, _AES_ENC_us23_n684, _AES_ENC_us23_n683, _AES_ENC_us23_n682, _AES_ENC_us23_n681, _AES_ENC_us23_n680, _AES_ENC_us23_n679, _AES_ENC_us23_n678, _AES_ENC_us23_n677, _AES_ENC_us23_n676, _AES_ENC_us23_n675, _AES_ENC_us23_n674, _AES_ENC_us23_n673, _AES_ENC_us23_n672, _AES_ENC_us23_n671, _AES_ENC_us23_n670, _AES_ENC_us23_n669, _AES_ENC_us23_n668, _AES_ENC_us23_n667, _AES_ENC_us23_n666, _AES_ENC_us23_n665, _AES_ENC_us23_n664, _AES_ENC_us23_n663, _AES_ENC_us23_n662, _AES_ENC_us23_n661, _AES_ENC_us23_n660, _AES_ENC_us23_n659, _AES_ENC_us23_n658, _AES_ENC_us23_n657, _AES_ENC_us23_n656, _AES_ENC_us23_n655, _AES_ENC_us23_n654, _AES_ENC_us23_n653, _AES_ENC_us23_n652, _AES_ENC_us23_n651, _AES_ENC_us23_n650, _AES_ENC_us23_n649, _AES_ENC_us23_n648, _AES_ENC_us23_n647, _AES_ENC_us23_n646, _AES_ENC_us23_n645, _AES_ENC_us23_n644, _AES_ENC_us23_n643, _AES_ENC_us23_n642, _AES_ENC_us23_n641, 
  _AES_ENC_us23_n640, _AES_ENC_us23_n639, _AES_ENC_us23_n638, _AES_ENC_us23_n637, _AES_ENC_us23_n636, _AES_ENC_us23_n635, _AES_ENC_us23_n634, _AES_ENC_us23_n633, _AES_ENC_us23_n632, _AES_ENC_us23_n631, _AES_ENC_us23_n630, _AES_ENC_us23_n629, _AES_ENC_us23_n628, _AES_ENC_us23_n627, _AES_ENC_us23_n626, _AES_ENC_us23_n625, _AES_ENC_us23_n624, _AES_ENC_us23_n623, _AES_ENC_us23_n622, _AES_ENC_us23_n621, _AES_ENC_us23_n620, _AES_ENC_us23_n619, _AES_ENC_us23_n618, _AES_ENC_us23_n617, _AES_ENC_us23_n616, _AES_ENC_us23_n615, _AES_ENC_us23_n614, _AES_ENC_us23_n613, _AES_ENC_us23_n612, _AES_ENC_us23_n611, _AES_ENC_us23_n610, _AES_ENC_us23_n609, _AES_ENC_us23_n608, _AES_ENC_us23_n607, _AES_ENC_us23_n606, _AES_ENC_us23_n605, _AES_ENC_us23_n604, _AES_ENC_us23_n603, _AES_ENC_us23_n602, _AES_ENC_us23_n601, _AES_ENC_us23_n600, _AES_ENC_us23_n599, _AES_ENC_us23_n598, _AES_ENC_us23_n597, _AES_ENC_us23_n596, _AES_ENC_us23_n595, _AES_ENC_us23_n594, _AES_ENC_us23_n593, _AES_ENC_us23_n592, _AES_ENC_us23_n591, 
  _AES_ENC_us23_n590, _AES_ENC_us23_n589, _AES_ENC_us23_n588, _AES_ENC_us23_n587, _AES_ENC_us23_n586, _AES_ENC_us23_n585, _AES_ENC_us23_n584, _AES_ENC_us23_n583, _AES_ENC_us23_n582, _AES_ENC_us23_n581, _AES_ENC_us23_n580, _AES_ENC_us23_n579, _AES_ENC_us23_n578, _AES_ENC_us23_n577, _AES_ENC_us23_n576, _AES_ENC_us23_n575, _AES_ENC_us23_n574, _AES_ENC_us23_n573, _AES_ENC_us23_n572, _AES_ENC_us23_n571, _AES_ENC_us23_n570, _AES_ENC_us23_n569, _AES_ENC_us30_n1135, _AES_ENC_us30_n1134, _AES_ENC_us30_n1133, _AES_ENC_us30_n1132, _AES_ENC_us30_n1131, _AES_ENC_us30_n1130, _AES_ENC_us30_n1129, _AES_ENC_us30_n1128, _AES_ENC_us30_n1127, _AES_ENC_us30_n1126, _AES_ENC_us30_n1125, _AES_ENC_us30_n1124, _AES_ENC_us30_n1123, _AES_ENC_us30_n1122, _AES_ENC_us30_n1121, _AES_ENC_us30_n1120, _AES_ENC_us30_n1119, _AES_ENC_us30_n1118, _AES_ENC_us30_n1117, _AES_ENC_us30_n1116, _AES_ENC_us30_n1115, _AES_ENC_us30_n1114, _AES_ENC_us30_n1113, _AES_ENC_us30_n1112, _AES_ENC_us30_n1111, _AES_ENC_us30_n1110, _AES_ENC_us30_n1109, _AES_ENC_us30_n1108, 
  _AES_ENC_us30_n1107, _AES_ENC_us30_n1106, _AES_ENC_us30_n1105, _AES_ENC_us30_n1104, _AES_ENC_us30_n1103, _AES_ENC_us30_n1102, _AES_ENC_us30_n1101, _AES_ENC_us30_n1100, _AES_ENC_us30_n1099, _AES_ENC_us30_n1098, _AES_ENC_us30_n1097, _AES_ENC_us30_n1096, _AES_ENC_us30_n1095, _AES_ENC_us30_n1094, _AES_ENC_us30_n1093, _AES_ENC_us30_n1092, _AES_ENC_us30_n1091, _AES_ENC_us30_n1090, _AES_ENC_us30_n1089, _AES_ENC_us30_n1088, _AES_ENC_us30_n1087, _AES_ENC_us30_n1086, _AES_ENC_us30_n1085, _AES_ENC_us30_n1084, _AES_ENC_us30_n1083, _AES_ENC_us30_n1082, _AES_ENC_us30_n1081, _AES_ENC_us30_n1080, _AES_ENC_us30_n1079, _AES_ENC_us30_n1078, _AES_ENC_us30_n1077, _AES_ENC_us30_n1076, _AES_ENC_us30_n1075, _AES_ENC_us30_n1074, _AES_ENC_us30_n1073, _AES_ENC_us30_n1072, _AES_ENC_us30_n1071, _AES_ENC_us30_n1070, _AES_ENC_us30_n1069, _AES_ENC_us30_n1068, _AES_ENC_us30_n1067, _AES_ENC_us30_n1066, _AES_ENC_us30_n1065, _AES_ENC_us30_n1064, _AES_ENC_us30_n1063, _AES_ENC_us30_n1062, _AES_ENC_us30_n1061, _AES_ENC_us30_n1060, _AES_ENC_us30_n1059, _AES_ENC_us30_n1058, 
  _AES_ENC_us30_n1057, _AES_ENC_us30_n1056, _AES_ENC_us30_n1055, _AES_ENC_us30_n1054, _AES_ENC_us30_n1053, _AES_ENC_us30_n1052, _AES_ENC_us30_n1051, _AES_ENC_us30_n1050, _AES_ENC_us30_n1049, _AES_ENC_us30_n1048, _AES_ENC_us30_n1047, _AES_ENC_us30_n1046, _AES_ENC_us30_n1045, _AES_ENC_us30_n1044, _AES_ENC_us30_n1043, _AES_ENC_us30_n1042, _AES_ENC_us30_n1041, _AES_ENC_us30_n1040, _AES_ENC_us30_n1039, _AES_ENC_us30_n1038, _AES_ENC_us30_n1037, _AES_ENC_us30_n1036, _AES_ENC_us30_n1035, _AES_ENC_us30_n1034, _AES_ENC_us30_n1033, _AES_ENC_us30_n1032, _AES_ENC_us30_n1031, _AES_ENC_us30_n1030, _AES_ENC_us30_n1029, _AES_ENC_us30_n1028, _AES_ENC_us30_n1027, _AES_ENC_us30_n1026, _AES_ENC_us30_n1025, _AES_ENC_us30_n1024, _AES_ENC_us30_n1023, _AES_ENC_us30_n1022, _AES_ENC_us30_n1021, _AES_ENC_us30_n1020, _AES_ENC_us30_n1019, _AES_ENC_us30_n1018, _AES_ENC_us30_n1017, _AES_ENC_us30_n1016, _AES_ENC_us30_n1015, _AES_ENC_us30_n1014, _AES_ENC_us30_n1013, _AES_ENC_us30_n1012, _AES_ENC_us30_n1011, _AES_ENC_us30_n1010, _AES_ENC_us30_n1009, _AES_ENC_us30_n1008, 
  _AES_ENC_us30_n1007, _AES_ENC_us30_n1006, _AES_ENC_us30_n1005, _AES_ENC_us30_n1004, _AES_ENC_us30_n1003, _AES_ENC_us30_n1002, _AES_ENC_us30_n1001, _AES_ENC_us30_n1000, _AES_ENC_us30_n999, _AES_ENC_us30_n998, _AES_ENC_us30_n997, _AES_ENC_us30_n996, _AES_ENC_us30_n995, _AES_ENC_us30_n994, _AES_ENC_us30_n993, _AES_ENC_us30_n992, _AES_ENC_us30_n991, _AES_ENC_us30_n990, _AES_ENC_us30_n989, _AES_ENC_us30_n988, _AES_ENC_us30_n987, _AES_ENC_us30_n986, _AES_ENC_us30_n985, _AES_ENC_us30_n984, _AES_ENC_us30_n983, _AES_ENC_us30_n982, _AES_ENC_us30_n981, _AES_ENC_us30_n980, _AES_ENC_us30_n979, _AES_ENC_us30_n978, _AES_ENC_us30_n977, _AES_ENC_us30_n976, _AES_ENC_us30_n975, _AES_ENC_us30_n974, _AES_ENC_us30_n973, _AES_ENC_us30_n972, _AES_ENC_us30_n971, _AES_ENC_us30_n970, _AES_ENC_us30_n969, _AES_ENC_us30_n968, _AES_ENC_us30_n967, _AES_ENC_us30_n966, _AES_ENC_us30_n965, _AES_ENC_us30_n964, _AES_ENC_us30_n963, _AES_ENC_us30_n962, _AES_ENC_us30_n961, _AES_ENC_us30_n960, _AES_ENC_us30_n959, _AES_ENC_us30_n958, 
  _AES_ENC_us30_n957, _AES_ENC_us30_n956, _AES_ENC_us30_n955, _AES_ENC_us30_n954, _AES_ENC_us30_n953, _AES_ENC_us30_n952, _AES_ENC_us30_n951, _AES_ENC_us30_n950, _AES_ENC_us30_n949, _AES_ENC_us30_n948, _AES_ENC_us30_n947, _AES_ENC_us30_n946, _AES_ENC_us30_n945, _AES_ENC_us30_n944, _AES_ENC_us30_n943, _AES_ENC_us30_n942, _AES_ENC_us30_n941, _AES_ENC_us30_n940, _AES_ENC_us30_n939, _AES_ENC_us30_n938, _AES_ENC_us30_n937, _AES_ENC_us30_n936, _AES_ENC_us30_n935, _AES_ENC_us30_n934, _AES_ENC_us30_n933, _AES_ENC_us30_n932, _AES_ENC_us30_n931, _AES_ENC_us30_n930, _AES_ENC_us30_n929, _AES_ENC_us30_n928, _AES_ENC_us30_n927, _AES_ENC_us30_n926, _AES_ENC_us30_n925, _AES_ENC_us30_n924, _AES_ENC_us30_n923, _AES_ENC_us30_n922, _AES_ENC_us30_n921, _AES_ENC_us30_n920, _AES_ENC_us30_n919, _AES_ENC_us30_n918, _AES_ENC_us30_n917, _AES_ENC_us30_n916, _AES_ENC_us30_n915, _AES_ENC_us30_n914, _AES_ENC_us30_n913, _AES_ENC_us30_n912, _AES_ENC_us30_n911, _AES_ENC_us30_n910, _AES_ENC_us30_n909, _AES_ENC_us30_n908, 
  _AES_ENC_us30_n907, _AES_ENC_us30_n906, _AES_ENC_us30_n905, _AES_ENC_us30_n904, _AES_ENC_us30_n903, _AES_ENC_us30_n902, _AES_ENC_us30_n901, _AES_ENC_us30_n900, _AES_ENC_us30_n899, _AES_ENC_us30_n898, _AES_ENC_us30_n897, _AES_ENC_us30_n896, _AES_ENC_us30_n895, _AES_ENC_us30_n894, _AES_ENC_us30_n893, _AES_ENC_us30_n892, _AES_ENC_us30_n891, _AES_ENC_us30_n890, _AES_ENC_us30_n889, _AES_ENC_us30_n888, _AES_ENC_us30_n887, _AES_ENC_us30_n886, _AES_ENC_us30_n885, _AES_ENC_us30_n884, _AES_ENC_us30_n883, _AES_ENC_us30_n882, _AES_ENC_us30_n881, _AES_ENC_us30_n880, _AES_ENC_us30_n879, _AES_ENC_us30_n878, _AES_ENC_us30_n877, _AES_ENC_us30_n876, _AES_ENC_us30_n875, _AES_ENC_us30_n874, _AES_ENC_us30_n873, _AES_ENC_us30_n872, _AES_ENC_us30_n871, _AES_ENC_us30_n870, _AES_ENC_us30_n869, _AES_ENC_us30_n868, _AES_ENC_us30_n867, _AES_ENC_us30_n866, _AES_ENC_us30_n865, _AES_ENC_us30_n864, _AES_ENC_us30_n863, _AES_ENC_us30_n862, _AES_ENC_us30_n861, _AES_ENC_us30_n860, _AES_ENC_us30_n859, _AES_ENC_us30_n858, 
  _AES_ENC_us30_n857, _AES_ENC_us30_n856, _AES_ENC_us30_n855, _AES_ENC_us30_n854, _AES_ENC_us30_n853, _AES_ENC_us30_n852, _AES_ENC_us30_n851, _AES_ENC_us30_n850, _AES_ENC_us30_n849, _AES_ENC_us30_n848, _AES_ENC_us30_n847, _AES_ENC_us30_n846, _AES_ENC_us30_n845, _AES_ENC_us30_n844, _AES_ENC_us30_n843, _AES_ENC_us30_n842, _AES_ENC_us30_n841, _AES_ENC_us30_n840, _AES_ENC_us30_n839, _AES_ENC_us30_n838, _AES_ENC_us30_n837, _AES_ENC_us30_n836, _AES_ENC_us30_n835, _AES_ENC_us30_n834, _AES_ENC_us30_n833, _AES_ENC_us30_n832, _AES_ENC_us30_n831, _AES_ENC_us30_n830, _AES_ENC_us30_n829, _AES_ENC_us30_n828, _AES_ENC_us30_n827, _AES_ENC_us30_n826, _AES_ENC_us30_n825, _AES_ENC_us30_n824, _AES_ENC_us30_n823, _AES_ENC_us30_n822, _AES_ENC_us30_n821, _AES_ENC_us30_n820, _AES_ENC_us30_n819, _AES_ENC_us30_n818, _AES_ENC_us30_n817, _AES_ENC_us30_n816, _AES_ENC_us30_n815, _AES_ENC_us30_n814, _AES_ENC_us30_n813, _AES_ENC_us30_n812, _AES_ENC_us30_n811, _AES_ENC_us30_n810, _AES_ENC_us30_n809, _AES_ENC_us30_n808, 
  _AES_ENC_us30_n807, _AES_ENC_us30_n806, _AES_ENC_us30_n805, _AES_ENC_us30_n804, _AES_ENC_us30_n803, _AES_ENC_us30_n802, _AES_ENC_us30_n801, _AES_ENC_us30_n800, _AES_ENC_us30_n799, _AES_ENC_us30_n798, _AES_ENC_us30_n797, _AES_ENC_us30_n796, _AES_ENC_us30_n795, _AES_ENC_us30_n794, _AES_ENC_us30_n793, _AES_ENC_us30_n792, _AES_ENC_us30_n791, _AES_ENC_us30_n790, _AES_ENC_us30_n789, _AES_ENC_us30_n788, _AES_ENC_us30_n787, _AES_ENC_us30_n786, _AES_ENC_us30_n785, _AES_ENC_us30_n784, _AES_ENC_us30_n783, _AES_ENC_us30_n782, _AES_ENC_us30_n781, _AES_ENC_us30_n780, _AES_ENC_us30_n779, _AES_ENC_us30_n778, _AES_ENC_us30_n777, _AES_ENC_us30_n776, _AES_ENC_us30_n775, _AES_ENC_us30_n774, _AES_ENC_us30_n773, _AES_ENC_us30_n772, _AES_ENC_us30_n771, _AES_ENC_us30_n770, _AES_ENC_us30_n769, _AES_ENC_us30_n768, _AES_ENC_us30_n767, _AES_ENC_us30_n766, _AES_ENC_us30_n765, _AES_ENC_us30_n764, _AES_ENC_us30_n763, _AES_ENC_us30_n762, _AES_ENC_us30_n761, _AES_ENC_us30_n760, _AES_ENC_us30_n759, _AES_ENC_us30_n758, 
  _AES_ENC_us30_n757, _AES_ENC_us30_n756, _AES_ENC_us30_n755, _AES_ENC_us30_n754, _AES_ENC_us30_n753, _AES_ENC_us30_n752, _AES_ENC_us30_n751, _AES_ENC_us30_n750, _AES_ENC_us30_n749, _AES_ENC_us30_n748, _AES_ENC_us30_n747, _AES_ENC_us30_n746, _AES_ENC_us30_n745, _AES_ENC_us30_n744, _AES_ENC_us30_n743, _AES_ENC_us30_n742, _AES_ENC_us30_n741, _AES_ENC_us30_n740, _AES_ENC_us30_n739, _AES_ENC_us30_n738, _AES_ENC_us30_n737, _AES_ENC_us30_n736, _AES_ENC_us30_n735, _AES_ENC_us30_n734, _AES_ENC_us30_n733, _AES_ENC_us30_n732, _AES_ENC_us30_n731, _AES_ENC_us30_n730, _AES_ENC_us30_n729, _AES_ENC_us30_n728, _AES_ENC_us30_n727, _AES_ENC_us30_n726, _AES_ENC_us30_n725, _AES_ENC_us30_n724, _AES_ENC_us30_n723, _AES_ENC_us30_n722, _AES_ENC_us30_n721, _AES_ENC_us30_n720, _AES_ENC_us30_n719, _AES_ENC_us30_n718, _AES_ENC_us30_n717, _AES_ENC_us30_n716, _AES_ENC_us30_n715, _AES_ENC_us30_n714, _AES_ENC_us30_n713, _AES_ENC_us30_n712, _AES_ENC_us30_n711, _AES_ENC_us30_n710, _AES_ENC_us30_n709, _AES_ENC_us30_n708, 
  _AES_ENC_us30_n707, _AES_ENC_us30_n706, _AES_ENC_us30_n705, _AES_ENC_us30_n704, _AES_ENC_us30_n703, _AES_ENC_us30_n702, _AES_ENC_us30_n701, _AES_ENC_us30_n700, _AES_ENC_us30_n699, _AES_ENC_us30_n698, _AES_ENC_us30_n697, _AES_ENC_us30_n696, _AES_ENC_us30_n695, _AES_ENC_us30_n694, _AES_ENC_us30_n693, _AES_ENC_us30_n692, _AES_ENC_us30_n691, _AES_ENC_us30_n690, _AES_ENC_us30_n689, _AES_ENC_us30_n688, _AES_ENC_us30_n687, _AES_ENC_us30_n686, _AES_ENC_us30_n685, _AES_ENC_us30_n684, _AES_ENC_us30_n683, _AES_ENC_us30_n682, _AES_ENC_us30_n681, _AES_ENC_us30_n680, _AES_ENC_us30_n679, _AES_ENC_us30_n678, _AES_ENC_us30_n677, _AES_ENC_us30_n676, _AES_ENC_us30_n675, _AES_ENC_us30_n674, _AES_ENC_us30_n673, _AES_ENC_us30_n672, _AES_ENC_us30_n671, _AES_ENC_us30_n670, _AES_ENC_us30_n669, _AES_ENC_us30_n668, _AES_ENC_us30_n667, _AES_ENC_us30_n666, _AES_ENC_us30_n665, _AES_ENC_us30_n664, _AES_ENC_us30_n663, _AES_ENC_us30_n662, _AES_ENC_us30_n661, _AES_ENC_us30_n660, _AES_ENC_us30_n659, _AES_ENC_us30_n658, 
  _AES_ENC_us30_n657, _AES_ENC_us30_n656, _AES_ENC_us30_n655, _AES_ENC_us30_n654, _AES_ENC_us30_n653, _AES_ENC_us30_n652, _AES_ENC_us30_n651, _AES_ENC_us30_n650, _AES_ENC_us30_n649, _AES_ENC_us30_n648, _AES_ENC_us30_n647, _AES_ENC_us30_n646, _AES_ENC_us30_n645, _AES_ENC_us30_n644, _AES_ENC_us30_n643, _AES_ENC_us30_n642, _AES_ENC_us30_n641, _AES_ENC_us30_n640, _AES_ENC_us30_n639, _AES_ENC_us30_n638, _AES_ENC_us30_n637, _AES_ENC_us30_n636, _AES_ENC_us30_n635, _AES_ENC_us30_n634, _AES_ENC_us30_n633, _AES_ENC_us30_n632, _AES_ENC_us30_n631, _AES_ENC_us30_n630, _AES_ENC_us30_n629, _AES_ENC_us30_n628, _AES_ENC_us30_n627, _AES_ENC_us30_n626, _AES_ENC_us30_n625, _AES_ENC_us30_n624, _AES_ENC_us30_n623, _AES_ENC_us30_n622, _AES_ENC_us30_n621, _AES_ENC_us30_n620, _AES_ENC_us30_n619, _AES_ENC_us30_n618, _AES_ENC_us30_n617, _AES_ENC_us30_n616, _AES_ENC_us30_n615, _AES_ENC_us30_n614, _AES_ENC_us30_n613, _AES_ENC_us30_n612, _AES_ENC_us30_n611, _AES_ENC_us30_n610, _AES_ENC_us30_n609, _AES_ENC_us30_n608, 
  _AES_ENC_us30_n607, _AES_ENC_us30_n606, _AES_ENC_us30_n605, _AES_ENC_us30_n604, _AES_ENC_us30_n603, _AES_ENC_us30_n602, _AES_ENC_us30_n601, _AES_ENC_us30_n600, _AES_ENC_us30_n599, _AES_ENC_us30_n598, _AES_ENC_us30_n597, _AES_ENC_us30_n596, _AES_ENC_us30_n595, _AES_ENC_us30_n594, _AES_ENC_us30_n593, _AES_ENC_us30_n592, _AES_ENC_us30_n591, _AES_ENC_us30_n590, _AES_ENC_us30_n589, _AES_ENC_us30_n588, _AES_ENC_us30_n587, _AES_ENC_us30_n586, _AES_ENC_us30_n585, _AES_ENC_us30_n584, _AES_ENC_us30_n583, _AES_ENC_us30_n582, _AES_ENC_us30_n581, _AES_ENC_us30_n580, _AES_ENC_us30_n579, _AES_ENC_us30_n578, _AES_ENC_us30_n577, _AES_ENC_us30_n576, _AES_ENC_us30_n575, _AES_ENC_us30_n574, _AES_ENC_us30_n573, _AES_ENC_us30_n572, _AES_ENC_us30_n571, _AES_ENC_us30_n570, _AES_ENC_us30_n569, _AES_ENC_us31_n1135, _AES_ENC_us31_n1134, _AES_ENC_us31_n1133, _AES_ENC_us31_n1132, _AES_ENC_us31_n1131, _AES_ENC_us31_n1130, _AES_ENC_us31_n1129, _AES_ENC_us31_n1128, _AES_ENC_us31_n1127, _AES_ENC_us31_n1126, _AES_ENC_us31_n1125, 
  _AES_ENC_us31_n1124, _AES_ENC_us31_n1123, _AES_ENC_us31_n1122, _AES_ENC_us31_n1121, _AES_ENC_us31_n1120, _AES_ENC_us31_n1119, _AES_ENC_us31_n1118, _AES_ENC_us31_n1117, _AES_ENC_us31_n1116, _AES_ENC_us31_n1115, _AES_ENC_us31_n1114, _AES_ENC_us31_n1113, _AES_ENC_us31_n1112, _AES_ENC_us31_n1111, _AES_ENC_us31_n1110, _AES_ENC_us31_n1109, _AES_ENC_us31_n1108, _AES_ENC_us31_n1107, _AES_ENC_us31_n1106, _AES_ENC_us31_n1105, _AES_ENC_us31_n1104, _AES_ENC_us31_n1103, _AES_ENC_us31_n1102, _AES_ENC_us31_n1101, _AES_ENC_us31_n1100, _AES_ENC_us31_n1099, _AES_ENC_us31_n1098, _AES_ENC_us31_n1097, _AES_ENC_us31_n1096, _AES_ENC_us31_n1095, _AES_ENC_us31_n1094, _AES_ENC_us31_n1093, _AES_ENC_us31_n1092, _AES_ENC_us31_n1091, _AES_ENC_us31_n1090, _AES_ENC_us31_n1089, _AES_ENC_us31_n1088, _AES_ENC_us31_n1087, _AES_ENC_us31_n1086, _AES_ENC_us31_n1085, _AES_ENC_us31_n1084, _AES_ENC_us31_n1083, _AES_ENC_us31_n1082, _AES_ENC_us31_n1081, _AES_ENC_us31_n1080, _AES_ENC_us31_n1079, _AES_ENC_us31_n1078, _AES_ENC_us31_n1077, _AES_ENC_us31_n1076, _AES_ENC_us31_n1075, 
  _AES_ENC_us31_n1074, _AES_ENC_us31_n1073, _AES_ENC_us31_n1072, _AES_ENC_us31_n1071, _AES_ENC_us31_n1070, _AES_ENC_us31_n1069, _AES_ENC_us31_n1068, _AES_ENC_us31_n1067, _AES_ENC_us31_n1066, _AES_ENC_us31_n1065, _AES_ENC_us31_n1064, _AES_ENC_us31_n1063, _AES_ENC_us31_n1062, _AES_ENC_us31_n1061, _AES_ENC_us31_n1060, _AES_ENC_us31_n1059, _AES_ENC_us31_n1058, _AES_ENC_us31_n1057, _AES_ENC_us31_n1056, _AES_ENC_us31_n1055, _AES_ENC_us31_n1054, _AES_ENC_us31_n1053, _AES_ENC_us31_n1052, _AES_ENC_us31_n1051, _AES_ENC_us31_n1050, _AES_ENC_us31_n1049, _AES_ENC_us31_n1048, _AES_ENC_us31_n1047, _AES_ENC_us31_n1046, _AES_ENC_us31_n1045, _AES_ENC_us31_n1044, _AES_ENC_us31_n1043, _AES_ENC_us31_n1042, _AES_ENC_us31_n1041, _AES_ENC_us31_n1040, _AES_ENC_us31_n1039, _AES_ENC_us31_n1038, _AES_ENC_us31_n1037, _AES_ENC_us31_n1036, _AES_ENC_us31_n1035, _AES_ENC_us31_n1034, _AES_ENC_us31_n1033, _AES_ENC_us31_n1032, _AES_ENC_us31_n1031, _AES_ENC_us31_n1030, _AES_ENC_us31_n1029, _AES_ENC_us31_n1028, _AES_ENC_us31_n1027, _AES_ENC_us31_n1026, _AES_ENC_us31_n1025, 
  _AES_ENC_us31_n1024, _AES_ENC_us31_n1023, _AES_ENC_us31_n1022, _AES_ENC_us31_n1021, _AES_ENC_us31_n1020, _AES_ENC_us31_n1019, _AES_ENC_us31_n1018, _AES_ENC_us31_n1017, _AES_ENC_us31_n1016, _AES_ENC_us31_n1015, _AES_ENC_us31_n1014, _AES_ENC_us31_n1013, _AES_ENC_us31_n1012, _AES_ENC_us31_n1011, _AES_ENC_us31_n1010, _AES_ENC_us31_n1009, _AES_ENC_us31_n1008, _AES_ENC_us31_n1007, _AES_ENC_us31_n1006, _AES_ENC_us31_n1005, _AES_ENC_us31_n1004, _AES_ENC_us31_n1003, _AES_ENC_us31_n1002, _AES_ENC_us31_n1001, _AES_ENC_us31_n1000, _AES_ENC_us31_n999, _AES_ENC_us31_n998, _AES_ENC_us31_n997, _AES_ENC_us31_n996, _AES_ENC_us31_n995, _AES_ENC_us31_n994, _AES_ENC_us31_n993, _AES_ENC_us31_n992, _AES_ENC_us31_n991, _AES_ENC_us31_n990, _AES_ENC_us31_n989, _AES_ENC_us31_n988, _AES_ENC_us31_n987, _AES_ENC_us31_n986, _AES_ENC_us31_n985, _AES_ENC_us31_n984, _AES_ENC_us31_n983, _AES_ENC_us31_n982, _AES_ENC_us31_n981, _AES_ENC_us31_n980, _AES_ENC_us31_n979, _AES_ENC_us31_n978, _AES_ENC_us31_n977, _AES_ENC_us31_n976, _AES_ENC_us31_n975, 
  _AES_ENC_us31_n974, _AES_ENC_us31_n973, _AES_ENC_us31_n972, _AES_ENC_us31_n971, _AES_ENC_us31_n970, _AES_ENC_us31_n969, _AES_ENC_us31_n968, _AES_ENC_us31_n967, _AES_ENC_us31_n966, _AES_ENC_us31_n965, _AES_ENC_us31_n964, _AES_ENC_us31_n963, _AES_ENC_us31_n962, _AES_ENC_us31_n961, _AES_ENC_us31_n960, _AES_ENC_us31_n959, _AES_ENC_us31_n958, _AES_ENC_us31_n957, _AES_ENC_us31_n956, _AES_ENC_us31_n955, _AES_ENC_us31_n954, _AES_ENC_us31_n953, _AES_ENC_us31_n952, _AES_ENC_us31_n951, _AES_ENC_us31_n950, _AES_ENC_us31_n949, _AES_ENC_us31_n948, _AES_ENC_us31_n947, _AES_ENC_us31_n946, _AES_ENC_us31_n945, _AES_ENC_us31_n944, _AES_ENC_us31_n943, _AES_ENC_us31_n942, _AES_ENC_us31_n941, _AES_ENC_us31_n940, _AES_ENC_us31_n939, _AES_ENC_us31_n938, _AES_ENC_us31_n937, _AES_ENC_us31_n936, _AES_ENC_us31_n935, _AES_ENC_us31_n934, _AES_ENC_us31_n933, _AES_ENC_us31_n932, _AES_ENC_us31_n931, _AES_ENC_us31_n930, _AES_ENC_us31_n929, _AES_ENC_us31_n928, _AES_ENC_us31_n927, _AES_ENC_us31_n926, _AES_ENC_us31_n925, 
  _AES_ENC_us31_n924, _AES_ENC_us31_n923, _AES_ENC_us31_n922, _AES_ENC_us31_n921, _AES_ENC_us31_n920, _AES_ENC_us31_n919, _AES_ENC_us31_n918, _AES_ENC_us31_n917, _AES_ENC_us31_n916, _AES_ENC_us31_n915, _AES_ENC_us31_n914, _AES_ENC_us31_n913, _AES_ENC_us31_n912, _AES_ENC_us31_n911, _AES_ENC_us31_n910, _AES_ENC_us31_n909, _AES_ENC_us31_n908, _AES_ENC_us31_n907, _AES_ENC_us31_n906, _AES_ENC_us31_n905, _AES_ENC_us31_n904, _AES_ENC_us31_n903, _AES_ENC_us31_n902, _AES_ENC_us31_n901, _AES_ENC_us31_n900, _AES_ENC_us31_n899, _AES_ENC_us31_n898, _AES_ENC_us31_n897, _AES_ENC_us31_n896, _AES_ENC_us31_n895, _AES_ENC_us31_n894, _AES_ENC_us31_n893, _AES_ENC_us31_n892, _AES_ENC_us31_n891, _AES_ENC_us31_n890, _AES_ENC_us31_n889, _AES_ENC_us31_n888, _AES_ENC_us31_n887, _AES_ENC_us31_n886, _AES_ENC_us31_n885, _AES_ENC_us31_n884, _AES_ENC_us31_n883, _AES_ENC_us31_n882, _AES_ENC_us31_n881, _AES_ENC_us31_n880, _AES_ENC_us31_n879, _AES_ENC_us31_n878, _AES_ENC_us31_n877, _AES_ENC_us31_n876, _AES_ENC_us31_n875, 
  _AES_ENC_us31_n874, _AES_ENC_us31_n873, _AES_ENC_us31_n872, _AES_ENC_us31_n871, _AES_ENC_us31_n870, _AES_ENC_us31_n869, _AES_ENC_us31_n868, _AES_ENC_us31_n867, _AES_ENC_us31_n866, _AES_ENC_us31_n865, _AES_ENC_us31_n864, _AES_ENC_us31_n863, _AES_ENC_us31_n862, _AES_ENC_us31_n861, _AES_ENC_us31_n860, _AES_ENC_us31_n859, _AES_ENC_us31_n858, _AES_ENC_us31_n857, _AES_ENC_us31_n856, _AES_ENC_us31_n855, _AES_ENC_us31_n854, _AES_ENC_us31_n853, _AES_ENC_us31_n852, _AES_ENC_us31_n851, _AES_ENC_us31_n850, _AES_ENC_us31_n849, _AES_ENC_us31_n848, _AES_ENC_us31_n847, _AES_ENC_us31_n846, _AES_ENC_us31_n845, _AES_ENC_us31_n844, _AES_ENC_us31_n843, _AES_ENC_us31_n842, _AES_ENC_us31_n841, _AES_ENC_us31_n840, _AES_ENC_us31_n839, _AES_ENC_us31_n838, _AES_ENC_us31_n837, _AES_ENC_us31_n836, _AES_ENC_us31_n835, _AES_ENC_us31_n834, _AES_ENC_us31_n833, _AES_ENC_us31_n832, _AES_ENC_us31_n831, _AES_ENC_us31_n830, _AES_ENC_us31_n829, _AES_ENC_us31_n828, _AES_ENC_us31_n827, _AES_ENC_us31_n826, _AES_ENC_us31_n825, 
  _AES_ENC_us31_n824, _AES_ENC_us31_n823, _AES_ENC_us31_n822, _AES_ENC_us31_n821, _AES_ENC_us31_n820, _AES_ENC_us31_n819, _AES_ENC_us31_n818, _AES_ENC_us31_n817, _AES_ENC_us31_n816, _AES_ENC_us31_n815, _AES_ENC_us31_n814, _AES_ENC_us31_n813, _AES_ENC_us31_n812, _AES_ENC_us31_n811, _AES_ENC_us31_n810, _AES_ENC_us31_n809, _AES_ENC_us31_n808, _AES_ENC_us31_n807, _AES_ENC_us31_n806, _AES_ENC_us31_n805, _AES_ENC_us31_n804, _AES_ENC_us31_n803, _AES_ENC_us31_n802, _AES_ENC_us31_n801, _AES_ENC_us31_n800, _AES_ENC_us31_n799, _AES_ENC_us31_n798, _AES_ENC_us31_n797, _AES_ENC_us31_n796, _AES_ENC_us31_n795, _AES_ENC_us31_n794, _AES_ENC_us31_n793, _AES_ENC_us31_n792, _AES_ENC_us31_n791, _AES_ENC_us31_n790, _AES_ENC_us31_n789, _AES_ENC_us31_n788, _AES_ENC_us31_n787, _AES_ENC_us31_n786, _AES_ENC_us31_n785, _AES_ENC_us31_n784, _AES_ENC_us31_n783, _AES_ENC_us31_n782, _AES_ENC_us31_n781, _AES_ENC_us31_n780, _AES_ENC_us31_n779, _AES_ENC_us31_n778, _AES_ENC_us31_n777, _AES_ENC_us31_n776, _AES_ENC_us31_n775, 
  _AES_ENC_us31_n774, _AES_ENC_us31_n773, _AES_ENC_us31_n772, _AES_ENC_us31_n771, _AES_ENC_us31_n770, _AES_ENC_us31_n769, _AES_ENC_us31_n768, _AES_ENC_us31_n767, _AES_ENC_us31_n766, _AES_ENC_us31_n765, _AES_ENC_us31_n764, _AES_ENC_us31_n763, _AES_ENC_us31_n762, _AES_ENC_us31_n761, _AES_ENC_us31_n760, _AES_ENC_us31_n759, _AES_ENC_us31_n758, _AES_ENC_us31_n757, _AES_ENC_us31_n756, _AES_ENC_us31_n755, _AES_ENC_us31_n754, _AES_ENC_us31_n753, _AES_ENC_us31_n752, _AES_ENC_us31_n751, _AES_ENC_us31_n750, _AES_ENC_us31_n749, _AES_ENC_us31_n748, _AES_ENC_us31_n747, _AES_ENC_us31_n746, _AES_ENC_us31_n745, _AES_ENC_us31_n744, _AES_ENC_us31_n743, _AES_ENC_us31_n742, _AES_ENC_us31_n741, _AES_ENC_us31_n740, _AES_ENC_us31_n739, _AES_ENC_us31_n738, _AES_ENC_us31_n737, _AES_ENC_us31_n736, _AES_ENC_us31_n735, _AES_ENC_us31_n734, _AES_ENC_us31_n733, _AES_ENC_us31_n732, _AES_ENC_us31_n731, _AES_ENC_us31_n730, _AES_ENC_us31_n729, _AES_ENC_us31_n728, _AES_ENC_us31_n727, _AES_ENC_us31_n726, _AES_ENC_us31_n725, 
  _AES_ENC_us31_n724, _AES_ENC_us31_n723, _AES_ENC_us31_n722, _AES_ENC_us31_n721, _AES_ENC_us31_n720, _AES_ENC_us31_n719, _AES_ENC_us31_n718, _AES_ENC_us31_n717, _AES_ENC_us31_n716, _AES_ENC_us31_n715, _AES_ENC_us31_n714, _AES_ENC_us31_n713, _AES_ENC_us31_n712, _AES_ENC_us31_n711, _AES_ENC_us31_n710, _AES_ENC_us31_n709, _AES_ENC_us31_n708, _AES_ENC_us31_n707, _AES_ENC_us31_n706, _AES_ENC_us31_n705, _AES_ENC_us31_n704, _AES_ENC_us31_n703, _AES_ENC_us31_n702, _AES_ENC_us31_n701, _AES_ENC_us31_n700, _AES_ENC_us31_n699, _AES_ENC_us31_n698, _AES_ENC_us31_n697, _AES_ENC_us31_n696, _AES_ENC_us31_n695, _AES_ENC_us31_n694, _AES_ENC_us31_n693, _AES_ENC_us31_n692, _AES_ENC_us31_n691, _AES_ENC_us31_n690, _AES_ENC_us31_n689, _AES_ENC_us31_n688, _AES_ENC_us31_n687, _AES_ENC_us31_n686, _AES_ENC_us31_n685, _AES_ENC_us31_n684, _AES_ENC_us31_n683, _AES_ENC_us31_n682, _AES_ENC_us31_n681, _AES_ENC_us31_n680, _AES_ENC_us31_n679, _AES_ENC_us31_n678, _AES_ENC_us31_n677, _AES_ENC_us31_n676, _AES_ENC_us31_n675, 
  _AES_ENC_us31_n674, _AES_ENC_us31_n673, _AES_ENC_us31_n672, _AES_ENC_us31_n671, _AES_ENC_us31_n670, _AES_ENC_us31_n669, _AES_ENC_us31_n668, _AES_ENC_us31_n667, _AES_ENC_us31_n666, _AES_ENC_us31_n665, _AES_ENC_us31_n664, _AES_ENC_us31_n663, _AES_ENC_us31_n662, _AES_ENC_us31_n661, _AES_ENC_us31_n660, _AES_ENC_us31_n659, _AES_ENC_us31_n658, _AES_ENC_us31_n657, _AES_ENC_us31_n656, _AES_ENC_us31_n655, _AES_ENC_us31_n654, _AES_ENC_us31_n653, _AES_ENC_us31_n652, _AES_ENC_us31_n651, _AES_ENC_us31_n650, _AES_ENC_us31_n649, _AES_ENC_us31_n648, _AES_ENC_us31_n647, _AES_ENC_us31_n646, _AES_ENC_us31_n645, _AES_ENC_us31_n644, _AES_ENC_us31_n643, _AES_ENC_us31_n642, _AES_ENC_us31_n641, _AES_ENC_us31_n640, _AES_ENC_us31_n639, _AES_ENC_us31_n638, _AES_ENC_us31_n637, _AES_ENC_us31_n636, _AES_ENC_us31_n635, _AES_ENC_us31_n634, _AES_ENC_us31_n633, _AES_ENC_us31_n632, _AES_ENC_us31_n631, _AES_ENC_us31_n630, _AES_ENC_us31_n629, _AES_ENC_us31_n628, _AES_ENC_us31_n627, _AES_ENC_us31_n626, _AES_ENC_us31_n625, 
  _AES_ENC_us31_n624, _AES_ENC_us31_n623, _AES_ENC_us31_n622, _AES_ENC_us31_n621, _AES_ENC_us31_n620, _AES_ENC_us31_n619, _AES_ENC_us31_n618, _AES_ENC_us31_n617, _AES_ENC_us31_n616, _AES_ENC_us31_n615, _AES_ENC_us31_n614, _AES_ENC_us31_n613, _AES_ENC_us31_n612, _AES_ENC_us31_n611, _AES_ENC_us31_n610, _AES_ENC_us31_n609, _AES_ENC_us31_n608, _AES_ENC_us31_n607, _AES_ENC_us31_n606, _AES_ENC_us31_n605, _AES_ENC_us31_n604, _AES_ENC_us31_n603, _AES_ENC_us31_n602, _AES_ENC_us31_n601, _AES_ENC_us31_n600, _AES_ENC_us31_n599, _AES_ENC_us31_n598, _AES_ENC_us31_n597, _AES_ENC_us31_n596, _AES_ENC_us31_n595, _AES_ENC_us31_n594, _AES_ENC_us31_n593, _AES_ENC_us31_n592, _AES_ENC_us31_n591, _AES_ENC_us31_n590, _AES_ENC_us31_n589, _AES_ENC_us31_n588, _AES_ENC_us31_n587, _AES_ENC_us31_n586, _AES_ENC_us31_n585, _AES_ENC_us31_n584, _AES_ENC_us31_n583, _AES_ENC_us31_n582, _AES_ENC_us31_n581, _AES_ENC_us31_n580, _AES_ENC_us31_n579, _AES_ENC_us31_n578, _AES_ENC_us31_n577, _AES_ENC_us31_n576, _AES_ENC_us31_n575, 
  _AES_ENC_us31_n574, _AES_ENC_us31_n573, _AES_ENC_us31_n572, _AES_ENC_us31_n571, _AES_ENC_us31_n570, _AES_ENC_us31_n569, _AES_ENC_us32_n1135, _AES_ENC_us32_n1134, _AES_ENC_us32_n1133, _AES_ENC_us32_n1132, _AES_ENC_us32_n1131, _AES_ENC_us32_n1130, _AES_ENC_us32_n1129, _AES_ENC_us32_n1128, _AES_ENC_us32_n1127, _AES_ENC_us32_n1126, _AES_ENC_us32_n1125, _AES_ENC_us32_n1124, _AES_ENC_us32_n1123, _AES_ENC_us32_n1122, _AES_ENC_us32_n1121, _AES_ENC_us32_n1120, _AES_ENC_us32_n1119, _AES_ENC_us32_n1118, _AES_ENC_us32_n1117, _AES_ENC_us32_n1116, _AES_ENC_us32_n1115, _AES_ENC_us32_n1114, _AES_ENC_us32_n1113, _AES_ENC_us32_n1112, _AES_ENC_us32_n1111, _AES_ENC_us32_n1110, _AES_ENC_us32_n1109, _AES_ENC_us32_n1108, _AES_ENC_us32_n1107, _AES_ENC_us32_n1106, _AES_ENC_us32_n1105, _AES_ENC_us32_n1104, _AES_ENC_us32_n1103, _AES_ENC_us32_n1102, _AES_ENC_us32_n1101, _AES_ENC_us32_n1100, _AES_ENC_us32_n1099, _AES_ENC_us32_n1098, _AES_ENC_us32_n1097, _AES_ENC_us32_n1096, _AES_ENC_us32_n1095, _AES_ENC_us32_n1094, _AES_ENC_us32_n1093, _AES_ENC_us32_n1092, 
  _AES_ENC_us32_n1091, _AES_ENC_us32_n1090, _AES_ENC_us32_n1089, _AES_ENC_us32_n1088, _AES_ENC_us32_n1087, _AES_ENC_us32_n1086, _AES_ENC_us32_n1085, _AES_ENC_us32_n1084, _AES_ENC_us32_n1083, _AES_ENC_us32_n1082, _AES_ENC_us32_n1081, _AES_ENC_us32_n1080, _AES_ENC_us32_n1079, _AES_ENC_us32_n1078, _AES_ENC_us32_n1077, _AES_ENC_us32_n1076, _AES_ENC_us32_n1075, _AES_ENC_us32_n1074, _AES_ENC_us32_n1073, _AES_ENC_us32_n1072, _AES_ENC_us32_n1071, _AES_ENC_us32_n1070, _AES_ENC_us32_n1069, _AES_ENC_us32_n1068, _AES_ENC_us32_n1067, _AES_ENC_us32_n1066, _AES_ENC_us32_n1065, _AES_ENC_us32_n1064, _AES_ENC_us32_n1063, _AES_ENC_us32_n1062, _AES_ENC_us32_n1061, _AES_ENC_us32_n1060, _AES_ENC_us32_n1059, _AES_ENC_us32_n1058, _AES_ENC_us32_n1057, _AES_ENC_us32_n1056, _AES_ENC_us32_n1055, _AES_ENC_us32_n1054, _AES_ENC_us32_n1053, _AES_ENC_us32_n1052, _AES_ENC_us32_n1051, _AES_ENC_us32_n1050, _AES_ENC_us32_n1049, _AES_ENC_us32_n1048, _AES_ENC_us32_n1047, _AES_ENC_us32_n1046, _AES_ENC_us32_n1045, _AES_ENC_us32_n1044, _AES_ENC_us32_n1043, _AES_ENC_us32_n1042, 
  _AES_ENC_us32_n1041, _AES_ENC_us32_n1040, _AES_ENC_us32_n1039, _AES_ENC_us32_n1038, _AES_ENC_us32_n1037, _AES_ENC_us32_n1036, _AES_ENC_us32_n1035, _AES_ENC_us32_n1034, _AES_ENC_us32_n1033, _AES_ENC_us32_n1032, _AES_ENC_us32_n1031, _AES_ENC_us32_n1030, _AES_ENC_us32_n1029, _AES_ENC_us32_n1028, _AES_ENC_us32_n1027, _AES_ENC_us32_n1026, _AES_ENC_us32_n1025, _AES_ENC_us32_n1024, _AES_ENC_us32_n1023, _AES_ENC_us32_n1022, _AES_ENC_us32_n1021, _AES_ENC_us32_n1020, _AES_ENC_us32_n1019, _AES_ENC_us32_n1018, _AES_ENC_us32_n1017, _AES_ENC_us32_n1016, _AES_ENC_us32_n1015, _AES_ENC_us32_n1014, _AES_ENC_us32_n1013, _AES_ENC_us32_n1012, _AES_ENC_us32_n1011, _AES_ENC_us32_n1010, _AES_ENC_us32_n1009, _AES_ENC_us32_n1008, _AES_ENC_us32_n1007, _AES_ENC_us32_n1006, _AES_ENC_us32_n1005, _AES_ENC_us32_n1004, _AES_ENC_us32_n1003, _AES_ENC_us32_n1002, _AES_ENC_us32_n1001, _AES_ENC_us32_n1000, _AES_ENC_us32_n999, _AES_ENC_us32_n998, _AES_ENC_us32_n997, _AES_ENC_us32_n996, _AES_ENC_us32_n995, _AES_ENC_us32_n994, _AES_ENC_us32_n993, _AES_ENC_us32_n992, 
  _AES_ENC_us32_n991, _AES_ENC_us32_n990, _AES_ENC_us32_n989, _AES_ENC_us32_n988, _AES_ENC_us32_n987, _AES_ENC_us32_n986, _AES_ENC_us32_n985, _AES_ENC_us32_n984, _AES_ENC_us32_n983, _AES_ENC_us32_n982, _AES_ENC_us32_n981, _AES_ENC_us32_n980, _AES_ENC_us32_n979, _AES_ENC_us32_n978, _AES_ENC_us32_n977, _AES_ENC_us32_n976, _AES_ENC_us32_n975, _AES_ENC_us32_n974, _AES_ENC_us32_n973, _AES_ENC_us32_n972, _AES_ENC_us32_n971, _AES_ENC_us32_n970, _AES_ENC_us32_n969, _AES_ENC_us32_n968, _AES_ENC_us32_n967, _AES_ENC_us32_n966, _AES_ENC_us32_n965, _AES_ENC_us32_n964, _AES_ENC_us32_n963, _AES_ENC_us32_n962, _AES_ENC_us32_n961, _AES_ENC_us32_n960, _AES_ENC_us32_n959, _AES_ENC_us32_n958, _AES_ENC_us32_n957, _AES_ENC_us32_n956, _AES_ENC_us32_n955, _AES_ENC_us32_n954, _AES_ENC_us32_n953, _AES_ENC_us32_n952, _AES_ENC_us32_n951, _AES_ENC_us32_n950, _AES_ENC_us32_n949, _AES_ENC_us32_n948, _AES_ENC_us32_n947, _AES_ENC_us32_n946, _AES_ENC_us32_n945, _AES_ENC_us32_n944, _AES_ENC_us32_n943, _AES_ENC_us32_n942, 
  _AES_ENC_us32_n941, _AES_ENC_us32_n940, _AES_ENC_us32_n939, _AES_ENC_us32_n938, _AES_ENC_us32_n937, _AES_ENC_us32_n936, _AES_ENC_us32_n935, _AES_ENC_us32_n934, _AES_ENC_us32_n933, _AES_ENC_us32_n932, _AES_ENC_us32_n931, _AES_ENC_us32_n930, _AES_ENC_us32_n929, _AES_ENC_us32_n928, _AES_ENC_us32_n927, _AES_ENC_us32_n926, _AES_ENC_us32_n925, _AES_ENC_us32_n924, _AES_ENC_us32_n923, _AES_ENC_us32_n922, _AES_ENC_us32_n921, _AES_ENC_us32_n920, _AES_ENC_us32_n919, _AES_ENC_us32_n918, _AES_ENC_us32_n917, _AES_ENC_us32_n916, _AES_ENC_us32_n915, _AES_ENC_us32_n914, _AES_ENC_us32_n913, _AES_ENC_us32_n912, _AES_ENC_us32_n911, _AES_ENC_us32_n910, _AES_ENC_us32_n909, _AES_ENC_us32_n908, _AES_ENC_us32_n907, _AES_ENC_us32_n906, _AES_ENC_us32_n905, _AES_ENC_us32_n904, _AES_ENC_us32_n903, _AES_ENC_us32_n902, _AES_ENC_us32_n901, _AES_ENC_us32_n900, _AES_ENC_us32_n899, _AES_ENC_us32_n898, _AES_ENC_us32_n897, _AES_ENC_us32_n896, _AES_ENC_us32_n895, _AES_ENC_us32_n894, _AES_ENC_us32_n893, _AES_ENC_us32_n892, 
  _AES_ENC_us32_n891, _AES_ENC_us32_n890, _AES_ENC_us32_n889, _AES_ENC_us32_n888, _AES_ENC_us32_n887, _AES_ENC_us32_n886, _AES_ENC_us32_n885, _AES_ENC_us32_n884, _AES_ENC_us32_n883, _AES_ENC_us32_n882, _AES_ENC_us32_n881, _AES_ENC_us32_n880, _AES_ENC_us32_n879, _AES_ENC_us32_n878, _AES_ENC_us32_n877, _AES_ENC_us32_n876, _AES_ENC_us32_n875, _AES_ENC_us32_n874, _AES_ENC_us32_n873, _AES_ENC_us32_n872, _AES_ENC_us32_n871, _AES_ENC_us32_n870, _AES_ENC_us32_n869, _AES_ENC_us32_n868, _AES_ENC_us32_n867, _AES_ENC_us32_n866, _AES_ENC_us32_n865, _AES_ENC_us32_n864, _AES_ENC_us32_n863, _AES_ENC_us32_n862, _AES_ENC_us32_n861, _AES_ENC_us32_n860, _AES_ENC_us32_n859, _AES_ENC_us32_n858, _AES_ENC_us32_n857, _AES_ENC_us32_n856, _AES_ENC_us32_n855, _AES_ENC_us32_n854, _AES_ENC_us32_n853, _AES_ENC_us32_n852, _AES_ENC_us32_n851, _AES_ENC_us32_n850, _AES_ENC_us32_n849, _AES_ENC_us32_n848, _AES_ENC_us32_n847, _AES_ENC_us32_n846, _AES_ENC_us32_n845, _AES_ENC_us32_n844, _AES_ENC_us32_n843, _AES_ENC_us32_n842, 
  _AES_ENC_us32_n841, _AES_ENC_us32_n840, _AES_ENC_us32_n839, _AES_ENC_us32_n838, _AES_ENC_us32_n837, _AES_ENC_us32_n836, _AES_ENC_us32_n835, _AES_ENC_us32_n834, _AES_ENC_us32_n833, _AES_ENC_us32_n832, _AES_ENC_us32_n831, _AES_ENC_us32_n830, _AES_ENC_us32_n829, _AES_ENC_us32_n828, _AES_ENC_us32_n827, _AES_ENC_us32_n826, _AES_ENC_us32_n825, _AES_ENC_us32_n824, _AES_ENC_us32_n823, _AES_ENC_us32_n822, _AES_ENC_us32_n821, _AES_ENC_us32_n820, _AES_ENC_us32_n819, _AES_ENC_us32_n818, _AES_ENC_us32_n817, _AES_ENC_us32_n816, _AES_ENC_us32_n815, _AES_ENC_us32_n814, _AES_ENC_us32_n813, _AES_ENC_us32_n812, _AES_ENC_us32_n811, _AES_ENC_us32_n810, _AES_ENC_us32_n809, _AES_ENC_us32_n808, _AES_ENC_us32_n807, _AES_ENC_us32_n806, _AES_ENC_us32_n805, _AES_ENC_us32_n804, _AES_ENC_us32_n803, _AES_ENC_us32_n802, _AES_ENC_us32_n801, _AES_ENC_us32_n800, _AES_ENC_us32_n799, _AES_ENC_us32_n798, _AES_ENC_us32_n797, _AES_ENC_us32_n796, _AES_ENC_us32_n795, _AES_ENC_us32_n794, _AES_ENC_us32_n793, _AES_ENC_us32_n792, 
  _AES_ENC_us32_n791, _AES_ENC_us32_n790, _AES_ENC_us32_n789, _AES_ENC_us32_n788, _AES_ENC_us32_n787, _AES_ENC_us32_n786, _AES_ENC_us32_n785, _AES_ENC_us32_n784, _AES_ENC_us32_n783, _AES_ENC_us32_n782, _AES_ENC_us32_n781, _AES_ENC_us32_n780, _AES_ENC_us32_n779, _AES_ENC_us32_n778, _AES_ENC_us32_n777, _AES_ENC_us32_n776, _AES_ENC_us32_n775, _AES_ENC_us32_n774, _AES_ENC_us32_n773, _AES_ENC_us32_n772, _AES_ENC_us32_n771, _AES_ENC_us32_n770, _AES_ENC_us32_n769, _AES_ENC_us32_n768, _AES_ENC_us32_n767, _AES_ENC_us32_n766, _AES_ENC_us32_n765, _AES_ENC_us32_n764, _AES_ENC_us32_n763, _AES_ENC_us32_n762, _AES_ENC_us32_n761, _AES_ENC_us32_n760, _AES_ENC_us32_n759, _AES_ENC_us32_n758, _AES_ENC_us32_n757, _AES_ENC_us32_n756, _AES_ENC_us32_n755, _AES_ENC_us32_n754, _AES_ENC_us32_n753, _AES_ENC_us32_n752, _AES_ENC_us32_n751, _AES_ENC_us32_n750, _AES_ENC_us32_n749, _AES_ENC_us32_n748, _AES_ENC_us32_n747, _AES_ENC_us32_n746, _AES_ENC_us32_n745, _AES_ENC_us32_n744, _AES_ENC_us32_n743, _AES_ENC_us32_n742, 
  _AES_ENC_us32_n741, _AES_ENC_us32_n740, _AES_ENC_us32_n739, _AES_ENC_us32_n738, _AES_ENC_us32_n737, _AES_ENC_us32_n736, _AES_ENC_us32_n735, _AES_ENC_us32_n734, _AES_ENC_us32_n733, _AES_ENC_us32_n732, _AES_ENC_us32_n731, _AES_ENC_us32_n730, _AES_ENC_us32_n729, _AES_ENC_us32_n728, _AES_ENC_us32_n727, _AES_ENC_us32_n726, _AES_ENC_us32_n725, _AES_ENC_us32_n724, _AES_ENC_us32_n723, _AES_ENC_us32_n722, _AES_ENC_us32_n721, _AES_ENC_us32_n720, _AES_ENC_us32_n719, _AES_ENC_us32_n718, _AES_ENC_us32_n717, _AES_ENC_us32_n716, _AES_ENC_us32_n715, _AES_ENC_us32_n714, _AES_ENC_us32_n713, _AES_ENC_us32_n712, _AES_ENC_us32_n711, _AES_ENC_us32_n710, _AES_ENC_us32_n709, _AES_ENC_us32_n708, _AES_ENC_us32_n707, _AES_ENC_us32_n706, _AES_ENC_us32_n705, _AES_ENC_us32_n704, _AES_ENC_us32_n703, _AES_ENC_us32_n702, _AES_ENC_us32_n701, _AES_ENC_us32_n700, _AES_ENC_us32_n699, _AES_ENC_us32_n698, _AES_ENC_us32_n697, _AES_ENC_us32_n696, _AES_ENC_us32_n695, _AES_ENC_us32_n694, _AES_ENC_us32_n693, _AES_ENC_us32_n692, 
  _AES_ENC_us32_n691, _AES_ENC_us32_n690, _AES_ENC_us32_n689, _AES_ENC_us32_n688, _AES_ENC_us32_n687, _AES_ENC_us32_n686, _AES_ENC_us32_n685, _AES_ENC_us32_n684, _AES_ENC_us32_n683, _AES_ENC_us32_n682, _AES_ENC_us32_n681, _AES_ENC_us32_n680, _AES_ENC_us32_n679, _AES_ENC_us32_n678, _AES_ENC_us32_n677, _AES_ENC_us32_n676, _AES_ENC_us32_n675, _AES_ENC_us32_n674, _AES_ENC_us32_n673, _AES_ENC_us32_n672, _AES_ENC_us32_n671, _AES_ENC_us32_n670, _AES_ENC_us32_n669, _AES_ENC_us32_n668, _AES_ENC_us32_n667, _AES_ENC_us32_n666, _AES_ENC_us32_n665, _AES_ENC_us32_n664, _AES_ENC_us32_n663, _AES_ENC_us32_n662, _AES_ENC_us32_n661, _AES_ENC_us32_n660, _AES_ENC_us32_n659, _AES_ENC_us32_n658, _AES_ENC_us32_n657, _AES_ENC_us32_n656, _AES_ENC_us32_n655, _AES_ENC_us32_n654, _AES_ENC_us32_n653, _AES_ENC_us32_n652, _AES_ENC_us32_n651, _AES_ENC_us32_n650, _AES_ENC_us32_n649, _AES_ENC_us32_n648, _AES_ENC_us32_n647, _AES_ENC_us32_n646, _AES_ENC_us32_n645, _AES_ENC_us32_n644, _AES_ENC_us32_n643, _AES_ENC_us32_n642, 
  _AES_ENC_us32_n641, _AES_ENC_us32_n640, _AES_ENC_us32_n639, _AES_ENC_us32_n638, _AES_ENC_us32_n637, _AES_ENC_us32_n636, _AES_ENC_us32_n635, _AES_ENC_us32_n634, _AES_ENC_us32_n633, _AES_ENC_us32_n632, _AES_ENC_us32_n631, _AES_ENC_us32_n630, _AES_ENC_us32_n629, _AES_ENC_us32_n628, _AES_ENC_us32_n627, _AES_ENC_us32_n626, _AES_ENC_us32_n625, _AES_ENC_us32_n624, _AES_ENC_us32_n623, _AES_ENC_us32_n622, _AES_ENC_us32_n621, _AES_ENC_us32_n620, _AES_ENC_us32_n619, _AES_ENC_us32_n618, _AES_ENC_us32_n617, _AES_ENC_us32_n616, _AES_ENC_us32_n615, _AES_ENC_us32_n614, _AES_ENC_us32_n613, _AES_ENC_us32_n612, _AES_ENC_us32_n611, _AES_ENC_us32_n610, _AES_ENC_us32_n609, _AES_ENC_us32_n608, _AES_ENC_us32_n607, _AES_ENC_us32_n606, _AES_ENC_us32_n605, _AES_ENC_us32_n604, _AES_ENC_us32_n603, _AES_ENC_us32_n602, _AES_ENC_us32_n601, _AES_ENC_us32_n600, _AES_ENC_us32_n599, _AES_ENC_us32_n598, _AES_ENC_us32_n597, _AES_ENC_us32_n596, _AES_ENC_us32_n595, _AES_ENC_us32_n594, _AES_ENC_us32_n593, _AES_ENC_us32_n592, 
  _AES_ENC_us32_n591, _AES_ENC_us32_n590, _AES_ENC_us32_n589, _AES_ENC_us32_n588, _AES_ENC_us32_n587, _AES_ENC_us32_n586, _AES_ENC_us32_n585, _AES_ENC_us32_n584, _AES_ENC_us32_n583, _AES_ENC_us32_n582, _AES_ENC_us32_n581, _AES_ENC_us32_n580, _AES_ENC_us32_n579, _AES_ENC_us32_n578, _AES_ENC_us32_n577, _AES_ENC_us32_n576, _AES_ENC_us32_n575, _AES_ENC_us32_n574, _AES_ENC_us32_n573, _AES_ENC_us32_n572, _AES_ENC_us32_n571, _AES_ENC_us32_n570, _AES_ENC_us32_n569, _AES_ENC_us33_n1135, _AES_ENC_us33_n1134, _AES_ENC_us33_n1133, _AES_ENC_us33_n1132, _AES_ENC_us33_n1131, _AES_ENC_us33_n1130, _AES_ENC_us33_n1129, _AES_ENC_us33_n1128, _AES_ENC_us33_n1127, _AES_ENC_us33_n1126, _AES_ENC_us33_n1125, _AES_ENC_us33_n1124, _AES_ENC_us33_n1123, _AES_ENC_us33_n1122, _AES_ENC_us33_n1121, _AES_ENC_us33_n1120, _AES_ENC_us33_n1119, _AES_ENC_us33_n1118, _AES_ENC_us33_n1117, _AES_ENC_us33_n1116, _AES_ENC_us33_n1115, _AES_ENC_us33_n1114, _AES_ENC_us33_n1113, _AES_ENC_us33_n1112, _AES_ENC_us33_n1111, _AES_ENC_us33_n1110, _AES_ENC_us33_n1109, 
  _AES_ENC_us33_n1108, _AES_ENC_us33_n1107, _AES_ENC_us33_n1106, _AES_ENC_us33_n1105, _AES_ENC_us33_n1104, _AES_ENC_us33_n1103, _AES_ENC_us33_n1102, _AES_ENC_us33_n1101, _AES_ENC_us33_n1100, _AES_ENC_us33_n1099, _AES_ENC_us33_n1098, _AES_ENC_us33_n1097, _AES_ENC_us33_n1096, _AES_ENC_us33_n1095, _AES_ENC_us33_n1094, _AES_ENC_us33_n1093, _AES_ENC_us33_n1092, _AES_ENC_us33_n1091, _AES_ENC_us33_n1090, _AES_ENC_us33_n1089, _AES_ENC_us33_n1088, _AES_ENC_us33_n1087, _AES_ENC_us33_n1086, _AES_ENC_us33_n1085, _AES_ENC_us33_n1084, _AES_ENC_us33_n1083, _AES_ENC_us33_n1082, _AES_ENC_us33_n1081, _AES_ENC_us33_n1080, _AES_ENC_us33_n1079, _AES_ENC_us33_n1078, _AES_ENC_us33_n1077, _AES_ENC_us33_n1076, _AES_ENC_us33_n1075, _AES_ENC_us33_n1074, _AES_ENC_us33_n1073, _AES_ENC_us33_n1072, _AES_ENC_us33_n1071, _AES_ENC_us33_n1070, _AES_ENC_us33_n1069, _AES_ENC_us33_n1068, _AES_ENC_us33_n1067, _AES_ENC_us33_n1066, _AES_ENC_us33_n1065, _AES_ENC_us33_n1064, _AES_ENC_us33_n1063, _AES_ENC_us33_n1062, _AES_ENC_us33_n1061, _AES_ENC_us33_n1060, _AES_ENC_us33_n1059, 
  _AES_ENC_us33_n1058, _AES_ENC_us33_n1057, _AES_ENC_us33_n1056, _AES_ENC_us33_n1055, _AES_ENC_us33_n1054, _AES_ENC_us33_n1053, _AES_ENC_us33_n1052, _AES_ENC_us33_n1051, _AES_ENC_us33_n1050, _AES_ENC_us33_n1049, _AES_ENC_us33_n1048, _AES_ENC_us33_n1047, _AES_ENC_us33_n1046, _AES_ENC_us33_n1045, _AES_ENC_us33_n1044, _AES_ENC_us33_n1043, _AES_ENC_us33_n1042, _AES_ENC_us33_n1041, _AES_ENC_us33_n1040, _AES_ENC_us33_n1039, _AES_ENC_us33_n1038, _AES_ENC_us33_n1037, _AES_ENC_us33_n1036, _AES_ENC_us33_n1035, _AES_ENC_us33_n1034, _AES_ENC_us33_n1033, _AES_ENC_us33_n1032, _AES_ENC_us33_n1031, _AES_ENC_us33_n1030, _AES_ENC_us33_n1029, _AES_ENC_us33_n1028, _AES_ENC_us33_n1027, _AES_ENC_us33_n1026, _AES_ENC_us33_n1025, _AES_ENC_us33_n1024, _AES_ENC_us33_n1023, _AES_ENC_us33_n1022, _AES_ENC_us33_n1021, _AES_ENC_us33_n1020, _AES_ENC_us33_n1019, _AES_ENC_us33_n1018, _AES_ENC_us33_n1017, _AES_ENC_us33_n1016, _AES_ENC_us33_n1015, _AES_ENC_us33_n1014, _AES_ENC_us33_n1013, _AES_ENC_us33_n1012, _AES_ENC_us33_n1011, _AES_ENC_us33_n1010, _AES_ENC_us33_n1009, 
  _AES_ENC_us33_n1008, _AES_ENC_us33_n1007, _AES_ENC_us33_n1006, _AES_ENC_us33_n1005, _AES_ENC_us33_n1004, _AES_ENC_us33_n1003, _AES_ENC_us33_n1002, _AES_ENC_us33_n1001, _AES_ENC_us33_n1000, _AES_ENC_us33_n999, _AES_ENC_us33_n998, _AES_ENC_us33_n997, _AES_ENC_us33_n996, _AES_ENC_us33_n995, _AES_ENC_us33_n994, _AES_ENC_us33_n993, _AES_ENC_us33_n992, _AES_ENC_us33_n991, _AES_ENC_us33_n990, _AES_ENC_us33_n989, _AES_ENC_us33_n988, _AES_ENC_us33_n987, _AES_ENC_us33_n986, _AES_ENC_us33_n985, _AES_ENC_us33_n984, _AES_ENC_us33_n983, _AES_ENC_us33_n982, _AES_ENC_us33_n981, _AES_ENC_us33_n980, _AES_ENC_us33_n979, _AES_ENC_us33_n978, _AES_ENC_us33_n977, _AES_ENC_us33_n976, _AES_ENC_us33_n975, _AES_ENC_us33_n974, _AES_ENC_us33_n973, _AES_ENC_us33_n972, _AES_ENC_us33_n971, _AES_ENC_us33_n970, _AES_ENC_us33_n969, _AES_ENC_us33_n968, _AES_ENC_us33_n967, _AES_ENC_us33_n966, _AES_ENC_us33_n965, _AES_ENC_us33_n964, _AES_ENC_us33_n963, _AES_ENC_us33_n962, _AES_ENC_us33_n961, _AES_ENC_us33_n960, _AES_ENC_us33_n959, 
  _AES_ENC_us33_n958, _AES_ENC_us33_n957, _AES_ENC_us33_n956, _AES_ENC_us33_n955, _AES_ENC_us33_n954, _AES_ENC_us33_n953, _AES_ENC_us33_n952, _AES_ENC_us33_n951, _AES_ENC_us33_n950, _AES_ENC_us33_n949, _AES_ENC_us33_n948, _AES_ENC_us33_n947, _AES_ENC_us33_n946, _AES_ENC_us33_n945, _AES_ENC_us33_n944, _AES_ENC_us33_n943, _AES_ENC_us33_n942, _AES_ENC_us33_n941, _AES_ENC_us33_n940, _AES_ENC_us33_n939, _AES_ENC_us33_n938, _AES_ENC_us33_n937, _AES_ENC_us33_n936, _AES_ENC_us33_n935, _AES_ENC_us33_n934, _AES_ENC_us33_n933, _AES_ENC_us33_n932, _AES_ENC_us33_n931, _AES_ENC_us33_n930, _AES_ENC_us33_n929, _AES_ENC_us33_n928, _AES_ENC_us33_n927, _AES_ENC_us33_n926, _AES_ENC_us33_n925, _AES_ENC_us33_n924, _AES_ENC_us33_n923, _AES_ENC_us33_n922, _AES_ENC_us33_n921, _AES_ENC_us33_n920, _AES_ENC_us33_n919, _AES_ENC_us33_n918, _AES_ENC_us33_n917, _AES_ENC_us33_n916, _AES_ENC_us33_n915, _AES_ENC_us33_n914, _AES_ENC_us33_n913, _AES_ENC_us33_n912, _AES_ENC_us33_n911, _AES_ENC_us33_n910, _AES_ENC_us33_n909, 
  _AES_ENC_us33_n908, _AES_ENC_us33_n907, _AES_ENC_us33_n906, _AES_ENC_us33_n905, _AES_ENC_us33_n904, _AES_ENC_us33_n903, _AES_ENC_us33_n902, _AES_ENC_us33_n901, _AES_ENC_us33_n900, _AES_ENC_us33_n899, _AES_ENC_us33_n898, _AES_ENC_us33_n897, _AES_ENC_us33_n896, _AES_ENC_us33_n895, _AES_ENC_us33_n894, _AES_ENC_us33_n893, _AES_ENC_us33_n892, _AES_ENC_us33_n891, _AES_ENC_us33_n890, _AES_ENC_us33_n889, _AES_ENC_us33_n888, _AES_ENC_us33_n887, _AES_ENC_us33_n886, _AES_ENC_us33_n885, _AES_ENC_us33_n884, _AES_ENC_us33_n883, _AES_ENC_us33_n882, _AES_ENC_us33_n881, _AES_ENC_us33_n880, _AES_ENC_us33_n879, _AES_ENC_us33_n878, _AES_ENC_us33_n877, _AES_ENC_us33_n876, _AES_ENC_us33_n875, _AES_ENC_us33_n874, _AES_ENC_us33_n873, _AES_ENC_us33_n872, _AES_ENC_us33_n871, _AES_ENC_us33_n870, _AES_ENC_us33_n869, _AES_ENC_us33_n868, _AES_ENC_us33_n867, _AES_ENC_us33_n866, _AES_ENC_us33_n865, _AES_ENC_us33_n864, _AES_ENC_us33_n863, _AES_ENC_us33_n862, _AES_ENC_us33_n861, _AES_ENC_us33_n860, _AES_ENC_us33_n859, 
  _AES_ENC_us33_n858, _AES_ENC_us33_n857, _AES_ENC_us33_n856, _AES_ENC_us33_n855, _AES_ENC_us33_n854, _AES_ENC_us33_n853, _AES_ENC_us33_n852, _AES_ENC_us33_n851, _AES_ENC_us33_n850, _AES_ENC_us33_n849, _AES_ENC_us33_n848, _AES_ENC_us33_n847, _AES_ENC_us33_n846, _AES_ENC_us33_n845, _AES_ENC_us33_n844, _AES_ENC_us33_n843, _AES_ENC_us33_n842, _AES_ENC_us33_n841, _AES_ENC_us33_n840, _AES_ENC_us33_n839, _AES_ENC_us33_n838, _AES_ENC_us33_n837, _AES_ENC_us33_n836, _AES_ENC_us33_n835, _AES_ENC_us33_n834, _AES_ENC_us33_n833, _AES_ENC_us33_n832, _AES_ENC_us33_n831, _AES_ENC_us33_n830, _AES_ENC_us33_n829, _AES_ENC_us33_n828, _AES_ENC_us33_n827, _AES_ENC_us33_n826, _AES_ENC_us33_n825, _AES_ENC_us33_n824, _AES_ENC_us33_n823, _AES_ENC_us33_n822, _AES_ENC_us33_n821, _AES_ENC_us33_n820, _AES_ENC_us33_n819, _AES_ENC_us33_n818, _AES_ENC_us33_n817, _AES_ENC_us33_n816, _AES_ENC_us33_n815, _AES_ENC_us33_n814, _AES_ENC_us33_n813, _AES_ENC_us33_n812, _AES_ENC_us33_n811, _AES_ENC_us33_n810, _AES_ENC_us33_n809, 
  _AES_ENC_us33_n808, _AES_ENC_us33_n807, _AES_ENC_us33_n806, _AES_ENC_us33_n805, _AES_ENC_us33_n804, _AES_ENC_us33_n803, _AES_ENC_us33_n802, _AES_ENC_us33_n801, _AES_ENC_us33_n800, _AES_ENC_us33_n799, _AES_ENC_us33_n798, _AES_ENC_us33_n797, _AES_ENC_us33_n796, _AES_ENC_us33_n795, _AES_ENC_us33_n794, _AES_ENC_us33_n793, _AES_ENC_us33_n792, _AES_ENC_us33_n791, _AES_ENC_us33_n790, _AES_ENC_us33_n789, _AES_ENC_us33_n788, _AES_ENC_us33_n787, _AES_ENC_us33_n786, _AES_ENC_us33_n785, _AES_ENC_us33_n784, _AES_ENC_us33_n783, _AES_ENC_us33_n782, _AES_ENC_us33_n781, _AES_ENC_us33_n780, _AES_ENC_us33_n779, _AES_ENC_us33_n778, _AES_ENC_us33_n777, _AES_ENC_us33_n776, _AES_ENC_us33_n775, _AES_ENC_us33_n774, _AES_ENC_us33_n773, _AES_ENC_us33_n772, _AES_ENC_us33_n771, _AES_ENC_us33_n770, _AES_ENC_us33_n769, _AES_ENC_us33_n768, _AES_ENC_us33_n767, _AES_ENC_us33_n766, _AES_ENC_us33_n765, _AES_ENC_us33_n764, _AES_ENC_us33_n763, _AES_ENC_us33_n762, _AES_ENC_us33_n761, _AES_ENC_us33_n760, _AES_ENC_us33_n759, 
  _AES_ENC_us33_n758, _AES_ENC_us33_n757, _AES_ENC_us33_n756, _AES_ENC_us33_n755, _AES_ENC_us33_n754, _AES_ENC_us33_n753, _AES_ENC_us33_n752, _AES_ENC_us33_n751, _AES_ENC_us33_n750, _AES_ENC_us33_n749, _AES_ENC_us33_n748, _AES_ENC_us33_n747, _AES_ENC_us33_n746, _AES_ENC_us33_n745, _AES_ENC_us33_n744, _AES_ENC_us33_n743, _AES_ENC_us33_n742, _AES_ENC_us33_n741, _AES_ENC_us33_n740, _AES_ENC_us33_n739, _AES_ENC_us33_n738, _AES_ENC_us33_n737, _AES_ENC_us33_n736, _AES_ENC_us33_n735, _AES_ENC_us33_n734, _AES_ENC_us33_n733, _AES_ENC_us33_n732, _AES_ENC_us33_n731, _AES_ENC_us33_n730, _AES_ENC_us33_n729, _AES_ENC_us33_n728, _AES_ENC_us33_n727, _AES_ENC_us33_n726, _AES_ENC_us33_n725, _AES_ENC_us33_n724, _AES_ENC_us33_n723, _AES_ENC_us33_n722, _AES_ENC_us33_n721, _AES_ENC_us33_n720, _AES_ENC_us33_n719, _AES_ENC_us33_n718, _AES_ENC_us33_n717, _AES_ENC_us33_n716, _AES_ENC_us33_n715, _AES_ENC_us33_n714, _AES_ENC_us33_n713, _AES_ENC_us33_n712, _AES_ENC_us33_n711, _AES_ENC_us33_n710, _AES_ENC_us33_n709, 
  _AES_ENC_us33_n708, _AES_ENC_us33_n707, _AES_ENC_us33_n706, _AES_ENC_us33_n705, _AES_ENC_us33_n704, _AES_ENC_us33_n703, _AES_ENC_us33_n702, _AES_ENC_us33_n701, _AES_ENC_us33_n700, _AES_ENC_us33_n699, _AES_ENC_us33_n698, _AES_ENC_us33_n697, _AES_ENC_us33_n696, _AES_ENC_us33_n695, _AES_ENC_us33_n694, _AES_ENC_us33_n693, _AES_ENC_us33_n692, _AES_ENC_us33_n691, _AES_ENC_us33_n690, _AES_ENC_us33_n689, _AES_ENC_us33_n688, _AES_ENC_us33_n687, _AES_ENC_us33_n686, _AES_ENC_us33_n685, _AES_ENC_us33_n684, _AES_ENC_us33_n683, _AES_ENC_us33_n682, _AES_ENC_us33_n681, _AES_ENC_us33_n680, _AES_ENC_us33_n679, _AES_ENC_us33_n678, _AES_ENC_us33_n677, _AES_ENC_us33_n676, _AES_ENC_us33_n675, _AES_ENC_us33_n674, _AES_ENC_us33_n673, _AES_ENC_us33_n672, _AES_ENC_us33_n671, _AES_ENC_us33_n670, _AES_ENC_us33_n669, _AES_ENC_us33_n668, _AES_ENC_us33_n667, _AES_ENC_us33_n666, _AES_ENC_us33_n665, _AES_ENC_us33_n664, _AES_ENC_us33_n663, _AES_ENC_us33_n662, _AES_ENC_us33_n661, _AES_ENC_us33_n660, _AES_ENC_us33_n659, 
  _AES_ENC_us33_n658, _AES_ENC_us33_n657, _AES_ENC_us33_n656, _AES_ENC_us33_n655, _AES_ENC_us33_n654, _AES_ENC_us33_n653, _AES_ENC_us33_n652, _AES_ENC_us33_n651, _AES_ENC_us33_n650, _AES_ENC_us33_n649, _AES_ENC_us33_n648, _AES_ENC_us33_n647, _AES_ENC_us33_n646, _AES_ENC_us33_n645, _AES_ENC_us33_n644, _AES_ENC_us33_n643, _AES_ENC_us33_n642, _AES_ENC_us33_n641, _AES_ENC_us33_n640, _AES_ENC_us33_n639, _AES_ENC_us33_n638, _AES_ENC_us33_n637, _AES_ENC_us33_n636, _AES_ENC_us33_n635, _AES_ENC_us33_n634, _AES_ENC_us33_n633, _AES_ENC_us33_n632, _AES_ENC_us33_n631, _AES_ENC_us33_n630, _AES_ENC_us33_n629, _AES_ENC_us33_n628, _AES_ENC_us33_n627, _AES_ENC_us33_n626, _AES_ENC_us33_n625, _AES_ENC_us33_n624, _AES_ENC_us33_n623, _AES_ENC_us33_n622, _AES_ENC_us33_n621, _AES_ENC_us33_n620, _AES_ENC_us33_n619, _AES_ENC_us33_n618, _AES_ENC_us33_n617, _AES_ENC_us33_n616, _AES_ENC_us33_n615, _AES_ENC_us33_n614, _AES_ENC_us33_n613, _AES_ENC_us33_n612, _AES_ENC_us33_n611, _AES_ENC_us33_n610, _AES_ENC_us33_n609, 
  _AES_ENC_us33_n608, _AES_ENC_us33_n607, _AES_ENC_us33_n606, _AES_ENC_us33_n605, _AES_ENC_us33_n604, _AES_ENC_us33_n603, _AES_ENC_us33_n602, _AES_ENC_us33_n601, _AES_ENC_us33_n600, _AES_ENC_us33_n599, _AES_ENC_us33_n598, _AES_ENC_us33_n597, _AES_ENC_us33_n596, _AES_ENC_us33_n595, _AES_ENC_us33_n594, _AES_ENC_us33_n593, _AES_ENC_us33_n592, _AES_ENC_us33_n591, _AES_ENC_us33_n590, _AES_ENC_us33_n589, _AES_ENC_us33_n588, _AES_ENC_us33_n587, _AES_ENC_us33_n586, _AES_ENC_us33_n585, _AES_ENC_us33_n584, _AES_ENC_us33_n583, _AES_ENC_us33_n582, _AES_ENC_us33_n581, _AES_ENC_us33_n580, _AES_ENC_us33_n579, _AES_ENC_us33_n578, _AES_ENC_us33_n577, _AES_ENC_us33_n576, _AES_ENC_us33_n575, _AES_ENC_us33_n574, _AES_ENC_us33_n573, _AES_ENC_us33_n572, _AES_ENC_us33_n571, _AES_ENC_us33_n570, _AES_ENC_us33_n569, _add_506_n647, _add_506_n646, _add_506_n645, _add_506_n644, _add_506_n643, _add_506_n642, _add_506_n641, _add_506_n640, _add_506_n639, _add_506_n638, 
  _add_506_n637, _add_506_n636, _add_506_n635, _add_506_n634, _add_506_n633, _add_506_n632, _add_506_n631, _add_506_n630, _add_506_n629, _add_506_n628, _add_506_n627, _add_506_n626, _add_506_n625, _add_506_n624, _add_506_n623, _add_506_n622, _add_506_n621, _add_506_n620, _add_506_n619, _add_506_n618, _add_506_n617, _add_506_n616, _add_506_n615, _add_506_n614, _add_506_n613, _add_506_n612, _add_506_n611, _add_506_n610, _add_506_n609, _add_506_n608, _add_506_n607, _add_506_n606, _add_506_n605, _add_506_n604, _add_506_n603, _add_506_n602, _add_506_n601, _add_506_n600, _add_506_n599, _add_506_n598, _add_506_n597, _add_506_n596, _add_506_n595, _add_506_n594, _add_506_n593, _add_506_n592, _add_506_n591, _add_506_n590, _add_506_n589, _add_506_n588, 
  _add_506_n587, _add_506_n586, _add_506_n585, _add_506_n584, _add_506_n583, _add_506_n582, _add_506_n581, _add_506_n580, _add_506_n579, _add_506_n578, _add_506_n577, _add_506_n576, _add_506_n575, _add_506_n574, _add_506_n573, _add_506_n572, _add_506_n571, _add_506_n570, _add_506_n569, _add_506_n568, _add_506_n567, _add_506_n566, _add_506_n565, _add_506_n564, _add_506_n563, _add_506_n562, _add_506_n561, _add_506_n560, _add_506_n559, _add_506_n558, _add_506_n557, _add_506_n556, _add_506_n555, _add_506_n554, _add_506_n553, _add_506_n552, _add_506_n551, _add_506_n550, _add_506_n549, _add_506_n548, _add_506_n547, _add_506_n546, _add_506_n545, _add_506_n544, _add_506_n543, _add_506_n542, _add_506_n541, _add_506_n540, _add_506_n539, _add_506_n538, 
  _add_506_n537, _add_506_n536, _add_506_n535, _add_506_n534, _add_506_n533, _add_506_n532, _add_506_n531, _add_506_n530, _add_506_n529, _add_506_n528, _add_506_n527, _add_506_n526, _add_506_n525, _add_506_n524, _add_506_n523, _add_506_n522, _add_506_n521, _add_506_n520, _add_506_n519, _add_506_n518, _add_506_n517, _add_506_n516, _add_506_n515, _add_506_n514, _add_506_n513, _add_506_n512, _add_506_n511, _add_506_n510, _add_506_n509, _add_506_n508, _add_506_n507, _add_506_n506, _add_506_n505, _add_506_n504, _add_506_n503, _add_506_n502, _add_506_n501, _add_506_n500, _add_506_n499, _add_506_n498, _add_506_n497, _add_506_n496, _add_506_n495, _add_506_n494, _add_506_n493, _add_506_n492, _add_506_n491, _add_506_n490, _add_506_n489, _add_506_n488, 
  _add_506_n487, _add_506_n486, _add_506_n485, _add_506_n484, _add_506_n483, _add_506_n482, _add_506_n481, _add_506_n480, _add_506_n479, _add_506_n478, _add_506_n477, _add_506_n476, _add_506_n475, _add_506_n474, _add_506_n473, _add_506_n472, _add_506_n471, _add_506_n470, _add_506_n469, _add_506_n468, _add_506_n467, _add_506_n466, _add_506_n465, _add_506_n464, _add_506_n463, _add_506_n462, _add_506_n461, _add_506_n460, _add_506_n459, _add_506_n458, _add_506_n457, _add_506_n456, _add_506_n455, _add_506_n454, _add_506_n453, _add_506_n452, _add_506_n451, _add_506_n450, _add_506_n449, _add_506_n448, _add_506_n447, _add_506_n446, _add_506_n445, _add_506_n444, _add_506_n443, _add_506_n442, _add_506_n441, _add_506_n440, _add_506_n439, _add_506_n438, 
  _add_506_n437, _add_506_n436, _add_506_n435, _add_506_n434, _add_506_n433, _add_506_n432, _add_506_n431, _add_506_n430, _add_506_n429, _add_506_n428, _add_506_n427, _add_506_n426, _add_506_n425, _add_506_n424, _add_506_n423, _add_506_n422, _add_506_n421, _add_506_n420, _add_506_n419, _add_506_n418, _add_506_n417, _add_506_n416, _add_506_n415, _add_506_n414, _add_506_n413, _add_506_n412, _add_506_n411, _add_506_n410, _add_506_n409, _add_506_n408, _add_506_n407, _add_506_n406, _add_506_n405, _add_506_n404, _add_506_n403, _add_506_n402, _add_506_n401, _add_506_n400, _add_506_n399, _add_506_n398, _add_506_n397, _add_506_n396, _add_506_n395, _add_506_n394, _add_506_n393, _add_506_n392, _add_506_n391, _add_506_n390, _add_506_n389, _add_506_n388, 
  _add_506_n387, _add_506_n386, _add_506_n385, _add_506_n384, _add_506_n383, _add_506_n382, _add_506_n381, _add_506_n380, _add_506_n379, _add_506_n378, _add_506_n377, _add_506_n376, _add_506_n375, _add_506_n374, _add_506_n373, _add_506_n372, _add_506_n371, _add_506_n370, _add_506_n369, _add_506_n368, _add_506_n367, _add_506_n366, _add_506_n365, _add_506_n364, _add_506_n363, _add_506_n362, _add_506_n361, _add_506_n360, _add_506_n359, _add_506_n358, _add_506_n357, _add_506_n356, _add_506_n355, _add_506_n354, _add_506_n353, _add_506_n352, _add_506_n351, _add_506_n350, _add_506_n349, _add_506_n348, _add_506_n347, _add_506_n346, _add_506_n345, _add_506_n344, _add_506_n343, _add_506_n342, _add_506_n341, _add_506_n340, _add_506_n339, _add_506_n338, 
  _add_506_n337, _add_506_n336, _add_506_n335, _add_506_n334, _add_506_n333, _add_506_n332, _add_506_n331, _add_506_n330, _add_506_n329, _add_506_n328, _add_506_n327, _add_506_n326, _add_506_n325, _add_506_n324, _add_506_n323, _add_506_n322, _add_506_n321, _add_506_n320, _add_506_n319, _add_506_n318, _add_506_n317, _add_506_n316, _add_506_n315, _add_506_n314, _add_506_n313, _add_506_n312, _add_506_n311, _add_506_n310, _add_506_n309, _add_506_n308, _add_506_n307, _add_506_n306, _add_506_n305, _add_506_n304, _add_506_n303, _add_506_n302, _add_506_n301, _add_506_n300, _add_506_n299, _add_506_n298, _add_506_n297, _add_506_n296, _add_506_n295, _add_506_n294, _add_506_n293, _add_506_n292, _add_506_n291, _add_506_n290, _add_506_n289, _add_506_n288, 
  _add_506_n287, _add_506_n286, _add_506_n285, _add_506_n284, _add_506_n283, _add_506_n282, _add_506_n281, _add_506_n280, _add_506_n279, _add_506_n278, _add_506_n277, _add_506_n276, _add_506_n275, _add_506_n274, _add_506_n273, _add_506_n272, _add_506_n271, _add_506_n270, _add_506_n269, _add_506_n268, _add_506_n267, _add_506_n266, _add_506_n265, _add_506_n264, _add_506_n263, _add_506_n262, _add_506_n261, _add_506_n260, _add_506_n259, _add_506_n258, _add_506_n257, _add_506_n256, _add_506_n255, _add_506_n254, _add_506_n253, _add_506_n252, _add_506_n251, _add_506_n250, _add_506_n249, _add_506_n248, _add_506_n247, _add_506_n246, _add_506_n245, _add_506_n244, _add_506_n243, _add_506_n242, _add_506_n241, _add_506_n240, _add_506_n239, _add_506_n238, 
  _add_506_n237, _add_506_n236, _add_506_n235, _add_506_n234, _add_506_n233, _add_506_n232, _add_506_n231, _add_506_n230, _add_506_n229, _add_506_n228, _add_506_n227, _add_506_n226, _add_506_n225, _add_506_n224, _add_506_n223, _add_506_n222, _add_506_n221, _add_506_n220, _add_506_n219, _add_506_n218, _add_506_n217, _add_506_n216, _add_506_n215, _add_506_n214, _add_506_n213, _add_506_n212, _add_506_n211, _add_506_n210, _add_506_n209, _add_506_n208, _add_506_n207, _add_506_n206, _add_506_n205, _add_506_n204, _add_506_n203, _add_506_n202, _add_506_n201, _add_506_n200, _add_506_n199, _add_506_n198, _add_506_n197, _add_506_n196, _add_506_n195, _add_506_n194, _add_506_n193, _add_506_n192, _add_506_n191, _add_506_n190, _add_506_n189, _add_506_n188, 
  _add_506_n187, _add_506_n186, _add_506_n185, _add_506_n184, _add_506_n183, _add_506_n182, _add_506_n181, _add_506_n180, _add_506_n179, _add_506_n178, _add_506_n177, _add_506_n176, _add_506_n175, _add_506_n174, _add_506_n173, _add_506_n172, _add_506_n171, _add_506_n170, _add_506_n169, _add_506_n168, _add_506_n167, _add_506_n166, _add_506_n165, _add_506_n164, _add_506_n163, _add_506_n162, _add_506_n161, _add_506_n160, _add_506_n159, _add_506_n158, _add_506_n157, _add_506_n156, _add_506_n155, _add_506_n154, _add_506_n153, _add_506_n152, _add_506_n151, _add_506_n150, _add_506_n149, _add_506_n148, _add_506_n147, _add_506_n146, _add_506_n145, _add_506_n144, _add_506_n143, _add_506_n142, _add_506_n141, _add_506_n140, _add_506_n139, _add_506_n138, 
  _add_506_n137, _add_506_n136, _add_506_n135, _add_506_n134, _add_506_n133, _add_506_n132, _add_506_n131, _add_506_n130, _add_506_n129, _add_506_n128, _add_506_n127, _add_506_n126, _add_506_n125, _add_506_n124, _add_506_n123, _add_506_n122, _add_506_n121, _add_506_n120, _add_506_n119, _add_506_n118, _add_506_n117, _add_506_n116, _add_506_n115, _add_506_n114, _add_506_n113, _add_506_n112, _add_506_n111, _add_506_n110, _add_506_n109, _add_506_n108, _add_506_n107, _add_506_n106, _add_506_n105, _add_506_n104, _add_506_n103, _add_506_n102, _add_506_n101, _add_506_n100, _add_506_n99, _add_506_n98, _add_506_n97, _add_506_n96, _add_506_n95, _add_506_n94, _add_506_n93, _add_506_n92, _add_506_n91, _add_506_n90, _add_506_n89, _add_506_n88, 
  _add_506_n87, _add_506_n86, _add_506_n85, _add_506_n84, _add_506_n83, _add_506_n82, _add_506_n81, _add_506_n80, _add_506_n79, _add_506_n78, _add_506_n77, _add_506_n76, _add_506_n75, _add_506_n74, _add_506_n73, _add_506_n72, _add_506_n71, _add_506_n70, _add_506_n69, _add_506_n68, _add_506_n67, _add_506_n66, _add_506_n65, _add_506_n64, _add_506_n63, _add_506_n62, _add_506_n61, _add_506_n60, _add_506_n59, _add_506_n58, _add_506_n57, _add_506_n56, _add_506_n55, _add_506_n54, _add_506_n53, _add_506_n52, _add_506_n51, _add_506_n50, _add_506_n49, _add_506_n48, _add_506_n47, _add_506_n46, _add_506_n45, _add_506_n44, _add_506_n43, _add_506_n42, _add_506_n41, _add_506_n40, _add_506_n39, _add_506_n38, 
  _add_506_n37, _add_506_n36, _add_506_n35, _add_506_n34, _add_506_n33, _add_506_n32, _add_506_n31, _add_506_n30, _add_506_n29, _add_506_n28, _add_506_n27, _add_506_n26, _add_506_n25, _add_506_n24, _add_506_n23, _add_506_n22, _add_506_n21, _add_506_n20, _add_506_n19, _add_506_n18, _add_506_n17, _add_506_n16, _add_506_n15, _add_506_n14, _add_506_n13, _add_506_n12, _add_506_n11, _add_506_n10, _add_506_n9, _add_506_n8, _add_506_n7, _add_506_n6, _add_506_n4, _add_506_n3, _add_506_n2, _add_506_n1, _add_1_root_add_519_2_n224, _add_1_root_add_519_2_n223, _add_1_root_add_519_2_n222, _add_1_root_add_519_2_n221, _add_1_root_add_519_2_n220, _add_1_root_add_519_2_n219, _add_1_root_add_519_2_n218, _add_1_root_add_519_2_n217, _add_1_root_add_519_2_n216, _add_1_root_add_519_2_n215, _add_1_root_add_519_2_n214, _add_1_root_add_519_2_n213, _add_1_root_add_519_2_n212, _add_1_root_add_519_2_n211, 
  _add_1_root_add_519_2_n210, _add_1_root_add_519_2_n209, _add_1_root_add_519_2_n208, _add_1_root_add_519_2_n207, _add_1_root_add_519_2_n206, _add_1_root_add_519_2_n205, _add_1_root_add_519_2_n204, _add_1_root_add_519_2_n203, _add_1_root_add_519_2_n202, _add_1_root_add_519_2_n201, _add_1_root_add_519_2_n200, _add_1_root_add_519_2_n199, _add_1_root_add_519_2_n198, _add_1_root_add_519_2_n197, _add_1_root_add_519_2_n196, _add_1_root_add_519_2_n195, _add_1_root_add_519_2_n194, _add_1_root_add_519_2_n193, _add_1_root_add_519_2_n192, _add_1_root_add_519_2_n191, _add_1_root_add_519_2_n190, _add_1_root_add_519_2_n189, _add_1_root_add_519_2_n188, _add_1_root_add_519_2_n187, _add_1_root_add_519_2_n186, _add_1_root_add_519_2_n185, _add_1_root_add_519_2_n184, _add_1_root_add_519_2_n183, _add_1_root_add_519_2_n182, _add_1_root_add_519_2_n181, _add_1_root_add_519_2_n180, _add_1_root_add_519_2_n179, _add_1_root_add_519_2_n178, _add_1_root_add_519_2_n177, _add_1_root_add_519_2_n176, _add_1_root_add_519_2_n175, _add_1_root_add_519_2_n174, _add_1_root_add_519_2_n173, _add_1_root_add_519_2_n172, _add_1_root_add_519_2_n171, _add_1_root_add_519_2_n170, _add_1_root_add_519_2_n169, _add_1_root_add_519_2_n168, _add_1_root_add_519_2_n167, _add_1_root_add_519_2_n166, _add_1_root_add_519_2_n165, _add_1_root_add_519_2_n164, _add_1_root_add_519_2_n163, _add_1_root_add_519_2_n162, _add_1_root_add_519_2_n161, 
  _add_1_root_add_519_2_n160, _add_1_root_add_519_2_n159, _add_1_root_add_519_2_n158, _add_1_root_add_519_2_n157, _add_1_root_add_519_2_n156, _add_1_root_add_519_2_n155, _add_1_root_add_519_2_n154, _add_1_root_add_519_2_n153, _add_1_root_add_519_2_n152, _add_1_root_add_519_2_n151, _add_1_root_add_519_2_n150, _add_1_root_add_519_2_n149, _add_1_root_add_519_2_n148, _add_1_root_add_519_2_n147, _add_1_root_add_519_2_n146, _add_1_root_add_519_2_n145, _add_1_root_add_519_2_n144, _add_1_root_add_519_2_n143, _add_1_root_add_519_2_n142, _add_1_root_add_519_2_n141, _add_1_root_add_519_2_n140, _add_1_root_add_519_2_n139, _add_1_root_add_519_2_n138, _add_1_root_add_519_2_n137, _add_1_root_add_519_2_n136, _add_1_root_add_519_2_n135, _add_1_root_add_519_2_n134, _add_1_root_add_519_2_n133, _add_1_root_add_519_2_n132, _add_1_root_add_519_2_n131, _add_1_root_add_519_2_n130, _add_1_root_add_519_2_n129, _add_1_root_add_519_2_n128, _add_1_root_add_519_2_n127, _add_1_root_add_519_2_n126, _add_1_root_add_519_2_n125, _add_1_root_add_519_2_n124, _add_1_root_add_519_2_n123, _add_1_root_add_519_2_n122, _add_1_root_add_519_2_n121, _add_1_root_add_519_2_n120, _add_1_root_add_519_2_n119, _add_1_root_add_519_2_n118, _add_1_root_add_519_2_n117, _add_1_root_add_519_2_n116, _add_1_root_add_519_2_n115, _add_1_root_add_519_2_n114, _add_1_root_add_519_2_n113, _add_1_root_add_519_2_n112, _add_1_root_add_519_2_n111, 
  _add_1_root_add_519_2_n110, _add_1_root_add_519_2_n109, _add_1_root_add_519_2_n108, _add_1_root_add_519_2_n107, _add_1_root_add_519_2_n106, _add_1_root_add_519_2_n105, _add_1_root_add_519_2_n104, _add_1_root_add_519_2_n103, _add_1_root_add_519_2_n102, _add_1_root_add_519_2_n101, _add_1_root_add_519_2_n100, _add_1_root_add_519_2_n99, _add_1_root_add_519_2_n98, _add_1_root_add_519_2_n97, _add_1_root_add_519_2_n96, _add_1_root_add_519_2_n95, _add_1_root_add_519_2_n94, _add_1_root_add_519_2_n93, _add_1_root_add_519_2_n92, _add_1_root_add_519_2_n91, _add_1_root_add_519_2_n90, _add_1_root_add_519_2_n89, _add_1_root_add_519_2_n88, _add_1_root_add_519_2_n87, _add_1_root_add_519_2_n86, _add_1_root_add_519_2_n85, _add_1_root_add_519_2_n84, _add_1_root_add_519_2_n83, _add_1_root_add_519_2_n82, _add_1_root_add_519_2_n81, _add_1_root_add_519_2_n80, _add_1_root_add_519_2_n79, _add_1_root_add_519_2_n78, _add_1_root_add_519_2_n77, _add_1_root_add_519_2_n76, _add_1_root_add_519_2_n75, _add_1_root_add_519_2_n74, _add_1_root_add_519_2_n73, _add_1_root_add_519_2_n72, _add_1_root_add_519_2_n71, _add_1_root_add_519_2_n70, _add_1_root_add_519_2_n69, _add_1_root_add_519_2_n68, _add_1_root_add_519_2_n67, _add_1_root_add_519_2_n66, _add_1_root_add_519_2_n65, _add_1_root_add_519_2_n64, _add_1_root_add_519_2_n63, _add_1_root_add_519_2_n62, _add_1_root_add_519_2_n61, 
  _add_1_root_add_519_2_n60, _add_1_root_add_519_2_n59, _add_1_root_add_519_2_n58, _add_1_root_add_519_2_n57, _add_1_root_add_519_2_n56, _add_1_root_add_519_2_n55, _add_1_root_add_519_2_n54, _add_1_root_add_519_2_n53, _add_1_root_add_519_2_n52, _add_1_root_add_519_2_n51, _add_1_root_add_519_2_n50, _add_1_root_add_519_2_n49, _add_1_root_add_519_2_n48, _add_1_root_add_519_2_n47, _add_1_root_add_519_2_n46, _add_1_root_add_519_2_n45, _add_1_root_add_519_2_n44, _add_1_root_add_519_2_n43, _add_1_root_add_519_2_n42, _add_1_root_add_519_2_n41, _add_1_root_add_519_2_n40, _add_1_root_add_519_2_n39, _add_1_root_add_519_2_n38, _add_1_root_add_519_2_n37, _add_1_root_add_519_2_n36, _add_1_root_add_519_2_n35, _add_1_root_add_519_2_n34, _add_1_root_add_519_2_n33, _add_1_root_add_519_2_n32, _add_1_root_add_519_2_n31, _add_1_root_add_519_2_n30, _add_1_root_add_519_2_n29, _add_1_root_add_519_2_n28, _add_1_root_add_519_2_n27, _add_1_root_add_519_2_n26, _add_1_root_add_519_2_n25, _add_1_root_add_519_2_n24, _add_1_root_add_519_2_n23, _add_1_root_add_519_2_n22, _add_1_root_add_519_2_n21, _add_1_root_add_519_2_n20, _add_1_root_add_519_2_n19, _add_1_root_add_519_2_n18, _add_1_root_add_519_2_n17, _add_1_root_add_519_2_n16, _add_1_root_add_519_2_n15, _add_1_root_add_519_2_n14, _add_1_root_add_519_2_n13, _add_1_root_add_519_2_n12, _add_1_root_add_519_2_n11, 
  _add_1_root_add_519_2_n10, _add_1_root_add_519_2_n9, _add_1_root_add_519_2_n8, _add_1_root_add_519_2_n7, _add_1_root_add_519_2_n6, _add_1_root_add_519_2_n5, _add_1_root_add_519_2_n4, _add_1_root_add_519_2_n3, _add_1_root_add_519_2_n2, _add_1_root_add_519_2_n1, _add_1_root_add_513_2_n224, _add_1_root_add_513_2_n223, _add_1_root_add_513_2_n222, _add_1_root_add_513_2_n221, _add_1_root_add_513_2_n220, _add_1_root_add_513_2_n219, _add_1_root_add_513_2_n218, _add_1_root_add_513_2_n217, _add_1_root_add_513_2_n216, _add_1_root_add_513_2_n215, _add_1_root_add_513_2_n214, _add_1_root_add_513_2_n213, _add_1_root_add_513_2_n212, _add_1_root_add_513_2_n211, _add_1_root_add_513_2_n210, _add_1_root_add_513_2_n209, _add_1_root_add_513_2_n208, _add_1_root_add_513_2_n207, _add_1_root_add_513_2_n206, _add_1_root_add_513_2_n205, _add_1_root_add_513_2_n204, _add_1_root_add_513_2_n203, _add_1_root_add_513_2_n202, _add_1_root_add_513_2_n201, _add_1_root_add_513_2_n200, _add_1_root_add_513_2_n199, _add_1_root_add_513_2_n198, _add_1_root_add_513_2_n197, _add_1_root_add_513_2_n196, _add_1_root_add_513_2_n195, _add_1_root_add_513_2_n194, _add_1_root_add_513_2_n193, _add_1_root_add_513_2_n192, _add_1_root_add_513_2_n191, _add_1_root_add_513_2_n190, _add_1_root_add_513_2_n189, _add_1_root_add_513_2_n188, _add_1_root_add_513_2_n187, _add_1_root_add_513_2_n186, _add_1_root_add_513_2_n185, 
  _add_1_root_add_513_2_n184, _add_1_root_add_513_2_n183, _add_1_root_add_513_2_n182, _add_1_root_add_513_2_n181, _add_1_root_add_513_2_n180, _add_1_root_add_513_2_n179, _add_1_root_add_513_2_n178, _add_1_root_add_513_2_n177, _add_1_root_add_513_2_n176, _add_1_root_add_513_2_n175, _add_1_root_add_513_2_n174, _add_1_root_add_513_2_n173, _add_1_root_add_513_2_n172, _add_1_root_add_513_2_n171, _add_1_root_add_513_2_n170, _add_1_root_add_513_2_n169, _add_1_root_add_513_2_n168, _add_1_root_add_513_2_n167, _add_1_root_add_513_2_n166, _add_1_root_add_513_2_n165, _add_1_root_add_513_2_n164, _add_1_root_add_513_2_n163, _add_1_root_add_513_2_n162, _add_1_root_add_513_2_n161, _add_1_root_add_513_2_n160, _add_1_root_add_513_2_n159, _add_1_root_add_513_2_n158, _add_1_root_add_513_2_n157, _add_1_root_add_513_2_n156, _add_1_root_add_513_2_n155, _add_1_root_add_513_2_n154, _add_1_root_add_513_2_n153, _add_1_root_add_513_2_n152, _add_1_root_add_513_2_n151, _add_1_root_add_513_2_n150, _add_1_root_add_513_2_n149, _add_1_root_add_513_2_n148, _add_1_root_add_513_2_n147, _add_1_root_add_513_2_n146, _add_1_root_add_513_2_n145, _add_1_root_add_513_2_n144, _add_1_root_add_513_2_n143, _add_1_root_add_513_2_n142, _add_1_root_add_513_2_n141, _add_1_root_add_513_2_n140, _add_1_root_add_513_2_n139, _add_1_root_add_513_2_n138, _add_1_root_add_513_2_n137, _add_1_root_add_513_2_n136, _add_1_root_add_513_2_n135, 
  _add_1_root_add_513_2_n134, _add_1_root_add_513_2_n133, _add_1_root_add_513_2_n132, _add_1_root_add_513_2_n131, _add_1_root_add_513_2_n130, _add_1_root_add_513_2_n129, _add_1_root_add_513_2_n128, _add_1_root_add_513_2_n127, _add_1_root_add_513_2_n126, _add_1_root_add_513_2_n125, _add_1_root_add_513_2_n124, _add_1_root_add_513_2_n123, _add_1_root_add_513_2_n122, _add_1_root_add_513_2_n121, _add_1_root_add_513_2_n120, _add_1_root_add_513_2_n119, _add_1_root_add_513_2_n118, _add_1_root_add_513_2_n117, _add_1_root_add_513_2_n116, _add_1_root_add_513_2_n115, _add_1_root_add_513_2_n114, _add_1_root_add_513_2_n113, _add_1_root_add_513_2_n112, _add_1_root_add_513_2_n111, _add_1_root_add_513_2_n110, _add_1_root_add_513_2_n109, _add_1_root_add_513_2_n108, _add_1_root_add_513_2_n107, _add_1_root_add_513_2_n106, _add_1_root_add_513_2_n105, _add_1_root_add_513_2_n104, _add_1_root_add_513_2_n103, _add_1_root_add_513_2_n102, _add_1_root_add_513_2_n101, _add_1_root_add_513_2_n100, _add_1_root_add_513_2_n99, _add_1_root_add_513_2_n98, _add_1_root_add_513_2_n97, _add_1_root_add_513_2_n96, _add_1_root_add_513_2_n95, _add_1_root_add_513_2_n94, _add_1_root_add_513_2_n93, _add_1_root_add_513_2_n92, _add_1_root_add_513_2_n91, _add_1_root_add_513_2_n90, _add_1_root_add_513_2_n89, _add_1_root_add_513_2_n88, _add_1_root_add_513_2_n87, _add_1_root_add_513_2_n86, _add_1_root_add_513_2_n85, 
  _add_1_root_add_513_2_n84, _add_1_root_add_513_2_n83, _add_1_root_add_513_2_n82, _add_1_root_add_513_2_n81, _add_1_root_add_513_2_n80, _add_1_root_add_513_2_n79, _add_1_root_add_513_2_n78, _add_1_root_add_513_2_n77, _add_1_root_add_513_2_n76, _add_1_root_add_513_2_n75, _add_1_root_add_513_2_n74, _add_1_root_add_513_2_n73, _add_1_root_add_513_2_n72, _add_1_root_add_513_2_n71, _add_1_root_add_513_2_n70, _add_1_root_add_513_2_n69, _add_1_root_add_513_2_n68, _add_1_root_add_513_2_n67, _add_1_root_add_513_2_n66, _add_1_root_add_513_2_n65, _add_1_root_add_513_2_n64, _add_1_root_add_513_2_n63, _add_1_root_add_513_2_n62, _add_1_root_add_513_2_n61, _add_1_root_add_513_2_n60, _add_1_root_add_513_2_n59, _add_1_root_add_513_2_n58, _add_1_root_add_513_2_n57, _add_1_root_add_513_2_n56, _add_1_root_add_513_2_n55, _add_1_root_add_513_2_n54, _add_1_root_add_513_2_n53, _add_1_root_add_513_2_n52, _add_1_root_add_513_2_n51, _add_1_root_add_513_2_n50, _add_1_root_add_513_2_n49, _add_1_root_add_513_2_n48, _add_1_root_add_513_2_n47, _add_1_root_add_513_2_n46, _add_1_root_add_513_2_n45, _add_1_root_add_513_2_n44, _add_1_root_add_513_2_n43, _add_1_root_add_513_2_n42, _add_1_root_add_513_2_n41, _add_1_root_add_513_2_n40, _add_1_root_add_513_2_n39, _add_1_root_add_513_2_n38, _add_1_root_add_513_2_n37, _add_1_root_add_513_2_n36, _add_1_root_add_513_2_n35, 
  _add_1_root_add_513_2_n34, _add_1_root_add_513_2_n33, _add_1_root_add_513_2_n32, _add_1_root_add_513_2_n31, _add_1_root_add_513_2_n30, _add_1_root_add_513_2_n29, _add_1_root_add_513_2_n28, _add_1_root_add_513_2_n27, _add_1_root_add_513_2_n26, _add_1_root_add_513_2_n25, _add_1_root_add_513_2_n24, _add_1_root_add_513_2_n23, _add_1_root_add_513_2_n22, _add_1_root_add_513_2_n21, _add_1_root_add_513_2_n20, _add_1_root_add_513_2_n19, _add_1_root_add_513_2_n18, _add_1_root_add_513_2_n17, _add_1_root_add_513_2_n16, _add_1_root_add_513_2_n15, _add_1_root_add_513_2_n14, _add_1_root_add_513_2_n13, _add_1_root_add_513_2_n12, _add_1_root_add_513_2_n11, _add_1_root_add_513_2_n10, _add_1_root_add_513_2_n9, _add_1_root_add_513_2_n8, _add_1_root_add_513_2_n7, _add_1_root_add_513_2_n6, _add_1_root_add_513_2_n5, _add_1_root_add_513_2_n4, _add_1_root_add_513_2_n3, _add_1_root_add_513_2_n2, _add_1_root_add_513_2_n1 ;
wire [9:0] state;
wire [127:0] aes_text_in;
wire [127:0] aes_text_out;
wire [63:0] aad_byte_cnt;
wire [63:0] enc_byte_cnt;
wire [127:0] z_out;
wire [127:0] v_in;
wire [127:0] z_in;
wire [127:0] b_in;
wire [127:0] v_out;
wire [7:0] _AES_ENC_sa00_next;
wire [7:0] _AES_ENC_sa00;
wire [7:0] _AES_ENC_sa10_next;
wire [7:0] _AES_ENC_sa10;
wire [7:0] _AES_ENC_sa20_next;
wire [7:0] _AES_ENC_sa20;
wire [7:0] _AES_ENC_sa30_next;
wire [7:0] _AES_ENC_sa30;
wire [7:0] _AES_ENC_sa01_next;
wire [7:0] _AES_ENC_sa01;
wire [7:0] _AES_ENC_sa11_next;
wire [7:0] _AES_ENC_sa11;
wire [7:0] _AES_ENC_sa21_next;
wire [7:0] _AES_ENC_sa21;
wire [7:0] _AES_ENC_sa31_next;
wire [7:0] _AES_ENC_sa31;
wire [7:0] _AES_ENC_sa02_next;
wire [7:0] _AES_ENC_sa02;
wire [7:0] _AES_ENC_sa12_next;
wire [7:0] _AES_ENC_sa12;
wire [7:0] _AES_ENC_sa22_next;
wire [7:0] _AES_ENC_sa22;
wire [7:0] _AES_ENC_sa32_next;
wire [7:0] _AES_ENC_sa32;
wire [7:0] _AES_ENC_sa03_next;
wire [7:0] _AES_ENC_sa03;
wire [7:0] _AES_ENC_sa13_next;
wire [7:0] _AES_ENC_sa13;
wire [7:0] _AES_ENC_sa23_next;
wire [7:0] _AES_ENC_sa23;
wire [7:0] __AES_ENC_sa33_next;
wire [7:0] _AES_ENC_sa33;
wire [31:24] _AES_ENC_u0_rcon;
CLKBUFX1 gbuf_d_1(.A(n6027), .Y(d_out_1));
CLKBUFX1 gbuf_q_1(.A(q_in_1), .Y(n17292));
CLKBUFX1 gbuf_d_2(.A(n6028), .Y(d_out_2));
CLKBUFX1 gbuf_q_2(.A(q_in_2), .Y(n17293));
CLKBUFX1 gbuf_d_3(.A(n6029), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(n17294));
CLKBUFX1 gbuf_d_4(.A(n6030), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(n17295));
CLKBUFX1 gbuf_d_5(.A(n6031), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(n17296));
CLKBUFX1 gbuf_d_6(.A(n6032), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(n17297));
CLKBUFX1 gbuf_d_7(.A(n6033), .Y(d_out_7));
CLKBUFX1 gbuf_q_7(.A(q_in_7), .Y(n17298));
CLKBUFX1 gbuf_d_8(.A(n6034), .Y(d_out_8));
CLKBUFX1 gbuf_q_8(.A(q_in_8), .Y(n17299));
CLKBUFX1 gbuf_d_9(.A(n6035), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(n17300));
CLKBUFX1 gbuf_d_10(.A(n6036), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(n17301));
CLKBUFX1 gbuf_d_11(.A(n6037), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(n17302));
CLKBUFX1 gbuf_d_12(.A(n6038), .Y(d_out_12));
CLKBUFX1 gbuf_q_12(.A(q_in_12), .Y(n17303));
CLKBUFX1 gbuf_d_13(.A(n6039), .Y(d_out_13));
CLKBUFX1 gbuf_q_13(.A(q_in_13), .Y(n17304));
CLKBUFX1 gbuf_d_14(.A(n6040), .Y(d_out_14));
CLKBUFX1 gbuf_q_14(.A(q_in_14), .Y(n17305));
CLKBUFX1 gbuf_d_15(.A(n6041), .Y(d_out_15));
CLKBUFX1 gbuf_q_15(.A(q_in_15), .Y(n17306));
CLKBUFX1 gbuf_d_16(.A(n6042), .Y(d_out_16));
CLKBUFX1 gbuf_q_16(.A(q_in_16), .Y(n17307));
CLKBUFX1 gbuf_d_17(.A(n6043), .Y(d_out_17));
CLKBUFX1 gbuf_q_17(.A(q_in_17), .Y(n17308));
CLKBUFX1 gbuf_d_18(.A(n6044), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(n17309));
CLKBUFX1 gbuf_d_19(.A(n6045), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(n17310));
CLKBUFX1 gbuf_d_20(.A(n6046), .Y(d_out_20));
CLKBUFX1 gbuf_q_20(.A(q_in_20), .Y(n17311));
CLKBUFX1 gbuf_d_21(.A(n6047), .Y(d_out_21));
CLKBUFX1 gbuf_q_21(.A(q_in_21), .Y(n17312));
CLKBUFX1 gbuf_d_22(.A(n6048), .Y(d_out_22));
CLKBUFX1 gbuf_q_22(.A(q_in_22), .Y(n17313));
CLKBUFX1 gbuf_d_23(.A(n6049), .Y(d_out_23));
CLKBUFX1 gbuf_q_23(.A(q_in_23), .Y(n17314));
CLKBUFX1 gbuf_d_24(.A(n6050), .Y(d_out_24));
CLKBUFX1 gbuf_q_24(.A(q_in_24), .Y(n17315));
CLKBUFX1 gbuf_d_25(.A(n6051), .Y(d_out_25));
CLKBUFX1 gbuf_q_25(.A(q_in_25), .Y(n17316));
CLKBUFX1 gbuf_d_26(.A(n6052), .Y(d_out_26));
CLKBUFX1 gbuf_q_26(.A(q_in_26), .Y(n17317));
CLKBUFX1 gbuf_d_27(.A(n6053), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(n17318));
CLKBUFX1 gbuf_d_28(.A(n6054), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(n17319));
CLKBUFX1 gbuf_d_29(.A(n6055), .Y(d_out_29));
CLKBUFX1 gbuf_q_29(.A(q_in_29), .Y(n17320));
CLKBUFX1 gbuf_d_30(.A(n6056), .Y(d_out_30));
CLKBUFX1 gbuf_q_30(.A(q_in_30), .Y(n17321));
CLKBUFX1 gbuf_d_31(.A(n6057), .Y(d_out_31));
CLKBUFX1 gbuf_q_31(.A(q_in_31), .Y(n17322));
CLKBUFX1 gbuf_d_32(.A(n6058), .Y(d_out_32));
CLKBUFX1 gbuf_q_32(.A(q_in_32), .Y(n17323));
CLKBUFX1 gbuf_d_33(.A(n6059), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(n17324));
CLKBUFX1 gbuf_d_34(.A(n6060), .Y(d_out_34));
CLKBUFX1 gbuf_q_34(.A(q_in_34), .Y(n17325));
CLKBUFX1 gbuf_d_35(.A(n6061), .Y(d_out_35));
CLKBUFX1 gbuf_q_35(.A(q_in_35), .Y(n17326));
CLKBUFX1 gbuf_d_36(.A(n6062), .Y(d_out_36));
CLKBUFX1 gbuf_q_36(.A(q_in_36), .Y(n17327));
CLKBUFX1 gbuf_d_37(.A(n6063), .Y(d_out_37));
CLKBUFX1 gbuf_q_37(.A(q_in_37), .Y(n17328));
CLKBUFX1 gbuf_d_38(.A(n6064), .Y(d_out_38));
CLKBUFX1 gbuf_q_38(.A(q_in_38), .Y(n17329));
CLKBUFX1 gbuf_d_39(.A(n6065), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(n17330));
CLKBUFX1 gbuf_d_40(.A(n6066), .Y(d_out_40));
CLKBUFX1 gbuf_q_40(.A(q_in_40), .Y(n17331));
CLKBUFX1 gbuf_d_41(.A(n6067), .Y(d_out_41));
CLKBUFX1 gbuf_q_41(.A(q_in_41), .Y(n17332));
CLKBUFX1 gbuf_d_42(.A(n6068), .Y(d_out_42));
CLKBUFX1 gbuf_q_42(.A(q_in_42), .Y(n17333));
CLKBUFX1 gbuf_d_43(.A(n6069), .Y(d_out_43));
CLKBUFX1 gbuf_q_43(.A(q_in_43), .Y(n17334));
CLKBUFX1 gbuf_d_44(.A(n6070), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(n17335));
CLKBUFX1 gbuf_d_45(.A(n6071), .Y(d_out_45));
CLKBUFX1 gbuf_q_45(.A(q_in_45), .Y(n17336));
CLKBUFX1 gbuf_d_46(.A(n6072), .Y(d_out_46));
CLKBUFX1 gbuf_q_46(.A(q_in_46), .Y(n17337));
CLKBUFX1 gbuf_d_47(.A(n6073), .Y(d_out_47));
CLKBUFX1 gbuf_q_47(.A(q_in_47), .Y(n17338));
CLKBUFX1 gbuf_d_48(.A(n6074), .Y(d_out_48));
CLKBUFX1 gbuf_q_48(.A(q_in_48), .Y(n17339));
CLKBUFX1 gbuf_d_49(.A(n6075), .Y(d_out_49));
CLKBUFX1 gbuf_q_49(.A(q_in_49), .Y(n17340));
CLKBUFX1 gbuf_d_50(.A(n6076), .Y(d_out_50));
CLKBUFX1 gbuf_q_50(.A(q_in_50), .Y(n17341));
CLKBUFX1 gbuf_d_51(.A(n6077), .Y(d_out_51));
CLKBUFX1 gbuf_q_51(.A(q_in_51), .Y(n17342));
CLKBUFX1 gbuf_d_52(.A(n6078), .Y(d_out_52));
CLKBUFX1 gbuf_q_52(.A(q_in_52), .Y(n17343));
CLKBUFX1 gbuf_d_53(.A(n6079), .Y(d_out_53));
CLKBUFX1 gbuf_q_53(.A(q_in_53), .Y(n17344));
CLKBUFX1 gbuf_d_54(.A(n6080), .Y(d_out_54));
CLKBUFX1 gbuf_q_54(.A(q_in_54), .Y(n17345));
CLKBUFX1 gbuf_d_55(.A(n6081), .Y(d_out_55));
CLKBUFX1 gbuf_q_55(.A(q_in_55), .Y(n17346));
CLKBUFX1 gbuf_d_56(.A(n6082), .Y(d_out_56));
CLKBUFX1 gbuf_q_56(.A(q_in_56), .Y(n17347));
CLKBUFX1 gbuf_d_57(.A(n6083), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(n17348));
CLKBUFX1 gbuf_d_58(.A(n6084), .Y(d_out_58));
CLKBUFX1 gbuf_q_58(.A(q_in_58), .Y(n17349));
CLKBUFX1 gbuf_d_59(.A(n6085), .Y(d_out_59));
CLKBUFX1 gbuf_q_59(.A(q_in_59), .Y(n17350));
CLKBUFX1 gbuf_d_60(.A(n6086), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(n17351));
CLKBUFX1 gbuf_d_61(.A(n6087), .Y(d_out_61));
CLKBUFX1 gbuf_q_61(.A(q_in_61), .Y(n17352));
CLKBUFX1 gbuf_d_62(.A(n6088), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(n17353));
CLKBUFX1 gbuf_d_63(.A(n6089), .Y(d_out_63));
CLKBUFX1 gbuf_q_63(.A(q_in_63), .Y(n17354));
CLKBUFX1 gbuf_d_64(.A(n6090), .Y(d_out_64));
CLKBUFX1 gbuf_q_64(.A(q_in_64), .Y(n17355));
CLKBUFX1 gbuf_d_65(.A(n6091), .Y(d_out_65));
CLKBUFX1 gbuf_q_65(.A(q_in_65), .Y(n17356));
CLKBUFX1 gbuf_d_66(.A(n6092), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(n17357));
CLKBUFX1 gbuf_d_67(.A(n6093), .Y(d_out_67));
CLKBUFX1 gbuf_q_67(.A(q_in_67), .Y(n17358));
CLKBUFX1 gbuf_d_68(.A(n6094), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(n17359));
CLKBUFX1 gbuf_d_69(.A(n6095), .Y(d_out_69));
CLKBUFX1 gbuf_q_69(.A(q_in_69), .Y(n17360));
CLKBUFX1 gbuf_d_70(.A(n6096), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(n17361));
CLKBUFX1 gbuf_d_71(.A(n6097), .Y(d_out_71));
CLKBUFX1 gbuf_q_71(.A(q_in_71), .Y(n17362));
CLKBUFX1 gbuf_d_72(.A(n6098), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(n17363));
CLKBUFX1 gbuf_d_73(.A(n6099), .Y(d_out_73));
CLKBUFX1 gbuf_q_73(.A(q_in_73), .Y(n17364));
CLKBUFX1 gbuf_d_74(.A(n6100), .Y(d_out_74));
CLKBUFX1 gbuf_q_74(.A(q_in_74), .Y(n17365));
CLKBUFX1 gbuf_d_75(.A(n6101), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(n17366));
CLKBUFX1 gbuf_d_76(.A(n6102), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(n17367));
CLKBUFX1 gbuf_d_77(.A(n6103), .Y(d_out_77));
CLKBUFX1 gbuf_q_77(.A(q_in_77), .Y(n17368));
CLKBUFX1 gbuf_d_78(.A(n6104), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(n17369));
CLKBUFX1 gbuf_d_79(.A(n6105), .Y(d_out_79));
CLKBUFX1 gbuf_q_79(.A(q_in_79), .Y(n17370));
CLKBUFX1 gbuf_d_80(.A(n6106), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(n17371));
CLKBUFX1 gbuf_d_81(.A(n6107), .Y(d_out_81));
CLKBUFX1 gbuf_q_81(.A(q_in_81), .Y(n17372));
CLKBUFX1 gbuf_d_82(.A(n6108), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(n17373));
CLKBUFX1 gbuf_d_83(.A(n6109), .Y(d_out_83));
CLKBUFX1 gbuf_q_83(.A(q_in_83), .Y(n17374));
CLKBUFX1 gbuf_d_84(.A(n6156), .Y(d_out_84));
CLKBUFX1 gbuf_qn_84(.A(qn_in_84), .Y(n17027));
CLKBUFX1 gbuf_d_85(.A(n6157), .Y(d_out_85));
CLKBUFX1 gbuf_qn_85(.A(qn_in_85), .Y(n17029));
CLKBUFX1 gbuf_d_86(.A(n6159), .Y(d_out_86));
CLKBUFX1 gbuf_qn_86(.A(qn_in_86), .Y(n17033));
CLKBUFX1 gbuf_d_87(.A(n6161), .Y(d_out_87));
CLKBUFX1 gbuf_qn_87(.A(qn_in_87), .Y(n17037));
CLKBUFX1 gbuf_d_88(.A(n6162), .Y(d_out_88));
CLKBUFX1 gbuf_qn_88(.A(qn_in_88), .Y(n17039));
CLKBUFX1 gbuf_d_89(.A(n6163), .Y(d_out_89));
CLKBUFX1 gbuf_qn_89(.A(qn_in_89), .Y(n17041));
CLKBUFX1 gbuf_d_90(.A(n6164), .Y(d_out_90));
CLKBUFX1 gbuf_qn_90(.A(qn_in_90), .Y(n17043));
CLKBUFX1 gbuf_d_91(.A(n6165), .Y(d_out_91));
CLKBUFX1 gbuf_qn_91(.A(qn_in_91), .Y(n17045));
CLKBUFX1 gbuf_d_92(.A(n6166), .Y(d_out_92));
CLKBUFX1 gbuf_qn_92(.A(qn_in_92), .Y(n17047));
CLKBUFX1 gbuf_d_93(.A(n6167), .Y(d_out_93));
CLKBUFX1 gbuf_qn_93(.A(qn_in_93), .Y(n17049));
CLKBUFX1 gbuf_d_94(.A(n6168), .Y(d_out_94));
CLKBUFX1 gbuf_qn_94(.A(qn_in_94), .Y(n17051));
CLKBUFX1 gbuf_d_95(.A(n6169), .Y(d_out_95));
CLKBUFX1 gbuf_qn_95(.A(qn_in_95), .Y(n17053));
CLKBUFX1 gbuf_d_96(.A(n6170), .Y(d_out_96));
CLKBUFX1 gbuf_qn_96(.A(qn_in_96), .Y(n17055));
CLKBUFX1 gbuf_d_97(.A(n6171), .Y(d_out_97));
CLKBUFX1 gbuf_qn_97(.A(qn_in_97), .Y(n17057));
CLKBUFX1 gbuf_d_98(.A(n6172), .Y(d_out_98));
CLKBUFX1 gbuf_qn_98(.A(qn_in_98), .Y(n17059));
CLKBUFX1 gbuf_d_99(.A(n6173), .Y(d_out_99));
CLKBUFX1 gbuf_qn_99(.A(qn_in_99), .Y(n17061));
CLKBUFX1 gbuf_d_100(.A(n6174), .Y(d_out_100));
CLKBUFX1 gbuf_qn_100(.A(qn_in_100), .Y(n17063));
CLKBUFX1 gbuf_d_101(.A(n6175), .Y(d_out_101));
CLKBUFX1 gbuf_qn_101(.A(qn_in_101), .Y(n17065));
CLKBUFX1 gbuf_d_102(.A(n6176), .Y(d_out_102));
CLKBUFX1 gbuf_qn_102(.A(qn_in_102), .Y(n17067));
CLKBUFX1 gbuf_d_103(.A(n6177), .Y(d_out_103));
CLKBUFX1 gbuf_qn_103(.A(qn_in_103), .Y(n17069));
CLKBUFX1 gbuf_d_104(.A(n6178), .Y(d_out_104));
CLKBUFX1 gbuf_qn_104(.A(qn_in_104), .Y(n17071));
CLKBUFX1 gbuf_d_105(.A(n6179), .Y(d_out_105));
CLKBUFX1 gbuf_qn_105(.A(qn_in_105), .Y(n17073));
CLKBUFX1 gbuf_d_106(.A(n6180), .Y(d_out_106));
CLKBUFX1 gbuf_qn_106(.A(qn_in_106), .Y(n17075));
CLKBUFX1 gbuf_d_107(.A(n6181), .Y(d_out_107));
CLKBUFX1 gbuf_qn_107(.A(qn_in_107), .Y(n17077));
CLKBUFX1 gbuf_d_108(.A(n6182), .Y(d_out_108));
CLKBUFX1 gbuf_qn_108(.A(qn_in_108), .Y(n17079));
CLKBUFX1 gbuf_d_109(.A(n6183), .Y(d_out_109));
CLKBUFX1 gbuf_qn_109(.A(qn_in_109), .Y(n17081));
CLKBUFX1 gbuf_d_110(.A(n6184), .Y(d_out_110));
CLKBUFX1 gbuf_qn_110(.A(qn_in_110), .Y(n17083));
CLKBUFX1 gbuf_d_111(.A(n6185), .Y(d_out_111));
CLKBUFX1 gbuf_qn_111(.A(qn_in_111), .Y(n17085));
CLKBUFX1 gbuf_d_112(.A(n6186), .Y(d_out_112));
CLKBUFX1 gbuf_qn_112(.A(qn_in_112), .Y(n17087));
CLKBUFX1 gbuf_d_113(.A(n6187), .Y(d_out_113));
CLKBUFX1 gbuf_qn_113(.A(qn_in_113), .Y(n17089));
CLKBUFX1 gbuf_d_114(.A(n6188), .Y(d_out_114));
CLKBUFX1 gbuf_qn_114(.A(qn_in_114), .Y(n17091));
CLKBUFX1 gbuf_d_115(.A(n6189), .Y(d_out_115));
CLKBUFX1 gbuf_qn_115(.A(qn_in_115), .Y(n17093));
CLKBUFX1 gbuf_d_116(.A(n6190), .Y(d_out_116));
CLKBUFX1 gbuf_qn_116(.A(qn_in_116), .Y(n17095));
CLKBUFX1 gbuf_d_117(.A(n6191), .Y(d_out_117));
CLKBUFX1 gbuf_qn_117(.A(qn_in_117), .Y(n17097));
CLKBUFX1 gbuf_d_118(.A(n6192), .Y(d_out_118));
CLKBUFX1 gbuf_qn_118(.A(qn_in_118), .Y(n17099));
CLKBUFX1 gbuf_d_119(.A(n6193), .Y(d_out_119));
CLKBUFX1 gbuf_qn_119(.A(qn_in_119), .Y(n17101));
CLKBUFX1 gbuf_d_120(.A(n6194), .Y(d_out_120));
CLKBUFX1 gbuf_qn_120(.A(qn_in_120), .Y(n17103));
CLKBUFX1 gbuf_d_121(.A(n6195), .Y(d_out_121));
CLKBUFX1 gbuf_qn_121(.A(qn_in_121), .Y(n17105));
CLKBUFX1 gbuf_d_122(.A(n6196), .Y(d_out_122));
CLKBUFX1 gbuf_qn_122(.A(qn_in_122), .Y(n17107));
CLKBUFX1 gbuf_d_123(.A(n6197), .Y(d_out_123));
CLKBUFX1 gbuf_qn_123(.A(qn_in_123), .Y(n17109));
CLKBUFX1 gbuf_d_124(.A(n6198), .Y(d_out_124));
CLKBUFX1 gbuf_qn_124(.A(qn_in_124), .Y(n17111));
CLKBUFX1 gbuf_d_125(.A(n6199), .Y(d_out_125));
CLKBUFX1 gbuf_qn_125(.A(qn_in_125), .Y(n17113));
CLKBUFX1 gbuf_d_126(.A(n6200), .Y(d_out_126));
CLKBUFX1 gbuf_qn_126(.A(qn_in_126), .Y(n17115));
CLKBUFX1 gbuf_d_127(.A(n6201), .Y(d_out_127));
CLKBUFX1 gbuf_qn_127(.A(qn_in_127), .Y(n17117));
CLKBUFX1 gbuf_d_128(.A(n6202), .Y(d_out_128));
CLKBUFX1 gbuf_qn_128(.A(qn_in_128), .Y(n17119));
CLKBUFX1 gbuf_d_129(.A(n6203), .Y(d_out_129));
CLKBUFX1 gbuf_qn_129(.A(qn_in_129), .Y(n17121));
CLKBUFX1 gbuf_d_130(.A(n6204), .Y(d_out_130));
CLKBUFX1 gbuf_qn_130(.A(qn_in_130), .Y(n17123));
CLKBUFX1 gbuf_d_131(.A(n6205), .Y(d_out_131));
CLKBUFX1 gbuf_qn_131(.A(qn_in_131), .Y(n17125));
CLKBUFX1 gbuf_d_132(.A(n6206), .Y(d_out_132));
CLKBUFX1 gbuf_qn_132(.A(qn_in_132), .Y(n17127));
CLKBUFX1 gbuf_d_133(.A(n6207), .Y(d_out_133));
CLKBUFX1 gbuf_qn_133(.A(qn_in_133), .Y(n17129));
CLKBUFX1 gbuf_d_134(.A(n6208), .Y(d_out_134));
CLKBUFX1 gbuf_qn_134(.A(qn_in_134), .Y(n17131));
CLKBUFX1 gbuf_d_135(.A(n6209), .Y(d_out_135));
CLKBUFX1 gbuf_qn_135(.A(qn_in_135), .Y(n17133));
CLKBUFX1 gbuf_d_136(.A(n6210), .Y(d_out_136));
CLKBUFX1 gbuf_qn_136(.A(qn_in_136), .Y(n17135));
CLKBUFX1 gbuf_d_137(.A(n6211), .Y(d_out_137));
CLKBUFX1 gbuf_qn_137(.A(qn_in_137), .Y(n17137));
CLKBUFX1 gbuf_d_138(.A(n6212), .Y(d_out_138));
CLKBUFX1 gbuf_qn_138(.A(qn_in_138), .Y(n17139));
CLKBUFX1 gbuf_d_139(.A(n6213), .Y(d_out_139));
CLKBUFX1 gbuf_qn_139(.A(qn_in_139), .Y(n17141));
CLKBUFX1 gbuf_d_140(.A(n6214), .Y(d_out_140));
CLKBUFX1 gbuf_qn_140(.A(qn_in_140), .Y(n17143));
CLKBUFX1 gbuf_d_141(.A(n6215), .Y(d_out_141));
CLKBUFX1 gbuf_qn_141(.A(qn_in_141), .Y(n17145));
CLKBUFX1 gbuf_d_142(.A(n6216), .Y(d_out_142));
CLKBUFX1 gbuf_qn_142(.A(qn_in_142), .Y(n17147));
CLKBUFX1 gbuf_d_143(.A(n6217), .Y(d_out_143));
CLKBUFX1 gbuf_qn_143(.A(qn_in_143), .Y(n17149));
CLKBUFX1 gbuf_d_144(.A(n6218), .Y(d_out_144));
CLKBUFX1 gbuf_qn_144(.A(qn_in_144), .Y(n17151));
CLKBUFX1 gbuf_d_145(.A(n6219), .Y(d_out_145));
CLKBUFX1 gbuf_qn_145(.A(qn_in_145), .Y(n17153));
CLKBUFX1 gbuf_d_146(.A(n6220), .Y(d_out_146));
CLKBUFX1 gbuf_qn_146(.A(qn_in_146), .Y(n17155));
CLKBUFX1 gbuf_d_147(.A(n6221), .Y(d_out_147));
CLKBUFX1 gbuf_qn_147(.A(qn_in_147), .Y(n17157));
CLKBUFX1 gbuf_d_148(.A(n6222), .Y(d_out_148));
CLKBUFX1 gbuf_qn_148(.A(qn_in_148), .Y(n17159));
CLKBUFX1 gbuf_d_149(.A(n6223), .Y(d_out_149));
CLKBUFX1 gbuf_qn_149(.A(qn_in_149), .Y(n17161));
CLKBUFX1 gbuf_d_150(.A(n6224), .Y(d_out_150));
CLKBUFX1 gbuf_qn_150(.A(qn_in_150), .Y(n17163));
CLKBUFX1 gbuf_d_151(.A(n6225), .Y(d_out_151));
CLKBUFX1 gbuf_qn_151(.A(qn_in_151), .Y(n17165));
CLKBUFX1 gbuf_d_152(.A(n6226), .Y(d_out_152));
CLKBUFX1 gbuf_qn_152(.A(qn_in_152), .Y(n17167));
CLKBUFX1 gbuf_d_153(.A(n6227), .Y(d_out_153));
CLKBUFX1 gbuf_qn_153(.A(qn_in_153), .Y(n17169));
CLKBUFX1 gbuf_d_154(.A(n6228), .Y(d_out_154));
CLKBUFX1 gbuf_qn_154(.A(qn_in_154), .Y(n17171));
CLKBUFX1 gbuf_d_155(.A(n6229), .Y(d_out_155));
CLKBUFX1 gbuf_qn_155(.A(qn_in_155), .Y(n17173));
CLKBUFX1 gbuf_d_156(.A(n6230), .Y(d_out_156));
CLKBUFX1 gbuf_qn_156(.A(qn_in_156), .Y(n17175));
CLKBUFX1 gbuf_d_157(.A(n6231), .Y(d_out_157));
CLKBUFX1 gbuf_qn_157(.A(qn_in_157), .Y(n17177));
CLKBUFX1 gbuf_d_158(.A(n6239), .Y(d_out_158));
CLKBUFX1 gbuf_qn_158(.A(qn_in_158), .Y(n17193));
CLKBUFX1 gbuf_d_159(.A(n6244), .Y(d_out_159));
CLKBUFX1 gbuf_qn_159(.A(qn_in_159), .Y(n17203));
CLKBUFX1 gbuf_d_160(.A(n6245), .Y(d_out_160));
CLKBUFX1 gbuf_qn_160(.A(qn_in_160), .Y(n17205));
CLKBUFX1 gbuf_d_161(.A(n6246), .Y(d_out_161));
CLKBUFX1 gbuf_qn_161(.A(qn_in_161), .Y(n17207));
CLKBUFX1 gbuf_d_162(.A(n6247), .Y(d_out_162));
CLKBUFX1 gbuf_qn_162(.A(qn_in_162), .Y(n17209));
CLKBUFX1 gbuf_d_163(.A(n6248), .Y(d_out_163));
CLKBUFX1 gbuf_qn_163(.A(qn_in_163), .Y(n17211));
CLKBUFX1 gbuf_d_164(.A(n6249), .Y(d_out_164));
CLKBUFX1 gbuf_qn_164(.A(qn_in_164), .Y(n17213));
CLKBUFX1 gbuf_d_165(.A(n6250), .Y(d_out_165));
CLKBUFX1 gbuf_qn_165(.A(qn_in_165), .Y(n17215));
CLKBUFX1 gbuf_d_166(.A(n6251), .Y(d_out_166));
CLKBUFX1 gbuf_qn_166(.A(qn_in_166), .Y(n17217));
CLKBUFX1 gbuf_d_167(.A(n6252), .Y(d_out_167));
CLKBUFX1 gbuf_qn_167(.A(qn_in_167), .Y(n17219));
CLKBUFX1 gbuf_d_168(.A(n6253), .Y(d_out_168));
CLKBUFX1 gbuf_qn_168(.A(qn_in_168), .Y(n17221));
CLKBUFX1 gbuf_d_169(.A(n6254), .Y(d_out_169));
CLKBUFX1 gbuf_qn_169(.A(qn_in_169), .Y(n17223));
CLKBUFX1 gbuf_d_170(.A(n6255), .Y(d_out_170));
CLKBUFX1 gbuf_qn_170(.A(qn_in_170), .Y(n17225));
CLKBUFX1 gbuf_d_171(.A(n6256), .Y(d_out_171));
CLKBUFX1 gbuf_qn_171(.A(qn_in_171), .Y(n17227));
CLKBUFX1 gbuf_d_172(.A(n6257), .Y(d_out_172));
CLKBUFX1 gbuf_qn_172(.A(qn_in_172), .Y(n17229));
CLKBUFX1 gbuf_d_173(.A(n6258), .Y(d_out_173));
CLKBUFX1 gbuf_qn_173(.A(qn_in_173), .Y(n17231));
CLKBUFX1 gbuf_d_174(.A(n6259), .Y(d_out_174));
CLKBUFX1 gbuf_qn_174(.A(qn_in_174), .Y(n17233));
CLKBUFX1 gbuf_d_175(.A(n6262), .Y(d_out_175));
CLKBUFX1 gbuf_qn_175(.A(qn_in_175), .Y(n17239));
CLKBUFX1 gbuf_d_176(.A(n6265), .Y(d_out_176));
CLKBUFX1 gbuf_qn_176(.A(qn_in_176), .Y(n17245));
CLKBUFX1 gbuf_d_177(.A(n6266), .Y(d_out_177));
CLKBUFX1 gbuf_qn_177(.A(qn_in_177), .Y(n17247));
CLKBUFX1 gbuf_d_178(.A(n6267), .Y(d_out_178));
CLKBUFX1 gbuf_qn_178(.A(qn_in_178), .Y(n17249));
CLKBUFX1 gbuf_d_179(.A(n6268), .Y(d_out_179));
CLKBUFX1 gbuf_qn_179(.A(qn_in_179), .Y(n17251));
CLKBUFX1 gbuf_d_180(.A(n6269), .Y(d_out_180));
CLKBUFX1 gbuf_qn_180(.A(qn_in_180), .Y(n17253));
CLKBUFX1 gbuf_d_181(.A(n6270), .Y(d_out_181));
CLKBUFX1 gbuf_qn_181(.A(qn_in_181), .Y(n17255));
CLKBUFX1 gbuf_d_182(.A(n6271), .Y(d_out_182));
CLKBUFX1 gbuf_qn_182(.A(qn_in_182), .Y(n17257));
CLKBUFX1 gbuf_d_183(.A(n6272), .Y(d_out_183));
CLKBUFX1 gbuf_qn_183(.A(qn_in_183), .Y(n17259));
CLKBUFX1 gbuf_d_184(.A(n6273), .Y(d_out_184));
CLKBUFX1 gbuf_qn_184(.A(qn_in_184), .Y(n17261));
CLKBUFX1 gbuf_d_185(.A(n6274), .Y(d_out_185));
CLKBUFX1 gbuf_qn_185(.A(qn_in_185), .Y(n17263));
CLKBUFX1 gbuf_d_186(.A(n6275), .Y(d_out_186));
CLKBUFX1 gbuf_qn_186(.A(qn_in_186), .Y(n17265));
CLKBUFX1 gbuf_d_187(.A(n6276), .Y(d_out_187));
CLKBUFX1 gbuf_qn_187(.A(qn_in_187), .Y(n17267));
CLKBUFX1 gbuf_d_188(.A(n6277), .Y(d_out_188));
CLKBUFX1 gbuf_qn_188(.A(qn_in_188), .Y(n17269));
CLKBUFX1 gbuf_d_189(.A(n6278), .Y(d_out_189));
CLKBUFX1 gbuf_qn_189(.A(qn_in_189), .Y(n17271));
CLKBUFX1 gbuf_d_190(.A(n6279), .Y(d_out_190));
CLKBUFX1 gbuf_qn_190(.A(qn_in_190), .Y(n17273));
CLKBUFX1 gbuf_d_191(.A(n6282), .Y(d_out_191));
CLKBUFX1 gbuf_qn_191(.A(qn_in_191), .Y(n17279));
CLKBUFX1 gbuf_d_1(.A(n17744), .Y(ddout__1));
CLKBUFX1 gbuf_q_1(.A(qq_in1), .Y(n18197));
CLKBUFX1 gbuf_qn_1(.A(qnn_in_1), .Y(n5473));
CLKBUFX1 gbuf_d_2(.A(n5956), .Y(ddout__2));
CLKBUFX1 gbuf_q_2(.A(qq_in2), .Y(n18589));
CLKBUFX1 gbuf_qn_2(.A(qnn_in_2), .Y(n5571));
CLKBUFX1 gbuf_d_3(.A(n5955), .Y(ddout__3));
CLKBUFX1 gbuf_q_3(.A(qq_in3), .Y(n18585));
CLKBUFX1 gbuf_qn_3(.A(qnn_in_3), .Y(n5570));
CLKBUFX1 gbuf_d_4(.A(n5954), .Y(ddout__4));
CLKBUFX1 gbuf_q_4(.A(qq_in4), .Y(n18581));
CLKBUFX1 gbuf_qn_4(.A(qnn_in_4), .Y(n5569));
CLKBUFX1 gbuf_d_5(.A(n5953), .Y(ddout__5));
CLKBUFX1 gbuf_q_5(.A(qq_in5), .Y(n18577));
CLKBUFX1 gbuf_qn_5(.A(qnn_in_5), .Y(n5568));
CLKBUFX1 gbuf_d_6(.A(n5952), .Y(ddout__6));
CLKBUFX1 gbuf_q_6(.A(qq_in6), .Y(n18573));
CLKBUFX1 gbuf_qn_6(.A(qnn_in_6), .Y(n5567));
CLKBUFX1 gbuf_d_7(.A(n5951), .Y(ddout__7));
CLKBUFX1 gbuf_q_7(.A(qq_in7), .Y(n18569));
CLKBUFX1 gbuf_qn_7(.A(qnn_in_7), .Y(n5566));
CLKBUFX1 gbuf_d_8(.A(n5950), .Y(ddout__8));
CLKBUFX1 gbuf_q_8(.A(qq_in8), .Y(n18565));
CLKBUFX1 gbuf_qn_8(.A(qnn_in_8), .Y(n5565));
CLKBUFX1 gbuf_d_9(.A(n5949), .Y(ddout__9));
CLKBUFX1 gbuf_q_9(.A(qq_in9), .Y(n18561));
CLKBUFX1 gbuf_qn_9(.A(qnn_in_9), .Y(n5564));
CLKBUFX1 gbuf_d_10(.A(n5948), .Y(ddout__10));
CLKBUFX1 gbuf_q_10(.A(qq_in10), .Y(n18557));
CLKBUFX1 gbuf_qn_10(.A(qnn_in_10), .Y(n5563));
CLKBUFX1 gbuf_d_11(.A(n5947), .Y(ddout__11));
CLKBUFX1 gbuf_q_11(.A(qq_in11), .Y(n18553));
CLKBUFX1 gbuf_qn_11(.A(qnn_in_11), .Y(n5562));
CLKBUFX1 gbuf_d_12(.A(n5946), .Y(ddout__12));
CLKBUFX1 gbuf_q_12(.A(qq_in12), .Y(n18549));
CLKBUFX1 gbuf_qn_12(.A(qnn_in_12), .Y(n5561));
CLKBUFX1 gbuf_d_13(.A(n5945), .Y(ddout__13));
CLKBUFX1 gbuf_q_13(.A(qq_in13), .Y(n18545));
CLKBUFX1 gbuf_qn_13(.A(qnn_in_13), .Y(n5560));
CLKBUFX1 gbuf_d_14(.A(n5944), .Y(ddout__14));
CLKBUFX1 gbuf_q_14(.A(qq_in14), .Y(n18541));
CLKBUFX1 gbuf_qn_14(.A(qnn_in_14), .Y(n5559));
CLKBUFX1 gbuf_d_15(.A(n5943), .Y(ddout__15));
CLKBUFX1 gbuf_q_15(.A(qq_in15), .Y(n18537));
CLKBUFX1 gbuf_qn_15(.A(qnn_in_15), .Y(n5558));
CLKBUFX1 gbuf_d_16(.A(n5942), .Y(ddout__16));
CLKBUFX1 gbuf_q_16(.A(qq_in16), .Y(n18533));
CLKBUFX1 gbuf_qn_16(.A(qnn_in_16), .Y(n5557));
CLKBUFX1 gbuf_d_17(.A(n5941), .Y(ddout__17));
CLKBUFX1 gbuf_q_17(.A(qq_in17), .Y(n18529));
CLKBUFX1 gbuf_qn_17(.A(qnn_in_17), .Y(n5556));
CLKBUFX1 gbuf_d_18(.A(n17726), .Y(ddout__18));
CLKBUFX1 gbuf_q_18(.A(qq_in18), .Y(n18525));
CLKBUFX1 gbuf_qn_18(.A(qnn_in_18), .Y(n5555));
CLKBUFX1 gbuf_d_19(.A(n17724), .Y(ddout__19));
CLKBUFX1 gbuf_q_19(.A(qq_in19), .Y(n18521));
CLKBUFX1 gbuf_qn_19(.A(qnn_in_19), .Y(n5554));
CLKBUFX1 gbuf_d_20(.A(n17722), .Y(ddout__20));
CLKBUFX1 gbuf_q_20(.A(qq_in20), .Y(n18517));
CLKBUFX1 gbuf_qn_20(.A(qnn_in_20), .Y(n5553));
CLKBUFX1 gbuf_d_21(.A(n17720), .Y(ddout__21));
CLKBUFX1 gbuf_q_21(.A(qq_in21), .Y(n18513));
CLKBUFX1 gbuf_qn_21(.A(qnn_in_21), .Y(n5552));
CLKBUFX1 gbuf_d_22(.A(n17718), .Y(ddout__22));
CLKBUFX1 gbuf_q_22(.A(qq_in22), .Y(n18509));
CLKBUFX1 gbuf_qn_22(.A(qnn_in_22), .Y(n5551));
CLKBUFX1 gbuf_d_23(.A(n17716), .Y(ddout__23));
CLKBUFX1 gbuf_q_23(.A(qq_in23), .Y(n18505));
CLKBUFX1 gbuf_qn_23(.A(qnn_in_23), .Y(n5550));
CLKBUFX1 gbuf_d_24(.A(n17714), .Y(ddout__24));
CLKBUFX1 gbuf_q_24(.A(qq_in24), .Y(n18501));
CLKBUFX1 gbuf_qn_24(.A(qnn_in_24), .Y(n5549));
CLKBUFX1 gbuf_d_25(.A(n17712), .Y(ddout__25));
CLKBUFX1 gbuf_q_25(.A(qq_in25), .Y(n18497));
CLKBUFX1 gbuf_qn_25(.A(qnn_in_25), .Y(n5548));
CLKBUFX1 gbuf_d_26(.A(n17710), .Y(ddout__26));
CLKBUFX1 gbuf_q_26(.A(qq_in26), .Y(n18493));
CLKBUFX1 gbuf_qn_26(.A(qnn_in_26), .Y(n5547));
CLKBUFX1 gbuf_d_27(.A(n17708), .Y(ddout__27));
CLKBUFX1 gbuf_q_27(.A(qq_in27), .Y(n18489));
CLKBUFX1 gbuf_qn_27(.A(qnn_in_27), .Y(n5546));
CLKBUFX1 gbuf_d_28(.A(n17706), .Y(ddout__28));
CLKBUFX1 gbuf_q_28(.A(qq_in28), .Y(n18485));
CLKBUFX1 gbuf_qn_28(.A(qnn_in_28), .Y(n5545));
CLKBUFX1 gbuf_d_29(.A(n17704), .Y(ddout__29));
CLKBUFX1 gbuf_q_29(.A(qq_in29), .Y(n18481));
CLKBUFX1 gbuf_qn_29(.A(qnn_in_29), .Y(n5544));
CLKBUFX1 gbuf_d_30(.A(n17702), .Y(ddout__30));
CLKBUFX1 gbuf_q_30(.A(qq_in30), .Y(n18477));
CLKBUFX1 gbuf_qn_30(.A(qnn_in_30), .Y(n5543));
CLKBUFX1 gbuf_d_31(.A(n17700), .Y(ddout__31));
CLKBUFX1 gbuf_q_31(.A(qq_in31), .Y(n18473));
CLKBUFX1 gbuf_qn_31(.A(qnn_in_31), .Y(n5542));
CLKBUFX1 gbuf_d_32(.A(n17698), .Y(ddout__32));
CLKBUFX1 gbuf_q_32(.A(qq_in32), .Y(n18469));
CLKBUFX1 gbuf_qn_32(.A(qnn_in_32), .Y(n5541));
CLKBUFX1 gbuf_d_33(.A(n17696), .Y(ddout__33));
CLKBUFX1 gbuf_q_33(.A(qq_in33), .Y(n18465));
CLKBUFX1 gbuf_qn_33(.A(qnn_in_33), .Y(n5540));
CLKBUFX1 gbuf_d_34(.A(n17694), .Y(ddout__34));
CLKBUFX1 gbuf_q_34(.A(qq_in34), .Y(n18461));
CLKBUFX1 gbuf_qn_34(.A(qnn_in_34), .Y(n5539));
CLKBUFX1 gbuf_d_35(.A(n17692), .Y(ddout__35));
CLKBUFX1 gbuf_q_35(.A(qq_in35), .Y(n18457));
CLKBUFX1 gbuf_qn_35(.A(qnn_in_35), .Y(n5538));
CLKBUFX1 gbuf_d_36(.A(n17690), .Y(ddout__36));
CLKBUFX1 gbuf_q_36(.A(qq_in36), .Y(n18453));
CLKBUFX1 gbuf_qn_36(.A(qnn_in_36), .Y(n5537));
CLKBUFX1 gbuf_d_37(.A(n17688), .Y(ddout__37));
CLKBUFX1 gbuf_q_37(.A(qq_in37), .Y(n18449));
CLKBUFX1 gbuf_qn_37(.A(qnn_in_37), .Y(n5536));
CLKBUFX1 gbuf_d_38(.A(n17686), .Y(ddout__38));
CLKBUFX1 gbuf_q_38(.A(qq_in38), .Y(n18445));
CLKBUFX1 gbuf_qn_38(.A(qnn_in_38), .Y(n5535));
CLKBUFX1 gbuf_d_39(.A(n17684), .Y(ddout__39));
CLKBUFX1 gbuf_q_39(.A(qq_in39), .Y(n18441));
CLKBUFX1 gbuf_qn_39(.A(qnn_in_39), .Y(n5534));
CLKBUFX1 gbuf_d_40(.A(n17682), .Y(ddout__40));
CLKBUFX1 gbuf_q_40(.A(qq_in40), .Y(n18437));
CLKBUFX1 gbuf_qn_40(.A(qnn_in_40), .Y(n5533));
CLKBUFX1 gbuf_d_41(.A(n17680), .Y(ddout__41));
CLKBUFX1 gbuf_q_41(.A(qq_in41), .Y(n18433));
CLKBUFX1 gbuf_qn_41(.A(qnn_in_41), .Y(n5532));
CLKBUFX1 gbuf_d_42(.A(n17678), .Y(ddout__42));
CLKBUFX1 gbuf_q_42(.A(qq_in42), .Y(n18429));
CLKBUFX1 gbuf_qn_42(.A(qnn_in_42), .Y(n5531));
CLKBUFX1 gbuf_d_43(.A(n17676), .Y(ddout__43));
CLKBUFX1 gbuf_q_43(.A(qq_in43), .Y(n18425));
CLKBUFX1 gbuf_qn_43(.A(qnn_in_43), .Y(n5530));
CLKBUFX1 gbuf_d_44(.A(n17674), .Y(ddout__44));
CLKBUFX1 gbuf_q_44(.A(qq_in44), .Y(n18421));
CLKBUFX1 gbuf_qn_44(.A(qnn_in_44), .Y(n5529));
CLKBUFX1 gbuf_d_45(.A(n17672), .Y(ddout__45));
CLKBUFX1 gbuf_q_45(.A(qq_in45), .Y(n18417));
CLKBUFX1 gbuf_qn_45(.A(qnn_in_45), .Y(n5528));
CLKBUFX1 gbuf_d_46(.A(n17670), .Y(ddout__46));
CLKBUFX1 gbuf_q_46(.A(qq_in46), .Y(n18413));
CLKBUFX1 gbuf_qn_46(.A(qnn_in_46), .Y(n5527));
CLKBUFX1 gbuf_d_47(.A(n17668), .Y(ddout__47));
CLKBUFX1 gbuf_q_47(.A(qq_in47), .Y(n18409));
CLKBUFX1 gbuf_qn_47(.A(qnn_in_47), .Y(n5526));
CLKBUFX1 gbuf_d_48(.A(n17666), .Y(ddout__48));
CLKBUFX1 gbuf_q_48(.A(qq_in48), .Y(n18405));
CLKBUFX1 gbuf_qn_48(.A(qnn_in_48), .Y(n5525));
CLKBUFX1 gbuf_d_49(.A(n17664), .Y(ddout__49));
CLKBUFX1 gbuf_q_49(.A(qq_in49), .Y(n18401));
CLKBUFX1 gbuf_qn_49(.A(qnn_in_49), .Y(n5524));
CLKBUFX1 gbuf_d_50(.A(n17662), .Y(ddout__50));
CLKBUFX1 gbuf_q_50(.A(qq_in50), .Y(n18397));
CLKBUFX1 gbuf_qn_50(.A(qnn_in_50), .Y(n5523));
CLKBUFX1 gbuf_d_51(.A(n17660), .Y(ddout__51));
CLKBUFX1 gbuf_q_51(.A(qq_in51), .Y(n18393));
CLKBUFX1 gbuf_qn_51(.A(qnn_in_51), .Y(n5522));
CLKBUFX1 gbuf_d_52(.A(n17658), .Y(ddout__52));
CLKBUFX1 gbuf_q_52(.A(qq_in52), .Y(n18389));
CLKBUFX1 gbuf_qn_52(.A(qnn_in_52), .Y(n5521));
CLKBUFX1 gbuf_d_53(.A(n17656), .Y(ddout__53));
CLKBUFX1 gbuf_q_53(.A(qq_in53), .Y(n18385));
CLKBUFX1 gbuf_qn_53(.A(qnn_in_53), .Y(n5520));
CLKBUFX1 gbuf_d_54(.A(n17654), .Y(ddout__54));
CLKBUFX1 gbuf_q_54(.A(qq_in54), .Y(n18381));
CLKBUFX1 gbuf_qn_54(.A(qnn_in_54), .Y(n5519));
CLKBUFX1 gbuf_d_55(.A(n17652), .Y(ddout__55));
CLKBUFX1 gbuf_q_55(.A(qq_in55), .Y(n18377));
CLKBUFX1 gbuf_qn_55(.A(qnn_in_55), .Y(n5518));
CLKBUFX1 gbuf_d_56(.A(n17650), .Y(ddout__56));
CLKBUFX1 gbuf_q_56(.A(qq_in56), .Y(n18373));
CLKBUFX1 gbuf_qn_56(.A(qnn_in_56), .Y(n5517));
CLKBUFX1 gbuf_d_57(.A(n17648), .Y(ddout__57));
CLKBUFX1 gbuf_q_57(.A(qq_in57), .Y(n18369));
CLKBUFX1 gbuf_qn_57(.A(qnn_in_57), .Y(n5516));
CLKBUFX1 gbuf_d_58(.A(n17646), .Y(ddout__58));
CLKBUFX1 gbuf_q_58(.A(qq_in58), .Y(n18365));
CLKBUFX1 gbuf_qn_58(.A(qnn_in_58), .Y(n5515));
CLKBUFX1 gbuf_d_59(.A(n17644), .Y(ddout__59));
CLKBUFX1 gbuf_q_59(.A(qq_in59), .Y(n18361));
CLKBUFX1 gbuf_qn_59(.A(qnn_in_59), .Y(n5514));
CLKBUFX1 gbuf_d_60(.A(n17642), .Y(ddout__60));
CLKBUFX1 gbuf_q_60(.A(qq_in60), .Y(n18357));
CLKBUFX1 gbuf_qn_60(.A(qnn_in_60), .Y(n5513));
CLKBUFX1 gbuf_d_61(.A(n17640), .Y(ddout__61));
CLKBUFX1 gbuf_q_61(.A(qq_in61), .Y(n18353));
CLKBUFX1 gbuf_qn_61(.A(qnn_in_61), .Y(n5512));
CLKBUFX1 gbuf_d_62(.A(n17638), .Y(ddout__62));
CLKBUFX1 gbuf_q_62(.A(qq_in62), .Y(n18349));
CLKBUFX1 gbuf_qn_62(.A(qnn_in_62), .Y(n5511));
CLKBUFX1 gbuf_d_63(.A(n17636), .Y(ddout__63));
CLKBUFX1 gbuf_q_63(.A(qq_in63), .Y(n18345));
CLKBUFX1 gbuf_qn_63(.A(qnn_in_63), .Y(n5510));
CLKBUFX1 gbuf_d_64(.A(n17634), .Y(ddout__64));
CLKBUFX1 gbuf_q_64(.A(qq_in64), .Y(n18341));
CLKBUFX1 gbuf_qn_64(.A(qnn_in_64), .Y(n5509));
CLKBUFX1 gbuf_d_65(.A(n17632), .Y(ddout__65));
CLKBUFX1 gbuf_q_65(.A(qq_in65), .Y(n18337));
CLKBUFX1 gbuf_qn_65(.A(qnn_in_65), .Y(n5508));
CLKBUFX1 gbuf_d_66(.A(n17630), .Y(ddout__66));
CLKBUFX1 gbuf_q_66(.A(qq_in66), .Y(n18333));
CLKBUFX1 gbuf_qn_66(.A(qnn_in_66), .Y(n5507));
CLKBUFX1 gbuf_d_67(.A(n17628), .Y(ddout__67));
CLKBUFX1 gbuf_q_67(.A(qq_in67), .Y(n18329));
CLKBUFX1 gbuf_qn_67(.A(qnn_in_67), .Y(n5506));
CLKBUFX1 gbuf_d_68(.A(n17626), .Y(ddout__68));
CLKBUFX1 gbuf_q_68(.A(qq_in68), .Y(n18325));
CLKBUFX1 gbuf_qn_68(.A(qnn_in_68), .Y(n5505));
CLKBUFX1 gbuf_d_69(.A(n5889), .Y(ddout__69));
CLKBUFX1 gbuf_q_69(.A(qq_in69), .Y(n18321));
CLKBUFX1 gbuf_qn_69(.A(qnn_in_69), .Y(n5504));
CLKBUFX1 gbuf_d_70(.A(n5888), .Y(ddout__70));
CLKBUFX1 gbuf_q_70(.A(qq_in70), .Y(n18317));
CLKBUFX1 gbuf_qn_70(.A(qnn_in_70), .Y(n5503));
CLKBUFX1 gbuf_d_71(.A(n5887), .Y(ddout__71));
CLKBUFX1 gbuf_q_71(.A(qq_in71), .Y(n18313));
CLKBUFX1 gbuf_qn_71(.A(qnn_in_71), .Y(n5502));
CLKBUFX1 gbuf_d_72(.A(n5886), .Y(ddout__72));
CLKBUFX1 gbuf_q_72(.A(qq_in72), .Y(n18309));
CLKBUFX1 gbuf_qn_72(.A(qnn_in_72), .Y(n5501));
CLKBUFX1 gbuf_d_73(.A(n5885), .Y(ddout__73));
CLKBUFX1 gbuf_q_73(.A(qq_in73), .Y(n18305));
CLKBUFX1 gbuf_qn_73(.A(qnn_in_73), .Y(n5500));
CLKBUFX1 gbuf_d_74(.A(n17614), .Y(ddout__74));
CLKBUFX1 gbuf_q_74(.A(qq_in74), .Y(n18301));
CLKBUFX1 gbuf_qn_74(.A(qnn_in_74), .Y(n5499));
CLKBUFX1 gbuf_d_75(.A(n17612), .Y(ddout__75));
CLKBUFX1 gbuf_q_75(.A(qq_in75), .Y(n18297));
CLKBUFX1 gbuf_qn_75(.A(qnn_in_75), .Y(n5498));
CLKBUFX1 gbuf_d_76(.A(n17610), .Y(ddout__76));
CLKBUFX1 gbuf_q_76(.A(qq_in76), .Y(n18293));
CLKBUFX1 gbuf_qn_76(.A(qnn_in_76), .Y(n5497));
CLKBUFX1 gbuf_d_77(.A(n17608), .Y(ddout__77));
CLKBUFX1 gbuf_q_77(.A(qq_in77), .Y(n18289));
CLKBUFX1 gbuf_qn_77(.A(qnn_in_77), .Y(n5496));
CLKBUFX1 gbuf_d_78(.A(n17606), .Y(ddout__78));
CLKBUFX1 gbuf_q_78(.A(qq_in78), .Y(n18285));
CLKBUFX1 gbuf_qn_78(.A(qnn_in_78), .Y(n5495));
CLKBUFX1 gbuf_d_79(.A(n17604), .Y(ddout__79));
CLKBUFX1 gbuf_q_79(.A(qq_in79), .Y(n18281));
CLKBUFX1 gbuf_qn_79(.A(qnn_in_79), .Y(n5494));
CLKBUFX1 gbuf_d_80(.A(n17602), .Y(ddout__80));
CLKBUFX1 gbuf_q_80(.A(qq_in80), .Y(n18277));
CLKBUFX1 gbuf_qn_80(.A(qnn_in_80), .Y(n5493));
CLKBUFX1 gbuf_d_81(.A(n17600), .Y(ddout__81));
CLKBUFX1 gbuf_q_81(.A(qq_in81), .Y(n18273));
CLKBUFX1 gbuf_qn_81(.A(qnn_in_81), .Y(n5492));
CLKBUFX1 gbuf_d_82(.A(n17598), .Y(ddout__82));
CLKBUFX1 gbuf_q_82(.A(qq_in82), .Y(n18269));
CLKBUFX1 gbuf_qn_82(.A(qnn_in_82), .Y(n5491));
CLKBUFX1 gbuf_d_83(.A(n17596), .Y(ddout__83));
CLKBUFX1 gbuf_q_83(.A(qq_in83), .Y(n18265));
CLKBUFX1 gbuf_qn_83(.A(qnn_in_83), .Y(n5490));
CLKBUFX1 gbuf_d_84(.A(n17594), .Y(ddout__84));
CLKBUFX1 gbuf_q_84(.A(qq_in84), .Y(n18261));
CLKBUFX1 gbuf_qn_84(.A(qnn_in_84), .Y(n5489));
CLKBUFX1 gbuf_d_85(.A(n17592), .Y(ddout__85));
CLKBUFX1 gbuf_q_85(.A(qq_in85), .Y(n18257));
CLKBUFX1 gbuf_qn_85(.A(qnn_in_85), .Y(n5488));
CLKBUFX1 gbuf_d_86(.A(n17590), .Y(ddout__86));
CLKBUFX1 gbuf_q_86(.A(qq_in86), .Y(n18253));
CLKBUFX1 gbuf_qn_86(.A(qnn_in_86), .Y(n5487));
CLKBUFX1 gbuf_d_87(.A(n17588), .Y(ddout__87));
CLKBUFX1 gbuf_q_87(.A(qq_in87), .Y(n18249));
CLKBUFX1 gbuf_qn_87(.A(qnn_in_87), .Y(n5486));
CLKBUFX1 gbuf_d_88(.A(n17586), .Y(ddout__88));
CLKBUFX1 gbuf_q_88(.A(qq_in88), .Y(n18245));
CLKBUFX1 gbuf_qn_88(.A(qnn_in_88), .Y(n5485));
CLKBUFX1 gbuf_d_89(.A(n17584), .Y(ddout__89));
CLKBUFX1 gbuf_q_89(.A(qq_in89), .Y(n18241));
CLKBUFX1 gbuf_qn_89(.A(qnn_in_89), .Y(n5484));
CLKBUFX1 gbuf_d_90(.A(n17582), .Y(ddout__90));
CLKBUFX1 gbuf_q_90(.A(qq_in90), .Y(n18237));
CLKBUFX1 gbuf_qn_90(.A(qnn_in_90), .Y(n5483));
CLKBUFX1 gbuf_d_91(.A(n17580), .Y(ddout__91));
CLKBUFX1 gbuf_q_91(.A(qq_in91), .Y(n18233));
CLKBUFX1 gbuf_qn_91(.A(qnn_in_91), .Y(n5482));
CLKBUFX1 gbuf_d_92(.A(n17578), .Y(ddout__92));
CLKBUFX1 gbuf_q_92(.A(qq_in92), .Y(n18229));
CLKBUFX1 gbuf_qn_92(.A(qnn_in_92), .Y(n5481));
CLKBUFX1 gbuf_d_93(.A(n17576), .Y(ddout__93));
CLKBUFX1 gbuf_q_93(.A(qq_in93), .Y(n18225));
CLKBUFX1 gbuf_qn_93(.A(qnn_in_93), .Y(n5480));
CLKBUFX1 gbuf_d_94(.A(n17574), .Y(ddout__94));
CLKBUFX1 gbuf_q_94(.A(qq_in94), .Y(n18221));
CLKBUFX1 gbuf_qn_94(.A(qnn_in_94), .Y(n5479));
CLKBUFX1 gbuf_d_95(.A(n17572), .Y(ddout__95));
CLKBUFX1 gbuf_q_95(.A(qq_in95), .Y(n18217));
CLKBUFX1 gbuf_qn_95(.A(qnn_in_95), .Y(n5478));
CLKBUFX1 gbuf_d_96(.A(n17570), .Y(ddout__96));
CLKBUFX1 gbuf_q_96(.A(qq_in96), .Y(n18213));
CLKBUFX1 gbuf_qn_96(.A(qnn_in_96), .Y(n5477));
CLKBUFX1 gbuf_d_97(.A(n17568), .Y(ddout__97));
CLKBUFX1 gbuf_q_97(.A(qq_in97), .Y(n18209));
CLKBUFX1 gbuf_qn_97(.A(qnn_in_97), .Y(n5476));
CLKBUFX1 gbuf_d_98(.A(n17566), .Y(ddout__98));
CLKBUFX1 gbuf_q_98(.A(qq_in98), .Y(n18205));
CLKBUFX1 gbuf_qn_98(.A(qnn_in_98), .Y(n5475));
CLKBUFX1 gbuf_d_99(.A(n17564), .Y(ddout__99));
CLKBUFX1 gbuf_q_99(.A(qq_in99), .Y(n18201));
CLKBUFX1 gbuf_qn_99(.A(qnn_in_99), .Y(n5474));
CLKBUFX1 gbuf_d_100(.A(n17562), .Y(ddout__100));
CLKBUFX1 gbuf_q_100(.A(qq_in100), .Y(n18193));
CLKBUFX1 gbuf_qn_100(.A(qnn_in_100), .Y(n5472));
CLKBUFX1 gbuf_d_101(.A(n17560), .Y(ddout__101));
CLKBUFX1 gbuf_q_101(.A(qq_in101), .Y(n18189));
CLKBUFX1 gbuf_qn_101(.A(qnn_in_101), .Y(n5471));
CLKBUFX1 gbuf_d_102(.A(n17558), .Y(ddout__102));
CLKBUFX1 gbuf_q_102(.A(qq_in102), .Y(n18185));
CLKBUFX1 gbuf_qn_102(.A(qnn_in_102), .Y(n5470));
CLKBUFX1 gbuf_d_103(.A(n17556), .Y(ddout__103));
CLKBUFX1 gbuf_q_103(.A(qq_in103), .Y(n18181));
CLKBUFX1 gbuf_qn_103(.A(qnn_in_103), .Y(n5469));
CLKBUFX1 gbuf_d_104(.A(n17554), .Y(ddout__104));
CLKBUFX1 gbuf_q_104(.A(qq_in104), .Y(n18177));
CLKBUFX1 gbuf_qn_104(.A(qnn_in_104), .Y(n5468));
CLKBUFX1 gbuf_d_105(.A(n17552), .Y(ddout__105));
CLKBUFX1 gbuf_q_105(.A(qq_in105), .Y(n18173));
CLKBUFX1 gbuf_qn_105(.A(qnn_in_105), .Y(n5467));
CLKBUFX1 gbuf_d_106(.A(n17550), .Y(ddout__106));
CLKBUFX1 gbuf_q_106(.A(qq_in106), .Y(n18169));
CLKBUFX1 gbuf_qn_106(.A(qnn_in_106), .Y(n5466));
CLKBUFX1 gbuf_d_107(.A(n17548), .Y(ddout__107));
CLKBUFX1 gbuf_q_107(.A(qq_in107), .Y(n18165));
CLKBUFX1 gbuf_qn_107(.A(qnn_in_107), .Y(n5465));
CLKBUFX1 gbuf_d_108(.A(n17546), .Y(ddout__108));
CLKBUFX1 gbuf_q_108(.A(qq_in108), .Y(n18161));
CLKBUFX1 gbuf_qn_108(.A(qnn_in_108), .Y(n5464));
CLKBUFX1 gbuf_d_109(.A(n17544), .Y(ddout__109));
CLKBUFX1 gbuf_q_109(.A(qq_in109), .Y(n18157));
CLKBUFX1 gbuf_qn_109(.A(qnn_in_109), .Y(n5463));
CLKBUFX1 gbuf_d_110(.A(n17542), .Y(ddout__110));
CLKBUFX1 gbuf_q_110(.A(qq_in110), .Y(n18153));
CLKBUFX1 gbuf_qn_110(.A(qnn_in_110), .Y(n5462));
CLKBUFX1 gbuf_d_111(.A(n17540), .Y(ddout__111));
CLKBUFX1 gbuf_q_111(.A(qq_in111), .Y(n18149));
CLKBUFX1 gbuf_qn_111(.A(qnn_in_111), .Y(n5461));
CLKBUFX1 gbuf_d_112(.A(n17538), .Y(ddout__112));
CLKBUFX1 gbuf_q_112(.A(qq_in112), .Y(n18145));
CLKBUFX1 gbuf_qn_112(.A(qnn_in_112), .Y(n5460));
CLKBUFX1 gbuf_d_113(.A(n5845), .Y(ddout__113));
CLKBUFX1 gbuf_q_113(.A(qq_in113), .Y(n18141));
CLKBUFX1 gbuf_qn_113(.A(qnn_in_113), .Y(n5459));
CLKBUFX1 gbuf_d_114(.A(n5844), .Y(ddout__114));
CLKBUFX1 gbuf_q_114(.A(qq_in114), .Y(n18137));
CLKBUFX1 gbuf_qn_114(.A(qnn_in_114), .Y(n5458));
CLKBUFX1 gbuf_d_115(.A(n5843), .Y(ddout__115));
CLKBUFX1 gbuf_q_115(.A(qq_in115), .Y(n18133));
CLKBUFX1 gbuf_qn_115(.A(qnn_in_115), .Y(n5457));
CLKBUFX1 gbuf_d_116(.A(n5842), .Y(ddout__116));
CLKBUFX1 gbuf_q_116(.A(qq_in116), .Y(n18129));
CLKBUFX1 gbuf_qn_116(.A(qnn_in_116), .Y(n5456));
CLKBUFX1 gbuf_d_117(.A(n5841), .Y(ddout__117));
CLKBUFX1 gbuf_q_117(.A(qq_in117), .Y(n18125));
CLKBUFX1 gbuf_qn_117(.A(qnn_in_117), .Y(n5455));
CLKBUFX1 gbuf_d_118(.A(n5840), .Y(ddout__118));
CLKBUFX1 gbuf_q_118(.A(qq_in118), .Y(n18121));
CLKBUFX1 gbuf_qn_118(.A(qnn_in_118), .Y(n5454));
CLKBUFX1 gbuf_d_119(.A(n5839), .Y(ddout__119));
CLKBUFX1 gbuf_q_119(.A(qq_in119), .Y(n18117));
CLKBUFX1 gbuf_qn_119(.A(qnn_in_119), .Y(n5453));
CLKBUFX1 gbuf_d_120(.A(n5838), .Y(ddout__120));
CLKBUFX1 gbuf_q_120(.A(qq_in120), .Y(n18113));
CLKBUFX1 gbuf_qn_120(.A(qnn_in_120), .Y(n5452));
CLKBUFX1 gbuf_d_121(.A(n17521), .Y(ddout__121));
CLKBUFX1 gbuf_q_121(.A(qq_in121), .Y(n18109));
CLKBUFX1 gbuf_qn_121(.A(qnn_in_121), .Y(n5451));
CLKBUFX1 gbuf_d_122(.A(n17519), .Y(ddout__122));
CLKBUFX1 gbuf_q_122(.A(qq_in122), .Y(n18105));
CLKBUFX1 gbuf_qn_122(.A(qnn_in_122), .Y(n5450));
CLKBUFX1 gbuf_d_123(.A(n17517), .Y(ddout__123));
CLKBUFX1 gbuf_q_123(.A(qq_in123), .Y(n18101));
CLKBUFX1 gbuf_qn_123(.A(qnn_in_123), .Y(n5449));
CLKBUFX1 gbuf_d_124(.A(n17515), .Y(ddout__124));
CLKBUFX1 gbuf_q_124(.A(qq_in124), .Y(n18097));
CLKBUFX1 gbuf_qn_124(.A(qnn_in_124), .Y(n5448));
CLKBUFX1 gbuf_d_125(.A(n17513), .Y(ddout__125));
CLKBUFX1 gbuf_q_125(.A(qq_in125), .Y(n18093));
CLKBUFX1 gbuf_qn_125(.A(qnn_in_125), .Y(n5447));
CLKBUFX1 gbuf_d_126(.A(n17511), .Y(ddout__126));
CLKBUFX1 gbuf_q_126(.A(qq_in126), .Y(n18089));
CLKBUFX1 gbuf_qn_126(.A(qnn_in_126), .Y(n5446));
CLKBUFX1 gbuf_d_127(.A(n17509), .Y(ddout__127));
CLKBUFX1 gbuf_q_127(.A(qq_in127), .Y(n18082));
CLKBUFX1 gbuf_qn_127(.A(qnn_in_127), .Y(n5445));
CLKBUFX1 gbuf_d_128(.A(n17507), .Y(ddout__128));
CLKBUFX1 gbuf_q_128(.A(qq_in128), .Y(n18593));
CLKBUFX1 gbuf_qn_128(.A(qnn_in_128), .Y(n5444));
CLKBUFX1 gbuf_d_129(.A(n17847), .Y(ddout__129));
CLKBUFX1 gbuf_q_129(.A(qq_in129), .Y(Tag_vld));
CLKBUFX1 gbuf_d_130(.A(n17505), .Y(ddout__130));
CLKBUFX1 gbuf_q_130(.A(qq_in130), .Y(Out_vld));
CLKBUFX1 gbuf_d_131(.A(n6022), .Y(ddout__131));
CLKBUFX1 gbuf_q_131(.A(qq_in131), .Y(Out_last_word));
CLKBUFX1 gbuf_d_132(.A(n6023), .Y(ddout__132));
CLKBUFX1 gbuf_q_132(.A(qq_in132), .Y(Out_data_size[3]));
CLKBUFX1 gbuf_d_133(.A(n17504), .Y(ddout__133));
CLKBUFX1 gbuf_q_133(.A(qq_in133), .Y(Out_data_size[2]));
CLKBUFX1 gbuf_d_134(.A(n17503), .Y(ddout__134));
CLKBUFX1 gbuf_q_134(.A(qq_in134), .Y(Out_data_size[1]));
CLKBUFX1 gbuf_d_135(.A(n6026), .Y(ddout__135));
CLKBUFX1 gbuf_q_135(.A(qq_in135), .Y(Out_data_size[0]));
CLKBUFX1 gbuf_d_136(.A(n6295), .Y(ddout__136));
CLKBUFX1 gbuf_q_136(.A(qq_in136), .Y(n16839));
CLKBUFX1 gbuf_d_137(.A(N2815), .Y(ddout__137));
CLKBUFX1 gbuf_q_137(.A(qq_in137), .Y(v_in[0]));
CLKBUFX1 gbuf_d_138(.A(n5701), .Y(ddout__138));
CLKBUFX1 gbuf_q_138(.A(qq_in138), .Y(Out_data[0]));
CLKBUFX1 gbuf_d_139(.A(N3071), .Y(ddout__139));
CLKBUFX1 gbuf_q_139(.A(qq_in139), .Y(b_in[0]));
CLKBUFX1 gbuf_d_140(.A(N2943), .Y(ddout__140));
CLKBUFX1 gbuf_q_140(.A(qq_in140), .Y(z_in[0]));
CLKBUFX1 gbuf_d_141(.A(n5700), .Y(ddout__141));
CLKBUFX1 gbuf_q_141(.A(qq_in141), .Y(Out_data[1]));
CLKBUFX1 gbuf_d_142(.A(N3072), .Y(ddout__142));
CLKBUFX1 gbuf_q_142(.A(qq_in142), .Y(b_in[1]));
CLKBUFX1 gbuf_d_143(.A(N2944), .Y(ddout__143));
CLKBUFX1 gbuf_q_143(.A(qq_in143), .Y(z_in[1]));
CLKBUFX1 gbuf_d_144(.A(n5699), .Y(ddout__144));
CLKBUFX1 gbuf_q_144(.A(qq_in144), .Y(Out_data[2]));
CLKBUFX1 gbuf_d_145(.A(N3073), .Y(ddout__145));
CLKBUFX1 gbuf_q_145(.A(qq_in145), .Y(b_in[2]));
CLKBUFX1 gbuf_d_146(.A(N2945), .Y(ddout__146));
CLKBUFX1 gbuf_q_146(.A(qq_in146), .Y(z_in[2]));
CLKBUFX1 gbuf_d_147(.A(n5698), .Y(ddout__147));
CLKBUFX1 gbuf_q_147(.A(qq_in147), .Y(Out_data[3]));
CLKBUFX1 gbuf_d_148(.A(N3074), .Y(ddout__148));
CLKBUFX1 gbuf_q_148(.A(qq_in148), .Y(b_in[3]));
CLKBUFX1 gbuf_d_149(.A(N2946), .Y(ddout__149));
CLKBUFX1 gbuf_q_149(.A(qq_in149), .Y(z_in[3]));
CLKBUFX1 gbuf_d_150(.A(n5697), .Y(ddout__150));
CLKBUFX1 gbuf_q_150(.A(qq_in150), .Y(Out_data[4]));
CLKBUFX1 gbuf_d_151(.A(N3075), .Y(ddout__151));
CLKBUFX1 gbuf_q_151(.A(qq_in151), .Y(b_in[4]));
CLKBUFX1 gbuf_d_152(.A(N2947), .Y(ddout__152));
CLKBUFX1 gbuf_q_152(.A(qq_in152), .Y(z_in[4]));
CLKBUFX1 gbuf_d_153(.A(n5696), .Y(ddout__153));
CLKBUFX1 gbuf_q_153(.A(qq_in153), .Y(Out_data[5]));
CLKBUFX1 gbuf_d_154(.A(N3076), .Y(ddout__154));
CLKBUFX1 gbuf_q_154(.A(qq_in154), .Y(b_in[5]));
CLKBUFX1 gbuf_d_155(.A(N2948), .Y(ddout__155));
CLKBUFX1 gbuf_q_155(.A(qq_in155), .Y(z_in[5]));
CLKBUFX1 gbuf_d_156(.A(n5695), .Y(ddout__156));
CLKBUFX1 gbuf_q_156(.A(qq_in156), .Y(Out_data[6]));
CLKBUFX1 gbuf_d_157(.A(N3077), .Y(ddout__157));
CLKBUFX1 gbuf_q_157(.A(qq_in157), .Y(b_in[6]));
CLKBUFX1 gbuf_d_158(.A(N2949), .Y(ddout__158));
CLKBUFX1 gbuf_q_158(.A(qq_in158), .Y(z_in[6]));
CLKBUFX1 gbuf_d_159(.A(n5694), .Y(ddout__159));
CLKBUFX1 gbuf_q_159(.A(qq_in159), .Y(Out_data[7]));
CLKBUFX1 gbuf_d_160(.A(N3078), .Y(ddout__160));
CLKBUFX1 gbuf_q_160(.A(qq_in160), .Y(b_in[7]));
CLKBUFX1 gbuf_d_161(.A(N2950), .Y(ddout__161));
CLKBUFX1 gbuf_q_161(.A(qq_in161), .Y(z_in[7]));
CLKBUFX1 gbuf_d_162(.A(n5693), .Y(ddout__162));
CLKBUFX1 gbuf_q_162(.A(qq_in162), .Y(Out_data[8]));
CLKBUFX1 gbuf_d_163(.A(N3079), .Y(ddout__163));
CLKBUFX1 gbuf_q_163(.A(qq_in163), .Y(b_in[8]));
CLKBUFX1 gbuf_d_164(.A(N2951), .Y(ddout__164));
CLKBUFX1 gbuf_q_164(.A(qq_in164), .Y(z_in[8]));
CLKBUFX1 gbuf_d_165(.A(n5692), .Y(ddout__165));
CLKBUFX1 gbuf_q_165(.A(qq_in165), .Y(Out_data[9]));
CLKBUFX1 gbuf_d_166(.A(N3080), .Y(ddout__166));
CLKBUFX1 gbuf_q_166(.A(qq_in166), .Y(b_in[9]));
CLKBUFX1 gbuf_d_167(.A(N2952), .Y(ddout__167));
CLKBUFX1 gbuf_q_167(.A(qq_in167), .Y(z_in[9]));
CLKBUFX1 gbuf_d_168(.A(n5691), .Y(ddout__168));
CLKBUFX1 gbuf_q_168(.A(qq_in168), .Y(Out_data[10]));
CLKBUFX1 gbuf_d_169(.A(N3081), .Y(ddout__169));
CLKBUFX1 gbuf_q_169(.A(qq_in169), .Y(b_in[10]));
CLKBUFX1 gbuf_d_170(.A(N2953), .Y(ddout__170));
CLKBUFX1 gbuf_q_170(.A(qq_in170), .Y(z_in[10]));
CLKBUFX1 gbuf_d_171(.A(n5690), .Y(ddout__171));
CLKBUFX1 gbuf_q_171(.A(qq_in171), .Y(Out_data[11]));
CLKBUFX1 gbuf_d_172(.A(N3082), .Y(ddout__172));
CLKBUFX1 gbuf_q_172(.A(qq_in172), .Y(b_in[11]));
CLKBUFX1 gbuf_d_173(.A(N2954), .Y(ddout__173));
CLKBUFX1 gbuf_q_173(.A(qq_in173), .Y(z_in[11]));
CLKBUFX1 gbuf_d_174(.A(n5689), .Y(ddout__174));
CLKBUFX1 gbuf_q_174(.A(qq_in174), .Y(Out_data[12]));
CLKBUFX1 gbuf_d_175(.A(N3083), .Y(ddout__175));
CLKBUFX1 gbuf_q_175(.A(qq_in175), .Y(b_in[12]));
CLKBUFX1 gbuf_d_176(.A(N2955), .Y(ddout__176));
CLKBUFX1 gbuf_q_176(.A(qq_in176), .Y(z_in[12]));
CLKBUFX1 gbuf_d_177(.A(n5688), .Y(ddout__177));
CLKBUFX1 gbuf_q_177(.A(qq_in177), .Y(Out_data[13]));
CLKBUFX1 gbuf_d_178(.A(N3084), .Y(ddout__178));
CLKBUFX1 gbuf_q_178(.A(qq_in178), .Y(b_in[13]));
CLKBUFX1 gbuf_d_179(.A(N2956), .Y(ddout__179));
CLKBUFX1 gbuf_q_179(.A(qq_in179), .Y(z_in[13]));
CLKBUFX1 gbuf_d_180(.A(n5687), .Y(ddout__180));
CLKBUFX1 gbuf_q_180(.A(qq_in180), .Y(Out_data[14]));
CLKBUFX1 gbuf_d_181(.A(N3085), .Y(ddout__181));
CLKBUFX1 gbuf_q_181(.A(qq_in181), .Y(b_in[14]));
CLKBUFX1 gbuf_d_182(.A(N2957), .Y(ddout__182));
CLKBUFX1 gbuf_q_182(.A(qq_in182), .Y(z_in[14]));
CLKBUFX1 gbuf_d_183(.A(n5686), .Y(ddout__183));
CLKBUFX1 gbuf_q_183(.A(qq_in183), .Y(Out_data[15]));
CLKBUFX1 gbuf_d_184(.A(N3086), .Y(ddout__184));
CLKBUFX1 gbuf_q_184(.A(qq_in184), .Y(b_in[15]));
CLKBUFX1 gbuf_d_185(.A(N2958), .Y(ddout__185));
CLKBUFX1 gbuf_q_185(.A(qq_in185), .Y(z_in[15]));
CLKBUFX1 gbuf_d_186(.A(n5685), .Y(ddout__186));
CLKBUFX1 gbuf_q_186(.A(qq_in186), .Y(Out_data[16]));
CLKBUFX1 gbuf_d_187(.A(N3087), .Y(ddout__187));
CLKBUFX1 gbuf_q_187(.A(qq_in187), .Y(b_in[16]));
CLKBUFX1 gbuf_d_188(.A(N2959), .Y(ddout__188));
CLKBUFX1 gbuf_q_188(.A(qq_in188), .Y(z_in[16]));
CLKBUFX1 gbuf_d_189(.A(n5684), .Y(ddout__189));
CLKBUFX1 gbuf_q_189(.A(qq_in189), .Y(Out_data[17]));
CLKBUFX1 gbuf_d_190(.A(N3088), .Y(ddout__190));
CLKBUFX1 gbuf_q_190(.A(qq_in190), .Y(b_in[17]));
CLKBUFX1 gbuf_d_191(.A(N2960), .Y(ddout__191));
CLKBUFX1 gbuf_q_191(.A(qq_in191), .Y(z_in[17]));
CLKBUFX1 gbuf_d_192(.A(n5683), .Y(ddout__192));
CLKBUFX1 gbuf_q_192(.A(qq_in192), .Y(Out_data[18]));
CLKBUFX1 gbuf_d_193(.A(N3089), .Y(ddout__193));
CLKBUFX1 gbuf_q_193(.A(qq_in193), .Y(b_in[18]));
CLKBUFX1 gbuf_d_194(.A(N2961), .Y(ddout__194));
CLKBUFX1 gbuf_q_194(.A(qq_in194), .Y(z_in[18]));
CLKBUFX1 gbuf_d_195(.A(n5682), .Y(ddout__195));
CLKBUFX1 gbuf_q_195(.A(qq_in195), .Y(Out_data[19]));
CLKBUFX1 gbuf_d_196(.A(N3090), .Y(ddout__196));
CLKBUFX1 gbuf_q_196(.A(qq_in196), .Y(b_in[19]));
CLKBUFX1 gbuf_d_197(.A(N2962), .Y(ddout__197));
CLKBUFX1 gbuf_q_197(.A(qq_in197), .Y(z_in[19]));
CLKBUFX1 gbuf_d_198(.A(n5681), .Y(ddout__198));
CLKBUFX1 gbuf_q_198(.A(qq_in198), .Y(Out_data[20]));
CLKBUFX1 gbuf_d_199(.A(N3091), .Y(ddout__199));
CLKBUFX1 gbuf_q_199(.A(qq_in199), .Y(b_in[20]));
CLKBUFX1 gbuf_d_200(.A(N2963), .Y(ddout__200));
CLKBUFX1 gbuf_q_200(.A(qq_in200), .Y(z_in[20]));
CLKBUFX1 gbuf_d_201(.A(n5680), .Y(ddout__201));
CLKBUFX1 gbuf_q_201(.A(qq_in201), .Y(Out_data[21]));
CLKBUFX1 gbuf_d_202(.A(N3092), .Y(ddout__202));
CLKBUFX1 gbuf_q_202(.A(qq_in202), .Y(b_in[21]));
CLKBUFX1 gbuf_d_203(.A(N2964), .Y(ddout__203));
CLKBUFX1 gbuf_q_203(.A(qq_in203), .Y(z_in[21]));
CLKBUFX1 gbuf_d_204(.A(n5679), .Y(ddout__204));
CLKBUFX1 gbuf_q_204(.A(qq_in204), .Y(Out_data[22]));
CLKBUFX1 gbuf_d_205(.A(N3093), .Y(ddout__205));
CLKBUFX1 gbuf_q_205(.A(qq_in205), .Y(b_in[22]));
CLKBUFX1 gbuf_d_206(.A(N2965), .Y(ddout__206));
CLKBUFX1 gbuf_q_206(.A(qq_in206), .Y(z_in[22]));
CLKBUFX1 gbuf_d_207(.A(n5678), .Y(ddout__207));
CLKBUFX1 gbuf_q_207(.A(qq_in207), .Y(Out_data[23]));
CLKBUFX1 gbuf_d_208(.A(N3094), .Y(ddout__208));
CLKBUFX1 gbuf_q_208(.A(qq_in208), .Y(b_in[23]));
CLKBUFX1 gbuf_d_209(.A(N2966), .Y(ddout__209));
CLKBUFX1 gbuf_q_209(.A(qq_in209), .Y(z_in[23]));
CLKBUFX1 gbuf_d_210(.A(n5677), .Y(ddout__210));
CLKBUFX1 gbuf_q_210(.A(qq_in210), .Y(Out_data[24]));
CLKBUFX1 gbuf_d_211(.A(N3095), .Y(ddout__211));
CLKBUFX1 gbuf_q_211(.A(qq_in211), .Y(b_in[24]));
CLKBUFX1 gbuf_d_212(.A(N2967), .Y(ddout__212));
CLKBUFX1 gbuf_q_212(.A(qq_in212), .Y(z_in[24]));
CLKBUFX1 gbuf_d_213(.A(n5676), .Y(ddout__213));
CLKBUFX1 gbuf_q_213(.A(qq_in213), .Y(Out_data[25]));
CLKBUFX1 gbuf_d_214(.A(N3096), .Y(ddout__214));
CLKBUFX1 gbuf_q_214(.A(qq_in214), .Y(b_in[25]));
CLKBUFX1 gbuf_d_215(.A(N2968), .Y(ddout__215));
CLKBUFX1 gbuf_q_215(.A(qq_in215), .Y(z_in[25]));
CLKBUFX1 gbuf_d_216(.A(n5675), .Y(ddout__216));
CLKBUFX1 gbuf_q_216(.A(qq_in216), .Y(Out_data[26]));
CLKBUFX1 gbuf_d_217(.A(N3097), .Y(ddout__217));
CLKBUFX1 gbuf_q_217(.A(qq_in217), .Y(b_in[26]));
CLKBUFX1 gbuf_d_218(.A(N2969), .Y(ddout__218));
CLKBUFX1 gbuf_q_218(.A(qq_in218), .Y(z_in[26]));
CLKBUFX1 gbuf_d_219(.A(n5674), .Y(ddout__219));
CLKBUFX1 gbuf_q_219(.A(qq_in219), .Y(Out_data[27]));
CLKBUFX1 gbuf_d_220(.A(N3098), .Y(ddout__220));
CLKBUFX1 gbuf_q_220(.A(qq_in220), .Y(b_in[27]));
CLKBUFX1 gbuf_d_221(.A(N2970), .Y(ddout__221));
CLKBUFX1 gbuf_q_221(.A(qq_in221), .Y(z_in[27]));
CLKBUFX1 gbuf_d_222(.A(n5673), .Y(ddout__222));
CLKBUFX1 gbuf_q_222(.A(qq_in222), .Y(Out_data[28]));
CLKBUFX1 gbuf_d_223(.A(N3099), .Y(ddout__223));
CLKBUFX1 gbuf_q_223(.A(qq_in223), .Y(b_in[28]));
CLKBUFX1 gbuf_d_224(.A(N2971), .Y(ddout__224));
CLKBUFX1 gbuf_q_224(.A(qq_in224), .Y(z_in[28]));
CLKBUFX1 gbuf_d_225(.A(n5672), .Y(ddout__225));
CLKBUFX1 gbuf_q_225(.A(qq_in225), .Y(Out_data[29]));
CLKBUFX1 gbuf_d_226(.A(N3100), .Y(ddout__226));
CLKBUFX1 gbuf_q_226(.A(qq_in226), .Y(b_in[29]));
CLKBUFX1 gbuf_d_227(.A(N2972), .Y(ddout__227));
CLKBUFX1 gbuf_q_227(.A(qq_in227), .Y(z_in[29]));
CLKBUFX1 gbuf_d_228(.A(n5671), .Y(ddout__228));
CLKBUFX1 gbuf_q_228(.A(qq_in228), .Y(Out_data[30]));
CLKBUFX1 gbuf_d_229(.A(N3101), .Y(ddout__229));
CLKBUFX1 gbuf_q_229(.A(qq_in229), .Y(b_in[30]));
CLKBUFX1 gbuf_d_230(.A(N2973), .Y(ddout__230));
CLKBUFX1 gbuf_q_230(.A(qq_in230), .Y(z_in[30]));
CLKBUFX1 gbuf_d_231(.A(n5670), .Y(ddout__231));
CLKBUFX1 gbuf_q_231(.A(qq_in231), .Y(Out_data[31]));
CLKBUFX1 gbuf_d_232(.A(N3102), .Y(ddout__232));
CLKBUFX1 gbuf_q_232(.A(qq_in232), .Y(b_in[31]));
CLKBUFX1 gbuf_d_233(.A(N2974), .Y(ddout__233));
CLKBUFX1 gbuf_q_233(.A(qq_in233), .Y(z_in[31]));
CLKBUFX1 gbuf_d_234(.A(n5669), .Y(ddout__234));
CLKBUFX1 gbuf_q_234(.A(qq_in234), .Y(Out_data[32]));
CLKBUFX1 gbuf_d_235(.A(N3103), .Y(ddout__235));
CLKBUFX1 gbuf_q_235(.A(qq_in235), .Y(b_in[32]));
CLKBUFX1 gbuf_d_236(.A(N2975), .Y(ddout__236));
CLKBUFX1 gbuf_q_236(.A(qq_in236), .Y(z_in[32]));
CLKBUFX1 gbuf_d_237(.A(n5668), .Y(ddout__237));
CLKBUFX1 gbuf_q_237(.A(qq_in237), .Y(Out_data[33]));
CLKBUFX1 gbuf_d_238(.A(N3104), .Y(ddout__238));
CLKBUFX1 gbuf_q_238(.A(qq_in238), .Y(b_in[33]));
CLKBUFX1 gbuf_d_239(.A(N2976), .Y(ddout__239));
CLKBUFX1 gbuf_q_239(.A(qq_in239), .Y(z_in[33]));
CLKBUFX1 gbuf_d_240(.A(n5667), .Y(ddout__240));
CLKBUFX1 gbuf_q_240(.A(qq_in240), .Y(Out_data[34]));
CLKBUFX1 gbuf_d_241(.A(N3105), .Y(ddout__241));
CLKBUFX1 gbuf_q_241(.A(qq_in241), .Y(b_in[34]));
CLKBUFX1 gbuf_d_242(.A(N2977), .Y(ddout__242));
CLKBUFX1 gbuf_q_242(.A(qq_in242), .Y(z_in[34]));
CLKBUFX1 gbuf_d_243(.A(n5666), .Y(ddout__243));
CLKBUFX1 gbuf_q_243(.A(qq_in243), .Y(Out_data[35]));
CLKBUFX1 gbuf_d_244(.A(N3106), .Y(ddout__244));
CLKBUFX1 gbuf_q_244(.A(qq_in244), .Y(b_in[35]));
CLKBUFX1 gbuf_d_245(.A(N2978), .Y(ddout__245));
CLKBUFX1 gbuf_q_245(.A(qq_in245), .Y(z_in[35]));
CLKBUFX1 gbuf_d_246(.A(n5665), .Y(ddout__246));
CLKBUFX1 gbuf_q_246(.A(qq_in246), .Y(Out_data[36]));
CLKBUFX1 gbuf_d_247(.A(N3107), .Y(ddout__247));
CLKBUFX1 gbuf_q_247(.A(qq_in247), .Y(b_in[36]));
CLKBUFX1 gbuf_d_248(.A(N2979), .Y(ddout__248));
CLKBUFX1 gbuf_q_248(.A(qq_in248), .Y(z_in[36]));
CLKBUFX1 gbuf_d_249(.A(n5664), .Y(ddout__249));
CLKBUFX1 gbuf_q_249(.A(qq_in249), .Y(Out_data[37]));
CLKBUFX1 gbuf_d_250(.A(N3108), .Y(ddout__250));
CLKBUFX1 gbuf_q_250(.A(qq_in250), .Y(b_in[37]));
CLKBUFX1 gbuf_d_251(.A(N2980), .Y(ddout__251));
CLKBUFX1 gbuf_q_251(.A(qq_in251), .Y(z_in[37]));
CLKBUFX1 gbuf_d_252(.A(n5663), .Y(ddout__252));
CLKBUFX1 gbuf_q_252(.A(qq_in252), .Y(Out_data[38]));
CLKBUFX1 gbuf_d_253(.A(N3109), .Y(ddout__253));
CLKBUFX1 gbuf_q_253(.A(qq_in253), .Y(b_in[38]));
CLKBUFX1 gbuf_d_254(.A(N2981), .Y(ddout__254));
CLKBUFX1 gbuf_q_254(.A(qq_in254), .Y(z_in[38]));
CLKBUFX1 gbuf_d_255(.A(n5662), .Y(ddout__255));
CLKBUFX1 gbuf_q_255(.A(qq_in255), .Y(Out_data[39]));
CLKBUFX1 gbuf_d_256(.A(N3110), .Y(ddout__256));
CLKBUFX1 gbuf_q_256(.A(qq_in256), .Y(b_in[39]));
CLKBUFX1 gbuf_d_257(.A(N2982), .Y(ddout__257));
CLKBUFX1 gbuf_q_257(.A(qq_in257), .Y(z_in[39]));
CLKBUFX1 gbuf_d_258(.A(n5661), .Y(ddout__258));
CLKBUFX1 gbuf_q_258(.A(qq_in258), .Y(Out_data[40]));
CLKBUFX1 gbuf_d_259(.A(N3111), .Y(ddout__259));
CLKBUFX1 gbuf_q_259(.A(qq_in259), .Y(b_in[40]));
CLKBUFX1 gbuf_d_260(.A(N2983), .Y(ddout__260));
CLKBUFX1 gbuf_q_260(.A(qq_in260), .Y(z_in[40]));
CLKBUFX1 gbuf_d_261(.A(n5660), .Y(ddout__261));
CLKBUFX1 gbuf_q_261(.A(qq_in261), .Y(Out_data[41]));
CLKBUFX1 gbuf_d_262(.A(N3112), .Y(ddout__262));
CLKBUFX1 gbuf_q_262(.A(qq_in262), .Y(b_in[41]));
CLKBUFX1 gbuf_d_263(.A(N2984), .Y(ddout__263));
CLKBUFX1 gbuf_q_263(.A(qq_in263), .Y(z_in[41]));
CLKBUFX1 gbuf_d_264(.A(n5659), .Y(ddout__264));
CLKBUFX1 gbuf_q_264(.A(qq_in264), .Y(Out_data[42]));
CLKBUFX1 gbuf_d_265(.A(N3113), .Y(ddout__265));
CLKBUFX1 gbuf_q_265(.A(qq_in265), .Y(b_in[42]));
CLKBUFX1 gbuf_d_266(.A(N2985), .Y(ddout__266));
CLKBUFX1 gbuf_q_266(.A(qq_in266), .Y(z_in[42]));
CLKBUFX1 gbuf_d_267(.A(n5658), .Y(ddout__267));
CLKBUFX1 gbuf_q_267(.A(qq_in267), .Y(Out_data[43]));
CLKBUFX1 gbuf_d_268(.A(N3114), .Y(ddout__268));
CLKBUFX1 gbuf_q_268(.A(qq_in268), .Y(b_in[43]));
CLKBUFX1 gbuf_d_269(.A(N2986), .Y(ddout__269));
CLKBUFX1 gbuf_q_269(.A(qq_in269), .Y(z_in[43]));
CLKBUFX1 gbuf_d_270(.A(n5657), .Y(ddout__270));
CLKBUFX1 gbuf_q_270(.A(qq_in270), .Y(Out_data[44]));
CLKBUFX1 gbuf_d_271(.A(N3115), .Y(ddout__271));
CLKBUFX1 gbuf_q_271(.A(qq_in271), .Y(b_in[44]));
CLKBUFX1 gbuf_d_272(.A(N2987), .Y(ddout__272));
CLKBUFX1 gbuf_q_272(.A(qq_in272), .Y(z_in[44]));
CLKBUFX1 gbuf_d_273(.A(n5656), .Y(ddout__273));
CLKBUFX1 gbuf_q_273(.A(qq_in273), .Y(Out_data[45]));
CLKBUFX1 gbuf_d_274(.A(N3116), .Y(ddout__274));
CLKBUFX1 gbuf_q_274(.A(qq_in274), .Y(b_in[45]));
CLKBUFX1 gbuf_d_275(.A(N2988), .Y(ddout__275));
CLKBUFX1 gbuf_q_275(.A(qq_in275), .Y(z_in[45]));
CLKBUFX1 gbuf_d_276(.A(n5655), .Y(ddout__276));
CLKBUFX1 gbuf_q_276(.A(qq_in276), .Y(Out_data[46]));
CLKBUFX1 gbuf_d_277(.A(N3117), .Y(ddout__277));
CLKBUFX1 gbuf_q_277(.A(qq_in277), .Y(b_in[46]));
CLKBUFX1 gbuf_d_278(.A(N2989), .Y(ddout__278));
CLKBUFX1 gbuf_q_278(.A(qq_in278), .Y(z_in[46]));
CLKBUFX1 gbuf_d_279(.A(n5654), .Y(ddout__279));
CLKBUFX1 gbuf_q_279(.A(qq_in279), .Y(Out_data[47]));
CLKBUFX1 gbuf_d_280(.A(N3118), .Y(ddout__280));
CLKBUFX1 gbuf_q_280(.A(qq_in280), .Y(b_in[47]));
CLKBUFX1 gbuf_d_281(.A(N2990), .Y(ddout__281));
CLKBUFX1 gbuf_q_281(.A(qq_in281), .Y(z_in[47]));
CLKBUFX1 gbuf_d_282(.A(n5653), .Y(ddout__282));
CLKBUFX1 gbuf_q_282(.A(qq_in282), .Y(Out_data[48]));
CLKBUFX1 gbuf_d_283(.A(N3119), .Y(ddout__283));
CLKBUFX1 gbuf_q_283(.A(qq_in283), .Y(b_in[48]));
CLKBUFX1 gbuf_d_284(.A(N2991), .Y(ddout__284));
CLKBUFX1 gbuf_q_284(.A(qq_in284), .Y(z_in[48]));
CLKBUFX1 gbuf_d_285(.A(n5652), .Y(ddout__285));
CLKBUFX1 gbuf_q_285(.A(qq_in285), .Y(Out_data[49]));
CLKBUFX1 gbuf_d_286(.A(N3120), .Y(ddout__286));
CLKBUFX1 gbuf_q_286(.A(qq_in286), .Y(b_in[49]));
CLKBUFX1 gbuf_d_287(.A(N2992), .Y(ddout__287));
CLKBUFX1 gbuf_q_287(.A(qq_in287), .Y(z_in[49]));
CLKBUFX1 gbuf_d_288(.A(n5651), .Y(ddout__288));
CLKBUFX1 gbuf_q_288(.A(qq_in288), .Y(Out_data[50]));
CLKBUFX1 gbuf_d_289(.A(N3121), .Y(ddout__289));
CLKBUFX1 gbuf_q_289(.A(qq_in289), .Y(b_in[50]));
CLKBUFX1 gbuf_d_290(.A(N2993), .Y(ddout__290));
CLKBUFX1 gbuf_q_290(.A(qq_in290), .Y(z_in[50]));
CLKBUFX1 gbuf_d_291(.A(n5650), .Y(ddout__291));
CLKBUFX1 gbuf_q_291(.A(qq_in291), .Y(Out_data[51]));
CLKBUFX1 gbuf_d_292(.A(N3122), .Y(ddout__292));
CLKBUFX1 gbuf_q_292(.A(qq_in292), .Y(b_in[51]));
CLKBUFX1 gbuf_d_293(.A(N2994), .Y(ddout__293));
CLKBUFX1 gbuf_q_293(.A(qq_in293), .Y(z_in[51]));
CLKBUFX1 gbuf_d_294(.A(n5649), .Y(ddout__294));
CLKBUFX1 gbuf_q_294(.A(qq_in294), .Y(Out_data[52]));
CLKBUFX1 gbuf_d_295(.A(N3123), .Y(ddout__295));
CLKBUFX1 gbuf_q_295(.A(qq_in295), .Y(b_in[52]));
CLKBUFX1 gbuf_d_296(.A(N2995), .Y(ddout__296));
CLKBUFX1 gbuf_q_296(.A(qq_in296), .Y(z_in[52]));
CLKBUFX1 gbuf_d_297(.A(n5648), .Y(ddout__297));
CLKBUFX1 gbuf_q_297(.A(qq_in297), .Y(Out_data[53]));
CLKBUFX1 gbuf_d_298(.A(N3124), .Y(ddout__298));
CLKBUFX1 gbuf_q_298(.A(qq_in298), .Y(b_in[53]));
CLKBUFX1 gbuf_d_299(.A(N2996), .Y(ddout__299));
CLKBUFX1 gbuf_q_299(.A(qq_in299), .Y(z_in[53]));
CLKBUFX1 gbuf_d_300(.A(n5647), .Y(ddout__300));
CLKBUFX1 gbuf_q_300(.A(qq_in300), .Y(Out_data[54]));
CLKBUFX1 gbuf_d_301(.A(N3125), .Y(ddout__301));
CLKBUFX1 gbuf_q_301(.A(qq_in301), .Y(b_in[54]));
CLKBUFX1 gbuf_d_302(.A(N2997), .Y(ddout__302));
CLKBUFX1 gbuf_q_302(.A(qq_in302), .Y(z_in[54]));
CLKBUFX1 gbuf_d_303(.A(n5646), .Y(ddout__303));
CLKBUFX1 gbuf_q_303(.A(qq_in303), .Y(Out_data[55]));
CLKBUFX1 gbuf_d_304(.A(N3126), .Y(ddout__304));
CLKBUFX1 gbuf_q_304(.A(qq_in304), .Y(b_in[55]));
CLKBUFX1 gbuf_d_305(.A(N2998), .Y(ddout__305));
CLKBUFX1 gbuf_q_305(.A(qq_in305), .Y(z_in[55]));
CLKBUFX1 gbuf_d_306(.A(n5645), .Y(ddout__306));
CLKBUFX1 gbuf_q_306(.A(qq_in306), .Y(Out_data[56]));
CLKBUFX1 gbuf_d_307(.A(N3127), .Y(ddout__307));
CLKBUFX1 gbuf_q_307(.A(qq_in307), .Y(b_in[56]));
CLKBUFX1 gbuf_d_308(.A(N2999), .Y(ddout__308));
CLKBUFX1 gbuf_q_308(.A(qq_in308), .Y(z_in[56]));
CLKBUFX1 gbuf_d_309(.A(n5644), .Y(ddout__309));
CLKBUFX1 gbuf_q_309(.A(qq_in309), .Y(Out_data[57]));
CLKBUFX1 gbuf_d_310(.A(N3128), .Y(ddout__310));
CLKBUFX1 gbuf_q_310(.A(qq_in310), .Y(b_in[57]));
CLKBUFX1 gbuf_d_311(.A(N3000), .Y(ddout__311));
CLKBUFX1 gbuf_q_311(.A(qq_in311), .Y(z_in[57]));
CLKBUFX1 gbuf_d_312(.A(n5643), .Y(ddout__312));
CLKBUFX1 gbuf_q_312(.A(qq_in312), .Y(Out_data[58]));
CLKBUFX1 gbuf_d_313(.A(N3129), .Y(ddout__313));
CLKBUFX1 gbuf_q_313(.A(qq_in313), .Y(b_in[58]));
CLKBUFX1 gbuf_d_314(.A(N3001), .Y(ddout__314));
CLKBUFX1 gbuf_q_314(.A(qq_in314), .Y(z_in[58]));
CLKBUFX1 gbuf_d_315(.A(n5642), .Y(ddout__315));
CLKBUFX1 gbuf_q_315(.A(qq_in315), .Y(Out_data[59]));
CLKBUFX1 gbuf_d_316(.A(N3130), .Y(ddout__316));
CLKBUFX1 gbuf_q_316(.A(qq_in316), .Y(b_in[59]));
CLKBUFX1 gbuf_d_317(.A(N3002), .Y(ddout__317));
CLKBUFX1 gbuf_q_317(.A(qq_in317), .Y(z_in[59]));
CLKBUFX1 gbuf_d_318(.A(n5641), .Y(ddout__318));
CLKBUFX1 gbuf_q_318(.A(qq_in318), .Y(Out_data[60]));
CLKBUFX1 gbuf_d_319(.A(N3131), .Y(ddout__319));
CLKBUFX1 gbuf_q_319(.A(qq_in319), .Y(b_in[60]));
CLKBUFX1 gbuf_d_320(.A(N3003), .Y(ddout__320));
CLKBUFX1 gbuf_q_320(.A(qq_in320), .Y(z_in[60]));
CLKBUFX1 gbuf_d_321(.A(n5640), .Y(ddout__321));
CLKBUFX1 gbuf_q_321(.A(qq_in321), .Y(Out_data[61]));
CLKBUFX1 gbuf_d_322(.A(N3132), .Y(ddout__322));
CLKBUFX1 gbuf_q_322(.A(qq_in322), .Y(b_in[61]));
CLKBUFX1 gbuf_d_323(.A(N3004), .Y(ddout__323));
CLKBUFX1 gbuf_q_323(.A(qq_in323), .Y(z_in[61]));
CLKBUFX1 gbuf_d_324(.A(n5639), .Y(ddout__324));
CLKBUFX1 gbuf_q_324(.A(qq_in324), .Y(Out_data[62]));
CLKBUFX1 gbuf_d_325(.A(N3133), .Y(ddout__325));
CLKBUFX1 gbuf_q_325(.A(qq_in325), .Y(b_in[62]));
CLKBUFX1 gbuf_d_326(.A(N3005), .Y(ddout__326));
CLKBUFX1 gbuf_q_326(.A(qq_in326), .Y(z_in[62]));
CLKBUFX1 gbuf_d_327(.A(n5638), .Y(ddout__327));
CLKBUFX1 gbuf_q_327(.A(qq_in327), .Y(Out_data[63]));
CLKBUFX1 gbuf_d_328(.A(N3134), .Y(ddout__328));
CLKBUFX1 gbuf_q_328(.A(qq_in328), .Y(b_in[63]));
CLKBUFX1 gbuf_d_329(.A(N3006), .Y(ddout__329));
CLKBUFX1 gbuf_q_329(.A(qq_in329), .Y(z_in[63]));
CLKBUFX1 gbuf_d_330(.A(n5637), .Y(ddout__330));
CLKBUFX1 gbuf_q_330(.A(qq_in330), .Y(Out_data[64]));
CLKBUFX1 gbuf_d_331(.A(N3135), .Y(ddout__331));
CLKBUFX1 gbuf_q_331(.A(qq_in331), .Y(b_in[64]));
CLKBUFX1 gbuf_d_332(.A(N3007), .Y(ddout__332));
CLKBUFX1 gbuf_q_332(.A(qq_in332), .Y(z_in[64]));
CLKBUFX1 gbuf_d_333(.A(n5636), .Y(ddout__333));
CLKBUFX1 gbuf_q_333(.A(qq_in333), .Y(Out_data[65]));
CLKBUFX1 gbuf_d_334(.A(N3136), .Y(ddout__334));
CLKBUFX1 gbuf_q_334(.A(qq_in334), .Y(b_in[65]));
CLKBUFX1 gbuf_d_335(.A(N3008), .Y(ddout__335));
CLKBUFX1 gbuf_q_335(.A(qq_in335), .Y(z_in[65]));
CLKBUFX1 gbuf_d_336(.A(n5635), .Y(ddout__336));
CLKBUFX1 gbuf_q_336(.A(qq_in336), .Y(Out_data[66]));
CLKBUFX1 gbuf_d_337(.A(N3137), .Y(ddout__337));
CLKBUFX1 gbuf_q_337(.A(qq_in337), .Y(b_in[66]));
CLKBUFX1 gbuf_d_338(.A(N3009), .Y(ddout__338));
CLKBUFX1 gbuf_q_338(.A(qq_in338), .Y(z_in[66]));
CLKBUFX1 gbuf_d_339(.A(n5634), .Y(ddout__339));
CLKBUFX1 gbuf_q_339(.A(qq_in339), .Y(Out_data[67]));
CLKBUFX1 gbuf_d_340(.A(N3138), .Y(ddout__340));
CLKBUFX1 gbuf_q_340(.A(qq_in340), .Y(b_in[67]));
CLKBUFX1 gbuf_d_341(.A(N3010), .Y(ddout__341));
CLKBUFX1 gbuf_q_341(.A(qq_in341), .Y(z_in[67]));
CLKBUFX1 gbuf_d_342(.A(n5633), .Y(ddout__342));
CLKBUFX1 gbuf_q_342(.A(qq_in342), .Y(Out_data[68]));
CLKBUFX1 gbuf_d_343(.A(N3139), .Y(ddout__343));
CLKBUFX1 gbuf_q_343(.A(qq_in343), .Y(b_in[68]));
CLKBUFX1 gbuf_d_344(.A(N3011), .Y(ddout__344));
CLKBUFX1 gbuf_q_344(.A(qq_in344), .Y(z_in[68]));
CLKBUFX1 gbuf_d_345(.A(n5632), .Y(ddout__345));
CLKBUFX1 gbuf_q_345(.A(qq_in345), .Y(Out_data[69]));
CLKBUFX1 gbuf_d_346(.A(N3140), .Y(ddout__346));
CLKBUFX1 gbuf_q_346(.A(qq_in346), .Y(b_in[69]));
CLKBUFX1 gbuf_d_347(.A(N3012), .Y(ddout__347));
CLKBUFX1 gbuf_q_347(.A(qq_in347), .Y(z_in[69]));
CLKBUFX1 gbuf_d_348(.A(n5631), .Y(ddout__348));
CLKBUFX1 gbuf_q_348(.A(qq_in348), .Y(Out_data[70]));
CLKBUFX1 gbuf_d_349(.A(N3141), .Y(ddout__349));
CLKBUFX1 gbuf_q_349(.A(qq_in349), .Y(b_in[70]));
CLKBUFX1 gbuf_d_350(.A(N3013), .Y(ddout__350));
CLKBUFX1 gbuf_q_350(.A(qq_in350), .Y(z_in[70]));
CLKBUFX1 gbuf_d_351(.A(n5630), .Y(ddout__351));
CLKBUFX1 gbuf_q_351(.A(qq_in351), .Y(Out_data[71]));
CLKBUFX1 gbuf_d_352(.A(N3142), .Y(ddout__352));
CLKBUFX1 gbuf_q_352(.A(qq_in352), .Y(b_in[71]));
CLKBUFX1 gbuf_d_353(.A(N3014), .Y(ddout__353));
CLKBUFX1 gbuf_q_353(.A(qq_in353), .Y(z_in[71]));
CLKBUFX1 gbuf_d_354(.A(n5629), .Y(ddout__354));
CLKBUFX1 gbuf_q_354(.A(qq_in354), .Y(Out_data[72]));
CLKBUFX1 gbuf_d_355(.A(N3143), .Y(ddout__355));
CLKBUFX1 gbuf_q_355(.A(qq_in355), .Y(b_in[72]));
CLKBUFX1 gbuf_d_356(.A(N3015), .Y(ddout__356));
CLKBUFX1 gbuf_q_356(.A(qq_in356), .Y(z_in[72]));
CLKBUFX1 gbuf_d_357(.A(n5628), .Y(ddout__357));
CLKBUFX1 gbuf_q_357(.A(qq_in357), .Y(Out_data[73]));
CLKBUFX1 gbuf_d_358(.A(N3144), .Y(ddout__358));
CLKBUFX1 gbuf_q_358(.A(qq_in358), .Y(b_in[73]));
CLKBUFX1 gbuf_d_359(.A(N3016), .Y(ddout__359));
CLKBUFX1 gbuf_q_359(.A(qq_in359), .Y(z_in[73]));
CLKBUFX1 gbuf_d_360(.A(n5627), .Y(ddout__360));
CLKBUFX1 gbuf_q_360(.A(qq_in360), .Y(Out_data[74]));
CLKBUFX1 gbuf_d_361(.A(N3145), .Y(ddout__361));
CLKBUFX1 gbuf_q_361(.A(qq_in361), .Y(b_in[74]));
CLKBUFX1 gbuf_d_362(.A(N3017), .Y(ddout__362));
CLKBUFX1 gbuf_q_362(.A(qq_in362), .Y(z_in[74]));
CLKBUFX1 gbuf_d_363(.A(n5626), .Y(ddout__363));
CLKBUFX1 gbuf_q_363(.A(qq_in363), .Y(Out_data[75]));
CLKBUFX1 gbuf_d_364(.A(N3146), .Y(ddout__364));
CLKBUFX1 gbuf_q_364(.A(qq_in364), .Y(b_in[75]));
CLKBUFX1 gbuf_d_365(.A(N3018), .Y(ddout__365));
CLKBUFX1 gbuf_q_365(.A(qq_in365), .Y(z_in[75]));
CLKBUFX1 gbuf_d_366(.A(n5625), .Y(ddout__366));
CLKBUFX1 gbuf_q_366(.A(qq_in366), .Y(Out_data[76]));
CLKBUFX1 gbuf_d_367(.A(N3147), .Y(ddout__367));
CLKBUFX1 gbuf_q_367(.A(qq_in367), .Y(b_in[76]));
CLKBUFX1 gbuf_d_368(.A(N3019), .Y(ddout__368));
CLKBUFX1 gbuf_q_368(.A(qq_in368), .Y(z_in[76]));
CLKBUFX1 gbuf_d_369(.A(n5624), .Y(ddout__369));
CLKBUFX1 gbuf_q_369(.A(qq_in369), .Y(Out_data[77]));
CLKBUFX1 gbuf_d_370(.A(N3148), .Y(ddout__370));
CLKBUFX1 gbuf_q_370(.A(qq_in370), .Y(b_in[77]));
CLKBUFX1 gbuf_d_371(.A(N3020), .Y(ddout__371));
CLKBUFX1 gbuf_q_371(.A(qq_in371), .Y(z_in[77]));
CLKBUFX1 gbuf_d_372(.A(n5623), .Y(ddout__372));
CLKBUFX1 gbuf_q_372(.A(qq_in372), .Y(Out_data[78]));
CLKBUFX1 gbuf_d_373(.A(N3149), .Y(ddout__373));
CLKBUFX1 gbuf_q_373(.A(qq_in373), .Y(b_in[78]));
CLKBUFX1 gbuf_d_374(.A(N3021), .Y(ddout__374));
CLKBUFX1 gbuf_q_374(.A(qq_in374), .Y(z_in[78]));
CLKBUFX1 gbuf_d_375(.A(n5622), .Y(ddout__375));
CLKBUFX1 gbuf_q_375(.A(qq_in375), .Y(Out_data[79]));
CLKBUFX1 gbuf_d_376(.A(N3150), .Y(ddout__376));
CLKBUFX1 gbuf_q_376(.A(qq_in376), .Y(b_in[79]));
CLKBUFX1 gbuf_d_377(.A(N3022), .Y(ddout__377));
CLKBUFX1 gbuf_q_377(.A(qq_in377), .Y(z_in[79]));
CLKBUFX1 gbuf_d_378(.A(n5621), .Y(ddout__378));
CLKBUFX1 gbuf_q_378(.A(qq_in378), .Y(Out_data[80]));
CLKBUFX1 gbuf_d_379(.A(N3151), .Y(ddout__379));
CLKBUFX1 gbuf_q_379(.A(qq_in379), .Y(b_in[80]));
CLKBUFX1 gbuf_d_380(.A(N3023), .Y(ddout__380));
CLKBUFX1 gbuf_q_380(.A(qq_in380), .Y(z_in[80]));
CLKBUFX1 gbuf_d_381(.A(n5620), .Y(ddout__381));
CLKBUFX1 gbuf_q_381(.A(qq_in381), .Y(Out_data[81]));
CLKBUFX1 gbuf_d_382(.A(N3152), .Y(ddout__382));
CLKBUFX1 gbuf_q_382(.A(qq_in382), .Y(b_in[81]));
CLKBUFX1 gbuf_d_383(.A(N3024), .Y(ddout__383));
CLKBUFX1 gbuf_q_383(.A(qq_in383), .Y(z_in[81]));
CLKBUFX1 gbuf_d_384(.A(n5619), .Y(ddout__384));
CLKBUFX1 gbuf_q_384(.A(qq_in384), .Y(Out_data[82]));
CLKBUFX1 gbuf_d_385(.A(N3153), .Y(ddout__385));
CLKBUFX1 gbuf_q_385(.A(qq_in385), .Y(b_in[82]));
CLKBUFX1 gbuf_d_386(.A(N3025), .Y(ddout__386));
CLKBUFX1 gbuf_q_386(.A(qq_in386), .Y(z_in[82]));
CLKBUFX1 gbuf_d_387(.A(n5618), .Y(ddout__387));
CLKBUFX1 gbuf_q_387(.A(qq_in387), .Y(Out_data[83]));
CLKBUFX1 gbuf_d_388(.A(N3154), .Y(ddout__388));
CLKBUFX1 gbuf_q_388(.A(qq_in388), .Y(b_in[83]));
CLKBUFX1 gbuf_d_389(.A(N3026), .Y(ddout__389));
CLKBUFX1 gbuf_q_389(.A(qq_in389), .Y(z_in[83]));
CLKBUFX1 gbuf_d_390(.A(n5617), .Y(ddout__390));
CLKBUFX1 gbuf_q_390(.A(qq_in390), .Y(Out_data[84]));
CLKBUFX1 gbuf_d_391(.A(N3155), .Y(ddout__391));
CLKBUFX1 gbuf_q_391(.A(qq_in391), .Y(b_in[84]));
CLKBUFX1 gbuf_d_392(.A(N3027), .Y(ddout__392));
CLKBUFX1 gbuf_q_392(.A(qq_in392), .Y(z_in[84]));
CLKBUFX1 gbuf_d_393(.A(n5616), .Y(ddout__393));
CLKBUFX1 gbuf_q_393(.A(qq_in393), .Y(Out_data[85]));
CLKBUFX1 gbuf_d_394(.A(N3156), .Y(ddout__394));
CLKBUFX1 gbuf_q_394(.A(qq_in394), .Y(b_in[85]));
CLKBUFX1 gbuf_d_395(.A(N3028), .Y(ddout__395));
CLKBUFX1 gbuf_q_395(.A(qq_in395), .Y(z_in[85]));
CLKBUFX1 gbuf_d_396(.A(n5615), .Y(ddout__396));
CLKBUFX1 gbuf_q_396(.A(qq_in396), .Y(Out_data[86]));
CLKBUFX1 gbuf_d_397(.A(N3157), .Y(ddout__397));
CLKBUFX1 gbuf_q_397(.A(qq_in397), .Y(b_in[86]));
CLKBUFX1 gbuf_d_398(.A(N3029), .Y(ddout__398));
CLKBUFX1 gbuf_q_398(.A(qq_in398), .Y(z_in[86]));
CLKBUFX1 gbuf_d_399(.A(n5614), .Y(ddout__399));
CLKBUFX1 gbuf_q_399(.A(qq_in399), .Y(Out_data[87]));
CLKBUFX1 gbuf_d_400(.A(N3158), .Y(ddout__400));
CLKBUFX1 gbuf_q_400(.A(qq_in400), .Y(b_in[87]));
CLKBUFX1 gbuf_d_401(.A(N3030), .Y(ddout__401));
CLKBUFX1 gbuf_q_401(.A(qq_in401), .Y(z_in[87]));
CLKBUFX1 gbuf_d_402(.A(n5613), .Y(ddout__402));
CLKBUFX1 gbuf_q_402(.A(qq_in402), .Y(Out_data[88]));
CLKBUFX1 gbuf_d_403(.A(N3159), .Y(ddout__403));
CLKBUFX1 gbuf_q_403(.A(qq_in403), .Y(b_in[88]));
CLKBUFX1 gbuf_d_404(.A(N3031), .Y(ddout__404));
CLKBUFX1 gbuf_q_404(.A(qq_in404), .Y(z_in[88]));
CLKBUFX1 gbuf_d_405(.A(n5612), .Y(ddout__405));
CLKBUFX1 gbuf_q_405(.A(qq_in405), .Y(Out_data[89]));
CLKBUFX1 gbuf_d_406(.A(N3160), .Y(ddout__406));
CLKBUFX1 gbuf_q_406(.A(qq_in406), .Y(b_in[89]));
CLKBUFX1 gbuf_d_407(.A(N3032), .Y(ddout__407));
CLKBUFX1 gbuf_q_407(.A(qq_in407), .Y(z_in[89]));
CLKBUFX1 gbuf_d_408(.A(n5611), .Y(ddout__408));
CLKBUFX1 gbuf_q_408(.A(qq_in408), .Y(Out_data[90]));
CLKBUFX1 gbuf_d_409(.A(N3161), .Y(ddout__409));
CLKBUFX1 gbuf_q_409(.A(qq_in409), .Y(b_in[90]));
CLKBUFX1 gbuf_d_410(.A(N3033), .Y(ddout__410));
CLKBUFX1 gbuf_q_410(.A(qq_in410), .Y(z_in[90]));
CLKBUFX1 gbuf_d_411(.A(n5610), .Y(ddout__411));
CLKBUFX1 gbuf_q_411(.A(qq_in411), .Y(Out_data[91]));
CLKBUFX1 gbuf_d_412(.A(N3162), .Y(ddout__412));
CLKBUFX1 gbuf_q_412(.A(qq_in412), .Y(b_in[91]));
CLKBUFX1 gbuf_d_413(.A(N3034), .Y(ddout__413));
CLKBUFX1 gbuf_q_413(.A(qq_in413), .Y(z_in[91]));
CLKBUFX1 gbuf_d_414(.A(n5609), .Y(ddout__414));
CLKBUFX1 gbuf_q_414(.A(qq_in414), .Y(Out_data[92]));
CLKBUFX1 gbuf_d_415(.A(N3163), .Y(ddout__415));
CLKBUFX1 gbuf_q_415(.A(qq_in415), .Y(b_in[92]));
CLKBUFX1 gbuf_d_416(.A(N3035), .Y(ddout__416));
CLKBUFX1 gbuf_q_416(.A(qq_in416), .Y(z_in[92]));
CLKBUFX1 gbuf_d_417(.A(n5608), .Y(ddout__417));
CLKBUFX1 gbuf_q_417(.A(qq_in417), .Y(Out_data[93]));
CLKBUFX1 gbuf_d_418(.A(N3164), .Y(ddout__418));
CLKBUFX1 gbuf_q_418(.A(qq_in418), .Y(b_in[93]));
CLKBUFX1 gbuf_d_419(.A(N3036), .Y(ddout__419));
CLKBUFX1 gbuf_q_419(.A(qq_in419), .Y(z_in[93]));
CLKBUFX1 gbuf_d_420(.A(n5607), .Y(ddout__420));
CLKBUFX1 gbuf_q_420(.A(qq_in420), .Y(Out_data[94]));
CLKBUFX1 gbuf_d_421(.A(N3165), .Y(ddout__421));
CLKBUFX1 gbuf_q_421(.A(qq_in421), .Y(b_in[94]));
CLKBUFX1 gbuf_d_422(.A(N3037), .Y(ddout__422));
CLKBUFX1 gbuf_q_422(.A(qq_in422), .Y(z_in[94]));
CLKBUFX1 gbuf_d_423(.A(n5606), .Y(ddout__423));
CLKBUFX1 gbuf_q_423(.A(qq_in423), .Y(Out_data[95]));
CLKBUFX1 gbuf_d_424(.A(N3166), .Y(ddout__424));
CLKBUFX1 gbuf_q_424(.A(qq_in424), .Y(b_in[95]));
CLKBUFX1 gbuf_d_425(.A(N3038), .Y(ddout__425));
CLKBUFX1 gbuf_q_425(.A(qq_in425), .Y(z_in[95]));
CLKBUFX1 gbuf_d_426(.A(n5605), .Y(ddout__426));
CLKBUFX1 gbuf_q_426(.A(qq_in426), .Y(Out_data[96]));
CLKBUFX1 gbuf_d_427(.A(N3167), .Y(ddout__427));
CLKBUFX1 gbuf_q_427(.A(qq_in427), .Y(b_in[96]));
CLKBUFX1 gbuf_d_428(.A(N3039), .Y(ddout__428));
CLKBUFX1 gbuf_q_428(.A(qq_in428), .Y(z_in[96]));
CLKBUFX1 gbuf_d_429(.A(n5604), .Y(ddout__429));
CLKBUFX1 gbuf_q_429(.A(qq_in429), .Y(Out_data[97]));
CLKBUFX1 gbuf_d_430(.A(N3168), .Y(ddout__430));
CLKBUFX1 gbuf_q_430(.A(qq_in430), .Y(b_in[97]));
CLKBUFX1 gbuf_d_431(.A(N3040), .Y(ddout__431));
CLKBUFX1 gbuf_q_431(.A(qq_in431), .Y(z_in[97]));
CLKBUFX1 gbuf_d_432(.A(n5603), .Y(ddout__432));
CLKBUFX1 gbuf_q_432(.A(qq_in432), .Y(Out_data[98]));
CLKBUFX1 gbuf_d_433(.A(N3169), .Y(ddout__433));
CLKBUFX1 gbuf_q_433(.A(qq_in433), .Y(b_in[98]));
CLKBUFX1 gbuf_d_434(.A(N3041), .Y(ddout__434));
CLKBUFX1 gbuf_q_434(.A(qq_in434), .Y(z_in[98]));
CLKBUFX1 gbuf_d_435(.A(n5602), .Y(ddout__435));
CLKBUFX1 gbuf_q_435(.A(qq_in435), .Y(Out_data[99]));
CLKBUFX1 gbuf_d_436(.A(N3170), .Y(ddout__436));
CLKBUFX1 gbuf_q_436(.A(qq_in436), .Y(b_in[99]));
CLKBUFX1 gbuf_d_437(.A(N3042), .Y(ddout__437));
CLKBUFX1 gbuf_q_437(.A(qq_in437), .Y(z_in[99]));
CLKBUFX1 gbuf_d_438(.A(n5601), .Y(ddout__438));
CLKBUFX1 gbuf_q_438(.A(qq_in438), .Y(Out_data[100]));
CLKBUFX1 gbuf_d_439(.A(N3171), .Y(ddout__439));
CLKBUFX1 gbuf_q_439(.A(qq_in439), .Y(b_in[100]));
CLKBUFX1 gbuf_d_440(.A(N3043), .Y(ddout__440));
CLKBUFX1 gbuf_q_440(.A(qq_in440), .Y(z_in[100]));
CLKBUFX1 gbuf_d_441(.A(n5600), .Y(ddout__441));
CLKBUFX1 gbuf_q_441(.A(qq_in441), .Y(Out_data[101]));
CLKBUFX1 gbuf_d_442(.A(N3172), .Y(ddout__442));
CLKBUFX1 gbuf_q_442(.A(qq_in442), .Y(b_in[101]));
CLKBUFX1 gbuf_d_443(.A(N3044), .Y(ddout__443));
CLKBUFX1 gbuf_q_443(.A(qq_in443), .Y(z_in[101]));
CLKBUFX1 gbuf_d_444(.A(n5599), .Y(ddout__444));
CLKBUFX1 gbuf_q_444(.A(qq_in444), .Y(Out_data[102]));
CLKBUFX1 gbuf_d_445(.A(N3173), .Y(ddout__445));
CLKBUFX1 gbuf_q_445(.A(qq_in445), .Y(b_in[102]));
CLKBUFX1 gbuf_d_446(.A(N3045), .Y(ddout__446));
CLKBUFX1 gbuf_q_446(.A(qq_in446), .Y(z_in[102]));
CLKBUFX1 gbuf_d_447(.A(n5598), .Y(ddout__447));
CLKBUFX1 gbuf_q_447(.A(qq_in447), .Y(Out_data[103]));
CLKBUFX1 gbuf_d_448(.A(N3174), .Y(ddout__448));
CLKBUFX1 gbuf_q_448(.A(qq_in448), .Y(b_in[103]));
CLKBUFX1 gbuf_d_449(.A(N3046), .Y(ddout__449));
CLKBUFX1 gbuf_q_449(.A(qq_in449), .Y(z_in[103]));
CLKBUFX1 gbuf_d_450(.A(n5597), .Y(ddout__450));
CLKBUFX1 gbuf_q_450(.A(qq_in450), .Y(Out_data[104]));
CLKBUFX1 gbuf_d_451(.A(N3175), .Y(ddout__451));
CLKBUFX1 gbuf_q_451(.A(qq_in451), .Y(b_in[104]));
CLKBUFX1 gbuf_d_452(.A(N3047), .Y(ddout__452));
CLKBUFX1 gbuf_q_452(.A(qq_in452), .Y(z_in[104]));
CLKBUFX1 gbuf_d_453(.A(n5596), .Y(ddout__453));
CLKBUFX1 gbuf_q_453(.A(qq_in453), .Y(Out_data[105]));
CLKBUFX1 gbuf_d_454(.A(N3176), .Y(ddout__454));
CLKBUFX1 gbuf_q_454(.A(qq_in454), .Y(b_in[105]));
CLKBUFX1 gbuf_d_455(.A(N3048), .Y(ddout__455));
CLKBUFX1 gbuf_q_455(.A(qq_in455), .Y(z_in[105]));
CLKBUFX1 gbuf_d_456(.A(n5595), .Y(ddout__456));
CLKBUFX1 gbuf_q_456(.A(qq_in456), .Y(Out_data[106]));
CLKBUFX1 gbuf_d_457(.A(N3177), .Y(ddout__457));
CLKBUFX1 gbuf_q_457(.A(qq_in457), .Y(b_in[106]));
CLKBUFX1 gbuf_d_458(.A(N3049), .Y(ddout__458));
CLKBUFX1 gbuf_q_458(.A(qq_in458), .Y(z_in[106]));
CLKBUFX1 gbuf_d_459(.A(n5594), .Y(ddout__459));
CLKBUFX1 gbuf_q_459(.A(qq_in459), .Y(Out_data[107]));
CLKBUFX1 gbuf_d_460(.A(N3178), .Y(ddout__460));
CLKBUFX1 gbuf_q_460(.A(qq_in460), .Y(b_in[107]));
CLKBUFX1 gbuf_d_461(.A(N3050), .Y(ddout__461));
CLKBUFX1 gbuf_q_461(.A(qq_in461), .Y(z_in[107]));
CLKBUFX1 gbuf_d_462(.A(n5593), .Y(ddout__462));
CLKBUFX1 gbuf_q_462(.A(qq_in462), .Y(Out_data[108]));
CLKBUFX1 gbuf_d_463(.A(N3179), .Y(ddout__463));
CLKBUFX1 gbuf_q_463(.A(qq_in463), .Y(b_in[108]));
CLKBUFX1 gbuf_d_464(.A(N3051), .Y(ddout__464));
CLKBUFX1 gbuf_q_464(.A(qq_in464), .Y(z_in[108]));
CLKBUFX1 gbuf_d_465(.A(n5592), .Y(ddout__465));
CLKBUFX1 gbuf_q_465(.A(qq_in465), .Y(Out_data[109]));
CLKBUFX1 gbuf_d_466(.A(N3180), .Y(ddout__466));
CLKBUFX1 gbuf_q_466(.A(qq_in466), .Y(b_in[109]));
CLKBUFX1 gbuf_d_467(.A(N3052), .Y(ddout__467));
CLKBUFX1 gbuf_q_467(.A(qq_in467), .Y(z_in[109]));
CLKBUFX1 gbuf_d_468(.A(n5591), .Y(ddout__468));
CLKBUFX1 gbuf_q_468(.A(qq_in468), .Y(Out_data[110]));
CLKBUFX1 gbuf_d_469(.A(N3181), .Y(ddout__469));
CLKBUFX1 gbuf_q_469(.A(qq_in469), .Y(b_in[110]));
CLKBUFX1 gbuf_d_470(.A(N3053), .Y(ddout__470));
CLKBUFX1 gbuf_q_470(.A(qq_in470), .Y(z_in[110]));
CLKBUFX1 gbuf_d_471(.A(n5590), .Y(ddout__471));
CLKBUFX1 gbuf_q_471(.A(qq_in471), .Y(Out_data[111]));
CLKBUFX1 gbuf_d_472(.A(N3182), .Y(ddout__472));
CLKBUFX1 gbuf_q_472(.A(qq_in472), .Y(b_in[111]));
CLKBUFX1 gbuf_d_473(.A(N3054), .Y(ddout__473));
CLKBUFX1 gbuf_q_473(.A(qq_in473), .Y(z_in[111]));
CLKBUFX1 gbuf_d_474(.A(n5589), .Y(ddout__474));
CLKBUFX1 gbuf_q_474(.A(qq_in474), .Y(Out_data[112]));
CLKBUFX1 gbuf_d_475(.A(N3183), .Y(ddout__475));
CLKBUFX1 gbuf_q_475(.A(qq_in475), .Y(b_in[112]));
CLKBUFX1 gbuf_d_476(.A(N3055), .Y(ddout__476));
CLKBUFX1 gbuf_q_476(.A(qq_in476), .Y(z_in[112]));
CLKBUFX1 gbuf_d_477(.A(n5588), .Y(ddout__477));
CLKBUFX1 gbuf_q_477(.A(qq_in477), .Y(Out_data[113]));
CLKBUFX1 gbuf_d_478(.A(N3184), .Y(ddout__478));
CLKBUFX1 gbuf_q_478(.A(qq_in478), .Y(b_in[113]));
CLKBUFX1 gbuf_d_479(.A(N3056), .Y(ddout__479));
CLKBUFX1 gbuf_q_479(.A(qq_in479), .Y(z_in[113]));
CLKBUFX1 gbuf_d_480(.A(n5587), .Y(ddout__480));
CLKBUFX1 gbuf_q_480(.A(qq_in480), .Y(Out_data[114]));
CLKBUFX1 gbuf_d_481(.A(N3185), .Y(ddout__481));
CLKBUFX1 gbuf_q_481(.A(qq_in481), .Y(b_in[114]));
CLKBUFX1 gbuf_d_482(.A(N3057), .Y(ddout__482));
CLKBUFX1 gbuf_q_482(.A(qq_in482), .Y(z_in[114]));
CLKBUFX1 gbuf_d_483(.A(n5586), .Y(ddout__483));
CLKBUFX1 gbuf_q_483(.A(qq_in483), .Y(Out_data[115]));
CLKBUFX1 gbuf_d_484(.A(N3186), .Y(ddout__484));
CLKBUFX1 gbuf_q_484(.A(qq_in484), .Y(b_in[115]));
CLKBUFX1 gbuf_d_485(.A(N3058), .Y(ddout__485));
CLKBUFX1 gbuf_q_485(.A(qq_in485), .Y(z_in[115]));
CLKBUFX1 gbuf_d_486(.A(n5585), .Y(ddout__486));
CLKBUFX1 gbuf_q_486(.A(qq_in486), .Y(Out_data[116]));
CLKBUFX1 gbuf_d_487(.A(N3187), .Y(ddout__487));
CLKBUFX1 gbuf_q_487(.A(qq_in487), .Y(b_in[116]));
CLKBUFX1 gbuf_d_488(.A(N3059), .Y(ddout__488));
CLKBUFX1 gbuf_q_488(.A(qq_in488), .Y(z_in[116]));
CLKBUFX1 gbuf_d_489(.A(n5584), .Y(ddout__489));
CLKBUFX1 gbuf_q_489(.A(qq_in489), .Y(Out_data[117]));
CLKBUFX1 gbuf_d_490(.A(N3188), .Y(ddout__490));
CLKBUFX1 gbuf_q_490(.A(qq_in490), .Y(b_in[117]));
CLKBUFX1 gbuf_d_491(.A(N3060), .Y(ddout__491));
CLKBUFX1 gbuf_q_491(.A(qq_in491), .Y(z_in[117]));
CLKBUFX1 gbuf_d_492(.A(n5583), .Y(ddout__492));
CLKBUFX1 gbuf_q_492(.A(qq_in492), .Y(Out_data[118]));
CLKBUFX1 gbuf_d_493(.A(N3189), .Y(ddout__493));
CLKBUFX1 gbuf_q_493(.A(qq_in493), .Y(b_in[118]));
CLKBUFX1 gbuf_d_494(.A(N3061), .Y(ddout__494));
CLKBUFX1 gbuf_q_494(.A(qq_in494), .Y(z_in[118]));
CLKBUFX1 gbuf_d_495(.A(n5582), .Y(ddout__495));
CLKBUFX1 gbuf_q_495(.A(qq_in495), .Y(Out_data[119]));
CLKBUFX1 gbuf_d_496(.A(N3190), .Y(ddout__496));
CLKBUFX1 gbuf_q_496(.A(qq_in496), .Y(b_in[119]));
CLKBUFX1 gbuf_d_497(.A(N3062), .Y(ddout__497));
CLKBUFX1 gbuf_q_497(.A(qq_in497), .Y(z_in[119]));
CLKBUFX1 gbuf_d_498(.A(n5581), .Y(ddout__498));
CLKBUFX1 gbuf_q_498(.A(qq_in498), .Y(Out_data[120]));
CLKBUFX1 gbuf_d_499(.A(N3191), .Y(ddout__499));
CLKBUFX1 gbuf_q_499(.A(qq_in499), .Y(b_in[120]));
CLKBUFX1 gbuf_d_500(.A(N3063), .Y(ddout__500));
CLKBUFX1 gbuf_q_500(.A(qq_in500), .Y(z_in[120]));
CLKBUFX1 gbuf_d_501(.A(n5580), .Y(ddout__501));
CLKBUFX1 gbuf_q_501(.A(qq_in501), .Y(Out_data[121]));
CLKBUFX1 gbuf_d_502(.A(N3192), .Y(ddout__502));
CLKBUFX1 gbuf_q_502(.A(qq_in502), .Y(b_in[121]));
CLKBUFX1 gbuf_d_503(.A(N3064), .Y(ddout__503));
CLKBUFX1 gbuf_q_503(.A(qq_in503), .Y(z_in[121]));
CLKBUFX1 gbuf_d_504(.A(n5579), .Y(ddout__504));
CLKBUFX1 gbuf_q_504(.A(qq_in504), .Y(Out_data[122]));
CLKBUFX1 gbuf_d_505(.A(N3193), .Y(ddout__505));
CLKBUFX1 gbuf_q_505(.A(qq_in505), .Y(b_in[122]));
CLKBUFX1 gbuf_d_506(.A(N3065), .Y(ddout__506));
CLKBUFX1 gbuf_q_506(.A(qq_in506), .Y(z_in[122]));
CLKBUFX1 gbuf_d_507(.A(n5578), .Y(ddout__507));
CLKBUFX1 gbuf_q_507(.A(qq_in507), .Y(Out_data[123]));
CLKBUFX1 gbuf_d_508(.A(N3194), .Y(ddout__508));
CLKBUFX1 gbuf_q_508(.A(qq_in508), .Y(b_in[123]));
CLKBUFX1 gbuf_d_509(.A(N3066), .Y(ddout__509));
CLKBUFX1 gbuf_q_509(.A(qq_in509), .Y(z_in[123]));
CLKBUFX1 gbuf_d_510(.A(n5577), .Y(ddout__510));
CLKBUFX1 gbuf_q_510(.A(qq_in510), .Y(Out_data[124]));
CLKBUFX1 gbuf_d_511(.A(N3195), .Y(ddout__511));
CLKBUFX1 gbuf_q_511(.A(qq_in511), .Y(b_in[124]));
CLKBUFX1 gbuf_d_512(.A(N3067), .Y(ddout__512));
CLKBUFX1 gbuf_q_512(.A(qq_in512), .Y(z_in[124]));
CLKBUFX1 gbuf_d_513(.A(n5576), .Y(ddout__513));
CLKBUFX1 gbuf_q_513(.A(qq_in513), .Y(Out_data[125]));
CLKBUFX1 gbuf_d_514(.A(N3196), .Y(ddout__514));
CLKBUFX1 gbuf_q_514(.A(qq_in514), .Y(b_in[125]));
CLKBUFX1 gbuf_d_515(.A(N3068), .Y(ddout__515));
CLKBUFX1 gbuf_q_515(.A(qq_in515), .Y(z_in[125]));
CLKBUFX1 gbuf_d_516(.A(n5575), .Y(ddout__516));
CLKBUFX1 gbuf_q_516(.A(qq_in516), .Y(Out_data[126]));
CLKBUFX1 gbuf_d_517(.A(N3197), .Y(ddout__517));
CLKBUFX1 gbuf_q_517(.A(qq_in517), .Y(b_in[126]));
CLKBUFX1 gbuf_d_518(.A(N3069), .Y(ddout__518));
CLKBUFX1 gbuf_q_518(.A(qq_in518), .Y(z_in[126]));
CLKBUFX1 gbuf_d_519(.A(n5574), .Y(ddout__519));
CLKBUFX1 gbuf_q_519(.A(qq_in519), .Y(Out_data[127]));
CLKBUFX1 gbuf_d_520(.A(N3198), .Y(ddout__520));
CLKBUFX1 gbuf_q_520(.A(qq_in520), .Y(b_in[127]));
CLKBUFX1 gbuf_d_521(.A(N3070), .Y(ddout__521));
CLKBUFX1 gbuf_q_521(.A(qq_in521), .Y(z_in[127]));
CLKBUFX1 gbuf_d_522(.A(N2816), .Y(ddout__522));
CLKBUFX1 gbuf_q_522(.A(qq_in522), .Y(v_in[1]));
CLKBUFX1 gbuf_d_523(.A(N2817), .Y(ddout__523));
CLKBUFX1 gbuf_q_523(.A(qq_in523), .Y(v_in[2]));
CLKBUFX1 gbuf_d_524(.A(N2818), .Y(ddout__524));
CLKBUFX1 gbuf_q_524(.A(qq_in524), .Y(v_in[3]));
CLKBUFX1 gbuf_d_525(.A(N2819), .Y(ddout__525));
CLKBUFX1 gbuf_q_525(.A(qq_in525), .Y(v_in[4]));
CLKBUFX1 gbuf_d_526(.A(N2820), .Y(ddout__526));
CLKBUFX1 gbuf_q_526(.A(qq_in526), .Y(v_in[5]));
CLKBUFX1 gbuf_d_527(.A(N2821), .Y(ddout__527));
CLKBUFX1 gbuf_q_527(.A(qq_in527), .Y(v_in[6]));
CLKBUFX1 gbuf_d_528(.A(N2822), .Y(ddout__528));
CLKBUFX1 gbuf_q_528(.A(qq_in528), .Y(v_in[7]));
CLKBUFX1 gbuf_d_529(.A(N2823), .Y(ddout__529));
CLKBUFX1 gbuf_q_529(.A(qq_in529), .Y(v_in[8]));
CLKBUFX1 gbuf_d_530(.A(N2824), .Y(ddout__530));
CLKBUFX1 gbuf_q_530(.A(qq_in530), .Y(v_in[9]));
CLKBUFX1 gbuf_d_531(.A(N2825), .Y(ddout__531));
CLKBUFX1 gbuf_q_531(.A(qq_in531), .Y(v_in[10]));
CLKBUFX1 gbuf_d_532(.A(N2826), .Y(ddout__532));
CLKBUFX1 gbuf_q_532(.A(qq_in532), .Y(v_in[11]));
CLKBUFX1 gbuf_d_533(.A(N2827), .Y(ddout__533));
CLKBUFX1 gbuf_q_533(.A(qq_in533), .Y(v_in[12]));
CLKBUFX1 gbuf_d_534(.A(N2828), .Y(ddout__534));
CLKBUFX1 gbuf_q_534(.A(qq_in534), .Y(v_in[13]));
CLKBUFX1 gbuf_d_535(.A(N2829), .Y(ddout__535));
CLKBUFX1 gbuf_q_535(.A(qq_in535), .Y(v_in[14]));
CLKBUFX1 gbuf_d_536(.A(N2830), .Y(ddout__536));
CLKBUFX1 gbuf_q_536(.A(qq_in536), .Y(v_in[15]));
CLKBUFX1 gbuf_d_537(.A(N2831), .Y(ddout__537));
CLKBUFX1 gbuf_q_537(.A(qq_in537), .Y(v_in[16]));
CLKBUFX1 gbuf_d_538(.A(N2832), .Y(ddout__538));
CLKBUFX1 gbuf_q_538(.A(qq_in538), .Y(v_in[17]));
CLKBUFX1 gbuf_d_539(.A(N2833), .Y(ddout__539));
CLKBUFX1 gbuf_q_539(.A(qq_in539), .Y(v_in[18]));
CLKBUFX1 gbuf_d_540(.A(N2834), .Y(ddout__540));
CLKBUFX1 gbuf_q_540(.A(qq_in540), .Y(v_in[19]));
CLKBUFX1 gbuf_d_541(.A(N2835), .Y(ddout__541));
CLKBUFX1 gbuf_q_541(.A(qq_in541), .Y(v_in[20]));
CLKBUFX1 gbuf_d_542(.A(N2836), .Y(ddout__542));
CLKBUFX1 gbuf_q_542(.A(qq_in542), .Y(v_in[21]));
CLKBUFX1 gbuf_d_543(.A(N2837), .Y(ddout__543));
CLKBUFX1 gbuf_q_543(.A(qq_in543), .Y(v_in[22]));
CLKBUFX1 gbuf_d_544(.A(N2838), .Y(ddout__544));
CLKBUFX1 gbuf_q_544(.A(qq_in544), .Y(v_in[23]));
CLKBUFX1 gbuf_d_545(.A(N2839), .Y(ddout__545));
CLKBUFX1 gbuf_q_545(.A(qq_in545), .Y(v_in[24]));
CLKBUFX1 gbuf_d_546(.A(N2840), .Y(ddout__546));
CLKBUFX1 gbuf_q_546(.A(qq_in546), .Y(v_in[25]));
CLKBUFX1 gbuf_d_547(.A(N2841), .Y(ddout__547));
CLKBUFX1 gbuf_q_547(.A(qq_in547), .Y(v_in[26]));
CLKBUFX1 gbuf_d_548(.A(N2842), .Y(ddout__548));
CLKBUFX1 gbuf_q_548(.A(qq_in548), .Y(v_in[27]));
CLKBUFX1 gbuf_d_549(.A(N2843), .Y(ddout__549));
CLKBUFX1 gbuf_q_549(.A(qq_in549), .Y(v_in[28]));
CLKBUFX1 gbuf_d_550(.A(N2844), .Y(ddout__550));
CLKBUFX1 gbuf_q_550(.A(qq_in550), .Y(v_in[29]));
CLKBUFX1 gbuf_d_551(.A(N2845), .Y(ddout__551));
CLKBUFX1 gbuf_q_551(.A(qq_in551), .Y(v_in[30]));
CLKBUFX1 gbuf_d_552(.A(N2846), .Y(ddout__552));
CLKBUFX1 gbuf_q_552(.A(qq_in552), .Y(v_in[31]));
CLKBUFX1 gbuf_d_553(.A(N2847), .Y(ddout__553));
CLKBUFX1 gbuf_q_553(.A(qq_in553), .Y(v_in[32]));
CLKBUFX1 gbuf_d_554(.A(N2848), .Y(ddout__554));
CLKBUFX1 gbuf_q_554(.A(qq_in554), .Y(v_in[33]));
CLKBUFX1 gbuf_d_555(.A(N2849), .Y(ddout__555));
CLKBUFX1 gbuf_q_555(.A(qq_in555), .Y(v_in[34]));
CLKBUFX1 gbuf_d_556(.A(N2850), .Y(ddout__556));
CLKBUFX1 gbuf_q_556(.A(qq_in556), .Y(v_in[35]));
CLKBUFX1 gbuf_d_557(.A(N2851), .Y(ddout__557));
CLKBUFX1 gbuf_q_557(.A(qq_in557), .Y(v_in[36]));
CLKBUFX1 gbuf_d_558(.A(N2852), .Y(ddout__558));
CLKBUFX1 gbuf_q_558(.A(qq_in558), .Y(v_in[37]));
CLKBUFX1 gbuf_d_559(.A(N2853), .Y(ddout__559));
CLKBUFX1 gbuf_q_559(.A(qq_in559), .Y(v_in[38]));
CLKBUFX1 gbuf_d_560(.A(N2854), .Y(ddout__560));
CLKBUFX1 gbuf_q_560(.A(qq_in560), .Y(v_in[39]));
CLKBUFX1 gbuf_d_561(.A(N2855), .Y(ddout__561));
CLKBUFX1 gbuf_q_561(.A(qq_in561), .Y(v_in[40]));
CLKBUFX1 gbuf_d_562(.A(N2856), .Y(ddout__562));
CLKBUFX1 gbuf_q_562(.A(qq_in562), .Y(v_in[41]));
CLKBUFX1 gbuf_d_563(.A(N2857), .Y(ddout__563));
CLKBUFX1 gbuf_q_563(.A(qq_in563), .Y(v_in[42]));
CLKBUFX1 gbuf_d_564(.A(N2858), .Y(ddout__564));
CLKBUFX1 gbuf_q_564(.A(qq_in564), .Y(v_in[43]));
CLKBUFX1 gbuf_d_565(.A(N2859), .Y(ddout__565));
CLKBUFX1 gbuf_q_565(.A(qq_in565), .Y(v_in[44]));
CLKBUFX1 gbuf_d_566(.A(N2860), .Y(ddout__566));
CLKBUFX1 gbuf_q_566(.A(qq_in566), .Y(v_in[45]));
CLKBUFX1 gbuf_d_567(.A(N2861), .Y(ddout__567));
CLKBUFX1 gbuf_q_567(.A(qq_in567), .Y(v_in[46]));
CLKBUFX1 gbuf_d_568(.A(N2862), .Y(ddout__568));
CLKBUFX1 gbuf_q_568(.A(qq_in568), .Y(v_in[47]));
CLKBUFX1 gbuf_d_569(.A(N2863), .Y(ddout__569));
CLKBUFX1 gbuf_q_569(.A(qq_in569), .Y(v_in[48]));
CLKBUFX1 gbuf_d_570(.A(N2864), .Y(ddout__570));
CLKBUFX1 gbuf_q_570(.A(qq_in570), .Y(v_in[49]));
CLKBUFX1 gbuf_d_571(.A(N2865), .Y(ddout__571));
CLKBUFX1 gbuf_q_571(.A(qq_in571), .Y(v_in[50]));
CLKBUFX1 gbuf_d_572(.A(N2866), .Y(ddout__572));
CLKBUFX1 gbuf_q_572(.A(qq_in572), .Y(v_in[51]));
CLKBUFX1 gbuf_d_573(.A(N2867), .Y(ddout__573));
CLKBUFX1 gbuf_q_573(.A(qq_in573), .Y(v_in[52]));
CLKBUFX1 gbuf_d_574(.A(N2868), .Y(ddout__574));
CLKBUFX1 gbuf_q_574(.A(qq_in574), .Y(v_in[53]));
CLKBUFX1 gbuf_d_575(.A(N2869), .Y(ddout__575));
CLKBUFX1 gbuf_q_575(.A(qq_in575), .Y(v_in[54]));
CLKBUFX1 gbuf_d_576(.A(N2870), .Y(ddout__576));
CLKBUFX1 gbuf_q_576(.A(qq_in576), .Y(v_in[55]));
CLKBUFX1 gbuf_d_577(.A(N2871), .Y(ddout__577));
CLKBUFX1 gbuf_q_577(.A(qq_in577), .Y(v_in[56]));
CLKBUFX1 gbuf_d_578(.A(N2872), .Y(ddout__578));
CLKBUFX1 gbuf_q_578(.A(qq_in578), .Y(v_in[57]));
CLKBUFX1 gbuf_d_579(.A(N2873), .Y(ddout__579));
CLKBUFX1 gbuf_q_579(.A(qq_in579), .Y(v_in[58]));
CLKBUFX1 gbuf_d_580(.A(N2874), .Y(ddout__580));
CLKBUFX1 gbuf_q_580(.A(qq_in580), .Y(v_in[59]));
CLKBUFX1 gbuf_d_581(.A(N2875), .Y(ddout__581));
CLKBUFX1 gbuf_q_581(.A(qq_in581), .Y(v_in[60]));
CLKBUFX1 gbuf_d_582(.A(N2876), .Y(ddout__582));
CLKBUFX1 gbuf_q_582(.A(qq_in582), .Y(v_in[61]));
CLKBUFX1 gbuf_d_583(.A(N2877), .Y(ddout__583));
CLKBUFX1 gbuf_q_583(.A(qq_in583), .Y(v_in[62]));
CLKBUFX1 gbuf_d_584(.A(N2878), .Y(ddout__584));
CLKBUFX1 gbuf_q_584(.A(qq_in584), .Y(v_in[63]));
CLKBUFX1 gbuf_d_585(.A(N2879), .Y(ddout__585));
CLKBUFX1 gbuf_q_585(.A(qq_in585), .Y(v_in[64]));
CLKBUFX1 gbuf_d_586(.A(N2880), .Y(ddout__586));
CLKBUFX1 gbuf_q_586(.A(qq_in586), .Y(v_in[65]));
CLKBUFX1 gbuf_d_587(.A(N2881), .Y(ddout__587));
CLKBUFX1 gbuf_q_587(.A(qq_in587), .Y(v_in[66]));
CLKBUFX1 gbuf_d_588(.A(N2882), .Y(ddout__588));
CLKBUFX1 gbuf_q_588(.A(qq_in588), .Y(v_in[67]));
CLKBUFX1 gbuf_d_589(.A(N2883), .Y(ddout__589));
CLKBUFX1 gbuf_q_589(.A(qq_in589), .Y(v_in[68]));
CLKBUFX1 gbuf_d_590(.A(N2884), .Y(ddout__590));
CLKBUFX1 gbuf_q_590(.A(qq_in590), .Y(v_in[69]));
CLKBUFX1 gbuf_d_591(.A(N2885), .Y(ddout__591));
CLKBUFX1 gbuf_q_591(.A(qq_in591), .Y(v_in[70]));
CLKBUFX1 gbuf_d_592(.A(N2886), .Y(ddout__592));
CLKBUFX1 gbuf_q_592(.A(qq_in592), .Y(v_in[71]));
CLKBUFX1 gbuf_d_593(.A(N2887), .Y(ddout__593));
CLKBUFX1 gbuf_q_593(.A(qq_in593), .Y(v_in[72]));
CLKBUFX1 gbuf_d_594(.A(N2888), .Y(ddout__594));
CLKBUFX1 gbuf_q_594(.A(qq_in594), .Y(v_in[73]));
CLKBUFX1 gbuf_d_595(.A(N2889), .Y(ddout__595));
CLKBUFX1 gbuf_q_595(.A(qq_in595), .Y(v_in[74]));
CLKBUFX1 gbuf_d_596(.A(N2890), .Y(ddout__596));
CLKBUFX1 gbuf_q_596(.A(qq_in596), .Y(v_in[75]));
CLKBUFX1 gbuf_d_597(.A(N2891), .Y(ddout__597));
CLKBUFX1 gbuf_q_597(.A(qq_in597), .Y(v_in[76]));
CLKBUFX1 gbuf_d_598(.A(N2892), .Y(ddout__598));
CLKBUFX1 gbuf_q_598(.A(qq_in598), .Y(v_in[77]));
CLKBUFX1 gbuf_d_599(.A(N2893), .Y(ddout__599));
CLKBUFX1 gbuf_q_599(.A(qq_in599), .Y(v_in[78]));
CLKBUFX1 gbuf_d_600(.A(N2894), .Y(ddout__600));
CLKBUFX1 gbuf_q_600(.A(qq_in600), .Y(v_in[79]));
CLKBUFX1 gbuf_d_601(.A(N2895), .Y(ddout__601));
CLKBUFX1 gbuf_q_601(.A(qq_in601), .Y(v_in[80]));
CLKBUFX1 gbuf_d_602(.A(N2896), .Y(ddout__602));
CLKBUFX1 gbuf_q_602(.A(qq_in602), .Y(v_in[81]));
CLKBUFX1 gbuf_d_603(.A(N2897), .Y(ddout__603));
CLKBUFX1 gbuf_q_603(.A(qq_in603), .Y(v_in[82]));
CLKBUFX1 gbuf_d_604(.A(N2898), .Y(ddout__604));
CLKBUFX1 gbuf_q_604(.A(qq_in604), .Y(v_in[83]));
CLKBUFX1 gbuf_d_605(.A(N2899), .Y(ddout__605));
CLKBUFX1 gbuf_q_605(.A(qq_in605), .Y(v_in[84]));
CLKBUFX1 gbuf_d_606(.A(N2900), .Y(ddout__606));
CLKBUFX1 gbuf_q_606(.A(qq_in606), .Y(v_in[85]));
CLKBUFX1 gbuf_d_607(.A(N2901), .Y(ddout__607));
CLKBUFX1 gbuf_q_607(.A(qq_in607), .Y(v_in[86]));
CLKBUFX1 gbuf_d_608(.A(N2902), .Y(ddout__608));
CLKBUFX1 gbuf_q_608(.A(qq_in608), .Y(v_in[87]));
CLKBUFX1 gbuf_d_609(.A(N2903), .Y(ddout__609));
CLKBUFX1 gbuf_q_609(.A(qq_in609), .Y(v_in[88]));
CLKBUFX1 gbuf_d_610(.A(N2904), .Y(ddout__610));
CLKBUFX1 gbuf_q_610(.A(qq_in610), .Y(v_in[89]));
CLKBUFX1 gbuf_d_611(.A(N2905), .Y(ddout__611));
CLKBUFX1 gbuf_q_611(.A(qq_in611), .Y(v_in[90]));
CLKBUFX1 gbuf_d_612(.A(N2906), .Y(ddout__612));
CLKBUFX1 gbuf_q_612(.A(qq_in612), .Y(v_in[91]));
CLKBUFX1 gbuf_d_613(.A(N2907), .Y(ddout__613));
CLKBUFX1 gbuf_q_613(.A(qq_in613), .Y(v_in[92]));
CLKBUFX1 gbuf_d_614(.A(N2908), .Y(ddout__614));
CLKBUFX1 gbuf_q_614(.A(qq_in614), .Y(v_in[93]));
CLKBUFX1 gbuf_d_615(.A(N2909), .Y(ddout__615));
CLKBUFX1 gbuf_q_615(.A(qq_in615), .Y(v_in[94]));
CLKBUFX1 gbuf_d_616(.A(N2910), .Y(ddout__616));
CLKBUFX1 gbuf_q_616(.A(qq_in616), .Y(v_in[95]));
CLKBUFX1 gbuf_d_617(.A(N2911), .Y(ddout__617));
CLKBUFX1 gbuf_q_617(.A(qq_in617), .Y(v_in[96]));
CLKBUFX1 gbuf_d_618(.A(N2912), .Y(ddout__618));
CLKBUFX1 gbuf_q_618(.A(qq_in618), .Y(v_in[97]));
CLKBUFX1 gbuf_d_619(.A(N2913), .Y(ddout__619));
CLKBUFX1 gbuf_q_619(.A(qq_in619), .Y(v_in[98]));
CLKBUFX1 gbuf_d_620(.A(N2914), .Y(ddout__620));
CLKBUFX1 gbuf_q_620(.A(qq_in620), .Y(v_in[99]));
CLKBUFX1 gbuf_d_621(.A(N2915), .Y(ddout__621));
CLKBUFX1 gbuf_q_621(.A(qq_in621), .Y(v_in[100]));
CLKBUFX1 gbuf_d_622(.A(N2916), .Y(ddout__622));
CLKBUFX1 gbuf_q_622(.A(qq_in622), .Y(v_in[101]));
CLKBUFX1 gbuf_d_623(.A(N2917), .Y(ddout__623));
CLKBUFX1 gbuf_q_623(.A(qq_in623), .Y(v_in[102]));
CLKBUFX1 gbuf_d_624(.A(N2918), .Y(ddout__624));
CLKBUFX1 gbuf_q_624(.A(qq_in624), .Y(v_in[103]));
CLKBUFX1 gbuf_d_625(.A(N2919), .Y(ddout__625));
CLKBUFX1 gbuf_q_625(.A(qq_in625), .Y(v_in[104]));
CLKBUFX1 gbuf_d_626(.A(N2920), .Y(ddout__626));
CLKBUFX1 gbuf_q_626(.A(qq_in626), .Y(v_in[105]));
CLKBUFX1 gbuf_d_627(.A(N2921), .Y(ddout__627));
CLKBUFX1 gbuf_q_627(.A(qq_in627), .Y(v_in[106]));
CLKBUFX1 gbuf_d_628(.A(N2922), .Y(ddout__628));
CLKBUFX1 gbuf_q_628(.A(qq_in628), .Y(v_in[107]));
CLKBUFX1 gbuf_d_629(.A(N2923), .Y(ddout__629));
CLKBUFX1 gbuf_q_629(.A(qq_in629), .Y(v_in[108]));
CLKBUFX1 gbuf_d_630(.A(N2924), .Y(ddout__630));
CLKBUFX1 gbuf_q_630(.A(qq_in630), .Y(v_in[109]));
CLKBUFX1 gbuf_d_631(.A(N2925), .Y(ddout__631));
CLKBUFX1 gbuf_q_631(.A(qq_in631), .Y(v_in[110]));
CLKBUFX1 gbuf_d_632(.A(N2926), .Y(ddout__632));
CLKBUFX1 gbuf_q_632(.A(qq_in632), .Y(v_in[111]));
CLKBUFX1 gbuf_d_633(.A(N2927), .Y(ddout__633));
CLKBUFX1 gbuf_q_633(.A(qq_in633), .Y(v_in[112]));
CLKBUFX1 gbuf_d_634(.A(N2928), .Y(ddout__634));
CLKBUFX1 gbuf_q_634(.A(qq_in634), .Y(v_in[113]));
CLKBUFX1 gbuf_d_635(.A(N2929), .Y(ddout__635));
CLKBUFX1 gbuf_q_635(.A(qq_in635), .Y(v_in[114]));
CLKBUFX1 gbuf_d_636(.A(N2930), .Y(ddout__636));
CLKBUFX1 gbuf_q_636(.A(qq_in636), .Y(v_in[115]));
CLKBUFX1 gbuf_d_637(.A(N2931), .Y(ddout__637));
CLKBUFX1 gbuf_q_637(.A(qq_in637), .Y(v_in[116]));
CLKBUFX1 gbuf_d_638(.A(N2932), .Y(ddout__638));
CLKBUFX1 gbuf_q_638(.A(qq_in638), .Y(v_in[117]));
CLKBUFX1 gbuf_d_639(.A(N2933), .Y(ddout__639));
CLKBUFX1 gbuf_q_639(.A(qq_in639), .Y(v_in[118]));
CLKBUFX1 gbuf_d_640(.A(N2934), .Y(ddout__640));
CLKBUFX1 gbuf_q_640(.A(qq_in640), .Y(v_in[119]));
CLKBUFX1 gbuf_d_641(.A(N2935), .Y(ddout__641));
CLKBUFX1 gbuf_q_641(.A(qq_in641), .Y(v_in[120]));
CLKBUFX1 gbuf_d_642(.A(N2936), .Y(ddout__642));
CLKBUFX1 gbuf_q_642(.A(qq_in642), .Y(v_in[121]));
CLKBUFX1 gbuf_d_643(.A(N2937), .Y(ddout__643));
CLKBUFX1 gbuf_q_643(.A(qq_in643), .Y(v_in[122]));
CLKBUFX1 gbuf_d_644(.A(N2938), .Y(ddout__644));
CLKBUFX1 gbuf_q_644(.A(qq_in644), .Y(v_in[123]));
CLKBUFX1 gbuf_d_645(.A(N2939), .Y(ddout__645));
CLKBUFX1 gbuf_q_645(.A(qq_in645), .Y(v_in[124]));
CLKBUFX1 gbuf_d_646(.A(N2940), .Y(ddout__646));
CLKBUFX1 gbuf_q_646(.A(qq_in646), .Y(v_in[125]));
CLKBUFX1 gbuf_d_647(.A(N2941), .Y(ddout__647));
CLKBUFX1 gbuf_q_647(.A(qq_in647), .Y(v_in[126]));
CLKBUFX1 gbuf_d_648(.A(N2942), .Y(ddout__648));
CLKBUFX1 gbuf_q_648(.A(qq_in648), .Y(v_in[127]));
NAND2_X2 U6736 ( .A1(n17747), .A2(n11931), .ZN(n6292) );
NAND2_X2 U6741 ( .A1(n11935), .A2(n11936), .ZN(n6290) );
NAND2_X2 U6743 ( .A1(n11923), .A2(n18893), .ZN(n11935) );
NAND2_X2 U6744 ( .A1(n18745), .A2(n11937), .ZN(n11923) );
NAND2_X2 U6749 ( .A1(n11939), .A2(n11940), .ZN(n6289) );
NAND2_X2 U6752 ( .A1(state[6]), .A2(n11926), .ZN(n11941) );
NAND2_X2 U6753 ( .A1(n11942), .A2(n11943), .ZN(n6287) );
NAND2_X2 U6755 ( .A1(n18747), .A2(n11944), .ZN(n11926) );
NAND2_X2 U6762 ( .A1(n11953), .A2(n11954), .ZN(n11948) );
NAND2_X2 U6763 ( .A1(n11955), .A2(n18892), .ZN(n11954) );
NAND2_X2 U6767 ( .A1(n11961), .A2(n11962), .ZN(n6283) );
NAND2_X2 U6768 ( .A1(state[0]), .A2(n11963), .ZN(n11962) );
NAND2_X2 U6769 ( .A1(n17375), .A2(n11953), .ZN(n11963) );
AND3_X2 U6770 ( .A1(n11964), .A2(n11965), .A3(n11966), .ZN(n11953) );
NAND2_X2 U6773 ( .A1(cii_IV_vld), .A2(aes_done), .ZN(n11968) );
NAND2_X2 U6774 ( .A1(n11960), .A2(dii_data_not_ready), .ZN(n11964) );
AND4_X2 U6775 ( .A1(n18844), .A2(n11957), .A3(n18014), .A4(n11970), .ZN(n11960) );
NAND4_X2 U6777 ( .A1(state[5]), .A2(n11973), .A3(n18627), .A4(n18601), .ZN(n11957) );
NAND2_X2 U6782 ( .A1(n11979), .A2(n11980), .ZN(n6282) );
OR2_X2 U6783 ( .A1(n18030), .A2(n17279), .ZN(n11980) );
NAND2_X2 U6784 ( .A1(aes_text_out[0]), .A2(n18022), .ZN(n11979) );
NAND2_X2 U6785 ( .A1(n11981), .A2(n11982), .ZN(n6281) );
OR2_X2 U6786 ( .A1(n18026), .A2(n17277), .ZN(n11982) );
NAND2_X2 U6787 ( .A1(aes_text_out[1]), .A2(n18022), .ZN(n11981) );
NAND2_X2 U6788 ( .A1(n11983), .A2(n11984), .ZN(n6280) );
OR2_X2 U6789 ( .A1(n18026), .A2(n17275), .ZN(n11984) );
NAND2_X2 U6790 ( .A1(aes_text_out[2]), .A2(n18023), .ZN(n11983) );
NAND2_X2 U6791 ( .A1(n11985), .A2(n11986), .ZN(n6279) );
OR2_X2 U6792 ( .A1(n18028), .A2(n17273), .ZN(n11986) );
NAND2_X2 U6793 ( .A1(aes_text_out[3]), .A2(n18023), .ZN(n11985) );
NAND2_X2 U6794 ( .A1(n11987), .A2(n11988), .ZN(n6278) );
OR2_X2 U6795 ( .A1(n18027), .A2(n17271), .ZN(n11988) );
NAND2_X2 U6796 ( .A1(aes_text_out[4]), .A2(n18023), .ZN(n11987) );
NAND2_X2 U6797 ( .A1(n11989), .A2(n11990), .ZN(n6277) );
OR2_X2 U6798 ( .A1(n18027), .A2(n17269), .ZN(n11990) );
NAND2_X2 U6799 ( .A1(aes_text_out[5]), .A2(n18024), .ZN(n11989) );
NAND2_X2 U6800 ( .A1(n11991), .A2(n11992), .ZN(n6276) );
OR2_X2 U6801 ( .A1(n18028), .A2(n17267), .ZN(n11992) );
NAND2_X2 U6802 ( .A1(aes_text_out[6]), .A2(n18024), .ZN(n11991) );
NAND2_X2 U6803 ( .A1(n11993), .A2(n11994), .ZN(n6275) );
OR2_X2 U6804 ( .A1(n18027), .A2(n17265), .ZN(n11994) );
NAND2_X2 U6805 ( .A1(aes_text_out[7]), .A2(n18023), .ZN(n11993) );
NAND2_X2 U6806 ( .A1(n11995), .A2(n11996), .ZN(n6274) );
OR2_X2 U6807 ( .A1(n18029), .A2(n17263), .ZN(n11996) );
NAND2_X2 U6808 ( .A1(aes_text_out[8]), .A2(n18025), .ZN(n11995) );
NAND2_X2 U6809 ( .A1(n11997), .A2(n11998), .ZN(n6273) );
OR2_X2 U6810 ( .A1(n18028), .A2(n17261), .ZN(n11998) );
NAND2_X2 U6811 ( .A1(aes_text_out[9]), .A2(n18025), .ZN(n11997) );
NAND2_X2 U6812 ( .A1(n11999), .A2(n12000), .ZN(n6272) );
OR2_X2 U6813 ( .A1(n18028), .A2(n17259), .ZN(n12000) );
NAND2_X2 U6814 ( .A1(aes_text_out[10]), .A2(n18023), .ZN(n11999) );
NAND2_X2 U6815 ( .A1(n12001), .A2(n12002), .ZN(n6271) );
OR2_X2 U6816 ( .A1(n18028), .A2(n17257), .ZN(n12002) );
NAND2_X2 U6817 ( .A1(aes_text_out[11]), .A2(n18025), .ZN(n12001) );
NAND2_X2 U6818 ( .A1(n12003), .A2(n12004), .ZN(n6270) );
OR2_X2 U6819 ( .A1(n18029), .A2(n17255), .ZN(n12004) );
NAND2_X2 U6820 ( .A1(aes_text_out[12]), .A2(n18025), .ZN(n12003) );
NAND2_X2 U6821 ( .A1(n12005), .A2(n12006), .ZN(n6269) );
OR2_X2 U6822 ( .A1(n18029), .A2(n17253), .ZN(n12006) );
NAND2_X2 U6823 ( .A1(aes_text_out[13]), .A2(n18023), .ZN(n12005) );
NAND2_X2 U6824 ( .A1(n12007), .A2(n12008), .ZN(n6268) );
OR2_X2 U6825 ( .A1(n18029), .A2(n17251), .ZN(n12008) );
NAND2_X2 U6826 ( .A1(aes_text_out[14]), .A2(n18026), .ZN(n12007) );
NAND2_X2 U6827 ( .A1(n12009), .A2(n12010), .ZN(n6267) );
OR2_X2 U6828 ( .A1(n18029), .A2(n17249), .ZN(n12010) );
NAND2_X2 U6829 ( .A1(aes_text_out[15]), .A2(n18026), .ZN(n12009) );
NAND2_X2 U6830 ( .A1(n12011), .A2(n12012), .ZN(n6266) );
OR2_X2 U6831 ( .A1(n18029), .A2(n17247), .ZN(n12012) );
NAND2_X2 U6832 ( .A1(aes_text_out[16]), .A2(n18024), .ZN(n12011) );
NAND2_X2 U6833 ( .A1(n12013), .A2(n12014), .ZN(n6265) );
OR2_X2 U6834 ( .A1(n18030), .A2(n17245), .ZN(n12014) );
NAND2_X2 U6835 ( .A1(aes_text_out[17]), .A2(n18026), .ZN(n12013) );
NAND2_X2 U6836 ( .A1(n12015), .A2(n12016), .ZN(n6264) );
OR2_X2 U6837 ( .A1(n18030), .A2(n17243), .ZN(n12016) );
NAND2_X2 U6838 ( .A1(aes_text_out[18]), .A2(n18026), .ZN(n12015) );
NAND2_X2 U6839 ( .A1(n12017), .A2(n12018), .ZN(n6263) );
OR2_X2 U6840 ( .A1(n18030), .A2(n17241), .ZN(n12018) );
NAND2_X2 U6841 ( .A1(aes_text_out[19]), .A2(n18026), .ZN(n12017) );
NAND2_X2 U6842 ( .A1(n12019), .A2(n12020), .ZN(n6262) );
OR2_X2 U6843 ( .A1(n18031), .A2(n17239), .ZN(n12020) );
NAND2_X2 U6844 ( .A1(aes_text_out[20]), .A2(n18024), .ZN(n12019) );
NAND2_X2 U6845 ( .A1(n12021), .A2(n12022), .ZN(n6261) );
OR2_X2 U6846 ( .A1(n18031), .A2(n17237), .ZN(n12022) );
NAND2_X2 U6847 ( .A1(aes_text_out[21]), .A2(n18026), .ZN(n12021) );
NAND2_X2 U6848 ( .A1(n12023), .A2(n12024), .ZN(n6260) );
OR2_X2 U6849 ( .A1(n18031), .A2(n17235), .ZN(n12024) );
NAND2_X2 U6850 ( .A1(aes_text_out[22]), .A2(n18026), .ZN(n12023) );
NAND2_X2 U6851 ( .A1(n12025), .A2(n12026), .ZN(n6259) );
OR2_X2 U6852 ( .A1(n18031), .A2(n17233), .ZN(n12026) );
NAND2_X2 U6853 ( .A1(aes_text_out[23]), .A2(n18025), .ZN(n12025) );
NAND2_X2 U6854 ( .A1(n12027), .A2(n12028), .ZN(n6258) );
OR2_X2 U6855 ( .A1(n18031), .A2(n17231), .ZN(n12028) );
NAND2_X2 U6856 ( .A1(aes_text_out[24]), .A2(n18025), .ZN(n12027) );
NAND2_X2 U6857 ( .A1(n12029), .A2(n12030), .ZN(n6257) );
OR2_X2 U6858 ( .A1(n18032), .A2(n17229), .ZN(n12030) );
NAND2_X2 U6859 ( .A1(aes_text_out[25]), .A2(n18025), .ZN(n12029) );
NAND2_X2 U6860 ( .A1(n12031), .A2(n12032), .ZN(n6256) );
OR2_X2 U6861 ( .A1(n18032), .A2(n17227), .ZN(n12032) );
NAND2_X2 U6862 ( .A1(aes_text_out[26]), .A2(n18025), .ZN(n12031) );
NAND2_X2 U6863 ( .A1(n12033), .A2(n12034), .ZN(n6255) );
OR2_X2 U6864 ( .A1(n18032), .A2(n17225), .ZN(n12034) );
NAND2_X2 U6865 ( .A1(aes_text_out[27]), .A2(n18025), .ZN(n12033) );
NAND2_X2 U6866 ( .A1(n12035), .A2(n12036), .ZN(n6254) );
OR2_X2 U6867 ( .A1(n18032), .A2(n17223), .ZN(n12036) );
NAND2_X2 U6868 ( .A1(aes_text_out[28]), .A2(n18025), .ZN(n12035) );
NAND2_X2 U6869 ( .A1(n12037), .A2(n12038), .ZN(n6253) );
OR2_X2 U6870 ( .A1(n18032), .A2(n17221), .ZN(n12038) );
NAND2_X2 U6871 ( .A1(aes_text_out[29]), .A2(n18023), .ZN(n12037) );
NAND2_X2 U6872 ( .A1(n12039), .A2(n12040), .ZN(n6252) );
OR2_X2 U6873 ( .A1(n18033), .A2(n17219), .ZN(n12040) );
NAND2_X2 U6874 ( .A1(aes_text_out[30]), .A2(n18025), .ZN(n12039) );
NAND2_X2 U6875 ( .A1(n12041), .A2(n12042), .ZN(n6251) );
OR2_X2 U6876 ( .A1(n18033), .A2(n17217), .ZN(n12042) );
NAND2_X2 U6877 ( .A1(aes_text_out[31]), .A2(n18024), .ZN(n12041) );
NAND2_X2 U6878 ( .A1(n12043), .A2(n12044), .ZN(n6250) );
OR2_X2 U6879 ( .A1(n18033), .A2(n17215), .ZN(n12044) );
NAND2_X2 U6880 ( .A1(aes_text_out[32]), .A2(n18024), .ZN(n12043) );
NAND2_X2 U6881 ( .A1(n12045), .A2(n12046), .ZN(n6249) );
OR2_X2 U6882 ( .A1(n18033), .A2(n17213), .ZN(n12046) );
NAND2_X2 U6883 ( .A1(aes_text_out[33]), .A2(n18024), .ZN(n12045) );
NAND2_X2 U6884 ( .A1(n12047), .A2(n12048), .ZN(n6248) );
OR2_X2 U6885 ( .A1(n18034), .A2(n17211), .ZN(n12048) );
NAND2_X2 U6886 ( .A1(aes_text_out[34]), .A2(n18024), .ZN(n12047) );
NAND2_X2 U6887 ( .A1(n12049), .A2(n12050), .ZN(n6247) );
OR2_X2 U6888 ( .A1(n18034), .A2(n17209), .ZN(n12050) );
NAND2_X2 U6889 ( .A1(aes_text_out[35]), .A2(n18024), .ZN(n12049) );
NAND2_X2 U6890 ( .A1(n12051), .A2(n12052), .ZN(n6246) );
OR2_X2 U6891 ( .A1(n18034), .A2(n17207), .ZN(n12052) );
NAND2_X2 U6892 ( .A1(aes_text_out[36]), .A2(n18024), .ZN(n12051) );
NAND2_X2 U6893 ( .A1(n12053), .A2(n12054), .ZN(n6245) );
OR2_X2 U6894 ( .A1(n18034), .A2(n17205), .ZN(n12054) );
NAND2_X2 U6895 ( .A1(aes_text_out[37]), .A2(n18024), .ZN(n12053) );
NAND2_X2 U6896 ( .A1(n12055), .A2(n12056), .ZN(n6244) );
OR2_X2 U6897 ( .A1(n18034), .A2(n17203), .ZN(n12056) );
NAND2_X2 U6898 ( .A1(aes_text_out[38]), .A2(n18023), .ZN(n12055) );
NAND2_X2 U6899 ( .A1(n12057), .A2(n12058), .ZN(n6243) );
OR2_X2 U6900 ( .A1(n18035), .A2(n17201), .ZN(n12058) );
NAND2_X2 U6901 ( .A1(aes_text_out[39]), .A2(n18023), .ZN(n12057) );
NAND2_X2 U6902 ( .A1(n12059), .A2(n12060), .ZN(n6242) );
OR2_X2 U6903 ( .A1(n18035), .A2(n17199), .ZN(n12060) );
NAND2_X2 U6904 ( .A1(aes_text_out[40]), .A2(n18023), .ZN(n12059) );
NAND2_X2 U6905 ( .A1(n12061), .A2(n12062), .ZN(n6241) );
OR2_X2 U6906 ( .A1(n18035), .A2(n17197), .ZN(n12062) );
NAND2_X2 U6907 ( .A1(aes_text_out[41]), .A2(n18023), .ZN(n12061) );
NAND2_X2 U6908 ( .A1(n12063), .A2(n12064), .ZN(n6240) );
OR2_X2 U6909 ( .A1(n18035), .A2(n17195), .ZN(n12064) );
NAND2_X2 U6910 ( .A1(aes_text_out[42]), .A2(n18022), .ZN(n12063) );
NAND2_X2 U6911 ( .A1(n12065), .A2(n12066), .ZN(n6239) );
OR2_X2 U6912 ( .A1(n18027), .A2(n17193), .ZN(n12066) );
NAND2_X2 U6913 ( .A1(aes_text_out[43]), .A2(n18022), .ZN(n12065) );
NAND2_X2 U6914 ( .A1(n12067), .A2(n12068), .ZN(n6238) );
OR2_X2 U6915 ( .A1(n18035), .A2(n17191), .ZN(n12068) );
NAND2_X2 U6916 ( .A1(aes_text_out[44]), .A2(n18022), .ZN(n12067) );
NAND2_X2 U6917 ( .A1(n12069), .A2(n12070), .ZN(n6237) );
OR2_X2 U6918 ( .A1(n18035), .A2(n17189), .ZN(n12070) );
NAND2_X2 U6919 ( .A1(aes_text_out[45]), .A2(n18022), .ZN(n12069) );
NAND2_X2 U6920 ( .A1(n12071), .A2(n12072), .ZN(n6236) );
OR2_X2 U6921 ( .A1(n18035), .A2(n17187), .ZN(n12072) );
NAND2_X2 U6922 ( .A1(aes_text_out[46]), .A2(n18022), .ZN(n12071) );
NAND2_X2 U6923 ( .A1(n12073), .A2(n12074), .ZN(n6235) );
OR2_X2 U6924 ( .A1(n18035), .A2(n17185), .ZN(n12074) );
NAND2_X2 U6925 ( .A1(aes_text_out[47]), .A2(n18022), .ZN(n12073) );
NAND2_X2 U6926 ( .A1(n12075), .A2(n12076), .ZN(n6234) );
OR2_X2 U6927 ( .A1(n18035), .A2(n17183), .ZN(n12076) );
NAND2_X2 U6928 ( .A1(aes_text_out[48]), .A2(n18022), .ZN(n12075) );
NAND2_X2 U6929 ( .A1(n12077), .A2(n12078), .ZN(n6233) );
OR2_X2 U6930 ( .A1(n18035), .A2(n17181), .ZN(n12078) );
NAND2_X2 U6931 ( .A1(aes_text_out[49]), .A2(n18022), .ZN(n12077) );
NAND2_X2 U6932 ( .A1(n12079), .A2(n12080), .ZN(n6232) );
OR2_X2 U6933 ( .A1(n18035), .A2(n17179), .ZN(n12080) );
NAND2_X2 U6934 ( .A1(aes_text_out[50]), .A2(n18021), .ZN(n12079) );
NAND2_X2 U6935 ( .A1(n12081), .A2(n12082), .ZN(n6231) );
OR2_X2 U6936 ( .A1(n18034), .A2(n17177), .ZN(n12082) );
NAND2_X2 U6937 ( .A1(aes_text_out[51]), .A2(n18021), .ZN(n12081) );
NAND2_X2 U6938 ( .A1(n12083), .A2(n12084), .ZN(n6230) );
OR2_X2 U6939 ( .A1(n18034), .A2(n17175), .ZN(n12084) );
NAND2_X2 U6940 ( .A1(aes_text_out[52]), .A2(n18021), .ZN(n12083) );
NAND2_X2 U6941 ( .A1(n12085), .A2(n12086), .ZN(n6229) );
OR2_X2 U6942 ( .A1(n18034), .A2(n17173), .ZN(n12086) );
NAND2_X2 U6943 ( .A1(aes_text_out[53]), .A2(n18021), .ZN(n12085) );
NAND2_X2 U6944 ( .A1(n12087), .A2(n12088), .ZN(n6228) );
OR2_X2 U6945 ( .A1(n18034), .A2(n17171), .ZN(n12088) );
NAND2_X2 U6946 ( .A1(aes_text_out[54]), .A2(n18021), .ZN(n12087) );
NAND2_X2 U6947 ( .A1(n12089), .A2(n12090), .ZN(n6227) );
OR2_X2 U6948 ( .A1(n18034), .A2(n17169), .ZN(n12090) );
NAND2_X2 U6949 ( .A1(aes_text_out[55]), .A2(n18021), .ZN(n12089) );
NAND2_X2 U6950 ( .A1(n12091), .A2(n12092), .ZN(n6226) );
OR2_X2 U6951 ( .A1(n18034), .A2(n17167), .ZN(n12092) );
NAND2_X2 U6952 ( .A1(aes_text_out[56]), .A2(n18021), .ZN(n12091) );
NAND2_X2 U6953 ( .A1(n12093), .A2(n12094), .ZN(n6225) );
OR2_X2 U6954 ( .A1(n18034), .A2(n17165), .ZN(n12094) );
NAND2_X2 U6955 ( .A1(aes_text_out[57]), .A2(n18021), .ZN(n12093) );
NAND2_X2 U6956 ( .A1(n12095), .A2(n12096), .ZN(n6224) );
OR2_X2 U6957 ( .A1(n18034), .A2(n17163), .ZN(n12096) );
NAND2_X2 U6958 ( .A1(aes_text_out[58]), .A2(n18021), .ZN(n12095) );
NAND2_X2 U6959 ( .A1(n12097), .A2(n12098), .ZN(n6223) );
OR2_X2 U6960 ( .A1(n18034), .A2(n17161), .ZN(n12098) );
NAND2_X2 U6961 ( .A1(aes_text_out[59]), .A2(n18021), .ZN(n12097) );
NAND2_X2 U6962 ( .A1(n12099), .A2(n12100), .ZN(n6222) );
OR2_X2 U6963 ( .A1(n18033), .A2(n17159), .ZN(n12100) );
NAND2_X2 U6964 ( .A1(aes_text_out[60]), .A2(n18021), .ZN(n12099) );
NAND2_X2 U6965 ( .A1(n12101), .A2(n12102), .ZN(n6221) );
OR2_X2 U6966 ( .A1(n18033), .A2(n17157), .ZN(n12102) );
NAND2_X2 U6967 ( .A1(aes_text_out[61]), .A2(n18020), .ZN(n12101) );
NAND2_X2 U6968 ( .A1(n12103), .A2(n12104), .ZN(n6220) );
OR2_X2 U6969 ( .A1(n18033), .A2(n17155), .ZN(n12104) );
NAND2_X2 U6970 ( .A1(aes_text_out[62]), .A2(n18020), .ZN(n12103) );
NAND2_X2 U6971 ( .A1(n12105), .A2(n12106), .ZN(n6219) );
OR2_X2 U6972 ( .A1(n18033), .A2(n17153), .ZN(n12106) );
NAND2_X2 U6973 ( .A1(aes_text_out[63]), .A2(n18022), .ZN(n12105) );
NAND2_X2 U6974 ( .A1(n12107), .A2(n12108), .ZN(n6218) );
OR2_X2 U6975 ( .A1(n18033), .A2(n17151), .ZN(n12108) );
NAND2_X2 U6976 ( .A1(aes_text_out[64]), .A2(n18020), .ZN(n12107) );
NAND2_X2 U6977 ( .A1(n12109), .A2(n12110), .ZN(n6217) );
OR2_X2 U6978 ( .A1(n18033), .A2(n17149), .ZN(n12110) );
NAND2_X2 U6979 ( .A1(aes_text_out[65]), .A2(n18020), .ZN(n12109) );
NAND2_X2 U6980 ( .A1(n12111), .A2(n12112), .ZN(n6216) );
OR2_X2 U6981 ( .A1(n18033), .A2(n17147), .ZN(n12112) );
NAND2_X2 U6982 ( .A1(aes_text_out[66]), .A2(n18020), .ZN(n12111) );
NAND2_X2 U6983 ( .A1(n12113), .A2(n12114), .ZN(n6215) );
OR2_X2 U6984 ( .A1(n18033), .A2(n17145), .ZN(n12114) );
NAND2_X2 U6985 ( .A1(aes_text_out[67]), .A2(n18020), .ZN(n12113) );
NAND2_X2 U6986 ( .A1(n12115), .A2(n12116), .ZN(n6214) );
OR2_X2 U6987 ( .A1(n18033), .A2(n17143), .ZN(n12116) );
NAND2_X2 U6988 ( .A1(aes_text_out[68]), .A2(n18020), .ZN(n12115) );
NAND2_X2 U6989 ( .A1(n12117), .A2(n12118), .ZN(n6213) );
OR2_X2 U6990 ( .A1(n18033), .A2(n17141), .ZN(n12118) );
NAND2_X2 U6991 ( .A1(aes_text_out[69]), .A2(n18020), .ZN(n12117) );
NAND2_X2 U6992 ( .A1(n12119), .A2(n12120), .ZN(n6212) );
OR2_X2 U6993 ( .A1(n18032), .A2(n17139), .ZN(n12120) );
NAND2_X2 U6994 ( .A1(aes_text_out[70]), .A2(n18020), .ZN(n12119) );
NAND2_X2 U6995 ( .A1(n12121), .A2(n12122), .ZN(n6211) );
OR2_X2 U6996 ( .A1(n18032), .A2(n17137), .ZN(n12122) );
NAND2_X2 U6997 ( .A1(aes_text_out[71]), .A2(n18020), .ZN(n12121) );
NAND2_X2 U6998 ( .A1(n12123), .A2(n12124), .ZN(n6210) );
OR2_X2 U6999 ( .A1(n18032), .A2(n17135), .ZN(n12124) );
NAND2_X2 U7000 ( .A1(aes_text_out[72]), .A2(n18019), .ZN(n12123) );
NAND2_X2 U7001 ( .A1(n12125), .A2(n12126), .ZN(n6209) );
OR2_X2 U7002 ( .A1(n18032), .A2(n17133), .ZN(n12126) );
NAND2_X2 U7003 ( .A1(aes_text_out[73]), .A2(n18019), .ZN(n12125) );
NAND2_X2 U7004 ( .A1(n12127), .A2(n12128), .ZN(n6208) );
OR2_X2 U7005 ( .A1(n18032), .A2(n17131), .ZN(n12128) );
NAND2_X2 U7006 ( .A1(aes_text_out[74]), .A2(n18019), .ZN(n12127) );
NAND2_X2 U7007 ( .A1(n12129), .A2(n12130), .ZN(n6207) );
OR2_X2 U7008 ( .A1(n18032), .A2(n17129), .ZN(n12130) );
NAND2_X2 U7009 ( .A1(aes_text_out[75]), .A2(n18019), .ZN(n12129) );
NAND2_X2 U7010 ( .A1(n12131), .A2(n12132), .ZN(n6206) );
OR2_X2 U7011 ( .A1(n18032), .A2(n17127), .ZN(n12132) );
NAND2_X2 U7012 ( .A1(aes_text_out[76]), .A2(n18019), .ZN(n12131) );
NAND2_X2 U7013 ( .A1(n12133), .A2(n12134), .ZN(n6205) );
OR2_X2 U7014 ( .A1(n18032), .A2(n17125), .ZN(n12134) );
NAND2_X2 U7015 ( .A1(aes_text_out[77]), .A2(n18019), .ZN(n12133) );
NAND2_X2 U7016 ( .A1(n12135), .A2(n12136), .ZN(n6204) );
OR2_X2 U7017 ( .A1(n18032), .A2(n17123), .ZN(n12136) );
NAND2_X2 U7018 ( .A1(aes_text_out[78]), .A2(n18019), .ZN(n12135) );
NAND2_X2 U7019 ( .A1(n12137), .A2(n12138), .ZN(n6203) );
OR2_X2 U7020 ( .A1(n18031), .A2(n17121), .ZN(n12138) );
NAND2_X2 U7021 ( .A1(aes_text_out[79]), .A2(n18019), .ZN(n12137) );
NAND2_X2 U7022 ( .A1(n12139), .A2(n12140), .ZN(n6202) );
OR2_X2 U7023 ( .A1(n18031), .A2(n17119), .ZN(n12140) );
NAND2_X2 U7024 ( .A1(aes_text_out[80]), .A2(n18019), .ZN(n12139) );
NAND2_X2 U7025 ( .A1(n12141), .A2(n12142), .ZN(n6201) );
OR2_X2 U7026 ( .A1(n18031), .A2(n17117), .ZN(n12142) );
NAND2_X2 U7027 ( .A1(aes_text_out[81]), .A2(n18019), .ZN(n12141) );
NAND2_X2 U7028 ( .A1(n12143), .A2(n12144), .ZN(n6200) );
OR2_X2 U7029 ( .A1(n18031), .A2(n17115), .ZN(n12144) );
NAND2_X2 U7030 ( .A1(aes_text_out[82]), .A2(n18019), .ZN(n12143) );
NAND2_X2 U7031 ( .A1(n12145), .A2(n12146), .ZN(n6199) );
OR2_X2 U7032 ( .A1(n18031), .A2(n17113), .ZN(n12146) );
NAND2_X2 U7033 ( .A1(aes_text_out[83]), .A2(n18018), .ZN(n12145) );
NAND2_X2 U7034 ( .A1(n12147), .A2(n12148), .ZN(n6198) );
OR2_X2 U7035 ( .A1(n18031), .A2(n17111), .ZN(n12148) );
NAND2_X2 U7036 ( .A1(aes_text_out[84]), .A2(n18018), .ZN(n12147) );
NAND2_X2 U7037 ( .A1(n12149), .A2(n12150), .ZN(n6197) );
OR2_X2 U7038 ( .A1(n18031), .A2(n17109), .ZN(n12150) );
NAND2_X2 U7039 ( .A1(aes_text_out[85]), .A2(n18018), .ZN(n12149) );
NAND2_X2 U7040 ( .A1(n12151), .A2(n12152), .ZN(n6196) );
OR2_X2 U7041 ( .A1(n18031), .A2(n17107), .ZN(n12152) );
NAND2_X2 U7042 ( .A1(aes_text_out[86]), .A2(n18018), .ZN(n12151) );
NAND2_X2 U7043 ( .A1(n12153), .A2(n12154), .ZN(n6195) );
OR2_X2 U7044 ( .A1(n18031), .A2(n17105), .ZN(n12154) );
NAND2_X2 U7045 ( .A1(aes_text_out[87]), .A2(n18018), .ZN(n12153) );
NAND2_X2 U7046 ( .A1(n12155), .A2(n12156), .ZN(n6194) );
OR2_X2 U7047 ( .A1(n18030), .A2(n17103), .ZN(n12156) );
NAND2_X2 U7048 ( .A1(aes_text_out[88]), .A2(n18018), .ZN(n12155) );
NAND2_X2 U7049 ( .A1(n12157), .A2(n12158), .ZN(n6193) );
OR2_X2 U7050 ( .A1(n18030), .A2(n17101), .ZN(n12158) );
NAND2_X2 U7051 ( .A1(aes_text_out[89]), .A2(n18018), .ZN(n12157) );
NAND2_X2 U7052 ( .A1(n12159), .A2(n12160), .ZN(n6192) );
OR2_X2 U7053 ( .A1(n18030), .A2(n17099), .ZN(n12160) );
NAND2_X2 U7054 ( .A1(aes_text_out[90]), .A2(n18018), .ZN(n12159) );
NAND2_X2 U7055 ( .A1(n12161), .A2(n12162), .ZN(n6191) );
OR2_X2 U7056 ( .A1(n18030), .A2(n17097), .ZN(n12162) );
NAND2_X2 U7057 ( .A1(aes_text_out[91]), .A2(n18018), .ZN(n12161) );
NAND2_X2 U7058 ( .A1(n12163), .A2(n12164), .ZN(n6190) );
OR2_X2 U7059 ( .A1(n18030), .A2(n17095), .ZN(n12164) );
NAND2_X2 U7060 ( .A1(aes_text_out[92]), .A2(n18018), .ZN(n12163) );
NAND2_X2 U7061 ( .A1(n12165), .A2(n12166), .ZN(n6189) );
OR2_X2 U7062 ( .A1(n18030), .A2(n17093), .ZN(n12166) );
NAND2_X2 U7063 ( .A1(aes_text_out[93]), .A2(n18018), .ZN(n12165) );
NAND2_X2 U7064 ( .A1(n12167), .A2(n12168), .ZN(n6188) );
OR2_X2 U7065 ( .A1(n18030), .A2(n17091), .ZN(n12168) );
NAND2_X2 U7066 ( .A1(aes_text_out[94]), .A2(n18017), .ZN(n12167) );
NAND2_X2 U7067 ( .A1(n12169), .A2(n12170), .ZN(n6187) );
OR2_X2 U7068 ( .A1(n18030), .A2(n17089), .ZN(n12170) );
NAND2_X2 U7069 ( .A1(aes_text_out[95]), .A2(n18017), .ZN(n12169) );
NAND2_X2 U7070 ( .A1(n12171), .A2(n12172), .ZN(n6186) );
OR2_X2 U7071 ( .A1(n18030), .A2(n17087), .ZN(n12172) );
NAND2_X2 U7072 ( .A1(aes_text_out[96]), .A2(n18017), .ZN(n12171) );
NAND2_X2 U7073 ( .A1(n12173), .A2(n12174), .ZN(n6185) );
OR2_X2 U7074 ( .A1(n18029), .A2(n17085), .ZN(n12174) );
NAND2_X2 U7075 ( .A1(aes_text_out[97]), .A2(n18017), .ZN(n12173) );
NAND2_X2 U7076 ( .A1(n12175), .A2(n12176), .ZN(n6184) );
OR2_X2 U7077 ( .A1(n18030), .A2(n17083), .ZN(n12176) );
NAND2_X2 U7078 ( .A1(aes_text_out[98]), .A2(n18017), .ZN(n12175) );
NAND2_X2 U7079 ( .A1(n12177), .A2(n12178), .ZN(n6183) );
OR2_X2 U7080 ( .A1(n18029), .A2(n17081), .ZN(n12178) );
NAND2_X2 U7081 ( .A1(aes_text_out[99]), .A2(n18017), .ZN(n12177) );
NAND2_X2 U7082 ( .A1(n12179), .A2(n12180), .ZN(n6182) );
OR2_X2 U7083 ( .A1(n18029), .A2(n17079), .ZN(n12180) );
NAND2_X2 U7084 ( .A1(aes_text_out[100]), .A2(n18017), .ZN(n12179) );
NAND2_X2 U7085 ( .A1(n12181), .A2(n12182), .ZN(n6181) );
OR2_X2 U7086 ( .A1(n18029), .A2(n17077), .ZN(n12182) );
NAND2_X2 U7087 ( .A1(aes_text_out[101]), .A2(n18017), .ZN(n12181) );
NAND2_X2 U7088 ( .A1(n12183), .A2(n12184), .ZN(n6180) );
OR2_X2 U7089 ( .A1(n18029), .A2(n17075), .ZN(n12184) );
NAND2_X2 U7090 ( .A1(aes_text_out[102]), .A2(n18017), .ZN(n12183) );
NAND2_X2 U7091 ( .A1(n12185), .A2(n12186), .ZN(n6179) );
OR2_X2 U7092 ( .A1(n18029), .A2(n17073), .ZN(n12186) );
NAND2_X2 U7093 ( .A1(aes_text_out[103]), .A2(n18017), .ZN(n12185) );
NAND2_X2 U7094 ( .A1(n12187), .A2(n12188), .ZN(n6178) );
OR2_X2 U7095 ( .A1(n18028), .A2(n17071), .ZN(n12188) );
NAND2_X2 U7096 ( .A1(aes_text_out[104]), .A2(n18017), .ZN(n12187) );
NAND2_X2 U7097 ( .A1(n12189), .A2(n12190), .ZN(n6177) );
OR2_X2 U7098 ( .A1(n18029), .A2(n17069), .ZN(n12190) );
NAND2_X2 U7099 ( .A1(aes_text_out[105]), .A2(n18016), .ZN(n12189) );
NAND2_X2 U7100 ( .A1(n12191), .A2(n12192), .ZN(n6176) );
OR2_X2 U7101 ( .A1(n18028), .A2(n17067), .ZN(n12192) );
NAND2_X2 U7102 ( .A1(aes_text_out[106]), .A2(n18016), .ZN(n12191) );
NAND2_X2 U7103 ( .A1(n12193), .A2(n12194), .ZN(n6175) );
OR2_X2 U7104 ( .A1(n18028), .A2(n17065), .ZN(n12194) );
NAND2_X2 U7105 ( .A1(aes_text_out[107]), .A2(n18016), .ZN(n12193) );
NAND2_X2 U7106 ( .A1(n12195), .A2(n12196), .ZN(n6174) );
OR2_X2 U7107 ( .A1(n18028), .A2(n17063), .ZN(n12196) );
NAND2_X2 U7108 ( .A1(aes_text_out[108]), .A2(n18016), .ZN(n12195) );
NAND2_X2 U7109 ( .A1(n12197), .A2(n12198), .ZN(n6173) );
OR2_X2 U7110 ( .A1(n18028), .A2(n17061), .ZN(n12198) );
NAND2_X2 U7111 ( .A1(aes_text_out[109]), .A2(n18016), .ZN(n12197) );
NAND2_X2 U7112 ( .A1(n12199), .A2(n12200), .ZN(n6172) );
OR2_X2 U7113 ( .A1(n18028), .A2(n17059), .ZN(n12200) );
NAND2_X2 U7114 ( .A1(aes_text_out[110]), .A2(n18016), .ZN(n12199) );
NAND2_X2 U7115 ( .A1(n12201), .A2(n12202), .ZN(n6171) );
OR2_X2 U7116 ( .A1(n18028), .A2(n17057), .ZN(n12202) );
NAND2_X2 U7117 ( .A1(aes_text_out[111]), .A2(n18016), .ZN(n12201) );
NAND2_X2 U7118 ( .A1(n12203), .A2(n12204), .ZN(n6170) );
OR2_X2 U7119 ( .A1(n18027), .A2(n17055), .ZN(n12204) );
NAND2_X2 U7120 ( .A1(aes_text_out[112]), .A2(n18016), .ZN(n12203) );
NAND2_X2 U7121 ( .A1(n12205), .A2(n12206), .ZN(n6169) );
OR2_X2 U7122 ( .A1(n18027), .A2(n17053), .ZN(n12206) );
NAND2_X2 U7123 ( .A1(aes_text_out[113]), .A2(n18016), .ZN(n12205) );
NAND2_X2 U7124 ( .A1(n12207), .A2(n12208), .ZN(n6168) );
OR2_X2 U7125 ( .A1(n18029), .A2(n17051), .ZN(n12208) );
NAND2_X2 U7126 ( .A1(aes_text_out[114]), .A2(n18016), .ZN(n12207) );
NAND2_X2 U7127 ( .A1(n12209), .A2(n12210), .ZN(n6167) );
OR2_X2 U7128 ( .A1(n18028), .A2(n17049), .ZN(n12210) );
NAND2_X2 U7129 ( .A1(aes_text_out[115]), .A2(n18016), .ZN(n12209) );
NAND2_X2 U7130 ( .A1(n12211), .A2(n12212), .ZN(n6166) );
OR2_X2 U7131 ( .A1(n18027), .A2(n17047), .ZN(n12212) );
NAND2_X2 U7132 ( .A1(aes_text_out[116]), .A2(n18015), .ZN(n12211) );
NAND2_X2 U7133 ( .A1(n12213), .A2(n12214), .ZN(n6165) );
OR2_X2 U7134 ( .A1(n18027), .A2(n17045), .ZN(n12214) );
NAND2_X2 U7135 ( .A1(aes_text_out[117]), .A2(n18015), .ZN(n12213) );
NAND2_X2 U7136 ( .A1(n12215), .A2(n12216), .ZN(n6164) );
OR2_X2 U7137 ( .A1(n18027), .A2(n17043), .ZN(n12216) );
NAND2_X2 U7138 ( .A1(aes_text_out[118]), .A2(n18015), .ZN(n12215) );
NAND2_X2 U7139 ( .A1(n12217), .A2(n12218), .ZN(n6163) );
OR2_X2 U7140 ( .A1(n18027), .A2(n17041), .ZN(n12218) );
NAND2_X2 U7141 ( .A1(aes_text_out[119]), .A2(n18015), .ZN(n12217) );
NAND2_X2 U7142 ( .A1(n12219), .A2(n12220), .ZN(n6162) );
OR2_X2 U7143 ( .A1(n18027), .A2(n17039), .ZN(n12220) );
NAND2_X2 U7144 ( .A1(aes_text_out[120]), .A2(n18015), .ZN(n12219) );
NAND2_X2 U7145 ( .A1(n12221), .A2(n12222), .ZN(n6161) );
OR2_X2 U7146 ( .A1(n18027), .A2(n17037), .ZN(n12222) );
NAND2_X2 U7147 ( .A1(aes_text_out[121]), .A2(n18015), .ZN(n12221) );
NAND2_X2 U7148 ( .A1(n12223), .A2(n12224), .ZN(n6160) );
OR2_X2 U7149 ( .A1(n18026), .A2(n17035), .ZN(n12224) );
NAND2_X2 U7150 ( .A1(aes_text_out[122]), .A2(n18015), .ZN(n12223) );
NAND2_X2 U7151 ( .A1(n12225), .A2(n12226), .ZN(n6159) );
OR2_X2 U7152 ( .A1(n18027), .A2(n17033), .ZN(n12226) );
NAND2_X2 U7153 ( .A1(aes_text_out[123]), .A2(n18015), .ZN(n12225) );
NAND2_X2 U7154 ( .A1(n12227), .A2(n12228), .ZN(n6158) );
OR2_X2 U7155 ( .A1(n18026), .A2(n17031), .ZN(n12228) );
NAND2_X2 U7156 ( .A1(aes_text_out[124]), .A2(n18015), .ZN(n12227) );
NAND2_X2 U7157 ( .A1(n12229), .A2(n12230), .ZN(n6157) );
OR2_X2 U7158 ( .A1(n18028), .A2(n17029), .ZN(n12230) );
NAND2_X2 U7159 ( .A1(aes_text_out[125]), .A2(n18015), .ZN(n12229) );
NAND2_X2 U7160 ( .A1(n12231), .A2(n12232), .ZN(n6156) );
OR2_X2 U7161 ( .A1(n18027), .A2(n17027), .ZN(n12232) );
NAND2_X2 U7162 ( .A1(aes_text_out[126]), .A2(n18015), .ZN(n12231) );
NAND2_X2 U7163 ( .A1(n12233), .A2(n12234), .ZN(n6155) );
OR2_X2 U7164 ( .A1(n18026), .A2(n17025), .ZN(n12234) );
NAND2_X2 U7165 ( .A1(aes_text_out[127]), .A2(n18020), .ZN(n12233) );
NAND2_X2 U7168 ( .A1(n12236), .A2(n12237), .ZN(n6154) );
NAND2_X2 U7169 ( .A1(aes_text_out[0]), .A2(n17989), .ZN(n12237) );
NAND2_X2 U7170 ( .A1(n17988), .A2(n18891), .ZN(n12236) );
NAND2_X2 U7171 ( .A1(n12239), .A2(n12240), .ZN(n6153) );
NAND2_X2 U7172 ( .A1(aes_text_out[1]), .A2(n17989), .ZN(n12240) );
NAND2_X2 U7173 ( .A1(n17988), .A2(n18890), .ZN(n12239) );
NAND2_X2 U7174 ( .A1(n12241), .A2(n12242), .ZN(n6152) );
NAND2_X2 U7175 ( .A1(aes_text_out[2]), .A2(n17989), .ZN(n12242) );
NAND2_X2 U7176 ( .A1(n17988), .A2(n18889), .ZN(n12241) );
NAND2_X2 U7177 ( .A1(n12243), .A2(n12244), .ZN(n6151) );
NAND2_X2 U7178 ( .A1(aes_text_out[3]), .A2(n17995), .ZN(n12244) );
NAND2_X2 U7179 ( .A1(n17988), .A2(n18888), .ZN(n12243) );
NAND2_X2 U7180 ( .A1(n12245), .A2(n12246), .ZN(n6150) );
NAND2_X2 U7181 ( .A1(aes_text_out[4]), .A2(n17995), .ZN(n12246) );
NAND2_X2 U7182 ( .A1(n17988), .A2(n18887), .ZN(n12245) );
NAND2_X2 U7183 ( .A1(n12247), .A2(n12248), .ZN(n6149) );
NAND2_X2 U7184 ( .A1(aes_text_out[5]), .A2(n17995), .ZN(n12248) );
NAND2_X2 U7185 ( .A1(n17988), .A2(n18886), .ZN(n12247) );
NAND2_X2 U7186 ( .A1(n12249), .A2(n12250), .ZN(n6148) );
NAND2_X2 U7187 ( .A1(aes_text_out[6]), .A2(n17995), .ZN(n12250) );
NAND2_X2 U7188 ( .A1(n17988), .A2(n18885), .ZN(n12249) );
NAND2_X2 U7189 ( .A1(n12251), .A2(n12252), .ZN(n6147) );
NAND2_X2 U7190 ( .A1(aes_text_out[7]), .A2(n17995), .ZN(n12252) );
NAND2_X2 U7191 ( .A1(n17987), .A2(n18884), .ZN(n12251) );
NAND2_X2 U7192 ( .A1(n12253), .A2(n12254), .ZN(n6146) );
NAND2_X2 U7193 ( .A1(aes_text_out[8]), .A2(n17995), .ZN(n12254) );
NAND2_X2 U7194 ( .A1(n17987), .A2(n18883), .ZN(n12253) );
NAND2_X2 U7195 ( .A1(n12255), .A2(n12256), .ZN(n6145) );
NAND2_X2 U7196 ( .A1(aes_text_out[9]), .A2(n17995), .ZN(n12256) );
NAND2_X2 U7197 ( .A1(n17987), .A2(n18882), .ZN(n12255) );
NAND2_X2 U7198 ( .A1(n12257), .A2(n12258), .ZN(n6144) );
NAND2_X2 U7199 ( .A1(aes_text_out[10]), .A2(n17995), .ZN(n12258) );
NAND2_X2 U7200 ( .A1(n17987), .A2(n18881), .ZN(n12257) );
NAND2_X2 U7201 ( .A1(n12259), .A2(n12260), .ZN(n6143) );
NAND2_X2 U7202 ( .A1(aes_text_out[11]), .A2(n17995), .ZN(n12260) );
NAND2_X2 U7203 ( .A1(n17987), .A2(n18880), .ZN(n12259) );
NAND2_X2 U7204 ( .A1(n12261), .A2(n12262), .ZN(n6142) );
NAND2_X2 U7205 ( .A1(aes_text_out[12]), .A2(n17995), .ZN(n12262) );
NAND2_X2 U7206 ( .A1(n17987), .A2(n18879), .ZN(n12261) );
NAND2_X2 U7207 ( .A1(n12263), .A2(n12264), .ZN(n6141) );
NAND2_X2 U7208 ( .A1(aes_text_out[13]), .A2(n17995), .ZN(n12264) );
NAND2_X2 U7209 ( .A1(n17987), .A2(n18878), .ZN(n12263) );
NAND2_X2 U7210 ( .A1(n12265), .A2(n12266), .ZN(n6140) );
NAND2_X2 U7211 ( .A1(aes_text_out[14]), .A2(n17995), .ZN(n12266) );
NAND2_X2 U7212 ( .A1(n17987), .A2(n18877), .ZN(n12265) );
NAND2_X2 U7213 ( .A1(n12267), .A2(n12268), .ZN(n6139) );
NAND2_X2 U7214 ( .A1(aes_text_out[15]), .A2(n17995), .ZN(n12268) );
NAND2_X2 U7215 ( .A1(n17987), .A2(n18876), .ZN(n12267) );
NAND2_X2 U7216 ( .A1(n12269), .A2(n12270), .ZN(n6138) );
NAND2_X2 U7217 ( .A1(aes_text_out[16]), .A2(n17995), .ZN(n12270) );
NAND2_X2 U7218 ( .A1(n17987), .A2(n18875), .ZN(n12269) );
NAND2_X2 U7219 ( .A1(n12271), .A2(n12272), .ZN(n6137) );
NAND2_X2 U7220 ( .A1(aes_text_out[17]), .A2(n17995), .ZN(n12272) );
NAND2_X2 U7221 ( .A1(n17987), .A2(n18874), .ZN(n12271) );
NAND2_X2 U7222 ( .A1(n12273), .A2(n12274), .ZN(n6136) );
NAND2_X2 U7223 ( .A1(aes_text_out[18]), .A2(n17995), .ZN(n12274) );
NAND2_X2 U7224 ( .A1(n17986), .A2(n18873), .ZN(n12273) );
NAND2_X2 U7225 ( .A1(n12275), .A2(n12276), .ZN(n6135) );
NAND2_X2 U7226 ( .A1(aes_text_out[19]), .A2(n17995), .ZN(n12276) );
NAND2_X2 U7227 ( .A1(n17986), .A2(n18872), .ZN(n12275) );
NAND2_X2 U7228 ( .A1(n12277), .A2(n12278), .ZN(n6134) );
NAND2_X2 U7229 ( .A1(aes_text_out[20]), .A2(n17995), .ZN(n12278) );
NAND2_X2 U7230 ( .A1(n17986), .A2(n18871), .ZN(n12277) );
NAND2_X2 U7231 ( .A1(n12279), .A2(n12280), .ZN(n6133) );
NAND2_X2 U7232 ( .A1(aes_text_out[21]), .A2(n17995), .ZN(n12280) );
NAND2_X2 U7233 ( .A1(n17986), .A2(n18870), .ZN(n12279) );
NAND2_X2 U7234 ( .A1(n12281), .A2(n12282), .ZN(n6132) );
NAND2_X2 U7235 ( .A1(aes_text_out[22]), .A2(n17995), .ZN(n12282) );
NAND2_X2 U7236 ( .A1(n17986), .A2(n18869), .ZN(n12281) );
NAND2_X2 U7237 ( .A1(n12283), .A2(n12284), .ZN(n6131) );
NAND2_X2 U7238 ( .A1(aes_text_out[23]), .A2(n17995), .ZN(n12284) );
NAND2_X2 U7239 ( .A1(n17986), .A2(n18868), .ZN(n12283) );
NAND2_X2 U7240 ( .A1(n12285), .A2(n12286), .ZN(n6130) );
NAND2_X2 U7241 ( .A1(aes_text_out[24]), .A2(n17994), .ZN(n12286) );
NAND2_X2 U7242 ( .A1(n17986), .A2(n18867), .ZN(n12285) );
NAND2_X2 U7243 ( .A1(n12287), .A2(n12288), .ZN(n6129) );
NAND2_X2 U7244 ( .A1(aes_text_out[25]), .A2(n17994), .ZN(n12288) );
NAND2_X2 U7245 ( .A1(n17986), .A2(n18866), .ZN(n12287) );
NAND2_X2 U7246 ( .A1(n12289), .A2(n12290), .ZN(n6128) );
NAND2_X2 U7247 ( .A1(aes_text_out[26]), .A2(n17994), .ZN(n12290) );
NAND2_X2 U7248 ( .A1(n17986), .A2(n18865), .ZN(n12289) );
NAND2_X2 U7249 ( .A1(n12291), .A2(n12292), .ZN(n6127) );
NAND2_X2 U7250 ( .A1(aes_text_out[27]), .A2(n17994), .ZN(n12292) );
NAND2_X2 U7251 ( .A1(n17986), .A2(n18864), .ZN(n12291) );
NAND2_X2 U7252 ( .A1(n12293), .A2(n12294), .ZN(n6126) );
NAND2_X2 U7253 ( .A1(aes_text_out[28]), .A2(n17994), .ZN(n12294) );
NAND2_X2 U7254 ( .A1(n17986), .A2(n18863), .ZN(n12293) );
NAND2_X2 U7255 ( .A1(n12295), .A2(n12296), .ZN(n6125) );
NAND2_X2 U7256 ( .A1(aes_text_out[29]), .A2(n17994), .ZN(n12296) );
NAND2_X2 U7257 ( .A1(n17985), .A2(n18862), .ZN(n12295) );
NAND2_X2 U7258 ( .A1(n12297), .A2(n12298), .ZN(n6124) );
NAND2_X2 U7259 ( .A1(aes_text_out[30]), .A2(n17994), .ZN(n12298) );
NAND2_X2 U7260 ( .A1(n17985), .A2(n18861), .ZN(n12297) );
NAND2_X2 U7261 ( .A1(n12299), .A2(n12300), .ZN(n6123) );
NAND2_X2 U7262 ( .A1(aes_text_out[31]), .A2(n17994), .ZN(n12300) );
NAND2_X2 U7263 ( .A1(n17985), .A2(n18860), .ZN(n12299) );
NAND2_X2 U7264 ( .A1(n12301), .A2(n12302), .ZN(n6122) );
NAND2_X2 U7265 ( .A1(aes_text_out[32]), .A2(n17994), .ZN(n12302) );
NAND2_X2 U7266 ( .A1(n17985), .A2(n18859), .ZN(n12301) );
NAND2_X2 U7267 ( .A1(n12303), .A2(n12304), .ZN(n6121) );
NAND2_X2 U7268 ( .A1(aes_text_out[33]), .A2(n17994), .ZN(n12304) );
NAND2_X2 U7269 ( .A1(n17985), .A2(n18858), .ZN(n12303) );
NAND2_X2 U7270 ( .A1(n12305), .A2(n12306), .ZN(n6120) );
NAND2_X2 U7271 ( .A1(aes_text_out[34]), .A2(n17994), .ZN(n12306) );
NAND2_X2 U7272 ( .A1(n17985), .A2(n18857), .ZN(n12305) );
NAND2_X2 U7273 ( .A1(n12307), .A2(n12308), .ZN(n6119) );
NAND2_X2 U7274 ( .A1(aes_text_out[35]), .A2(n17994), .ZN(n12308) );
NAND2_X2 U7275 ( .A1(n17985), .A2(n18856), .ZN(n12307) );
NAND2_X2 U7276 ( .A1(n12309), .A2(n12310), .ZN(n6118) );
NAND2_X2 U7277 ( .A1(aes_text_out[36]), .A2(n17994), .ZN(n12310) );
NAND2_X2 U7278 ( .A1(n17985), .A2(n18855), .ZN(n12309) );
NAND2_X2 U7279 ( .A1(n12311), .A2(n12312), .ZN(n6117) );
NAND2_X2 U7280 ( .A1(aes_text_out[37]), .A2(n17994), .ZN(n12312) );
NAND2_X2 U7281 ( .A1(n17985), .A2(n18854), .ZN(n12311) );
NAND2_X2 U7282 ( .A1(n12313), .A2(n12314), .ZN(n6116) );
NAND2_X2 U7283 ( .A1(aes_text_out[38]), .A2(n17994), .ZN(n12314) );
NAND2_X2 U7284 ( .A1(n17985), .A2(n18853), .ZN(n12313) );
NAND2_X2 U7285 ( .A1(n12315), .A2(n12316), .ZN(n6115) );
NAND2_X2 U7286 ( .A1(aes_text_out[39]), .A2(n17994), .ZN(n12316) );
NAND2_X2 U7287 ( .A1(n17985), .A2(n18852), .ZN(n12315) );
NAND2_X2 U7288 ( .A1(n12317), .A2(n12318), .ZN(n6114) );
NAND2_X2 U7289 ( .A1(aes_text_out[40]), .A2(n17994), .ZN(n12318) );
NAND2_X2 U7290 ( .A1(n17984), .A2(n18851), .ZN(n12317) );
NAND2_X2 U7291 ( .A1(n12319), .A2(n12320), .ZN(n6113) );
NAND2_X2 U7292 ( .A1(aes_text_out[41]), .A2(n17994), .ZN(n12320) );
NAND2_X2 U7293 ( .A1(n17984), .A2(n18850), .ZN(n12319) );
NAND2_X2 U7294 ( .A1(n12321), .A2(n12322), .ZN(n6112) );
NAND2_X2 U7295 ( .A1(aes_text_out[42]), .A2(n17994), .ZN(n12322) );
NAND2_X2 U7296 ( .A1(n17984), .A2(n18849), .ZN(n12321) );
NAND2_X2 U7297 ( .A1(n12323), .A2(n12324), .ZN(n6111) );
NAND2_X2 U7298 ( .A1(aes_text_out[43]), .A2(n17994), .ZN(n12324) );
NAND2_X2 U7299 ( .A1(n17984), .A2(n18848), .ZN(n12323) );
NAND2_X2 U7300 ( .A1(n12325), .A2(n12326), .ZN(n6110) );
NAND2_X2 U7301 ( .A1(aes_text_out[44]), .A2(n17994), .ZN(n12326) );
NAND2_X2 U7302 ( .A1(n17984), .A2(n18847), .ZN(n12325) );
NAND2_X2 U7303 ( .A1(n12327), .A2(n12328), .ZN(n6109) );
NAND2_X2 U7304 ( .A1(aes_text_out[45]), .A2(n17993), .ZN(n12328) );
NAND2_X2 U7305 ( .A1(n17984), .A2(n17374), .ZN(n12327) );
NAND2_X2 U7306 ( .A1(n12329), .A2(n12330), .ZN(n6108) );
NAND2_X2 U7307 ( .A1(aes_text_out[46]), .A2(n17993), .ZN(n12330) );
NAND2_X2 U7308 ( .A1(n17984), .A2(n17373), .ZN(n12329) );
NAND2_X2 U7309 ( .A1(n12331), .A2(n12332), .ZN(n6107) );
NAND2_X2 U7310 ( .A1(aes_text_out[47]), .A2(n17993), .ZN(n12332) );
NAND2_X2 U7311 ( .A1(n17984), .A2(n17372), .ZN(n12331) );
NAND2_X2 U7312 ( .A1(n12333), .A2(n12334), .ZN(n6106) );
NAND2_X2 U7313 ( .A1(aes_text_out[48]), .A2(n17993), .ZN(n12334) );
NAND2_X2 U7314 ( .A1(n17984), .A2(n17371), .ZN(n12333) );
NAND2_X2 U7315 ( .A1(n12335), .A2(n12336), .ZN(n6105) );
NAND2_X2 U7316 ( .A1(aes_text_out[49]), .A2(n17993), .ZN(n12336) );
NAND2_X2 U7317 ( .A1(n17984), .A2(n17370), .ZN(n12335) );
NAND2_X2 U7318 ( .A1(n12337), .A2(n12338), .ZN(n6104) );
NAND2_X2 U7319 ( .A1(aes_text_out[50]), .A2(n17993), .ZN(n12338) );
NAND2_X2 U7320 ( .A1(n17984), .A2(n17369), .ZN(n12337) );
NAND2_X2 U7321 ( .A1(n12339), .A2(n12340), .ZN(n6103) );
NAND2_X2 U7322 ( .A1(aes_text_out[51]), .A2(n17993), .ZN(n12340) );
NAND2_X2 U7323 ( .A1(n17983), .A2(n17368), .ZN(n12339) );
NAND2_X2 U7324 ( .A1(n12341), .A2(n12342), .ZN(n6102) );
NAND2_X2 U7325 ( .A1(aes_text_out[52]), .A2(n17993), .ZN(n12342) );
NAND2_X2 U7326 ( .A1(n17983), .A2(n17367), .ZN(n12341) );
NAND2_X2 U7327 ( .A1(n12343), .A2(n12344), .ZN(n6101) );
NAND2_X2 U7328 ( .A1(aes_text_out[53]), .A2(n17993), .ZN(n12344) );
NAND2_X2 U7329 ( .A1(n17983), .A2(n17366), .ZN(n12343) );
NAND2_X2 U7330 ( .A1(n12345), .A2(n12346), .ZN(n6100) );
NAND2_X2 U7331 ( .A1(aes_text_out[54]), .A2(n17993), .ZN(n12346) );
NAND2_X2 U7332 ( .A1(n17983), .A2(n17365), .ZN(n12345) );
NAND2_X2 U7333 ( .A1(n12347), .A2(n12348), .ZN(n6099) );
NAND2_X2 U7334 ( .A1(aes_text_out[55]), .A2(n17993), .ZN(n12348) );
NAND2_X2 U7335 ( .A1(n17983), .A2(n17364), .ZN(n12347) );
NAND2_X2 U7336 ( .A1(n12349), .A2(n12350), .ZN(n6098) );
NAND2_X2 U7337 ( .A1(aes_text_out[56]), .A2(n17993), .ZN(n12350) );
NAND2_X2 U7338 ( .A1(n17983), .A2(n17363), .ZN(n12349) );
NAND2_X2 U7339 ( .A1(n12351), .A2(n12352), .ZN(n6097) );
NAND2_X2 U7340 ( .A1(aes_text_out[57]), .A2(n17993), .ZN(n12352) );
NAND2_X2 U7341 ( .A1(n17983), .A2(n17362), .ZN(n12351) );
NAND2_X2 U7342 ( .A1(n12353), .A2(n12354), .ZN(n6096) );
NAND2_X2 U7343 ( .A1(aes_text_out[58]), .A2(n17993), .ZN(n12354) );
NAND2_X2 U7344 ( .A1(n17983), .A2(n17361), .ZN(n12353) );
NAND2_X2 U7345 ( .A1(n12355), .A2(n12356), .ZN(n6095) );
NAND2_X2 U7346 ( .A1(aes_text_out[59]), .A2(n17993), .ZN(n12356) );
NAND2_X2 U7347 ( .A1(n17983), .A2(n17360), .ZN(n12355) );
NAND2_X2 U7348 ( .A1(n12357), .A2(n12358), .ZN(n6094) );
NAND2_X2 U7349 ( .A1(aes_text_out[60]), .A2(n17993), .ZN(n12358) );
NAND2_X2 U7350 ( .A1(n17983), .A2(n17359), .ZN(n12357) );
NAND2_X2 U7351 ( .A1(n12359), .A2(n12360), .ZN(n6093) );
NAND2_X2 U7352 ( .A1(aes_text_out[61]), .A2(n17993), .ZN(n12360) );
NAND2_X2 U7353 ( .A1(n17983), .A2(n17358), .ZN(n12359) );
NAND2_X2 U7354 ( .A1(n12361), .A2(n12362), .ZN(n6092) );
NAND2_X2 U7355 ( .A1(aes_text_out[62]), .A2(n17993), .ZN(n12362) );
NAND2_X2 U7356 ( .A1(n17982), .A2(n17357), .ZN(n12361) );
NAND2_X2 U7357 ( .A1(n12363), .A2(n12364), .ZN(n6091) );
NAND2_X2 U7358 ( .A1(aes_text_out[63]), .A2(n17993), .ZN(n12364) );
NAND2_X2 U7359 ( .A1(n17982), .A2(n17356), .ZN(n12363) );
NAND2_X2 U7360 ( .A1(n12365), .A2(n12366), .ZN(n6090) );
NAND2_X2 U7361 ( .A1(aes_text_out[64]), .A2(n17993), .ZN(n12366) );
NAND2_X2 U7362 ( .A1(n17982), .A2(n17355), .ZN(n12365) );
NAND2_X2 U7363 ( .A1(n12367), .A2(n12368), .ZN(n6089) );
NAND2_X2 U7364 ( .A1(aes_text_out[65]), .A2(n17993), .ZN(n12368) );
NAND2_X2 U7365 ( .A1(n17982), .A2(n17354), .ZN(n12367) );
NAND2_X2 U7366 ( .A1(n12369), .A2(n12370), .ZN(n6088) );
NAND2_X2 U7367 ( .A1(aes_text_out[66]), .A2(n17992), .ZN(n12370) );
NAND2_X2 U7368 ( .A1(n17982), .A2(n17353), .ZN(n12369) );
NAND2_X2 U7369 ( .A1(n12371), .A2(n12372), .ZN(n6087) );
NAND2_X2 U7370 ( .A1(aes_text_out[67]), .A2(n17992), .ZN(n12372) );
NAND2_X2 U7371 ( .A1(n17982), .A2(n17352), .ZN(n12371) );
NAND2_X2 U7372 ( .A1(n12373), .A2(n12374), .ZN(n6086) );
NAND2_X2 U7373 ( .A1(aes_text_out[68]), .A2(n17992), .ZN(n12374) );
NAND2_X2 U7374 ( .A1(n17982), .A2(n17351), .ZN(n12373) );
NAND2_X2 U7375 ( .A1(n12375), .A2(n12376), .ZN(n6085) );
NAND2_X2 U7376 ( .A1(aes_text_out[69]), .A2(n17992), .ZN(n12376) );
NAND2_X2 U7377 ( .A1(n17982), .A2(n17350), .ZN(n12375) );
NAND2_X2 U7378 ( .A1(n12377), .A2(n12378), .ZN(n6084) );
NAND2_X2 U7379 ( .A1(aes_text_out[70]), .A2(n17992), .ZN(n12378) );
NAND2_X2 U7380 ( .A1(n17982), .A2(n17349), .ZN(n12377) );
NAND2_X2 U7381 ( .A1(n12379), .A2(n12380), .ZN(n6083) );
NAND2_X2 U7382 ( .A1(aes_text_out[71]), .A2(n17992), .ZN(n12380) );
NAND2_X2 U7383 ( .A1(n17982), .A2(n17348), .ZN(n12379) );
NAND2_X2 U7384 ( .A1(n12381), .A2(n12382), .ZN(n6082) );
NAND2_X2 U7385 ( .A1(aes_text_out[72]), .A2(n17992), .ZN(n12382) );
NAND2_X2 U7386 ( .A1(n17982), .A2(n17347), .ZN(n12381) );
NAND2_X2 U7387 ( .A1(n12383), .A2(n12384), .ZN(n6081) );
NAND2_X2 U7388 ( .A1(aes_text_out[73]), .A2(n17992), .ZN(n12384) );
NAND2_X2 U7389 ( .A1(n17981), .A2(n17346), .ZN(n12383) );
NAND2_X2 U7390 ( .A1(n12385), .A2(n12386), .ZN(n6080) );
NAND2_X2 U7391 ( .A1(aes_text_out[74]), .A2(n17992), .ZN(n12386) );
NAND2_X2 U7392 ( .A1(n17981), .A2(n17345), .ZN(n12385) );
NAND2_X2 U7393 ( .A1(n12387), .A2(n12388), .ZN(n6079) );
NAND2_X2 U7394 ( .A1(aes_text_out[75]), .A2(n17992), .ZN(n12388) );
NAND2_X2 U7395 ( .A1(n17981), .A2(n17344), .ZN(n12387) );
NAND2_X2 U7396 ( .A1(n12389), .A2(n12390), .ZN(n6078) );
NAND2_X2 U7397 ( .A1(aes_text_out[76]), .A2(n17992), .ZN(n12390) );
NAND2_X2 U7398 ( .A1(n17981), .A2(n17343), .ZN(n12389) );
NAND2_X2 U7399 ( .A1(n12391), .A2(n12392), .ZN(n6077) );
NAND2_X2 U7400 ( .A1(aes_text_out[77]), .A2(n17992), .ZN(n12392) );
NAND2_X2 U7401 ( .A1(n17981), .A2(n17342), .ZN(n12391) );
NAND2_X2 U7402 ( .A1(n12393), .A2(n12394), .ZN(n6076) );
NAND2_X2 U7403 ( .A1(aes_text_out[78]), .A2(n17992), .ZN(n12394) );
NAND2_X2 U7404 ( .A1(n17981), .A2(n17341), .ZN(n12393) );
NAND2_X2 U7405 ( .A1(n12395), .A2(n12396), .ZN(n6075) );
NAND2_X2 U7406 ( .A1(aes_text_out[79]), .A2(n17992), .ZN(n12396) );
NAND2_X2 U7407 ( .A1(n17981), .A2(n17340), .ZN(n12395) );
NAND2_X2 U7408 ( .A1(n12397), .A2(n12398), .ZN(n6074) );
NAND2_X2 U7409 ( .A1(aes_text_out[80]), .A2(n17992), .ZN(n12398) );
NAND2_X2 U7410 ( .A1(n17981), .A2(n17339), .ZN(n12397) );
NAND2_X2 U7411 ( .A1(n12399), .A2(n12400), .ZN(n6073) );
NAND2_X2 U7412 ( .A1(aes_text_out[81]), .A2(n17992), .ZN(n12400) );
NAND2_X2 U7413 ( .A1(n17981), .A2(n17338), .ZN(n12399) );
NAND2_X2 U7414 ( .A1(n12401), .A2(n12402), .ZN(n6072) );
NAND2_X2 U7415 ( .A1(aes_text_out[82]), .A2(n17992), .ZN(n12402) );
NAND2_X2 U7416 ( .A1(n17981), .A2(n17337), .ZN(n12401) );
NAND2_X2 U7417 ( .A1(n12403), .A2(n12404), .ZN(n6071) );
NAND2_X2 U7418 ( .A1(aes_text_out[83]), .A2(n17992), .ZN(n12404) );
NAND2_X2 U7419 ( .A1(n17981), .A2(n17336), .ZN(n12403) );
NAND2_X2 U7420 ( .A1(n12405), .A2(n12406), .ZN(n6070) );
NAND2_X2 U7421 ( .A1(aes_text_out[84]), .A2(n17992), .ZN(n12406) );
NAND2_X2 U7422 ( .A1(n17980), .A2(n17335), .ZN(n12405) );
NAND2_X2 U7423 ( .A1(n12407), .A2(n12408), .ZN(n6069) );
NAND2_X2 U7424 ( .A1(aes_text_out[85]), .A2(n17992), .ZN(n12408) );
NAND2_X2 U7425 ( .A1(n17980), .A2(n17334), .ZN(n12407) );
NAND2_X2 U7426 ( .A1(n12409), .A2(n12410), .ZN(n6068) );
NAND2_X2 U7427 ( .A1(aes_text_out[86]), .A2(n17992), .ZN(n12410) );
NAND2_X2 U7428 ( .A1(n17980), .A2(n17333), .ZN(n12409) );
NAND2_X2 U7429 ( .A1(n12411), .A2(n12412), .ZN(n6067) );
NAND2_X2 U7430 ( .A1(aes_text_out[87]), .A2(n17991), .ZN(n12412) );
NAND2_X2 U7431 ( .A1(n17980), .A2(n17332), .ZN(n12411) );
NAND2_X2 U7432 ( .A1(n12413), .A2(n12414), .ZN(n6066) );
NAND2_X2 U7433 ( .A1(aes_text_out[88]), .A2(n17991), .ZN(n12414) );
NAND2_X2 U7434 ( .A1(n17980), .A2(n17331), .ZN(n12413) );
NAND2_X2 U7435 ( .A1(n12415), .A2(n12416), .ZN(n6065) );
NAND2_X2 U7436 ( .A1(aes_text_out[89]), .A2(n17991), .ZN(n12416) );
NAND2_X2 U7437 ( .A1(n17980), .A2(n17330), .ZN(n12415) );
NAND2_X2 U7438 ( .A1(n12417), .A2(n12418), .ZN(n6064) );
NAND2_X2 U7439 ( .A1(aes_text_out[90]), .A2(n17991), .ZN(n12418) );
NAND2_X2 U7440 ( .A1(n17980), .A2(n17329), .ZN(n12417) );
NAND2_X2 U7441 ( .A1(n12419), .A2(n12420), .ZN(n6063) );
NAND2_X2 U7442 ( .A1(aes_text_out[91]), .A2(n17991), .ZN(n12420) );
NAND2_X2 U7443 ( .A1(n17980), .A2(n17328), .ZN(n12419) );
NAND2_X2 U7444 ( .A1(n12421), .A2(n12422), .ZN(n6062) );
NAND2_X2 U7445 ( .A1(aes_text_out[92]), .A2(n17991), .ZN(n12422) );
NAND2_X2 U7446 ( .A1(n17980), .A2(n17327), .ZN(n12421) );
NAND2_X2 U7447 ( .A1(n12423), .A2(n12424), .ZN(n6061) );
NAND2_X2 U7448 ( .A1(aes_text_out[93]), .A2(n17991), .ZN(n12424) );
NAND2_X2 U7449 ( .A1(n17980), .A2(n17326), .ZN(n12423) );
NAND2_X2 U7450 ( .A1(n12425), .A2(n12426), .ZN(n6060) );
NAND2_X2 U7451 ( .A1(aes_text_out[94]), .A2(n17991), .ZN(n12426) );
NAND2_X2 U7452 ( .A1(n17980), .A2(n17325), .ZN(n12425) );
NAND2_X2 U7453 ( .A1(n12427), .A2(n12428), .ZN(n6059) );
NAND2_X2 U7454 ( .A1(aes_text_out[95]), .A2(n17991), .ZN(n12428) );
NAND2_X2 U7455 ( .A1(n17979), .A2(n17324), .ZN(n12427) );
NAND2_X2 U7456 ( .A1(n12429), .A2(n12430), .ZN(n6058) );
NAND2_X2 U7457 ( .A1(aes_text_out[96]), .A2(n17991), .ZN(n12430) );
NAND2_X2 U7458 ( .A1(n17979), .A2(n17323), .ZN(n12429) );
NAND2_X2 U7459 ( .A1(n12431), .A2(n12432), .ZN(n6057) );
NAND2_X2 U7460 ( .A1(aes_text_out[97]), .A2(n17991), .ZN(n12432) );
NAND2_X2 U7461 ( .A1(n17979), .A2(n17322), .ZN(n12431) );
NAND2_X2 U7462 ( .A1(n12433), .A2(n12434), .ZN(n6056) );
NAND2_X2 U7463 ( .A1(aes_text_out[98]), .A2(n17991), .ZN(n12434) );
NAND2_X2 U7464 ( .A1(n17979), .A2(n17321), .ZN(n12433) );
NAND2_X2 U7465 ( .A1(n12435), .A2(n12436), .ZN(n6055) );
NAND2_X2 U7466 ( .A1(aes_text_out[99]), .A2(n17991), .ZN(n12436) );
NAND2_X2 U7467 ( .A1(n17979), .A2(n17320), .ZN(n12435) );
NAND2_X2 U7468 ( .A1(n12437), .A2(n12438), .ZN(n6054) );
NAND2_X2 U7469 ( .A1(aes_text_out[100]), .A2(n17991), .ZN(n12438) );
NAND2_X2 U7470 ( .A1(n17979), .A2(n17319), .ZN(n12437) );
NAND2_X2 U7471 ( .A1(n12439), .A2(n12440), .ZN(n6053) );
NAND2_X2 U7472 ( .A1(aes_text_out[101]), .A2(n17991), .ZN(n12440) );
NAND2_X2 U7473 ( .A1(n17979), .A2(n17318), .ZN(n12439) );
NAND2_X2 U7474 ( .A1(n12441), .A2(n12442), .ZN(n6052) );
NAND2_X2 U7475 ( .A1(aes_text_out[102]), .A2(n17991), .ZN(n12442) );
NAND2_X2 U7476 ( .A1(n17979), .A2(n17317), .ZN(n12441) );
NAND2_X2 U7477 ( .A1(n12443), .A2(n12444), .ZN(n6051) );
NAND2_X2 U7478 ( .A1(aes_text_out[103]), .A2(n17991), .ZN(n12444) );
NAND2_X2 U7479 ( .A1(n17979), .A2(n17316), .ZN(n12443) );
NAND2_X2 U7480 ( .A1(n12445), .A2(n12446), .ZN(n6050) );
NAND2_X2 U7481 ( .A1(aes_text_out[104]), .A2(n17991), .ZN(n12446) );
NAND2_X2 U7482 ( .A1(n17979), .A2(n17315), .ZN(n12445) );
NAND2_X2 U7483 ( .A1(n12447), .A2(n12448), .ZN(n6049) );
NAND2_X2 U7484 ( .A1(aes_text_out[105]), .A2(n17991), .ZN(n12448) );
NAND2_X2 U7485 ( .A1(n17979), .A2(n17314), .ZN(n12447) );
NAND2_X2 U7486 ( .A1(n12449), .A2(n12450), .ZN(n6048) );
NAND2_X2 U7487 ( .A1(aes_text_out[106]), .A2(n17991), .ZN(n12450) );
NAND2_X2 U7488 ( .A1(n17978), .A2(n17313), .ZN(n12449) );
NAND2_X2 U7489 ( .A1(n12451), .A2(n12452), .ZN(n6047) );
NAND2_X2 U7490 ( .A1(aes_text_out[107]), .A2(n17991), .ZN(n12452) );
NAND2_X2 U7491 ( .A1(n17978), .A2(n17312), .ZN(n12451) );
NAND2_X2 U7492 ( .A1(n12453), .A2(n12454), .ZN(n6046) );
NAND2_X2 U7493 ( .A1(aes_text_out[108]), .A2(n17990), .ZN(n12454) );
NAND2_X2 U7494 ( .A1(n17978), .A2(n17311), .ZN(n12453) );
NAND2_X2 U7495 ( .A1(n12455), .A2(n12456), .ZN(n6045) );
NAND2_X2 U7496 ( .A1(aes_text_out[109]), .A2(n17990), .ZN(n12456) );
NAND2_X2 U7497 ( .A1(n17978), .A2(n17310), .ZN(n12455) );
NAND2_X2 U7498 ( .A1(n12457), .A2(n12458), .ZN(n6044) );
NAND2_X2 U7499 ( .A1(aes_text_out[110]), .A2(n17990), .ZN(n12458) );
NAND2_X2 U7500 ( .A1(n17978), .A2(n17309), .ZN(n12457) );
NAND2_X2 U7501 ( .A1(n12459), .A2(n12460), .ZN(n6043) );
NAND2_X2 U7502 ( .A1(aes_text_out[111]), .A2(n17990), .ZN(n12460) );
NAND2_X2 U7503 ( .A1(n17978), .A2(n17308), .ZN(n12459) );
NAND2_X2 U7504 ( .A1(n12461), .A2(n12462), .ZN(n6042) );
NAND2_X2 U7505 ( .A1(aes_text_out[112]), .A2(n17990), .ZN(n12462) );
NAND2_X2 U7506 ( .A1(n17978), .A2(n17307), .ZN(n12461) );
NAND2_X2 U7507 ( .A1(n12463), .A2(n12464), .ZN(n6041) );
NAND2_X2 U7508 ( .A1(aes_text_out[113]), .A2(n17990), .ZN(n12464) );
NAND2_X2 U7509 ( .A1(n17978), .A2(n17306), .ZN(n12463) );
NAND2_X2 U7510 ( .A1(n12465), .A2(n12466), .ZN(n6040) );
NAND2_X2 U7511 ( .A1(aes_text_out[114]), .A2(n17990), .ZN(n12466) );
NAND2_X2 U7512 ( .A1(n17978), .A2(n17305), .ZN(n12465) );
NAND2_X2 U7513 ( .A1(n12467), .A2(n12468), .ZN(n6039) );
NAND2_X2 U7514 ( .A1(aes_text_out[115]), .A2(n17990), .ZN(n12468) );
NAND2_X2 U7515 ( .A1(n17978), .A2(n17304), .ZN(n12467) );
NAND2_X2 U7516 ( .A1(n12469), .A2(n12470), .ZN(n6038) );
NAND2_X2 U7517 ( .A1(aes_text_out[116]), .A2(n17990), .ZN(n12470) );
NAND2_X2 U7518 ( .A1(n17978), .A2(n17303), .ZN(n12469) );
NAND2_X2 U7519 ( .A1(n12471), .A2(n12472), .ZN(n6037) );
NAND2_X2 U7520 ( .A1(aes_text_out[117]), .A2(n17990), .ZN(n12472) );
NAND2_X2 U7521 ( .A1(n17977), .A2(n17302), .ZN(n12471) );
NAND2_X2 U7522 ( .A1(n12473), .A2(n12474), .ZN(n6036) );
NAND2_X2 U7523 ( .A1(aes_text_out[118]), .A2(n17990), .ZN(n12474) );
NAND2_X2 U7524 ( .A1(n17977), .A2(n17301), .ZN(n12473) );
NAND2_X2 U7525 ( .A1(n12475), .A2(n12476), .ZN(n6035) );
NAND2_X2 U7526 ( .A1(aes_text_out[119]), .A2(n17990), .ZN(n12476) );
NAND2_X2 U7527 ( .A1(n17977), .A2(n17300), .ZN(n12475) );
NAND2_X2 U7528 ( .A1(n12477), .A2(n12478), .ZN(n6034) );
NAND2_X2 U7529 ( .A1(aes_text_out[120]), .A2(n17990), .ZN(n12478) );
NAND2_X2 U7530 ( .A1(n17977), .A2(n17299), .ZN(n12477) );
NAND2_X2 U7531 ( .A1(n12479), .A2(n12480), .ZN(n6033) );
NAND2_X2 U7532 ( .A1(aes_text_out[121]), .A2(n17990), .ZN(n12480) );
NAND2_X2 U7533 ( .A1(n17977), .A2(n17298), .ZN(n12479) );
NAND2_X2 U7534 ( .A1(n12481), .A2(n12482), .ZN(n6032) );
NAND2_X2 U7535 ( .A1(aes_text_out[122]), .A2(n17990), .ZN(n12482) );
NAND2_X2 U7536 ( .A1(n17977), .A2(n17297), .ZN(n12481) );
NAND2_X2 U7537 ( .A1(n12483), .A2(n12484), .ZN(n6031) );
NAND2_X2 U7538 ( .A1(aes_text_out[123]), .A2(n17990), .ZN(n12484) );
NAND2_X2 U7539 ( .A1(n17977), .A2(n17296), .ZN(n12483) );
NAND2_X2 U7540 ( .A1(n12485), .A2(n12486), .ZN(n6030) );
NAND2_X2 U7541 ( .A1(aes_text_out[124]), .A2(n17990), .ZN(n12486) );
NAND2_X2 U7542 ( .A1(n17977), .A2(n17295), .ZN(n12485) );
NAND2_X2 U7543 ( .A1(n12487), .A2(n12488), .ZN(n6029) );
NAND2_X2 U7544 ( .A1(aes_text_out[125]), .A2(n17990), .ZN(n12488) );
NAND2_X2 U7545 ( .A1(n17977), .A2(n17294), .ZN(n12487) );
NAND2_X2 U7546 ( .A1(n12489), .A2(n12490), .ZN(n6028) );
NAND2_X2 U7547 ( .A1(aes_text_out[126]), .A2(n17990), .ZN(n12490) );
NAND2_X2 U7548 ( .A1(n17977), .A2(n17293), .ZN(n12489) );
NAND2_X2 U7549 ( .A1(n12491), .A2(n12492), .ZN(n6027) );
NAND2_X2 U7550 ( .A1(aes_text_out[127]), .A2(n17990), .ZN(n12492) );
NAND2_X2 U7551 ( .A1(n17977), .A2(n17292), .ZN(n12491) );
NAND2_X2 U7552 ( .A1(n12493), .A2(n12494), .ZN(n6026) );
NAND2_X2 U7553 ( .A1(n17750), .A2(n17281), .ZN(n12494) );
NAND2_X2 U7554 ( .A1(n18744), .A2(Out_data_size[0]), .ZN(n12493) );
NAND2_X2 U7557 ( .A1(n18744), .A2(Out_data_size[1]), .ZN(n12495) );
NAND2_X2 U7560 ( .A1(n18744), .A2(Out_data_size[2]), .ZN(n12497) );
NAND2_X2 U7561 ( .A1(n12499), .A2(n12500), .ZN(n6023) );
NAND2_X2 U7562 ( .A1(n18074), .A2(n17281), .ZN(n12500) );
NAND2_X2 U7563 ( .A1(n18744), .A2(Out_data_size[3]), .ZN(n12499) );
NAND2_X2 U7564 ( .A1(n12501), .A2(n12502), .ZN(n6022) );
NAND2_X2 U7565 ( .A1(n17281), .A2(n17748), .ZN(n12502) );
NAND2_X2 U7566 ( .A1(n18744), .A2(Out_last_word), .ZN(n12501) );
NAND2_X2 U8275 ( .A1(n11967), .A2(aes_done), .ZN(n12238) );
AND4_X2 U8276 ( .A1(state[1]), .A2(n18628), .A3(n18625), .A4(n18629), .ZN(n11967) );
NAND2_X2 U8277 ( .A1(n13019), .A2(n13020), .ZN(n5829) );
NAND2_X2 U8278 ( .A1(n17976), .A2(n18895), .ZN(n13020) );
NAND2_X2 U8279 ( .A1(z_out[0]), .A2(n17961), .ZN(n13019) );
NAND2_X2 U8280 ( .A1(n13023), .A2(n13024), .ZN(n5828) );
NAND2_X2 U8281 ( .A1(n17976), .A2(n18896), .ZN(n13024) );
NAND2_X2 U8282 ( .A1(z_out[1]), .A2(n17958), .ZN(n13023) );
NAND2_X2 U8283 ( .A1(n13025), .A2(n13026), .ZN(n5827) );
NAND2_X2 U8284 ( .A1(n17976), .A2(n18897), .ZN(n13026) );
NAND2_X2 U8285 ( .A1(z_out[2]), .A2(n17958), .ZN(n13025) );
NAND2_X2 U8286 ( .A1(n13027), .A2(n13028), .ZN(n5826) );
NAND2_X2 U8287 ( .A1(n17976), .A2(n18898), .ZN(n13028) );
NAND2_X2 U8288 ( .A1(z_out[3]), .A2(n17958), .ZN(n13027) );
NAND2_X2 U8289 ( .A1(n13029), .A2(n13030), .ZN(n5825) );
NAND2_X2 U8290 ( .A1(n17976), .A2(n18899), .ZN(n13030) );
NAND2_X2 U8291 ( .A1(z_out[4]), .A2(n17958), .ZN(n13029) );
NAND2_X2 U8292 ( .A1(n13031), .A2(n13032), .ZN(n5824) );
NAND2_X2 U8293 ( .A1(n17976), .A2(n18900), .ZN(n13032) );
NAND2_X2 U8294 ( .A1(z_out[5]), .A2(n17958), .ZN(n13031) );
NAND2_X2 U8295 ( .A1(n13033), .A2(n13034), .ZN(n5823) );
NAND2_X2 U8296 ( .A1(n17976), .A2(n18901), .ZN(n13034) );
NAND2_X2 U8297 ( .A1(z_out[6]), .A2(n17958), .ZN(n13033) );
NAND2_X2 U8298 ( .A1(n13035), .A2(n13036), .ZN(n5822) );
NAND2_X2 U8299 ( .A1(n17975), .A2(n18902), .ZN(n13036) );
NAND2_X2 U8300 ( .A1(z_out[7]), .A2(n17958), .ZN(n13035) );
NAND2_X2 U8301 ( .A1(n13037), .A2(n13038), .ZN(n5821) );
NAND2_X2 U8302 ( .A1(n17975), .A2(n18903), .ZN(n13038) );
NAND2_X2 U8303 ( .A1(z_out[8]), .A2(n17958), .ZN(n13037) );
NAND2_X2 U8304 ( .A1(n13039), .A2(n13040), .ZN(n5820) );
NAND2_X2 U8305 ( .A1(n17975), .A2(n18904), .ZN(n13040) );
NAND2_X2 U8306 ( .A1(z_out[9]), .A2(n17958), .ZN(n13039) );
NAND2_X2 U8307 ( .A1(n13041), .A2(n13042), .ZN(n5819) );
NAND2_X2 U8308 ( .A1(n17975), .A2(n18905), .ZN(n13042) );
NAND2_X2 U8309 ( .A1(z_out[10]), .A2(n17958), .ZN(n13041) );
NAND2_X2 U8310 ( .A1(n13043), .A2(n13044), .ZN(n5818) );
NAND2_X2 U8311 ( .A1(n17975), .A2(n18906), .ZN(n13044) );
NAND2_X2 U8312 ( .A1(z_out[11]), .A2(n17958), .ZN(n13043) );
NAND2_X2 U8313 ( .A1(n13045), .A2(n13046), .ZN(n5817) );
NAND2_X2 U8314 ( .A1(n17975), .A2(n18907), .ZN(n13046) );
NAND2_X2 U8315 ( .A1(z_out[12]), .A2(n17958), .ZN(n13045) );
NAND2_X2 U8316 ( .A1(n13047), .A2(n13048), .ZN(n5816) );
NAND2_X2 U8317 ( .A1(n17975), .A2(n18908), .ZN(n13048) );
NAND2_X2 U8318 ( .A1(z_out[13]), .A2(n17958), .ZN(n13047) );
NAND2_X2 U8319 ( .A1(n13049), .A2(n13050), .ZN(n5815) );
NAND2_X2 U8320 ( .A1(n17975), .A2(n18909), .ZN(n13050) );
NAND2_X2 U8321 ( .A1(z_out[14]), .A2(n17958), .ZN(n13049) );
NAND2_X2 U8322 ( .A1(n13051), .A2(n13052), .ZN(n5814) );
NAND2_X2 U8323 ( .A1(n17975), .A2(n18910), .ZN(n13052) );
NAND2_X2 U8324 ( .A1(z_out[15]), .A2(n17958), .ZN(n13051) );
NAND2_X2 U8325 ( .A1(n13053), .A2(n13054), .ZN(n5813) );
NAND2_X2 U8326 ( .A1(n17975), .A2(n18911), .ZN(n13054) );
NAND2_X2 U8327 ( .A1(z_out[16]), .A2(n17958), .ZN(n13053) );
NAND2_X2 U8328 ( .A1(n13055), .A2(n13056), .ZN(n5812) );
NAND2_X2 U8329 ( .A1(n17975), .A2(n18912), .ZN(n13056) );
NAND2_X2 U8330 ( .A1(z_out[17]), .A2(n17958), .ZN(n13055) );
NAND2_X2 U8331 ( .A1(n13057), .A2(n13058), .ZN(n5811) );
NAND2_X2 U8332 ( .A1(n17974), .A2(n18913), .ZN(n13058) );
NAND2_X2 U8333 ( .A1(z_out[18]), .A2(n17959), .ZN(n13057) );
NAND2_X2 U8334 ( .A1(n13059), .A2(n13060), .ZN(n5810) );
NAND2_X2 U8335 ( .A1(n17974), .A2(n18914), .ZN(n13060) );
NAND2_X2 U8336 ( .A1(z_out[19]), .A2(n17959), .ZN(n13059) );
NAND2_X2 U8337 ( .A1(n13061), .A2(n13062), .ZN(n5809) );
NAND2_X2 U8338 ( .A1(n17974), .A2(n18915), .ZN(n13062) );
NAND2_X2 U8339 ( .A1(z_out[20]), .A2(n17959), .ZN(n13061) );
NAND2_X2 U8340 ( .A1(n13063), .A2(n13064), .ZN(n5808) );
NAND2_X2 U8341 ( .A1(n17974), .A2(n18916), .ZN(n13064) );
NAND2_X2 U8342 ( .A1(z_out[21]), .A2(n17959), .ZN(n13063) );
NAND2_X2 U8343 ( .A1(n13065), .A2(n13066), .ZN(n5807) );
NAND2_X2 U8344 ( .A1(n17974), .A2(n18917), .ZN(n13066) );
NAND2_X2 U8345 ( .A1(z_out[22]), .A2(n17959), .ZN(n13065) );
NAND2_X2 U8346 ( .A1(n13067), .A2(n13068), .ZN(n5806) );
NAND2_X2 U8347 ( .A1(n17974), .A2(n18918), .ZN(n13068) );
NAND2_X2 U8348 ( .A1(z_out[23]), .A2(n17959), .ZN(n13067) );
NAND2_X2 U8349 ( .A1(n13069), .A2(n13070), .ZN(n5805) );
NAND2_X2 U8350 ( .A1(n17974), .A2(n18919), .ZN(n13070) );
NAND2_X2 U8351 ( .A1(z_out[24]), .A2(n17959), .ZN(n13069) );
NAND2_X2 U8352 ( .A1(n13071), .A2(n13072), .ZN(n5804) );
NAND2_X2 U8353 ( .A1(n17974), .A2(n18920), .ZN(n13072) );
NAND2_X2 U8354 ( .A1(z_out[25]), .A2(n17959), .ZN(n13071) );
NAND2_X2 U8355 ( .A1(n13073), .A2(n13074), .ZN(n5803) );
NAND2_X2 U8356 ( .A1(n17974), .A2(n18921), .ZN(n13074) );
NAND2_X2 U8357 ( .A1(z_out[26]), .A2(n17959), .ZN(n13073) );
NAND2_X2 U8358 ( .A1(n13075), .A2(n13076), .ZN(n5802) );
NAND2_X2 U8359 ( .A1(n17974), .A2(n18922), .ZN(n13076) );
NAND2_X2 U8360 ( .A1(z_out[27]), .A2(n17959), .ZN(n13075) );
NAND2_X2 U8361 ( .A1(n13077), .A2(n13078), .ZN(n5801) );
NAND2_X2 U8362 ( .A1(n17974), .A2(n18923), .ZN(n13078) );
NAND2_X2 U8363 ( .A1(z_out[28]), .A2(n17959), .ZN(n13077) );
NAND2_X2 U8364 ( .A1(n13079), .A2(n13080), .ZN(n5800) );
NAND2_X2 U8365 ( .A1(n17973), .A2(n18924), .ZN(n13080) );
NAND2_X2 U8366 ( .A1(z_out[29]), .A2(n17959), .ZN(n13079) );
NAND2_X2 U8367 ( .A1(n13081), .A2(n13082), .ZN(n5799) );
NAND2_X2 U8368 ( .A1(n17973), .A2(n18925), .ZN(n13082) );
NAND2_X2 U8369 ( .A1(z_out[30]), .A2(n17959), .ZN(n13081) );
NAND2_X2 U8370 ( .A1(n13083), .A2(n13084), .ZN(n5798) );
NAND2_X2 U8371 ( .A1(n17973), .A2(n18926), .ZN(n13084) );
NAND2_X2 U8372 ( .A1(z_out[31]), .A2(n17959), .ZN(n13083) );
NAND2_X2 U8373 ( .A1(n13085), .A2(n13086), .ZN(n5797) );
NAND2_X2 U8374 ( .A1(n17973), .A2(n18927), .ZN(n13086) );
NAND2_X2 U8375 ( .A1(z_out[32]), .A2(n17959), .ZN(n13085) );
NAND2_X2 U8376 ( .A1(n13087), .A2(n13088), .ZN(n5796) );
NAND2_X2 U8377 ( .A1(n17973), .A2(n18928), .ZN(n13088) );
NAND2_X2 U8378 ( .A1(z_out[33]), .A2(n17959), .ZN(n13087) );
NAND2_X2 U8379 ( .A1(n13089), .A2(n13090), .ZN(n5795) );
NAND2_X2 U8380 ( .A1(n17973), .A2(n18929), .ZN(n13090) );
NAND2_X2 U8381 ( .A1(z_out[34]), .A2(n17959), .ZN(n13089) );
NAND2_X2 U8382 ( .A1(n13091), .A2(n13092), .ZN(n5794) );
NAND2_X2 U8383 ( .A1(n17973), .A2(n18930), .ZN(n13092) );
NAND2_X2 U8384 ( .A1(z_out[35]), .A2(n17959), .ZN(n13091) );
NAND2_X2 U8385 ( .A1(n13093), .A2(n13094), .ZN(n5793) );
NAND2_X2 U8386 ( .A1(n17973), .A2(n18931), .ZN(n13094) );
NAND2_X2 U8387 ( .A1(z_out[36]), .A2(n17959), .ZN(n13093) );
NAND2_X2 U8388 ( .A1(n13095), .A2(n13096), .ZN(n5792) );
NAND2_X2 U8389 ( .A1(n17973), .A2(n18932), .ZN(n13096) );
NAND2_X2 U8390 ( .A1(z_out[37]), .A2(n17960), .ZN(n13095) );
NAND2_X2 U8391 ( .A1(n13097), .A2(n13098), .ZN(n5791) );
NAND2_X2 U8392 ( .A1(n17973), .A2(n18933), .ZN(n13098) );
NAND2_X2 U8393 ( .A1(z_out[38]), .A2(n17960), .ZN(n13097) );
NAND2_X2 U8394 ( .A1(n13099), .A2(n13100), .ZN(n5790) );
NAND2_X2 U8395 ( .A1(n17973), .A2(n18934), .ZN(n13100) );
NAND2_X2 U8396 ( .A1(z_out[39]), .A2(n17960), .ZN(n13099) );
NAND2_X2 U8397 ( .A1(n13101), .A2(n13102), .ZN(n5789) );
NAND2_X2 U8398 ( .A1(n17972), .A2(n18935), .ZN(n13102) );
NAND2_X2 U8399 ( .A1(z_out[40]), .A2(n17960), .ZN(n13101) );
NAND2_X2 U8400 ( .A1(n13103), .A2(n13104), .ZN(n5788) );
NAND2_X2 U8401 ( .A1(n17972), .A2(n18936), .ZN(n13104) );
NAND2_X2 U8402 ( .A1(z_out[41]), .A2(n17960), .ZN(n13103) );
NAND2_X2 U8403 ( .A1(n13105), .A2(n13106), .ZN(n5787) );
NAND2_X2 U8404 ( .A1(n17972), .A2(n18937), .ZN(n13106) );
NAND2_X2 U8405 ( .A1(z_out[42]), .A2(n17960), .ZN(n13105) );
NAND2_X2 U8406 ( .A1(n13107), .A2(n13108), .ZN(n5786) );
NAND2_X2 U8407 ( .A1(n17972), .A2(n18938), .ZN(n13108) );
NAND2_X2 U8408 ( .A1(z_out[43]), .A2(n17960), .ZN(n13107) );
NAND2_X2 U8409 ( .A1(n13109), .A2(n13110), .ZN(n5785) );
NAND2_X2 U8410 ( .A1(n17972), .A2(n18939), .ZN(n13110) );
NAND2_X2 U8411 ( .A1(z_out[44]), .A2(n17960), .ZN(n13109) );
NAND2_X2 U8412 ( .A1(n13111), .A2(n13112), .ZN(n5784) );
NAND2_X2 U8413 ( .A1(n17972), .A2(n18940), .ZN(n13112) );
NAND2_X2 U8414 ( .A1(z_out[45]), .A2(n17960), .ZN(n13111) );
NAND2_X2 U8415 ( .A1(n13113), .A2(n13114), .ZN(n5783) );
NAND2_X2 U8416 ( .A1(n17972), .A2(n18941), .ZN(n13114) );
NAND2_X2 U8417 ( .A1(z_out[46]), .A2(n17960), .ZN(n13113) );
NAND2_X2 U8418 ( .A1(n13115), .A2(n13116), .ZN(n5782) );
NAND2_X2 U8419 ( .A1(n17972), .A2(n18942), .ZN(n13116) );
NAND2_X2 U8420 ( .A1(z_out[47]), .A2(n17960), .ZN(n13115) );
NAND2_X2 U8421 ( .A1(n13117), .A2(n13118), .ZN(n5781) );
NAND2_X2 U8422 ( .A1(n17972), .A2(n18943), .ZN(n13118) );
NAND2_X2 U8423 ( .A1(z_out[48]), .A2(n17960), .ZN(n13117) );
NAND2_X2 U8424 ( .A1(n13119), .A2(n13120), .ZN(n5780) );
NAND2_X2 U8425 ( .A1(n17972), .A2(n18944), .ZN(n13120) );
NAND2_X2 U8426 ( .A1(z_out[49]), .A2(n17960), .ZN(n13119) );
NAND2_X2 U8427 ( .A1(n13121), .A2(n13122), .ZN(n5779) );
NAND2_X2 U8428 ( .A1(n17972), .A2(n18945), .ZN(n13122) );
NAND2_X2 U8429 ( .A1(z_out[50]), .A2(n17960), .ZN(n13121) );
NAND2_X2 U8430 ( .A1(n13123), .A2(n13124), .ZN(n5778) );
NAND2_X2 U8431 ( .A1(n17971), .A2(n18946), .ZN(n13124) );
NAND2_X2 U8432 ( .A1(z_out[51]), .A2(n17960), .ZN(n13123) );
NAND2_X2 U8433 ( .A1(n13125), .A2(n13126), .ZN(n5777) );
NAND2_X2 U8434 ( .A1(n17971), .A2(n18947), .ZN(n13126) );
NAND2_X2 U8435 ( .A1(z_out[52]), .A2(n17960), .ZN(n13125) );
NAND2_X2 U8436 ( .A1(n13127), .A2(n13128), .ZN(n5776) );
NAND2_X2 U8437 ( .A1(n17971), .A2(n18948), .ZN(n13128) );
NAND2_X2 U8438 ( .A1(z_out[53]), .A2(n17960), .ZN(n13127) );
NAND2_X2 U8439 ( .A1(n13129), .A2(n13130), .ZN(n5775) );
NAND2_X2 U8440 ( .A1(n17971), .A2(n18949), .ZN(n13130) );
NAND2_X2 U8441 ( .A1(z_out[54]), .A2(n17960), .ZN(n13129) );
NAND2_X2 U8442 ( .A1(n13131), .A2(n13132), .ZN(n5774) );
NAND2_X2 U8443 ( .A1(n17971), .A2(n18950), .ZN(n13132) );
NAND2_X2 U8444 ( .A1(z_out[55]), .A2(n17960), .ZN(n13131) );
NAND2_X2 U8445 ( .A1(n13133), .A2(n13134), .ZN(n5773) );
NAND2_X2 U8446 ( .A1(n17971), .A2(n18951), .ZN(n13134) );
NAND2_X2 U8447 ( .A1(z_out[56]), .A2(n17961), .ZN(n13133) );
NAND2_X2 U8448 ( .A1(n13135), .A2(n13136), .ZN(n5772) );
NAND2_X2 U8449 ( .A1(n17971), .A2(n18952), .ZN(n13136) );
NAND2_X2 U8450 ( .A1(z_out[57]), .A2(n17961), .ZN(n13135) );
NAND2_X2 U8451 ( .A1(n13137), .A2(n13138), .ZN(n5771) );
NAND2_X2 U8452 ( .A1(n17971), .A2(n18953), .ZN(n13138) );
NAND2_X2 U8453 ( .A1(z_out[58]), .A2(n17961), .ZN(n13137) );
NAND2_X2 U8454 ( .A1(n13139), .A2(n13140), .ZN(n5770) );
NAND2_X2 U8455 ( .A1(n17971), .A2(n18954), .ZN(n13140) );
NAND2_X2 U8456 ( .A1(z_out[59]), .A2(n17961), .ZN(n13139) );
NAND2_X2 U8457 ( .A1(n13141), .A2(n13142), .ZN(n5769) );
NAND2_X2 U8458 ( .A1(n17971), .A2(n18955), .ZN(n13142) );
NAND2_X2 U8459 ( .A1(z_out[60]), .A2(n17961), .ZN(n13141) );
NAND2_X2 U8460 ( .A1(n13143), .A2(n13144), .ZN(n5768) );
NAND2_X2 U8461 ( .A1(n17971), .A2(n18956), .ZN(n13144) );
NAND2_X2 U8462 ( .A1(z_out[61]), .A2(n17961), .ZN(n13143) );
NAND2_X2 U8463 ( .A1(n13145), .A2(n13146), .ZN(n5767) );
NAND2_X2 U8464 ( .A1(n17970), .A2(n18957), .ZN(n13146) );
NAND2_X2 U8465 ( .A1(z_out[62]), .A2(n17961), .ZN(n13145) );
NAND2_X2 U8466 ( .A1(n13147), .A2(n13148), .ZN(n5766) );
NAND2_X2 U8467 ( .A1(n17970), .A2(n18958), .ZN(n13148) );
NAND2_X2 U8468 ( .A1(z_out[63]), .A2(n17961), .ZN(n13147) );
NAND2_X2 U8469 ( .A1(n13149), .A2(n13150), .ZN(n5765) );
NAND2_X2 U8470 ( .A1(n17970), .A2(n18959), .ZN(n13150) );
NAND2_X2 U8471 ( .A1(z_out[64]), .A2(n17961), .ZN(n13149) );
NAND2_X2 U8472 ( .A1(n13151), .A2(n13152), .ZN(n5764) );
NAND2_X2 U8473 ( .A1(n17970), .A2(n18960), .ZN(n13152) );
NAND2_X2 U8474 ( .A1(z_out[65]), .A2(n17961), .ZN(n13151) );
NAND2_X2 U8475 ( .A1(n13153), .A2(n13154), .ZN(n5763) );
NAND2_X2 U8476 ( .A1(n17970), .A2(n18961), .ZN(n13154) );
NAND2_X2 U8477 ( .A1(z_out[66]), .A2(n17961), .ZN(n13153) );
NAND2_X2 U8478 ( .A1(n13155), .A2(n13156), .ZN(n5762) );
NAND2_X2 U8479 ( .A1(n17970), .A2(n18962), .ZN(n13156) );
NAND2_X2 U8480 ( .A1(z_out[67]), .A2(n17961), .ZN(n13155) );
NAND2_X2 U8481 ( .A1(n13157), .A2(n13158), .ZN(n5761) );
NAND2_X2 U8482 ( .A1(n17970), .A2(n18963), .ZN(n13158) );
NAND2_X2 U8483 ( .A1(z_out[68]), .A2(n17961), .ZN(n13157) );
NAND2_X2 U8484 ( .A1(n13159), .A2(n13160), .ZN(n5760) );
NAND2_X2 U8485 ( .A1(n17970), .A2(n18964), .ZN(n13160) );
NAND2_X2 U8486 ( .A1(z_out[69]), .A2(n17961), .ZN(n13159) );
NAND2_X2 U8487 ( .A1(n13161), .A2(n13162), .ZN(n5759) );
NAND2_X2 U8488 ( .A1(n17970), .A2(n18965), .ZN(n13162) );
NAND2_X2 U8489 ( .A1(z_out[70]), .A2(n17961), .ZN(n13161) );
NAND2_X2 U8490 ( .A1(n13163), .A2(n13164), .ZN(n5758) );
NAND2_X2 U8491 ( .A1(n17970), .A2(n18966), .ZN(n13164) );
NAND2_X2 U8492 ( .A1(z_out[71]), .A2(n17961), .ZN(n13163) );
NAND2_X2 U8493 ( .A1(n13165), .A2(n13166), .ZN(n5757) );
NAND2_X2 U8494 ( .A1(n17970), .A2(n18967), .ZN(n13166) );
NAND2_X2 U8495 ( .A1(z_out[72]), .A2(n17961), .ZN(n13165) );
NAND2_X2 U8496 ( .A1(n13167), .A2(n13168), .ZN(n5756) );
NAND2_X2 U8497 ( .A1(n17969), .A2(n18968), .ZN(n13168) );
NAND2_X2 U8498 ( .A1(z_out[73]), .A2(n17961), .ZN(n13167) );
NAND2_X2 U8499 ( .A1(n13169), .A2(n13170), .ZN(n5755) );
NAND2_X2 U8500 ( .A1(n17969), .A2(n18969), .ZN(n13170) );
NAND2_X2 U8501 ( .A1(z_out[74]), .A2(n17962), .ZN(n13169) );
NAND2_X2 U8502 ( .A1(n13171), .A2(n13172), .ZN(n5754) );
NAND2_X2 U8503 ( .A1(n17969), .A2(n18970), .ZN(n13172) );
NAND2_X2 U8504 ( .A1(z_out[75]), .A2(n17962), .ZN(n13171) );
NAND2_X2 U8505 ( .A1(n13173), .A2(n13174), .ZN(n5753) );
NAND2_X2 U8506 ( .A1(n17969), .A2(n18971), .ZN(n13174) );
NAND2_X2 U8507 ( .A1(z_out[76]), .A2(n17962), .ZN(n13173) );
NAND2_X2 U8508 ( .A1(n13175), .A2(n13176), .ZN(n5752) );
NAND2_X2 U8509 ( .A1(n17969), .A2(n18972), .ZN(n13176) );
NAND2_X2 U8510 ( .A1(z_out[77]), .A2(n17962), .ZN(n13175) );
NAND2_X2 U8511 ( .A1(n13177), .A2(n13178), .ZN(n5751) );
NAND2_X2 U8512 ( .A1(n17969), .A2(n18973), .ZN(n13178) );
NAND2_X2 U8513 ( .A1(z_out[78]), .A2(n17962), .ZN(n13177) );
NAND2_X2 U8514 ( .A1(n13179), .A2(n13180), .ZN(n5750) );
NAND2_X2 U8515 ( .A1(n17969), .A2(n18974), .ZN(n13180) );
NAND2_X2 U8516 ( .A1(z_out[79]), .A2(n17962), .ZN(n13179) );
NAND2_X2 U8517 ( .A1(n13181), .A2(n13182), .ZN(n5749) );
NAND2_X2 U8518 ( .A1(n17969), .A2(n18975), .ZN(n13182) );
NAND2_X2 U8519 ( .A1(z_out[80]), .A2(n17962), .ZN(n13181) );
NAND2_X2 U8520 ( .A1(n13183), .A2(n13184), .ZN(n5748) );
NAND2_X2 U8521 ( .A1(n17969), .A2(n18976), .ZN(n13184) );
NAND2_X2 U8522 ( .A1(z_out[81]), .A2(n17962), .ZN(n13183) );
NAND2_X2 U8523 ( .A1(n13185), .A2(n13186), .ZN(n5747) );
NAND2_X2 U8524 ( .A1(n17969), .A2(n18977), .ZN(n13186) );
NAND2_X2 U8525 ( .A1(z_out[82]), .A2(n17962), .ZN(n13185) );
NAND2_X2 U8526 ( .A1(n13187), .A2(n13188), .ZN(n5746) );
NAND2_X2 U8527 ( .A1(n17969), .A2(n18978), .ZN(n13188) );
NAND2_X2 U8528 ( .A1(z_out[83]), .A2(n17962), .ZN(n13187) );
NAND2_X2 U8529 ( .A1(n13189), .A2(n13190), .ZN(n5745) );
NAND2_X2 U8530 ( .A1(n17968), .A2(n18979), .ZN(n13190) );
NAND2_X2 U8531 ( .A1(z_out[84]), .A2(n17962), .ZN(n13189) );
NAND2_X2 U8532 ( .A1(n13191), .A2(n13192), .ZN(n5744) );
NAND2_X2 U8533 ( .A1(n17968), .A2(n18980), .ZN(n13192) );
NAND2_X2 U8534 ( .A1(z_out[85]), .A2(n17962), .ZN(n13191) );
NAND2_X2 U8535 ( .A1(n13193), .A2(n13194), .ZN(n5743) );
NAND2_X2 U8536 ( .A1(n17968), .A2(n18981), .ZN(n13194) );
NAND2_X2 U8537 ( .A1(z_out[86]), .A2(n17962), .ZN(n13193) );
NAND2_X2 U8538 ( .A1(n13195), .A2(n13196), .ZN(n5742) );
NAND2_X2 U8539 ( .A1(n17968), .A2(n18982), .ZN(n13196) );
NAND2_X2 U8540 ( .A1(z_out[87]), .A2(n17962), .ZN(n13195) );
NAND2_X2 U8541 ( .A1(n13197), .A2(n13198), .ZN(n5741) );
NAND2_X2 U8542 ( .A1(n17968), .A2(n18983), .ZN(n13198) );
NAND2_X2 U8543 ( .A1(z_out[88]), .A2(n17962), .ZN(n13197) );
NAND2_X2 U8544 ( .A1(n13199), .A2(n13200), .ZN(n5740) );
NAND2_X2 U8545 ( .A1(n17968), .A2(n18984), .ZN(n13200) );
NAND2_X2 U8546 ( .A1(z_out[89]), .A2(n17962), .ZN(n13199) );
NAND2_X2 U8547 ( .A1(n13201), .A2(n13202), .ZN(n5739) );
NAND2_X2 U8548 ( .A1(n17968), .A2(n18985), .ZN(n13202) );
NAND2_X2 U8549 ( .A1(z_out[90]), .A2(n17962), .ZN(n13201) );
NAND2_X2 U8550 ( .A1(n13203), .A2(n13204), .ZN(n5738) );
NAND2_X2 U8551 ( .A1(n17968), .A2(n18986), .ZN(n13204) );
NAND2_X2 U8552 ( .A1(z_out[91]), .A2(n17962), .ZN(n13203) );
NAND2_X2 U8553 ( .A1(n13205), .A2(n13206), .ZN(n5737) );
NAND2_X2 U8554 ( .A1(n17968), .A2(n18987), .ZN(n13206) );
NAND2_X2 U8555 ( .A1(z_out[92]), .A2(n17962), .ZN(n13205) );
NAND2_X2 U8556 ( .A1(n13207), .A2(n13208), .ZN(n5736) );
NAND2_X2 U8557 ( .A1(n17968), .A2(n18988), .ZN(n13208) );
NAND2_X2 U8558 ( .A1(z_out[93]), .A2(n17963), .ZN(n13207) );
NAND2_X2 U8559 ( .A1(n13209), .A2(n13210), .ZN(n5735) );
NAND2_X2 U8560 ( .A1(n17968), .A2(n18989), .ZN(n13210) );
NAND2_X2 U8561 ( .A1(z_out[94]), .A2(n17963), .ZN(n13209) );
NAND2_X2 U8562 ( .A1(n13211), .A2(n13212), .ZN(n5734) );
NAND2_X2 U8563 ( .A1(n17967), .A2(n18990), .ZN(n13212) );
NAND2_X2 U8564 ( .A1(z_out[95]), .A2(n17963), .ZN(n13211) );
NAND2_X2 U8565 ( .A1(n13213), .A2(n13214), .ZN(n5733) );
NAND2_X2 U8566 ( .A1(n17967), .A2(n18991), .ZN(n13214) );
NAND2_X2 U8567 ( .A1(z_out[96]), .A2(n17963), .ZN(n13213) );
NAND2_X2 U8568 ( .A1(n13215), .A2(n13216), .ZN(n5732) );
NAND2_X2 U8569 ( .A1(n17967), .A2(n18992), .ZN(n13216) );
NAND2_X2 U8570 ( .A1(z_out[97]), .A2(n17963), .ZN(n13215) );
NAND2_X2 U8571 ( .A1(n13217), .A2(n13218), .ZN(n5731) );
NAND2_X2 U8572 ( .A1(n17967), .A2(n18993), .ZN(n13218) );
NAND2_X2 U8573 ( .A1(z_out[98]), .A2(n17963), .ZN(n13217) );
NAND2_X2 U8574 ( .A1(n13219), .A2(n13220), .ZN(n5730) );
NAND2_X2 U8575 ( .A1(n17967), .A2(n18994), .ZN(n13220) );
NAND2_X2 U8576 ( .A1(z_out[99]), .A2(n17963), .ZN(n13219) );
NAND2_X2 U8577 ( .A1(n13221), .A2(n13222), .ZN(n5729) );
NAND2_X2 U8578 ( .A1(n17967), .A2(n18995), .ZN(n13222) );
NAND2_X2 U8579 ( .A1(z_out[100]), .A2(n17963), .ZN(n13221) );
NAND2_X2 U8580 ( .A1(n13223), .A2(n13224), .ZN(n5728) );
NAND2_X2 U8581 ( .A1(n17967), .A2(n18996), .ZN(n13224) );
NAND2_X2 U8582 ( .A1(z_out[101]), .A2(n17963), .ZN(n13223) );
NAND2_X2 U8583 ( .A1(n13225), .A2(n13226), .ZN(n5727) );
NAND2_X2 U8584 ( .A1(n17967), .A2(n18997), .ZN(n13226) );
NAND2_X2 U8585 ( .A1(z_out[102]), .A2(n17963), .ZN(n13225) );
NAND2_X2 U8586 ( .A1(n13227), .A2(n13228), .ZN(n5726) );
NAND2_X2 U8587 ( .A1(n17967), .A2(n18998), .ZN(n13228) );
NAND2_X2 U8588 ( .A1(z_out[103]), .A2(n17963), .ZN(n13227) );
NAND2_X2 U8589 ( .A1(n13229), .A2(n13230), .ZN(n5725) );
NAND2_X2 U8590 ( .A1(n17967), .A2(n18999), .ZN(n13230) );
NAND2_X2 U8591 ( .A1(z_out[104]), .A2(n17963), .ZN(n13229) );
NAND2_X2 U8592 ( .A1(n13231), .A2(n13232), .ZN(n5724) );
NAND2_X2 U8593 ( .A1(n17967), .A2(n19000), .ZN(n13232) );
NAND2_X2 U8594 ( .A1(z_out[105]), .A2(n17963), .ZN(n13231) );
NAND2_X2 U8595 ( .A1(n13233), .A2(n13234), .ZN(n5723) );
NAND2_X2 U8596 ( .A1(n17966), .A2(n19001), .ZN(n13234) );
NAND2_X2 U8597 ( .A1(z_out[106]), .A2(n17963), .ZN(n13233) );
NAND2_X2 U8598 ( .A1(n13235), .A2(n13236), .ZN(n5722) );
NAND2_X2 U8599 ( .A1(n17966), .A2(n19002), .ZN(n13236) );
NAND2_X2 U8600 ( .A1(z_out[107]), .A2(n17963), .ZN(n13235) );
NAND2_X2 U8601 ( .A1(n13237), .A2(n13238), .ZN(n5721) );
NAND2_X2 U8602 ( .A1(n17966), .A2(n19003), .ZN(n13238) );
NAND2_X2 U8603 ( .A1(z_out[108]), .A2(n17963), .ZN(n13237) );
NAND2_X2 U8604 ( .A1(n13239), .A2(n13240), .ZN(n5720) );
NAND2_X2 U8605 ( .A1(n17966), .A2(n19004), .ZN(n13240) );
NAND2_X2 U8606 ( .A1(z_out[109]), .A2(n17963), .ZN(n13239) );
NAND2_X2 U8607 ( .A1(n13241), .A2(n13242), .ZN(n5719) );
NAND2_X2 U8608 ( .A1(n17966), .A2(n19005), .ZN(n13242) );
NAND2_X2 U8609 ( .A1(z_out[110]), .A2(n17963), .ZN(n13241) );
NAND2_X2 U8610 ( .A1(n13243), .A2(n13244), .ZN(n5718) );
NAND2_X2 U8611 ( .A1(n17966), .A2(n19006), .ZN(n13244) );
NAND2_X2 U8612 ( .A1(z_out[111]), .A2(n17963), .ZN(n13243) );
NAND2_X2 U8613 ( .A1(n13245), .A2(n13246), .ZN(n5717) );
NAND2_X2 U8614 ( .A1(n17966), .A2(n19007), .ZN(n13246) );
NAND2_X2 U8615 ( .A1(z_out[112]), .A2(n17964), .ZN(n13245) );
NAND2_X2 U8616 ( .A1(n13247), .A2(n13248), .ZN(n5716) );
NAND2_X2 U8617 ( .A1(n17966), .A2(n19008), .ZN(n13248) );
NAND2_X2 U8618 ( .A1(z_out[113]), .A2(n17964), .ZN(n13247) );
NAND2_X2 U8619 ( .A1(n13249), .A2(n13250), .ZN(n5715) );
NAND2_X2 U8620 ( .A1(n17966), .A2(n19009), .ZN(n13250) );
NAND2_X2 U8621 ( .A1(z_out[114]), .A2(n17964), .ZN(n13249) );
NAND2_X2 U8622 ( .A1(n13251), .A2(n13252), .ZN(n5714) );
NAND2_X2 U8623 ( .A1(n17966), .A2(n19010), .ZN(n13252) );
NAND2_X2 U8624 ( .A1(z_out[115]), .A2(n17964), .ZN(n13251) );
NAND2_X2 U8625 ( .A1(n13253), .A2(n13254), .ZN(n5713) );
NAND2_X2 U8626 ( .A1(n17966), .A2(n19011), .ZN(n13254) );
NAND2_X2 U8627 ( .A1(z_out[116]), .A2(n17964), .ZN(n13253) );
NAND2_X2 U8628 ( .A1(n13255), .A2(n13256), .ZN(n5712) );
NAND2_X2 U8629 ( .A1(n17965), .A2(n19012), .ZN(n13256) );
NAND2_X2 U8630 ( .A1(z_out[117]), .A2(n17964), .ZN(n13255) );
NAND2_X2 U8631 ( .A1(n13257), .A2(n13258), .ZN(n5711) );
NAND2_X2 U8632 ( .A1(n17965), .A2(n19013), .ZN(n13258) );
NAND2_X2 U8633 ( .A1(z_out[118]), .A2(n17964), .ZN(n13257) );
NAND2_X2 U8634 ( .A1(n13259), .A2(n13260), .ZN(n5710) );
NAND2_X2 U8635 ( .A1(n17965), .A2(n19014), .ZN(n13260) );
NAND2_X2 U8636 ( .A1(z_out[119]), .A2(n17964), .ZN(n13259) );
NAND2_X2 U8637 ( .A1(n13261), .A2(n13262), .ZN(n5709) );
NAND2_X2 U8638 ( .A1(n17965), .A2(n19015), .ZN(n13262) );
NAND2_X2 U8639 ( .A1(z_out[120]), .A2(n17964), .ZN(n13261) );
NAND2_X2 U8640 ( .A1(n13263), .A2(n13264), .ZN(n5708) );
NAND2_X2 U8641 ( .A1(n17965), .A2(n19016), .ZN(n13264) );
NAND2_X2 U8642 ( .A1(z_out[121]), .A2(n17964), .ZN(n13263) );
NAND2_X2 U8643 ( .A1(n13265), .A2(n13266), .ZN(n5707) );
NAND2_X2 U8644 ( .A1(n17965), .A2(n19017), .ZN(n13266) );
NAND2_X2 U8645 ( .A1(z_out[122]), .A2(n17964), .ZN(n13265) );
NAND2_X2 U8646 ( .A1(n13267), .A2(n13268), .ZN(n5706) );
NAND2_X2 U8647 ( .A1(n17965), .A2(n19018), .ZN(n13268) );
NAND2_X2 U8648 ( .A1(z_out[123]), .A2(n17964), .ZN(n13267) );
NAND2_X2 U8649 ( .A1(n13269), .A2(n13270), .ZN(n5705) );
NAND2_X2 U8650 ( .A1(n17965), .A2(n19019), .ZN(n13270) );
NAND2_X2 U8651 ( .A1(z_out[124]), .A2(n17964), .ZN(n13269) );
NAND2_X2 U8652 ( .A1(n13271), .A2(n13272), .ZN(n5704) );
NAND2_X2 U8653 ( .A1(n17965), .A2(n19020), .ZN(n13272) );
NAND2_X2 U8654 ( .A1(z_out[125]), .A2(n17964), .ZN(n13271) );
NAND2_X2 U8655 ( .A1(n13273), .A2(n13274), .ZN(n5703) );
NAND2_X2 U8656 ( .A1(n17965), .A2(n19021), .ZN(n13274) );
NAND2_X2 U8657 ( .A1(z_out[126]), .A2(n17964), .ZN(n13273) );
NAND2_X2 U8658 ( .A1(n13275), .A2(n13276), .ZN(n5702) );
NAND2_X2 U8659 ( .A1(n17965), .A2(n19022), .ZN(n13276) );
NAND2_X2 U8661 ( .A1(z_out[127]), .A2(n17958), .ZN(n13275) );
NAND4_X2 U8663 ( .A1(n13277), .A2(n13278), .A3(n13279), .A4(n13280), .ZN(n5701) );
NAND2_X2 U8664 ( .A1(n13281), .A2(n17847), .ZN(n13279) );
XNOR2_X2 U8665 ( .A(n17279), .B(z_out[0]), .ZN(n13281) );
NAND2_X2 U8666 ( .A1(n17957), .A2(Out_data[0]), .ZN(n13278) );
NAND2_X2 U8667 ( .A1(n17935), .A2(aes_text_out[0]), .ZN(n13277) );
NAND4_X2 U8668 ( .A1(n13284), .A2(n13285), .A3(n13286), .A4(n13287), .ZN(n5700) );
NAND2_X2 U8669 ( .A1(n13288), .A2(n17847), .ZN(n13286) );
XNOR2_X2 U8670 ( .A(n17277), .B(z_out[1]), .ZN(n13288) );
NAND2_X2 U8671 ( .A1(n17957), .A2(Out_data[1]), .ZN(n13285) );
NAND2_X2 U8672 ( .A1(n17933), .A2(aes_text_out[1]), .ZN(n13284) );
NAND4_X2 U8673 ( .A1(n13289), .A2(n13290), .A3(n13291), .A4(n13292), .ZN(n5699) );
NAND2_X2 U8674 ( .A1(n13293), .A2(n17847), .ZN(n13291) );
XNOR2_X2 U8675 ( .A(n17275), .B(z_out[2]), .ZN(n13293) );
NAND2_X2 U8676 ( .A1(n17957), .A2(Out_data[2]), .ZN(n13290) );
NAND2_X2 U8677 ( .A1(n17934), .A2(aes_text_out[2]), .ZN(n13289) );
NAND4_X2 U8678 ( .A1(n13294), .A2(n13295), .A3(n13296), .A4(n13297), .ZN(n5698) );
NAND2_X2 U8679 ( .A1(n13298), .A2(n17847), .ZN(n13296) );
XNOR2_X2 U8680 ( .A(n17273), .B(z_out[3]), .ZN(n13298) );
NAND2_X2 U8681 ( .A1(n17957), .A2(Out_data[3]), .ZN(n13295) );
NAND2_X2 U8682 ( .A1(n17933), .A2(aes_text_out[3]), .ZN(n13294) );
NAND4_X2 U8683 ( .A1(n13299), .A2(n13300), .A3(n13301), .A4(n13302), .ZN(n5697) );
NAND2_X2 U8684 ( .A1(n13303), .A2(n17847), .ZN(n13301) );
XNOR2_X2 U8685 ( .A(n17271), .B(z_out[4]), .ZN(n13303) );
NAND2_X2 U8686 ( .A1(n17957), .A2(Out_data[4]), .ZN(n13300) );
NAND2_X2 U8687 ( .A1(n17934), .A2(aes_text_out[4]), .ZN(n13299) );
NAND4_X2 U8688 ( .A1(n13304), .A2(n13305), .A3(n13306), .A4(n13307), .ZN(n5696) );
NAND2_X2 U8689 ( .A1(n13308), .A2(n17847), .ZN(n13306) );
XNOR2_X2 U8690 ( .A(n17269), .B(z_out[5]), .ZN(n13308) );
NAND2_X2 U8691 ( .A1(n17957), .A2(Out_data[5]), .ZN(n13305) );
NAND2_X2 U8692 ( .A1(n17934), .A2(aes_text_out[5]), .ZN(n13304) );
NAND4_X2 U8693 ( .A1(n13309), .A2(n13310), .A3(n13311), .A4(n13312), .ZN(n5695) );
NAND2_X2 U8694 ( .A1(n13313), .A2(n17847), .ZN(n13311) );
XNOR2_X2 U8695 ( .A(n17267), .B(z_out[6]), .ZN(n13313) );
NAND2_X2 U8696 ( .A1(n17957), .A2(Out_data[6]), .ZN(n13310) );
NAND2_X2 U8697 ( .A1(n17935), .A2(aes_text_out[6]), .ZN(n13309) );
NAND4_X2 U8698 ( .A1(n13314), .A2(n13315), .A3(n13316), .A4(n13317), .ZN(n5694) );
NAND2_X2 U8699 ( .A1(n13318), .A2(n17847), .ZN(n13316) );
XNOR2_X2 U8700 ( .A(n17265), .B(z_out[7]), .ZN(n13318) );
NAND2_X2 U8701 ( .A1(n17956), .A2(Out_data[7]), .ZN(n13315) );
NAND2_X2 U8702 ( .A1(n17935), .A2(aes_text_out[7]), .ZN(n13314) );
NAND4_X2 U8703 ( .A1(n13319), .A2(n13320), .A3(n13321), .A4(n13322), .ZN(n5693) );
NAND2_X2 U8704 ( .A1(aes_text_out[8]), .A2(n13323), .ZN(n13321) );
NAND2_X2 U8705 ( .A1(n13324), .A2(n17847), .ZN(n13320) );
XNOR2_X2 U8706 ( .A(n17263), .B(z_out[8]), .ZN(n13324) );
NAND2_X2 U8707 ( .A1(n17956), .A2(Out_data[8]), .ZN(n13319) );
NAND4_X2 U8708 ( .A1(n13325), .A2(n13326), .A3(n13327), .A4(n13328), .ZN(n5692) );
NAND2_X2 U8709 ( .A1(aes_text_out[9]), .A2(n13329), .ZN(n13327) );
NAND2_X2 U8710 ( .A1(n13330), .A2(n17847), .ZN(n13326) );
XNOR2_X2 U8711 ( .A(n17261), .B(z_out[9]), .ZN(n13330) );
NAND2_X2 U8712 ( .A1(n17956), .A2(Out_data[9]), .ZN(n13325) );
NAND4_X2 U8713 ( .A1(n13331), .A2(n13332), .A3(n13333), .A4(n13334), .ZN(n5691) );
NAND2_X2 U8714 ( .A1(aes_text_out[10]), .A2(n13335), .ZN(n13333) );
NAND2_X2 U8715 ( .A1(n13336), .A2(n17847), .ZN(n13332) );
XNOR2_X2 U8716 ( .A(n17259), .B(z_out[10]), .ZN(n13336) );
NAND2_X2 U8717 ( .A1(n17956), .A2(Out_data[10]), .ZN(n13331) );
NAND4_X2 U8718 ( .A1(n13337), .A2(n13338), .A3(n13339), .A4(n13340), .ZN(n5690) );
NAND2_X2 U8719 ( .A1(aes_text_out[11]), .A2(n13341), .ZN(n13339) );
NAND2_X2 U8720 ( .A1(n13342), .A2(n17847), .ZN(n13338) );
XNOR2_X2 U8721 ( .A(n17257), .B(z_out[11]), .ZN(n13342) );
NAND2_X2 U8722 ( .A1(n17956), .A2(Out_data[11]), .ZN(n13337) );
NAND4_X2 U8723 ( .A1(n13343), .A2(n13344), .A3(n13345), .A4(n13346), .ZN(n5689) );
NAND2_X2 U8724 ( .A1(aes_text_out[12]), .A2(n13347), .ZN(n13345) );
NAND2_X2 U8725 ( .A1(n13348), .A2(n17847), .ZN(n13344) );
XNOR2_X2 U8726 ( .A(n17255), .B(z_out[12]), .ZN(n13348) );
NAND2_X2 U8727 ( .A1(n17956), .A2(Out_data[12]), .ZN(n13343) );
NAND4_X2 U8728 ( .A1(n13349), .A2(n13350), .A3(n13351), .A4(n13352), .ZN(n5688) );
NAND2_X2 U8729 ( .A1(aes_text_out[13]), .A2(n13353), .ZN(n13351) );
NAND2_X2 U8730 ( .A1(n13354), .A2(n17847), .ZN(n13350) );
XNOR2_X2 U8731 ( .A(n17253), .B(z_out[13]), .ZN(n13354) );
NAND2_X2 U8732 ( .A1(n17956), .A2(Out_data[13]), .ZN(n13349) );
NAND4_X2 U8733 ( .A1(n13355), .A2(n13356), .A3(n13357), .A4(n13358), .ZN(n5687) );
NAND2_X2 U8734 ( .A1(aes_text_out[14]), .A2(n13359), .ZN(n13357) );
NAND2_X2 U8735 ( .A1(n13360), .A2(n17847), .ZN(n13356) );
XNOR2_X2 U8736 ( .A(n17251), .B(z_out[14]), .ZN(n13360) );
NAND2_X2 U8737 ( .A1(n17956), .A2(Out_data[14]), .ZN(n13355) );
NAND4_X2 U8738 ( .A1(n13361), .A2(n13362), .A3(n13363), .A4(n13364), .ZN(n5686) );
NAND2_X2 U8739 ( .A1(aes_text_out[15]), .A2(n13365), .ZN(n13363) );
NAND2_X2 U8740 ( .A1(n13366), .A2(n17846), .ZN(n13362) );
XNOR2_X2 U8741 ( .A(n17249), .B(z_out[15]), .ZN(n13366) );
NAND2_X2 U8742 ( .A1(n17956), .A2(Out_data[15]), .ZN(n13361) );
NAND4_X2 U8743 ( .A1(n13367), .A2(n13368), .A3(n13369), .A4(n13370), .ZN(n5685) );
NAND2_X2 U8744 ( .A1(n13371), .A2(n17846), .ZN(n13369) );
XNOR2_X2 U8745 ( .A(n17247), .B(z_out[16]), .ZN(n13371) );
NAND2_X2 U8746 ( .A1(n17956), .A2(Out_data[16]), .ZN(n13368) );
NAND2_X2 U8747 ( .A1(n13372), .A2(n17936), .ZN(n13367) );
NAND4_X2 U8748 ( .A1(n13373), .A2(n13374), .A3(n13375), .A4(n13376), .ZN(n5684) );
NAND2_X2 U8749 ( .A1(n13377), .A2(n17846), .ZN(n13375) );
XNOR2_X2 U8750 ( .A(n17245), .B(z_out[17]), .ZN(n13377) );
NAND2_X2 U8751 ( .A1(n17956), .A2(Out_data[17]), .ZN(n13374) );
NAND2_X2 U8752 ( .A1(n13378), .A2(n17936), .ZN(n13373) );
NAND4_X2 U8753 ( .A1(n13379), .A2(n13380), .A3(n13381), .A4(n13382), .ZN(n5683) );
NAND2_X2 U8754 ( .A1(n13383), .A2(n17846), .ZN(n13381) );
XNOR2_X2 U8755 ( .A(n17243), .B(z_out[18]), .ZN(n13383) );
NAND2_X2 U8756 ( .A1(n17955), .A2(Out_data[18]), .ZN(n13380) );
NAND2_X2 U8757 ( .A1(n13384), .A2(n17936), .ZN(n13379) );
NAND4_X2 U8758 ( .A1(n13385), .A2(n13386), .A3(n13387), .A4(n13388), .ZN(n5682) );
NAND2_X2 U8759 ( .A1(n13389), .A2(n17846), .ZN(n13387) );
XNOR2_X2 U8760 ( .A(n17241), .B(z_out[19]), .ZN(n13389) );
NAND2_X2 U8761 ( .A1(n17955), .A2(Out_data[19]), .ZN(n13386) );
NAND2_X2 U8762 ( .A1(n13390), .A2(n17936), .ZN(n13385) );
NAND4_X2 U8763 ( .A1(n13391), .A2(n13392), .A3(n13393), .A4(n13394), .ZN(n5681) );
NAND2_X2 U8764 ( .A1(n13395), .A2(n17846), .ZN(n13393) );
XNOR2_X2 U8765 ( .A(n17239), .B(z_out[20]), .ZN(n13395) );
NAND2_X2 U8766 ( .A1(n17955), .A2(Out_data[20]), .ZN(n13392) );
NAND2_X2 U8767 ( .A1(n13396), .A2(n17936), .ZN(n13391) );
NAND4_X2 U8768 ( .A1(n13397), .A2(n13398), .A3(n13399), .A4(n13400), .ZN(n5680) );
NAND2_X2 U8769 ( .A1(n13401), .A2(n17846), .ZN(n13399) );
XNOR2_X2 U8770 ( .A(n17237), .B(z_out[21]), .ZN(n13401) );
NAND2_X2 U8771 ( .A1(n17955), .A2(Out_data[21]), .ZN(n13398) );
NAND2_X2 U8772 ( .A1(n13402), .A2(n17936), .ZN(n13397) );
NAND4_X2 U8773 ( .A1(n13403), .A2(n13404), .A3(n13405), .A4(n13406), .ZN(n5679) );
NAND2_X2 U8774 ( .A1(n13407), .A2(n17846), .ZN(n13405) );
XNOR2_X2 U8775 ( .A(n17235), .B(z_out[22]), .ZN(n13407) );
NAND2_X2 U8776 ( .A1(n17955), .A2(Out_data[22]), .ZN(n13404) );
NAND2_X2 U8777 ( .A1(n13408), .A2(n17936), .ZN(n13403) );
NAND4_X2 U8778 ( .A1(n13409), .A2(n13410), .A3(n13411), .A4(n13412), .ZN(n5678) );
NAND2_X2 U8779 ( .A1(n13413), .A2(n17846), .ZN(n13411) );
XNOR2_X2 U8780 ( .A(n17233), .B(z_out[23]), .ZN(n13413) );
NAND2_X2 U8781 ( .A1(n17955), .A2(Out_data[23]), .ZN(n13410) );
NAND2_X2 U8782 ( .A1(n13414), .A2(n17936), .ZN(n13409) );
NAND4_X2 U8783 ( .A1(n13415), .A2(n13416), .A3(n13417), .A4(n13418), .ZN(n5677) );
NAND2_X2 U8784 ( .A1(n13419), .A2(n17846), .ZN(n13417) );
XNOR2_X2 U8785 ( .A(n17231), .B(z_out[24]), .ZN(n13419) );
NAND2_X2 U8786 ( .A1(n17955), .A2(Out_data[24]), .ZN(n13416) );
NAND2_X2 U8787 ( .A1(n18835), .A2(n17936), .ZN(n13415) );
NAND4_X2 U8788 ( .A1(n13421), .A2(n13422), .A3(n13423), .A4(n13424), .ZN(n5676) );
NAND2_X2 U8789 ( .A1(n13425), .A2(n17846), .ZN(n13423) );
XNOR2_X2 U8790 ( .A(n17229), .B(z_out[25]), .ZN(n13425) );
NAND2_X2 U8791 ( .A1(n17955), .A2(Out_data[25]), .ZN(n13422) );
NAND2_X2 U8792 ( .A1(n18834), .A2(n17936), .ZN(n13421) );
NAND4_X2 U8793 ( .A1(n13427), .A2(n13428), .A3(n13429), .A4(n13430), .ZN(n5675) );
NAND2_X2 U8794 ( .A1(n13431), .A2(n17846), .ZN(n13429) );
XNOR2_X2 U8795 ( .A(n17227), .B(z_out[26]), .ZN(n13431) );
NAND2_X2 U8796 ( .A1(n17955), .A2(Out_data[26]), .ZN(n13428) );
NAND2_X2 U8797 ( .A1(n18833), .A2(n17936), .ZN(n13427) );
NAND4_X2 U8798 ( .A1(n13433), .A2(n13434), .A3(n13435), .A4(n13436), .ZN(n5674) );
NAND2_X2 U8799 ( .A1(n13437), .A2(n17846), .ZN(n13435) );
XNOR2_X2 U8800 ( .A(n17225), .B(z_out[27]), .ZN(n13437) );
NAND2_X2 U8801 ( .A1(n17955), .A2(Out_data[27]), .ZN(n13434) );
NAND2_X2 U8802 ( .A1(n18832), .A2(n17937), .ZN(n13433) );
NAND4_X2 U8803 ( .A1(n13439), .A2(n13440), .A3(n13441), .A4(n13442), .ZN(n5673) );
NAND2_X2 U8804 ( .A1(n13443), .A2(n17846), .ZN(n13441) );
XNOR2_X2 U8805 ( .A(n17223), .B(z_out[28]), .ZN(n13443) );
NAND2_X2 U8806 ( .A1(n17955), .A2(Out_data[28]), .ZN(n13440) );
NAND2_X2 U8807 ( .A1(n18831), .A2(n17937), .ZN(n13439) );
NAND4_X2 U8808 ( .A1(n13445), .A2(n13446), .A3(n13447), .A4(n13448), .ZN(n5672) );
NAND2_X2 U8809 ( .A1(n13449), .A2(n17846), .ZN(n13447) );
XNOR2_X2 U8810 ( .A(n17221), .B(z_out[29]), .ZN(n13449) );
NAND2_X2 U8811 ( .A1(n17954), .A2(Out_data[29]), .ZN(n13446) );
NAND2_X2 U8812 ( .A1(n18830), .A2(n17937), .ZN(n13445) );
NAND4_X2 U8813 ( .A1(n13451), .A2(n13452), .A3(n13453), .A4(n13454), .ZN(n5671) );
NAND2_X2 U8814 ( .A1(n13455), .A2(n17846), .ZN(n13453) );
XNOR2_X2 U8815 ( .A(n17219), .B(z_out[30]), .ZN(n13455) );
NAND2_X2 U8816 ( .A1(n17954), .A2(Out_data[30]), .ZN(n13452) );
NAND2_X2 U8817 ( .A1(n18829), .A2(n17937), .ZN(n13451) );
NAND4_X2 U8818 ( .A1(n13457), .A2(n13458), .A3(n13459), .A4(n13460), .ZN(n5670) );
NAND2_X2 U8819 ( .A1(n13461), .A2(n17846), .ZN(n13459) );
XNOR2_X2 U8820 ( .A(n17217), .B(z_out[31]), .ZN(n13461) );
NAND2_X2 U8821 ( .A1(n17954), .A2(Out_data[31]), .ZN(n13458) );
NAND2_X2 U8822 ( .A1(n18828), .A2(n17937), .ZN(n13457) );
NAND4_X2 U8823 ( .A1(n13463), .A2(n13464), .A3(n13465), .A4(n13466), .ZN(n5669) );
NAND2_X2 U8824 ( .A1(n13467), .A2(n17846), .ZN(n13465) );
XNOR2_X2 U8825 ( .A(n17215), .B(z_out[32]), .ZN(n13467) );
NAND2_X2 U8826 ( .A1(n17954), .A2(Out_data[32]), .ZN(n13464) );
NAND2_X2 U8827 ( .A1(n13468), .A2(n17937), .ZN(n13463) );
NAND4_X2 U8828 ( .A1(n13469), .A2(n13470), .A3(n13471), .A4(n13472), .ZN(n5668) );
NAND2_X2 U8829 ( .A1(n13473), .A2(n17846), .ZN(n13471) );
XNOR2_X2 U8830 ( .A(n17213), .B(z_out[33]), .ZN(n13473) );
NAND2_X2 U8831 ( .A1(n17954), .A2(Out_data[33]), .ZN(n13470) );
NAND2_X2 U8832 ( .A1(n13474), .A2(n17937), .ZN(n13469) );
NAND4_X2 U8833 ( .A1(n13475), .A2(n13476), .A3(n13477), .A4(n13478), .ZN(n5667) );
NAND2_X2 U8834 ( .A1(n13479), .A2(n17845), .ZN(n13477) );
XNOR2_X2 U8835 ( .A(n17211), .B(z_out[34]), .ZN(n13479) );
NAND2_X2 U8836 ( .A1(n17954), .A2(Out_data[34]), .ZN(n13476) );
NAND2_X2 U8837 ( .A1(n13480), .A2(n17937), .ZN(n13475) );
NAND4_X2 U8838 ( .A1(n13481), .A2(n13482), .A3(n13483), .A4(n13484), .ZN(n5666) );
NAND2_X2 U8839 ( .A1(n13485), .A2(n17845), .ZN(n13483) );
XNOR2_X2 U8840 ( .A(n17209), .B(z_out[35]), .ZN(n13485) );
NAND2_X2 U8841 ( .A1(n17954), .A2(Out_data[35]), .ZN(n13482) );
NAND2_X2 U8842 ( .A1(n13486), .A2(n17937), .ZN(n13481) );
NAND4_X2 U8843 ( .A1(n13487), .A2(n13488), .A3(n13489), .A4(n13490), .ZN(n5665) );
NAND2_X2 U8844 ( .A1(n13491), .A2(n17845), .ZN(n13489) );
XNOR2_X2 U8845 ( .A(n17207), .B(z_out[36]), .ZN(n13491) );
NAND2_X2 U8846 ( .A1(n17954), .A2(Out_data[36]), .ZN(n13488) );
NAND2_X2 U8847 ( .A1(n13492), .A2(n17937), .ZN(n13487) );
NAND4_X2 U8848 ( .A1(n13493), .A2(n13494), .A3(n13495), .A4(n13496), .ZN(n5664) );
NAND2_X2 U8849 ( .A1(n13497), .A2(n17845), .ZN(n13495) );
XNOR2_X2 U8850 ( .A(n17205), .B(z_out[37]), .ZN(n13497) );
NAND2_X2 U8851 ( .A1(n17954), .A2(Out_data[37]), .ZN(n13494) );
NAND2_X2 U8852 ( .A1(n13498), .A2(n17937), .ZN(n13493) );
NAND4_X2 U8853 ( .A1(n13499), .A2(n13500), .A3(n13501), .A4(n13502), .ZN(n5663) );
NAND2_X2 U8854 ( .A1(n13503), .A2(n17845), .ZN(n13501) );
XNOR2_X2 U8855 ( .A(n17203), .B(z_out[38]), .ZN(n13503) );
NAND2_X2 U8856 ( .A1(n17954), .A2(Out_data[38]), .ZN(n13500) );
NAND2_X2 U8857 ( .A1(n13504), .A2(n17937), .ZN(n13499) );
NAND4_X2 U8858 ( .A1(n13505), .A2(n13506), .A3(n13507), .A4(n13508), .ZN(n5662) );
NAND2_X2 U8859 ( .A1(n13509), .A2(n17845), .ZN(n13507) );
XNOR2_X2 U8860 ( .A(n17201), .B(z_out[39]), .ZN(n13509) );
NAND2_X2 U8861 ( .A1(n17954), .A2(Out_data[39]), .ZN(n13506) );
NAND2_X2 U8862 ( .A1(n13510), .A2(n17938), .ZN(n13505) );
NAND4_X2 U8863 ( .A1(n13511), .A2(n13512), .A3(n13513), .A4(n13514), .ZN(n5661) );
NAND2_X2 U8864 ( .A1(n13515), .A2(n17845), .ZN(n13513) );
XNOR2_X2 U8865 ( .A(n17199), .B(z_out[40]), .ZN(n13515) );
NAND2_X2 U8866 ( .A1(n17953), .A2(Out_data[40]), .ZN(n13512) );
NAND2_X2 U8867 ( .A1(n18827), .A2(n17938), .ZN(n13511) );
NAND4_X2 U8868 ( .A1(n13517), .A2(n13518), .A3(n13519), .A4(n13520), .ZN(n5660) );
NAND2_X2 U8869 ( .A1(n13521), .A2(n17845), .ZN(n13519) );
XNOR2_X2 U8870 ( .A(n17197), .B(z_out[41]), .ZN(n13521) );
NAND2_X2 U8871 ( .A1(n17953), .A2(Out_data[41]), .ZN(n13518) );
NAND2_X2 U8872 ( .A1(n18826), .A2(n17938), .ZN(n13517) );
NAND4_X2 U8873 ( .A1(n13523), .A2(n13524), .A3(n13525), .A4(n13526), .ZN(n5659) );
NAND2_X2 U8874 ( .A1(n13527), .A2(n17845), .ZN(n13525) );
XNOR2_X2 U8875 ( .A(n17195), .B(z_out[42]), .ZN(n13527) );
NAND2_X2 U8876 ( .A1(n17953), .A2(Out_data[42]), .ZN(n13524) );
NAND2_X2 U8877 ( .A1(n18825), .A2(n17938), .ZN(n13523) );
NAND4_X2 U8878 ( .A1(n13529), .A2(n13530), .A3(n13531), .A4(n13532), .ZN(n5658) );
NAND2_X2 U8879 ( .A1(n13533), .A2(n17845), .ZN(n13531) );
XNOR2_X2 U8880 ( .A(n17193), .B(z_out[43]), .ZN(n13533) );
NAND2_X2 U8881 ( .A1(n17953), .A2(Out_data[43]), .ZN(n13530) );
NAND2_X2 U8882 ( .A1(n18824), .A2(n17938), .ZN(n13529) );
NAND4_X2 U8883 ( .A1(n13535), .A2(n13536), .A3(n13537), .A4(n13538), .ZN(n5657) );
NAND2_X2 U8884 ( .A1(n13539), .A2(n17845), .ZN(n13537) );
XNOR2_X2 U8885 ( .A(n17191), .B(z_out[44]), .ZN(n13539) );
NAND2_X2 U8886 ( .A1(n17953), .A2(Out_data[44]), .ZN(n13536) );
NAND2_X2 U8887 ( .A1(n18823), .A2(n17940), .ZN(n13535) );
NAND4_X2 U8888 ( .A1(n13541), .A2(n13542), .A3(n13543), .A4(n13544), .ZN(n5656) );
NAND2_X2 U8889 ( .A1(n13545), .A2(n17845), .ZN(n13543) );
XNOR2_X2 U8890 ( .A(n17189), .B(z_out[45]), .ZN(n13545) );
NAND2_X2 U8891 ( .A1(n17953), .A2(Out_data[45]), .ZN(n13542) );
NAND2_X2 U8892 ( .A1(n18822), .A2(n17938), .ZN(n13541) );
NAND4_X2 U8893 ( .A1(n13547), .A2(n13548), .A3(n13549), .A4(n13550), .ZN(n5655) );
NAND2_X2 U8894 ( .A1(n13551), .A2(n17845), .ZN(n13549) );
XNOR2_X2 U8895 ( .A(n17187), .B(z_out[46]), .ZN(n13551) );
NAND2_X2 U8896 ( .A1(n17953), .A2(Out_data[46]), .ZN(n13548) );
NAND2_X2 U8897 ( .A1(n18821), .A2(n17938), .ZN(n13547) );
NAND4_X2 U8898 ( .A1(n13553), .A2(n13554), .A3(n13555), .A4(n13556), .ZN(n5654) );
NAND2_X2 U8899 ( .A1(n13557), .A2(n17845), .ZN(n13555) );
XNOR2_X2 U8900 ( .A(n17185), .B(z_out[47]), .ZN(n13557) );
NAND2_X2 U8901 ( .A1(n17953), .A2(Out_data[47]), .ZN(n13554) );
NAND2_X2 U8902 ( .A1(n18820), .A2(n17938), .ZN(n13553) );
NAND4_X2 U8903 ( .A1(n13559), .A2(n13560), .A3(n13561), .A4(n13562), .ZN(n5653) );
NAND2_X2 U8904 ( .A1(n13563), .A2(n17845), .ZN(n13561) );
XNOR2_X2 U8905 ( .A(n17183), .B(z_out[48]), .ZN(n13563) );
NAND2_X2 U8906 ( .A1(n17953), .A2(Out_data[48]), .ZN(n13560) );
NAND2_X2 U8907 ( .A1(n13564), .A2(n17938), .ZN(n13559) );
NAND4_X2 U8908 ( .A1(n13565), .A2(n13566), .A3(n13567), .A4(n13568), .ZN(n5652) );
NAND2_X2 U8909 ( .A1(n13569), .A2(n17845), .ZN(n13567) );
XNOR2_X2 U8910 ( .A(n17181), .B(z_out[49]), .ZN(n13569) );
NAND2_X2 U8911 ( .A1(n17953), .A2(Out_data[49]), .ZN(n13566) );
NAND2_X2 U8912 ( .A1(n13570), .A2(n17938), .ZN(n13565) );
NAND4_X2 U8913 ( .A1(n13571), .A2(n13572), .A3(n13573), .A4(n13574), .ZN(n5651) );
NAND2_X2 U8914 ( .A1(n13575), .A2(n17845), .ZN(n13573) );
XNOR2_X2 U8915 ( .A(n17179), .B(z_out[50]), .ZN(n13575) );
NAND2_X2 U8916 ( .A1(n17953), .A2(Out_data[50]), .ZN(n13572) );
NAND2_X2 U8917 ( .A1(n13576), .A2(n17938), .ZN(n13571) );
NAND4_X2 U8918 ( .A1(n13577), .A2(n13578), .A3(n13579), .A4(n13580), .ZN(n5650) );
NAND2_X2 U8919 ( .A1(n13581), .A2(n17845), .ZN(n13579) );
XNOR2_X2 U8920 ( .A(n17177), .B(z_out[51]), .ZN(n13581) );
NAND2_X2 U8921 ( .A1(n17952), .A2(Out_data[51]), .ZN(n13578) );
NAND2_X2 U8922 ( .A1(n13582), .A2(n17938), .ZN(n13577) );
NAND4_X2 U8923 ( .A1(n13583), .A2(n13584), .A3(n13585), .A4(n13586), .ZN(n5649) );
NAND2_X2 U8924 ( .A1(n13587), .A2(n17845), .ZN(n13585) );
XNOR2_X2 U8925 ( .A(n17175), .B(z_out[52]), .ZN(n13587) );
NAND2_X2 U8926 ( .A1(n17952), .A2(Out_data[52]), .ZN(n13584) );
NAND2_X2 U8927 ( .A1(n13588), .A2(n17939), .ZN(n13583) );
NAND4_X2 U8928 ( .A1(n13589), .A2(n13590), .A3(n13591), .A4(n13592), .ZN(n5648) );
NAND2_X2 U8929 ( .A1(n13593), .A2(n17844), .ZN(n13591) );
XNOR2_X2 U8930 ( .A(n17173), .B(z_out[53]), .ZN(n13593) );
NAND2_X2 U8931 ( .A1(n17952), .A2(Out_data[53]), .ZN(n13590) );
NAND2_X2 U8932 ( .A1(n13594), .A2(n17939), .ZN(n13589) );
NAND4_X2 U8933 ( .A1(n13595), .A2(n13596), .A3(n13597), .A4(n13598), .ZN(n5647) );
NAND2_X2 U8934 ( .A1(n13599), .A2(n17844), .ZN(n13597) );
XNOR2_X2 U8935 ( .A(n17171), .B(z_out[54]), .ZN(n13599) );
NAND2_X2 U8936 ( .A1(n17952), .A2(Out_data[54]), .ZN(n13596) );
NAND2_X2 U8937 ( .A1(n13600), .A2(n17939), .ZN(n13595) );
NAND4_X2 U8938 ( .A1(n13601), .A2(n13602), .A3(n13603), .A4(n13604), .ZN(n5646) );
NAND2_X2 U8939 ( .A1(n13605), .A2(n17844), .ZN(n13603) );
XNOR2_X2 U8940 ( .A(n17169), .B(z_out[55]), .ZN(n13605) );
NAND2_X2 U8941 ( .A1(n17952), .A2(Out_data[55]), .ZN(n13602) );
NAND2_X2 U8942 ( .A1(n13606), .A2(n17939), .ZN(n13601) );
NAND4_X2 U8943 ( .A1(n13607), .A2(n13608), .A3(n13609), .A4(n13610), .ZN(n5645) );
NAND2_X2 U8944 ( .A1(n13611), .A2(n17844), .ZN(n13609) );
XNOR2_X2 U8945 ( .A(n17167), .B(z_out[56]), .ZN(n13611) );
NAND2_X2 U8946 ( .A1(n17952), .A2(Out_data[56]), .ZN(n13608) );
NAND2_X2 U8947 ( .A1(n18819), .A2(n17939), .ZN(n13607) );
NAND4_X2 U8948 ( .A1(n13613), .A2(n13614), .A3(n13615), .A4(n13616), .ZN(n5644) );
NAND2_X2 U8949 ( .A1(n13617), .A2(n17844), .ZN(n13615) );
XNOR2_X2 U8950 ( .A(n17165), .B(z_out[57]), .ZN(n13617) );
NAND2_X2 U8951 ( .A1(n17952), .A2(Out_data[57]), .ZN(n13614) );
NAND2_X2 U8952 ( .A1(n18818), .A2(n17939), .ZN(n13613) );
NAND4_X2 U8953 ( .A1(n13619), .A2(n13620), .A3(n13621), .A4(n13622), .ZN(n5643) );
NAND2_X2 U8954 ( .A1(n13623), .A2(n17844), .ZN(n13621) );
XNOR2_X2 U8955 ( .A(n17163), .B(z_out[58]), .ZN(n13623) );
NAND2_X2 U8956 ( .A1(n17952), .A2(Out_data[58]), .ZN(n13620) );
NAND2_X2 U8957 ( .A1(n18817), .A2(n17939), .ZN(n13619) );
NAND4_X2 U8958 ( .A1(n13625), .A2(n13626), .A3(n13627), .A4(n13628), .ZN(n5642) );
NAND2_X2 U8959 ( .A1(n13629), .A2(n17844), .ZN(n13627) );
XNOR2_X2 U8960 ( .A(n17161), .B(z_out[59]), .ZN(n13629) );
NAND2_X2 U8961 ( .A1(n17952), .A2(Out_data[59]), .ZN(n13626) );
NAND2_X2 U8962 ( .A1(n18816), .A2(n17939), .ZN(n13625) );
NAND4_X2 U8963 ( .A1(n13631), .A2(n13632), .A3(n13633), .A4(n13634), .ZN(n5641) );
NAND2_X2 U8964 ( .A1(n13635), .A2(n17844), .ZN(n13633) );
XNOR2_X2 U8965 ( .A(n17159), .B(z_out[60]), .ZN(n13635) );
NAND2_X2 U8966 ( .A1(n17952), .A2(Out_data[60]), .ZN(n13632) );
NAND2_X2 U8967 ( .A1(n18815), .A2(n17939), .ZN(n13631) );
NAND4_X2 U8968 ( .A1(n13637), .A2(n13638), .A3(n13639), .A4(n13640), .ZN(n5640) );
NAND2_X2 U8969 ( .A1(n13641), .A2(n17844), .ZN(n13639) );
XNOR2_X2 U8970 ( .A(n17157), .B(z_out[61]), .ZN(n13641) );
NAND2_X2 U8971 ( .A1(n17952), .A2(Out_data[61]), .ZN(n13638) );
NAND2_X2 U8972 ( .A1(n18814), .A2(n17939), .ZN(n13637) );
NAND4_X2 U8973 ( .A1(n13643), .A2(n13644), .A3(n13645), .A4(n13646), .ZN(n5639) );
NAND2_X2 U8974 ( .A1(n13647), .A2(n17844), .ZN(n13645) );
XNOR2_X2 U8975 ( .A(n17155), .B(z_out[62]), .ZN(n13647) );
NAND2_X2 U8976 ( .A1(n17951), .A2(Out_data[62]), .ZN(n13644) );
NAND2_X2 U8977 ( .A1(n18813), .A2(n17939), .ZN(n13643) );
NAND4_X2 U8978 ( .A1(n13649), .A2(n13650), .A3(n13651), .A4(n13652), .ZN(n5638) );
NAND2_X2 U8979 ( .A1(n13653), .A2(n17844), .ZN(n13651) );
XNOR2_X2 U8980 ( .A(n17153), .B(z_out[63]), .ZN(n13653) );
NAND2_X2 U8981 ( .A1(n17951), .A2(Out_data[63]), .ZN(n13650) );
NAND2_X2 U8982 ( .A1(n18812), .A2(n17939), .ZN(n13649) );
NAND4_X2 U8983 ( .A1(n13655), .A2(n13656), .A3(n13657), .A4(n13658), .ZN(n5637) );
NAND2_X2 U8984 ( .A1(n13659), .A2(n17844), .ZN(n13658) );
XNOR2_X2 U8985 ( .A(n17151), .B(z_out[64]), .ZN(n13659) );
NAND2_X2 U8986 ( .A1(n17951), .A2(Out_data[64]), .ZN(n13657) );
NAND2_X2 U8988 ( .A1(n18811), .A2(n17940), .ZN(n13655) );
NAND4_X2 U8989 ( .A1(n13663), .A2(n13664), .A3(n13665), .A4(n13666), .ZN(n5636) );
NAND2_X2 U8990 ( .A1(n13667), .A2(n17844), .ZN(n13666) );
XNOR2_X2 U8991 ( .A(n17149), .B(z_out[65]), .ZN(n13667) );
NAND2_X2 U8992 ( .A1(n17951), .A2(Out_data[65]), .ZN(n13665) );
NAND2_X2 U8993 ( .A1(n17930), .A2(n13668), .ZN(n13664) );
NAND2_X2 U8994 ( .A1(n18810), .A2(n17940), .ZN(n13663) );
NAND4_X2 U8995 ( .A1(n13670), .A2(n13671), .A3(n13672), .A4(n13673), .ZN(n5635) );
NAND2_X2 U8996 ( .A1(n13674), .A2(n17844), .ZN(n13673) );
XNOR2_X2 U8997 ( .A(n17147), .B(z_out[66]), .ZN(n13674) );
NAND2_X2 U8998 ( .A1(n17951), .A2(Out_data[66]), .ZN(n13672) );
NAND2_X2 U9000 ( .A1(n18809), .A2(n17940), .ZN(n13670) );
NAND4_X2 U9001 ( .A1(n13677), .A2(n13678), .A3(n13679), .A4(n13680), .ZN(n5634) );
NAND2_X2 U9002 ( .A1(n13681), .A2(n17844), .ZN(n13679) );
XNOR2_X2 U9003 ( .A(n17145), .B(z_out[67]), .ZN(n13681) );
NAND2_X2 U9004 ( .A1(n17951), .A2(Out_data[67]), .ZN(n13678) );
NAND2_X2 U9005 ( .A1(n18808), .A2(n17940), .ZN(n13677) );
NAND4_X2 U9006 ( .A1(n13683), .A2(n13684), .A3(n13685), .A4(n13686), .ZN(n5633) );
NAND2_X2 U9007 ( .A1(n13687), .A2(n17844), .ZN(n13685) );
XNOR2_X2 U9008 ( .A(n17143), .B(z_out[68]), .ZN(n13687) );
NAND2_X2 U9009 ( .A1(n17951), .A2(Out_data[68]), .ZN(n13684) );
NAND2_X2 U9010 ( .A1(n18807), .A2(n17940), .ZN(n13683) );
NAND4_X2 U9011 ( .A1(n13689), .A2(n13690), .A3(n13691), .A4(n13692), .ZN(n5632) );
NAND2_X2 U9012 ( .A1(n13693), .A2(n17844), .ZN(n13691) );
XNOR2_X2 U9013 ( .A(n17141), .B(z_out[69]), .ZN(n13693) );
NAND2_X2 U9014 ( .A1(n17951), .A2(Out_data[69]), .ZN(n13690) );
NAND2_X2 U9015 ( .A1(n18806), .A2(n17940), .ZN(n13689) );
NAND4_X2 U9016 ( .A1(n13695), .A2(n13696), .A3(n13697), .A4(n13698), .ZN(n5631) );
NAND2_X2 U9017 ( .A1(n13699), .A2(n17844), .ZN(n13697) );
XNOR2_X2 U9018 ( .A(n17139), .B(z_out[70]), .ZN(n13699) );
NAND2_X2 U9019 ( .A1(n17951), .A2(Out_data[70]), .ZN(n13696) );
NAND2_X2 U9020 ( .A1(n18805), .A2(n17940), .ZN(n13695) );
NAND4_X2 U9021 ( .A1(n13701), .A2(n13702), .A3(n13703), .A4(n13704), .ZN(n5630) );
NAND2_X2 U9022 ( .A1(n13705), .A2(n17844), .ZN(n13703) );
XNOR2_X2 U9023 ( .A(n17137), .B(z_out[71]), .ZN(n13705) );
NAND2_X2 U9024 ( .A1(n17951), .A2(Out_data[71]), .ZN(n13702) );
NAND2_X2 U9025 ( .A1(n18804), .A2(n17940), .ZN(n13701) );
NAND4_X2 U9026 ( .A1(n13707), .A2(n13708), .A3(n13709), .A4(n13710), .ZN(n5629) );
NAND2_X2 U9027 ( .A1(n13711), .A2(n17843), .ZN(n13709) );
XNOR2_X2 U9028 ( .A(n17135), .B(z_out[72]), .ZN(n13711) );
NAND2_X2 U9029 ( .A1(n17951), .A2(Out_data[72]), .ZN(n13708) );
NAND2_X2 U9030 ( .A1(n18803), .A2(n17940), .ZN(n13707) );
NAND4_X2 U9031 ( .A1(n13713), .A2(n13714), .A3(n13715), .A4(n13716), .ZN(n5628) );
NAND2_X2 U9032 ( .A1(n13717), .A2(n17843), .ZN(n13715) );
XNOR2_X2 U9033 ( .A(n17133), .B(z_out[73]), .ZN(n13717) );
NAND2_X2 U9034 ( .A1(n17950), .A2(Out_data[73]), .ZN(n13714) );
NAND2_X2 U9035 ( .A1(n18802), .A2(n17940), .ZN(n13713) );
NAND4_X2 U9036 ( .A1(n13719), .A2(n13720), .A3(n13721), .A4(n13722), .ZN(n5627) );
NAND2_X2 U9037 ( .A1(n13723), .A2(n17843), .ZN(n13721) );
XNOR2_X2 U9038 ( .A(n17131), .B(z_out[74]), .ZN(n13723) );
NAND2_X2 U9039 ( .A1(n17950), .A2(Out_data[74]), .ZN(n13720) );
NAND2_X2 U9040 ( .A1(n18801), .A2(n17940), .ZN(n13719) );
NAND4_X2 U9041 ( .A1(n13725), .A2(n13726), .A3(n13727), .A4(n13728), .ZN(n5626) );
NAND2_X2 U9042 ( .A1(n13729), .A2(n17843), .ZN(n13727) );
XNOR2_X2 U9043 ( .A(n17129), .B(z_out[75]), .ZN(n13729) );
NAND2_X2 U9044 ( .A1(n17950), .A2(Out_data[75]), .ZN(n13726) );
NAND2_X2 U9045 ( .A1(n18800), .A2(n17941), .ZN(n13725) );
NAND4_X2 U9046 ( .A1(n13731), .A2(n13732), .A3(n13733), .A4(n13734), .ZN(n5625) );
NAND2_X2 U9047 ( .A1(n13735), .A2(n17843), .ZN(n13733) );
XNOR2_X2 U9048 ( .A(n17127), .B(z_out[76]), .ZN(n13735) );
NAND2_X2 U9049 ( .A1(n17950), .A2(Out_data[76]), .ZN(n13732) );
NAND2_X2 U9050 ( .A1(n18799), .A2(n17941), .ZN(n13731) );
NAND4_X2 U9051 ( .A1(n13737), .A2(n13738), .A3(n13739), .A4(n13740), .ZN(n5624) );
NAND2_X2 U9052 ( .A1(n13741), .A2(n17843), .ZN(n13739) );
XNOR2_X2 U9053 ( .A(n17125), .B(z_out[77]), .ZN(n13741) );
NAND2_X2 U9054 ( .A1(n17950), .A2(Out_data[77]), .ZN(n13738) );
NAND2_X2 U9055 ( .A1(n18798), .A2(n17941), .ZN(n13737) );
NAND4_X2 U9056 ( .A1(n13743), .A2(n13744), .A3(n13745), .A4(n13746), .ZN(n5623) );
NAND2_X2 U9057 ( .A1(n13747), .A2(n17843), .ZN(n13745) );
XNOR2_X2 U9058 ( .A(n17123), .B(z_out[78]), .ZN(n13747) );
NAND2_X2 U9059 ( .A1(n17950), .A2(Out_data[78]), .ZN(n13744) );
NAND2_X2 U9060 ( .A1(n18797), .A2(n17941), .ZN(n13743) );
NAND4_X2 U9061 ( .A1(n13749), .A2(n13750), .A3(n13751), .A4(n13752), .ZN(n5622) );
NAND2_X2 U9062 ( .A1(n13753), .A2(n17843), .ZN(n13751) );
XNOR2_X2 U9063 ( .A(n17121), .B(z_out[79]), .ZN(n13753) );
NAND2_X2 U9064 ( .A1(n17950), .A2(Out_data[79]), .ZN(n13750) );
NAND2_X2 U9065 ( .A1(n18796), .A2(n17941), .ZN(n13749) );
NAND4_X2 U9066 ( .A1(n13755), .A2(n13756), .A3(n13757), .A4(n13758), .ZN(n5621) );
NAND2_X2 U9067 ( .A1(n13759), .A2(n17843), .ZN(n13757) );
XNOR2_X2 U9068 ( .A(n17119), .B(z_out[80]), .ZN(n13759) );
NAND2_X2 U9069 ( .A1(n17950), .A2(Out_data[80]), .ZN(n13756) );
NAND2_X2 U9070 ( .A1(n18795), .A2(n17941), .ZN(n13755) );
NAND4_X2 U9071 ( .A1(n13761), .A2(n13762), .A3(n13763), .A4(n13764), .ZN(n5620) );
NAND2_X2 U9072 ( .A1(n13765), .A2(n17843), .ZN(n13763) );
XNOR2_X2 U9073 ( .A(n17117), .B(z_out[81]), .ZN(n13765) );
NAND2_X2 U9074 ( .A1(n17950), .A2(Out_data[81]), .ZN(n13762) );
NAND2_X2 U9075 ( .A1(n18794), .A2(n17941), .ZN(n13761) );
NAND4_X2 U9076 ( .A1(n13767), .A2(n13768), .A3(n13769), .A4(n13770), .ZN(n5619) );
NAND2_X2 U9077 ( .A1(n13771), .A2(n17843), .ZN(n13769) );
XNOR2_X2 U9078 ( .A(n17115), .B(z_out[82]), .ZN(n13771) );
NAND2_X2 U9079 ( .A1(n17950), .A2(Out_data[82]), .ZN(n13768) );
NAND2_X2 U9080 ( .A1(n18793), .A2(n17941), .ZN(n13767) );
NAND4_X2 U9081 ( .A1(n13773), .A2(n13774), .A3(n13775), .A4(n13776), .ZN(n5618) );
NAND2_X2 U9082 ( .A1(n13777), .A2(n17843), .ZN(n13775) );
XNOR2_X2 U9083 ( .A(n17113), .B(z_out[83]), .ZN(n13777) );
NAND2_X2 U9084 ( .A1(n17950), .A2(Out_data[83]), .ZN(n13774) );
NAND2_X2 U9085 ( .A1(n18792), .A2(n17941), .ZN(n13773) );
NAND4_X2 U9086 ( .A1(n13779), .A2(n13780), .A3(n13781), .A4(n13782), .ZN(n5617) );
NAND2_X2 U9087 ( .A1(n13783), .A2(n17843), .ZN(n13781) );
XNOR2_X2 U9088 ( .A(n17111), .B(z_out[84]), .ZN(n13783) );
NAND2_X2 U9089 ( .A1(n17949), .A2(Out_data[84]), .ZN(n13780) );
NAND2_X2 U9090 ( .A1(n18791), .A2(n17941), .ZN(n13779) );
NAND4_X2 U9091 ( .A1(n13785), .A2(n13786), .A3(n13787), .A4(n13788), .ZN(n5616) );
NAND2_X2 U9092 ( .A1(n13789), .A2(n17843), .ZN(n13787) );
XNOR2_X2 U9093 ( .A(n17109), .B(z_out[85]), .ZN(n13789) );
NAND2_X2 U9094 ( .A1(n17949), .A2(Out_data[85]), .ZN(n13786) );
NAND2_X2 U9095 ( .A1(n18790), .A2(n17941), .ZN(n13785) );
NAND4_X2 U9096 ( .A1(n13791), .A2(n13792), .A3(n13793), .A4(n13794), .ZN(n5615) );
NAND2_X2 U9097 ( .A1(n13795), .A2(n17843), .ZN(n13793) );
XNOR2_X2 U9098 ( .A(n17107), .B(z_out[86]), .ZN(n13795) );
NAND2_X2 U9099 ( .A1(n17949), .A2(Out_data[86]), .ZN(n13792) );
NAND2_X2 U9100 ( .A1(n18789), .A2(n17941), .ZN(n13791) );
NAND4_X2 U9101 ( .A1(n13797), .A2(n13798), .A3(n13799), .A4(n13800), .ZN(n5614) );
NAND2_X2 U9102 ( .A1(n13801), .A2(n17843), .ZN(n13799) );
XNOR2_X2 U9103 ( .A(n17105), .B(z_out[87]), .ZN(n13801) );
NAND2_X2 U9104 ( .A1(n17949), .A2(Out_data[87]), .ZN(n13798) );
NAND2_X2 U9105 ( .A1(n18788), .A2(n17942), .ZN(n13797) );
NAND4_X2 U9106 ( .A1(n13803), .A2(n13804), .A3(n13805), .A4(n13806), .ZN(n5613) );
NAND2_X2 U9107 ( .A1(n13807), .A2(n17843), .ZN(n13805) );
XNOR2_X2 U9108 ( .A(n17103), .B(z_out[88]), .ZN(n13807) );
NAND2_X2 U9109 ( .A1(n17949), .A2(Out_data[88]), .ZN(n13804) );
NAND2_X2 U9110 ( .A1(n18787), .A2(n17942), .ZN(n13803) );
NAND4_X2 U9111 ( .A1(n13809), .A2(n13810), .A3(n13811), .A4(n13812), .ZN(n5612) );
NAND2_X2 U9112 ( .A1(n13813), .A2(n17843), .ZN(n13811) );
XNOR2_X2 U9113 ( .A(n17101), .B(z_out[89]), .ZN(n13813) );
NAND2_X2 U9114 ( .A1(n17949), .A2(Out_data[89]), .ZN(n13810) );
NAND2_X2 U9115 ( .A1(n18786), .A2(n17942), .ZN(n13809) );
NAND4_X2 U9116 ( .A1(n13815), .A2(n13816), .A3(n13817), .A4(n13818), .ZN(n5611) );
NAND2_X2 U9117 ( .A1(n13819), .A2(n17843), .ZN(n13817) );
XNOR2_X2 U9118 ( .A(n17099), .B(z_out[90]), .ZN(n13819) );
NAND2_X2 U9119 ( .A1(n17949), .A2(Out_data[90]), .ZN(n13816) );
NAND2_X2 U9120 ( .A1(n18785), .A2(n17942), .ZN(n13815) );
NAND4_X2 U9121 ( .A1(n13821), .A2(n13822), .A3(n13823), .A4(n13824), .ZN(n5610) );
NAND2_X2 U9122 ( .A1(n13825), .A2(n17842), .ZN(n13823) );
XNOR2_X2 U9123 ( .A(n17097), .B(z_out[91]), .ZN(n13825) );
NAND2_X2 U9124 ( .A1(n17949), .A2(Out_data[91]), .ZN(n13822) );
NAND2_X2 U9125 ( .A1(n18784), .A2(n17942), .ZN(n13821) );
NAND4_X2 U9126 ( .A1(n13827), .A2(n13828), .A3(n13829), .A4(n13830), .ZN(n5609) );
NAND2_X2 U9127 ( .A1(n13831), .A2(n17842), .ZN(n13829) );
XNOR2_X2 U9128 ( .A(n17095), .B(z_out[92]), .ZN(n13831) );
NAND2_X2 U9129 ( .A1(n17949), .A2(Out_data[92]), .ZN(n13828) );
NAND2_X2 U9130 ( .A1(n18783), .A2(n17942), .ZN(n13827) );
NAND4_X2 U9131 ( .A1(n13833), .A2(n13834), .A3(n13835), .A4(n13836), .ZN(n5608) );
NAND2_X2 U9132 ( .A1(n13837), .A2(n17842), .ZN(n13835) );
XNOR2_X2 U9133 ( .A(n17093), .B(z_out[93]), .ZN(n13837) );
NAND2_X2 U9134 ( .A1(n17949), .A2(Out_data[93]), .ZN(n13834) );
NAND2_X2 U9135 ( .A1(n18782), .A2(n17942), .ZN(n13833) );
NAND4_X2 U9136 ( .A1(n13839), .A2(n13840), .A3(n13841), .A4(n13842), .ZN(n5607) );
NAND2_X2 U9137 ( .A1(n13843), .A2(n17842), .ZN(n13841) );
XNOR2_X2 U9138 ( .A(n17091), .B(z_out[94]), .ZN(n13843) );
NAND2_X2 U9139 ( .A1(n17949), .A2(Out_data[94]), .ZN(n13840) );
NAND2_X2 U9140 ( .A1(n18781), .A2(n17942), .ZN(n13839) );
NAND4_X2 U9141 ( .A1(n13845), .A2(n13846), .A3(n13847), .A4(n13848), .ZN(n5606) );
NAND2_X2 U9142 ( .A1(n13849), .A2(n17842), .ZN(n13847) );
XNOR2_X2 U9143 ( .A(n17089), .B(z_out[95]), .ZN(n13849) );
NAND2_X2 U9144 ( .A1(n17948), .A2(Out_data[95]), .ZN(n13846) );
NAND2_X2 U9145 ( .A1(n18780), .A2(n17942), .ZN(n13845) );
NAND4_X2 U9146 ( .A1(n13851), .A2(n13852), .A3(n13853), .A4(n13854), .ZN(n5605) );
NAND2_X2 U9147 ( .A1(n13855), .A2(n17842), .ZN(n13853) );
XNOR2_X2 U9148 ( .A(n17087), .B(z_out[96]), .ZN(n13855) );
NAND2_X2 U9149 ( .A1(n17948), .A2(Out_data[96]), .ZN(n13852) );
NAND2_X2 U9150 ( .A1(n18779), .A2(n17942), .ZN(n13851) );
NAND4_X2 U9151 ( .A1(n13857), .A2(n13858), .A3(n13859), .A4(n13860), .ZN(n5604) );
NAND2_X2 U9152 ( .A1(n13861), .A2(n17842), .ZN(n13859) );
XNOR2_X2 U9153 ( .A(n17085), .B(z_out[97]), .ZN(n13861) );
NAND2_X2 U9154 ( .A1(n17948), .A2(Out_data[97]), .ZN(n13858) );
NAND2_X2 U9155 ( .A1(n18778), .A2(n17942), .ZN(n13857) );
NAND4_X2 U9156 ( .A1(n13863), .A2(n13864), .A3(n13865), .A4(n13866), .ZN(n5603) );
NAND2_X2 U9157 ( .A1(n13867), .A2(n17842), .ZN(n13865) );
XNOR2_X2 U9158 ( .A(n17083), .B(z_out[98]), .ZN(n13867) );
NAND2_X2 U9159 ( .A1(n17948), .A2(Out_data[98]), .ZN(n13864) );
NAND2_X2 U9160 ( .A1(n18777), .A2(n17942), .ZN(n13863) );
NAND4_X2 U9161 ( .A1(n13869), .A2(n13870), .A3(n13871), .A4(n13872), .ZN(n5602) );
NAND2_X2 U9162 ( .A1(n13873), .A2(n17842), .ZN(n13871) );
XNOR2_X2 U9163 ( .A(n17081), .B(z_out[99]), .ZN(n13873) );
NAND2_X2 U9164 ( .A1(n17948), .A2(Out_data[99]), .ZN(n13870) );
NAND2_X2 U9165 ( .A1(n18776), .A2(n17943), .ZN(n13869) );
NAND4_X2 U9166 ( .A1(n13875), .A2(n13876), .A3(n13877), .A4(n13878), .ZN(n5601) );
NAND2_X2 U9167 ( .A1(n13879), .A2(n17842), .ZN(n13877) );
XNOR2_X2 U9168 ( .A(n17079), .B(z_out[100]), .ZN(n13879) );
NAND2_X2 U9169 ( .A1(n17948), .A2(Out_data[100]), .ZN(n13876) );
NAND2_X2 U9170 ( .A1(n18775), .A2(n17943), .ZN(n13875) );
NAND4_X2 U9171 ( .A1(n13881), .A2(n13882), .A3(n13883), .A4(n13884), .ZN(n5600) );
NAND2_X2 U9172 ( .A1(n13885), .A2(n17842), .ZN(n13883) );
XNOR2_X2 U9173 ( .A(n17077), .B(z_out[101]), .ZN(n13885) );
NAND2_X2 U9174 ( .A1(n17948), .A2(Out_data[101]), .ZN(n13882) );
NAND2_X2 U9175 ( .A1(n18774), .A2(n17943), .ZN(n13881) );
NAND4_X2 U9176 ( .A1(n13887), .A2(n13888), .A3(n13889), .A4(n13890), .ZN(n5599) );
NAND2_X2 U9177 ( .A1(n13891), .A2(n17842), .ZN(n13889) );
XNOR2_X2 U9178 ( .A(n17075), .B(z_out[102]), .ZN(n13891) );
NAND2_X2 U9179 ( .A1(n17948), .A2(Out_data[102]), .ZN(n13888) );
NAND2_X2 U9180 ( .A1(n18773), .A2(n17943), .ZN(n13887) );
NAND4_X2 U9181 ( .A1(n13893), .A2(n13894), .A3(n13895), .A4(n13896), .ZN(n5598) );
NAND2_X2 U9182 ( .A1(n13897), .A2(n17842), .ZN(n13895) );
XNOR2_X2 U9183 ( .A(n17073), .B(z_out[103]), .ZN(n13897) );
NAND2_X2 U9184 ( .A1(n17948), .A2(Out_data[103]), .ZN(n13894) );
NAND2_X2 U9185 ( .A1(n18772), .A2(n17943), .ZN(n13893) );
NAND4_X2 U9186 ( .A1(n13899), .A2(n13900), .A3(n13901), .A4(n13902), .ZN(n5597) );
NAND2_X2 U9187 ( .A1(n13903), .A2(n17842), .ZN(n13901) );
XNOR2_X2 U9188 ( .A(n17071), .B(z_out[104]), .ZN(n13903) );
NAND2_X2 U9189 ( .A1(n17948), .A2(Out_data[104]), .ZN(n13900) );
NAND2_X2 U9190 ( .A1(n18771), .A2(n17943), .ZN(n13899) );
NAND4_X2 U9191 ( .A1(n13905), .A2(n13906), .A3(n13907), .A4(n13908), .ZN(n5596) );
NAND2_X2 U9192 ( .A1(n13909), .A2(n17842), .ZN(n13907) );
XNOR2_X2 U9193 ( .A(n17069), .B(z_out[105]), .ZN(n13909) );
NAND2_X2 U9194 ( .A1(n17948), .A2(Out_data[105]), .ZN(n13906) );
NAND2_X2 U9195 ( .A1(n18770), .A2(n17943), .ZN(n13905) );
NAND4_X2 U9196 ( .A1(n13911), .A2(n13912), .A3(n13913), .A4(n13914), .ZN(n5595) );
NAND2_X2 U9197 ( .A1(n13915), .A2(n17842), .ZN(n13913) );
XNOR2_X2 U9198 ( .A(n17067), .B(z_out[106]), .ZN(n13915) );
NAND2_X2 U9199 ( .A1(n17947), .A2(Out_data[106]), .ZN(n13912) );
NAND2_X2 U9200 ( .A1(n18769), .A2(n17943), .ZN(n13911) );
NAND4_X2 U9201 ( .A1(n13917), .A2(n13918), .A3(n13919), .A4(n13920), .ZN(n5594) );
NAND2_X2 U9202 ( .A1(n13921), .A2(n17842), .ZN(n13919) );
XNOR2_X2 U9203 ( .A(n17065), .B(z_out[107]), .ZN(n13921) );
NAND2_X2 U9204 ( .A1(n17947), .A2(Out_data[107]), .ZN(n13918) );
NAND2_X2 U9205 ( .A1(n18768), .A2(n17943), .ZN(n13917) );
NAND4_X2 U9206 ( .A1(n13923), .A2(n13924), .A3(n13925), .A4(n13926), .ZN(n5593) );
NAND2_X2 U9207 ( .A1(n13927), .A2(n17842), .ZN(n13925) );
XNOR2_X2 U9208 ( .A(n17063), .B(z_out[108]), .ZN(n13927) );
NAND2_X2 U9209 ( .A1(n17947), .A2(Out_data[108]), .ZN(n13924) );
NAND2_X2 U9210 ( .A1(n18767), .A2(n17943), .ZN(n13923) );
NAND4_X2 U9211 ( .A1(n13929), .A2(n13930), .A3(n13931), .A4(n13932), .ZN(n5592) );
NAND2_X2 U9212 ( .A1(n13933), .A2(n17842), .ZN(n13931) );
XNOR2_X2 U9213 ( .A(n17061), .B(z_out[109]), .ZN(n13933) );
NAND2_X2 U9214 ( .A1(n17947), .A2(Out_data[109]), .ZN(n13930) );
NAND2_X2 U9215 ( .A1(n18766), .A2(n17943), .ZN(n13929) );
NAND4_X2 U9216 ( .A1(n13935), .A2(n13936), .A3(n13937), .A4(n13938), .ZN(n5591) );
NAND2_X2 U9217 ( .A1(n13939), .A2(n17841), .ZN(n13937) );
XNOR2_X2 U9218 ( .A(n17059), .B(z_out[110]), .ZN(n13939) );
NAND2_X2 U9219 ( .A1(n17947), .A2(Out_data[110]), .ZN(n13936) );
NAND2_X2 U9220 ( .A1(n18765), .A2(n17943), .ZN(n13935) );
NAND4_X2 U9221 ( .A1(n13941), .A2(n13942), .A3(n13943), .A4(n13944), .ZN(n5590) );
NAND2_X2 U9222 ( .A1(n13945), .A2(n17841), .ZN(n13943) );
XNOR2_X2 U9223 ( .A(n17057), .B(z_out[111]), .ZN(n13945) );
NAND2_X2 U9224 ( .A1(n17947), .A2(Out_data[111]), .ZN(n13942) );
NAND2_X2 U9225 ( .A1(n18764), .A2(n17944), .ZN(n13941) );
NAND4_X2 U9226 ( .A1(n13947), .A2(n13948), .A3(n13949), .A4(n13950), .ZN(n5589) );
NAND2_X2 U9227 ( .A1(n13951), .A2(n17841), .ZN(n13949) );
XNOR2_X2 U9228 ( .A(n17055), .B(z_out[112]), .ZN(n13951) );
NAND2_X2 U9229 ( .A1(n17947), .A2(Out_data[112]), .ZN(n13948) );
NAND2_X2 U9230 ( .A1(n18763), .A2(n17944), .ZN(n13947) );
NAND4_X2 U9231 ( .A1(n13953), .A2(n13954), .A3(n13955), .A4(n13956), .ZN(n5588) );
NAND2_X2 U9232 ( .A1(n13957), .A2(n17841), .ZN(n13955) );
XNOR2_X2 U9233 ( .A(n17053), .B(z_out[113]), .ZN(n13957) );
NAND2_X2 U9234 ( .A1(n17947), .A2(Out_data[113]), .ZN(n13954) );
NAND2_X2 U9235 ( .A1(n18762), .A2(n17944), .ZN(n13953) );
NAND4_X2 U9236 ( .A1(n13959), .A2(n13960), .A3(n13961), .A4(n13962), .ZN(n5587) );
NAND2_X2 U9237 ( .A1(n13963), .A2(n17841), .ZN(n13961) );
XNOR2_X2 U9238 ( .A(n17051), .B(z_out[114]), .ZN(n13963) );
NAND2_X2 U9239 ( .A1(n17947), .A2(Out_data[114]), .ZN(n13960) );
NAND2_X2 U9240 ( .A1(n18761), .A2(n17944), .ZN(n13959) );
NAND4_X2 U9241 ( .A1(n13965), .A2(n13966), .A3(n13967), .A4(n13968), .ZN(n5586) );
NAND2_X2 U9242 ( .A1(n13969), .A2(n17841), .ZN(n13967) );
XNOR2_X2 U9243 ( .A(n17049), .B(z_out[115]), .ZN(n13969) );
NAND2_X2 U9244 ( .A1(n17947), .A2(Out_data[115]), .ZN(n13966) );
NAND2_X2 U9245 ( .A1(n18760), .A2(n17944), .ZN(n13965) );
NAND4_X2 U9246 ( .A1(n13971), .A2(n13972), .A3(n13973), .A4(n13974), .ZN(n5585) );
NAND2_X2 U9247 ( .A1(n13975), .A2(n17841), .ZN(n13973) );
XNOR2_X2 U9248 ( .A(n17047), .B(z_out[116]), .ZN(n13975) );
NAND2_X2 U9249 ( .A1(n17947), .A2(Out_data[116]), .ZN(n13972) );
NAND2_X2 U9250 ( .A1(n18759), .A2(n17944), .ZN(n13971) );
NAND4_X2 U9251 ( .A1(n13977), .A2(n13978), .A3(n13979), .A4(n13980), .ZN(n5584) );
NAND2_X2 U9252 ( .A1(n13981), .A2(n17841), .ZN(n13979) );
XNOR2_X2 U9253 ( .A(n17045), .B(z_out[117]), .ZN(n13981) );
NAND2_X2 U9254 ( .A1(n17946), .A2(Out_data[117]), .ZN(n13978) );
NAND2_X2 U9255 ( .A1(n18758), .A2(n17944), .ZN(n13977) );
NAND4_X2 U9256 ( .A1(n13983), .A2(n13984), .A3(n13985), .A4(n13986), .ZN(n5583) );
NAND2_X2 U9257 ( .A1(n13987), .A2(n17841), .ZN(n13985) );
XNOR2_X2 U9258 ( .A(n17043), .B(z_out[118]), .ZN(n13987) );
NAND2_X2 U9259 ( .A1(n17946), .A2(Out_data[118]), .ZN(n13984) );
NAND2_X2 U9260 ( .A1(n18757), .A2(n17944), .ZN(n13983) );
NAND4_X2 U9261 ( .A1(n13989), .A2(n13990), .A3(n13991), .A4(n13992), .ZN(n5582) );
NAND2_X2 U9262 ( .A1(n13993), .A2(n17841), .ZN(n13991) );
XNOR2_X2 U9263 ( .A(n17041), .B(z_out[119]), .ZN(n13993) );
NAND2_X2 U9264 ( .A1(n17946), .A2(Out_data[119]), .ZN(n13990) );
NAND2_X2 U9265 ( .A1(n18756), .A2(n17944), .ZN(n13989) );
NAND2_X2 U9267 ( .A1(n13998), .A2(n17841), .ZN(n13996) );
XNOR2_X2 U9268 ( .A(n17039), .B(z_out[120]), .ZN(n13998) );
NAND2_X2 U9269 ( .A1(n17946), .A2(Out_data[120]), .ZN(n13995) );
NAND2_X2 U9271 ( .A1(n14002), .A2(n17841), .ZN(n14000) );
XNOR2_X2 U9272 ( .A(n17037), .B(z_out[121]), .ZN(n14002) );
NAND2_X2 U9273 ( .A1(n17946), .A2(Out_data[121]), .ZN(n13999) );
NAND2_X2 U9275 ( .A1(n14006), .A2(n17841), .ZN(n14004) );
XNOR2_X2 U9276 ( .A(n17035), .B(z_out[122]), .ZN(n14006) );
NAND2_X2 U9277 ( .A1(n17946), .A2(Out_data[122]), .ZN(n14003) );
NAND2_X2 U9279 ( .A1(n14010), .A2(n17841), .ZN(n14008) );
XNOR2_X2 U9280 ( .A(n17033), .B(z_out[123]), .ZN(n14010) );
NAND2_X2 U9281 ( .A1(n17946), .A2(Out_data[123]), .ZN(n14007) );
NAND2_X2 U9283 ( .A1(n14014), .A2(n17841), .ZN(n14012) );
XNOR2_X2 U9284 ( .A(n17031), .B(z_out[124]), .ZN(n14014) );
NAND2_X2 U9285 ( .A1(n17946), .A2(Out_data[124]), .ZN(n14011) );
NAND2_X2 U9287 ( .A1(n14018), .A2(n17841), .ZN(n14016) );
XNOR2_X2 U9288 ( .A(n17029), .B(z_out[125]), .ZN(n14018) );
NAND2_X2 U9289 ( .A1(n17946), .A2(Out_data[125]), .ZN(n14015) );
NAND2_X2 U9291 ( .A1(n14022), .A2(n17841), .ZN(n14020) );
XNOR2_X2 U9292 ( .A(n17027), .B(z_out[126]), .ZN(n14022) );
NAND2_X2 U9293 ( .A1(n17946), .A2(Out_data[126]), .ZN(n14019) );
NAND2_X2 U9295 ( .A1(n14026), .A2(n17841), .ZN(n14024) );
XNOR2_X2 U9296 ( .A(n17025), .B(z_out[127]), .ZN(n14026) );
NAND2_X2 U9297 ( .A1(n17946), .A2(Out_data[127]), .ZN(n14023) );
AND4_X2 U9301 ( .A1(state[9]), .A2(n18845), .A3(n18601), .A4(n18079), .ZN(n11955) );
NAND2_X2 U9622 ( .A1(n18014), .A2(n17747), .ZN(aes_kld) );
AND4_X2 U9624 ( .A1(n18078), .A2(n18629), .A3(n18630), .A4(n14155), .ZN(n11971) );
NAND2_X2 U9631 ( .A1(n14158), .A2(n14159), .ZN(N3198) );
NAND2_X2 U9632 ( .A1(n14160), .A2(n18064), .ZN(n14159) );
XNOR2_X2 U9633 ( .A(n17024), .B(n14161), .ZN(n14160) );
NAND4_X2 U9634 ( .A1(n14025), .A2(n14162), .A3(n14163), .A4(n14164), .ZN(n14161) );
NAND2_X2 U9635 ( .A1(n17916), .A2(n14166), .ZN(n14164) );
NAND2_X2 U9636 ( .A1(n17906), .A2(dii_data[127]), .ZN(n14163) );
AND2_X2 U9638 ( .A1(n14168), .A2(n14169), .ZN(n14025) );
NAND2_X2 U9639 ( .A1(n14170), .A2(n18748), .ZN(n14169) );
NAND2_X2 U9640 ( .A1(n14171), .A2(n14172), .ZN(n14170) );
NAND2_X2 U9641 ( .A1(n17935), .A2(n14166), .ZN(n14172) );
NAND2_X2 U9642 ( .A1(n17288), .A2(dii_data[127]), .ZN(n14171) );
NAND2_X2 U9643 ( .A1(aes_text_out[127]), .A2(n14173), .ZN(n14168) );
NAND2_X2 U9644 ( .A1(n14174), .A2(n14175), .ZN(n14173) );
NAND2_X2 U9645 ( .A1(n19023), .A2(n17944), .ZN(n14175) );
NAND4_X2 U9646 ( .A1(n14176), .A2(n14177), .A3(n14178), .A4(n14179), .ZN(n14166) );
NAND2_X2 U9655 ( .A1(n17877), .A2(dii_data[95]), .ZN(n14177) );
NAND2_X2 U9656 ( .A1(n17849), .A2(dii_data[119]), .ZN(n14176) );
OR2_X2 U9657 ( .A1(n17932), .A2(dii_data[127]), .ZN(n14174) );
NAND2_X2 U9658 ( .A1(n18037), .A2(b_in[111]), .ZN(n14158) );
NAND2_X2 U9659 ( .A1(n14192), .A2(n14193), .ZN(N3197) );
NAND2_X2 U9660 ( .A1(n14194), .A2(n18064), .ZN(n14193) );
XNOR2_X2 U9661 ( .A(n17026), .B(n14195), .ZN(n14194) );
NAND4_X2 U9662 ( .A1(n14021), .A2(n14196), .A3(n14197), .A4(n14198), .ZN(n14195) );
NAND2_X2 U9663 ( .A1(n17916), .A2(n14199), .ZN(n14198) );
NAND2_X2 U9664 ( .A1(n17906), .A2(dii_data[126]), .ZN(n14197) );
AND2_X2 U9666 ( .A1(n14200), .A2(n14201), .ZN(n14021) );
NAND2_X2 U9667 ( .A1(n14202), .A2(n18749), .ZN(n14201) );
NAND2_X2 U9668 ( .A1(n14203), .A2(n14204), .ZN(n14202) );
NAND2_X2 U9669 ( .A1(n17935), .A2(n14199), .ZN(n14204) );
NAND2_X2 U9670 ( .A1(n17288), .A2(dii_data[126]), .ZN(n14203) );
NAND2_X2 U9671 ( .A1(aes_text_out[126]), .A2(n14205), .ZN(n14200) );
NAND2_X2 U9672 ( .A1(n14206), .A2(n14207), .ZN(n14205) );
NAND2_X2 U9673 ( .A1(n19024), .A2(n17944), .ZN(n14207) );
NAND4_X2 U9674 ( .A1(n14208), .A2(n14209), .A3(n14210), .A4(n14211), .ZN(n14199) );
NAND2_X2 U9683 ( .A1(n17873), .A2(dii_data[94]), .ZN(n14209) );
NAND2_X2 U9684 ( .A1(n17848), .A2(dii_data[118]), .ZN(n14208) );
OR2_X2 U9685 ( .A1(n17932), .A2(dii_data[126]), .ZN(n14206) );
NAND2_X2 U9686 ( .A1(n18043), .A2(b_in[110]), .ZN(n14192) );
NAND2_X2 U9687 ( .A1(n14221), .A2(n14222), .ZN(N3196) );
NAND2_X2 U9688 ( .A1(n14223), .A2(n18064), .ZN(n14222) );
XNOR2_X2 U9689 ( .A(n17028), .B(n14224), .ZN(n14223) );
NAND4_X2 U9690 ( .A1(n14017), .A2(n14225), .A3(n14226), .A4(n14227), .ZN(n14224) );
NAND2_X2 U9691 ( .A1(n17916), .A2(n14228), .ZN(n14227) );
NAND2_X2 U9692 ( .A1(n17906), .A2(dii_data[125]), .ZN(n14226) );
AND2_X2 U9694 ( .A1(n14229), .A2(n14230), .ZN(n14017) );
NAND2_X2 U9695 ( .A1(n14231), .A2(n18750), .ZN(n14230) );
NAND2_X2 U9696 ( .A1(n14232), .A2(n14233), .ZN(n14231) );
NAND2_X2 U9697 ( .A1(n17935), .A2(n14228), .ZN(n14233) );
NAND2_X2 U9698 ( .A1(n17288), .A2(dii_data[125]), .ZN(n14232) );
NAND2_X2 U9699 ( .A1(aes_text_out[125]), .A2(n14234), .ZN(n14229) );
NAND2_X2 U9700 ( .A1(n14235), .A2(n14236), .ZN(n14234) );
NAND2_X2 U9701 ( .A1(n19025), .A2(n17944), .ZN(n14236) );
NAND4_X2 U9702 ( .A1(n14237), .A2(n14238), .A3(n14239), .A4(n14240), .ZN(n14228) );
NAND2_X2 U9711 ( .A1(n17873), .A2(dii_data[93]), .ZN(n14238) );
NAND2_X2 U9712 ( .A1(n17848), .A2(dii_data[117]), .ZN(n14237) );
OR2_X2 U9713 ( .A1(n17932), .A2(dii_data[125]), .ZN(n14235) );
NAND2_X2 U9714 ( .A1(n18043), .A2(b_in[109]), .ZN(n14221) );
NAND2_X2 U9715 ( .A1(n14250), .A2(n14251), .ZN(N3195) );
NAND2_X2 U9716 ( .A1(n14252), .A2(n18064), .ZN(n14251) );
XNOR2_X2 U9717 ( .A(n17030), .B(n14253), .ZN(n14252) );
NAND4_X2 U9718 ( .A1(n14013), .A2(n14254), .A3(n14255), .A4(n14256), .ZN(n14253) );
NAND2_X2 U9719 ( .A1(n17916), .A2(n14257), .ZN(n14256) );
NAND2_X2 U9720 ( .A1(n17906), .A2(dii_data[124]), .ZN(n14255) );
AND2_X2 U9722 ( .A1(n14258), .A2(n14259), .ZN(n14013) );
NAND2_X2 U9723 ( .A1(n14260), .A2(n18751), .ZN(n14259) );
NAND2_X2 U9724 ( .A1(n14261), .A2(n14262), .ZN(n14260) );
NAND2_X2 U9725 ( .A1(n17935), .A2(n14257), .ZN(n14262) );
NAND2_X2 U9726 ( .A1(n17288), .A2(dii_data[124]), .ZN(n14261) );
NAND2_X2 U9727 ( .A1(aes_text_out[124]), .A2(n14263), .ZN(n14258) );
NAND2_X2 U9728 ( .A1(n14264), .A2(n14265), .ZN(n14263) );
NAND2_X2 U9729 ( .A1(n19026), .A2(n17945), .ZN(n14265) );
NAND4_X2 U9730 ( .A1(n14266), .A2(n14267), .A3(n14268), .A4(n14269), .ZN(n14257) );
NAND2_X2 U9739 ( .A1(n17873), .A2(dii_data[92]), .ZN(n14267) );
NAND2_X2 U9740 ( .A1(n17848), .A2(dii_data[116]), .ZN(n14266) );
OR2_X2 U9741 ( .A1(n17932), .A2(dii_data[124]), .ZN(n14264) );
NAND2_X2 U9742 ( .A1(n18043), .A2(b_in[108]), .ZN(n14250) );
NAND2_X2 U9743 ( .A1(n14279), .A2(n14280), .ZN(N3194) );
NAND2_X2 U9744 ( .A1(n14281), .A2(n18064), .ZN(n14280) );
XNOR2_X2 U9745 ( .A(n17032), .B(n14282), .ZN(n14281) );
NAND4_X2 U9746 ( .A1(n14009), .A2(n14283), .A3(n14284), .A4(n14285), .ZN(n14282) );
NAND2_X2 U9747 ( .A1(n17915), .A2(n14286), .ZN(n14285) );
NAND2_X2 U9748 ( .A1(n17906), .A2(dii_data[123]), .ZN(n14284) );
AND2_X2 U9750 ( .A1(n14287), .A2(n14288), .ZN(n14009) );
NAND2_X2 U9751 ( .A1(n14289), .A2(n18752), .ZN(n14288) );
NAND2_X2 U9752 ( .A1(n14290), .A2(n14291), .ZN(n14289) );
NAND2_X2 U9753 ( .A1(n17935), .A2(n14286), .ZN(n14291) );
NAND2_X2 U9754 ( .A1(n17288), .A2(dii_data[123]), .ZN(n14290) );
NAND2_X2 U9755 ( .A1(aes_text_out[123]), .A2(n14292), .ZN(n14287) );
NAND2_X2 U9756 ( .A1(n14293), .A2(n14294), .ZN(n14292) );
NAND2_X2 U9757 ( .A1(n19027), .A2(n17945), .ZN(n14294) );
NAND4_X2 U9758 ( .A1(n14295), .A2(n14296), .A3(n14297), .A4(n14298), .ZN(n14286) );
NAND2_X2 U9767 ( .A1(n17873), .A2(dii_data[91]), .ZN(n14296) );
NAND2_X2 U9768 ( .A1(n17848), .A2(dii_data[115]), .ZN(n14295) );
OR2_X2 U9769 ( .A1(n17932), .A2(dii_data[123]), .ZN(n14293) );
NAND2_X2 U9770 ( .A1(n18043), .A2(b_in[107]), .ZN(n14279) );
NAND2_X2 U9771 ( .A1(n14308), .A2(n14309), .ZN(N3193) );
NAND2_X2 U9772 ( .A1(n14310), .A2(n18064), .ZN(n14309) );
XNOR2_X2 U9773 ( .A(n17034), .B(n14311), .ZN(n14310) );
NAND4_X2 U9774 ( .A1(n14005), .A2(n14312), .A3(n14313), .A4(n14314), .ZN(n14311) );
NAND2_X2 U9775 ( .A1(n17915), .A2(n14315), .ZN(n14314) );
NAND2_X2 U9776 ( .A1(n17906), .A2(dii_data[122]), .ZN(n14313) );
AND2_X2 U9778 ( .A1(n14316), .A2(n14317), .ZN(n14005) );
NAND2_X2 U9779 ( .A1(n14318), .A2(n18753), .ZN(n14317) );
NAND2_X2 U9780 ( .A1(n14319), .A2(n14320), .ZN(n14318) );
NAND2_X2 U9781 ( .A1(n17935), .A2(n14315), .ZN(n14320) );
NAND2_X2 U9782 ( .A1(n17288), .A2(dii_data[122]), .ZN(n14319) );
NAND2_X2 U9783 ( .A1(aes_text_out[122]), .A2(n14321), .ZN(n14316) );
NAND2_X2 U9784 ( .A1(n14322), .A2(n14323), .ZN(n14321) );
NAND2_X2 U9785 ( .A1(n19028), .A2(n17945), .ZN(n14323) );
NAND4_X2 U9786 ( .A1(n14324), .A2(n14325), .A3(n14326), .A4(n14327), .ZN(n14315) );
NAND2_X2 U9795 ( .A1(n17873), .A2(dii_data[90]), .ZN(n14325) );
NAND2_X2 U9796 ( .A1(n17848), .A2(dii_data[114]), .ZN(n14324) );
OR2_X2 U9797 ( .A1(n17932), .A2(dii_data[122]), .ZN(n14322) );
NAND2_X2 U9798 ( .A1(n18043), .A2(b_in[106]), .ZN(n14308) );
NAND2_X2 U9799 ( .A1(n14337), .A2(n14338), .ZN(N3192) );
NAND2_X2 U9800 ( .A1(n14339), .A2(n18064), .ZN(n14338) );
XNOR2_X2 U9801 ( .A(n17036), .B(n14340), .ZN(n14339) );
NAND4_X2 U9802 ( .A1(n14001), .A2(n14341), .A3(n14342), .A4(n14343), .ZN(n14340) );
NAND2_X2 U9803 ( .A1(n17915), .A2(n14344), .ZN(n14343) );
NAND2_X2 U9804 ( .A1(n17906), .A2(dii_data[121]), .ZN(n14342) );
AND2_X2 U9806 ( .A1(n14345), .A2(n14346), .ZN(n14001) );
NAND2_X2 U9807 ( .A1(n14347), .A2(n18754), .ZN(n14346) );
NAND2_X2 U9808 ( .A1(n14348), .A2(n14349), .ZN(n14347) );
NAND2_X2 U9809 ( .A1(n17935), .A2(n14344), .ZN(n14349) );
NAND2_X2 U9810 ( .A1(n17288), .A2(dii_data[121]), .ZN(n14348) );
NAND2_X2 U9811 ( .A1(aes_text_out[121]), .A2(n14350), .ZN(n14345) );
NAND2_X2 U9812 ( .A1(n14351), .A2(n14352), .ZN(n14350) );
NAND2_X2 U9813 ( .A1(n19029), .A2(n17945), .ZN(n14352) );
NAND4_X2 U9814 ( .A1(n14353), .A2(n14354), .A3(n14355), .A4(n14356), .ZN(n14344) );
NAND2_X2 U9823 ( .A1(n17873), .A2(dii_data[89]), .ZN(n14354) );
NAND2_X2 U9824 ( .A1(n17848), .A2(dii_data[113]), .ZN(n14353) );
OR2_X2 U9825 ( .A1(n17932), .A2(dii_data[121]), .ZN(n14351) );
NAND2_X2 U9826 ( .A1(n18043), .A2(b_in[105]), .ZN(n14337) );
NAND2_X2 U9827 ( .A1(n14366), .A2(n14367), .ZN(N3191) );
NAND2_X2 U9828 ( .A1(n14368), .A2(n18064), .ZN(n14367) );
XNOR2_X2 U9829 ( .A(n17038), .B(n14369), .ZN(n14368) );
NAND4_X2 U9830 ( .A1(n13997), .A2(n14370), .A3(n14371), .A4(n14372), .ZN(n14369) );
NAND2_X2 U9831 ( .A1(n17915), .A2(n14373), .ZN(n14372) );
NAND2_X2 U9832 ( .A1(n17907), .A2(dii_data[120]), .ZN(n14371) );
AND2_X2 U9834 ( .A1(n14374), .A2(n14375), .ZN(n13997) );
NAND2_X2 U9835 ( .A1(n14376), .A2(n18755), .ZN(n14375) );
NAND2_X2 U9836 ( .A1(n14377), .A2(n14378), .ZN(n14376) );
NAND2_X2 U9837 ( .A1(n17934), .A2(n14373), .ZN(n14378) );
NAND2_X2 U9838 ( .A1(n17288), .A2(dii_data[120]), .ZN(n14377) );
NAND2_X2 U9839 ( .A1(aes_text_out[120]), .A2(n14379), .ZN(n14374) );
NAND2_X2 U9840 ( .A1(n14380), .A2(n14381), .ZN(n14379) );
NAND2_X2 U9841 ( .A1(n19030), .A2(n17945), .ZN(n14381) );
NAND4_X2 U9842 ( .A1(n14382), .A2(n14383), .A3(n14384), .A4(n14385), .ZN(n14373) );
NAND2_X2 U9846 ( .A1(n17897), .A2(n18076), .ZN(n14184) );
NAND2_X2 U9848 ( .A1(n17892), .A2(n18072), .ZN(n14186) );
NAND2_X2 U9850 ( .A1(n14393), .A2(n17892), .ZN(n14187) );
NAND2_X2 U9854 ( .A1(n17873), .A2(dii_data[88]), .ZN(n14383) );
NAND2_X2 U9855 ( .A1(n17848), .A2(dii_data[112]), .ZN(n14382) );
OR2_X2 U9856 ( .A1(n17932), .A2(dii_data[120]), .ZN(n14380) );
NAND2_X2 U9857 ( .A1(n18043), .A2(b_in[104]), .ZN(n14366) );
NAND2_X2 U9858 ( .A1(n14398), .A2(n14399), .ZN(N3190) );
NAND2_X2 U9859 ( .A1(n14400), .A2(n18064), .ZN(n14399) );
XNOR2_X2 U9860 ( .A(n19014), .B(n14401), .ZN(n14400) );
NAND2_X2 U9862 ( .A1(n17919), .A2(n14405), .ZN(n13992) );
XOR2_X2 U9863 ( .A(n17523), .B(aes_text_out[119]), .Z(n14405) );
XNOR2_X2 U9865 ( .A(n14407), .B(aes_text_out[119]), .ZN(n13994) );
AND2_X2 U9866 ( .A1(dii_data[119]), .A2(n17908), .ZN(n14403) );
NAND2_X2 U9867 ( .A1(n14408), .A2(n14409), .ZN(n14402) );
NAND2_X2 U9869 ( .A1(n17915), .A2(n14407), .ZN(n14408) );
NAND4_X2 U9870 ( .A1(n14410), .A2(n14411), .A3(n14412), .A4(n14413), .ZN(n14407) );
NAND2_X2 U9871 ( .A1(n19047), .A2(n17890), .ZN(n14413) );
NAND2_X2 U9875 ( .A1(n19031), .A2(n17896), .ZN(n14411) );
NAND2_X2 U9877 ( .A1(n14421), .A2(n18071), .ZN(n14420) );
NAND2_X2 U9878 ( .A1(n14393), .A2(n19151), .ZN(n14419) );
NAND2_X2 U9879 ( .A1(n17882), .A2(n19032), .ZN(n14418) );
NAND2_X2 U9880 ( .A1(n19079), .A2(n17898), .ZN(n14410) );
NAND2_X2 U9881 ( .A1(n18043), .A2(b_in[103]), .ZN(n14398) );
NAND2_X2 U9882 ( .A1(n14423), .A2(n14424), .ZN(N3189) );
NAND2_X2 U9883 ( .A1(n14425), .A2(n18064), .ZN(n14424) );
XNOR2_X2 U9884 ( .A(n19013), .B(n14426), .ZN(n14425) );
NAND2_X2 U9886 ( .A1(n17919), .A2(n14430), .ZN(n13986) );
XOR2_X2 U9887 ( .A(n17525), .B(aes_text_out[118]), .Z(n14430) );
XNOR2_X2 U9889 ( .A(n14431), .B(aes_text_out[118]), .ZN(n13988) );
AND2_X2 U9890 ( .A1(dii_data[118]), .A2(n17908), .ZN(n14428) );
NAND2_X2 U9891 ( .A1(n14432), .A2(n14433), .ZN(n14427) );
NAND2_X2 U9893 ( .A1(n17915), .A2(n14431), .ZN(n14432) );
NAND4_X2 U9894 ( .A1(n14434), .A2(n14435), .A3(n14436), .A4(n14437), .ZN(n14431) );
NAND2_X2 U9895 ( .A1(n19049), .A2(n17890), .ZN(n14437) );
NAND2_X2 U9899 ( .A1(n19033), .A2(n17896), .ZN(n14435) );
NAND2_X2 U9901 ( .A1(n14444), .A2(n18071), .ZN(n14443) );
NAND2_X2 U9902 ( .A1(n14393), .A2(n19152), .ZN(n14442) );
NAND2_X2 U9903 ( .A1(n17884), .A2(n19034), .ZN(n14441) );
NAND2_X2 U9904 ( .A1(n19082), .A2(n17899), .ZN(n14434) );
NAND2_X2 U9905 ( .A1(n18043), .A2(b_in[102]), .ZN(n14423) );
NAND2_X2 U9906 ( .A1(n14445), .A2(n14446), .ZN(N3188) );
NAND2_X2 U9907 ( .A1(n14447), .A2(n18064), .ZN(n14446) );
XNOR2_X2 U9908 ( .A(n19012), .B(n14448), .ZN(n14447) );
NAND2_X2 U9910 ( .A1(n17919), .A2(n14452), .ZN(n13980) );
XOR2_X2 U9911 ( .A(n17527), .B(aes_text_out[117]), .Z(n14452) );
XNOR2_X2 U9913 ( .A(n14453), .B(aes_text_out[117]), .ZN(n13982) );
AND2_X2 U9914 ( .A1(dii_data[117]), .A2(n17908), .ZN(n14450) );
NAND2_X2 U9915 ( .A1(n14454), .A2(n14455), .ZN(n14449) );
NAND2_X2 U9917 ( .A1(n17915), .A2(n14453), .ZN(n14454) );
NAND4_X2 U9918 ( .A1(n14456), .A2(n14457), .A3(n14458), .A4(n14459), .ZN(n14453) );
NAND2_X2 U9919 ( .A1(n19051), .A2(n17890), .ZN(n14459) );
NAND2_X2 U9923 ( .A1(n19035), .A2(n17896), .ZN(n14457) );
NAND2_X2 U9925 ( .A1(n14466), .A2(n18071), .ZN(n14465) );
NAND2_X2 U9926 ( .A1(n14393), .A2(n19153), .ZN(n14464) );
NAND2_X2 U9927 ( .A1(n17884), .A2(n19036), .ZN(n14463) );
NAND2_X2 U9928 ( .A1(n19085), .A2(n17899), .ZN(n14456) );
NAND2_X2 U9929 ( .A1(n18043), .A2(b_in[101]), .ZN(n14445) );
NAND2_X2 U9930 ( .A1(n14467), .A2(n14468), .ZN(N3187) );
NAND2_X2 U9931 ( .A1(n14469), .A2(n18064), .ZN(n14468) );
XNOR2_X2 U9932 ( .A(n19011), .B(n14470), .ZN(n14469) );
NAND2_X2 U9934 ( .A1(n17919), .A2(n14474), .ZN(n13974) );
XOR2_X2 U9935 ( .A(n17529), .B(aes_text_out[116]), .Z(n14474) );
XNOR2_X2 U9937 ( .A(n14475), .B(aes_text_out[116]), .ZN(n13976) );
AND2_X2 U9938 ( .A1(dii_data[116]), .A2(n17908), .ZN(n14472) );
NAND2_X2 U9939 ( .A1(n14476), .A2(n14477), .ZN(n14471) );
NAND2_X2 U9940 ( .A1(n17998), .A2(aad_byte_cnt[49]), .ZN(n14477) );
NAND2_X2 U9941 ( .A1(n17915), .A2(n14475), .ZN(n14476) );
NAND4_X2 U9942 ( .A1(n14478), .A2(n14479), .A3(n14480), .A4(n14481), .ZN(n14475) );
NAND2_X2 U9943 ( .A1(n19053), .A2(n17890), .ZN(n14481) );
NAND2_X2 U9947 ( .A1(n19037), .A2(n17896), .ZN(n14479) );
NAND2_X2 U9949 ( .A1(n14488), .A2(n18071), .ZN(n14487) );
NAND2_X2 U9950 ( .A1(n14393), .A2(n19154), .ZN(n14486) );
NAND2_X2 U9951 ( .A1(n17884), .A2(n19038), .ZN(n14485) );
NAND2_X2 U9952 ( .A1(n19088), .A2(n17899), .ZN(n14478) );
NAND2_X2 U9953 ( .A1(n18043), .A2(b_in[100]), .ZN(n14467) );
NAND2_X2 U9954 ( .A1(n14489), .A2(n14490), .ZN(N3186) );
NAND2_X2 U9955 ( .A1(n14491), .A2(n18064), .ZN(n14490) );
XNOR2_X2 U9956 ( .A(n19010), .B(n14492), .ZN(n14491) );
NAND2_X2 U9958 ( .A1(n17919), .A2(n14496), .ZN(n13968) );
XOR2_X2 U9959 ( .A(n17531), .B(aes_text_out[115]), .Z(n14496) );
XNOR2_X2 U9961 ( .A(n14497), .B(aes_text_out[115]), .ZN(n13970) );
AND2_X2 U9962 ( .A1(dii_data[115]), .A2(n17908), .ZN(n14494) );
NAND2_X2 U9963 ( .A1(n14498), .A2(n14499), .ZN(n14493) );
NAND2_X2 U9964 ( .A1(n17996), .A2(aad_byte_cnt[48]), .ZN(n14499) );
NAND2_X2 U9965 ( .A1(n17915), .A2(n14497), .ZN(n14498) );
NAND4_X2 U9966 ( .A1(n14500), .A2(n14501), .A3(n14502), .A4(n14503), .ZN(n14497) );
NAND2_X2 U9967 ( .A1(n19055), .A2(n17890), .ZN(n14503) );
NAND2_X2 U9971 ( .A1(n19039), .A2(n17896), .ZN(n14501) );
NAND2_X2 U9973 ( .A1(n14510), .A2(n18071), .ZN(n14509) );
NAND2_X2 U9974 ( .A1(n14393), .A2(n19155), .ZN(n14508) );
NAND2_X2 U9975 ( .A1(n17884), .A2(n19040), .ZN(n14507) );
NAND2_X2 U9976 ( .A1(n19091), .A2(n17899), .ZN(n14500) );
NAND2_X2 U9977 ( .A1(n18043), .A2(b_in[99]), .ZN(n14489) );
NAND2_X2 U9978 ( .A1(n14511), .A2(n14512), .ZN(N3185) );
NAND2_X2 U9979 ( .A1(n14513), .A2(n18064), .ZN(n14512) );
XNOR2_X2 U9980 ( .A(n19009), .B(n14514), .ZN(n14513) );
NAND2_X2 U9982 ( .A1(n17919), .A2(n14518), .ZN(n13962) );
XOR2_X2 U9983 ( .A(n17533), .B(aes_text_out[114]), .Z(n14518) );
XNOR2_X2 U9985 ( .A(n14519), .B(aes_text_out[114]), .ZN(n13964) );
AND2_X2 U9986 ( .A1(dii_data[114]), .A2(n17908), .ZN(n14516) );
NAND2_X2 U9987 ( .A1(n14520), .A2(n14521), .ZN(n14515) );
NAND2_X2 U9988 ( .A1(n17996), .A2(aad_byte_cnt[47]), .ZN(n14521) );
NAND2_X2 U9989 ( .A1(n17915), .A2(n14519), .ZN(n14520) );
NAND4_X2 U9990 ( .A1(n14522), .A2(n14523), .A3(n14524), .A4(n14525), .ZN(n14519) );
NAND2_X2 U9991 ( .A1(n19057), .A2(n17890), .ZN(n14525) );
NAND2_X2 U9995 ( .A1(n19041), .A2(n17896), .ZN(n14523) );
NAND2_X2 U9997 ( .A1(n14532), .A2(n18071), .ZN(n14531) );
NAND2_X2 U9998 ( .A1(n14393), .A2(n19156), .ZN(n14530) );
NAND2_X2 U9999 ( .A1(n17884), .A2(n19042), .ZN(n14529) );
NAND2_X2 U10000 ( .A1(n19094), .A2(n17898), .ZN(n14522) );
NAND2_X2 U10001 ( .A1(n18043), .A2(b_in[98]), .ZN(n14511) );
NAND2_X2 U10002 ( .A1(n14533), .A2(n14534), .ZN(N3184) );
NAND2_X2 U10003 ( .A1(n14535), .A2(n18064), .ZN(n14534) );
XNOR2_X2 U10004 ( .A(n19008), .B(n14536), .ZN(n14535) );
NAND2_X2 U10006 ( .A1(n17919), .A2(n14540), .ZN(n13956) );
XOR2_X2 U10007 ( .A(n17535), .B(aes_text_out[113]), .Z(n14540) );
XNOR2_X2 U10009 ( .A(n14541), .B(aes_text_out[113]), .ZN(n13958) );
AND2_X2 U10010 ( .A1(dii_data[113]), .A2(n17908), .ZN(n14538) );
NAND2_X2 U10011 ( .A1(n14542), .A2(n14543), .ZN(n14537) );
NAND2_X2 U10012 ( .A1(n17996), .A2(aad_byte_cnt[46]), .ZN(n14543) );
NAND2_X2 U10013 ( .A1(n17915), .A2(n14541), .ZN(n14542) );
NAND4_X2 U10014 ( .A1(n14544), .A2(n14545), .A3(n14546), .A4(n14547), .ZN(n14541) );
NAND2_X2 U10015 ( .A1(n19059), .A2(n17889), .ZN(n14547) );
NAND2_X2 U10019 ( .A1(n19043), .A2(n17895), .ZN(n14545) );
NAND2_X2 U10021 ( .A1(n14554), .A2(n18071), .ZN(n14553) );
NAND2_X2 U10022 ( .A1(n14393), .A2(n19157), .ZN(n14552) );
NAND2_X2 U10023 ( .A1(n17884), .A2(n19044), .ZN(n14551) );
NAND2_X2 U10024 ( .A1(n19097), .A2(n17898), .ZN(n14544) );
NAND2_X2 U10025 ( .A1(n18043), .A2(b_in[97]), .ZN(n14533) );
NAND2_X2 U10026 ( .A1(n14555), .A2(n14556), .ZN(N3183) );
NAND2_X2 U10027 ( .A1(n14557), .A2(n18064), .ZN(n14556) );
XNOR2_X2 U10028 ( .A(n19007), .B(n14558), .ZN(n14557) );
NAND2_X2 U10030 ( .A1(n17919), .A2(n14562), .ZN(n13950) );
XOR2_X2 U10031 ( .A(n17537), .B(aes_text_out[112]), .Z(n14562) );
NAND2_X2 U10033 ( .A1(n17935), .A2(n14563), .ZN(n14406) );
NAND2_X2 U10034 ( .A1(n19200), .A2(n14564), .ZN(n14563) );
XNOR2_X2 U10035 ( .A(n14565), .B(aes_text_out[112]), .ZN(n13952) );
AND2_X2 U10036 ( .A1(dii_data[112]), .A2(n17908), .ZN(n14560) );
NAND2_X2 U10037 ( .A1(n14566), .A2(n14567), .ZN(n14559) );
NAND2_X2 U10038 ( .A1(n17996), .A2(aad_byte_cnt[45]), .ZN(n14567) );
NAND2_X2 U10039 ( .A1(n17914), .A2(n14565), .ZN(n14566) );
NAND4_X2 U10040 ( .A1(n14568), .A2(n14569), .A3(n14570), .A4(n14571), .ZN(n14565) );
NAND2_X2 U10041 ( .A1(n19061), .A2(n17889), .ZN(n14571) );
NAND2_X2 U10045 ( .A1(n19045), .A2(n17895), .ZN(n14569) );
NAND2_X2 U10047 ( .A1(n14578), .A2(n18071), .ZN(n14577) );
NAND2_X2 U10048 ( .A1(n14393), .A2(n19158), .ZN(n14576) );
NAND2_X2 U10049 ( .A1(n17884), .A2(n19046), .ZN(n14575) );
NAND2_X2 U10050 ( .A1(n19100), .A2(n17898), .ZN(n14568) );
NAND2_X2 U10051 ( .A1(n18043), .A2(b_in[96]), .ZN(n14555) );
NAND2_X2 U10052 ( .A1(n14579), .A2(n14580), .ZN(N3182) );
NAND2_X2 U10053 ( .A1(n14581), .A2(n18065), .ZN(n14580) );
XNOR2_X2 U10054 ( .A(n19006), .B(n14582), .ZN(n14581) );
NAND2_X2 U10056 ( .A1(n17919), .A2(n14586), .ZN(n13944) );
XNOR2_X2 U10057 ( .A(n19032), .B(aes_text_out[111]), .ZN(n14586) );
XNOR2_X2 U10059 ( .A(n14588), .B(aes_text_out[111]), .ZN(n13946) );
NAND2_X2 U10061 ( .A1(n14589), .A2(n14590), .ZN(n14583) );
NAND2_X2 U10062 ( .A1(n17996), .A2(aad_byte_cnt[44]), .ZN(n14590) );
NAND2_X2 U10063 ( .A1(n17914), .A2(n14588), .ZN(n14589) );
NAND4_X2 U10064 ( .A1(n14591), .A2(n14592), .A3(n14593), .A4(n14594), .ZN(n14588) );
NAND2_X2 U10065 ( .A1(n19063), .A2(n17889), .ZN(n14594) );
NAND2_X2 U10069 ( .A1(n19047), .A2(n17895), .ZN(n14592) );
NAND2_X2 U10071 ( .A1(n19127), .A2(n18071), .ZN(n14600) );
NAND2_X2 U10072 ( .A1(n14393), .A2(n19159), .ZN(n14599) );
NAND2_X2 U10073 ( .A1(n17884), .A2(n19048), .ZN(n14598) );
NAND2_X2 U10074 ( .A1(n19103), .A2(n17898), .ZN(n14591) );
NAND2_X2 U10075 ( .A1(n18043), .A2(b_in[95]), .ZN(n14579) );
NAND2_X2 U10076 ( .A1(n14601), .A2(n14602), .ZN(N3181) );
NAND2_X2 U10077 ( .A1(n14603), .A2(n18065), .ZN(n14602) );
XNOR2_X2 U10078 ( .A(n19005), .B(n14604), .ZN(n14603) );
NAND2_X2 U10080 ( .A1(n17919), .A2(n14608), .ZN(n13938) );
XNOR2_X2 U10081 ( .A(n19034), .B(aes_text_out[110]), .ZN(n14608) );
XNOR2_X2 U10083 ( .A(n14609), .B(aes_text_out[110]), .ZN(n13940) );
NAND2_X2 U10085 ( .A1(n14610), .A2(n14611), .ZN(n14605) );
NAND2_X2 U10086 ( .A1(n17996), .A2(aad_byte_cnt[43]), .ZN(n14611) );
NAND2_X2 U10087 ( .A1(n17914), .A2(n14609), .ZN(n14610) );
NAND4_X2 U10088 ( .A1(n14612), .A2(n14613), .A3(n14614), .A4(n14615), .ZN(n14609) );
NAND2_X2 U10089 ( .A1(n19065), .A2(n17889), .ZN(n14615) );
NAND2_X2 U10093 ( .A1(n19049), .A2(n17895), .ZN(n14613) );
NAND2_X2 U10095 ( .A1(n19128), .A2(n18071), .ZN(n14621) );
NAND2_X2 U10096 ( .A1(n14393), .A2(n19160), .ZN(n14620) );
NAND2_X2 U10097 ( .A1(n17884), .A2(n19050), .ZN(n14619) );
NAND2_X2 U10098 ( .A1(n19106), .A2(n17898), .ZN(n14612) );
NAND2_X2 U10099 ( .A1(n18042), .A2(b_in[94]), .ZN(n14601) );
NAND2_X2 U10100 ( .A1(n14622), .A2(n14623), .ZN(N3180) );
NAND2_X2 U10101 ( .A1(n14624), .A2(n18065), .ZN(n14623) );
XNOR2_X2 U10102 ( .A(n19004), .B(n14625), .ZN(n14624) );
NAND2_X2 U10104 ( .A1(n17919), .A2(n14629), .ZN(n13932) );
XNOR2_X2 U10105 ( .A(n19036), .B(aes_text_out[109]), .ZN(n14629) );
XNOR2_X2 U10107 ( .A(n14630), .B(aes_text_out[109]), .ZN(n13934) );
NAND2_X2 U10109 ( .A1(n14631), .A2(n14632), .ZN(n14626) );
NAND2_X2 U10110 ( .A1(n17996), .A2(aad_byte_cnt[42]), .ZN(n14632) );
NAND2_X2 U10111 ( .A1(n17914), .A2(n14630), .ZN(n14631) );
NAND4_X2 U10112 ( .A1(n14633), .A2(n14634), .A3(n14635), .A4(n14636), .ZN(n14630) );
NAND2_X2 U10113 ( .A1(n19067), .A2(n17889), .ZN(n14636) );
NAND2_X2 U10117 ( .A1(n19051), .A2(n17895), .ZN(n14634) );
NAND2_X2 U10119 ( .A1(n19129), .A2(n18071), .ZN(n14642) );
NAND2_X2 U10120 ( .A1(n14393), .A2(n19161), .ZN(n14641) );
NAND2_X2 U10121 ( .A1(n17884), .A2(n19052), .ZN(n14640) );
NAND2_X2 U10122 ( .A1(n19109), .A2(n17898), .ZN(n14633) );
NAND2_X2 U10123 ( .A1(n18042), .A2(b_in[93]), .ZN(n14622) );
NAND2_X2 U10124 ( .A1(n14643), .A2(n14644), .ZN(N3179) );
NAND2_X2 U10125 ( .A1(n14645), .A2(n18065), .ZN(n14644) );
XNOR2_X2 U10126 ( .A(n19003), .B(n14646), .ZN(n14645) );
NAND2_X2 U10128 ( .A1(n17920), .A2(n14650), .ZN(n13926) );
XNOR2_X2 U10129 ( .A(n19038), .B(aes_text_out[108]), .ZN(n14650) );
XNOR2_X2 U10131 ( .A(n14651), .B(aes_text_out[108]), .ZN(n13928) );
NAND2_X2 U10133 ( .A1(n14652), .A2(n14653), .ZN(n14647) );
NAND2_X2 U10134 ( .A1(n17996), .A2(aad_byte_cnt[41]), .ZN(n14653) );
NAND2_X2 U10135 ( .A1(n17914), .A2(n14651), .ZN(n14652) );
NAND4_X2 U10136 ( .A1(n14654), .A2(n14655), .A3(n14656), .A4(n14657), .ZN(n14651) );
NAND2_X2 U10137 ( .A1(n19069), .A2(n17889), .ZN(n14657) );
NAND2_X2 U10141 ( .A1(n19053), .A2(n17895), .ZN(n14655) );
NAND2_X2 U10143 ( .A1(n19130), .A2(n18071), .ZN(n14663) );
NAND2_X2 U10144 ( .A1(n14393), .A2(n19162), .ZN(n14662) );
NAND2_X2 U10145 ( .A1(n17884), .A2(n19054), .ZN(n14661) );
NAND2_X2 U10146 ( .A1(n19112), .A2(n17898), .ZN(n14654) );
NAND2_X2 U10147 ( .A1(n18042), .A2(b_in[92]), .ZN(n14643) );
NAND2_X2 U10148 ( .A1(n14664), .A2(n14665), .ZN(N3178) );
NAND2_X2 U10149 ( .A1(n14666), .A2(n18065), .ZN(n14665) );
XNOR2_X2 U10150 ( .A(n19002), .B(n14667), .ZN(n14666) );
NAND2_X2 U10152 ( .A1(n17920), .A2(n14671), .ZN(n13920) );
XNOR2_X2 U10153 ( .A(n19040), .B(aes_text_out[107]), .ZN(n14671) );
XNOR2_X2 U10155 ( .A(n14672), .B(aes_text_out[107]), .ZN(n13922) );
NAND2_X2 U10157 ( .A1(n14673), .A2(n14674), .ZN(n14668) );
NAND2_X2 U10158 ( .A1(n17996), .A2(aad_byte_cnt[40]), .ZN(n14674) );
NAND2_X2 U10159 ( .A1(n17914), .A2(n14672), .ZN(n14673) );
NAND4_X2 U10160 ( .A1(n14675), .A2(n14676), .A3(n14677), .A4(n14678), .ZN(n14672) );
NAND2_X2 U10161 ( .A1(n19071), .A2(n17889), .ZN(n14678) );
NAND2_X2 U10165 ( .A1(n19055), .A2(n17895), .ZN(n14676) );
NAND2_X2 U10167 ( .A1(n19131), .A2(n18072), .ZN(n14684) );
NAND2_X2 U10168 ( .A1(n14393), .A2(n19163), .ZN(n14683) );
NAND2_X2 U10169 ( .A1(n17883), .A2(n19056), .ZN(n14682) );
NAND2_X2 U10170 ( .A1(n19115), .A2(n17898), .ZN(n14675) );
NAND2_X2 U10171 ( .A1(n18042), .A2(b_in[91]), .ZN(n14664) );
NAND2_X2 U10172 ( .A1(n14685), .A2(n14686), .ZN(N3177) );
NAND2_X2 U10173 ( .A1(n14687), .A2(n18065), .ZN(n14686) );
XNOR2_X2 U10174 ( .A(n19001), .B(n14688), .ZN(n14687) );
NAND2_X2 U10176 ( .A1(n17920), .A2(n14692), .ZN(n13914) );
XNOR2_X2 U10177 ( .A(n19042), .B(aes_text_out[106]), .ZN(n14692) );
XNOR2_X2 U10179 ( .A(n14693), .B(aes_text_out[106]), .ZN(n13916) );
NAND2_X2 U10181 ( .A1(n14694), .A2(n14695), .ZN(n14689) );
NAND2_X2 U10182 ( .A1(n17996), .A2(aad_byte_cnt[39]), .ZN(n14695) );
NAND2_X2 U10183 ( .A1(n17914), .A2(n14693), .ZN(n14694) );
NAND4_X2 U10184 ( .A1(n14696), .A2(n14697), .A3(n14698), .A4(n14699), .ZN(n14693) );
NAND2_X2 U10185 ( .A1(n19073), .A2(n17889), .ZN(n14699) );
NAND2_X2 U10189 ( .A1(n19057), .A2(n17895), .ZN(n14697) );
NAND2_X2 U10191 ( .A1(n19132), .A2(n18071), .ZN(n14705) );
NAND2_X2 U10192 ( .A1(n14393), .A2(n19164), .ZN(n14704) );
NAND2_X2 U10193 ( .A1(n17883), .A2(n19058), .ZN(n14703) );
NAND2_X2 U10194 ( .A1(n19118), .A2(n17898), .ZN(n14696) );
NAND2_X2 U10195 ( .A1(n18042), .A2(b_in[90]), .ZN(n14685) );
NAND2_X2 U10196 ( .A1(n14706), .A2(n14707), .ZN(N3176) );
NAND2_X2 U10197 ( .A1(n14708), .A2(n18065), .ZN(n14707) );
XNOR2_X2 U10198 ( .A(n19000), .B(n14709), .ZN(n14708) );
NAND2_X2 U10200 ( .A1(n17920), .A2(n14713), .ZN(n13908) );
XNOR2_X2 U10201 ( .A(n19044), .B(aes_text_out[105]), .ZN(n14713) );
XNOR2_X2 U10203 ( .A(n14714), .B(aes_text_out[105]), .ZN(n13910) );
NAND2_X2 U10205 ( .A1(n14715), .A2(n14716), .ZN(n14710) );
NAND2_X2 U10206 ( .A1(n17996), .A2(aad_byte_cnt[38]), .ZN(n14716) );
NAND2_X2 U10207 ( .A1(n17914), .A2(n14714), .ZN(n14715) );
NAND4_X2 U10208 ( .A1(n14717), .A2(n14718), .A3(n14719), .A4(n14720), .ZN(n14714) );
NAND2_X2 U10209 ( .A1(n19075), .A2(n17889), .ZN(n14720) );
NAND2_X2 U10213 ( .A1(n19059), .A2(n17895), .ZN(n14718) );
NAND2_X2 U10215 ( .A1(n19133), .A2(n18071), .ZN(n14726) );
NAND2_X2 U10216 ( .A1(n14393), .A2(n19165), .ZN(n14725) );
NAND2_X2 U10217 ( .A1(n17883), .A2(n19060), .ZN(n14724) );
NAND2_X2 U10218 ( .A1(n19121), .A2(n17898), .ZN(n14717) );
NAND2_X2 U10219 ( .A1(n18042), .A2(b_in[89]), .ZN(n14706) );
NAND2_X2 U10220 ( .A1(n14727), .A2(n14728), .ZN(N3175) );
NAND2_X2 U10221 ( .A1(n14729), .A2(n18065), .ZN(n14728) );
XNOR2_X2 U10222 ( .A(n18999), .B(n14730), .ZN(n14729) );
NAND2_X2 U10224 ( .A1(n17920), .A2(n14734), .ZN(n13902) );
XNOR2_X2 U10225 ( .A(n19046), .B(aes_text_out[104]), .ZN(n14734) );
NAND2_X2 U10227 ( .A1(n17934), .A2(n14735), .ZN(n14587) );
NAND2_X2 U10228 ( .A1(n19200), .A2(n19204), .ZN(n14735) );
XNOR2_X2 U10229 ( .A(n14737), .B(aes_text_out[104]), .ZN(n13904) );
NAND2_X2 U10231 ( .A1(n14738), .A2(n14739), .ZN(n14731) );
NAND2_X2 U10232 ( .A1(n17996), .A2(aad_byte_cnt[37]), .ZN(n14739) );
NAND2_X2 U10233 ( .A1(n17914), .A2(n14737), .ZN(n14738) );
NAND4_X2 U10234 ( .A1(n14740), .A2(n14741), .A3(n14742), .A4(n14743), .ZN(n14737) );
NAND2_X2 U10235 ( .A1(n19077), .A2(n17889), .ZN(n14743) );
NAND2_X2 U10239 ( .A1(n19061), .A2(n17895), .ZN(n14741) );
NAND2_X2 U10241 ( .A1(n19134), .A2(n18071), .ZN(n14749) );
NAND2_X2 U10242 ( .A1(n14393), .A2(n19166), .ZN(n14748) );
NAND2_X2 U10244 ( .A1(n17883), .A2(n19062), .ZN(n14747) );
NAND2_X2 U10245 ( .A1(n19124), .A2(n17898), .ZN(n14740) );
NAND2_X2 U10246 ( .A1(n18042), .A2(b_in[88]), .ZN(n14727) );
NAND2_X2 U10247 ( .A1(n14750), .A2(n14751), .ZN(N3174) );
NAND2_X2 U10248 ( .A1(n14752), .A2(n18065), .ZN(n14751) );
XNOR2_X2 U10249 ( .A(n18998), .B(n14753), .ZN(n14752) );
NAND2_X2 U10251 ( .A1(n17920), .A2(n14757), .ZN(n13896) );
XNOR2_X2 U10252 ( .A(n19048), .B(aes_text_out[103]), .ZN(n14757) );
XNOR2_X2 U10254 ( .A(n14759), .B(aes_text_out[103]), .ZN(n13898) );
NAND2_X2 U10256 ( .A1(n14760), .A2(n14761), .ZN(n14754) );
NAND2_X2 U10257 ( .A1(n17996), .A2(aad_byte_cnt[36]), .ZN(n14761) );
NAND2_X2 U10258 ( .A1(n17914), .A2(n14759), .ZN(n14760) );
NAND4_X2 U10259 ( .A1(n14762), .A2(n14763), .A3(n14764), .A4(n14765), .ZN(n14759) );
NAND2_X2 U10260 ( .A1(n19080), .A2(n17889), .ZN(n14765) );
NAND2_X2 U10264 ( .A1(n19063), .A2(n17895), .ZN(n14763) );
NAND4_X2 U10265 ( .A1(n14769), .A2(n14770), .A3(n14771), .A4(n17881), .ZN(n14417) );
NAND2_X2 U10266 ( .A1(n17883), .A2(n19064), .ZN(n14771) );
NAND2_X2 U10267 ( .A1(n19167), .A2(n18076), .ZN(n14770) );
NAND2_X2 U10268 ( .A1(n19135), .A2(n18071), .ZN(n14769) );
NAND2_X2 U10269 ( .A1(n17897), .A2(n14773), .ZN(n14762) );
NAND2_X2 U10270 ( .A1(n18042), .A2(b_in[87]), .ZN(n14750) );
NAND2_X2 U10271 ( .A1(n14774), .A2(n14775), .ZN(N3173) );
NAND2_X2 U10272 ( .A1(n14776), .A2(n18065), .ZN(n14775) );
XNOR2_X2 U10273 ( .A(n18997), .B(n14777), .ZN(n14776) );
NAND2_X2 U10275 ( .A1(n17920), .A2(n14781), .ZN(n13890) );
XNOR2_X2 U10276 ( .A(n19050), .B(aes_text_out[102]), .ZN(n14781) );
XNOR2_X2 U10278 ( .A(n14782), .B(aes_text_out[102]), .ZN(n13892) );
NAND2_X2 U10280 ( .A1(n14783), .A2(n14784), .ZN(n14778) );
NAND2_X2 U10281 ( .A1(n17996), .A2(aad_byte_cnt[35]), .ZN(n14784) );
NAND2_X2 U10282 ( .A1(n17914), .A2(n14782), .ZN(n14783) );
NAND4_X2 U10283 ( .A1(n14785), .A2(n14786), .A3(n14787), .A4(n14788), .ZN(n14782) );
NAND2_X2 U10284 ( .A1(n19083), .A2(n17889), .ZN(n14788) );
NAND2_X2 U10288 ( .A1(n19065), .A2(n17895), .ZN(n14786) );
NAND4_X2 U10289 ( .A1(n14792), .A2(n14793), .A3(n14794), .A4(n17881), .ZN(n14440) );
NAND2_X2 U10290 ( .A1(n17883), .A2(n19066), .ZN(n14794) );
NAND2_X2 U10291 ( .A1(n19168), .A2(n18076), .ZN(n14793) );
NAND2_X2 U10292 ( .A1(n19136), .A2(n18072), .ZN(n14792) );
NAND2_X2 U10293 ( .A1(n17897), .A2(n14795), .ZN(n14785) );
NAND2_X2 U10294 ( .A1(n18042), .A2(b_in[86]), .ZN(n14774) );
NAND2_X2 U10295 ( .A1(n14796), .A2(n14797), .ZN(N3172) );
NAND2_X2 U10296 ( .A1(n14798), .A2(n18065), .ZN(n14797) );
XNOR2_X2 U10297 ( .A(n18996), .B(n14799), .ZN(n14798) );
NAND2_X2 U10299 ( .A1(n17920), .A2(n14803), .ZN(n13884) );
XNOR2_X2 U10300 ( .A(n19052), .B(aes_text_out[101]), .ZN(n14803) );
XNOR2_X2 U10302 ( .A(n14804), .B(aes_text_out[101]), .ZN(n13886) );
NAND2_X2 U10304 ( .A1(n14805), .A2(n14806), .ZN(n14800) );
NAND2_X2 U10305 ( .A1(n17997), .A2(aad_byte_cnt[34]), .ZN(n14806) );
NAND2_X2 U10306 ( .A1(n17913), .A2(n14804), .ZN(n14805) );
NAND4_X2 U10307 ( .A1(n14807), .A2(n14808), .A3(n14809), .A4(n14810), .ZN(n14804) );
NAND2_X2 U10308 ( .A1(n19086), .A2(n17888), .ZN(n14810) );
NAND2_X2 U10312 ( .A1(n19067), .A2(n17894), .ZN(n14808) );
NAND4_X2 U10313 ( .A1(n14814), .A2(n14815), .A3(n14816), .A4(n17881), .ZN(n14462) );
NAND2_X2 U10314 ( .A1(n17883), .A2(n19068), .ZN(n14816) );
NAND2_X2 U10315 ( .A1(n19169), .A2(n18076), .ZN(n14815) );
NAND2_X2 U10316 ( .A1(n19137), .A2(n18072), .ZN(n14814) );
NAND2_X2 U10317 ( .A1(n17897), .A2(n14817), .ZN(n14807) );
NAND2_X2 U10318 ( .A1(n18042), .A2(b_in[85]), .ZN(n14796) );
NAND2_X2 U10319 ( .A1(n14818), .A2(n14819), .ZN(N3171) );
NAND2_X2 U10320 ( .A1(n14820), .A2(n18065), .ZN(n14819) );
XNOR2_X2 U10321 ( .A(n18995), .B(n14821), .ZN(n14820) );
NAND2_X2 U10323 ( .A1(n17920), .A2(n14825), .ZN(n13878) );
XNOR2_X2 U10324 ( .A(n19054), .B(aes_text_out[100]), .ZN(n14825) );
XNOR2_X2 U10326 ( .A(n14826), .B(aes_text_out[100]), .ZN(n13880) );
NAND2_X2 U10328 ( .A1(n14827), .A2(n14828), .ZN(n14822) );
NAND2_X2 U10329 ( .A1(n17996), .A2(aad_byte_cnt[33]), .ZN(n14828) );
NAND2_X2 U10330 ( .A1(n17913), .A2(n14826), .ZN(n14827) );
NAND4_X2 U10331 ( .A1(n14829), .A2(n14830), .A3(n14831), .A4(n14832), .ZN(n14826) );
NAND2_X2 U10332 ( .A1(n19089), .A2(n17888), .ZN(n14832) );
NAND2_X2 U10336 ( .A1(n19069), .A2(n17894), .ZN(n14830) );
NAND4_X2 U10337 ( .A1(n14836), .A2(n14837), .A3(n14838), .A4(n17881), .ZN(n14484) );
NAND2_X2 U10338 ( .A1(n17883), .A2(n19070), .ZN(n14838) );
NAND2_X2 U10339 ( .A1(n19170), .A2(n18076), .ZN(n14837) );
NAND2_X2 U10340 ( .A1(n19138), .A2(n18072), .ZN(n14836) );
NAND2_X2 U10341 ( .A1(n17897), .A2(n14839), .ZN(n14829) );
NAND2_X2 U10342 ( .A1(n18042), .A2(b_in[84]), .ZN(n14818) );
NAND2_X2 U10343 ( .A1(n14840), .A2(n14841), .ZN(N3170) );
NAND2_X2 U10344 ( .A1(n14842), .A2(n18065), .ZN(n14841) );
XNOR2_X2 U10345 ( .A(n18994), .B(n14843), .ZN(n14842) );
NAND2_X2 U10347 ( .A1(n17920), .A2(n14847), .ZN(n13872) );
XNOR2_X2 U10348 ( .A(n19056), .B(aes_text_out[99]), .ZN(n14847) );
XNOR2_X2 U10350 ( .A(n14848), .B(aes_text_out[99]), .ZN(n13874) );
NAND2_X2 U10352 ( .A1(n14849), .A2(n14850), .ZN(n14844) );
NAND2_X2 U10353 ( .A1(n17996), .A2(aad_byte_cnt[32]), .ZN(n14850) );
NAND2_X2 U10354 ( .A1(n17913), .A2(n14848), .ZN(n14849) );
NAND4_X2 U10355 ( .A1(n14851), .A2(n14852), .A3(n14853), .A4(n14854), .ZN(n14848) );
NAND2_X2 U10356 ( .A1(n19092), .A2(n17888), .ZN(n14854) );
NAND2_X2 U10360 ( .A1(n19071), .A2(n17894), .ZN(n14852) );
NAND4_X2 U10361 ( .A1(n14858), .A2(n14859), .A3(n14860), .A4(n17881), .ZN(n14506) );
NAND2_X2 U10362 ( .A1(n17883), .A2(n19072), .ZN(n14860) );
NAND2_X2 U10363 ( .A1(n19171), .A2(n18076), .ZN(n14859) );
NAND2_X2 U10364 ( .A1(n19139), .A2(n18072), .ZN(n14858) );
NAND2_X2 U10365 ( .A1(n17897), .A2(n14861), .ZN(n14851) );
NAND2_X2 U10366 ( .A1(n18042), .A2(b_in[83]), .ZN(n14840) );
NAND2_X2 U10367 ( .A1(n14862), .A2(n14863), .ZN(N3169) );
NAND2_X2 U10368 ( .A1(n14864), .A2(n18065), .ZN(n14863) );
XNOR2_X2 U10369 ( .A(n18993), .B(n14865), .ZN(n14864) );
NAND2_X2 U10371 ( .A1(n17920), .A2(n14869), .ZN(n13866) );
XNOR2_X2 U10372 ( .A(n19058), .B(aes_text_out[98]), .ZN(n14869) );
XNOR2_X2 U10374 ( .A(n14870), .B(aes_text_out[98]), .ZN(n13868) );
NAND2_X2 U10376 ( .A1(n14871), .A2(n14872), .ZN(n14866) );
NAND2_X2 U10377 ( .A1(n17996), .A2(aad_byte_cnt[31]), .ZN(n14872) );
NAND2_X2 U10378 ( .A1(n17913), .A2(n14870), .ZN(n14871) );
NAND4_X2 U10379 ( .A1(n14873), .A2(n14874), .A3(n14875), .A4(n14876), .ZN(n14870) );
NAND2_X2 U10380 ( .A1(n19095), .A2(n17888), .ZN(n14876) );
NAND2_X2 U10384 ( .A1(n19073), .A2(n17894), .ZN(n14874) );
NAND4_X2 U10385 ( .A1(n14880), .A2(n14881), .A3(n14882), .A4(n17881), .ZN(n14528) );
NAND2_X2 U10386 ( .A1(n17883), .A2(n19074), .ZN(n14882) );
NAND2_X2 U10387 ( .A1(n19172), .A2(n18076), .ZN(n14881) );
NAND2_X2 U10388 ( .A1(n19140), .A2(n18072), .ZN(n14880) );
NAND2_X2 U10389 ( .A1(n17897), .A2(n14883), .ZN(n14873) );
NAND2_X2 U10390 ( .A1(n18042), .A2(b_in[82]), .ZN(n14862) );
NAND2_X2 U10391 ( .A1(n14884), .A2(n14885), .ZN(N3168) );
NAND2_X2 U10392 ( .A1(n14886), .A2(n18065), .ZN(n14885) );
XNOR2_X2 U10393 ( .A(n18992), .B(n14887), .ZN(n14886) );
NAND2_X2 U10395 ( .A1(n17921), .A2(n14891), .ZN(n13860) );
XNOR2_X2 U10396 ( .A(n19060), .B(aes_text_out[97]), .ZN(n14891) );
XNOR2_X2 U10398 ( .A(n14892), .B(aes_text_out[97]), .ZN(n13862) );
NAND2_X2 U10400 ( .A1(n14893), .A2(n14894), .ZN(n14888) );
NAND2_X2 U10401 ( .A1(n17997), .A2(aad_byte_cnt[30]), .ZN(n14894) );
NAND2_X2 U10402 ( .A1(n17913), .A2(n14892), .ZN(n14893) );
NAND4_X2 U10403 ( .A1(n14895), .A2(n14896), .A3(n14897), .A4(n14898), .ZN(n14892) );
NAND2_X2 U10404 ( .A1(n19098), .A2(n17888), .ZN(n14898) );
NAND2_X2 U10408 ( .A1(n19075), .A2(n17894), .ZN(n14896) );
NAND4_X2 U10409 ( .A1(n14902), .A2(n14903), .A3(n14904), .A4(n17881), .ZN(n14550) );
NAND2_X2 U10410 ( .A1(n17882), .A2(n19076), .ZN(n14904) );
NAND2_X2 U10411 ( .A1(n19173), .A2(n18076), .ZN(n14903) );
NAND2_X2 U10412 ( .A1(n19141), .A2(n18072), .ZN(n14902) );
NAND2_X2 U10413 ( .A1(n17897), .A2(n14905), .ZN(n14895) );
NAND2_X2 U10414 ( .A1(n18042), .A2(b_in[81]), .ZN(n14884) );
NAND2_X2 U10415 ( .A1(n14906), .A2(n14907), .ZN(N3167) );
NAND2_X2 U10416 ( .A1(n14908), .A2(n18065), .ZN(n14907) );
XNOR2_X2 U10417 ( .A(n18991), .B(n14909), .ZN(n14908) );
NAND2_X2 U10419 ( .A1(n17921), .A2(n14913), .ZN(n13854) );
XNOR2_X2 U10420 ( .A(n19062), .B(aes_text_out[96]), .ZN(n14913) );
NAND2_X2 U10422 ( .A1(n17934), .A2(n14736), .ZN(n14758) );
NAND2_X2 U10424 ( .A1(dii_data_size[1]), .A2(dii_data_size[0]), .ZN(n14914));
XNOR2_X2 U10425 ( .A(n14915), .B(aes_text_out[96]), .ZN(n13856) );
NAND2_X2 U10427 ( .A1(n14916), .A2(n14917), .ZN(n14910) );
NAND2_X2 U10428 ( .A1(n17997), .A2(aad_byte_cnt[29]), .ZN(n14917) );
NAND2_X2 U10429 ( .A1(n17913), .A2(n14915), .ZN(n14916) );
NAND4_X2 U10430 ( .A1(n14918), .A2(n14919), .A3(n14920), .A4(n14921), .ZN(n14915) );
NAND2_X2 U10431 ( .A1(n19101), .A2(n17888), .ZN(n14921) );
NAND2_X2 U10435 ( .A1(n19077), .A2(n17894), .ZN(n14919) );
NAND4_X2 U10436 ( .A1(n14925), .A2(n14926), .A3(n14927), .A4(n17881), .ZN(n14574) );
NAND2_X2 U10437 ( .A1(n17882), .A2(n19078), .ZN(n14927) );
NAND2_X2 U10438 ( .A1(n19174), .A2(n18076), .ZN(n14926) );
NAND2_X2 U10439 ( .A1(n19142), .A2(n18072), .ZN(n14925) );
NAND2_X2 U10440 ( .A1(n17897), .A2(n14928), .ZN(n14918) );
NAND2_X2 U10441 ( .A1(n18042), .A2(b_in[80]), .ZN(n14906) );
NAND2_X2 U10442 ( .A1(n14929), .A2(n14930), .ZN(N3166) );
NAND2_X2 U10443 ( .A1(n14931), .A2(n18065), .ZN(n14930) );
XNOR2_X2 U10444 ( .A(n18990), .B(n14932), .ZN(n14931) );
NAND2_X2 U10446 ( .A1(n17921), .A2(n14936), .ZN(n13848) );
XNOR2_X2 U10447 ( .A(n19064), .B(aes_text_out[95]), .ZN(n14936) );
XNOR2_X2 U10449 ( .A(n14938), .B(aes_text_out[95]), .ZN(n13850) );
NAND2_X2 U10451 ( .A1(n14939), .A2(n14940), .ZN(n14933) );
NAND2_X2 U10452 ( .A1(n17997), .A2(aad_byte_cnt[28]), .ZN(n14940) );
NAND2_X2 U10453 ( .A1(n17913), .A2(n14938), .ZN(n14939) );
NAND4_X2 U10454 ( .A1(n14941), .A2(n14942), .A3(n14943), .A4(n14944), .ZN(n14938) );
NAND2_X2 U10455 ( .A1(n14945), .A2(n14564), .ZN(n14944) );
NAND2_X2 U10459 ( .A1(n19104), .A2(n17888), .ZN(n14942) );
NAND2_X2 U10460 ( .A1(n19080), .A2(n17894), .ZN(n14941) );
NAND2_X2 U10462 ( .A1(n19143), .A2(n18072), .ZN(n14950) );
NAND2_X2 U10463 ( .A1(dii_data_size[2]), .A2(n14185), .ZN(n14949) );
NAND2_X2 U10464 ( .A1(n14951), .A2(n14952), .ZN(n14185) );
NAND2_X2 U10465 ( .A1(n19175), .A2(n18076), .ZN(n14952) );
NAND2_X2 U10466 ( .A1(n18074), .A2(n19081), .ZN(n14951) );
NAND2_X2 U10467 ( .A1(n18042), .A2(b_in[79]), .ZN(n14929) );
NAND2_X2 U10468 ( .A1(n14953), .A2(n14954), .ZN(N3165) );
NAND2_X2 U10469 ( .A1(n14955), .A2(n18065), .ZN(n14954) );
XNOR2_X2 U10470 ( .A(n18989), .B(n14956), .ZN(n14955) );
NAND2_X2 U10472 ( .A1(n17921), .A2(n14960), .ZN(n13842) );
XNOR2_X2 U10473 ( .A(n19066), .B(aes_text_out[94]), .ZN(n14960) );
XNOR2_X2 U10475 ( .A(n14961), .B(aes_text_out[94]), .ZN(n13844) );
NAND2_X2 U10477 ( .A1(n14962), .A2(n14963), .ZN(n14957) );
NAND2_X2 U10478 ( .A1(n17997), .A2(aad_byte_cnt[27]), .ZN(n14963) );
NAND2_X2 U10479 ( .A1(n17913), .A2(n14961), .ZN(n14962) );
NAND4_X2 U10480 ( .A1(n14964), .A2(n14965), .A3(n14966), .A4(n14967), .ZN(n14961) );
NAND2_X2 U10481 ( .A1(n14968), .A2(n14564), .ZN(n14967) );
NAND2_X2 U10485 ( .A1(n19107), .A2(n17888), .ZN(n14965) );
NAND2_X2 U10486 ( .A1(n19083), .A2(n17894), .ZN(n14964) );
NAND2_X2 U10488 ( .A1(n19144), .A2(n18072), .ZN(n14972) );
NAND2_X2 U10489 ( .A1(dii_data_size[2]), .A2(n14216), .ZN(n14971) );
NAND2_X2 U10490 ( .A1(n14973), .A2(n14974), .ZN(n14216) );
NAND2_X2 U10491 ( .A1(n19176), .A2(n18076), .ZN(n14974) );
NAND2_X2 U10492 ( .A1(n18074), .A2(n19084), .ZN(n14973) );
NAND2_X2 U10493 ( .A1(n18042), .A2(b_in[78]), .ZN(n14953) );
NAND2_X2 U10494 ( .A1(n14975), .A2(n14976), .ZN(N3164) );
NAND2_X2 U10495 ( .A1(n14977), .A2(n18065), .ZN(n14976) );
XNOR2_X2 U10496 ( .A(n18988), .B(n14978), .ZN(n14977) );
NAND2_X2 U10498 ( .A1(n17921), .A2(n14982), .ZN(n13836) );
XNOR2_X2 U10499 ( .A(n19068), .B(aes_text_out[93]), .ZN(n14982) );
XNOR2_X2 U10501 ( .A(n14983), .B(aes_text_out[93]), .ZN(n13838) );
NAND2_X2 U10503 ( .A1(n14984), .A2(n14985), .ZN(n14979) );
NAND2_X2 U10504 ( .A1(n17997), .A2(aad_byte_cnt[26]), .ZN(n14985) );
NAND2_X2 U10505 ( .A1(n17913), .A2(n14983), .ZN(n14984) );
NAND4_X2 U10506 ( .A1(n14986), .A2(n14987), .A3(n14988), .A4(n14989), .ZN(n14983) );
NAND2_X2 U10507 ( .A1(n14990), .A2(n14564), .ZN(n14989) );
NAND2_X2 U10511 ( .A1(n19110), .A2(n17888), .ZN(n14987) );
NAND2_X2 U10512 ( .A1(n19086), .A2(n17894), .ZN(n14986) );
NAND2_X2 U10514 ( .A1(n19145), .A2(n18072), .ZN(n14994) );
NAND2_X2 U10515 ( .A1(dii_data_size[2]), .A2(n14245), .ZN(n14993) );
NAND2_X2 U10516 ( .A1(n14995), .A2(n14996), .ZN(n14245) );
NAND2_X2 U10517 ( .A1(n19177), .A2(n18076), .ZN(n14996) );
NAND2_X2 U10518 ( .A1(n18074), .A2(n19087), .ZN(n14995) );
NAND2_X2 U10519 ( .A1(n18041), .A2(b_in[77]), .ZN(n14975) );
NAND2_X2 U10520 ( .A1(n14997), .A2(n14998), .ZN(N3163) );
NAND2_X2 U10521 ( .A1(n14999), .A2(n18065), .ZN(n14998) );
XNOR2_X2 U10522 ( .A(n18987), .B(n15000), .ZN(n14999) );
NAND2_X2 U10524 ( .A1(n17921), .A2(n15004), .ZN(n13830) );
XNOR2_X2 U10525 ( .A(n19070), .B(aes_text_out[92]), .ZN(n15004) );
XNOR2_X2 U10527 ( .A(n15005), .B(aes_text_out[92]), .ZN(n13832) );
NAND2_X2 U10529 ( .A1(n15006), .A2(n15007), .ZN(n15001) );
NAND2_X2 U10530 ( .A1(n17997), .A2(aad_byte_cnt[25]), .ZN(n15007) );
NAND2_X2 U10531 ( .A1(n17913), .A2(n15005), .ZN(n15006) );
NAND4_X2 U10532 ( .A1(n15008), .A2(n15009), .A3(n15010), .A4(n15011), .ZN(n15005) );
NAND2_X2 U10533 ( .A1(n15012), .A2(n14564), .ZN(n15011) );
NAND2_X2 U10537 ( .A1(n19113), .A2(n17888), .ZN(n15009) );
NAND2_X2 U10538 ( .A1(n19089), .A2(n17894), .ZN(n15008) );
NAND2_X2 U10540 ( .A1(n19146), .A2(n18072), .ZN(n15016) );
NAND2_X2 U10541 ( .A1(dii_data_size[2]), .A2(n14274), .ZN(n15015) );
NAND2_X2 U10542 ( .A1(n15017), .A2(n15018), .ZN(n14274) );
NAND2_X2 U10543 ( .A1(n19178), .A2(n18076), .ZN(n15018) );
NAND2_X2 U10544 ( .A1(n18074), .A2(n19090), .ZN(n15017) );
NAND2_X2 U10545 ( .A1(n18041), .A2(b_in[76]), .ZN(n14997) );
NAND2_X2 U10546 ( .A1(n15019), .A2(n15020), .ZN(N3162) );
NAND2_X2 U10547 ( .A1(n15021), .A2(n18065), .ZN(n15020) );
XNOR2_X2 U10548 ( .A(n18986), .B(n15022), .ZN(n15021) );
NAND2_X2 U10550 ( .A1(n17921), .A2(n15026), .ZN(n13824) );
XNOR2_X2 U10551 ( .A(n19072), .B(aes_text_out[91]), .ZN(n15026) );
XNOR2_X2 U10553 ( .A(n15027), .B(aes_text_out[91]), .ZN(n13826) );
NAND2_X2 U10555 ( .A1(n15028), .A2(n15029), .ZN(n15023) );
NAND2_X2 U10556 ( .A1(n17997), .A2(aad_byte_cnt[24]), .ZN(n15029) );
NAND2_X2 U10557 ( .A1(n17913), .A2(n15027), .ZN(n15028) );
NAND4_X2 U10558 ( .A1(n15030), .A2(n15031), .A3(n15032), .A4(n15033), .ZN(n15027) );
NAND2_X2 U10559 ( .A1(n15034), .A2(n14564), .ZN(n15033) );
NAND2_X2 U10563 ( .A1(n19116), .A2(n17888), .ZN(n15031) );
NAND2_X2 U10564 ( .A1(n19092), .A2(n17894), .ZN(n15030) );
NAND2_X2 U10566 ( .A1(n19147), .A2(n18072), .ZN(n15038) );
NAND2_X2 U10567 ( .A1(dii_data_size[2]), .A2(n14303), .ZN(n15037) );
NAND2_X2 U10568 ( .A1(n15039), .A2(n15040), .ZN(n14303) );
NAND2_X2 U10569 ( .A1(n19179), .A2(n18076), .ZN(n15040) );
NAND2_X2 U10570 ( .A1(n18074), .A2(n19093), .ZN(n15039) );
NAND2_X2 U10571 ( .A1(n18041), .A2(b_in[75]), .ZN(n15019) );
NAND2_X2 U10572 ( .A1(n15041), .A2(n15042), .ZN(N3161) );
NAND2_X2 U10573 ( .A1(n15043), .A2(n18066), .ZN(n15042) );
XNOR2_X2 U10574 ( .A(n18985), .B(n15044), .ZN(n15043) );
NAND2_X2 U10576 ( .A1(n17921), .A2(n15048), .ZN(n13818) );
XNOR2_X2 U10577 ( .A(n19074), .B(aes_text_out[90]), .ZN(n15048) );
XNOR2_X2 U10579 ( .A(n15049), .B(aes_text_out[90]), .ZN(n13820) );
NAND2_X2 U10581 ( .A1(n15050), .A2(n15051), .ZN(n15045) );
NAND2_X2 U10582 ( .A1(n17997), .A2(aad_byte_cnt[23]), .ZN(n15051) );
NAND2_X2 U10583 ( .A1(n17912), .A2(n15049), .ZN(n15050) );
NAND4_X2 U10584 ( .A1(n15052), .A2(n15053), .A3(n15054), .A4(n15055), .ZN(n15049) );
NAND2_X2 U10585 ( .A1(n15056), .A2(n14564), .ZN(n15055) );
NAND2_X2 U10589 ( .A1(n19119), .A2(n17888), .ZN(n15053) );
NAND2_X2 U10590 ( .A1(n19095), .A2(n17893), .ZN(n15052) );
NAND2_X2 U10592 ( .A1(n19148), .A2(n18072), .ZN(n15060) );
NAND2_X2 U10593 ( .A1(dii_data_size[2]), .A2(n14332), .ZN(n15059) );
NAND2_X2 U10594 ( .A1(n15061), .A2(n15062), .ZN(n14332) );
NAND2_X2 U10595 ( .A1(n19180), .A2(n18076), .ZN(n15062) );
NAND2_X2 U10596 ( .A1(n18074), .A2(n19096), .ZN(n15061) );
NAND2_X2 U10597 ( .A1(n18041), .A2(b_in[74]), .ZN(n15041) );
NAND2_X2 U10598 ( .A1(n15063), .A2(n15064), .ZN(N3160) );
NAND2_X2 U10599 ( .A1(n15065), .A2(n18066), .ZN(n15064) );
XNOR2_X2 U10600 ( .A(n18984), .B(n15066), .ZN(n15065) );
NAND2_X2 U10602 ( .A1(n17921), .A2(n15070), .ZN(n13812) );
XNOR2_X2 U10603 ( .A(n19076), .B(aes_text_out[89]), .ZN(n15070) );
XNOR2_X2 U10605 ( .A(n15071), .B(aes_text_out[89]), .ZN(n13814) );
NAND2_X2 U10607 ( .A1(n15072), .A2(n15073), .ZN(n15067) );
NAND2_X2 U10608 ( .A1(n17997), .A2(aad_byte_cnt[22]), .ZN(n15073) );
NAND2_X2 U10609 ( .A1(n17912), .A2(n15071), .ZN(n15072) );
NAND4_X2 U10610 ( .A1(n15074), .A2(n15075), .A3(n15076), .A4(n15077), .ZN(n15071) );
NAND2_X2 U10611 ( .A1(n15078), .A2(n14564), .ZN(n15077) );
NAND2_X2 U10615 ( .A1(n19122), .A2(n17887), .ZN(n15075) );
NAND2_X2 U10616 ( .A1(n19098), .A2(n17893), .ZN(n15074) );
NAND2_X2 U10618 ( .A1(n19149), .A2(n18072), .ZN(n15082) );
NAND2_X2 U10619 ( .A1(dii_data_size[2]), .A2(n14361), .ZN(n15081) );
NAND2_X2 U10620 ( .A1(n15083), .A2(n15084), .ZN(n14361) );
NAND2_X2 U10621 ( .A1(n19181), .A2(n18076), .ZN(n15084) );
NAND2_X2 U10622 ( .A1(n18074), .A2(n19099), .ZN(n15083) );
NAND2_X2 U10623 ( .A1(n18041), .A2(b_in[73]), .ZN(n15063) );
NAND2_X2 U10624 ( .A1(n15085), .A2(n15086), .ZN(N3159) );
NAND2_X2 U10625 ( .A1(n15087), .A2(n18066), .ZN(n15086) );
XNOR2_X2 U10626 ( .A(n18983), .B(n15088), .ZN(n15087) );
NAND2_X2 U10628 ( .A1(n17921), .A2(n15092), .ZN(n13806) );
XNOR2_X2 U10629 ( .A(n19078), .B(aes_text_out[88]), .ZN(n15092) );
NAND2_X2 U10631 ( .A1(n17934), .A2(n15093), .ZN(n14937) );
NAND2_X2 U10632 ( .A1(n19201), .A2(n18072), .ZN(n15093) );
XNOR2_X2 U10633 ( .A(n15095), .B(aes_text_out[88]), .ZN(n13808) );
NAND2_X2 U10635 ( .A1(n15096), .A2(n15097), .ZN(n15089) );
NAND2_X2 U10636 ( .A1(n17997), .A2(aad_byte_cnt[21]), .ZN(n15097) );
NAND2_X2 U10637 ( .A1(n17912), .A2(n15095), .ZN(n15096) );
NAND4_X2 U10638 ( .A1(n15098), .A2(n15099), .A3(n15100), .A4(n15101), .ZN(n15095) );
NAND2_X2 U10639 ( .A1(n15102), .A2(n14564), .ZN(n15101) );
NAND2_X2 U10643 ( .A1(n19125), .A2(n17887), .ZN(n15099) );
NAND2_X2 U10644 ( .A1(n19101), .A2(n17893), .ZN(n15098) );
NAND2_X2 U10646 ( .A1(n19150), .A2(n18072), .ZN(n15106) );
NAND2_X2 U10647 ( .A1(dii_data_size[2]), .A2(n14391), .ZN(n15105) );
NAND2_X2 U10648 ( .A1(n15107), .A2(n15108), .ZN(n14391) );
NAND2_X2 U10649 ( .A1(n19182), .A2(n18076), .ZN(n15108) );
NAND2_X2 U10650 ( .A1(n18074), .A2(n19102), .ZN(n15107) );
NAND2_X2 U10651 ( .A1(n18041), .A2(b_in[72]), .ZN(n15085) );
NAND2_X2 U10652 ( .A1(n15109), .A2(n15110), .ZN(N3158) );
NAND2_X2 U10653 ( .A1(n15111), .A2(n18066), .ZN(n15110) );
XNOR2_X2 U10654 ( .A(n18982), .B(n15112), .ZN(n15111) );
NAND2_X2 U10656 ( .A1(n17921), .A2(n15116), .ZN(n13800) );
XNOR2_X2 U10657 ( .A(n19081), .B(aes_text_out[87]), .ZN(n15116) );
XNOR2_X2 U10659 ( .A(n15118), .B(aes_text_out[87]), .ZN(n13802) );
NAND2_X2 U10661 ( .A1(n15119), .A2(n15120), .ZN(n15113) );
NAND2_X2 U10662 ( .A1(n17997), .A2(aad_byte_cnt[20]), .ZN(n15120) );
NAND2_X2 U10663 ( .A1(n17912), .A2(n15118), .ZN(n15119) );
NAND2_X2 U10669 ( .A1(n14945), .A2(n17887), .ZN(n15122) );
NAND2_X2 U10670 ( .A1(n19104), .A2(n17893), .ZN(n15121) );
NAND2_X2 U10672 ( .A1(n19151), .A2(n18072), .ZN(n15129) );
NAND2_X2 U10673 ( .A1(dii_data_size[2]), .A2(n14421), .ZN(n15128) );
NAND2_X2 U10674 ( .A1(n15130), .A2(n15131), .ZN(n14421) );
NAND2_X2 U10675 ( .A1(n19183), .A2(n18076), .ZN(n15131) );
NAND2_X2 U10676 ( .A1(n18074), .A2(n19105), .ZN(n15130) );
NAND2_X2 U10677 ( .A1(n18041), .A2(b_in[71]), .ZN(n15109) );
NAND2_X2 U10678 ( .A1(n15132), .A2(n15133), .ZN(N3157) );
NAND2_X2 U10679 ( .A1(n15134), .A2(n18066), .ZN(n15133) );
XNOR2_X2 U10680 ( .A(n18981), .B(n15135), .ZN(n15134) );
NAND2_X2 U10682 ( .A1(n17922), .A2(n15139), .ZN(n13794) );
XNOR2_X2 U10683 ( .A(n19084), .B(aes_text_out[86]), .ZN(n15139) );
XNOR2_X2 U10685 ( .A(n15140), .B(aes_text_out[86]), .ZN(n13796) );
NAND2_X2 U10687 ( .A1(n15141), .A2(n15142), .ZN(n15136) );
NAND2_X2 U10688 ( .A1(n17997), .A2(aad_byte_cnt[19]), .ZN(n15142) );
NAND2_X2 U10689 ( .A1(n17912), .A2(n15140), .ZN(n15141) );
NAND2_X2 U10695 ( .A1(n14968), .A2(n17887), .ZN(n15144) );
NAND2_X2 U10696 ( .A1(n19107), .A2(n17893), .ZN(n15143) );
NAND2_X2 U10698 ( .A1(n19152), .A2(n18072), .ZN(n15151) );
NAND2_X2 U10699 ( .A1(dii_data_size[2]), .A2(n14444), .ZN(n15150) );
NAND2_X2 U10700 ( .A1(n15152), .A2(n15153), .ZN(n14444) );
NAND2_X2 U10701 ( .A1(n19184), .A2(n18076), .ZN(n15153) );
NAND2_X2 U10702 ( .A1(n18074), .A2(n19108), .ZN(n15152) );
NAND2_X2 U10703 ( .A1(n18041), .A2(b_in[70]), .ZN(n15132) );
NAND2_X2 U10704 ( .A1(n15154), .A2(n15155), .ZN(N3156) );
NAND2_X2 U10705 ( .A1(n15156), .A2(n18066), .ZN(n15155) );
XNOR2_X2 U10706 ( .A(n18980), .B(n15157), .ZN(n15156) );
NAND2_X2 U10708 ( .A1(n17922), .A2(n15161), .ZN(n13788) );
XNOR2_X2 U10709 ( .A(n19087), .B(aes_text_out[85]), .ZN(n15161) );
XNOR2_X2 U10711 ( .A(n15162), .B(aes_text_out[85]), .ZN(n13790) );
NAND2_X2 U10713 ( .A1(n15163), .A2(n15164), .ZN(n15158) );
NAND2_X2 U10714 ( .A1(n17997), .A2(aad_byte_cnt[18]), .ZN(n15164) );
NAND2_X2 U10715 ( .A1(n17912), .A2(n15162), .ZN(n15163) );
NAND2_X2 U10721 ( .A1(n14990), .A2(n17887), .ZN(n15166) );
NAND2_X2 U10722 ( .A1(n19110), .A2(n17893), .ZN(n15165) );
NAND2_X2 U10724 ( .A1(n19153), .A2(n18072), .ZN(n15173) );
NAND2_X2 U10725 ( .A1(dii_data_size[2]), .A2(n14466), .ZN(n15172) );
NAND2_X2 U10726 ( .A1(n15174), .A2(n15175), .ZN(n14466) );
NAND2_X2 U10727 ( .A1(n19185), .A2(n18076), .ZN(n15175) );
NAND2_X2 U10728 ( .A1(n18074), .A2(n19111), .ZN(n15174) );
NAND2_X2 U10729 ( .A1(n18041), .A2(b_in[69]), .ZN(n15154) );
NAND2_X2 U10730 ( .A1(n15176), .A2(n15177), .ZN(N3155) );
NAND2_X2 U10731 ( .A1(n15178), .A2(n18066), .ZN(n15177) );
XNOR2_X2 U10732 ( .A(n18979), .B(n15179), .ZN(n15178) );
NAND2_X2 U10734 ( .A1(n17922), .A2(n15183), .ZN(n13782) );
XNOR2_X2 U10735 ( .A(n19090), .B(aes_text_out[84]), .ZN(n15183) );
XNOR2_X2 U10737 ( .A(n15184), .B(aes_text_out[84]), .ZN(n13784) );
NAND2_X2 U10739 ( .A1(n15185), .A2(n15186), .ZN(n15180) );
NAND2_X2 U10740 ( .A1(n17997), .A2(aad_byte_cnt[17]), .ZN(n15186) );
NAND2_X2 U10741 ( .A1(n17912), .A2(n15184), .ZN(n15185) );
NAND2_X2 U10747 ( .A1(n15012), .A2(n17887), .ZN(n15188) );
NAND2_X2 U10748 ( .A1(n19113), .A2(n17893), .ZN(n15187) );
NAND2_X2 U10750 ( .A1(n19154), .A2(n18072), .ZN(n15195) );
NAND2_X2 U10751 ( .A1(dii_data_size[2]), .A2(n14488), .ZN(n15194) );
NAND2_X2 U10752 ( .A1(n15196), .A2(n15197), .ZN(n14488) );
NAND2_X2 U10753 ( .A1(n19186), .A2(n18076), .ZN(n15197) );
NAND2_X2 U10754 ( .A1(n18074), .A2(n19114), .ZN(n15196) );
NAND2_X2 U10755 ( .A1(n18041), .A2(b_in[68]), .ZN(n15176) );
NAND2_X2 U10756 ( .A1(n15198), .A2(n15199), .ZN(N3154) );
NAND2_X2 U10757 ( .A1(n15200), .A2(n18066), .ZN(n15199) );
XNOR2_X2 U10758 ( .A(n18978), .B(n15201), .ZN(n15200) );
NAND2_X2 U10760 ( .A1(n17922), .A2(n15205), .ZN(n13776) );
XNOR2_X2 U10761 ( .A(n19093), .B(aes_text_out[83]), .ZN(n15205) );
XNOR2_X2 U10763 ( .A(n15206), .B(aes_text_out[83]), .ZN(n13778) );
NAND2_X2 U10765 ( .A1(n15207), .A2(n15208), .ZN(n15202) );
NAND2_X2 U10766 ( .A1(n17997), .A2(aad_byte_cnt[16]), .ZN(n15208) );
NAND2_X2 U10767 ( .A1(n17912), .A2(n15206), .ZN(n15207) );
NAND2_X2 U10773 ( .A1(n15034), .A2(n17887), .ZN(n15210) );
NAND2_X2 U10774 ( .A1(n19116), .A2(n17893), .ZN(n15209) );
NAND2_X2 U10776 ( .A1(n19155), .A2(n18072), .ZN(n15217) );
NAND2_X2 U10777 ( .A1(dii_data_size[2]), .A2(n14510), .ZN(n15216) );
NAND2_X2 U10778 ( .A1(n15218), .A2(n15219), .ZN(n14510) );
NAND2_X2 U10779 ( .A1(n19187), .A2(n18076), .ZN(n15219) );
NAND2_X2 U10780 ( .A1(n18074), .A2(n19117), .ZN(n15218) );
NAND2_X2 U10781 ( .A1(n18041), .A2(b_in[67]), .ZN(n15198) );
NAND2_X2 U10782 ( .A1(n15220), .A2(n15221), .ZN(N3153) );
NAND2_X2 U10783 ( .A1(n15222), .A2(n18066), .ZN(n15221) );
XNOR2_X2 U10784 ( .A(n18977), .B(n15223), .ZN(n15222) );
NAND2_X2 U10786 ( .A1(n17922), .A2(n15227), .ZN(n13770) );
XNOR2_X2 U10787 ( .A(n19096), .B(aes_text_out[82]), .ZN(n15227) );
XNOR2_X2 U10789 ( .A(n15228), .B(aes_text_out[82]), .ZN(n13772) );
NAND2_X2 U10791 ( .A1(n15229), .A2(n15230), .ZN(n15224) );
NAND2_X2 U10792 ( .A1(n17997), .A2(aad_byte_cnt[15]), .ZN(n15230) );
NAND2_X2 U10793 ( .A1(n17912), .A2(n15228), .ZN(n15229) );
NAND2_X2 U10799 ( .A1(n15056), .A2(n17887), .ZN(n15232) );
NAND2_X2 U10800 ( .A1(n19119), .A2(n17893), .ZN(n15231) );
NAND2_X2 U10802 ( .A1(n19156), .A2(n18072), .ZN(n15239) );
NAND2_X2 U10803 ( .A1(dii_data_size[2]), .A2(n14532), .ZN(n15238) );
NAND2_X2 U10804 ( .A1(n15240), .A2(n15241), .ZN(n14532) );
NAND2_X2 U10805 ( .A1(n19188), .A2(n18076), .ZN(n15241) );
NAND2_X2 U10806 ( .A1(n18074), .A2(n19120), .ZN(n15240) );
NAND2_X2 U10807 ( .A1(n18041), .A2(b_in[66]), .ZN(n15220) );
NAND2_X2 U10808 ( .A1(n15242), .A2(n15243), .ZN(N3152) );
NAND2_X2 U10809 ( .A1(n15244), .A2(n18066), .ZN(n15243) );
XNOR2_X2 U10810 ( .A(n18976), .B(n15245), .ZN(n15244) );
NAND2_X2 U10812 ( .A1(n17922), .A2(n15249), .ZN(n13764) );
XNOR2_X2 U10813 ( .A(n19099), .B(aes_text_out[81]), .ZN(n15249) );
XNOR2_X2 U10815 ( .A(n15250), .B(aes_text_out[81]), .ZN(n13766) );
NAND2_X2 U10817 ( .A1(n15251), .A2(n15252), .ZN(n15246) );
NAND2_X2 U10818 ( .A1(n17997), .A2(aad_byte_cnt[14]), .ZN(n15252) );
NAND2_X2 U10819 ( .A1(n17912), .A2(n15250), .ZN(n15251) );
NAND2_X2 U10825 ( .A1(n15078), .A2(n17887), .ZN(n15254) );
NAND2_X2 U10826 ( .A1(n19122), .A2(n17894), .ZN(n15253) );
NAND2_X2 U10828 ( .A1(n19157), .A2(n18072), .ZN(n15261) );
NAND2_X2 U10829 ( .A1(dii_data_size[2]), .A2(n14554), .ZN(n15260) );
NAND2_X2 U10830 ( .A1(n15262), .A2(n15263), .ZN(n14554) );
NAND2_X2 U10831 ( .A1(n18074), .A2(n19123), .ZN(n15263) );
NAND2_X2 U10832 ( .A1(n19189), .A2(n18076), .ZN(n15262) );
NAND2_X2 U10833 ( .A1(n18041), .A2(b_in[65]), .ZN(n15242) );
NAND2_X2 U10834 ( .A1(n15264), .A2(n15265), .ZN(N3151) );
NAND2_X2 U10835 ( .A1(n15266), .A2(n18066), .ZN(n15265) );
XNOR2_X2 U10836 ( .A(n18975), .B(n15267), .ZN(n15266) );
NAND2_X2 U10838 ( .A1(n17922), .A2(n15271), .ZN(n13758) );
XNOR2_X2 U10839 ( .A(n19102), .B(aes_text_out[80]), .ZN(n15271) );
NAND2_X2 U10841 ( .A1(n17934), .A2(n15094), .ZN(n15117) );
NAND2_X2 U10842 ( .A1(n15272), .A2(n15273), .ZN(n15094) );
NAND2_X2 U10843 ( .A1(dii_data_size[2]), .A2(n17865), .ZN(n15273) );
XNOR2_X2 U10844 ( .A(n15274), .B(aes_text_out[80]), .ZN(n13760) );
NAND2_X2 U10846 ( .A1(n15275), .A2(n15276), .ZN(n15268) );
NAND2_X2 U10847 ( .A1(n17997), .A2(aad_byte_cnt[13]), .ZN(n15276) );
NAND2_X2 U10848 ( .A1(n17912), .A2(n15274), .ZN(n15275) );
NAND2_X2 U10854 ( .A1(n15102), .A2(n17887), .ZN(n15278) );
NAND2_X2 U10855 ( .A1(n19125), .A2(n17893), .ZN(n15277) );
NAND2_X2 U10857 ( .A1(n19158), .A2(n18073), .ZN(n15285) );
NAND2_X2 U10858 ( .A1(dii_data_size[2]), .A2(n14578), .ZN(n15284) );
NAND2_X2 U10859 ( .A1(n15286), .A2(n15287), .ZN(n14578) );
NAND2_X2 U10860 ( .A1(n18074), .A2(n19126), .ZN(n15287) );
NAND2_X2 U10861 ( .A1(n19190), .A2(n18075), .ZN(n15286) );
NAND2_X2 U10862 ( .A1(n18041), .A2(b_in[64]), .ZN(n15264) );
NAND2_X2 U10863 ( .A1(n15288), .A2(n15289), .ZN(N3150) );
NAND2_X2 U10864 ( .A1(n15290), .A2(n18066), .ZN(n15289) );
XNOR2_X2 U10865 ( .A(n18974), .B(n15291), .ZN(n15290) );
NAND2_X2 U10867 ( .A1(n17922), .A2(n15295), .ZN(n13752) );
XNOR2_X2 U10868 ( .A(n19105), .B(aes_text_out[79]), .ZN(n15295) );
XNOR2_X2 U10870 ( .A(n15297), .B(aes_text_out[79]), .ZN(n13754) );
NAND2_X2 U10872 ( .A1(n15298), .A2(n15299), .ZN(n15292) );
NAND2_X2 U10873 ( .A1(n17997), .A2(aad_byte_cnt[12]), .ZN(n15299) );
NAND2_X2 U10874 ( .A1(n17911), .A2(n15297), .ZN(n15298) );
NAND4_X2 U10875 ( .A1(n15300), .A2(n15301), .A3(n15302), .A4(n15303), .ZN(n15297) );
AND2_X2 U10880 ( .A1(n15307), .A2(n15308), .ZN(n15127) );
NAND2_X2 U10881 ( .A1(dii_data[31]), .A2(n15309), .ZN(n15308) );
NAND2_X2 U10882 ( .A1(n17882), .A2(dii_data[63]), .ZN(n15307) );
NAND2_X2 U10883 ( .A1(n17857), .A2(dii_data[55]), .ZN(n15302) );
NAND2_X2 U10884 ( .A1(n14945), .A2(n17893), .ZN(n15301) );
AND3_X2 U10885 ( .A1(n15310), .A2(n17881), .A3(n15311), .ZN(n14945) );
NAND2_X2 U10886 ( .A1(n19159), .A2(n18073), .ZN(n15311) );
NAND2_X2 U10887 ( .A1(n19127), .A2(dii_data_size[2]), .ZN(n15310) );
NAND2_X2 U10888 ( .A1(n15312), .A2(n15313), .ZN(n14773) );
NAND2_X2 U10889 ( .A1(dii_data[71]), .A2(n18074), .ZN(n15313) );
NAND2_X2 U10890 ( .A1(dii_data[7]), .A2(n18075), .ZN(n15312) );
NAND2_X2 U10891 ( .A1(n19202), .A2(n17713), .ZN(n15300) );
NAND2_X2 U10892 ( .A1(n18041), .A2(b_in[63]), .ZN(n15288) );
NAND2_X2 U10893 ( .A1(n15314), .A2(n15315), .ZN(N3149) );
NAND2_X2 U10894 ( .A1(n15316), .A2(n18066), .ZN(n15315) );
XNOR2_X2 U10895 ( .A(n18973), .B(n15317), .ZN(n15316) );
NAND2_X2 U10897 ( .A1(n17922), .A2(n15321), .ZN(n13746) );
XNOR2_X2 U10898 ( .A(n19108), .B(aes_text_out[78]), .ZN(n15321) );
XNOR2_X2 U10900 ( .A(n15322), .B(aes_text_out[78]), .ZN(n13748) );
NAND2_X2 U10902 ( .A1(n15323), .A2(n15324), .ZN(n15318) );
NAND2_X2 U10903 ( .A1(n17997), .A2(aad_byte_cnt[11]), .ZN(n15324) );
NAND2_X2 U10904 ( .A1(n17911), .A2(n15322), .ZN(n15323) );
NAND4_X2 U10905 ( .A1(n15325), .A2(n15326), .A3(n15327), .A4(n15328), .ZN(n15322) );
AND2_X2 U10910 ( .A1(n15332), .A2(n15333), .ZN(n15149) );
NAND2_X2 U10911 ( .A1(dii_data[30]), .A2(n15309), .ZN(n15333) );
NAND2_X2 U10912 ( .A1(n17882), .A2(dii_data[62]), .ZN(n15332) );
NAND2_X2 U10913 ( .A1(n17859), .A2(dii_data[54]), .ZN(n15327) );
NAND2_X2 U10914 ( .A1(n14968), .A2(n17893), .ZN(n15326) );
AND3_X2 U10915 ( .A1(n15334), .A2(n17881), .A3(n15335), .ZN(n14968) );
NAND2_X2 U10916 ( .A1(n19160), .A2(n18073), .ZN(n15335) );
NAND2_X2 U10917 ( .A1(n19128), .A2(dii_data_size[2]), .ZN(n15334) );
NAND2_X2 U10918 ( .A1(n15336), .A2(n15337), .ZN(n14795) );
NAND2_X2 U10919 ( .A1(dii_data[6]), .A2(n18075), .ZN(n15337) );
NAND2_X2 U10920 ( .A1(dii_data[70]), .A2(n18074), .ZN(n15336) );
NAND2_X2 U10921 ( .A1(n19202), .A2(n17715), .ZN(n15325) );
NAND2_X2 U10922 ( .A1(n18041), .A2(b_in[62]), .ZN(n15314) );
NAND2_X2 U10923 ( .A1(n15338), .A2(n15339), .ZN(N3148) );
NAND2_X2 U10924 ( .A1(n15340), .A2(n18066), .ZN(n15339) );
XNOR2_X2 U10925 ( .A(n18972), .B(n15341), .ZN(n15340) );
NAND2_X2 U10927 ( .A1(n17922), .A2(n15345), .ZN(n13740) );
XNOR2_X2 U10928 ( .A(n19111), .B(aes_text_out[77]), .ZN(n15345) );
XNOR2_X2 U10930 ( .A(n15346), .B(aes_text_out[77]), .ZN(n13742) );
NAND2_X2 U10932 ( .A1(n15347), .A2(n15348), .ZN(n15342) );
NAND2_X2 U10933 ( .A1(n17998), .A2(aad_byte_cnt[10]), .ZN(n15348) );
NAND2_X2 U10934 ( .A1(n17911), .A2(n15346), .ZN(n15347) );
NAND4_X2 U10935 ( .A1(n15349), .A2(n15350), .A3(n15351), .A4(n15352), .ZN(n15346) );
AND2_X2 U10940 ( .A1(n15356), .A2(n15357), .ZN(n15171) );
NAND2_X2 U10941 ( .A1(dii_data[29]), .A2(n15309), .ZN(n15357) );
NAND2_X2 U10942 ( .A1(n17883), .A2(dii_data[61]), .ZN(n15356) );
NAND2_X2 U10943 ( .A1(n17859), .A2(dii_data[53]), .ZN(n15351) );
NAND2_X2 U10944 ( .A1(n14990), .A2(n17892), .ZN(n15350) );
AND3_X2 U10945 ( .A1(n15358), .A2(n17881), .A3(n15359), .ZN(n14990) );
NAND2_X2 U10946 ( .A1(n19161), .A2(n18073), .ZN(n15359) );
NAND2_X2 U10947 ( .A1(n19129), .A2(dii_data_size[2]), .ZN(n15358) );
NAND2_X2 U10948 ( .A1(n15360), .A2(n15361), .ZN(n14817) );
NAND2_X2 U10949 ( .A1(dii_data[5]), .A2(n18075), .ZN(n15361) );
NAND2_X2 U10950 ( .A1(dii_data[69]), .A2(n18074), .ZN(n15360) );
NAND2_X2 U10951 ( .A1(n19202), .A2(n17717), .ZN(n15349) );
NAND2_X2 U10952 ( .A1(n18041), .A2(b_in[61]), .ZN(n15338) );
NAND2_X2 U10953 ( .A1(n15362), .A2(n15363), .ZN(N3147) );
NAND2_X2 U10954 ( .A1(n15364), .A2(n18066), .ZN(n15363) );
XNOR2_X2 U10955 ( .A(n18971), .B(n15365), .ZN(n15364) );
NAND2_X2 U10957 ( .A1(n17922), .A2(n15369), .ZN(n13734) );
XNOR2_X2 U10958 ( .A(n19114), .B(aes_text_out[76]), .ZN(n15369) );
XNOR2_X2 U10960 ( .A(n15370), .B(aes_text_out[76]), .ZN(n13736) );
NAND2_X2 U10962 ( .A1(n15371), .A2(n15372), .ZN(n15366) );
NAND2_X2 U10963 ( .A1(n17998), .A2(aad_byte_cnt[9]), .ZN(n15372) );
NAND2_X2 U10964 ( .A1(n17911), .A2(n15370), .ZN(n15371) );
NAND4_X2 U10965 ( .A1(n15373), .A2(n15374), .A3(n15375), .A4(n15376), .ZN(n15370) );
AND2_X2 U10970 ( .A1(n15380), .A2(n15381), .ZN(n15193) );
NAND2_X2 U10971 ( .A1(dii_data[28]), .A2(n15309), .ZN(n15381) );
NAND2_X2 U10972 ( .A1(n17882), .A2(dii_data[60]), .ZN(n15380) );
NAND2_X2 U10973 ( .A1(n17859), .A2(dii_data[52]), .ZN(n15375) );
NAND2_X2 U10974 ( .A1(n15012), .A2(n17892), .ZN(n15374) );
AND3_X2 U10975 ( .A1(n15382), .A2(n17881), .A3(n15383), .ZN(n15012) );
NAND2_X2 U10976 ( .A1(n19162), .A2(n18073), .ZN(n15383) );
NAND2_X2 U10977 ( .A1(n19130), .A2(dii_data_size[2]), .ZN(n15382) );
NAND2_X2 U10978 ( .A1(n15384), .A2(n15385), .ZN(n14839) );
NAND2_X2 U10979 ( .A1(dii_data[4]), .A2(n18075), .ZN(n15385) );
NAND2_X2 U10980 ( .A1(dii_data[68]), .A2(n18074), .ZN(n15384) );
NAND2_X2 U10981 ( .A1(n19202), .A2(n17719), .ZN(n15373) );
NAND2_X2 U10982 ( .A1(n18040), .A2(b_in[60]), .ZN(n15362) );
NAND2_X2 U10983 ( .A1(n15386), .A2(n15387), .ZN(N3146) );
NAND2_X2 U10984 ( .A1(n15388), .A2(n18066), .ZN(n15387) );
XNOR2_X2 U10985 ( .A(n18970), .B(n15389), .ZN(n15388) );
NAND2_X2 U10987 ( .A1(n17923), .A2(n15393), .ZN(n13728) );
XNOR2_X2 U10988 ( .A(n19117), .B(aes_text_out[75]), .ZN(n15393) );
XNOR2_X2 U10990 ( .A(n15394), .B(aes_text_out[75]), .ZN(n13730) );
NAND2_X2 U10992 ( .A1(n15395), .A2(n15396), .ZN(n15390) );
NAND2_X2 U10993 ( .A1(n17998), .A2(aad_byte_cnt[8]), .ZN(n15396) );
NAND2_X2 U10994 ( .A1(n17911), .A2(n15394), .ZN(n15395) );
NAND4_X2 U10995 ( .A1(n15397), .A2(n15398), .A3(n15399), .A4(n15400), .ZN(n15394) );
AND2_X2 U11000 ( .A1(n15404), .A2(n15405), .ZN(n15215) );
NAND2_X2 U11001 ( .A1(dii_data[27]), .A2(n15309), .ZN(n15405) );
NAND2_X2 U11002 ( .A1(n17882), .A2(dii_data[59]), .ZN(n15404) );
NAND2_X2 U11003 ( .A1(n17859), .A2(dii_data[51]), .ZN(n15399) );
NAND2_X2 U11004 ( .A1(n15034), .A2(n17892), .ZN(n15398) );
AND3_X2 U11005 ( .A1(n15406), .A2(n17881), .A3(n15407), .ZN(n15034) );
NAND2_X2 U11006 ( .A1(n19163), .A2(n18073), .ZN(n15407) );
NAND2_X2 U11007 ( .A1(n19131), .A2(dii_data_size[2]), .ZN(n15406) );
NAND2_X2 U11008 ( .A1(n15408), .A2(n15409), .ZN(n14861) );
NAND2_X2 U11009 ( .A1(dii_data[3]), .A2(n18075), .ZN(n15409) );
NAND2_X2 U11010 ( .A1(dii_data[67]), .A2(n18074), .ZN(n15408) );
NAND2_X2 U11011 ( .A1(n19202), .A2(n17721), .ZN(n15397) );
NAND2_X2 U11012 ( .A1(n18040), .A2(b_in[59]), .ZN(n15386) );
NAND2_X2 U11013 ( .A1(n15410), .A2(n15411), .ZN(N3145) );
NAND2_X2 U11014 ( .A1(n15412), .A2(n18066), .ZN(n15411) );
XNOR2_X2 U11015 ( .A(n18969), .B(n15413), .ZN(n15412) );
NAND2_X2 U11017 ( .A1(n17923), .A2(n15417), .ZN(n13722) );
XNOR2_X2 U11018 ( .A(n19120), .B(aes_text_out[74]), .ZN(n15417) );
XNOR2_X2 U11020 ( .A(n15418), .B(aes_text_out[74]), .ZN(n13724) );
NAND2_X2 U11022 ( .A1(n15419), .A2(n15420), .ZN(n15414) );
NAND2_X2 U11023 ( .A1(n17998), .A2(aad_byte_cnt[7]), .ZN(n15420) );
NAND2_X2 U11024 ( .A1(n17911), .A2(n15418), .ZN(n15419) );
NAND4_X2 U11025 ( .A1(n15421), .A2(n15422), .A3(n15423), .A4(n15424), .ZN(n15418) );
AND2_X2 U11030 ( .A1(n15428), .A2(n15429), .ZN(n15237) );
NAND2_X2 U11031 ( .A1(dii_data[26]), .A2(n15309), .ZN(n15429) );
NAND2_X2 U11032 ( .A1(n17882), .A2(dii_data[58]), .ZN(n15428) );
NAND2_X2 U11033 ( .A1(n17859), .A2(dii_data[50]), .ZN(n15423) );
NAND2_X2 U11034 ( .A1(n15056), .A2(n17892), .ZN(n15422) );
AND3_X2 U11035 ( .A1(n15430), .A2(n17881), .A3(n15431), .ZN(n15056) );
NAND2_X2 U11036 ( .A1(n19164), .A2(n18073), .ZN(n15431) );
NAND2_X2 U11037 ( .A1(n19132), .A2(dii_data_size[2]), .ZN(n15430) );
NAND2_X2 U11038 ( .A1(n15432), .A2(n15433), .ZN(n14883) );
NAND2_X2 U11039 ( .A1(dii_data[2]), .A2(n18075), .ZN(n15433) );
NAND2_X2 U11040 ( .A1(dii_data[66]), .A2(n18074), .ZN(n15432) );
NAND2_X2 U11041 ( .A1(n19202), .A2(n17723), .ZN(n15421) );
NAND2_X2 U11042 ( .A1(n18040), .A2(b_in[58]), .ZN(n15410) );
NAND2_X2 U11043 ( .A1(n15434), .A2(n15435), .ZN(N3144) );
NAND2_X2 U11044 ( .A1(n15436), .A2(n18066), .ZN(n15435) );
XNOR2_X2 U11045 ( .A(n18968), .B(n15437), .ZN(n15436) );
NAND2_X2 U11047 ( .A1(n17923), .A2(n15441), .ZN(n13716) );
XNOR2_X2 U11048 ( .A(n19123), .B(aes_text_out[73]), .ZN(n15441) );
XNOR2_X2 U11050 ( .A(n15442), .B(aes_text_out[73]), .ZN(n13718) );
NAND2_X2 U11052 ( .A1(n15443), .A2(n15444), .ZN(n15438) );
NAND2_X2 U11053 ( .A1(n17998), .A2(aad_byte_cnt[6]), .ZN(n15444) );
NAND2_X2 U11054 ( .A1(n17911), .A2(n15442), .ZN(n15443) );
NAND4_X2 U11055 ( .A1(n15445), .A2(n15446), .A3(n15447), .A4(n15448), .ZN(n15442) );
AND2_X2 U11060 ( .A1(n15452), .A2(n15453), .ZN(n15259) );
NAND2_X2 U11061 ( .A1(dii_data[25]), .A2(n15309), .ZN(n15453) );
NAND2_X2 U11062 ( .A1(n17882), .A2(dii_data[57]), .ZN(n15452) );
NAND2_X2 U11063 ( .A1(n17859), .A2(dii_data[49]), .ZN(n15447) );
NAND2_X2 U11064 ( .A1(n15078), .A2(n17892), .ZN(n15446) );
AND3_X2 U11065 ( .A1(n15454), .A2(n17881), .A3(n15455), .ZN(n15078) );
NAND2_X2 U11066 ( .A1(n19165), .A2(n18073), .ZN(n15455) );
NAND2_X2 U11067 ( .A1(n19133), .A2(dii_data_size[2]), .ZN(n15454) );
NAND2_X2 U11068 ( .A1(n15456), .A2(n15457), .ZN(n14905) );
NAND2_X2 U11069 ( .A1(dii_data[1]), .A2(n18075), .ZN(n15457) );
NAND2_X2 U11070 ( .A1(dii_data[65]), .A2(n18074), .ZN(n15456) );
NAND2_X2 U11071 ( .A1(n19202), .A2(n17725), .ZN(n15445) );
NAND2_X2 U11072 ( .A1(n18040), .A2(b_in[57]), .ZN(n15434) );
NAND2_X2 U11073 ( .A1(n15458), .A2(n15459), .ZN(N3143) );
NAND2_X2 U11074 ( .A1(n15460), .A2(n18066), .ZN(n15459) );
XNOR2_X2 U11075 ( .A(n18967), .B(n15461), .ZN(n15460) );
NAND2_X2 U11077 ( .A1(n17923), .A2(n15465), .ZN(n13710) );
XNOR2_X2 U11078 ( .A(n19126), .B(aes_text_out[72]), .ZN(n15465) );
NAND2_X2 U11080 ( .A1(n17934), .A2(n15466), .ZN(n15296) );
NAND2_X2 U11081 ( .A1(n15272), .A2(n15467), .ZN(n15466) );
NAND2_X2 U11082 ( .A1(n17892), .A2(dii_data_size[2]), .ZN(n15467) );
XNOR2_X2 U11083 ( .A(n15468), .B(aes_text_out[72]), .ZN(n13712) );
NAND2_X2 U11085 ( .A1(n15469), .A2(n15470), .ZN(n15462) );
NAND2_X2 U11086 ( .A1(n17998), .A2(aad_byte_cnt[5]), .ZN(n15470) );
NAND2_X2 U11087 ( .A1(n17911), .A2(n15468), .ZN(n15469) );
NAND4_X2 U11088 ( .A1(n15471), .A2(n15472), .A3(n15473), .A4(n15474), .ZN(n15468) );
AND2_X2 U11094 ( .A1(n15478), .A2(n15479), .ZN(n15283) );
NAND2_X2 U11095 ( .A1(dii_data[24]), .A2(n15309), .ZN(n15479) );
NAND2_X2 U11096 ( .A1(n17882), .A2(dii_data[56]), .ZN(n15478) );
NAND2_X2 U11097 ( .A1(n17859), .A2(dii_data[48]), .ZN(n15473) );
NAND2_X2 U11098 ( .A1(n15102), .A2(n17892), .ZN(n15472) );
AND3_X2 U11099 ( .A1(n15480), .A2(n17881), .A3(n15481), .ZN(n15102) );
NAND2_X2 U11100 ( .A1(n19166), .A2(n18071), .ZN(n15481) );
NAND2_X2 U11102 ( .A1(n19134), .A2(dii_data_size[2]), .ZN(n15480) );
NAND2_X2 U11103 ( .A1(n15482), .A2(n15483), .ZN(n14928) );
NAND2_X2 U11104 ( .A1(dii_data[0]), .A2(n18075), .ZN(n15483) );
NAND2_X2 U11105 ( .A1(dii_data[64]), .A2(n18074), .ZN(n15482) );
NAND2_X2 U11106 ( .A1(n19202), .A2(n17727), .ZN(n15471) );
NAND2_X2 U11107 ( .A1(n18040), .A2(b_in[56]), .ZN(n15458) );
NAND2_X2 U11108 ( .A1(n15484), .A2(n15485), .ZN(N3142) );
NAND2_X2 U11109 ( .A1(n15486), .A2(n18066), .ZN(n15485) );
XNOR2_X2 U11110 ( .A(n18966), .B(n15487), .ZN(n15486) );
XOR2_X2 U11114 ( .A(aes_text_out[71]), .B(n15491), .Z(n13706) );
AND4_X2 U11115 ( .A1(n15493), .A2(n15494), .A3(n15495), .A4(n15496), .ZN(n15491) );
NAND2_X2 U11124 ( .A1(n17848), .A2(dii_data[63]), .ZN(n15494) );
NAND2_X2 U11125 ( .A1(n15509), .A2(dii_data[7]), .ZN(n15493) );
NAND2_X2 U11126 ( .A1(n15510), .A2(n15511), .ZN(n15488) );
NAND2_X2 U11127 ( .A1(n17906), .A2(dii_data[71]), .ZN(n15511) );
NAND2_X2 U11128 ( .A1(n17998), .A2(aad_byte_cnt[4]), .ZN(n15510) );
NAND2_X2 U11129 ( .A1(n17923), .A2(n15512), .ZN(n13704) );
XOR2_X2 U11130 ( .A(n17617), .B(aes_text_out[71]), .Z(n15512) );
NAND2_X2 U11131 ( .A1(n18040), .A2(b_in[55]), .ZN(n15484) );
NAND2_X2 U11132 ( .A1(n15513), .A2(n15514), .ZN(N3141) );
NAND2_X2 U11133 ( .A1(n15515), .A2(n18066), .ZN(n15514) );
XNOR2_X2 U11134 ( .A(n18965), .B(n15516), .ZN(n15515) );
XOR2_X2 U11138 ( .A(aes_text_out[70]), .B(n15520), .Z(n13700) );
AND4_X2 U11139 ( .A1(n15521), .A2(n15522), .A3(n15523), .A4(n15524), .ZN(n15520) );
NAND2_X2 U11148 ( .A1(n17848), .A2(dii_data[62]), .ZN(n15522) );
NAND2_X2 U11149 ( .A1(n15509), .A2(dii_data[6]), .ZN(n15521) );
NAND2_X2 U11151 ( .A1(n17906), .A2(dii_data[70]), .ZN(n15532) );
NAND2_X2 U11153 ( .A1(n17923), .A2(n15533), .ZN(n13698) );
XOR2_X2 U11154 ( .A(n17619), .B(aes_text_out[70]), .Z(n15533) );
NAND2_X2 U11155 ( .A1(n18040), .A2(b_in[54]), .ZN(n15513) );
NAND2_X2 U11156 ( .A1(n15534), .A2(n15535), .ZN(N3140) );
NAND2_X2 U11157 ( .A1(n15536), .A2(n18067), .ZN(n15535) );
XNOR2_X2 U11158 ( .A(n18964), .B(n15537), .ZN(n15536) );
XOR2_X2 U11162 ( .A(aes_text_out[69]), .B(n15541), .Z(n13694) );
AND4_X2 U11163 ( .A1(n15542), .A2(n15543), .A3(n15544), .A4(n15545), .ZN(n15541) );
NAND2_X2 U11172 ( .A1(n17848), .A2(dii_data[61]), .ZN(n15543) );
NAND2_X2 U11173 ( .A1(n15509), .A2(dii_data[5]), .ZN(n15542) );
NAND2_X2 U11175 ( .A1(n17906), .A2(dii_data[69]), .ZN(n15553) );
NAND2_X2 U11177 ( .A1(n17923), .A2(n15554), .ZN(n13692) );
XOR2_X2 U11178 ( .A(n17621), .B(aes_text_out[69]), .Z(n15554) );
NAND2_X2 U11179 ( .A1(n18040), .A2(b_in[53]), .ZN(n15534) );
NAND2_X2 U11180 ( .A1(n15555), .A2(n15556), .ZN(N3139) );
NAND2_X2 U11181 ( .A1(n15557), .A2(n18067), .ZN(n15556) );
XNOR2_X2 U11182 ( .A(n18963), .B(n15558), .ZN(n15557) );
XOR2_X2 U11186 ( .A(aes_text_out[68]), .B(n15562), .Z(n13688) );
AND4_X2 U11187 ( .A1(n15563), .A2(n15564), .A3(n15565), .A4(n15566), .ZN(n15562) );
NAND2_X2 U11196 ( .A1(n17848), .A2(dii_data[60]), .ZN(n15564) );
NAND2_X2 U11197 ( .A1(n15509), .A2(dii_data[4]), .ZN(n15563) );
NAND2_X2 U11199 ( .A1(n17906), .A2(dii_data[68]), .ZN(n15574) );
NAND2_X2 U11201 ( .A1(n17923), .A2(n15575), .ZN(n13686) );
XOR2_X2 U11202 ( .A(n17623), .B(aes_text_out[68]), .Z(n15575) );
NAND2_X2 U11203 ( .A1(n18040), .A2(b_in[52]), .ZN(n15555) );
NAND2_X2 U11204 ( .A1(n15576), .A2(n15577), .ZN(N3138) );
NAND2_X2 U11205 ( .A1(n15578), .A2(n18067), .ZN(n15577) );
XNOR2_X2 U11206 ( .A(n18962), .B(n15579), .ZN(n15578) );
XOR2_X2 U11210 ( .A(aes_text_out[67]), .B(n15583), .Z(n13682) );
AND4_X2 U11211 ( .A1(n15584), .A2(n15585), .A3(n15586), .A4(n15587), .ZN(n15583) );
NAND2_X2 U11220 ( .A1(n17848), .A2(dii_data[59]), .ZN(n15585) );
NAND2_X2 U11221 ( .A1(n15509), .A2(dii_data[3]), .ZN(n15584) );
NAND2_X2 U11223 ( .A1(n17906), .A2(dii_data[67]), .ZN(n15595) );
NAND2_X2 U11225 ( .A1(n17923), .A2(n15596), .ZN(n13680) );
XOR2_X2 U11226 ( .A(n17625), .B(aes_text_out[67]), .Z(n15596) );
NAND2_X2 U11227 ( .A1(n18040), .A2(b_in[51]), .ZN(n15576) );
NAND2_X2 U11228 ( .A1(n15597), .A2(n15598), .ZN(N3137) );
NAND2_X2 U11229 ( .A1(n15599), .A2(n18067), .ZN(n15598) );
XNOR2_X2 U11230 ( .A(n18961), .B(n15600), .ZN(n15599) );
AND2_X2 U11233 ( .A1(dii_data[66]), .A2(n17908), .ZN(n15603) );
XOR2_X2 U11235 ( .A(aes_text_out[66]), .B(n15605), .Z(n13676) );
AND4_X2 U11236 ( .A1(n15606), .A2(n15607), .A3(n15608), .A4(n15609), .ZN(n15605) );
OR2_X2 U11245 ( .A1(n17872), .A2(n19172), .ZN(n15607) );
NAND2_X2 U11246 ( .A1(n17848), .A2(dii_data[58]), .ZN(n15606) );
AND2_X2 U11247 ( .A1(n13675), .A2(n17930), .ZN(n15601) );
XOR2_X2 U11248 ( .A(aes_text_out[66]), .B(n17627), .Z(n13675) );
NAND2_X2 U11249 ( .A1(n18040), .A2(b_in[50]), .ZN(n15597) );
NAND2_X2 U11250 ( .A1(n15616), .A2(n15617), .ZN(N3136) );
NAND2_X2 U11251 ( .A1(n15618), .A2(n18067), .ZN(n15617) );
XNOR2_X2 U11252 ( .A(n18960), .B(n15619), .ZN(n15618) );
AND2_X2 U11255 ( .A1(dii_data[65]), .A2(n17908), .ZN(n15622) );
XOR2_X2 U11257 ( .A(aes_text_out[65]), .B(n15624), .Z(n13669) );
AND4_X2 U11258 ( .A1(n15625), .A2(n15626), .A3(n15627), .A4(n15628), .ZN(n15624) );
NAND2_X2 U11267 ( .A1(n17848), .A2(dii_data[57]), .ZN(n15626) );
NAND2_X2 U11268 ( .A1(n15509), .A2(dii_data[1]), .ZN(n15625) );
AND2_X2 U11269 ( .A1(n13668), .A2(n17930), .ZN(n15620) );
NAND2_X2 U11271 ( .A1(n18040), .A2(b_in[49]), .ZN(n15616) );
NAND2_X2 U11272 ( .A1(n15635), .A2(n15636), .ZN(N3135) );
NAND2_X2 U11273 ( .A1(n15637), .A2(n18067), .ZN(n15636) );
XNOR2_X2 U11274 ( .A(n18959), .B(n15638), .ZN(n15637) );
AND2_X2 U11277 ( .A1(dii_data[64]), .A2(n17908), .ZN(n15641) );
NAND2_X2 U11279 ( .A1(n17934), .A2(n19199), .ZN(n15492) );
XOR2_X2 U11281 ( .A(aes_text_out[64]), .B(n15643), .Z(n13662) );
AND4_X2 U11282 ( .A1(n15645), .A2(n15646), .A3(n15647), .A4(n15648), .ZN(n15643) );
NAND2_X2 U11291 ( .A1(n17848), .A2(dii_data[56]), .ZN(n15646) );
NAND2_X2 U11292 ( .A1(n15509), .A2(dii_data[0]), .ZN(n15645) );
AND2_X2 U11293 ( .A1(n13661), .A2(n17930), .ZN(n15639) );
XOR2_X2 U11294 ( .A(aes_text_out[64]), .B(n17631), .Z(n13661) );
NAND2_X2 U11295 ( .A1(n18040), .A2(b_in[48]), .ZN(n15635) );
NAND2_X2 U11296 ( .A1(n15655), .A2(n15656), .ZN(N3134) );
NAND2_X2 U11297 ( .A1(n15657), .A2(n18067), .ZN(n15656) );
XNOR2_X2 U11298 ( .A(n18958), .B(n15658), .ZN(n15657) );
XOR2_X2 U11302 ( .A(n15662), .B(aes_text_out[63]), .Z(n13654) );
AND4_X2 U11303 ( .A1(n15664), .A2(n15665), .A3(n15666), .A4(n15667), .ZN(n15662) );
NAND2_X2 U11309 ( .A1(n17848), .A2(dii_data[55]), .ZN(n15666) );
NAND2_X2 U11310 ( .A1(n17859), .A2(dii_data[39]), .ZN(n15665) );
NAND2_X2 U11311 ( .A1(n17852), .A2(dii_data[47]), .ZN(n15664) );
NAND2_X2 U11312 ( .A1(n15672), .A2(n15673), .ZN(n15659) );
NAND2_X2 U11313 ( .A1(n17906), .A2(dii_data[63]), .ZN(n15673) );
NAND2_X2 U11315 ( .A1(n17923), .A2(n15674), .ZN(n13652) );
XNOR2_X2 U11316 ( .A(n19135), .B(aes_text_out[63]), .ZN(n15674) );
NAND2_X2 U11317 ( .A1(n18040), .A2(b_in[47]), .ZN(n15655) );
NAND2_X2 U11318 ( .A1(n15675), .A2(n15676), .ZN(N3133) );
NAND2_X2 U11319 ( .A1(n15677), .A2(n18067), .ZN(n15676) );
XNOR2_X2 U11320 ( .A(n18957), .B(n15678), .ZN(n15677) );
XOR2_X2 U11324 ( .A(n15682), .B(aes_text_out[62]), .Z(n13648) );
AND4_X2 U11325 ( .A1(n15683), .A2(n15684), .A3(n15685), .A4(n15686), .ZN(n15682) );
NAND2_X2 U11331 ( .A1(n17849), .A2(dii_data[54]), .ZN(n15685) );
NAND2_X2 U11332 ( .A1(n17859), .A2(dii_data[38]), .ZN(n15684) );
NAND2_X2 U11333 ( .A1(n17852), .A2(dii_data[46]), .ZN(n15683) );
NAND2_X2 U11334 ( .A1(n15691), .A2(n15692), .ZN(n15679) );
NAND2_X2 U11335 ( .A1(n17906), .A2(dii_data[62]), .ZN(n15692) );
NAND2_X2 U11337 ( .A1(n17923), .A2(n15693), .ZN(n13646) );
XNOR2_X2 U11338 ( .A(n19136), .B(aes_text_out[62]), .ZN(n15693) );
NAND2_X2 U11339 ( .A1(n18040), .A2(b_in[46]), .ZN(n15675) );
NAND2_X2 U11340 ( .A1(n15694), .A2(n15695), .ZN(N3132) );
NAND2_X2 U11341 ( .A1(n15696), .A2(n18067), .ZN(n15695) );
XNOR2_X2 U11342 ( .A(n18956), .B(n15697), .ZN(n15696) );
XOR2_X2 U11346 ( .A(n15701), .B(aes_text_out[61]), .Z(n13642) );
AND4_X2 U11347 ( .A1(n15702), .A2(n15703), .A3(n15704), .A4(n15705), .ZN(n15701) );
NAND2_X2 U11353 ( .A1(n17849), .A2(dii_data[53]), .ZN(n15704) );
NAND2_X2 U11354 ( .A1(n17859), .A2(dii_data[37]), .ZN(n15703) );
NAND2_X2 U11355 ( .A1(n17852), .A2(dii_data[45]), .ZN(n15702) );
NAND2_X2 U11356 ( .A1(n15710), .A2(n15711), .ZN(n15698) );
NAND2_X2 U11357 ( .A1(n17906), .A2(dii_data[61]), .ZN(n15711) );
NAND2_X2 U11359 ( .A1(n17924), .A2(n15712), .ZN(n13640) );
XNOR2_X2 U11360 ( .A(n19137), .B(aes_text_out[61]), .ZN(n15712) );
NAND2_X2 U11361 ( .A1(n18040), .A2(b_in[45]), .ZN(n15694) );
NAND2_X2 U11362 ( .A1(n15713), .A2(n15714), .ZN(N3131) );
NAND2_X2 U11363 ( .A1(n15715), .A2(n18067), .ZN(n15714) );
XNOR2_X2 U11364 ( .A(n18955), .B(n15716), .ZN(n15715) );
XOR2_X2 U11368 ( .A(n15720), .B(aes_text_out[60]), .Z(n13636) );
AND4_X2 U11369 ( .A1(n15721), .A2(n15722), .A3(n15723), .A4(n15724), .ZN(n15720) );
NAND2_X2 U11375 ( .A1(n17849), .A2(dii_data[52]), .ZN(n15723) );
NAND2_X2 U11376 ( .A1(n17859), .A2(dii_data[36]), .ZN(n15722) );
NAND2_X2 U11377 ( .A1(n17852), .A2(dii_data[44]), .ZN(n15721) );
NAND2_X2 U11378 ( .A1(n15729), .A2(n15730), .ZN(n15717) );
NAND2_X2 U11379 ( .A1(n17906), .A2(dii_data[60]), .ZN(n15730) );
NAND2_X2 U11381 ( .A1(n17924), .A2(n15731), .ZN(n13634) );
XNOR2_X2 U11382 ( .A(n19138), .B(aes_text_out[60]), .ZN(n15731) );
NAND2_X2 U11383 ( .A1(n18039), .A2(b_in[44]), .ZN(n15713) );
NAND2_X2 U11384 ( .A1(n15732), .A2(n15733), .ZN(N3130) );
NAND2_X2 U11385 ( .A1(n15734), .A2(n18067), .ZN(n15733) );
XNOR2_X2 U11386 ( .A(n18954), .B(n15735), .ZN(n15734) );
XOR2_X2 U11390 ( .A(n15739), .B(aes_text_out[59]), .Z(n13630) );
AND4_X2 U11391 ( .A1(n15740), .A2(n15741), .A3(n15742), .A4(n15743), .ZN(n15739) );
NAND2_X2 U11397 ( .A1(n17849), .A2(dii_data[51]), .ZN(n15742) );
NAND2_X2 U11398 ( .A1(n17859), .A2(dii_data[35]), .ZN(n15741) );
NAND2_X2 U11399 ( .A1(n17852), .A2(dii_data[43]), .ZN(n15740) );
NAND2_X2 U11400 ( .A1(n15748), .A2(n15749), .ZN(n15736) );
NAND2_X2 U11401 ( .A1(n17906), .A2(dii_data[59]), .ZN(n15749) );
NAND2_X2 U11403 ( .A1(n17924), .A2(n15750), .ZN(n13628) );
XNOR2_X2 U11404 ( .A(n19139), .B(aes_text_out[59]), .ZN(n15750) );
NAND2_X2 U11405 ( .A1(n18039), .A2(b_in[43]), .ZN(n15732) );
NAND2_X2 U11406 ( .A1(n15751), .A2(n15752), .ZN(N3129) );
NAND2_X2 U11407 ( .A1(n15753), .A2(n18067), .ZN(n15752) );
XNOR2_X2 U11408 ( .A(n18953), .B(n15754), .ZN(n15753) );
XOR2_X2 U11412 ( .A(n15758), .B(aes_text_out[58]), .Z(n13624) );
AND4_X2 U11413 ( .A1(n15759), .A2(n15760), .A3(n15761), .A4(n15762), .ZN(n15758) );
NAND2_X2 U11419 ( .A1(n17849), .A2(dii_data[50]), .ZN(n15761) );
NAND2_X2 U11420 ( .A1(n17858), .A2(dii_data[34]), .ZN(n15760) );
NAND2_X2 U11421 ( .A1(n17852), .A2(dii_data[42]), .ZN(n15759) );
NAND2_X2 U11422 ( .A1(n15767), .A2(n15768), .ZN(n15755) );
NAND2_X2 U11423 ( .A1(n17906), .A2(dii_data[58]), .ZN(n15768) );
NAND2_X2 U11425 ( .A1(n17924), .A2(n15769), .ZN(n13622) );
XNOR2_X2 U11426 ( .A(n19140), .B(aes_text_out[58]), .ZN(n15769) );
NAND2_X2 U11427 ( .A1(n18039), .A2(b_in[42]), .ZN(n15751) );
NAND2_X2 U11428 ( .A1(n15770), .A2(n15771), .ZN(N3128) );
NAND2_X2 U11429 ( .A1(n15772), .A2(n18067), .ZN(n15771) );
XNOR2_X2 U11430 ( .A(n18952), .B(n15773), .ZN(n15772) );
XOR2_X2 U11434 ( .A(n15777), .B(aes_text_out[57]), .Z(n13618) );
AND4_X2 U11435 ( .A1(n15778), .A2(n15779), .A3(n15780), .A4(n15781), .ZN(n15777) );
NAND2_X2 U11441 ( .A1(n17849), .A2(dii_data[49]), .ZN(n15780) );
NAND2_X2 U11442 ( .A1(n17858), .A2(dii_data[33]), .ZN(n15779) );
NAND2_X2 U11443 ( .A1(n17852), .A2(dii_data[41]), .ZN(n15778) );
NAND2_X2 U11444 ( .A1(n15786), .A2(n15787), .ZN(n15774) );
NAND2_X2 U11445 ( .A1(n17906), .A2(dii_data[57]), .ZN(n15787) );
NAND2_X2 U11447 ( .A1(n17924), .A2(n15788), .ZN(n13616) );
XNOR2_X2 U11448 ( .A(n19141), .B(aes_text_out[57]), .ZN(n15788) );
NAND2_X2 U11449 ( .A1(n18039), .A2(b_in[41]), .ZN(n15770) );
NAND2_X2 U11450 ( .A1(n15789), .A2(n15790), .ZN(N3127) );
NAND2_X2 U11451 ( .A1(n15791), .A2(n18067), .ZN(n15790) );
XNOR2_X2 U11452 ( .A(n18951), .B(n15792), .ZN(n15791) );
XOR2_X2 U11456 ( .A(n15796), .B(aes_text_out[56]), .Z(n13612) );
AND4_X2 U11457 ( .A1(n15797), .A2(n15798), .A3(n15799), .A4(n15800), .ZN(n15796) );
NAND2_X2 U11463 ( .A1(n17849), .A2(dii_data[48]), .ZN(n15799) );
NAND2_X2 U11464 ( .A1(n17858), .A2(dii_data[32]), .ZN(n15798) );
NAND2_X2 U11465 ( .A1(n17852), .A2(dii_data[40]), .ZN(n15797) );
AND2_X2 U11467 ( .A1(n19202), .A2(n17945), .ZN(n15806) );
NAND2_X2 U11469 ( .A1(n15807), .A2(n15808), .ZN(n15793) );
NAND2_X2 U11470 ( .A1(n17906), .A2(dii_data[56]), .ZN(n15808) );
NAND2_X2 U11472 ( .A1(n17924), .A2(n15809), .ZN(n13610) );
XNOR2_X2 U11473 ( .A(n19142), .B(aes_text_out[56]), .ZN(n15809) );
NAND2_X2 U11474 ( .A1(n18039), .A2(b_in[40]), .ZN(n15789) );
NAND2_X2 U11475 ( .A1(n15810), .A2(n15811), .ZN(N3126) );
NAND2_X2 U11476 ( .A1(n15812), .A2(n18067), .ZN(n15811) );
XNOR2_X2 U11477 ( .A(n18950), .B(n15813), .ZN(n15812) );
NAND2_X2 U11481 ( .A1(n17924), .A2(n15817), .ZN(n13604) );
XNOR2_X2 U11482 ( .A(n19143), .B(aes_text_out[55]), .ZN(n15817) );
NAND2_X2 U11483 ( .A1(n15818), .A2(n15819), .ZN(n15814) );
NAND2_X2 U11484 ( .A1(n13606), .A2(n15805), .ZN(n15819) );
XOR2_X2 U11485 ( .A(n15820), .B(aes_text_out[55]), .Z(n13606) );
NAND2_X2 U11486 ( .A1(n17911), .A2(n15820), .ZN(n15818) );
NAND4_X2 U11487 ( .A1(n15821), .A2(n15822), .A3(n15823), .A4(n15824), .ZN(n15820) );
NAND2_X2 U11492 ( .A1(n17849), .A2(dii_data[47]), .ZN(n15823) );
NAND2_X2 U11493 ( .A1(n17858), .A2(dii_data[31]), .ZN(n15822) );
NAND2_X2 U11494 ( .A1(n17852), .A2(n17681), .ZN(n15821) );
NAND2_X2 U11495 ( .A1(n18039), .A2(b_in[39]), .ZN(n15810) );
NAND2_X2 U11496 ( .A1(n15828), .A2(n15829), .ZN(N3125) );
NAND2_X2 U11497 ( .A1(n15830), .A2(n18067), .ZN(n15829) );
XNOR2_X2 U11498 ( .A(n18949), .B(n15831), .ZN(n15830) );
NAND2_X2 U11502 ( .A1(n17924), .A2(n15835), .ZN(n13598) );
XNOR2_X2 U11503 ( .A(n19144), .B(aes_text_out[54]), .ZN(n15835) );
NAND2_X2 U11504 ( .A1(n15836), .A2(n15837), .ZN(n15832) );
NAND2_X2 U11505 ( .A1(n13600), .A2(n15805), .ZN(n15837) );
XOR2_X2 U11506 ( .A(n15838), .B(aes_text_out[54]), .Z(n13600) );
NAND2_X2 U11507 ( .A1(n17911), .A2(n15838), .ZN(n15836) );
NAND4_X2 U11508 ( .A1(n15839), .A2(n15840), .A3(n15841), .A4(n15842), .ZN(n15838) );
NAND2_X2 U11513 ( .A1(n17849), .A2(dii_data[46]), .ZN(n15841) );
NAND2_X2 U11514 ( .A1(n17858), .A2(dii_data[30]), .ZN(n15840) );
NAND2_X2 U11515 ( .A1(n17852), .A2(n17683), .ZN(n15839) );
NAND2_X2 U11516 ( .A1(n18039), .A2(b_in[38]), .ZN(n15828) );
NAND2_X2 U11517 ( .A1(n15846), .A2(n15847), .ZN(N3124) );
NAND2_X2 U11518 ( .A1(n15848), .A2(n18067), .ZN(n15847) );
XNOR2_X2 U11519 ( .A(n18948), .B(n15849), .ZN(n15848) );
NAND2_X2 U11523 ( .A1(n17924), .A2(n15853), .ZN(n13592) );
XNOR2_X2 U11524 ( .A(n19145), .B(aes_text_out[53]), .ZN(n15853) );
NAND2_X2 U11525 ( .A1(n15854), .A2(n15855), .ZN(n15850) );
NAND2_X2 U11526 ( .A1(n13594), .A2(n15805), .ZN(n15855) );
XOR2_X2 U11527 ( .A(n15856), .B(aes_text_out[53]), .Z(n13594) );
NAND2_X2 U11528 ( .A1(n17911), .A2(n15856), .ZN(n15854) );
NAND4_X2 U11529 ( .A1(n15857), .A2(n15858), .A3(n15859), .A4(n15860), .ZN(n15856) );
NAND2_X2 U11534 ( .A1(n17849), .A2(dii_data[45]), .ZN(n15859) );
NAND2_X2 U11535 ( .A1(n17858), .A2(dii_data[29]), .ZN(n15858) );
NAND2_X2 U11536 ( .A1(n17852), .A2(n17685), .ZN(n15857) );
NAND2_X2 U11537 ( .A1(n18039), .A2(b_in[37]), .ZN(n15846) );
NAND2_X2 U11538 ( .A1(n15864), .A2(n15865), .ZN(N3123) );
NAND2_X2 U11539 ( .A1(n15866), .A2(n18067), .ZN(n15865) );
XNOR2_X2 U11540 ( .A(n18947), .B(n15867), .ZN(n15866) );
NAND2_X2 U11544 ( .A1(n17925), .A2(n15871), .ZN(n13586) );
XNOR2_X2 U11545 ( .A(n19146), .B(aes_text_out[52]), .ZN(n15871) );
NAND2_X2 U11546 ( .A1(n15872), .A2(n15873), .ZN(n15868) );
NAND2_X2 U11547 ( .A1(n13588), .A2(n15805), .ZN(n15873) );
XOR2_X2 U11548 ( .A(n15874), .B(aes_text_out[52]), .Z(n13588) );
NAND2_X2 U11549 ( .A1(n17910), .A2(n15874), .ZN(n15872) );
NAND4_X2 U11550 ( .A1(n15875), .A2(n15876), .A3(n15877), .A4(n15878), .ZN(n15874) );
NAND2_X2 U11555 ( .A1(n17849), .A2(dii_data[44]), .ZN(n15877) );
NAND2_X2 U11556 ( .A1(n17858), .A2(dii_data[28]), .ZN(n15876) );
NAND2_X2 U11557 ( .A1(n17853), .A2(n17687), .ZN(n15875) );
NAND2_X2 U11558 ( .A1(n18039), .A2(b_in[36]), .ZN(n15864) );
NAND2_X2 U11559 ( .A1(n15882), .A2(n15883), .ZN(N3122) );
NAND2_X2 U11560 ( .A1(n15884), .A2(n18067), .ZN(n15883) );
XNOR2_X2 U11561 ( .A(n18946), .B(n15885), .ZN(n15884) );
NAND2_X2 U11565 ( .A1(n17925), .A2(n15889), .ZN(n13580) );
XNOR2_X2 U11566 ( .A(n19147), .B(aes_text_out[51]), .ZN(n15889) );
NAND2_X2 U11567 ( .A1(n15890), .A2(n15891), .ZN(n15886) );
NAND2_X2 U11568 ( .A1(n13582), .A2(n15805), .ZN(n15891) );
XOR2_X2 U11569 ( .A(n15892), .B(aes_text_out[51]), .Z(n13582) );
NAND2_X2 U11570 ( .A1(n17910), .A2(n15892), .ZN(n15890) );
NAND4_X2 U11571 ( .A1(n15893), .A2(n15894), .A3(n15895), .A4(n15896), .ZN(n15892) );
NAND2_X2 U11576 ( .A1(n17849), .A2(dii_data[43]), .ZN(n15895) );
NAND2_X2 U11577 ( .A1(n17858), .A2(dii_data[27]), .ZN(n15894) );
NAND2_X2 U11578 ( .A1(n17853), .A2(n17689), .ZN(n15893) );
NAND2_X2 U11579 ( .A1(n18039), .A2(b_in[35]), .ZN(n15882) );
NAND2_X2 U11580 ( .A1(n15900), .A2(n15901), .ZN(N3121) );
NAND2_X2 U11581 ( .A1(n15902), .A2(n18067), .ZN(n15901) );
XNOR2_X2 U11582 ( .A(n18945), .B(n15903), .ZN(n15902) );
NAND2_X2 U11586 ( .A1(n17925), .A2(n15907), .ZN(n13574) );
XNOR2_X2 U11587 ( .A(n19148), .B(aes_text_out[50]), .ZN(n15907) );
NAND2_X2 U11588 ( .A1(n15908), .A2(n15909), .ZN(n15904) );
NAND2_X2 U11589 ( .A1(n13576), .A2(n15805), .ZN(n15909) );
XOR2_X2 U11590 ( .A(n15910), .B(aes_text_out[50]), .Z(n13576) );
NAND2_X2 U11591 ( .A1(n17910), .A2(n15910), .ZN(n15908) );
NAND4_X2 U11592 ( .A1(n15911), .A2(n15912), .A3(n15913), .A4(n15914), .ZN(n15910) );
NAND2_X2 U11597 ( .A1(n17849), .A2(dii_data[42]), .ZN(n15913) );
NAND2_X2 U11598 ( .A1(n17858), .A2(dii_data[26]), .ZN(n15912) );
NAND2_X2 U11599 ( .A1(n17853), .A2(n17691), .ZN(n15911) );
NAND2_X2 U11600 ( .A1(n18039), .A2(b_in[34]), .ZN(n15900) );
NAND2_X2 U11601 ( .A1(n15918), .A2(n15919), .ZN(N3120) );
NAND2_X2 U11602 ( .A1(n15920), .A2(n18067), .ZN(n15919) );
XNOR2_X2 U11603 ( .A(n18944), .B(n15921), .ZN(n15920) );
NAND2_X2 U11607 ( .A1(n17925), .A2(n15925), .ZN(n13568) );
XNOR2_X2 U11608 ( .A(n19149), .B(aes_text_out[49]), .ZN(n15925) );
NAND2_X2 U11609 ( .A1(n15926), .A2(n15927), .ZN(n15922) );
NAND2_X2 U11610 ( .A1(n13570), .A2(n15805), .ZN(n15927) );
XOR2_X2 U11611 ( .A(n15928), .B(aes_text_out[49]), .Z(n13570) );
NAND2_X2 U11612 ( .A1(n17910), .A2(n15928), .ZN(n15926) );
NAND4_X2 U11613 ( .A1(n15929), .A2(n15930), .A3(n15931), .A4(n15932), .ZN(n15928) );
NAND2_X2 U11618 ( .A1(n17849), .A2(dii_data[41]), .ZN(n15931) );
NAND2_X2 U11619 ( .A1(n17858), .A2(dii_data[25]), .ZN(n15930) );
NAND2_X2 U11620 ( .A1(n17853), .A2(n17693), .ZN(n15929) );
NAND2_X2 U11621 ( .A1(n18039), .A2(b_in[33]), .ZN(n15918) );
NAND2_X2 U11622 ( .A1(n15936), .A2(n15937), .ZN(N3119) );
NAND2_X2 U11623 ( .A1(n15938), .A2(n18068), .ZN(n15937) );
XNOR2_X2 U11624 ( .A(n18943), .B(n15939), .ZN(n15938) );
NAND2_X2 U11628 ( .A1(n17925), .A2(n15943), .ZN(n13562) );
XNOR2_X2 U11629 ( .A(n19150), .B(aes_text_out[48]), .ZN(n15943) );
NAND2_X2 U11630 ( .A1(n15944), .A2(n15945), .ZN(n15940) );
NAND2_X2 U11631 ( .A1(n13564), .A2(n15805), .ZN(n15945) );
NAND2_X2 U11633 ( .A1(n17755), .A2(n17945), .ZN(n15947) );
XOR2_X2 U11634 ( .A(n15948), .B(aes_text_out[48]), .Z(n13564) );
NAND2_X2 U11635 ( .A1(n17910), .A2(n15948), .ZN(n15944) );
NAND4_X2 U11636 ( .A1(n15949), .A2(n15950), .A3(n15951), .A4(n15952), .ZN(n15948) );
NAND2_X2 U11643 ( .A1(n17849), .A2(dii_data[40]), .ZN(n15951) );
NAND2_X2 U11644 ( .A1(n17858), .A2(dii_data[24]), .ZN(n15950) );
NAND2_X2 U11645 ( .A1(n17853), .A2(n17695), .ZN(n15949) );
NAND2_X2 U11646 ( .A1(n18039), .A2(b_in[32]), .ZN(n15936) );
NAND2_X2 U11647 ( .A1(n15956), .A2(n15957), .ZN(N3118) );
NAND2_X2 U11648 ( .A1(n15958), .A2(n18068), .ZN(n15957) );
XNOR2_X2 U11649 ( .A(n18942), .B(n15959), .ZN(n15958) );
XOR2_X2 U11653 ( .A(n15963), .B(aes_text_out[47]), .Z(n13558) );
AND4_X2 U11654 ( .A1(n15964), .A2(n15965), .A3(n15966), .A4(n15967), .ZN(n15963) );
NAND2_X2 U11655 ( .A1(n17858), .A2(dii_data[23]), .ZN(n15967) );
NAND2_X2 U11659 ( .A1(n17853), .A2(dii_data[31]), .ZN(n15965) );
NAND2_X2 U11660 ( .A1(n17849), .A2(dii_data[39]), .ZN(n15964) );
NAND2_X2 U11661 ( .A1(n15970), .A2(n15971), .ZN(n15960) );
NAND2_X2 U11662 ( .A1(n17907), .A2(dii_data[47]), .ZN(n15971) );
NAND2_X2 U11663 ( .A1(n17998), .A2(enc_byte_cnt[44]), .ZN(n15970) );
NAND2_X2 U11664 ( .A1(n17924), .A2(n15972), .ZN(n13556) );
XNOR2_X2 U11665 ( .A(n19151), .B(aes_text_out[47]), .ZN(n15972) );
NAND2_X2 U11666 ( .A1(n18039), .A2(b_in[31]), .ZN(n15956) );
NAND2_X2 U11667 ( .A1(n15973), .A2(n15974), .ZN(N3117) );
NAND2_X2 U11668 ( .A1(n15975), .A2(n18068), .ZN(n15974) );
XNOR2_X2 U11669 ( .A(n18941), .B(n15976), .ZN(n15975) );
XOR2_X2 U11673 ( .A(n15980), .B(aes_text_out[46]), .Z(n13552) );
AND4_X2 U11674 ( .A1(n15981), .A2(n15982), .A3(n15983), .A4(n15984), .ZN(n15980) );
NAND2_X2 U11675 ( .A1(n17858), .A2(dii_data[22]), .ZN(n15984) );
NAND2_X2 U11679 ( .A1(n17853), .A2(dii_data[30]), .ZN(n15982) );
NAND2_X2 U11680 ( .A1(n17850), .A2(dii_data[38]), .ZN(n15981) );
NAND2_X2 U11681 ( .A1(n15987), .A2(n15988), .ZN(n15977) );
NAND2_X2 U11682 ( .A1(n17907), .A2(dii_data[46]), .ZN(n15988) );
NAND2_X2 U11683 ( .A1(n17998), .A2(enc_byte_cnt[43]), .ZN(n15987) );
NAND2_X2 U11684 ( .A1(n17925), .A2(n15989), .ZN(n13550) );
XNOR2_X2 U11685 ( .A(n19152), .B(aes_text_out[46]), .ZN(n15989) );
NAND2_X2 U11686 ( .A1(n18039), .A2(b_in[30]), .ZN(n15973) );
NAND2_X2 U11687 ( .A1(n15990), .A2(n15991), .ZN(N3116) );
NAND2_X2 U11688 ( .A1(n15992), .A2(n18068), .ZN(n15991) );
XNOR2_X2 U11689 ( .A(n18940), .B(n15993), .ZN(n15992) );
XOR2_X2 U11693 ( .A(n15997), .B(aes_text_out[45]), .Z(n13546) );
AND4_X2 U11694 ( .A1(n15998), .A2(n15999), .A3(n16000), .A4(n16001), .ZN(n15997) );
NAND2_X2 U11695 ( .A1(n17858), .A2(dii_data[21]), .ZN(n16001) );
NAND2_X2 U11699 ( .A1(n17853), .A2(dii_data[29]), .ZN(n15999) );
NAND2_X2 U11700 ( .A1(n17850), .A2(dii_data[37]), .ZN(n15998) );
NAND2_X2 U11701 ( .A1(n16004), .A2(n16005), .ZN(n15994) );
NAND2_X2 U11702 ( .A1(n17907), .A2(dii_data[45]), .ZN(n16005) );
NAND2_X2 U11703 ( .A1(n17998), .A2(enc_byte_cnt[42]), .ZN(n16004) );
NAND2_X2 U11704 ( .A1(n17925), .A2(n16006), .ZN(n13544) );
XNOR2_X2 U11705 ( .A(n19153), .B(aes_text_out[45]), .ZN(n16006) );
NAND2_X2 U11706 ( .A1(n18039), .A2(b_in[29]), .ZN(n15990) );
NAND2_X2 U11707 ( .A1(n16007), .A2(n16008), .ZN(N3115) );
NAND2_X2 U11708 ( .A1(n16009), .A2(n18068), .ZN(n16008) );
XNOR2_X2 U11709 ( .A(n18939), .B(n16010), .ZN(n16009) );
XOR2_X2 U11713 ( .A(n16014), .B(aes_text_out[44]), .Z(n13540) );
AND4_X2 U11714 ( .A1(n16015), .A2(n16016), .A3(n16017), .A4(n16018), .ZN(n16014) );
NAND2_X2 U11715 ( .A1(n17858), .A2(dii_data[20]), .ZN(n16018) );
NAND2_X2 U11719 ( .A1(n17853), .A2(dii_data[28]), .ZN(n16016) );
NAND2_X2 U11720 ( .A1(n17850), .A2(dii_data[36]), .ZN(n16015) );
NAND2_X2 U11721 ( .A1(n16021), .A2(n16022), .ZN(n16011) );
NAND2_X2 U11722 ( .A1(n17907), .A2(dii_data[44]), .ZN(n16022) );
NAND2_X2 U11723 ( .A1(n17998), .A2(enc_byte_cnt[41]), .ZN(n16021) );
NAND2_X2 U11724 ( .A1(n17925), .A2(n16023), .ZN(n13538) );
XNOR2_X2 U11725 ( .A(n19154), .B(aes_text_out[44]), .ZN(n16023) );
NAND2_X2 U11726 ( .A1(n18039), .A2(b_in[28]), .ZN(n16007) );
NAND2_X2 U11727 ( .A1(n16024), .A2(n16025), .ZN(N3114) );
NAND2_X2 U11728 ( .A1(n16026), .A2(n18068), .ZN(n16025) );
XNOR2_X2 U11729 ( .A(n18938), .B(n16027), .ZN(n16026) );
XOR2_X2 U11733 ( .A(n16031), .B(aes_text_out[43]), .Z(n13534) );
AND4_X2 U11734 ( .A1(n16032), .A2(n16033), .A3(n16034), .A4(n16035), .ZN(n16031) );
NAND2_X2 U11735 ( .A1(n17858), .A2(dii_data[19]), .ZN(n16035) );
NAND2_X2 U11739 ( .A1(n17853), .A2(dii_data[27]), .ZN(n16033) );
NAND2_X2 U11740 ( .A1(n17850), .A2(dii_data[35]), .ZN(n16032) );
NAND2_X2 U11741 ( .A1(n16038), .A2(n16039), .ZN(n16028) );
NAND2_X2 U11742 ( .A1(n17907), .A2(dii_data[43]), .ZN(n16039) );
NAND2_X2 U11743 ( .A1(n17998), .A2(enc_byte_cnt[40]), .ZN(n16038) );
NAND2_X2 U11744 ( .A1(n17925), .A2(n16040), .ZN(n13532) );
XNOR2_X2 U11745 ( .A(n19155), .B(aes_text_out[43]), .ZN(n16040) );
NAND2_X2 U11746 ( .A1(n18038), .A2(b_in[27]), .ZN(n16024) );
NAND2_X2 U11747 ( .A1(n16041), .A2(n16042), .ZN(N3113) );
NAND2_X2 U11748 ( .A1(n16043), .A2(n18068), .ZN(n16042) );
XNOR2_X2 U11749 ( .A(n18937), .B(n16044), .ZN(n16043) );
XOR2_X2 U11753 ( .A(n16048), .B(aes_text_out[42]), .Z(n13528) );
AND4_X2 U11754 ( .A1(n16049), .A2(n16050), .A3(n16051), .A4(n16052), .ZN(n16048) );
NAND2_X2 U11755 ( .A1(n17858), .A2(dii_data[18]), .ZN(n16052) );
NAND2_X2 U11759 ( .A1(n17853), .A2(dii_data[26]), .ZN(n16050) );
NAND2_X2 U11760 ( .A1(n17850), .A2(dii_data[34]), .ZN(n16049) );
NAND2_X2 U11761 ( .A1(n16055), .A2(n16056), .ZN(n16045) );
NAND2_X2 U11762 ( .A1(n17907), .A2(dii_data[42]), .ZN(n16056) );
NAND2_X2 U11763 ( .A1(n17998), .A2(enc_byte_cnt[39]), .ZN(n16055) );
NAND2_X2 U11764 ( .A1(n17926), .A2(n16057), .ZN(n13526) );
XNOR2_X2 U11765 ( .A(n19156), .B(aes_text_out[42]), .ZN(n16057) );
NAND2_X2 U11766 ( .A1(n18038), .A2(b_in[26]), .ZN(n16041) );
NAND2_X2 U11767 ( .A1(n16058), .A2(n16059), .ZN(N3112) );
NAND2_X2 U11768 ( .A1(n16060), .A2(n18068), .ZN(n16059) );
XNOR2_X2 U11769 ( .A(n18936), .B(n16061), .ZN(n16060) );
XOR2_X2 U11773 ( .A(n16065), .B(aes_text_out[41]), .Z(n13522) );
AND4_X2 U11774 ( .A1(n16066), .A2(n16067), .A3(n16068), .A4(n16069), .ZN(n16065) );
NAND2_X2 U11775 ( .A1(n17858), .A2(dii_data[17]), .ZN(n16069) );
NAND2_X2 U11779 ( .A1(n17854), .A2(dii_data[25]), .ZN(n16067) );
NAND2_X2 U11780 ( .A1(n17850), .A2(dii_data[33]), .ZN(n16066) );
NAND2_X2 U11781 ( .A1(n16072), .A2(n16073), .ZN(n16062) );
NAND2_X2 U11782 ( .A1(n17907), .A2(dii_data[41]), .ZN(n16073) );
NAND2_X2 U11783 ( .A1(n17998), .A2(enc_byte_cnt[38]), .ZN(n16072) );
NAND2_X2 U11784 ( .A1(n17925), .A2(n16074), .ZN(n13520) );
XNOR2_X2 U11785 ( .A(n19157), .B(aes_text_out[41]), .ZN(n16074) );
NAND2_X2 U11786 ( .A1(n18038), .A2(b_in[25]), .ZN(n16058) );
NAND2_X2 U11787 ( .A1(n16075), .A2(n16076), .ZN(N3111) );
NAND2_X2 U11788 ( .A1(n16077), .A2(n18068), .ZN(n16076) );
XNOR2_X2 U11789 ( .A(n18935), .B(n16078), .ZN(n16077) );
NAND4_X2 U11794 ( .A1(n17872), .A2(n17876), .A3(n16083), .A4(n15507), .ZN(n15644) );
XOR2_X2 U11796 ( .A(n16082), .B(aes_text_out[40]), .Z(n13516) );
AND4_X2 U11797 ( .A1(n16084), .A2(n16085), .A3(n16086), .A4(n16087), .ZN(n16082) );
NAND2_X2 U11798 ( .A1(n17857), .A2(dii_data[16]), .ZN(n16087) );
NAND2_X2 U11804 ( .A1(n17854), .A2(dii_data[24]), .ZN(n16085) );
NAND2_X2 U11805 ( .A1(n17850), .A2(dii_data[32]), .ZN(n16084) );
NAND2_X2 U11806 ( .A1(n16090), .A2(n16091), .ZN(n16079) );
NAND2_X2 U11807 ( .A1(n17907), .A2(dii_data[40]), .ZN(n16091) );
NAND2_X2 U11808 ( .A1(n17998), .A2(enc_byte_cnt[37]), .ZN(n16090) );
NAND2_X2 U11809 ( .A1(n17926), .A2(n16092), .ZN(n13514) );
XNOR2_X2 U11810 ( .A(n19158), .B(aes_text_out[40]), .ZN(n16092) );
NAND2_X2 U11811 ( .A1(n18038), .A2(b_in[24]), .ZN(n16075) );
NAND2_X2 U11812 ( .A1(n16093), .A2(n16094), .ZN(N3110) );
NAND2_X2 U11813 ( .A1(n16095), .A2(n18068), .ZN(n16094) );
XNOR2_X2 U11814 ( .A(n18934), .B(n16096), .ZN(n16095) );
NAND2_X2 U11818 ( .A1(n17926), .A2(n16100), .ZN(n13508) );
XNOR2_X2 U11819 ( .A(n19159), .B(aes_text_out[39]), .ZN(n16100) );
NAND2_X2 U11820 ( .A1(n16101), .A2(n16102), .ZN(n16097) );
NAND2_X2 U11821 ( .A1(n13510), .A2(n16103), .ZN(n16102) );
XOR2_X2 U11822 ( .A(n16104), .B(aes_text_out[39]), .Z(n13510) );
NAND2_X2 U11823 ( .A1(n17910), .A2(n16104), .ZN(n16101) );
NAND4_X2 U11824 ( .A1(n16105), .A2(n16106), .A3(n16107), .A4(n16108), .ZN(n16104) );
NAND2_X2 U11825 ( .A1(n17873), .A2(dii_data[7]), .ZN(n16108) );
NAND2_X2 U11826 ( .A1(n17857), .A2(dii_data[15]), .ZN(n16107) );
NAND2_X2 U11827 ( .A1(n17854), .A2(dii_data[23]), .ZN(n16106) );
NAND2_X2 U11828 ( .A1(n17850), .A2(n17697), .ZN(n16105) );
NAND2_X2 U11829 ( .A1(n18038), .A2(b_in[23]), .ZN(n16093) );
NAND2_X2 U11830 ( .A1(n16109), .A2(n16110), .ZN(N3109) );
NAND2_X2 U11831 ( .A1(n16111), .A2(n18068), .ZN(n16110) );
XNOR2_X2 U11832 ( .A(n18933), .B(n16112), .ZN(n16111) );
NAND2_X2 U11836 ( .A1(n17926), .A2(n16116), .ZN(n13502) );
XNOR2_X2 U11837 ( .A(n19160), .B(aes_text_out[38]), .ZN(n16116) );
NAND2_X2 U11838 ( .A1(n16117), .A2(n16118), .ZN(n16113) );
NAND2_X2 U11839 ( .A1(n13504), .A2(n16103), .ZN(n16118) );
XOR2_X2 U11840 ( .A(n16119), .B(aes_text_out[38]), .Z(n13504) );
NAND2_X2 U11841 ( .A1(n17910), .A2(n16119), .ZN(n16117) );
NAND4_X2 U11842 ( .A1(n16120), .A2(n16121), .A3(n16122), .A4(n16123), .ZN(n16119) );
NAND2_X2 U11843 ( .A1(n17873), .A2(dii_data[6]), .ZN(n16123) );
NAND2_X2 U11844 ( .A1(n17857), .A2(dii_data[14]), .ZN(n16122) );
NAND2_X2 U11845 ( .A1(n17854), .A2(dii_data[22]), .ZN(n16121) );
NAND2_X2 U11846 ( .A1(n17850), .A2(n17699), .ZN(n16120) );
NAND2_X2 U11847 ( .A1(n18038), .A2(b_in[22]), .ZN(n16109) );
NAND2_X2 U11848 ( .A1(n16124), .A2(n16125), .ZN(N3108) );
NAND2_X2 U11849 ( .A1(n16126), .A2(n18068), .ZN(n16125) );
XNOR2_X2 U11850 ( .A(n18932), .B(n16127), .ZN(n16126) );
NAND2_X2 U11854 ( .A1(n17926), .A2(n16131), .ZN(n13496) );
XNOR2_X2 U11855 ( .A(n19161), .B(aes_text_out[37]), .ZN(n16131) );
NAND2_X2 U11856 ( .A1(n16132), .A2(n16133), .ZN(n16128) );
NAND2_X2 U11857 ( .A1(n13498), .A2(n16103), .ZN(n16133) );
XOR2_X2 U11858 ( .A(n16134), .B(aes_text_out[37]), .Z(n13498) );
NAND2_X2 U11859 ( .A1(n17910), .A2(n16134), .ZN(n16132) );
NAND4_X2 U11860 ( .A1(n16135), .A2(n16136), .A3(n16137), .A4(n16138), .ZN(n16134) );
NAND2_X2 U11861 ( .A1(n17873), .A2(dii_data[5]), .ZN(n16138) );
NAND2_X2 U11862 ( .A1(n17857), .A2(dii_data[13]), .ZN(n16137) );
NAND2_X2 U11863 ( .A1(n17854), .A2(dii_data[21]), .ZN(n16136) );
NAND2_X2 U11864 ( .A1(n17850), .A2(n17701), .ZN(n16135) );
NAND2_X2 U11865 ( .A1(n18038), .A2(b_in[21]), .ZN(n16124) );
NAND2_X2 U11866 ( .A1(n16139), .A2(n16140), .ZN(N3107) );
NAND2_X2 U11867 ( .A1(n16141), .A2(n18068), .ZN(n16140) );
XNOR2_X2 U11868 ( .A(n18931), .B(n16142), .ZN(n16141) );
NAND2_X2 U11872 ( .A1(n17926), .A2(n16146), .ZN(n13490) );
XNOR2_X2 U11873 ( .A(n19162), .B(aes_text_out[36]), .ZN(n16146) );
NAND2_X2 U11874 ( .A1(n16147), .A2(n16148), .ZN(n16143) );
NAND2_X2 U11875 ( .A1(n13492), .A2(n16103), .ZN(n16148) );
XOR2_X2 U11876 ( .A(n16149), .B(aes_text_out[36]), .Z(n13492) );
NAND2_X2 U11877 ( .A1(n17910), .A2(n16149), .ZN(n16147) );
NAND4_X2 U11878 ( .A1(n16150), .A2(n16151), .A3(n16152), .A4(n16153), .ZN(n16149) );
NAND2_X2 U11879 ( .A1(n17873), .A2(dii_data[4]), .ZN(n16153) );
NAND2_X2 U11880 ( .A1(n17857), .A2(dii_data[12]), .ZN(n16152) );
NAND2_X2 U11881 ( .A1(n17854), .A2(dii_data[20]), .ZN(n16151) );
NAND2_X2 U11882 ( .A1(n17850), .A2(n17703), .ZN(n16150) );
NAND2_X2 U11883 ( .A1(n18038), .A2(b_in[20]), .ZN(n16139) );
NAND2_X2 U11884 ( .A1(n16154), .A2(n16155), .ZN(N3106) );
NAND2_X2 U11885 ( .A1(n16156), .A2(n18068), .ZN(n16155) );
XNOR2_X2 U11886 ( .A(n18930), .B(n16157), .ZN(n16156) );
NAND2_X2 U11890 ( .A1(n17925), .A2(n16161), .ZN(n13484) );
XNOR2_X2 U11891 ( .A(n19163), .B(aes_text_out[35]), .ZN(n16161) );
NAND2_X2 U11892 ( .A1(n16162), .A2(n16163), .ZN(n16158) );
NAND2_X2 U11893 ( .A1(n13486), .A2(n16103), .ZN(n16163) );
XOR2_X2 U11894 ( .A(n16164), .B(aes_text_out[35]), .Z(n13486) );
NAND2_X2 U11895 ( .A1(n17910), .A2(n16164), .ZN(n16162) );
NAND4_X2 U11896 ( .A1(n16165), .A2(n16166), .A3(n16167), .A4(n16168), .ZN(n16164) );
NAND2_X2 U11897 ( .A1(n17873), .A2(dii_data[3]), .ZN(n16168) );
NAND2_X2 U11898 ( .A1(n17858), .A2(dii_data[11]), .ZN(n16167) );
NAND2_X2 U11899 ( .A1(n17854), .A2(dii_data[19]), .ZN(n16166) );
NAND2_X2 U11900 ( .A1(n17850), .A2(n17705), .ZN(n16165) );
NAND2_X2 U11901 ( .A1(n18038), .A2(b_in[19]), .ZN(n16154) );
NAND2_X2 U11902 ( .A1(n16169), .A2(n16170), .ZN(N3105) );
NAND2_X2 U11903 ( .A1(n16171), .A2(n18068), .ZN(n16170) );
XNOR2_X2 U11904 ( .A(n18929), .B(n16172), .ZN(n16171) );
NAND2_X2 U11908 ( .A1(n17926), .A2(n16176), .ZN(n13478) );
XNOR2_X2 U11909 ( .A(n19164), .B(aes_text_out[34]), .ZN(n16176) );
NAND2_X2 U11910 ( .A1(n16177), .A2(n16178), .ZN(n16173) );
NAND2_X2 U11911 ( .A1(n13480), .A2(n16103), .ZN(n16178) );
XOR2_X2 U11912 ( .A(n16179), .B(aes_text_out[34]), .Z(n13480) );
NAND2_X2 U11913 ( .A1(n17910), .A2(n16179), .ZN(n16177) );
NAND4_X2 U11914 ( .A1(n16180), .A2(n16181), .A3(n16182), .A4(n16183), .ZN(n16179) );
NAND2_X2 U11915 ( .A1(n17873), .A2(dii_data[2]), .ZN(n16183) );
NAND2_X2 U11916 ( .A1(n17857), .A2(dii_data[10]), .ZN(n16182) );
NAND2_X2 U11917 ( .A1(n17854), .A2(dii_data[18]), .ZN(n16181) );
NAND2_X2 U11918 ( .A1(n17850), .A2(n17707), .ZN(n16180) );
NAND2_X2 U11919 ( .A1(n18038), .A2(b_in[18]), .ZN(n16169) );
NAND2_X2 U11920 ( .A1(n16184), .A2(n16185), .ZN(N3104) );
NAND2_X2 U11921 ( .A1(n16186), .A2(n18068), .ZN(n16185) );
XNOR2_X2 U11922 ( .A(n18928), .B(n16187), .ZN(n16186) );
NAND2_X2 U11926 ( .A1(n17926), .A2(n16191), .ZN(n13472) );
XNOR2_X2 U11927 ( .A(n19165), .B(aes_text_out[33]), .ZN(n16191) );
NAND2_X2 U11928 ( .A1(n16192), .A2(n16193), .ZN(n16188) );
NAND2_X2 U11929 ( .A1(n13474), .A2(n16103), .ZN(n16193) );
XOR2_X2 U11930 ( .A(n16194), .B(aes_text_out[33]), .Z(n13474) );
NAND2_X2 U11931 ( .A1(n17909), .A2(n16194), .ZN(n16192) );
NAND4_X2 U11932 ( .A1(n16195), .A2(n16196), .A3(n16197), .A4(n16198), .ZN(n16194) );
NAND2_X2 U11933 ( .A1(n17873), .A2(dii_data[1]), .ZN(n16198) );
NAND2_X2 U11934 ( .A1(n17857), .A2(dii_data[9]), .ZN(n16197) );
NAND2_X2 U11935 ( .A1(n17854), .A2(dii_data[17]), .ZN(n16196) );
NAND2_X2 U11936 ( .A1(n17850), .A2(n17709), .ZN(n16195) );
NAND2_X2 U11937 ( .A1(n18038), .A2(b_in[17]), .ZN(n16184) );
NAND2_X2 U11938 ( .A1(n16199), .A2(n16200), .ZN(N3103) );
NAND2_X2 U11939 ( .A1(n16201), .A2(n18068), .ZN(n16200) );
XNOR2_X2 U11940 ( .A(n18927), .B(n16202), .ZN(n16201) );
NAND2_X2 U11944 ( .A1(n17926), .A2(n16206), .ZN(n13466) );
XNOR2_X2 U11945 ( .A(n19166), .B(aes_text_out[32]), .ZN(n16206) );
NAND2_X2 U11946 ( .A1(n16207), .A2(n16208), .ZN(n16203) );
NAND2_X2 U11947 ( .A1(n13468), .A2(n16103), .ZN(n16208) );
NAND2_X2 U11948 ( .A1(n16209), .A2(n16210), .ZN(n16103) );
NAND2_X2 U11949 ( .A1(n17873), .A2(n17945), .ZN(n16210) );
XOR2_X2 U11950 ( .A(n16211), .B(aes_text_out[32]), .Z(n13468) );
NAND2_X2 U11951 ( .A1(n17909), .A2(n16211), .ZN(n16207) );
NAND4_X2 U11952 ( .A1(n16212), .A2(n16213), .A3(n16214), .A4(n16215), .ZN(n16211) );
NAND2_X2 U11953 ( .A1(n17873), .A2(dii_data[0]), .ZN(n16215) );
NAND2_X2 U11954 ( .A1(n17897), .A2(n18074), .ZN(n15501) );
NAND2_X2 U11956 ( .A1(n17857), .A2(dii_data[8]), .ZN(n16214) );
NAND2_X2 U11957 ( .A1(n17854), .A2(dii_data[16]), .ZN(n16213) );
NAND2_X2 U11958 ( .A1(n17850), .A2(n17711), .ZN(n16212) );
NAND2_X2 U11959 ( .A1(n18040), .A2(b_in[16]), .ZN(n16199) );
NAND2_X2 U11960 ( .A1(n16216), .A2(n16217), .ZN(N3102) );
NAND2_X2 U11961 ( .A1(n16218), .A2(n18068), .ZN(n16217) );
XNOR2_X2 U11962 ( .A(n18926), .B(n16219), .ZN(n16218) );
XOR2_X2 U11966 ( .A(n16223), .B(aes_text_out[31]), .Z(n13462) );
AND3_X2 U11967 ( .A1(n16224), .A2(n16225), .A3(n16226), .ZN(n16223) );
NAND2_X2 U11968 ( .A1(n17850), .A2(dii_data[23]), .ZN(n16226) );
NAND2_X2 U11969 ( .A1(n17857), .A2(dii_data[7]), .ZN(n16225) );
NAND2_X2 U11970 ( .A1(n17854), .A2(dii_data[15]), .ZN(n16224) );
NAND2_X2 U11971 ( .A1(n16227), .A2(n16228), .ZN(n16220) );
NAND2_X2 U11972 ( .A1(n17907), .A2(dii_data[31]), .ZN(n16228) );
NAND2_X2 U11973 ( .A1(n17998), .A2(enc_byte_cnt[28]), .ZN(n16227) );
NAND2_X2 U11974 ( .A1(n17926), .A2(n16229), .ZN(n13460) );
XNOR2_X2 U11975 ( .A(n19167), .B(aes_text_out[31]), .ZN(n16229) );
NAND2_X2 U11976 ( .A1(n18038), .A2(b_in[15]), .ZN(n16216) );
NAND2_X2 U11977 ( .A1(n16230), .A2(n16231), .ZN(N3101) );
NAND2_X2 U11978 ( .A1(n16232), .A2(n18068), .ZN(n16231) );
XNOR2_X2 U11979 ( .A(n18925), .B(n16233), .ZN(n16232) );
XOR2_X2 U11983 ( .A(n16237), .B(aes_text_out[30]), .Z(n13456) );
AND3_X2 U11984 ( .A1(n16238), .A2(n16239), .A3(n16240), .ZN(n16237) );
NAND2_X2 U11985 ( .A1(n17850), .A2(dii_data[22]), .ZN(n16240) );
NAND2_X2 U11986 ( .A1(n17857), .A2(dii_data[6]), .ZN(n16239) );
NAND2_X2 U11987 ( .A1(n17855), .A2(dii_data[14]), .ZN(n16238) );
NAND2_X2 U11988 ( .A1(n16241), .A2(n16242), .ZN(n16234) );
NAND2_X2 U11989 ( .A1(n17907), .A2(dii_data[30]), .ZN(n16242) );
NAND2_X2 U11990 ( .A1(n17998), .A2(enc_byte_cnt[27]), .ZN(n16241) );
NAND2_X2 U11991 ( .A1(n17927), .A2(n16243), .ZN(n13454) );
XNOR2_X2 U11992 ( .A(n19168), .B(aes_text_out[30]), .ZN(n16243) );
NAND2_X2 U11993 ( .A1(n18038), .A2(b_in[14]), .ZN(n16230) );
NAND2_X2 U11994 ( .A1(n16244), .A2(n16245), .ZN(N3100) );
NAND2_X2 U11995 ( .A1(n16246), .A2(n18068), .ZN(n16245) );
XNOR2_X2 U11996 ( .A(n18924), .B(n16247), .ZN(n16246) );
XOR2_X2 U12000 ( .A(n16251), .B(aes_text_out[29]), .Z(n13450) );
AND3_X2 U12001 ( .A1(n16252), .A2(n16253), .A3(n16254), .ZN(n16251) );
NAND2_X2 U12002 ( .A1(n17851), .A2(dii_data[21]), .ZN(n16254) );
NAND2_X2 U12003 ( .A1(n17857), .A2(dii_data[5]), .ZN(n16253) );
NAND2_X2 U12004 ( .A1(n17855), .A2(dii_data[13]), .ZN(n16252) );
NAND2_X2 U12005 ( .A1(n16255), .A2(n16256), .ZN(n16248) );
NAND2_X2 U12006 ( .A1(n17907), .A2(dii_data[29]), .ZN(n16256) );
NAND2_X2 U12007 ( .A1(n17998), .A2(enc_byte_cnt[26]), .ZN(n16255) );
NAND2_X2 U12008 ( .A1(n17926), .A2(n16257), .ZN(n13448) );
XNOR2_X2 U12009 ( .A(n19169), .B(aes_text_out[29]), .ZN(n16257) );
NAND2_X2 U12010 ( .A1(n18038), .A2(b_in[13]), .ZN(n16244) );
NAND2_X2 U12011 ( .A1(n16258), .A2(n16259), .ZN(N3099) );
NAND2_X2 U12012 ( .A1(n16260), .A2(n18068), .ZN(n16259) );
XNOR2_X2 U12013 ( .A(n18923), .B(n16261), .ZN(n16260) );
XOR2_X2 U12017 ( .A(n16265), .B(aes_text_out[28]), .Z(n13444) );
AND3_X2 U12018 ( .A1(n16266), .A2(n16267), .A3(n16268), .ZN(n16265) );
NAND2_X2 U12019 ( .A1(n17851), .A2(dii_data[20]), .ZN(n16268) );
NAND2_X2 U12020 ( .A1(n17857), .A2(dii_data[4]), .ZN(n16267) );
NAND2_X2 U12021 ( .A1(n17855), .A2(dii_data[12]), .ZN(n16266) );
NAND2_X2 U12022 ( .A1(n16269), .A2(n16270), .ZN(n16262) );
NAND2_X2 U12023 ( .A1(n17907), .A2(dii_data[28]), .ZN(n16270) );
NAND2_X2 U12024 ( .A1(n17998), .A2(enc_byte_cnt[25]), .ZN(n16269) );
NAND2_X2 U12025 ( .A1(n17927), .A2(n16271), .ZN(n13442) );
XNOR2_X2 U12026 ( .A(n19170), .B(aes_text_out[28]), .ZN(n16271) );
NAND2_X2 U12027 ( .A1(n18038), .A2(b_in[12]), .ZN(n16258) );
NAND2_X2 U12028 ( .A1(n16272), .A2(n16273), .ZN(N3098) );
NAND2_X2 U12029 ( .A1(n16274), .A2(n18069), .ZN(n16273) );
XNOR2_X2 U12030 ( .A(n18922), .B(n16275), .ZN(n16274) );
XOR2_X2 U12034 ( .A(n16279), .B(aes_text_out[27]), .Z(n13438) );
AND3_X2 U12035 ( .A1(n16280), .A2(n16281), .A3(n16282), .ZN(n16279) );
NAND2_X2 U12036 ( .A1(n17851), .A2(dii_data[19]), .ZN(n16282) );
NAND2_X2 U12037 ( .A1(n17857), .A2(dii_data[3]), .ZN(n16281) );
NAND2_X2 U12038 ( .A1(n17855), .A2(dii_data[11]), .ZN(n16280) );
NAND2_X2 U12039 ( .A1(n16283), .A2(n16284), .ZN(n16276) );
NAND2_X2 U12040 ( .A1(n17907), .A2(dii_data[27]), .ZN(n16284) );
NAND2_X2 U12041 ( .A1(n17998), .A2(enc_byte_cnt[24]), .ZN(n16283) );
NAND2_X2 U12042 ( .A1(n17927), .A2(n16285), .ZN(n13436) );
XNOR2_X2 U12043 ( .A(n19171), .B(aes_text_out[27]), .ZN(n16285) );
NAND2_X2 U12044 ( .A1(n18038), .A2(b_in[11]), .ZN(n16272) );
NAND2_X2 U12045 ( .A1(n16286), .A2(n16287), .ZN(N3097) );
NAND2_X2 U12046 ( .A1(n16288), .A2(n18069), .ZN(n16287) );
XNOR2_X2 U12047 ( .A(n18921), .B(n16289), .ZN(n16288) );
XOR2_X2 U12051 ( .A(n16293), .B(aes_text_out[26]), .Z(n13432) );
AND3_X2 U12052 ( .A1(n16294), .A2(n16295), .A3(n16296), .ZN(n16293) );
NAND2_X2 U12053 ( .A1(n17851), .A2(dii_data[18]), .ZN(n16296) );
NAND2_X2 U12054 ( .A1(n17857), .A2(dii_data[2]), .ZN(n16295) );
NAND2_X2 U12055 ( .A1(n17855), .A2(dii_data[10]), .ZN(n16294) );
NAND2_X2 U12056 ( .A1(n16297), .A2(n16298), .ZN(n16290) );
NAND2_X2 U12057 ( .A1(n17907), .A2(dii_data[26]), .ZN(n16298) );
NAND2_X2 U12058 ( .A1(n17999), .A2(enc_byte_cnt[23]), .ZN(n16297) );
NAND2_X2 U12059 ( .A1(n17927), .A2(n16299), .ZN(n13430) );
XNOR2_X2 U12060 ( .A(n19172), .B(aes_text_out[26]), .ZN(n16299) );
NAND2_X2 U12061 ( .A1(n18038), .A2(b_in[10]), .ZN(n16286) );
NAND2_X2 U12062 ( .A1(n16300), .A2(n16301), .ZN(N3096) );
NAND2_X2 U12063 ( .A1(n16302), .A2(n18069), .ZN(n16301) );
XNOR2_X2 U12064 ( .A(n18920), .B(n16303), .ZN(n16302) );
XOR2_X2 U12068 ( .A(n16307), .B(aes_text_out[25]), .Z(n13426) );
AND3_X2 U12069 ( .A1(n16308), .A2(n16309), .A3(n16310), .ZN(n16307) );
NAND2_X2 U12070 ( .A1(n17851), .A2(dii_data[17]), .ZN(n16310) );
NAND2_X2 U12071 ( .A1(n17857), .A2(dii_data[1]), .ZN(n16309) );
NAND2_X2 U12072 ( .A1(n17855), .A2(dii_data[9]), .ZN(n16308) );
NAND2_X2 U12073 ( .A1(n16311), .A2(n16312), .ZN(n16304) );
NAND2_X2 U12074 ( .A1(n17907), .A2(dii_data[25]), .ZN(n16312) );
NAND2_X2 U12075 ( .A1(n17999), .A2(enc_byte_cnt[22]), .ZN(n16311) );
NAND2_X2 U12076 ( .A1(n17927), .A2(n16313), .ZN(n13424) );
XNOR2_X2 U12077 ( .A(n19173), .B(aes_text_out[25]), .ZN(n16313) );
NAND2_X2 U12078 ( .A1(n18037), .A2(b_in[9]), .ZN(n16300) );
NAND2_X2 U12079 ( .A1(n16314), .A2(n16315), .ZN(N3095) );
NAND2_X2 U12080 ( .A1(n16316), .A2(n18069), .ZN(n16315) );
XNOR2_X2 U12081 ( .A(n18919), .B(n16317), .ZN(n16316) );
XOR2_X2 U12085 ( .A(n16321), .B(aes_text_out[24]), .Z(n13420) );
AND3_X2 U12086 ( .A1(n16322), .A2(n16323), .A3(n16324), .ZN(n16321) );
NAND2_X2 U12087 ( .A1(n17851), .A2(dii_data[16]), .ZN(n16324) );
NAND2_X2 U12088 ( .A1(n17857), .A2(dii_data[0]), .ZN(n16323) );
NAND2_X2 U12089 ( .A1(n17855), .A2(dii_data[8]), .ZN(n16322) );
AND2_X2 U12091 ( .A1(n17859), .A2(n17945), .ZN(n16326) );
NAND2_X2 U12094 ( .A1(n16327), .A2(n16328), .ZN(n16318) );
NAND2_X2 U12095 ( .A1(n17907), .A2(dii_data[24]), .ZN(n16328) );
NAND2_X2 U12096 ( .A1(n17999), .A2(enc_byte_cnt[21]), .ZN(n16327) );
NAND2_X2 U12097 ( .A1(n17927), .A2(n16329), .ZN(n13418) );
XNOR2_X2 U12098 ( .A(n19174), .B(aes_text_out[24]), .ZN(n16329) );
NAND2_X2 U12099 ( .A1(n18037), .A2(b_in[8]), .ZN(n16314) );
NAND2_X2 U12100 ( .A1(n16330), .A2(n16331), .ZN(N3094) );
NAND2_X2 U12101 ( .A1(n16332), .A2(n18069), .ZN(n16331) );
XNOR2_X2 U12102 ( .A(n18918), .B(n16333), .ZN(n16332) );
NAND2_X2 U12106 ( .A1(n17927), .A2(n16337), .ZN(n13412) );
XNOR2_X2 U12107 ( .A(n19175), .B(aes_text_out[23]), .ZN(n16337) );
NAND2_X2 U12108 ( .A1(n16338), .A2(n16339), .ZN(n16334) );
NAND2_X2 U12109 ( .A1(n13414), .A2(n16325), .ZN(n16339) );
XOR2_X2 U12110 ( .A(n16340), .B(aes_text_out[23]), .Z(n13414) );
NAND2_X2 U12111 ( .A1(n17909), .A2(n16340), .ZN(n16338) );
NAND2_X2 U12112 ( .A1(n16341), .A2(n16342), .ZN(n16340) );
NAND2_X2 U12113 ( .A1(n17855), .A2(n17736), .ZN(n16342) );
NAND2_X2 U12114 ( .A1(n17851), .A2(n17728), .ZN(n16341) );
NAND2_X2 U12115 ( .A1(n18037), .A2(b_in[7]), .ZN(n16330) );
NAND2_X2 U12116 ( .A1(n16343), .A2(n16344), .ZN(N3093) );
NAND2_X2 U12117 ( .A1(n16345), .A2(n18069), .ZN(n16344) );
XNOR2_X2 U12118 ( .A(n18917), .B(n16346), .ZN(n16345) );
NAND2_X2 U12122 ( .A1(n17927), .A2(n16350), .ZN(n13406) );
XNOR2_X2 U12123 ( .A(n19176), .B(aes_text_out[22]), .ZN(n16350) );
NAND2_X2 U12124 ( .A1(n16351), .A2(n16352), .ZN(n16347) );
NAND2_X2 U12125 ( .A1(n13408), .A2(n16325), .ZN(n16352) );
XOR2_X2 U12126 ( .A(n16353), .B(aes_text_out[22]), .Z(n13408) );
NAND2_X2 U12127 ( .A1(n17909), .A2(n16353), .ZN(n16351) );
NAND2_X2 U12128 ( .A1(n16354), .A2(n16355), .ZN(n16353) );
NAND2_X2 U12129 ( .A1(n17855), .A2(n17737), .ZN(n16355) );
NAND2_X2 U12130 ( .A1(n17851), .A2(n17729), .ZN(n16354) );
NAND2_X2 U12131 ( .A1(n18037), .A2(b_in[6]), .ZN(n16343) );
NAND2_X2 U12132 ( .A1(n16356), .A2(n16357), .ZN(N3092) );
NAND2_X2 U12133 ( .A1(n16358), .A2(n18069), .ZN(n16357) );
XNOR2_X2 U12134 ( .A(n18916), .B(n16359), .ZN(n16358) );
NAND2_X2 U12138 ( .A1(n17927), .A2(n16363), .ZN(n13400) );
XNOR2_X2 U12139 ( .A(n19177), .B(aes_text_out[21]), .ZN(n16363) );
NAND2_X2 U12140 ( .A1(n16364), .A2(n16365), .ZN(n16360) );
NAND2_X2 U12141 ( .A1(n13402), .A2(n16325), .ZN(n16365) );
XOR2_X2 U12142 ( .A(n16366), .B(aes_text_out[21]), .Z(n13402) );
NAND2_X2 U12143 ( .A1(n17909), .A2(n16366), .ZN(n16364) );
NAND2_X2 U12144 ( .A1(n16367), .A2(n16368), .ZN(n16366) );
NAND2_X2 U12145 ( .A1(n17855), .A2(n17738), .ZN(n16368) );
NAND2_X2 U12146 ( .A1(n17851), .A2(n17730), .ZN(n16367) );
NAND2_X2 U12147 ( .A1(n18037), .A2(b_in[5]), .ZN(n16356) );
NAND2_X2 U12148 ( .A1(n16369), .A2(n16370), .ZN(N3091) );
NAND2_X2 U12149 ( .A1(n16371), .A2(n18069), .ZN(n16370) );
XNOR2_X2 U12150 ( .A(n18915), .B(n16372), .ZN(n16371) );
NAND2_X2 U12154 ( .A1(n17928), .A2(n16376), .ZN(n13394) );
XNOR2_X2 U12155 ( .A(n19178), .B(aes_text_out[20]), .ZN(n16376) );
NAND2_X2 U12156 ( .A1(n16377), .A2(n16378), .ZN(n16373) );
NAND2_X2 U12157 ( .A1(n13396), .A2(n16325), .ZN(n16378) );
XOR2_X2 U12158 ( .A(n16379), .B(aes_text_out[20]), .Z(n13396) );
NAND2_X2 U12159 ( .A1(n17909), .A2(n16379), .ZN(n16377) );
NAND2_X2 U12160 ( .A1(n16380), .A2(n16381), .ZN(n16379) );
NAND2_X2 U12161 ( .A1(n17855), .A2(n17739), .ZN(n16381) );
NAND2_X2 U12162 ( .A1(n17851), .A2(n17731), .ZN(n16380) );
NAND2_X2 U12163 ( .A1(n18037), .A2(b_in[4]), .ZN(n16369) );
NAND2_X2 U12164 ( .A1(n16382), .A2(n16383), .ZN(N3090) );
NAND2_X2 U12165 ( .A1(n16384), .A2(n18069), .ZN(n16383) );
XNOR2_X2 U12166 ( .A(n18914), .B(n16385), .ZN(n16384) );
NAND2_X2 U12170 ( .A1(n17927), .A2(n16389), .ZN(n13388) );
XNOR2_X2 U12171 ( .A(n19179), .B(aes_text_out[19]), .ZN(n16389) );
NAND2_X2 U12172 ( .A1(n16390), .A2(n16391), .ZN(n16386) );
NAND2_X2 U12173 ( .A1(n13390), .A2(n16325), .ZN(n16391) );
XOR2_X2 U12174 ( .A(n16392), .B(aes_text_out[19]), .Z(n13390) );
NAND2_X2 U12175 ( .A1(n17909), .A2(n16392), .ZN(n16390) );
NAND2_X2 U12176 ( .A1(n16393), .A2(n16394), .ZN(n16392) );
NAND2_X2 U12177 ( .A1(n17856), .A2(n17740), .ZN(n16394) );
NAND2_X2 U12178 ( .A1(n17851), .A2(n17732), .ZN(n16393) );
NAND2_X2 U12179 ( .A1(n18037), .A2(b_in[3]), .ZN(n16382) );
NAND2_X2 U12180 ( .A1(n16395), .A2(n16396), .ZN(N3089) );
NAND2_X2 U12181 ( .A1(n16397), .A2(n18069), .ZN(n16396) );
XNOR2_X2 U12182 ( .A(n18913), .B(n16398), .ZN(n16397) );
NAND2_X2 U12186 ( .A1(n17928), .A2(n16402), .ZN(n13382) );
XNOR2_X2 U12187 ( .A(n19180), .B(aes_text_out[18]), .ZN(n16402) );
NAND2_X2 U12188 ( .A1(n16403), .A2(n16404), .ZN(n16399) );
NAND2_X2 U12189 ( .A1(n13384), .A2(n16325), .ZN(n16404) );
XOR2_X2 U12190 ( .A(n16405), .B(aes_text_out[18]), .Z(n13384) );
NAND2_X2 U12191 ( .A1(n17909), .A2(n16405), .ZN(n16403) );
NAND2_X2 U12192 ( .A1(n16406), .A2(n16407), .ZN(n16405) );
NAND2_X2 U12193 ( .A1(n17856), .A2(n17741), .ZN(n16407) );
NAND2_X2 U12194 ( .A1(n17851), .A2(n17733), .ZN(n16406) );
NAND2_X2 U12195 ( .A1(n18037), .A2(b_in[2]), .ZN(n16395) );
NAND2_X2 U12196 ( .A1(n16408), .A2(n16409), .ZN(N3088) );
NAND2_X2 U12197 ( .A1(n16410), .A2(n18069), .ZN(n16409) );
XNOR2_X2 U12198 ( .A(n18912), .B(n16411), .ZN(n16410) );
NAND2_X2 U12202 ( .A1(n17927), .A2(n16415), .ZN(n13376) );
XNOR2_X2 U12203 ( .A(n19181), .B(aes_text_out[17]), .ZN(n16415) );
NAND2_X2 U12204 ( .A1(n16416), .A2(n16417), .ZN(n16412) );
NAND2_X2 U12205 ( .A1(n13378), .A2(n16325), .ZN(n16417) );
XOR2_X2 U12206 ( .A(n16418), .B(aes_text_out[17]), .Z(n13378) );
NAND2_X2 U12207 ( .A1(n17909), .A2(n16418), .ZN(n16416) );
NAND2_X2 U12208 ( .A1(n16419), .A2(n16420), .ZN(n16418) );
NAND2_X2 U12209 ( .A1(n17856), .A2(n17742), .ZN(n16420) );
NAND2_X2 U12210 ( .A1(n17851), .A2(n17734), .ZN(n16419) );
NAND2_X2 U12211 ( .A1(n18037), .A2(b_in[1]), .ZN(n16408) );
NAND2_X2 U12212 ( .A1(n16421), .A2(n16422), .ZN(N3087) );
NAND2_X2 U12213 ( .A1(n16423), .A2(n18064), .ZN(n16422) );
XNOR2_X2 U12214 ( .A(n18911), .B(n16424), .ZN(n16423) );
NAND2_X2 U12218 ( .A1(n17928), .A2(n16428), .ZN(n13370) );
XNOR2_X2 U12219 ( .A(n19182), .B(aes_text_out[16]), .ZN(n16428) );
NAND2_X2 U12220 ( .A1(n16429), .A2(n16430), .ZN(n16425) );
NAND2_X2 U12221 ( .A1(n13372), .A2(n16325), .ZN(n16430) );
NAND2_X2 U12223 ( .A1(n17856), .A2(n17945), .ZN(n16432) );
XOR2_X2 U12224 ( .A(n16433), .B(aes_text_out[16]), .Z(n13372) );
NAND2_X2 U12225 ( .A1(n17909), .A2(n16433), .ZN(n16429) );
NAND2_X2 U12226 ( .A1(n16434), .A2(n16435), .ZN(n16433) );
NAND2_X2 U12227 ( .A1(n17856), .A2(n17743), .ZN(n16435) );
NAND2_X2 U12229 ( .A1(n17851), .A2(n17735), .ZN(n16434) );
NAND2_X2 U12230 ( .A1(n18037), .A2(b_in[0]), .ZN(n16421) );
XNOR2_X2 U12232 ( .A(n16437), .B(n18910), .ZN(n16436) );
NAND2_X2 U12236 ( .A1(n16443), .A2(n16444), .ZN(n13365) );
NAND2_X2 U12237 ( .A1(n17933), .A2(n19191), .ZN(n16444) );
NAND2_X2 U12238 ( .A1(n16445), .A2(n16446), .ZN(n13364) );
NAND2_X2 U12240 ( .A1(n18634), .A2(n17736), .ZN(n16448) );
NAND2_X2 U12241 ( .A1(n17928), .A2(n17728), .ZN(n16447) );
NAND2_X2 U12242 ( .A1(aes_text_out[15]), .A2(n16449), .ZN(n16445) );
NAND2_X2 U12243 ( .A1(n17928), .A2(n19183), .ZN(n16449) );
NAND2_X2 U12245 ( .A1(n17907), .A2(n17728), .ZN(n16439) );
NAND2_X2 U12246 ( .A1(n17999), .A2(enc_byte_cnt[12]), .ZN(n16438) );
XNOR2_X2 U12248 ( .A(n16452), .B(n18909), .ZN(n16451) );
NAND2_X2 U12252 ( .A1(n16443), .A2(n16458), .ZN(n13359) );
NAND2_X2 U12253 ( .A1(n17933), .A2(n19192), .ZN(n16458) );
NAND2_X2 U12254 ( .A1(n16459), .A2(n16460), .ZN(n13358) );
NAND2_X2 U12256 ( .A1(n18634), .A2(n17737), .ZN(n16462) );
NAND2_X2 U12257 ( .A1(n17928), .A2(n17729), .ZN(n16461) );
NAND2_X2 U12258 ( .A1(aes_text_out[14]), .A2(n16463), .ZN(n16459) );
NAND2_X2 U12259 ( .A1(n17928), .A2(n19184), .ZN(n16463) );
NAND2_X2 U12261 ( .A1(n17908), .A2(n17729), .ZN(n16454) );
NAND2_X2 U12262 ( .A1(n17999), .A2(enc_byte_cnt[11]), .ZN(n16453) );
XNOR2_X2 U12264 ( .A(n16465), .B(n18908), .ZN(n16464) );
NAND2_X2 U12268 ( .A1(n16443), .A2(n16471), .ZN(n13353) );
NAND2_X2 U12269 ( .A1(n17933), .A2(n19193), .ZN(n16471) );
NAND2_X2 U12270 ( .A1(n16472), .A2(n16473), .ZN(n13352) );
NAND2_X2 U12272 ( .A1(n18634), .A2(n17738), .ZN(n16475) );
NAND2_X2 U12273 ( .A1(n17928), .A2(n17730), .ZN(n16474) );
NAND2_X2 U12274 ( .A1(aes_text_out[13]), .A2(n16476), .ZN(n16472) );
NAND2_X2 U12275 ( .A1(n17928), .A2(n19185), .ZN(n16476) );
NAND2_X2 U12277 ( .A1(n17907), .A2(n17730), .ZN(n16467) );
NAND2_X2 U12278 ( .A1(n17999), .A2(enc_byte_cnt[10]), .ZN(n16466) );
XNOR2_X2 U12280 ( .A(n16478), .B(n18907), .ZN(n16477) );
NAND2_X2 U12284 ( .A1(n16443), .A2(n16484), .ZN(n13347) );
NAND2_X2 U12285 ( .A1(n17933), .A2(n19194), .ZN(n16484) );
NAND2_X2 U12286 ( .A1(n16485), .A2(n16486), .ZN(n13346) );
NAND2_X2 U12288 ( .A1(n18634), .A2(n17739), .ZN(n16488) );
NAND2_X2 U12289 ( .A1(n17928), .A2(n17731), .ZN(n16487) );
NAND2_X2 U12290 ( .A1(aes_text_out[12]), .A2(n16489), .ZN(n16485) );
NAND2_X2 U12291 ( .A1(n17929), .A2(n19186), .ZN(n16489) );
NAND2_X2 U12293 ( .A1(n17908), .A2(n17731), .ZN(n16480) );
NAND2_X2 U12294 ( .A1(n17999), .A2(enc_byte_cnt[9]), .ZN(n16479) );
XNOR2_X2 U12296 ( .A(n16491), .B(n18906), .ZN(n16490) );
NAND2_X2 U12300 ( .A1(n16443), .A2(n16497), .ZN(n13341) );
NAND2_X2 U12301 ( .A1(n17933), .A2(n19195), .ZN(n16497) );
NAND2_X2 U12302 ( .A1(n16498), .A2(n16499), .ZN(n13340) );
NAND2_X2 U12304 ( .A1(n18634), .A2(n17740), .ZN(n16501) );
NAND2_X2 U12305 ( .A1(n17929), .A2(n17732), .ZN(n16500) );
NAND2_X2 U12306 ( .A1(aes_text_out[11]), .A2(n16502), .ZN(n16498) );
NAND2_X2 U12307 ( .A1(n17929), .A2(n19187), .ZN(n16502) );
NAND2_X2 U12309 ( .A1(n17907), .A2(n17732), .ZN(n16493) );
NAND2_X2 U12310 ( .A1(n17999), .A2(enc_byte_cnt[8]), .ZN(n16492) );
XNOR2_X2 U12312 ( .A(n16504), .B(n18905), .ZN(n16503) );
NAND2_X2 U12316 ( .A1(n16443), .A2(n16510), .ZN(n13335) );
NAND2_X2 U12317 ( .A1(n17933), .A2(n19196), .ZN(n16510) );
NAND2_X2 U12318 ( .A1(n16511), .A2(n16512), .ZN(n13334) );
NAND2_X2 U12320 ( .A1(n18634), .A2(n17741), .ZN(n16514) );
NAND2_X2 U12321 ( .A1(n17928), .A2(n17733), .ZN(n16513) );
NAND2_X2 U12322 ( .A1(aes_text_out[10]), .A2(n16515), .ZN(n16511) );
NAND2_X2 U12323 ( .A1(n17929), .A2(n19188), .ZN(n16515) );
NAND2_X2 U12325 ( .A1(n17908), .A2(n17733), .ZN(n16506) );
NAND2_X2 U12326 ( .A1(n17999), .A2(enc_byte_cnt[7]), .ZN(n16505) );
XNOR2_X2 U12328 ( .A(n16517), .B(n18904), .ZN(n16516) );
NAND2_X2 U12332 ( .A1(n16443), .A2(n16523), .ZN(n13329) );
NAND2_X2 U12333 ( .A1(n17933), .A2(n19197), .ZN(n16523) );
NAND2_X2 U12334 ( .A1(n16524), .A2(n16525), .ZN(n13328) );
NAND2_X2 U12336 ( .A1(n18634), .A2(n17742), .ZN(n16527) );
NAND2_X2 U12337 ( .A1(n17929), .A2(n17734), .ZN(n16526) );
NAND2_X2 U12338 ( .A1(aes_text_out[9]), .A2(n16528), .ZN(n16524) );
NAND2_X2 U12339 ( .A1(n17929), .A2(n19189), .ZN(n16528) );
NAND2_X2 U12341 ( .A1(n17907), .A2(n17734), .ZN(n16519) );
NAND2_X2 U12342 ( .A1(n17999), .A2(enc_byte_cnt[6]), .ZN(n16518) );
XNOR2_X2 U12344 ( .A(n16530), .B(n18903), .ZN(n16529) );
NAND2_X2 U12348 ( .A1(n16443), .A2(n16536), .ZN(n13323) );
NAND2_X2 U12349 ( .A1(n17933), .A2(n19198), .ZN(n16536) );
NAND2_X2 U12350 ( .A1(n17933), .A2(n16537), .ZN(n16443) );
NAND2_X2 U12351 ( .A1(n16538), .A2(n16539), .ZN(n13322) );
NAND2_X2 U12353 ( .A1(n18634), .A2(n17743), .ZN(n16541) );
NAND2_X2 U12354 ( .A1(n17851), .A2(n17936), .ZN(n16431) );
NAND2_X2 U12356 ( .A1(n17929), .A2(n17735), .ZN(n16540) );
NAND2_X2 U12357 ( .A1(aes_text_out[8]), .A2(n16543), .ZN(n16538) );
NAND2_X2 U12358 ( .A1(n17929), .A2(n19190), .ZN(n16543) );
NAND2_X2 U12360 ( .A1(n17909), .A2(n17851), .ZN(n16450) );
NAND2_X2 U12361 ( .A1(n17892), .A2(n17882), .ZN(n16537) );
NAND2_X2 U12365 ( .A1(n17906), .A2(n17735), .ZN(n16532) );
NAND2_X2 U12366 ( .A1(n17999), .A2(enc_byte_cnt[5]), .ZN(n16531) );
XNOR2_X2 U12368 ( .A(n17264), .B(n16545), .ZN(n16544) );
NAND2_X2 U12370 ( .A1(n17929), .A2(n16548), .ZN(n13317) );
XNOR2_X2 U12371 ( .A(n19191), .B(aes_text_out[7]), .ZN(n16548) );
XNOR2_X2 U12375 ( .A(n17266), .B(n16550), .ZN(n16549) );
NAND2_X2 U12377 ( .A1(n17930), .A2(n16553), .ZN(n13312) );
XNOR2_X2 U12378 ( .A(n19192), .B(aes_text_out[6]), .ZN(n16553) );
XNOR2_X2 U12382 ( .A(n17268), .B(n16555), .ZN(n16554) );
NAND2_X2 U12384 ( .A1(n17929), .A2(n16558), .ZN(n13307) );
XNOR2_X2 U12385 ( .A(n19193), .B(aes_text_out[5]), .ZN(n16558) );
XNOR2_X2 U12389 ( .A(n17270), .B(n16560), .ZN(n16559) );
NAND2_X2 U12391 ( .A1(n17930), .A2(n16563), .ZN(n13302) );
XNOR2_X2 U12392 ( .A(n19194), .B(aes_text_out[4]), .ZN(n16563) );
XNOR2_X2 U12396 ( .A(n17272), .B(n16565), .ZN(n16564) );
NAND2_X2 U12398 ( .A1(n17930), .A2(n16568), .ZN(n13297) );
XNOR2_X2 U12399 ( .A(n19195), .B(aes_text_out[3]), .ZN(n16568) );
XNOR2_X2 U12403 ( .A(n17274), .B(n16570), .ZN(n16569) );
NAND2_X2 U12406 ( .A1(n17930), .A2(n16572), .ZN(n13292) );
XNOR2_X2 U12407 ( .A(n19196), .B(aes_text_out[2]), .ZN(n16572) );
XNOR2_X2 U12409 ( .A(n17276), .B(n16574), .ZN(n16573) );
NAND2_X2 U12412 ( .A1(n17929), .A2(n16576), .ZN(n13287) );
XNOR2_X2 U12413 ( .A(n19197), .B(aes_text_out[1]), .ZN(n16576) );
XNOR2_X2 U12415 ( .A(n17278), .B(n16578), .ZN(n16577) );
NAND2_X2 U12419 ( .A1(n17930), .A2(n16580), .ZN(n13280) );
XNOR2_X2 U12420 ( .A(n19198), .B(aes_text_out[0]), .ZN(n16580) );
AND2_X2 U12424 ( .A1(n18056), .A2(z_out[127]), .ZN(N3070) );
AND2_X2 U12425 ( .A1(n18056), .A2(z_out[126]), .ZN(N3069) );
AND2_X2 U12426 ( .A1(n18056), .A2(z_out[125]), .ZN(N3068) );
AND2_X2 U12427 ( .A1(n18056), .A2(z_out[124]), .ZN(N3067) );
AND2_X2 U12428 ( .A1(n18056), .A2(z_out[123]), .ZN(N3066) );
AND2_X2 U12429 ( .A1(n18056), .A2(z_out[122]), .ZN(N3065) );
AND2_X2 U12430 ( .A1(n18056), .A2(z_out[121]), .ZN(N3064) );
AND2_X2 U12431 ( .A1(n18056), .A2(z_out[120]), .ZN(N3063) );
AND2_X2 U12432 ( .A1(n18056), .A2(z_out[119]), .ZN(N3062) );
AND2_X2 U12433 ( .A1(n18056), .A2(z_out[118]), .ZN(N3061) );
AND2_X2 U12434 ( .A1(n18056), .A2(z_out[117]), .ZN(N3060) );
AND2_X2 U12435 ( .A1(n18056), .A2(z_out[116]), .ZN(N3059) );
AND2_X2 U12436 ( .A1(n18056), .A2(z_out[115]), .ZN(N3058) );
AND2_X2 U12437 ( .A1(n18056), .A2(z_out[114]), .ZN(N3057) );
AND2_X2 U12438 ( .A1(n18056), .A2(z_out[113]), .ZN(N3056) );
AND2_X2 U12439 ( .A1(n18055), .A2(z_out[112]), .ZN(N3055) );
AND2_X2 U12440 ( .A1(n18055), .A2(z_out[111]), .ZN(N3054) );
AND2_X2 U12441 ( .A1(n18055), .A2(z_out[110]), .ZN(N3053) );
AND2_X2 U12442 ( .A1(n18055), .A2(z_out[109]), .ZN(N3052) );
AND2_X2 U12443 ( .A1(n18055), .A2(z_out[108]), .ZN(N3051) );
AND2_X2 U12444 ( .A1(n18055), .A2(z_out[107]), .ZN(N3050) );
AND2_X2 U12445 ( .A1(n18055), .A2(z_out[106]), .ZN(N3049) );
AND2_X2 U12446 ( .A1(n18055), .A2(z_out[105]), .ZN(N3048) );
AND2_X2 U12447 ( .A1(n18055), .A2(z_out[104]), .ZN(N3047) );
AND2_X2 U12448 ( .A1(n18055), .A2(z_out[103]), .ZN(N3046) );
AND2_X2 U12449 ( .A1(n18055), .A2(z_out[102]), .ZN(N3045) );
AND2_X2 U12450 ( .A1(n18055), .A2(z_out[101]), .ZN(N3044) );
AND2_X2 U12451 ( .A1(n18055), .A2(z_out[100]), .ZN(N3043) );
AND2_X2 U12452 ( .A1(n18055), .A2(z_out[99]), .ZN(N3042) );
AND2_X2 U12453 ( .A1(n18055), .A2(z_out[98]), .ZN(N3041) );
AND2_X2 U12454 ( .A1(n18055), .A2(z_out[97]), .ZN(N3040) );
AND2_X2 U12455 ( .A1(n18055), .A2(z_out[96]), .ZN(N3039) );
AND2_X2 U12456 ( .A1(n18055), .A2(z_out[95]), .ZN(N3038) );
AND2_X2 U12457 ( .A1(n18055), .A2(z_out[94]), .ZN(N3037) );
AND2_X2 U12458 ( .A1(n18055), .A2(z_out[93]), .ZN(N3036) );
AND2_X2 U12459 ( .A1(n18055), .A2(z_out[92]), .ZN(N3035) );
AND2_X2 U12460 ( .A1(n18055), .A2(z_out[91]), .ZN(N3034) );
AND2_X2 U12461 ( .A1(n18055), .A2(z_out[90]), .ZN(N3033) );
AND2_X2 U12462 ( .A1(n18054), .A2(z_out[89]), .ZN(N3032) );
AND2_X2 U12463 ( .A1(n18054), .A2(z_out[88]), .ZN(N3031) );
AND2_X2 U12464 ( .A1(n18054), .A2(z_out[87]), .ZN(N3030) );
AND2_X2 U12465 ( .A1(n18054), .A2(z_out[86]), .ZN(N3029) );
AND2_X2 U12466 ( .A1(n18054), .A2(z_out[85]), .ZN(N3028) );
AND2_X2 U12467 ( .A1(n18054), .A2(z_out[84]), .ZN(N3027) );
AND2_X2 U12468 ( .A1(n18054), .A2(z_out[83]), .ZN(N3026) );
AND2_X2 U12469 ( .A1(n18054), .A2(z_out[82]), .ZN(N3025) );
AND2_X2 U12470 ( .A1(n18054), .A2(z_out[81]), .ZN(N3024) );
AND2_X2 U12471 ( .A1(n18054), .A2(z_out[80]), .ZN(N3023) );
AND2_X2 U12472 ( .A1(n18054), .A2(z_out[79]), .ZN(N3022) );
AND2_X2 U12473 ( .A1(n18054), .A2(z_out[78]), .ZN(N3021) );
AND2_X2 U12474 ( .A1(n18054), .A2(z_out[77]), .ZN(N3020) );
AND2_X2 U12475 ( .A1(n18054), .A2(z_out[76]), .ZN(N3019) );
AND2_X2 U12476 ( .A1(n18054), .A2(z_out[75]), .ZN(N3018) );
AND2_X2 U12477 ( .A1(n18054), .A2(z_out[74]), .ZN(N3017) );
AND2_X2 U12478 ( .A1(n18054), .A2(z_out[73]), .ZN(N3016) );
AND2_X2 U12479 ( .A1(n18054), .A2(z_out[72]), .ZN(N3015) );
AND2_X2 U12480 ( .A1(n18054), .A2(z_out[71]), .ZN(N3014) );
AND2_X2 U12481 ( .A1(n18054), .A2(z_out[70]), .ZN(N3013) );
AND2_X2 U12482 ( .A1(n18054), .A2(z_out[69]), .ZN(N3012) );
AND2_X2 U12483 ( .A1(n18054), .A2(z_out[68]), .ZN(N3011) );
AND2_X2 U12484 ( .A1(n18054), .A2(z_out[67]), .ZN(N3010) );
AND2_X2 U12485 ( .A1(n18053), .A2(z_out[66]), .ZN(N3009) );
AND2_X2 U12486 ( .A1(n18053), .A2(z_out[65]), .ZN(N3008) );
AND2_X2 U12487 ( .A1(n18051), .A2(z_out[64]), .ZN(N3007) );
AND2_X2 U12488 ( .A1(n18053), .A2(z_out[63]), .ZN(N3006) );
AND2_X2 U12489 ( .A1(n18053), .A2(z_out[62]), .ZN(N3005) );
AND2_X2 U12490 ( .A1(n18053), .A2(z_out[61]), .ZN(N3004) );
AND2_X2 U12491 ( .A1(n18053), .A2(z_out[60]), .ZN(N3003) );
AND2_X2 U12492 ( .A1(n18053), .A2(z_out[59]), .ZN(N3002) );
AND2_X2 U12493 ( .A1(n18053), .A2(z_out[58]), .ZN(N3001) );
AND2_X2 U12494 ( .A1(n18053), .A2(z_out[57]), .ZN(N3000) );
AND2_X2 U12495 ( .A1(n18053), .A2(z_out[56]), .ZN(N2999) );
AND2_X2 U12496 ( .A1(n18053), .A2(z_out[55]), .ZN(N2998) );
AND2_X2 U12497 ( .A1(n18053), .A2(z_out[54]), .ZN(N2997) );
AND2_X2 U12498 ( .A1(n18053), .A2(z_out[53]), .ZN(N2996) );
AND2_X2 U12499 ( .A1(n18053), .A2(z_out[52]), .ZN(N2995) );
AND2_X2 U12500 ( .A1(n18053), .A2(z_out[51]), .ZN(N2994) );
AND2_X2 U12501 ( .A1(n18053), .A2(z_out[50]), .ZN(N2993) );
AND2_X2 U12502 ( .A1(n18053), .A2(z_out[49]), .ZN(N2992) );
AND2_X2 U12503 ( .A1(n18053), .A2(z_out[48]), .ZN(N2991) );
AND2_X2 U12504 ( .A1(n18053), .A2(z_out[47]), .ZN(N2990) );
AND2_X2 U12505 ( .A1(n18053), .A2(z_out[46]), .ZN(N2989) );
AND2_X2 U12506 ( .A1(n18053), .A2(z_out[45]), .ZN(N2988) );
AND2_X2 U12507 ( .A1(n18053), .A2(z_out[44]), .ZN(N2987) );
AND2_X2 U12508 ( .A1(n18052), .A2(z_out[43]), .ZN(N2986) );
AND2_X2 U12509 ( .A1(n18052), .A2(z_out[42]), .ZN(N2985) );
AND2_X2 U12510 ( .A1(n18052), .A2(z_out[41]), .ZN(N2984) );
AND2_X2 U12511 ( .A1(n18052), .A2(z_out[40]), .ZN(N2983) );
AND2_X2 U12512 ( .A1(n18052), .A2(z_out[39]), .ZN(N2982) );
AND2_X2 U12513 ( .A1(n18052), .A2(z_out[38]), .ZN(N2981) );
AND2_X2 U12514 ( .A1(n18052), .A2(z_out[37]), .ZN(N2980) );
AND2_X2 U12515 ( .A1(n18052), .A2(z_out[36]), .ZN(N2979) );
AND2_X2 U12516 ( .A1(n18052), .A2(z_out[35]), .ZN(N2978) );
AND2_X2 U12517 ( .A1(n18052), .A2(z_out[34]), .ZN(N2977) );
AND2_X2 U12518 ( .A1(n18052), .A2(z_out[33]), .ZN(N2976) );
AND2_X2 U12519 ( .A1(n18052), .A2(z_out[32]), .ZN(N2975) );
AND2_X2 U12520 ( .A1(n18052), .A2(z_out[31]), .ZN(N2974) );
AND2_X2 U12521 ( .A1(n18052), .A2(z_out[30]), .ZN(N2973) );
AND2_X2 U12522 ( .A1(n18052), .A2(z_out[29]), .ZN(N2972) );
AND2_X2 U12523 ( .A1(n18052), .A2(z_out[28]), .ZN(N2971) );
AND2_X2 U12524 ( .A1(n18052), .A2(z_out[27]), .ZN(N2970) );
AND2_X2 U12525 ( .A1(n18052), .A2(z_out[26]), .ZN(N2969) );
AND2_X2 U12526 ( .A1(n18052), .A2(z_out[25]), .ZN(N2968) );
AND2_X2 U12527 ( .A1(n18052), .A2(z_out[24]), .ZN(N2967) );
AND2_X2 U12528 ( .A1(n18052), .A2(z_out[23]), .ZN(N2966) );
AND2_X2 U12529 ( .A1(n18052), .A2(z_out[22]), .ZN(N2965) );
AND2_X2 U12530 ( .A1(n18052), .A2(z_out[21]), .ZN(N2964) );
AND2_X2 U12531 ( .A1(n18051), .A2(z_out[20]), .ZN(N2963) );
AND2_X2 U12532 ( .A1(n18051), .A2(z_out[19]), .ZN(N2962) );
AND2_X2 U12533 ( .A1(n18051), .A2(z_out[18]), .ZN(N2961) );
AND2_X2 U12534 ( .A1(n18051), .A2(z_out[17]), .ZN(N2960) );
AND2_X2 U12535 ( .A1(n18051), .A2(z_out[16]), .ZN(N2959) );
AND2_X2 U12536 ( .A1(n18051), .A2(z_out[15]), .ZN(N2958) );
AND2_X2 U12537 ( .A1(n18051), .A2(z_out[14]), .ZN(N2957) );
AND2_X2 U12538 ( .A1(n18051), .A2(z_out[13]), .ZN(N2956) );
AND2_X2 U12539 ( .A1(n18051), .A2(z_out[12]), .ZN(N2955) );
AND2_X2 U12540 ( .A1(n18051), .A2(z_out[11]), .ZN(N2954) );
AND2_X2 U12541 ( .A1(n18051), .A2(z_out[10]), .ZN(N2953) );
AND2_X2 U12542 ( .A1(n18051), .A2(z_out[9]), .ZN(N2952) );
AND2_X2 U12543 ( .A1(n18051), .A2(z_out[8]), .ZN(N2951) );
AND2_X2 U12544 ( .A1(n18051), .A2(z_out[7]), .ZN(N2950) );
AND2_X2 U12545 ( .A1(n18051), .A2(z_out[6]), .ZN(N2949) );
AND2_X2 U12546 ( .A1(n18051), .A2(z_out[5]), .ZN(N2948) );
AND2_X2 U12547 ( .A1(n18051), .A2(z_out[4]), .ZN(N2947) );
AND2_X2 U12548 ( .A1(n18051), .A2(z_out[3]), .ZN(N2946) );
AND2_X2 U12549 ( .A1(n18053), .A2(z_out[2]), .ZN(N2945) );
AND2_X2 U12550 ( .A1(n18051), .A2(z_out[1]), .ZN(N2944) );
AND2_X2 U12551 ( .A1(n18056), .A2(z_out[0]), .ZN(N2943) );
NAND2_X2 U12552 ( .A1(n16581), .A2(n16582), .ZN(N2942) );
NAND2_X2 U12553 ( .A1(v_out[127]), .A2(n18047), .ZN(n16582) );
NAND2_X2 U12554 ( .A1(n18059), .A2(n17292), .ZN(n16581) );
NAND2_X2 U12555 ( .A1(n16583), .A2(n16584), .ZN(N2941) );
NAND2_X2 U12556 ( .A1(v_out[126]), .A2(n18044), .ZN(n16584) );
NAND2_X2 U12557 ( .A1(n18059), .A2(n17293), .ZN(n16583) );
NAND2_X2 U12558 ( .A1(n16585), .A2(n16586), .ZN(N2940) );
NAND2_X2 U12559 ( .A1(v_out[125]), .A2(n18044), .ZN(n16586) );
NAND2_X2 U12560 ( .A1(n18059), .A2(n17294), .ZN(n16585) );
NAND2_X2 U12561 ( .A1(n16587), .A2(n16588), .ZN(N2939) );
NAND2_X2 U12562 ( .A1(v_out[124]), .A2(n18044), .ZN(n16588) );
NAND2_X2 U12563 ( .A1(n18059), .A2(n17295), .ZN(n16587) );
NAND2_X2 U12564 ( .A1(n16589), .A2(n16590), .ZN(N2938) );
NAND2_X2 U12565 ( .A1(v_out[123]), .A2(n18044), .ZN(n16590) );
NAND2_X2 U12566 ( .A1(n18059), .A2(n17296), .ZN(n16589) );
NAND2_X2 U12567 ( .A1(n16591), .A2(n16592), .ZN(N2937) );
NAND2_X2 U12568 ( .A1(v_out[122]), .A2(n18044), .ZN(n16592) );
NAND2_X2 U12569 ( .A1(n18059), .A2(n17297), .ZN(n16591) );
NAND2_X2 U12570 ( .A1(n16593), .A2(n16594), .ZN(N2936) );
NAND2_X2 U12571 ( .A1(v_out[121]), .A2(n18044), .ZN(n16594) );
NAND2_X2 U12572 ( .A1(n18059), .A2(n17298), .ZN(n16593) );
NAND2_X2 U12573 ( .A1(n16595), .A2(n16596), .ZN(N2935) );
NAND2_X2 U12574 ( .A1(v_out[120]), .A2(n18044), .ZN(n16596) );
NAND2_X2 U12575 ( .A1(n18059), .A2(n17299), .ZN(n16595) );
NAND2_X2 U12576 ( .A1(n16597), .A2(n16598), .ZN(N2934) );
NAND2_X2 U12577 ( .A1(v_out[119]), .A2(n18044), .ZN(n16598) );
NAND2_X2 U12578 ( .A1(n18059), .A2(n17300), .ZN(n16597) );
NAND2_X2 U12579 ( .A1(n16599), .A2(n16600), .ZN(N2933) );
NAND2_X2 U12580 ( .A1(v_out[118]), .A2(n18044), .ZN(n16600) );
NAND2_X2 U12581 ( .A1(n18059), .A2(n17301), .ZN(n16599) );
NAND2_X2 U12582 ( .A1(n16601), .A2(n16602), .ZN(N2932) );
NAND2_X2 U12583 ( .A1(v_out[117]), .A2(n18044), .ZN(n16602) );
NAND2_X2 U12584 ( .A1(n18059), .A2(n17302), .ZN(n16601) );
NAND2_X2 U12585 ( .A1(n16603), .A2(n16604), .ZN(N2931) );
NAND2_X2 U12586 ( .A1(v_out[116]), .A2(n18044), .ZN(n16604) );
NAND2_X2 U12587 ( .A1(n18059), .A2(n17303), .ZN(n16603) );
NAND2_X2 U12588 ( .A1(n16605), .A2(n16606), .ZN(N2930) );
NAND2_X2 U12589 ( .A1(v_out[115]), .A2(n18044), .ZN(n16606) );
NAND2_X2 U12590 ( .A1(n18059), .A2(n17304), .ZN(n16605) );
NAND2_X2 U12591 ( .A1(n16607), .A2(n16608), .ZN(N2929) );
NAND2_X2 U12592 ( .A1(v_out[114]), .A2(n18044), .ZN(n16608) );
NAND2_X2 U12593 ( .A1(n18059), .A2(n17305), .ZN(n16607) );
NAND2_X2 U12594 ( .A1(n16609), .A2(n16610), .ZN(N2928) );
NAND2_X2 U12595 ( .A1(v_out[113]), .A2(n18044), .ZN(n16610) );
NAND2_X2 U12596 ( .A1(n18060), .A2(n17306), .ZN(n16609) );
NAND2_X2 U12597 ( .A1(n16611), .A2(n16612), .ZN(N2927) );
NAND2_X2 U12598 ( .A1(v_out[112]), .A2(n18044), .ZN(n16612) );
NAND2_X2 U12599 ( .A1(n18059), .A2(n17307), .ZN(n16611) );
NAND2_X2 U12600 ( .A1(n16613), .A2(n16614), .ZN(N2926) );
NAND2_X2 U12601 ( .A1(v_out[111]), .A2(n18044), .ZN(n16614) );
NAND2_X2 U12602 ( .A1(n18059), .A2(n17308), .ZN(n16613) );
NAND2_X2 U12603 ( .A1(n16615), .A2(n16616), .ZN(N2925) );
NAND2_X2 U12604 ( .A1(v_out[110]), .A2(n18044), .ZN(n16616) );
NAND2_X2 U12605 ( .A1(n18059), .A2(n17309), .ZN(n16615) );
NAND2_X2 U12606 ( .A1(n16617), .A2(n16618), .ZN(N2924) );
NAND2_X2 U12607 ( .A1(v_out[109]), .A2(n18045), .ZN(n16618) );
NAND2_X2 U12608 ( .A1(n18059), .A2(n17310), .ZN(n16617) );
NAND2_X2 U12609 ( .A1(n16619), .A2(n16620), .ZN(N2923) );
NAND2_X2 U12610 ( .A1(v_out[108]), .A2(n18045), .ZN(n16620) );
NAND2_X2 U12611 ( .A1(n18060), .A2(n17311), .ZN(n16619) );
NAND2_X2 U12612 ( .A1(n16621), .A2(n16622), .ZN(N2922) );
NAND2_X2 U12613 ( .A1(v_out[107]), .A2(n18045), .ZN(n16622) );
NAND2_X2 U12614 ( .A1(n18060), .A2(n17312), .ZN(n16621) );
NAND2_X2 U12615 ( .A1(n16623), .A2(n16624), .ZN(N2921) );
NAND2_X2 U12616 ( .A1(v_out[106]), .A2(n18045), .ZN(n16624) );
NAND2_X2 U12617 ( .A1(n18060), .A2(n17313), .ZN(n16623) );
NAND2_X2 U12618 ( .A1(n16625), .A2(n16626), .ZN(N2920) );
NAND2_X2 U12619 ( .A1(v_out[105]), .A2(n18045), .ZN(n16626) );
NAND2_X2 U12620 ( .A1(n18060), .A2(n17314), .ZN(n16625) );
NAND2_X2 U12621 ( .A1(n16627), .A2(n16628), .ZN(N2919) );
NAND2_X2 U12622 ( .A1(v_out[104]), .A2(n18045), .ZN(n16628) );
NAND2_X2 U12623 ( .A1(n18060), .A2(n17315), .ZN(n16627) );
NAND2_X2 U12624 ( .A1(n16629), .A2(n16630), .ZN(N2918) );
NAND2_X2 U12625 ( .A1(v_out[103]), .A2(n18045), .ZN(n16630) );
NAND2_X2 U12626 ( .A1(n18060), .A2(n17316), .ZN(n16629) );
NAND2_X2 U12627 ( .A1(n16631), .A2(n16632), .ZN(N2917) );
NAND2_X2 U12628 ( .A1(v_out[102]), .A2(n18045), .ZN(n16632) );
NAND2_X2 U12629 ( .A1(n18060), .A2(n17317), .ZN(n16631) );
NAND2_X2 U12630 ( .A1(n16633), .A2(n16634), .ZN(N2916) );
NAND2_X2 U12631 ( .A1(v_out[101]), .A2(n18045), .ZN(n16634) );
NAND2_X2 U12632 ( .A1(n18060), .A2(n17318), .ZN(n16633) );
NAND2_X2 U12633 ( .A1(n16635), .A2(n16636), .ZN(N2915) );
NAND2_X2 U12634 ( .A1(v_out[100]), .A2(n18045), .ZN(n16636) );
NAND2_X2 U12635 ( .A1(n18060), .A2(n17319), .ZN(n16635) );
NAND2_X2 U12636 ( .A1(n16637), .A2(n16638), .ZN(N2914) );
NAND2_X2 U12637 ( .A1(v_out[99]), .A2(n18045), .ZN(n16638) );
NAND2_X2 U12638 ( .A1(n18060), .A2(n17320), .ZN(n16637) );
NAND2_X2 U12639 ( .A1(n16639), .A2(n16640), .ZN(N2913) );
NAND2_X2 U12640 ( .A1(v_out[98]), .A2(n18045), .ZN(n16640) );
NAND2_X2 U12641 ( .A1(n18060), .A2(n17321), .ZN(n16639) );
NAND2_X2 U12642 ( .A1(n16641), .A2(n16642), .ZN(N2912) );
NAND2_X2 U12643 ( .A1(v_out[97]), .A2(n18045), .ZN(n16642) );
NAND2_X2 U12644 ( .A1(n18060), .A2(n17322), .ZN(n16641) );
NAND2_X2 U12645 ( .A1(n16643), .A2(n16644), .ZN(N2911) );
NAND2_X2 U12646 ( .A1(v_out[96]), .A2(n18045), .ZN(n16644) );
NAND2_X2 U12647 ( .A1(n18060), .A2(n17323), .ZN(n16643) );
NAND2_X2 U12648 ( .A1(n16645), .A2(n16646), .ZN(N2910) );
NAND2_X2 U12649 ( .A1(v_out[95]), .A2(n18045), .ZN(n16646) );
NAND2_X2 U12650 ( .A1(n18060), .A2(n17324), .ZN(n16645) );
NAND2_X2 U12651 ( .A1(n16647), .A2(n16648), .ZN(N2909) );
NAND2_X2 U12652 ( .A1(v_out[94]), .A2(n18045), .ZN(n16648) );
NAND2_X2 U12653 ( .A1(n18060), .A2(n17325), .ZN(n16647) );
NAND2_X2 U12654 ( .A1(n16649), .A2(n16650), .ZN(N2908) );
NAND2_X2 U12655 ( .A1(v_out[93]), .A2(n18045), .ZN(n16650) );
NAND2_X2 U12656 ( .A1(n18060), .A2(n17326), .ZN(n16649) );
NAND2_X2 U12657 ( .A1(n16651), .A2(n16652), .ZN(N2907) );
NAND2_X2 U12658 ( .A1(v_out[92]), .A2(n18045), .ZN(n16652) );
NAND2_X2 U12659 ( .A1(n18058), .A2(n17327), .ZN(n16651) );
NAND2_X2 U12660 ( .A1(n16653), .A2(n16654), .ZN(N2906) );
NAND2_X2 U12661 ( .A1(v_out[91]), .A2(n18046), .ZN(n16654) );
NAND2_X2 U12662 ( .A1(n18060), .A2(n17328), .ZN(n16653) );
NAND2_X2 U12663 ( .A1(n16655), .A2(n16656), .ZN(N2905) );
NAND2_X2 U12664 ( .A1(v_out[90]), .A2(n18046), .ZN(n16656) );
NAND2_X2 U12665 ( .A1(n18060), .A2(n17329), .ZN(n16655) );
NAND2_X2 U12666 ( .A1(n16657), .A2(n16658), .ZN(N2904) );
NAND2_X2 U12667 ( .A1(v_out[89]), .A2(n18046), .ZN(n16658) );
NAND2_X2 U12668 ( .A1(n18060), .A2(n17330), .ZN(n16657) );
NAND2_X2 U12669 ( .A1(n16659), .A2(n16660), .ZN(N2903) );
NAND2_X2 U12670 ( .A1(v_out[88]), .A2(n18046), .ZN(n16660) );
NAND2_X2 U12671 ( .A1(n18060), .A2(n17331), .ZN(n16659) );
NAND2_X2 U12672 ( .A1(n16661), .A2(n16662), .ZN(N2902) );
NAND2_X2 U12673 ( .A1(v_out[87]), .A2(n18046), .ZN(n16662) );
NAND2_X2 U12674 ( .A1(n18058), .A2(n17332), .ZN(n16661) );
NAND2_X2 U12675 ( .A1(n16663), .A2(n16664), .ZN(N2901) );
NAND2_X2 U12676 ( .A1(v_out[86]), .A2(n18046), .ZN(n16664) );
NAND2_X2 U12677 ( .A1(n18057), .A2(n17333), .ZN(n16663) );
NAND2_X2 U12678 ( .A1(n16665), .A2(n16666), .ZN(N2900) );
NAND2_X2 U12679 ( .A1(v_out[85]), .A2(n18046), .ZN(n16666) );
NAND2_X2 U12680 ( .A1(n18064), .A2(n17334), .ZN(n16665) );
NAND2_X2 U12681 ( .A1(n16667), .A2(n16668), .ZN(N2899) );
NAND2_X2 U12682 ( .A1(v_out[84]), .A2(n18046), .ZN(n16668) );
NAND2_X2 U12683 ( .A1(n18066), .A2(n17335), .ZN(n16667) );
NAND2_X2 U12684 ( .A1(n16669), .A2(n16670), .ZN(N2898) );
NAND2_X2 U12685 ( .A1(v_out[83]), .A2(n18046), .ZN(n16670) );
NAND2_X2 U12686 ( .A1(n18068), .A2(n17336), .ZN(n16669) );
NAND2_X2 U12687 ( .A1(n16671), .A2(n16672), .ZN(N2897) );
NAND2_X2 U12688 ( .A1(v_out[82]), .A2(n18046), .ZN(n16672) );
NAND2_X2 U12689 ( .A1(n18067), .A2(n17337), .ZN(n16671) );
NAND2_X2 U12690 ( .A1(n16673), .A2(n16674), .ZN(N2896) );
NAND2_X2 U12691 ( .A1(v_out[81]), .A2(n18046), .ZN(n16674) );
NAND2_X2 U12692 ( .A1(n18065), .A2(n17338), .ZN(n16673) );
NAND2_X2 U12693 ( .A1(n16675), .A2(n16676), .ZN(N2895) );
NAND2_X2 U12694 ( .A1(v_out[80]), .A2(n18046), .ZN(n16676) );
NAND2_X2 U12695 ( .A1(n18069), .A2(n17339), .ZN(n16675) );
NAND2_X2 U12696 ( .A1(n16677), .A2(n16678), .ZN(N2894) );
NAND2_X2 U12697 ( .A1(v_out[79]), .A2(n18046), .ZN(n16678) );
NAND2_X2 U12698 ( .A1(n18057), .A2(n17340), .ZN(n16677) );
NAND2_X2 U12699 ( .A1(n16679), .A2(n16680), .ZN(N2893) );
NAND2_X2 U12700 ( .A1(v_out[78]), .A2(n18046), .ZN(n16680) );
NAND2_X2 U12701 ( .A1(n18064), .A2(n17341), .ZN(n16679) );
NAND2_X2 U12702 ( .A1(n16681), .A2(n16682), .ZN(N2892) );
NAND2_X2 U12703 ( .A1(v_out[77]), .A2(n18046), .ZN(n16682) );
NAND2_X2 U12704 ( .A1(n18066), .A2(n17342), .ZN(n16681) );
NAND2_X2 U12705 ( .A1(n16683), .A2(n16684), .ZN(N2891) );
NAND2_X2 U12706 ( .A1(v_out[76]), .A2(n18046), .ZN(n16684) );
NAND2_X2 U12707 ( .A1(n18068), .A2(n17343), .ZN(n16683) );
NAND2_X2 U12708 ( .A1(n16685), .A2(n16686), .ZN(N2890) );
NAND2_X2 U12709 ( .A1(v_out[75]), .A2(n18046), .ZN(n16686) );
NAND2_X2 U12710 ( .A1(n18067), .A2(n17344), .ZN(n16685) );
NAND2_X2 U12711 ( .A1(n16687), .A2(n16688), .ZN(N2889) );
NAND2_X2 U12712 ( .A1(v_out[74]), .A2(n18046), .ZN(n16688) );
NAND2_X2 U12713 ( .A1(n18065), .A2(n17345), .ZN(n16687) );
NAND2_X2 U12714 ( .A1(n16689), .A2(n16690), .ZN(N2888) );
NAND2_X2 U12715 ( .A1(v_out[73]), .A2(n18047), .ZN(n16690) );
NAND2_X2 U12716 ( .A1(n18069), .A2(n17346), .ZN(n16689) );
NAND2_X2 U12717 ( .A1(n16691), .A2(n16692), .ZN(N2887) );
NAND2_X2 U12718 ( .A1(v_out[72]), .A2(n18047), .ZN(n16692) );
NAND2_X2 U12719 ( .A1(n18069), .A2(n17347), .ZN(n16691) );
NAND2_X2 U12720 ( .A1(n16693), .A2(n16694), .ZN(N2886) );
NAND2_X2 U12721 ( .A1(v_out[71]), .A2(n18047), .ZN(n16694) );
NAND2_X2 U12722 ( .A1(n18069), .A2(n17348), .ZN(n16693) );
NAND2_X2 U12723 ( .A1(n16695), .A2(n16696), .ZN(N2885) );
NAND2_X2 U12724 ( .A1(v_out[70]), .A2(n18047), .ZN(n16696) );
NAND2_X2 U12725 ( .A1(n18069), .A2(n17349), .ZN(n16695) );
NAND2_X2 U12726 ( .A1(n16697), .A2(n16698), .ZN(N2884) );
NAND2_X2 U12727 ( .A1(v_out[69]), .A2(n18047), .ZN(n16698) );
NAND2_X2 U12728 ( .A1(n18069), .A2(n17350), .ZN(n16697) );
NAND2_X2 U12729 ( .A1(n16699), .A2(n16700), .ZN(N2883) );
NAND2_X2 U12730 ( .A1(v_out[68]), .A2(n18047), .ZN(n16700) );
NAND2_X2 U12731 ( .A1(n18069), .A2(n17351), .ZN(n16699) );
NAND2_X2 U12732 ( .A1(n16701), .A2(n16702), .ZN(N2882) );
NAND2_X2 U12733 ( .A1(v_out[67]), .A2(n18047), .ZN(n16702) );
NAND2_X2 U12734 ( .A1(n18061), .A2(n17352), .ZN(n16701) );
NAND2_X2 U12735 ( .A1(n16703), .A2(n16704), .ZN(N2881) );
NAND2_X2 U12736 ( .A1(v_out[66]), .A2(n18047), .ZN(n16704) );
NAND2_X2 U12737 ( .A1(n18061), .A2(n17353), .ZN(n16703) );
NAND2_X2 U12738 ( .A1(n16705), .A2(n16706), .ZN(N2880) );
NAND2_X2 U12739 ( .A1(v_out[65]), .A2(n18047), .ZN(n16706) );
NAND2_X2 U12740 ( .A1(n18061), .A2(n17354), .ZN(n16705) );
NAND2_X2 U12741 ( .A1(n16707), .A2(n16708), .ZN(N2879) );
NAND2_X2 U12742 ( .A1(v_out[64]), .A2(n18047), .ZN(n16708) );
NAND2_X2 U12743 ( .A1(n18064), .A2(n17355), .ZN(n16707) );
NAND2_X2 U12744 ( .A1(n16709), .A2(n16710), .ZN(N2878) );
NAND2_X2 U12745 ( .A1(v_out[63]), .A2(n18047), .ZN(n16710) );
NAND2_X2 U12746 ( .A1(n18064), .A2(n17356), .ZN(n16709) );
NAND2_X2 U12747 ( .A1(n16711), .A2(n16712), .ZN(N2877) );
NAND2_X2 U12748 ( .A1(v_out[62]), .A2(n18047), .ZN(n16712) );
NAND2_X2 U12749 ( .A1(n18064), .A2(n17357), .ZN(n16711) );
NAND2_X2 U12750 ( .A1(n16713), .A2(n16714), .ZN(N2876) );
NAND2_X2 U12751 ( .A1(v_out[61]), .A2(n18047), .ZN(n16714) );
NAND2_X2 U12752 ( .A1(n18064), .A2(n17358), .ZN(n16713) );
NAND2_X2 U12753 ( .A1(n16715), .A2(n16716), .ZN(N2875) );
NAND2_X2 U12754 ( .A1(v_out[60]), .A2(n18047), .ZN(n16716) );
NAND2_X2 U12755 ( .A1(n18063), .A2(n17359), .ZN(n16715) );
NAND2_X2 U12756 ( .A1(n16717), .A2(n16718), .ZN(N2874) );
NAND2_X2 U12757 ( .A1(v_out[59]), .A2(n18047), .ZN(n16718) );
NAND2_X2 U12758 ( .A1(n18063), .A2(n17360), .ZN(n16717) );
NAND2_X2 U12759 ( .A1(n16719), .A2(n16720), .ZN(N2873) );
NAND2_X2 U12760 ( .A1(v_out[58]), .A2(n18047), .ZN(n16720) );
NAND2_X2 U12761 ( .A1(n18063), .A2(n17361), .ZN(n16719) );
NAND2_X2 U12762 ( .A1(n16721), .A2(n16722), .ZN(N2872) );
NAND2_X2 U12763 ( .A1(v_out[57]), .A2(n18048), .ZN(n16722) );
NAND2_X2 U12764 ( .A1(n18063), .A2(n17362), .ZN(n16721) );
NAND2_X2 U12765 ( .A1(n16723), .A2(n16724), .ZN(N2871) );
NAND2_X2 U12766 ( .A1(v_out[56]), .A2(n18048), .ZN(n16724) );
NAND2_X2 U12767 ( .A1(n18063), .A2(n17363), .ZN(n16723) );
NAND2_X2 U12768 ( .A1(n16725), .A2(n16726), .ZN(N2870) );
NAND2_X2 U12769 ( .A1(v_out[55]), .A2(n18048), .ZN(n16726) );
NAND2_X2 U12770 ( .A1(n18063), .A2(n17364), .ZN(n16725) );
NAND2_X2 U12771 ( .A1(n16727), .A2(n16728), .ZN(N2869) );
NAND2_X2 U12772 ( .A1(v_out[54]), .A2(n18048), .ZN(n16728) );
NAND2_X2 U12773 ( .A1(n18063), .A2(n17365), .ZN(n16727) );
NAND2_X2 U12774 ( .A1(n16729), .A2(n16730), .ZN(N2868) );
NAND2_X2 U12775 ( .A1(v_out[53]), .A2(n18048), .ZN(n16730) );
NAND2_X2 U12776 ( .A1(n18063), .A2(n17366), .ZN(n16729) );
NAND2_X2 U12777 ( .A1(n16731), .A2(n16732), .ZN(N2867) );
NAND2_X2 U12778 ( .A1(v_out[52]), .A2(n18048), .ZN(n16732) );
NAND2_X2 U12779 ( .A1(n18063), .A2(n17367), .ZN(n16731) );
NAND2_X2 U12780 ( .A1(n16733), .A2(n16734), .ZN(N2866) );
NAND2_X2 U12781 ( .A1(v_out[51]), .A2(n18048), .ZN(n16734) );
NAND2_X2 U12782 ( .A1(n18063), .A2(n17368), .ZN(n16733) );
NAND2_X2 U12783 ( .A1(n16735), .A2(n16736), .ZN(N2865) );
NAND2_X2 U12784 ( .A1(v_out[50]), .A2(n18048), .ZN(n16736) );
NAND2_X2 U12785 ( .A1(n18063), .A2(n17369), .ZN(n16735) );
NAND2_X2 U12786 ( .A1(n16737), .A2(n16738), .ZN(N2864) );
NAND2_X2 U12787 ( .A1(v_out[49]), .A2(n18048), .ZN(n16738) );
NAND2_X2 U12788 ( .A1(n18063), .A2(n17370), .ZN(n16737) );
NAND2_X2 U12789 ( .A1(n16739), .A2(n16740), .ZN(N2863) );
NAND2_X2 U12790 ( .A1(v_out[48]), .A2(n18048), .ZN(n16740) );
NAND2_X2 U12791 ( .A1(n18063), .A2(n17371), .ZN(n16739) );
NAND2_X2 U12792 ( .A1(n16741), .A2(n16742), .ZN(N2862) );
NAND2_X2 U12793 ( .A1(v_out[47]), .A2(n18048), .ZN(n16742) );
NAND2_X2 U12794 ( .A1(n18063), .A2(n17372), .ZN(n16741) );
NAND2_X2 U12795 ( .A1(n16743), .A2(n16744), .ZN(N2861) );
NAND2_X2 U12796 ( .A1(v_out[46]), .A2(n18048), .ZN(n16744) );
NAND2_X2 U12797 ( .A1(n18063), .A2(n17373), .ZN(n16743) );
NAND2_X2 U12798 ( .A1(n16745), .A2(n16746), .ZN(N2860) );
NAND2_X2 U12799 ( .A1(v_out[45]), .A2(n18048), .ZN(n16746) );
NAND2_X2 U12800 ( .A1(n18063), .A2(n17374), .ZN(n16745) );
NAND2_X2 U12801 ( .A1(n16747), .A2(n16748), .ZN(N2859) );
NAND2_X2 U12802 ( .A1(v_out[44]), .A2(n18048), .ZN(n16748) );
NAND2_X2 U12803 ( .A1(n18063), .A2(n18847), .ZN(n16747) );
NAND2_X2 U12804 ( .A1(n16749), .A2(n16750), .ZN(N2858) );
NAND2_X2 U12805 ( .A1(v_out[43]), .A2(n18048), .ZN(n16750) );
NAND2_X2 U12806 ( .A1(n18062), .A2(n18848), .ZN(n16749) );
NAND2_X2 U12807 ( .A1(n16751), .A2(n16752), .ZN(N2857) );
NAND2_X2 U12808 ( .A1(v_out[42]), .A2(n18048), .ZN(n16752) );
NAND2_X2 U12809 ( .A1(n18063), .A2(n18849), .ZN(n16751) );
NAND2_X2 U12810 ( .A1(n16753), .A2(n16754), .ZN(N2856) );
NAND2_X2 U12811 ( .A1(v_out[41]), .A2(n18048), .ZN(n16754) );
NAND2_X2 U12812 ( .A1(n18063), .A2(n18850), .ZN(n16753) );
NAND2_X2 U12813 ( .A1(n16755), .A2(n16756), .ZN(N2855) );
NAND2_X2 U12814 ( .A1(v_out[40]), .A2(n18048), .ZN(n16756) );
NAND2_X2 U12815 ( .A1(n18063), .A2(n18851), .ZN(n16755) );
NAND2_X2 U12816 ( .A1(n16757), .A2(n16758), .ZN(N2854) );
NAND2_X2 U12817 ( .A1(v_out[39]), .A2(n18049), .ZN(n16758) );
NAND2_X2 U12818 ( .A1(n18063), .A2(n18852), .ZN(n16757) );
NAND2_X2 U12819 ( .A1(n16759), .A2(n16760), .ZN(N2853) );
NAND2_X2 U12820 ( .A1(v_out[38]), .A2(n18049), .ZN(n16760) );
NAND2_X2 U12821 ( .A1(n18062), .A2(n18853), .ZN(n16759) );
NAND2_X2 U12822 ( .A1(n16761), .A2(n16762), .ZN(N2852) );
NAND2_X2 U12823 ( .A1(v_out[37]), .A2(n18049), .ZN(n16762) );
NAND2_X2 U12824 ( .A1(n18062), .A2(n18854), .ZN(n16761) );
NAND2_X2 U12825 ( .A1(n16763), .A2(n16764), .ZN(N2851) );
NAND2_X2 U12826 ( .A1(v_out[36]), .A2(n18049), .ZN(n16764) );
NAND2_X2 U12827 ( .A1(n18062), .A2(n18855), .ZN(n16763) );
NAND2_X2 U12828 ( .A1(n16765), .A2(n16766), .ZN(N2850) );
NAND2_X2 U12829 ( .A1(v_out[35]), .A2(n18049), .ZN(n16766) );
NAND2_X2 U12830 ( .A1(n18062), .A2(n18856), .ZN(n16765) );
NAND2_X2 U12831 ( .A1(n16767), .A2(n16768), .ZN(N2849) );
NAND2_X2 U12832 ( .A1(v_out[34]), .A2(n18049), .ZN(n16768) );
NAND2_X2 U12833 ( .A1(n18062), .A2(n18857), .ZN(n16767) );
NAND2_X2 U12834 ( .A1(n16769), .A2(n16770), .ZN(N2848) );
NAND2_X2 U12835 ( .A1(v_out[33]), .A2(n18049), .ZN(n16770) );
NAND2_X2 U12836 ( .A1(n18062), .A2(n18858), .ZN(n16769) );
NAND2_X2 U12837 ( .A1(n16771), .A2(n16772), .ZN(N2847) );
NAND2_X2 U12838 ( .A1(v_out[32]), .A2(n18049), .ZN(n16772) );
NAND2_X2 U12839 ( .A1(n18062), .A2(n18859), .ZN(n16771) );
NAND2_X2 U12840 ( .A1(n16773), .A2(n16774), .ZN(N2846) );
NAND2_X2 U12841 ( .A1(v_out[31]), .A2(n18049), .ZN(n16774) );
NAND2_X2 U12842 ( .A1(n18062), .A2(n18860), .ZN(n16773) );
NAND2_X2 U12843 ( .A1(n16775), .A2(n16776), .ZN(N2845) );
NAND2_X2 U12844 ( .A1(v_out[30]), .A2(n18049), .ZN(n16776) );
NAND2_X2 U12845 ( .A1(n18062), .A2(n18861), .ZN(n16775) );
NAND2_X2 U12846 ( .A1(n16777), .A2(n16778), .ZN(N2844) );
NAND2_X2 U12847 ( .A1(v_out[29]), .A2(n18049), .ZN(n16778) );
NAND2_X2 U12848 ( .A1(n18062), .A2(n18862), .ZN(n16777) );
NAND2_X2 U12849 ( .A1(n16779), .A2(n16780), .ZN(N2843) );
NAND2_X2 U12850 ( .A1(v_out[28]), .A2(n18049), .ZN(n16780) );
NAND2_X2 U12851 ( .A1(n18062), .A2(n18863), .ZN(n16779) );
NAND2_X2 U12852 ( .A1(n16781), .A2(n16782), .ZN(N2842) );
NAND2_X2 U12853 ( .A1(v_out[27]), .A2(n18049), .ZN(n16782) );
NAND2_X2 U12854 ( .A1(n18062), .A2(n18864), .ZN(n16781) );
NAND2_X2 U12855 ( .A1(n16783), .A2(n16784), .ZN(N2841) );
NAND2_X2 U12856 ( .A1(v_out[26]), .A2(n18049), .ZN(n16784) );
NAND2_X2 U12857 ( .A1(n18062), .A2(n18865), .ZN(n16783) );
NAND2_X2 U12858 ( .A1(n16785), .A2(n16786), .ZN(N2840) );
NAND2_X2 U12859 ( .A1(v_out[25]), .A2(n18049), .ZN(n16786) );
NAND2_X2 U12860 ( .A1(n18062), .A2(n18866), .ZN(n16785) );
NAND2_X2 U12861 ( .A1(n16787), .A2(n16788), .ZN(N2839) );
NAND2_X2 U12862 ( .A1(v_out[24]), .A2(n18049), .ZN(n16788) );
NAND2_X2 U12863 ( .A1(n18062), .A2(n18867), .ZN(n16787) );
NAND2_X2 U12864 ( .A1(n16789), .A2(n16790), .ZN(N2838) );
NAND2_X2 U12865 ( .A1(v_out[23]), .A2(n18049), .ZN(n16790) );
NAND2_X2 U12866 ( .A1(n18062), .A2(n18868), .ZN(n16789) );
NAND2_X2 U12867 ( .A1(n16791), .A2(n16792), .ZN(N2837) );
NAND2_X2 U12868 ( .A1(v_out[22]), .A2(n18049), .ZN(n16792) );
NAND2_X2 U12869 ( .A1(n18062), .A2(n18869), .ZN(n16791) );
NAND2_X2 U12870 ( .A1(n16793), .A2(n16794), .ZN(N2836) );
NAND2_X2 U12871 ( .A1(v_out[21]), .A2(n18050), .ZN(n16794) );
NAND2_X2 U12872 ( .A1(n18062), .A2(n18870), .ZN(n16793) );
NAND2_X2 U12873 ( .A1(n16795), .A2(n16796), .ZN(N2835) );
NAND2_X2 U12874 ( .A1(v_out[20]), .A2(n18050), .ZN(n16796) );
NAND2_X2 U12875 ( .A1(n18062), .A2(n18871), .ZN(n16795) );
NAND2_X2 U12876 ( .A1(n16797), .A2(n16798), .ZN(N2834) );
NAND2_X2 U12877 ( .A1(v_out[19]), .A2(n18050), .ZN(n16798) );
NAND2_X2 U12878 ( .A1(n18062), .A2(n18872), .ZN(n16797) );
NAND2_X2 U12879 ( .A1(n16799), .A2(n16800), .ZN(N2833) );
NAND2_X2 U12880 ( .A1(v_out[18]), .A2(n18050), .ZN(n16800) );
NAND2_X2 U12881 ( .A1(n18061), .A2(n18873), .ZN(n16799) );
NAND2_X2 U12882 ( .A1(n16801), .A2(n16802), .ZN(N2832) );
NAND2_X2 U12883 ( .A1(v_out[17]), .A2(n18050), .ZN(n16802) );
NAND2_X2 U12884 ( .A1(n18061), .A2(n18874), .ZN(n16801) );
NAND2_X2 U12885 ( .A1(n16803), .A2(n16804), .ZN(N2831) );
NAND2_X2 U12886 ( .A1(v_out[16]), .A2(n18050), .ZN(n16804) );
NAND2_X2 U12887 ( .A1(n18061), .A2(n18875), .ZN(n16803) );
NAND2_X2 U12888 ( .A1(n16805), .A2(n16806), .ZN(N2830) );
NAND2_X2 U12889 ( .A1(v_out[15]), .A2(n18050), .ZN(n16806) );
NAND2_X2 U12890 ( .A1(n18061), .A2(n18876), .ZN(n16805) );
NAND2_X2 U12891 ( .A1(n16807), .A2(n16808), .ZN(N2829) );
NAND2_X2 U12892 ( .A1(v_out[14]), .A2(n18050), .ZN(n16808) );
NAND2_X2 U12893 ( .A1(n18061), .A2(n18877), .ZN(n16807) );
NAND2_X2 U12894 ( .A1(n16809), .A2(n16810), .ZN(N2828) );
NAND2_X2 U12895 ( .A1(v_out[13]), .A2(n18050), .ZN(n16810) );
NAND2_X2 U12896 ( .A1(n18061), .A2(n18878), .ZN(n16809) );
NAND2_X2 U12897 ( .A1(n16811), .A2(n16812), .ZN(N2827) );
NAND2_X2 U12898 ( .A1(v_out[12]), .A2(n18050), .ZN(n16812) );
NAND2_X2 U12899 ( .A1(n18061), .A2(n18879), .ZN(n16811) );
NAND2_X2 U12900 ( .A1(n16813), .A2(n16814), .ZN(N2826) );
NAND2_X2 U12901 ( .A1(v_out[11]), .A2(n18050), .ZN(n16814) );
NAND2_X2 U12902 ( .A1(n18061), .A2(n18880), .ZN(n16813) );
NAND2_X2 U12903 ( .A1(n16815), .A2(n16816), .ZN(N2825) );
NAND2_X2 U12904 ( .A1(v_out[10]), .A2(n18050), .ZN(n16816) );
NAND2_X2 U12905 ( .A1(n18061), .A2(n18881), .ZN(n16815) );
NAND2_X2 U12906 ( .A1(n16817), .A2(n16818), .ZN(N2824) );
NAND2_X2 U12907 ( .A1(v_out[9]), .A2(n18050), .ZN(n16818) );
NAND2_X2 U12908 ( .A1(n18061), .A2(n18882), .ZN(n16817) );
NAND2_X2 U12909 ( .A1(n16819), .A2(n16820), .ZN(N2823) );
NAND2_X2 U12910 ( .A1(v_out[8]), .A2(n18050), .ZN(n16820) );
NAND2_X2 U12911 ( .A1(n18061), .A2(n18883), .ZN(n16819) );
NAND2_X2 U12912 ( .A1(n16821), .A2(n16822), .ZN(N2822) );
NAND2_X2 U12913 ( .A1(v_out[7]), .A2(n18050), .ZN(n16822) );
NAND2_X2 U12914 ( .A1(n18061), .A2(n18884), .ZN(n16821) );
NAND2_X2 U12915 ( .A1(n16823), .A2(n16824), .ZN(N2821) );
NAND2_X2 U12916 ( .A1(v_out[6]), .A2(n18050), .ZN(n16824) );
NAND2_X2 U12917 ( .A1(n18061), .A2(n18885), .ZN(n16823) );
NAND2_X2 U12918 ( .A1(n16825), .A2(n16826), .ZN(N2820) );
NAND2_X2 U12919 ( .A1(v_out[5]), .A2(n18050), .ZN(n16826) );
NAND2_X2 U12920 ( .A1(n18061), .A2(n18886), .ZN(n16825) );
NAND2_X2 U12921 ( .A1(n16827), .A2(n16828), .ZN(N2819) );
NAND2_X2 U12922 ( .A1(v_out[4]), .A2(n18050), .ZN(n16828) );
NAND2_X2 U12923 ( .A1(n18061), .A2(n18887), .ZN(n16827) );
NAND2_X2 U12924 ( .A1(n16829), .A2(n16830), .ZN(N2818) );
NAND2_X2 U12925 ( .A1(v_out[3]), .A2(n18051), .ZN(n16830) );
NAND2_X2 U12926 ( .A1(n18061), .A2(n18888), .ZN(n16829) );
NAND2_X2 U12927 ( .A1(n16831), .A2(n16832), .ZN(N2817) );
NAND2_X2 U12928 ( .A1(v_out[2]), .A2(n18051), .ZN(n16832) );
NAND2_X2 U12929 ( .A1(n18061), .A2(n18889), .ZN(n16831) );
NAND2_X2 U12930 ( .A1(n16833), .A2(n16834), .ZN(N2816) );
NAND2_X2 U12931 ( .A1(v_out[1]), .A2(n18047), .ZN(n16834) );
NAND2_X2 U12932 ( .A1(n18061), .A2(n18890), .ZN(n16833) );
NAND2_X2 U12933 ( .A1(n16835), .A2(n16836), .ZN(N2815) );
NAND2_X2 U12934 ( .A1(v_out[0]), .A2(n18043), .ZN(n16836) );
NAND2_X2 U12935 ( .A1(n18059), .A2(n18891), .ZN(n16835) );
NAND2_X2 U12942 ( .A1(n18845), .A2(n18627), .ZN(n11976) );
NAND2_X2 U12944 ( .A1(n11973), .A2(n18600), .ZN(n16837) );
AND4_X2 U12945 ( .A1(n18628), .A2(n18631), .A3(n18629), .A4(n18626), .ZN(n11973) );
CLKBUFX1 gbuf_d_192(.A(n5437), .Y(d_out_192));
CLKBUFX1 gbuf_q_192(.A(q_in_192), .Y(enc_byte_cnt[4]));
CLKBUFX1 gbuf_qn_192(.A(qn_in_192), .Y(n5374));
CLKBUFX1 gbuf_d_193(.A(n5439), .Y(d_out_193));
CLKBUFX1 gbuf_q_193(.A(q_in_193), .Y(enc_byte_cnt[2]));
CLKBUFX1 gbuf_qn_193(.A(qn_in_193), .Y(n5376));
CLKBUFX1 gbuf_d_194(.A(n5440), .Y(d_out_194));
CLKBUFX1 gbuf_q_194(.A(q_in_194), .Y(enc_byte_cnt[1]));
CLKBUFX1 gbuf_qn_194(.A(qn_in_194), .Y(n5377));
CLKBUFX1 gbuf_d_195(.A(n5438), .Y(d_out_195));
CLKBUFX1 gbuf_q_195(.A(q_in_195), .Y(enc_byte_cnt[3]));
CLKBUFX1 gbuf_qn_195(.A(qn_in_195), .Y(n5375));
CLKBUFX1 gbuf_d_196(.A(n5436), .Y(d_out_196));
CLKBUFX1 gbuf_q_196(.A(q_in_196), .Y(enc_byte_cnt[5]));
CLKBUFX1 gbuf_d_197(.A(n5441), .Y(d_out_197));
CLKBUFX1 gbuf_q_197(.A(q_in_197), .Y(enc_byte_cnt[0]));
CLKBUFX1 gbuf_qn_197(.A(qn_in_197), .Y(n5378));
CLKBUFX1 gbuf_d_198(.A(n5425), .Y(d_out_198));
CLKBUFX1 gbuf_q_198(.A(q_in_198), .Y(enc_byte_cnt[16]));
CLKBUFX1 gbuf_qn_198(.A(qn_in_198), .Y(n5362));
CLKBUFX1 gbuf_d_199(.A(n5433), .Y(d_out_199));
CLKBUFX1 gbuf_q_199(.A(q_in_199), .Y(enc_byte_cnt[8]));
CLKBUFX1 gbuf_d_200(.A(n5435), .Y(d_out_200));
CLKBUFX1 gbuf_q_200(.A(q_in_200), .Y(enc_byte_cnt[6]));
CLKBUFX1 gbuf_d_201(.A(n5432), .Y(d_out_201));
CLKBUFX1 gbuf_q_201(.A(q_in_201), .Y(enc_byte_cnt[9]));
CLKBUFX1 gbuf_d_202(.A(n5429), .Y(d_out_202));
CLKBUFX1 gbuf_q_202(.A(q_in_202), .Y(enc_byte_cnt[12]));
CLKBUFX1 gbuf_d_203(.A(n5434), .Y(d_out_203));
CLKBUFX1 gbuf_q_203(.A(q_in_203), .Y(enc_byte_cnt[7]));
CLKBUFX1 gbuf_d_204(.A(n5417), .Y(d_out_204));
CLKBUFX1 gbuf_q_204(.A(q_in_204), .Y(enc_byte_cnt[24]));
CLKBUFX1 gbuf_d_205(.A(n5431), .Y(d_out_205));
CLKBUFX1 gbuf_q_205(.A(q_in_205), .Y(enc_byte_cnt[10]));
CLKBUFX1 gbuf_d_206(.A(n5428), .Y(d_out_206));
CLKBUFX1 gbuf_q_206(.A(q_in_206), .Y(enc_byte_cnt[13]));
CLKBUFX1 gbuf_qn_206(.A(qn_in_206), .Y(n5365));
CLKBUFX1 gbuf_d_207(.A(n5424), .Y(d_out_207));
CLKBUFX1 gbuf_q_207(.A(q_in_207), .Y(enc_byte_cnt[17]));
CLKBUFX1 gbuf_qn_207(.A(qn_in_207), .Y(n5361));
CLKBUFX1 gbuf_d_208(.A(n5421), .Y(d_out_208));
CLKBUFX1 gbuf_q_208(.A(q_in_208), .Y(enc_byte_cnt[20]));
CLKBUFX1 gbuf_qn_208(.A(qn_in_208), .Y(n5358));
CLKBUFX1 gbuf_d_209(.A(n5420), .Y(d_out_209));
CLKBUFX1 gbuf_q_209(.A(q_in_209), .Y(enc_byte_cnt[21]));
CLKBUFX1 gbuf_d_210(.A(n5423), .Y(d_out_210));
CLKBUFX1 gbuf_q_210(.A(q_in_210), .Y(enc_byte_cnt[18]));
CLKBUFX1 gbuf_qn_210(.A(qn_in_210), .Y(n5360));
CLKBUFX1 gbuf_d_211(.A(n6016), .Y(d_out_211));
CLKBUFX1 gbuf_q_211(.A(q_in_211), .Y(aad_byte_cnt[4]));
CLKBUFX1 gbuf_d_212(.A(n6018), .Y(d_out_212));
CLKBUFX1 gbuf_q_212(.A(q_in_212), .Y(aad_byte_cnt[2]));
CLKBUFX1 gbuf_d_213(.A(n6019), .Y(d_out_213));
CLKBUFX1 gbuf_q_213(.A(q_in_213), .Y(aad_byte_cnt[1]));
CLKBUFX1 gbuf_d_214(.A(n6017), .Y(d_out_214));
CLKBUFX1 gbuf_q_214(.A(q_in_214), .Y(aad_byte_cnt[3]));
CLKBUFX1 gbuf_d_215(.A(n6008), .Y(d_out_215));
CLKBUFX1 gbuf_q_215(.A(q_in_215), .Y(aad_byte_cnt[12]));
CLKBUFX1 gbuf_d_216(.A(n6010), .Y(d_out_216));
CLKBUFX1 gbuf_q_216(.A(q_in_216), .Y(aad_byte_cnt[10]));
CLKBUFX1 gbuf_d_217(.A(n6011), .Y(d_out_217));
CLKBUFX1 gbuf_q_217(.A(q_in_217), .Y(aad_byte_cnt[9]));
CLKBUFX1 gbuf_d_218(.A(n6012), .Y(d_out_218));
CLKBUFX1 gbuf_q_218(.A(q_in_218), .Y(aad_byte_cnt[8]));
CLKBUFX1 gbuf_d_219(.A(n6013), .Y(d_out_219));
CLKBUFX1 gbuf_q_219(.A(q_in_219), .Y(aad_byte_cnt[7]));
CLKBUFX1 gbuf_d_220(.A(n6014), .Y(d_out_220));
CLKBUFX1 gbuf_q_220(.A(q_in_220), .Y(aad_byte_cnt[6]));
CLKBUFX1 gbuf_d_221(.A(n6015), .Y(d_out_221));
CLKBUFX1 gbuf_q_221(.A(q_in_221), .Y(aad_byte_cnt[5]));
CLKBUFX1 gbuf_d_222(.A(n6020), .Y(d_out_222));
CLKBUFX1 gbuf_q_222(.A(q_in_222), .Y(aad_byte_cnt[0]));
CLKBUFX1 gbuf_d_223(.A(n5427), .Y(d_out_223));
CLKBUFX1 gbuf_q_223(.A(q_in_223), .Y(enc_byte_cnt[14]));
CLKBUFX1 gbuf_qn_223(.A(qn_in_223), .Y(n5364));
CLKBUFX1 gbuf_d_224(.A(n6004), .Y(d_out_224));
CLKBUFX1 gbuf_q_224(.A(q_in_224), .Y(aad_byte_cnt[16]));
CLKBUFX1 gbuf_d_225(.A(n5996), .Y(d_out_225));
CLKBUFX1 gbuf_q_225(.A(q_in_225), .Y(aad_byte_cnt[24]));
CLKBUFX1 gbuf_d_226(.A(n5999), .Y(d_out_226));
CLKBUFX1 gbuf_q_226(.A(q_in_226), .Y(aad_byte_cnt[21]));
CLKBUFX1 gbuf_d_227(.A(n6000), .Y(d_out_227));
CLKBUFX1 gbuf_q_227(.A(q_in_227), .Y(aad_byte_cnt[20]));
CLKBUFX1 gbuf_d_228(.A(n6002), .Y(d_out_228));
CLKBUFX1 gbuf_q_228(.A(q_in_228), .Y(aad_byte_cnt[18]));
CLKBUFX1 gbuf_d_229(.A(n6003), .Y(d_out_229));
CLKBUFX1 gbuf_q_229(.A(q_in_229), .Y(aad_byte_cnt[17]));
CLKBUFX1 gbuf_d_230(.A(n6006), .Y(d_out_230));
CLKBUFX1 gbuf_q_230(.A(q_in_230), .Y(aad_byte_cnt[14]));
CLKBUFX1 gbuf_d_231(.A(n6007), .Y(d_out_231));
CLKBUFX1 gbuf_q_231(.A(q_in_231), .Y(aad_byte_cnt[13]));
CLKBUFX1 gbuf_d_232(.A(n5413), .Y(d_out_232));
CLKBUFX1 gbuf_q_232(.A(q_in_232), .Y(enc_byte_cnt[28]));
CLKBUFX1 gbuf_d_233(.A(n5430), .Y(d_out_233));
CLKBUFX1 gbuf_q_233(.A(q_in_233), .Y(enc_byte_cnt[11]));
CLKBUFX1 gbuf_d_234(.A(n6009), .Y(d_out_234));
CLKBUFX1 gbuf_q_234(.A(q_in_234), .Y(aad_byte_cnt[11]));
CLKBUFX1 gbuf_d_235(.A(n5992), .Y(d_out_235));
CLKBUFX1 gbuf_q_235(.A(q_in_235), .Y(aad_byte_cnt[28]));
CLKBUFX1 gbuf_d_236(.A(n5416), .Y(d_out_236));
CLKBUFX1 gbuf_q_236(.A(q_in_236), .Y(enc_byte_cnt[25]));
CLKBUFX1 gbuf_d_237(.A(n5995), .Y(d_out_237));
CLKBUFX1 gbuf_q_237(.A(q_in_237), .Y(aad_byte_cnt[25]));
CLKBUFX1 gbuf_d_238(.A(n5426), .Y(d_out_238));
CLKBUFX1 gbuf_q_238(.A(q_in_238), .Y(enc_byte_cnt[15]));
CLKBUFX1 gbuf_qn_238(.A(qn_in_238), .Y(n5363));
CLKBUFX1 gbuf_d_239(.A(n6005), .Y(d_out_239));
CLKBUFX1 gbuf_q_239(.A(q_in_239), .Y(aad_byte_cnt[15]));
CLKBUFX1 gbuf_d_240(.A(n5405), .Y(d_out_240));
CLKBUFX1 gbuf_q_240(.A(q_in_240), .Y(enc_byte_cnt[36]));
CLKBUFX1 gbuf_qn_240(.A(qn_in_240), .Y(n5342));
CLKBUFX1 gbuf_d_241(.A(n5984), .Y(d_out_241));
CLKBUFX1 gbuf_q_241(.A(q_in_241), .Y(aad_byte_cnt[36]));
CLKBUFX1 gbuf_d_242(.A(n6001), .Y(d_out_242));
CLKBUFX1 gbuf_q_242(.A(q_in_242), .Y(aad_byte_cnt[19]));
CLKBUFX1 gbuf_d_243(.A(n5387), .Y(d_out_243));
CLKBUFX1 gbuf_q_243(.A(q_in_243), .Y(enc_byte_cnt[54]));
CLKBUFX1 gbuf_d_244(.A(n5966), .Y(d_out_244));
CLKBUFX1 gbuf_q_244(.A(q_in_244), .Y(aad_byte_cnt[54]));
CLKBUFX1 gbuf_d_245(.A(n5422), .Y(d_out_245));
CLKBUFX1 gbuf_q_245(.A(q_in_245), .Y(enc_byte_cnt[19]));
CLKBUFX1 gbuf_qn_245(.A(qn_in_245), .Y(n5359));
CLKBUFX1 gbuf_d_246(.A(n5419), .Y(d_out_246));
CLKBUFX1 gbuf_q_246(.A(q_in_246), .Y(enc_byte_cnt[22]));
CLKBUFX1 gbuf_d_247(.A(n5998), .Y(d_out_247));
CLKBUFX1 gbuf_q_247(.A(q_in_247), .Y(aad_byte_cnt[22]));
CLKBUFX1 gbuf_d_248(.A(n5991), .Y(d_out_248));
CLKBUFX1 gbuf_q_248(.A(q_in_248), .Y(aad_byte_cnt[29]));
CLKBUFX1 gbuf_d_249(.A(n5392), .Y(d_out_249));
CLKBUFX1 gbuf_q_249(.A(q_in_249), .Y(enc_byte_cnt[49]));
CLKBUFX1 gbuf_qn_249(.A(qn_in_249), .Y(n5329));
CLKBUFX1 gbuf_d_250(.A(n5412), .Y(d_out_250));
CLKBUFX1 gbuf_q_250(.A(q_in_250), .Y(enc_byte_cnt[29]));
CLKBUFX1 gbuf_qn_250(.A(qn_in_250), .Y(n5349));
CLKBUFX1 gbuf_d_251(.A(n5388), .Y(d_out_251));
CLKBUFX1 gbuf_q_251(.A(q_in_251), .Y(enc_byte_cnt[53]));
CLKBUFX1 gbuf_d_252(.A(n5381), .Y(d_out_252));
CLKBUFX1 gbuf_q_252(.A(q_in_252), .Y(enc_byte_cnt[60]));
CLKBUFX1 gbuf_d_253(.A(n5960), .Y(d_out_253));
CLKBUFX1 gbuf_q_253(.A(q_in_253), .Y(aad_byte_cnt[60]));
CLKBUFX1 gbuf_d_254(.A(n5971), .Y(d_out_254));
CLKBUFX1 gbuf_q_254(.A(q_in_254), .Y(aad_byte_cnt[49]));
CLKBUFX1 gbuf_d_255(.A(n5967), .Y(d_out_255));
CLKBUFX1 gbuf_q_255(.A(q_in_255), .Y(aad_byte_cnt[53]));
CLKBUFX1 gbuf_d_256(.A(n5968), .Y(d_out_256));
CLKBUFX1 gbuf_q_256(.A(q_in_256), .Y(aad_byte_cnt[52]));
CLKBUFX1 gbuf_d_257(.A(n5969), .Y(d_out_257));
CLKBUFX1 gbuf_q_257(.A(q_in_257), .Y(aad_byte_cnt[51]));
CLKBUFX1 gbuf_d_258(.A(n5411), .Y(d_out_258));
CLKBUFX1 gbuf_q_258(.A(q_in_258), .Y(enc_byte_cnt[30]));
CLKBUFX1 gbuf_qn_258(.A(qn_in_258), .Y(n5348));
CLKBUFX1 gbuf_d_259(.A(n5389), .Y(d_out_259));
CLKBUFX1 gbuf_q_259(.A(q_in_259), .Y(enc_byte_cnt[52]));
CLKBUFX1 gbuf_qn_259(.A(qn_in_259), .Y(n5326));
CLKBUFX1 gbuf_d_260(.A(n5390), .Y(d_out_260));
CLKBUFX1 gbuf_q_260(.A(q_in_260), .Y(enc_byte_cnt[51]));
CLKBUFX1 gbuf_qn_260(.A(qn_in_260), .Y(n5327));
CLKBUFX1 gbuf_d_261(.A(n5415), .Y(d_out_261));
CLKBUFX1 gbuf_q_261(.A(q_in_261), .Y(enc_byte_cnt[26]));
CLKBUFX1 gbuf_d_262(.A(n5994), .Y(d_out_262));
CLKBUFX1 gbuf_q_262(.A(q_in_262), .Y(aad_byte_cnt[26]));
CLKBUFX1 gbuf_d_263(.A(n5990), .Y(d_out_263));
CLKBUFX1 gbuf_q_263(.A(q_in_263), .Y(aad_byte_cnt[30]));
CLKBUFX1 gbuf_d_264(.A(n5382), .Y(d_out_264));
CLKBUFX1 gbuf_q_264(.A(q_in_264), .Y(enc_byte_cnt[59]));
CLKBUFX1 gbuf_d_265(.A(n5383), .Y(d_out_265));
CLKBUFX1 gbuf_q_265(.A(q_in_265), .Y(enc_byte_cnt[58]));
CLKBUFX1 gbuf_d_266(.A(n5384), .Y(d_out_266));
CLKBUFX1 gbuf_q_266(.A(q_in_266), .Y(enc_byte_cnt[57]));
CLKBUFX1 gbuf_d_267(.A(n5385), .Y(d_out_267));
CLKBUFX1 gbuf_q_267(.A(q_in_267), .Y(enc_byte_cnt[56]));
CLKBUFX1 gbuf_d_268(.A(n5961), .Y(d_out_268));
CLKBUFX1 gbuf_q_268(.A(q_in_268), .Y(aad_byte_cnt[59]));
CLKBUFX1 gbuf_d_269(.A(n5962), .Y(d_out_269));
CLKBUFX1 gbuf_q_269(.A(q_in_269), .Y(aad_byte_cnt[58]));
CLKBUFX1 gbuf_d_270(.A(n5963), .Y(d_out_270));
CLKBUFX1 gbuf_q_270(.A(q_in_270), .Y(aad_byte_cnt[57]));
CLKBUFX1 gbuf_d_271(.A(n5964), .Y(d_out_271));
CLKBUFX1 gbuf_q_271(.A(q_in_271), .Y(aad_byte_cnt[56]));
CLKBUFX1 gbuf_d_272(.A(n5404), .Y(d_out_272));
CLKBUFX1 gbuf_q_272(.A(q_in_272), .Y(enc_byte_cnt[37]));
CLKBUFX1 gbuf_d_273(.A(n5983), .Y(d_out_273));
CLKBUFX1 gbuf_q_273(.A(q_in_273), .Y(aad_byte_cnt[37]));
CLKBUFX1 gbuf_d_274(.A(n5409), .Y(d_out_274));
CLKBUFX1 gbuf_q_274(.A(q_in_274), .Y(enc_byte_cnt[32]));
CLKBUFX1 gbuf_qn_274(.A(qn_in_274), .Y(n5346));
CLKBUFX1 gbuf_d_275(.A(n5988), .Y(d_out_275));
CLKBUFX1 gbuf_q_275(.A(q_in_275), .Y(aad_byte_cnt[32]));
CLKBUFX1 gbuf_d_276(.A(n5386), .Y(d_out_276));
CLKBUFX1 gbuf_q_276(.A(q_in_276), .Y(enc_byte_cnt[55]));
CLKBUFX1 gbuf_d_277(.A(n5965), .Y(d_out_277));
CLKBUFX1 gbuf_q_277(.A(q_in_277), .Y(aad_byte_cnt[55]));
CLKBUFX1 gbuf_d_278(.A(n5407), .Y(d_out_278));
CLKBUFX1 gbuf_q_278(.A(q_in_278), .Y(enc_byte_cnt[34]));
CLKBUFX1 gbuf_qn_278(.A(qn_in_278), .Y(n5344));
CLKBUFX1 gbuf_d_279(.A(n5408), .Y(d_out_279));
CLKBUFX1 gbuf_q_279(.A(q_in_279), .Y(enc_byte_cnt[33]));
CLKBUFX1 gbuf_qn_279(.A(qn_in_279), .Y(n5345));
CLKBUFX1 gbuf_d_280(.A(n5986), .Y(d_out_280));
CLKBUFX1 gbuf_q_280(.A(q_in_280), .Y(aad_byte_cnt[34]));
CLKBUFX1 gbuf_d_281(.A(n5987), .Y(d_out_281));
CLKBUFX1 gbuf_q_281(.A(q_in_281), .Y(aad_byte_cnt[33]));
CLKBUFX1 gbuf_d_282(.A(n5403), .Y(d_out_282));
CLKBUFX1 gbuf_q_282(.A(q_in_282), .Y(enc_byte_cnt[38]));
CLKBUFX1 gbuf_d_283(.A(n5982), .Y(d_out_283));
CLKBUFX1 gbuf_q_283(.A(q_in_283), .Y(aad_byte_cnt[38]));
CLKBUFX1 gbuf_d_284(.A(n5418), .Y(d_out_284));
CLKBUFX1 gbuf_q_284(.A(q_in_284), .Y(enc_byte_cnt[23]));
CLKBUFX1 gbuf_d_285(.A(n5997), .Y(d_out_285));
CLKBUFX1 gbuf_q_285(.A(q_in_285), .Y(aad_byte_cnt[23]));
CLKBUFX1 gbuf_d_286(.A(n5391), .Y(d_out_286));
CLKBUFX1 gbuf_q_286(.A(q_in_286), .Y(enc_byte_cnt[50]));
CLKBUFX1 gbuf_qn_286(.A(qn_in_286), .Y(n5328));
CLKBUFX1 gbuf_d_287(.A(n5410), .Y(d_out_287));
CLKBUFX1 gbuf_q_287(.A(q_in_287), .Y(enc_byte_cnt[31]));
CLKBUFX1 gbuf_qn_287(.A(qn_in_287), .Y(n5347));
CLKBUFX1 gbuf_d_288(.A(n5970), .Y(d_out_288));
CLKBUFX1 gbuf_q_288(.A(q_in_288), .Y(aad_byte_cnt[50]));
CLKBUFX1 gbuf_d_289(.A(n5406), .Y(d_out_289));
CLKBUFX1 gbuf_q_289(.A(q_in_289), .Y(enc_byte_cnt[35]));
CLKBUFX1 gbuf_qn_289(.A(qn_in_289), .Y(n5343));
CLKBUFX1 gbuf_d_290(.A(n5985), .Y(d_out_290));
CLKBUFX1 gbuf_q_290(.A(q_in_290), .Y(aad_byte_cnt[35]));
CLKBUFX1 gbuf_d_291(.A(n5989), .Y(d_out_291));
CLKBUFX1 gbuf_q_291(.A(q_in_291), .Y(aad_byte_cnt[31]));
CLKBUFX1 gbuf_d_292(.A(n5414), .Y(d_out_292));
CLKBUFX1 gbuf_q_292(.A(q_in_292), .Y(enc_byte_cnt[27]));
CLKBUFX1 gbuf_d_293(.A(n5993), .Y(d_out_293));
CLKBUFX1 gbuf_q_293(.A(q_in_293), .Y(aad_byte_cnt[27]));
CLKBUFX1 gbuf_d_294(.A(n5972), .Y(d_out_294));
CLKBUFX1 gbuf_q_294(.A(q_in_294), .Y(aad_byte_cnt[48]));
CLKBUFX1 gbuf_d_295(.A(n5395), .Y(d_out_295));
CLKBUFX1 gbuf_q_295(.A(q_in_295), .Y(enc_byte_cnt[46]));
CLKBUFX1 gbuf_qn_295(.A(qn_in_295), .Y(n5332));
CLKBUFX1 gbuf_d_296(.A(n5974), .Y(d_out_296));
CLKBUFX1 gbuf_q_296(.A(q_in_296), .Y(aad_byte_cnt[46]));
CLKBUFX1 gbuf_d_297(.A(n5393), .Y(d_out_297));
CLKBUFX1 gbuf_q_297(.A(q_in_297), .Y(enc_byte_cnt[48]));
CLKBUFX1 gbuf_qn_297(.A(qn_in_297), .Y(n5330));
CLKBUFX1 gbuf_d_298(.A(n5394), .Y(d_out_298));
CLKBUFX1 gbuf_q_298(.A(q_in_298), .Y(enc_byte_cnt[47]));
CLKBUFX1 gbuf_qn_298(.A(qn_in_298), .Y(n5331));
CLKBUFX1 gbuf_d_299(.A(n5398), .Y(d_out_299));
CLKBUFX1 gbuf_q_299(.A(q_in_299), .Y(enc_byte_cnt[43]));
CLKBUFX1 gbuf_d_300(.A(n5973), .Y(d_out_300));
CLKBUFX1 gbuf_q_300(.A(q_in_300), .Y(aad_byte_cnt[47]));
CLKBUFX1 gbuf_d_301(.A(n5977), .Y(d_out_301));
CLKBUFX1 gbuf_q_301(.A(q_in_301), .Y(aad_byte_cnt[43]));
CLKBUFX1 gbuf_d_302(.A(n5402), .Y(d_out_302));
CLKBUFX1 gbuf_q_302(.A(q_in_302), .Y(enc_byte_cnt[39]));
CLKBUFX1 gbuf_d_303(.A(n5981), .Y(d_out_303));
CLKBUFX1 gbuf_q_303(.A(q_in_303), .Y(aad_byte_cnt[39]));
CLKBUFX1 gbuf_d_304(.A(n5399), .Y(d_out_304));
CLKBUFX1 gbuf_q_304(.A(q_in_304), .Y(enc_byte_cnt[42]));
CLKBUFX1 gbuf_d_305(.A(n5978), .Y(d_out_305));
CLKBUFX1 gbuf_q_305(.A(q_in_305), .Y(aad_byte_cnt[42]));
CLKBUFX1 gbuf_d_306(.A(n5397), .Y(d_out_306));
CLKBUFX1 gbuf_q_306(.A(q_in_306), .Y(enc_byte_cnt[44]));
CLKBUFX1 gbuf_d_307(.A(n5400), .Y(d_out_307));
CLKBUFX1 gbuf_q_307(.A(q_in_307), .Y(enc_byte_cnt[41]));
CLKBUFX1 gbuf_d_308(.A(n5401), .Y(d_out_308));
CLKBUFX1 gbuf_q_308(.A(q_in_308), .Y(enc_byte_cnt[40]));
CLKBUFX1 gbuf_d_309(.A(n5975), .Y(d_out_309));
CLKBUFX1 gbuf_q_309(.A(q_in_309), .Y(aad_byte_cnt[45]));
CLKBUFX1 gbuf_d_310(.A(n5976), .Y(d_out_310));
CLKBUFX1 gbuf_q_310(.A(q_in_310), .Y(aad_byte_cnt[44]));
CLKBUFX1 gbuf_d_311(.A(n5979), .Y(d_out_311));
CLKBUFX1 gbuf_q_311(.A(q_in_311), .Y(aad_byte_cnt[41]));
CLKBUFX1 gbuf_d_312(.A(n5980), .Y(d_out_312));
CLKBUFX1 gbuf_q_312(.A(q_in_312), .Y(aad_byte_cnt[40]));
CLKBUFX1 gbuf_d_313(.A(n5396), .Y(d_out_313));
CLKBUFX1 gbuf_q_313(.A(q_in_313), .Y(enc_byte_cnt[45]));
CLKBUFX1 gbuf_qn_313(.A(qn_in_313), .Y(n5333));
CLKBUFX1 gbuf_d_314(.A(n6283), .Y(d_out_314));
CLKBUFX1 gbuf_q_314(.A(q_in_314), .Y(state[0]));
CLKBUFX1 gbuf_qn_314(.A(qn_in_314), .Y(n18611));
CLKBUFX1 gbuf_d_315(.A(n6284), .Y(d_out_315));
CLKBUFX1 gbuf_q_315(.A(q_in_315), .Y(state[2]));
CLKBUFX1 gbuf_qn_315(.A(qn_in_315), .Y(n18630));
CLKBUFX1 gbuf_d_316(.A(n5442), .Y(d_out_316));
CLKBUFX1 gbuf_q_316(.A(q_in_316), .Y(enc_byte_cnt[63]));
CLKBUFX1 gbuf_d_317(.A(n6021), .Y(d_out_317));
CLKBUFX1 gbuf_q_317(.A(q_in_317), .Y(aad_byte_cnt[63]));
CLKBUFX1 gbuf_d_318(.A(n5379), .Y(d_out_318));
CLKBUFX1 gbuf_q_318(.A(q_in_318), .Y(enc_byte_cnt[62]));
CLKBUFX1 gbuf_d_319(.A(n5380), .Y(d_out_319));
CLKBUFX1 gbuf_q_319(.A(q_in_319), .Y(enc_byte_cnt[61]));
CLKBUFX1 gbuf_d_320(.A(n5958), .Y(d_out_320));
CLKBUFX1 gbuf_q_320(.A(q_in_320), .Y(aad_byte_cnt[62]));
CLKBUFX1 gbuf_d_321(.A(n5959), .Y(d_out_321));
CLKBUFX1 gbuf_q_321(.A(q_in_321), .Y(aad_byte_cnt[61]));
CLKBUFX1 gbuf_d_322(.A(n6286), .Y(d_out_322));
CLKBUFX1 gbuf_q_322(.A(q_in_322), .Y(state[5]));
CLKBUFX1 gbuf_qn_322(.A(qn_in_322), .Y(n18600));
CLKBUFX1 gbuf_d_323(.A(n6285), .Y(d_out_323));
CLKBUFX1 gbuf_q_323(.A(q_in_323), .Y(state[4]));
CLKBUFX1 gbuf_qn_323(.A(qn_in_323), .Y(n18629));
CLKBUFX1 gbuf_d_324(.A(n6292), .Y(d_out_324));
CLKBUFX1 gbuf_q_324(.A(q_in_324), .Y(state[1]));
CLKBUFX1 gbuf_qn_324(.A(qn_in_324), .Y(n18631));
CLKBUFX1 gbuf_d_325(.A(n6287), .Y(d_out_325));
CLKBUFX1 gbuf_q_325(.A(q_in_325), .Y(state[3]));
CLKBUFX1 gbuf_qn_325(.A(qn_in_325), .Y(n18078));
CLKBUFX1 gbuf_d_326(.A(n6293), .Y(d_out_326));
CLKBUFX1 gbuf_q_326(.A(q_in_326), .Y(state[8]));
CLKBUFX1 gbuf_qn_326(.A(qn_in_326), .Y(n18079));
CLKBUFX1 gbuf_d_327(.A(n6288), .Y(d_out_327));
CLKBUFX1 gbuf_q_327(.A(q_in_327), .Y(state[6]));
CLKBUFX1 gbuf_qn_327(.A(qn_in_327), .Y(n18626));
CLKBUFX1 gbuf_d_328(.A(n6294), .Y(d_out_328));
CLKBUFX1 gbuf_q_328(.A(q_in_328), .Y(state[9]));
CLKBUFX1 gbuf_qn_328(.A(qn_in_328), .Y(n18080));
CLKBUFX1 gbuf_d_329(.A(n6289), .Y(d_out_329));
CLKBUFX1 gbuf_q_329(.A(q_in_329), .Y(state[7]));
CLKBUFX1 gbuf_qn_329(.A(qn_in_329), .Y(n18601));
CLKBUFX1 gbuf_d_330(.A(n6152), .Y(d_out_330));
CLKBUFX1 gbuf_q_330(.A(q_in_330), .Y(n18889));
CLKBUFX1 gbuf_d_331(.A(n6153), .Y(d_out_331));
CLKBUFX1 gbuf_q_331(.A(q_in_331), .Y(n18890));
CLKBUFX1 gbuf_d_332(.A(n6154), .Y(d_out_332));
CLKBUFX1 gbuf_q_332(.A(q_in_332), .Y(n18891));
CLKBUFX1 gbuf_d_333(.A(n6110), .Y(d_out_333));
CLKBUFX1 gbuf_q_333(.A(q_in_333), .Y(n18847));
CLKBUFX1 gbuf_d_334(.A(n6111), .Y(d_out_334));
CLKBUFX1 gbuf_q_334(.A(q_in_334), .Y(n18848));
CLKBUFX1 gbuf_d_335(.A(n6112), .Y(d_out_335));
CLKBUFX1 gbuf_q_335(.A(q_in_335), .Y(n18849));
CLKBUFX1 gbuf_d_336(.A(n6113), .Y(d_out_336));
CLKBUFX1 gbuf_q_336(.A(q_in_336), .Y(n18850));
CLKBUFX1 gbuf_d_337(.A(n6114), .Y(d_out_337));
CLKBUFX1 gbuf_q_337(.A(q_in_337), .Y(n18851));
CLKBUFX1 gbuf_d_338(.A(n6115), .Y(d_out_338));
CLKBUFX1 gbuf_q_338(.A(q_in_338), .Y(n18852));
CLKBUFX1 gbuf_d_339(.A(n6116), .Y(d_out_339));
CLKBUFX1 gbuf_q_339(.A(q_in_339), .Y(n18853));
CLKBUFX1 gbuf_d_340(.A(n6117), .Y(d_out_340));
CLKBUFX1 gbuf_q_340(.A(q_in_340), .Y(n18854));
CLKBUFX1 gbuf_d_341(.A(n6118), .Y(d_out_341));
CLKBUFX1 gbuf_q_341(.A(q_in_341), .Y(n18855));
CLKBUFX1 gbuf_d_342(.A(n6119), .Y(d_out_342));
CLKBUFX1 gbuf_q_342(.A(q_in_342), .Y(n18856));
CLKBUFX1 gbuf_d_343(.A(n6120), .Y(d_out_343));
CLKBUFX1 gbuf_q_343(.A(q_in_343), .Y(n18857));
CLKBUFX1 gbuf_d_344(.A(n6121), .Y(d_out_344));
CLKBUFX1 gbuf_q_344(.A(q_in_344), .Y(n18858));
CLKBUFX1 gbuf_d_345(.A(n6122), .Y(d_out_345));
CLKBUFX1 gbuf_q_345(.A(q_in_345), .Y(n18859));
CLKBUFX1 gbuf_d_346(.A(n6123), .Y(d_out_346));
CLKBUFX1 gbuf_q_346(.A(q_in_346), .Y(n18860));
CLKBUFX1 gbuf_d_347(.A(n6124), .Y(d_out_347));
CLKBUFX1 gbuf_q_347(.A(q_in_347), .Y(n18861));
CLKBUFX1 gbuf_d_348(.A(n6125), .Y(d_out_348));
CLKBUFX1 gbuf_q_348(.A(q_in_348), .Y(n18862));
CLKBUFX1 gbuf_d_349(.A(n6126), .Y(d_out_349));
CLKBUFX1 gbuf_q_349(.A(q_in_349), .Y(n18863));
CLKBUFX1 gbuf_d_350(.A(n6127), .Y(d_out_350));
CLKBUFX1 gbuf_q_350(.A(q_in_350), .Y(n18864));
CLKBUFX1 gbuf_d_351(.A(n6128), .Y(d_out_351));
CLKBUFX1 gbuf_q_351(.A(q_in_351), .Y(n18865));
CLKBUFX1 gbuf_d_352(.A(n6129), .Y(d_out_352));
CLKBUFX1 gbuf_q_352(.A(q_in_352), .Y(n18866));
CLKBUFX1 gbuf_d_353(.A(n6130), .Y(d_out_353));
CLKBUFX1 gbuf_q_353(.A(q_in_353), .Y(n18867));
CLKBUFX1 gbuf_d_354(.A(n6131), .Y(d_out_354));
CLKBUFX1 gbuf_q_354(.A(q_in_354), .Y(n18868));
CLKBUFX1 gbuf_d_355(.A(n6132), .Y(d_out_355));
CLKBUFX1 gbuf_q_355(.A(q_in_355), .Y(n18869));
CLKBUFX1 gbuf_d_356(.A(n6133), .Y(d_out_356));
CLKBUFX1 gbuf_q_356(.A(q_in_356), .Y(n18870));
CLKBUFX1 gbuf_d_357(.A(n6134), .Y(d_out_357));
CLKBUFX1 gbuf_q_357(.A(q_in_357), .Y(n18871));
CLKBUFX1 gbuf_d_358(.A(n6135), .Y(d_out_358));
CLKBUFX1 gbuf_q_358(.A(q_in_358), .Y(n18872));
CLKBUFX1 gbuf_d_359(.A(n6136), .Y(d_out_359));
CLKBUFX1 gbuf_q_359(.A(q_in_359), .Y(n18873));
CLKBUFX1 gbuf_d_360(.A(n6137), .Y(d_out_360));
CLKBUFX1 gbuf_q_360(.A(q_in_360), .Y(n18874));
CLKBUFX1 gbuf_d_361(.A(n6138), .Y(d_out_361));
CLKBUFX1 gbuf_q_361(.A(q_in_361), .Y(n18875));
CLKBUFX1 gbuf_d_362(.A(n6139), .Y(d_out_362));
CLKBUFX1 gbuf_q_362(.A(q_in_362), .Y(n18876));
CLKBUFX1 gbuf_d_363(.A(n6140), .Y(d_out_363));
CLKBUFX1 gbuf_q_363(.A(q_in_363), .Y(n18877));
CLKBUFX1 gbuf_d_364(.A(n6141), .Y(d_out_364));
CLKBUFX1 gbuf_q_364(.A(q_in_364), .Y(n18878));
CLKBUFX1 gbuf_d_365(.A(n6142), .Y(d_out_365));
CLKBUFX1 gbuf_q_365(.A(q_in_365), .Y(n18879));
CLKBUFX1 gbuf_d_366(.A(n6143), .Y(d_out_366));
CLKBUFX1 gbuf_q_366(.A(q_in_366), .Y(n18880));
CLKBUFX1 gbuf_d_367(.A(n6144), .Y(d_out_367));
CLKBUFX1 gbuf_q_367(.A(q_in_367), .Y(n18881));
CLKBUFX1 gbuf_d_368(.A(n6145), .Y(d_out_368));
CLKBUFX1 gbuf_q_368(.A(q_in_368), .Y(n18882));
CLKBUFX1 gbuf_d_369(.A(n6146), .Y(d_out_369));
CLKBUFX1 gbuf_q_369(.A(q_in_369), .Y(n18883));
CLKBUFX1 gbuf_d_370(.A(n6147), .Y(d_out_370));
CLKBUFX1 gbuf_q_370(.A(q_in_370), .Y(n18884));
CLKBUFX1 gbuf_d_371(.A(n6148), .Y(d_out_371));
CLKBUFX1 gbuf_q_371(.A(q_in_371), .Y(n18885));
CLKBUFX1 gbuf_d_372(.A(n6149), .Y(d_out_372));
CLKBUFX1 gbuf_q_372(.A(q_in_372), .Y(n18886));
CLKBUFX1 gbuf_d_373(.A(n6150), .Y(d_out_373));
CLKBUFX1 gbuf_q_373(.A(q_in_373), .Y(n18887));
CLKBUFX1 gbuf_d_374(.A(n6151), .Y(d_out_374));
CLKBUFX1 gbuf_q_374(.A(q_in_374), .Y(n18888));
CLKBUFX1 gbuf_d_375(.A(n6232), .Y(d_out_375));
CLKBUFX1 gbuf_qn_375(.A(qn_in_375), .Y(n17179));
CLKBUFX1 gbuf_d_376(.A(n6233), .Y(d_out_376));
CLKBUFX1 gbuf_qn_376(.A(qn_in_376), .Y(n17181));
CLKBUFX1 gbuf_d_377(.A(n6234), .Y(d_out_377));
CLKBUFX1 gbuf_qn_377(.A(qn_in_377), .Y(n17183));
CLKBUFX1 gbuf_d_378(.A(n6235), .Y(d_out_378));
CLKBUFX1 gbuf_qn_378(.A(qn_in_378), .Y(n17185));
CLKBUFX1 gbuf_d_379(.A(n6236), .Y(d_out_379));
CLKBUFX1 gbuf_qn_379(.A(qn_in_379), .Y(n17187));
CLKBUFX1 gbuf_d_380(.A(n6237), .Y(d_out_380));
CLKBUFX1 gbuf_qn_380(.A(qn_in_380), .Y(n17189));
CLKBUFX1 gbuf_d_381(.A(n6238), .Y(d_out_381));
CLKBUFX1 gbuf_qn_381(.A(qn_in_381), .Y(n17191));
CLKBUFX1 gbuf_d_382(.A(n6240), .Y(d_out_382));
CLKBUFX1 gbuf_qn_382(.A(qn_in_382), .Y(n17195));
CLKBUFX1 gbuf_d_383(.A(n6241), .Y(d_out_383));
CLKBUFX1 gbuf_qn_383(.A(qn_in_383), .Y(n17197));
CLKBUFX1 gbuf_d_384(.A(n6242), .Y(d_out_384));
CLKBUFX1 gbuf_qn_384(.A(qn_in_384), .Y(n17199));
CLKBUFX1 gbuf_d_385(.A(n6243), .Y(d_out_385));
CLKBUFX1 gbuf_qn_385(.A(qn_in_385), .Y(n17201));
CLKBUFX1 gbuf_d_386(.A(n6155), .Y(d_out_386));
CLKBUFX1 gbuf_qn_386(.A(qn_in_386), .Y(n17025));
CLKBUFX1 gbuf_d_387(.A(n6158), .Y(d_out_387));
CLKBUFX1 gbuf_qn_387(.A(qn_in_387), .Y(n17031));
CLKBUFX1 gbuf_d_388(.A(n6160), .Y(d_out_388));
CLKBUFX1 gbuf_qn_388(.A(qn_in_388), .Y(n17035));
CLKBUFX1 gbuf_d_389(.A(n6280), .Y(d_out_389));
CLKBUFX1 gbuf_qn_389(.A(qn_in_389), .Y(n17275));
CLKBUFX1 gbuf_d_390(.A(n6281), .Y(d_out_390));
CLKBUFX1 gbuf_qn_390(.A(qn_in_390), .Y(n17277));
CLKBUFX1 gbuf_d_391(.A(n6260), .Y(d_out_391));
CLKBUFX1 gbuf_qn_391(.A(qn_in_391), .Y(n17235));
CLKBUFX1 gbuf_d_392(.A(n6261), .Y(d_out_392));
CLKBUFX1 gbuf_qn_392(.A(qn_in_392), .Y(n17237));
CLKBUFX1 gbuf_d_393(.A(n6263), .Y(d_out_393));
CLKBUFX1 gbuf_qn_393(.A(qn_in_393), .Y(n17241));
CLKBUFX1 gbuf_d_394(.A(n6264), .Y(d_out_394));
CLKBUFX1 gbuf_qn_394(.A(qn_in_394), .Y(n17243));
CLKBUFX1 gbuf_d_649(.A(n5827), .Y(ddout__649));
CLKBUFX1 gbuf_q_649(.A(qq_in649), .Y(n18897));
CLKBUFX1 gbuf_qn_649(.A(qnn_in_649), .Y(n17274));
CLKBUFX1 gbuf_d_650(.A(n5829), .Y(ddout__650));
CLKBUFX1 gbuf_q_650(.A(qq_in650), .Y(n18895));
CLKBUFX1 gbuf_qn_650(.A(qnn_in_650), .Y(n17278));
CLKBUFX1 gbuf_d_651(.A(n5826), .Y(ddout__651));
CLKBUFX1 gbuf_q_651(.A(qq_in651), .Y(n18898));
CLKBUFX1 gbuf_qn_651(.A(qnn_in_651), .Y(n17272));
CLKBUFX1 gbuf_d_652(.A(n5796), .Y(ddout__652));
CLKBUFX1 gbuf_q_652(.A(qq_in652), .Y(n18928));
CLKBUFX1 gbuf_d_653(.A(n5815), .Y(ddout__653));
CLKBUFX1 gbuf_q_653(.A(qq_in653), .Y(n18909));
CLKBUFX1 gbuf_d_654(.A(n5825), .Y(ddout__654));
CLKBUFX1 gbuf_q_654(.A(qq_in654), .Y(n18899));
CLKBUFX1 gbuf_qn_654(.A(qnn_in_654), .Y(n17270));
CLKBUFX1 gbuf_d_655(.A(n5793), .Y(ddout__655));
CLKBUFX1 gbuf_q_655(.A(qq_in655), .Y(n18931));
CLKBUFX1 gbuf_d_656(.A(n5789), .Y(ddout__656));
CLKBUFX1 gbuf_q_656(.A(qq_in656), .Y(n18935));
CLKBUFX1 gbuf_d_657(.A(n5790), .Y(ddout__657));
CLKBUFX1 gbuf_q_657(.A(qq_in657), .Y(n18934));
CLKBUFX1 gbuf_d_658(.A(n5788), .Y(ddout__658));
CLKBUFX1 gbuf_q_658(.A(qq_in658), .Y(n18936));
CLKBUFX1 gbuf_d_659(.A(n5791), .Y(ddout__659));
CLKBUFX1 gbuf_q_659(.A(qq_in659), .Y(n18933));
CLKBUFX1 gbuf_d_660(.A(n5792), .Y(ddout__660));
CLKBUFX1 gbuf_q_660(.A(qq_in660), .Y(n18932));
CLKBUFX1 gbuf_d_661(.A(n5786), .Y(ddout__661));
CLKBUFX1 gbuf_q_661(.A(qq_in661), .Y(n18938));
CLKBUFX1 gbuf_d_662(.A(n5787), .Y(ddout__662));
CLKBUFX1 gbuf_q_662(.A(qq_in662), .Y(n18937));
CLKBUFX1 gbuf_d_663(.A(n5785), .Y(ddout__663));
CLKBUFX1 gbuf_q_663(.A(qq_in663), .Y(n18939));
CLKBUFX1 gbuf_d_664(.A(n5784), .Y(ddout__664));
CLKBUFX1 gbuf_q_664(.A(qq_in664), .Y(n18940));
CLKBUFX1 gbuf_d_665(.A(n5794), .Y(ddout__665));
CLKBUFX1 gbuf_q_665(.A(qq_in665), .Y(n18930));
CLKBUFX1 gbuf_d_666(.A(n5816), .Y(ddout__666));
CLKBUFX1 gbuf_q_666(.A(qq_in666), .Y(n18908));
CLKBUFX1 gbuf_d_667(.A(n5828), .Y(ddout__667));
CLKBUFX1 gbuf_q_667(.A(qq_in667), .Y(n18896));
CLKBUFX1 gbuf_qn_667(.A(qnn_in_667), .Y(n17276));
CLKBUFX1 gbuf_d_668(.A(n5823), .Y(ddout__668));
CLKBUFX1 gbuf_q_668(.A(qq_in668), .Y(n18901));
CLKBUFX1 gbuf_qn_668(.A(qnn_in_668), .Y(n17266));
CLKBUFX1 gbuf_d_669(.A(n5824), .Y(ddout__669));
CLKBUFX1 gbuf_q_669(.A(qq_in669), .Y(n18900));
CLKBUFX1 gbuf_qn_669(.A(qnn_in_669), .Y(n17268));
CLKBUFX1 gbuf_d_670(.A(n5822), .Y(ddout__670));
CLKBUFX1 gbuf_q_670(.A(qq_in670), .Y(n18902));
CLKBUFX1 gbuf_qn_670(.A(qnn_in_670), .Y(n17264));
CLKBUFX1 gbuf_d_671(.A(n5821), .Y(ddout__671));
CLKBUFX1 gbuf_q_671(.A(qq_in671), .Y(n18903));
CLKBUFX1 gbuf_d_672(.A(n5820), .Y(ddout__672));
CLKBUFX1 gbuf_q_672(.A(qq_in672), .Y(n18904));
CLKBUFX1 gbuf_d_673(.A(n5799), .Y(ddout__673));
CLKBUFX1 gbuf_q_673(.A(qq_in673), .Y(n18925));
CLKBUFX1 gbuf_d_674(.A(n5800), .Y(ddout__674));
CLKBUFX1 gbuf_q_674(.A(qq_in674), .Y(n18924));
CLKBUFX1 gbuf_d_675(.A(n5801), .Y(ddout__675));
CLKBUFX1 gbuf_q_675(.A(qq_in675), .Y(n18923));
CLKBUFX1 gbuf_d_676(.A(n5803), .Y(ddout__676));
CLKBUFX1 gbuf_q_676(.A(qq_in676), .Y(n18921));
CLKBUFX1 gbuf_d_677(.A(n5804), .Y(ddout__677));
CLKBUFX1 gbuf_q_677(.A(qq_in677), .Y(n18920));
CLKBUFX1 gbuf_d_678(.A(n5805), .Y(ddout__678));
CLKBUFX1 gbuf_q_678(.A(qq_in678), .Y(n18919));
CLKBUFX1 gbuf_d_679(.A(n5806), .Y(ddout__679));
CLKBUFX1 gbuf_q_679(.A(qq_in679), .Y(n18918));
CLKBUFX1 gbuf_d_680(.A(n5808), .Y(ddout__680));
CLKBUFX1 gbuf_q_680(.A(qq_in680), .Y(n18916));
CLKBUFX1 gbuf_d_681(.A(n5809), .Y(ddout__681));
CLKBUFX1 gbuf_q_681(.A(qq_in681), .Y(n18915));
CLKBUFX1 gbuf_d_682(.A(n5813), .Y(ddout__682));
CLKBUFX1 gbuf_q_682(.A(qq_in682), .Y(n18911));
CLKBUFX1 gbuf_d_683(.A(n5795), .Y(ddout__683));
CLKBUFX1 gbuf_q_683(.A(qq_in683), .Y(n18929));
CLKBUFX1 gbuf_d_684(.A(n5819), .Y(ddout__684));
CLKBUFX1 gbuf_q_684(.A(qq_in684), .Y(n18905));
CLKBUFX1 gbuf_d_685(.A(n5783), .Y(ddout__685));
CLKBUFX1 gbuf_q_685(.A(qq_in685), .Y(n18941));
CLKBUFX1 gbuf_d_686(.A(n5719), .Y(ddout__686));
CLKBUFX1 gbuf_q_686(.A(qq_in686), .Y(n19005));
CLKBUFX1 gbuf_d_687(.A(n5720), .Y(ddout__687));
CLKBUFX1 gbuf_q_687(.A(qq_in687), .Y(n19004));
CLKBUFX1 gbuf_d_688(.A(n5721), .Y(ddout__688));
CLKBUFX1 gbuf_q_688(.A(qq_in688), .Y(n19003));
CLKBUFX1 gbuf_d_689(.A(n5722), .Y(ddout__689));
CLKBUFX1 gbuf_q_689(.A(qq_in689), .Y(n19002));
CLKBUFX1 gbuf_d_690(.A(n5723), .Y(ddout__690));
CLKBUFX1 gbuf_q_690(.A(qq_in690), .Y(n19001));
CLKBUFX1 gbuf_d_691(.A(n5724), .Y(ddout__691));
CLKBUFX1 gbuf_q_691(.A(qq_in691), .Y(n19000));
CLKBUFX1 gbuf_d_692(.A(n5725), .Y(ddout__692));
CLKBUFX1 gbuf_q_692(.A(qq_in692), .Y(n18999));
CLKBUFX1 gbuf_d_693(.A(n5726), .Y(ddout__693));
CLKBUFX1 gbuf_q_693(.A(qq_in693), .Y(n18998));
CLKBUFX1 gbuf_d_694(.A(n5727), .Y(ddout__694));
CLKBUFX1 gbuf_q_694(.A(qq_in694), .Y(n18997));
CLKBUFX1 gbuf_d_695(.A(n5728), .Y(ddout__695));
CLKBUFX1 gbuf_q_695(.A(qq_in695), .Y(n18996));
CLKBUFX1 gbuf_d_696(.A(n5729), .Y(ddout__696));
CLKBUFX1 gbuf_q_696(.A(qq_in696), .Y(n18995));
CLKBUFX1 gbuf_d_697(.A(n5730), .Y(ddout__697));
CLKBUFX1 gbuf_q_697(.A(qq_in697), .Y(n18994));
CLKBUFX1 gbuf_d_698(.A(n5731), .Y(ddout__698));
CLKBUFX1 gbuf_q_698(.A(qq_in698), .Y(n18993));
CLKBUFX1 gbuf_d_699(.A(n5732), .Y(ddout__699));
CLKBUFX1 gbuf_q_699(.A(qq_in699), .Y(n18992));
CLKBUFX1 gbuf_d_700(.A(n5733), .Y(ddout__700));
CLKBUFX1 gbuf_q_700(.A(qq_in700), .Y(n18991));
CLKBUFX1 gbuf_d_701(.A(n5734), .Y(ddout__701));
CLKBUFX1 gbuf_q_701(.A(qq_in701), .Y(n18990));
CLKBUFX1 gbuf_d_702(.A(n5735), .Y(ddout__702));
CLKBUFX1 gbuf_q_702(.A(qq_in702), .Y(n18989));
CLKBUFX1 gbuf_d_703(.A(n5736), .Y(ddout__703));
CLKBUFX1 gbuf_q_703(.A(qq_in703), .Y(n18988));
CLKBUFX1 gbuf_d_704(.A(n5737), .Y(ddout__704));
CLKBUFX1 gbuf_q_704(.A(qq_in704), .Y(n18987));
CLKBUFX1 gbuf_d_705(.A(n5738), .Y(ddout__705));
CLKBUFX1 gbuf_q_705(.A(qq_in705), .Y(n18986));
CLKBUFX1 gbuf_d_706(.A(n5739), .Y(ddout__706));
CLKBUFX1 gbuf_q_706(.A(qq_in706), .Y(n18985));
CLKBUFX1 gbuf_d_707(.A(n5740), .Y(ddout__707));
CLKBUFX1 gbuf_q_707(.A(qq_in707), .Y(n18984));
CLKBUFX1 gbuf_d_708(.A(n5741), .Y(ddout__708));
CLKBUFX1 gbuf_q_708(.A(qq_in708), .Y(n18983));
CLKBUFX1 gbuf_d_709(.A(n5742), .Y(ddout__709));
CLKBUFX1 gbuf_q_709(.A(qq_in709), .Y(n18982));
CLKBUFX1 gbuf_d_710(.A(n5743), .Y(ddout__710));
CLKBUFX1 gbuf_q_710(.A(qq_in710), .Y(n18981));
CLKBUFX1 gbuf_d_711(.A(n5744), .Y(ddout__711));
CLKBUFX1 gbuf_q_711(.A(qq_in711), .Y(n18980));
CLKBUFX1 gbuf_d_712(.A(n5745), .Y(ddout__712));
CLKBUFX1 gbuf_q_712(.A(qq_in712), .Y(n18979));
CLKBUFX1 gbuf_d_713(.A(n5746), .Y(ddout__713));
CLKBUFX1 gbuf_q_713(.A(qq_in713), .Y(n18978));
CLKBUFX1 gbuf_d_714(.A(n5747), .Y(ddout__714));
CLKBUFX1 gbuf_q_714(.A(qq_in714), .Y(n18977));
CLKBUFX1 gbuf_d_715(.A(n5748), .Y(ddout__715));
CLKBUFX1 gbuf_q_715(.A(qq_in715), .Y(n18976));
CLKBUFX1 gbuf_d_716(.A(n5749), .Y(ddout__716));
CLKBUFX1 gbuf_q_716(.A(qq_in716), .Y(n18975));
CLKBUFX1 gbuf_d_717(.A(n5750), .Y(ddout__717));
CLKBUFX1 gbuf_q_717(.A(qq_in717), .Y(n18974));
CLKBUFX1 gbuf_d_718(.A(n5751), .Y(ddout__718));
CLKBUFX1 gbuf_q_718(.A(qq_in718), .Y(n18973));
CLKBUFX1 gbuf_d_719(.A(n5752), .Y(ddout__719));
CLKBUFX1 gbuf_q_719(.A(qq_in719), .Y(n18972));
CLKBUFX1 gbuf_d_720(.A(n5753), .Y(ddout__720));
CLKBUFX1 gbuf_q_720(.A(qq_in720), .Y(n18971));
CLKBUFX1 gbuf_d_721(.A(n5754), .Y(ddout__721));
CLKBUFX1 gbuf_q_721(.A(qq_in721), .Y(n18970));
CLKBUFX1 gbuf_d_722(.A(n5755), .Y(ddout__722));
CLKBUFX1 gbuf_q_722(.A(qq_in722), .Y(n18969));
CLKBUFX1 gbuf_d_723(.A(n5756), .Y(ddout__723));
CLKBUFX1 gbuf_q_723(.A(qq_in723), .Y(n18968));
CLKBUFX1 gbuf_d_724(.A(n5757), .Y(ddout__724));
CLKBUFX1 gbuf_q_724(.A(qq_in724), .Y(n18967));
CLKBUFX1 gbuf_d_725(.A(n5758), .Y(ddout__725));
CLKBUFX1 gbuf_q_725(.A(qq_in725), .Y(n18966));
CLKBUFX1 gbuf_d_726(.A(n5759), .Y(ddout__726));
CLKBUFX1 gbuf_q_726(.A(qq_in726), .Y(n18965));
CLKBUFX1 gbuf_d_727(.A(n5760), .Y(ddout__727));
CLKBUFX1 gbuf_q_727(.A(qq_in727), .Y(n18964));
CLKBUFX1 gbuf_d_728(.A(n5761), .Y(ddout__728));
CLKBUFX1 gbuf_q_728(.A(qq_in728), .Y(n18963));
CLKBUFX1 gbuf_d_729(.A(n5762), .Y(ddout__729));
CLKBUFX1 gbuf_q_729(.A(qq_in729), .Y(n18962));
CLKBUFX1 gbuf_d_730(.A(n5763), .Y(ddout__730));
CLKBUFX1 gbuf_q_730(.A(qq_in730), .Y(n18961));
CLKBUFX1 gbuf_d_731(.A(n5764), .Y(ddout__731));
CLKBUFX1 gbuf_q_731(.A(qq_in731), .Y(n18960));
CLKBUFX1 gbuf_d_732(.A(n5765), .Y(ddout__732));
CLKBUFX1 gbuf_q_732(.A(qq_in732), .Y(n18959));
CLKBUFX1 gbuf_d_733(.A(n5766), .Y(ddout__733));
CLKBUFX1 gbuf_q_733(.A(qq_in733), .Y(n18958));
CLKBUFX1 gbuf_d_734(.A(n5767), .Y(ddout__734));
CLKBUFX1 gbuf_q_734(.A(qq_in734), .Y(n18957));
CLKBUFX1 gbuf_d_735(.A(n5768), .Y(ddout__735));
CLKBUFX1 gbuf_q_735(.A(qq_in735), .Y(n18956));
CLKBUFX1 gbuf_d_736(.A(n5769), .Y(ddout__736));
CLKBUFX1 gbuf_q_736(.A(qq_in736), .Y(n18955));
CLKBUFX1 gbuf_d_737(.A(n5770), .Y(ddout__737));
CLKBUFX1 gbuf_q_737(.A(qq_in737), .Y(n18954));
CLKBUFX1 gbuf_d_738(.A(n5771), .Y(ddout__738));
CLKBUFX1 gbuf_q_738(.A(qq_in738), .Y(n18953));
CLKBUFX1 gbuf_d_739(.A(n5772), .Y(ddout__739));
CLKBUFX1 gbuf_q_739(.A(qq_in739), .Y(n18952));
CLKBUFX1 gbuf_d_740(.A(n5773), .Y(ddout__740));
CLKBUFX1 gbuf_q_740(.A(qq_in740), .Y(n18951));
CLKBUFX1 gbuf_d_741(.A(n5774), .Y(ddout__741));
CLKBUFX1 gbuf_q_741(.A(qq_in741), .Y(n18950));
CLKBUFX1 gbuf_d_742(.A(n5775), .Y(ddout__742));
CLKBUFX1 gbuf_q_742(.A(qq_in742), .Y(n18949));
CLKBUFX1 gbuf_d_743(.A(n5776), .Y(ddout__743));
CLKBUFX1 gbuf_q_743(.A(qq_in743), .Y(n18948));
CLKBUFX1 gbuf_d_744(.A(n5777), .Y(ddout__744));
CLKBUFX1 gbuf_q_744(.A(qq_in744), .Y(n18947));
CLKBUFX1 gbuf_d_745(.A(n5778), .Y(ddout__745));
CLKBUFX1 gbuf_q_745(.A(qq_in745), .Y(n18946));
CLKBUFX1 gbuf_d_746(.A(n5779), .Y(ddout__746));
CLKBUFX1 gbuf_q_746(.A(qq_in746), .Y(n18945));
CLKBUFX1 gbuf_d_747(.A(n5780), .Y(ddout__747));
CLKBUFX1 gbuf_q_747(.A(qq_in747), .Y(n18944));
CLKBUFX1 gbuf_d_748(.A(n5781), .Y(ddout__748));
CLKBUFX1 gbuf_q_748(.A(qq_in748), .Y(n18943));
CLKBUFX1 gbuf_d_749(.A(n5782), .Y(ddout__749));
CLKBUFX1 gbuf_q_749(.A(qq_in749), .Y(n18942));
CLKBUFX1 gbuf_d_750(.A(n5802), .Y(ddout__750));
CLKBUFX1 gbuf_q_750(.A(qq_in750), .Y(n18922));
CLKBUFX1 gbuf_d_751(.A(n5807), .Y(ddout__751));
CLKBUFX1 gbuf_q_751(.A(qq_in751), .Y(n18917));
CLKBUFX1 gbuf_d_752(.A(n5810), .Y(ddout__752));
CLKBUFX1 gbuf_q_752(.A(qq_in752), .Y(n18914));
CLKBUFX1 gbuf_d_753(.A(n5811), .Y(ddout__753));
CLKBUFX1 gbuf_q_753(.A(qq_in753), .Y(n18913));
CLKBUFX1 gbuf_d_754(.A(n5812), .Y(ddout__754));
CLKBUFX1 gbuf_q_754(.A(qq_in754), .Y(n18912));
CLKBUFX1 gbuf_d_755(.A(n5814), .Y(ddout__755));
CLKBUFX1 gbuf_q_755(.A(qq_in755), .Y(n18910));
CLKBUFX1 gbuf_d_756(.A(n5818), .Y(ddout__756));
CLKBUFX1 gbuf_q_756(.A(qq_in756), .Y(n18906));
CLKBUFX1 gbuf_d_757(.A(n5798), .Y(ddout__757));
CLKBUFX1 gbuf_q_757(.A(qq_in757), .Y(n18926));
CLKBUFX1 gbuf_d_758(.A(n5797), .Y(ddout__758));
CLKBUFX1 gbuf_q_758(.A(qq_in758), .Y(n18927));
CLKBUFX1 gbuf_d_759(.A(n5817), .Y(ddout__759));
CLKBUFX1 gbuf_q_759(.A(qq_in759), .Y(n18907));
CLKBUFX1 gbuf_d_760(.A(n5702), .Y(ddout__760));
CLKBUFX1 gbuf_q_760(.A(qq_in760), .Y(n19022));
CLKBUFX1 gbuf_qn_760(.A(qnn_in_760), .Y(n17024));
CLKBUFX1 gbuf_d_761(.A(n5705), .Y(ddout__761));
CLKBUFX1 gbuf_q_761(.A(qq_in761), .Y(n19019));
CLKBUFX1 gbuf_qn_761(.A(qnn_in_761), .Y(n17030));
CLKBUFX1 gbuf_d_762(.A(n5708), .Y(ddout__762));
CLKBUFX1 gbuf_q_762(.A(qq_in762), .Y(n19016));
CLKBUFX1 gbuf_qn_762(.A(qnn_in_762), .Y(n17036));
CLKBUFX1 gbuf_d_763(.A(n5706), .Y(ddout__763));
CLKBUFX1 gbuf_q_763(.A(qq_in763), .Y(n19018));
CLKBUFX1 gbuf_qn_763(.A(qnn_in_763), .Y(n17032));
CLKBUFX1 gbuf_d_764(.A(n5707), .Y(ddout__764));
CLKBUFX1 gbuf_q_764(.A(qq_in764), .Y(n19017));
CLKBUFX1 gbuf_qn_764(.A(qnn_in_764), .Y(n17034));
CLKBUFX1 gbuf_d_765(.A(n5718), .Y(ddout__765));
CLKBUFX1 gbuf_q_765(.A(qq_in765), .Y(n19006));
CLKBUFX1 gbuf_d_766(.A(n5703), .Y(ddout__766));
CLKBUFX1 gbuf_q_766(.A(qq_in766), .Y(n19021));
CLKBUFX1 gbuf_qn_766(.A(qnn_in_766), .Y(n17026));
CLKBUFX1 gbuf_d_767(.A(n5704), .Y(ddout__767));
CLKBUFX1 gbuf_q_767(.A(qq_in767), .Y(n19020));
CLKBUFX1 gbuf_qn_767(.A(qnn_in_767), .Y(n17028));
CLKBUFX1 gbuf_d_768(.A(n5709), .Y(ddout__768));
CLKBUFX1 gbuf_q_768(.A(qq_in768), .Y(n19015));
CLKBUFX1 gbuf_qn_768(.A(qnn_in_768), .Y(n17038));
CLKBUFX1 gbuf_d_769(.A(n5713), .Y(ddout__769));
CLKBUFX1 gbuf_q_769(.A(qq_in769), .Y(n19011));
CLKBUFX1 gbuf_d_770(.A(n5714), .Y(ddout__770));
CLKBUFX1 gbuf_q_770(.A(qq_in770), .Y(n19010));
CLKBUFX1 gbuf_d_771(.A(n5712), .Y(ddout__771));
CLKBUFX1 gbuf_q_771(.A(qq_in771), .Y(n19012));
CLKBUFX1 gbuf_d_772(.A(n5717), .Y(ddout__772));
CLKBUFX1 gbuf_q_772(.A(qq_in772), .Y(n19007));
CLKBUFX1 gbuf_d_773(.A(n5710), .Y(ddout__773));
CLKBUFX1 gbuf_q_773(.A(qq_in773), .Y(n19014));
CLKBUFX1 gbuf_d_774(.A(n5715), .Y(ddout__774));
CLKBUFX1 gbuf_q_774(.A(qq_in774), .Y(n19009));
CLKBUFX1 gbuf_d_775(.A(n5711), .Y(ddout__775));
CLKBUFX1 gbuf_q_775(.A(qq_in775), .Y(n19013));
CLKBUFX1 gbuf_d_776(.A(n5716), .Y(ddout__776));
CLKBUFX1 gbuf_q_776(.A(qq_in776), .Y(n19008));
CLKBUFX1 gbuf_d_777(.A(n17280), .Y(ddout__777));
CLKBUFX1 gbuf_q_777(.A(qq_in777), .Y(n18622));
CLKBUFX1 gbuf_qn_777(.A(qnn_in_777), .Y(n6859));
CLKBUFX1 gbuf_d_778(.A(n6291), .Y(ddout__778));
CLKBUFX1 gbuf_q_778(.A(qq_in778), .Y(n18624));
CLKBUFX1 gbuf_qn_778(.A(qnn_in_778), .Y(n6850));
CLKBUFX1 gbuf_d_779(.A(n6290), .Y(ddout__779));
CLKBUFX1 gbuf_q_779(.A(qq_in779), .Y(n18893));
CLKBUFX1 gbuf_qn_779(.A(qnn_in_779), .Y(n16838));
OR3_X4 U13738 ( .A1(n17281), .A2(n17837), .A3(n17996), .ZN(n17282) );
NOR4_X2 U13739 ( .A1(n18079), .A2(n16837), .A3(state[7]), .A4(state[9]),.ZN(n17283) );
OR2_X4 U13740 ( .A1(n11946), .A2(n16542), .ZN(n17284) );
OR2_X4 U13741 ( .A1(n17281), .A2(n17841), .ZN(n17285) );
OR2_X4 U13742 ( .A1(cii_ctl_vld), .A2(n17958), .ZN(n17286) );
NAND3_X2 U13743 ( .A1(dii_data_vld), .A2(n18617), .A3(n18081), .ZN(n18085));
OR2_X4 U13744 ( .A1(n19204), .A2(dii_data_size[0]), .ZN(n17287) );
NOR2_X2 U13745 ( .A1(n19203), .A2(n18744), .ZN(n17288) );
OR2_X4 U13746 ( .A1(n18892), .A2(cii_ctl_vld), .ZN(n17289) );
AND2_X4 U13747 ( .A1(n12235), .A2(state[3]), .ZN(n17290) );
AND2_X4 U13748 ( .A1(n18623), .A2(n18622), .ZN(n17291) );
AND2_X4 U13749 ( .A1(n18619), .A2(n18618), .ZN(n17375) );
BUF_X32 U13750 ( .A(cii_K[64]), .Z(n17376) );
BUF_X32 U13751 ( .A(cii_K[32]), .Z(n17377) );
BUF_X32 U13752 ( .A(cii_K[79]), .Z(n17378) );
BUF_X32 U13753 ( .A(cii_K[47]), .Z(n17379) );
BUF_X32 U13754 ( .A(cii_K[87]), .Z(n17380) );
BUF_X32 U13755 ( .A(cii_K[55]), .Z(n17381) );
BUF_X32 U13756 ( .A(cii_K[95]), .Z(n17382) );
BUF_X32 U13757 ( .A(cii_K[63]), .Z(n17383) );
BUF_X32 U13758 ( .A(cii_K[71]), .Z(n17384) );
BUF_X32 U13759 ( .A(cii_K[39]), .Z(n17385) );
BUF_X32 U13760 ( .A(cii_K[7]), .Z(n17386) );
BUF_X32 U13761 ( .A(cii_K[103]), .Z(n17387) );
BUF_X32 U13762 ( .A(cii_K[70]), .Z(n17388) );
BUF_X32 U13763 ( .A(cii_K[38]), .Z(n17389) );
BUF_X32 U13764 ( .A(cii_K[6]), .Z(n17390) );
BUF_X32 U13765 ( .A(cii_K[102]), .Z(n17391) );
BUF_X32 U13766 ( .A(cii_K[69]), .Z(n17392) );
BUF_X32 U13767 ( .A(cii_K[37]), .Z(n17393) );
BUF_X32 U13768 ( .A(cii_K[5]), .Z(n17394) );
BUF_X32 U13769 ( .A(cii_K[101]), .Z(n17395) );
BUF_X32 U13770 ( .A(cii_K[68]), .Z(n17396) );
BUF_X32 U13771 ( .A(cii_K[36]), .Z(n17397) );
BUF_X32 U13772 ( .A(cii_K[4]), .Z(n17398) );
BUF_X32 U13773 ( .A(cii_K[100]), .Z(n17399) );
BUF_X32 U13774 ( .A(cii_K[67]), .Z(n17400) );
BUF_X32 U13775 ( .A(cii_K[35]), .Z(n17401) );
BUF_X32 U13776 ( .A(cii_K[3]), .Z(n17402) );
BUF_X32 U13777 ( .A(cii_K[99]), .Z(n17403) );
BUF_X32 U13778 ( .A(cii_K[66]), .Z(n17404) );
BUF_X32 U13779 ( .A(cii_K[34]), .Z(n17405) );
BUF_X32 U13780 ( .A(cii_K[2]), .Z(n17406) );
BUF_X32 U13781 ( .A(cii_K[98]), .Z(n17407) );
BUF_X32 U13782 ( .A(cii_K[65]), .Z(n17408) );
BUF_X32 U13783 ( .A(cii_K[33]), .Z(n17409) );
BUF_X32 U13784 ( .A(cii_K[1]), .Z(n17410) );
BUF_X32 U13785 ( .A(cii_K[97]), .Z(n17411) );
BUF_X32 U13786 ( .A(cii_K[31]), .Z(n17412) );
BUF_X32 U13787 ( .A(cii_K[126]), .Z(n17413) );
BUF_X32 U13788 ( .A(cii_K[94]), .Z(n17414) );
BUF_X32 U13789 ( .A(cii_K[62]), .Z(n17415) );
BUF_X32 U13790 ( .A(cii_K[30]), .Z(n17416) );
BUF_X32 U13791 ( .A(cii_K[125]), .Z(n17417) );
BUF_X32 U13792 ( .A(cii_K[93]), .Z(n17418) );
BUF_X32 U13793 ( .A(cii_K[61]), .Z(n17419) );
BUF_X32 U13794 ( .A(cii_K[29]), .Z(n17420) );
BUF_X32 U13795 ( .A(cii_K[124]), .Z(n17421) );
BUF_X32 U13796 ( .A(cii_K[92]), .Z(n17422) );
BUF_X32 U13797 ( .A(cii_K[60]), .Z(n17423) );
BUF_X32 U13798 ( .A(cii_K[28]), .Z(n17424) );
BUF_X32 U13799 ( .A(cii_K[123]), .Z(n17425) );
BUF_X32 U13800 ( .A(cii_K[91]), .Z(n17426) );
BUF_X32 U13801 ( .A(cii_K[59]), .Z(n17427) );
BUF_X32 U13802 ( .A(cii_K[27]), .Z(n17428) );
BUF_X32 U13803 ( .A(cii_K[122]), .Z(n17429) );
BUF_X32 U13804 ( .A(cii_K[90]), .Z(n17430) );
BUF_X32 U13805 ( .A(cii_K[58]), .Z(n17431) );
BUF_X32 U13806 ( .A(cii_K[26]), .Z(n17432) );
BUF_X32 U13807 ( .A(cii_K[121]), .Z(n17433) );
BUF_X32 U13808 ( .A(cii_K[89]), .Z(n17434) );
BUF_X32 U13809 ( .A(cii_K[57]), .Z(n17435) );
BUF_X32 U13810 ( .A(cii_K[25]), .Z(n17436) );
BUF_X32 U13811 ( .A(cii_K[120]), .Z(n17437) );
BUF_X32 U13812 ( .A(cii_K[88]), .Z(n17438) );
BUF_X32 U13813 ( .A(cii_K[56]), .Z(n17439) );
BUF_X32 U13814 ( .A(cii_K[24]), .Z(n17440) );
BUF_X32 U13815 ( .A(cii_K[23]), .Z(n17441) );
BUF_X32 U13816 ( .A(cii_K[119]), .Z(n17442) );
BUF_X32 U13817 ( .A(cii_K[86]), .Z(n17443) );
BUF_X32 U13818 ( .A(cii_K[54]), .Z(n17444) );
BUF_X32 U13819 ( .A(cii_K[22]), .Z(n17445) );
BUF_X32 U13820 ( .A(cii_K[118]), .Z(n17446) );
BUF_X32 U13821 ( .A(cii_K[85]), .Z(n17447) );
BUF_X32 U13822 ( .A(cii_K[53]), .Z(n17448) );
BUF_X32 U13823 ( .A(cii_K[21]), .Z(n17449) );
BUF_X32 U13824 ( .A(cii_K[117]), .Z(n17450) );
BUF_X32 U13825 ( .A(cii_K[84]), .Z(n17451) );
BUF_X32 U13826 ( .A(cii_K[52]), .Z(n17452) );
BUF_X32 U13827 ( .A(cii_K[20]), .Z(n17453) );
BUF_X32 U13828 ( .A(cii_K[116]), .Z(n17454) );
BUF_X32 U13829 ( .A(cii_K[83]), .Z(n17455) );
BUF_X32 U13830 ( .A(cii_K[51]), .Z(n17456) );
BUF_X32 U13831 ( .A(cii_K[19]), .Z(n17457) );
BUF_X32 U13832 ( .A(cii_K[115]), .Z(n17458) );
BUF_X32 U13833 ( .A(cii_K[82]), .Z(n17459) );
BUF_X32 U13834 ( .A(cii_K[50]), .Z(n17460) );
BUF_X32 U13835 ( .A(cii_K[18]), .Z(n17461) );
BUF_X32 U13836 ( .A(cii_K[114]), .Z(n17462) );
BUF_X32 U13837 ( .A(cii_K[81]), .Z(n17463) );
BUF_X32 U13838 ( .A(cii_K[49]), .Z(n17464) );
BUF_X32 U13839 ( .A(cii_K[17]), .Z(n17465) );
BUF_X32 U13840 ( .A(cii_K[113]), .Z(n17466) );
BUF_X32 U13841 ( .A(cii_K[80]), .Z(n17467) );
BUF_X32 U13842 ( .A(cii_K[48]), .Z(n17468) );
BUF_X32 U13843 ( .A(cii_K[16]), .Z(n17469) );
BUF_X32 U13844 ( .A(cii_K[112]), .Z(n17470) );
BUF_X32 U13845 ( .A(cii_K[15]), .Z(n17471) );
BUF_X32 U13846 ( .A(cii_K[111]), .Z(n17472) );
BUF_X32 U13847 ( .A(cii_K[78]), .Z(n17473) );
BUF_X32 U13848 ( .A(cii_K[46]), .Z(n17474) );
BUF_X32 U13849 ( .A(cii_K[14]), .Z(n17475) );
BUF_X32 U13850 ( .A(cii_K[110]), .Z(n17476) );
BUF_X32 U13851 ( .A(cii_K[77]), .Z(n17477) );
BUF_X32 U13852 ( .A(cii_K[45]), .Z(n17478) );
BUF_X32 U13853 ( .A(cii_K[13]), .Z(n17479) );
BUF_X32 U13854 ( .A(cii_K[109]), .Z(n17480) );
BUF_X32 U13855 ( .A(cii_K[76]), .Z(n17481) );
BUF_X32 U13856 ( .A(cii_K[44]), .Z(n17482) );
BUF_X32 U13857 ( .A(cii_K[12]), .Z(n17483) );
BUF_X32 U13858 ( .A(cii_K[108]), .Z(n17484) );
BUF_X32 U13859 ( .A(cii_K[75]), .Z(n17485) );
BUF_X32 U13860 ( .A(cii_K[43]), .Z(n17486) );
BUF_X32 U13861 ( .A(cii_K[11]), .Z(n17487) );
BUF_X32 U13862 ( .A(cii_K[107]), .Z(n17488) );
BUF_X32 U13863 ( .A(cii_K[74]), .Z(n17489) );
BUF_X32 U13864 ( .A(cii_K[42]), .Z(n17490) );
BUF_X32 U13865 ( .A(cii_K[10]), .Z(n17491) );
BUF_X32 U13866 ( .A(cii_K[106]), .Z(n17492) );
BUF_X32 U13867 ( .A(cii_K[73]), .Z(n17493) );
BUF_X32 U13868 ( .A(cii_K[41]), .Z(n17494) );
BUF_X32 U13869 ( .A(cii_K[9]), .Z(n17495) );
BUF_X32 U13870 ( .A(cii_K[105]), .Z(n17496) );
BUF_X32 U13871 ( .A(cii_K[72]), .Z(n17497) );
BUF_X32 U13872 ( .A(cii_K[40]), .Z(n17498) );
BUF_X32 U13873 ( .A(cii_K[8]), .Z(n17499) );
BUF_X32 U13874 ( .A(cii_K[104]), .Z(n17500) );
BUF_X32 U13875 ( .A(cii_K[0]), .Z(n17501) );
BUF_X32 U13876 ( .A(cii_K[96]), .Z(n17502) );
NAND2_X1 U13877 ( .A1(n17930), .A2(n13675), .ZN(n13671) );
XOR2_X1 U13878 ( .A(aes_text_out[65]), .B(n17629), .Z(n13668) );
NAND2_X1 U13879 ( .A1(n17924), .A2(n13661), .ZN(n13656) );
BUF_X32 U13880 ( .A(n6025), .Z(n17503) );
NAND2_X1 U13881 ( .A1(n12495), .A2(n12496), .ZN(n6025) );
NAND2_X1 U13882 ( .A1(dii_data_size[1]), .A2(n17281), .ZN(n12496) );
BUF_X32 U13883 ( .A(n6024), .Z(n17504) );
NAND2_X1 U13884 ( .A1(n12497), .A2(n12498), .ZN(n6024) );
NAND2_X1 U13885 ( .A1(dii_data_size[2]), .A2(n17281), .ZN(n12498) );
NOR3_X1 U13886 ( .A1(n18746), .A2(n11976), .A3(n18601), .ZN(n17281) );
CLKBUF_X2 U13887 ( .A(n17281), .Z(n17505) );
NAND3_X1 U13888 ( .A1(n18596), .A2(n17506), .A3(n18594), .ZN(n5830) );
BUF_X8 U13889 ( .A(n18595), .Z(n17506) );
CLKBUF_X2 U13890 ( .A(n5830), .Z(n17507) );
NAND2_X1 U13891 ( .A1(dii_data[127]), .A2(n17799), .ZN(n18595) );
NAND3_X1 U13892 ( .A1(n18088), .A2(n17508), .A3(n18086), .ZN(n5831) );
BUF_X8 U13893 ( .A(n18087), .Z(n17508) );
CLKBUF_X2 U13894 ( .A(n5831), .Z(n17509) );
NAND2_X1 U13895 ( .A1(dii_data[126]), .A2(n17788), .ZN(n18087) );
NAND3_X1 U13896 ( .A1(n18092), .A2(n17510), .A3(n18090), .ZN(n5832) );
BUF_X8 U13897 ( .A(n18091), .Z(n17510) );
CLKBUF_X2 U13898 ( .A(n5832), .Z(n17511) );
NAND2_X1 U13899 ( .A1(dii_data[125]), .A2(n17788), .ZN(n18091) );
NAND3_X1 U13900 ( .A1(n18096), .A2(n17512), .A3(n18094), .ZN(n5833) );
BUF_X8 U13901 ( .A(n18095), .Z(n17512) );
CLKBUF_X2 U13902 ( .A(n5833), .Z(n17513) );
NAND2_X1 U13903 ( .A1(dii_data[124]), .A2(n17788), .ZN(n18095) );
NAND3_X1 U13904 ( .A1(n18100), .A2(n17514), .A3(n18098), .ZN(n5834) );
BUF_X8 U13905 ( .A(n18099), .Z(n17514) );
CLKBUF_X2 U13906 ( .A(n5834), .Z(n17515) );
NAND2_X1 U13907 ( .A1(dii_data[123]), .A2(n17788), .ZN(n18099) );
NAND3_X1 U13908 ( .A1(n18104), .A2(n17516), .A3(n18102), .ZN(n5835) );
BUF_X8 U13909 ( .A(n18103), .Z(n17516) );
CLKBUF_X2 U13910 ( .A(n5835), .Z(n17517) );
NAND2_X1 U13911 ( .A1(dii_data[122]), .A2(n17788), .ZN(n18103) );
NAND3_X1 U13912 ( .A1(n18108), .A2(n17518), .A3(n18106), .ZN(n5836) );
BUF_X8 U13913 ( .A(n18107), .Z(n17518) );
CLKBUF_X2 U13914 ( .A(n5836), .Z(n17519) );
NAND2_X1 U13915 ( .A1(dii_data[121]), .A2(n17788), .ZN(n18107) );
NAND3_X1 U13916 ( .A1(n18112), .A2(n17520), .A3(n18110), .ZN(n5837) );
BUF_X8 U13917 ( .A(n18111), .Z(n17520) );
CLKBUF_X2 U13918 ( .A(n5837), .Z(n17521) );
NAND2_X1 U13919 ( .A1(dii_data[120]), .A2(n17788), .ZN(n18111) );
CLKBUF_X1 U13920 ( .A(dii_data[119]), .Z(n17523) );
CLKBUF_X2 U13921 ( .A(n17523), .Z(n17522) );
NAND2_X1 U13922 ( .A1(n17522), .A2(n17788), .ZN(n18115) );
CLKBUF_X1 U13923 ( .A(dii_data[118]), .Z(n17525) );
CLKBUF_X2 U13924 ( .A(n17525), .Z(n17524) );
NAND2_X1 U13925 ( .A1(n17524), .A2(n17788), .ZN(n18119) );
CLKBUF_X1 U13926 ( .A(dii_data[117]), .Z(n17527) );
CLKBUF_X2 U13927 ( .A(n17527), .Z(n17526) );
NAND2_X1 U13928 ( .A1(n17526), .A2(n17788), .ZN(n18123) );
CLKBUF_X1 U13929 ( .A(dii_data[116]), .Z(n17529) );
CLKBUF_X2 U13930 ( .A(n17529), .Z(n17528) );
NAND2_X1 U13931 ( .A1(n17528), .A2(n17788), .ZN(n18127) );
CLKBUF_X1 U13932 ( .A(dii_data[115]), .Z(n17531) );
CLKBUF_X2 U13933 ( .A(n17531), .Z(n17530) );
NAND2_X1 U13934 ( .A1(n17530), .A2(n17789), .ZN(n18131) );
CLKBUF_X1 U13935 ( .A(dii_data[114]), .Z(n17533) );
CLKBUF_X2 U13936 ( .A(n17533), .Z(n17532) );
NAND2_X1 U13937 ( .A1(n17532), .A2(n17789), .ZN(n18135) );
CLKBUF_X1 U13938 ( .A(dii_data[113]), .Z(n17535) );
CLKBUF_X2 U13939 ( .A(n17535), .Z(n17534) );
NAND2_X1 U13940 ( .A1(n17534), .A2(n17789), .ZN(n18139) );
CLKBUF_X1 U13941 ( .A(dii_data[112]), .Z(n17537) );
CLKBUF_X2 U13942 ( .A(n17537), .Z(n17536) );
NAND2_X1 U13943 ( .A1(n17536), .A2(n17789), .ZN(n18143) );
NAND3_X1 U13944 ( .A1(n18148), .A2(n18147), .A3(n18146), .ZN(n5846) );
CLKBUF_X2 U13945 ( .A(n5846), .Z(n17538) );
CLKBUF_X2 U13946 ( .A(dii_data[111]), .Z(n17539) );
NAND2_X1 U13947 ( .A1(n17539), .A2(n17789), .ZN(n18147) );
NAND3_X1 U13948 ( .A1(n18152), .A2(n18151), .A3(n18150), .ZN(n5847) );
CLKBUF_X2 U13949 ( .A(n5847), .Z(n17540) );
CLKBUF_X2 U13950 ( .A(dii_data[110]), .Z(n17541) );
NAND2_X1 U13951 ( .A1(n17541), .A2(n17789), .ZN(n18151) );
NAND3_X1 U13952 ( .A1(n18156), .A2(n18155), .A3(n18154), .ZN(n5848) );
CLKBUF_X2 U13953 ( .A(n5848), .Z(n17542) );
CLKBUF_X2 U13954 ( .A(dii_data[109]), .Z(n17543) );
NAND2_X1 U13955 ( .A1(n17543), .A2(n17789), .ZN(n18155) );
NAND3_X1 U13956 ( .A1(n18160), .A2(n18159), .A3(n18158), .ZN(n5849) );
CLKBUF_X2 U13957 ( .A(n5849), .Z(n17544) );
CLKBUF_X2 U13958 ( .A(dii_data[108]), .Z(n17545) );
NAND2_X1 U13959 ( .A1(n17545), .A2(n17789), .ZN(n18159) );
NAND3_X1 U13960 ( .A1(n18164), .A2(n18163), .A3(n18162), .ZN(n5850) );
CLKBUF_X2 U13961 ( .A(n5850), .Z(n17546) );
CLKBUF_X2 U13962 ( .A(dii_data[107]), .Z(n17547) );
NAND2_X1 U13963 ( .A1(n17547), .A2(n17789), .ZN(n18163) );
NAND3_X1 U13964 ( .A1(n18168), .A2(n18167), .A3(n18166), .ZN(n5851) );
CLKBUF_X2 U13965 ( .A(n5851), .Z(n17548) );
CLKBUF_X2 U13966 ( .A(dii_data[106]), .Z(n17549) );
NAND2_X1 U13967 ( .A1(n17549), .A2(n17789), .ZN(n18167) );
NAND3_X1 U13968 ( .A1(n18172), .A2(n18171), .A3(n18170), .ZN(n5852) );
CLKBUF_X2 U13969 ( .A(n5852), .Z(n17550) );
CLKBUF_X2 U13970 ( .A(dii_data[105]), .Z(n17551) );
NAND2_X1 U13971 ( .A1(n17551), .A2(n17789), .ZN(n18171) );
NAND3_X1 U13972 ( .A1(n18176), .A2(n18175), .A3(n18174), .ZN(n5853) );
CLKBUF_X2 U13973 ( .A(n5853), .Z(n17552) );
CLKBUF_X2 U13974 ( .A(dii_data[104]), .Z(n17553) );
NAND2_X1 U13975 ( .A1(n17553), .A2(n17790), .ZN(n18175) );
NAND3_X1 U13976 ( .A1(n18180), .A2(n18179), .A3(n18178), .ZN(n5854) );
CLKBUF_X2 U13977 ( .A(n5854), .Z(n17554) );
CLKBUF_X2 U13978 ( .A(dii_data[103]), .Z(n17555) );
NAND2_X1 U13979 ( .A1(n17555), .A2(n17790), .ZN(n18179) );
NAND3_X1 U13980 ( .A1(n18184), .A2(n18183), .A3(n18182), .ZN(n5855) );
CLKBUF_X2 U13981 ( .A(n5855), .Z(n17556) );
CLKBUF_X2 U13982 ( .A(dii_data[102]), .Z(n17557) );
NAND2_X1 U13983 ( .A1(n17557), .A2(n17790), .ZN(n18183) );
NAND3_X1 U13984 ( .A1(n18188), .A2(n18187), .A3(n18186), .ZN(n5856) );
CLKBUF_X2 U13985 ( .A(n5856), .Z(n17558) );
CLKBUF_X2 U13986 ( .A(dii_data[101]), .Z(n17559) );
NAND2_X1 U13987 ( .A1(n17559), .A2(n17790), .ZN(n18187) );
NAND3_X1 U13988 ( .A1(n18192), .A2(n18191), .A3(n18190), .ZN(n5857) );
CLKBUF_X2 U13989 ( .A(n5857), .Z(n17560) );
CLKBUF_X2 U13990 ( .A(dii_data[100]), .Z(n17561) );
NAND2_X1 U13991 ( .A1(n17561), .A2(n17790), .ZN(n18191) );
NAND3_X1 U13992 ( .A1(n18196), .A2(n18195), .A3(n18194), .ZN(n5858) );
CLKBUF_X2 U13993 ( .A(n5858), .Z(n17562) );
CLKBUF_X2 U13994 ( .A(dii_data[99]), .Z(n17563) );
NAND2_X1 U13995 ( .A1(n17563), .A2(n17790), .ZN(n18195) );
NAND3_X1 U13996 ( .A1(n18204), .A2(n18203), .A3(n18202), .ZN(n5859) );
CLKBUF_X2 U13997 ( .A(n5859), .Z(n17564) );
CLKBUF_X2 U13998 ( .A(dii_data[97]), .Z(n17565) );
NAND2_X1 U13999 ( .A1(n17565), .A2(n17790), .ZN(n18203) );
NAND3_X1 U14000 ( .A1(n18208), .A2(n18207), .A3(n18206), .ZN(n5860) );
CLKBUF_X2 U14001 ( .A(n5860), .Z(n17566) );
CLKBUF_X2 U14002 ( .A(dii_data[96]), .Z(n17567) );
NAND2_X1 U14003 ( .A1(n17567), .A2(n17790), .ZN(n18207) );
NAND3_X1 U14004 ( .A1(n18212), .A2(n18211), .A3(n18210), .ZN(n5861) );
CLKBUF_X2 U14005 ( .A(n5861), .Z(n17568) );
CLKBUF_X2 U14006 ( .A(dii_data[95]), .Z(n17569) );
NAND2_X1 U14007 ( .A1(n17569), .A2(n17790), .ZN(n18211) );
NAND3_X1 U14008 ( .A1(n18216), .A2(n18215), .A3(n18214), .ZN(n5862) );
CLKBUF_X2 U14009 ( .A(n5862), .Z(n17570) );
CLKBUF_X2 U14010 ( .A(dii_data[94]), .Z(n17571) );
NAND2_X1 U14011 ( .A1(n17571), .A2(n17790), .ZN(n18215) );
NAND3_X1 U14012 ( .A1(n18220), .A2(n18219), .A3(n18218), .ZN(n5863) );
CLKBUF_X2 U14013 ( .A(n5863), .Z(n17572) );
CLKBUF_X2 U14014 ( .A(dii_data[93]), .Z(n17573) );
NAND2_X1 U14015 ( .A1(n17573), .A2(n17791), .ZN(n18219) );
NAND3_X1 U14016 ( .A1(n18224), .A2(n18223), .A3(n18222), .ZN(n5864) );
CLKBUF_X2 U14017 ( .A(n5864), .Z(n17574) );
CLKBUF_X2 U14018 ( .A(dii_data[92]), .Z(n17575) );
NAND2_X1 U14019 ( .A1(n17575), .A2(n17791), .ZN(n18223) );
NAND3_X1 U14020 ( .A1(n18228), .A2(n18227), .A3(n18226), .ZN(n5865) );
CLKBUF_X2 U14021 ( .A(n5865), .Z(n17576) );
CLKBUF_X2 U14022 ( .A(dii_data[91]), .Z(n17577) );
NAND2_X1 U14023 ( .A1(n17577), .A2(n17791), .ZN(n18227) );
NAND3_X1 U14024 ( .A1(n18232), .A2(n18231), .A3(n18230), .ZN(n5866) );
CLKBUF_X2 U14025 ( .A(n5866), .Z(n17578) );
CLKBUF_X2 U14026 ( .A(dii_data[90]), .Z(n17579) );
NAND2_X1 U14027 ( .A1(n17579), .A2(n17791), .ZN(n18231) );
NAND3_X1 U14028 ( .A1(n18236), .A2(n18235), .A3(n18234), .ZN(n5867) );
CLKBUF_X2 U14029 ( .A(n5867), .Z(n17580) );
CLKBUF_X2 U14030 ( .A(dii_data[89]), .Z(n17581) );
NAND2_X1 U14031 ( .A1(n17581), .A2(n17791), .ZN(n18235) );
NAND3_X1 U14032 ( .A1(n18240), .A2(n18239), .A3(n18238), .ZN(n5868) );
CLKBUF_X2 U14033 ( .A(n5868), .Z(n17582) );
CLKBUF_X2 U14034 ( .A(dii_data[88]), .Z(n17583) );
NAND2_X1 U14035 ( .A1(n17583), .A2(n17791), .ZN(n18239) );
NAND3_X1 U14036 ( .A1(n18244), .A2(n18243), .A3(n18242), .ZN(n5869) );
CLKBUF_X2 U14037 ( .A(n5869), .Z(n17584) );
CLKBUF_X2 U14038 ( .A(dii_data[87]), .Z(n17585) );
NAND2_X1 U14039 ( .A1(n17585), .A2(n17791), .ZN(n18243) );
NAND3_X1 U14040 ( .A1(n18248), .A2(n18247), .A3(n18246), .ZN(n5870) );
CLKBUF_X2 U14041 ( .A(n5870), .Z(n17586) );
CLKBUF_X2 U14042 ( .A(dii_data[86]), .Z(n17587) );
NAND2_X1 U14043 ( .A1(n17587), .A2(n17791), .ZN(n18247) );
NAND3_X1 U14044 ( .A1(n18252), .A2(n18251), .A3(n18250), .ZN(n5871) );
CLKBUF_X2 U14045 ( .A(n5871), .Z(n17588) );
CLKBUF_X2 U14046 ( .A(dii_data[85]), .Z(n17589) );
NAND2_X1 U14047 ( .A1(n17589), .A2(n17791), .ZN(n18251) );
NAND3_X1 U14048 ( .A1(n18256), .A2(n18255), .A3(n18254), .ZN(n5872) );
CLKBUF_X2 U14049 ( .A(n5872), .Z(n17590) );
CLKBUF_X2 U14050 ( .A(dii_data[84]), .Z(n17591) );
NAND2_X1 U14051 ( .A1(n17591), .A2(n17791), .ZN(n18255) );
NAND3_X1 U14052 ( .A1(n18260), .A2(n18259), .A3(n18258), .ZN(n5873) );
CLKBUF_X2 U14053 ( .A(n5873), .Z(n17592) );
CLKBUF_X2 U14054 ( .A(dii_data[83]), .Z(n17593) );
NAND2_X1 U14055 ( .A1(n17593), .A2(n17791), .ZN(n18259) );
NAND3_X1 U14056 ( .A1(n18264), .A2(n18263), .A3(n18262), .ZN(n5874) );
CLKBUF_X2 U14057 ( .A(n5874), .Z(n17594) );
CLKBUF_X2 U14058 ( .A(dii_data[82]), .Z(n17595) );
NAND2_X1 U14059 ( .A1(n17595), .A2(n17792), .ZN(n18263) );
NAND3_X1 U14060 ( .A1(n18268), .A2(n18267), .A3(n18266), .ZN(n5875) );
CLKBUF_X2 U14061 ( .A(n5875), .Z(n17596) );
CLKBUF_X2 U14062 ( .A(dii_data[81]), .Z(n17597) );
NAND2_X1 U14063 ( .A1(n17597), .A2(n17792), .ZN(n18267) );
NAND3_X1 U14064 ( .A1(n18272), .A2(n18271), .A3(n18270), .ZN(n5876) );
CLKBUF_X2 U14065 ( .A(n5876), .Z(n17598) );
CLKBUF_X2 U14066 ( .A(dii_data[80]), .Z(n17599) );
NAND2_X1 U14067 ( .A1(n17599), .A2(n17792), .ZN(n18271) );
NAND3_X1 U14068 ( .A1(n18276), .A2(n18275), .A3(n18274), .ZN(n5877) );
CLKBUF_X2 U14069 ( .A(n5877), .Z(n17600) );
CLKBUF_X2 U14070 ( .A(dii_data[79]), .Z(n17601) );
NAND2_X1 U14071 ( .A1(n17601), .A2(n17792), .ZN(n18275) );
NAND3_X1 U14072 ( .A1(n18280), .A2(n18279), .A3(n18278), .ZN(n5878) );
CLKBUF_X2 U14073 ( .A(n5878), .Z(n17602) );
CLKBUF_X2 U14074 ( .A(dii_data[78]), .Z(n17603) );
NAND2_X1 U14075 ( .A1(n17603), .A2(n17792), .ZN(n18279) );
NAND3_X1 U14076 ( .A1(n18284), .A2(n18283), .A3(n18282), .ZN(n5879) );
CLKBUF_X2 U14077 ( .A(n5879), .Z(n17604) );
CLKBUF_X2 U14078 ( .A(dii_data[77]), .Z(n17605) );
NAND2_X1 U14079 ( .A1(n17605), .A2(n17792), .ZN(n18283) );
NAND3_X1 U14080 ( .A1(n18288), .A2(n18287), .A3(n18286), .ZN(n5880) );
CLKBUF_X2 U14081 ( .A(n5880), .Z(n17606) );
CLKBUF_X2 U14082 ( .A(dii_data[76]), .Z(n17607) );
NAND2_X1 U14083 ( .A1(n17607), .A2(n17792), .ZN(n18287) );
NAND3_X1 U14084 ( .A1(n18292), .A2(n18291), .A3(n18290), .ZN(n5881) );
CLKBUF_X2 U14085 ( .A(n5881), .Z(n17608) );
CLKBUF_X2 U14086 ( .A(dii_data[75]), .Z(n17609) );
NAND2_X1 U14087 ( .A1(n17609), .A2(n17792), .ZN(n18291) );
NAND3_X1 U14088 ( .A1(n18296), .A2(n18295), .A3(n18294), .ZN(n5882) );
CLKBUF_X2 U14089 ( .A(n5882), .Z(n17610) );
CLKBUF_X2 U14090 ( .A(dii_data[74]), .Z(n17611) );
NAND2_X1 U14091 ( .A1(n17611), .A2(n17792), .ZN(n18295) );
NAND3_X1 U14092 ( .A1(n18300), .A2(n18299), .A3(n18298), .ZN(n5883) );
CLKBUF_X2 U14093 ( .A(n5883), .Z(n17612) );
CLKBUF_X2 U14094 ( .A(dii_data[73]), .Z(n17613) );
NAND2_X1 U14095 ( .A1(n17613), .A2(n17792), .ZN(n18299) );
NAND3_X1 U14096 ( .A1(n18304), .A2(n18303), .A3(n18302), .ZN(n5884) );
CLKBUF_X2 U14097 ( .A(n5884), .Z(n17614) );
CLKBUF_X2 U14098 ( .A(dii_data[72]), .Z(n17615) );
NAND2_X1 U14099 ( .A1(n17615), .A2(n17792), .ZN(n18303) );
CLKBUF_X1 U14100 ( .A(dii_data[71]), .Z(n17617) );
CLKBUF_X2 U14101 ( .A(n17617), .Z(n17616) );
NAND2_X1 U14102 ( .A1(n17616), .A2(n17793), .ZN(n18307) );
CLKBUF_X1 U14103 ( .A(dii_data[70]), .Z(n17619) );
CLKBUF_X2 U14104 ( .A(n17619), .Z(n17618) );
NAND2_X1 U14105 ( .A1(n17618), .A2(n17793), .ZN(n18311) );
CLKBUF_X1 U14106 ( .A(dii_data[69]), .Z(n17621) );
CLKBUF_X2 U14107 ( .A(n17621), .Z(n17620) );
NAND2_X1 U14108 ( .A1(n17620), .A2(n17793), .ZN(n18315) );
CLKBUF_X1 U14109 ( .A(dii_data[68]), .Z(n17623) );
CLKBUF_X2 U14110 ( .A(n17623), .Z(n17622) );
NAND2_X1 U14111 ( .A1(n17622), .A2(n17793), .ZN(n18319) );
CLKBUF_X1 U14112 ( .A(dii_data[67]), .Z(n17625) );
CLKBUF_X2 U14113 ( .A(n17625), .Z(n17624) );
NAND2_X1 U14114 ( .A1(n17624), .A2(n17793), .ZN(n18323) );
CLKBUF_X1 U14115 ( .A(n5890), .Z(n17626) );
NAND3_X1 U14116 ( .A1(n18328), .A2(n18327), .A3(n18326), .ZN(n5890) );
CLKBUF_X2 U14117 ( .A(dii_data[66]), .Z(n17627) );
NAND2_X1 U14118 ( .A1(n17627), .A2(n17793), .ZN(n18327) );
CLKBUF_X1 U14119 ( .A(n5891), .Z(n17628) );
NAND3_X1 U14120 ( .A1(n18332), .A2(n18331), .A3(n18330), .ZN(n5891) );
CLKBUF_X2 U14121 ( .A(dii_data[65]), .Z(n17629) );
NAND2_X1 U14122 ( .A1(n17629), .A2(n17793), .ZN(n18331) );
CLKBUF_X1 U14123 ( .A(n5892), .Z(n17630) );
NAND3_X1 U14124 ( .A1(n18336), .A2(n18335), .A3(n18334), .ZN(n5892) );
CLKBUF_X2 U14125 ( .A(dii_data[64]), .Z(n17631) );
NAND2_X1 U14126 ( .A1(n17631), .A2(n17793), .ZN(n18335) );
NAND3_X1 U14127 ( .A1(n18340), .A2(n18339), .A3(n18338), .ZN(n5893) );
CLKBUF_X2 U14128 ( .A(n5893), .Z(n17632) );
CLKBUF_X2 U14129 ( .A(dii_data[63]), .Z(n17633) );
NAND2_X1 U14130 ( .A1(n17633), .A2(n17793), .ZN(n18339) );
NAND3_X1 U14131 ( .A1(n18344), .A2(n18343), .A3(n18342), .ZN(n5894) );
CLKBUF_X2 U14132 ( .A(n5894), .Z(n17634) );
CLKBUF_X2 U14133 ( .A(dii_data[62]), .Z(n17635) );
NAND2_X1 U14134 ( .A1(n17635), .A2(n17793), .ZN(n18343) );
NAND3_X1 U14135 ( .A1(n18348), .A2(n18347), .A3(n18346), .ZN(n5895) );
CLKBUF_X2 U14136 ( .A(n5895), .Z(n17636) );
CLKBUF_X2 U14137 ( .A(dii_data[61]), .Z(n17637) );
NAND2_X1 U14138 ( .A1(n17637), .A2(n17793), .ZN(n18347) );
NAND3_X1 U14139 ( .A1(n18352), .A2(n18351), .A3(n18350), .ZN(n5896) );
CLKBUF_X2 U14140 ( .A(n5896), .Z(n17638) );
CLKBUF_X2 U14141 ( .A(dii_data[60]), .Z(n17639) );
NAND2_X1 U14142 ( .A1(n17639), .A2(n17794), .ZN(n18351) );
NAND3_X1 U14143 ( .A1(n18356), .A2(n18355), .A3(n18354), .ZN(n5897) );
CLKBUF_X2 U14144 ( .A(n5897), .Z(n17640) );
CLKBUF_X2 U14145 ( .A(dii_data[59]), .Z(n17641) );
NAND2_X1 U14146 ( .A1(n17641), .A2(n17794), .ZN(n18355) );
NAND3_X1 U14147 ( .A1(n18360), .A2(n18359), .A3(n18358), .ZN(n5898) );
CLKBUF_X2 U14148 ( .A(n5898), .Z(n17642) );
CLKBUF_X2 U14149 ( .A(dii_data[58]), .Z(n17643) );
NAND2_X1 U14150 ( .A1(n17643), .A2(n17794), .ZN(n18359) );
NAND3_X1 U14151 ( .A1(n18364), .A2(n18363), .A3(n18362), .ZN(n5899) );
CLKBUF_X2 U14152 ( .A(n5899), .Z(n17644) );
CLKBUF_X2 U14153 ( .A(dii_data[57]), .Z(n17645) );
NAND2_X1 U14154 ( .A1(n17645), .A2(n17794), .ZN(n18363) );
NAND3_X1 U14155 ( .A1(n18368), .A2(n18367), .A3(n18366), .ZN(n5900) );
CLKBUF_X2 U14156 ( .A(n5900), .Z(n17646) );
CLKBUF_X2 U14157 ( .A(dii_data[56]), .Z(n17647) );
NAND2_X1 U14158 ( .A1(n17647), .A2(n17794), .ZN(n18367) );
NAND3_X1 U14159 ( .A1(n18372), .A2(n18371), .A3(n18370), .ZN(n5901) );
CLKBUF_X2 U14160 ( .A(n5901), .Z(n17648) );
CLKBUF_X2 U14161 ( .A(dii_data[55]), .Z(n17649) );
NAND2_X1 U14162 ( .A1(n17649), .A2(n17794), .ZN(n18371) );
NAND3_X1 U14163 ( .A1(n18376), .A2(n18375), .A3(n18374), .ZN(n5902) );
CLKBUF_X2 U14164 ( .A(n5902), .Z(n17650) );
CLKBUF_X2 U14165 ( .A(dii_data[54]), .Z(n17651) );
NAND2_X1 U14166 ( .A1(n17651), .A2(n17794), .ZN(n18375) );
NAND3_X1 U14167 ( .A1(n18380), .A2(n18379), .A3(n18378), .ZN(n5903) );
CLKBUF_X2 U14168 ( .A(n5903), .Z(n17652) );
CLKBUF_X2 U14169 ( .A(dii_data[53]), .Z(n17653) );
NAND2_X1 U14170 ( .A1(n17653), .A2(n17794), .ZN(n18379) );
NAND3_X1 U14171 ( .A1(n18384), .A2(n18383), .A3(n18382), .ZN(n5904) );
CLKBUF_X2 U14172 ( .A(n5904), .Z(n17654) );
CLKBUF_X2 U14173 ( .A(dii_data[52]), .Z(n17655) );
NAND2_X1 U14174 ( .A1(n17655), .A2(n17794), .ZN(n18383) );
NAND3_X1 U14175 ( .A1(n18388), .A2(n18387), .A3(n18386), .ZN(n5905) );
CLKBUF_X2 U14176 ( .A(n5905), .Z(n17656) );
CLKBUF_X2 U14177 ( .A(dii_data[51]), .Z(n17657) );
NAND2_X1 U14178 ( .A1(n17657), .A2(n17794), .ZN(n18387) );
NAND3_X1 U14179 ( .A1(n18392), .A2(n18391), .A3(n18390), .ZN(n5906) );
CLKBUF_X2 U14180 ( .A(n5906), .Z(n17658) );
CLKBUF_X2 U14181 ( .A(dii_data[50]), .Z(n17659) );
NAND2_X1 U14182 ( .A1(n17659), .A2(n17794), .ZN(n18391) );
NAND3_X1 U14183 ( .A1(n18396), .A2(n18395), .A3(n18394), .ZN(n5907) );
CLKBUF_X2 U14184 ( .A(n5907), .Z(n17660) );
CLKBUF_X2 U14185 ( .A(dii_data[49]), .Z(n17661) );
NAND2_X1 U14186 ( .A1(n17661), .A2(n17795), .ZN(n18395) );
NAND3_X1 U14187 ( .A1(n18400), .A2(n18399), .A3(n18398), .ZN(n5908) );
CLKBUF_X2 U14188 ( .A(n5908), .Z(n17662) );
CLKBUF_X2 U14189 ( .A(dii_data[48]), .Z(n17663) );
NAND2_X1 U14190 ( .A1(n17663), .A2(n17795), .ZN(n18399) );
NAND3_X1 U14191 ( .A1(n18404), .A2(n18403), .A3(n18402), .ZN(n5909) );
CLKBUF_X2 U14192 ( .A(n5909), .Z(n17664) );
CLKBUF_X2 U14193 ( .A(dii_data[47]), .Z(n17665) );
NAND2_X1 U14194 ( .A1(n17665), .A2(n17795), .ZN(n18403) );
NAND3_X1 U14195 ( .A1(n18408), .A2(n18407), .A3(n18406), .ZN(n5910) );
CLKBUF_X2 U14196 ( .A(n5910), .Z(n17666) );
CLKBUF_X2 U14197 ( .A(dii_data[46]), .Z(n17667) );
NAND2_X1 U14198 ( .A1(n17667), .A2(n17795), .ZN(n18407) );
NAND3_X1 U14199 ( .A1(n18412), .A2(n18411), .A3(n18410), .ZN(n5911) );
CLKBUF_X2 U14200 ( .A(n5911), .Z(n17668) );
CLKBUF_X2 U14201 ( .A(dii_data[45]), .Z(n17669) );
NAND2_X1 U14202 ( .A1(n17669), .A2(n17795), .ZN(n18411) );
NAND3_X1 U14203 ( .A1(n18416), .A2(n18415), .A3(n18414), .ZN(n5912) );
CLKBUF_X2 U14204 ( .A(n5912), .Z(n17670) );
CLKBUF_X2 U14205 ( .A(dii_data[44]), .Z(n17671) );
NAND2_X1 U14206 ( .A1(n17671), .A2(n17795), .ZN(n18415) );
NAND3_X1 U14207 ( .A1(n18420), .A2(n18419), .A3(n18418), .ZN(n5913) );
CLKBUF_X2 U14208 ( .A(n5913), .Z(n17672) );
CLKBUF_X2 U14209 ( .A(dii_data[43]), .Z(n17673) );
NAND2_X1 U14210 ( .A1(n17673), .A2(n17795), .ZN(n18419) );
NAND3_X1 U14211 ( .A1(n18424), .A2(n18423), .A3(n18422), .ZN(n5914) );
CLKBUF_X2 U14212 ( .A(n5914), .Z(n17674) );
CLKBUF_X2 U14213 ( .A(dii_data[42]), .Z(n17675) );
NAND2_X1 U14214 ( .A1(n17675), .A2(n17795), .ZN(n18423) );
NAND3_X1 U14215 ( .A1(n18428), .A2(n18427), .A3(n18426), .ZN(n5915) );
CLKBUF_X2 U14216 ( .A(n5915), .Z(n17676) );
CLKBUF_X2 U14217 ( .A(dii_data[41]), .Z(n17677) );
NAND2_X1 U14218 ( .A1(n17677), .A2(n17795), .ZN(n18427) );
NAND3_X1 U14219 ( .A1(n18432), .A2(n18431), .A3(n18430), .ZN(n5916) );
CLKBUF_X2 U14220 ( .A(n5916), .Z(n17678) );
CLKBUF_X2 U14221 ( .A(dii_data[40]), .Z(n17679) );
NAND2_X1 U14222 ( .A1(n17679), .A2(n17795), .ZN(n18431) );
CLKBUF_X2 U14223 ( .A(n5917), .Z(n17680) );
CLKBUF_X2 U14224 ( .A(dii_data[39]), .Z(n17681) );
NAND2_X1 U14225 ( .A1(n17681), .A2(n17795), .ZN(n18435) );
CLKBUF_X2 U14226 ( .A(n5918), .Z(n17682) );
CLKBUF_X2 U14227 ( .A(dii_data[38]), .Z(n17683) );
NAND2_X1 U14228 ( .A1(n17683), .A2(n17796), .ZN(n18439) );
CLKBUF_X2 U14229 ( .A(n5919), .Z(n17684) );
CLKBUF_X2 U14230 ( .A(dii_data[37]), .Z(n17685) );
NAND2_X1 U14231 ( .A1(n17685), .A2(n17796), .ZN(n18443) );
CLKBUF_X2 U14232 ( .A(n5920), .Z(n17686) );
CLKBUF_X2 U14233 ( .A(dii_data[36]), .Z(n17687) );
NAND2_X1 U14234 ( .A1(n17687), .A2(n17796), .ZN(n18447) );
CLKBUF_X2 U14235 ( .A(n5921), .Z(n17688) );
CLKBUF_X2 U14236 ( .A(dii_data[35]), .Z(n17689) );
NAND2_X1 U14237 ( .A1(n17689), .A2(n17796), .ZN(n18451) );
CLKBUF_X2 U14238 ( .A(n5922), .Z(n17690) );
CLKBUF_X2 U14239 ( .A(dii_data[34]), .Z(n17691) );
NAND2_X1 U14240 ( .A1(n17691), .A2(n17796), .ZN(n18455) );
CLKBUF_X2 U14241 ( .A(n5923), .Z(n17692) );
CLKBUF_X2 U14242 ( .A(dii_data[33]), .Z(n17693) );
NAND2_X1 U14243 ( .A1(n17693), .A2(n17796), .ZN(n18459) );
CLKBUF_X2 U14244 ( .A(n5924), .Z(n17694) );
CLKBUF_X2 U14245 ( .A(dii_data[32]), .Z(n17695) );
NAND2_X1 U14246 ( .A1(n17695), .A2(n17796), .ZN(n18463) );
CLKBUF_X2 U14247 ( .A(n5925), .Z(n17696) );
CLKBUF_X2 U14248 ( .A(dii_data[31]), .Z(n17697) );
NAND2_X1 U14249 ( .A1(n17697), .A2(n17796), .ZN(n18467) );
CLKBUF_X2 U14250 ( .A(n5926), .Z(n17698) );
CLKBUF_X2 U14251 ( .A(dii_data[30]), .Z(n17699) );
NAND2_X1 U14252 ( .A1(n17699), .A2(n17796), .ZN(n18471) );
CLKBUF_X2 U14253 ( .A(n5927), .Z(n17700) );
CLKBUF_X2 U14254 ( .A(dii_data[29]), .Z(n17701) );
NAND2_X1 U14255 ( .A1(n17701), .A2(n17796), .ZN(n18475) );
CLKBUF_X2 U14256 ( .A(n5928), .Z(n17702) );
CLKBUF_X2 U14257 ( .A(dii_data[28]), .Z(n17703) );
NAND2_X1 U14258 ( .A1(n17703), .A2(n17796), .ZN(n18479) );
CLKBUF_X2 U14259 ( .A(n5929), .Z(n17704) );
CLKBUF_X2 U14260 ( .A(dii_data[27]), .Z(n17705) );
NAND2_X1 U14261 ( .A1(n17705), .A2(n17797), .ZN(n18483) );
CLKBUF_X2 U14262 ( .A(n5930), .Z(n17706) );
CLKBUF_X2 U14263 ( .A(dii_data[26]), .Z(n17707) );
NAND2_X1 U14264 ( .A1(n17707), .A2(n17797), .ZN(n18487) );
CLKBUF_X2 U14265 ( .A(n5931), .Z(n17708) );
CLKBUF_X2 U14266 ( .A(dii_data[25]), .Z(n17709) );
NAND2_X1 U14267 ( .A1(n17709), .A2(n17797), .ZN(n18491) );
CLKBUF_X2 U14268 ( .A(n5932), .Z(n17710) );
CLKBUF_X2 U14269 ( .A(dii_data[24]), .Z(n17711) );
NAND2_X1 U14270 ( .A1(n17711), .A2(n17797), .ZN(n18495) );
CLKBUF_X2 U14271 ( .A(n5933), .Z(n17712) );
CLKBUF_X2 U14272 ( .A(dii_data[23]), .Z(n17713) );
NAND2_X1 U14273 ( .A1(n17713), .A2(n17797), .ZN(n18499) );
CLKBUF_X2 U14274 ( .A(n5934), .Z(n17714) );
CLKBUF_X2 U14275 ( .A(dii_data[22]), .Z(n17715) );
NAND2_X1 U14276 ( .A1(n17715), .A2(n17797), .ZN(n18503) );
CLKBUF_X2 U14277 ( .A(n5935), .Z(n17716) );
CLKBUF_X2 U14278 ( .A(dii_data[21]), .Z(n17717) );
NAND2_X1 U14279 ( .A1(n17717), .A2(n17797), .ZN(n18507) );
CLKBUF_X2 U14280 ( .A(n5936), .Z(n17718) );
CLKBUF_X2 U14281 ( .A(dii_data[20]), .Z(n17719) );
NAND2_X1 U14282 ( .A1(n17719), .A2(n17797), .ZN(n18511) );
CLKBUF_X2 U14283 ( .A(n5937), .Z(n17720) );
CLKBUF_X2 U14284 ( .A(dii_data[19]), .Z(n17721) );
NAND2_X1 U14285 ( .A1(n17721), .A2(n17797), .ZN(n18515) );
CLKBUF_X2 U14286 ( .A(n5938), .Z(n17722) );
CLKBUF_X2 U14287 ( .A(dii_data[18]), .Z(n17723) );
NAND2_X1 U14288 ( .A1(n17723), .A2(n17797), .ZN(n18519) );
CLKBUF_X2 U14289 ( .A(n5939), .Z(n17724) );
CLKBUF_X2 U14290 ( .A(dii_data[17]), .Z(n17725) );
NAND2_X1 U14291 ( .A1(n17725), .A2(n17797), .ZN(n18523) );
CLKBUF_X2 U14292 ( .A(n5940), .Z(n17726) );
CLKBUF_X2 U14293 ( .A(dii_data[16]), .Z(n17727) );
NAND2_X1 U14294 ( .A1(n17727), .A2(n17798), .ZN(n18527) );
CLKBUF_X1 U14295 ( .A(dii_data[15]), .Z(n17728) );
NAND2_X1 U14296 ( .A1(n17728), .A2(n17798), .ZN(n18531) );
CLKBUF_X1 U14297 ( .A(dii_data[14]), .Z(n17729) );
NAND2_X1 U14298 ( .A1(n17729), .A2(n17798), .ZN(n18535) );
CLKBUF_X1 U14299 ( .A(dii_data[13]), .Z(n17730) );
NAND2_X1 U14300 ( .A1(n17730), .A2(n17798), .ZN(n18539) );
CLKBUF_X1 U14301 ( .A(dii_data[12]), .Z(n17731) );
NAND2_X1 U14302 ( .A1(n17731), .A2(n17798), .ZN(n18543) );
CLKBUF_X1 U14303 ( .A(dii_data[11]), .Z(n17732) );
NAND2_X1 U14304 ( .A1(n17732), .A2(n17798), .ZN(n18547) );
CLKBUF_X1 U14305 ( .A(dii_data[10]), .Z(n17733) );
NAND2_X1 U14306 ( .A1(n17733), .A2(n17798), .ZN(n18551) );
CLKBUF_X1 U14307 ( .A(dii_data[9]), .Z(n17734) );
NAND2_X1 U14308 ( .A1(n17734), .A2(n17798), .ZN(n18555) );
CLKBUF_X1 U14309 ( .A(dii_data[8]), .Z(n17735) );
NAND2_X1 U14310 ( .A1(n17735), .A2(n17798), .ZN(n18559) );
CLKBUF_X1 U14311 ( .A(dii_data[7]), .Z(n17736) );
NAND2_X1 U14312 ( .A1(n17736), .A2(n17798), .ZN(n18563) );
CLKBUF_X1 U14313 ( .A(dii_data[6]), .Z(n17737) );
NAND2_X1 U14314 ( .A1(n17737), .A2(n17798), .ZN(n18567) );
CLKBUF_X1 U14315 ( .A(dii_data[5]), .Z(n17738) );
NAND2_X1 U14316 ( .A1(n17738), .A2(n17799), .ZN(n18571) );
CLKBUF_X1 U14317 ( .A(dii_data[4]), .Z(n17739) );
NAND2_X1 U14318 ( .A1(n17739), .A2(n17799), .ZN(n18575) );
CLKBUF_X1 U14319 ( .A(dii_data[3]), .Z(n17740) );
NAND2_X1 U14320 ( .A1(n17740), .A2(n17799), .ZN(n18579) );
CLKBUF_X1 U14321 ( .A(dii_data[2]), .Z(n17741) );
NAND2_X1 U14322 ( .A1(n17741), .A2(n17799), .ZN(n18583) );
CLKBUF_X1 U14323 ( .A(dii_data[1]), .Z(n17742) );
NAND2_X1 U14324 ( .A1(n17742), .A2(n17799), .ZN(n18587) );
CLKBUF_X1 U14325 ( .A(dii_data[0]), .Z(n17743) );
NAND2_X1 U14326 ( .A1(n17743), .A2(n17799), .ZN(n18591) );
NAND3_X1 U14327 ( .A1(n18200), .A2(n18199), .A3(n18198), .ZN(n5957) );
CLKBUF_X2 U14328 ( .A(n5957), .Z(n17744) );
CLKBUF_X2 U14329 ( .A(dii_data[98]), .Z(n17745) );
NAND2_X1 U14330 ( .A1(n17745), .A2(n17790), .ZN(n18199) );
BUF_X16 U14331 ( .A(n11958), .Z(n17746) );
NAND2_X1 U14332 ( .A1(n17746), .A2(n11959), .ZN(n6284) );
NAND2_X1 U14333 ( .A1(n17990), .A2(cii_IV_vld), .ZN(n11958) );
BUF_X32 U14334 ( .A(n11930), .Z(n17747) );
NAND2_X1 U14335 ( .A1(cii_ctl_vld), .A2(n11971), .ZN(n11930) );
BUF_X16 U14336 ( .A(dii_last_word), .Z(n17749) );
NAND2_X1 U14337 ( .A1(n11927), .A2(n11928), .ZN(n6293) );
CLKBUF_X2 U14338 ( .A(n17749), .Z(n17748) );
OR3_X1 U14339 ( .A1(n18892), .A2(n17748), .A3(n11957), .ZN(n11949) );
NAND3_X1 U14340 ( .A1(n18744), .A2(n11946), .A3(n11947), .ZN(n6286) );
NAND3_X1 U14341 ( .A1(dii_data_type), .A2(dii_data_vld), .A3(n18617), .ZN(n11946) );
NAND2_X1 U14342 ( .A1(n11941), .A2(n18085), .ZN(n6288) );
MUX2_X1 U14343 ( .A(aad_byte_cnt[1]), .B(N2480), .S(n17837), .Z(n6019) );
CLKBUF_X1 U14344 ( .A(dii_data_size[0]), .Z(n17750) );
MUX2_X1 U14345 ( .A(enc_byte_cnt[0]), .B(N2349), .S(n17817), .Z(n5441) );
MUX2_X1 U14346 ( .A(enc_byte_cnt[1]), .B(N2350), .S(n17817), .Z(n5440) );
INV_X8 U14347 ( .A(rst), .ZN(n17751) );
INV_X8 U14348 ( .A(rst), .ZN(n17752) );
INV_X8 U14349 ( .A(rst), .ZN(n17753) );
INV_X4 U14350 ( .A(n16431), .ZN(n18634) );
INV_X4 U14351 ( .A(n18057), .ZN(n18036) );
INV_X4 U14352 ( .A(n18057), .ZN(n18037) );
INV_X4 U14353 ( .A(n17282), .ZN(n18044) );
INV_X4 U14354 ( .A(n18058), .ZN(n18045) );
INV_X4 U14355 ( .A(n18058), .ZN(n18046) );
INV_X4 U14356 ( .A(n18058), .ZN(n18048) );
INV_X4 U14357 ( .A(n18058), .ZN(n18049) );
INV_X4 U14358 ( .A(n18058), .ZN(n18050) );
INV_X4 U14359 ( .A(n18058), .ZN(n18047) );
INV_X4 U14360 ( .A(n17282), .ZN(n18042) );
INV_X4 U14361 ( .A(n18058), .ZN(n18041) );
INV_X4 U14362 ( .A(n18057), .ZN(n18039) );
INV_X4 U14363 ( .A(n18058), .ZN(n18040) );
INV_X4 U14364 ( .A(n18058), .ZN(n18038) );
INV_X4 U14365 ( .A(n17282), .ZN(n18043) );
INV_X4 U14366 ( .A(n18057), .ZN(n18052) );
INV_X4 U14367 ( .A(n18057), .ZN(n18053) );
INV_X4 U14368 ( .A(n18057), .ZN(n18051) );
INV_X4 U14369 ( .A(n17931), .ZN(n17928) );
INV_X4 U14370 ( .A(n17931), .ZN(n17922) );
INV_X4 U14371 ( .A(n17931), .ZN(n17923) );
INV_X4 U14372 ( .A(n17931), .ZN(n17924) );
INV_X4 U14373 ( .A(n17931), .ZN(n17925) );
INV_X4 U14374 ( .A(n17931), .ZN(n17926) );
INV_X4 U14375 ( .A(n17931), .ZN(n17927) );
INV_X4 U14376 ( .A(n17931), .ZN(n17929) );
INV_X4 U14377 ( .A(n17931), .ZN(n17919) );
INV_X4 U14378 ( .A(n17931), .ZN(n17920) );
INV_X4 U14379 ( .A(n17931), .ZN(n17921) );
INV_X4 U14380 ( .A(n17931), .ZN(n17930) );
INV_X4 U14381 ( .A(n16537), .ZN(n17849) );
INV_X4 U14382 ( .A(n16537), .ZN(n17850) );
INV_X4 U14383 ( .A(n16537), .ZN(n17851) );
INV_X4 U14384 ( .A(n18070), .ZN(n18058) );
INV_X4 U14385 ( .A(n17288), .ZN(n17931) );
INV_X4 U14386 ( .A(n18042), .ZN(n18060) );
INV_X4 U14387 ( .A(n18042), .ZN(n18063) );
INV_X4 U14388 ( .A(n18043), .ZN(n18062) );
INV_X4 U14389 ( .A(n18042), .ZN(n18061) );
INV_X4 U14390 ( .A(n18070), .ZN(n18059) );
INV_X4 U14391 ( .A(n18070), .ZN(n18064) );
INV_X4 U14392 ( .A(n18070), .ZN(n18065) );
INV_X4 U14393 ( .A(n18070), .ZN(n18066) );
INV_X4 U14394 ( .A(n16537), .ZN(n17848) );
INV_X4 U14395 ( .A(n18057), .ZN(n18055) );
INV_X4 U14396 ( .A(n18057), .ZN(n18054) );
INV_X4 U14397 ( .A(n17288), .ZN(n17932) );
INV_X4 U14398 ( .A(n17754), .ZN(n17944) );
INV_X4 U14399 ( .A(n17754), .ZN(n17943) );
INV_X4 U14400 ( .A(n17754), .ZN(n17942) );
INV_X4 U14401 ( .A(n17754), .ZN(n17941) );
INV_X4 U14402 ( .A(n17754), .ZN(n17939) );
INV_X4 U14403 ( .A(n17754), .ZN(n17940) );
INV_X4 U14404 ( .A(n17754), .ZN(n17938) );
INV_X4 U14405 ( .A(n17754), .ZN(n17937) );
INV_X4 U14406 ( .A(n17754), .ZN(n17936) );
INV_X4 U14407 ( .A(n17754), .ZN(n17934) );
INV_X4 U14408 ( .A(n18057), .ZN(n18056) );
INV_X4 U14409 ( .A(n17285), .ZN(n17949) );
INV_X4 U14410 ( .A(n17285), .ZN(n17950) );
INV_X4 U14411 ( .A(n17285), .ZN(n17951) );
INV_X4 U14412 ( .A(n17285), .ZN(n17952) );
INV_X4 U14413 ( .A(n17285), .ZN(n17953) );
INV_X4 U14414 ( .A(n17285), .ZN(n17954) );
INV_X4 U14415 ( .A(n17285), .ZN(n17955) );
INV_X4 U14416 ( .A(n17285), .ZN(n17956) );
INV_X4 U14417 ( .A(n18083), .ZN(n17779) );
INV_X4 U14418 ( .A(n18083), .ZN(n17780) );
INV_X4 U14419 ( .A(n18083), .ZN(n17781) );
INV_X4 U14420 ( .A(n18083), .ZN(n17782) );
INV_X4 U14421 ( .A(n18083), .ZN(n17783) );
INV_X4 U14422 ( .A(n18083), .ZN(n17784) );
INV_X4 U14423 ( .A(n18083), .ZN(n17785) );
INV_X4 U14424 ( .A(n18083), .ZN(n17786) );
INV_X4 U14425 ( .A(n17754), .ZN(n17935) );
INV_X4 U14426 ( .A(n17754), .ZN(n17945) );
INV_X4 U14427 ( .A(n17285), .ZN(n17957) );
INV_X4 U14428 ( .A(n18083), .ZN(n17787) );
NOR2_X2 U14429 ( .A1(n16325), .A2(n16326), .ZN(n16209) );
NAND2_X2 U14430 ( .A1(n16431), .A2(n16432), .ZN(n16325) );
INV_X4 U14431 ( .A(n17282), .ZN(n18070) );
INV_X4 U14432 ( .A(n18070), .ZN(n18067) );
INV_X4 U14433 ( .A(n18070), .ZN(n18068) );
INV_X4 U14434 ( .A(n14167), .ZN(n17900) );
INV_X4 U14435 ( .A(n14167), .ZN(n17901) );
INV_X4 U14436 ( .A(n14167), .ZN(n17902) );
INV_X4 U14437 ( .A(n14167), .ZN(n17903) );
INV_X4 U14438 ( .A(n14167), .ZN(n17904) );
INV_X4 U14439 ( .A(n14167), .ZN(n17905) );
INV_X4 U14440 ( .A(n15509), .ZN(n17864) );
INV_X4 U14441 ( .A(n17877), .ZN(n17876) );
INV_X4 U14442 ( .A(n17284), .ZN(n17910) );
INV_X4 U14443 ( .A(n17284), .ZN(n17909) );
INV_X4 U14444 ( .A(n17284), .ZN(n17914) );
INV_X4 U14445 ( .A(n17284), .ZN(n17913) );
INV_X4 U14446 ( .A(n17284), .ZN(n17912) );
INV_X4 U14447 ( .A(n17284), .ZN(n17911) );
INV_X4 U14448 ( .A(n17284), .ZN(n17915) );
INV_X4 U14449 ( .A(n17285), .ZN(n17946) );
INV_X4 U14450 ( .A(n17285), .ZN(n17947) );
INV_X4 U14451 ( .A(n17285), .ZN(n17948) );
INV_X4 U14452 ( .A(n18083), .ZN(n17776) );
INV_X4 U14453 ( .A(n18083), .ZN(n17777) );
INV_X4 U14454 ( .A(n18083), .ZN(n17778) );
INV_X4 U14455 ( .A(n18084), .ZN(n17791) );
INV_X4 U14456 ( .A(n18084), .ZN(n17792) );
INV_X4 U14457 ( .A(n18084), .ZN(n17793) );
INV_X4 U14458 ( .A(n18084), .ZN(n17794) );
INV_X4 U14459 ( .A(n18084), .ZN(n17795) );
INV_X4 U14460 ( .A(n18084), .ZN(n17796) );
INV_X4 U14461 ( .A(n18084), .ZN(n17797) );
INV_X4 U14462 ( .A(n18084), .ZN(n17798) );
INV_X4 U14463 ( .A(n18043), .ZN(n18069) );
INV_X4 U14464 ( .A(n17754), .ZN(n17933) );
INV_X4 U14465 ( .A(n18602), .ZN(n18014) );
INV_X4 U14466 ( .A(n18070), .ZN(n18057) );
INV_X4 U14467 ( .A(n18084), .ZN(n17799) );
INV_X4 U14468 ( .A(n17284), .ZN(n17916) );
INV_X4 U14469 ( .A(n17877), .ZN(n17875) );
INV_X4 U14470 ( .A(n17877), .ZN(n17874) );
INV_X4 U14471 ( .A(n15509), .ZN(n17862) );
INV_X4 U14472 ( .A(n15509), .ZN(n17863) );
INV_X4 U14473 ( .A(n15509), .ZN(n17861) );
INV_X4 U14474 ( .A(n15509), .ZN(n17860) );
INV_X4 U14475 ( .A(n11961), .ZN(n17842) );
INV_X4 U14476 ( .A(n11961), .ZN(n17843) );
INV_X4 U14477 ( .A(n11961), .ZN(n17844) );
INV_X4 U14478 ( .A(n11961), .ZN(n17845) );
INV_X4 U14479 ( .A(n11961), .ZN(n17846) );
INV_X4 U14480 ( .A(n11961), .ZN(n17847) );
INV_X4 U14481 ( .A(n17989), .ZN(n17982) );
INV_X4 U14482 ( .A(n17989), .ZN(n17981) );
INV_X4 U14483 ( .A(n17989), .ZN(n17980) );
INV_X4 U14484 ( .A(n17989), .ZN(n17979) );
INV_X4 U14485 ( .A(n17989), .ZN(n17978) );
INV_X4 U14486 ( .A(n17989), .ZN(n17977) );
INV_X4 U14487 ( .A(n18602), .ZN(n18006) );
INV_X4 U14488 ( .A(n18602), .ZN(n18007) );
INV_X4 U14489 ( .A(n18602), .ZN(n18008) );
INV_X4 U14490 ( .A(n18602), .ZN(n18009) );
INV_X4 U14491 ( .A(n18602), .ZN(n18010) );
INV_X4 U14492 ( .A(n18602), .ZN(n18011) );
INV_X4 U14493 ( .A(n18602), .ZN(n18012) );
INV_X4 U14494 ( .A(n18602), .ZN(n18013) );
INV_X4 U14495 ( .A(n17989), .ZN(n17987) );
INV_X4 U14496 ( .A(n17989), .ZN(n17986) );
INV_X4 U14497 ( .A(n17989), .ZN(n17985) );
INV_X4 U14498 ( .A(n17989), .ZN(n17984) );
INV_X4 U14499 ( .A(n17989), .ZN(n17983) );
INV_X4 U14500 ( .A(n18085), .ZN(n17803) );
INV_X4 U14501 ( .A(n18085), .ZN(n17804) );
INV_X4 U14502 ( .A(n18085), .ZN(n17805) );
INV_X4 U14503 ( .A(n18085), .ZN(n17806) );
INV_X4 U14504 ( .A(n18085), .ZN(n17807) );
INV_X4 U14505 ( .A(n18085), .ZN(n17808) );
INV_X4 U14506 ( .A(n18085), .ZN(n17809) );
INV_X4 U14507 ( .A(n18085), .ZN(n17810) );
INV_X4 U14508 ( .A(n18085), .ZN(n17811) );
INV_X4 U14509 ( .A(n17989), .ZN(n17988) );
NOR2_X2 U14510 ( .A1(n15805), .A2(n15806), .ZN(n15663) );
BUF_X4 U14511 ( .A(n11956), .Z(n18026) );
BUF_X4 U14512 ( .A(n11956), .Z(n18034) );
BUF_X4 U14513 ( .A(n11956), .Z(n18033) );
BUF_X4 U14514 ( .A(n11956), .Z(n18032) );
BUF_X4 U14515 ( .A(n11956), .Z(n18031) );
BUF_X4 U14516 ( .A(n11956), .Z(n18030) );
BUF_X4 U14517 ( .A(n11956), .Z(n18029) );
BUF_X4 U14518 ( .A(n11956), .Z(n18028) );
BUF_X4 U14519 ( .A(n11956), .Z(n18027) );
BUF_X4 U14520 ( .A(n11956), .Z(n18035) );
INV_X4 U14521 ( .A(n15501), .ZN(n17877) );
INV_X4 U14522 ( .A(n17916), .ZN(n17918) );
INV_X4 U14523 ( .A(n17916), .ZN(n17917) );
INV_X4 U14524 ( .A(n18000), .ZN(n17996) );
INV_X4 U14525 ( .A(n18001), .ZN(n17999) );
INV_X4 U14526 ( .A(n17905), .ZN(n17906) );
INV_X4 U14527 ( .A(n17903), .ZN(n17907) );
INV_X4 U14528 ( .A(n12238), .ZN(n17990) );
INV_X4 U14529 ( .A(n15508), .ZN(n17857) );
INV_X4 U14530 ( .A(n17904), .ZN(n17908) );
INV_X4 U14531 ( .A(n18084), .ZN(n17788) );
INV_X4 U14532 ( .A(n18084), .ZN(n17789) );
INV_X4 U14533 ( .A(n18084), .ZN(n17790) );
INV_X4 U14534 ( .A(n11961), .ZN(n17841) );
BUF_X4 U14535 ( .A(n11956), .Z(n18025) );
BUF_X4 U14536 ( .A(n11956), .Z(n18024) );
BUF_X4 U14537 ( .A(n11956), .Z(n18023) );
BUF_X4 U14538 ( .A(n11956), .Z(n18021) );
BUF_X4 U14539 ( .A(n11956), .Z(n18022) );
BUF_X4 U14540 ( .A(n11956), .Z(n18019) );
BUF_X4 U14541 ( .A(n11956), .Z(n18018) );
BUF_X4 U14542 ( .A(n11956), .Z(n18017) );
BUF_X4 U14543 ( .A(n11956), .Z(n18016) );
BUF_X4 U14544 ( .A(n11956), .Z(n18015) );
BUF_X4 U14545 ( .A(n11956), .Z(n18020) );
INV_X4 U14546 ( .A(n12238), .ZN(n17989) );
INV_X4 U14547 ( .A(n14564), .ZN(n17867) );
INV_X4 U14548 ( .A(n14564), .ZN(n17866) );
INV_X4 U14549 ( .A(n18000), .ZN(n17997) );
INV_X4 U14550 ( .A(n18001), .ZN(n17998) );
INV_X4 U14551 ( .A(n11946), .ZN(n17839) );
INV_X4 U14552 ( .A(n11946), .ZN(n17838) );
INV_X4 U14553 ( .A(n17988), .ZN(n17993) );
INV_X4 U14554 ( .A(n17988), .ZN(n17992) );
INV_X4 U14555 ( .A(n17988), .ZN(n17991) );
INV_X4 U14556 ( .A(n15508), .ZN(n17858) );
INV_X4 U14557 ( .A(n11946), .ZN(n17840) );
INV_X4 U14558 ( .A(n15508), .ZN(n17859) );
INV_X4 U14559 ( .A(n11939), .ZN(n17812) );
INV_X4 U14560 ( .A(n11939), .ZN(n17813) );
INV_X4 U14561 ( .A(n11939), .ZN(n17814) );
INV_X4 U14562 ( .A(n11939), .ZN(n17815) );
INV_X4 U14563 ( .A(n11939), .ZN(n17816) );
INV_X4 U14564 ( .A(n11939), .ZN(n17817) );
INV_X4 U14565 ( .A(n17286), .ZN(n17968) );
INV_X4 U14566 ( .A(n17286), .ZN(n17969) );
INV_X4 U14567 ( .A(n17286), .ZN(n17970) );
INV_X4 U14568 ( .A(n17286), .ZN(n17971) );
INV_X4 U14569 ( .A(n17286), .ZN(n17972) );
INV_X4 U14570 ( .A(n17286), .ZN(n17973) );
INV_X4 U14571 ( .A(n17286), .ZN(n17974) );
INV_X4 U14572 ( .A(n17286), .ZN(n17975) );
INV_X4 U14573 ( .A(n17885), .ZN(n17884) );
INV_X4 U14574 ( .A(n17885), .ZN(n17883) );
INV_X4 U14575 ( .A(n15507), .ZN(n17854) );
INV_X4 U14576 ( .A(n15507), .ZN(n17855) );
INV_X4 U14577 ( .A(n18602), .ZN(n18004) );
INV_X4 U14578 ( .A(n18602), .ZN(n18005) );
INV_X4 U14579 ( .A(n18602), .ZN(n18003) );
INV_X4 U14580 ( .A(n15507), .ZN(n17852) );
INV_X4 U14581 ( .A(n15507), .ZN(n17853) );
INV_X4 U14582 ( .A(n18085), .ZN(n17800) );
INV_X4 U14583 ( .A(n18085), .ZN(n17801) );
INV_X4 U14584 ( .A(n18085), .ZN(n17802) );
INV_X4 U14585 ( .A(n17286), .ZN(n17976) );
INV_X4 U14586 ( .A(n15507), .ZN(n17856) );
NAND2_X2 U14587 ( .A1(n17934), .A2(n15644), .ZN(n15946) );
OR2_X2 U14588 ( .A1(n18744), .A2(n16542), .ZN(n17754) );
NAND2_X2 U14589 ( .A1(n15946), .A2(n15947), .ZN(n15805) );
NOR4_X2 U14590 ( .A1(n15644), .A2(n19202), .A3(n17755), .A4(n15509), .ZN(n15272) );
INV_X4 U14591 ( .A(n18633), .ZN(n11956) );
NOR2_X2 U14592 ( .A1(n17291), .A2(n18059), .ZN(n17280) );
INV_X4 U14593 ( .A(n17283), .ZN(n18000) );
INV_X4 U14594 ( .A(n14422), .ZN(n17885) );
INV_X4 U14595 ( .A(n11946), .ZN(n17837) );
INV_X4 U14596 ( .A(n17756), .ZN(n17872) );
INV_X4 U14597 ( .A(n15501), .ZN(n17873) );
INV_X4 U14598 ( .A(n17891), .ZN(n17887) );
INV_X4 U14599 ( .A(n17287), .ZN(n17892) );
INV_X4 U14600 ( .A(n17757), .ZN(n17880) );
NOR2_X2 U14601 ( .A1(n17886), .A2(n14190), .ZN(n14189) );
NOR2_X2 U14602 ( .A1(n17886), .A2(n14219), .ZN(n14218) );
NOR2_X2 U14603 ( .A1(n17886), .A2(n14248), .ZN(n14247) );
NOR2_X2 U14604 ( .A1(n17886), .A2(n14277), .ZN(n14276) );
NOR2_X2 U14605 ( .A1(n17886), .A2(n14306), .ZN(n14305) );
NOR2_X2 U14606 ( .A1(n17886), .A2(n14335), .ZN(n14334) );
NOR2_X2 U14607 ( .A1(n17886), .A2(n14364), .ZN(n14363) );
NOR2_X2 U14608 ( .A1(n17891), .A2(n14396), .ZN(n14395) );
NOR2_X2 U14609 ( .A1(n17866), .A2(n14191), .ZN(n14188) );
NOR2_X2 U14610 ( .A1(n17865), .A2(n14220), .ZN(n14217) );
NOR2_X2 U14611 ( .A1(n17865), .A2(n14249), .ZN(n14246) );
NOR2_X2 U14612 ( .A1(n17865), .A2(n14278), .ZN(n14275) );
NOR2_X2 U14613 ( .A1(n17865), .A2(n14307), .ZN(n14304) );
NOR2_X2 U14614 ( .A1(n17866), .A2(n14336), .ZN(n14333) );
NOR2_X2 U14615 ( .A1(n17866), .A2(n14365), .ZN(n14362) );
NOR2_X2 U14616 ( .A1(n17866), .A2(n14397), .ZN(n14394) );
INV_X4 U14617 ( .A(n17757), .ZN(n17881) );
INV_X4 U14618 ( .A(n17756), .ZN(n17871) );
INV_X4 U14619 ( .A(n17756), .ZN(n17870) );
INV_X4 U14620 ( .A(n17755), .ZN(n17869) );
INV_X4 U14621 ( .A(n17755), .ZN(n17868) );
INV_X4 U14622 ( .A(n17758), .ZN(n17879) );
INV_X4 U14623 ( .A(n17758), .ZN(n17878) );
INV_X4 U14624 ( .A(n17283), .ZN(n18001) );
INV_X4 U14625 ( .A(n17988), .ZN(n17995) );
INV_X4 U14626 ( .A(n17985), .ZN(n17994) );
INV_X4 U14627 ( .A(n14564), .ZN(n17865) );
INV_X4 U14628 ( .A(n17289), .ZN(n17963) );
INV_X4 U14629 ( .A(n17289), .ZN(n17962) );
INV_X4 U14630 ( .A(n17289), .ZN(n17960) );
INV_X4 U14631 ( .A(n17289), .ZN(n17959) );
INV_X4 U14632 ( .A(n17289), .ZN(n17961) );
INV_X4 U14633 ( .A(n17289), .ZN(n17964) );
INV_X4 U14634 ( .A(n15504), .ZN(n19202) );
INV_X4 U14635 ( .A(n17891), .ZN(n17889) );
INV_X4 U14636 ( .A(n17886), .ZN(n17888) );
INV_X4 U14637 ( .A(n17287), .ZN(n17895) );
INV_X4 U14638 ( .A(n17287), .ZN(n17894) );
INV_X4 U14639 ( .A(n17287), .ZN(n17893) );
INV_X4 U14640 ( .A(n17286), .ZN(n17965) );
INV_X4 U14641 ( .A(n17286), .ZN(n17966) );
INV_X4 U14642 ( .A(n17286), .ZN(n17967) );
INV_X4 U14643 ( .A(n17885), .ZN(n17882) );
INV_X4 U14644 ( .A(n17886), .ZN(n17890) );
INV_X4 U14645 ( .A(n17287), .ZN(n17896) );
NOR3_X2 U14646 ( .A1(n19204), .A2(n19205), .A3(n18071), .ZN(n15509) );
AND2_X2 U14647 ( .A1(n17887), .A2(n15309), .ZN(n17755) );
NAND2_X2 U14648 ( .A1(n14564), .A2(n14422), .ZN(n15508) );
NOR2_X2 U14649 ( .A1(n17848), .A2(n17857), .ZN(n16083) );
NOR2_X2 U14650 ( .A1(n17864), .A2(n18075), .ZN(n16542) );
NOR4_X2 U14651 ( .A1(n14583), .A2(n14584), .A3(n14585), .A4(n18735), .ZN(n14582) );
NOR2_X2 U14652 ( .A1(n19032), .A2(n17900), .ZN(n14584) );
NOR4_X2 U14653 ( .A1(n14605), .A2(n14606), .A3(n14607), .A4(n18734), .ZN(n14604) );
NOR2_X2 U14654 ( .A1(n19034), .A2(n17900), .ZN(n14606) );
NOR4_X2 U14655 ( .A1(n14626), .A2(n14627), .A3(n14628), .A4(n18733), .ZN(n14625) );
NOR2_X2 U14656 ( .A1(n19036), .A2(n17900), .ZN(n14627) );
NOR4_X2 U14657 ( .A1(n14647), .A2(n14648), .A3(n14649), .A4(n18732), .ZN(n14646) );
NOR2_X2 U14658 ( .A1(n19038), .A2(n17900), .ZN(n14648) );
NOR4_X2 U14659 ( .A1(n14668), .A2(n14669), .A3(n14670), .A4(n18731), .ZN(n14667) );
NOR2_X2 U14660 ( .A1(n19040), .A2(n17900), .ZN(n14669) );
NOR4_X2 U14661 ( .A1(n14689), .A2(n14690), .A3(n14691), .A4(n18730), .ZN(n14688) );
NOR2_X2 U14662 ( .A1(n19042), .A2(n17900), .ZN(n14690) );
NOR4_X2 U14663 ( .A1(n14710), .A2(n14711), .A3(n14712), .A4(n18729), .ZN(n14709) );
NOR2_X2 U14664 ( .A1(n19044), .A2(n17900), .ZN(n14711) );
NOR4_X2 U14665 ( .A1(n14731), .A2(n14732), .A3(n14733), .A4(n18728), .ZN(n14730) );
NOR2_X2 U14666 ( .A1(n19046), .A2(n17900), .ZN(n14732) );
NOR4_X2 U14667 ( .A1(n14754), .A2(n14755), .A3(n14756), .A4(n18727), .ZN(n14753) );
NOR2_X2 U14668 ( .A1(n19048), .A2(n17900), .ZN(n14755) );
NOR4_X2 U14669 ( .A1(n14778), .A2(n14779), .A3(n14780), .A4(n18726), .ZN(n14777) );
NOR2_X2 U14670 ( .A1(n19050), .A2(n17900), .ZN(n14779) );
NOR4_X2 U14671 ( .A1(n14800), .A2(n14801), .A3(n14802), .A4(n18725), .ZN(n14799) );
NOR2_X2 U14672 ( .A1(n19052), .A2(n17900), .ZN(n14801) );
NOR4_X2 U14673 ( .A1(n14822), .A2(n14823), .A3(n14824), .A4(n18724), .ZN(n14821) );
NOR2_X2 U14674 ( .A1(n19054), .A2(n17900), .ZN(n14823) );
NOR4_X2 U14675 ( .A1(n14844), .A2(n14845), .A3(n14846), .A4(n18723), .ZN(n14843) );
NOR2_X2 U14676 ( .A1(n19056), .A2(n17901), .ZN(n14845) );
NOR4_X2 U14677 ( .A1(n14866), .A2(n14867), .A3(n14868), .A4(n18722), .ZN(n14865) );
NOR2_X2 U14678 ( .A1(n19058), .A2(n17901), .ZN(n14867) );
NOR4_X2 U14679 ( .A1(n14888), .A2(n14889), .A3(n14890), .A4(n18721), .ZN(n14887) );
NOR2_X2 U14680 ( .A1(n19060), .A2(n17901), .ZN(n14889) );
NOR4_X2 U14681 ( .A1(n14910), .A2(n14911), .A3(n14912), .A4(n18720), .ZN(n14909) );
NOR2_X2 U14682 ( .A1(n19062), .A2(n17901), .ZN(n14911) );
NOR4_X2 U14683 ( .A1(n14933), .A2(n14934), .A3(n14935), .A4(n18719), .ZN(n14932) );
NOR2_X2 U14684 ( .A1(n19064), .A2(n17901), .ZN(n14934) );
NOR4_X2 U14685 ( .A1(n14957), .A2(n14958), .A3(n14959), .A4(n18718), .ZN(n14956) );
NOR2_X2 U14686 ( .A1(n19066), .A2(n17901), .ZN(n14958) );
NOR4_X2 U14687 ( .A1(n14979), .A2(n14980), .A3(n14981), .A4(n18717), .ZN(n14978) );
NOR2_X2 U14688 ( .A1(n19068), .A2(n17901), .ZN(n14980) );
NOR4_X2 U14689 ( .A1(n15001), .A2(n15002), .A3(n15003), .A4(n18716), .ZN(n15000) );
NOR2_X2 U14690 ( .A1(n19070), .A2(n17901), .ZN(n15002) );
NOR4_X2 U14691 ( .A1(n15023), .A2(n15024), .A3(n15025), .A4(n18715), .ZN(n15022) );
NOR2_X2 U14692 ( .A1(n19072), .A2(n17901), .ZN(n15024) );
NOR4_X2 U14693 ( .A1(n15045), .A2(n15046), .A3(n15047), .A4(n18714), .ZN(n15044) );
NOR2_X2 U14694 ( .A1(n19074), .A2(n17901), .ZN(n15046) );
NOR4_X2 U14695 ( .A1(n15067), .A2(n15068), .A3(n15069), .A4(n18713), .ZN(n15066) );
NOR2_X2 U14696 ( .A1(n19076), .A2(n17901), .ZN(n15068) );
NOR4_X2 U14697 ( .A1(n15089), .A2(n15090), .A3(n15091), .A4(n18712), .ZN(n15088) );
NOR2_X2 U14698 ( .A1(n19078), .A2(n17901), .ZN(n15090) );
NOR4_X2 U14699 ( .A1(n15113), .A2(n15114), .A3(n15115), .A4(n18711), .ZN(n15112) );
NOR2_X2 U14700 ( .A1(n19081), .A2(n17902), .ZN(n15114) );
NOR4_X2 U14701 ( .A1(n15136), .A2(n15137), .A3(n15138), .A4(n18710), .ZN(n15135) );
NOR2_X2 U14702 ( .A1(n19084), .A2(n17902), .ZN(n15137) );
NOR4_X2 U14703 ( .A1(n15158), .A2(n15159), .A3(n15160), .A4(n18709), .ZN(n15157) );
NOR2_X2 U14704 ( .A1(n19087), .A2(n17902), .ZN(n15159) );
NOR4_X2 U14705 ( .A1(n15180), .A2(n15181), .A3(n15182), .A4(n18708), .ZN(n15179) );
NOR2_X2 U14706 ( .A1(n19090), .A2(n17902), .ZN(n15181) );
NOR4_X2 U14707 ( .A1(n15202), .A2(n15203), .A3(n15204), .A4(n18707), .ZN(n15201) );
NOR2_X2 U14708 ( .A1(n19093), .A2(n17902), .ZN(n15203) );
NOR4_X2 U14709 ( .A1(n15224), .A2(n15225), .A3(n15226), .A4(n18706), .ZN(n15223) );
NOR2_X2 U14710 ( .A1(n19096), .A2(n17902), .ZN(n15225) );
NOR4_X2 U14711 ( .A1(n15246), .A2(n15247), .A3(n15248), .A4(n18705), .ZN(n15245) );
NOR2_X2 U14712 ( .A1(n19099), .A2(n17902), .ZN(n15247) );
NOR4_X2 U14713 ( .A1(n15268), .A2(n15269), .A3(n15270), .A4(n18704), .ZN(n15267) );
NOR2_X2 U14714 ( .A1(n19102), .A2(n17902), .ZN(n15269) );
NOR4_X2 U14715 ( .A1(n15292), .A2(n15293), .A3(n15294), .A4(n18703), .ZN(n15291) );
NOR2_X2 U14716 ( .A1(n19105), .A2(n17902), .ZN(n15293) );
NOR4_X2 U14717 ( .A1(n15318), .A2(n15319), .A3(n15320), .A4(n18702), .ZN(n15317) );
NOR2_X2 U14718 ( .A1(n19108), .A2(n17902), .ZN(n15319) );
NOR4_X2 U14719 ( .A1(n15342), .A2(n15343), .A3(n15344), .A4(n18701), .ZN(n15341) );
NOR2_X2 U14720 ( .A1(n19111), .A2(n17902), .ZN(n15343) );
NOR4_X2 U14721 ( .A1(n15366), .A2(n15367), .A3(n15368), .A4(n18700), .ZN(n15365) );
NOR2_X2 U14722 ( .A1(n19114), .A2(n17902), .ZN(n15367) );
NOR4_X2 U14723 ( .A1(n15390), .A2(n15391), .A3(n15392), .A4(n18699), .ZN(n15389) );
NOR2_X2 U14724 ( .A1(n19117), .A2(n17903), .ZN(n15391) );
NOR4_X2 U14725 ( .A1(n15414), .A2(n15415), .A3(n15416), .A4(n18698), .ZN(n15413) );
NOR2_X2 U14726 ( .A1(n19120), .A2(n17903), .ZN(n15415) );
NOR4_X2 U14727 ( .A1(n15438), .A2(n15439), .A3(n15440), .A4(n18697), .ZN(n15437) );
NOR2_X2 U14728 ( .A1(n19123), .A2(n17903), .ZN(n15439) );
NOR4_X2 U14729 ( .A1(n15462), .A2(n15463), .A3(n15464), .A4(n18696), .ZN(n15461) );
NOR2_X2 U14730 ( .A1(n19126), .A2(n17903), .ZN(n15463) );
NOR4_X2 U14731 ( .A1(n18695), .A2(n15488), .A3(n15489), .A4(n15490), .ZN(n15487) );
NOR2_X2 U14732 ( .A1(n15491), .A2(n17284), .ZN(n15490) );
NOR4_X2 U14733 ( .A1(n18694), .A2(n15517), .A3(n15518), .A4(n15519), .ZN(n15516) );
NOR2_X2 U14734 ( .A1(n15520), .A2(n17918), .ZN(n15519) );
NOR4_X2 U14735 ( .A1(n18693), .A2(n15538), .A3(n15539), .A4(n15540), .ZN(n15537) );
NOR2_X2 U14736 ( .A1(n15541), .A2(n17918), .ZN(n15540) );
NOR4_X2 U14737 ( .A1(n18692), .A2(n15559), .A3(n15560), .A4(n15561), .ZN(n15558) );
NOR2_X2 U14738 ( .A1(n15562), .A2(n17918), .ZN(n15561) );
NOR4_X2 U14739 ( .A1(n18691), .A2(n15580), .A3(n15581), .A4(n15582), .ZN(n15579) );
NOR2_X2 U14740 ( .A1(n15583), .A2(n17918), .ZN(n15582) );
NOR4_X2 U14741 ( .A1(n18658), .A2(n16220), .A3(n16221), .A4(n16222), .ZN(n16219) );
NOR2_X2 U14742 ( .A1(n16223), .A2(n17917), .ZN(n16222) );
NOR4_X2 U14743 ( .A1(n18657), .A2(n16234), .A3(n16235), .A4(n16236), .ZN(n16233) );
NOR2_X2 U14744 ( .A1(n16237), .A2(n17917), .ZN(n16236) );
NOR4_X2 U14745 ( .A1(n18656), .A2(n16248), .A3(n16249), .A4(n16250), .ZN(n16247) );
NOR2_X2 U14746 ( .A1(n16251), .A2(n17917), .ZN(n16250) );
NOR4_X2 U14747 ( .A1(n18655), .A2(n16262), .A3(n16263), .A4(n16264), .ZN(n16261) );
NOR2_X2 U14748 ( .A1(n16265), .A2(n17284), .ZN(n16264) );
NOR4_X2 U14749 ( .A1(n18654), .A2(n16276), .A3(n16277), .A4(n16278), .ZN(n16275) );
NOR2_X2 U14750 ( .A1(n16279), .A2(n17284), .ZN(n16278) );
NOR4_X2 U14751 ( .A1(n18653), .A2(n16290), .A3(n16291), .A4(n16292), .ZN(n16289) );
NOR2_X2 U14752 ( .A1(n16293), .A2(n17284), .ZN(n16292) );
NOR4_X2 U14753 ( .A1(n18652), .A2(n16304), .A3(n16305), .A4(n16306), .ZN(n16303) );
NOR2_X2 U14754 ( .A1(n16307), .A2(n17284), .ZN(n16306) );
NOR4_X2 U14755 ( .A1(n18651), .A2(n16318), .A3(n16319), .A4(n16320), .ZN(n16317) );
NOR2_X2 U14756 ( .A1(n16321), .A2(n17284), .ZN(n16320) );
NOR4_X2 U14757 ( .A1(n18690), .A2(n15659), .A3(n15660), .A4(n15661), .ZN(n15658) );
NOR2_X2 U14758 ( .A1(n15662), .A2(n17918), .ZN(n15661) );
NOR4_X2 U14759 ( .A1(n18689), .A2(n15679), .A3(n15680), .A4(n15681), .ZN(n15678) );
NOR2_X2 U14760 ( .A1(n15682), .A2(n17918), .ZN(n15681) );
NOR4_X2 U14761 ( .A1(n18688), .A2(n15698), .A3(n15699), .A4(n15700), .ZN(n15697) );
NOR2_X2 U14762 ( .A1(n15701), .A2(n17918), .ZN(n15700) );
NOR4_X2 U14763 ( .A1(n18687), .A2(n15717), .A3(n15718), .A4(n15719), .ZN(n15716) );
NOR2_X2 U14764 ( .A1(n15720), .A2(n17918), .ZN(n15719) );
NOR4_X2 U14765 ( .A1(n18686), .A2(n15736), .A3(n15737), .A4(n15738), .ZN(n15735) );
NOR2_X2 U14766 ( .A1(n15739), .A2(n17918), .ZN(n15738) );
NOR4_X2 U14767 ( .A1(n18685), .A2(n15755), .A3(n15756), .A4(n15757), .ZN(n15754) );
NOR2_X2 U14768 ( .A1(n15758), .A2(n17918), .ZN(n15757) );
NOR4_X2 U14769 ( .A1(n18684), .A2(n15774), .A3(n15775), .A4(n15776), .ZN(n15773) );
NOR2_X2 U14770 ( .A1(n15777), .A2(n17917), .ZN(n15776) );
NOR4_X2 U14771 ( .A1(n18683), .A2(n15793), .A3(n15794), .A4(n15795), .ZN(n15792) );
NOR2_X2 U14772 ( .A1(n15796), .A2(n17917), .ZN(n15795) );
NOR4_X2 U14773 ( .A1(n18674), .A2(n15960), .A3(n15961), .A4(n15962), .ZN(n15959) );
NOR2_X2 U14774 ( .A1(n15963), .A2(n17917), .ZN(n15962) );
NOR4_X2 U14775 ( .A1(n18673), .A2(n15977), .A3(n15978), .A4(n15979), .ZN(n15976) );
NOR2_X2 U14776 ( .A1(n15980), .A2(n17917), .ZN(n15979) );
NOR4_X2 U14777 ( .A1(n18672), .A2(n15994), .A3(n15995), .A4(n15996), .ZN(n15993) );
NOR2_X2 U14778 ( .A1(n15997), .A2(n17917), .ZN(n15996) );
NOR4_X2 U14779 ( .A1(n18671), .A2(n16011), .A3(n16012), .A4(n16013), .ZN(n16010) );
NOR2_X2 U14780 ( .A1(n16014), .A2(n17917), .ZN(n16013) );
NOR4_X2 U14781 ( .A1(n18670), .A2(n16028), .A3(n16029), .A4(n16030), .ZN(n16027) );
NOR2_X2 U14782 ( .A1(n16031), .A2(n17917), .ZN(n16030) );
NOR4_X2 U14783 ( .A1(n18669), .A2(n16045), .A3(n16046), .A4(n16047), .ZN(n16044) );
NOR2_X2 U14784 ( .A1(n16048), .A2(n17917), .ZN(n16047) );
NOR4_X2 U14785 ( .A1(n18668), .A2(n16062), .A3(n16063), .A4(n16064), .ZN(n16061) );
NOR2_X2 U14786 ( .A1(n16065), .A2(n17917), .ZN(n16064) );
NOR4_X2 U14787 ( .A1(n18667), .A2(n16079), .A3(n16080), .A4(n16081), .ZN(n16078) );
NOR2_X2 U14788 ( .A1(n16082), .A2(n17917), .ZN(n16081) );
NOR2_X2 U14789 ( .A1(n13802), .A2(n15117), .ZN(n15115) );
NOR2_X2 U14790 ( .A1(n13796), .A2(n15117), .ZN(n15138) );
NOR2_X2 U14791 ( .A1(n13790), .A2(n15117), .ZN(n15160) );
NOR2_X2 U14792 ( .A1(n13784), .A2(n15117), .ZN(n15182) );
NOR2_X2 U14793 ( .A1(n13778), .A2(n15117), .ZN(n15204) );
NOR2_X2 U14794 ( .A1(n13772), .A2(n15117), .ZN(n15226) );
NOR2_X2 U14795 ( .A1(n13766), .A2(n15117), .ZN(n15248) );
NOR2_X2 U14796 ( .A1(n13760), .A2(n15117), .ZN(n15270) );
NOR2_X2 U14797 ( .A1(n13898), .A2(n14758), .ZN(n14756) );
NOR2_X2 U14798 ( .A1(n13892), .A2(n14758), .ZN(n14780) );
NOR2_X2 U14799 ( .A1(n13886), .A2(n14758), .ZN(n14802) );
NOR2_X2 U14800 ( .A1(n13880), .A2(n14758), .ZN(n14824) );
NOR2_X2 U14801 ( .A1(n13874), .A2(n14758), .ZN(n14846) );
NOR2_X2 U14802 ( .A1(n13868), .A2(n14758), .ZN(n14868) );
NOR2_X2 U14803 ( .A1(n13862), .A2(n14758), .ZN(n14890) );
NOR2_X2 U14804 ( .A1(n13856), .A2(n14758), .ZN(n14912) );
NOR2_X2 U14805 ( .A1(n13754), .A2(n15296), .ZN(n15294) );
NOR2_X2 U14806 ( .A1(n13748), .A2(n15296), .ZN(n15320) );
NOR2_X2 U14807 ( .A1(n13742), .A2(n15296), .ZN(n15344) );
NOR2_X2 U14808 ( .A1(n13736), .A2(n15296), .ZN(n15368) );
NOR2_X2 U14809 ( .A1(n13730), .A2(n15296), .ZN(n15392) );
NOR2_X2 U14810 ( .A1(n13724), .A2(n15296), .ZN(n15416) );
NOR2_X2 U14811 ( .A1(n13718), .A2(n15296), .ZN(n15440) );
NOR2_X2 U14812 ( .A1(n13712), .A2(n15296), .ZN(n15464) );
NOR2_X2 U14813 ( .A1(n13706), .A2(n15492), .ZN(n15489) );
NOR2_X2 U14814 ( .A1(n13700), .A2(n15492), .ZN(n15518) );
NOR2_X2 U14815 ( .A1(n13694), .A2(n15492), .ZN(n15539) );
NOR2_X2 U14816 ( .A1(n13688), .A2(n15492), .ZN(n15560) );
NOR2_X2 U14817 ( .A1(n13682), .A2(n15492), .ZN(n15581) );
NOR2_X2 U14818 ( .A1(n13946), .A2(n14587), .ZN(n14585) );
NOR2_X2 U14819 ( .A1(n13940), .A2(n14587), .ZN(n14607) );
NOR2_X2 U14820 ( .A1(n13934), .A2(n14587), .ZN(n14628) );
NOR2_X2 U14821 ( .A1(n13928), .A2(n14587), .ZN(n14649) );
NOR2_X2 U14822 ( .A1(n13922), .A2(n14587), .ZN(n14670) );
NOR2_X2 U14823 ( .A1(n13916), .A2(n14587), .ZN(n14691) );
NOR2_X2 U14824 ( .A1(n13910), .A2(n14587), .ZN(n14712) );
NOR2_X2 U14825 ( .A1(n13904), .A2(n14587), .ZN(n14733) );
NOR2_X2 U14826 ( .A1(n13850), .A2(n14937), .ZN(n14935) );
NOR2_X2 U14827 ( .A1(n13844), .A2(n14937), .ZN(n14959) );
NOR2_X2 U14828 ( .A1(n13838), .A2(n14937), .ZN(n14981) );
NOR2_X2 U14829 ( .A1(n13832), .A2(n14937), .ZN(n15003) );
NOR2_X2 U14830 ( .A1(n13826), .A2(n14937), .ZN(n15025) );
NOR2_X2 U14831 ( .A1(n13820), .A2(n14937), .ZN(n15047) );
NOR2_X2 U14832 ( .A1(n13814), .A2(n14937), .ZN(n15069) );
NOR2_X2 U14833 ( .A1(n13808), .A2(n14937), .ZN(n15091) );
NOR2_X2 U14834 ( .A1(n13994), .A2(n14406), .ZN(n14404) );
NOR2_X2 U14835 ( .A1(n13988), .A2(n14406), .ZN(n14429) );
NOR2_X2 U14836 ( .A1(n13982), .A2(n14406), .ZN(n14451) );
NOR2_X2 U14837 ( .A1(n13976), .A2(n14406), .ZN(n14473) );
NOR2_X2 U14838 ( .A1(n13970), .A2(n14406), .ZN(n14495) );
NOR2_X2 U14839 ( .A1(n13964), .A2(n14406), .ZN(n14517) );
NOR2_X2 U14840 ( .A1(n13958), .A2(n14406), .ZN(n14539) );
NOR2_X2 U14841 ( .A1(n13952), .A2(n14406), .ZN(n14561) );
NOR2_X2 U14842 ( .A1(n13676), .A2(n15492), .ZN(n15602) );
NOR2_X2 U14843 ( .A1(n13669), .A2(n15492), .ZN(n15621) );
NOR2_X2 U14844 ( .A1(n13662), .A2(n15492), .ZN(n15640) );
NOR2_X2 U14845 ( .A1(n16209), .A2(n13462), .ZN(n16221) );
NOR2_X2 U14846 ( .A1(n16209), .A2(n13456), .ZN(n16235) );
NOR2_X2 U14847 ( .A1(n16209), .A2(n13450), .ZN(n16249) );
NOR2_X2 U14848 ( .A1(n16209), .A2(n13444), .ZN(n16263) );
NOR2_X2 U14849 ( .A1(n16209), .A2(n13438), .ZN(n16277) );
NOR2_X2 U14850 ( .A1(n16209), .A2(n13432), .ZN(n16291) );
NOR2_X2 U14851 ( .A1(n16209), .A2(n13426), .ZN(n16305) );
NOR2_X2 U14852 ( .A1(n16209), .A2(n13420), .ZN(n16319) );
NOR2_X2 U14853 ( .A1(n15663), .A2(n13654), .ZN(n15660) );
NOR2_X2 U14854 ( .A1(n15663), .A2(n13648), .ZN(n15680) );
NOR2_X2 U14855 ( .A1(n15663), .A2(n13642), .ZN(n15699) );
NOR2_X2 U14856 ( .A1(n15663), .A2(n13636), .ZN(n15718) );
NOR2_X2 U14857 ( .A1(n15663), .A2(n13630), .ZN(n15737) );
NOR2_X2 U14858 ( .A1(n15663), .A2(n13624), .ZN(n15756) );
NOR2_X2 U14859 ( .A1(n15663), .A2(n13618), .ZN(n15775) );
NOR2_X2 U14860 ( .A1(n15663), .A2(n13612), .ZN(n15794) );
NOR2_X2 U14861 ( .A1(n13558), .A2(n15946), .ZN(n15961) );
NOR2_X2 U14862 ( .A1(n13552), .A2(n15946), .ZN(n15978) );
NOR2_X2 U14863 ( .A1(n13546), .A2(n15946), .ZN(n15995) );
NOR2_X2 U14864 ( .A1(n13540), .A2(n15946), .ZN(n16012) );
NOR2_X2 U14865 ( .A1(n13534), .A2(n15946), .ZN(n16029) );
NOR2_X2 U14866 ( .A1(n13528), .A2(n15946), .ZN(n16046) );
NOR2_X2 U14867 ( .A1(n13522), .A2(n15946), .ZN(n16063) );
NOR2_X2 U14868 ( .A1(n13516), .A2(n15946), .ZN(n16080) );
AND2_X2 U14869 ( .A1(n17892), .A2(n15309), .ZN(n17756) );
NOR2_X2 U14870 ( .A1(n19191), .A2(n17905), .ZN(n16546) );
NOR2_X2 U14871 ( .A1(n19192), .A2(n17905), .ZN(n16551) );
NOR2_X2 U14872 ( .A1(n19193), .A2(n17905), .ZN(n16556) );
NOR2_X2 U14873 ( .A1(n19194), .A2(n17905), .ZN(n16561) );
NOR2_X2 U14874 ( .A1(n19195), .A2(n17905), .ZN(n16566) );
INV_X4 U14875 ( .A(n14414), .ZN(n17891) );
NOR2_X2 U14876 ( .A1(n18037), .A2(n16436), .ZN(N3086) );
NAND3_X2 U14877 ( .A1(n16438), .A2(n16439), .A3(n16440), .ZN(n16437) );
NOR2_X2 U14878 ( .A1(n18037), .A2(n16451), .ZN(N3085) );
NAND3_X2 U14879 ( .A1(n16453), .A2(n16454), .A3(n16455), .ZN(n16452) );
NOR2_X2 U14880 ( .A1(n18037), .A2(n16464), .ZN(N3084) );
NAND3_X2 U14881 ( .A1(n16466), .A2(n16467), .A3(n16468), .ZN(n16465) );
NOR2_X2 U14882 ( .A1(n18036), .A2(n16477), .ZN(N3083) );
NAND3_X2 U14883 ( .A1(n16479), .A2(n16480), .A3(n16481), .ZN(n16478) );
NOR2_X2 U14884 ( .A1(n18036), .A2(n16490), .ZN(N3082) );
NAND3_X2 U14885 ( .A1(n16492), .A2(n16493), .A3(n16494), .ZN(n16491) );
NOR2_X2 U14886 ( .A1(n18036), .A2(n16503), .ZN(N3081) );
NAND3_X2 U14887 ( .A1(n16505), .A2(n16506), .A3(n16507), .ZN(n16504) );
NOR2_X2 U14888 ( .A1(n18036), .A2(n16516), .ZN(N3080) );
NAND3_X2 U14889 ( .A1(n16518), .A2(n16519), .A3(n16520), .ZN(n16517) );
NOR2_X2 U14890 ( .A1(n18036), .A2(n16529), .ZN(N3079) );
NAND3_X2 U14891 ( .A1(n16531), .A2(n16532), .A3(n16533), .ZN(n16530) );
NOR2_X2 U14892 ( .A1(n19203), .A2(n11946), .ZN(n14167) );
NOR2_X2 U14893 ( .A1(n18075), .A2(n18071), .ZN(n14422) );
INV_X4 U14894 ( .A(n17775), .ZN(n17897) );
NOR4_X2 U14895 ( .A1(n14180), .A2(n14181), .A3(n14182), .A4(n14183), .ZN(n14179) );
NOR2_X2 U14896 ( .A1(n19135), .A2(n17860), .ZN(n14183) );
NOR2_X2 U14897 ( .A1(n19143), .A2(n14187), .ZN(n14180) );
NOR2_X2 U14898 ( .A1(n14185), .A2(n14186), .ZN(n14181) );
NOR4_X2 U14899 ( .A1(n14212), .A2(n14213), .A3(n14214), .A4(n14215), .ZN(n14211) );
NOR2_X2 U14900 ( .A1(n19136), .A2(n17860), .ZN(n14215) );
NOR2_X2 U14901 ( .A1(n19144), .A2(n14187), .ZN(n14212) );
NOR2_X2 U14902 ( .A1(n14216), .A2(n14186), .ZN(n14213) );
NOR4_X2 U14903 ( .A1(n14241), .A2(n14242), .A3(n14243), .A4(n14244), .ZN(n14240) );
NOR2_X2 U14904 ( .A1(n19137), .A2(n17860), .ZN(n14244) );
NOR2_X2 U14905 ( .A1(n19145), .A2(n14187), .ZN(n14241) );
NOR2_X2 U14906 ( .A1(n14245), .A2(n14186), .ZN(n14242) );
NOR4_X2 U14907 ( .A1(n14270), .A2(n14271), .A3(n14272), .A4(n14273), .ZN(n14269) );
NOR2_X2 U14908 ( .A1(n19138), .A2(n17860), .ZN(n14273) );
NOR2_X2 U14909 ( .A1(n19146), .A2(n14187), .ZN(n14270) );
NOR2_X2 U14910 ( .A1(n14274), .A2(n14186), .ZN(n14271) );
NOR4_X2 U14911 ( .A1(n14299), .A2(n14300), .A3(n14301), .A4(n14302), .ZN(n14298) );
NOR2_X2 U14912 ( .A1(n19139), .A2(n17860), .ZN(n14302) );
NOR2_X2 U14913 ( .A1(n19147), .A2(n14187), .ZN(n14299) );
NOR2_X2 U14914 ( .A1(n14303), .A2(n14186), .ZN(n14300) );
NOR4_X2 U14915 ( .A1(n14328), .A2(n14329), .A3(n14330), .A4(n14331), .ZN(n14327) );
NOR2_X2 U14916 ( .A1(n19140), .A2(n17860), .ZN(n14331) );
NOR2_X2 U14917 ( .A1(n19148), .A2(n14187), .ZN(n14328) );
NOR2_X2 U14918 ( .A1(n14332), .A2(n14186), .ZN(n14329) );
NOR4_X2 U14919 ( .A1(n14357), .A2(n14358), .A3(n14359), .A4(n14360), .ZN(n14356) );
NOR2_X2 U14920 ( .A1(n19141), .A2(n17860), .ZN(n14360) );
NOR2_X2 U14921 ( .A1(n19149), .A2(n14187), .ZN(n14357) );
NOR2_X2 U14922 ( .A1(n14361), .A2(n14186), .ZN(n14358) );
NOR4_X2 U14923 ( .A1(n14386), .A2(n14387), .A3(n14388), .A4(n14389), .ZN(n14385) );
NOR2_X2 U14924 ( .A1(n19142), .A2(n17860), .ZN(n14389) );
NOR2_X2 U14925 ( .A1(n19150), .A2(n14187), .ZN(n14386) );
NOR2_X2 U14926 ( .A1(n14391), .A2(n14186), .ZN(n14387) );
NOR4_X2 U14927 ( .A1(n15610), .A2(n15611), .A3(n15612), .A4(n15613), .ZN(n15609) );
NOR2_X2 U14928 ( .A1(n19148), .A2(n15507), .ZN(n15610) );
NOR2_X2 U14929 ( .A1(n19156), .A2(n15508), .ZN(n15611) );
NOR2_X2 U14930 ( .A1(n19180), .A2(n17869), .ZN(n15612) );
NOR4_X2 U14931 ( .A1(n15629), .A2(n15630), .A3(n15631), .A4(n15632), .ZN(n15628) );
NOR2_X2 U14932 ( .A1(n19149), .A2(n15507), .ZN(n15629) );
NOR2_X2 U14933 ( .A1(n19157), .A2(n15508), .ZN(n15630) );
NOR2_X2 U14934 ( .A1(n19181), .A2(n17869), .ZN(n15631) );
NOR4_X2 U14935 ( .A1(n15649), .A2(n15650), .A3(n15651), .A4(n15652), .ZN(n15648) );
NOR2_X2 U14936 ( .A1(n19150), .A2(n15507), .ZN(n15649) );
NOR2_X2 U14937 ( .A1(n19158), .A2(n15508), .ZN(n15650) );
NOR2_X2 U14938 ( .A1(n19182), .A2(n17869), .ZN(n15651) );
NOR4_X2 U14939 ( .A1(n15668), .A2(n15669), .A3(n15670), .A4(n15671), .ZN(n15667) );
NOR2_X2 U14940 ( .A1(n19191), .A2(n15504), .ZN(n15668) );
NOR2_X2 U14941 ( .A1(n19183), .A2(n17869), .ZN(n15669) );
NOR2_X2 U14942 ( .A1(n19175), .A2(n17870), .ZN(n15670) );
NOR4_X2 U14943 ( .A1(n15687), .A2(n15688), .A3(n15689), .A4(n15690), .ZN(n15686) );
NOR2_X2 U14944 ( .A1(n19192), .A2(n15504), .ZN(n15687) );
NOR2_X2 U14945 ( .A1(n19184), .A2(n17869), .ZN(n15688) );
NOR2_X2 U14946 ( .A1(n19176), .A2(n17870), .ZN(n15689) );
NOR4_X2 U14947 ( .A1(n15706), .A2(n15707), .A3(n15708), .A4(n15709), .ZN(n15705) );
NOR2_X2 U14948 ( .A1(n19193), .A2(n15504), .ZN(n15706) );
NOR2_X2 U14949 ( .A1(n19185), .A2(n17869), .ZN(n15707) );
NOR2_X2 U14950 ( .A1(n19177), .A2(n17870), .ZN(n15708) );
NOR4_X2 U14951 ( .A1(n15725), .A2(n15726), .A3(n15727), .A4(n15728), .ZN(n15724) );
NOR2_X2 U14952 ( .A1(n19194), .A2(n15504), .ZN(n15725) );
NOR2_X2 U14953 ( .A1(n19186), .A2(n17869), .ZN(n15726) );
NOR2_X2 U14954 ( .A1(n19178), .A2(n17870), .ZN(n15727) );
NOR4_X2 U14955 ( .A1(n15744), .A2(n15745), .A3(n15746), .A4(n15747), .ZN(n15743) );
NOR2_X2 U14956 ( .A1(n19195), .A2(n15504), .ZN(n15744) );
NOR2_X2 U14957 ( .A1(n19187), .A2(n17868), .ZN(n15745) );
NOR2_X2 U14958 ( .A1(n19179), .A2(n17870), .ZN(n15746) );
NOR4_X2 U14959 ( .A1(n15763), .A2(n15764), .A3(n15765), .A4(n15766), .ZN(n15762) );
NOR2_X2 U14960 ( .A1(n19196), .A2(n15504), .ZN(n15763) );
NOR2_X2 U14961 ( .A1(n19188), .A2(n17868), .ZN(n15764) );
NOR2_X2 U14962 ( .A1(n19180), .A2(n17871), .ZN(n15765) );
NOR4_X2 U14963 ( .A1(n15782), .A2(n15783), .A3(n15784), .A4(n15785), .ZN(n15781) );
NOR2_X2 U14964 ( .A1(n19197), .A2(n15504), .ZN(n15782) );
NOR2_X2 U14965 ( .A1(n19189), .A2(n17868), .ZN(n15783) );
NOR2_X2 U14966 ( .A1(n19181), .A2(n17871), .ZN(n15784) );
NOR4_X2 U14967 ( .A1(n15801), .A2(n15802), .A3(n15803), .A4(n15804), .ZN(n15800) );
NOR2_X2 U14968 ( .A1(n19198), .A2(n15504), .ZN(n15801) );
NOR2_X2 U14969 ( .A1(n19190), .A2(n17868), .ZN(n15802) );
NOR2_X2 U14970 ( .A1(n19182), .A2(n17871), .ZN(n15803) );
NOR4_X2 U14971 ( .A1(n15497), .A2(n15498), .A3(n15499), .A4(n15500), .ZN(n15496) );
NOR2_X2 U14972 ( .A1(n19183), .A2(n15504), .ZN(n15497) );
NOR2_X2 U14973 ( .A1(n19175), .A2(n17869), .ZN(n15498) );
NOR2_X2 U14974 ( .A1(n19167), .A2(n17871), .ZN(n15499) );
NOR4_X2 U14975 ( .A1(n15525), .A2(n15526), .A3(n15527), .A4(n15528), .ZN(n15524) );
NOR2_X2 U14976 ( .A1(n19184), .A2(n15504), .ZN(n15525) );
NOR2_X2 U14977 ( .A1(n19176), .A2(n17869), .ZN(n15526) );
NOR2_X2 U14978 ( .A1(n19168), .A2(n17870), .ZN(n15527) );
NOR4_X2 U14979 ( .A1(n15546), .A2(n15547), .A3(n15548), .A4(n15549), .ZN(n15545) );
NOR2_X2 U14980 ( .A1(n19185), .A2(n15504), .ZN(n15546) );
NOR2_X2 U14981 ( .A1(n19177), .A2(n17869), .ZN(n15547) );
NOR2_X2 U14982 ( .A1(n19169), .A2(n17870), .ZN(n15548) );
NOR4_X2 U14983 ( .A1(n15567), .A2(n15568), .A3(n15569), .A4(n15570), .ZN(n15566) );
NOR2_X2 U14984 ( .A1(n19186), .A2(n15504), .ZN(n15567) );
NOR2_X2 U14985 ( .A1(n19178), .A2(n17869), .ZN(n15568) );
NOR2_X2 U14986 ( .A1(n19170), .A2(n17870), .ZN(n15569) );
NOR4_X2 U14987 ( .A1(n15588), .A2(n15589), .A3(n15590), .A4(n15591), .ZN(n15587) );
NOR2_X2 U14988 ( .A1(n19187), .A2(n15504), .ZN(n15588) );
NOR2_X2 U14989 ( .A1(n19179), .A2(n17869), .ZN(n15589) );
NOR2_X2 U14990 ( .A1(n19171), .A2(n17870), .ZN(n15590) );
NAND3_X2 U14991 ( .A1(n14418), .A2(n14419), .A3(n14420), .ZN(n14190) );
NAND3_X2 U14992 ( .A1(n14441), .A2(n14442), .A3(n14443), .ZN(n14219) );
NAND3_X2 U14993 ( .A1(n14463), .A2(n14464), .A3(n14465), .ZN(n14248) );
NAND3_X2 U14994 ( .A1(n14485), .A2(n14486), .A3(n14487), .ZN(n14277) );
NAND3_X2 U14995 ( .A1(n14507), .A2(n14508), .A3(n14509), .ZN(n14306) );
NAND3_X2 U14996 ( .A1(n14529), .A2(n14530), .A3(n14531), .ZN(n14335) );
NAND3_X2 U14997 ( .A1(n14551), .A2(n14552), .A3(n14553), .ZN(n14364) );
NAND3_X2 U14998 ( .A1(n14575), .A2(n14576), .A3(n14577), .ZN(n14396) );
NOR2_X2 U14999 ( .A1(n19167), .A2(n14184), .ZN(n14182) );
NOR2_X2 U15000 ( .A1(n19168), .A2(n14184), .ZN(n14214) );
NOR2_X2 U15001 ( .A1(n19169), .A2(n14184), .ZN(n14243) );
NOR2_X2 U15002 ( .A1(n19170), .A2(n14184), .ZN(n14272) );
NOR2_X2 U15003 ( .A1(n19171), .A2(n14184), .ZN(n14301) );
NOR2_X2 U15004 ( .A1(n19172), .A2(n14184), .ZN(n14330) );
NOR2_X2 U15005 ( .A1(n19173), .A2(n14184), .ZN(n14359) );
NOR2_X2 U15006 ( .A1(n19174), .A2(n14184), .ZN(n14388) );
INV_X4 U15007 ( .A(n18075), .ZN(n18074) );
NOR2_X2 U15008 ( .A1(n19159), .A2(n17875), .ZN(n15500) );
NOR2_X2 U15009 ( .A1(n19160), .A2(n17874), .ZN(n15528) );
NOR2_X2 U15010 ( .A1(n19161), .A2(n17874), .ZN(n15549) );
NOR2_X2 U15011 ( .A1(n19162), .A2(n17874), .ZN(n15570) );
NOR2_X2 U15012 ( .A1(n19163), .A2(n17874), .ZN(n15591) );
NOR2_X2 U15013 ( .A1(n19164), .A2(n17874), .ZN(n15613) );
NOR2_X2 U15014 ( .A1(n19165), .A2(n17874), .ZN(n15632) );
NOR2_X2 U15015 ( .A1(n19166), .A2(n17874), .ZN(n15652) );
NOR2_X2 U15016 ( .A1(n19167), .A2(n17874), .ZN(n15671) );
NOR2_X2 U15017 ( .A1(n19168), .A2(n17874), .ZN(n15690) );
NOR2_X2 U15018 ( .A1(n19169), .A2(n17874), .ZN(n15709) );
NOR2_X2 U15019 ( .A1(n19170), .A2(n17874), .ZN(n15728) );
NOR2_X2 U15020 ( .A1(n19171), .A2(n17875), .ZN(n15747) );
NOR2_X2 U15021 ( .A1(n19172), .A2(n17875), .ZN(n15766) );
NOR2_X2 U15022 ( .A1(n19173), .A2(n17875), .ZN(n15785) );
NOR2_X2 U15023 ( .A1(n19174), .A2(n17875), .ZN(n15804) );
NAND2_X2 U15024 ( .A1(n14564), .A2(n15309), .ZN(n15504) );
NOR3_X2 U15025 ( .A1(n15915), .A2(n15916), .A3(n15917), .ZN(n15914) );
NOR2_X2 U15026 ( .A1(n19188), .A2(n17871), .ZN(n15917) );
NOR2_X2 U15027 ( .A1(n19196), .A2(n17868), .ZN(n15916) );
NOR2_X2 U15028 ( .A1(n19180), .A2(n17875), .ZN(n15915) );
NOR3_X2 U15029 ( .A1(n15825), .A2(n15826), .A3(n15827), .ZN(n15824) );
NOR2_X2 U15030 ( .A1(n19183), .A2(n17871), .ZN(n15827) );
NOR2_X2 U15031 ( .A1(n19191), .A2(n17868), .ZN(n15826) );
NOR2_X2 U15032 ( .A1(n19175), .A2(n17875), .ZN(n15825) );
NOR3_X2 U15033 ( .A1(n15843), .A2(n15844), .A3(n15845), .ZN(n15842) );
NOR2_X2 U15034 ( .A1(n19184), .A2(n17871), .ZN(n15845) );
NOR2_X2 U15035 ( .A1(n19192), .A2(n17868), .ZN(n15844) );
NOR2_X2 U15036 ( .A1(n19176), .A2(n17875), .ZN(n15843) );
NOR3_X2 U15037 ( .A1(n15861), .A2(n15862), .A3(n15863), .ZN(n15860) );
NOR2_X2 U15038 ( .A1(n19185), .A2(n17871), .ZN(n15863) );
NOR2_X2 U15039 ( .A1(n19193), .A2(n17868), .ZN(n15862) );
NOR2_X2 U15040 ( .A1(n19177), .A2(n17875), .ZN(n15861) );
NOR3_X2 U15041 ( .A1(n15879), .A2(n15880), .A3(n15881), .ZN(n15878) );
NOR2_X2 U15042 ( .A1(n19186), .A2(n17871), .ZN(n15881) );
NOR2_X2 U15043 ( .A1(n19194), .A2(n17868), .ZN(n15880) );
NOR2_X2 U15044 ( .A1(n19178), .A2(n17875), .ZN(n15879) );
NOR3_X2 U15045 ( .A1(n15897), .A2(n15898), .A3(n15899), .ZN(n15896) );
NOR2_X2 U15046 ( .A1(n19187), .A2(n17871), .ZN(n15899) );
NOR2_X2 U15047 ( .A1(n19195), .A2(n17868), .ZN(n15898) );
NOR2_X2 U15048 ( .A1(n19179), .A2(n17875), .ZN(n15897) );
NOR3_X2 U15049 ( .A1(n15933), .A2(n15934), .A3(n15935), .ZN(n15932) );
NOR2_X2 U15050 ( .A1(n19189), .A2(n17871), .ZN(n15935) );
NOR2_X2 U15051 ( .A1(n19197), .A2(n17868), .ZN(n15934) );
NOR2_X2 U15052 ( .A1(n19181), .A2(n17875), .ZN(n15933) );
NOR3_X2 U15053 ( .A1(n15953), .A2(n15954), .A3(n15955), .ZN(n15952) );
NOR2_X2 U15054 ( .A1(n19190), .A2(n17871), .ZN(n15955) );
NOR2_X2 U15055 ( .A1(n19198), .A2(n17868), .ZN(n15954) );
NOR2_X2 U15056 ( .A1(n19182), .A2(n17876), .ZN(n15953) );
NOR3_X2 U15057 ( .A1(n15304), .A2(n15305), .A3(n15306), .ZN(n15303) );
NOR2_X2 U15058 ( .A1(n15127), .A2(n17891), .ZN(n15304) );
NOR2_X2 U15059 ( .A1(n19183), .A2(n17864), .ZN(n15306) );
NOR2_X2 U15060 ( .A1(n19151), .A2(n17878), .ZN(n15305) );
NOR3_X2 U15061 ( .A1(n15329), .A2(n15330), .A3(n15331), .ZN(n15328) );
NOR2_X2 U15062 ( .A1(n15149), .A2(n17891), .ZN(n15329) );
NOR2_X2 U15063 ( .A1(n19184), .A2(n17864), .ZN(n15331) );
NOR2_X2 U15064 ( .A1(n19152), .A2(n17878), .ZN(n15330) );
NOR3_X2 U15065 ( .A1(n15353), .A2(n15354), .A3(n15355), .ZN(n15352) );
NOR2_X2 U15066 ( .A1(n15171), .A2(n17891), .ZN(n15353) );
NOR2_X2 U15067 ( .A1(n19185), .A2(n17864), .ZN(n15355) );
NOR2_X2 U15068 ( .A1(n19153), .A2(n17878), .ZN(n15354) );
NOR3_X2 U15069 ( .A1(n15377), .A2(n15378), .A3(n15379), .ZN(n15376) );
NOR2_X2 U15070 ( .A1(n15193), .A2(n17891), .ZN(n15377) );
NOR2_X2 U15071 ( .A1(n19186), .A2(n17864), .ZN(n15379) );
NOR2_X2 U15072 ( .A1(n19154), .A2(n17878), .ZN(n15378) );
NOR3_X2 U15073 ( .A1(n15401), .A2(n15402), .A3(n15403), .ZN(n15400) );
NOR2_X2 U15074 ( .A1(n15215), .A2(n17891), .ZN(n15401) );
NOR2_X2 U15075 ( .A1(n19187), .A2(n17864), .ZN(n15403) );
NOR2_X2 U15076 ( .A1(n19155), .A2(n17878), .ZN(n15402) );
NOR3_X2 U15077 ( .A1(n15425), .A2(n15426), .A3(n15427), .ZN(n15424) );
NOR2_X2 U15078 ( .A1(n15237), .A2(n17891), .ZN(n15425) );
NOR2_X2 U15079 ( .A1(n19188), .A2(n17864), .ZN(n15427) );
NOR2_X2 U15080 ( .A1(n19156), .A2(n17878), .ZN(n15426) );
NOR3_X2 U15081 ( .A1(n15449), .A2(n15450), .A3(n15451), .ZN(n15448) );
NOR2_X2 U15082 ( .A1(n15259), .A2(n17891), .ZN(n15449) );
NOR2_X2 U15083 ( .A1(n19189), .A2(n17864), .ZN(n15451) );
NOR2_X2 U15084 ( .A1(n19157), .A2(n17878), .ZN(n15450) );
NOR3_X2 U15085 ( .A1(n15475), .A2(n15476), .A3(n15477), .ZN(n15474) );
NOR2_X2 U15086 ( .A1(n15283), .A2(n17891), .ZN(n15475) );
NOR2_X2 U15087 ( .A1(n19190), .A2(n17864), .ZN(n15477) );
NOR2_X2 U15088 ( .A1(n19158), .A2(n17878), .ZN(n15476) );
NOR2_X2 U15089 ( .A1(n19143), .A2(n17879), .ZN(n15125) );
NOR2_X2 U15090 ( .A1(n19144), .A2(n17879), .ZN(n15147) );
NOR2_X2 U15091 ( .A1(n19145), .A2(n17879), .ZN(n15169) );
NOR2_X2 U15092 ( .A1(n19146), .A2(n17879), .ZN(n15191) );
NOR2_X2 U15093 ( .A1(n19147), .A2(n17878), .ZN(n15213) );
NOR2_X2 U15094 ( .A1(n19148), .A2(n17878), .ZN(n15235) );
NOR2_X2 U15095 ( .A1(n19149), .A2(n17878), .ZN(n15257) );
NOR2_X2 U15096 ( .A1(n19150), .A2(n17878), .ZN(n15281) );
NOR2_X2 U15097 ( .A1(n15127), .A2(n17865), .ZN(n15124) );
NOR2_X2 U15098 ( .A1(n15149), .A2(n17865), .ZN(n15146) );
NOR2_X2 U15099 ( .A1(n15171), .A2(n17865), .ZN(n15168) );
NOR2_X2 U15100 ( .A1(n15193), .A2(n17865), .ZN(n15190) );
NOR2_X2 U15101 ( .A1(n15215), .A2(n17865), .ZN(n15212) );
NOR2_X2 U15102 ( .A1(n15237), .A2(n17865), .ZN(n15234) );
NOR2_X2 U15103 ( .A1(n15259), .A2(n17865), .ZN(n15256) );
NOR2_X2 U15104 ( .A1(n15283), .A2(n17865), .ZN(n15280) );
NOR2_X2 U15105 ( .A1(n19175), .A2(n17863), .ZN(n15126) );
NOR2_X2 U15106 ( .A1(n19176), .A2(n17863), .ZN(n15148) );
NOR2_X2 U15107 ( .A1(n19177), .A2(n17863), .ZN(n15170) );
NOR2_X2 U15108 ( .A1(n19178), .A2(n17863), .ZN(n15192) );
NOR2_X2 U15109 ( .A1(n19179), .A2(n17863), .ZN(n15214) );
NOR2_X2 U15110 ( .A1(n19180), .A2(n17863), .ZN(n15236) );
NOR2_X2 U15111 ( .A1(n19181), .A2(n17863), .ZN(n15258) );
NOR2_X2 U15112 ( .A1(n19182), .A2(n17863), .ZN(n15282) );
NOR2_X2 U15113 ( .A1(n19151), .A2(n15508), .ZN(n15505) );
NOR2_X2 U15114 ( .A1(n19152), .A2(n15508), .ZN(n15529) );
NOR2_X2 U15115 ( .A1(n19153), .A2(n15508), .ZN(n15550) );
NOR2_X2 U15116 ( .A1(n19154), .A2(n15508), .ZN(n15571) );
NOR2_X2 U15117 ( .A1(n19155), .A2(n15508), .ZN(n15592) );
NOR2_X2 U15118 ( .A1(n19196), .A2(n17864), .ZN(n15615) );
AND2_X2 U15119 ( .A1(n18071), .A2(n18075), .ZN(n17757) );
AND2_X2 U15120 ( .A1(n17897), .A2(n15309), .ZN(n17758) );
NOR2_X2 U15121 ( .A1(n19143), .A2(n15507), .ZN(n15506) );
NOR2_X2 U15122 ( .A1(n19144), .A2(n15507), .ZN(n15530) );
NOR2_X2 U15123 ( .A1(n19145), .A2(n15507), .ZN(n15551) );
NOR2_X2 U15124 ( .A1(n19146), .A2(n15507), .ZN(n15572) );
NOR2_X2 U15125 ( .A1(n19147), .A2(n15507), .ZN(n15593) );
NOR2_X2 U15126 ( .A1(n14415), .A2(n14416), .ZN(n14412) );
NOR2_X2 U15127 ( .A1(n17866), .A2(n14417), .ZN(n14416) );
NOR2_X2 U15128 ( .A1(n19143), .A2(n17860), .ZN(n14415) );
NOR2_X2 U15129 ( .A1(n14438), .A2(n14439), .ZN(n14436) );
NOR2_X2 U15130 ( .A1(n17866), .A2(n14440), .ZN(n14439) );
NOR2_X2 U15131 ( .A1(n19144), .A2(n17860), .ZN(n14438) );
NOR2_X2 U15132 ( .A1(n14460), .A2(n14461), .ZN(n14458) );
NOR2_X2 U15133 ( .A1(n17866), .A2(n14462), .ZN(n14461) );
NOR2_X2 U15134 ( .A1(n19145), .A2(n17860), .ZN(n14460) );
NOR2_X2 U15135 ( .A1(n14482), .A2(n14483), .ZN(n14480) );
NOR2_X2 U15136 ( .A1(n17866), .A2(n14484), .ZN(n14483) );
NOR2_X2 U15137 ( .A1(n19146), .A2(n17860), .ZN(n14482) );
NOR2_X2 U15138 ( .A1(n14504), .A2(n14505), .ZN(n14502) );
NOR2_X2 U15139 ( .A1(n17866), .A2(n14506), .ZN(n14505) );
NOR2_X2 U15140 ( .A1(n19147), .A2(n17861), .ZN(n14504) );
NOR2_X2 U15141 ( .A1(n14526), .A2(n14527), .ZN(n14524) );
NOR2_X2 U15142 ( .A1(n17866), .A2(n14528), .ZN(n14527) );
NOR2_X2 U15143 ( .A1(n19148), .A2(n17861), .ZN(n14526) );
NOR2_X2 U15144 ( .A1(n14548), .A2(n14549), .ZN(n14546) );
NOR2_X2 U15145 ( .A1(n17866), .A2(n14550), .ZN(n14549) );
NOR2_X2 U15146 ( .A1(n19149), .A2(n17861), .ZN(n14548) );
NOR2_X2 U15147 ( .A1(n14572), .A2(n14573), .ZN(n14570) );
NOR2_X2 U15148 ( .A1(n17866), .A2(n14574), .ZN(n14573) );
NOR2_X2 U15149 ( .A1(n19150), .A2(n17861), .ZN(n14572) );
NOR2_X2 U15150 ( .A1(n19189), .A2(n15504), .ZN(n15634) );
NOR2_X2 U15151 ( .A1(n19190), .A2(n15504), .ZN(n15654) );
NOR2_X2 U15152 ( .A1(n16088), .A2(n16089), .ZN(n16086) );
NOR2_X2 U15153 ( .A1(n19198), .A2(n17870), .ZN(n16088) );
NOR2_X2 U15154 ( .A1(n19190), .A2(n17874), .ZN(n16089) );
NOR2_X2 U15155 ( .A1(n19188), .A2(n15504), .ZN(n15614) );
NOR2_X2 U15156 ( .A1(n19173), .A2(n17870), .ZN(n15633) );
NOR2_X2 U15157 ( .A1(n19174), .A2(n17870), .ZN(n15653) );
NOR2_X2 U15158 ( .A1(n14595), .A2(n14596), .ZN(n14593) );
NOR2_X2 U15159 ( .A1(n17866), .A2(n14597), .ZN(n14596) );
NOR2_X2 U15160 ( .A1(n19151), .A2(n17861), .ZN(n14595) );
NOR2_X2 U15161 ( .A1(n14616), .A2(n14617), .ZN(n14614) );
NOR2_X2 U15162 ( .A1(n17867), .A2(n14618), .ZN(n14617) );
NOR2_X2 U15163 ( .A1(n19152), .A2(n17861), .ZN(n14616) );
NOR2_X2 U15164 ( .A1(n14637), .A2(n14638), .ZN(n14635) );
NOR2_X2 U15165 ( .A1(n17867), .A2(n14639), .ZN(n14638) );
NOR2_X2 U15166 ( .A1(n19153), .A2(n17861), .ZN(n14637) );
NOR2_X2 U15167 ( .A1(n14658), .A2(n14659), .ZN(n14656) );
NOR2_X2 U15168 ( .A1(n17867), .A2(n14660), .ZN(n14659) );
NOR2_X2 U15169 ( .A1(n19154), .A2(n17861), .ZN(n14658) );
NOR2_X2 U15170 ( .A1(n14679), .A2(n14680), .ZN(n14677) );
NOR2_X2 U15171 ( .A1(n17867), .A2(n14681), .ZN(n14680) );
NOR2_X2 U15172 ( .A1(n19155), .A2(n17861), .ZN(n14679) );
NOR2_X2 U15173 ( .A1(n14700), .A2(n14701), .ZN(n14698) );
NOR2_X2 U15174 ( .A1(n17867), .A2(n14702), .ZN(n14701) );
NOR2_X2 U15175 ( .A1(n19156), .A2(n17861), .ZN(n14700) );
NOR2_X2 U15176 ( .A1(n14721), .A2(n14722), .ZN(n14719) );
NOR2_X2 U15177 ( .A1(n17867), .A2(n14723), .ZN(n14722) );
NOR2_X2 U15178 ( .A1(n19157), .A2(n17861), .ZN(n14721) );
NOR2_X2 U15179 ( .A1(n14744), .A2(n14745), .ZN(n14742) );
NOR2_X2 U15180 ( .A1(n17867), .A2(n14746), .ZN(n14745) );
NOR2_X2 U15181 ( .A1(n19158), .A2(n17861), .ZN(n14744) );
NOR2_X2 U15182 ( .A1(n14766), .A2(n14767), .ZN(n14764) );
NOR2_X2 U15183 ( .A1(n17867), .A2(n14768), .ZN(n14767) );
NOR2_X2 U15184 ( .A1(n19159), .A2(n17862), .ZN(n14766) );
NOR2_X2 U15185 ( .A1(n14789), .A2(n14790), .ZN(n14787) );
NOR2_X2 U15186 ( .A1(n17867), .A2(n14791), .ZN(n14790) );
NOR2_X2 U15187 ( .A1(n19160), .A2(n17862), .ZN(n14789) );
NOR2_X2 U15188 ( .A1(n14811), .A2(n14812), .ZN(n14809) );
NOR2_X2 U15189 ( .A1(n17867), .A2(n14813), .ZN(n14812) );
NOR2_X2 U15190 ( .A1(n19161), .A2(n17862), .ZN(n14811) );
NOR2_X2 U15191 ( .A1(n14833), .A2(n14834), .ZN(n14831) );
NOR2_X2 U15192 ( .A1(n17867), .A2(n14835), .ZN(n14834) );
NOR2_X2 U15193 ( .A1(n19162), .A2(n17862), .ZN(n14833) );
NOR2_X2 U15194 ( .A1(n14855), .A2(n14856), .ZN(n14853) );
NOR2_X2 U15195 ( .A1(n17867), .A2(n14857), .ZN(n14856) );
NOR2_X2 U15196 ( .A1(n19163), .A2(n17862), .ZN(n14855) );
NOR2_X2 U15197 ( .A1(n14877), .A2(n14878), .ZN(n14875) );
NOR2_X2 U15198 ( .A1(n17867), .A2(n14879), .ZN(n14878) );
NOR2_X2 U15199 ( .A1(n19164), .A2(n17862), .ZN(n14877) );
NOR2_X2 U15200 ( .A1(n14899), .A2(n14900), .ZN(n14897) );
NOR2_X2 U15201 ( .A1(n17867), .A2(n14901), .ZN(n14900) );
NOR2_X2 U15202 ( .A1(n19165), .A2(n17862), .ZN(n14899) );
NOR2_X2 U15203 ( .A1(n14922), .A2(n14923), .ZN(n14920) );
NOR2_X2 U15204 ( .A1(n17866), .A2(n14924), .ZN(n14923) );
NOR2_X2 U15205 ( .A1(n19166), .A2(n17862), .ZN(n14922) );
NAND3_X2 U15206 ( .A1(n14598), .A2(n14599), .A3(n14600), .ZN(n14191) );
NAND3_X2 U15207 ( .A1(n14619), .A2(n14620), .A3(n14621), .ZN(n14220) );
NAND3_X2 U15208 ( .A1(n14640), .A2(n14641), .A3(n14642), .ZN(n14249) );
NAND3_X2 U15209 ( .A1(n14661), .A2(n14662), .A3(n14663), .ZN(n14278) );
NAND3_X2 U15210 ( .A1(n14682), .A2(n14683), .A3(n14684), .ZN(n14307) );
NAND3_X2 U15211 ( .A1(n14703), .A2(n14704), .A3(n14705), .ZN(n14336) );
NAND3_X2 U15212 ( .A1(n14724), .A2(n14725), .A3(n14726), .ZN(n14365) );
NAND3_X2 U15213 ( .A1(n14747), .A2(n14748), .A3(n14749), .ZN(n14397) );
NAND3_X2 U15214 ( .A1(n15121), .A2(n15122), .A3(n15123), .ZN(n15118) );
NOR3_X2 U15215 ( .A1(n15124), .A2(n15125), .A3(n15126), .ZN(n15123) );
NAND3_X2 U15216 ( .A1(n15143), .A2(n15144), .A3(n15145), .ZN(n15140) );
NOR3_X2 U15217 ( .A1(n15146), .A2(n15147), .A3(n15148), .ZN(n15145) );
NAND3_X2 U15218 ( .A1(n15165), .A2(n15166), .A3(n15167), .ZN(n15162) );
NOR3_X2 U15219 ( .A1(n15168), .A2(n15169), .A3(n15170), .ZN(n15167) );
NAND3_X2 U15220 ( .A1(n15187), .A2(n15188), .A3(n15189), .ZN(n15184) );
NOR3_X2 U15221 ( .A1(n15190), .A2(n15191), .A3(n15192), .ZN(n15189) );
NAND3_X2 U15222 ( .A1(n15209), .A2(n15210), .A3(n15211), .ZN(n15206) );
NOR3_X2 U15223 ( .A1(n15212), .A2(n15213), .A3(n15214), .ZN(n15211) );
NAND3_X2 U15224 ( .A1(n15231), .A2(n15232), .A3(n15233), .ZN(n15228) );
NOR3_X2 U15225 ( .A1(n15234), .A2(n15235), .A3(n15236), .ZN(n15233) );
NAND3_X2 U15226 ( .A1(n15253), .A2(n15254), .A3(n15255), .ZN(n15250) );
NOR3_X2 U15227 ( .A1(n15256), .A2(n15257), .A3(n15258), .ZN(n15255) );
NAND3_X2 U15228 ( .A1(n15277), .A2(n15278), .A3(n15279), .ZN(n15274) );
NOR3_X2 U15229 ( .A1(n15280), .A2(n15281), .A3(n15282), .ZN(n15279) );
NOR2_X2 U15230 ( .A1(n14946), .A2(n14947), .ZN(n14943) );
NOR2_X2 U15231 ( .A1(n19167), .A2(n17862), .ZN(n14947) );
NOR2_X2 U15232 ( .A1(n19135), .A2(n17879), .ZN(n14946) );
NOR2_X2 U15233 ( .A1(n14969), .A2(n14970), .ZN(n14966) );
NOR2_X2 U15234 ( .A1(n19168), .A2(n17862), .ZN(n14970) );
NOR2_X2 U15235 ( .A1(n19136), .A2(n17879), .ZN(n14969) );
NOR2_X2 U15236 ( .A1(n14991), .A2(n14992), .ZN(n14988) );
NOR2_X2 U15237 ( .A1(n19169), .A2(n17862), .ZN(n14992) );
NOR2_X2 U15238 ( .A1(n19137), .A2(n17879), .ZN(n14991) );
NOR2_X2 U15239 ( .A1(n15013), .A2(n15014), .ZN(n15010) );
NOR2_X2 U15240 ( .A1(n19170), .A2(n17862), .ZN(n15014) );
NOR2_X2 U15241 ( .A1(n19138), .A2(n17879), .ZN(n15013) );
NOR2_X2 U15242 ( .A1(n15035), .A2(n15036), .ZN(n15032) );
NOR2_X2 U15243 ( .A1(n19171), .A2(n17863), .ZN(n15036) );
NOR2_X2 U15244 ( .A1(n19139), .A2(n17879), .ZN(n15035) );
NOR2_X2 U15245 ( .A1(n15079), .A2(n15080), .ZN(n15076) );
NOR2_X2 U15246 ( .A1(n19173), .A2(n17863), .ZN(n15080) );
NOR2_X2 U15247 ( .A1(n19141), .A2(n17879), .ZN(n15079) );
NOR2_X2 U15248 ( .A1(n15103), .A2(n15104), .ZN(n15100) );
NOR2_X2 U15249 ( .A1(n19174), .A2(n17863), .ZN(n15104) );
NOR2_X2 U15250 ( .A1(n19142), .A2(n17879), .ZN(n15103) );
NOR2_X2 U15251 ( .A1(n15057), .A2(n15058), .ZN(n15054) );
NOR2_X2 U15252 ( .A1(n19172), .A2(n17863), .ZN(n15058) );
NOR2_X2 U15253 ( .A1(n19140), .A2(n17879), .ZN(n15057) );
INV_X4 U15254 ( .A(n17289), .ZN(n17958) );
NOR2_X2 U15255 ( .A1(n16053), .A2(n16054), .ZN(n16051) );
NOR2_X2 U15256 ( .A1(n19196), .A2(n17872), .ZN(n16053) );
NOR2_X2 U15257 ( .A1(n19188), .A2(n17876), .ZN(n16054) );
NOR2_X2 U15258 ( .A1(n15968), .A2(n15969), .ZN(n15966) );
NOR2_X2 U15259 ( .A1(n19191), .A2(n17872), .ZN(n15968) );
NOR2_X2 U15260 ( .A1(n19183), .A2(n17876), .ZN(n15969) );
NOR2_X2 U15261 ( .A1(n15985), .A2(n15986), .ZN(n15983) );
NOR2_X2 U15262 ( .A1(n19192), .A2(n17872), .ZN(n15985) );
NOR2_X2 U15263 ( .A1(n19184), .A2(n17876), .ZN(n15986) );
NOR2_X2 U15264 ( .A1(n16002), .A2(n16003), .ZN(n16000) );
NOR2_X2 U15265 ( .A1(n19193), .A2(n17872), .ZN(n16002) );
NOR2_X2 U15266 ( .A1(n19185), .A2(n17876), .ZN(n16003) );
NOR2_X2 U15267 ( .A1(n16019), .A2(n16020), .ZN(n16017) );
NOR2_X2 U15268 ( .A1(n19194), .A2(n17872), .ZN(n16019) );
NOR2_X2 U15269 ( .A1(n19186), .A2(n17876), .ZN(n16020) );
NOR2_X2 U15270 ( .A1(n16036), .A2(n16037), .ZN(n16034) );
NOR2_X2 U15271 ( .A1(n19195), .A2(n17872), .ZN(n16036) );
NOR2_X2 U15272 ( .A1(n19187), .A2(n17876), .ZN(n16037) );
NOR2_X2 U15273 ( .A1(n16070), .A2(n16071), .ZN(n16068) );
NOR2_X2 U15274 ( .A1(n19197), .A2(n17872), .ZN(n16070) );
NOR2_X2 U15275 ( .A1(n19189), .A2(n17876), .ZN(n16071) );
NOR2_X2 U15276 ( .A1(n18071), .A2(n18074), .ZN(n14393) );
INV_X4 U15277 ( .A(n17775), .ZN(n17898) );
INV_X4 U15278 ( .A(n17283), .ZN(n18002) );
INV_X4 U15279 ( .A(n17775), .ZN(n17899) );
BUF_X4 U15280 ( .A(n17752), .Z(n17823) );
BUF_X4 U15281 ( .A(n17753), .Z(n17822) );
BUF_X4 U15282 ( .A(n17818), .Z(n17821) );
BUF_X4 U15283 ( .A(n17751), .Z(n17820) );
BUF_X4 U15284 ( .A(n17752), .Z(n17819) );
BUF_X4 U15285 ( .A(n18632), .Z(n17835) );
BUF_X4 U15286 ( .A(n17753), .Z(n17834) );
BUF_X4 U15287 ( .A(n17752), .Z(n17833) );
BUF_X4 U15288 ( .A(n17751), .Z(n17832) );
BUF_X4 U15289 ( .A(n17826), .Z(n17831) );
BUF_X4 U15290 ( .A(n17751), .Z(n17830) );
BUF_X4 U15291 ( .A(n17752), .Z(n17829) );
BUF_X4 U15292 ( .A(n17753), .Z(n17828) );
BUF_X4 U15293 ( .A(n17830), .Z(n17827) );
BUF_X4 U15294 ( .A(n17751), .Z(n17826) );
BUF_X4 U15295 ( .A(n17752), .Z(n17825) );
BUF_X4 U15296 ( .A(n17753), .Z(n17824) );
BUF_X4 U15297 ( .A(n17751), .Z(n17818) );
BUF_X4 U15298 ( .A(n17752), .Z(n17836) );
NOR4_X2 U15299 ( .A1(n14157), .A2(state[0]), .A3(state[1]), .A4(state[4]),.ZN(n12235) );
NOR4_X2 U15300 ( .A1(n14402), .A2(n14403), .A3(n14404), .A4(n18743), .ZN(n14401) );
NOR4_X2 U15301 ( .A1(n14427), .A2(n14428), .A3(n14429), .A4(n18742), .ZN(n14426) );
NOR4_X2 U15302 ( .A1(n14449), .A2(n14450), .A3(n14451), .A4(n18741), .ZN(n14448) );
NOR4_X2 U15303 ( .A1(n14471), .A2(n14472), .A3(n14473), .A4(n18740), .ZN(n14470) );
NOR4_X2 U15304 ( .A1(n14493), .A2(n14494), .A3(n14495), .A4(n18739), .ZN(n14492) );
NOR4_X2 U15305 ( .A1(n14515), .A2(n14516), .A3(n14517), .A4(n18738), .ZN(n14514) );
NOR4_X2 U15306 ( .A1(n14537), .A2(n14538), .A3(n14539), .A4(n18737), .ZN(n14536) );
NOR4_X2 U15307 ( .A1(n14559), .A2(n14560), .A3(n14561), .A4(n18736), .ZN(n14558) );
NOR4_X2 U15308 ( .A1(n15814), .A2(n18682), .A3(n15815), .A4(n15816), .ZN(n15813) );
NOR2_X2 U15309 ( .A1(n19143), .A2(n17903), .ZN(n15815) );
NOR4_X2 U15310 ( .A1(n15832), .A2(n18681), .A3(n15833), .A4(n15834), .ZN(n15831) );
NOR2_X2 U15311 ( .A1(n19144), .A2(n17903), .ZN(n15833) );
NOR4_X2 U15312 ( .A1(n15850), .A2(n18680), .A3(n15851), .A4(n15852), .ZN(n15849) );
NOR2_X2 U15313 ( .A1(n19145), .A2(n17903), .ZN(n15851) );
NOR4_X2 U15314 ( .A1(n15868), .A2(n18679), .A3(n15869), .A4(n15870), .ZN(n15867) );
NOR2_X2 U15315 ( .A1(n5329), .A2(n18001), .ZN(n15870) );
NOR2_X2 U15316 ( .A1(n19146), .A2(n17903), .ZN(n15869) );
NOR4_X2 U15317 ( .A1(n15886), .A2(n18678), .A3(n15887), .A4(n15888), .ZN(n15885) );
NOR2_X2 U15318 ( .A1(n5330), .A2(n18000), .ZN(n15888) );
NOR2_X2 U15319 ( .A1(n19147), .A2(n17903), .ZN(n15887) );
NOR4_X2 U15320 ( .A1(n15904), .A2(n18677), .A3(n15905), .A4(n15906), .ZN(n15903) );
NOR2_X2 U15321 ( .A1(n5331), .A2(n18000), .ZN(n15906) );
NOR2_X2 U15322 ( .A1(n19148), .A2(n17903), .ZN(n15905) );
NOR4_X2 U15323 ( .A1(n15922), .A2(n18676), .A3(n15923), .A4(n15924), .ZN(n15921) );
NOR2_X2 U15324 ( .A1(n5332), .A2(n18000), .ZN(n15924) );
NOR2_X2 U15325 ( .A1(n19149), .A2(n17903), .ZN(n15923) );
NOR4_X2 U15326 ( .A1(n15940), .A2(n18675), .A3(n15941), .A4(n15942), .ZN(n15939) );
NOR2_X2 U15327 ( .A1(n5333), .A2(n18000), .ZN(n15942) );
NOR2_X2 U15328 ( .A1(n19150), .A2(n17903), .ZN(n15941) );
NOR4_X2 U15329 ( .A1(n16334), .A2(n18650), .A3(n16335), .A4(n16336), .ZN(n16333) );
NOR2_X2 U15330 ( .A1(n5358), .A2(n18001), .ZN(n16336) );
NOR2_X2 U15331 ( .A1(n19175), .A2(n17904), .ZN(n16335) );
NOR4_X2 U15332 ( .A1(n16347), .A2(n18649), .A3(n16348), .A4(n16349), .ZN(n16346) );
NOR2_X2 U15333 ( .A1(n5359), .A2(n18001), .ZN(n16349) );
NOR2_X2 U15334 ( .A1(n19176), .A2(n17904), .ZN(n16348) );
NOR4_X2 U15335 ( .A1(n16360), .A2(n18648), .A3(n16361), .A4(n16362), .ZN(n16359) );
NOR2_X2 U15336 ( .A1(n5360), .A2(n18001), .ZN(n16362) );
NOR2_X2 U15337 ( .A1(n19177), .A2(n17904), .ZN(n16361) );
NOR4_X2 U15338 ( .A1(n16373), .A2(n18647), .A3(n16374), .A4(n16375), .ZN(n16372) );
NOR2_X2 U15339 ( .A1(n5361), .A2(n18001), .ZN(n16375) );
NOR2_X2 U15340 ( .A1(n19178), .A2(n17904), .ZN(n16374) );
NOR4_X2 U15341 ( .A1(n16386), .A2(n18646), .A3(n16387), .A4(n16388), .ZN(n16385) );
NOR2_X2 U15342 ( .A1(n5362), .A2(n18001), .ZN(n16388) );
NOR2_X2 U15343 ( .A1(n19179), .A2(n17905), .ZN(n16387) );
NOR4_X2 U15344 ( .A1(n16399), .A2(n18645), .A3(n16400), .A4(n16401), .ZN(n16398) );
NOR2_X2 U15345 ( .A1(n5363), .A2(n18002), .ZN(n16401) );
NOR2_X2 U15346 ( .A1(n19180), .A2(n17905), .ZN(n16400) );
NOR4_X2 U15347 ( .A1(n16412), .A2(n18644), .A3(n16413), .A4(n16414), .ZN(n16411) );
NOR2_X2 U15348 ( .A1(n5364), .A2(n18002), .ZN(n16414) );
NOR2_X2 U15349 ( .A1(n19181), .A2(n17905), .ZN(n16413) );
NOR4_X2 U15350 ( .A1(n16425), .A2(n18643), .A3(n16426), .A4(n16427), .ZN(n16424) );
NOR2_X2 U15351 ( .A1(n5365), .A2(n18002), .ZN(n16427) );
NOR2_X2 U15352 ( .A1(n19182), .A2(n17905), .ZN(n16426) );
NOR4_X2 U15353 ( .A1(n15601), .A2(n15602), .A3(n15603), .A4(n15604), .ZN(n15600) );
NOR2_X2 U15354 ( .A1(n15605), .A2(n17918), .ZN(n15604) );
NOR4_X2 U15355 ( .A1(n15620), .A2(n15621), .A3(n15622), .A4(n15623), .ZN(n15619) );
NOR2_X2 U15356 ( .A1(n15624), .A2(n17918), .ZN(n15623) );
NOR4_X2 U15357 ( .A1(n15639), .A2(n15640), .A3(n15641), .A4(n15642), .ZN(n15638) );
NOR2_X2 U15358 ( .A1(n15643), .A2(n17918), .ZN(n15642) );
NOR4_X2 U15359 ( .A1(n16097), .A2(n18666), .A3(n16098), .A4(n16099), .ZN(n16096) );
NOR2_X2 U15360 ( .A1(n5342), .A2(n18000), .ZN(n16099) );
NOR2_X2 U15361 ( .A1(n19159), .A2(n17904), .ZN(n16098) );
NOR4_X2 U15362 ( .A1(n16113), .A2(n18665), .A3(n16114), .A4(n16115), .ZN(n16112) );
NOR2_X2 U15363 ( .A1(n5343), .A2(n18001), .ZN(n16115) );
NOR2_X2 U15364 ( .A1(n19160), .A2(n17904), .ZN(n16114) );
NOR4_X2 U15365 ( .A1(n16128), .A2(n18664), .A3(n16129), .A4(n16130), .ZN(n16127) );
NOR2_X2 U15366 ( .A1(n5344), .A2(n18001), .ZN(n16130) );
NOR2_X2 U15367 ( .A1(n19161), .A2(n17904), .ZN(n16129) );
NOR4_X2 U15368 ( .A1(n16143), .A2(n18663), .A3(n16144), .A4(n16145), .ZN(n16142) );
NOR2_X2 U15369 ( .A1(n5345), .A2(n18001), .ZN(n16145) );
NOR2_X2 U15370 ( .A1(n19162), .A2(n17904), .ZN(n16144) );
NOR4_X2 U15371 ( .A1(n16158), .A2(n18662), .A3(n16159), .A4(n16160), .ZN(n16157) );
NOR2_X2 U15372 ( .A1(n5346), .A2(n18001), .ZN(n16160) );
NOR2_X2 U15373 ( .A1(n19163), .A2(n17904), .ZN(n16159) );
NOR4_X2 U15374 ( .A1(n16173), .A2(n18661), .A3(n16174), .A4(n16175), .ZN(n16172) );
NOR2_X2 U15375 ( .A1(n5347), .A2(n18001), .ZN(n16175) );
NOR2_X2 U15376 ( .A1(n19164), .A2(n17904), .ZN(n16174) );
NOR4_X2 U15377 ( .A1(n16188), .A2(n18660), .A3(n16189), .A4(n16190), .ZN(n16187) );
NOR2_X2 U15378 ( .A1(n5348), .A2(n18001), .ZN(n16190) );
NOR2_X2 U15379 ( .A1(n19165), .A2(n17904), .ZN(n16189) );
NOR4_X2 U15380 ( .A1(n16203), .A2(n18659), .A3(n16204), .A4(n16205), .ZN(n16202) );
NOR2_X2 U15381 ( .A1(n5349), .A2(n18001), .ZN(n16205) );
NOR2_X2 U15382 ( .A1(n19166), .A2(n17904), .ZN(n16204) );
NOR2_X2 U15383 ( .A1(n18036), .A2(n16549), .ZN(N3077) );
NOR2_X2 U15384 ( .A1(n18036), .A2(n16554), .ZN(N3076) );
NOR2_X2 U15385 ( .A1(n18036), .A2(n16559), .ZN(N3075) );
NOR2_X2 U15386 ( .A1(n18036), .A2(n16564), .ZN(N3074) );
AND3_X2 U15387 ( .A1(n17759), .A2(n13364), .A3(n17760), .ZN(n16440) );
OR2_X4 U15388 ( .A1(n19191), .A2(n16450), .ZN(n17759) );
NAND3_X2 U15389 ( .A1(n18634), .A2(n13365), .A3(aes_text_out[15]), .ZN(n17760) );
AND3_X2 U15390 ( .A1(n17761), .A2(n13358), .A3(n17762), .ZN(n16455) );
OR2_X4 U15391 ( .A1(n19192), .A2(n16450), .ZN(n17761) );
NAND3_X2 U15392 ( .A1(n18634), .A2(n13359), .A3(aes_text_out[14]), .ZN(n17762) );
AND3_X2 U15393 ( .A1(n17763), .A2(n13352), .A3(n17764), .ZN(n16468) );
OR2_X4 U15394 ( .A1(n19193), .A2(n16450), .ZN(n17763) );
NAND3_X2 U15395 ( .A1(n18634), .A2(n13353), .A3(aes_text_out[13]), .ZN(n17764) );
AND3_X2 U15396 ( .A1(n17765), .A2(n13346), .A3(n17766), .ZN(n16481) );
OR2_X4 U15397 ( .A1(n19194), .A2(n16450), .ZN(n17765) );
NAND3_X2 U15398 ( .A1(n18634), .A2(n13347), .A3(aes_text_out[12]), .ZN(n17766) );
AND3_X2 U15399 ( .A1(n17767), .A2(n13340), .A3(n17768), .ZN(n16494) );
OR2_X4 U15400 ( .A1(n19195), .A2(n16450), .ZN(n17767) );
NAND3_X2 U15401 ( .A1(n18634), .A2(n13341), .A3(aes_text_out[11]), .ZN(n17768) );
AND3_X2 U15402 ( .A1(n17769), .A2(n13334), .A3(n17770), .ZN(n16507) );
OR2_X4 U15403 ( .A1(n19196), .A2(n16450), .ZN(n17769) );
NAND3_X2 U15404 ( .A1(n18634), .A2(n13335), .A3(aes_text_out[10]), .ZN(n17770) );
AND3_X2 U15405 ( .A1(n17771), .A2(n13328), .A3(n17772), .ZN(n16520) );
OR2_X4 U15406 ( .A1(n19197), .A2(n16450), .ZN(n17771) );
NAND3_X2 U15407 ( .A1(n18634), .A2(n13329), .A3(aes_text_out[9]), .ZN(n17772) );
AND3_X2 U15408 ( .A1(n17773), .A2(n13322), .A3(n17774), .ZN(n16533) );
OR2_X4 U15409 ( .A1(n19198), .A2(n16450), .ZN(n17773) );
NAND3_X2 U15410 ( .A1(n18634), .A2(n13323), .A3(aes_text_out[8]), .ZN(n17774) );
NAND3_X2 U15411 ( .A1(n16447), .A2(n18836), .A3(n16448), .ZN(n16446) );
NAND3_X2 U15412 ( .A1(n16461), .A2(n18837), .A3(n16462), .ZN(n16460) );
NAND3_X2 U15413 ( .A1(n16474), .A2(n18838), .A3(n16475), .ZN(n16473) );
NAND3_X2 U15414 ( .A1(n16487), .A2(n18839), .A3(n16488), .ZN(n16486) );
NAND3_X2 U15415 ( .A1(n16500), .A2(n18840), .A3(n16501), .ZN(n16499) );
NAND3_X2 U15416 ( .A1(n16513), .A2(n18841), .A3(n16514), .ZN(n16512) );
NAND3_X2 U15417 ( .A1(n16526), .A2(n18842), .A3(n16527), .ZN(n16525) );
NAND3_X2 U15418 ( .A1(n16540), .A2(n18843), .A3(n16541), .ZN(n16539) );
NOR2_X2 U15419 ( .A1(n18036), .A2(n16544), .ZN(N3078) );
NOR3_X2 U15420 ( .A1(n16546), .A2(n16547), .A3(n18642), .ZN(n16545) );
NOR2_X2 U15421 ( .A1(n5374), .A2(n18002), .ZN(n16547) );
OR3_X2 U15422 ( .A1(n19205), .A2(dii_data_size[2]), .A3(n19204), .ZN(n17775));
NAND3_X2 U15423 ( .A1(n12235), .A2(n18078), .A3(state[2]), .ZN(n11942) );
INV_X4 U15424 ( .A(dii_data_size[2]), .ZN(n18071) );
NOR2_X2 U15425 ( .A1(n18036), .A2(n16573), .ZN(N3072) );
NOR2_X2 U15426 ( .A1(n18636), .A2(n16575), .ZN(n16574) );
NOR2_X2 U15427 ( .A1(n19197), .A2(n17905), .ZN(n16575) );
NOR2_X2 U15428 ( .A1(n18037), .A2(n16577), .ZN(N3071) );
NOR2_X2 U15429 ( .A1(n18635), .A2(n16579), .ZN(n16578) );
NOR2_X2 U15430 ( .A1(n19198), .A2(n17905), .ZN(n16579) );
NAND3_X2 U15431 ( .A1(n11949), .A2(n18633), .A3(n11950), .ZN(n6285) );
INV_X4 U15432 ( .A(n14414), .ZN(n17886) );
NOR2_X2 U15433 ( .A1(n19205), .A2(dii_data_size[1]), .ZN(n14414) );
NAND3_X2 U15434 ( .A1(n14914), .A2(n18071), .A3(n19201), .ZN(n14736) );
NAND3_X2 U15435 ( .A1(n18846), .A2(n11929), .A3(n17748), .ZN(n11928) );
INV_X4 U15436 ( .A(dii_data_size[3]), .ZN(n18075) );
NOR2_X2 U15437 ( .A1(n11921), .A2(n18894), .ZN(n6295) );
NOR2_X2 U15438 ( .A1(n11922), .A2(n11923), .ZN(n11921) );
NOR2_X2 U15439 ( .A1(n11924), .A2(n18893), .ZN(n11922) );
NOR2_X2 U15440 ( .A1(n18036), .A2(n16569), .ZN(N3073) );
NOR2_X2 U15441 ( .A1(n18637), .A2(n16571), .ZN(n16570) );
NOR2_X2 U15442 ( .A1(n19196), .A2(n17905), .ZN(n16571) );
NAND3_X2 U15443 ( .A1(n14023), .A2(n14024), .A3(n14025), .ZN(n5574) );
NAND3_X2 U15444 ( .A1(n14019), .A2(n14020), .A3(n14021), .ZN(n5575) );
NAND3_X2 U15445 ( .A1(n14015), .A2(n14016), .A3(n14017), .ZN(n5576) );
NAND3_X2 U15446 ( .A1(n14011), .A2(n14012), .A3(n14013), .ZN(n5577) );
NAND3_X2 U15447 ( .A1(n14007), .A2(n14008), .A3(n14009), .ZN(n5578) );
NAND3_X2 U15448 ( .A1(n14003), .A2(n14004), .A3(n14005), .ZN(n5579) );
NAND3_X2 U15449 ( .A1(n13999), .A2(n14000), .A3(n14001), .ZN(n5580) );
NAND3_X2 U15450 ( .A1(n13995), .A2(n13996), .A3(n13997), .ZN(n5581) );
NOR2_X2 U15451 ( .A1(dii_data_size[0]), .A2(dii_data_size[1]), .ZN(n14564));
NOR2_X2 U15452 ( .A1(n18075), .A2(dii_data_size[2]), .ZN(n15309) );
NOR4_X2 U15453 ( .A1(n6850), .A2(n6859), .A3(n16839), .A4(n16838), .ZN(n11929) );
NOR2_X2 U15454 ( .A1(n14188), .A2(n14189), .ZN(n14178) );
NOR2_X2 U15455 ( .A1(n14217), .A2(n14218), .ZN(n14210) );
NOR2_X2 U15456 ( .A1(n14246), .A2(n14247), .ZN(n14239) );
NOR2_X2 U15457 ( .A1(n14275), .A2(n14276), .ZN(n14268) );
NOR2_X2 U15458 ( .A1(n14304), .A2(n14305), .ZN(n14297) );
NOR2_X2 U15459 ( .A1(n14333), .A2(n14334), .ZN(n14326) );
NOR2_X2 U15460 ( .A1(n14362), .A2(n14363), .ZN(n14355) );
NOR2_X2 U15461 ( .A1(n14394), .A2(n14395), .ZN(n14384) );
NOR2_X2 U15462 ( .A1(n15505), .A2(n15506), .ZN(n15495) );
NOR2_X2 U15463 ( .A1(n15529), .A2(n15530), .ZN(n15523) );
NOR2_X2 U15464 ( .A1(n15550), .A2(n15551), .ZN(n15544) );
NOR2_X2 U15465 ( .A1(n15571), .A2(n15572), .ZN(n15565) );
NOR2_X2 U15466 ( .A1(n15592), .A2(n15593), .ZN(n15586) );
NOR2_X2 U15467 ( .A1(n15614), .A2(n15615), .ZN(n15608) );
NOR2_X2 U15468 ( .A1(n15633), .A2(n15634), .ZN(n15627) );
NOR2_X2 U15469 ( .A1(n15653), .A2(n15654), .ZN(n15647) );
NAND3_X2 U15470 ( .A1(n14949), .A2(n17880), .A3(n14950), .ZN(n14597) );
NAND3_X2 U15471 ( .A1(n14971), .A2(n17880), .A3(n14972), .ZN(n14618) );
NAND3_X2 U15472 ( .A1(n14993), .A2(n17881), .A3(n14994), .ZN(n14639) );
NAND3_X2 U15473 ( .A1(n15015), .A2(n17881), .A3(n15016), .ZN(n14660) );
NAND3_X2 U15474 ( .A1(n15037), .A2(n17881), .A3(n15038), .ZN(n14681) );
NAND3_X2 U15475 ( .A1(n15059), .A2(n17880), .A3(n15060), .ZN(n14702) );
NAND3_X2 U15476 ( .A1(n15081), .A2(n17881), .A3(n15082), .ZN(n14723) );
NAND3_X2 U15477 ( .A1(n15105), .A2(n17880), .A3(n15106), .ZN(n14746) );
NAND3_X2 U15478 ( .A1(n15128), .A2(n17880), .A3(n15129), .ZN(n14768) );
NAND3_X2 U15479 ( .A1(n15150), .A2(n17880), .A3(n15151), .ZN(n14791) );
NAND3_X2 U15480 ( .A1(n15172), .A2(n17880), .A3(n15173), .ZN(n14813) );
NAND3_X2 U15481 ( .A1(n15194), .A2(n17880), .A3(n15195), .ZN(n14835) );
NAND3_X2 U15482 ( .A1(n15216), .A2(n17880), .A3(n15217), .ZN(n14857) );
NAND3_X2 U15483 ( .A1(n15238), .A2(n17880), .A3(n15239), .ZN(n14879) );
NAND3_X2 U15484 ( .A1(n15260), .A2(n17880), .A3(n15261), .ZN(n14901) );
NAND3_X2 U15485 ( .A1(n15284), .A2(n17880), .A3(n15285), .ZN(n14924) );
INV_X4 U15486 ( .A(dii_data_size[2]), .ZN(n18072) );
INV_X4 U15487 ( .A(dii_data_size[3]), .ZN(n18076) );
NAND2_X2 U15488 ( .A1(n17882), .A2(dii_data_size[0]), .ZN(n15507) );
INV_X4 U15489 ( .A(dii_data_size[2]), .ZN(n18073) );
INV_X4 U15490 ( .A(rst), .ZN(n18632) );
NAND2_X2 U15491 ( .A1(state[9]), .A2(n11926), .ZN(n18077) );
NAND2_X2 U15492 ( .A1(n18002), .A2(n18077), .ZN(n6294) );
NAND3_X2 U15493 ( .A1(n18630), .A2(n18078), .A3(n18611), .ZN(n18598) );
INV_X4 U15494 ( .A(n18598), .ZN(n18628) );
NAND2_X2 U15495 ( .A1(n18080), .A2(n18079), .ZN(n18597) );
INV_X4 U15496 ( .A(n18597), .ZN(n18627) );
NAND4_X2 U15497 ( .A1(n18600), .A2(n18601), .A3(n18627), .A4(n18626), .ZN(n14157) );
INV_X4 U15498 ( .A(n14157), .ZN(n18625) );
NAND4_X2 U15499 ( .A1(n18628), .A2(state[4]), .A3(n18625), .A4(n18631), .ZN(dii_data_not_ready) );
INV_X4 U15500 ( .A(dii_data_not_ready), .ZN(n18617) );
INV_X4 U15501 ( .A(dii_data_type), .ZN(n18081) );
NAND2_X2 U15502 ( .A1(n11958), .A2(n18085), .ZN(n18083) );
NAND2_X2 U15503 ( .A1(n17776), .A2(n18082), .ZN(n18088) );
NAND2_X2 U15504 ( .A1(n18083), .A2(n18085), .ZN(n18084) );
NAND2_X2 U15505 ( .A1(N2153), .A2(n17800), .ZN(n18086) );
NAND2_X2 U15506 ( .A1(n17776), .A2(n18089), .ZN(n18092) );
NAND2_X2 U15507 ( .A1(N2152), .A2(n17800), .ZN(n18090) );
NAND2_X2 U15508 ( .A1(n17776), .A2(n18093), .ZN(n18096) );
NAND2_X2 U15509 ( .A1(N2151), .A2(n17800), .ZN(n18094) );
NAND2_X2 U15510 ( .A1(n17776), .A2(n18097), .ZN(n18100) );
NAND2_X2 U15511 ( .A1(N2150), .A2(n17800), .ZN(n18098) );
NAND2_X2 U15512 ( .A1(n17776), .A2(n18101), .ZN(n18104) );
NAND2_X2 U15513 ( .A1(N2149), .A2(n17800), .ZN(n18102) );
NAND2_X2 U15514 ( .A1(n17776), .A2(n18105), .ZN(n18108) );
NAND2_X2 U15515 ( .A1(N2148), .A2(n17800), .ZN(n18106) );
NAND2_X2 U15516 ( .A1(n17776), .A2(n18109), .ZN(n18112) );
NAND2_X2 U15517 ( .A1(N2147), .A2(n17800), .ZN(n18110) );
NAND2_X2 U15518 ( .A1(n17776), .A2(n18113), .ZN(n18116) );
NAND2_X2 U15519 ( .A1(N2146), .A2(n17800), .ZN(n18114) );
NAND3_X2 U15520 ( .A1(n18116), .A2(n18115), .A3(n18114), .ZN(n5838) );
NAND2_X2 U15521 ( .A1(n17776), .A2(n18117), .ZN(n18120) );
NAND2_X2 U15522 ( .A1(N2145), .A2(n17800), .ZN(n18118) );
NAND3_X2 U15523 ( .A1(n18120), .A2(n18119), .A3(n18118), .ZN(n5839) );
NAND2_X2 U15524 ( .A1(n17776), .A2(n18121), .ZN(n18124) );
NAND2_X2 U15525 ( .A1(N2144), .A2(n17800), .ZN(n18122) );
NAND3_X2 U15526 ( .A1(n18124), .A2(n18123), .A3(n18122), .ZN(n5840) );
NAND2_X2 U15527 ( .A1(n17776), .A2(n18125), .ZN(n18128) );
NAND2_X2 U15528 ( .A1(N2143), .A2(n17800), .ZN(n18126) );
NAND3_X2 U15529 ( .A1(n18128), .A2(n18127), .A3(n18126), .ZN(n5841) );
NAND2_X2 U15530 ( .A1(n17777), .A2(n18129), .ZN(n18132) );
NAND2_X2 U15531 ( .A1(N2142), .A2(n17801), .ZN(n18130) );
NAND3_X2 U15532 ( .A1(n18132), .A2(n18131), .A3(n18130), .ZN(n5842) );
NAND2_X2 U15533 ( .A1(n17777), .A2(n18133), .ZN(n18136) );
NAND2_X2 U15534 ( .A1(N2141), .A2(n17801), .ZN(n18134) );
NAND3_X2 U15535 ( .A1(n18136), .A2(n18135), .A3(n18134), .ZN(n5843) );
NAND2_X2 U15536 ( .A1(n17777), .A2(n18137), .ZN(n18140) );
NAND2_X2 U15537 ( .A1(N2140), .A2(n17801), .ZN(n18138) );
NAND3_X2 U15538 ( .A1(n18140), .A2(n18139), .A3(n18138), .ZN(n5844) );
NAND2_X2 U15539 ( .A1(n17777), .A2(n18141), .ZN(n18144) );
NAND2_X2 U15540 ( .A1(N2139), .A2(n17801), .ZN(n18142) );
NAND3_X2 U15541 ( .A1(n18144), .A2(n18143), .A3(n18142), .ZN(n5845) );
NAND2_X2 U15542 ( .A1(n17777), .A2(n18145), .ZN(n18148) );
NAND2_X2 U15543 ( .A1(N2138), .A2(n17801), .ZN(n18146) );
NAND2_X2 U15544 ( .A1(n17777), .A2(n18149), .ZN(n18152) );
NAND2_X2 U15545 ( .A1(N2137), .A2(n17801), .ZN(n18150) );
NAND2_X2 U15546 ( .A1(n17777), .A2(n18153), .ZN(n18156) );
NAND2_X2 U15547 ( .A1(N2136), .A2(n17801), .ZN(n18154) );
NAND2_X2 U15548 ( .A1(n17777), .A2(n18157), .ZN(n18160) );
NAND2_X2 U15549 ( .A1(N2135), .A2(n17801), .ZN(n18158) );
NAND2_X2 U15550 ( .A1(n17777), .A2(n18161), .ZN(n18164) );
NAND2_X2 U15551 ( .A1(N2134), .A2(n17801), .ZN(n18162) );
NAND2_X2 U15552 ( .A1(n17777), .A2(n18165), .ZN(n18168) );
NAND2_X2 U15553 ( .A1(N2133), .A2(n17801), .ZN(n18166) );
NAND2_X2 U15554 ( .A1(n17777), .A2(n18169), .ZN(n18172) );
NAND2_X2 U15555 ( .A1(N2132), .A2(n17801), .ZN(n18170) );
NAND2_X2 U15556 ( .A1(n17778), .A2(n18173), .ZN(n18176) );
NAND2_X2 U15557 ( .A1(N2131), .A2(n17802), .ZN(n18174) );
NAND2_X2 U15558 ( .A1(n17778), .A2(n18177), .ZN(n18180) );
NAND2_X2 U15559 ( .A1(N2130), .A2(n17802), .ZN(n18178) );
NAND2_X2 U15560 ( .A1(n17778), .A2(n18181), .ZN(n18184) );
NAND2_X2 U15561 ( .A1(N2129), .A2(n17802), .ZN(n18182) );
NAND2_X2 U15562 ( .A1(n17778), .A2(n18185), .ZN(n18188) );
NAND2_X2 U15563 ( .A1(N2128), .A2(n17802), .ZN(n18186) );
NAND2_X2 U15564 ( .A1(n17778), .A2(n18189), .ZN(n18192) );
NAND2_X2 U15565 ( .A1(N2127), .A2(n17802), .ZN(n18190) );
NAND2_X2 U15566 ( .A1(n17778), .A2(n18193), .ZN(n18196) );
NAND2_X2 U15567 ( .A1(N2126), .A2(n17802), .ZN(n18194) );
NAND2_X2 U15568 ( .A1(n17778), .A2(n18197), .ZN(n18200) );
NAND2_X2 U15569 ( .A1(N2125), .A2(n17802), .ZN(n18198) );
NAND2_X2 U15570 ( .A1(n17778), .A2(n18201), .ZN(n18204) );
NAND2_X2 U15571 ( .A1(N2124), .A2(n17802), .ZN(n18202) );
NAND2_X2 U15572 ( .A1(n17778), .A2(n18205), .ZN(n18208) );
NAND2_X2 U15573 ( .A1(N2123), .A2(n17802), .ZN(n18206) );
NAND2_X2 U15574 ( .A1(n17778), .A2(n18209), .ZN(n18212) );
NAND2_X2 U15575 ( .A1(N2122), .A2(n17802), .ZN(n18210) );
NAND2_X2 U15576 ( .A1(n17778), .A2(n18213), .ZN(n18216) );
NAND2_X2 U15577 ( .A1(N2121), .A2(n17802), .ZN(n18214) );
NAND2_X2 U15578 ( .A1(n17779), .A2(n18217), .ZN(n18220) );
NAND2_X2 U15579 ( .A1(N2120), .A2(n17803), .ZN(n18218) );
NAND2_X2 U15580 ( .A1(n17779), .A2(n18221), .ZN(n18224) );
NAND2_X2 U15581 ( .A1(N2119), .A2(n17803), .ZN(n18222) );
NAND2_X2 U15582 ( .A1(n17779), .A2(n18225), .ZN(n18228) );
NAND2_X2 U15583 ( .A1(N2118), .A2(n17803), .ZN(n18226) );
NAND2_X2 U15584 ( .A1(n17779), .A2(n18229), .ZN(n18232) );
NAND2_X2 U15585 ( .A1(N2117), .A2(n17803), .ZN(n18230) );
NAND2_X2 U15586 ( .A1(n17779), .A2(n18233), .ZN(n18236) );
NAND2_X2 U15587 ( .A1(N2116), .A2(n17803), .ZN(n18234) );
NAND2_X2 U15588 ( .A1(n17779), .A2(n18237), .ZN(n18240) );
NAND2_X2 U15589 ( .A1(N2115), .A2(n17803), .ZN(n18238) );
NAND2_X2 U15590 ( .A1(n17779), .A2(n18241), .ZN(n18244) );
NAND2_X2 U15591 ( .A1(N2114), .A2(n17803), .ZN(n18242) );
NAND2_X2 U15592 ( .A1(n17779), .A2(n18245), .ZN(n18248) );
NAND2_X2 U15593 ( .A1(N2113), .A2(n17803), .ZN(n18246) );
NAND2_X2 U15594 ( .A1(n17779), .A2(n18249), .ZN(n18252) );
NAND2_X2 U15595 ( .A1(N2112), .A2(n17803), .ZN(n18250) );
NAND2_X2 U15596 ( .A1(n17779), .A2(n18253), .ZN(n18256) );
NAND2_X2 U15597 ( .A1(N2111), .A2(n17803), .ZN(n18254) );
NAND2_X2 U15598 ( .A1(n17779), .A2(n18257), .ZN(n18260) );
NAND2_X2 U15599 ( .A1(N2110), .A2(n17803), .ZN(n18258) );
NAND2_X2 U15600 ( .A1(n17780), .A2(n18261), .ZN(n18264) );
NAND2_X2 U15601 ( .A1(N2109), .A2(n17804), .ZN(n18262) );
NAND2_X2 U15602 ( .A1(n17780), .A2(n18265), .ZN(n18268) );
NAND2_X2 U15603 ( .A1(N2108), .A2(n17804), .ZN(n18266) );
NAND2_X2 U15604 ( .A1(n17780), .A2(n18269), .ZN(n18272) );
NAND2_X2 U15605 ( .A1(N2107), .A2(n17804), .ZN(n18270) );
NAND2_X2 U15606 ( .A1(n17780), .A2(n18273), .ZN(n18276) );
NAND2_X2 U15607 ( .A1(N2106), .A2(n17804), .ZN(n18274) );
NAND2_X2 U15608 ( .A1(n17780), .A2(n18277), .ZN(n18280) );
NAND2_X2 U15609 ( .A1(N2105), .A2(n17804), .ZN(n18278) );
NAND2_X2 U15610 ( .A1(n17780), .A2(n18281), .ZN(n18284) );
NAND2_X2 U15611 ( .A1(N2104), .A2(n17804), .ZN(n18282) );
NAND2_X2 U15612 ( .A1(n17780), .A2(n18285), .ZN(n18288) );
NAND2_X2 U15613 ( .A1(N2103), .A2(n17804), .ZN(n18286) );
NAND2_X2 U15614 ( .A1(n17780), .A2(n18289), .ZN(n18292) );
NAND2_X2 U15615 ( .A1(N2102), .A2(n17804), .ZN(n18290) );
NAND2_X2 U15616 ( .A1(n17780), .A2(n18293), .ZN(n18296) );
NAND2_X2 U15617 ( .A1(N2101), .A2(n17804), .ZN(n18294) );
NAND2_X2 U15618 ( .A1(n17780), .A2(n18297), .ZN(n18300) );
NAND2_X2 U15619 ( .A1(N2100), .A2(n17804), .ZN(n18298) );
NAND2_X2 U15620 ( .A1(n17780), .A2(n18301), .ZN(n18304) );
NAND2_X2 U15621 ( .A1(N2099), .A2(n17804), .ZN(n18302) );
NAND2_X2 U15622 ( .A1(n17781), .A2(n18305), .ZN(n18308) );
NAND2_X2 U15623 ( .A1(N2098), .A2(n17805), .ZN(n18306) );
NAND3_X2 U15624 ( .A1(n18308), .A2(n18307), .A3(n18306), .ZN(n5885) );
NAND2_X2 U15625 ( .A1(n17781), .A2(n18309), .ZN(n18312) );
NAND2_X2 U15626 ( .A1(N2097), .A2(n17805), .ZN(n18310) );
NAND3_X2 U15627 ( .A1(n18312), .A2(n18311), .A3(n18310), .ZN(n5886) );
NAND2_X2 U15628 ( .A1(n17781), .A2(n18313), .ZN(n18316) );
NAND2_X2 U15629 ( .A1(N2096), .A2(n17805), .ZN(n18314) );
NAND3_X2 U15630 ( .A1(n18316), .A2(n18315), .A3(n18314), .ZN(n5887) );
NAND2_X2 U15631 ( .A1(n17781), .A2(n18317), .ZN(n18320) );
NAND2_X2 U15632 ( .A1(N2095), .A2(n17805), .ZN(n18318) );
NAND3_X2 U15633 ( .A1(n18320), .A2(n18319), .A3(n18318), .ZN(n5888) );
NAND2_X2 U15634 ( .A1(n17781), .A2(n18321), .ZN(n18324) );
NAND2_X2 U15635 ( .A1(N2094), .A2(n17805), .ZN(n18322) );
NAND3_X2 U15636 ( .A1(n18324), .A2(n18323), .A3(n18322), .ZN(n5889) );
NAND2_X2 U15637 ( .A1(n17781), .A2(n18325), .ZN(n18328) );
NAND2_X2 U15638 ( .A1(N2093), .A2(n17805), .ZN(n18326) );
NAND2_X2 U15639 ( .A1(n17781), .A2(n18329), .ZN(n18332) );
NAND2_X2 U15640 ( .A1(N2092), .A2(n17805), .ZN(n18330) );
NAND2_X2 U15641 ( .A1(n17781), .A2(n18333), .ZN(n18336) );
NAND2_X2 U15642 ( .A1(N2091), .A2(n17805), .ZN(n18334) );
NAND2_X2 U15643 ( .A1(n17781), .A2(n18337), .ZN(n18340) );
NAND2_X2 U15644 ( .A1(N2090), .A2(n17805), .ZN(n18338) );
NAND2_X2 U15645 ( .A1(n17781), .A2(n18341), .ZN(n18344) );
NAND2_X2 U15646 ( .A1(N2089), .A2(n17805), .ZN(n18342) );
NAND2_X2 U15647 ( .A1(n17781), .A2(n18345), .ZN(n18348) );
NAND2_X2 U15648 ( .A1(N2088), .A2(n17805), .ZN(n18346) );
NAND2_X2 U15649 ( .A1(n17782), .A2(n18349), .ZN(n18352) );
NAND2_X2 U15650 ( .A1(N2087), .A2(n17806), .ZN(n18350) );
NAND2_X2 U15651 ( .A1(n17782), .A2(n18353), .ZN(n18356) );
NAND2_X2 U15652 ( .A1(N2086), .A2(n17806), .ZN(n18354) );
NAND2_X2 U15653 ( .A1(n17782), .A2(n18357), .ZN(n18360) );
NAND2_X2 U15654 ( .A1(N2085), .A2(n17806), .ZN(n18358) );
NAND2_X2 U15655 ( .A1(n17782), .A2(n18361), .ZN(n18364) );
NAND2_X2 U15656 ( .A1(N2084), .A2(n17806), .ZN(n18362) );
NAND2_X2 U15657 ( .A1(n17782), .A2(n18365), .ZN(n18368) );
NAND2_X2 U15658 ( .A1(N2083), .A2(n17806), .ZN(n18366) );
NAND2_X2 U15659 ( .A1(n17782), .A2(n18369), .ZN(n18372) );
NAND2_X2 U15660 ( .A1(N2082), .A2(n17806), .ZN(n18370) );
NAND2_X2 U15661 ( .A1(n17782), .A2(n18373), .ZN(n18376) );
NAND2_X2 U15662 ( .A1(N2081), .A2(n17806), .ZN(n18374) );
NAND2_X2 U15663 ( .A1(n17782), .A2(n18377), .ZN(n18380) );
NAND2_X2 U15664 ( .A1(N2080), .A2(n17806), .ZN(n18378) );
NAND2_X2 U15665 ( .A1(n17782), .A2(n18381), .ZN(n18384) );
NAND2_X2 U15666 ( .A1(N2079), .A2(n17806), .ZN(n18382) );
NAND2_X2 U15667 ( .A1(n17782), .A2(n18385), .ZN(n18388) );
NAND2_X2 U15668 ( .A1(N2078), .A2(n17806), .ZN(n18386) );
NAND2_X2 U15669 ( .A1(n17782), .A2(n18389), .ZN(n18392) );
NAND2_X2 U15670 ( .A1(N2077), .A2(n17806), .ZN(n18390) );
NAND2_X2 U15671 ( .A1(n17783), .A2(n18393), .ZN(n18396) );
NAND2_X2 U15672 ( .A1(N2076), .A2(n17807), .ZN(n18394) );
NAND2_X2 U15673 ( .A1(n17783), .A2(n18397), .ZN(n18400) );
NAND2_X2 U15674 ( .A1(N2075), .A2(n17807), .ZN(n18398) );
NAND2_X2 U15675 ( .A1(n17783), .A2(n18401), .ZN(n18404) );
NAND2_X2 U15676 ( .A1(N2074), .A2(n17807), .ZN(n18402) );
NAND2_X2 U15677 ( .A1(n17783), .A2(n18405), .ZN(n18408) );
NAND2_X2 U15678 ( .A1(N2073), .A2(n17807), .ZN(n18406) );
NAND2_X2 U15679 ( .A1(n17783), .A2(n18409), .ZN(n18412) );
NAND2_X2 U15680 ( .A1(N2072), .A2(n17807), .ZN(n18410) );
NAND2_X2 U15681 ( .A1(n17783), .A2(n18413), .ZN(n18416) );
NAND2_X2 U15682 ( .A1(N2071), .A2(n17807), .ZN(n18414) );
NAND2_X2 U15683 ( .A1(n17783), .A2(n18417), .ZN(n18420) );
NAND2_X2 U15684 ( .A1(N2070), .A2(n17807), .ZN(n18418) );
NAND2_X2 U15685 ( .A1(n17783), .A2(n18421), .ZN(n18424) );
NAND2_X2 U15686 ( .A1(N2069), .A2(n17807), .ZN(n18422) );
NAND2_X2 U15687 ( .A1(n17783), .A2(n18425), .ZN(n18428) );
NAND2_X2 U15688 ( .A1(N2068), .A2(n17807), .ZN(n18426) );
NAND2_X2 U15689 ( .A1(n17783), .A2(n18429), .ZN(n18432) );
NAND2_X2 U15690 ( .A1(N2067), .A2(n17807), .ZN(n18430) );
NAND2_X2 U15691 ( .A1(n17783), .A2(n18433), .ZN(n18436) );
NAND2_X2 U15692 ( .A1(N2066), .A2(n17807), .ZN(n18434) );
NAND3_X2 U15693 ( .A1(n18436), .A2(n18435), .A3(n18434), .ZN(n5917) );
NAND2_X2 U15694 ( .A1(n17784), .A2(n18437), .ZN(n18440) );
NAND2_X2 U15695 ( .A1(N2065), .A2(n17808), .ZN(n18438) );
NAND3_X2 U15696 ( .A1(n18440), .A2(n18439), .A3(n18438), .ZN(n5918) );
NAND2_X2 U15697 ( .A1(n17784), .A2(n18441), .ZN(n18444) );
NAND2_X2 U15698 ( .A1(N2064), .A2(n17808), .ZN(n18442) );
NAND3_X2 U15699 ( .A1(n18444), .A2(n18443), .A3(n18442), .ZN(n5919) );
NAND2_X2 U15700 ( .A1(n17784), .A2(n18445), .ZN(n18448) );
NAND2_X2 U15701 ( .A1(N2063), .A2(n17808), .ZN(n18446) );
NAND3_X2 U15702 ( .A1(n18448), .A2(n18447), .A3(n18446), .ZN(n5920) );
NAND2_X2 U15703 ( .A1(n17784), .A2(n18449), .ZN(n18452) );
NAND2_X2 U15704 ( .A1(N2062), .A2(n17808), .ZN(n18450) );
NAND3_X2 U15705 ( .A1(n18452), .A2(n18451), .A3(n18450), .ZN(n5921) );
NAND2_X2 U15706 ( .A1(n17784), .A2(n18453), .ZN(n18456) );
NAND2_X2 U15707 ( .A1(N2061), .A2(n17808), .ZN(n18454) );
NAND3_X2 U15708 ( .A1(n18456), .A2(n18455), .A3(n18454), .ZN(n5922) );
NAND2_X2 U15709 ( .A1(n17784), .A2(n18457), .ZN(n18460) );
NAND2_X2 U15710 ( .A1(N2060), .A2(n17808), .ZN(n18458) );
NAND3_X2 U15711 ( .A1(n18460), .A2(n18459), .A3(n18458), .ZN(n5923) );
NAND2_X2 U15712 ( .A1(n17784), .A2(n18461), .ZN(n18464) );
NAND2_X2 U15713 ( .A1(N2059), .A2(n17808), .ZN(n18462) );
NAND3_X2 U15714 ( .A1(n18464), .A2(n18463), .A3(n18462), .ZN(n5924) );
NAND2_X2 U15715 ( .A1(n17784), .A2(n18465), .ZN(n18468) );
NAND2_X2 U15716 ( .A1(N2058), .A2(n17808), .ZN(n18466) );
NAND3_X2 U15717 ( .A1(n18468), .A2(n18467), .A3(n18466), .ZN(n5925) );
NAND2_X2 U15718 ( .A1(n17784), .A2(n18469), .ZN(n18472) );
NAND2_X2 U15719 ( .A1(N2057), .A2(n17808), .ZN(n18470) );
NAND3_X2 U15720 ( .A1(n18472), .A2(n18471), .A3(n18470), .ZN(n5926) );
NAND2_X2 U15721 ( .A1(n17784), .A2(n18473), .ZN(n18476) );
NAND2_X2 U15722 ( .A1(N2056), .A2(n17808), .ZN(n18474) );
NAND3_X2 U15723 ( .A1(n18476), .A2(n18475), .A3(n18474), .ZN(n5927) );
NAND2_X2 U15724 ( .A1(n17784), .A2(n18477), .ZN(n18480) );
NAND2_X2 U15725 ( .A1(N2055), .A2(n17808), .ZN(n18478) );
NAND3_X2 U15726 ( .A1(n18480), .A2(n18479), .A3(n18478), .ZN(n5928) );
NAND2_X2 U15727 ( .A1(n17785), .A2(n18481), .ZN(n18484) );
NAND2_X2 U15728 ( .A1(N2054), .A2(n17809), .ZN(n18482) );
NAND3_X2 U15729 ( .A1(n18484), .A2(n18483), .A3(n18482), .ZN(n5929) );
NAND2_X2 U15730 ( .A1(n17785), .A2(n18485), .ZN(n18488) );
NAND2_X2 U15731 ( .A1(N2053), .A2(n17809), .ZN(n18486) );
NAND3_X2 U15732 ( .A1(n18488), .A2(n18487), .A3(n18486), .ZN(n5930) );
NAND2_X2 U15733 ( .A1(n17785), .A2(n18489), .ZN(n18492) );
NAND2_X2 U15734 ( .A1(N2052), .A2(n17809), .ZN(n18490) );
NAND3_X2 U15735 ( .A1(n18492), .A2(n18491), .A3(n18490), .ZN(n5931) );
NAND2_X2 U15736 ( .A1(n17785), .A2(n18493), .ZN(n18496) );
NAND2_X2 U15737 ( .A1(N2051), .A2(n17809), .ZN(n18494) );
NAND3_X2 U15738 ( .A1(n18496), .A2(n18495), .A3(n18494), .ZN(n5932) );
NAND2_X2 U15739 ( .A1(n17785), .A2(n18497), .ZN(n18500) );
NAND2_X2 U15740 ( .A1(N2050), .A2(n17809), .ZN(n18498) );
NAND3_X2 U15741 ( .A1(n18500), .A2(n18499), .A3(n18498), .ZN(n5933) );
NAND2_X2 U15742 ( .A1(n17785), .A2(n18501), .ZN(n18504) );
NAND2_X2 U15743 ( .A1(N2049), .A2(n17809), .ZN(n18502) );
NAND3_X2 U15744 ( .A1(n18504), .A2(n18503), .A3(n18502), .ZN(n5934) );
NAND2_X2 U15745 ( .A1(n17785), .A2(n18505), .ZN(n18508) );
NAND2_X2 U15746 ( .A1(N2048), .A2(n17809), .ZN(n18506) );
NAND3_X2 U15747 ( .A1(n18508), .A2(n18507), .A3(n18506), .ZN(n5935) );
NAND2_X2 U15748 ( .A1(n17785), .A2(n18509), .ZN(n18512) );
NAND2_X2 U15749 ( .A1(N2047), .A2(n17809), .ZN(n18510) );
NAND3_X2 U15750 ( .A1(n18512), .A2(n18511), .A3(n18510), .ZN(n5936) );
NAND2_X2 U15751 ( .A1(n17785), .A2(n18513), .ZN(n18516) );
NAND2_X2 U15752 ( .A1(N2046), .A2(n17809), .ZN(n18514) );
NAND3_X2 U15753 ( .A1(n18516), .A2(n18515), .A3(n18514), .ZN(n5937) );
NAND2_X2 U15754 ( .A1(n17785), .A2(n18517), .ZN(n18520) );
NAND2_X2 U15755 ( .A1(N2045), .A2(n17809), .ZN(n18518) );
NAND3_X2 U15756 ( .A1(n18520), .A2(n18519), .A3(n18518), .ZN(n5938) );
NAND2_X2 U15757 ( .A1(n17785), .A2(n18521), .ZN(n18524) );
NAND2_X2 U15758 ( .A1(N2044), .A2(n17809), .ZN(n18522) );
NAND3_X2 U15759 ( .A1(n18524), .A2(n18523), .A3(n18522), .ZN(n5939) );
NAND2_X2 U15760 ( .A1(n17786), .A2(n18525), .ZN(n18528) );
NAND2_X2 U15761 ( .A1(N2043), .A2(n17810), .ZN(n18526) );
NAND3_X2 U15762 ( .A1(n18528), .A2(n18527), .A3(n18526), .ZN(n5940) );
NAND2_X2 U15763 ( .A1(n17786), .A2(n18529), .ZN(n18532) );
NAND2_X2 U15764 ( .A1(N2042), .A2(n17810), .ZN(n18530) );
NAND3_X2 U15765 ( .A1(n18532), .A2(n18531), .A3(n18530), .ZN(n5941) );
NAND2_X2 U15766 ( .A1(n17786), .A2(n18533), .ZN(n18536) );
NAND2_X2 U15767 ( .A1(N2041), .A2(n17810), .ZN(n18534) );
NAND3_X2 U15768 ( .A1(n18536), .A2(n18535), .A3(n18534), .ZN(n5942) );
NAND2_X2 U15769 ( .A1(n17786), .A2(n18537), .ZN(n18540) );
NAND2_X2 U15770 ( .A1(N2040), .A2(n17810), .ZN(n18538) );
NAND3_X2 U15771 ( .A1(n18540), .A2(n18539), .A3(n18538), .ZN(n5943) );
NAND2_X2 U15772 ( .A1(n17786), .A2(n18541), .ZN(n18544) );
NAND2_X2 U15773 ( .A1(N2039), .A2(n17810), .ZN(n18542) );
NAND3_X2 U15774 ( .A1(n18544), .A2(n18543), .A3(n18542), .ZN(n5944) );
NAND2_X2 U15775 ( .A1(n17786), .A2(n18545), .ZN(n18548) );
NAND2_X2 U15776 ( .A1(N2038), .A2(n17810), .ZN(n18546) );
NAND3_X2 U15777 ( .A1(n18548), .A2(n18547), .A3(n18546), .ZN(n5945) );
NAND2_X2 U15778 ( .A1(n17786), .A2(n18549), .ZN(n18552) );
NAND2_X2 U15779 ( .A1(N2037), .A2(n17810), .ZN(n18550) );
NAND3_X2 U15780 ( .A1(n18552), .A2(n18551), .A3(n18550), .ZN(n5946) );
NAND2_X2 U15781 ( .A1(n17786), .A2(n18553), .ZN(n18556) );
NAND2_X2 U15782 ( .A1(N2036), .A2(n17810), .ZN(n18554) );
NAND3_X2 U15783 ( .A1(n18556), .A2(n18555), .A3(n18554), .ZN(n5947) );
NAND2_X2 U15784 ( .A1(n17786), .A2(n18557), .ZN(n18560) );
NAND2_X2 U15785 ( .A1(N2035), .A2(n17810), .ZN(n18558) );
NAND3_X2 U15786 ( .A1(n18560), .A2(n18559), .A3(n18558), .ZN(n5948) );
NAND2_X2 U15787 ( .A1(n17786), .A2(n18561), .ZN(n18564) );
NAND2_X2 U15788 ( .A1(N2034), .A2(n17810), .ZN(n18562) );
NAND3_X2 U15789 ( .A1(n18564), .A2(n18563), .A3(n18562), .ZN(n5949) );
NAND2_X2 U15790 ( .A1(n17786), .A2(n18565), .ZN(n18568) );
NAND2_X2 U15791 ( .A1(N2033), .A2(n17810), .ZN(n18566) );
NAND3_X2 U15792 ( .A1(n18568), .A2(n18567), .A3(n18566), .ZN(n5950) );
NAND2_X2 U15793 ( .A1(n17787), .A2(n18569), .ZN(n18572) );
NAND2_X2 U15794 ( .A1(N2032), .A2(n17811), .ZN(n18570) );
NAND3_X2 U15795 ( .A1(n18572), .A2(n18571), .A3(n18570), .ZN(n5951) );
NAND2_X2 U15796 ( .A1(n17787), .A2(n18573), .ZN(n18576) );
NAND2_X2 U15797 ( .A1(N2031), .A2(n17811), .ZN(n18574) );
NAND3_X2 U15798 ( .A1(n18576), .A2(n18575), .A3(n18574), .ZN(n5952) );
NAND2_X2 U15799 ( .A1(n17787), .A2(n18577), .ZN(n18580) );
NAND2_X2 U15800 ( .A1(N2030), .A2(n17811), .ZN(n18578) );
NAND3_X2 U15801 ( .A1(n18580), .A2(n18579), .A3(n18578), .ZN(n5953) );
NAND2_X2 U15802 ( .A1(n17787), .A2(n18581), .ZN(n18584) );
NAND2_X2 U15803 ( .A1(N2029), .A2(n17811), .ZN(n18582) );
NAND3_X2 U15804 ( .A1(n18584), .A2(n18583), .A3(n18582), .ZN(n5954) );
NAND2_X2 U15805 ( .A1(n17787), .A2(n18585), .ZN(n18588) );
NAND2_X2 U15806 ( .A1(N2028), .A2(n17811), .ZN(n18586) );
NAND3_X2 U15807 ( .A1(n18588), .A2(n18587), .A3(n18586), .ZN(n5955) );
NAND2_X2 U15808 ( .A1(n17787), .A2(n18589), .ZN(n18592) );
NAND2_X2 U15809 ( .A1(N2027), .A2(n17811), .ZN(n18590) );
NAND3_X2 U15810 ( .A1(n18592), .A2(n18591), .A3(n18590), .ZN(n5956) );
NAND2_X2 U15811 ( .A1(n17787), .A2(n18593), .ZN(n18596) );
NAND2_X2 U15812 ( .A1(N2154), .A2(n17811), .ZN(n18594) );
NOR4_X2 U15813 ( .A1(state[4]), .A2(n18598), .A3(n18626), .A4(n18597), .ZN(n18599) );
NAND4_X2 U15814 ( .A1(n18631), .A2(n18601), .A3(n18600), .A4(n18599), .ZN(n11939) );
NAND2_X2 U15815 ( .A1(n11942), .A2(n11939), .ZN(n18602) );
NOR2_X2 U15816 ( .A1(n5444), .A2(n18003), .ZN(aes_text_in[127]) );
NOR2_X2 U15817 ( .A1(n5445), .A2(n18014), .ZN(aes_text_in[126]) );
NOR2_X2 U15818 ( .A1(n5446), .A2(n18014), .ZN(aes_text_in[125]) );
NOR2_X2 U15819 ( .A1(n5447), .A2(n18014), .ZN(aes_text_in[124]) );
NOR2_X2 U15820 ( .A1(n5448), .A2(n18014), .ZN(aes_text_in[123]) );
NOR2_X2 U15821 ( .A1(n5449), .A2(n18014), .ZN(aes_text_in[122]) );
NOR2_X2 U15822 ( .A1(n5450), .A2(n18014), .ZN(aes_text_in[121]) );
NOR2_X2 U15823 ( .A1(n5451), .A2(n18014), .ZN(aes_text_in[120]) );
NOR2_X2 U15824 ( .A1(n5452), .A2(n18013), .ZN(aes_text_in[119]) );
NOR2_X2 U15825 ( .A1(n5453), .A2(n18013), .ZN(aes_text_in[118]) );
NOR2_X2 U15826 ( .A1(n5454), .A2(n18013), .ZN(aes_text_in[117]) );
NOR2_X2 U15827 ( .A1(n5455), .A2(n18013), .ZN(aes_text_in[116]) );
NOR2_X2 U15828 ( .A1(n5456), .A2(n18013), .ZN(aes_text_in[115]) );
NOR2_X2 U15829 ( .A1(n5457), .A2(n18013), .ZN(aes_text_in[114]) );
NOR2_X2 U15830 ( .A1(n5458), .A2(n18013), .ZN(aes_text_in[113]) );
NOR2_X2 U15831 ( .A1(n5459), .A2(n18013), .ZN(aes_text_in[112]) );
NOR2_X2 U15832 ( .A1(n5460), .A2(n18013), .ZN(aes_text_in[111]) );
NOR2_X2 U15833 ( .A1(n5461), .A2(n18013), .ZN(aes_text_in[110]) );
NOR2_X2 U15834 ( .A1(n5462), .A2(n18012), .ZN(aes_text_in[109]) );
NOR2_X2 U15835 ( .A1(n5463), .A2(n18013), .ZN(aes_text_in[108]) );
NOR2_X2 U15836 ( .A1(n5464), .A2(n18012), .ZN(aes_text_in[107]) );
NOR2_X2 U15837 ( .A1(n5465), .A2(n18012), .ZN(aes_text_in[106]) );
NOR2_X2 U15838 ( .A1(n5466), .A2(n18012), .ZN(aes_text_in[105]) );
NOR2_X2 U15839 ( .A1(n5467), .A2(n18012), .ZN(aes_text_in[104]) );
NOR2_X2 U15840 ( .A1(n5468), .A2(n18012), .ZN(aes_text_in[103]) );
NOR2_X2 U15841 ( .A1(n5469), .A2(n18012), .ZN(aes_text_in[102]) );
NOR2_X2 U15842 ( .A1(n5470), .A2(n18012), .ZN(aes_text_in[101]) );
NOR2_X2 U15843 ( .A1(n5471), .A2(n18012), .ZN(aes_text_in[100]) );
NOR2_X2 U15844 ( .A1(n5472), .A2(n18012), .ZN(aes_text_in[99]) );
NOR2_X2 U15845 ( .A1(n5473), .A2(n18012), .ZN(aes_text_in[98]) );
NOR2_X2 U15846 ( .A1(n5474), .A2(n18011), .ZN(aes_text_in[97]) );
NOR2_X2 U15847 ( .A1(n5475), .A2(n18011), .ZN(aes_text_in[96]) );
NOR2_X2 U15848 ( .A1(n5476), .A2(n18011), .ZN(aes_text_in[95]) );
NOR2_X2 U15849 ( .A1(n5477), .A2(n18011), .ZN(aes_text_in[94]) );
NOR2_X2 U15850 ( .A1(n5478), .A2(n18011), .ZN(aes_text_in[93]) );
NOR2_X2 U15851 ( .A1(n5479), .A2(n18011), .ZN(aes_text_in[92]) );
NOR2_X2 U15852 ( .A1(n5480), .A2(n18011), .ZN(aes_text_in[91]) );
NOR2_X2 U15853 ( .A1(n5481), .A2(n18011), .ZN(aes_text_in[90]) );
NOR2_X2 U15854 ( .A1(n5482), .A2(n18011), .ZN(aes_text_in[89]) );
NOR2_X2 U15855 ( .A1(n5483), .A2(n18011), .ZN(aes_text_in[88]) );
NOR2_X2 U15856 ( .A1(n5484), .A2(n18011), .ZN(aes_text_in[87]) );
NOR2_X2 U15857 ( .A1(n5485), .A2(n18010), .ZN(aes_text_in[86]) );
NOR2_X2 U15858 ( .A1(n5486), .A2(n18010), .ZN(aes_text_in[85]) );
NOR2_X2 U15859 ( .A1(n5487), .A2(n18010), .ZN(aes_text_in[84]) );
NOR2_X2 U15860 ( .A1(n5488), .A2(n18010), .ZN(aes_text_in[83]) );
NOR2_X2 U15861 ( .A1(n5489), .A2(n18010), .ZN(aes_text_in[82]) );
NOR2_X2 U15862 ( .A1(n5490), .A2(n18010), .ZN(aes_text_in[81]) );
NOR2_X2 U15863 ( .A1(n5491), .A2(n18010), .ZN(aes_text_in[80]) );
NOR2_X2 U15864 ( .A1(n5492), .A2(n18010), .ZN(aes_text_in[79]) );
NOR2_X2 U15865 ( .A1(n5493), .A2(n18010), .ZN(aes_text_in[78]) );
NOR2_X2 U15866 ( .A1(n5494), .A2(n18010), .ZN(aes_text_in[77]) );
NOR2_X2 U15867 ( .A1(n5495), .A2(n18010), .ZN(aes_text_in[76]) );
NOR2_X2 U15868 ( .A1(n5496), .A2(n18009), .ZN(aes_text_in[75]) );
NOR2_X2 U15869 ( .A1(n5497), .A2(n18009), .ZN(aes_text_in[74]) );
NOR2_X2 U15870 ( .A1(n5498), .A2(n18009), .ZN(aes_text_in[73]) );
NOR2_X2 U15871 ( .A1(n5499), .A2(n18009), .ZN(aes_text_in[72]) );
NOR2_X2 U15872 ( .A1(n5500), .A2(n18009), .ZN(aes_text_in[71]) );
NOR2_X2 U15873 ( .A1(n5501), .A2(n18009), .ZN(aes_text_in[70]) );
NOR2_X2 U15874 ( .A1(n5502), .A2(n18009), .ZN(aes_text_in[69]) );
NOR2_X2 U15875 ( .A1(n5503), .A2(n18009), .ZN(aes_text_in[68]) );
NOR2_X2 U15876 ( .A1(n5504), .A2(n18009), .ZN(aes_text_in[67]) );
NOR2_X2 U15877 ( .A1(n5505), .A2(n18009), .ZN(aes_text_in[66]) );
NOR2_X2 U15878 ( .A1(n5506), .A2(n18009), .ZN(aes_text_in[65]) );
NOR2_X2 U15879 ( .A1(n5507), .A2(n18008), .ZN(aes_text_in[64]) );
NOR2_X2 U15880 ( .A1(n5508), .A2(n18008), .ZN(aes_text_in[63]) );
NOR2_X2 U15881 ( .A1(n5509), .A2(n18008), .ZN(aes_text_in[62]) );
NOR2_X2 U15882 ( .A1(n5510), .A2(n18008), .ZN(aes_text_in[61]) );
NOR2_X2 U15883 ( .A1(n5511), .A2(n18008), .ZN(aes_text_in[60]) );
NOR2_X2 U15884 ( .A1(n5512), .A2(n18008), .ZN(aes_text_in[59]) );
NOR2_X2 U15885 ( .A1(n5513), .A2(n18008), .ZN(aes_text_in[58]) );
NOR2_X2 U15886 ( .A1(n5514), .A2(n18008), .ZN(aes_text_in[57]) );
NOR2_X2 U15887 ( .A1(n5515), .A2(n18008), .ZN(aes_text_in[56]) );
NOR2_X2 U15888 ( .A1(n5516), .A2(n18008), .ZN(aes_text_in[55]) );
NOR2_X2 U15889 ( .A1(n5517), .A2(n18007), .ZN(aes_text_in[54]) );
NOR2_X2 U15890 ( .A1(n5518), .A2(n18007), .ZN(aes_text_in[53]) );
NOR2_X2 U15891 ( .A1(n5519), .A2(n18007), .ZN(aes_text_in[52]) );
NOR2_X2 U15892 ( .A1(n5520), .A2(n18007), .ZN(aes_text_in[51]) );
NOR2_X2 U15893 ( .A1(n5521), .A2(n18007), .ZN(aes_text_in[50]) );
NOR2_X2 U15894 ( .A1(n5522), .A2(n18007), .ZN(aes_text_in[49]) );
NOR2_X2 U15895 ( .A1(n5523), .A2(n18007), .ZN(aes_text_in[48]) );
NOR2_X2 U15896 ( .A1(n5524), .A2(n18007), .ZN(aes_text_in[47]) );
NOR2_X2 U15897 ( .A1(n5525), .A2(n18007), .ZN(aes_text_in[46]) );
NOR2_X2 U15898 ( .A1(n5526), .A2(n18007), .ZN(aes_text_in[45]) );
NOR2_X2 U15899 ( .A1(n5527), .A2(n18007), .ZN(aes_text_in[44]) );
NOR2_X2 U15900 ( .A1(n5528), .A2(n18006), .ZN(aes_text_in[43]) );
NOR2_X2 U15901 ( .A1(n5529), .A2(n18006), .ZN(aes_text_in[42]) );
NOR2_X2 U15902 ( .A1(n5530), .A2(n18006), .ZN(aes_text_in[41]) );
NOR2_X2 U15903 ( .A1(n5531), .A2(n18006), .ZN(aes_text_in[40]) );
NOR2_X2 U15904 ( .A1(n5532), .A2(n18006), .ZN(aes_text_in[39]) );
NOR2_X2 U15905 ( .A1(n5533), .A2(n18006), .ZN(aes_text_in[38]) );
NOR2_X2 U15906 ( .A1(n5534), .A2(n18006), .ZN(aes_text_in[37]) );
NOR2_X2 U15907 ( .A1(n5535), .A2(n18006), .ZN(aes_text_in[36]) );
NOR2_X2 U15908 ( .A1(n5536), .A2(n18006), .ZN(aes_text_in[35]) );
NOR2_X2 U15909 ( .A1(n5537), .A2(n18006), .ZN(aes_text_in[34]) );
NOR2_X2 U15910 ( .A1(n5538), .A2(n18006), .ZN(aes_text_in[33]) );
NOR2_X2 U15911 ( .A1(n5539), .A2(n18005), .ZN(aes_text_in[32]) );
NOR2_X2 U15912 ( .A1(n5540), .A2(n18005), .ZN(aes_text_in[31]) );
NOR2_X2 U15913 ( .A1(n5541), .A2(n18008), .ZN(aes_text_in[30]) );
NOR2_X2 U15914 ( .A1(n5542), .A2(n18005), .ZN(aes_text_in[29]) );
NOR2_X2 U15915 ( .A1(n5543), .A2(n18005), .ZN(aes_text_in[28]) );
NOR2_X2 U15916 ( .A1(n5544), .A2(n18005), .ZN(aes_text_in[27]) );
NOR2_X2 U15917 ( .A1(n5545), .A2(n18005), .ZN(aes_text_in[26]) );
NOR2_X2 U15918 ( .A1(n5546), .A2(n18005), .ZN(aes_text_in[25]) );
NOR2_X2 U15919 ( .A1(n5547), .A2(n18005), .ZN(aes_text_in[24]) );
NOR2_X2 U15920 ( .A1(n5548), .A2(n18005), .ZN(aes_text_in[23]) );
NOR2_X2 U15921 ( .A1(n5549), .A2(n18005), .ZN(aes_text_in[22]) );
NOR2_X2 U15922 ( .A1(n5550), .A2(n18005), .ZN(aes_text_in[21]) );
NOR2_X2 U15923 ( .A1(n5551), .A2(n18004), .ZN(aes_text_in[20]) );
NOR2_X2 U15924 ( .A1(n5552), .A2(n18004), .ZN(aes_text_in[19]) );
NOR2_X2 U15925 ( .A1(n5553), .A2(n18004), .ZN(aes_text_in[18]) );
NOR2_X2 U15926 ( .A1(n5554), .A2(n18004), .ZN(aes_text_in[17]) );
NOR2_X2 U15927 ( .A1(n5555), .A2(n18004), .ZN(aes_text_in[16]) );
NOR2_X2 U15928 ( .A1(n5556), .A2(n18004), .ZN(aes_text_in[15]) );
NOR2_X2 U15929 ( .A1(n5557), .A2(n18004), .ZN(aes_text_in[14]) );
NOR2_X2 U15930 ( .A1(n5558), .A2(n18004), .ZN(aes_text_in[13]) );
NOR2_X2 U15931 ( .A1(n5559), .A2(n18004), .ZN(aes_text_in[12]) );
NOR2_X2 U15932 ( .A1(n5560), .A2(n18004), .ZN(aes_text_in[11]) );
NOR2_X2 U15933 ( .A1(n5561), .A2(n18004), .ZN(aes_text_in[10]) );
NOR2_X2 U15934 ( .A1(n5562), .A2(n18003), .ZN(aes_text_in[9]) );
NOR2_X2 U15935 ( .A1(n5563), .A2(n18003), .ZN(aes_text_in[8]) );
NOR2_X2 U15936 ( .A1(n5564), .A2(n18003), .ZN(aes_text_in[7]) );
NOR2_X2 U15937 ( .A1(n5565), .A2(n18003), .ZN(aes_text_in[6]) );
NOR2_X2 U15938 ( .A1(n5566), .A2(n18003), .ZN(aes_text_in[5]) );
NOR2_X2 U15939 ( .A1(n5567), .A2(n18003), .ZN(aes_text_in[4]) );
NOR2_X2 U15940 ( .A1(n5568), .A2(n18003), .ZN(aes_text_in[3]) );
NOR2_X2 U15941 ( .A1(n5569), .A2(n18003), .ZN(aes_text_in[2]) );
NOR2_X2 U15942 ( .A1(n5570), .A2(n18003), .ZN(aes_text_in[1]) );
NOR2_X2 U15943 ( .A1(n5571), .A2(n18003), .ZN(aes_text_in[0]) );
NAND2_X2 U15944 ( .A1(n11955), .A2(n11929), .ZN(n11961) );
MUX2_X2 U15945 ( .A(enc_byte_cnt[60]), .B(N2409), .S(n17812), .Z(n5381) );
MUX2_X2 U15946 ( .A(enc_byte_cnt[59]), .B(N2408), .S(n17812), .Z(n5382) );
MUX2_X2 U15947 ( .A(enc_byte_cnt[58]), .B(N2407), .S(n17812), .Z(n5383) );
MUX2_X2 U15948 ( .A(enc_byte_cnt[57]), .B(N2406), .S(n17812), .Z(n5384) );
MUX2_X2 U15949 ( .A(enc_byte_cnt[56]), .B(N2405), .S(n17812), .Z(n5385) );
MUX2_X2 U15950 ( .A(enc_byte_cnt[55]), .B(N2404), .S(n17812), .Z(n5386) );
MUX2_X2 U15951 ( .A(enc_byte_cnt[54]), .B(N2403), .S(n17812), .Z(n5387) );
MUX2_X2 U15952 ( .A(enc_byte_cnt[53]), .B(N2402), .S(n17812), .Z(n5388) );
MUX2_X2 U15953 ( .A(enc_byte_cnt[52]), .B(N2401), .S(n17812), .Z(n5389) );
MUX2_X2 U15954 ( .A(enc_byte_cnt[51]), .B(N2400), .S(n17812), .Z(n5390) );
MUX2_X2 U15955 ( .A(enc_byte_cnt[50]), .B(N2399), .S(n17812), .Z(n5391) );
MUX2_X2 U15956 ( .A(enc_byte_cnt[49]), .B(N2398), .S(n17813), .Z(n5392) );
MUX2_X2 U15957 ( .A(enc_byte_cnt[48]), .B(N2397), .S(n17813), .Z(n5393) );
MUX2_X2 U15958 ( .A(enc_byte_cnt[47]), .B(N2396), .S(n17813), .Z(n5394) );
MUX2_X2 U15959 ( .A(enc_byte_cnt[46]), .B(N2395), .S(n17813), .Z(n5395) );
MUX2_X2 U15960 ( .A(enc_byte_cnt[45]), .B(N2394), .S(n17813), .Z(n5396) );
MUX2_X2 U15961 ( .A(enc_byte_cnt[44]), .B(N2393), .S(n17813), .Z(n5397) );
MUX2_X2 U15962 ( .A(enc_byte_cnt[43]), .B(N2392), .S(n17813), .Z(n5398) );
MUX2_X2 U15963 ( .A(enc_byte_cnt[42]), .B(N2391), .S(n17813), .Z(n5399) );
MUX2_X2 U15964 ( .A(enc_byte_cnt[41]), .B(N2390), .S(n17813), .Z(n5400) );
MUX2_X2 U15965 ( .A(enc_byte_cnt[40]), .B(N2389), .S(n17813), .Z(n5401) );
MUX2_X2 U15966 ( .A(enc_byte_cnt[39]), .B(N2388), .S(n17813), .Z(n5402) );
MUX2_X2 U15967 ( .A(enc_byte_cnt[38]), .B(N2387), .S(n17814), .Z(n5403) );
MUX2_X2 U15968 ( .A(enc_byte_cnt[37]), .B(N2386), .S(n17814), .Z(n5404) );
MUX2_X2 U15969 ( .A(enc_byte_cnt[36]), .B(N2385), .S(n17814), .Z(n5405) );
MUX2_X2 U15970 ( .A(enc_byte_cnt[35]), .B(N2384), .S(n17814), .Z(n5406) );
MUX2_X2 U15971 ( .A(enc_byte_cnt[34]), .B(N2383), .S(n17814), .Z(n5407) );
MUX2_X2 U15972 ( .A(enc_byte_cnt[33]), .B(N2382), .S(n17814), .Z(n5408) );
MUX2_X2 U15973 ( .A(enc_byte_cnt[32]), .B(N2381), .S(n17814), .Z(n5409) );
MUX2_X2 U15974 ( .A(enc_byte_cnt[31]), .B(N2380), .S(n17814), .Z(n5410) );
MUX2_X2 U15975 ( .A(enc_byte_cnt[30]), .B(N2379), .S(n17814), .Z(n5411) );
MUX2_X2 U15976 ( .A(enc_byte_cnt[29]), .B(N2378), .S(n17814), .Z(n5412) );
MUX2_X2 U15977 ( .A(enc_byte_cnt[28]), .B(N2377), .S(n17814), .Z(n5413) );
MUX2_X2 U15978 ( .A(enc_byte_cnt[27]), .B(N2376), .S(n17815), .Z(n5414) );
MUX2_X2 U15979 ( .A(enc_byte_cnt[26]), .B(N2375), .S(n17815), .Z(n5415) );
MUX2_X2 U15980 ( .A(enc_byte_cnt[25]), .B(N2374), .S(n17815), .Z(n5416) );
MUX2_X2 U15981 ( .A(enc_byte_cnt[24]), .B(N2373), .S(n17815), .Z(n5417) );
MUX2_X2 U15982 ( .A(enc_byte_cnt[23]), .B(N2372), .S(n17815), .Z(n5418) );
MUX2_X2 U15983 ( .A(enc_byte_cnt[22]), .B(N2371), .S(n17815), .Z(n5419) );
MUX2_X2 U15984 ( .A(enc_byte_cnt[21]), .B(N2370), .S(n17815), .Z(n5420) );
MUX2_X2 U15985 ( .A(enc_byte_cnt[20]), .B(N2369), .S(n17815), .Z(n5421) );
MUX2_X2 U15986 ( .A(enc_byte_cnt[19]), .B(N2368), .S(n17815), .Z(n5422) );
MUX2_X2 U15987 ( .A(enc_byte_cnt[18]), .B(N2367), .S(n17815), .Z(n5423) );
MUX2_X2 U15988 ( .A(enc_byte_cnt[17]), .B(N2366), .S(n17815), .Z(n5424) );
MUX2_X2 U15989 ( .A(enc_byte_cnt[16]), .B(N2365), .S(n17816), .Z(n5425) );
MUX2_X2 U15990 ( .A(enc_byte_cnt[15]), .B(N2364), .S(n17816), .Z(n5426) );
MUX2_X2 U15991 ( .A(enc_byte_cnt[14]), .B(N2363), .S(n17816), .Z(n5427) );
MUX2_X2 U15992 ( .A(enc_byte_cnt[13]), .B(N2362), .S(n17816), .Z(n5428) );
MUX2_X2 U15993 ( .A(enc_byte_cnt[12]), .B(N2361), .S(n17816), .Z(n5429) );
MUX2_X2 U15994 ( .A(enc_byte_cnt[11]), .B(N2360), .S(n17816), .Z(n5430) );
MUX2_X2 U15995 ( .A(enc_byte_cnt[10]), .B(N2359), .S(n17816), .Z(n5431) );
MUX2_X2 U15996 ( .A(enc_byte_cnt[9]), .B(N2358), .S(n17816), .Z(n5432) );
MUX2_X2 U15997 ( .A(enc_byte_cnt[8]), .B(N2357), .S(n17816), .Z(n5433) );
MUX2_X2 U15998 ( .A(enc_byte_cnt[7]), .B(N2356), .S(n17816), .Z(n5434) );
MUX2_X2 U15999 ( .A(enc_byte_cnt[6]), .B(N2355), .S(n17816), .Z(n5435) );
MUX2_X2 U16000 ( .A(enc_byte_cnt[5]), .B(N2354), .S(n17817), .Z(n5436) );
MUX2_X2 U16001 ( .A(enc_byte_cnt[4]), .B(N2353), .S(n17817), .Z(n5437) );
MUX2_X2 U16002 ( .A(enc_byte_cnt[3]), .B(N2352), .S(n17817), .Z(n5438) );
MUX2_X2 U16003 ( .A(enc_byte_cnt[2]), .B(N2351), .S(n17817), .Z(n5439) );
NOR2_X2 U16004 ( .A1(n5378), .A2(n18002), .ZN(n18603) );
NOR3_X2 U16005 ( .A1(n16566), .A2(n18638), .A3(n18603), .ZN(n16565) );
NOR2_X2 U16006 ( .A1(n5377), .A2(n18002), .ZN(n18604) );
NOR3_X2 U16007 ( .A1(n16561), .A2(n18639), .A3(n18604), .ZN(n16560) );
NOR2_X2 U16008 ( .A1(n5376), .A2(n18002), .ZN(n18605) );
NOR3_X2 U16009 ( .A1(n16556), .A2(n18640), .A3(n18605), .ZN(n16555) );
NOR2_X2 U16010 ( .A1(n5375), .A2(n18002), .ZN(n18606) );
NOR3_X2 U16011 ( .A1(n16551), .A2(n18641), .A3(n18606), .ZN(n16550) );
NOR2_X2 U16012 ( .A1(n5328), .A2(n18002), .ZN(n15852) );
NOR2_X2 U16013 ( .A1(n5327), .A2(n18002), .ZN(n15834) );
NOR2_X2 U16014 ( .A1(n5326), .A2(n18002), .ZN(n15816) );
NAND2_X2 U16015 ( .A1(n17996), .A2(enc_byte_cnt[53]), .ZN(n15807) );
NAND2_X2 U16016 ( .A1(n17999), .A2(enc_byte_cnt[54]), .ZN(n15786) );
NAND2_X2 U16017 ( .A1(n17283), .A2(enc_byte_cnt[55]), .ZN(n15767) );
NAND2_X2 U16018 ( .A1(n17999), .A2(enc_byte_cnt[56]), .ZN(n15748) );
NAND2_X2 U16019 ( .A1(n17999), .A2(enc_byte_cnt[57]), .ZN(n15729) );
NAND2_X2 U16020 ( .A1(n17999), .A2(enc_byte_cnt[58]), .ZN(n15710) );
NAND2_X2 U16021 ( .A1(n17999), .A2(enc_byte_cnt[59]), .ZN(n15691) );
NAND2_X2 U16022 ( .A1(n17999), .A2(enc_byte_cnt[60]), .ZN(n15672) );
MUX2_X2 U16023 ( .A(aad_byte_cnt[60]), .B(N2539), .S(n17840), .Z(n5960) );
MUX2_X2 U16024 ( .A(aad_byte_cnt[59]), .B(N2538), .S(n17840), .Z(n5961) );
MUX2_X2 U16025 ( .A(aad_byte_cnt[58]), .B(N2537), .S(n17840), .Z(n5962) );
MUX2_X2 U16026 ( .A(aad_byte_cnt[57]), .B(N2536), .S(n17840), .Z(n5963) );
MUX2_X2 U16027 ( .A(aad_byte_cnt[56]), .B(N2535), .S(n17840), .Z(n5964) );
MUX2_X2 U16028 ( .A(aad_byte_cnt[55]), .B(N2534), .S(n17840), .Z(n5965) );
MUX2_X2 U16029 ( .A(aad_byte_cnt[54]), .B(N2533), .S(n17840), .Z(n5966) );
MUX2_X2 U16030 ( .A(aad_byte_cnt[53]), .B(N2532), .S(n17840), .Z(n5967) );
MUX2_X2 U16031 ( .A(aad_byte_cnt[52]), .B(N2531), .S(n17840), .Z(n5968) );
MUX2_X2 U16032 ( .A(aad_byte_cnt[51]), .B(N2530), .S(n17840), .Z(n5969) );
MUX2_X2 U16033 ( .A(aad_byte_cnt[50]), .B(N2529), .S(n17840), .Z(n5970) );
MUX2_X2 U16034 ( .A(aad_byte_cnt[49]), .B(N2528), .S(n17840), .Z(n5971) );
MUX2_X2 U16035 ( .A(aad_byte_cnt[48]), .B(N2527), .S(n17840), .Z(n5972) );
MUX2_X2 U16036 ( .A(aad_byte_cnt[47]), .B(N2526), .S(n17840), .Z(n5973) );
MUX2_X2 U16037 ( .A(aad_byte_cnt[46]), .B(N2525), .S(n17839), .Z(n5974) );
MUX2_X2 U16038 ( .A(aad_byte_cnt[45]), .B(N2524), .S(n17839), .Z(n5975) );
MUX2_X2 U16039 ( .A(aad_byte_cnt[44]), .B(N2523), .S(n17839), .Z(n5976) );
MUX2_X2 U16040 ( .A(aad_byte_cnt[43]), .B(N2522), .S(n17839), .Z(n5977) );
MUX2_X2 U16041 ( .A(aad_byte_cnt[42]), .B(N2521), .S(n17839), .Z(n5978) );
MUX2_X2 U16042 ( .A(aad_byte_cnt[41]), .B(N2520), .S(n17839), .Z(n5979) );
MUX2_X2 U16043 ( .A(aad_byte_cnt[40]), .B(N2519), .S(n17839), .Z(n5980) );
MUX2_X2 U16044 ( .A(aad_byte_cnt[39]), .B(N2518), .S(n17839), .Z(n5981) );
MUX2_X2 U16045 ( .A(aad_byte_cnt[38]), .B(N2517), .S(n17839), .Z(n5982) );
MUX2_X2 U16046 ( .A(aad_byte_cnt[37]), .B(N2516), .S(n17839), .Z(n5983) );
MUX2_X2 U16047 ( .A(aad_byte_cnt[36]), .B(N2515), .S(n17839), .Z(n5984) );
MUX2_X2 U16048 ( .A(aad_byte_cnt[35]), .B(N2514), .S(n17839), .Z(n5985) );
MUX2_X2 U16049 ( .A(aad_byte_cnt[34]), .B(N2513), .S(n17839), .Z(n5986) );
MUX2_X2 U16050 ( .A(aad_byte_cnt[33]), .B(N2512), .S(n17839), .Z(n5987) );
MUX2_X2 U16051 ( .A(aad_byte_cnt[32]), .B(N2511), .S(n17839), .Z(n5988) );
MUX2_X2 U16052 ( .A(aad_byte_cnt[31]), .B(N2510), .S(n17839), .Z(n5989) );
MUX2_X2 U16053 ( .A(aad_byte_cnt[30]), .B(N2509), .S(n17839), .Z(n5990) );
MUX2_X2 U16054 ( .A(aad_byte_cnt[29]), .B(N2508), .S(n17838), .Z(n5991) );
MUX2_X2 U16055 ( .A(aad_byte_cnt[28]), .B(N2507), .S(n17838), .Z(n5992) );
MUX2_X2 U16056 ( .A(aad_byte_cnt[27]), .B(N2506), .S(n17838), .Z(n5993) );
MUX2_X2 U16057 ( .A(aad_byte_cnt[26]), .B(N2505), .S(n17838), .Z(n5994) );
MUX2_X2 U16058 ( .A(aad_byte_cnt[25]), .B(N2504), .S(n17838), .Z(n5995) );
MUX2_X2 U16059 ( .A(aad_byte_cnt[24]), .B(N2503), .S(n17838), .Z(n5996) );
MUX2_X2 U16060 ( .A(aad_byte_cnt[23]), .B(N2502), .S(n17838), .Z(n5997) );
MUX2_X2 U16061 ( .A(aad_byte_cnt[22]), .B(N2501), .S(n17838), .Z(n5998) );
MUX2_X2 U16062 ( .A(aad_byte_cnt[21]), .B(N2500), .S(n17838), .Z(n5999) );
MUX2_X2 U16063 ( .A(aad_byte_cnt[20]), .B(N2499), .S(n17838), .Z(n6000) );
MUX2_X2 U16064 ( .A(aad_byte_cnt[19]), .B(N2498), .S(n17838), .Z(n6001) );
MUX2_X2 U16065 ( .A(aad_byte_cnt[18]), .B(N2497), .S(n17838), .Z(n6002) );
MUX2_X2 U16066 ( .A(aad_byte_cnt[17]), .B(N2496), .S(n17838), .Z(n6003) );
MUX2_X2 U16067 ( .A(aad_byte_cnt[16]), .B(N2495), .S(n17838), .Z(n6004) );
MUX2_X2 U16068 ( .A(aad_byte_cnt[15]), .B(N2494), .S(n17838), .Z(n6005) );
MUX2_X2 U16069 ( .A(aad_byte_cnt[14]), .B(N2493), .S(n17838), .Z(n6006) );
MUX2_X2 U16070 ( .A(aad_byte_cnt[13]), .B(N2492), .S(n17838), .Z(n6007) );
MUX2_X2 U16071 ( .A(aad_byte_cnt[12]), .B(N2491), .S(n17837), .Z(n6008) );
MUX2_X2 U16072 ( .A(aad_byte_cnt[11]), .B(N2490), .S(n17837), .Z(n6009) );
MUX2_X2 U16073 ( .A(aad_byte_cnt[10]), .B(N2489), .S(n17837), .Z(n6010) );
MUX2_X2 U16074 ( .A(aad_byte_cnt[9]), .B(N2488), .S(n17837), .Z(n6011) );
MUX2_X2 U16075 ( .A(aad_byte_cnt[8]), .B(N2487), .S(n17837), .Z(n6012) );
MUX2_X2 U16076 ( .A(aad_byte_cnt[7]), .B(N2486), .S(n17837), .Z(n6013) );
MUX2_X2 U16077 ( .A(aad_byte_cnt[6]), .B(N2485), .S(n17837), .Z(n6014) );
MUX2_X2 U16078 ( .A(aad_byte_cnt[5]), .B(N2484), .S(n17837), .Z(n6015) );
MUX2_X2 U16079 ( .A(aad_byte_cnt[4]), .B(N2483), .S(n17837), .Z(n6016) );
MUX2_X2 U16080 ( .A(aad_byte_cnt[3]), .B(N2482), .S(n17837), .Z(n6017) );
MUX2_X2 U16081 ( .A(aad_byte_cnt[2]), .B(N2481), .S(n17837), .Z(n6018) );
MUX2_X2 U16082 ( .A(aad_byte_cnt[0]), .B(N2479), .S(n17837), .Z(n6020) );
NAND2_X2 U16083 ( .A1(n17999), .A2(aad_byte_cnt[0]), .ZN(n18607) );
NAND2_X2 U16084 ( .A1(n15595), .A2(n18607), .ZN(n15580) );
NAND2_X2 U16085 ( .A1(n17999), .A2(aad_byte_cnt[1]), .ZN(n18608) );
NAND2_X2 U16086 ( .A1(n15574), .A2(n18608), .ZN(n15559) );
NAND2_X2 U16087 ( .A1(n17999), .A2(aad_byte_cnt[2]), .ZN(n18609) );
NAND2_X2 U16088 ( .A1(n15553), .A2(n18609), .ZN(n15538) );
NAND2_X2 U16089 ( .A1(n17999), .A2(aad_byte_cnt[3]), .ZN(n18610) );
NAND2_X2 U16090 ( .A1(n15532), .A2(n18610), .ZN(n15517) );
NAND2_X2 U16091 ( .A1(aad_byte_cnt[50]), .A2(n17283), .ZN(n14455) );
NAND2_X2 U16092 ( .A1(aad_byte_cnt[51]), .A2(n17283), .ZN(n14433) );
NAND2_X2 U16093 ( .A1(aad_byte_cnt[52]), .A2(n17283), .ZN(n14409) );
NAND2_X2 U16094 ( .A1(aad_byte_cnt[53]), .A2(n17283), .ZN(n14370) );
NAND2_X2 U16095 ( .A1(aad_byte_cnt[54]), .A2(n17283), .ZN(n14341) );
NAND2_X2 U16096 ( .A1(aad_byte_cnt[55]), .A2(n17283), .ZN(n14312) );
NAND2_X2 U16097 ( .A1(aad_byte_cnt[56]), .A2(n17283), .ZN(n14283) );
NAND2_X2 U16098 ( .A1(aad_byte_cnt[57]), .A2(n17283), .ZN(n14254) );
NAND2_X2 U16099 ( .A1(aad_byte_cnt[58]), .A2(n17283), .ZN(n14225) );
NAND2_X2 U16100 ( .A1(aad_byte_cnt[59]), .A2(n17283), .ZN(n14196) );
NAND2_X2 U16101 ( .A1(aad_byte_cnt[60]), .A2(n17283), .ZN(n14162) );
NOR3_X2 U16102 ( .A1(n14157), .A2(state[1]), .A3(n18611), .ZN(n14155) );
NAND2_X2 U16103 ( .A1(n18892), .A2(n18044), .ZN(n11924) );
INV_X4 U16104 ( .A(n11924), .ZN(n18623) );
NAND2_X2 U16105 ( .A1(n6850), .A2(n18623), .ZN(n11937) );
INV_X4 U16106 ( .A(n11937), .ZN(n18612) );
NAND2_X2 U16107 ( .A1(n18612), .A2(n18622), .ZN(n18614) );
NAND2_X2 U16108 ( .A1(n17280), .A2(n18624), .ZN(n18613) );
NAND2_X2 U16109 ( .A1(n18614), .A2(n18613), .ZN(n6291) );
NAND3_X2 U16110 ( .A1(n18630), .A2(aes_done), .A3(n17290), .ZN(n18633) );
NAND2_X2 U16111 ( .A1(n17290), .A2(n18630), .ZN(n18615) );
NAND2_X2 U16112 ( .A1(n11976), .A2(n18615), .ZN(n18621) );
INV_X4 U16113 ( .A(n18621), .ZN(n18844) );
NOR4_X2 U16114 ( .A1(n11967), .A2(n11955), .A3(n11971), .A4(n17996), .ZN(n11970) );
NAND2_X2 U16115 ( .A1(n11968), .A2(n11967), .ZN(n11965) );
NAND2_X2 U16116 ( .A1(n18846), .A2(n18892), .ZN(n11966) );
INV_X4 U16117 ( .A(dii_data_vld), .ZN(n18616) );
NAND2_X2 U16118 ( .A1(n18617), .A2(n18616), .ZN(n18619) );
NAND2_X2 U16119 ( .A1(n19206), .A2(n11971), .ZN(n18618) );
NAND2_X2 U16120 ( .A1(n11960), .A2(state[2]), .ZN(n11959) );
NAND2_X2 U16121 ( .A1(n18747), .A2(n17375), .ZN(n18620) );
NAND2_X2 U16122 ( .A1(state[4]), .A2(n18620), .ZN(n11950) );
NAND2_X2 U16123 ( .A1(n11948), .A2(state[5]), .ZN(n11947) );
NAND2_X2 U16124 ( .A1(n18746), .A2(n18621), .ZN(n11944) );
NAND2_X2 U16125 ( .A1(n11926), .A2(state[3]), .ZN(n11943) );
NAND2_X2 U16126 ( .A1(state[7]), .A2(n11926), .ZN(n11940) );
NAND3_X2 U16127 ( .A1(n16838), .A2(n17291), .A3(n18624), .ZN(n11936) );
NAND2_X2 U16128 ( .A1(n11926), .A2(state[1]), .ZN(n11931) );
NAND2_X2 U16129 ( .A1(state[8]), .A2(n11926), .ZN(n11927) );
INV_X4 U16130 ( .A(n16839), .ZN(n18894) );
MUX2_X2 U16131 ( .A(aad_byte_cnt[62]), .B(N2541), .S(n17837), .Z(n5958) );
MUX2_X2 U16132 ( .A(aad_byte_cnt[61]), .B(N2540), .S(n17837), .Z(n5959) );
MUX2_X2 U16133 ( .A(aad_byte_cnt[63]), .B(N2542), .S(n17837), .Z(n6021) );
MUX2_X2 U16134 ( .A(enc_byte_cnt[62]), .B(N2411), .S(n17817), .Z(n5379) );
MUX2_X2 U16135 ( .A(enc_byte_cnt[61]), .B(N2410), .S(n17817), .Z(n5380) );
MUX2_X2 U16136 ( .A(enc_byte_cnt[63]), .B(N2412), .S(n17817), .Z(n5442) );
INV_X4 U16137 ( .A(n13280), .ZN(n18635) );
INV_X4 U16138 ( .A(n13287), .ZN(n18636) );
INV_X4 U16139 ( .A(n13292), .ZN(n18637) );
INV_X4 U16140 ( .A(n13297), .ZN(n18638) );
INV_X4 U16141 ( .A(n13302), .ZN(n18639) );
INV_X4 U16142 ( .A(n13307), .ZN(n18640) );
INV_X4 U16143 ( .A(n13312), .ZN(n18641) );
INV_X4 U16144 ( .A(n13317), .ZN(n18642) );
INV_X4 U16145 ( .A(n13370), .ZN(n18643) );
INV_X4 U16146 ( .A(n13376), .ZN(n18644) );
INV_X4 U16147 ( .A(n13382), .ZN(n18645) );
INV_X4 U16148 ( .A(n13388), .ZN(n18646) );
INV_X4 U16149 ( .A(n13394), .ZN(n18647) );
INV_X4 U16150 ( .A(n13400), .ZN(n18648) );
INV_X4 U16151 ( .A(n13406), .ZN(n18649) );
INV_X4 U16152 ( .A(n13412), .ZN(n18650) );
INV_X4 U16153 ( .A(n13418), .ZN(n18651) );
INV_X4 U16154 ( .A(n13424), .ZN(n18652) );
INV_X4 U16155 ( .A(n13430), .ZN(n18653) );
INV_X4 U16156 ( .A(n13436), .ZN(n18654) );
INV_X4 U16157 ( .A(n13442), .ZN(n18655) );
INV_X4 U16158 ( .A(n13448), .ZN(n18656) );
INV_X4 U16159 ( .A(n13454), .ZN(n18657) );
INV_X4 U16160 ( .A(n13460), .ZN(n18658) );
INV_X4 U16161 ( .A(n13466), .ZN(n18659) );
INV_X4 U16162 ( .A(n13472), .ZN(n18660) );
INV_X4 U16163 ( .A(n13478), .ZN(n18661) );
INV_X4 U16164 ( .A(n13484), .ZN(n18662) );
INV_X4 U16165 ( .A(n13490), .ZN(n18663) );
INV_X4 U16166 ( .A(n13496), .ZN(n18664) );
INV_X4 U16167 ( .A(n13502), .ZN(n18665) );
INV_X4 U16168 ( .A(n13508), .ZN(n18666) );
INV_X4 U16169 ( .A(n13514), .ZN(n18667) );
INV_X4 U16170 ( .A(n13520), .ZN(n18668) );
INV_X4 U16171 ( .A(n13526), .ZN(n18669) );
INV_X4 U16172 ( .A(n13532), .ZN(n18670) );
INV_X4 U16173 ( .A(n13538), .ZN(n18671) );
INV_X4 U16174 ( .A(n13544), .ZN(n18672) );
INV_X4 U16175 ( .A(n13550), .ZN(n18673) );
INV_X4 U16176 ( .A(n13556), .ZN(n18674) );
INV_X4 U16177 ( .A(n13562), .ZN(n18675) );
INV_X4 U16178 ( .A(n13568), .ZN(n18676) );
INV_X4 U16179 ( .A(n13574), .ZN(n18677) );
INV_X4 U16180 ( .A(n13580), .ZN(n18678) );
INV_X4 U16181 ( .A(n13586), .ZN(n18679) );
INV_X4 U16182 ( .A(n13592), .ZN(n18680) );
INV_X4 U16183 ( .A(n13598), .ZN(n18681) );
INV_X4 U16184 ( .A(n13604), .ZN(n18682) );
INV_X4 U16185 ( .A(n13610), .ZN(n18683) );
INV_X4 U16186 ( .A(n13616), .ZN(n18684) );
INV_X4 U16187 ( .A(n13622), .ZN(n18685) );
INV_X4 U16188 ( .A(n13628), .ZN(n18686) );
INV_X4 U16189 ( .A(n13634), .ZN(n18687) );
INV_X4 U16190 ( .A(n13640), .ZN(n18688) );
INV_X4 U16191 ( .A(n13646), .ZN(n18689) );
INV_X4 U16192 ( .A(n13652), .ZN(n18690) );
INV_X4 U16193 ( .A(n13680), .ZN(n18691) );
INV_X4 U16194 ( .A(n13686), .ZN(n18692) );
INV_X4 U16195 ( .A(n13692), .ZN(n18693) );
INV_X4 U16196 ( .A(n13698), .ZN(n18694) );
INV_X4 U16197 ( .A(n13704), .ZN(n18695) );
INV_X4 U16198 ( .A(n13710), .ZN(n18696) );
INV_X4 U16199 ( .A(n13716), .ZN(n18697) );
INV_X4 U16200 ( .A(n13722), .ZN(n18698) );
INV_X4 U16201 ( .A(n13728), .ZN(n18699) );
INV_X4 U16202 ( .A(n13734), .ZN(n18700) );
INV_X4 U16203 ( .A(n13740), .ZN(n18701) );
INV_X4 U16204 ( .A(n13746), .ZN(n18702) );
INV_X4 U16205 ( .A(n13752), .ZN(n18703) );
INV_X4 U16206 ( .A(n13758), .ZN(n18704) );
INV_X4 U16207 ( .A(n13764), .ZN(n18705) );
INV_X4 U16208 ( .A(n13770), .ZN(n18706) );
INV_X4 U16209 ( .A(n13776), .ZN(n18707) );
INV_X4 U16210 ( .A(n13782), .ZN(n18708) );
INV_X4 U16211 ( .A(n13788), .ZN(n18709) );
INV_X4 U16212 ( .A(n13794), .ZN(n18710) );
INV_X4 U16213 ( .A(n13800), .ZN(n18711) );
INV_X4 U16214 ( .A(n13806), .ZN(n18712) );
INV_X4 U16215 ( .A(n13812), .ZN(n18713) );
INV_X4 U16216 ( .A(n13818), .ZN(n18714) );
INV_X4 U16217 ( .A(n13824), .ZN(n18715) );
INV_X4 U16218 ( .A(n13830), .ZN(n18716) );
INV_X4 U16219 ( .A(n13836), .ZN(n18717) );
INV_X4 U16220 ( .A(n13842), .ZN(n18718) );
INV_X4 U16221 ( .A(n13848), .ZN(n18719) );
INV_X4 U16222 ( .A(n13854), .ZN(n18720) );
INV_X4 U16223 ( .A(n13860), .ZN(n18721) );
INV_X4 U16224 ( .A(n13866), .ZN(n18722) );
INV_X4 U16225 ( .A(n13872), .ZN(n18723) );
INV_X4 U16226 ( .A(n13878), .ZN(n18724) );
INV_X4 U16227 ( .A(n13884), .ZN(n18725) );
INV_X4 U16228 ( .A(n13890), .ZN(n18726) );
INV_X4 U16229 ( .A(n13896), .ZN(n18727) );
INV_X4 U16230 ( .A(n13902), .ZN(n18728) );
INV_X4 U16231 ( .A(n13908), .ZN(n18729) );
INV_X4 U16232 ( .A(n13914), .ZN(n18730) );
INV_X4 U16233 ( .A(n13920), .ZN(n18731) );
INV_X4 U16234 ( .A(n13926), .ZN(n18732) );
INV_X4 U16235 ( .A(n13932), .ZN(n18733) );
INV_X4 U16236 ( .A(n13938), .ZN(n18734) );
INV_X4 U16237 ( .A(n13944), .ZN(n18735) );
INV_X4 U16238 ( .A(n13950), .ZN(n18736) );
INV_X4 U16239 ( .A(n13956), .ZN(n18737) );
INV_X4 U16240 ( .A(n13962), .ZN(n18738) );
INV_X4 U16241 ( .A(n13968), .ZN(n18739) );
INV_X4 U16242 ( .A(n13974), .ZN(n18740) );
INV_X4 U16243 ( .A(n13980), .ZN(n18741) );
INV_X4 U16244 ( .A(n13986), .ZN(n18742) );
INV_X4 U16245 ( .A(n13992), .ZN(n18743) );
INV_X4 U16246 ( .A(n17281), .ZN(n18744) );
INV_X4 U16247 ( .A(n17280), .ZN(n18745) );
INV_X4 U16248 ( .A(aes_done), .ZN(n18746) );
INV_X4 U16249 ( .A(n11948), .ZN(n18747) );
INV_X4 U16250 ( .A(aes_text_out[127]), .ZN(n18748) );
INV_X4 U16251 ( .A(aes_text_out[126]), .ZN(n18749) );
INV_X4 U16252 ( .A(aes_text_out[125]), .ZN(n18750) );
INV_X4 U16253 ( .A(aes_text_out[124]), .ZN(n18751) );
INV_X4 U16254 ( .A(aes_text_out[123]), .ZN(n18752) );
INV_X4 U16255 ( .A(aes_text_out[122]), .ZN(n18753) );
INV_X4 U16256 ( .A(aes_text_out[121]), .ZN(n18754) );
INV_X4 U16257 ( .A(aes_text_out[120]), .ZN(n18755) );
INV_X4 U16258 ( .A(n13994), .ZN(n18756) );
INV_X4 U16259 ( .A(n13988), .ZN(n18757) );
INV_X4 U16260 ( .A(n13982), .ZN(n18758) );
INV_X4 U16261 ( .A(n13976), .ZN(n18759) );
INV_X4 U16262 ( .A(n13970), .ZN(n18760) );
INV_X4 U16263 ( .A(n13964), .ZN(n18761) );
INV_X4 U16264 ( .A(n13958), .ZN(n18762) );
INV_X4 U16265 ( .A(n13952), .ZN(n18763) );
INV_X4 U16266 ( .A(n13946), .ZN(n18764) );
INV_X4 U16267 ( .A(n13940), .ZN(n18765) );
INV_X4 U16268 ( .A(n13934), .ZN(n18766) );
INV_X4 U16269 ( .A(n13928), .ZN(n18767) );
INV_X4 U16270 ( .A(n13922), .ZN(n18768) );
INV_X4 U16271 ( .A(n13916), .ZN(n18769) );
INV_X4 U16272 ( .A(n13910), .ZN(n18770) );
INV_X4 U16273 ( .A(n13904), .ZN(n18771) );
INV_X4 U16274 ( .A(n13898), .ZN(n18772) );
INV_X4 U16275 ( .A(n13892), .ZN(n18773) );
INV_X4 U16276 ( .A(n13886), .ZN(n18774) );
INV_X4 U16277 ( .A(n13880), .ZN(n18775) );
INV_X4 U16278 ( .A(n13874), .ZN(n18776) );
INV_X4 U16279 ( .A(n13868), .ZN(n18777) );
INV_X4 U16280 ( .A(n13862), .ZN(n18778) );
INV_X4 U16281 ( .A(n13856), .ZN(n18779) );
INV_X4 U16282 ( .A(n13850), .ZN(n18780) );
INV_X4 U16283 ( .A(n13844), .ZN(n18781) );
INV_X4 U16284 ( .A(n13838), .ZN(n18782) );
INV_X4 U16285 ( .A(n13832), .ZN(n18783) );
INV_X4 U16286 ( .A(n13826), .ZN(n18784) );
INV_X4 U16287 ( .A(n13820), .ZN(n18785) );
INV_X4 U16288 ( .A(n13814), .ZN(n18786) );
INV_X4 U16289 ( .A(n13808), .ZN(n18787) );
INV_X4 U16290 ( .A(n13802), .ZN(n18788) );
INV_X4 U16291 ( .A(n13796), .ZN(n18789) );
INV_X4 U16292 ( .A(n13790), .ZN(n18790) );
INV_X4 U16293 ( .A(n13784), .ZN(n18791) );
INV_X4 U16294 ( .A(n13778), .ZN(n18792) );
INV_X4 U16295 ( .A(n13772), .ZN(n18793) );
INV_X4 U16296 ( .A(n13766), .ZN(n18794) );
INV_X4 U16297 ( .A(n13760), .ZN(n18795) );
INV_X4 U16298 ( .A(n13754), .ZN(n18796) );
INV_X4 U16299 ( .A(n13748), .ZN(n18797) );
INV_X4 U16300 ( .A(n13742), .ZN(n18798) );
INV_X4 U16301 ( .A(n13736), .ZN(n18799) );
INV_X4 U16302 ( .A(n13730), .ZN(n18800) );
INV_X4 U16303 ( .A(n13724), .ZN(n18801) );
INV_X4 U16304 ( .A(n13718), .ZN(n18802) );
INV_X4 U16305 ( .A(n13712), .ZN(n18803) );
INV_X4 U16306 ( .A(n13706), .ZN(n18804) );
INV_X4 U16307 ( .A(n13700), .ZN(n18805) );
INV_X4 U16308 ( .A(n13694), .ZN(n18806) );
INV_X4 U16309 ( .A(n13688), .ZN(n18807) );
INV_X4 U16310 ( .A(n13682), .ZN(n18808) );
INV_X4 U16311 ( .A(n13676), .ZN(n18809) );
INV_X4 U16312 ( .A(n13669), .ZN(n18810) );
INV_X4 U16313 ( .A(n13662), .ZN(n18811) );
INV_X4 U16314 ( .A(n13654), .ZN(n18812) );
INV_X4 U16315 ( .A(n13648), .ZN(n18813) );
INV_X4 U16316 ( .A(n13642), .ZN(n18814) );
INV_X4 U16317 ( .A(n13636), .ZN(n18815) );
INV_X4 U16318 ( .A(n13630), .ZN(n18816) );
INV_X4 U16319 ( .A(n13624), .ZN(n18817) );
INV_X4 U16320 ( .A(n13618), .ZN(n18818) );
INV_X4 U16321 ( .A(n13612), .ZN(n18819) );
INV_X4 U16322 ( .A(n13558), .ZN(n18820) );
INV_X4 U16323 ( .A(n13552), .ZN(n18821) );
INV_X4 U16324 ( .A(n13546), .ZN(n18822) );
INV_X4 U16325 ( .A(n13540), .ZN(n18823) );
INV_X4 U16326 ( .A(n13534), .ZN(n18824) );
INV_X4 U16327 ( .A(n13528), .ZN(n18825) );
INV_X4 U16328 ( .A(n13522), .ZN(n18826) );
INV_X4 U16329 ( .A(n13516), .ZN(n18827) );
INV_X4 U16330 ( .A(n13462), .ZN(n18828) );
INV_X4 U16331 ( .A(n13456), .ZN(n18829) );
INV_X4 U16332 ( .A(n13450), .ZN(n18830) );
INV_X4 U16333 ( .A(n13444), .ZN(n18831) );
INV_X4 U16334 ( .A(n13438), .ZN(n18832) );
INV_X4 U16335 ( .A(n13432), .ZN(n18833) );
INV_X4 U16336 ( .A(n13426), .ZN(n18834) );
INV_X4 U16337 ( .A(n13420), .ZN(n18835) );
INV_X4 U16338 ( .A(aes_text_out[15]), .ZN(n18836) );
INV_X4 U16339 ( .A(aes_text_out[14]), .ZN(n18837) );
INV_X4 U16340 ( .A(aes_text_out[13]), .ZN(n18838) );
INV_X4 U16341 ( .A(aes_text_out[12]), .ZN(n18839) );
INV_X4 U16342 ( .A(aes_text_out[11]), .ZN(n18840) );
INV_X4 U16343 ( .A(aes_text_out[10]), .ZN(n18841) );
INV_X4 U16344 ( .A(aes_text_out[9]), .ZN(n18842) );
INV_X4 U16345 ( .A(aes_text_out[8]), .ZN(n18843) );
INV_X4 U16346 ( .A(n16837), .ZN(n18845) );
INV_X4 U16347 ( .A(n11957), .ZN(n18846) );
INV_X4 U16348 ( .A(n11929), .ZN(n18892) );
INV_X4 U16349 ( .A(n14166), .ZN(n19023) );
INV_X4 U16350 ( .A(n14199), .ZN(n19024) );
INV_X4 U16351 ( .A(n14228), .ZN(n19025) );
INV_X4 U16352 ( .A(n14257), .ZN(n19026) );
INV_X4 U16353 ( .A(n14286), .ZN(n19027) );
INV_X4 U16354 ( .A(n14315), .ZN(n19028) );
INV_X4 U16355 ( .A(n14344), .ZN(n19029) );
INV_X4 U16356 ( .A(n14373), .ZN(n19030) );
INV_X4 U16357 ( .A(n14190), .ZN(n19031) );
INV_X4 U16358 ( .A(n17539), .ZN(n19032) );
INV_X4 U16359 ( .A(n14219), .ZN(n19033) );
INV_X4 U16360 ( .A(n17541), .ZN(n19034) );
INV_X4 U16361 ( .A(n14248), .ZN(n19035) );
INV_X4 U16362 ( .A(n17543), .ZN(n19036) );
INV_X4 U16363 ( .A(n14277), .ZN(n19037) );
INV_X4 U16364 ( .A(n17545), .ZN(n19038) );
INV_X4 U16365 ( .A(n14306), .ZN(n19039) );
INV_X4 U16366 ( .A(n17547), .ZN(n19040) );
INV_X4 U16367 ( .A(n14335), .ZN(n19041) );
INV_X4 U16368 ( .A(n17549), .ZN(n19042) );
INV_X4 U16369 ( .A(n14364), .ZN(n19043) );
INV_X4 U16370 ( .A(n17551), .ZN(n19044) );
INV_X4 U16371 ( .A(n14396), .ZN(n19045) );
INV_X4 U16372 ( .A(n17553), .ZN(n19046) );
INV_X4 U16373 ( .A(n14191), .ZN(n19047) );
INV_X4 U16374 ( .A(n17555), .ZN(n19048) );
INV_X4 U16375 ( .A(n14220), .ZN(n19049) );
INV_X4 U16376 ( .A(n17557), .ZN(n19050) );
INV_X4 U16377 ( .A(n14249), .ZN(n19051) );
INV_X4 U16378 ( .A(n17559), .ZN(n19052) );
INV_X4 U16379 ( .A(n14278), .ZN(n19053) );
INV_X4 U16380 ( .A(n17561), .ZN(n19054) );
INV_X4 U16381 ( .A(n14307), .ZN(n19055) );
INV_X4 U16382 ( .A(n17563), .ZN(n19056) );
INV_X4 U16383 ( .A(n14336), .ZN(n19057) );
INV_X4 U16384 ( .A(n17745), .ZN(n19058) );
INV_X4 U16385 ( .A(n14365), .ZN(n19059) );
INV_X4 U16386 ( .A(n17565), .ZN(n19060) );
INV_X4 U16387 ( .A(n14397), .ZN(n19061) );
INV_X4 U16388 ( .A(n17567), .ZN(n19062) );
INV_X4 U16389 ( .A(n14417), .ZN(n19063) );
INV_X4 U16390 ( .A(n17569), .ZN(n19064) );
INV_X4 U16391 ( .A(n14440), .ZN(n19065) );
INV_X4 U16392 ( .A(n17571), .ZN(n19066) );
INV_X4 U16393 ( .A(n14462), .ZN(n19067) );
INV_X4 U16394 ( .A(n17573), .ZN(n19068) );
INV_X4 U16395 ( .A(n14484), .ZN(n19069) );
INV_X4 U16396 ( .A(n17575), .ZN(n19070) );
INV_X4 U16397 ( .A(n14506), .ZN(n19071) );
INV_X4 U16398 ( .A(n17577), .ZN(n19072) );
INV_X4 U16399 ( .A(n14528), .ZN(n19073) );
INV_X4 U16400 ( .A(n17579), .ZN(n19074) );
INV_X4 U16401 ( .A(n14550), .ZN(n19075) );
INV_X4 U16402 ( .A(n17581), .ZN(n19076) );
INV_X4 U16403 ( .A(n14574), .ZN(n19077) );
INV_X4 U16404 ( .A(n17583), .ZN(n19078) );
INV_X4 U16405 ( .A(n14185), .ZN(n19079) );
INV_X4 U16406 ( .A(n14597), .ZN(n19080) );
INV_X4 U16407 ( .A(n17585), .ZN(n19081) );
INV_X4 U16408 ( .A(n14216), .ZN(n19082) );
INV_X4 U16409 ( .A(n14618), .ZN(n19083) );
INV_X4 U16410 ( .A(n17587), .ZN(n19084) );
INV_X4 U16411 ( .A(n14245), .ZN(n19085) );
INV_X4 U16412 ( .A(n14639), .ZN(n19086) );
INV_X4 U16413 ( .A(n17589), .ZN(n19087) );
INV_X4 U16414 ( .A(n14274), .ZN(n19088) );
INV_X4 U16415 ( .A(n14660), .ZN(n19089) );
INV_X4 U16416 ( .A(n17591), .ZN(n19090) );
INV_X4 U16417 ( .A(n14303), .ZN(n19091) );
INV_X4 U16418 ( .A(n14681), .ZN(n19092) );
INV_X4 U16419 ( .A(n17593), .ZN(n19093) );
INV_X4 U16420 ( .A(n14332), .ZN(n19094) );
INV_X4 U16421 ( .A(n14702), .ZN(n19095) );
INV_X4 U16422 ( .A(n17595), .ZN(n19096) );
INV_X4 U16423 ( .A(n14361), .ZN(n19097) );
INV_X4 U16424 ( .A(n14723), .ZN(n19098) );
INV_X4 U16425 ( .A(n17597), .ZN(n19099) );
INV_X4 U16426 ( .A(n14391), .ZN(n19100) );
INV_X4 U16427 ( .A(n14746), .ZN(n19101) );
INV_X4 U16428 ( .A(n17599), .ZN(n19102) );
INV_X4 U16429 ( .A(n14421), .ZN(n19103) );
INV_X4 U16430 ( .A(n14768), .ZN(n19104) );
INV_X4 U16431 ( .A(n17601), .ZN(n19105) );
INV_X4 U16432 ( .A(n14444), .ZN(n19106) );
INV_X4 U16433 ( .A(n14791), .ZN(n19107) );
INV_X4 U16434 ( .A(n17603), .ZN(n19108) );
INV_X4 U16435 ( .A(n14466), .ZN(n19109) );
INV_X4 U16436 ( .A(n14813), .ZN(n19110) );
INV_X4 U16437 ( .A(n17605), .ZN(n19111) );
INV_X4 U16438 ( .A(n14488), .ZN(n19112) );
INV_X4 U16439 ( .A(n14835), .ZN(n19113) );
INV_X4 U16440 ( .A(n17607), .ZN(n19114) );
INV_X4 U16441 ( .A(n14510), .ZN(n19115) );
INV_X4 U16442 ( .A(n14857), .ZN(n19116) );
INV_X4 U16443 ( .A(n17609), .ZN(n19117) );
INV_X4 U16444 ( .A(n14532), .ZN(n19118) );
INV_X4 U16445 ( .A(n14879), .ZN(n19119) );
INV_X4 U16446 ( .A(n17611), .ZN(n19120) );
INV_X4 U16447 ( .A(n14554), .ZN(n19121) );
INV_X4 U16448 ( .A(n14901), .ZN(n19122) );
INV_X4 U16449 ( .A(n17613), .ZN(n19123) );
INV_X4 U16450 ( .A(n14578), .ZN(n19124) );
INV_X4 U16451 ( .A(n14924), .ZN(n19125) );
INV_X4 U16452 ( .A(n17615), .ZN(n19126) );
INV_X4 U16453 ( .A(n14773), .ZN(n19127) );
INV_X4 U16454 ( .A(n14795), .ZN(n19128) );
INV_X4 U16455 ( .A(n14817), .ZN(n19129) );
INV_X4 U16456 ( .A(n14839), .ZN(n19130) );
INV_X4 U16457 ( .A(n14861), .ZN(n19131) );
INV_X4 U16458 ( .A(n14883), .ZN(n19132) );
INV_X4 U16459 ( .A(n14905), .ZN(n19133) );
INV_X4 U16460 ( .A(n14928), .ZN(n19134) );
INV_X4 U16461 ( .A(n17633), .ZN(n19135) );
INV_X4 U16462 ( .A(n17635), .ZN(n19136) );
INV_X4 U16463 ( .A(n17637), .ZN(n19137) );
INV_X4 U16464 ( .A(n17639), .ZN(n19138) );
INV_X4 U16465 ( .A(n17641), .ZN(n19139) );
INV_X4 U16466 ( .A(n17643), .ZN(n19140) );
INV_X4 U16467 ( .A(n17645), .ZN(n19141) );
INV_X4 U16468 ( .A(n17647), .ZN(n19142) );
INV_X4 U16469 ( .A(n17649), .ZN(n19143) );
INV_X4 U16470 ( .A(n17651), .ZN(n19144) );
INV_X4 U16471 ( .A(n17653), .ZN(n19145) );
INV_X4 U16472 ( .A(n17655), .ZN(n19146) );
INV_X4 U16473 ( .A(n17657), .ZN(n19147) );
INV_X4 U16474 ( .A(n17659), .ZN(n19148) );
INV_X4 U16475 ( .A(n17661), .ZN(n19149) );
INV_X4 U16476 ( .A(n17663), .ZN(n19150) );
INV_X4 U16477 ( .A(n17665), .ZN(n19151) );
INV_X4 U16478 ( .A(n17667), .ZN(n19152) );
INV_X4 U16479 ( .A(n17669), .ZN(n19153) );
INV_X4 U16480 ( .A(n17671), .ZN(n19154) );
INV_X4 U16481 ( .A(n17673), .ZN(n19155) );
INV_X4 U16482 ( .A(n17675), .ZN(n19156) );
INV_X4 U16483 ( .A(n17677), .ZN(n19157) );
INV_X4 U16484 ( .A(n17679), .ZN(n19158) );
INV_X4 U16485 ( .A(n17681), .ZN(n19159) );
INV_X4 U16486 ( .A(n17683), .ZN(n19160) );
INV_X4 U16487 ( .A(n17685), .ZN(n19161) );
INV_X4 U16488 ( .A(n17687), .ZN(n19162) );
INV_X4 U16489 ( .A(n17689), .ZN(n19163) );
INV_X4 U16490 ( .A(n17691), .ZN(n19164) );
INV_X4 U16491 ( .A(n17693), .ZN(n19165) );
INV_X4 U16492 ( .A(n17695), .ZN(n19166) );
INV_X4 U16493 ( .A(n17697), .ZN(n19167) );
INV_X4 U16494 ( .A(n17699), .ZN(n19168) );
INV_X4 U16495 ( .A(n17701), .ZN(n19169) );
INV_X4 U16496 ( .A(n17703), .ZN(n19170) );
INV_X4 U16497 ( .A(n17705), .ZN(n19171) );
INV_X4 U16498 ( .A(n17707), .ZN(n19172) );
INV_X4 U16499 ( .A(n17709), .ZN(n19173) );
INV_X4 U16500 ( .A(n17711), .ZN(n19174) );
INV_X4 U16501 ( .A(n17713), .ZN(n19175) );
INV_X4 U16502 ( .A(n17715), .ZN(n19176) );
INV_X4 U16503 ( .A(n17717), .ZN(n19177) );
INV_X4 U16504 ( .A(n17719), .ZN(n19178) );
INV_X4 U16505 ( .A(n17721), .ZN(n19179) );
INV_X4 U16506 ( .A(n17723), .ZN(n19180) );
INV_X4 U16507 ( .A(n17725), .ZN(n19181) );
INV_X4 U16508 ( .A(n17727), .ZN(n19182) );
INV_X4 U16509 ( .A(n17728), .ZN(n19183) );
INV_X4 U16510 ( .A(n17729), .ZN(n19184) );
INV_X4 U16511 ( .A(n17730), .ZN(n19185) );
INV_X4 U16512 ( .A(n17731), .ZN(n19186) );
INV_X4 U16513 ( .A(n17732), .ZN(n19187) );
INV_X4 U16514 ( .A(n17733), .ZN(n19188) );
INV_X4 U16515 ( .A(n17734), .ZN(n19189) );
INV_X4 U16516 ( .A(n17735), .ZN(n19190) );
INV_X4 U16517 ( .A(n17736), .ZN(n19191) );
INV_X4 U16518 ( .A(n17737), .ZN(n19192) );
INV_X4 U16519 ( .A(n17738), .ZN(n19193) );
INV_X4 U16520 ( .A(n17739), .ZN(n19194) );
INV_X4 U16521 ( .A(n17740), .ZN(n19195) );
INV_X4 U16522 ( .A(n17741), .ZN(n19196) );
INV_X4 U16523 ( .A(n17742), .ZN(n19197) );
INV_X4 U16524 ( .A(n17743), .ZN(n19198) );
INV_X4 U16525 ( .A(n15272), .ZN(n19199) );
INV_X4 U16526 ( .A(n14736), .ZN(n19200) );
INV_X4 U16527 ( .A(n15094), .ZN(n19201) );
INV_X4 U16528 ( .A(n16542), .ZN(n19203) );
INV_X4 U16529 ( .A(dii_data_size[1]), .ZN(n19204) );
INV_X4 U16530 ( .A(dii_data_size[0]), .ZN(n19205) );
INV_X4 U16531 ( .A(cii_ctl_vld), .ZN(n19206) );
INV_X4 _GFM_U4594  ( .A(v_in[127]), .ZN(_GFM_n2699 ) );
INV_X4 _GFM_U4593  ( .A(v_in[125]), .ZN(_GFM_n26980 ) );
INV_X4 _GFM_U4592  ( .A(v_in[124]), .ZN(_GFM_n2697 ) );
INV_X4 _GFM_U4591  ( .A(v_in[123]), .ZN(_GFM_n2696 ) );
INV_X4 _GFM_U4590  ( .A(v_in[122]), .ZN(_GFM_n2695 ) );
INV_X4 _GFM_U4589  ( .A(v_out[123]), .ZN(_GFM_n2585 ) );
INV_X4 _GFM_U4588  ( .A(v_out[122]), .ZN(_GFM_n25830 ) );
INV_X4 _GFM_U4587  ( .A(v_out[121]), .ZN(_GFM_n25810 ) );
INV_X4 _GFM_U4586  ( .A(_GFM_N4250 ), .ZN(_GFM_n2579 ) );
INV_X4 _GFM_U4585  ( .A(_GFM_N4248 ), .ZN(_GFM_n25770 ) );
INV_X4 _GFM_U4584  ( .A(v_out[118]), .ZN(_GFM_n2575 ) );
INV_X4 _GFM_U4583  ( .A(_GFM_N4254 ), .ZN(_GFM_n25740 ) );
INV_X4 _GFM_U4582  ( .A(v_out[117]), .ZN(_GFM_n2572 ) );
INV_X4 _GFM_U4581  ( .A(_GFM_N4257 ), .ZN(_GFM_n2571 ) );
INV_X4 _GFM_U4580  ( .A(v_out[116]), .ZN(_GFM_n25690 ) );
INV_X4 _GFM_U4579  ( .A(_GFM_N4242 ), .ZN(_GFM_n2568 ) );
INV_X4 _GFM_U4578  ( .A(v_in[4]), .ZN(_GFM_n25660 ) );
INV_X4 _GFM_U4577  ( .A(v_out[115]), .ZN(_GFM_n2565 ) );
INV_X4 _GFM_U4576  ( .A(_GFM_N4239 ), .ZN(_GFM_n2564 ) );
INV_X4 _GFM_U4575  ( .A(v_in[3]), .ZN(_GFM_n25620 ) );
INV_X4 _GFM_U4574  ( .A(v_out[114]), .ZN(_GFM_n25611 ) );
INV_X4 _GFM_U4573  ( .A(_GFM_N4232 ), .ZN(_GFM_n25600 ) );
INV_X4 _GFM_U4572  ( .A(v_in[2]), .ZN(_GFM_n25580 ) );
INV_X4 _GFM_U4571  ( .A(v_out[113]), .ZN(_GFM_n25570 ) );
INV_X4 _GFM_U4570  ( .A(_GFM_N4235 ), .ZN(_GFM_n2556 ) );
INV_X4 _GFM_U4569  ( .A(v_in[1]), .ZN(_GFM_n2554 ) );
INV_X4 _GFM_U4568  ( .A(b_in[115]), .ZN(_GFM_n25530 ) );
INV_X4 _GFM_U4567  ( .A(_GFM_N4224 ), .ZN(_GFM_n25500 ) );
INV_X4 _GFM_U4566  ( .A(v_out[112]), .ZN(_GFM_n25490 ) );
INV_X4 _GFM_U4565  ( .A(_GFM_N4227 ), .ZN(_GFM_n2548 ) );
INV_X4 _GFM_U4564  ( .A(v_in[0]), .ZN(_GFM_n25460 ) );
BUF_X4 _GFM_U4563  ( .A(v_in[98]), .Z(v_out[82]) );
BUF_X4 _GFM_U4562  ( .A(v_in[99]), .Z(v_out[83]) );
BUF_X4 _GFM_U4561  ( .A(v_in[100]), .Z(v_out[84]) );
BUF_X4 _GFM_U4560  ( .A(v_in[101]), .Z(v_out[85]) );
BUF_X4 _GFM_U4559  ( .A(v_in[102]), .Z(v_out[86]) );
BUF_X4 _GFM_U4558  ( .A(v_in[103]), .Z(v_out[87]) );
BUF_X4 _GFM_U4557  ( .A(v_in[104]), .Z(v_out[88]) );
BUF_X4 _GFM_U4556  ( .A(v_in[105]), .Z(v_out[89]) );
BUF_X4 _GFM_U4555  ( .A(v_in[106]), .Z(v_out[90]) );
BUF_X4 _GFM_U4554  ( .A(v_in[107]), .Z(v_out[91]) );
BUF_X4 _GFM_U4553  ( .A(v_in[108]), .Z(v_out[92]) );
BUF_X4 _GFM_U4552  ( .A(v_in[109]), .Z(v_out[93]) );
BUF_X4 _GFM_U4551  ( .A(v_in[110]), .Z(v_out[94]) );
BUF_X4 _GFM_U4550  ( .A(v_in[111]), .Z(v_out[95]) );
BUF_X4 _GFM_U4549  ( .A(v_in[112]), .Z(v_out[96]) );
BUF_X4 _GFM_U4548  ( .A(v_in[113]), .Z(v_out[97]) );
BUF_X4 _GFM_U4547  ( .A(v_in[114]), .Z(v_out[98]) );
BUF_X4 _GFM_U4546  ( .A(v_in[115]), .Z(v_out[99]) );
BUF_X4 _GFM_U4545  ( .A(v_in[116]), .Z(v_out[100]) );
BUF_X4 _GFM_U4544  ( .A(v_in[117]), .Z(v_out[101]) );
BUF_X4 _GFM_U4543  ( .A(v_in[118]), .Z(v_out[102]) );
BUF_X4 _GFM_U4542  ( .A(v_in[119]), .Z(v_out[103]) );
BUF_X4 _GFM_U4541  ( .A(v_in[120]), .Z(v_out[104]) );
INV_X4 _GFM_U4540  ( .A(v_in[36]), .ZN(_GFM_n2610 ) );
INV_X4 _GFM_U4539  ( .A(v_in[34]), .ZN(_GFM_n26080 ) );
INV_X4 _GFM_U4538  ( .A(v_in[33]), .ZN(_GFM_n26070 ) );
INV_X4 _GFM_U4537  ( .A(v_in[32]), .ZN(_GFM_n2606 ) );
INV_X4 _GFM_U4536  ( .A(v_in[46]), .ZN(_GFM_n26200 ) );
INV_X4 _GFM_U4535  ( .A(v_in[45]), .ZN(_GFM_n26190 ) );
INV_X4 _GFM_U4534  ( .A(v_in[43]), .ZN(_GFM_n2617 ) );
INV_X4 _GFM_U4533  ( .A(v_in[44]), .ZN(_GFM_n2618 ) );
INV_X4 _GFM_U4532  ( .A(v_in[38]), .ZN(_GFM_n26120 ) );
INV_X4 _GFM_U4531  ( .A(v_in[39]), .ZN(_GFM_n2613 ) );
INV_X4 _GFM_U4530  ( .A(v_in[42]), .ZN(_GFM_n2616 ) );
INV_X4 _GFM_U4529  ( .A(v_in[40]), .ZN(_GFM_n26140 ) );
INV_X4 _GFM_U4528  ( .A(v_in[41]), .ZN(_GFM_n26150 ) );
INV_X4 _GFM_U4527  ( .A(v_in[37]), .ZN(_GFM_n26110 ) );
INV_X4 _GFM_U4526  ( .A(v_in[16]), .ZN(_GFM_n25901 ) );
INV_X4 _GFM_U4525  ( .A(v_in[17]), .ZN(_GFM_n25910 ) );
INV_X4 _GFM_U4524  ( .A(v_in[18]), .ZN(_GFM_n2592 ) );
INV_X4 _GFM_U4523  ( .A(v_in[19]), .ZN(_GFM_n25930 ) );
INV_X4 _GFM_U4522  ( .A(v_in[20]), .ZN(_GFM_n25940 ) );
INV_X4 _GFM_U4521  ( .A(v_in[21]), .ZN(_GFM_n2595 ) );
INV_X4 _GFM_U4520  ( .A(v_in[22]), .ZN(_GFM_n2596 ) );
INV_X4 _GFM_U4519  ( .A(v_in[23]), .ZN(_GFM_n25970 ) );
INV_X4 _GFM_U4518  ( .A(v_in[24]), .ZN(_GFM_n25980 ) );
INV_X4 _GFM_U4517  ( .A(v_in[25]), .ZN(_GFM_n2599 ) );
INV_X4 _GFM_U4516  ( .A(v_in[26]), .ZN(_GFM_n26000 ) );
INV_X4 _GFM_U4515  ( .A(v_in[27]), .ZN(_GFM_n26010 ) );
INV_X4 _GFM_U4514  ( .A(v_in[28]), .ZN(_GFM_n2602 ) );
INV_X4 _GFM_U4513  ( .A(v_in[29]), .ZN(_GFM_n2603 ) );
INV_X4 _GFM_U4512  ( .A(v_in[30]), .ZN(_GFM_n2604 ) );
INV_X4 _GFM_U4511  ( .A(v_in[31]), .ZN(_GFM_n26050 ) );
INV_X4 _GFM_U4510  ( .A(v_in[35]), .ZN(_GFM_n2609 ) );
INV_X4 _GFM_U4509  ( .A(v_in[47]), .ZN(_GFM_n2621 ) );
INV_X4 _GFM_U4508  ( .A(v_in[48]), .ZN(_GFM_n26220 ) );
INV_X4 _GFM_U4507  ( .A(v_in[49]), .ZN(_GFM_n2623 ) );
INV_X4 _GFM_U4506  ( .A(v_in[50]), .ZN(_GFM_n26240 ) );
INV_X4 _GFM_U4505  ( .A(v_in[51]), .ZN(_GFM_n26250 ) );
INV_X4 _GFM_U4504  ( .A(v_in[52]), .ZN(_GFM_n2626 ) );
INV_X4 _GFM_U4503  ( .A(v_in[53]), .ZN(_GFM_n2627 ) );
INV_X4 _GFM_U4502  ( .A(v_in[54]), .ZN(_GFM_n26280 ) );
INV_X4 _GFM_U4501  ( .A(v_in[55]), .ZN(_GFM_n26290 ) );
INV_X4 _GFM_U4500  ( .A(v_in[56]), .ZN(_GFM_n26301 ) );
INV_X4 _GFM_U4499  ( .A(v_in[57]), .ZN(_GFM_n26310 ) );
INV_X4 _GFM_U4498  ( .A(v_in[58]), .ZN(_GFM_n26320 ) );
INV_X4 _GFM_U4497  ( .A(v_in[59]), .ZN(_GFM_n2633 ) );
INV_X4 _GFM_U4496  ( .A(v_in[60]), .ZN(_GFM_n2634 ) );
INV_X4 _GFM_U4495  ( .A(v_in[61]), .ZN(_GFM_n2635 ) );
INV_X4 _GFM_U4494  ( .A(v_in[62]), .ZN(_GFM_n26360 ) );
INV_X4 _GFM_U4493  ( .A(v_in[63]), .ZN(_GFM_n2637 ) );
INV_X4 _GFM_U4492  ( .A(v_in[64]), .ZN(_GFM_n26380 ) );
INV_X4 _GFM_U4491  ( .A(v_in[68]), .ZN(_GFM_n26420 ) );
INV_X4 _GFM_U4490  ( .A(v_in[69]), .ZN(_GFM_n26430 ) );
INV_X4 _GFM_U4489  ( .A(v_in[70]), .ZN(_GFM_n2644 ) );
INV_X4 _GFM_U4488  ( .A(v_in[71]), .ZN(_GFM_n26450 ) );
INV_X4 _GFM_U4487  ( .A(v_in[72]), .ZN(_GFM_n26460 ) );
INV_X4 _GFM_U4486  ( .A(v_in[73]), .ZN(_GFM_n2647 ) );
INV_X4 _GFM_U4485  ( .A(v_in[74]), .ZN(_GFM_n2648 ) );
INV_X4 _GFM_U4484  ( .A(v_in[75]), .ZN(_GFM_n2649 ) );
INV_X4 _GFM_U4483  ( .A(v_in[76]), .ZN(_GFM_n26500 ) );
INV_X4 _GFM_U4482  ( .A(v_in[77]), .ZN(_GFM_n26510 ) );
INV_X4 _GFM_U4481  ( .A(v_in[78]), .ZN(_GFM_n2652 ) );
INV_X4 _GFM_U4480  ( .A(v_in[79]), .ZN(_GFM_n26530 ) );
INV_X4 _GFM_U4479  ( .A(v_in[80]), .ZN(_GFM_n2654 ) );
INV_X4 _GFM_U4478  ( .A(v_in[81]), .ZN(_GFM_n26550 ) );
INV_X4 _GFM_U4477  ( .A(v_in[82]), .ZN(_GFM_n26560 ) );
INV_X4 _GFM_U4476  ( .A(v_in[83]), .ZN(_GFM_n2657 ) );
INV_X4 _GFM_U4475  ( .A(v_in[84]), .ZN(_GFM_n2658 ) );
INV_X4 _GFM_U4474  ( .A(v_in[85]), .ZN(_GFM_n26590 ) );
INV_X4 _GFM_U4473  ( .A(v_in[86]), .ZN(_GFM_n26600 ) );
INV_X4 _GFM_U4472  ( .A(v_in[87]), .ZN(_GFM_n26611 ) );
INV_X4 _GFM_U4471  ( .A(v_in[88]), .ZN(_GFM_n26620 ) );
INV_X4 _GFM_U4470  ( .A(v_in[89]), .ZN(_GFM_n26630 ) );
INV_X4 _GFM_U4469  ( .A(v_in[90]), .ZN(_GFM_n2664 ) );
INV_X4 _GFM_U4468  ( .A(v_in[91]), .ZN(_GFM_n2665 ) );
INV_X4 _GFM_U4467  ( .A(v_in[92]), .ZN(_GFM_n2666 ) );
INV_X4 _GFM_U4466  ( .A(v_in[93]), .ZN(_GFM_n26670 ) );
INV_X4 _GFM_U4465  ( .A(v_in[94]), .ZN(_GFM_n2668 ) );
INV_X4 _GFM_U4464  ( .A(v_in[95]), .ZN(_GFM_n26690 ) );
INV_X4 _GFM_U4463  ( .A(v_in[96]), .ZN(_GFM_n26700 ) );
INV_X4 _GFM_U4462  ( .A(v_in[97]), .ZN(_GFM_n2671 ) );
INV_X4 _GFM_U4461  ( .A(v_in[98]), .ZN(_GFM_n2672 ) );
INV_X4 _GFM_U4460  ( .A(v_in[99]), .ZN(_GFM_n26730 ) );
INV_X4 _GFM_U4459  ( .A(v_in[100]), .ZN(_GFM_n26740 ) );
INV_X4 _GFM_U4458  ( .A(v_in[101]), .ZN(_GFM_n2675 ) );
INV_X4 _GFM_U4457  ( .A(v_in[102]), .ZN(_GFM_n26760 ) );
INV_X4 _GFM_U4456  ( .A(v_in[103]), .ZN(_GFM_n26770 ) );
INV_X4 _GFM_U4455  ( .A(v_in[104]), .ZN(_GFM_n2678 ) );
INV_X4 _GFM_U4454  ( .A(v_in[105]), .ZN(_GFM_n2679 ) );
INV_X4 _GFM_U4453  ( .A(v_in[106]), .ZN(_GFM_n26801 ) );
INV_X4 _GFM_U4452  ( .A(v_in[107]), .ZN(_GFM_n26810 ) );
INV_X4 _GFM_U4451  ( .A(v_in[108]), .ZN(_GFM_n26820 ) );
INV_X4 _GFM_U4450  ( .A(v_in[109]), .ZN(_GFM_n2683 ) );
INV_X4 _GFM_U4449  ( .A(v_in[110]), .ZN(_GFM_n26840 ) );
INV_X4 _GFM_U4448  ( .A(v_in[111]), .ZN(_GFM_n2685 ) );
INV_X4 _GFM_U4447  ( .A(v_in[112]), .ZN(_GFM_n26860 ) );
INV_X4 _GFM_U4446  ( .A(v_in[113]), .ZN(_GFM_n26870 ) );
INV_X4 _GFM_U4445  ( .A(v_in[114]), .ZN(_GFM_n2688 ) );
INV_X4 _GFM_U4444  ( .A(v_in[115]), .ZN(_GFM_n2689 ) );
INV_X4 _GFM_U4443  ( .A(v_in[116]), .ZN(_GFM_n26900 ) );
INV_X4 _GFM_U4442  ( .A(v_in[117]), .ZN(_GFM_n26910 ) );
INV_X4 _GFM_U4441  ( .A(v_in[118]), .ZN(_GFM_n26921 ) );
INV_X4 _GFM_U4440  ( .A(v_in[119]), .ZN(_GFM_n26930 ) );
INV_X4 _GFM_U4439  ( .A(v_in[120]), .ZN(_GFM_n26940 ) );
BUF_X4 _GFM_U4438  ( .A(v_in[16]), .Z(v_out[0]) );
BUF_X4 _GFM_U4437  ( .A(v_in[17]), .Z(v_out[1]) );
BUF_X4 _GFM_U4436  ( .A(v_in[18]), .Z(v_out[2]) );
BUF_X4 _GFM_U4435  ( .A(v_in[19]), .Z(v_out[3]) );
BUF_X4 _GFM_U4434  ( .A(v_in[20]), .Z(v_out[4]) );
BUF_X4 _GFM_U4433  ( .A(v_in[21]), .Z(v_out[5]) );
BUF_X4 _GFM_U4432  ( .A(v_in[22]), .Z(v_out[6]) );
BUF_X4 _GFM_U4431  ( .A(v_in[23]), .Z(v_out[7]) );
BUF_X4 _GFM_U4430  ( .A(v_in[24]), .Z(v_out[8]) );
BUF_X4 _GFM_U4429  ( .A(v_in[25]), .Z(v_out[9]) );
BUF_X4 _GFM_U4428  ( .A(v_in[26]), .Z(v_out[10]) );
BUF_X4 _GFM_U4427  ( .A(v_in[27]), .Z(v_out[11]) );
BUF_X4 _GFM_U4426  ( .A(v_in[28]), .Z(v_out[12]) );
BUF_X4 _GFM_U4425  ( .A(v_in[29]), .Z(v_out[13]) );
BUF_X4 _GFM_U4424  ( .A(v_in[30]), .Z(v_out[14]) );
BUF_X4 _GFM_U4423  ( .A(v_in[31]), .Z(v_out[15]) );
BUF_X4 _GFM_U4422  ( .A(v_in[32]), .Z(v_out[16]) );
BUF_X4 _GFM_U4421  ( .A(v_in[33]), .Z(v_out[17]) );
BUF_X4 _GFM_U4420  ( .A(v_in[34]), .Z(v_out[18]) );
BUF_X4 _GFM_U4419  ( .A(v_in[35]), .Z(v_out[19]) );
BUF_X4 _GFM_U4418  ( .A(v_in[36]), .Z(v_out[20]) );
BUF_X4 _GFM_U4417  ( .A(v_in[37]), .Z(v_out[21]) );
BUF_X4 _GFM_U4416  ( .A(v_in[38]), .Z(v_out[22]) );
BUF_X4 _GFM_U4415  ( .A(v_in[39]), .Z(v_out[23]) );
BUF_X4 _GFM_U4414  ( .A(v_in[40]), .Z(v_out[24]) );
BUF_X4 _GFM_U4413  ( .A(v_in[41]), .Z(v_out[25]) );
BUF_X4 _GFM_U4412  ( .A(v_in[42]), .Z(v_out[26]) );
BUF_X4 _GFM_U4411  ( .A(v_in[43]), .Z(v_out[27]) );
BUF_X4 _GFM_U4410  ( .A(v_in[44]), .Z(v_out[28]) );
BUF_X4 _GFM_U4409  ( .A(v_in[45]), .Z(v_out[29]) );
BUF_X4 _GFM_U4408  ( .A(v_in[46]), .Z(v_out[30]) );
BUF_X4 _GFM_U4407  ( .A(v_in[47]), .Z(v_out[31]) );
BUF_X4 _GFM_U4406  ( .A(v_in[48]), .Z(v_out[32]) );
BUF_X4 _GFM_U4405  ( .A(v_in[49]), .Z(v_out[33]) );
BUF_X4 _GFM_U4404  ( .A(v_in[50]), .Z(v_out[34]) );
BUF_X4 _GFM_U4403  ( .A(v_in[51]), .Z(v_out[35]) );
BUF_X4 _GFM_U4402  ( .A(v_in[52]), .Z(v_out[36]) );
BUF_X4 _GFM_U4401  ( .A(v_in[53]), .Z(v_out[37]) );
BUF_X4 _GFM_U4400  ( .A(v_in[54]), .Z(v_out[38]) );
BUF_X4 _GFM_U4399  ( .A(v_in[55]), .Z(v_out[39]) );
BUF_X4 _GFM_U4398  ( .A(v_in[56]), .Z(v_out[40]) );
BUF_X4 _GFM_U4397  ( .A(v_in[57]), .Z(v_out[41]) );
BUF_X4 _GFM_U4396  ( .A(v_in[58]), .Z(v_out[42]) );
BUF_X4 _GFM_U4395  ( .A(v_in[59]), .Z(v_out[43]) );
BUF_X4 _GFM_U4394  ( .A(v_in[60]), .Z(v_out[44]) );
BUF_X4 _GFM_U4393  ( .A(v_in[61]), .Z(v_out[45]) );
BUF_X4 _GFM_U4392  ( .A(v_in[62]), .Z(v_out[46]) );
BUF_X4 _GFM_U4391  ( .A(v_in[63]), .Z(v_out[47]) );
BUF_X4 _GFM_U4390  ( .A(v_in[64]), .Z(v_out[48]) );
BUF_X4 _GFM_U4389  ( .A(v_in[65]), .Z(v_out[49]) );
BUF_X4 _GFM_U4388  ( .A(v_in[66]), .Z(v_out[50]) );
BUF_X4 _GFM_U4387  ( .A(v_in[67]), .Z(v_out[51]) );
BUF_X4 _GFM_U4386  ( .A(v_in[68]), .Z(v_out[52]) );
BUF_X4 _GFM_U4385  ( .A(v_in[69]), .Z(v_out[53]) );
BUF_X4 _GFM_U4384  ( .A(v_in[70]), .Z(v_out[54]) );
BUF_X4 _GFM_U4383  ( .A(v_in[71]), .Z(v_out[55]) );
BUF_X4 _GFM_U4382  ( .A(v_in[72]), .Z(v_out[56]) );
BUF_X4 _GFM_U4381  ( .A(v_in[73]), .Z(v_out[57]) );
BUF_X4 _GFM_U4380  ( .A(v_in[74]), .Z(v_out[58]) );
BUF_X4 _GFM_U4379  ( .A(v_in[75]), .Z(v_out[59]) );
BUF_X4 _GFM_U4378  ( .A(v_in[76]), .Z(v_out[60]) );
BUF_X4 _GFM_U4377  ( .A(v_in[77]), .Z(v_out[61]) );
BUF_X4 _GFM_U4376  ( .A(v_in[78]), .Z(v_out[62]) );
BUF_X4 _GFM_U4375  ( .A(v_in[79]), .Z(v_out[63]) );
BUF_X4 _GFM_U4374  ( .A(v_in[80]), .Z(v_out[64]) );
BUF_X4 _GFM_U4373  ( .A(v_in[81]), .Z(v_out[65]) );
BUF_X4 _GFM_U4372  ( .A(v_in[82]), .Z(v_out[66]) );
BUF_X4 _GFM_U4371  ( .A(v_in[83]), .Z(v_out[67]) );
BUF_X4 _GFM_U4370  ( .A(v_in[84]), .Z(v_out[68]) );
BUF_X4 _GFM_U4369  ( .A(v_in[85]), .Z(v_out[69]) );
BUF_X4 _GFM_U4368  ( .A(v_in[86]), .Z(v_out[70]) );
BUF_X4 _GFM_U4367  ( .A(v_in[87]), .Z(v_out[71]) );
BUF_X4 _GFM_U4366  ( .A(v_in[88]), .Z(v_out[72]) );
BUF_X4 _GFM_U4365  ( .A(v_in[89]), .Z(v_out[73]) );
BUF_X4 _GFM_U4364  ( .A(v_in[90]), .Z(v_out[74]) );
BUF_X4 _GFM_U4363  ( .A(v_in[91]), .Z(v_out[75]) );
BUF_X4 _GFM_U4362  ( .A(v_in[92]), .Z(v_out[76]) );
BUF_X4 _GFM_U4361  ( .A(v_in[93]), .Z(v_out[77]) );
BUF_X4 _GFM_U4360  ( .A(v_in[94]), .Z(v_out[78]) );
BUF_X4 _GFM_U4359  ( .A(v_in[95]), .Z(v_out[79]) );
BUF_X4 _GFM_U4358  ( .A(v_in[96]), .Z(v_out[80]) );
BUF_X4 _GFM_U4357  ( .A(v_in[97]), .Z(v_out[81]) );
NOR2_X2 _GFM_U4356  ( .A1(_GFM_n2409 ), .A2(_GFM_n2572 ), .ZN(_GFM_N3985 ));
NOR2_X2 _GFM_U4355  ( .A1(_GFM_n2697 ), .A2(_GFM_n2516 ), .ZN(_GFM_N4049 ));
NOR2_X2 _GFM_U4354  ( .A1(_GFM_n2695 ), .A2(_GFM_n25360 ), .ZN(_GFM_N4047 ));
NAND3_X2 _GFM_U4353  ( .A1(b_in[119]), .A2(_GFM_n25760 ), .A3(v_in[6]), .ZN(_GFM_n17911 ) );
BUF_X4 _GFM_U4352  ( .A(v_in[15]), .Z(v_out[127]) );
NAND3_X2 _GFM_U4351  ( .A1(b_in[115]), .A2(_GFM_n25840 ), .A3(v_in[10]),.ZN(_GFM_n17511 ) );
NAND3_X2 _GFM_U4350  ( .A1(b_in[116]), .A2(_GFM_n25821 ), .A3(v_in[9]), .ZN(_GFM_n18310 ) );
NAND3_X2 _GFM_U4349  ( .A1(b_in[117]), .A2(_GFM_n25800 ), .A3(v_in[8]), .ZN(_GFM_n2121 ) );
NAND3_X2 _GFM_U4348  ( .A1(b_in[118]), .A2(_GFM_n2578 ), .A3(v_in[7]), .ZN(_GFM_n181 ) );
NAND3_X2 _GFM_U4347  ( .A1(b_in[113]), .A2(_GFM_n2587 ), .A3(v_in[12]), .ZN(_GFM_n17310 ) );
NAND3_X2 _GFM_U4346  ( .A1(b_in[120]), .A2(_GFM_n2573 ), .A3(v_in[5]), .ZN(_GFM_n21230 ) );
NAND3_X2 _GFM_U4345  ( .A1(b_in[114]), .A2(_GFM_n2586 ), .A3(v_in[11]), .ZN(_GFM_n177 ) );
NAND3_X2 _GFM_U4344  ( .A1(b_in[126]), .A2(_GFM_n25460 ), .A3(v_in[127]),.ZN(_GFM_n21350 ) );
NAND3_X2 _GFM_U4343  ( .A1(v_in[3]), .A2(_GFM_n25660 ), .A3(b_in[122]), .ZN(_GFM_n21290 ) );
NAND3_X2 _GFM_U4342  ( .A1(b_in[112]), .A2(_GFM_n25880 ), .A3(v_in[13]),.ZN(_GFM_n17110 ) );
NAND3_X2 _GFM_U4341  ( .A1(v_in[4]), .A2(_GFM_n25700 ), .A3(b_in[121]), .ZN(_GFM_n2125 ) );
NAND3_X2 _GFM_U4340  ( .A1(v_in[2]), .A2(_GFM_n25620 ), .A3(b_in[123]), .ZN(_GFM_n2127 ) );
NAND3_X2 _GFM_U4339  ( .A1(v_in[1]), .A2(_GFM_n25580 ), .A3(b_in[124]), .ZN(_GFM_n2131 ) );
NAND3_X2 _GFM_U4338  ( .A1(v_in[0]), .A2(_GFM_n2554 ), .A3(b_in[125]), .ZN(_GFM_n21330 ) );
INV_X4 _GFM_U4337  ( .A(v_in[5]), .ZN(_GFM_n25700 ) );
INV_X4 _GFM_U4336  ( .A(v_in[6]), .ZN(_GFM_n2573 ) );
INV_X4 _GFM_U4335  ( .A(v_in[7]), .ZN(_GFM_n25760 ) );
INV_X4 _GFM_U4334  ( .A(v_in[8]), .ZN(_GFM_n2578 ) );
INV_X4 _GFM_U4333  ( .A(v_in[9]), .ZN(_GFM_n25800 ) );
INV_X4 _GFM_U4332  ( .A(v_in[65]), .ZN(_GFM_n26390 ) );
INV_X4 _GFM_U4331  ( .A(v_in[66]), .ZN(_GFM_n26401 ) );
INV_X4 _GFM_U4330  ( .A(v_in[67]), .ZN(_GFM_n2641 ) );
INV_X4 _GFM_U4329  ( .A(v_in[10]), .ZN(_GFM_n25821 ) );
INV_X4 _GFM_U2238  ( .A(v_in[15]), .ZN(_GFM_n25890 ) );
INV_X4 _GFM_U2237  ( .A(v_in[11]), .ZN(_GFM_n25840 ) );
NOR2_X2 _GFM_U2236  ( .A1(_GFM_n25890 ), .A2(_GFM_n2387 ), .ZN(_GFM_N28 ) );
NOR2_X2 _GFM_U2235  ( .A1(_GFM_n25890 ), .A2(_GFM_n23970 ), .ZN(_GFM_N58 ));
NOR2_X2 _GFM_U2234  ( .A1(_GFM_n23980 ), .A2(_GFM_n25901 ), .ZN(_GFM_N89 ));
NOR2_X2 _GFM_U2233  ( .A1(_GFM_n2406 ), .A2(_GFM_n25910 ), .ZN(_GFM_N120 ));
NOR2_X2 _GFM_U2232  ( .A1(_GFM_n24050 ), .A2(_GFM_n2592 ), .ZN(_GFM_N151 ));
NOR2_X2 _GFM_U2231  ( .A1(_GFM_n2404 ), .A2(_GFM_n25930 ), .ZN(_GFM_N182 ));
NOR2_X2 _GFM_U2230  ( .A1(_GFM_n24030 ), .A2(_GFM_n25940 ), .ZN(_GFM_N213 ));
NOR2_X2 _GFM_U2229  ( .A1(_GFM_n24030 ), .A2(_GFM_n2595 ), .ZN(_GFM_N244 ));
NOR2_X2 _GFM_U2228  ( .A1(_GFM_n24020 ), .A2(_GFM_n2596 ), .ZN(_GFM_N275 ));
NOR2_X2 _GFM_U2227  ( .A1(_GFM_n2401 ), .A2(_GFM_n25970 ), .ZN(_GFM_N306 ));
NOR2_X2 _GFM_U2226  ( .A1(_GFM_n2400 ), .A2(_GFM_n25980 ), .ZN(_GFM_N337 ));
NOR2_X2 _GFM_U2225  ( .A1(_GFM_n2400 ), .A2(_GFM_n2599 ), .ZN(_GFM_N368 ) );
NOR2_X2 _GFM_U2224  ( .A1(_GFM_n2399 ), .A2(_GFM_n26000 ), .ZN(_GFM_N399 ));
NOR2_X2 _GFM_U2223  ( .A1(_GFM_n2399 ), .A2(_GFM_n26010 ), .ZN(_GFM_N430 ));
NOR2_X2 _GFM_U2222  ( .A1(_GFM_n23980 ), .A2(_GFM_n2602 ), .ZN(_GFM_N461 ));
NOR2_X2 _GFM_U2221  ( .A1(_GFM_n2399 ), .A2(_GFM_n2603 ), .ZN(_GFM_N492 ) );
NOR2_X2 _GFM_U2220  ( .A1(_GFM_n23980 ), .A2(_GFM_n2604 ), .ZN(_GFM_N523 ));
NOR2_X2 _GFM_U2219  ( .A1(_GFM_n2606 ), .A2(_GFM_n2387 ), .ZN(_GFM_N555 ) );
NOR2_X2 _GFM_U2218  ( .A1(_GFM_n2606 ), .A2(_GFM_n23970 ), .ZN(_GFM_N585 ));
NOR2_X2 _GFM_U2217  ( .A1(_GFM_n26070 ), .A2(_GFM_n23970 ), .ZN(_GFM_N616 ));
NOR2_X2 _GFM_U2216  ( .A1(_GFM_n26080 ), .A2(_GFM_n23970 ), .ZN(_GFM_N647 ));
NOR2_X2 _GFM_U2215  ( .A1(_GFM_n2610 ), .A2(_GFM_n2387 ), .ZN(_GFM_N679 ) );
NOR2_X2 _GFM_U2214  ( .A1(_GFM_n2610 ), .A2(_GFM_n23970 ), .ZN(_GFM_N709 ));
NOR2_X2 _GFM_U2213  ( .A1(_GFM_n23980 ), .A2(_GFM_n26110 ), .ZN(_GFM_N740 ));
NOR2_X2 _GFM_U2212  ( .A1(_GFM_n23980 ), .A2(_GFM_n26120 ), .ZN(_GFM_N771 ));
NOR2_X2 _GFM_U2211  ( .A1(_GFM_n23980 ), .A2(_GFM_n2613 ), .ZN(_GFM_N802 ));
NOR2_X2 _GFM_U2210  ( .A1(_GFM_n23980 ), .A2(_GFM_n26140 ), .ZN(_GFM_N833 ));
NOR2_X2 _GFM_U2209  ( .A1(_GFM_n23980 ), .A2(_GFM_n26150 ), .ZN(_GFM_N864 ));
NOR2_X2 _GFM_U2208  ( .A1(_GFM_n23980 ), .A2(_GFM_n2616 ), .ZN(_GFM_N895 ));
NOR2_X2 _GFM_U2207  ( .A1(_GFM_n2387 ), .A2(_GFM_n2618 ), .ZN(_GFM_N927 ) );
NOR2_X2 _GFM_U2206  ( .A1(_GFM_n23980 ), .A2(_GFM_n2618 ), .ZN(_GFM_N957 ));
NOR2_X2 _GFM_U2205  ( .A1(_GFM_n24020 ), .A2(_GFM_n26190 ), .ZN(_GFM_N988 ));
NOR2_X2 _GFM_U2204  ( .A1(_GFM_n26200 ), .A2(_GFM_n23970 ), .ZN(_GFM_N1019 ));
NOR2_X2 _GFM_U2203  ( .A1(_GFM_n23980 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1050 ));
NOR2_X2 _GFM_U2202  ( .A1(_GFM_n2406 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1081 ));
NOR2_X2 _GFM_U2201  ( .A1(_GFM_n2406 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1112 ));
NOR2_X2 _GFM_U2200  ( .A1(_GFM_n2406 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1143 ));
NOR2_X2 _GFM_U2199  ( .A1(_GFM_n2406 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1174 ));
NOR2_X2 _GFM_U2198  ( .A1(_GFM_n2406 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1205 ));
NOR2_X2 _GFM_U2197  ( .A1(_GFM_n2406 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1236 ));
NOR2_X2 _GFM_U2196  ( .A1(_GFM_n2406 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1267 ));
NOR2_X2 _GFM_U2195  ( .A1(_GFM_n2406 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1298 ));
NOR2_X2 _GFM_U2194  ( .A1(_GFM_n2406 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1329 ));
NOR2_X2 _GFM_U2193  ( .A1(_GFM_n2406 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1360 ));
NOR2_X2 _GFM_U2192  ( .A1(_GFM_n24050 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1391 ));
NOR2_X2 _GFM_U2191  ( .A1(_GFM_n24050 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1422 ));
NOR2_X2 _GFM_U2190  ( .A1(_GFM_n24050 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1453 ));
NOR2_X2 _GFM_U2189  ( .A1(_GFM_n24050 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1484 ));
NOR2_X2 _GFM_U2188  ( .A1(_GFM_n24050 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1515 ));
NOR2_X2 _GFM_U2187  ( .A1(_GFM_n24050 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1546 ));
NOR2_X2 _GFM_U2186  ( .A1(_GFM_n24050 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1577 ));
NOR2_X2 _GFM_U2185  ( .A1(_GFM_n24050 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1608 ));
NOR2_X2 _GFM_U2184  ( .A1(_GFM_n24050 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1639 ));
NOR2_X2 _GFM_U2183  ( .A1(_GFM_n24050 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1670 ));
NOR2_X2 _GFM_U2182  ( .A1(_GFM_n24050 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1701 ));
NOR2_X2 _GFM_U2181  ( .A1(_GFM_n24050 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1732 ));
NOR2_X2 _GFM_U2180  ( .A1(_GFM_n2404 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1763 ));
NOR2_X2 _GFM_U2179  ( .A1(_GFM_n2404 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1794 ));
NOR2_X2 _GFM_U2178  ( .A1(_GFM_n2404 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1825 ));
NOR2_X2 _GFM_U2177  ( .A1(_GFM_n2404 ), .A2(_GFM_n2647 ), .ZN(_GFM_N1856 ));
NOR2_X2 _GFM_U2176  ( .A1(_GFM_n2404 ), .A2(_GFM_n2648 ), .ZN(_GFM_N1887 ));
NOR2_X2 _GFM_U2175  ( .A1(_GFM_n2404 ), .A2(_GFM_n2649 ), .ZN(_GFM_N1918 ));
NOR2_X2 _GFM_U2174  ( .A1(_GFM_n2404 ), .A2(_GFM_n26500 ), .ZN(_GFM_N1949 ));
NOR2_X2 _GFM_U2173  ( .A1(_GFM_n2404 ), .A2(_GFM_n26510 ), .ZN(_GFM_N1980 ));
NOR2_X2 _GFM_U2172  ( .A1(_GFM_n2404 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2011 ));
NOR2_X2 _GFM_U2171  ( .A1(_GFM_n2404 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2042 ));
NOR2_X2 _GFM_U2170  ( .A1(_GFM_n2404 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2073 ));
NOR2_X2 _GFM_U2169  ( .A1(_GFM_n2404 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2104 ));
NOR2_X2 _GFM_U2168  ( .A1(_GFM_n24030 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2135 ));
NOR2_X2 _GFM_U2167  ( .A1(_GFM_n24030 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2166 ));
NOR2_X2 _GFM_U2166  ( .A1(_GFM_n24030 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2197 ));
NOR2_X2 _GFM_U2165  ( .A1(_GFM_n24030 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2228 ));
NOR2_X2 _GFM_U2164  ( .A1(_GFM_n24030 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2259 ));
NOR2_X2 _GFM_U2163  ( .A1(_GFM_n24030 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2290 ));
NOR2_X2 _GFM_U2162  ( .A1(_GFM_n24030 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2321 ));
NOR2_X2 _GFM_U2161  ( .A1(_GFM_n24030 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2352 ));
NOR2_X2 _GFM_U2160  ( .A1(_GFM_n24030 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2383 ));
NOR2_X2 _GFM_U2159  ( .A1(_GFM_n24030 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2414 ));
NOR2_X2 _GFM_U2158  ( .A1(_GFM_n24030 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2445 ));
NOR2_X2 _GFM_U2157  ( .A1(_GFM_n24020 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2476 ));
NOR2_X2 _GFM_U2156  ( .A1(_GFM_n24020 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2507 ));
NOR2_X2 _GFM_U2155  ( .A1(_GFM_n24020 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2538 ));
NOR2_X2 _GFM_U2154  ( .A1(_GFM_n24020 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2569 ));
NOR2_X2 _GFM_U2153  ( .A1(_GFM_n24020 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2600 ));
NOR2_X2 _GFM_U2152  ( .A1(_GFM_n24020 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2631 ));
NOR2_X2 _GFM_U2151  ( .A1(_GFM_n24020 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2662 ));
NOR2_X2 _GFM_U2150  ( .A1(_GFM_n24020 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2693 ));
NOR2_X2 _GFM_U2149  ( .A1(_GFM_n24020 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2724 ));
NOR2_X2 _GFM_U2148  ( .A1(_GFM_n24020 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2755 ));
NOR2_X2 _GFM_U2147  ( .A1(_GFM_n24020 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2786 ));
NOR2_X2 _GFM_U2146  ( .A1(_GFM_n2401 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2817 ));
NOR2_X2 _GFM_U2145  ( .A1(_GFM_n2401 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2848 ));
NOR2_X2 _GFM_U2144  ( .A1(_GFM_n2401 ), .A2(_GFM_n26801 ), .ZN(_GFM_N2879 ));
NOR2_X2 _GFM_U2143  ( .A1(_GFM_n2401 ), .A2(_GFM_n26810 ), .ZN(_GFM_N2910 ));
NOR2_X2 _GFM_U2142  ( .A1(_GFM_n2401 ), .A2(_GFM_n26820 ), .ZN(_GFM_N2941 ));
NOR2_X2 _GFM_U2141  ( .A1(_GFM_n2401 ), .A2(_GFM_n2683 ), .ZN(_GFM_N2972 ));
NOR2_X2 _GFM_U2140  ( .A1(_GFM_n2401 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3003 ));
NOR2_X2 _GFM_U2139  ( .A1(_GFM_n2401 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3034 ));
NOR2_X2 _GFM_U2138  ( .A1(_GFM_n2401 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3065 ));
NOR2_X2 _GFM_U2137  ( .A1(_GFM_n2401 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3096 ));
NOR2_X2 _GFM_U2136  ( .A1(_GFM_n2401 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3127 ));
NOR2_X2 _GFM_U2135  ( .A1(_GFM_n2401 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3158 ));
NOR2_X2 _GFM_U2134  ( .A1(_GFM_n2400 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3189 ));
NOR2_X2 _GFM_U2133  ( .A1(_GFM_n2400 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3220 ));
NOR2_X2 _GFM_U2132  ( .A1(_GFM_n2400 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3251 ));
NOR2_X2 _GFM_U2131  ( .A1(_GFM_n2400 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3282 ));
NOR2_X2 _GFM_U2130  ( .A1(_GFM_n25180 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3747 ));
NOR2_X2 _GFM_U2129  ( .A1(_GFM_n25380 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3745 ));
NOR2_X2 _GFM_U2128  ( .A1(_GFM_n2547 ), .A2(_GFM_n25270 ), .ZN(_GFM_N3931 ));
NOR2_X2 _GFM_U2127  ( .A1(_GFM_n25380 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3928 ));
INV_X4 _GFM_U2126  ( .A(v_in[12]), .ZN(_GFM_n2586 ) );
INV_X4 _GFM_U2125  ( .A(v_in[14]), .ZN(_GFM_n25880 ) );
INV_X4 _GFM_U2124  ( .A(v_in[13]), .ZN(_GFM_n2587 ) );
INV_X4 _GFM_U2123  ( .A(b_in[123]), .ZN(_GFM_n24960 ) );
INV_X4 _GFM_U2122  ( .A(b_in[112]), .ZN(_GFM_n2387 ) );
INV_X4 _GFM_U2121  ( .A(b_in[114]), .ZN(_GFM_n24070 ) );
INV_X4 _GFM_U2120  ( .A(b_in[113]), .ZN(_GFM_n23970 ) );
INV_X4 _GFM_U2119  ( .A(b_in[117]), .ZN(_GFM_n24360 ) );
INV_X4 _GFM_U2118  ( .A(b_in[118]), .ZN(_GFM_n24460 ) );
INV_X4 _GFM_U2117  ( .A(b_in[120]), .ZN(_GFM_n2466 ) );
INV_X4 _GFM_U2116  ( .A(b_in[119]), .ZN(_GFM_n24560 ) );
INV_X4 _GFM_U2115  ( .A(b_in[122]), .ZN(_GFM_n2486 ) );
INV_X4 _GFM_U2114  ( .A(b_in[121]), .ZN(_GFM_n24760 ) );
INV_X4 _GFM_U2113  ( .A(b_in[124]), .ZN(_GFM_n2506 ) );
NOR2_X2 _GFM_U2112  ( .A1(_GFM_n25210 ), .A2(_GFM_n26080 ), .ZN(_GFM_N996 ));
NOR2_X2 _GFM_U2111  ( .A1(_GFM_n25180 ), .A2(_GFM_n26070 ), .ZN(_GFM_N965 ));
NOR2_X2 _GFM_U2110  ( .A1(_GFM_n2525 ), .A2(_GFM_n26200 ), .ZN(_GFM_N1368 ));
NOR2_X2 _GFM_U2109  ( .A1(_GFM_n2525 ), .A2(_GFM_n26190 ), .ZN(_GFM_N1337 ));
NOR2_X2 _GFM_U2108  ( .A1(_GFM_n2399 ), .A2(_GFM_n2617 ), .ZN(_GFM_N926 ) );
NOR2_X2 _GFM_U2107  ( .A1(_GFM_n24120 ), .A2(_GFM_n2618 ), .ZN(_GFM_N985 ));
NOR2_X2 _GFM_U2106  ( .A1(_GFM_n24080 ), .A2(_GFM_n26120 ), .ZN(_GFM_N799 ));
NOR2_X2 _GFM_U2105  ( .A1(_GFM_n2409 ), .A2(_GFM_n2613 ), .ZN(_GFM_N830 ) );
NOR2_X2 _GFM_U2104  ( .A1(_GFM_n24080 ), .A2(_GFM_n2616 ), .ZN(_GFM_N923 ));
NOR2_X2 _GFM_U2103  ( .A1(_GFM_n24650 ), .A2(_GFM_n2616 ), .ZN(_GFM_N1074 ));
NOR2_X2 _GFM_U2102  ( .A1(_GFM_n24080 ), .A2(_GFM_n26140 ), .ZN(_GFM_N861 ));
NOR2_X2 _GFM_U2101  ( .A1(_GFM_n24080 ), .A2(_GFM_n26150 ), .ZN(_GFM_N892 ));
NOR2_X2 _GFM_U2100  ( .A1(_GFM_n24650 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1043 ));
NOR2_X2 _GFM_U2099  ( .A1(_GFM_n24080 ), .A2(_GFM_n26110 ), .ZN(_GFM_N768 ));
NOR2_X2 _GFM_U2098  ( .A1(_GFM_n24570 ), .A2(_GFM_n26110 ), .ZN(_GFM_N919 ));
NOR2_X2 _GFM_U2097  ( .A1(_GFM_n2525 ), .A2(_GFM_n26110 ), .ZN(_GFM_N1089 ));
NOR2_X2 _GFM_U2096  ( .A1(_GFM_n2416 ), .A2(_GFM_n25901 ), .ZN(_GFM_N117 ));
NOR2_X2 _GFM_U2095  ( .A1(_GFM_n2461 ), .A2(_GFM_n25901 ), .ZN(_GFM_N268 ));
NOR2_X2 _GFM_U2094  ( .A1(_GFM_n24120 ), .A2(_GFM_n2595 ), .ZN(_GFM_N272 ));
NOR2_X2 _GFM_U2093  ( .A1(_GFM_n24110 ), .A2(_GFM_n2596 ), .ZN(_GFM_N303 ));
NOR2_X2 _GFM_U2092  ( .A1(_GFM_n24101 ), .A2(_GFM_n25970 ), .ZN(_GFM_N334 ));
NOR2_X2 _GFM_U2091  ( .A1(_GFM_n24101 ), .A2(_GFM_n25980 ), .ZN(_GFM_N365 ));
NOR2_X2 _GFM_U2090  ( .A1(_GFM_n2409 ), .A2(_GFM_n2599 ), .ZN(_GFM_N396 ) );
NOR2_X2 _GFM_U2089  ( .A1(_GFM_n2509 ), .A2(_GFM_n25901 ), .ZN(_GFM_N411 ));
NOR2_X2 _GFM_U2088  ( .A1(_GFM_n2409 ), .A2(_GFM_n26000 ), .ZN(_GFM_N427 ));
NOR2_X2 _GFM_U2087  ( .A1(_GFM_n25080 ), .A2(_GFM_n25910 ), .ZN(_GFM_N442 ));
NOR2_X2 _GFM_U2086  ( .A1(_GFM_n2409 ), .A2(_GFM_n26010 ), .ZN(_GFM_N458 ));
NOR2_X2 _GFM_U2085  ( .A1(_GFM_n2509 ), .A2(_GFM_n2592 ), .ZN(_GFM_N473 ) );
NOR2_X2 _GFM_U2084  ( .A1(_GFM_n24080 ), .A2(_GFM_n2602 ), .ZN(_GFM_N489 ));
NOR2_X2 _GFM_U2083  ( .A1(_GFM_n2509 ), .A2(_GFM_n25930 ), .ZN(_GFM_N504 ));
NOR2_X2 _GFM_U2082  ( .A1(_GFM_n2409 ), .A2(_GFM_n2603 ), .ZN(_GFM_N520 ) );
NOR2_X2 _GFM_U2081  ( .A1(_GFM_n2509 ), .A2(_GFM_n25940 ), .ZN(_GFM_N535 ));
NOR2_X2 _GFM_U2080  ( .A1(_GFM_n24080 ), .A2(_GFM_n2604 ), .ZN(_GFM_N551 ));
NOR2_X2 _GFM_U2079  ( .A1(_GFM_n2399 ), .A2(_GFM_n26050 ), .ZN(_GFM_N554 ));
NOR2_X2 _GFM_U2078  ( .A1(_GFM_n25080 ), .A2(_GFM_n2595 ), .ZN(_GFM_N566 ));
NOR2_X2 _GFM_U2077  ( .A1(_GFM_n24080 ), .A2(_GFM_n26050 ), .ZN(_GFM_N582 ));
NOR2_X2 _GFM_U2076  ( .A1(_GFM_n2509 ), .A2(_GFM_n2596 ), .ZN(_GFM_N597 ) );
NOR2_X2 _GFM_U2075  ( .A1(_GFM_n25080 ), .A2(_GFM_n25970 ), .ZN(_GFM_N628 ));
NOR2_X2 _GFM_U2074  ( .A1(_GFM_n24570 ), .A2(_GFM_n2602 ), .ZN(_GFM_N640 ));
NOR2_X2 _GFM_U2073  ( .A1(_GFM_n25080 ), .A2(_GFM_n25980 ), .ZN(_GFM_N659 ));
NOR2_X2 _GFM_U2072  ( .A1(_GFM_n2458 ), .A2(_GFM_n2603 ), .ZN(_GFM_N671 ) );
NOR2_X2 _GFM_U2071  ( .A1(_GFM_n23980 ), .A2(_GFM_n2609 ), .ZN(_GFM_N678 ));
NOR2_X2 _GFM_U2070  ( .A1(_GFM_n25080 ), .A2(_GFM_n2599 ), .ZN(_GFM_N690 ));
NOR2_X2 _GFM_U2069  ( .A1(_GFM_n24080 ), .A2(_GFM_n2609 ), .ZN(_GFM_N706 ));
NOR2_X2 _GFM_U2068  ( .A1(_GFM_n24570 ), .A2(_GFM_n2604 ), .ZN(_GFM_N702 ));
NOR2_X2 _GFM_U2067  ( .A1(_GFM_n25080 ), .A2(_GFM_n26000 ), .ZN(_GFM_N721 ));
NOR2_X2 _GFM_U2066  ( .A1(_GFM_n2517 ), .A2(_GFM_n26000 ), .ZN(_GFM_N748 ));
NOR2_X2 _GFM_U2065  ( .A1(_GFM_n25080 ), .A2(_GFM_n2602 ), .ZN(_GFM_N783 ));
NOR2_X2 _GFM_U2064  ( .A1(_GFM_n25180 ), .A2(_GFM_n2602 ), .ZN(_GFM_N810 ));
NOR2_X2 _GFM_U2063  ( .A1(_GFM_n24570 ), .A2(_GFM_n2609 ), .ZN(_GFM_N857 ));
NOR2_X2 _GFM_U2062  ( .A1(_GFM_n25080 ), .A2(_GFM_n26050 ), .ZN(_GFM_N876 ));
NOR2_X2 _GFM_U2061  ( .A1(_GFM_n24770 ), .A2(_GFM_n2609 ), .ZN(_GFM_N910 ));
NOR2_X2 _GFM_U2060  ( .A1(_GFM_n2511 ), .A2(_GFM_n2609 ), .ZN(_GFM_N1000 ));
NOR2_X2 _GFM_U2059  ( .A1(_GFM_n2517 ), .A2(_GFM_n2609 ), .ZN(_GFM_N1027 ));
NOR2_X2 _GFM_U2058  ( .A1(_GFM_n24080 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1078 ));
NOR2_X2 _GFM_U2057  ( .A1(_GFM_n2416 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1109 ));
NOR2_X2 _GFM_U2056  ( .A1(_GFM_n2416 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1140 ));
NOR2_X2 _GFM_U2055  ( .A1(_GFM_n2416 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1171 ));
NOR2_X2 _GFM_U2054  ( .A1(_GFM_n2455 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1194 ));
NOR2_X2 _GFM_U2053  ( .A1(_GFM_n2416 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1202 ));
NOR2_X2 _GFM_U2052  ( .A1(_GFM_n2455 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1225 ));
NOR2_X2 _GFM_U2051  ( .A1(_GFM_n24650 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1229 ));
NOR2_X2 _GFM_U2050  ( .A1(_GFM_n2416 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1233 ));
NOR2_X2 _GFM_U2049  ( .A1(_GFM_n2455 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1256 ));
NOR2_X2 _GFM_U2048  ( .A1(_GFM_n2416 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1264 ));
NOR2_X2 _GFM_U2047  ( .A1(_GFM_n2455 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1287 ));
NOR2_X2 _GFM_U2046  ( .A1(_GFM_n2416 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1295 ));
NOR2_X2 _GFM_U2045  ( .A1(_GFM_n2416 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1326 ));
NOR2_X2 _GFM_U2044  ( .A1(_GFM_n2416 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1357 ));
NOR2_X2 _GFM_U2043  ( .A1(_GFM_n2416 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1388 ));
NOR2_X2 _GFM_U2042  ( .A1(_GFM_n2524 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1399 ));
NOR2_X2 _GFM_U2041  ( .A1(_GFM_n24150 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1419 ));
NOR2_X2 _GFM_U2040  ( .A1(_GFM_n2524 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1430 ));
NOR2_X2 _GFM_U2039  ( .A1(_GFM_n24150 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1450 ));
NOR2_X2 _GFM_U2038  ( .A1(_GFM_n2524 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1461 ));
NOR2_X2 _GFM_U2037  ( .A1(_GFM_n24150 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1481 ));
NOR2_X2 _GFM_U2036  ( .A1(_GFM_n2524 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1492 ));
NOR2_X2 _GFM_U2035  ( .A1(_GFM_n24150 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1512 ));
NOR2_X2 _GFM_U2034  ( .A1(_GFM_n2524 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1523 ));
NOR2_X2 _GFM_U2033  ( .A1(_GFM_n24150 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1543 ));
NOR2_X2 _GFM_U2032  ( .A1(_GFM_n2524 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1554 ));
NOR2_X2 _GFM_U2031  ( .A1(_GFM_n24150 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1574 ));
NOR2_X2 _GFM_U2030  ( .A1(_GFM_n2524 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1585 ));
NOR2_X2 _GFM_U2029  ( .A1(_GFM_n24150 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1605 ));
NOR2_X2 _GFM_U2028  ( .A1(_GFM_n25150 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1620 ));
NOR2_X2 _GFM_U2027  ( .A1(_GFM_n24150 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1636 ));
NOR2_X2 _GFM_U2026  ( .A1(_GFM_n25150 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1651 ));
NOR2_X2 _GFM_U2025  ( .A1(_GFM_n24150 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1667 ));
NOR2_X2 _GFM_U2024  ( .A1(_GFM_n25140 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1682 ));
NOR2_X2 _GFM_U2023  ( .A1(_GFM_n24150 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1698 ));
NOR2_X2 _GFM_U2022  ( .A1(_GFM_n25140 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1713 ));
NOR2_X2 _GFM_U2021  ( .A1(_GFM_n24150 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1729 ));
NOR2_X2 _GFM_U2020  ( .A1(_GFM_n25140 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1744 ));
NOR2_X2 _GFM_U2019  ( .A1(_GFM_n24150 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1760 ));
NOR2_X2 _GFM_U2018  ( .A1(_GFM_n25140 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1775 ));
NOR2_X2 _GFM_U2017  ( .A1(_GFM_n24140 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1791 ));
NOR2_X2 _GFM_U2016  ( .A1(_GFM_n25140 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1806 ));
NOR2_X2 _GFM_U2015  ( .A1(_GFM_n24140 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1822 ));
NOR2_X2 _GFM_U2014  ( .A1(_GFM_n25140 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1837 ));
NOR2_X2 _GFM_U2013  ( .A1(_GFM_n24140 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1853 ));
NOR2_X2 _GFM_U2012  ( .A1(_GFM_n25140 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1868 ));
NOR2_X2 _GFM_U2011  ( .A1(_GFM_n24140 ), .A2(_GFM_n2647 ), .ZN(_GFM_N1884 ));
NOR2_X2 _GFM_U2010  ( .A1(_GFM_n25140 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1899 ));
NOR2_X2 _GFM_U2009  ( .A1(_GFM_n24140 ), .A2(_GFM_n2648 ), .ZN(_GFM_N1915 ));
NOR2_X2 _GFM_U2008  ( .A1(_GFM_n25140 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1930 ));
NOR2_X2 _GFM_U2007  ( .A1(_GFM_n24140 ), .A2(_GFM_n2649 ), .ZN(_GFM_N1946 ));
NOR2_X2 _GFM_U2006  ( .A1(_GFM_n25140 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1961 ));
NOR2_X2 _GFM_U2005  ( .A1(_GFM_n24140 ), .A2(_GFM_n26500 ), .ZN(_GFM_N1977 ));
NOR2_X2 _GFM_U2004  ( .A1(_GFM_n25140 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1992 ));
NOR2_X2 _GFM_U2003  ( .A1(_GFM_n24140 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2008 ));
NOR2_X2 _GFM_U2002  ( .A1(_GFM_n25140 ), .A2(_GFM_n26420 ), .ZN(_GFM_N2023 ));
NOR2_X2 _GFM_U2001  ( .A1(_GFM_n24140 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2039 ));
NOR2_X2 _GFM_U2000  ( .A1(_GFM_n2513 ), .A2(_GFM_n26430 ), .ZN(_GFM_N2054 ));
NOR2_X2 _GFM_U1999  ( .A1(_GFM_n24140 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2070 ));
NOR2_X2 _GFM_U1998  ( .A1(_GFM_n2513 ), .A2(_GFM_n2644 ), .ZN(_GFM_N2085 ));
NOR2_X2 _GFM_U1997  ( .A1(_GFM_n24140 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2101 ));
NOR2_X2 _GFM_U1996  ( .A1(_GFM_n2513 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2116 ));
NOR2_X2 _GFM_U1995  ( .A1(_GFM_n2413 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2132 ));
NOR2_X2 _GFM_U1994  ( .A1(_GFM_n2513 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2147 ));
NOR2_X2 _GFM_U1993  ( .A1(_GFM_n2413 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2163 ));
NOR2_X2 _GFM_U1992  ( .A1(_GFM_n2513 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2178 ));
NOR2_X2 _GFM_U1991  ( .A1(_GFM_n2413 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2194 ));
NOR2_X2 _GFM_U1990  ( .A1(_GFM_n2513 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2209 ));
NOR2_X2 _GFM_U1989  ( .A1(_GFM_n2413 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2225 ));
NOR2_X2 _GFM_U1988  ( .A1(_GFM_n2513 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2240 ));
NOR2_X2 _GFM_U1987  ( .A1(_GFM_n2413 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2256 ));
NOR2_X2 _GFM_U1986  ( .A1(_GFM_n2513 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2271 ));
NOR2_X2 _GFM_U1985  ( .A1(_GFM_n2413 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2287 ));
NOR2_X2 _GFM_U1984  ( .A1(_GFM_n2513 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2302 ));
NOR2_X2 _GFM_U1983  ( .A1(_GFM_n2413 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2318 ));
NOR2_X2 _GFM_U1982  ( .A1(_GFM_n2513 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2333 ));
NOR2_X2 _GFM_U1981  ( .A1(_GFM_n2413 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2349 ));
NOR2_X2 _GFM_U1980  ( .A1(_GFM_n2513 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2364 ));
NOR2_X2 _GFM_U1979  ( .A1(_GFM_n2413 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2380 ));
NOR2_X2 _GFM_U1978  ( .A1(_GFM_n2513 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2395 ));
NOR2_X2 _GFM_U1977  ( .A1(_GFM_n2413 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2411 ));
NOR2_X2 _GFM_U1976  ( .A1(_GFM_n25120 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2426 ));
NOR2_X2 _GFM_U1975  ( .A1(_GFM_n2413 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2442 ));
NOR2_X2 _GFM_U1974  ( .A1(_GFM_n25120 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2457 ));
NOR2_X2 _GFM_U1973  ( .A1(_GFM_n24120 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2473 ));
NOR2_X2 _GFM_U1972  ( .A1(_GFM_n25120 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2488 ));
NOR2_X2 _GFM_U1971  ( .A1(_GFM_n24120 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2504 ));
NOR2_X2 _GFM_U1970  ( .A1(_GFM_n25120 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2519 ));
NOR2_X2 _GFM_U1969  ( .A1(_GFM_n24120 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2535 ));
NOR2_X2 _GFM_U1968  ( .A1(_GFM_n25120 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2550 ));
NOR2_X2 _GFM_U1967  ( .A1(_GFM_n24120 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2566 ));
NOR2_X2 _GFM_U1966  ( .A1(_GFM_n25120 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2581 ));
NOR2_X2 _GFM_U1965  ( .A1(_GFM_n24120 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2597 ));
NOR2_X2 _GFM_U1964  ( .A1(_GFM_n25120 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2612 ));
NOR2_X2 _GFM_U1963  ( .A1(_GFM_n24120 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2628 ));
NOR2_X2 _GFM_U1962  ( .A1(_GFM_n25120 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2643 ));
NOR2_X2 _GFM_U1961  ( .A1(_GFM_n25120 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2674 ));
NOR2_X2 _GFM_U1960  ( .A1(_GFM_n25120 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2705 ));
NOR2_X2 _GFM_U1959  ( .A1(_GFM_n25120 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2736 ));
NOR2_X2 _GFM_U1958  ( .A1(_GFM_n25120 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2767 ));
NOR2_X2 _GFM_U1957  ( .A1(_GFM_n2511 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2798 ));
NOR2_X2 _GFM_U1956  ( .A1(_GFM_n2511 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2829 ));
NOR2_X2 _GFM_U1955  ( .A1(_GFM_n2511 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2860 ));
NOR2_X2 _GFM_U1954  ( .A1(_GFM_n2511 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2891 ));
NOR2_X2 _GFM_U1953  ( .A1(_GFM_n2511 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2922 ));
NOR2_X2 _GFM_U1952  ( .A1(_GFM_n24120 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2659 ));
NOR2_X2 _GFM_U1951  ( .A1(_GFM_n24120 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2690 ));
NOR2_X2 _GFM_U1950  ( .A1(_GFM_n24120 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2721 ));
NOR2_X2 _GFM_U1949  ( .A1(_GFM_n24120 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2752 ));
NOR2_X2 _GFM_U1948  ( .A1(_GFM_n24120 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2783 ));
NOR2_X2 _GFM_U1947  ( .A1(_GFM_n24110 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2814 ));
NOR2_X2 _GFM_U1946  ( .A1(_GFM_n24110 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2845 ));
NOR2_X2 _GFM_U1945  ( .A1(_GFM_n24110 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2876 ));
NOR2_X2 _GFM_U1944  ( .A1(_GFM_n24110 ), .A2(_GFM_n26801 ), .ZN(_GFM_N2907 ));
NOR2_X2 _GFM_U1943  ( .A1(_GFM_n24110 ), .A2(_GFM_n26810 ), .ZN(_GFM_N2938 ));
NOR2_X2 _GFM_U1942  ( .A1(_GFM_n2511 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2953 ));
NOR2_X2 _GFM_U1941  ( .A1(_GFM_n24110 ), .A2(_GFM_n26820 ), .ZN(_GFM_N2969 ));
NOR2_X2 _GFM_U1940  ( .A1(_GFM_n2511 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2984 ));
NOR2_X2 _GFM_U1939  ( .A1(_GFM_n24110 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3000 ));
NOR2_X2 _GFM_U1938  ( .A1(_GFM_n2511 ), .A2(_GFM_n26740 ), .ZN(_GFM_N3015 ));
NOR2_X2 _GFM_U1937  ( .A1(_GFM_n24110 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3031 ));
NOR2_X2 _GFM_U1936  ( .A1(_GFM_n2511 ), .A2(_GFM_n2675 ), .ZN(_GFM_N3046 ));
NOR2_X2 _GFM_U1935  ( .A1(_GFM_n24110 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3062 ));
NOR2_X2 _GFM_U1934  ( .A1(_GFM_n2511 ), .A2(_GFM_n26760 ), .ZN(_GFM_N3077 ));
NOR2_X2 _GFM_U1933  ( .A1(_GFM_n24110 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3093 ));
NOR2_X2 _GFM_U1932  ( .A1(_GFM_n2511 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3108 ));
NOR2_X2 _GFM_U1931  ( .A1(_GFM_n24110 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3124 ));
NOR2_X2 _GFM_U1930  ( .A1(_GFM_n25101 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3139 ));
NOR2_X2 _GFM_U1929  ( .A1(_GFM_n24110 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3155 ));
NOR2_X2 _GFM_U1928  ( .A1(_GFM_n25101 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3170 ));
NOR2_X2 _GFM_U1927  ( .A1(_GFM_n24101 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3186 ));
NOR2_X2 _GFM_U1926  ( .A1(_GFM_n25101 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3201 ));
NOR2_X2 _GFM_U1925  ( .A1(_GFM_n24101 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3217 ));
NOR2_X2 _GFM_U1924  ( .A1(_GFM_n25101 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3232 ));
NOR2_X2 _GFM_U1923  ( .A1(_GFM_n24101 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3248 ));
NOR2_X2 _GFM_U1922  ( .A1(_GFM_n25101 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3263 ));
NOR2_X2 _GFM_U1921  ( .A1(_GFM_n24101 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3279 ));
NOR2_X2 _GFM_U1920  ( .A1(_GFM_n24900 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3294 ));
NOR2_X2 _GFM_U1919  ( .A1(_GFM_n24590 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3309 ));
NOR2_X2 _GFM_U1918  ( .A1(_GFM_n24101 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3313 ));
NOR2_X2 _GFM_U1917  ( .A1(_GFM_n24900 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3326 ));
NOR2_X2 _GFM_U1916  ( .A1(_GFM_n24101 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3346 ));
NOR2_X2 _GFM_U1915  ( .A1(_GFM_n24590 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3341 ));
NOR2_X2 _GFM_U1914  ( .A1(_GFM_n24900 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3359 ));
NOR2_X2 _GFM_U1913  ( .A1(_GFM_n24590 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3374 ));
NOR2_X2 _GFM_U1912  ( .A1(_GFM_n24900 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3393 ));
NOR2_X2 _GFM_U1911  ( .A1(_GFM_n24290 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3402 ));
NOR2_X2 _GFM_U1910  ( .A1(_GFM_n24900 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3429 ));
NOR2_X2 _GFM_U1909  ( .A1(_GFM_n24590 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3514 ));
NOR2_X2 _GFM_U1908  ( .A1(_GFM_n25000 ), .A2(_GFM_n2610 ), .ZN(_GFM_N999 ));
NOR2_X2 _GFM_U1907  ( .A1(_GFM_n2497 ), .A2(_GFM_n26080 ), .ZN(_GFM_N937 ));
NOR2_X2 _GFM_U1906  ( .A1(_GFM_n2497 ), .A2(_GFM_n2606 ), .ZN(_GFM_N875 ) );
NOR2_X2 _GFM_U1905  ( .A1(_GFM_n25050 ), .A2(_GFM_n26200 ), .ZN(_GFM_N1309 ));
NOR2_X2 _GFM_U1904  ( .A1(_GFM_n25050 ), .A2(_GFM_n26190 ), .ZN(_GFM_N1278 ));
NOR2_X2 _GFM_U1903  ( .A1(_GFM_n2525 ), .A2(_GFM_n2617 ), .ZN(_GFM_N1275 ));
NOR2_X2 _GFM_U1902  ( .A1(_GFM_n25050 ), .A2(_GFM_n2617 ), .ZN(_GFM_N1216 ));
NOR2_X2 _GFM_U1901  ( .A1(_GFM_n2525 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1213 ));
NOR2_X2 _GFM_U1900  ( .A1(_GFM_n24210 ), .A2(_GFM_n2617 ), .ZN(_GFM_N986 ));
NOR2_X2 _GFM_U1899  ( .A1(_GFM_n2417 ), .A2(_GFM_n2618 ), .ZN(_GFM_N1017 ));
NOR2_X2 _GFM_U1898  ( .A1(_GFM_n2417 ), .A2(_GFM_n26120 ), .ZN(_GFM_N831 ));
NOR2_X2 _GFM_U1897  ( .A1(_GFM_n2471 ), .A2(_GFM_n26120 ), .ZN(_GFM_N982 ));
NOR2_X2 _GFM_U1896  ( .A1(_GFM_n25050 ), .A2(_GFM_n26120 ), .ZN(_GFM_N1061 ));
NOR2_X2 _GFM_U1895  ( .A1(_GFM_n2417 ), .A2(_GFM_n2613 ), .ZN(_GFM_N862 ) );
NOR2_X2 _GFM_U1894  ( .A1(_GFM_n24670 ), .A2(_GFM_n2613 ), .ZN(_GFM_N1013 ));
NOR2_X2 _GFM_U1893  ( .A1(_GFM_n25050 ), .A2(_GFM_n2613 ), .ZN(_GFM_N1092 ));
NOR2_X2 _GFM_U1892  ( .A1(_GFM_n2431 ), .A2(_GFM_n2616 ), .ZN(_GFM_N979 ) );
NOR2_X2 _GFM_U1891  ( .A1(_GFM_n24511 ), .A2(_GFM_n26140 ), .ZN(_GFM_N977 ));
NOR2_X2 _GFM_U1890  ( .A1(_GFM_n25050 ), .A2(_GFM_n2616 ), .ZN(_GFM_N1185 ));
NOR2_X2 _GFM_U1889  ( .A1(_GFM_n2525 ), .A2(_GFM_n26140 ), .ZN(_GFM_N1182 ));
NOR2_X2 _GFM_U1888  ( .A1(_GFM_n2417 ), .A2(_GFM_n2616 ), .ZN(_GFM_N955 ) );
NOR2_X2 _GFM_U1887  ( .A1(_GFM_n2475 ), .A2(_GFM_n2616 ), .ZN(_GFM_N1106 ));
NOR2_X2 _GFM_U1886  ( .A1(_GFM_n25050 ), .A2(_GFM_n26140 ), .ZN(_GFM_N1123 ));
NOR2_X2 _GFM_U1885  ( .A1(_GFM_n2525 ), .A2(_GFM_n26120 ), .ZN(_GFM_N1120 ));
NOR2_X2 _GFM_U1884  ( .A1(_GFM_n2417 ), .A2(_GFM_n26140 ), .ZN(_GFM_N893 ));
NOR2_X2 _GFM_U1883  ( .A1(_GFM_n2427 ), .A2(_GFM_n26140 ), .ZN(_GFM_N917 ));
NOR2_X2 _GFM_U1882  ( .A1(_GFM_n2475 ), .A2(_GFM_n26140 ), .ZN(_GFM_N1044 ));
NOR2_X2 _GFM_U1881  ( .A1(_GFM_n26980 ), .A2(_GFM_n25070 ), .ZN(_GFM_N4052 ));
NOR2_X2 _GFM_U1880  ( .A1(_GFM_n2427 ), .A2(_GFM_n26150 ), .ZN(_GFM_N948 ));
NOR2_X2 _GFM_U1879  ( .A1(_GFM_n2613 ), .A2(_GFM_n24460 ), .ZN(_GFM_N946 ));
NOR2_X2 _GFM_U1878  ( .A1(_GFM_n25050 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1154 ));
NOR2_X2 _GFM_U1877  ( .A1(_GFM_n2525 ), .A2(_GFM_n2613 ), .ZN(_GFM_N1151 ));
NOR2_X2 _GFM_U1876  ( .A1(_GFM_n2417 ), .A2(_GFM_n26150 ), .ZN(_GFM_N924 ));
NOR2_X2 _GFM_U1875  ( .A1(_GFM_n2475 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1075 ));
NOR2_X2 _GFM_U1874  ( .A1(_GFM_n2417 ), .A2(_GFM_n26110 ), .ZN(_GFM_N800 ));
NOR2_X2 _GFM_U1873  ( .A1(_GFM_n2437 ), .A2(_GFM_n26110 ), .ZN(_GFM_N852 ));
NOR2_X2 _GFM_U1872  ( .A1(_GFM_n24670 ), .A2(_GFM_n26110 ), .ZN(_GFM_N951 ));
NOR2_X2 _GFM_U1871  ( .A1(_GFM_n25050 ), .A2(_GFM_n26110 ), .ZN(_GFM_N1030 ));
NOR2_X2 _GFM_U1870  ( .A1(_GFM_n24330 ), .A2(_GFM_n25910 ), .ZN(_GFM_N204 ));
NOR2_X2 _GFM_U1869  ( .A1(_GFM_n25890 ), .A2(_GFM_n2447 ), .ZN(_GFM_N202 ));
NOR2_X2 _GFM_U1868  ( .A1(_GFM_n2427 ), .A2(_GFM_n2604 ), .ZN(_GFM_N607 ) );
NOR2_X2 _GFM_U1867  ( .A1(_GFM_n2448 ), .A2(_GFM_n2602 ), .ZN(_GFM_N605 ) );
NOR2_X2 _GFM_U1866  ( .A1(_GFM_n2427 ), .A2(_GFM_n26050 ), .ZN(_GFM_N638 ));
NOR2_X2 _GFM_U1865  ( .A1(_GFM_n2447 ), .A2(_GFM_n2603 ), .ZN(_GFM_N636 ) );
NOR2_X2 _GFM_U1864  ( .A1(_GFM_n2435 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1320 ));
NOR2_X2 _GFM_U1863  ( .A1(_GFM_n2455 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1318 ));
NOR2_X2 _GFM_U1862  ( .A1(_GFM_n2435 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1351 ));
NOR2_X2 _GFM_U1861  ( .A1(_GFM_n2455 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1349 ));
NOR2_X2 _GFM_U1860  ( .A1(_GFM_n2435 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1382 ));
NOR2_X2 _GFM_U1859  ( .A1(_GFM_n2455 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1380 ));
NOR2_X2 _GFM_U1858  ( .A1(_GFM_n2435 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1413 ));
NOR2_X2 _GFM_U1857  ( .A1(_GFM_n2455 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1411 ));
NOR2_X2 _GFM_U1856  ( .A1(_GFM_n2435 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1444 ));
NOR2_X2 _GFM_U1855  ( .A1(_GFM_n2455 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1442 ));
NOR2_X2 _GFM_U1854  ( .A1(_GFM_n2435 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1475 ));
NOR2_X2 _GFM_U1853  ( .A1(_GFM_n2455 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1473 ));
NOR2_X2 _GFM_U1852  ( .A1(_GFM_n2435 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1506 ));
NOR2_X2 _GFM_U1851  ( .A1(_GFM_n2454 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1504 ));
NOR2_X2 _GFM_U1850  ( .A1(_GFM_n24330 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2002 ));
NOR2_X2 _GFM_U1849  ( .A1(_GFM_n24530 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2000 ));
NOR2_X2 _GFM_U1848  ( .A1(_GFM_n24330 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2033 ));
NOR2_X2 _GFM_U1847  ( .A1(_GFM_n24530 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2031 ));
NOR2_X2 _GFM_U1846  ( .A1(_GFM_n24330 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2064 ));
NOR2_X2 _GFM_U1845  ( .A1(_GFM_n24530 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2062 ));
NOR2_X2 _GFM_U1844  ( .A1(_GFM_n2396 ), .A2(_GFM_n2592 ), .ZN(_GFM_N121 ) );
NOR2_X2 _GFM_U1843  ( .A1(_GFM_n2424 ), .A2(_GFM_n25901 ), .ZN(_GFM_N149 ));
NOR2_X2 _GFM_U1842  ( .A1(_GFM_n2423 ), .A2(_GFM_n25910 ), .ZN(_GFM_N180 ));
NOR2_X2 _GFM_U1841  ( .A1(_GFM_n2423 ), .A2(_GFM_n2592 ), .ZN(_GFM_N211 ) );
NOR2_X2 _GFM_U1840  ( .A1(_GFM_n24220 ), .A2(_GFM_n25930 ), .ZN(_GFM_N242 ));
NOR2_X2 _GFM_U1839  ( .A1(_GFM_n24210 ), .A2(_GFM_n25940 ), .ZN(_GFM_N273 ));
NOR2_X2 _GFM_U1838  ( .A1(_GFM_n23910 ), .A2(_GFM_n25970 ), .ZN(_GFM_N276 ));
NOR2_X2 _GFM_U1837  ( .A1(_GFM_n24700 ), .A2(_GFM_n25901 ), .ZN(_GFM_N300 ));
NOR2_X2 _GFM_U1836  ( .A1(_GFM_n24201 ), .A2(_GFM_n2595 ), .ZN(_GFM_N304 ));
NOR2_X2 _GFM_U1835  ( .A1(_GFM_n23910 ), .A2(_GFM_n25980 ), .ZN(_GFM_N307 ));
NOR2_X2 _GFM_U1834  ( .A1(_GFM_n24690 ), .A2(_GFM_n25910 ), .ZN(_GFM_N331 ));
NOR2_X2 _GFM_U1833  ( .A1(_GFM_n24190 ), .A2(_GFM_n2596 ), .ZN(_GFM_N335 ));
NOR2_X2 _GFM_U1832  ( .A1(_GFM_n23900 ), .A2(_GFM_n2599 ), .ZN(_GFM_N338 ));
NOR2_X2 _GFM_U1831  ( .A1(_GFM_n2489 ), .A2(_GFM_n25901 ), .ZN(_GFM_N351 ));
NOR2_X2 _GFM_U1830  ( .A1(_GFM_n24690 ), .A2(_GFM_n2592 ), .ZN(_GFM_N362 ));
NOR2_X2 _GFM_U1829  ( .A1(_GFM_n24190 ), .A2(_GFM_n25970 ), .ZN(_GFM_N366 ));
NOR2_X2 _GFM_U1828  ( .A1(_GFM_n23900 ), .A2(_GFM_n26000 ), .ZN(_GFM_N369 ));
NOR2_X2 _GFM_U1827  ( .A1(_GFM_n24980 ), .A2(_GFM_n25901 ), .ZN(_GFM_N379 ));
NOR2_X2 _GFM_U1826  ( .A1(_GFM_n24910 ), .A2(_GFM_n25910 ), .ZN(_GFM_N382 ));
NOR2_X2 _GFM_U1825  ( .A1(_GFM_n2468 ), .A2(_GFM_n25930 ), .ZN(_GFM_N393 ));
NOR2_X2 _GFM_U1824  ( .A1(_GFM_n2418 ), .A2(_GFM_n25980 ), .ZN(_GFM_N397 ));
NOR2_X2 _GFM_U1823  ( .A1(_GFM_n2389 ), .A2(_GFM_n26010 ), .ZN(_GFM_N400 ));
NOR2_X2 _GFM_U1822  ( .A1(_GFM_n24980 ), .A2(_GFM_n25910 ), .ZN(_GFM_N410 ));
NOR2_X2 _GFM_U1821  ( .A1(_GFM_n2489 ), .A2(_GFM_n2592 ), .ZN(_GFM_N413 ) );
NOR2_X2 _GFM_U1820  ( .A1(_GFM_n24690 ), .A2(_GFM_n25940 ), .ZN(_GFM_N424 ));
NOR2_X2 _GFM_U1819  ( .A1(_GFM_n2418 ), .A2(_GFM_n2599 ), .ZN(_GFM_N428 ) );
NOR2_X2 _GFM_U1818  ( .A1(_GFM_n2389 ), .A2(_GFM_n2602 ), .ZN(_GFM_N431 ) );
NOR2_X2 _GFM_U1817  ( .A1(_GFM_n24980 ), .A2(_GFM_n2592 ), .ZN(_GFM_N441 ));
NOR2_X2 _GFM_U1816  ( .A1(_GFM_n2489 ), .A2(_GFM_n25930 ), .ZN(_GFM_N444 ));
NOR2_X2 _GFM_U1815  ( .A1(_GFM_n2468 ), .A2(_GFM_n2595 ), .ZN(_GFM_N455 ) );
NOR2_X2 _GFM_U1814  ( .A1(_GFM_n2418 ), .A2(_GFM_n26000 ), .ZN(_GFM_N459 ));
NOR2_X2 _GFM_U1813  ( .A1(_GFM_n23880 ), .A2(_GFM_n2603 ), .ZN(_GFM_N462 ));
NOR2_X2 _GFM_U1812  ( .A1(_GFM_n2497 ), .A2(_GFM_n25930 ), .ZN(_GFM_N472 ));
NOR2_X2 _GFM_U1811  ( .A1(_GFM_n24880 ), .A2(_GFM_n25940 ), .ZN(_GFM_N475 ));
NOR2_X2 _GFM_U1810  ( .A1(_GFM_n2468 ), .A2(_GFM_n2596 ), .ZN(_GFM_N486 ) );
NOR2_X2 _GFM_U1809  ( .A1(_GFM_n2417 ), .A2(_GFM_n26010 ), .ZN(_GFM_N490 ));
NOR2_X2 _GFM_U1808  ( .A1(_GFM_n23880 ), .A2(_GFM_n2604 ), .ZN(_GFM_N493 ));
NOR2_X2 _GFM_U1807  ( .A1(_GFM_n24980 ), .A2(_GFM_n25940 ), .ZN(_GFM_N503 ));
NOR2_X2 _GFM_U1806  ( .A1(_GFM_n24880 ), .A2(_GFM_n2595 ), .ZN(_GFM_N506 ));
NOR2_X2 _GFM_U1805  ( .A1(_GFM_n2468 ), .A2(_GFM_n25970 ), .ZN(_GFM_N517 ));
NOR2_X2 _GFM_U1804  ( .A1(_GFM_n2418 ), .A2(_GFM_n2602 ), .ZN(_GFM_N521 ) );
NOR2_X2 _GFM_U1803  ( .A1(_GFM_n24980 ), .A2(_GFM_n2595 ), .ZN(_GFM_N534 ));
NOR2_X2 _GFM_U1802  ( .A1(_GFM_n24880 ), .A2(_GFM_n2596 ), .ZN(_GFM_N537 ));
NOR2_X2 _GFM_U1801  ( .A1(_GFM_n2468 ), .A2(_GFM_n25980 ), .ZN(_GFM_N548 ));
NOR2_X2 _GFM_U1800  ( .A1(_GFM_n2418 ), .A2(_GFM_n2603 ), .ZN(_GFM_N552 ) );
NOR2_X2 _GFM_U1799  ( .A1(_GFM_n2497 ), .A2(_GFM_n2596 ), .ZN(_GFM_N565 ) );
NOR2_X2 _GFM_U1798  ( .A1(_GFM_n24880 ), .A2(_GFM_n25970 ), .ZN(_GFM_N568 ));
NOR2_X2 _GFM_U1797  ( .A1(_GFM_n24670 ), .A2(_GFM_n2599 ), .ZN(_GFM_N579 ));
NOR2_X2 _GFM_U1796  ( .A1(_GFM_n2417 ), .A2(_GFM_n2604 ), .ZN(_GFM_N583 ) );
NOR2_X2 _GFM_U1795  ( .A1(_GFM_n2497 ), .A2(_GFM_n25970 ), .ZN(_GFM_N596 ));
NOR2_X2 _GFM_U1794  ( .A1(_GFM_n24880 ), .A2(_GFM_n25980 ), .ZN(_GFM_N599 ));
NOR2_X2 _GFM_U1793  ( .A1(_GFM_n24670 ), .A2(_GFM_n26000 ), .ZN(_GFM_N610 ));
NOR2_X2 _GFM_U1792  ( .A1(_GFM_n2417 ), .A2(_GFM_n26050 ), .ZN(_GFM_N614 ));
NOR2_X2 _GFM_U1791  ( .A1(_GFM_n24980 ), .A2(_GFM_n25980 ), .ZN(_GFM_N627 ));
NOR2_X2 _GFM_U1790  ( .A1(_GFM_n24880 ), .A2(_GFM_n2599 ), .ZN(_GFM_N630 ));
NOR2_X2 _GFM_U1789  ( .A1(_GFM_n24670 ), .A2(_GFM_n26010 ), .ZN(_GFM_N641 ));
NOR2_X2 _GFM_U1788  ( .A1(_GFM_n2497 ), .A2(_GFM_n2599 ), .ZN(_GFM_N658 ) );
NOR2_X2 _GFM_U1787  ( .A1(_GFM_n24880 ), .A2(_GFM_n26000 ), .ZN(_GFM_N661 ));
NOR2_X2 _GFM_U1786  ( .A1(_GFM_n2468 ), .A2(_GFM_n2602 ), .ZN(_GFM_N672 ) );
NOR2_X2 _GFM_U1785  ( .A1(_GFM_n2497 ), .A2(_GFM_n26000 ), .ZN(_GFM_N689 ));
NOR2_X2 _GFM_U1784  ( .A1(_GFM_n24880 ), .A2(_GFM_n26010 ), .ZN(_GFM_N692 ));
NOR2_X2 _GFM_U1783  ( .A1(_GFM_n24670 ), .A2(_GFM_n2603 ), .ZN(_GFM_N703 ));
NOR2_X2 _GFM_U1782  ( .A1(_GFM_n2497 ), .A2(_GFM_n26010 ), .ZN(_GFM_N720 ));
NOR2_X2 _GFM_U1781  ( .A1(_GFM_n24880 ), .A2(_GFM_n2602 ), .ZN(_GFM_N723 ));
NOR2_X2 _GFM_U1780  ( .A1(_GFM_n2468 ), .A2(_GFM_n2604 ), .ZN(_GFM_N734 ) );
NOR2_X2 _GFM_U1779  ( .A1(_GFM_n2417 ), .A2(_GFM_n2609 ), .ZN(_GFM_N738 ) );
NOR2_X2 _GFM_U1778  ( .A1(_GFM_n24870 ), .A2(_GFM_n2603 ), .ZN(_GFM_N754 ));
NOR2_X2 _GFM_U1777  ( .A1(_GFM_n2497 ), .A2(_GFM_n2602 ), .ZN(_GFM_N751 ) );
NOR2_X2 _GFM_U1776  ( .A1(_GFM_n24670 ), .A2(_GFM_n26050 ), .ZN(_GFM_N765 ));
NOR2_X2 _GFM_U1775  ( .A1(_GFM_n2497 ), .A2(_GFM_n2603 ), .ZN(_GFM_N782 ) );
NOR2_X2 _GFM_U1774  ( .A1(_GFM_n2489 ), .A2(_GFM_n2604 ), .ZN(_GFM_N785 ) );
NOR2_X2 _GFM_U1773  ( .A1(_GFM_n24870 ), .A2(_GFM_n26050 ), .ZN(_GFM_N816 ));
NOR2_X2 _GFM_U1772  ( .A1(_GFM_n2497 ), .A2(_GFM_n2604 ), .ZN(_GFM_N813 ) );
NOR2_X2 _GFM_U1771  ( .A1(_GFM_n24670 ), .A2(_GFM_n2609 ), .ZN(_GFM_N889 ));
NOR2_X2 _GFM_U1770  ( .A1(_GFM_n24880 ), .A2(_GFM_n2609 ), .ZN(_GFM_N940 ));
NOR2_X2 _GFM_U1769  ( .A1(_GFM_n2387 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1020 ));
NOR2_X2 _GFM_U1768  ( .A1(_GFM_n2396 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1051 ));
NOR2_X2 _GFM_U1767  ( .A1(_GFM_n2396 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1082 ));
NOR2_X2 _GFM_U1766  ( .A1(_GFM_n24250 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1110 ));
NOR2_X2 _GFM_U1765  ( .A1(_GFM_n2396 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1113 ));
NOR2_X2 _GFM_U1764  ( .A1(_GFM_n2427 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1134 ));
NOR2_X2 _GFM_U1763  ( .A1(_GFM_n24250 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1141 ));
NOR2_X2 _GFM_U1762  ( .A1(_GFM_n2396 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1144 ));
NOR2_X2 _GFM_U1761  ( .A1(_GFM_n24450 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1162 ));
NOR2_X2 _GFM_U1760  ( .A1(_GFM_n2435 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1165 ));
NOR2_X2 _GFM_U1759  ( .A1(_GFM_n24250 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1172 ));
NOR2_X2 _GFM_U1758  ( .A1(_GFM_n2396 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1175 ));
NOR2_X2 _GFM_U1757  ( .A1(_GFM_n24450 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1193 ));
NOR2_X2 _GFM_U1756  ( .A1(_GFM_n2435 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1196 ));
NOR2_X2 _GFM_U1755  ( .A1(_GFM_n24250 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1203 ));
NOR2_X2 _GFM_U1754  ( .A1(_GFM_n2396 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1206 ));
NOR2_X2 _GFM_U1753  ( .A1(_GFM_n24450 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1224 ));
NOR2_X2 _GFM_U1752  ( .A1(_GFM_n2435 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1227 ));
NOR2_X2 _GFM_U1751  ( .A1(_GFM_n24250 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1234 ));
NOR2_X2 _GFM_U1750  ( .A1(_GFM_n2396 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1237 ));
NOR2_X2 _GFM_U1749  ( .A1(_GFM_n24450 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1255 ));
NOR2_X2 _GFM_U1748  ( .A1(_GFM_n2435 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1258 ));
NOR2_X2 _GFM_U1747  ( .A1(_GFM_n2475 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1261 ));
NOR2_X2 _GFM_U1746  ( .A1(_GFM_n24250 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1265 ));
NOR2_X2 _GFM_U1745  ( .A1(_GFM_n2396 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1268 ));
NOR2_X2 _GFM_U1744  ( .A1(_GFM_n24450 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1286 ));
NOR2_X2 _GFM_U1743  ( .A1(_GFM_n2435 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1289 ));
NOR2_X2 _GFM_U1742  ( .A1(_GFM_n2475 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1292 ));
NOR2_X2 _GFM_U1741  ( .A1(_GFM_n24250 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1296 ));
NOR2_X2 _GFM_U1740  ( .A1(_GFM_n24950 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1312 ));
NOR2_X2 _GFM_U1739  ( .A1(_GFM_n2475 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1323 ));
NOR2_X2 _GFM_U1738  ( .A1(_GFM_n24250 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1327 ));
NOR2_X2 _GFM_U1737  ( .A1(_GFM_n24950 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1343 ));
NOR2_X2 _GFM_U1736  ( .A1(_GFM_n25040 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1340 ));
NOR2_X2 _GFM_U1735  ( .A1(_GFM_n2475 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1354 ));
NOR2_X2 _GFM_U1734  ( .A1(_GFM_n24250 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1358 ));
NOR2_X2 _GFM_U1733  ( .A1(_GFM_n24950 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1374 ));
NOR2_X2 _GFM_U1732  ( .A1(_GFM_n25040 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1371 ));
NOR2_X2 _GFM_U1731  ( .A1(_GFM_n2475 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1385 ));
NOR2_X2 _GFM_U1730  ( .A1(_GFM_n24250 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1389 ));
NOR2_X2 _GFM_U1729  ( .A1(_GFM_n24950 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1405 ));
NOR2_X2 _GFM_U1728  ( .A1(_GFM_n25040 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1402 ));
NOR2_X2 _GFM_U1727  ( .A1(_GFM_n2475 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1416 ));
NOR2_X2 _GFM_U1726  ( .A1(_GFM_n24250 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1420 ));
NOR2_X2 _GFM_U1725  ( .A1(_GFM_n24950 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1436 ));
NOR2_X2 _GFM_U1724  ( .A1(_GFM_n25040 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1433 ));
NOR2_X2 _GFM_U1723  ( .A1(_GFM_n2475 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1447 ));
NOR2_X2 _GFM_U1722  ( .A1(_GFM_n2424 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1451 ));
NOR2_X2 _GFM_U1721  ( .A1(_GFM_n24950 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1467 ));
NOR2_X2 _GFM_U1720  ( .A1(_GFM_n25040 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1464 ));
NOR2_X2 _GFM_U1719  ( .A1(_GFM_n24740 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1478 ));
NOR2_X2 _GFM_U1718  ( .A1(_GFM_n2424 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1482 ));
NOR2_X2 _GFM_U1717  ( .A1(_GFM_n24950 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1498 ));
NOR2_X2 _GFM_U1716  ( .A1(_GFM_n25040 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1495 ));
NOR2_X2 _GFM_U1715  ( .A1(_GFM_n24740 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1509 ));
NOR2_X2 _GFM_U1714  ( .A1(_GFM_n2424 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1513 ));
NOR2_X2 _GFM_U1713  ( .A1(_GFM_n24950 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1529 ));
NOR2_X2 _GFM_U1712  ( .A1(_GFM_n25040 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1526 ));
NOR2_X2 _GFM_U1711  ( .A1(_GFM_n24740 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1540 ));
NOR2_X2 _GFM_U1710  ( .A1(_GFM_n2424 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1544 ));
NOR2_X2 _GFM_U1709  ( .A1(_GFM_n24950 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1560 ));
NOR2_X2 _GFM_U1708  ( .A1(_GFM_n25040 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1557 ));
NOR2_X2 _GFM_U1707  ( .A1(_GFM_n24740 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1571 ));
NOR2_X2 _GFM_U1706  ( .A1(_GFM_n2424 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1575 ));
NOR2_X2 _GFM_U1705  ( .A1(_GFM_n24950 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1591 ));
NOR2_X2 _GFM_U1704  ( .A1(_GFM_n25040 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1588 ));
NOR2_X2 _GFM_U1703  ( .A1(_GFM_n24740 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1602 ));
NOR2_X2 _GFM_U1702  ( .A1(_GFM_n2424 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1606 ));
NOR2_X2 _GFM_U1701  ( .A1(_GFM_n25040 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1619 ));
NOR2_X2 _GFM_U1700  ( .A1(_GFM_n2494 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1622 ));
NOR2_X2 _GFM_U1699  ( .A1(_GFM_n24740 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1633 ));
NOR2_X2 _GFM_U1698  ( .A1(_GFM_n2424 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1637 ));
NOR2_X2 _GFM_U1697  ( .A1(_GFM_n25040 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1650 ));
NOR2_X2 _GFM_U1696  ( .A1(_GFM_n2494 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1653 ));
NOR2_X2 _GFM_U1695  ( .A1(_GFM_n24740 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1664 ));
NOR2_X2 _GFM_U1694  ( .A1(_GFM_n2424 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1668 ));
NOR2_X2 _GFM_U1693  ( .A1(_GFM_n25040 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1681 ));
NOR2_X2 _GFM_U1692  ( .A1(_GFM_n2494 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1684 ));
NOR2_X2 _GFM_U1691  ( .A1(_GFM_n24740 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1695 ));
NOR2_X2 _GFM_U1690  ( .A1(_GFM_n2424 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1699 ));
NOR2_X2 _GFM_U1689  ( .A1(_GFM_n2503 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1712 ));
NOR2_X2 _GFM_U1688  ( .A1(_GFM_n2494 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1715 ));
NOR2_X2 _GFM_U1687  ( .A1(_GFM_n24740 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1726 ));
NOR2_X2 _GFM_U1686  ( .A1(_GFM_n2424 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1730 ));
NOR2_X2 _GFM_U1685  ( .A1(_GFM_n2503 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1743 ));
NOR2_X2 _GFM_U1684  ( .A1(_GFM_n2494 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1746 ));
NOR2_X2 _GFM_U1683  ( .A1(_GFM_n24740 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1757 ));
NOR2_X2 _GFM_U1682  ( .A1(_GFM_n2424 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1761 ));
NOR2_X2 _GFM_U1681  ( .A1(_GFM_n2503 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1774 ));
NOR2_X2 _GFM_U1680  ( .A1(_GFM_n2494 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1777 ));
NOR2_X2 _GFM_U1679  ( .A1(_GFM_n24740 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1788 ));
NOR2_X2 _GFM_U1678  ( .A1(_GFM_n2424 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1792 ));
NOR2_X2 _GFM_U1677  ( .A1(_GFM_n2503 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1805 ));
NOR2_X2 _GFM_U1676  ( .A1(_GFM_n2494 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1808 ));
NOR2_X2 _GFM_U1675  ( .A1(_GFM_n24730 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1819 ));
NOR2_X2 _GFM_U1674  ( .A1(_GFM_n2423 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1823 ));
NOR2_X2 _GFM_U1673  ( .A1(_GFM_n2503 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1836 ));
NOR2_X2 _GFM_U1672  ( .A1(_GFM_n2494 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1839 ));
NOR2_X2 _GFM_U1671  ( .A1(_GFM_n24730 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1850 ));
NOR2_X2 _GFM_U1670  ( .A1(_GFM_n2423 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1854 ));
NOR2_X2 _GFM_U1669  ( .A1(_GFM_n2503 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1867 ));
NOR2_X2 _GFM_U1668  ( .A1(_GFM_n2494 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1870 ));
NOR2_X2 _GFM_U1667  ( .A1(_GFM_n24730 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1881 ));
NOR2_X2 _GFM_U1666  ( .A1(_GFM_n2423 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1885 ));
NOR2_X2 _GFM_U1665  ( .A1(_GFM_n2503 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1898 ));
NOR2_X2 _GFM_U1664  ( .A1(_GFM_n2494 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1901 ));
NOR2_X2 _GFM_U1663  ( .A1(_GFM_n24730 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1912 ));
NOR2_X2 _GFM_U1662  ( .A1(_GFM_n2423 ), .A2(_GFM_n2647 ), .ZN(_GFM_N1916 ));
NOR2_X2 _GFM_U1661  ( .A1(_GFM_n2503 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1929 ));
NOR2_X2 _GFM_U1660  ( .A1(_GFM_n2494 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1932 ));
NOR2_X2 _GFM_U1659  ( .A1(_GFM_n24730 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1943 ));
NOR2_X2 _GFM_U1658  ( .A1(_GFM_n2423 ), .A2(_GFM_n2648 ), .ZN(_GFM_N1947 ));
NOR2_X2 _GFM_U1657  ( .A1(_GFM_n2503 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1960 ));
NOR2_X2 _GFM_U1656  ( .A1(_GFM_n2493 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1963 ));
NOR2_X2 _GFM_U1655  ( .A1(_GFM_n24730 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1974 ));
NOR2_X2 _GFM_U1654  ( .A1(_GFM_n2423 ), .A2(_GFM_n2649 ), .ZN(_GFM_N1978 ));
NOR2_X2 _GFM_U1653  ( .A1(_GFM_n2503 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1991 ));
NOR2_X2 _GFM_U1652  ( .A1(_GFM_n2493 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1994 ));
NOR2_X2 _GFM_U1651  ( .A1(_GFM_n24730 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2005 ));
NOR2_X2 _GFM_U1650  ( .A1(_GFM_n2423 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2009 ));
NOR2_X2 _GFM_U1649  ( .A1(_GFM_n2503 ), .A2(_GFM_n26430 ), .ZN(_GFM_N2022 ));
NOR2_X2 _GFM_U1648  ( .A1(_GFM_n2493 ), .A2(_GFM_n2644 ), .ZN(_GFM_N2025 ));
NOR2_X2 _GFM_U1647  ( .A1(_GFM_n24730 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2036 ));
NOR2_X2 _GFM_U1646  ( .A1(_GFM_n2423 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2040 ));
NOR2_X2 _GFM_U1645  ( .A1(_GFM_n2503 ), .A2(_GFM_n2644 ), .ZN(_GFM_N2053 ));
NOR2_X2 _GFM_U1644  ( .A1(_GFM_n2493 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2056 ));
NOR2_X2 _GFM_U1643  ( .A1(_GFM_n24730 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2067 ));
NOR2_X2 _GFM_U1642  ( .A1(_GFM_n2423 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2071 ));
NOR2_X2 _GFM_U1641  ( .A1(_GFM_n2502 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2084 ));
NOR2_X2 _GFM_U1640  ( .A1(_GFM_n2493 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2087 ));
NOR2_X2 _GFM_U1639  ( .A1(_GFM_n24730 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2098 ));
NOR2_X2 _GFM_U1638  ( .A1(_GFM_n2423 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2102 ));
NOR2_X2 _GFM_U1637  ( .A1(_GFM_n2502 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2115 ));
NOR2_X2 _GFM_U1636  ( .A1(_GFM_n2493 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2118 ));
NOR2_X2 _GFM_U1635  ( .A1(_GFM_n24730 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2129 ));
NOR2_X2 _GFM_U1634  ( .A1(_GFM_n2423 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2133 ));
NOR2_X2 _GFM_U1633  ( .A1(_GFM_n2502 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2146 ));
NOR2_X2 _GFM_U1632  ( .A1(_GFM_n2493 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2149 ));
NOR2_X2 _GFM_U1631  ( .A1(_GFM_n2472 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2160 ));
NOR2_X2 _GFM_U1630  ( .A1(_GFM_n24220 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2164 ));
NOR2_X2 _GFM_U1629  ( .A1(_GFM_n2502 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2177 ));
NOR2_X2 _GFM_U1628  ( .A1(_GFM_n2493 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2180 ));
NOR2_X2 _GFM_U1627  ( .A1(_GFM_n2472 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2191 ));
NOR2_X2 _GFM_U1626  ( .A1(_GFM_n24220 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2195 ));
NOR2_X2 _GFM_U1625  ( .A1(_GFM_n2502 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2208 ));
NOR2_X2 _GFM_U1624  ( .A1(_GFM_n2493 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2211 ));
NOR2_X2 _GFM_U1623  ( .A1(_GFM_n2472 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2222 ));
NOR2_X2 _GFM_U1622  ( .A1(_GFM_n24220 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2226 ));
NOR2_X2 _GFM_U1621  ( .A1(_GFM_n2502 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2239 ));
NOR2_X2 _GFM_U1620  ( .A1(_GFM_n2493 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2242 ));
NOR2_X2 _GFM_U1619  ( .A1(_GFM_n2472 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2253 ));
NOR2_X2 _GFM_U1618  ( .A1(_GFM_n24220 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2257 ));
NOR2_X2 _GFM_U1617  ( .A1(_GFM_n2502 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2270 ));
NOR2_X2 _GFM_U1616  ( .A1(_GFM_n2493 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2273 ));
NOR2_X2 _GFM_U1615  ( .A1(_GFM_n2472 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2284 ));
NOR2_X2 _GFM_U1614  ( .A1(_GFM_n24220 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2288 ));
NOR2_X2 _GFM_U1613  ( .A1(_GFM_n2502 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2301 ));
NOR2_X2 _GFM_U1612  ( .A1(_GFM_n2493 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2304 ));
NOR2_X2 _GFM_U1611  ( .A1(_GFM_n2472 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2315 ));
NOR2_X2 _GFM_U1610  ( .A1(_GFM_n24220 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2319 ));
NOR2_X2 _GFM_U1609  ( .A1(_GFM_n2502 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2332 ));
NOR2_X2 _GFM_U1608  ( .A1(_GFM_n24921 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2335 ));
NOR2_X2 _GFM_U1607  ( .A1(_GFM_n2472 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2346 ));
NOR2_X2 _GFM_U1606  ( .A1(_GFM_n24220 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2350 ));
NOR2_X2 _GFM_U1605  ( .A1(_GFM_n2502 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2363 ));
NOR2_X2 _GFM_U1604  ( .A1(_GFM_n24921 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2366 ));
NOR2_X2 _GFM_U1603  ( .A1(_GFM_n2472 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2377 ));
NOR2_X2 _GFM_U1602  ( .A1(_GFM_n24220 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2381 ));
NOR2_X2 _GFM_U1601  ( .A1(_GFM_n2502 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2394 ));
NOR2_X2 _GFM_U1600  ( .A1(_GFM_n24921 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2397 ));
NOR2_X2 _GFM_U1599  ( .A1(_GFM_n2472 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2408 ));
NOR2_X2 _GFM_U1598  ( .A1(_GFM_n24220 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2412 ));
NOR2_X2 _GFM_U1597  ( .A1(_GFM_n2502 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2425 ));
NOR2_X2 _GFM_U1596  ( .A1(_GFM_n24921 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2428 ));
NOR2_X2 _GFM_U1595  ( .A1(_GFM_n2472 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2439 ));
NOR2_X2 _GFM_U1594  ( .A1(_GFM_n24220 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2443 ));
NOR2_X2 _GFM_U1593  ( .A1(_GFM_n25010 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2456 ));
NOR2_X2 _GFM_U1592  ( .A1(_GFM_n24921 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2459 ));
NOR2_X2 _GFM_U1591  ( .A1(_GFM_n2472 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2470 ));
NOR2_X2 _GFM_U1590  ( .A1(_GFM_n24220 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2474 ));
NOR2_X2 _GFM_U1589  ( .A1(_GFM_n25010 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2487 ));
NOR2_X2 _GFM_U1588  ( .A1(_GFM_n24921 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2490 ));
NOR2_X2 _GFM_U1587  ( .A1(_GFM_n2472 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2501 ));
NOR2_X2 _GFM_U1586  ( .A1(_GFM_n24210 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2505 ));
NOR2_X2 _GFM_U1585  ( .A1(_GFM_n25010 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2518 ));
NOR2_X2 _GFM_U1584  ( .A1(_GFM_n24921 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2521 ));
NOR2_X2 _GFM_U1583  ( .A1(_GFM_n2472 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2532 ));
NOR2_X2 _GFM_U1582  ( .A1(_GFM_n24210 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2536 ));
NOR2_X2 _GFM_U1581  ( .A1(_GFM_n25010 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2549 ));
NOR2_X2 _GFM_U1580  ( .A1(_GFM_n24921 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2552 ));
NOR2_X2 _GFM_U1579  ( .A1(_GFM_n2471 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2563 ));
NOR2_X2 _GFM_U1578  ( .A1(_GFM_n24210 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2567 ));
NOR2_X2 _GFM_U1577  ( .A1(_GFM_n25010 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2580 ));
NOR2_X2 _GFM_U1576  ( .A1(_GFM_n24921 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2583 ));
NOR2_X2 _GFM_U1575  ( .A1(_GFM_n2471 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2594 ));
NOR2_X2 _GFM_U1574  ( .A1(_GFM_n24210 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2598 ));
NOR2_X2 _GFM_U1573  ( .A1(_GFM_n25010 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2611 ));
NOR2_X2 _GFM_U1572  ( .A1(_GFM_n24921 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2614 ));
NOR2_X2 _GFM_U1571  ( .A1(_GFM_n2471 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2625 ));
NOR2_X2 _GFM_U1570  ( .A1(_GFM_n24210 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2629 ));
NOR2_X2 _GFM_U1569  ( .A1(_GFM_n25010 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2642 ));
NOR2_X2 _GFM_U1568  ( .A1(_GFM_n24921 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2645 ));
NOR2_X2 _GFM_U1567  ( .A1(_GFM_n2471 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2656 ));
NOR2_X2 _GFM_U1566  ( .A1(_GFM_n24210 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2660 ));
NOR2_X2 _GFM_U1565  ( .A1(_GFM_n25010 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2673 ));
NOR2_X2 _GFM_U1564  ( .A1(_GFM_n24921 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2676 ));
NOR2_X2 _GFM_U1563  ( .A1(_GFM_n2471 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2687 ));
NOR2_X2 _GFM_U1562  ( .A1(_GFM_n25010 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2704 ));
NOR2_X2 _GFM_U1561  ( .A1(_GFM_n24910 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2707 ));
NOR2_X2 _GFM_U1560  ( .A1(_GFM_n2471 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2718 ));
NOR2_X2 _GFM_U1559  ( .A1(_GFM_n25010 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2735 ));
NOR2_X2 _GFM_U1558  ( .A1(_GFM_n24910 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2738 ));
NOR2_X2 _GFM_U1557  ( .A1(_GFM_n2471 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2749 ));
NOR2_X2 _GFM_U1556  ( .A1(_GFM_n25010 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2766 ));
NOR2_X2 _GFM_U1555  ( .A1(_GFM_n24910 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2769 ));
NOR2_X2 _GFM_U1554  ( .A1(_GFM_n2471 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2780 ));
NOR2_X2 _GFM_U1553  ( .A1(_GFM_n25010 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2797 ));
NOR2_X2 _GFM_U1552  ( .A1(_GFM_n24910 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2800 ));
NOR2_X2 _GFM_U1551  ( .A1(_GFM_n2471 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2811 ));
NOR2_X2 _GFM_U1550  ( .A1(_GFM_n25000 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2828 ));
NOR2_X2 _GFM_U1549  ( .A1(_GFM_n24910 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2831 ));
NOR2_X2 _GFM_U1548  ( .A1(_GFM_n25000 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2859 ));
NOR2_X2 _GFM_U1547  ( .A1(_GFM_n24910 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2862 ));
NOR2_X2 _GFM_U1546  ( .A1(_GFM_n25000 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2890 ));
NOR2_X2 _GFM_U1545  ( .A1(_GFM_n24210 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2691 ));
NOR2_X2 _GFM_U1544  ( .A1(_GFM_n24210 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2722 ));
NOR2_X2 _GFM_U1543  ( .A1(_GFM_n24210 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2753 ));
NOR2_X2 _GFM_U1542  ( .A1(_GFM_n24210 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2784 ));
NOR2_X2 _GFM_U1541  ( .A1(_GFM_n24210 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2815 ));
NOR2_X2 _GFM_U1540  ( .A1(_GFM_n2471 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2842 ));
NOR2_X2 _GFM_U1539  ( .A1(_GFM_n24201 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2846 ));
NOR2_X2 _GFM_U1538  ( .A1(_GFM_n2471 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2873 ));
NOR2_X2 _GFM_U1537  ( .A1(_GFM_n24201 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2877 ));
NOR2_X2 _GFM_U1536  ( .A1(_GFM_n24910 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2893 ));
NOR2_X2 _GFM_U1535  ( .A1(_GFM_n2471 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2904 ));
NOR2_X2 _GFM_U1534  ( .A1(_GFM_n24201 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2908 ));
NOR2_X2 _GFM_U1533  ( .A1(_GFM_n25000 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2921 ));
NOR2_X2 _GFM_U1532  ( .A1(_GFM_n24910 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2924 ));
NOR2_X2 _GFM_U1531  ( .A1(_GFM_n24700 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2935 ));
NOR2_X2 _GFM_U1530  ( .A1(_GFM_n24201 ), .A2(_GFM_n26801 ), .ZN(_GFM_N2939 ));
NOR2_X2 _GFM_U1529  ( .A1(_GFM_n25000 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2952 ));
NOR2_X2 _GFM_U1528  ( .A1(_GFM_n24910 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2955 ));
NOR2_X2 _GFM_U1527  ( .A1(_GFM_n24700 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2966 ));
NOR2_X2 _GFM_U1526  ( .A1(_GFM_n24201 ), .A2(_GFM_n26810 ), .ZN(_GFM_N2970 ));
NOR2_X2 _GFM_U1525  ( .A1(_GFM_n25000 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2983 ));
NOR2_X2 _GFM_U1524  ( .A1(_GFM_n24910 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2986 ));
NOR2_X2 _GFM_U1523  ( .A1(_GFM_n24700 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2997 ));
NOR2_X2 _GFM_U1522  ( .A1(_GFM_n24201 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3001 ));
NOR2_X2 _GFM_U1521  ( .A1(_GFM_n25000 ), .A2(_GFM_n2675 ), .ZN(_GFM_N3014 ));
NOR2_X2 _GFM_U1520  ( .A1(_GFM_n24910 ), .A2(_GFM_n26760 ), .ZN(_GFM_N3017 ));
NOR2_X2 _GFM_U1519  ( .A1(_GFM_n24700 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3028 ));
NOR2_X2 _GFM_U1518  ( .A1(_GFM_n24201 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3032 ));
NOR2_X2 _GFM_U1517  ( .A1(_GFM_n25000 ), .A2(_GFM_n26760 ), .ZN(_GFM_N3045 ));
NOR2_X2 _GFM_U1516  ( .A1(_GFM_n24900 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3048 ));
NOR2_X2 _GFM_U1515  ( .A1(_GFM_n24700 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3059 ));
NOR2_X2 _GFM_U1514  ( .A1(_GFM_n24201 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3063 ));
NOR2_X2 _GFM_U1513  ( .A1(_GFM_n25000 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3076 ));
NOR2_X2 _GFM_U1512  ( .A1(_GFM_n24900 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3079 ));
NOR2_X2 _GFM_U1511  ( .A1(_GFM_n24700 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3090 ));
NOR2_X2 _GFM_U1510  ( .A1(_GFM_n24201 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3094 ));
NOR2_X2 _GFM_U1509  ( .A1(_GFM_n25000 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3107 ));
NOR2_X2 _GFM_U1508  ( .A1(_GFM_n24900 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3110 ));
NOR2_X2 _GFM_U1507  ( .A1(_GFM_n24700 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3121 ));
NOR2_X2 _GFM_U1506  ( .A1(_GFM_n24201 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3125 ));
NOR2_X2 _GFM_U1505  ( .A1(_GFM_n25000 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3138 ));
NOR2_X2 _GFM_U1504  ( .A1(_GFM_n24900 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3141 ));
NOR2_X2 _GFM_U1503  ( .A1(_GFM_n24700 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3152 ));
NOR2_X2 _GFM_U1502  ( .A1(_GFM_n24201 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3156 ));
NOR2_X2 _GFM_U1501  ( .A1(_GFM_n2499 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3169 ));
NOR2_X2 _GFM_U1500  ( .A1(_GFM_n24900 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3172 ));
NOR2_X2 _GFM_U1499  ( .A1(_GFM_n24700 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3183 ));
NOR2_X2 _GFM_U1498  ( .A1(_GFM_n24201 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3187 ));
NOR2_X2 _GFM_U1497  ( .A1(_GFM_n2499 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3200 ));
NOR2_X2 _GFM_U1496  ( .A1(_GFM_n24900 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3203 ));
NOR2_X2 _GFM_U1495  ( .A1(_GFM_n24700 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3214 ));
NOR2_X2 _GFM_U1494  ( .A1(_GFM_n24190 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3218 ));
NOR2_X2 _GFM_U1493  ( .A1(_GFM_n2499 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3231 ));
NOR2_X2 _GFM_U1492  ( .A1(_GFM_n24910 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3234 ));
NOR2_X2 _GFM_U1491  ( .A1(_GFM_n24700 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3245 ));
NOR2_X2 _GFM_U1490  ( .A1(_GFM_n24190 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3249 ));
NOR2_X2 _GFM_U1489  ( .A1(_GFM_n2499 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3262 ));
NOR2_X2 _GFM_U1488  ( .A1(_GFM_n24900 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3265 ));
NOR2_X2 _GFM_U1487  ( .A1(_GFM_n24700 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3276 ));
NOR2_X2 _GFM_U1486  ( .A1(_GFM_n24190 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3280 ));
NOR2_X2 _GFM_U1485  ( .A1(_GFM_n2499 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3293 ));
NOR2_X2 _GFM_U1484  ( .A1(_GFM_n25101 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3296 ));
NOR2_X2 _GFM_U1483  ( .A1(_GFM_n24500 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3308 ));
NOR2_X2 _GFM_U1482  ( .A1(_GFM_n2400 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3312 ));
NOR2_X2 _GFM_U1481  ( .A1(_GFM_n2499 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3325 ));
NOR2_X2 _GFM_U1480  ( .A1(_GFM_n25101 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3328 ));
NOR2_X2 _GFM_U1479  ( .A1(_GFM_n2449 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3340 ));
NOR2_X2 _GFM_U1478  ( .A1(_GFM_n2499 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3358 ));
NOR2_X2 _GFM_U1477  ( .A1(_GFM_n25101 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3361 ));
NOR2_X2 _GFM_U1476  ( .A1(_GFM_n2449 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3373 ));
NOR2_X2 _GFM_U1475  ( .A1(_GFM_n2499 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3392 ));
NOR2_X2 _GFM_U1474  ( .A1(_GFM_n25101 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3395 ));
NOR2_X2 _GFM_U1473  ( .A1(_GFM_n24690 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3398 ));
NOR2_X2 _GFM_U1472  ( .A1(_GFM_n2499 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3428 ));
NOR2_X2 _GFM_U1471  ( .A1(_GFM_n25101 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3431 ));
NOR2_X2 _GFM_U1470  ( .A1(_GFM_n24690 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3434 ));
NOR2_X2 _GFM_U1469  ( .A1(_GFM_n24690 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3472 ));
NOR2_X2 _GFM_U1468  ( .A1(_GFM_n2449 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3483 ));
NOR2_X2 _GFM_U1467  ( .A1(_GFM_n24690 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3513 ));
NOR2_X2 _GFM_U1466  ( .A1(_GFM_n24690 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3556 ));
NOR2_X2 _GFM_U1465  ( .A1(_GFM_n2509 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3750 ));
NOR2_X2 _GFM_U1464  ( .A1(_GFM_n2610 ), .A2(_GFM_n24070 ), .ZN(_GFM_N737 ));
NOR2_X2 _GFM_U1463  ( .A1(_GFM_n2610 ), .A2(_GFM_n2516 ), .ZN(_GFM_N1058 ));
NOR2_X2 _GFM_U1462  ( .A1(_GFM_n26080 ), .A2(_GFM_n2506 ), .ZN(_GFM_N969 ));
NOR2_X2 _GFM_U1461  ( .A1(_GFM_n26070 ), .A2(_GFM_n24760 ), .ZN(_GFM_N848 ));
NOR2_X2 _GFM_U1460  ( .A1(_GFM_n26070 ), .A2(_GFM_n2506 ), .ZN(_GFM_N938 ));
NOR2_X2 _GFM_U1459  ( .A1(_GFM_n2606 ), .A2(_GFM_n24070 ), .ZN(_GFM_N613 ));
NOR2_X2 _GFM_U1458  ( .A1(_GFM_n2606 ), .A2(_GFM_n24560 ), .ZN(_GFM_N764 ));
NOR2_X2 _GFM_U1457  ( .A1(_GFM_n26200 ), .A2(_GFM_n24460 ), .ZN(_GFM_N1163 ));
NOR2_X2 _GFM_U1456  ( .A1(_GFM_n26190 ), .A2(_GFM_n24070 ), .ZN(_GFM_N1016 ));
NOR2_X2 _GFM_U1455  ( .A1(_GFM_n26190 ), .A2(_GFM_n24460 ), .ZN(_GFM_N1132 ));
NOR2_X2 _GFM_U1454  ( .A1(_GFM_n26190 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1310 ));
NOR2_X2 _GFM_U1453  ( .A1(_GFM_n2617 ), .A2(_GFM_n24070 ), .ZN(_GFM_N954 ));
NOR2_X2 _GFM_U1452  ( .A1(_GFM_n26120 ), .A2(_GFM_n24460 ), .ZN(_GFM_N915 ));
NOR2_X2 _GFM_U1451  ( .A1(_GFM_n2517 ), .A2(_GFM_n25700 ), .ZN(_GFM_N97 ) );
NOR2_X2 _GFM_U1450  ( .A1(_GFM_n25150 ), .A2(_GFM_n25760 ), .ZN(_GFM_N132 ));
NOR2_X2 _GFM_U1449  ( .A1(_GFM_n25150 ), .A2(_GFM_n2578 ), .ZN(_GFM_N163 ));
NOR2_X2 _GFM_U1448  ( .A1(_GFM_n2610 ), .A2(_GFM_n24870 ), .ZN(_GFM_N971 ));
NOR2_X2 _GFM_U1447  ( .A1(_GFM_n26080 ), .A2(_GFM_n2427 ), .ZN(_GFM_N731 ));
NOR2_X2 _GFM_U1446  ( .A1(_GFM_n2606 ), .A2(_GFM_n24460 ), .ZN(_GFM_N729 ));
NOR2_X2 _GFM_U1445  ( .A1(_GFM_n26080 ), .A2(_GFM_n2387 ), .ZN(_GFM_N617 ));
NOR2_X2 _GFM_U1444  ( .A1(_GFM_n26070 ), .A2(_GFM_n2437 ), .ZN(_GFM_N728 ));
NOR2_X2 _GFM_U1443  ( .A1(_GFM_n24770 ), .A2(_GFM_n2603 ), .ZN(_GFM_N724 ));
NOR2_X2 _GFM_U1442  ( .A1(_GFM_n26070 ), .A2(_GFM_n2387 ), .ZN(_GFM_N586 ));
NOR2_X2 _GFM_U1441  ( .A1(_GFM_n26070 ), .A2(_GFM_n25530 ), .ZN(_GFM_N676 ));
NOR2_X2 _GFM_U1440  ( .A1(_GFM_n26070 ), .A2(_GFM_n2466 ), .ZN(_GFM_N827 ));
NOR2_X2 _GFM_U1439  ( .A1(_GFM_n26070 ), .A2(_GFM_n24870 ), .ZN(_GFM_N878 ));
NOR2_X2 _GFM_U1438  ( .A1(_GFM_n2606 ), .A2(_GFM_n2427 ), .ZN(_GFM_N669 ) );
NOR2_X2 _GFM_U1437  ( .A1(_GFM_n2448 ), .A2(_GFM_n2604 ), .ZN(_GFM_N667 ) );
NOR2_X2 _GFM_U1436  ( .A1(_GFM_n2606 ), .A2(_GFM_n25530 ), .ZN(_GFM_N645 ));
NOR2_X2 _GFM_U1435  ( .A1(_GFM_n2606 ), .A2(_GFM_n2466 ), .ZN(_GFM_N796 ) );
NOR2_X2 _GFM_U1434  ( .A1(_GFM_n26200 ), .A2(_GFM_n24360 ), .ZN(_GFM_N1131 ));
NOR2_X2 _GFM_U1433  ( .A1(_GFM_n26190 ), .A2(_GFM_n24260 ), .ZN(_GFM_N1072 ));
NOR2_X2 _GFM_U1432  ( .A1(_GFM_n2617 ), .A2(_GFM_n24460 ), .ZN(_GFM_N1070 ));
NOR2_X2 _GFM_U1431  ( .A1(_GFM_n26190 ), .A2(_GFM_n24360 ), .ZN(_GFM_N1100 ));
NOR2_X2 _GFM_U1430  ( .A1(_GFM_n26150 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1096 ));
NOR2_X2 _GFM_U1429  ( .A1(_GFM_n26190 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1250 ));
NOR2_X2 _GFM_U1428  ( .A1(_GFM_n2617 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1248 ));
NOR2_X2 _GFM_U1427  ( .A1(_GFM_n26190 ), .A2(_GFM_n25530 ), .ZN(_GFM_N1048 ));
NOR2_X2 _GFM_U1426  ( .A1(_GFM_n26190 ), .A2(_GFM_n2466 ), .ZN(_GFM_N1199 ));
NOR2_X2 _GFM_U1425  ( .A1(_GFM_n2617 ), .A2(_GFM_n2466 ), .ZN(_GFM_N1137 ));
NOR2_X2 _GFM_U1424  ( .A1(_GFM_n2618 ), .A2(_GFM_n2466 ), .ZN(_GFM_N1168 ));
NOR2_X2 _GFM_U1423  ( .A1(_GFM_n26120 ), .A2(_GFM_n24260 ), .ZN(_GFM_N855 ));
NOR2_X2 _GFM_U1422  ( .A1(_GFM_n26120 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1033 ));
NOR2_X2 _GFM_U1421  ( .A1(_GFM_n2613 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1064 ));
NOR2_X2 _GFM_U1420  ( .A1(_GFM_n26140 ), .A2(_GFM_n24360 ), .ZN(_GFM_N945 ));
NOR2_X2 _GFM_U1419  ( .A1(_GFM_n2610 ), .A2(_GFM_n24760 ), .ZN(_GFM_N941 ));
NOR2_X2 _GFM_U1418  ( .A1(_GFM_n26140 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1095 ));
NOR2_X2 _GFM_U1417  ( .A1(_GFM_n26150 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1126 ));
NOR2_X2 _GFM_U1416  ( .A1(_GFM_n2613 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1124 ));
NOR2_X2 _GFM_U1415  ( .A1(_GFM_n25140 ), .A2(_GFM_n25800 ), .ZN(_GFM_N194 ));
NOR2_X2 _GFM_U1414  ( .A1(_GFM_n24880 ), .A2(_GFM_n25700 ), .ZN(_GFM_N10 ));
NOR2_X2 _GFM_U1413  ( .A1(_GFM_n24980 ), .A2(_GFM_n25700 ), .ZN(_GFM_N38 ));
NOR2_X2 _GFM_U1412  ( .A1(_GFM_n24570 ), .A2(_GFM_n25821 ), .ZN(_GFM_N82 ));
NOR2_X2 _GFM_U1411  ( .A1(_GFM_n2513 ), .A2(_GFM_n25821 ), .ZN(_GFM_N225 ));
NOR2_X2 _GFM_U1410  ( .A1(_GFM_n2489 ), .A2(_GFM_n2573 ), .ZN(_GFM_N41 ) );
NOR2_X2 _GFM_U1409  ( .A1(_GFM_n2497 ), .A2(_GFM_n2573 ), .ZN(_GFM_N69 ) );
NOR2_X2 _GFM_U1408  ( .A1(_GFM_n24730 ), .A2(_GFM_n25760 ), .ZN(_GFM_N21 ));
NOR2_X2 _GFM_U1407  ( .A1(_GFM_n24880 ), .A2(_GFM_n25760 ), .ZN(_GFM_N72 ));
NOR2_X2 _GFM_U1406  ( .A1(_GFM_n2497 ), .A2(_GFM_n25760 ), .ZN(_GFM_N100 ));
NOR2_X2 _GFM_U1405  ( .A1(_GFM_n24650 ), .A2(_GFM_n25840 ), .ZN(_GFM_N113 ));
NOR2_X2 _GFM_U1404  ( .A1(_GFM_n25120 ), .A2(_GFM_n25840 ), .ZN(_GFM_N256 ));
NOR2_X2 _GFM_U1403  ( .A1(_GFM_n2468 ), .A2(_GFM_n2578 ), .ZN(_GFM_N52 ) );
NOR2_X2 _GFM_U1402  ( .A1(_GFM_n24950 ), .A2(_GFM_n2578 ), .ZN(_GFM_N103 ));
NOR2_X2 _GFM_U1401  ( .A1(_GFM_n25050 ), .A2(_GFM_n2578 ), .ZN(_GFM_N131 ));
NOR2_X2 _GFM_U1400  ( .A1(_GFM_n24650 ), .A2(_GFM_n2586 ), .ZN(_GFM_N144 ));
NOR2_X2 _GFM_U1399  ( .A1(_GFM_n2511 ), .A2(_GFM_n2586 ), .ZN(_GFM_N287 ) );
NOR2_X2 _GFM_U1398  ( .A1(_GFM_n25201 ), .A2(_GFM_n2586 ), .ZN(_GFM_N314 ));
NOR2_X2 _GFM_U1397  ( .A1(_GFM_n24670 ), .A2(_GFM_n25800 ), .ZN(_GFM_N83 ));
NOR2_X2 _GFM_U1396  ( .A1(_GFM_n24950 ), .A2(_GFM_n25800 ), .ZN(_GFM_N134 ));
NOR2_X2 _GFM_U1395  ( .A1(_GFM_n25040 ), .A2(_GFM_n25800 ), .ZN(_GFM_N162 ));
NOR2_X2 _GFM_U1394  ( .A1(_GFM_n2475 ), .A2(_GFM_n25821 ), .ZN(_GFM_N114 ));
NOR2_X2 _GFM_U1393  ( .A1(_GFM_n2494 ), .A2(_GFM_n25821 ), .ZN(_GFM_N165 ));
NOR2_X2 _GFM_U1392  ( .A1(_GFM_n2503 ), .A2(_GFM_n25821 ), .ZN(_GFM_N193 ));
NOR2_X2 _GFM_U1391  ( .A1(_GFM_n2413 ), .A2(_GFM_n2587 ), .ZN(_GFM_N24 ) );
NOR2_X2 _GFM_U1390  ( .A1(_GFM_n24640 ), .A2(_GFM_n2587 ), .ZN(_GFM_N175 ));
NOR2_X2 _GFM_U1389  ( .A1(_GFM_n25101 ), .A2(_GFM_n2587 ), .ZN(_GFM_N318 ));
NOR2_X2 _GFM_U1388  ( .A1(_GFM_n25190 ), .A2(_GFM_n2587 ), .ZN(_GFM_N345 ));
NOR2_X2 _GFM_U1387  ( .A1(_GFM_n24340 ), .A2(_GFM_n25840 ), .ZN(_GFM_N18 ));
NOR2_X2 _GFM_U1386  ( .A1(_GFM_n2454 ), .A2(_GFM_n25800 ), .ZN(_GFM_N16 ) );
NOR2_X2 _GFM_U1385  ( .A1(_GFM_n24740 ), .A2(_GFM_n25840 ), .ZN(_GFM_N145 ));
NOR2_X2 _GFM_U1384  ( .A1(_GFM_n2494 ), .A2(_GFM_n25840 ), .ZN(_GFM_N196 ));
NOR2_X2 _GFM_U1383  ( .A1(_GFM_n2502 ), .A2(_GFM_n25840 ), .ZN(_GFM_N224 ));
NOR2_X2 _GFM_U1382  ( .A1(_GFM_n24380 ), .A2(_GFM_n2586 ), .ZN(_GFM_N77 ) );
NOR2_X2 _GFM_U1381  ( .A1(_GFM_n2478 ), .A2(_GFM_n2578 ), .ZN(_GFM_N73 ) );
NOR2_X2 _GFM_U1380  ( .A1(_GFM_n24220 ), .A2(_GFM_n2586 ), .ZN(_GFM_N25 ) );
NOR2_X2 _GFM_U1379  ( .A1(_GFM_n24740 ), .A2(_GFM_n2586 ), .ZN(_GFM_N176 ));
NOR2_X2 _GFM_U1378  ( .A1(_GFM_n2493 ), .A2(_GFM_n2586 ), .ZN(_GFM_N227 ) );
NOR2_X2 _GFM_U1377  ( .A1(_GFM_n25010 ), .A2(_GFM_n2586 ), .ZN(_GFM_N255 ));
NOR2_X2 _GFM_U1376  ( .A1(_GFM_n2427 ), .A2(_GFM_n2587 ), .ZN(_GFM_N80 ) );
NOR2_X2 _GFM_U1375  ( .A1(_GFM_n2448 ), .A2(_GFM_n25840 ), .ZN(_GFM_N78 ) );
NOR2_X2 _GFM_U1374  ( .A1(_GFM_n2418 ), .A2(_GFM_n2587 ), .ZN(_GFM_N56 ) );
NOR2_X2 _GFM_U1373  ( .A1(_GFM_n24730 ), .A2(_GFM_n2587 ), .ZN(_GFM_N207 ));
NOR2_X2 _GFM_U1372  ( .A1(_GFM_n24921 ), .A2(_GFM_n2587 ), .ZN(_GFM_N258 ));
NOR2_X2 _GFM_U1371  ( .A1(_GFM_n25000 ), .A2(_GFM_n2587 ), .ZN(_GFM_N286 ));
NOR2_X2 _GFM_U1370  ( .A1(_GFM_n25890 ), .A2(_GFM_n24570 ), .ZN(_GFM_N237 ));
NOR2_X2 _GFM_U1369  ( .A1(_GFM_n25890 ), .A2(_GFM_n25070 ), .ZN(_GFM_N380 ));
NOR2_X2 _GFM_U1368  ( .A1(_GFM_n25700 ), .A2(_GFM_n25070 ), .ZN(_GFM_N70 ));
NOR2_X2 _GFM_U1367  ( .A1(_GFM_n25890 ), .A2(_GFM_n24870 ), .ZN(_GFM_N320 ));
NOR2_X2 _GFM_U1366  ( .A1(_GFM_n25880 ), .A2(_GFM_n23980 ), .ZN(_GFM_N27 ));
NOR2_X2 _GFM_U1365  ( .A1(_GFM_n25880 ), .A2(_GFM_n24070 ), .ZN(_GFM_N55 ));
NOR2_X2 _GFM_U1364  ( .A1(_GFM_n25880 ), .A2(_GFM_n24570 ), .ZN(_GFM_N206 ));
NOR2_X2 _GFM_U1363  ( .A1(_GFM_n25880 ), .A2(_GFM_n25070 ), .ZN(_GFM_N349 ));
NOR2_X2 _GFM_U1362  ( .A1(_GFM_n25880 ), .A2(_GFM_n25530 ), .ZN(_GFM_N87 ));
NOR2_X2 _GFM_U1361  ( .A1(_GFM_n25880 ), .A2(_GFM_n24670 ), .ZN(_GFM_N238 ));
NOR2_X2 _GFM_U1360  ( .A1(_GFM_n25880 ), .A2(_GFM_n24870 ), .ZN(_GFM_N289 ));
NOR2_X2 _GFM_U1359  ( .A1(_GFM_n25620 ), .A2(_GFM_n25070 ), .ZN(_GFM_N8 ) );
NOR2_X2 _GFM_U1358  ( .A1(_GFM_n25660 ), .A2(_GFM_n25070 ), .ZN(_GFM_N39 ));
NOR2_X2 _GFM_U1357  ( .A1(_GFM_n25660 ), .A2(_GFM_n24960 ), .ZN(_GFM_N7 ) );
NOR2_X2 _GFM_U1356  ( .A1(_GFM_n25700 ), .A2(_GFM_n24760 ), .ZN(_GFM_N4332 ));
NOR2_X2 _GFM_U1355  ( .A1(_GFM_n25580 ), .A2(_GFM_n2516 ), .ZN(_GFM_N4 ) );
NOR2_X2 _GFM_U1354  ( .A1(_GFM_n25620 ), .A2(_GFM_n2516 ), .ZN(_GFM_N35 ) );
NOR2_X2 _GFM_U1353  ( .A1(_GFM_n26070 ), .A2(_GFM_n24070 ), .ZN(_GFM_N644 ));
NOR2_X2 _GFM_U1352  ( .A1(_GFM_n26080 ), .A2(_GFM_n24070 ), .ZN(_GFM_N675 ));
NOR2_X2 _GFM_U1351  ( .A1(_GFM_n26080 ), .A2(_GFM_n24250 ), .ZN(_GFM_N707 ));
NOR2_X2 _GFM_U1350  ( .A1(_GFM_n25080 ), .A2(_GFM_n26010 ), .ZN(_GFM_N752 ));
NOR2_X2 _GFM_U1349  ( .A1(_GFM_n2610 ), .A2(_GFM_n24250 ), .ZN(_GFM_N769 ));
NOR2_X2 _GFM_U1348  ( .A1(_GFM_n25080 ), .A2(_GFM_n2603 ), .ZN(_GFM_N814 ));
NOR2_X2 _GFM_U1347  ( .A1(_GFM_n2610 ), .A2(_GFM_n24460 ), .ZN(_GFM_N853 ));
NOR2_X2 _GFM_U1346  ( .A1(_GFM_n26110 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1002 ));
NOR2_X2 _GFM_U1345  ( .A1(_GFM_n2610 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1031 ));
NOR2_X2 _GFM_U1344  ( .A1(_GFM_n26200 ), .A2(_GFM_n24070 ), .ZN(_GFM_N1047 ));
NOR2_X2 _GFM_U1343  ( .A1(_GFM_n26110 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1062 ));
NOR2_X2 _GFM_U1342  ( .A1(_GFM_n26200 ), .A2(_GFM_n25530 ), .ZN(_GFM_N1079 ));
NOR2_X2 _GFM_U1341  ( .A1(_GFM_n26120 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1093 ));
NOR2_X2 _GFM_U1340  ( .A1(_GFM_n26200 ), .A2(_GFM_n25070 ), .ZN(_GFM_N1341 ));
NOR2_X2 _GFM_U1339  ( .A1(_GFM_n25150 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1372 ));
NOR2_X2 _GFM_U1338  ( .A1(_GFM_n25150 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1403 ));
NOR2_X2 _GFM_U1337  ( .A1(_GFM_n25150 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1434 ));
NOR2_X2 _GFM_U1336  ( .A1(_GFM_n25150 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1465 ));
NOR2_X2 _GFM_U1335  ( .A1(_GFM_n25150 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1496 ));
NOR2_X2 _GFM_U1334  ( .A1(_GFM_n25150 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1527 ));
NOR2_X2 _GFM_U1333  ( .A1(_GFM_n25150 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1558 ));
NOR2_X2 _GFM_U1332  ( .A1(_GFM_n25150 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1589 ));
NOR2_X2 _GFM_U1331  ( .A1(_GFM_n24401 ), .A2(_GFM_n25940 ), .ZN(_GFM_N325 ));
NOR2_X2 _GFM_U1330  ( .A1(_GFM_n2480 ), .A2(_GFM_n25901 ), .ZN(_GFM_N321 ));
NOR2_X2 _GFM_U1329  ( .A1(_GFM_n24390 ), .A2(_GFM_n2595 ), .ZN(_GFM_N356 ));
NOR2_X2 _GFM_U1328  ( .A1(_GFM_n2479 ), .A2(_GFM_n25910 ), .ZN(_GFM_N352 ));
NOR2_X2 _GFM_U1327  ( .A1(_GFM_n24390 ), .A2(_GFM_n2596 ), .ZN(_GFM_N387 ));
NOR2_X2 _GFM_U1326  ( .A1(_GFM_n2479 ), .A2(_GFM_n2592 ), .ZN(_GFM_N383 ) );
NOR2_X2 _GFM_U1325  ( .A1(_GFM_n24390 ), .A2(_GFM_n25970 ), .ZN(_GFM_N418 ));
NOR2_X2 _GFM_U1324  ( .A1(_GFM_n2479 ), .A2(_GFM_n25930 ), .ZN(_GFM_N414 ));
NOR2_X2 _GFM_U1323  ( .A1(_GFM_n24380 ), .A2(_GFM_n25980 ), .ZN(_GFM_N449 ));
NOR2_X2 _GFM_U1322  ( .A1(_GFM_n2479 ), .A2(_GFM_n25940 ), .ZN(_GFM_N445 ));
NOR2_X2 _GFM_U1321  ( .A1(_GFM_n24380 ), .A2(_GFM_n2599 ), .ZN(_GFM_N480 ));
NOR2_X2 _GFM_U1320  ( .A1(_GFM_n2478 ), .A2(_GFM_n2595 ), .ZN(_GFM_N476 ) );
NOR2_X2 _GFM_U1319  ( .A1(_GFM_n24380 ), .A2(_GFM_n26000 ), .ZN(_GFM_N511 ));
NOR2_X2 _GFM_U1318  ( .A1(_GFM_n2478 ), .A2(_GFM_n2596 ), .ZN(_GFM_N507 ) );
NOR2_X2 _GFM_U1317  ( .A1(_GFM_n24380 ), .A2(_GFM_n26010 ), .ZN(_GFM_N542 ));
NOR2_X2 _GFM_U1316  ( .A1(_GFM_n2478 ), .A2(_GFM_n25970 ), .ZN(_GFM_N538 ));
NOR2_X2 _GFM_U1315  ( .A1(_GFM_n24380 ), .A2(_GFM_n2602 ), .ZN(_GFM_N573 ));
NOR2_X2 _GFM_U1314  ( .A1(_GFM_n2478 ), .A2(_GFM_n25980 ), .ZN(_GFM_N569 ));
NOR2_X2 _GFM_U1313  ( .A1(_GFM_n2437 ), .A2(_GFM_n2603 ), .ZN(_GFM_N604 ) );
NOR2_X2 _GFM_U1312  ( .A1(_GFM_n2478 ), .A2(_GFM_n2599 ), .ZN(_GFM_N600 ) );
NOR2_X2 _GFM_U1311  ( .A1(_GFM_n24380 ), .A2(_GFM_n2604 ), .ZN(_GFM_N635 ));
NOR2_X2 _GFM_U1310  ( .A1(_GFM_n2478 ), .A2(_GFM_n26000 ), .ZN(_GFM_N631 ));
NOR2_X2 _GFM_U1309  ( .A1(_GFM_n2437 ), .A2(_GFM_n26050 ), .ZN(_GFM_N666 ));
NOR2_X2 _GFM_U1308  ( .A1(_GFM_n2478 ), .A2(_GFM_n26010 ), .ZN(_GFM_N662 ));
NOR2_X2 _GFM_U1307  ( .A1(_GFM_n2478 ), .A2(_GFM_n2602 ), .ZN(_GFM_N693 ) );
NOR2_X2 _GFM_U1306  ( .A1(_GFM_n2606 ), .A2(_GFM_n24360 ), .ZN(_GFM_N697 ));
NOR2_X2 _GFM_U1305  ( .A1(_GFM_n24770 ), .A2(_GFM_n2604 ), .ZN(_GFM_N755 ));
NOR2_X2 _GFM_U1304  ( .A1(_GFM_n26080 ), .A2(_GFM_n24360 ), .ZN(_GFM_N759 ));
NOR2_X2 _GFM_U1303  ( .A1(_GFM_n24380 ), .A2(_GFM_n2609 ), .ZN(_GFM_N790 ));
NOR2_X2 _GFM_U1302  ( .A1(_GFM_n2480 ), .A2(_GFM_n26050 ), .ZN(_GFM_N786 ));
NOR2_X2 _GFM_U1301  ( .A1(_GFM_n2606 ), .A2(_GFM_n24770 ), .ZN(_GFM_N817 ));
NOR2_X2 _GFM_U1300  ( .A1(_GFM_n2610 ), .A2(_GFM_n24360 ), .ZN(_GFM_N821 ));
NOR2_X2 _GFM_U1299  ( .A1(_GFM_n2517 ), .A2(_GFM_n2603 ), .ZN(_GFM_N841 ) );
NOR2_X2 _GFM_U1298  ( .A1(_GFM_n24960 ), .A2(_GFM_n26050 ), .ZN(_GFM_N844 ));
NOR2_X2 _GFM_U1297  ( .A1(_GFM_n26080 ), .A2(_GFM_n24770 ), .ZN(_GFM_N879 ));
NOR2_X2 _GFM_U1296  ( .A1(_GFM_n26120 ), .A2(_GFM_n24360 ), .ZN(_GFM_N883 ));
NOR2_X2 _GFM_U1295  ( .A1(_GFM_n2517 ), .A2(_GFM_n26050 ), .ZN(_GFM_N903 ));
NOR2_X2 _GFM_U1294  ( .A1(_GFM_n24960 ), .A2(_GFM_n26070 ), .ZN(_GFM_N906 ));
NOR2_X2 _GFM_U1293  ( .A1(_GFM_n2441 ), .A2(_GFM_n26150 ), .ZN(_GFM_N976 ));
NOR2_X2 _GFM_U1292  ( .A1(_GFM_n24810 ), .A2(_GFM_n26110 ), .ZN(_GFM_N972 ));
NOR2_X2 _GFM_U1291  ( .A1(_GFM_n24450 ), .A2(_GFM_n25821 ), .ZN(_GFM_N15 ));
NOR2_X2 _GFM_U1290  ( .A1(_GFM_n2485 ), .A2(_GFM_n2573 ), .ZN(_GFM_N11 ) );
NOR2_X2 _GFM_U1289  ( .A1(_GFM_n24380 ), .A2(_GFM_n25840 ), .ZN(_GFM_N46 ));
NOR2_X2 _GFM_U1288  ( .A1(_GFM_n2478 ), .A2(_GFM_n25760 ), .ZN(_GFM_N42 ) );
NOR2_X2 _GFM_U1287  ( .A1(_GFM_n2437 ), .A2(_GFM_n2587 ), .ZN(_GFM_N108 ) );
NOR2_X2 _GFM_U1286  ( .A1(_GFM_n2479 ), .A2(_GFM_n25800 ), .ZN(_GFM_N104 ));
NOR2_X2 _GFM_U1285  ( .A1(_GFM_n2485 ), .A2(_GFM_n25821 ), .ZN(_GFM_N135 ));
NOR2_X2 _GFM_U1284  ( .A1(_GFM_n25880 ), .A2(_GFM_n24360 ), .ZN(_GFM_N139 ));
NOR2_X2 _GFM_U1283  ( .A1(_GFM_n25890 ), .A2(_GFM_n2437 ), .ZN(_GFM_N170 ));
NOR2_X2 _GFM_U1282  ( .A1(_GFM_n24840 ), .A2(_GFM_n25840 ), .ZN(_GFM_N166 ));
NOR2_X2 _GFM_U1281  ( .A1(_GFM_n2616 ), .A2(_GFM_n24360 ), .ZN(_GFM_N1007 ));
NOR2_X2 _GFM_U1280  ( .A1(_GFM_n26120 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1003 ));
NOR2_X2 _GFM_U1279  ( .A1(_GFM_n2617 ), .A2(_GFM_n24360 ), .ZN(_GFM_N1038 ));
NOR2_X2 _GFM_U1278  ( .A1(_GFM_n2613 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1034 ));
NOR2_X2 _GFM_U1277  ( .A1(_GFM_n2618 ), .A2(_GFM_n24360 ), .ZN(_GFM_N1069 ));
NOR2_X2 _GFM_U1276  ( .A1(_GFM_n26140 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1065 ));
NOR2_X2 _GFM_U1275  ( .A1(_GFM_n25050 ), .A2(_GFM_n2618 ), .ZN(_GFM_N1247 ));
NOR2_X2 _GFM_U1274  ( .A1(_GFM_n2525 ), .A2(_GFM_n2616 ), .ZN(_GFM_N1244 ));
NOR2_X2 _GFM_U1273  ( .A1(_GFM_n24450 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1317 ));
NOR2_X2 _GFM_U1272  ( .A1(_GFM_n2485 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1313 ));
NOR2_X2 _GFM_U1271  ( .A1(_GFM_n24450 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1348 ));
NOR2_X2 _GFM_U1270  ( .A1(_GFM_n2485 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1344 ));
NOR2_X2 _GFM_U1269  ( .A1(_GFM_n24450 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1379 ));
NOR2_X2 _GFM_U1268  ( .A1(_GFM_n2485 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1375 ));
NOR2_X2 _GFM_U1267  ( .A1(_GFM_n24450 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1410 ));
NOR2_X2 _GFM_U1266  ( .A1(_GFM_n2485 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1406 ));
NOR2_X2 _GFM_U1265  ( .A1(_GFM_n24450 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1441 ));
NOR2_X2 _GFM_U1264  ( .A1(_GFM_n2485 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1437 ));
NOR2_X2 _GFM_U1263  ( .A1(_GFM_n24450 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1472 ));
NOR2_X2 _GFM_U1262  ( .A1(_GFM_n2485 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1468 ));
NOR2_X2 _GFM_U1261  ( .A1(_GFM_n2444 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1503 ));
NOR2_X2 _GFM_U1260  ( .A1(_GFM_n2485 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1499 ));
NOR2_X2 _GFM_U1259  ( .A1(_GFM_n2444 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1534 ));
NOR2_X2 _GFM_U1258  ( .A1(_GFM_n2485 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1530 ));
NOR2_X2 _GFM_U1257  ( .A1(_GFM_n2444 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1565 ));
NOR2_X2 _GFM_U1256  ( .A1(_GFM_n2485 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1561 ));
NOR2_X2 _GFM_U1255  ( .A1(_GFM_n2444 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1596 ));
NOR2_X2 _GFM_U1254  ( .A1(_GFM_n24840 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1592 ));
NOR2_X2 _GFM_U1253  ( .A1(_GFM_n2444 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1627 ));
NOR2_X2 _GFM_U1252  ( .A1(_GFM_n24840 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1623 ));
NOR2_X2 _GFM_U1251  ( .A1(_GFM_n2444 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1658 ));
NOR2_X2 _GFM_U1250  ( .A1(_GFM_n24840 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1654 ));
NOR2_X2 _GFM_U1249  ( .A1(_GFM_n2444 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1689 ));
NOR2_X2 _GFM_U1248  ( .A1(_GFM_n24840 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1685 ));
NOR2_X2 _GFM_U1247  ( .A1(_GFM_n2444 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1720 ));
NOR2_X2 _GFM_U1246  ( .A1(_GFM_n24840 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1716 ));
NOR2_X2 _GFM_U1245  ( .A1(_GFM_n2444 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1751 ));
NOR2_X2 _GFM_U1244  ( .A1(_GFM_n24840 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1747 ));
NOR2_X2 _GFM_U1243  ( .A1(_GFM_n2444 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1782 ));
NOR2_X2 _GFM_U1242  ( .A1(_GFM_n24840 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1778 ));
NOR2_X2 _GFM_U1241  ( .A1(_GFM_n2444 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1813 ));
NOR2_X2 _GFM_U1240  ( .A1(_GFM_n24840 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1809 ));
NOR2_X2 _GFM_U1239  ( .A1(_GFM_n2444 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1844 ));
NOR2_X2 _GFM_U1238  ( .A1(_GFM_n24840 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1840 ));
NOR2_X2 _GFM_U1237  ( .A1(_GFM_n2444 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1875 ));
NOR2_X2 _GFM_U1236  ( .A1(_GFM_n24840 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1871 ));
NOR2_X2 _GFM_U1235  ( .A1(_GFM_n24430 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1906 ));
NOR2_X2 _GFM_U1234  ( .A1(_GFM_n24840 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1902 ));
NOR2_X2 _GFM_U1233  ( .A1(_GFM_n24430 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1937 ));
NOR2_X2 _GFM_U1232  ( .A1(_GFM_n24840 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1933 ));
NOR2_X2 _GFM_U1231  ( .A1(_GFM_n24430 ), .A2(_GFM_n2647 ), .ZN(_GFM_N1968 ));
NOR2_X2 _GFM_U1230  ( .A1(_GFM_n24830 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1964 ));
NOR2_X2 _GFM_U1229  ( .A1(_GFM_n24430 ), .A2(_GFM_n2648 ), .ZN(_GFM_N1999 ));
NOR2_X2 _GFM_U1228  ( .A1(_GFM_n24830 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1995 ));
NOR2_X2 _GFM_U1227  ( .A1(_GFM_n24430 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2030 ));
NOR2_X2 _GFM_U1226  ( .A1(_GFM_n24830 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2026 ));
NOR2_X2 _GFM_U1225  ( .A1(_GFM_n24430 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2061 ));
NOR2_X2 _GFM_U1224  ( .A1(_GFM_n24830 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2057 ));
NOR2_X2 _GFM_U1223  ( .A1(_GFM_n24430 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2092 ));
NOR2_X2 _GFM_U1222  ( .A1(_GFM_n24830 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2088 ));
NOR2_X2 _GFM_U1221  ( .A1(_GFM_n24430 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2123 ));
NOR2_X2 _GFM_U1220  ( .A1(_GFM_n24830 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2119 ));
NOR2_X2 _GFM_U1219  ( .A1(_GFM_n24430 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2154 ));
NOR2_X2 _GFM_U1218  ( .A1(_GFM_n24830 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2150 ));
NOR2_X2 _GFM_U1217  ( .A1(_GFM_n24430 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2185 ));
NOR2_X2 _GFM_U1216  ( .A1(_GFM_n24830 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2181 ));
NOR2_X2 _GFM_U1215  ( .A1(_GFM_n24430 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2216 ));
NOR2_X2 _GFM_U1214  ( .A1(_GFM_n24830 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2212 ));
NOR2_X2 _GFM_U1213  ( .A1(_GFM_n24430 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2247 ));
NOR2_X2 _GFM_U1212  ( .A1(_GFM_n24830 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2243 ));
NOR2_X2 _GFM_U1211  ( .A1(_GFM_n24420 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2278 ));
NOR2_X2 _GFM_U1210  ( .A1(_GFM_n24830 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2274 ));
NOR2_X2 _GFM_U1209  ( .A1(_GFM_n24420 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2309 ));
NOR2_X2 _GFM_U1208  ( .A1(_GFM_n2482 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2305 ));
NOR2_X2 _GFM_U1207  ( .A1(_GFM_n24420 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2340 ));
NOR2_X2 _GFM_U1206  ( .A1(_GFM_n2482 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2336 ));
NOR2_X2 _GFM_U1205  ( .A1(_GFM_n24420 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2371 ));
NOR2_X2 _GFM_U1204  ( .A1(_GFM_n2482 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2367 ));
NOR2_X2 _GFM_U1203  ( .A1(_GFM_n24420 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2402 ));
NOR2_X2 _GFM_U1202  ( .A1(_GFM_n2482 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2398 ));
NOR2_X2 _GFM_U1201  ( .A1(_GFM_n24420 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2433 ));
NOR2_X2 _GFM_U1200  ( .A1(_GFM_n2482 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2429 ));
NOR2_X2 _GFM_U1199  ( .A1(_GFM_n24420 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2464 ));
NOR2_X2 _GFM_U1198  ( .A1(_GFM_n2482 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2460 ));
NOR2_X2 _GFM_U1197  ( .A1(_GFM_n24420 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2495 ));
NOR2_X2 _GFM_U1196  ( .A1(_GFM_n2482 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2491 ));
NOR2_X2 _GFM_U1195  ( .A1(_GFM_n24420 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2526 ));
NOR2_X2 _GFM_U1194  ( .A1(_GFM_n2482 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2522 ));
NOR2_X2 _GFM_U1193  ( .A1(_GFM_n24420 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2557 ));
NOR2_X2 _GFM_U1192  ( .A1(_GFM_n2482 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2553 ));
NOR2_X2 _GFM_U1191  ( .A1(_GFM_n24420 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2588 ));
NOR2_X2 _GFM_U1190  ( .A1(_GFM_n2482 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2584 ));
NOR2_X2 _GFM_U1189  ( .A1(_GFM_n24420 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2619 ));
NOR2_X2 _GFM_U1188  ( .A1(_GFM_n2482 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2615 ));
NOR2_X2 _GFM_U1187  ( .A1(_GFM_n2441 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2650 ));
NOR2_X2 _GFM_U1186  ( .A1(_GFM_n2482 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2646 ));
NOR2_X2 _GFM_U1185  ( .A1(_GFM_n2441 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2681 ));
NOR2_X2 _GFM_U1184  ( .A1(_GFM_n2482 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2677 ));
NOR2_X2 _GFM_U1183  ( .A1(_GFM_n2441 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2712 ));
NOR2_X2 _GFM_U1182  ( .A1(_GFM_n24810 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2708 ));
NOR2_X2 _GFM_U1181  ( .A1(_GFM_n2441 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2743 ));
NOR2_X2 _GFM_U1180  ( .A1(_GFM_n24810 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2739 ));
NOR2_X2 _GFM_U1179  ( .A1(_GFM_n2441 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2774 ));
NOR2_X2 _GFM_U1178  ( .A1(_GFM_n24810 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2770 ));
NOR2_X2 _GFM_U1177  ( .A1(_GFM_n2441 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2805 ));
NOR2_X2 _GFM_U1176  ( .A1(_GFM_n24810 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2801 ));
NOR2_X2 _GFM_U1175  ( .A1(_GFM_n2441 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2836 ));
NOR2_X2 _GFM_U1174  ( .A1(_GFM_n24810 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2832 ));
NOR2_X2 _GFM_U1173  ( .A1(_GFM_n2441 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2867 ));
NOR2_X2 _GFM_U1172  ( .A1(_GFM_n24810 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2863 ));
NOR2_X2 _GFM_U1171  ( .A1(_GFM_n2441 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2898 ));
NOR2_X2 _GFM_U1170  ( .A1(_GFM_n24810 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2894 ));
NOR2_X2 _GFM_U1169  ( .A1(_GFM_n2441 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2929 ));
NOR2_X2 _GFM_U1168  ( .A1(_GFM_n24810 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2925 ));
NOR2_X2 _GFM_U1167  ( .A1(_GFM_n24401 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2960 ));
NOR2_X2 _GFM_U1166  ( .A1(_GFM_n24810 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2956 ));
NOR2_X2 _GFM_U1165  ( .A1(_GFM_n24401 ), .A2(_GFM_n26801 ), .ZN(_GFM_N2991 ));
NOR2_X2 _GFM_U1164  ( .A1(_GFM_n24810 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2987 ));
NOR2_X2 _GFM_U1163  ( .A1(_GFM_n24401 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3022 ));
NOR2_X2 _GFM_U1162  ( .A1(_GFM_n24810 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3018 ));
NOR2_X2 _GFM_U1161  ( .A1(_GFM_n24401 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3053 ));
NOR2_X2 _GFM_U1160  ( .A1(_GFM_n2480 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3049 ));
NOR2_X2 _GFM_U1159  ( .A1(_GFM_n24401 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3084 ));
NOR2_X2 _GFM_U1158  ( .A1(_GFM_n2480 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3080 ));
NOR2_X2 _GFM_U1157  ( .A1(_GFM_n24401 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3115 ));
NOR2_X2 _GFM_U1156  ( .A1(_GFM_n2480 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3111 ));
NOR2_X2 _GFM_U1155  ( .A1(_GFM_n24401 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3146 ));
NOR2_X2 _GFM_U1154  ( .A1(_GFM_n2480 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3142 ));
NOR2_X2 _GFM_U1153  ( .A1(_GFM_n24401 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3177 ));
NOR2_X2 _GFM_U1152  ( .A1(_GFM_n2480 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3173 ));
NOR2_X2 _GFM_U1151  ( .A1(_GFM_n24401 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3208 ));
NOR2_X2 _GFM_U1150  ( .A1(_GFM_n2480 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3204 ));
NOR2_X2 _GFM_U1149  ( .A1(_GFM_n24401 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3239 ));
NOR2_X2 _GFM_U1148  ( .A1(_GFM_n24810 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3235 ));
NOR2_X2 _GFM_U1147  ( .A1(_GFM_n24401 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3270 ));
NOR2_X2 _GFM_U1146  ( .A1(_GFM_n2480 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3266 ));
NOR2_X2 _GFM_U1145  ( .A1(_GFM_n24690 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3299 ));
NOR2_X2 _GFM_U1144  ( .A1(_GFM_n2480 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3298 ));
NOR2_X2 _GFM_U1143  ( .A1(_GFM_n24690 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3331 ));
NOR2_X2 _GFM_U1142  ( .A1(_GFM_n2480 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3330 ));
NOR2_X2 _GFM_U1141  ( .A1(_GFM_n24690 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3364 ));
NOR2_X2 _GFM_U1140  ( .A1(_GFM_n2480 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3363 ));
NOR2_X2 _GFM_U1139  ( .A1(_GFM_n24390 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3407 ));
NOR2_X2 _GFM_U1138  ( .A1(_GFM_n2449 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3406 ));
NOR2_X2 _GFM_U1137  ( .A1(_GFM_n24390 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3444 ));
NOR2_X2 _GFM_U1136  ( .A1(_GFM_n2449 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3443 ));
NOR2_X2 _GFM_U1135  ( .A1(_GFM_n2499 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3466 ));
NOR2_X2 _GFM_U1134  ( .A1(_GFM_n25190 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3463 ));
NOR2_X2 _GFM_U1133  ( .A1(_GFM_n2509 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3505 ));
NOR2_X2 _GFM_U1132  ( .A1(_GFM_n25290 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3503 ));
NOR2_X2 _GFM_U1131  ( .A1(_GFM_n25101 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3548 ));
NOR2_X2 _GFM_U1130  ( .A1(_GFM_n25290 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3546 ));
NOR2_X2 _GFM_U1129  ( .A1(_GFM_n2509 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3594 ));
NOR2_X2 _GFM_U1128  ( .A1(_GFM_n2528 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3592 ));
NOR2_X2 _GFM_U1127  ( .A1(_GFM_n2509 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3643 ));
NOR2_X2 _GFM_U1126  ( .A1(_GFM_n2528 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3641 ));
NOR2_X2 _GFM_U1125  ( .A1(_GFM_n2509 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3695 ));
NOR2_X2 _GFM_U1124  ( .A1(_GFM_n2528 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3693 ));
NOR2_X2 _GFM_U1123  ( .A1(_GFM_n2697 ), .A2(_GFM_n25070 ), .ZN(_GFM_N3999 ));
NOR2_X2 _GFM_U1122  ( .A1(_GFM_n2695 ), .A2(_GFM_n25260 ), .ZN(_GFM_N3997 ));
NOR2_X2 _GFM_U1121  ( .A1(_GFM_n25890 ), .A2(_GFM_n24070 ), .ZN(_GFM_N86 ));
NOR2_X2 _GFM_U1120  ( .A1(_GFM_n25080 ), .A2(_GFM_n2573 ), .ZN(_GFM_N101 ));
NOR2_X2 _GFM_U1119  ( .A1(_GFM_n25890 ), .A2(_GFM_n25530 ), .ZN(_GFM_N118 ));
NOR2_X2 _GFM_U1118  ( .A1(_GFM_n24150 ), .A2(_GFM_n25910 ), .ZN(_GFM_N148 ));
NOR2_X2 _GFM_U1117  ( .A1(_GFM_n24140 ), .A2(_GFM_n2592 ), .ZN(_GFM_N179 ));
NOR2_X2 _GFM_U1116  ( .A1(_GFM_n24140 ), .A2(_GFM_n25930 ), .ZN(_GFM_N210 ));
NOR2_X2 _GFM_U1115  ( .A1(_GFM_n2413 ), .A2(_GFM_n25940 ), .ZN(_GFM_N241 ));
NOR2_X2 _GFM_U1114  ( .A1(_GFM_n24430 ), .A2(_GFM_n25901 ), .ZN(_GFM_N201 ));
NOR2_X2 _GFM_U1113  ( .A1(_GFM_n24830 ), .A2(_GFM_n2586 ), .ZN(_GFM_N197 ));
NOR2_X2 _GFM_U1112  ( .A1(_GFM_n24420 ), .A2(_GFM_n25910 ), .ZN(_GFM_N232 ));
NOR2_X2 _GFM_U1111  ( .A1(_GFM_n24830 ), .A2(_GFM_n2587 ), .ZN(_GFM_N228 ));
NOR2_X2 _GFM_U1110  ( .A1(_GFM_n2441 ), .A2(_GFM_n2592 ), .ZN(_GFM_N263 ) );
NOR2_X2 _GFM_U1109  ( .A1(_GFM_n25880 ), .A2(_GFM_n24770 ), .ZN(_GFM_N259 ));
NOR2_X2 _GFM_U1108  ( .A1(_GFM_n2441 ), .A2(_GFM_n25930 ), .ZN(_GFM_N294 ));
NOR2_X2 _GFM_U1107  ( .A1(_GFM_n25890 ), .A2(_GFM_n24770 ), .ZN(_GFM_N290 ));
NOR2_X2 _GFM_U1106  ( .A1(_GFM_n25890 ), .A2(_GFM_n2466 ), .ZN(_GFM_N269 ));
NOR2_X2 _GFM_U1105  ( .A1(_GFM_n24600 ), .A2(_GFM_n25910 ), .ZN(_GFM_N299 ));
NOR2_X2 _GFM_U1104  ( .A1(_GFM_n24600 ), .A2(_GFM_n2592 ), .ZN(_GFM_N330 ));
NOR2_X2 _GFM_U1103  ( .A1(_GFM_n24590 ), .A2(_GFM_n25930 ), .ZN(_GFM_N361 ));
NOR2_X2 _GFM_U1102  ( .A1(_GFM_n2458 ), .A2(_GFM_n25940 ), .ZN(_GFM_N392 ));
NOR2_X2 _GFM_U1101  ( .A1(_GFM_n25890 ), .A2(_GFM_n2516 ), .ZN(_GFM_N407 ));
NOR2_X2 _GFM_U1100  ( .A1(_GFM_n2458 ), .A2(_GFM_n2595 ), .ZN(_GFM_N423 ) );
NOR2_X2 _GFM_U1099  ( .A1(_GFM_n25180 ), .A2(_GFM_n25901 ), .ZN(_GFM_N438 ));
NOR2_X2 _GFM_U1098  ( .A1(_GFM_n2458 ), .A2(_GFM_n2596 ), .ZN(_GFM_N454 ) );
NOR2_X2 _GFM_U1097  ( .A1(_GFM_n2517 ), .A2(_GFM_n25910 ), .ZN(_GFM_N469 ));
NOR2_X2 _GFM_U1096  ( .A1(_GFM_n2458 ), .A2(_GFM_n25970 ), .ZN(_GFM_N485 ));
NOR2_X2 _GFM_U1095  ( .A1(_GFM_n25180 ), .A2(_GFM_n2592 ), .ZN(_GFM_N500 ));
NOR2_X2 _GFM_U1094  ( .A1(_GFM_n2458 ), .A2(_GFM_n25980 ), .ZN(_GFM_N516 ));
NOR2_X2 _GFM_U1093  ( .A1(_GFM_n25180 ), .A2(_GFM_n25930 ), .ZN(_GFM_N531 ));
NOR2_X2 _GFM_U1092  ( .A1(_GFM_n2458 ), .A2(_GFM_n2599 ), .ZN(_GFM_N547 ) );
NOR2_X2 _GFM_U1091  ( .A1(_GFM_n25180 ), .A2(_GFM_n25940 ), .ZN(_GFM_N562 ));
NOR2_X2 _GFM_U1090  ( .A1(_GFM_n24570 ), .A2(_GFM_n26000 ), .ZN(_GFM_N578 ));
NOR2_X2 _GFM_U1089  ( .A1(_GFM_n2517 ), .A2(_GFM_n2595 ), .ZN(_GFM_N593 ) );
NOR2_X2 _GFM_U1088  ( .A1(_GFM_n2458 ), .A2(_GFM_n26010 ), .ZN(_GFM_N609 ));
NOR2_X2 _GFM_U1087  ( .A1(_GFM_n25180 ), .A2(_GFM_n2596 ), .ZN(_GFM_N624 ));
NOR2_X2 _GFM_U1086  ( .A1(_GFM_n2517 ), .A2(_GFM_n25970 ), .ZN(_GFM_N655 ));
NOR2_X2 _GFM_U1085  ( .A1(_GFM_n2517 ), .A2(_GFM_n25980 ), .ZN(_GFM_N686 ));
NOR2_X2 _GFM_U1084  ( .A1(_GFM_n2517 ), .A2(_GFM_n2599 ), .ZN(_GFM_N717 ) );
NOR2_X2 _GFM_U1083  ( .A1(_GFM_n24570 ), .A2(_GFM_n26050 ), .ZN(_GFM_N733 ));
NOR2_X2 _GFM_U1082  ( .A1(_GFM_n2517 ), .A2(_GFM_n26010 ), .ZN(_GFM_N779 ));
NOR2_X2 _GFM_U1081  ( .A1(_GFM_n26070 ), .A2(_GFM_n24560 ), .ZN(_GFM_N795 ));
NOR2_X2 _GFM_U1080  ( .A1(_GFM_n26080 ), .A2(_GFM_n24560 ), .ZN(_GFM_N826 ));
NOR2_X2 _GFM_U1079  ( .A1(_GFM_n26080 ), .A2(_GFM_n2466 ), .ZN(_GFM_N858 ));
NOR2_X2 _GFM_U1078  ( .A1(_GFM_n2517 ), .A2(_GFM_n2604 ), .ZN(_GFM_N872 ) );
NOR2_X2 _GFM_U1077  ( .A1(_GFM_n2610 ), .A2(_GFM_n24560 ), .ZN(_GFM_N888 ));
NOR2_X2 _GFM_U1076  ( .A1(_GFM_n2610 ), .A2(_GFM_n2466 ), .ZN(_GFM_N920 ) );
NOR2_X2 _GFM_U1075  ( .A1(_GFM_n2525 ), .A2(_GFM_n2573 ), .ZN(_GFM_N128 ) );
NOR2_X2 _GFM_U1074  ( .A1(_GFM_n2524 ), .A2(_GFM_n25760 ), .ZN(_GFM_N159 ));
NOR2_X2 _GFM_U1073  ( .A1(_GFM_n2523 ), .A2(_GFM_n2578 ), .ZN(_GFM_N190 ) );
NOR2_X2 _GFM_U1072  ( .A1(_GFM_n25220 ), .A2(_GFM_n25800 ), .ZN(_GFM_N221 ));
NOR2_X2 _GFM_U1071  ( .A1(_GFM_n2613 ), .A2(_GFM_n24360 ), .ZN(_GFM_N914 ));
NOR2_X2 _GFM_U1070  ( .A1(_GFM_n2517 ), .A2(_GFM_n2606 ), .ZN(_GFM_N934 ) );
NOR2_X2 _GFM_U1069  ( .A1(_GFM_n26120 ), .A2(_GFM_n24560 ), .ZN(_GFM_N950 ));
NOR2_X2 _GFM_U1068  ( .A1(_GFM_n24960 ), .A2(_GFM_n2609 ), .ZN(_GFM_N968 ));
NOR2_X2 _GFM_U1067  ( .A1(_GFM_n2461 ), .A2(_GFM_n2613 ), .ZN(_GFM_N981 ) );
NOR2_X2 _GFM_U1066  ( .A1(_GFM_n2458 ), .A2(_GFM_n26140 ), .ZN(_GFM_N1012 ));
NOR2_X2 _GFM_U1065  ( .A1(_GFM_n2617 ), .A2(_GFM_n24560 ), .ZN(_GFM_N1105 ));
NOR2_X2 _GFM_U1064  ( .A1(_GFM_n2616 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1127 ));
NOR2_X2 _GFM_U1063  ( .A1(_GFM_n2618 ), .A2(_GFM_n24560 ), .ZN(_GFM_N1136 ));
NOR2_X2 _GFM_U1062  ( .A1(_GFM_n2617 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1158 ));
NOR2_X2 _GFM_U1061  ( .A1(_GFM_n26190 ), .A2(_GFM_n24560 ), .ZN(_GFM_N1167 ));
NOR2_X2 _GFM_U1060  ( .A1(_GFM_n2618 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1189 ));
NOR2_X2 _GFM_U1059  ( .A1(_GFM_n26200 ), .A2(_GFM_n24560 ), .ZN(_GFM_N1198 ));
NOR2_X2 _GFM_U1058  ( .A1(_GFM_n26190 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1220 ));
NOR2_X2 _GFM_U1057  ( .A1(_GFM_n26200 ), .A2(_GFM_n2466 ), .ZN(_GFM_N1230 ));
NOR2_X2 _GFM_U1056  ( .A1(_GFM_n26200 ), .A2(_GFM_n24760 ), .ZN(_GFM_N1251 ));
NOR2_X2 _GFM_U1055  ( .A1(_GFM_n24650 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1260 ));
NOR2_X2 _GFM_U1054  ( .A1(_GFM_n2485 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1282 ));
NOR2_X2 _GFM_U1053  ( .A1(_GFM_n24650 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1291 ));
NOR2_X2 _GFM_U1052  ( .A1(_GFM_n2525 ), .A2(_GFM_n2618 ), .ZN(_GFM_N1306 ));
NOR2_X2 _GFM_U1051  ( .A1(_GFM_n24650 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1322 ));
NOR2_X2 _GFM_U1050  ( .A1(_GFM_n24650 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1353 ));
NOR2_X2 _GFM_U1049  ( .A1(_GFM_n24650 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1384 ));
NOR2_X2 _GFM_U1048  ( .A1(_GFM_n24650 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1415 ));
NOR2_X2 _GFM_U1047  ( .A1(_GFM_n24650 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1446 ));
NOR2_X2 _GFM_U1046  ( .A1(_GFM_n24640 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1477 ));
NOR2_X2 _GFM_U1045  ( .A1(_GFM_n24640 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1508 ));
NOR2_X2 _GFM_U1044  ( .A1(_GFM_n24640 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1539 ));
NOR2_X2 _GFM_U1043  ( .A1(_GFM_n24640 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1570 ));
NOR2_X2 _GFM_U1042  ( .A1(_GFM_n24640 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1601 ));
NOR2_X2 _GFM_U1041  ( .A1(_GFM_n2524 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1616 ));
NOR2_X2 _GFM_U1040  ( .A1(_GFM_n24640 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1632 ));
NOR2_X2 _GFM_U1039  ( .A1(_GFM_n2524 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1647 ));
NOR2_X2 _GFM_U1038  ( .A1(_GFM_n24640 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1663 ));
NOR2_X2 _GFM_U1037  ( .A1(_GFM_n2524 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1678 ));
NOR2_X2 _GFM_U1036  ( .A1(_GFM_n24640 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1694 ));
NOR2_X2 _GFM_U1035  ( .A1(_GFM_n2524 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1709 ));
NOR2_X2 _GFM_U1034  ( .A1(_GFM_n24640 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1725 ));
NOR2_X2 _GFM_U1033  ( .A1(_GFM_n2524 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1740 ));
NOR2_X2 _GFM_U1032  ( .A1(_GFM_n24640 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1756 ));
NOR2_X2 _GFM_U1031  ( .A1(_GFM_n2523 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1771 ));
NOR2_X2 _GFM_U1030  ( .A1(_GFM_n24640 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1787 ));
NOR2_X2 _GFM_U1029  ( .A1(_GFM_n2523 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1802 ));
NOR2_X2 _GFM_U1028  ( .A1(_GFM_n24640 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1818 ));
NOR2_X2 _GFM_U1027  ( .A1(_GFM_n2523 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1833 ));
NOR2_X2 _GFM_U1026  ( .A1(_GFM_n2463 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1849 ));
NOR2_X2 _GFM_U1025  ( .A1(_GFM_n2523 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1864 ));
NOR2_X2 _GFM_U1024  ( .A1(_GFM_n2463 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1880 ));
NOR2_X2 _GFM_U1023  ( .A1(_GFM_n2523 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1895 ));
NOR2_X2 _GFM_U1022  ( .A1(_GFM_n2463 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1911 ));
NOR2_X2 _GFM_U1021  ( .A1(_GFM_n2523 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1926 ));
NOR2_X2 _GFM_U1020  ( .A1(_GFM_n2463 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1942 ));
NOR2_X2 _GFM_U1019  ( .A1(_GFM_n2523 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1957 ));
NOR2_X2 _GFM_U1018  ( .A1(_GFM_n2463 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1973 ));
NOR2_X2 _GFM_U1017  ( .A1(_GFM_n2523 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1988 ));
NOR2_X2 _GFM_U1016  ( .A1(_GFM_n2463 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2004 ));
NOR2_X2 _GFM_U1015  ( .A1(_GFM_n2523 ), .A2(_GFM_n2641 ), .ZN(_GFM_N2019 ));
NOR2_X2 _GFM_U1014  ( .A1(_GFM_n2463 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2035 ));
NOR2_X2 _GFM_U1013  ( .A1(_GFM_n2523 ), .A2(_GFM_n26420 ), .ZN(_GFM_N2050 ));
NOR2_X2 _GFM_U1012  ( .A1(_GFM_n2463 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2066 ));
NOR2_X2 _GFM_U1011  ( .A1(_GFM_n2523 ), .A2(_GFM_n26430 ), .ZN(_GFM_N2081 ));
NOR2_X2 _GFM_U1010  ( .A1(_GFM_n2463 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2097 ));
NOR2_X2 _GFM_U1009  ( .A1(_GFM_n2523 ), .A2(_GFM_n2644 ), .ZN(_GFM_N2112 ));
NOR2_X2 _GFM_U1008  ( .A1(_GFM_n2463 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2128 ));
NOR2_X2 _GFM_U1007  ( .A1(_GFM_n25220 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2143 ));
NOR2_X2 _GFM_U1006  ( .A1(_GFM_n2463 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2159 ));
NOR2_X2 _GFM_U1005  ( .A1(_GFM_n25220 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2174 ));
NOR2_X2 _GFM_U1004  ( .A1(_GFM_n2463 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2190 ));
NOR2_X2 _GFM_U1003  ( .A1(_GFM_n25220 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2205 ));
NOR2_X2 _GFM_U1002  ( .A1(_GFM_n2462 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2221 ));
NOR2_X2 _GFM_U1001  ( .A1(_GFM_n25220 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2236 ));
NOR2_X2 _GFM_U1000  ( .A1(_GFM_n2462 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2252 ));
NOR2_X2 _GFM_U999  ( .A1(_GFM_n25220 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2267 ));
NOR2_X2 _GFM_U998  ( .A1(_GFM_n2462 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2283 ));
NOR2_X2 _GFM_U997  ( .A1(_GFM_n25220 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2298 ));
NOR2_X2 _GFM_U996  ( .A1(_GFM_n2462 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2314 ));
NOR2_X2 _GFM_U995  ( .A1(_GFM_n25220 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2329 ));
NOR2_X2 _GFM_U994  ( .A1(_GFM_n2462 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2345 ) );
NOR2_X2 _GFM_U993  ( .A1(_GFM_n25220 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2360 ));
NOR2_X2 _GFM_U992  ( .A1(_GFM_n2462 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2376 ) );
NOR2_X2 _GFM_U991  ( .A1(_GFM_n25220 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2391 ));
NOR2_X2 _GFM_U990  ( .A1(_GFM_n2462 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2407 ));
NOR2_X2 _GFM_U989  ( .A1(_GFM_n25220 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2422 ));
NOR2_X2 _GFM_U988  ( .A1(_GFM_n2462 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2438 ));
NOR2_X2 _GFM_U987  ( .A1(_GFM_n25220 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2453 ));
NOR2_X2 _GFM_U986  ( .A1(_GFM_n2462 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2469 ));
NOR2_X2 _GFM_U985  ( .A1(_GFM_n25220 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2484 ));
NOR2_X2 _GFM_U984  ( .A1(_GFM_n2462 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2500 ));
NOR2_X2 _GFM_U983  ( .A1(_GFM_n25210 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2515 ));
NOR2_X2 _GFM_U982  ( .A1(_GFM_n2462 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2531 ));
NOR2_X2 _GFM_U981  ( .A1(_GFM_n25210 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2546 ));
NOR2_X2 _GFM_U980  ( .A1(_GFM_n2462 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2562 ) );
NOR2_X2 _GFM_U979  ( .A1(_GFM_n25210 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2577 ));
NOR2_X2 _GFM_U978  ( .A1(_GFM_n2462 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2593 ) );
NOR2_X2 _GFM_U977  ( .A1(_GFM_n25210 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2608 ));
NOR2_X2 _GFM_U976  ( .A1(_GFM_n2461 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2624 ) );
NOR2_X2 _GFM_U975  ( .A1(_GFM_n25210 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2639 ));
NOR2_X2 _GFM_U974  ( .A1(_GFM_n2461 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2655 ));
NOR2_X2 _GFM_U973  ( .A1(_GFM_n25210 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2670 ));
NOR2_X2 _GFM_U972  ( .A1(_GFM_n2461 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2686 ) );
NOR2_X2 _GFM_U971  ( .A1(_GFM_n25210 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2701 ));
NOR2_X2 _GFM_U970  ( .A1(_GFM_n2461 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2717 ));
NOR2_X2 _GFM_U969  ( .A1(_GFM_n25210 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2732 ));
NOR2_X2 _GFM_U968  ( .A1(_GFM_n2461 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2748 ));
NOR2_X2 _GFM_U967  ( .A1(_GFM_n25210 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2763 ));
NOR2_X2 _GFM_U966  ( .A1(_GFM_n2461 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2779 ) );
NOR2_X2 _GFM_U965  ( .A1(_GFM_n25210 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2794 ));
NOR2_X2 _GFM_U964  ( .A1(_GFM_n2461 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2810 ) );
NOR2_X2 _GFM_U963  ( .A1(_GFM_n25210 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2825 ));
NOR2_X2 _GFM_U962  ( .A1(_GFM_n2461 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2841 ));
NOR2_X2 _GFM_U961  ( .A1(_GFM_n25201 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2856 ));
NOR2_X2 _GFM_U960  ( .A1(_GFM_n2461 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2872 ));
NOR2_X2 _GFM_U959  ( .A1(_GFM_n25201 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2887 ));
NOR2_X2 _GFM_U958  ( .A1(_GFM_n2461 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2903 ) );
NOR2_X2 _GFM_U957  ( .A1(_GFM_n25201 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2918 ));
NOR2_X2 _GFM_U956  ( .A1(_GFM_n2461 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2934 ));
NOR2_X2 _GFM_U955  ( .A1(_GFM_n25201 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2949 ));
NOR2_X2 _GFM_U954  ( .A1(_GFM_n24600 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2965 ));
NOR2_X2 _GFM_U953  ( .A1(_GFM_n25201 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2980 ));
NOR2_X2 _GFM_U952  ( .A1(_GFM_n24600 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2996 ));
NOR2_X2 _GFM_U951  ( .A1(_GFM_n25201 ), .A2(_GFM_n26730 ), .ZN(_GFM_N3011 ));
NOR2_X2 _GFM_U950  ( .A1(_GFM_n24600 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3027 ));
NOR2_X2 _GFM_U949  ( .A1(_GFM_n25201 ), .A2(_GFM_n26740 ), .ZN(_GFM_N3042 ));
NOR2_X2 _GFM_U948  ( .A1(_GFM_n24600 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3058 ));
NOR2_X2 _GFM_U947  ( .A1(_GFM_n25201 ), .A2(_GFM_n2675 ), .ZN(_GFM_N3073 ));
NOR2_X2 _GFM_U946  ( .A1(_GFM_n24600 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3089 ));
NOR2_X2 _GFM_U945  ( .A1(_GFM_n25201 ), .A2(_GFM_n26760 ), .ZN(_GFM_N3104 ));
NOR2_X2 _GFM_U944  ( .A1(_GFM_n24600 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3120 ));
NOR2_X2 _GFM_U943  ( .A1(_GFM_n25201 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3135 ));
NOR2_X2 _GFM_U942  ( .A1(_GFM_n24600 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3151 ));
NOR2_X2 _GFM_U941  ( .A1(_GFM_n25201 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3166 ));
NOR2_X2 _GFM_U940  ( .A1(_GFM_n24600 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3182 ));
NOR2_X2 _GFM_U939  ( .A1(_GFM_n25190 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3197 ));
NOR2_X2 _GFM_U938  ( .A1(_GFM_n24600 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3213 ));
NOR2_X2 _GFM_U937  ( .A1(_GFM_n25190 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3228 ));
NOR2_X2 _GFM_U936  ( .A1(_GFM_n24600 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3244 ));
NOR2_X2 _GFM_U935  ( .A1(_GFM_n25190 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3259 ));
NOR2_X2 _GFM_U934  ( .A1(_GFM_n24600 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3275 ));
NOR2_X2 _GFM_U933  ( .A1(_GFM_n25190 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3290 ));
NOR2_X2 _GFM_U932  ( .A1(_GFM_n24190 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3306 ));
NOR2_X2 _GFM_U931  ( .A1(_GFM_n25190 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3322 ));
NOR2_X2 _GFM_U930  ( .A1(_GFM_n25190 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3355 ));
NOR2_X2 _GFM_U929  ( .A1(_GFM_n25190 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3389 ));
NOR2_X2 _GFM_U928  ( .A1(_GFM_n25190 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3425 ));
NOR2_X2 _GFM_U927  ( .A1(_GFM_n2432 ), .A2(_GFM_n2592 ), .ZN(_GFM_N235 ) );
NOR2_X2 _GFM_U926  ( .A1(_GFM_n24520 ), .A2(_GFM_n25901 ), .ZN(_GFM_N233 ));
NOR2_X2 _GFM_U925  ( .A1(_GFM_n2431 ), .A2(_GFM_n25930 ), .ZN(_GFM_N266 ) );
NOR2_X2 _GFM_U924  ( .A1(_GFM_n24511 ), .A2(_GFM_n25910 ), .ZN(_GFM_N264 ));
NOR2_X2 _GFM_U923  ( .A1(_GFM_n2430 ), .A2(_GFM_n25940 ), .ZN(_GFM_N297 ) );
NOR2_X2 _GFM_U922  ( .A1(_GFM_n24511 ), .A2(_GFM_n2592 ), .ZN(_GFM_N295 ) );
NOR2_X2 _GFM_U921  ( .A1(_GFM_n2430 ), .A2(_GFM_n2595 ), .ZN(_GFM_N328 ) );
NOR2_X2 _GFM_U920  ( .A1(_GFM_n24500 ), .A2(_GFM_n25930 ), .ZN(_GFM_N326 ));
NOR2_X2 _GFM_U919  ( .A1(_GFM_n24290 ), .A2(_GFM_n2596 ), .ZN(_GFM_N359 ) );
NOR2_X2 _GFM_U918  ( .A1(_GFM_n2449 ), .A2(_GFM_n25940 ), .ZN(_GFM_N357 ) );
NOR2_X2 _GFM_U917  ( .A1(_GFM_n24280 ), .A2(_GFM_n25970 ), .ZN(_GFM_N390 ));
NOR2_X2 _GFM_U916  ( .A1(_GFM_n2449 ), .A2(_GFM_n2595 ), .ZN(_GFM_N388 ) );
NOR2_X2 _GFM_U915  ( .A1(_GFM_n24280 ), .A2(_GFM_n25980 ), .ZN(_GFM_N421 ));
NOR2_X2 _GFM_U914  ( .A1(_GFM_n2448 ), .A2(_GFM_n2596 ), .ZN(_GFM_N419 ) );
NOR2_X2 _GFM_U913  ( .A1(_GFM_n24290 ), .A2(_GFM_n2599 ), .ZN(_GFM_N452 ) );
NOR2_X2 _GFM_U912  ( .A1(_GFM_n2448 ), .A2(_GFM_n25970 ), .ZN(_GFM_N450 ) );
NOR2_X2 _GFM_U911  ( .A1(_GFM_n24280 ), .A2(_GFM_n26000 ), .ZN(_GFM_N483 ));
NOR2_X2 _GFM_U910  ( .A1(_GFM_n2448 ), .A2(_GFM_n25980 ), .ZN(_GFM_N481 ) );
NOR2_X2 _GFM_U909  ( .A1(_GFM_n24280 ), .A2(_GFM_n26010 ), .ZN(_GFM_N514 ));
NOR2_X2 _GFM_U908  ( .A1(_GFM_n2448 ), .A2(_GFM_n2599 ), .ZN(_GFM_N512 ) );
NOR2_X2 _GFM_U907  ( .A1(_GFM_n24280 ), .A2(_GFM_n2602 ), .ZN(_GFM_N545 ) );
NOR2_X2 _GFM_U906  ( .A1(_GFM_n2448 ), .A2(_GFM_n26000 ), .ZN(_GFM_N543 ) );
NOR2_X2 _GFM_U905  ( .A1(_GFM_n24280 ), .A2(_GFM_n2603 ), .ZN(_GFM_N576 ) );
NOR2_X2 _GFM_U904  ( .A1(_GFM_n2448 ), .A2(_GFM_n26010 ), .ZN(_GFM_N574 ) );
NOR2_X2 _GFM_U903  ( .A1(_GFM_n26070 ), .A2(_GFM_n2427 ), .ZN(_GFM_N700 ) );
NOR2_X2 _GFM_U902  ( .A1(_GFM_n2447 ), .A2(_GFM_n26050 ), .ZN(_GFM_N698 ) );
NOR2_X2 _GFM_U901  ( .A1(_GFM_n24280 ), .A2(_GFM_n2609 ), .ZN(_GFM_N762 ) );
NOR2_X2 _GFM_U900  ( .A1(_GFM_n26070 ), .A2(_GFM_n2447 ), .ZN(_GFM_N760 ) );
NOR2_X2 _GFM_U899  ( .A1(_GFM_n2610 ), .A2(_GFM_n24260 ), .ZN(_GFM_N793 ) );
NOR2_X2 _GFM_U898  ( .A1(_GFM_n26080 ), .A2(_GFM_n24460 ), .ZN(_GFM_N791 ));
NOR2_X2 _GFM_U897  ( .A1(_GFM_n24280 ), .A2(_GFM_n26110 ), .ZN(_GFM_N824 ));
NOR2_X2 _GFM_U896  ( .A1(_GFM_n2447 ), .A2(_GFM_n2609 ), .ZN(_GFM_N822 ) );
NOR2_X2 _GFM_U895  ( .A1(_GFM_n25080 ), .A2(_GFM_n2604 ), .ZN(_GFM_N845 ) );
NOR2_X2 _GFM_U894  ( .A1(_GFM_n2606 ), .A2(_GFM_n2486 ), .ZN(_GFM_N847 ) );
NOR2_X2 _GFM_U893  ( .A1(_GFM_n2447 ), .A2(_GFM_n26110 ), .ZN(_GFM_N884 ) );
NOR2_X2 _GFM_U892  ( .A1(_GFM_n2613 ), .A2(_GFM_n24260 ), .ZN(_GFM_N886 ) );
NOR2_X2 _GFM_U891  ( .A1(_GFM_n2606 ), .A2(_GFM_n25070 ), .ZN(_GFM_N907 ) );
NOR2_X2 _GFM_U890  ( .A1(_GFM_n26080 ), .A2(_GFM_n2486 ), .ZN(_GFM_N909 ) );
NOR2_X2 _GFM_U889  ( .A1(_GFM_n2447 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1008 ));
NOR2_X2 _GFM_U888  ( .A1(_GFM_n2617 ), .A2(_GFM_n24260 ), .ZN(_GFM_N1010 ));
NOR2_X2 _GFM_U887  ( .A1(_GFM_n2618 ), .A2(_GFM_n24260 ), .ZN(_GFM_N1041 ));
NOR2_X2 _GFM_U886  ( .A1(_GFM_n2616 ), .A2(_GFM_n24460 ), .ZN(_GFM_N1039 ));
NOR2_X2 _GFM_U885  ( .A1(_GFM_n26200 ), .A2(_GFM_n24260 ), .ZN(_GFM_N1103 ));
NOR2_X2 _GFM_U884  ( .A1(_GFM_n2618 ), .A2(_GFM_n24460 ), .ZN(_GFM_N1101 ));
NOR2_X2 _GFM_U883  ( .A1(_GFM_n2616 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1157 ) );
NOR2_X2 _GFM_U882  ( .A1(_GFM_n26140 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1155 ));
NOR2_X2 _GFM_U881  ( .A1(_GFM_n2618 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1219 ) );
NOR2_X2 _GFM_U880  ( .A1(_GFM_n2616 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1217 ) );
NOR2_X2 _GFM_U879  ( .A1(_GFM_n26200 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1281 ));
NOR2_X2 _GFM_U878  ( .A1(_GFM_n2618 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1279 ) );
NOR2_X2 _GFM_U877  ( .A1(_GFM_n24340 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1537 ));
NOR2_X2 _GFM_U876  ( .A1(_GFM_n2454 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1535 ));
NOR2_X2 _GFM_U875  ( .A1(_GFM_n24340 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1568 ));
NOR2_X2 _GFM_U874  ( .A1(_GFM_n2454 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1566 ) );
NOR2_X2 _GFM_U873  ( .A1(_GFM_n24340 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1599 ));
NOR2_X2 _GFM_U872  ( .A1(_GFM_n2454 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1597 ) );
NOR2_X2 _GFM_U871  ( .A1(_GFM_n24340 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1630 ));
NOR2_X2 _GFM_U870  ( .A1(_GFM_n2454 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1628 ) );
NOR2_X2 _GFM_U869  ( .A1(_GFM_n24340 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1661 ));
NOR2_X2 _GFM_U868  ( .A1(_GFM_n2454 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1659 ));
NOR2_X2 _GFM_U867  ( .A1(_GFM_n24340 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1692 ));
NOR2_X2 _GFM_U866  ( .A1(_GFM_n2454 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1690 ) );
NOR2_X2 _GFM_U865  ( .A1(_GFM_n24340 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1723 ));
NOR2_X2 _GFM_U864  ( .A1(_GFM_n2454 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1721 ));
NOR2_X2 _GFM_U863  ( .A1(_GFM_n24340 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1754 ));
NOR2_X2 _GFM_U862  ( .A1(_GFM_n2454 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1752 ));
NOR2_X2 _GFM_U861  ( .A1(_GFM_n24340 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1785 ));
NOR2_X2 _GFM_U860  ( .A1(_GFM_n2454 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1783 ));
NOR2_X2 _GFM_U859  ( .A1(_GFM_n24340 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1816 ));
NOR2_X2 _GFM_U858  ( .A1(_GFM_n2454 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1814 ) );
NOR2_X2 _GFM_U857  ( .A1(_GFM_n24340 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1847 ));
NOR2_X2 _GFM_U856  ( .A1(_GFM_n2454 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1845 ));
NOR2_X2 _GFM_U855  ( .A1(_GFM_n24330 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1878 ));
NOR2_X2 _GFM_U854  ( .A1(_GFM_n24530 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1876 ));
NOR2_X2 _GFM_U853  ( .A1(_GFM_n24330 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1909 ));
NOR2_X2 _GFM_U852  ( .A1(_GFM_n24530 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1907 ));
NOR2_X2 _GFM_U851  ( .A1(_GFM_n24330 ), .A2(_GFM_n2647 ), .ZN(_GFM_N1940 ));
NOR2_X2 _GFM_U850  ( .A1(_GFM_n24530 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1938 ));
NOR2_X2 _GFM_U849  ( .A1(_GFM_n24330 ), .A2(_GFM_n2648 ), .ZN(_GFM_N1971 ));
NOR2_X2 _GFM_U848  ( .A1(_GFM_n24530 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1969 ));
NOR2_X2 _GFM_U847  ( .A1(_GFM_n24330 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2095 ));
NOR2_X2 _GFM_U846  ( .A1(_GFM_n24530 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2093 ));
NOR2_X2 _GFM_U845  ( .A1(_GFM_n24330 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2126 ));
NOR2_X2 _GFM_U844  ( .A1(_GFM_n24530 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2124 ));
NOR2_X2 _GFM_U843  ( .A1(_GFM_n24330 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2157 ));
NOR2_X2 _GFM_U842  ( .A1(_GFM_n24530 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2155 ));
NOR2_X2 _GFM_U841  ( .A1(_GFM_n24330 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2188 ));
NOR2_X2 _GFM_U840  ( .A1(_GFM_n24530 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2186 ));
NOR2_X2 _GFM_U839  ( .A1(_GFM_n24330 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2219 ));
NOR2_X2 _GFM_U838  ( .A1(_GFM_n24530 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2217 ));
NOR2_X2 _GFM_U837  ( .A1(_GFM_n2432 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2250 ) );
NOR2_X2 _GFM_U836  ( .A1(_GFM_n24530 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2248 ));
NOR2_X2 _GFM_U835  ( .A1(_GFM_n2432 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2281 ) );
NOR2_X2 _GFM_U834  ( .A1(_GFM_n24520 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2279 ));
NOR2_X2 _GFM_U833  ( .A1(_GFM_n2432 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2312 ));
NOR2_X2 _GFM_U832  ( .A1(_GFM_n24520 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2310 ));
NOR2_X2 _GFM_U831  ( .A1(_GFM_n2432 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2343 ));
NOR2_X2 _GFM_U830  ( .A1(_GFM_n24520 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2341 ));
NOR2_X2 _GFM_U829  ( .A1(_GFM_n2432 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2374 ));
NOR2_X2 _GFM_U828  ( .A1(_GFM_n24520 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2372 ));
NOR2_X2 _GFM_U827  ( .A1(_GFM_n2432 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2405 ));
NOR2_X2 _GFM_U826  ( .A1(_GFM_n24520 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2403 ));
NOR2_X2 _GFM_U825  ( .A1(_GFM_n2432 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2436 ));
NOR2_X2 _GFM_U824  ( .A1(_GFM_n24520 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2434 ));
NOR2_X2 _GFM_U823  ( .A1(_GFM_n2432 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2467 ) );
NOR2_X2 _GFM_U822  ( .A1(_GFM_n24520 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2465 ));
NOR2_X2 _GFM_U821  ( .A1(_GFM_n2432 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2498 ) );
NOR2_X2 _GFM_U820  ( .A1(_GFM_n24520 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2496 ));
NOR2_X2 _GFM_U819  ( .A1(_GFM_n2432 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2529 ) );
NOR2_X2 _GFM_U818  ( .A1(_GFM_n24520 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2527 ));
NOR2_X2 _GFM_U817  ( .A1(_GFM_n2432 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2560 ));
NOR2_X2 _GFM_U816  ( .A1(_GFM_n24520 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2558 ));
NOR2_X2 _GFM_U815  ( .A1(_GFM_n2432 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2591 ) );
NOR2_X2 _GFM_U814  ( .A1(_GFM_n24520 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2589 ));
NOR2_X2 _GFM_U813  ( .A1(_GFM_n2431 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2622 ));
NOR2_X2 _GFM_U812  ( .A1(_GFM_n24520 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2620 ));
NOR2_X2 _GFM_U811  ( .A1(_GFM_n2431 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2653 ));
NOR2_X2 _GFM_U810  ( .A1(_GFM_n24511 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2651 ));
NOR2_X2 _GFM_U809  ( .A1(_GFM_n2431 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2684 ) );
NOR2_X2 _GFM_U808  ( .A1(_GFM_n24511 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2682 ));
NOR2_X2 _GFM_U807  ( .A1(_GFM_n2431 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2715 ) );
NOR2_X2 _GFM_U806  ( .A1(_GFM_n24511 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2713 ));
NOR2_X2 _GFM_U805  ( .A1(_GFM_n2431 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2746 ));
NOR2_X2 _GFM_U804  ( .A1(_GFM_n24511 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2744 ));
NOR2_X2 _GFM_U803  ( .A1(_GFM_n2463 ), .A2(_GFM_n2578 ), .ZN(_GFM_N20 ) );
NOR2_X2 _GFM_U802  ( .A1(_GFM_n25210 ), .A2(_GFM_n25821 ), .ZN(_GFM_N252 ));
NOR2_X2 _GFM_U801  ( .A1(_GFM_n2617 ), .A2(_GFM_n2486 ), .ZN(_GFM_N1188 ) );
NOR2_X2 _GFM_U800  ( .A1(_GFM_n26150 ), .A2(_GFM_n2506 ), .ZN(_GFM_N1186 ));
NOR2_X2 _GFM_U799  ( .A1(_GFM_n2431 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2777 ));
NOR2_X2 _GFM_U798  ( .A1(_GFM_n24511 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2775 ));
NOR2_X2 _GFM_U797  ( .A1(_GFM_n2431 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2808 ) );
NOR2_X2 _GFM_U796  ( .A1(_GFM_n24511 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2806 ));
NOR2_X2 _GFM_U795  ( .A1(_GFM_n2431 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2839 ));
NOR2_X2 _GFM_U794  ( .A1(_GFM_n24511 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2837 ));
NOR2_X2 _GFM_U793  ( .A1(_GFM_n2431 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2870 ));
NOR2_X2 _GFM_U792  ( .A1(_GFM_n24511 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2868 ));
NOR2_X2 _GFM_U791  ( .A1(_GFM_n2431 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2901 ) );
NOR2_X2 _GFM_U790  ( .A1(_GFM_n24511 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2899 ));
NOR2_X2 _GFM_U789  ( .A1(_GFM_n2431 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2932 ) );
NOR2_X2 _GFM_U788  ( .A1(_GFM_n24511 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2930 ));
NOR2_X2 _GFM_U787  ( .A1(_GFM_n2430 ), .A2(_GFM_n26801 ), .ZN(_GFM_N2963 ));
NOR2_X2 _GFM_U786  ( .A1(_GFM_n24500 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2961 ));
NOR2_X2 _GFM_U785  ( .A1(_GFM_n2430 ), .A2(_GFM_n26810 ), .ZN(_GFM_N2994 ));
NOR2_X2 _GFM_U784  ( .A1(_GFM_n24500 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2992 ));
NOR2_X2 _GFM_U783  ( .A1(_GFM_n2430 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3025 ));
NOR2_X2 _GFM_U782  ( .A1(_GFM_n24500 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3023 ));
NOR2_X2 _GFM_U781  ( .A1(_GFM_n2430 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3056 ) );
NOR2_X2 _GFM_U780  ( .A1(_GFM_n24500 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3054 ));
NOR2_X2 _GFM_U779  ( .A1(_GFM_n2430 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3087 ));
NOR2_X2 _GFM_U778  ( .A1(_GFM_n24500 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3085 ));
NOR2_X2 _GFM_U777  ( .A1(_GFM_n2430 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3118 ) );
NOR2_X2 _GFM_U776  ( .A1(_GFM_n24500 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3116 ));
NOR2_X2 _GFM_U775  ( .A1(_GFM_n2430 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3149 ));
NOR2_X2 _GFM_U774  ( .A1(_GFM_n24500 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3147 ));
NOR2_X2 _GFM_U773  ( .A1(_GFM_n2430 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3180 ));
NOR2_X2 _GFM_U772  ( .A1(_GFM_n24500 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3178 ));
NOR2_X2 _GFM_U771  ( .A1(_GFM_n2430 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3211 ) );
NOR2_X2 _GFM_U770  ( .A1(_GFM_n24500 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3209 ));
NOR2_X2 _GFM_U769  ( .A1(_GFM_n2430 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3242 ) );
NOR2_X2 _GFM_U768  ( .A1(_GFM_n24500 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3240 ));
NOR2_X2 _GFM_U767  ( .A1(_GFM_n2430 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3273 ));
NOR2_X2 _GFM_U766  ( .A1(_GFM_n24500 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3271 ));
NOR2_X2 _GFM_U765  ( .A1(_GFM_n24401 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3304 ));
NOR2_X2 _GFM_U764  ( .A1(_GFM_n24290 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3303 ));
NOR2_X2 _GFM_U763  ( .A1(_GFM_n24390 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3336 ));
NOR2_X2 _GFM_U762  ( .A1(_GFM_n24290 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3335 ));
NOR2_X2 _GFM_U761  ( .A1(_GFM_n24390 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3369 ));
NOR2_X2 _GFM_U760  ( .A1(_GFM_n24290 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3368 ));
NOR2_X2 _GFM_U759  ( .A1(_GFM_n25101 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3469 ));
NOR2_X2 _GFM_U758  ( .A1(_GFM_n2489 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3467 ));
NOR2_X2 _GFM_U757  ( .A1(_GFM_n2479 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3509 ));
NOR2_X2 _GFM_U756  ( .A1(_GFM_n2489 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3508 ));
NOR2_X2 _GFM_U754  ( .A1(_GFM_n2479 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3552 ));
NOR2_X2 _GFM_U753  ( .A1(_GFM_n2489 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3551 ));
NOR2_X2 _GFM_U752  ( .A1(_GFM_n2479 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3598 ));
NOR2_X2 _GFM_U751  ( .A1(_GFM_n2489 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3597 ));
NOR2_X2 _GFM_U750  ( .A1(_GFM_n25201 ), .A2(_GFM_n25840 ), .ZN(_GFM_N283 ));
NOR2_X2 _GFM_U749  ( .A1(_GFM_n2458 ), .A2(_GFM_n25800 ), .ZN(_GFM_N51 ) );
NOR2_X2 _GFM_U748  ( .A1(_GFM_n25660 ), .A2(_GFM_n2516 ), .ZN(_GFM_N66 ) );
NOR2_X2 _GFM_U747  ( .A1(_GFM_n25880 ), .A2(_GFM_n24960 ), .ZN(_GFM_N317 ));
NOR2_X2 _GFM_U746  ( .A1(_GFM_n24280 ), .A2(_GFM_n2586 ), .ZN(_GFM_N49 ) );
NOR2_X2 _GFM_U745  ( .A1(_GFM_n2448 ), .A2(_GFM_n25821 ), .ZN(_GFM_N47 ) );
NOR2_X2 _GFM_U744  ( .A1(_GFM_n2455 ), .A2(_GFM_n2586 ), .ZN(_GFM_N109 ) );
NOR2_X2 _GFM_U743  ( .A1(_GFM_n25880 ), .A2(_GFM_n24260 ), .ZN(_GFM_N111 ));
NOR2_X2 _GFM_U742  ( .A1(_GFM_n25890 ), .A2(_GFM_n24960 ), .ZN(_GFM_N348 ));
NOR2_X2 _GFM_U741  ( .A1(_GFM_n25880 ), .A2(_GFM_n2516 ), .ZN(_GFM_N376 ) );
NOR2_X2 _GFM_U740  ( .A1(_GFM_n2455 ), .A2(_GFM_n2587 ), .ZN(_GFM_N140 ) );
NOR2_X2 _GFM_U739  ( .A1(_GFM_n25890 ), .A2(_GFM_n24260 ), .ZN(_GFM_N142 ));
NOR2_X2 _GFM_U738  ( .A1(_GFM_n24340 ), .A2(_GFM_n25901 ), .ZN(_GFM_N173 ));
NOR2_X2 _GFM_U736  ( .A1(_GFM_n25880 ), .A2(_GFM_n24460 ), .ZN(_GFM_N171 ));
INV_X4 _GFM_U735  ( .A(b_in[127]), .ZN(_GFM_n25360 ) );
INV_X4 _GFM_U734  ( .A(b_in[125]), .ZN(_GFM_n2516 ) );
INV_X4 _GFM_U733  ( .A(b_in[116]), .ZN(_GFM_n24260 ) );
INV_X4 _GFM_U732  ( .A(b_in[126]), .ZN(_GFM_n25260 ) );
NOR2_X2 _GFM_U731  ( .A1(_GFM_n25380 ), .A2(_GFM_n2699 ), .ZN(_GFM_N4322 ));
NOR2_X2 _GFM_U730  ( .A1(_GFM_n2696 ), .A2(_GFM_n25360 ), .ZN(_GFM_N4102 ));
NOR2_X2 _GFM_U729  ( .A1(_GFM_n2697 ), .A2(_GFM_n25360 ), .ZN(_GFM_N4159 ));
NOR2_X2 _GFM_U728  ( .A1(_GFM_n2696 ), .A2(_GFM_n2516 ), .ZN(_GFM_N3996 ) );
NOR2_X2 _GFM_U727  ( .A1(_GFM_n25390 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3287 ));
NOR2_X2 _GFM_U726  ( .A1(_GFM_n25390 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3319 ));
NOR2_X2 _GFM_U725  ( .A1(_GFM_n25390 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3352 ));
NOR2_X2 _GFM_U724  ( .A1(_GFM_n25390 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3386 ));
NOR2_X2 _GFM_U723  ( .A1(_GFM_n25390 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3422 ));
NOR2_X2 _GFM_U722  ( .A1(_GFM_n25390 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3460 ));
NOR2_X2 _GFM_U721  ( .A1(_GFM_n25390 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3500 ));
NOR2_X2 _GFM_U720  ( .A1(_GFM_n25390 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3543 ));
NOR2_X2 _GFM_U719  ( .A1(_GFM_n25390 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3589 ));
NOR2_X2 _GFM_U718  ( .A1(_GFM_n2540 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3638 ) );
NOR2_X2 _GFM_U716  ( .A1(_GFM_n25380 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3690 ));
NOR2_X2 _GFM_U715  ( .A1(_GFM_n25380 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3803 ));
NOR2_X2 _GFM_U714  ( .A1(_GFM_n25380 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3864 ));
NOR2_X2 _GFM_U713  ( .A1(_GFM_n2697 ), .A2(_GFM_n25270 ), .ZN(_GFM_N4103 ));
NOR2_X2 _GFM_U712  ( .A1(_GFM_n2479 ), .A2(_GFM_n25500 ), .ZN(_GFM_N4004 ));
NOR2_X2 _GFM_U711  ( .A1(_GFM_n21360 ), .A2(_GFM_n24870 ), .ZN(_GFM_N4006 ));
NOR2_X2 _GFM_U710  ( .A1(_GFM_n25310 ), .A2(_GFM_n26070 ), .ZN(_GFM_N995 ));
NOR2_X2 _GFM_U709  ( .A1(_GFM_n2541 ), .A2(_GFM_n2606 ), .ZN(_GFM_N993 ) );
NOR2_X2 _GFM_U708  ( .A1(_GFM_n23910 ), .A2(_GFM_n26200 ), .ZN(_GFM_N989 ));
NOR2_X2 _GFM_U707  ( .A1(_GFM_n25350 ), .A2(_GFM_n26200 ), .ZN(_GFM_N1398 ));
NOR2_X2 _GFM_U706  ( .A1(_GFM_n25450 ), .A2(_GFM_n26190 ), .ZN(_GFM_N1396 ));
NOR2_X2 _GFM_U705  ( .A1(_GFM_n2389 ), .A2(_GFM_n26190 ), .ZN(_GFM_N958 ) );
NOR2_X2 _GFM_U704  ( .A1(_GFM_n23880 ), .A2(_GFM_n2617 ), .ZN(_GFM_N896 ) );
NOR2_X2 _GFM_U703  ( .A1(_GFM_n25350 ), .A2(_GFM_n2617 ), .ZN(_GFM_N1305 ));
NOR2_X2 _GFM_U702  ( .A1(_GFM_n25450 ), .A2(_GFM_n2616 ), .ZN(_GFM_N1303 ));
NOR2_X2 _GFM_U701  ( .A1(_GFM_n23880 ), .A2(_GFM_n26120 ), .ZN(_GFM_N741 ));
NOR2_X2 _GFM_U700  ( .A1(_GFM_n25350 ), .A2(_GFM_n26120 ), .ZN(_GFM_N1150 ));
NOR2_X2 _GFM_U698  ( .A1(_GFM_n25450 ), .A2(_GFM_n26110 ), .ZN(_GFM_N1148 ));
NOR2_X2 _GFM_U697  ( .A1(_GFM_n23880 ), .A2(_GFM_n2613 ), .ZN(_GFM_N772 ) );
NOR2_X2 _GFM_U696  ( .A1(_GFM_n23880 ), .A2(_GFM_n2616 ), .ZN(_GFM_N865 ) );
NOR2_X2 _GFM_U695  ( .A1(_GFM_n25350 ), .A2(_GFM_n2616 ), .ZN(_GFM_N1274 ));
NOR2_X2 _GFM_U694  ( .A1(_GFM_n25450 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1272 ));
NOR2_X2 _GFM_U693  ( .A1(_GFM_n23880 ), .A2(_GFM_n26140 ), .ZN(_GFM_N803 ));
NOR2_X2 _GFM_U692  ( .A1(_GFM_n26980 ), .A2(_GFM_n25260 ), .ZN(_GFM_N4160 ));
NOR2_X2 _GFM_U691  ( .A1(_GFM_n2389 ), .A2(_GFM_n26150 ), .ZN(_GFM_N834 ) );
NOR2_X2 _GFM_U690  ( .A1(_GFM_n25350 ), .A2(_GFM_n26150 ), .ZN(_GFM_N1243 ));
NOR2_X2 _GFM_U689  ( .A1(_GFM_n25450 ), .A2(_GFM_n26140 ), .ZN(_GFM_N1241 ));
NOR2_X2 _GFM_U688  ( .A1(_GFM_n23880 ), .A2(_GFM_n26110 ), .ZN(_GFM_N710 ));
NOR2_X2 _GFM_U687  ( .A1(_GFM_n23880 ), .A2(_GFM_n25901 ), .ZN(_GFM_N59 ) );
NOR2_X2 _GFM_U686  ( .A1(_GFM_n23880 ), .A2(_GFM_n25910 ), .ZN(_GFM_N90 ) );
NOR2_X2 _GFM_U685  ( .A1(_GFM_n23950 ), .A2(_GFM_n25930 ), .ZN(_GFM_N152 ));
NOR2_X2 _GFM_U684  ( .A1(_GFM_n23940 ), .A2(_GFM_n25940 ), .ZN(_GFM_N183 ));
NOR2_X2 _GFM_U683  ( .A1(_GFM_n2393 ), .A2(_GFM_n2595 ), .ZN(_GFM_N214 ) );
NOR2_X2 _GFM_U682  ( .A1(_GFM_n2392 ), .A2(_GFM_n2596 ), .ZN(_GFM_N245 ) );
NOR2_X2 _GFM_U681  ( .A1(_GFM_n2528 ), .A2(_GFM_n25901 ), .ZN(_GFM_N468 ) );
NOR2_X2 _GFM_U680  ( .A1(_GFM_n25890 ), .A2(_GFM_n25360 ), .ZN(_GFM_N466 ));
NOR2_X2 _GFM_U678  ( .A1(_GFM_n23880 ), .A2(_GFM_n26050 ), .ZN(_GFM_N524 ));
NOR2_X2 _GFM_U677  ( .A1(_GFM_n25270 ), .A2(_GFM_n25910 ), .ZN(_GFM_N499 ));
NOR2_X2 _GFM_U676  ( .A1(_GFM_n25380 ), .A2(_GFM_n25901 ), .ZN(_GFM_N497 ));
NOR2_X2 _GFM_U675  ( .A1(_GFM_n2528 ), .A2(_GFM_n2592 ), .ZN(_GFM_N530 ) );
NOR2_X2 _GFM_U674  ( .A1(_GFM_n25380 ), .A2(_GFM_n25910 ), .ZN(_GFM_N528 ));
NOR2_X2 _GFM_U673  ( .A1(_GFM_n2528 ), .A2(_GFM_n25930 ), .ZN(_GFM_N561 ) );
NOR2_X2 _GFM_U672  ( .A1(_GFM_n2537 ), .A2(_GFM_n2592 ), .ZN(_GFM_N559 ) );
NOR2_X2 _GFM_U671  ( .A1(_GFM_n2528 ), .A2(_GFM_n25940 ), .ZN(_GFM_N592 ) );
NOR2_X2 _GFM_U670  ( .A1(_GFM_n25380 ), .A2(_GFM_n25930 ), .ZN(_GFM_N590 ));
NOR2_X2 _GFM_U669  ( .A1(_GFM_n23880 ), .A2(_GFM_n2609 ), .ZN(_GFM_N648 ) );
NOR2_X2 _GFM_U668  ( .A1(_GFM_n25270 ), .A2(_GFM_n2595 ), .ZN(_GFM_N623 ) );
NOR2_X2 _GFM_U667  ( .A1(_GFM_n25380 ), .A2(_GFM_n25940 ), .ZN(_GFM_N621 ));
NOR2_X2 _GFM_U666  ( .A1(_GFM_n25270 ), .A2(_GFM_n2596 ), .ZN(_GFM_N654 ) );
NOR2_X2 _GFM_U665  ( .A1(_GFM_n2537 ), .A2(_GFM_n2595 ), .ZN(_GFM_N652 ) );
NOR2_X2 _GFM_U664  ( .A1(_GFM_n2528 ), .A2(_GFM_n25970 ), .ZN(_GFM_N685 ) );
NOR2_X2 _GFM_U663  ( .A1(_GFM_n2537 ), .A2(_GFM_n2596 ), .ZN(_GFM_N683 ) );
NOR2_X2 _GFM_U662  ( .A1(_GFM_n25270 ), .A2(_GFM_n25980 ), .ZN(_GFM_N716 ));
NOR2_X2 _GFM_U661  ( .A1(_GFM_n2537 ), .A2(_GFM_n25970 ), .ZN(_GFM_N714 ) );
NOR2_X2 _GFM_U660  ( .A1(_GFM_n25270 ), .A2(_GFM_n2599 ), .ZN(_GFM_N747 ) );
NOR2_X2 _GFM_U659  ( .A1(_GFM_n25380 ), .A2(_GFM_n25980 ), .ZN(_GFM_N745 ));
NOR2_X2 _GFM_U658  ( .A1(_GFM_n25270 ), .A2(_GFM_n26000 ), .ZN(_GFM_N778 ));
NOR2_X2 _GFM_U657  ( .A1(_GFM_n2537 ), .A2(_GFM_n2599 ), .ZN(_GFM_N776 ) );
NOR2_X2 _GFM_U656  ( .A1(_GFM_n25270 ), .A2(_GFM_n26010 ), .ZN(_GFM_N809 ));
NOR2_X2 _GFM_U655  ( .A1(_GFM_n25390 ), .A2(_GFM_n26000 ), .ZN(_GFM_N807 ));
NOR2_X2 _GFM_U654  ( .A1(_GFM_n2528 ), .A2(_GFM_n2602 ), .ZN(_GFM_N840 ) );
NOR2_X2 _GFM_U653  ( .A1(_GFM_n2537 ), .A2(_GFM_n26010 ), .ZN(_GFM_N838 ) );
NOR2_X2 _GFM_U652  ( .A1(_GFM_n25270 ), .A2(_GFM_n2603 ), .ZN(_GFM_N871 ) );
NOR2_X2 _GFM_U651  ( .A1(_GFM_n2537 ), .A2(_GFM_n2602 ), .ZN(_GFM_N869 ) );
NOR2_X2 _GFM_U650  ( .A1(_GFM_n25270 ), .A2(_GFM_n2604 ), .ZN(_GFM_N902 ) );
NOR2_X2 _GFM_U649  ( .A1(_GFM_n2537 ), .A2(_GFM_n2603 ), .ZN(_GFM_N900 ) );
NOR2_X2 _GFM_U648  ( .A1(_GFM_n25270 ), .A2(_GFM_n26050 ), .ZN(_GFM_N933 ));
NOR2_X2 _GFM_U647  ( .A1(_GFM_n2537 ), .A2(_GFM_n2604 ), .ZN(_GFM_N931 ) );
NOR2_X2 _GFM_U646  ( .A1(_GFM_n25270 ), .A2(_GFM_n2609 ), .ZN(_GFM_N1057 ));
NOR2_X2 _GFM_U645  ( .A1(_GFM_n26080 ), .A2(_GFM_n25360 ), .ZN(_GFM_N1055 ));
NOR2_X2 _GFM_U644  ( .A1(_GFM_n23950 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1299 ));
NOR2_X2 _GFM_U643  ( .A1(_GFM_n23950 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1330 ));
NOR2_X2 _GFM_U642  ( .A1(_GFM_n23950 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1361 ));
NOR2_X2 _GFM_U641  ( .A1(_GFM_n23950 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1392 ));
NOR2_X2 _GFM_U640  ( .A1(_GFM_n23950 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1423 ));
NOR2_X2 _GFM_U639  ( .A1(_GFM_n23950 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1454 ));
NOR2_X2 _GFM_U638  ( .A1(_GFM_n2534 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1429 ) );
NOR2_X2 _GFM_U637  ( .A1(_GFM_n25450 ), .A2(_GFM_n26200 ), .ZN(_GFM_N1427 ));
NOR2_X2 _GFM_U636  ( .A1(_GFM_n23950 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1485 ));
NOR2_X2 _GFM_U635  ( .A1(_GFM_n2534 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1460 ));
NOR2_X2 _GFM_U634  ( .A1(_GFM_n2544 ), .A2(_GFM_n2621 ), .ZN(_GFM_N1458 ) );
NOR2_X2 _GFM_U633  ( .A1(_GFM_n23950 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1516 ));
NOR2_X2 _GFM_U632  ( .A1(_GFM_n2534 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1491 ) );
NOR2_X2 _GFM_U631  ( .A1(_GFM_n2544 ), .A2(_GFM_n26220 ), .ZN(_GFM_N1489 ));
NOR2_X2 _GFM_U630  ( .A1(_GFM_n23950 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1547 ));
NOR2_X2 _GFM_U629  ( .A1(_GFM_n2534 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1522 ));
NOR2_X2 _GFM_U628  ( .A1(_GFM_n2544 ), .A2(_GFM_n2623 ), .ZN(_GFM_N1520 ) );
NOR2_X2 _GFM_U627  ( .A1(_GFM_n23950 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1578 ));
NOR2_X2 _GFM_U626  ( .A1(_GFM_n2534 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1553 ));
NOR2_X2 _GFM_U625  ( .A1(_GFM_n2544 ), .A2(_GFM_n26240 ), .ZN(_GFM_N1551 ));
NOR2_X2 _GFM_U624  ( .A1(_GFM_n23950 ), .A2(_GFM_n26401 ), .ZN(_GFM_N1609 ));
NOR2_X2 _GFM_U623  ( .A1(_GFM_n2534 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1584 ) );
NOR2_X2 _GFM_U622  ( .A1(_GFM_n2544 ), .A2(_GFM_n26250 ), .ZN(_GFM_N1582 ));
NOR2_X2 _GFM_U621  ( .A1(_GFM_n23950 ), .A2(_GFM_n2641 ), .ZN(_GFM_N1640 ));
NOR2_X2 _GFM_U620  ( .A1(_GFM_n2534 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1615 ) );
NOR2_X2 _GFM_U619  ( .A1(_GFM_n2544 ), .A2(_GFM_n2626 ), .ZN(_GFM_N1613 ) );
NOR2_X2 _GFM_U618  ( .A1(_GFM_n23940 ), .A2(_GFM_n26420 ), .ZN(_GFM_N1671 ));
NOR2_X2 _GFM_U617  ( .A1(_GFM_n2534 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1646 ));
NOR2_X2 _GFM_U616  ( .A1(_GFM_n2544 ), .A2(_GFM_n2627 ), .ZN(_GFM_N1644 ) );
NOR2_X2 _GFM_U615  ( .A1(_GFM_n23940 ), .A2(_GFM_n26430 ), .ZN(_GFM_N1702 ));
NOR2_X2 _GFM_U614  ( .A1(_GFM_n2534 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1677 ));
NOR2_X2 _GFM_U613  ( .A1(_GFM_n2544 ), .A2(_GFM_n26280 ), .ZN(_GFM_N1675 ));
NOR2_X2 _GFM_U612  ( .A1(_GFM_n23940 ), .A2(_GFM_n2644 ), .ZN(_GFM_N1733 ));
NOR2_X2 _GFM_U611  ( .A1(_GFM_n2534 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1708 ));
NOR2_X2 _GFM_U610  ( .A1(_GFM_n2544 ), .A2(_GFM_n26290 ), .ZN(_GFM_N1706 ));
NOR2_X2 _GFM_U609  ( .A1(_GFM_n23940 ), .A2(_GFM_n26450 ), .ZN(_GFM_N1764 ));
NOR2_X2 _GFM_U608  ( .A1(_GFM_n2534 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1739 ));
NOR2_X2 _GFM_U607  ( .A1(_GFM_n2544 ), .A2(_GFM_n26301 ), .ZN(_GFM_N1737 ));
NOR2_X2 _GFM_U606  ( .A1(_GFM_n23940 ), .A2(_GFM_n26460 ), .ZN(_GFM_N1795 ));
NOR2_X2 _GFM_U605  ( .A1(_GFM_n2534 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1770 ));
NOR2_X2 _GFM_U604  ( .A1(_GFM_n2544 ), .A2(_GFM_n26310 ), .ZN(_GFM_N1768 ));
NOR2_X2 _GFM_U603  ( .A1(_GFM_n23940 ), .A2(_GFM_n2647 ), .ZN(_GFM_N1826 ));
NOR2_X2 _GFM_U602  ( .A1(_GFM_n2533 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1801 ) );
NOR2_X2 _GFM_U601  ( .A1(_GFM_n2544 ), .A2(_GFM_n26320 ), .ZN(_GFM_N1799 ));
NOR2_X2 _GFM_U600  ( .A1(_GFM_n23940 ), .A2(_GFM_n2648 ), .ZN(_GFM_N1857 ));
NOR2_X2 _GFM_U599  ( .A1(_GFM_n2533 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1832 ) );
NOR2_X2 _GFM_U598  ( .A1(_GFM_n25430 ), .A2(_GFM_n2633 ), .ZN(_GFM_N1830 ));
NOR2_X2 _GFM_U597  ( .A1(_GFM_n23940 ), .A2(_GFM_n2649 ), .ZN(_GFM_N1888 ));
NOR2_X2 _GFM_U596  ( .A1(_GFM_n2533 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1863 ) );
NOR2_X2 _GFM_U595  ( .A1(_GFM_n25430 ), .A2(_GFM_n2634 ), .ZN(_GFM_N1861 ));
NOR2_X2 _GFM_U594  ( .A1(_GFM_n23940 ), .A2(_GFM_n26500 ), .ZN(_GFM_N1919 ));
NOR2_X2 _GFM_U593  ( .A1(_GFM_n2533 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1894 ));
NOR2_X2 _GFM_U592  ( .A1(_GFM_n25430 ), .A2(_GFM_n2635 ), .ZN(_GFM_N1892 ));
NOR2_X2 _GFM_U591  ( .A1(_GFM_n23940 ), .A2(_GFM_n26510 ), .ZN(_GFM_N1950 ));
NOR2_X2 _GFM_U590  ( .A1(_GFM_n2533 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1925 ) );
NOR2_X2 _GFM_U589  ( .A1(_GFM_n25430 ), .A2(_GFM_n26360 ), .ZN(_GFM_N1923 ));
NOR2_X2 _GFM_U588  ( .A1(_GFM_n23940 ), .A2(_GFM_n2652 ), .ZN(_GFM_N1981 ));
NOR2_X2 _GFM_U587  ( .A1(_GFM_n2533 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1956 ));
NOR2_X2 _GFM_U586  ( .A1(_GFM_n25430 ), .A2(_GFM_n2637 ), .ZN(_GFM_N1954 ));
NOR2_X2 _GFM_U585  ( .A1(_GFM_n23940 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2012 ));
NOR2_X2 _GFM_U584  ( .A1(_GFM_n2533 ), .A2(_GFM_n26390 ), .ZN(_GFM_N1987 ));
NOR2_X2 _GFM_U583  ( .A1(_GFM_n25430 ), .A2(_GFM_n26380 ), .ZN(_GFM_N1985 ));
NOR2_X2 _GFM_U582  ( .A1(_GFM_n2393 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2043 ) );
NOR2_X2 _GFM_U581  ( .A1(_GFM_n2533 ), .A2(_GFM_n26401 ), .ZN(_GFM_N2018 ));
NOR2_X2 _GFM_U580  ( .A1(_GFM_n25430 ), .A2(_GFM_n26390 ), .ZN(_GFM_N2016 ));
NOR2_X2 _GFM_U579  ( .A1(_GFM_n2393 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2074 ));
NOR2_X2 _GFM_U578  ( .A1(_GFM_n2533 ), .A2(_GFM_n2641 ), .ZN(_GFM_N2049 ) );
NOR2_X2 _GFM_U577  ( .A1(_GFM_n25430 ), .A2(_GFM_n26401 ), .ZN(_GFM_N2047 ));
NOR2_X2 _GFM_U576  ( .A1(_GFM_n2393 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2105 ));
NOR2_X2 _GFM_U575  ( .A1(_GFM_n2533 ), .A2(_GFM_n26420 ), .ZN(_GFM_N2080 ));
NOR2_X2 _GFM_U574  ( .A1(_GFM_n25430 ), .A2(_GFM_n2641 ), .ZN(_GFM_N2078 ));
NOR2_X2 _GFM_U573  ( .A1(_GFM_n2393 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2136 ) );
NOR2_X2 _GFM_U572  ( .A1(_GFM_n2533 ), .A2(_GFM_n26430 ), .ZN(_GFM_N2111 ));
NOR2_X2 _GFM_U571  ( .A1(_GFM_n25430 ), .A2(_GFM_n26420 ), .ZN(_GFM_N2109 ));
NOR2_X2 _GFM_U570  ( .A1(_GFM_n2393 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2167 ) );
NOR2_X2 _GFM_U569  ( .A1(_GFM_n2533 ), .A2(_GFM_n2644 ), .ZN(_GFM_N2142 ) );
NOR2_X2 _GFM_U568  ( .A1(_GFM_n25430 ), .A2(_GFM_n26430 ), .ZN(_GFM_N2140 ));
NOR2_X2 _GFM_U567  ( .A1(_GFM_n2393 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2198 ));
NOR2_X2 _GFM_U566  ( .A1(_GFM_n25320 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2173 ));
NOR2_X2 _GFM_U565  ( .A1(_GFM_n25430 ), .A2(_GFM_n2644 ), .ZN(_GFM_N2171 ));
NOR2_X2 _GFM_U564  ( .A1(_GFM_n2393 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2229 ));
NOR2_X2 _GFM_U563  ( .A1(_GFM_n25320 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2204 ));
NOR2_X2 _GFM_U562  ( .A1(_GFM_n2542 ), .A2(_GFM_n26450 ), .ZN(_GFM_N2202 ));
NOR2_X2 _GFM_U561  ( .A1(_GFM_n2393 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2260 ));
NOR2_X2 _GFM_U560  ( .A1(_GFM_n25320 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2235 ));
NOR2_X2 _GFM_U559  ( .A1(_GFM_n2542 ), .A2(_GFM_n26460 ), .ZN(_GFM_N2233 ));
NOR2_X2 _GFM_U558  ( .A1(_GFM_n2393 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2291 ));
NOR2_X2 _GFM_U557  ( .A1(_GFM_n25320 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2266 ));
NOR2_X2 _GFM_U556  ( .A1(_GFM_n2542 ), .A2(_GFM_n2647 ), .ZN(_GFM_N2264 ) );
NOR2_X2 _GFM_U555  ( .A1(_GFM_n2393 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2322 ));
NOR2_X2 _GFM_U554  ( .A1(_GFM_n25320 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2297 ));
NOR2_X2 _GFM_U553  ( .A1(_GFM_n2542 ), .A2(_GFM_n2648 ), .ZN(_GFM_N2295 ) );
NOR2_X2 _GFM_U552  ( .A1(_GFM_n2393 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2353 ) );
NOR2_X2 _GFM_U551  ( .A1(_GFM_n25320 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2328 ));
NOR2_X2 _GFM_U550  ( .A1(_GFM_n2542 ), .A2(_GFM_n2649 ), .ZN(_GFM_N2326 ) );
NOR2_X2 _GFM_U549  ( .A1(_GFM_n2393 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2384 ) );
NOR2_X2 _GFM_U548  ( .A1(_GFM_n25320 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2359 ));
NOR2_X2 _GFM_U547  ( .A1(_GFM_n2542 ), .A2(_GFM_n26500 ), .ZN(_GFM_N2357 ));
NOR2_X2 _GFM_U546  ( .A1(_GFM_n2392 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2415 ) );
NOR2_X2 _GFM_U545  ( .A1(_GFM_n25320 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2390 ));
NOR2_X2 _GFM_U544  ( .A1(_GFM_n2542 ), .A2(_GFM_n26510 ), .ZN(_GFM_N2388 ));
NOR2_X2 _GFM_U543  ( .A1(_GFM_n2392 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2446 ));
NOR2_X2 _GFM_U542  ( .A1(_GFM_n25320 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2421 ));
NOR2_X2 _GFM_U541  ( .A1(_GFM_n2542 ), .A2(_GFM_n2652 ), .ZN(_GFM_N2419 ) );
NOR2_X2 _GFM_U540  ( .A1(_GFM_n2392 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2477 ) );
NOR2_X2 _GFM_U539  ( .A1(_GFM_n25320 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2452 ));
NOR2_X2 _GFM_U538  ( .A1(_GFM_n2542 ), .A2(_GFM_n26530 ), .ZN(_GFM_N2450 ));
NOR2_X2 _GFM_U537  ( .A1(_GFM_n2392 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2508 ));
NOR2_X2 _GFM_U536  ( .A1(_GFM_n25320 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2483 ));
NOR2_X2 _GFM_U535  ( .A1(_GFM_n2542 ), .A2(_GFM_n2654 ), .ZN(_GFM_N2481 ) );
NOR2_X2 _GFM_U534  ( .A1(_GFM_n2392 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2539 ));
NOR2_X2 _GFM_U533  ( .A1(_GFM_n25310 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2514 ));
NOR2_X2 _GFM_U532  ( .A1(_GFM_n2542 ), .A2(_GFM_n26550 ), .ZN(_GFM_N2512 ));
NOR2_X2 _GFM_U531  ( .A1(_GFM_n2392 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2570 ) );
NOR2_X2 _GFM_U530  ( .A1(_GFM_n25310 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2545 ));
NOR2_X2 _GFM_U529  ( .A1(_GFM_n2541 ), .A2(_GFM_n26560 ), .ZN(_GFM_N2543 ));
NOR2_X2 _GFM_U528  ( .A1(_GFM_n25310 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2576 ));
NOR2_X2 _GFM_U527  ( .A1(_GFM_n2541 ), .A2(_GFM_n2657 ), .ZN(_GFM_N2574 ) );
NOR2_X2 _GFM_U526  ( .A1(_GFM_n25310 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2607 ));
NOR2_X2 _GFM_U525  ( .A1(_GFM_n2541 ), .A2(_GFM_n2658 ), .ZN(_GFM_N2605 ) );
NOR2_X2 _GFM_U524  ( .A1(_GFM_n25310 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2638 ));
NOR2_X2 _GFM_U523  ( .A1(_GFM_n2541 ), .A2(_GFM_n26590 ), .ZN(_GFM_N2636 ));
NOR2_X2 _GFM_U522  ( .A1(_GFM_n25310 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2669 ));
NOR2_X2 _GFM_U521  ( .A1(_GFM_n2541 ), .A2(_GFM_n26600 ), .ZN(_GFM_N2667 ));
NOR2_X2 _GFM_U520  ( .A1(_GFM_n25310 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2700 ));
NOR2_X2 _GFM_U519  ( .A1(_GFM_n2541 ), .A2(_GFM_n26611 ), .ZN(_GFM_N2698 ));
NOR2_X2 _GFM_U518  ( .A1(_GFM_n25310 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2731 ));
NOR2_X2 _GFM_U517  ( .A1(_GFM_n2541 ), .A2(_GFM_n26620 ), .ZN(_GFM_N2729 ));
NOR2_X2 _GFM_U516  ( .A1(_GFM_n25310 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2762 ));
NOR2_X2 _GFM_U515  ( .A1(_GFM_n2541 ), .A2(_GFM_n26630 ), .ZN(_GFM_N2760 ));
NOR2_X2 _GFM_U514  ( .A1(_GFM_n25310 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2793 ));
NOR2_X2 _GFM_U513  ( .A1(_GFM_n2541 ), .A2(_GFM_n2664 ), .ZN(_GFM_N2791 ) );
NOR2_X2 _GFM_U512  ( .A1(_GFM_n25310 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2824 ));
NOR2_X2 _GFM_U511  ( .A1(_GFM_n2541 ), .A2(_GFM_n2665 ), .ZN(_GFM_N2822 ) );
NOR2_X2 _GFM_U510  ( .A1(_GFM_n2530 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2855 ));
NOR2_X2 _GFM_U509  ( .A1(_GFM_n2541 ), .A2(_GFM_n2666 ), .ZN(_GFM_N2853 ) );
NOR2_X2 _GFM_U508  ( .A1(_GFM_n2530 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2886 ) );
NOR2_X2 _GFM_U507  ( .A1(_GFM_n2540 ), .A2(_GFM_n26670 ), .ZN(_GFM_N2884 ));
NOR2_X2 _GFM_U506  ( .A1(_GFM_n2530 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2917 ));
NOR2_X2 _GFM_U505  ( .A1(_GFM_n2540 ), .A2(_GFM_n2668 ), .ZN(_GFM_N2915 ) );
NOR2_X2 _GFM_U504  ( .A1(_GFM_n2530 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2948 ));
NOR2_X2 _GFM_U503  ( .A1(_GFM_n2540 ), .A2(_GFM_n26690 ), .ZN(_GFM_N2946 ));
NOR2_X2 _GFM_U502  ( .A1(_GFM_n2530 ), .A2(_GFM_n2671 ), .ZN(_GFM_N2979 ) );
NOR2_X2 _GFM_U501  ( .A1(_GFM_n2540 ), .A2(_GFM_n26700 ), .ZN(_GFM_N2977 ));
NOR2_X2 _GFM_U500  ( .A1(_GFM_n2392 ), .A2(_GFM_n2672 ), .ZN(_GFM_N2601 ) );
NOR2_X2 _GFM_U499  ( .A1(_GFM_n2392 ), .A2(_GFM_n26730 ), .ZN(_GFM_N2632 ));
NOR2_X2 _GFM_U498  ( .A1(_GFM_n2392 ), .A2(_GFM_n26740 ), .ZN(_GFM_N2663 ));
NOR2_X2 _GFM_U497  ( .A1(_GFM_n2392 ), .A2(_GFM_n2675 ), .ZN(_GFM_N2694 ) );
NOR2_X2 _GFM_U496  ( .A1(_GFM_n2392 ), .A2(_GFM_n26760 ), .ZN(_GFM_N2725 ));
NOR2_X2 _GFM_U495  ( .A1(_GFM_n2392 ), .A2(_GFM_n26770 ), .ZN(_GFM_N2756 ));
NOR2_X2 _GFM_U494  ( .A1(_GFM_n23910 ), .A2(_GFM_n2678 ), .ZN(_GFM_N2787 ));
NOR2_X2 _GFM_U493  ( .A1(_GFM_n23910 ), .A2(_GFM_n2679 ), .ZN(_GFM_N2818 ));
NOR2_X2 _GFM_U492  ( .A1(_GFM_n23910 ), .A2(_GFM_n26801 ), .ZN(_GFM_N2849 ));
NOR2_X2 _GFM_U491  ( .A1(_GFM_n23910 ), .A2(_GFM_n26810 ), .ZN(_GFM_N2880 ));
NOR2_X2 _GFM_U490  ( .A1(_GFM_n23910 ), .A2(_GFM_n26820 ), .ZN(_GFM_N2911 ));
NOR2_X2 _GFM_U489  ( .A1(_GFM_n23910 ), .A2(_GFM_n2683 ), .ZN(_GFM_N2942 ));
NOR2_X2 _GFM_U488  ( .A1(_GFM_n23910 ), .A2(_GFM_n26840 ), .ZN(_GFM_N2973 ));
NOR2_X2 _GFM_U485  ( .A1(_GFM_n23910 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3004 ));
NOR2_X2 _GFM_U484  ( .A1(_GFM_n23910 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3035 ));
NOR2_X2 _GFM_U483  ( .A1(_GFM_n23910 ), .A2(_GFM_n26870 ), .ZN(_GFM_N3066 ));
NOR2_X2 _GFM_U482  ( .A1(_GFM_n23900 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3097 ));
NOR2_X2 _GFM_U481  ( .A1(_GFM_n23900 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3128 ));
NOR2_X2 _GFM_U480  ( .A1(_GFM_n23900 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3159 ));
NOR2_X2 _GFM_U478  ( .A1(_GFM_n23900 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3190 ));
NOR2_X2 _GFM_U477  ( .A1(_GFM_n23900 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3221 ));
NOR2_X2 _GFM_U476  ( .A1(_GFM_n23900 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3252 ));
NOR2_X2 _GFM_U475  ( .A1(_GFM_n23900 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3283 ));
NOR2_X2 _GFM_U474  ( .A1(_GFM_n25290 ), .A2(_GFM_n26810 ), .ZN(_GFM_N3289 ));
NOR2_X2 _GFM_U473  ( .A1(_GFM_n25290 ), .A2(_GFM_n26820 ), .ZN(_GFM_N3321 ));
NOR2_X2 _GFM_U472  ( .A1(_GFM_n25290 ), .A2(_GFM_n2683 ), .ZN(_GFM_N3354 ));
NOR2_X2 _GFM_U471  ( .A1(_GFM_n25290 ), .A2(_GFM_n26840 ), .ZN(_GFM_N3388 ));
NOR2_X2 _GFM_U470  ( .A1(_GFM_n25290 ), .A2(_GFM_n2685 ), .ZN(_GFM_N3424 ));
NOR2_X2 _GFM_U469  ( .A1(_GFM_n25290 ), .A2(_GFM_n26860 ), .ZN(_GFM_N3462 ));
NOR2_X2 _GFM_U468  ( .A1(_GFM_n25190 ), .A2(_GFM_n2688 ), .ZN(_GFM_N3502 ));
NOR2_X2 _GFM_U467  ( .A1(_GFM_n25190 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3545 ));
NOR2_X2 _GFM_U466  ( .A1(_GFM_n25190 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3591 ));
NOR2_X2 _GFM_U465  ( .A1(_GFM_n25180 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3640 ));
NOR2_X2 _GFM_U464  ( .A1(_GFM_n25180 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3692 ));
NOR2_X2 _GFM_U463  ( .A1(_GFM_n2528 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3804 ));
NOR2_X2 _GFM_U462  ( .A1(_GFM_n2528 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3865 ));
NOR2_X2 _GFM_U461  ( .A1(_GFM_n26080 ), .A2(_GFM_n25260 ), .ZN(_GFM_N1026 ));
NOR2_X2 _GFM_U460  ( .A1(_GFM_n26070 ), .A2(_GFM_n25360 ), .ZN(_GFM_N1024 ));
NOR2_X2 _GFM_U459  ( .A1(_GFM_n2534 ), .A2(_GFM_n2573 ), .ZN(_GFM_N158 ) );
NOR2_X2 _GFM_U458  ( .A1(_GFM_n2544 ), .A2(_GFM_n25700 ), .ZN(_GFM_N156 ) );
NOR2_X2 _GFM_U457  ( .A1(_GFM_n25320 ), .A2(_GFM_n2578 ), .ZN(_GFM_N220 ) );
NOR2_X2 _GFM_U456  ( .A1(_GFM_n2542 ), .A2(_GFM_n25760 ), .ZN(_GFM_N218 ) );
NOR2_X2 _GFM_U455  ( .A1(_GFM_n25320 ), .A2(_GFM_n25800 ), .ZN(_GFM_N251 ));
NOR2_X2 _GFM_U454  ( .A1(_GFM_n2542 ), .A2(_GFM_n2578 ), .ZN(_GFM_N249 ) );
NOR2_X2 _GFM_U453  ( .A1(_GFM_n2530 ), .A2(_GFM_n25840 ), .ZN(_GFM_N313 ) );
NOR2_X2 _GFM_U452  ( .A1(_GFM_n2540 ), .A2(_GFM_n25821 ), .ZN(_GFM_N311 ) );
NOR2_X2 _GFM_U451  ( .A1(_GFM_n25290 ), .A2(_GFM_n2586 ), .ZN(_GFM_N344 ) );
NOR2_X2 _GFM_U450  ( .A1(_GFM_n25390 ), .A2(_GFM_n25840 ), .ZN(_GFM_N342 ));
NOR2_X2 _GFM_U449  ( .A1(_GFM_n25290 ), .A2(_GFM_n2587 ), .ZN(_GFM_N375 ) );
NOR2_X2 _GFM_U448  ( .A1(_GFM_n25380 ), .A2(_GFM_n2586 ), .ZN(_GFM_N373 ) );
NOR2_X2 _GFM_U447  ( .A1(_GFM_n2547 ), .A2(_GFM_n24770 ), .ZN(_GFM_N3647 ));
NOR2_X2 _GFM_U446  ( .A1(_GFM_n2489 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3648 ));
NOR2_X2 _GFM_U445  ( .A1(_GFM_n25890 ), .A2(_GFM_n25260 ), .ZN(_GFM_N437 ));
NOR2_X2 _GFM_U444  ( .A1(_GFM_n25880 ), .A2(_GFM_n25360 ), .ZN(_GFM_N435 ));
NOR2_X2 _GFM_U443  ( .A1(_GFM_n2554 ), .A2(_GFM_n25260 ), .ZN(_GFM_N3 ) );
NOR2_X2 _GFM_U442  ( .A1(_GFM_n25460 ), .A2(_GFM_n25360 ), .ZN(_GFM_N1 ) );
NOR2_X2 _GFM_U441  ( .A1(_GFM_n25620 ), .A2(_GFM_n25260 ), .ZN(_GFM_N65 ) );
NOR2_X2 _GFM_U440  ( .A1(_GFM_n25580 ), .A2(_GFM_n25360 ), .ZN(_GFM_N63 ) );
NOR2_X2 _GFM_U439  ( .A1(_GFM_n25660 ), .A2(_GFM_n25260 ), .ZN(_GFM_N96 ) );
NOR2_X2 _GFM_U438  ( .A1(_GFM_n25620 ), .A2(_GFM_n25360 ), .ZN(_GFM_N94 ) );
NOR2_X2 _GFM_U437  ( .A1(_GFM_n25180 ), .A2(_GFM_n2554 ), .ZN(_GFM_N4325 ));
NOR2_X2 _GFM_U436  ( .A1(_GFM_n2509 ), .A2(_GFM_n25580 ), .ZN(_GFM_N4329 ));
NOR2_X2 _GFM_U435  ( .A1(_GFM_n25290 ), .A2(_GFM_n25460 ), .ZN(_GFM_N4324 ));
NOR2_X2 _GFM_U434  ( .A1(_GFM_n23880 ), .A2(_GFM_n25880 ), .ZN(_GFM_N4349 ));
NOR2_X2 _GFM_U433  ( .A1(_GFM_n24980 ), .A2(_GFM_n25620 ), .ZN(_GFM_N4328 ));
NOR2_X2 _GFM_U432  ( .A1(_GFM_n25760 ), .A2(_GFM_n24570 ), .ZN(_GFM_N4341 ));
NOR2_X2 _GFM_U431  ( .A1(_GFM_n2578 ), .A2(_GFM_n2447 ), .ZN(_GFM_N4337 ) );
NOR2_X2 _GFM_U430  ( .A1(_GFM_n2573 ), .A2(_GFM_n24670 ), .ZN(_GFM_N4342 ));
NOR2_X2 _GFM_U429  ( .A1(_GFM_n24900 ), .A2(_GFM_n25660 ), .ZN(_GFM_N4331 ));
NOR2_X2 _GFM_U428  ( .A1(_GFM_n25800 ), .A2(_GFM_n2437 ), .ZN(_GFM_N4336 ));
NOR2_X2 _GFM_U427  ( .A1(_GFM_n25821 ), .A2(_GFM_n24260 ), .ZN(_GFM_N4339 ));
NOR2_X2 _GFM_U426  ( .A1(_GFM_n2586 ), .A2(_GFM_n24080 ), .ZN(_GFM_N4345 ));
NOR2_X2 _GFM_U425  ( .A1(_GFM_n25840 ), .A2(_GFM_n25530 ), .ZN(_GFM_N4346 ));
NOR2_X2 _GFM_U424  ( .A1(_GFM_n2587 ), .A2(_GFM_n23970 ), .ZN(_GFM_N4348 ));
NOR2_X2 _GFM_U423  ( .A1(_GFM_n21360 ), .A2(_GFM_n25070 ), .ZN(_GFM_N4108 ));
NOR2_X2 _GFM_U422  ( .A1(_GFM_n26980 ), .A2(_GFM_n2516 ), .ZN(_GFM_N4106 ));
NOR2_X2 _GFM_U421  ( .A1(_GFM_n21360 ), .A2(_GFM_n24960 ), .ZN(_GFM_N4059 ));
INV_X4 _GFM_U420  ( .A(v_out[109]), .ZN(_GFM_n25670 ) );
INV_X4 _GFM_U419  ( .A(v_out[108]), .ZN(_GFM_n25630 ) );
INV_X4 _GFM_U418  ( .A(v_out[107]), .ZN(_GFM_n2559 ) );
INV_X4 _GFM_U417  ( .A(v_out[106]), .ZN(_GFM_n2555 ) );
INV_X4 _GFM_U416  ( .A(v_out[105]), .ZN(_GFM_n2547 ) );
NOR2_X2 _GFM_U415  ( .A1(_GFM_n2696 ), .A2(_GFM_n25260 ), .ZN(_GFM_N4050 ));
NOR2_X2 _GFM_U414  ( .A1(_GFM_n24590 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3484 ));
NOR2_X2 _GFM_U413  ( .A1(_GFM_n2547 ), .A2(_GFM_n25070 ), .ZN(_GFM_N3808 ));
NOR2_X2 _GFM_U412  ( .A1(_GFM_n25180 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3809 ));
NOR2_X2 _GFM_U411  ( .A1(_GFM_n2509 ), .A2(_GFM_n25500 ), .ZN(_GFM_N4167 ));
NOR2_X2 _GFM_U410  ( .A1(_GFM_n21360 ), .A2(_GFM_n2516 ), .ZN(_GFM_N4164 ));
NOR2_X2 _GFM_U409  ( .A1(_GFM_n26980 ), .A2(_GFM_n24960 ), .ZN(_GFM_N4007 ));
NOR2_X2 _GFM_U408  ( .A1(_GFM_n24190 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3338 ));
NOR2_X2 _GFM_U407  ( .A1(_GFM_n24190 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3371 ));
NOR2_X2 _GFM_U406  ( .A1(_GFM_n2480 ), .A2(_GFM_n2689 ), .ZN(_GFM_N3397 ) );
NOR2_X2 _GFM_U405  ( .A1(_GFM_n2499 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3511 ));
NOR2_X2 _GFM_U404  ( .A1(_GFM_n2559 ), .A2(_GFM_n23970 ), .ZN(_GFM_N3413 ));
NOR2_X2 _GFM_U403  ( .A1(_GFM_n24590 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3409 ));
NOR2_X2 _GFM_U402  ( .A1(_GFM_n25630 ), .A2(_GFM_n23970 ), .ZN(_GFM_N3450 ));
NOR2_X2 _GFM_U401  ( .A1(_GFM_n24590 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3446 ));
NOR2_X2 _GFM_U400  ( .A1(_GFM_n2528 ), .A2(_GFM_n2606 ), .ZN(_GFM_N964 ) );
NOR2_X2 _GFM_U399  ( .A1(_GFM_n2537 ), .A2(_GFM_n26050 ), .ZN(_GFM_N962 ) );
NOR2_X2 _GFM_U398  ( .A1(_GFM_n2537 ), .A2(_GFM_n2609 ), .ZN(_GFM_N1086 ) );
NOR2_X2 _GFM_U397  ( .A1(_GFM_n2610 ), .A2(_GFM_n25260 ), .ZN(_GFM_N1088 ));
NOR2_X2 _GFM_U396  ( .A1(_GFM_n25350 ), .A2(_GFM_n26110 ), .ZN(_GFM_N1119 ));
NOR2_X2 _GFM_U395  ( .A1(_GFM_n2610 ), .A2(_GFM_n25360 ), .ZN(_GFM_N1117 ));
NOR2_X2 _GFM_U394  ( .A1(_GFM_n25350 ), .A2(_GFM_n2613 ), .ZN(_GFM_N1181 ));
NOR2_X2 _GFM_U393  ( .A1(_GFM_n25450 ), .A2(_GFM_n26120 ), .ZN(_GFM_N1179 ));
NOR2_X2 _GFM_U392  ( .A1(_GFM_n25350 ), .A2(_GFM_n26140 ), .ZN(_GFM_N1212 ));
NOR2_X2 _GFM_U391  ( .A1(_GFM_n25450 ), .A2(_GFM_n2613 ), .ZN(_GFM_N1210 ));
NOR2_X2 _GFM_U390  ( .A1(_GFM_n25350 ), .A2(_GFM_n2618 ), .ZN(_GFM_N1336 ));
NOR2_X2 _GFM_U387  ( .A1(_GFM_n25450 ), .A2(_GFM_n2617 ), .ZN(_GFM_N1334 ));
NOR2_X2 _GFM_U385  ( .A1(_GFM_n25350 ), .A2(_GFM_n26190 ), .ZN(_GFM_N1367 ));
NOR2_X2 _GFM_U383  ( .A1(_GFM_n25450 ), .A2(_GFM_n2618 ), .ZN(_GFM_N1365 ));
NOR2_X2 _GFM_U382  ( .A1(_GFM_n2530 ), .A2(_GFM_n2672 ), .ZN(_GFM_N3010 ) );
NOR2_X2 _GFM_U380  ( .A1(_GFM_n2540 ), .A2(_GFM_n2671 ), .ZN(_GFM_N3008 ) );
NOR2_X2 _GFM_U378  ( .A1(_GFM_n2530 ), .A2(_GFM_n26730 ), .ZN(_GFM_N3041 ));
NOR2_X2 _GFM_U376  ( .A1(_GFM_n2540 ), .A2(_GFM_n2672 ), .ZN(_GFM_N3039 ) );
NOR2_X2 _GFM_U374  ( .A1(_GFM_n2530 ), .A2(_GFM_n26740 ), .ZN(_GFM_N3072 ));
NOR2_X2 _GFM_U372  ( .A1(_GFM_n2540 ), .A2(_GFM_n26730 ), .ZN(_GFM_N3070 ));
NOR2_X2 _GFM_U370  ( .A1(_GFM_n2530 ), .A2(_GFM_n2675 ), .ZN(_GFM_N3103 ) );
NOR2_X2 _GFM_U368  ( .A1(_GFM_n2540 ), .A2(_GFM_n26740 ), .ZN(_GFM_N3101 ));
NOR2_X2 _GFM_U366  ( .A1(_GFM_n2530 ), .A2(_GFM_n26760 ), .ZN(_GFM_N3134 ));
NOR2_X2 _GFM_U364  ( .A1(_GFM_n2540 ), .A2(_GFM_n2675 ), .ZN(_GFM_N3132 ) );
NOR2_X2 _GFM_U362  ( .A1(_GFM_n2530 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3165 ));
NOR2_X2 _GFM_U360  ( .A1(_GFM_n2540 ), .A2(_GFM_n26760 ), .ZN(_GFM_N3163 ));
NOR2_X2 _GFM_U358  ( .A1(_GFM_n25290 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3196 ));
NOR2_X2 _GFM_U357  ( .A1(_GFM_n2540 ), .A2(_GFM_n26770 ), .ZN(_GFM_N3194 ));
NOR2_X2 _GFM_U355  ( .A1(_GFM_n25290 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3227 ));
NOR2_X2 _GFM_U353  ( .A1(_GFM_n25390 ), .A2(_GFM_n2678 ), .ZN(_GFM_N3225 ));
NOR2_X2 _GFM_U351  ( .A1(_GFM_n2530 ), .A2(_GFM_n26801 ), .ZN(_GFM_N3258 ));
NOR2_X2 _GFM_U349  ( .A1(_GFM_n25390 ), .A2(_GFM_n2679 ), .ZN(_GFM_N3256 ));
NOR2_X2 _GFM_U347  ( .A1(_GFM_n21360 ), .A2(_GFM_n25260 ), .ZN(_GFM_N4221 ));
NOR2_X2 _GFM_U345  ( .A1(_GFM_n26980 ), .A2(_GFM_n2537 ), .ZN(_GFM_N4218 ));
NOR2_X2 _GFM_U343  ( .A1(_GFM_n2479 ), .A2(_GFM_n26900 ), .ZN(_GFM_N3433 ));
NOR2_X2 _GFM_U341  ( .A1(_GFM_n2479 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3471 ));
NOR2_X2 _GFM_U340  ( .A1(_GFM_n2499 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3600 ));
NOR2_X2 _GFM_U338  ( .A1(_GFM_n24980 ), .A2(_GFM_n26930 ), .ZN(_GFM_N3649 ));
NOR2_X2 _GFM_U336  ( .A1(_GFM_n24980 ), .A2(_GFM_n26940 ), .ZN(_GFM_N3703 ));
NOR2_X2 _GFM_U334  ( .A1(_GFM_n2499 ), .A2(_GFM_n26910 ), .ZN(_GFM_N3554 ));
NOR2_X2 _GFM_U332  ( .A1(_GFM_n2528 ), .A2(_GFM_n26921 ), .ZN(_GFM_N3748 ));
NOR2_X2 _GFM_U330  ( .A1(_GFM_n2533 ), .A2(_GFM_n25760 ), .ZN(_GFM_N189 ) );
NOR2_X2 _GFM_U328  ( .A1(_GFM_n25430 ), .A2(_GFM_n2573 ), .ZN(_GFM_N187 ) );
NOR2_X2 _GFM_U326  ( .A1(_GFM_n25310 ), .A2(_GFM_n25821 ), .ZN(_GFM_N282 ));
NOR2_X2 _GFM_U324  ( .A1(_GFM_n2541 ), .A2(_GFM_n25800 ), .ZN(_GFM_N280 ) );
NOR2_X2 _GFM_U323  ( .A1(_GFM_n25380 ), .A2(_GFM_n2587 ), .ZN(_GFM_N404 ) );
NOR2_X2 _GFM_U322  ( .A1(_GFM_n25880 ), .A2(_GFM_n25260 ), .ZN(_GFM_N406 ));
NOR2_X2 _GFM_U321  ( .A1(_GFM_n2554 ), .A2(_GFM_n2537 ), .ZN(_GFM_N32 ) );
NOR2_X2 _GFM_U320  ( .A1(_GFM_n25580 ), .A2(_GFM_n25260 ), .ZN(_GFM_N34 ) );
NOR2_X2 _GFM_U319  ( .A1(_GFM_n25350 ), .A2(_GFM_n25700 ), .ZN(_GFM_N127 ));
NOR2_X2 _GFM_U318  ( .A1(_GFM_n25660 ), .A2(_GFM_n25360 ), .ZN(_GFM_N125 ));
INV_X4 _GFM_U317  ( .A(v_out[111]), .ZN(_GFM_n25511 ) );
INV_X4 _GFM_U316  ( .A(v_out[110]), .ZN(_GFM_n25520 ) );
NOR2_X2 _GFM_U315  ( .A1(_GFM_n2399 ), .A2(_GFM_n2585 ), .ZN(_GFM_N4269 ) );
NOR2_X2 _GFM_U314  ( .A1(_GFM_n2399 ), .A2(_GFM_n25830 ), .ZN(_GFM_N4210 ));
NOR2_X2 _GFM_U313  ( .A1(_GFM_n2389 ), .A2(_GFM_n2575 ), .ZN(_GFM_N3923 ) );
NOR2_X2 _GFM_U312  ( .A1(_GFM_n2389 ), .A2(_GFM_n2585 ), .ZN(_GFM_N4213 ) );
NOR2_X2 _GFM_U311  ( .A1(_GFM_n2409 ), .A2(_GFM_n25690 ), .ZN(_GFM_N3918 ));
NOR2_X2 _GFM_U310  ( .A1(_GFM_n2418 ), .A2(_GFM_n25690 ), .ZN(_GFM_N3966 ));
NOR2_X2 _GFM_U309  ( .A1(_GFM_n2399 ), .A2(_GFM_n25810 ), .ZN(_GFM_N4151 ));
NOR2_X2 _GFM_U308  ( .A1(_GFM_n2409 ), .A2(_GFM_n25810 ), .ZN(_GFM_N4203 ));
NOR2_X2 _GFM_U307  ( .A1(_GFM_n2389 ), .A2(_GFM_n25830 ), .ZN(_GFM_N4154 ));
NOR2_X2 _GFM_U306  ( .A1(_GFM_n2389 ), .A2(_GFM_n2572 ), .ZN(_GFM_N3859 ) );
NOR2_X2 _GFM_U305  ( .A1(_GFM_n2399 ), .A2(_GFM_n2572 ), .ZN(_GFM_N3914 ) );
NOR2_X2 _GFM_U304  ( .A1(_GFM_n2409 ), .A2(_GFM_n2565 ), .ZN(_GFM_N3854 ) );
NOR2_X2 _GFM_U303  ( .A1(_GFM_n24190 ), .A2(_GFM_n2565 ), .ZN(_GFM_N3899 ));
NOR2_X2 _GFM_U302  ( .A1(_GFM_n2399 ), .A2(_GFM_n2579 ), .ZN(_GFM_N4094 ) );
NOR2_X2 _GFM_U301  ( .A1(_GFM_n2389 ), .A2(_GFM_n25810 ), .ZN(_GFM_N4097 ));
NOR2_X2 _GFM_U300  ( .A1(_GFM_n2489 ), .A2(_GFM_n2548 ), .ZN(_GFM_N4113 ) );
NOR2_X2 _GFM_U299  ( .A1(_GFM_n24980 ), .A2(_GFM_n25500 ), .ZN(_GFM_N4116 ));
NOR2_X2 _GFM_U298  ( .A1(_GFM_n24880 ), .A2(_GFM_n2556 ), .ZN(_GFM_N4172 ));
NOR2_X2 _GFM_U297  ( .A1(_GFM_n24980 ), .A2(_GFM_n2548 ), .ZN(_GFM_N4175 ));
NOR2_X2 _GFM_U296  ( .A1(_GFM_n2489 ), .A2(_GFM_n25600 ), .ZN(_GFM_N4233 ));
NOR2_X2 _GFM_U295  ( .A1(_GFM_n24980 ), .A2(_GFM_n2556 ), .ZN(_GFM_N4236 ));
NOR2_X2 _GFM_U294  ( .A1(_GFM_n24380 ), .A2(_GFM_n2564 ), .ZN(_GFM_N4017 ));
NOR2_X2 _GFM_U293  ( .A1(_GFM_n2400 ), .A2(_GFM_n25770 ), .ZN(_GFM_N4039 ));
NOR2_X2 _GFM_U292  ( .A1(_GFM_n2449 ), .A2(_GFM_n25600 ), .ZN(_GFM_N4024 ));
NOR2_X2 _GFM_U291  ( .A1(_GFM_n2409 ), .A2(_GFM_n25740 ), .ZN(_GFM_N4032 ));
NOR2_X2 _GFM_U290  ( .A1(_GFM_n2449 ), .A2(_GFM_n2564 ), .ZN(_GFM_N4079 ) );
NOR2_X2 _GFM_U289  ( .A1(_GFM_n24101 ), .A2(_GFM_n25770 ), .ZN(_GFM_N4087 ));
NOR2_X2 _GFM_U288  ( .A1(_GFM_n2478 ), .A2(_GFM_n2548 ), .ZN(_GFM_N4063 ) );
NOR2_X2 _GFM_U287  ( .A1(_GFM_n24390 ), .A2(_GFM_n2568 ), .ZN(_GFM_N4072 ));
NOR2_X2 _GFM_U286  ( .A1(_GFM_n2479 ), .A2(_GFM_n2556 ), .ZN(_GFM_N4120 ) );
NOR2_X2 _GFM_U285  ( .A1(_GFM_n24390 ), .A2(_GFM_n2571 ), .ZN(_GFM_N4129 ));
NOR2_X2 _GFM_U284  ( .A1(_GFM_n2448 ), .A2(_GFM_n2568 ), .ZN(_GFM_N4136 ) );
NOR2_X2 _GFM_U283  ( .A1(_GFM_n2409 ), .A2(_GFM_n2579 ), .ZN(_GFM_N4144 ) );
NOR2_X2 _GFM_U282  ( .A1(_GFM_n24380 ), .A2(_GFM_n25740 ), .ZN(_GFM_N4188 ));
NOR2_X2 _GFM_U281  ( .A1(_GFM_n2448 ), .A2(_GFM_n2571 ), .ZN(_GFM_N4195 ) );
NOR2_X2 _GFM_U280  ( .A1(_GFM_n24380 ), .A2(_GFM_n25770 ), .ZN(_GFM_N4249 ));
NOR2_X2 _GFM_U279  ( .A1(_GFM_n2449 ), .A2(_GFM_n25740 ), .ZN(_GFM_N4255 ));
NOR2_X2 _GFM_U278  ( .A1(_GFM_n25180 ), .A2(_GFM_n25500 ), .ZN(_GFM_N4225 ));
NOR2_X2 _GFM_U277  ( .A1(_GFM_n2509 ), .A2(_GFM_n2548 ), .ZN(_GFM_N4228 ) );
NOR2_X2 _GFM_U276  ( .A1(_GFM_n2489 ), .A2(_GFM_n25500 ), .ZN(_GFM_N4057 ));
NOR2_X2 _GFM_U275  ( .A1(_GFM_n2418 ), .A2(_GFM_n25810 ), .ZN(_GFM_N4265 ));
NOR2_X2 _GFM_U274  ( .A1(_GFM_n2400 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3580 ));
NOR2_X2 _GFM_U273  ( .A1(_GFM_n24101 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3615 ));
NOR2_X2 _GFM_U272  ( .A1(_GFM_n2449 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3844 ));
NOR2_X2 _GFM_U271  ( .A1(_GFM_n24590 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3889 ));
NOR2_X2 _GFM_U270  ( .A1(_GFM_n2418 ), .A2(_GFM_n25611 ), .ZN(_GFM_N3835 ));
NOR2_X2 _GFM_U269  ( .A1(_GFM_n2400 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3534 ));
NOR2_X2 _GFM_U268  ( .A1(_GFM_n24101 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3566 ));
NOR2_X2 _GFM_U267  ( .A1(_GFM_n2449 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3783 ));
NOR2_X2 _GFM_U266  ( .A1(_GFM_n2458 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3825 ));
NOR2_X2 _GFM_U265  ( .A1(_GFM_n2389 ), .A2(_GFM_n2565 ), .ZN(_GFM_N3740 ) );
NOR2_X2 _GFM_U264  ( .A1(_GFM_n2399 ), .A2(_GFM_n2565 ), .ZN(_GFM_N3789 ) );
NOR2_X2 _GFM_U263  ( .A1(_GFM_n24290 ), .A2(_GFM_n2565 ), .ZN(_GFM_N3962 ));
NOR2_X2 _GFM_U262  ( .A1(_GFM_n2400 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3681 ));
NOR2_X2 _GFM_U261  ( .A1(_GFM_n2409 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3735 ));
NOR2_X2 _GFM_U260  ( .A1(_GFM_n2448 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3975 ));
NOR2_X2 _GFM_U259  ( .A1(_GFM_n24690 ), .A2(_GFM_n2548 ), .ZN(_GFM_N4012 ));
NOR2_X2 _GFM_U258  ( .A1(_GFM_n24280 ), .A2(_GFM_n2568 ), .ZN(_GFM_N4020 ));
NOR2_X2 _GFM_U257  ( .A1(_GFM_n23900 ), .A2(_GFM_n2579 ), .ZN(_GFM_N4042 ));
NOR2_X2 _GFM_U256  ( .A1(_GFM_n24190 ), .A2(_GFM_n2571 ), .ZN(_GFM_N4035 ));
NOR2_X2 _GFM_U255  ( .A1(_GFM_n2418 ), .A2(_GFM_n25740 ), .ZN(_GFM_N4090 ));
NOR2_X2 _GFM_U254  ( .A1(_GFM_n24280 ), .A2(_GFM_n2571 ), .ZN(_GFM_N4075 ));
NOR2_X2 _GFM_U253  ( .A1(_GFM_n24290 ), .A2(_GFM_n25740 ), .ZN(_GFM_N4132 ));
NOR2_X2 _GFM_U252  ( .A1(_GFM_n2418 ), .A2(_GFM_n25770 ), .ZN(_GFM_N4147 ));
NOR2_X2 _GFM_U251  ( .A1(_GFM_n2468 ), .A2(_GFM_n2564 ), .ZN(_GFM_N4182 ) );
NOR2_X2 _GFM_U250  ( .A1(_GFM_n24280 ), .A2(_GFM_n25770 ), .ZN(_GFM_N4191 ));
NOR2_X2 _GFM_U249  ( .A1(_GFM_n2418 ), .A2(_GFM_n2579 ), .ZN(_GFM_N4206 ) );
NOR2_X2 _GFM_U248  ( .A1(_GFM_n24690 ), .A2(_GFM_n2568 ), .ZN(_GFM_N4243 ));
NOR2_X2 _GFM_U247  ( .A1(_GFM_n24280 ), .A2(_GFM_n2579 ), .ZN(_GFM_N4251 ));
NOR2_X2 _GFM_U246  ( .A1(_GFM_n24590 ), .A2(_GFM_n2571 ), .ZN(_GFM_N4258 ));
NOR2_X2 _GFM_U245  ( .A1(_GFM_n23900 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3538 ));
NOR2_X2 _GFM_U244  ( .A1(_GFM_n24190 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3662 ));
NOR2_X2 _GFM_U243  ( .A1(_GFM_n24290 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3715 ));
NOR2_X2 _GFM_U242  ( .A1(_GFM_n24390 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3780 ));
NOR2_X2 _GFM_U241  ( .A1(_GFM_n2468 ), .A2(_GFM_n25511 ), .ZN(_GFM_N3951 ));
NOR2_X2 _GFM_U240  ( .A1(_GFM_n2389 ), .A2(_GFM_n25611 ), .ZN(_GFM_N3685 ));
NOR2_X2 _GFM_U239  ( .A1(_GFM_n2400 ), .A2(_GFM_n25611 ), .ZN(_GFM_N3731 ));
NOR2_X2 _GFM_U238  ( .A1(_GFM_n24290 ), .A2(_GFM_n25611 ), .ZN(_GFM_N3895 ));
NOR2_X2 _GFM_U237  ( .A1(_GFM_n24390 ), .A2(_GFM_n25611 ), .ZN(_GFM_N3971 ));
NOR2_X2 _GFM_U236  ( .A1(_GFM_n23900 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3495 ));
NOR2_X2 _GFM_U235  ( .A1(_GFM_n24190 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3611 ));
NOR2_X2 _GFM_U234  ( .A1(_GFM_n24290 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3670 ));
NOR2_X2 _GFM_U233  ( .A1(_GFM_n24390 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3723 ));
NOR2_X2 _GFM_U232  ( .A1(_GFM_n2479 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3944 ));
NOR2_X2 _GFM_U231  ( .A1(_GFM_n2400 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3629 ));
NOR2_X2 _GFM_U230  ( .A1(_GFM_n24101 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3666 ));
NOR2_X2 _GFM_U229  ( .A1(_GFM_n2418 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3719 ));
NOR2_X2 _GFM_U228  ( .A1(_GFM_n2449 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3908 ));
NOR2_X2 _GFM_U227  ( .A1(_GFM_n24590 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3955 ));
NOR2_X2 _GFM_U226  ( .A1(_GFM_n23900 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3633 ));
NOR2_X2 _GFM_U225  ( .A1(_GFM_n24290 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3831 ));
NOR2_X2 _GFM_U224  ( .A1(_GFM_n25670 ), .A2(_GFM_n24260 ), .ZN(_GFM_N3620 ));
NOR2_X2 _GFM_U223  ( .A1(_GFM_n25670 ), .A2(_GFM_n2437 ), .ZN(_GFM_N3672 ));
NOR2_X2 _GFM_U222  ( .A1(_GFM_n25670 ), .A2(_GFM_n24560 ), .ZN(_GFM_N3764 ));
NOR2_X2 _GFM_U221  ( .A1(_GFM_n25670 ), .A2(_GFM_n24670 ), .ZN(_GFM_N3818 ));
NOR2_X2 _GFM_U220  ( .A1(_GFM_n25670 ), .A2(_GFM_n24770 ), .ZN(_GFM_N3881 ));
NOR2_X2 _GFM_U219  ( .A1(_GFM_n2389 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3584 ));
NOR2_X2 _GFM_U218  ( .A1(_GFM_n24290 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3771 ));
NOR2_X2 _GFM_U217  ( .A1(_GFM_n24390 ), .A2(_GFM_n25490 ), .ZN(_GFM_N3840 ));
NOR2_X2 _GFM_U216  ( .A1(_GFM_n25630 ), .A2(_GFM_n24080 ), .ZN(_GFM_N3491 ));
NOR2_X2 _GFM_U215  ( .A1(_GFM_n25630 ), .A2(_GFM_n24570 ), .ZN(_GFM_N3708 ));
NOR2_X2 _GFM_U214  ( .A1(_GFM_n25630 ), .A2(_GFM_n24960 ), .ZN(_GFM_N3939 ));
NOR2_X2 _GFM_U213  ( .A1(_GFM_n2559 ), .A2(_GFM_n24070 ), .ZN(_GFM_N3452 ));
NOR2_X2 _GFM_U212  ( .A1(_GFM_n2559 ), .A2(_GFM_n2427 ), .ZN(_GFM_N3521 ) );
NOR2_X2 _GFM_U211  ( .A1(_GFM_n2559 ), .A2(_GFM_n24560 ), .ZN(_GFM_N3655 ));
NOR2_X2 _GFM_U210  ( .A1(_GFM_n25670 ), .A2(_GFM_n2387 ), .ZN(_GFM_N3455 ));
NOR2_X2 _GFM_U209  ( .A1(_GFM_n25670 ), .A2(_GFM_n23970 ), .ZN(_GFM_N3489 ));
NOR2_X2 _GFM_U208  ( .A1(_GFM_n25670 ), .A2(_GFM_n25530 ), .ZN(_GFM_N3563 ));
NOR2_X2 _GFM_U207  ( .A1(_GFM_n2555 ), .A2(_GFM_n24080 ), .ZN(_GFM_N3415 ));
NOR2_X2 _GFM_U206  ( .A1(_GFM_n2555 ), .A2(_GFM_n2427 ), .ZN(_GFM_N3477 ) );
NOR2_X2 _GFM_U205  ( .A1(_GFM_n2555 ), .A2(_GFM_n2437 ), .ZN(_GFM_N3527 ) );
NOR2_X2 _GFM_U204  ( .A1(_GFM_n2555 ), .A2(_GFM_n24560 ), .ZN(_GFM_N3605 ));
NOR2_X2 _GFM_U203  ( .A1(_GFM_n2555 ), .A2(_GFM_n24870 ), .ZN(_GFM_N3754 ));
NOR2_X2 _GFM_U202  ( .A1(_GFM_n25630 ), .A2(_GFM_n2387 ), .ZN(_GFM_N3418 ));
NOR2_X2 _GFM_U201  ( .A1(_GFM_n25630 ), .A2(_GFM_n25530 ), .ZN(_GFM_N3519 ));
NOR2_X2 _GFM_U200  ( .A1(_GFM_n25630 ), .A2(_GFM_n2437 ), .ZN(_GFM_N3618 ));
NOR2_X2 _GFM_U199  ( .A1(_GFM_n2559 ), .A2(_GFM_n2387 ), .ZN(_GFM_N3383 ) );
NOR2_X2 _GFM_U198  ( .A1(_GFM_n2559 ), .A2(_GFM_n2417 ), .ZN(_GFM_N3479 ) );
NOR2_X2 _GFM_U197  ( .A1(_GFM_n2559 ), .A2(_GFM_n2437 ), .ZN(_GFM_N3569 ) );
NOR2_X2 _GFM_U196  ( .A1(_GFM_n2559 ), .A2(_GFM_n24670 ), .ZN(_GFM_N3706 ));
NOR2_X2 _GFM_U195  ( .A1(_GFM_n2559 ), .A2(_GFM_n24770 ), .ZN(_GFM_N3756 ));
NOR2_X2 _GFM_U194  ( .A1(_GFM_n2547 ), .A2(_GFM_n24870 ), .ZN(_GFM_N3699 ));
NOR2_X2 _GFM_U193  ( .A1(_GFM_n2555 ), .A2(_GFM_n24770 ), .ZN(_GFM_N3701 ));
NOR2_X2 _GFM_U192  ( .A1(_GFM_n2547 ), .A2(_GFM_n24070 ), .ZN(_GFM_N3380 ));
NOR2_X2 _GFM_U191  ( .A1(_GFM_n2547 ), .A2(_GFM_n24260 ), .ZN(_GFM_N3439 ));
NOR2_X2 _GFM_U190  ( .A1(_GFM_n2547 ), .A2(_GFM_n2437 ), .ZN(_GFM_N3482 ) );
NOR2_X2 _GFM_U189  ( .A1(_GFM_n2547 ), .A2(_GFM_n24570 ), .ZN(_GFM_N3558 ));
NOR2_X2 _GFM_U188  ( .A1(_GFM_n2547 ), .A2(_GFM_n24960 ), .ZN(_GFM_N3759 ));
NOR2_X2 _GFM_U187  ( .A1(_GFM_n2555 ), .A2(_GFM_n2387 ), .ZN(_GFM_N3349 ) );
NOR2_X2 _GFM_U186  ( .A1(_GFM_n2555 ), .A2(_GFM_n23970 ), .ZN(_GFM_N3378 ));
NOR2_X2 _GFM_U185  ( .A1(_GFM_n2555 ), .A2(_GFM_n25530 ), .ZN(_GFM_N3441 ));
NOR2_X2 _GFM_U184  ( .A1(_GFM_n2555 ), .A2(_GFM_n24460 ), .ZN(_GFM_N3574 ));
NOR2_X2 _GFM_U183  ( .A1(_GFM_n2555 ), .A2(_GFM_n2466 ), .ZN(_GFM_N3653 ) );
NOR2_X2 _GFM_U182  ( .A1(_GFM_n2555 ), .A2(_GFM_n2516 ), .ZN(_GFM_N3936 ) );
NOR2_X2 _GFM_U181  ( .A1(_GFM_n2547 ), .A2(_GFM_n2387 ), .ZN(_GFM_N3316 ) );
NOR2_X2 _GFM_U180  ( .A1(_GFM_n2547 ), .A2(_GFM_n23970 ), .ZN(_GFM_N3345 ));
NOR2_X2 _GFM_U179  ( .A1(_GFM_n2547 ), .A2(_GFM_n2417 ), .ZN(_GFM_N3404 ) );
NOR2_X2 _GFM_U178  ( .A1(_GFM_n2547 ), .A2(_GFM_n2447 ), .ZN(_GFM_N3529 ) );
NOR2_X2 _GFM_U177  ( .A1(_GFM_n2547 ), .A2(_GFM_n2466 ), .ZN(_GFM_N3603 ) );
NOR2_X2 _GFM_U176  ( .A1(_GFM_n25670 ), .A2(_GFM_n24070 ), .ZN(_GFM_N3524 ));
NOR2_X2 _GFM_U175  ( .A1(_GFM_n25630 ), .A2(_GFM_n2447 ), .ZN(_GFM_N3674 ));
NOR2_X2 _GFM_U174  ( .A1(_GFM_n25670 ), .A2(_GFM_n2447 ), .ZN(_GFM_N3725 ));
NOR2_X2 _GFM_U173  ( .A1(_GFM_n24380 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3904 ));
NOR2_X2 _GFM_U172  ( .A1(_GFM_n2409 ), .A2(_GFM_n25830 ), .ZN(_GFM_N4263 ));
NOR2_X2 _GFM_U171  ( .A1(_GFM_n2399 ), .A2(_GFM_n2575 ), .ZN(_GFM_N3981 ) );
NOR2_X2 _GFM_U170  ( .A1(_GFM_n25630 ), .A2(_GFM_n2427 ), .ZN(_GFM_N3571 ));
NOR2_X2 _GFM_U169  ( .A1(_GFM_n2559 ), .A2(_GFM_n2447 ), .ZN(_GFM_N3623 ) );
NOR2_X2 _GFM_U168  ( .A1(_GFM_n2399 ), .A2(_GFM_n25690 ), .ZN(_GFM_N3850 ));
NOR2_X2 _GFM_U167  ( .A1(_GFM_n2389 ), .A2(_GFM_n25690 ), .ZN(_GFM_N3798 ));
NOR2_X2 _GFM_U166  ( .A1(_GFM_n24101 ), .A2(_GFM_n25611 ), .ZN(_GFM_N3793 ));
NOR2_X2 _GFM_U165  ( .A1(_GFM_n2547 ), .A2(_GFM_n2516 ), .ZN(_GFM_N3871 ) );
NOR2_X2 _GFM_U164  ( .A1(_GFM_n2555 ), .A2(_GFM_n25080 ), .ZN(_GFM_N3869 ));
NOR2_X2 _GFM_U163  ( .A1(_GFM_n25670 ), .A2(_GFM_n24870 ), .ZN(_GFM_N3946 ));
NOR2_X2 _GFM_U162  ( .A1(_GFM_n24190 ), .A2(_GFM_n25570 ), .ZN(_GFM_N3775 ));
NOR2_X2 _GFM_U161  ( .A1(_GFM_n2559 ), .A2(_GFM_n24870 ), .ZN(_GFM_N3821 ));
NOR2_X2 _GFM_U160  ( .A1(_GFM_n25630 ), .A2(_GFM_n24870 ), .ZN(_GFM_N3883 ));
NOR2_X2 _GFM_U159  ( .A1(_GFM_n24590 ), .A2(_GFM_n2556 ), .ZN(_GFM_N4027 ));
NOR2_X2 _GFM_U158  ( .A1(_GFM_n24590 ), .A2(_GFM_n25600 ), .ZN(_GFM_N4082 ));
NOR2_X2 _GFM_U157  ( .A1(_GFM_n2468 ), .A2(_GFM_n2556 ), .ZN(_GFM_N4066 ) );
NOR2_X2 _GFM_U156  ( .A1(_GFM_n2468 ), .A2(_GFM_n25600 ), .ZN(_GFM_N4123 ));
NOR2_X2 _GFM_U155  ( .A1(_GFM_n2458 ), .A2(_GFM_n2564 ), .ZN(_GFM_N4139 ) );
NOR2_X2 _GFM_U154  ( .A1(_GFM_n2478 ), .A2(_GFM_n25600 ), .ZN(_GFM_N4179 ));
NOR2_X2 _GFM_U153  ( .A1(_GFM_n2458 ), .A2(_GFM_n2568 ), .ZN(_GFM_N4198 ) );
NOR2_X2 _GFM_U152  ( .A1(_GFM_n2478 ), .A2(_GFM_n2564 ), .ZN(_GFM_N4240 ) );
NOR2_X2 _GFM_U151  ( .A1(_GFM_n25630 ), .A2(_GFM_n2466 ), .ZN(_GFM_N3762 ));
NOR2_X2 _GFM_U150  ( .A1(_GFM_n2559 ), .A2(_GFM_n25070 ), .ZN(_GFM_N3934 ));
NOR2_X2 _GFM_U149  ( .A1(_GFM_n2555 ), .A2(_GFM_n24960 ), .ZN(_GFM_N3812 ));
NOR2_X2 _GFM_U148  ( .A1(_GFM_n25630 ), .A2(_GFM_n24770 ), .ZN(_GFM_N3816 ));
NOR2_X2 _GFM_U147  ( .A1(_GFM_n2468 ), .A2(_GFM_n25520 ), .ZN(_GFM_N3879 ));
NOR2_X2 _GFM_U146  ( .A1(_GFM_n2559 ), .A2(_GFM_n24960 ), .ZN(_GFM_N3874 ));
INV_X4 _GFM_U145  ( .A(b_in[112]), .ZN(_GFM_n2396 ) );
INV_X4 _GFM_U144  ( .A(b_in[114]), .ZN(_GFM_n2416 ) );
INV_X4 _GFM_U143  ( .A(b_in[120]), .ZN(_GFM_n2475 ) );
INV_X4 _GFM_U142  ( .A(b_in[113]), .ZN(_GFM_n2406 ) );
INV_X4 _GFM_U141  ( .A(b_in[125]), .ZN(_GFM_n2525 ) );
INV_X4 _GFM_U140  ( .A(b_in[123]), .ZN(_GFM_n25050 ) );
INV_X4 _GFM_U139  ( .A(b_in[115]), .ZN(_GFM_n24250 ) );
INV_X4 _GFM_U138  ( .A(b_in[121]), .ZN(_GFM_n2485 ) );
INV_X4 _GFM_U137  ( .A(b_in[117]), .ZN(_GFM_n24450 ) );
INV_X4 _GFM_U136  ( .A(b_in[118]), .ZN(_GFM_n2455 ) );
INV_X4 _GFM_U135  ( .A(b_in[122]), .ZN(_GFM_n24950 ) );
INV_X4 _GFM_U134  ( .A(b_in[119]), .ZN(_GFM_n24650 ) );
INV_X4 _GFM_U133  ( .A(b_in[124]), .ZN(_GFM_n25150 ) );
INV_X4 _GFM_U132  ( .A(b_in[116]), .ZN(_GFM_n2435 ) );
INV_X4 _GFM_U131  ( .A(b_in[116]), .ZN(_GFM_n2427 ) );
INV_X4 _GFM_U130  ( .A(b_in[121]), .ZN(_GFM_n24770 ) );
INV_X4 _GFM_U129  ( .A(b_in[122]), .ZN(_GFM_n24870 ) );
INV_X4 _GFM_U128  ( .A(b_in[124]), .ZN(_GFM_n25070 ) );
INV_X4 _GFM_U127  ( .A(b_in[118]), .ZN(_GFM_n2454 ) );
INV_X4 _GFM_U126  ( .A(b_in[116]), .ZN(_GFM_n24340 ) );
INV_X4 _GFM_U125  ( .A(b_in[122]), .ZN(_GFM_n24880 ) );
INV_X4 _GFM_U124  ( .A(b_in[119]), .ZN(_GFM_n2463 ) );
INV_X4 _GFM_U123  ( .A(b_in[120]), .ZN(_GFM_n24730 ) );
INV_X4 _GFM_U122  ( .A(b_in[114]), .ZN(_GFM_n2413 ) );
INV_X4 _GFM_U121  ( .A(b_in[115]), .ZN(_GFM_n24220 ) );
INV_X4 _GFM_U120  ( .A(b_in[121]), .ZN(_GFM_n2478 ) );
INV_X4 _GFM_U119  ( .A(b_in[117]), .ZN(_GFM_n24380 ) );
INV_X4 _GFM_U118  ( .A(b_in[118]), .ZN(_GFM_n2448 ) );
INV_X4 _GFM_U117  ( .A(b_in[116]), .ZN(_GFM_n24280 ) );
INV_X4 _GFM_U116  ( .A(b_in[122]), .ZN(_GFM_n2489 ) );
INV_X4 _GFM_U115  ( .A(b_in[119]), .ZN(_GFM_n2458 ) );
INV_X4 _GFM_U114  ( .A(b_in[120]), .ZN(_GFM_n2468 ) );
INV_X4 _GFM_U113  ( .A(b_in[115]), .ZN(_GFM_n2418 ) );
INV_X4 _GFM_U112  ( .A(b_in[123]), .ZN(_GFM_n2497 ) );
INV_X4 _GFM_U111  ( .A(b_in[121]), .ZN(_GFM_n2479 ) );
INV_X4 _GFM_U110  ( .A(b_in[125]), .ZN(_GFM_n2517 ) );
INV_X4 _GFM_U109  ( .A(b_in[114]), .ZN(_GFM_n24150 ) );
INV_X4 _GFM_U108  ( .A(b_in[115]), .ZN(_GFM_n2424 ) );
INV_X4 _GFM_U107  ( .A(b_in[120]), .ZN(_GFM_n24740 ) );
INV_X4 _GFM_U106  ( .A(b_in[113]), .ZN(_GFM_n24050 ) );
INV_X4 _GFM_U105  ( .A(b_in[121]), .ZN(_GFM_n24840 ) );
INV_X4 _GFM_U104  ( .A(b_in[125]), .ZN(_GFM_n2524 ) );
INV_X4 _GFM_U103  ( .A(b_in[123]), .ZN(_GFM_n25040 ) );
INV_X4 _GFM_U102  ( .A(b_in[122]), .ZN(_GFM_n2494 ) );
INV_X4 _GFM_U101  ( .A(b_in[114]), .ZN(_GFM_n24140 ) );
INV_X4 _GFM_U100  ( .A(b_in[115]), .ZN(_GFM_n2423 ) );
INV_X4 _GFM_U99  ( .A(b_in[119]), .ZN(_GFM_n24640 ) );
INV_X4 _GFM_U98  ( .A(b_in[113]), .ZN(_GFM_n2404 ) );
INV_X4 _GFM_U97  ( .A(b_in[121]), .ZN(_GFM_n24830 ) );
INV_X4 _GFM_U96  ( .A(b_in[117]), .ZN(_GFM_n24430 ) );
INV_X4 _GFM_U95  ( .A(b_in[116]), .ZN(_GFM_n24330 ) );
INV_X4 _GFM_U94  ( .A(b_in[125]), .ZN(_GFM_n2523 ) );
INV_X4 _GFM_U93  ( .A(b_in[123]), .ZN(_GFM_n2503 ) );
INV_X4 _GFM_U92  ( .A(b_in[124]), .ZN(_GFM_n25140 ) );
INV_X4 _GFM_U91  ( .A(b_in[113]), .ZN(_GFM_n24030 ) );
INV_X4 _GFM_U90  ( .A(b_in[117]), .ZN(_GFM_n24420 ) );
INV_X4 _GFM_U89  ( .A(b_in[118]), .ZN(_GFM_n24520 ) );
INV_X4 _GFM_U88  ( .A(b_in[116]), .ZN(_GFM_n2432 ) );
INV_X4 _GFM_U87  ( .A(b_in[125]), .ZN(_GFM_n25220 ) );
INV_X4 _GFM_U86  ( .A(b_in[123]), .ZN(_GFM_n2502 ) );
INV_X4 _GFM_U85  ( .A(b_in[124]), .ZN(_GFM_n2513 ) );
INV_X4 _GFM_U84  ( .A(b_in[122]), .ZN(_GFM_n2493 ) );
INV_X4 _GFM_U83  ( .A(b_in[117]), .ZN(_GFM_n2441 ) );
INV_X4 _GFM_U82  ( .A(b_in[118]), .ZN(_GFM_n24511 ) );
INV_X4 _GFM_U81  ( .A(b_in[116]), .ZN(_GFM_n2431 ) );
INV_X4 _GFM_U80  ( .A(b_in[125]), .ZN(_GFM_n25210 ) );
INV_X4 _GFM_U79  ( .A(b_in[123]), .ZN(_GFM_n25010 ) );
INV_X4 _GFM_U78  ( .A(b_in[124]), .ZN(_GFM_n25120 ) );
INV_X4 _GFM_U77  ( .A(b_in[122]), .ZN(_GFM_n24921 ) );
INV_X4 _GFM_U76  ( .A(b_in[119]), .ZN(_GFM_n2461 ) );
INV_X4 _GFM_U75  ( .A(b_in[114]), .ZN(_GFM_n24120 ) );
INV_X4 _GFM_U74  ( .A(b_in[115]), .ZN(_GFM_n24210 ) );
INV_X4 _GFM_U73  ( .A(b_in[113]), .ZN(_GFM_n24020 ) );
INV_X4 _GFM_U72  ( .A(b_in[116]), .ZN(_GFM_n2430 ) );
INV_X4 _GFM_U71  ( .A(b_in[125]), .ZN(_GFM_n25201 ) );
INV_X4 _GFM_U70  ( .A(b_in[123]), .ZN(_GFM_n25000 ) );
INV_X4 _GFM_U69  ( .A(b_in[124]), .ZN(_GFM_n2511 ) );
INV_X4 _GFM_U68  ( .A(b_in[119]), .ZN(_GFM_n24600 ) );
INV_X4 _GFM_U67  ( .A(b_in[120]), .ZN(_GFM_n24700 ) );
INV_X4 _GFM_U66  ( .A(b_in[114]), .ZN(_GFM_n24110 ) );
INV_X4 _GFM_U65  ( .A(b_in[115]), .ZN(_GFM_n24201 ) );
INV_X4 _GFM_U64  ( .A(b_in[113]), .ZN(_GFM_n2401 ) );
INV_X4 _GFM_U63  ( .A(b_in[121]), .ZN(_GFM_n2480 ) );
INV_X4 _GFM_U62  ( .A(b_in[117]), .ZN(_GFM_n24401 ) );
INV_X4 _GFM_U61  ( .A(b_in[118]), .ZN(_GFM_n24500 ) );
INV_X4 _GFM_U60  ( .A(b_in[124]), .ZN(_GFM_n25101 ) );
INV_X4 _GFM_U59  ( .A(b_in[120]), .ZN(_GFM_n24690 ) );
INV_X4 _GFM_U58  ( .A(b_in[114]), .ZN(_GFM_n24101 ) );
INV_X4 _GFM_U57  ( .A(b_in[115]), .ZN(_GFM_n24190 ) );
INV_X4 _GFM_U56  ( .A(b_in[113]), .ZN(_GFM_n2400 ) );
INV_X4 _GFM_U55  ( .A(b_in[117]), .ZN(_GFM_n24390 ) );
INV_X4 _GFM_U54  ( .A(b_in[118]), .ZN(_GFM_n2449 ) );
INV_X4 _GFM_U53  ( .A(b_in[116]), .ZN(_GFM_n24290 ) );
INV_X4 _GFM_U52  ( .A(b_in[119]), .ZN(_GFM_n24590 ) );
INV_X4 _GFM_U51  ( .A(b_in[122]), .ZN(_GFM_n24910 ) );
INV_X4 _GFM_U50  ( .A(b_in[114]), .ZN(_GFM_n2409 ) );
INV_X4 _GFM_U49  ( .A(b_in[113]), .ZN(_GFM_n2399 ) );
INV_X4 _GFM_U48  ( .A(b_in[121]), .ZN(_GFM_n24810 ) );
INV_X4 _GFM_U47  ( .A(b_in[120]), .ZN(_GFM_n2471 ) );
INV_X4 _GFM_U46  ( .A(b_in[117]), .ZN(_GFM_n2444 ) );
INV_X4 _GFM_U45  ( .A(b_in[118]), .ZN(_GFM_n24530 ) );
INV_X4 _GFM_U44  ( .A(b_in[120]), .ZN(_GFM_n2472 ) );
INV_X4 _GFM_U43  ( .A(b_in[119]), .ZN(_GFM_n2462 ) );
INV_X4 _GFM_U42  ( .A(b_in[121]), .ZN(_GFM_n2482 ) );
INV_X4 _GFM_U41  ( .A(b_in[123]), .ZN(_GFM_n2499 ) );
INV_X4 _GFM_U40  ( .A(b_in[113]), .ZN(_GFM_n23980 ) );
INV_X4 _GFM_U39  ( .A(b_in[124]), .ZN(_GFM_n25080 ) );
INV_X4 _GFM_U38  ( .A(b_in[115]), .ZN(_GFM_n2417 ) );
INV_X4 _GFM_U37  ( .A(b_in[127]), .ZN(_GFM_n25450 ) );
INV_X4 _GFM_U36  ( .A(b_in[126]), .ZN(_GFM_n25350 ) );
INV_X4 _GFM_U35  ( .A(b_in[119]), .ZN(_GFM_n24570 ) );
INV_X4 _GFM_U34  ( .A(b_in[118]), .ZN(_GFM_n2447 ) );
INV_X4 _GFM_U33  ( .A(b_in[117]), .ZN(_GFM_n2437 ) );
INV_X4 _GFM_U32  ( .A(b_in[123]), .ZN(_GFM_n24980 ) );
INV_X4 _GFM_U31  ( .A(b_in[112]), .ZN(_GFM_n23880 ) );
INV_X4 _GFM_U30  ( .A(b_in[112]), .ZN(_GFM_n23950 ) );
INV_X4 _GFM_U29  ( .A(b_in[112]), .ZN(_GFM_n23940 ) );
INV_X4 _GFM_U28  ( .A(b_in[112]), .ZN(_GFM_n2393 ) );
INV_X4 _GFM_U27  ( .A(b_in[112]), .ZN(_GFM_n2392 ) );
INV_X4 _GFM_U26  ( .A(b_in[112]), .ZN(_GFM_n23910 ) );
INV_X4 _GFM_U25  ( .A(b_in[112]), .ZN(_GFM_n23900 ) );
INV_X4 _GFM_U24  ( .A(b_in[125]), .ZN(_GFM_n25190 ) );
INV_X4 _GFM_U23  ( .A(b_in[112]), .ZN(_GFM_n2389 ) );
INV_X4 _GFM_U22  ( .A(b_in[124]), .ZN(_GFM_n2509 ) );
INV_X4 _GFM_U21  ( .A(b_in[125]), .ZN(_GFM_n25180 ) );
INV_X4 _GFM_U20  ( .A(b_in[122]), .ZN(_GFM_n24900 ) );
INV_X4 _GFM_U19  ( .A(b_in[126]), .ZN(_GFM_n25290 ) );
INV_X4 _GFM_U18  ( .A(b_in[126]), .ZN(_GFM_n2528 ) );
INV_X4 _GFM_U17  ( .A(b_in[127]), .ZN(_GFM_n2544 ) );
INV_X4 _GFM_U16  ( .A(b_in[126]), .ZN(_GFM_n2534 ) );
INV_X4 _GFM_U15  ( .A(b_in[127]), .ZN(_GFM_n25430 ) );
INV_X4 _GFM_U14  ( .A(b_in[126]), .ZN(_GFM_n2533 ) );
INV_X4 _GFM_U13  ( .A(b_in[127]), .ZN(_GFM_n2542 ) );
INV_X4 _GFM_U12  ( .A(b_in[126]), .ZN(_GFM_n25320 ) );
INV_X4 _GFM_U11  ( .A(b_in[127]), .ZN(_GFM_n2541 ) );
INV_X4 _GFM_U10  ( .A(b_in[126]), .ZN(_GFM_n25310 ) );
INV_X4 _GFM_U9  ( .A(b_in[127]), .ZN(_GFM_n2540 ) );
INV_X4 _GFM_U8  ( .A(b_in[126]), .ZN(_GFM_n2530 ) );
INV_X4 _GFM_U7  ( .A(b_in[127]), .ZN(_GFM_n25390 ) );
INV_X4 _GFM_U6  ( .A(b_in[127]), .ZN(_GFM_n25380 ) );
INV_X4 _GFM_U5  ( .A(b_in[127]), .ZN(_GFM_n2537 ) );
INV_X4 _GFM_U4  ( .A(b_in[126]), .ZN(_GFM_n25270 ) );
INV_X4 _GFM_U3  ( .A(b_in[114]), .ZN(_GFM_n24080 ) );
INV_X4 _GFM_U2  ( .A(b_in[120]), .ZN(_GFM_n24670 ) );
XOR2_X2 _GFM_U755  ( .A(v_in[121]), .B(v_in[0]), .Z(v_out[105]) );
XNOR2_X2 _GFM_U737  ( .A(_GFM_n2695 ), .B(v_in[1]), .ZN(v_out[106]) );
XNOR2_X2 _GFM_U717  ( .A(_GFM_n2696 ), .B(v_in[2]), .ZN(v_out[107]) );
XNOR2_X2 _GFM_U699  ( .A(_GFM_n2697 ), .B(v_in[3]), .ZN(v_out[108]) );
XNOR2_X2 _GFM_U679  ( .A(_GFM_n26980 ), .B(v_in[4]), .ZN(v_out[109]) );
AND2_X2 _GFM_U487  ( .A1(v_out[119]), .A2(b_in[112]), .ZN(_GFM_N3990 ) );
AND2_X2 _GFM_U486  ( .A1(v_in[121]), .A2(b_in[127]), .ZN(_GFM_N3994 ) );
XOR2_X2 _GFM_U479  ( .A(v_in[126]), .B(_GFM_n25460 ), .Z(_GFM_n21360 ) );
AND2_X2 _GFM_U389  ( .A1(v_out[124]), .A2(b_in[112]), .ZN(_GFM_N4272 ) );
AND2_X2 _GFM_U388  ( .A1(b_in[127]), .A2(v_in[126]), .ZN(_GFM_N4276 ) );
NAND2_X2 _GFM_U386  ( .A1(_GFM_N4324 ), .A2(_GFM_n2699 ), .ZN(_GFM_n2134 ));
NAND2_X2 _GFM_U384  ( .A1(_GFM_n2134 ), .A2(_GFM_n21350 ), .ZN(_GFM_N4279 ));
NAND2_X2 _GFM_U381  ( .A1(_GFM_N4325 ), .A2(_GFM_n25460 ), .ZN(_GFM_n21320 ));
NAND2_X2 _GFM_U379  ( .A1(_GFM_n21320 ), .A2(_GFM_n21330 ), .ZN(_GFM_N4282 ));
NAND2_X2 _GFM_U377  ( .A1(_GFM_N4329 ), .A2(_GFM_n2554 ), .ZN(_GFM_n21301 ));
NAND2_X2 _GFM_U375  ( .A1(_GFM_n21301 ), .A2(_GFM_n2131 ), .ZN(_GFM_N4284 ));
NAND2_X2 _GFM_U373  ( .A1(_GFM_N4331 ), .A2(_GFM_n25620 ), .ZN(_GFM_n21280 ));
NAND2_X2 _GFM_U371  ( .A1(_GFM_n21280 ), .A2(_GFM_n21290 ), .ZN(_GFM_N4288 ));
NAND2_X2 _GFM_U369  ( .A1(_GFM_N4328 ), .A2(_GFM_n25580 ), .ZN(_GFM_n21260 ));
NAND2_X2 _GFM_U367  ( .A1(_GFM_n21260 ), .A2(_GFM_n2127 ), .ZN(_GFM_N4290 ));
NAND2_X2 _GFM_U365  ( .A1(_GFM_N4332 ), .A2(_GFM_n25660 ), .ZN(_GFM_n21240 ));
NAND2_X2 _GFM_U363  ( .A1(_GFM_n21240 ), .A2(_GFM_n2125 ), .ZN(_GFM_N4293 ));
NAND2_X2 _GFM_U361  ( .A1(_GFM_N4342 ), .A2(_GFM_n25700 ), .ZN(_GFM_n2122 ));
NAND2_X2 _GFM_U359  ( .A1(_GFM_n2122 ), .A2(_GFM_n21230 ), .ZN(_GFM_N4295 ));
NAND2_X2 _GFM_U356  ( .A1(_GFM_N4336 ), .A2(_GFM_n2578 ), .ZN(_GFM_n184 ) );
NAND2_X2 _GFM_U354  ( .A1(_GFM_n184 ), .A2(_GFM_n2121 ), .ZN(_GFM_N4300 ) );
NAND2_X2 _GFM_U352  ( .A1(_GFM_N4339 ), .A2(_GFM_n25800 ), .ZN(_GFM_n18210 ));
NAND2_X2 _GFM_U350  ( .A1(_GFM_n18210 ), .A2(_GFM_n18310 ), .ZN(_GFM_N4302 ));
NAND2_X2 _GFM_U348  ( .A1(_GFM_N4337 ), .A2(_GFM_n25760 ), .ZN(_GFM_n18011 ));
NAND2_X2 _GFM_U346  ( .A1(_GFM_n18011 ), .A2(_GFM_n181 ), .ZN(_GFM_N4305 ));
NAND2_X2 _GFM_U344  ( .A1(_GFM_N4341 ), .A2(_GFM_n2573 ), .ZN(_GFM_n178 ) );
NAND2_X2 _GFM_U342  ( .A1(_GFM_n178 ), .A2(_GFM_n17911 ), .ZN(_GFM_N4307 ));
NAND2_X2 _GFM_U339  ( .A1(_GFM_N4345 ), .A2(_GFM_n25840 ), .ZN(_GFM_n17611 ));
NAND2_X2 _GFM_U337  ( .A1(_GFM_n17611 ), .A2(_GFM_n177 ), .ZN(_GFM_N4311 ));
NAND2_X2 _GFM_U335  ( .A1(_GFM_N4346 ), .A2(_GFM_n25821 ), .ZN(_GFM_n174 ));
NAND2_X2 _GFM_U333  ( .A1(_GFM_n174 ), .A2(_GFM_n17511 ), .ZN(_GFM_N4313 ));
NAND2_X2 _GFM_U331  ( .A1(_GFM_N4348 ), .A2(_GFM_n2586 ), .ZN(_GFM_n172 ) );
NAND2_X2 _GFM_U329  ( .A1(_GFM_n172 ), .A2(_GFM_n17310 ), .ZN(_GFM_N4316 ));
NAND2_X2 _GFM_U327  ( .A1(_GFM_N4349 ), .A2(_GFM_n2587 ), .ZN(_GFM_n17011 ));
NAND2_X2 _GFM_U325  ( .A1(_GFM_n17011 ), .A2(_GFM_n17110 ), .ZN(_GFM_N4318 ));
XOR2_X2 _GFM_U1  ( .A(v_in[15]), .B(v_in[14]), .Z(v_out[126]) );
XOR2_X2 _GFM_U4328  ( .A(_GFM_n186 ), .B(_GFM_n185 ), .Z(z_out[0]) );
XOR2_X2 _GFM_U4327  ( .A(_GFM_n188 ), .B(_GFM_n18720 ), .Z(_GFM_n185 ) );
XOR2_X2 _GFM_U4326  ( .A(_GFM_n19000 ), .B(_GFM_n18900 ), .Z(_GFM_n186 ) );
XOR2_X2 _GFM_U4325  ( .A(_GFM_n192 ), .B(_GFM_n191 ), .Z(_GFM_n18720 ) );
XOR2_X2 _GFM_U4324  ( .A(_GFM_n19410 ), .B(_GFM_n19310 ), .Z(_GFM_n188 ) );
XOR2_X2 _GFM_U4323  ( .A(_GFM_n19620 ), .B(_GFM_n195 ), .Z(_GFM_n18900 ) );
XOR2_X2 _GFM_U4322  ( .A(_GFM_n198 ), .B(_GFM_n19700 ), .Z(_GFM_n19000 ) );
XOR2_X2 _GFM_U4321  ( .A(z_in[0]), .B(_GFM_n199 ), .Z(_GFM_n191 ) );
XOR2_X2 _GFM_U4320  ( .A(_GFM_N27 ), .B(_GFM_N28 ), .Z(_GFM_n192 ) );
XOR2_X2 _GFM_U4319  ( .A(_GFM_N24 ), .B(_GFM_N25 ), .Z(_GFM_n19310 ) );
XOR2_X2 _GFM_U4318  ( .A(_GFM_N20 ), .B(_GFM_N21 ), .Z(_GFM_n19410 ) );
XOR2_X2 _GFM_U4317  ( .A(_GFM_N16 ), .B(_GFM_N18 ), .Z(_GFM_n195 ) );
XOR2_X2 _GFM_U4316  ( .A(_GFM_N11 ), .B(_GFM_N15 ), .Z(_GFM_n19620 ) );
XOR2_X2 _GFM_U4315  ( .A(_GFM_N8 ), .B(_GFM_N10 ), .Z(_GFM_n19700 ) );
XOR2_X2 _GFM_U4314  ( .A(_GFM_N4 ), .B(_GFM_N7 ), .Z(_GFM_n198 ) );
XOR2_X2 _GFM_U4313  ( .A(_GFM_N1 ), .B(_GFM_N3 ), .Z(_GFM_n199 ) );
XOR2_X2 _GFM_U4312  ( .A(_GFM_n20100 ), .B(_GFM_n200 ), .Z(z_out[1]) );
XOR2_X2 _GFM_U4311  ( .A(_GFM_n203 ), .B(_GFM_n20200 ), .Z(_GFM_n200 ) );
XOR2_X2 _GFM_U4310  ( .A(_GFM_n205 ), .B(_GFM_n20410 ), .Z(_GFM_n20100 ) );
XOR2_X2 _GFM_U4309  ( .A(_GFM_n20720 ), .B(_GFM_n20600 ), .Z(_GFM_n20200 ));
XOR2_X2 _GFM_U4308  ( .A(_GFM_n209 ), .B(_GFM_n208 ), .Z(_GFM_n203 ) );
XOR2_X2 _GFM_U4307  ( .A(_GFM_n21100 ), .B(_GFM_n21000 ), .Z(_GFM_n20410 ));
XOR2_X2 _GFM_U4306  ( .A(_GFM_n21300 ), .B(_GFM_n212 ), .Z(_GFM_n205 ) );
XOR2_X2 _GFM_U4305  ( .A(z_in[1]), .B(_GFM_n2141 ), .Z(_GFM_n20600 ) );
XOR2_X2 _GFM_U4304  ( .A(_GFM_N58 ), .B(_GFM_N59 ), .Z(_GFM_n20720 ) );
XOR2_X2 _GFM_U4303  ( .A(_GFM_N55 ), .B(_GFM_N56 ), .Z(_GFM_n208 ) );
XOR2_X2 _GFM_U4302  ( .A(_GFM_N51 ), .B(_GFM_N52 ), .Z(_GFM_n209 ) );
XOR2_X2 _GFM_U4301  ( .A(_GFM_N47 ), .B(_GFM_N49 ), .Z(_GFM_n21000 ) );
XOR2_X2 _GFM_U4300  ( .A(_GFM_N42 ), .B(_GFM_N46 ), .Z(_GFM_n21100 ) );
XOR2_X2 _GFM_U4299  ( .A(_GFM_N39 ), .B(_GFM_N41 ), .Z(_GFM_n212 ) );
XOR2_X2 _GFM_U4298  ( .A(_GFM_N35 ), .B(_GFM_N38 ), .Z(_GFM_n21300 ) );
XOR2_X2 _GFM_U4297  ( .A(_GFM_N32 ), .B(_GFM_N34 ), .Z(_GFM_n2141 ) );
XOR2_X2 _GFM_U4296  ( .A(_GFM_n216 ), .B(_GFM_n215 ), .Z(z_out[2]) );
XOR2_X2 _GFM_U4295  ( .A(_GFM_n2182 ), .B(_GFM_n217 ), .Z(_GFM_n215 ) );
XOR2_X2 _GFM_U4294  ( .A(_GFM_n2200 ), .B(_GFM_n219 ), .Z(_GFM_n216 ) );
XOR2_X2 _GFM_U4293  ( .A(_GFM_n222 ), .B(_GFM_n2210 ), .Z(_GFM_n217 ) );
XOR2_X2 _GFM_U4292  ( .A(_GFM_n2241 ), .B(_GFM_n223 ), .Z(_GFM_n2182 ) );
XOR2_X2 _GFM_U4291  ( .A(_GFM_n226 ), .B(_GFM_n2251 ), .Z(_GFM_n219 ) );
XOR2_X2 _GFM_U4290  ( .A(_GFM_n2280 ), .B(_GFM_n2272 ), .Z(_GFM_n2200 ) );
XOR2_X2 _GFM_U4289  ( .A(z_in[2]), .B(_GFM_n229 ), .Z(_GFM_n2210 ) );
XOR2_X2 _GFM_U4288  ( .A(_GFM_N89 ), .B(_GFM_N90 ), .Z(_GFM_n222 ) );
XOR2_X2 _GFM_U4287  ( .A(_GFM_N86 ), .B(_GFM_N87 ), .Z(_GFM_n223 ) );
XOR2_X2 _GFM_U4286  ( .A(_GFM_N82 ), .B(_GFM_N83 ), .Z(_GFM_n2241 ) );
XOR2_X2 _GFM_U4285  ( .A(_GFM_N78 ), .B(_GFM_N80 ), .Z(_GFM_n2251 ) );
XOR2_X2 _GFM_U4284  ( .A(_GFM_N73 ), .B(_GFM_N77 ), .Z(_GFM_n226 ) );
XOR2_X2 _GFM_U4283  ( .A(_GFM_N70 ), .B(_GFM_N72 ), .Z(_GFM_n2272 ) );
XOR2_X2 _GFM_U4282  ( .A(_GFM_N66 ), .B(_GFM_N69 ), .Z(_GFM_n2280 ) );
XOR2_X2 _GFM_U4281  ( .A(_GFM_N63 ), .B(_GFM_N65 ), .Z(_GFM_n229 ) );
XOR2_X2 _GFM_U4280  ( .A(_GFM_n231 ), .B(_GFM_n230 ), .Z(z_out[3]) );
XOR2_X2 _GFM_U4279  ( .A(_GFM_n2330 ), .B(_GFM_n2320 ), .Z(_GFM_n230 ) );
XOR2_X2 _GFM_U4278  ( .A(_GFM_n2351 ), .B(_GFM_n234 ), .Z(_GFM_n231 ) );
XOR2_X2 _GFM_U4277  ( .A(_GFM_n2370 ), .B(_GFM_n236 ), .Z(_GFM_n2320 ) );
XOR2_X2 _GFM_U4276  ( .A(_GFM_n239 ), .B(_GFM_n2382 ), .Z(_GFM_n2330 ) );
XOR2_X2 _GFM_U4275  ( .A(_GFM_n24100 ), .B(_GFM_n240 ), .Z(_GFM_n234 ) );
XOR2_X2 _GFM_U4274  ( .A(_GFM_n243 ), .B(_GFM_n24200 ), .Z(_GFM_n2351 ) );
XOR2_X2 _GFM_U4273  ( .A(z_in[3]), .B(_GFM_n24400 ), .Z(_GFM_n236 ) );
XOR2_X2 _GFM_U4272  ( .A(_GFM_N120 ), .B(_GFM_N121 ), .Z(_GFM_n2370 ) );
XOR2_X2 _GFM_U4271  ( .A(_GFM_N117 ), .B(_GFM_N118 ), .Z(_GFM_n2382 ) );
XOR2_X2 _GFM_U4270  ( .A(_GFM_N113 ), .B(_GFM_N114 ), .Z(_GFM_n239 ) );
XOR2_X2 _GFM_U4269  ( .A(_GFM_N109 ), .B(_GFM_N111 ), .Z(_GFM_n240 ) );
XOR2_X2 _GFM_U4268  ( .A(_GFM_N104 ), .B(_GFM_N108 ), .Z(_GFM_n24100 ) );
XOR2_X2 _GFM_U4267  ( .A(_GFM_N101 ), .B(_GFM_N103 ), .Z(_GFM_n24200 ) );
XOR2_X2 _GFM_U4266  ( .A(_GFM_N97 ), .B(_GFM_N100 ), .Z(_GFM_n243 ) );
XOR2_X2 _GFM_U4265  ( .A(_GFM_N94 ), .B(_GFM_N96 ), .Z(_GFM_n24400 ) );
XOR2_X2 _GFM_U4264  ( .A(_GFM_n246 ), .B(_GFM_n24510 ), .Z(z_out[4]) );
XOR2_X2 _GFM_U4263  ( .A(_GFM_n248 ), .B(_GFM_n247 ), .Z(_GFM_n24510 ) );
XOR2_X2 _GFM_U4262  ( .A(_GFM_n250 ), .B(_GFM_n24920 ), .Z(_GFM_n246 ) );
XOR2_X2 _GFM_U4261  ( .A(_GFM_n25200 ), .B(_GFM_n25100 ), .Z(_GFM_n247 ) );
XOR2_X2 _GFM_U4260  ( .A(_GFM_n254 ), .B(_GFM_n253 ), .Z(_GFM_n248 ) );
XOR2_X2 _GFM_U4259  ( .A(_GFM_n25610 ), .B(_GFM_n25510 ), .Z(_GFM_n24920 ));
XOR2_X2 _GFM_U4258  ( .A(_GFM_n25820 ), .B(_GFM_n257 ), .Z(_GFM_n250 ) );
XOR2_X2 _GFM_U4257  ( .A(z_in[4]), .B(_GFM_n25900 ), .Z(_GFM_n25100 ) );
XOR2_X2 _GFM_U4256  ( .A(_GFM_N151 ), .B(_GFM_N152 ), .Z(_GFM_n25200 ) );
XOR2_X2 _GFM_U4255  ( .A(_GFM_N148 ), .B(_GFM_N149 ), .Z(_GFM_n253 ) );
XOR2_X2 _GFM_U4254  ( .A(_GFM_N144 ), .B(_GFM_N145 ), .Z(_GFM_n254 ) );
XOR2_X2 _GFM_U4253  ( .A(_GFM_N140 ), .B(_GFM_N142 ), .Z(_GFM_n25510 ) );
XOR2_X2 _GFM_U4252  ( .A(_GFM_N135 ), .B(_GFM_N139 ), .Z(_GFM_n25610 ) );
XOR2_X2 _GFM_U4251  ( .A(_GFM_N132 ), .B(_GFM_N134 ), .Z(_GFM_n257 ) );
XOR2_X2 _GFM_U4250  ( .A(_GFM_N128 ), .B(_GFM_N131 ), .Z(_GFM_n25820 ) );
XOR2_X2 _GFM_U4249  ( .A(_GFM_N125 ), .B(_GFM_N127 ), .Z(_GFM_n25900 ) );
XOR2_X2 _GFM_U4248  ( .A(_GFM_n261 ), .B(_GFM_n260 ), .Z(z_out[5]) );
XOR2_X2 _GFM_U4247  ( .A(_GFM_n26300 ), .B(_GFM_n262 ), .Z(_GFM_n260 ) );
XOR2_X2 _GFM_U4246  ( .A(_GFM_n265 ), .B(_GFM_n26400 ), .Z(_GFM_n261 ) );
XOR2_X2 _GFM_U4245  ( .A(_GFM_n267 ), .B(_GFM_n26610 ), .Z(_GFM_n262 ) );
XOR2_X2 _GFM_U4244  ( .A(_GFM_n26920 ), .B(_GFM_n26800 ), .Z(_GFM_n26300 ));
XOR2_X2 _GFM_U4243  ( .A(_GFM_n271 ), .B(_GFM_n270 ), .Z(_GFM_n26400 ) );
XOR2_X2 _GFM_U4242  ( .A(_GFM_n2730 ), .B(_GFM_n2720 ), .Z(_GFM_n265 ) );
XOR2_X2 _GFM_U4241  ( .A(z_in[5]), .B(_GFM_n274 ), .Z(_GFM_n26610 ) );
XOR2_X2 _GFM_U4240  ( .A(_GFM_N182 ), .B(_GFM_N183 ), .Z(_GFM_n267 ) );
XOR2_X2 _GFM_U4239  ( .A(_GFM_N179 ), .B(_GFM_N180 ), .Z(_GFM_n26800 ) );
XOR2_X2 _GFM_U4238  ( .A(_GFM_N175 ), .B(_GFM_N176 ), .Z(_GFM_n26920 ) );
XOR2_X2 _GFM_U4237  ( .A(_GFM_N171 ), .B(_GFM_N173 ), .Z(_GFM_n270 ) );
XOR2_X2 _GFM_U4236  ( .A(_GFM_N166 ), .B(_GFM_N170 ), .Z(_GFM_n271 ) );
XOR2_X2 _GFM_U4235  ( .A(_GFM_N163 ), .B(_GFM_N165 ), .Z(_GFM_n2720 ) );
XOR2_X2 _GFM_U4234  ( .A(_GFM_N159 ), .B(_GFM_N162 ), .Z(_GFM_n2730 ) );
XOR2_X2 _GFM_U4233  ( .A(_GFM_N156 ), .B(_GFM_N158 ), .Z(_GFM_n274 ) );
XOR2_X2 _GFM_U4232  ( .A(_GFM_n2761 ), .B(_GFM_n2750 ), .Z(z_out[6]) );
XOR2_X2 _GFM_U4231  ( .A(_GFM_n278 ), .B(_GFM_n277 ), .Z(_GFM_n2750 ) );
XOR2_X2 _GFM_U4230  ( .A(_GFM_n2802 ), .B(_GFM_n279 ), .Z(_GFM_n2761 ) );
XOR2_X2 _GFM_U4229  ( .A(_GFM_n2820 ), .B(_GFM_n281 ), .Z(_GFM_n277 ) );
XOR2_X2 _GFM_U4228  ( .A(_GFM_n284 ), .B(_GFM_n2830 ), .Z(_GFM_n278 ) );
XOR2_X2 _GFM_U4227  ( .A(_GFM_n2861 ), .B(_GFM_n285 ), .Z(_GFM_n279 ) );
XOR2_X2 _GFM_U4226  ( .A(_GFM_n288 ), .B(_GFM_n2871 ), .Z(_GFM_n2802 ) );
XOR2_X2 _GFM_U4225  ( .A(z_in[6]), .B(_GFM_n2892 ), .Z(_GFM_n281 ) );
XOR2_X2 _GFM_U4224  ( .A(_GFM_N213 ), .B(_GFM_N214 ), .Z(_GFM_n2820 ) );
XOR2_X2 _GFM_U4223  ( .A(_GFM_N210 ), .B(_GFM_N211 ), .Z(_GFM_n2830 ) );
XOR2_X2 _GFM_U4222  ( .A(_GFM_N206 ), .B(_GFM_N207 ), .Z(_GFM_n284 ) );
XOR2_X2 _GFM_U4221  ( .A(_GFM_N202 ), .B(_GFM_N204 ), .Z(_GFM_n285 ) );
XOR2_X2 _GFM_U4220  ( .A(_GFM_N197 ), .B(_GFM_N201 ), .Z(_GFM_n2861 ) );
XOR2_X2 _GFM_U4219  ( .A(_GFM_N194 ), .B(_GFM_N196 ), .Z(_GFM_n2871 ) );
XOR2_X2 _GFM_U4218  ( .A(_GFM_N190 ), .B(_GFM_N193 ), .Z(_GFM_n288 ) );
XOR2_X2 _GFM_U4217  ( .A(_GFM_N187 ), .B(_GFM_N189 ), .Z(_GFM_n2892 ) );
XOR2_X2 _GFM_U4216  ( .A(_GFM_n291 ), .B(_GFM_n2900 ), .Z(z_out[7]) );
XOR2_X2 _GFM_U4215  ( .A(_GFM_n293 ), .B(_GFM_n292 ), .Z(_GFM_n2900 ) );
XOR2_X2 _GFM_U4214  ( .A(_GFM_n2950 ), .B(_GFM_n2940 ), .Z(_GFM_n291 ) );
XOR2_X2 _GFM_U4213  ( .A(_GFM_n2971 ), .B(_GFM_n296 ), .Z(_GFM_n292 ) );
XOR2_X2 _GFM_U4212  ( .A(_GFM_n2990 ), .B(_GFM_n298 ), .Z(_GFM_n293 ) );
XOR2_X2 _GFM_U4211  ( .A(_GFM_n301 ), .B(_GFM_n3002 ), .Z(_GFM_n2940 ) );
XOR2_X2 _GFM_U4210  ( .A(_GFM_n3030 ), .B(_GFM_n302 ), .Z(_GFM_n2950 ) );
XOR2_X2 _GFM_U4209  ( .A(z_in[7]), .B(_GFM_n3040 ), .Z(_GFM_n296 ) );
XOR2_X2 _GFM_U4208  ( .A(_GFM_N244 ), .B(_GFM_N245 ), .Z(_GFM_n2971 ) );
XOR2_X2 _GFM_U4207  ( .A(_GFM_N241 ), .B(_GFM_N242 ), .Z(_GFM_n298 ) );
XOR2_X2 _GFM_U4206  ( .A(_GFM_N237 ), .B(_GFM_N238 ), .Z(_GFM_n2990 ) );
XOR2_X2 _GFM_U4205  ( .A(_GFM_N233 ), .B(_GFM_N235 ), .Z(_GFM_n3002 ) );
XOR2_X2 _GFM_U4204  ( .A(_GFM_N228 ), .B(_GFM_N232 ), .Z(_GFM_n301 ) );
XOR2_X2 _GFM_U4203  ( .A(_GFM_N225 ), .B(_GFM_N227 ), .Z(_GFM_n302 ) );
XOR2_X2 _GFM_U4202  ( .A(_GFM_N221 ), .B(_GFM_N224 ), .Z(_GFM_n3030 ) );
XOR2_X2 _GFM_U4201  ( .A(_GFM_N218 ), .B(_GFM_N220 ), .Z(_GFM_n3040 ) );
XOR2_X2 _GFM_U4200  ( .A(_GFM_n3060 ), .B(_GFM_n305 ), .Z(z_out[8]) );
XOR2_X2 _GFM_U4199  ( .A(_GFM_n308 ), .B(_GFM_n3071 ), .Z(_GFM_n305 ) );
XOR2_X2 _GFM_U4198  ( .A(_GFM_n310 ), .B(_GFM_n309 ), .Z(_GFM_n3060 ) );
XOR2_X2 _GFM_U4197  ( .A(_GFM_n312 ), .B(_GFM_n3112 ), .Z(_GFM_n3071 ) );
XOR2_X2 _GFM_U4196  ( .A(_GFM_n3140 ), .B(_GFM_n3130 ), .Z(_GFM_n308 ) );
XOR2_X2 _GFM_U4195  ( .A(_GFM_n316 ), .B(_GFM_n315 ), .Z(_GFM_n309 ) );
XOR2_X2 _GFM_U4194  ( .A(_GFM_n3181 ), .B(_GFM_n3171 ), .Z(_GFM_n310 ) );
XOR2_X2 _GFM_U4193  ( .A(z_in[8]), .B(_GFM_n319 ), .Z(_GFM_n3112 ) );
XOR2_X2 _GFM_U4192  ( .A(_GFM_N275 ), .B(_GFM_N276 ), .Z(_GFM_n312 ) );
XOR2_X2 _GFM_U4191  ( .A(_GFM_N272 ), .B(_GFM_N273 ), .Z(_GFM_n3130 ) );
XOR2_X2 _GFM_U4190  ( .A(_GFM_N268 ), .B(_GFM_N269 ), .Z(_GFM_n3140 ) );
XOR2_X2 _GFM_U4189  ( .A(_GFM_N264 ), .B(_GFM_N266 ), .Z(_GFM_n315 ) );
XOR2_X2 _GFM_U4188  ( .A(_GFM_N259 ), .B(_GFM_N263 ), .Z(_GFM_n316 ) );
XOR2_X2 _GFM_U4187  ( .A(_GFM_N256 ), .B(_GFM_N258 ), .Z(_GFM_n3171 ) );
XOR2_X2 _GFM_U4186  ( .A(_GFM_N252 ), .B(_GFM_N255 ), .Z(_GFM_n3181 ) );
XOR2_X2 _GFM_U4185  ( .A(_GFM_N249 ), .B(_GFM_N251 ), .Z(_GFM_n319 ) );
XOR2_X2 _GFM_U4184  ( .A(_GFM_n3210 ), .B(_GFM_n3202 ), .Z(z_out[9]) );
XOR2_X2 _GFM_U4183  ( .A(_GFM_n323 ), .B(_GFM_n322 ), .Z(_GFM_n3202 ) );
XOR2_X2 _GFM_U4182  ( .A(_GFM_n3250 ), .B(_GFM_n324 ), .Z(_GFM_n3210 ) );
XOR2_X2 _GFM_U4181  ( .A(_GFM_n327 ), .B(_GFM_n3260 ), .Z(_GFM_n322 ) );
XOR2_X2 _GFM_U4180  ( .A(_GFM_n329 ), .B(_GFM_n3281 ), .Z(_GFM_n323 ) );
XOR2_X2 _GFM_U4179  ( .A(_GFM_n3310 ), .B(_GFM_n3300 ), .Z(_GFM_n324 ) );
XOR2_X2 _GFM_U4178  ( .A(_GFM_n333 ), .B(_GFM_n332 ), .Z(_GFM_n3250 ) );
XOR2_X2 _GFM_U4177  ( .A(z_in[9]), .B(_GFM_n3342 ), .Z(_GFM_n3260 ) );
XOR2_X2 _GFM_U4176  ( .A(_GFM_N306 ), .B(_GFM_N307 ), .Z(_GFM_n327 ) );
XOR2_X2 _GFM_U4175  ( .A(_GFM_N303 ), .B(_GFM_N304 ), .Z(_GFM_n3281 ) );
XOR2_X2 _GFM_U4174  ( .A(_GFM_N299 ), .B(_GFM_N300 ), .Z(_GFM_n329 ) );
XOR2_X2 _GFM_U4173  ( .A(_GFM_N295 ), .B(_GFM_N297 ), .Z(_GFM_n3300 ) );
XOR2_X2 _GFM_U4172  ( .A(_GFM_N290 ), .B(_GFM_N294 ), .Z(_GFM_n3310 ) );
XOR2_X2 _GFM_U4171  ( .A(_GFM_N287 ), .B(_GFM_N289 ), .Z(_GFM_n332 ) );
XOR2_X2 _GFM_U4170  ( .A(_GFM_N283 ), .B(_GFM_N286 ), .Z(_GFM_n333 ) );
XOR2_X2 _GFM_U4169  ( .A(_GFM_N280 ), .B(_GFM_N282 ), .Z(_GFM_n3342 ) );
XOR2_X2 _GFM_U4168  ( .A(_GFM_n336 ), .B(_GFM_n3350 ), .Z(z_out[10]) );
XOR2_X2 _GFM_U4167  ( .A(_GFM_n3381 ), .B(_GFM_n3370 ), .Z(_GFM_n3350 ) );
XOR2_X2 _GFM_U4166  ( .A(_GFM_n340 ), .B(_GFM_n339 ), .Z(_GFM_n336 ) );
XOR2_X2 _GFM_U4165  ( .A(_GFM_n3420 ), .B(_GFM_n341 ), .Z(_GFM_n3370 ) );
XOR2_X2 _GFM_U4164  ( .A(_GFM_n3440 ), .B(_GFM_n343 ), .Z(_GFM_n3381 ) );
XOR2_X2 _GFM_U4163  ( .A(_GFM_n346 ), .B(_GFM_n3451 ), .Z(_GFM_n339 ) );
XOR2_X2 _GFM_U4162  ( .A(_GFM_n3480 ), .B(_GFM_n347 ), .Z(_GFM_n340 ) );
XOR2_X2 _GFM_U4161  ( .A(z_in[10]), .B(_GFM_n3490 ), .Z(_GFM_n341 ) );
XOR2_X2 _GFM_U4160  ( .A(_GFM_N337 ), .B(_GFM_N338 ), .Z(_GFM_n3420 ) );
XOR2_X2 _GFM_U4159  ( .A(_GFM_N334 ), .B(_GFM_N335 ), .Z(_GFM_n343 ) );
XOR2_X2 _GFM_U4158  ( .A(_GFM_N330 ), .B(_GFM_N331 ), .Z(_GFM_n3440 ) );
XOR2_X2 _GFM_U4157  ( .A(_GFM_N326 ), .B(_GFM_N328 ), .Z(_GFM_n3451 ) );
XOR2_X2 _GFM_U4156  ( .A(_GFM_N321 ), .B(_GFM_N325 ), .Z(_GFM_n346 ) );
XOR2_X2 _GFM_U4155  ( .A(_GFM_N318 ), .B(_GFM_N320 ), .Z(_GFM_n347 ) );
XOR2_X2 _GFM_U4154  ( .A(_GFM_N314 ), .B(_GFM_N317 ), .Z(_GFM_n3480 ) );
XOR2_X2 _GFM_U4153  ( .A(_GFM_N311 ), .B(_GFM_N313 ), .Z(_GFM_n3490 ) );
XOR2_X2 _GFM_U4152  ( .A(_GFM_n3510 ), .B(_GFM_n350 ), .Z(z_out[11]) );
XOR2_X2 _GFM_U4151  ( .A(_GFM_n353 ), .B(_GFM_n3520 ), .Z(_GFM_n350 ) );
XOR2_X2 _GFM_U4150  ( .A(_GFM_n355 ), .B(_GFM_n354 ), .Z(_GFM_n3510 ) );
XOR2_X2 _GFM_U4149  ( .A(_GFM_n3570 ), .B(_GFM_n3560 ), .Z(_GFM_n3520 ) );
XOR2_X2 _GFM_U4148  ( .A(_GFM_n3590 ), .B(_GFM_n358 ), .Z(_GFM_n353 ) );
XOR2_X2 _GFM_U4147  ( .A(_GFM_n3610 ), .B(_GFM_n360 ), .Z(_GFM_n354 ) );
XOR2_X2 _GFM_U4146  ( .A(_GFM_n363 ), .B(_GFM_n3621 ), .Z(_GFM_n355 ) );
XOR2_X2 _GFM_U4145  ( .A(z_in[11]), .B(_GFM_n364 ), .Z(_GFM_n3560 ) );
XOR2_X2 _GFM_U4144  ( .A(_GFM_N368 ), .B(_GFM_N369 ), .Z(_GFM_n3570 ) );
XOR2_X2 _GFM_U4143  ( .A(_GFM_N365 ), .B(_GFM_N366 ), .Z(_GFM_n358 ) );
XOR2_X2 _GFM_U4142  ( .A(_GFM_N361 ), .B(_GFM_N362 ), .Z(_GFM_n3590 ) );
XOR2_X2 _GFM_U4141  ( .A(_GFM_N357 ), .B(_GFM_N359 ), .Z(_GFM_n360 ) );
XOR2_X2 _GFM_U4140  ( .A(_GFM_N352 ), .B(_GFM_N356 ), .Z(_GFM_n3610 ) );
XOR2_X2 _GFM_U4139  ( .A(_GFM_N349 ), .B(_GFM_N351 ), .Z(_GFM_n3621 ) );
XOR2_X2 _GFM_U4138  ( .A(_GFM_N345 ), .B(_GFM_N348 ), .Z(_GFM_n363 ) );
XOR2_X2 _GFM_U4137  ( .A(_GFM_N342 ), .B(_GFM_N344 ), .Z(_GFM_n364 ) );
XOR2_X2 _GFM_U4136  ( .A(_GFM_n3660 ), .B(_GFM_n3650 ), .Z(z_out[12]) );
XOR2_X2 _GFM_U4135  ( .A(_GFM_n3680 ), .B(_GFM_n367 ), .Z(_GFM_n3650 ) );
XOR2_X2 _GFM_U4134  ( .A(_GFM_n370 ), .B(_GFM_n3691 ), .Z(_GFM_n3660 ) );
XOR2_X2 _GFM_U4133  ( .A(_GFM_n372 ), .B(_GFM_n371 ), .Z(_GFM_n367 ) );
XOR2_X2 _GFM_U4132  ( .A(_GFM_n374 ), .B(_GFM_n3730 ), .Z(_GFM_n3680 ) );
XOR2_X2 _GFM_U4131  ( .A(_GFM_n3760 ), .B(_GFM_n3751 ), .Z(_GFM_n3691 ) );
XOR2_X2 _GFM_U4130  ( .A(_GFM_n378 ), .B(_GFM_n377 ), .Z(_GFM_n370 ) );
XOR2_X2 _GFM_U4129  ( .A(z_in[12]), .B(_GFM_n3790 ), .Z(_GFM_n371 ) );
XOR2_X2 _GFM_U4128  ( .A(_GFM_N399 ), .B(_GFM_N400 ), .Z(_GFM_n372 ) );
XOR2_X2 _GFM_U4127  ( .A(_GFM_N396 ), .B(_GFM_N397 ), .Z(_GFM_n3730 ) );
XOR2_X2 _GFM_U4126  ( .A(_GFM_N392 ), .B(_GFM_N393 ), .Z(_GFM_n374 ) );
XOR2_X2 _GFM_U4125  ( .A(_GFM_N388 ), .B(_GFM_N390 ), .Z(_GFM_n3751 ) );
XOR2_X2 _GFM_U4124  ( .A(_GFM_N383 ), .B(_GFM_N387 ), .Z(_GFM_n3760 ) );
XOR2_X2 _GFM_U4123  ( .A(_GFM_N380 ), .B(_GFM_N382 ), .Z(_GFM_n377 ) );
XOR2_X2 _GFM_U4122  ( .A(_GFM_N376 ), .B(_GFM_N379 ), .Z(_GFM_n378 ) );
XOR2_X2 _GFM_U4121  ( .A(_GFM_N373 ), .B(_GFM_N375 ), .Z(_GFM_n3790 ) );
XOR2_X2 _GFM_U4120  ( .A(_GFM_n381 ), .B(_GFM_n3800 ), .Z(z_out[13]) );
XOR2_X2 _GFM_U4119  ( .A(_GFM_n3830 ), .B(_GFM_n3820 ), .Z(_GFM_n3800 ) );
XOR2_X2 _GFM_U4118  ( .A(_GFM_n385 ), .B(_GFM_n384 ), .Z(_GFM_n381 ) );
XOR2_X2 _GFM_U4117  ( .A(_GFM_n3870 ), .B(_GFM_n386 ), .Z(_GFM_n3820 ) );
XOR2_X2 _GFM_U4116  ( .A(_GFM_n389 ), .B(_GFM_n3880 ), .Z(_GFM_n3830 ) );
XOR2_X2 _GFM_U4115  ( .A(_GFM_n391 ), .B(_GFM_n3900 ), .Z(_GFM_n384 ) );
XOR2_X2 _GFM_U4114  ( .A(_GFM_n3930 ), .B(_GFM_n3920 ), .Z(_GFM_n385 ) );
XOR2_X2 _GFM_U4113  ( .A(z_in[13]), .B(_GFM_n394 ), .Z(_GFM_n386 ) );
XOR2_X2 _GFM_U4112  ( .A(_GFM_N430 ), .B(_GFM_N431 ), .Z(_GFM_n3870 ) );
XOR2_X2 _GFM_U4111  ( .A(_GFM_N427 ), .B(_GFM_N428 ), .Z(_GFM_n3880 ) );
XOR2_X2 _GFM_U4110  ( .A(_GFM_N423 ), .B(_GFM_N424 ), .Z(_GFM_n389 ) );
XOR2_X2 _GFM_U4109  ( .A(_GFM_N419 ), .B(_GFM_N421 ), .Z(_GFM_n3900 ) );
XOR2_X2 _GFM_U4108  ( .A(_GFM_N414 ), .B(_GFM_N418 ), .Z(_GFM_n391 ) );
XOR2_X2 _GFM_U4107  ( .A(_GFM_N411 ), .B(_GFM_N413 ), .Z(_GFM_n3920 ) );
XOR2_X2 _GFM_U4106  ( .A(_GFM_N407 ), .B(_GFM_N410 ), .Z(_GFM_n3930 ) );
XOR2_X2 _GFM_U4105  ( .A(_GFM_N404 ), .B(_GFM_N406 ), .Z(_GFM_n394 ) );
XOR2_X2 _GFM_U4104  ( .A(_GFM_n3960 ), .B(_GFM_n395 ), .Z(z_out[14]) );
XOR2_X2 _GFM_U4103  ( .A(_GFM_n398 ), .B(_GFM_n3970 ), .Z(_GFM_n395 ) );
XOR2_X2 _GFM_U4102  ( .A(_GFM_n4000 ), .B(_GFM_n3991 ), .Z(_GFM_n3960 ) );
XOR2_X2 _GFM_U4101  ( .A(_GFM_n402 ), .B(_GFM_n401 ), .Z(_GFM_n3970 ) );
XOR2_X2 _GFM_U4100  ( .A(_GFM_n4040 ), .B(_GFM_n403 ), .Z(_GFM_n398 ) );
XOR2_X2 _GFM_U4099  ( .A(_GFM_n4060 ), .B(_GFM_n405 ), .Z(_GFM_n3991 ) );
XOR2_X2 _GFM_U4098  ( .A(_GFM_n408 ), .B(_GFM_n4070 ), .Z(_GFM_n4000 ) );
XOR2_X2 _GFM_U4097  ( .A(z_in[14]), .B(_GFM_n409 ), .Z(_GFM_n401 ) );
XOR2_X2 _GFM_U4096  ( .A(_GFM_N461 ), .B(_GFM_N462 ), .Z(_GFM_n402 ) );
XOR2_X2 _GFM_U4095  ( .A(_GFM_N458 ), .B(_GFM_N459 ), .Z(_GFM_n403 ) );
XOR2_X2 _GFM_U4094  ( .A(_GFM_N454 ), .B(_GFM_N455 ), .Z(_GFM_n4040 ) );
XOR2_X2 _GFM_U4093  ( .A(_GFM_N450 ), .B(_GFM_N452 ), .Z(_GFM_n405 ) );
XOR2_X2 _GFM_U4092  ( .A(_GFM_N445 ), .B(_GFM_N449 ), .Z(_GFM_n4060 ) );
XOR2_X2 _GFM_U4091  ( .A(_GFM_N442 ), .B(_GFM_N444 ), .Z(_GFM_n4070 ) );
XOR2_X2 _GFM_U4090  ( .A(_GFM_N438 ), .B(_GFM_N441 ), .Z(_GFM_n408 ) );
XOR2_X2 _GFM_U4089  ( .A(_GFM_N435 ), .B(_GFM_N437 ), .Z(_GFM_n409 ) );
XOR2_X2 _GFM_U4088  ( .A(_GFM_n4110 ), .B(_GFM_n4100 ), .Z(z_out[15]) );
XOR2_X2 _GFM_U4087  ( .A(_GFM_n4130 ), .B(_GFM_n412 ), .Z(_GFM_n4100 ) );
XOR2_X2 _GFM_U4086  ( .A(_GFM_n415 ), .B(_GFM_n4140 ), .Z(_GFM_n4110 ) );
XOR2_X2 _GFM_U4085  ( .A(_GFM_n417 ), .B(_GFM_n416 ), .Z(_GFM_n412 ) );
XOR2_X2 _GFM_U4084  ( .A(_GFM_n4190 ), .B(_GFM_n4180 ), .Z(_GFM_n4130 ) );
XOR2_X2 _GFM_U4083  ( .A(_GFM_n4211 ), .B(_GFM_n420 ), .Z(_GFM_n4140 ) );
XOR2_X2 _GFM_U4082  ( .A(_GFM_n4230 ), .B(_GFM_n422 ), .Z(_GFM_n415 ) );
XOR2_X2 _GFM_U4081  ( .A(z_in[15]), .B(_GFM_n4241 ), .Z(_GFM_n416 ) );
XOR2_X2 _GFM_U4080  ( .A(_GFM_N492 ), .B(_GFM_N493 ), .Z(_GFM_n417 ) );
XOR2_X2 _GFM_U4079  ( .A(_GFM_N489 ), .B(_GFM_N490 ), .Z(_GFM_n4180 ) );
XOR2_X2 _GFM_U4078  ( .A(_GFM_N485 ), .B(_GFM_N486 ), .Z(_GFM_n4190 ) );
XOR2_X2 _GFM_U4077  ( .A(_GFM_N481 ), .B(_GFM_N483 ), .Z(_GFM_n420 ) );
XOR2_X2 _GFM_U4076  ( .A(_GFM_N476 ), .B(_GFM_N480 ), .Z(_GFM_n4211 ) );
XOR2_X2 _GFM_U4075  ( .A(_GFM_N473 ), .B(_GFM_N475 ), .Z(_GFM_n422 ) );
XOR2_X2 _GFM_U4074  ( .A(_GFM_N469 ), .B(_GFM_N472 ), .Z(_GFM_n4230 ) );
XOR2_X2 _GFM_U4073  ( .A(_GFM_N466 ), .B(_GFM_N468 ), .Z(_GFM_n4241 ) );
XOR2_X2 _GFM_U4072  ( .A(_GFM_n426 ), .B(_GFM_n425 ), .Z(z_out[16]) );
XOR2_X2 _GFM_U4071  ( .A(_GFM_n4280 ), .B(_GFM_n4270 ), .Z(_GFM_n425 ) );
XOR2_X2 _GFM_U4070  ( .A(_GFM_n4301 ), .B(_GFM_n429 ), .Z(_GFM_n426 ) );
XOR2_X2 _GFM_U4069  ( .A(_GFM_n432 ), .B(_GFM_n4310 ), .Z(_GFM_n4270 ) );
XOR2_X2 _GFM_U4068  ( .A(_GFM_n434 ), .B(_GFM_n433 ), .Z(_GFM_n4280 ) );
XOR2_X2 _GFM_U4067  ( .A(_GFM_n436 ), .B(_GFM_n4350 ), .Z(_GFM_n429 ) );
XOR2_X2 _GFM_U4066  ( .A(_GFM_n4380 ), .B(_GFM_n4370 ), .Z(_GFM_n4301 ) );
XOR2_X2 _GFM_U4065  ( .A(z_in[16]), .B(_GFM_n439 ), .Z(_GFM_n4310 ) );
XOR2_X2 _GFM_U4064  ( .A(_GFM_N523 ), .B(_GFM_N524 ), .Z(_GFM_n432 ) );
XOR2_X2 _GFM_U4063  ( .A(_GFM_N520 ), .B(_GFM_N521 ), .Z(_GFM_n433 ) );
XOR2_X2 _GFM_U4062  ( .A(_GFM_N516 ), .B(_GFM_N517 ), .Z(_GFM_n434 ) );
XOR2_X2 _GFM_U4061  ( .A(_GFM_N512 ), .B(_GFM_N514 ), .Z(_GFM_n4350 ) );
XOR2_X2 _GFM_U4060  ( .A(_GFM_N507 ), .B(_GFM_N511 ), .Z(_GFM_n436 ) );
XOR2_X2 _GFM_U4059  ( .A(_GFM_N504 ), .B(_GFM_N506 ), .Z(_GFM_n4370 ) );
XOR2_X2 _GFM_U4058  ( .A(_GFM_N500 ), .B(_GFM_N503 ), .Z(_GFM_n4380 ) );
XOR2_X2 _GFM_U4057  ( .A(_GFM_N497 ), .B(_GFM_N499 ), .Z(_GFM_n439 ) );
XOR2_X2 _GFM_U4056  ( .A(_GFM_n4410 ), .B(_GFM_n440 ), .Z(z_out[17]) );
XOR2_X2 _GFM_U4055  ( .A(_GFM_n443 ), .B(_GFM_n4420 ), .Z(_GFM_n440 ) );
XOR2_X2 _GFM_U4054  ( .A(_GFM_n4450 ), .B(_GFM_n4440 ), .Z(_GFM_n4410 ) );
XOR2_X2 _GFM_U4053  ( .A(_GFM_n447 ), .B(_GFM_n446 ), .Z(_GFM_n4420 ) );
XOR2_X2 _GFM_U4052  ( .A(_GFM_n4490 ), .B(_GFM_n448 ), .Z(_GFM_n443 ) );
XOR2_X2 _GFM_U4051  ( .A(_GFM_n451 ), .B(_GFM_n4500 ), .Z(_GFM_n4440 ) );
XOR2_X2 _GFM_U4050  ( .A(_GFM_n453 ), .B(_GFM_n4520 ), .Z(_GFM_n4450 ) );
XOR2_X2 _GFM_U4049  ( .A(z_in[17]), .B(_GFM_n4540 ), .Z(_GFM_n446 ) );
XOR2_X2 _GFM_U4048  ( .A(_GFM_N554 ), .B(_GFM_N555 ), .Z(_GFM_n447 ) );
XOR2_X2 _GFM_U4047  ( .A(_GFM_N551 ), .B(_GFM_N552 ), .Z(_GFM_n448 ) );
XOR2_X2 _GFM_U4046  ( .A(_GFM_N547 ), .B(_GFM_N548 ), .Z(_GFM_n4490 ) );
XOR2_X2 _GFM_U4045  ( .A(_GFM_N543 ), .B(_GFM_N545 ), .Z(_GFM_n4500 ) );
XOR2_X2 _GFM_U4044  ( .A(_GFM_N538 ), .B(_GFM_N542 ), .Z(_GFM_n451 ) );
XOR2_X2 _GFM_U4043  ( .A(_GFM_N535 ), .B(_GFM_N537 ), .Z(_GFM_n4520 ) );
XOR2_X2 _GFM_U4042  ( .A(_GFM_N531 ), .B(_GFM_N534 ), .Z(_GFM_n453 ) );
XOR2_X2 _GFM_U4041  ( .A(_GFM_N528 ), .B(_GFM_N530 ), .Z(_GFM_n4540 ) );
XOR2_X2 _GFM_U4040  ( .A(_GFM_n456 ), .B(_GFM_n4550 ), .Z(z_out[18]) );
XOR2_X2 _GFM_U4039  ( .A(_GFM_n4580 ), .B(_GFM_n457 ), .Z(_GFM_n4550 ) );
XOR2_X2 _GFM_U4038  ( .A(_GFM_n460 ), .B(_GFM_n4590 ), .Z(_GFM_n456 ) );
XOR2_X2 _GFM_U4037  ( .A(_GFM_n4620 ), .B(_GFM_n4610 ), .Z(_GFM_n457 ) );
XOR2_X2 _GFM_U4036  ( .A(_GFM_n464 ), .B(_GFM_n463 ), .Z(_GFM_n4580 ) );
XOR2_X2 _GFM_U4035  ( .A(_GFM_n4660 ), .B(_GFM_n465 ), .Z(_GFM_n4590 ) );
XOR2_X2 _GFM_U4034  ( .A(_GFM_n4680 ), .B(_GFM_n467 ), .Z(_GFM_n460 ) );
XOR2_X2 _GFM_U4033  ( .A(z_in[18]), .B(_GFM_n4690 ), .Z(_GFM_n4610 ) );
XOR2_X2 _GFM_U4032  ( .A(_GFM_N585 ), .B(_GFM_N586 ), .Z(_GFM_n4620 ) );
XOR2_X2 _GFM_U4031  ( .A(_GFM_N582 ), .B(_GFM_N583 ), .Z(_GFM_n463 ) );
XOR2_X2 _GFM_U4030  ( .A(_GFM_N578 ), .B(_GFM_N579 ), .Z(_GFM_n464 ) );
XOR2_X2 _GFM_U4029  ( .A(_GFM_N574 ), .B(_GFM_N576 ), .Z(_GFM_n465 ) );
XOR2_X2 _GFM_U4028  ( .A(_GFM_N569 ), .B(_GFM_N573 ), .Z(_GFM_n4660 ) );
XOR2_X2 _GFM_U4027  ( .A(_GFM_N566 ), .B(_GFM_N568 ), .Z(_GFM_n467 ) );
XOR2_X2 _GFM_U4026  ( .A(_GFM_N562 ), .B(_GFM_N565 ), .Z(_GFM_n4680 ) );
XOR2_X2 _GFM_U4025  ( .A(_GFM_N559 ), .B(_GFM_N561 ), .Z(_GFM_n4690 ) );
XOR2_X2 _GFM_U4024  ( .A(_GFM_n471 ), .B(_GFM_n470 ), .Z(z_out[19]) );
XOR2_X2 _GFM_U4023  ( .A(_GFM_n4730 ), .B(_GFM_n4720 ), .Z(_GFM_n470 ) );
XOR2_X2 _GFM_U4022  ( .A(_GFM_n4750 ), .B(_GFM_n474 ), .Z(_GFM_n471 ) );
XOR2_X2 _GFM_U4021  ( .A(_GFM_n477 ), .B(_GFM_n4760 ), .Z(_GFM_n4720 ) );
XOR2_X2 _GFM_U4020  ( .A(_GFM_n479 ), .B(_GFM_n478 ), .Z(_GFM_n4730 ) );
XOR2_X2 _GFM_U4019  ( .A(_GFM_n4810 ), .B(_GFM_n4800 ), .Z(_GFM_n474 ) );
XOR2_X2 _GFM_U4018  ( .A(_GFM_n4830 ), .B(_GFM_n482 ), .Z(_GFM_n4750 ) );
XOR2_X2 _GFM_U4017  ( .A(z_in[19]), .B(_GFM_n484 ), .Z(_GFM_n4760 ) );
XOR2_X2 _GFM_U4016  ( .A(_GFM_N616 ), .B(_GFM_N617 ), .Z(_GFM_n477 ) );
XOR2_X2 _GFM_U4015  ( .A(_GFM_N613 ), .B(_GFM_N614 ), .Z(_GFM_n478 ) );
XOR2_X2 _GFM_U4014  ( .A(_GFM_N609 ), .B(_GFM_N610 ), .Z(_GFM_n479 ) );
XOR2_X2 _GFM_U4013  ( .A(_GFM_N605 ), .B(_GFM_N607 ), .Z(_GFM_n4800 ) );
XOR2_X2 _GFM_U4012  ( .A(_GFM_N600 ), .B(_GFM_N604 ), .Z(_GFM_n4810 ) );
XOR2_X2 _GFM_U4011  ( .A(_GFM_N597 ), .B(_GFM_N599 ), .Z(_GFM_n482 ) );
XOR2_X2 _GFM_U4010  ( .A(_GFM_N593 ), .B(_GFM_N596 ), .Z(_GFM_n4830 ) );
XOR2_X2 _GFM_U4009  ( .A(_GFM_N590 ), .B(_GFM_N592 ), .Z(_GFM_n484 ) );
XOR2_X2 _GFM_U4008  ( .A(_GFM_n4860 ), .B(_GFM_n4850 ), .Z(z_out[20]) );
XOR2_X2 _GFM_U4007  ( .A(_GFM_n488 ), .B(_GFM_n487 ), .Z(_GFM_n4850 ) );
XOR2_X2 _GFM_U4006  ( .A(_GFM_n4900 ), .B(_GFM_n4890 ), .Z(_GFM_n4860 ) );
XOR2_X2 _GFM_U4005  ( .A(_GFM_n4920 ), .B(_GFM_n491 ), .Z(_GFM_n487 ) );
XOR2_X2 _GFM_U4004  ( .A(_GFM_n494 ), .B(_GFM_n4930 ), .Z(_GFM_n488 ) );
XOR2_X2 _GFM_U4003  ( .A(_GFM_n496 ), .B(_GFM_n495 ), .Z(_GFM_n4890 ) );
XOR2_X2 _GFM_U4002  ( .A(_GFM_n498 ), .B(_GFM_n4970 ), .Z(_GFM_n4900 ) );
XOR2_X2 _GFM_U4001  ( .A(z_in[20]), .B(_GFM_n4990 ), .Z(_GFM_n491 ) );
XOR2_X2 _GFM_U4000  ( .A(_GFM_N647 ), .B(_GFM_N648 ), .Z(_GFM_n4920 ) );
XOR2_X2 _GFM_U3999  ( .A(_GFM_N644 ), .B(_GFM_N645 ), .Z(_GFM_n4930 ) );
XOR2_X2 _GFM_U3998  ( .A(_GFM_N640 ), .B(_GFM_N641 ), .Z(_GFM_n494 ) );
XOR2_X2 _GFM_U3997  ( .A(_GFM_N636 ), .B(_GFM_N638 ), .Z(_GFM_n495 ) );
XOR2_X2 _GFM_U3996  ( .A(_GFM_N631 ), .B(_GFM_N635 ), .Z(_GFM_n496 ) );
XOR2_X2 _GFM_U3995  ( .A(_GFM_N628 ), .B(_GFM_N630 ), .Z(_GFM_n4970 ) );
XOR2_X2 _GFM_U3994  ( .A(_GFM_N624 ), .B(_GFM_N627 ), .Z(_GFM_n498 ) );
XOR2_X2 _GFM_U3993  ( .A(_GFM_N621 ), .B(_GFM_N623 ), .Z(_GFM_n4990 ) );
XOR2_X2 _GFM_U3992  ( .A(_GFM_n501 ), .B(_GFM_n5000 ), .Z(z_out[21]) );
XOR2_X2 _GFM_U3991  ( .A(_GFM_n5030 ), .B(_GFM_n502 ), .Z(_GFM_n5000 ) );
XOR2_X2 _GFM_U3990  ( .A(_GFM_n505 ), .B(_GFM_n5040 ), .Z(_GFM_n501 ) );
XOR2_X2 _GFM_U3989  ( .A(_GFM_n5070 ), .B(_GFM_n5060 ), .Z(_GFM_n502 ) );
XOR2_X2 _GFM_U3988  ( .A(_GFM_n509 ), .B(_GFM_n508 ), .Z(_GFM_n5030 ) );
XOR2_X2 _GFM_U3987  ( .A(_GFM_n5110 ), .B(_GFM_n510 ), .Z(_GFM_n5040 ) );
XOR2_X2 _GFM_U3986  ( .A(_GFM_n513 ), .B(_GFM_n5120 ), .Z(_GFM_n505 ) );
XOR2_X2 _GFM_U3985  ( .A(z_in[21]), .B(_GFM_n5140 ), .Z(_GFM_n5060 ) );
XOR2_X2 _GFM_U3984  ( .A(_GFM_N678 ), .B(_GFM_N679 ), .Z(_GFM_n5070 ) );
XOR2_X2 _GFM_U3983  ( .A(_GFM_N675 ), .B(_GFM_N676 ), .Z(_GFM_n508 ) );
XOR2_X2 _GFM_U3982  ( .A(_GFM_N671 ), .B(_GFM_N672 ), .Z(_GFM_n509 ) );
XOR2_X2 _GFM_U3981  ( .A(_GFM_N667 ), .B(_GFM_N669 ), .Z(_GFM_n510 ) );
XOR2_X2 _GFM_U3980  ( .A(_GFM_N662 ), .B(_GFM_N666 ), .Z(_GFM_n5110 ) );
XOR2_X2 _GFM_U3979  ( .A(_GFM_N659 ), .B(_GFM_N661 ), .Z(_GFM_n5120 ) );
XOR2_X2 _GFM_U3978  ( .A(_GFM_N655 ), .B(_GFM_N658 ), .Z(_GFM_n513 ) );
XOR2_X2 _GFM_U3977  ( .A(_GFM_N652 ), .B(_GFM_N654 ), .Z(_GFM_n5140 ) );
XOR2_X2 _GFM_U3976  ( .A(_GFM_n5160 ), .B(_GFM_n515 ), .Z(z_out[22]) );
XOR2_X2 _GFM_U3975  ( .A(_GFM_n518 ), .B(_GFM_n5170 ), .Z(_GFM_n515 ) );
XOR2_X2 _GFM_U3974  ( .A(_GFM_n5200 ), .B(_GFM_n519 ), .Z(_GFM_n5160 ) );
XOR2_X2 _GFM_U3973  ( .A(_GFM_n522 ), .B(_GFM_n5210 ), .Z(_GFM_n5170 ) );
XOR2_X2 _GFM_U3972  ( .A(_GFM_n5240 ), .B(_GFM_n5230 ), .Z(_GFM_n518 ) );
XOR2_X2 _GFM_U3971  ( .A(_GFM_n526 ), .B(_GFM_n525 ), .Z(_GFM_n519 ) );
XOR2_X2 _GFM_U3970  ( .A(_GFM_n5280 ), .B(_GFM_n527 ), .Z(_GFM_n5200 ) );
XOR2_X2 _GFM_U3969  ( .A(z_in[22]), .B(_GFM_n529 ), .Z(_GFM_n5210 ) );
XOR2_X2 _GFM_U3968  ( .A(_GFM_N709 ), .B(_GFM_N710 ), .Z(_GFM_n522 ) );
XOR2_X2 _GFM_U3967  ( .A(_GFM_N706 ), .B(_GFM_N707 ), .Z(_GFM_n5230 ) );
XOR2_X2 _GFM_U3966  ( .A(_GFM_N702 ), .B(_GFM_N703 ), .Z(_GFM_n5240 ) );
XOR2_X2 _GFM_U3965  ( .A(_GFM_N698 ), .B(_GFM_N700 ), .Z(_GFM_n525 ) );
XOR2_X2 _GFM_U3964  ( .A(_GFM_N693 ), .B(_GFM_N697 ), .Z(_GFM_n526 ) );
XOR2_X2 _GFM_U3963  ( .A(_GFM_N690 ), .B(_GFM_N692 ), .Z(_GFM_n527 ) );
XOR2_X2 _GFM_U3962  ( .A(_GFM_N686 ), .B(_GFM_N689 ), .Z(_GFM_n5280 ) );
XOR2_X2 _GFM_U3961  ( .A(_GFM_N683 ), .B(_GFM_N685 ), .Z(_GFM_n529 ) );
XOR2_X2 _GFM_U3960  ( .A(_GFM_n5310 ), .B(_GFM_n5300 ), .Z(z_out[23]) );
XOR2_X2 _GFM_U3959  ( .A(_GFM_n533 ), .B(_GFM_n532 ), .Z(_GFM_n5300 ) );
XOR2_X2 _GFM_U3958  ( .A(_GFM_n5350 ), .B(_GFM_n5340 ), .Z(_GFM_n5310 ) );
XOR2_X2 _GFM_U3957  ( .A(_GFM_n5370 ), .B(_GFM_n536 ), .Z(_GFM_n532 ) );
XOR2_X2 _GFM_U3956  ( .A(_GFM_n539 ), .B(_GFM_n5380 ), .Z(_GFM_n533 ) );
XOR2_X2 _GFM_U3955  ( .A(_GFM_n541 ), .B(_GFM_n540 ), .Z(_GFM_n5340 ) );
XOR2_X2 _GFM_U3954  ( .A(_GFM_n5430 ), .B(_GFM_n5420 ), .Z(_GFM_n5350 ) );
XOR2_X2 _GFM_U3953  ( .A(z_in[23]), .B(_GFM_n544 ), .Z(_GFM_n536 ) );
XOR2_X2 _GFM_U3952  ( .A(_GFM_N740 ), .B(_GFM_N741 ), .Z(_GFM_n5370 ) );
XOR2_X2 _GFM_U3951  ( .A(_GFM_N737 ), .B(_GFM_N738 ), .Z(_GFM_n5380 ) );
XOR2_X2 _GFM_U3950  ( .A(_GFM_N733 ), .B(_GFM_N734 ), .Z(_GFM_n539 ) );
XOR2_X2 _GFM_U3949  ( .A(_GFM_N729 ), .B(_GFM_N731 ), .Z(_GFM_n540 ) );
XOR2_X2 _GFM_U3948  ( .A(_GFM_N724 ), .B(_GFM_N728 ), .Z(_GFM_n541 ) );
XOR2_X2 _GFM_U3947  ( .A(_GFM_N721 ), .B(_GFM_N723 ), .Z(_GFM_n5420 ) );
XOR2_X2 _GFM_U3946  ( .A(_GFM_N717 ), .B(_GFM_N720 ), .Z(_GFM_n5430 ) );
XOR2_X2 _GFM_U3945  ( .A(_GFM_N714 ), .B(_GFM_N716 ), .Z(_GFM_n544 ) );
XOR2_X2 _GFM_U3944  ( .A(_GFM_n546 ), .B(_GFM_n5450 ), .Z(z_out[24]) );
XOR2_X2 _GFM_U3943  ( .A(_GFM_n5480 ), .B(_GFM_n5470 ), .Z(_GFM_n5450 ) );
XOR2_X2 _GFM_U3942  ( .A(_GFM_n550 ), .B(_GFM_n549 ), .Z(_GFM_n546 ) );
XOR2_X2 _GFM_U3941  ( .A(_GFM_n5520 ), .B(_GFM_n5510 ), .Z(_GFM_n5470 ) );
XOR2_X2 _GFM_U3940  ( .A(_GFM_n5540 ), .B(_GFM_n553 ), .Z(_GFM_n5480 ) );
XOR2_X2 _GFM_U3939  ( .A(_GFM_n556 ), .B(_GFM_n5550 ), .Z(_GFM_n549 ) );
XOR2_X2 _GFM_U3938  ( .A(_GFM_n558 ), .B(_GFM_n557 ), .Z(_GFM_n550 ) );
XOR2_X2 _GFM_U3937  ( .A(z_in[24]), .B(_GFM_n5590 ), .Z(_GFM_n5510 ) );
XOR2_X2 _GFM_U3936  ( .A(_GFM_N771 ), .B(_GFM_N772 ), .Z(_GFM_n5520 ) );
XOR2_X2 _GFM_U3935  ( .A(_GFM_N768 ), .B(_GFM_N769 ), .Z(_GFM_n553 ) );
XOR2_X2 _GFM_U3934  ( .A(_GFM_N764 ), .B(_GFM_N765 ), .Z(_GFM_n5540 ) );
XOR2_X2 _GFM_U3933  ( .A(_GFM_N760 ), .B(_GFM_N762 ), .Z(_GFM_n5550 ) );
XOR2_X2 _GFM_U3932  ( .A(_GFM_N755 ), .B(_GFM_N759 ), .Z(_GFM_n556 ) );
XOR2_X2 _GFM_U3931  ( .A(_GFM_N752 ), .B(_GFM_N754 ), .Z(_GFM_n557 ) );
XOR2_X2 _GFM_U3930  ( .A(_GFM_N748 ), .B(_GFM_N751 ), .Z(_GFM_n558 ) );
XOR2_X2 _GFM_U3929  ( .A(_GFM_N745 ), .B(_GFM_N747 ), .Z(_GFM_n5590 ) );
XOR2_X2 _GFM_U3928  ( .A(_GFM_n5610 ), .B(_GFM_n560 ), .Z(z_out[25]) );
XOR2_X2 _GFM_U3927  ( .A(_GFM_n563 ), .B(_GFM_n5620 ), .Z(_GFM_n560 ) );
XOR2_X2 _GFM_U3926  ( .A(_GFM_n5650 ), .B(_GFM_n564 ), .Z(_GFM_n5610 ) );
XOR2_X2 _GFM_U3925  ( .A(_GFM_n567 ), .B(_GFM_n5660 ), .Z(_GFM_n5620 ) );
XOR2_X2 _GFM_U3924  ( .A(_GFM_n5690 ), .B(_GFM_n5680 ), .Z(_GFM_n563 ) );
XOR2_X2 _GFM_U3923  ( .A(_GFM_n571 ), .B(_GFM_n570 ), .Z(_GFM_n564 ) );
XOR2_X2 _GFM_U3922  ( .A(_GFM_n5730 ), .B(_GFM_n572 ), .Z(_GFM_n5650 ) );
XOR2_X2 _GFM_U3921  ( .A(z_in[25]), .B(_GFM_n5740 ), .Z(_GFM_n5660 ) );
XOR2_X2 _GFM_U3920  ( .A(_GFM_N802 ), .B(_GFM_N803 ), .Z(_GFM_n567 ) );
XOR2_X2 _GFM_U3919  ( .A(_GFM_N799 ), .B(_GFM_N800 ), .Z(_GFM_n5680 ) );
XOR2_X2 _GFM_U3918  ( .A(_GFM_N795 ), .B(_GFM_N796 ), .Z(_GFM_n5690 ) );
XOR2_X2 _GFM_U3917  ( .A(_GFM_N791 ), .B(_GFM_N793 ), .Z(_GFM_n570 ) );
XOR2_X2 _GFM_U3916  ( .A(_GFM_N786 ), .B(_GFM_N790 ), .Z(_GFM_n571 ) );
XOR2_X2 _GFM_U3915  ( .A(_GFM_N783 ), .B(_GFM_N785 ), .Z(_GFM_n572 ) );
XOR2_X2 _GFM_U3914  ( .A(_GFM_N779 ), .B(_GFM_N782 ), .Z(_GFM_n5730 ) );
XOR2_X2 _GFM_U3913  ( .A(_GFM_N776 ), .B(_GFM_N778 ), .Z(_GFM_n5740 ) );
XOR2_X2 _GFM_U3912  ( .A(_GFM_n5760 ), .B(_GFM_n575 ), .Z(z_out[26]) );
XOR2_X2 _GFM_U3911  ( .A(_GFM_n5780 ), .B(_GFM_n577 ), .Z(_GFM_n575 ) );
XOR2_X2 _GFM_U3910  ( .A(_GFM_n580 ), .B(_GFM_n5790 ), .Z(_GFM_n5760 ) );
XOR2_X2 _GFM_U3909  ( .A(_GFM_n5820 ), .B(_GFM_n581 ), .Z(_GFM_n577 ) );
XOR2_X2 _GFM_U3908  ( .A(_GFM_n584 ), .B(_GFM_n5830 ), .Z(_GFM_n5780 ) );
XOR2_X2 _GFM_U3907  ( .A(_GFM_n5860 ), .B(_GFM_n5850 ), .Z(_GFM_n5790 ) );
XOR2_X2 _GFM_U3906  ( .A(_GFM_n588 ), .B(_GFM_n587 ), .Z(_GFM_n580 ) );
XOR2_X2 _GFM_U3905  ( .A(z_in[26]), .B(_GFM_n589 ), .Z(_GFM_n581 ) );
XOR2_X2 _GFM_U3904  ( .A(_GFM_N833 ), .B(_GFM_N834 ), .Z(_GFM_n5820 ) );
XOR2_X2 _GFM_U3903  ( .A(_GFM_N830 ), .B(_GFM_N831 ), .Z(_GFM_n5830 ) );
XOR2_X2 _GFM_U3902  ( .A(_GFM_N826 ), .B(_GFM_N827 ), .Z(_GFM_n584 ) );
XOR2_X2 _GFM_U3901  ( .A(_GFM_N822 ), .B(_GFM_N824 ), .Z(_GFM_n5850 ) );
XOR2_X2 _GFM_U3900  ( .A(_GFM_N817 ), .B(_GFM_N821 ), .Z(_GFM_n5860 ) );
XOR2_X2 _GFM_U3899  ( .A(_GFM_N814 ), .B(_GFM_N816 ), .Z(_GFM_n587 ) );
XOR2_X2 _GFM_U3898  ( .A(_GFM_N810 ), .B(_GFM_N813 ), .Z(_GFM_n588 ) );
XOR2_X2 _GFM_U3897  ( .A(_GFM_N807 ), .B(_GFM_N809 ), .Z(_GFM_n589 ) );
XOR2_X2 _GFM_U3896  ( .A(_GFM_n591 ), .B(_GFM_n5900 ), .Z(z_out[27]) );
XOR2_X2 _GFM_U3895  ( .A(_GFM_n5930 ), .B(_GFM_n5920 ), .Z(_GFM_n5900 ) );
XOR2_X2 _GFM_U3894  ( .A(_GFM_n595 ), .B(_GFM_n594 ), .Z(_GFM_n591 ) );
XOR2_X2 _GFM_U3893  ( .A(_GFM_n5970 ), .B(_GFM_n5960 ), .Z(_GFM_n5920 ) );
XOR2_X2 _GFM_U3892  ( .A(_GFM_n5990 ), .B(_GFM_n598 ), .Z(_GFM_n5930 ) );
XOR2_X2 _GFM_U3891  ( .A(_GFM_n601 ), .B(_GFM_n6000 ), .Z(_GFM_n594 ) );
XOR2_X2 _GFM_U3890  ( .A(_GFM_n603 ), .B(_GFM_n602 ), .Z(_GFM_n595 ) );
XOR2_X2 _GFM_U3889  ( .A(z_in[27]), .B(_GFM_n6040 ), .Z(_GFM_n5960 ) );
XOR2_X2 _GFM_U3888  ( .A(_GFM_N864 ), .B(_GFM_N865 ), .Z(_GFM_n5970 ) );
XOR2_X2 _GFM_U3887  ( .A(_GFM_N861 ), .B(_GFM_N862 ), .Z(_GFM_n598 ) );
XOR2_X2 _GFM_U3886  ( .A(_GFM_N857 ), .B(_GFM_N858 ), .Z(_GFM_n5990 ) );
XOR2_X2 _GFM_U3885  ( .A(_GFM_N853 ), .B(_GFM_N855 ), .Z(_GFM_n6000 ) );
XOR2_X2 _GFM_U3884  ( .A(_GFM_N848 ), .B(_GFM_N852 ), .Z(_GFM_n601 ) );
XOR2_X2 _GFM_U3883  ( .A(_GFM_N845 ), .B(_GFM_N847 ), .Z(_GFM_n602 ) );
XOR2_X2 _GFM_U3882  ( .A(_GFM_N841 ), .B(_GFM_N844 ), .Z(_GFM_n603 ) );
XOR2_X2 _GFM_U3881  ( .A(_GFM_N838 ), .B(_GFM_N840 ), .Z(_GFM_n6040 ) );
XOR2_X2 _GFM_U3880  ( .A(_GFM_n606 ), .B(_GFM_n6050 ), .Z(z_out[28]) );
XOR2_X2 _GFM_U3879  ( .A(_GFM_n608 ), .B(_GFM_n6070 ), .Z(_GFM_n6050 ) );
XOR2_X2 _GFM_U3878  ( .A(_GFM_n6100 ), .B(_GFM_n6090 ), .Z(_GFM_n606 ) );
XOR2_X2 _GFM_U3877  ( .A(_GFM_n612 ), .B(_GFM_n611 ), .Z(_GFM_n6070 ) );
XOR2_X2 _GFM_U3876  ( .A(_GFM_n6140 ), .B(_GFM_n6130 ), .Z(_GFM_n608 ) );
XOR2_X2 _GFM_U3875  ( .A(_GFM_n6160 ), .B(_GFM_n615 ), .Z(_GFM_n6090 ) );
XOR2_X2 _GFM_U3874  ( .A(_GFM_n618 ), .B(_GFM_n6170 ), .Z(_GFM_n6100 ) );
XOR2_X2 _GFM_U3873  ( .A(z_in[28]), .B(_GFM_n619 ), .Z(_GFM_n611 ) );
XOR2_X2 _GFM_U3872  ( .A(_GFM_N895 ), .B(_GFM_N896 ), .Z(_GFM_n612 ) );
XOR2_X2 _GFM_U3871  ( .A(_GFM_N892 ), .B(_GFM_N893 ), .Z(_GFM_n6130 ) );
XOR2_X2 _GFM_U3870  ( .A(_GFM_N888 ), .B(_GFM_N889 ), .Z(_GFM_n6140 ) );
XOR2_X2 _GFM_U3869  ( .A(_GFM_N884 ), .B(_GFM_N886 ), .Z(_GFM_n615 ) );
XOR2_X2 _GFM_U3868  ( .A(_GFM_N879 ), .B(_GFM_N883 ), .Z(_GFM_n6160 ) );
XOR2_X2 _GFM_U3867  ( .A(_GFM_N876 ), .B(_GFM_N878 ), .Z(_GFM_n6170 ) );
XOR2_X2 _GFM_U3866  ( .A(_GFM_N872 ), .B(_GFM_N875 ), .Z(_GFM_n618 ) );
XOR2_X2 _GFM_U3865  ( .A(_GFM_N869 ), .B(_GFM_N871 ), .Z(_GFM_n619 ) );
XOR2_X2 _GFM_U3864  ( .A(_GFM_n6210 ), .B(_GFM_n620 ), .Z(z_out[29]) );
XOR2_X2 _GFM_U3863  ( .A(_GFM_n6230 ), .B(_GFM_n622 ), .Z(_GFM_n620 ) );
XOR2_X2 _GFM_U3862  ( .A(_GFM_n625 ), .B(_GFM_n6240 ), .Z(_GFM_n6210 ) );
XOR2_X2 _GFM_U3861  ( .A(_GFM_n6270 ), .B(_GFM_n626 ), .Z(_GFM_n622 ) );
XOR2_X2 _GFM_U3860  ( .A(_GFM_n629 ), .B(_GFM_n6280 ), .Z(_GFM_n6230 ) );
XOR2_X2 _GFM_U3859  ( .A(_GFM_n6310 ), .B(_GFM_n6300 ), .Z(_GFM_n6240 ) );
XOR2_X2 _GFM_U3858  ( .A(_GFM_n633 ), .B(_GFM_n632 ), .Z(_GFM_n625 ) );
XOR2_X2 _GFM_U3857  ( .A(z_in[29]), .B(_GFM_n634 ), .Z(_GFM_n626 ) );
XOR2_X2 _GFM_U3856  ( .A(_GFM_N926 ), .B(_GFM_N927 ), .Z(_GFM_n6270 ) );
XOR2_X2 _GFM_U3855  ( .A(_GFM_N923 ), .B(_GFM_N924 ), .Z(_GFM_n6280 ) );
XOR2_X2 _GFM_U3854  ( .A(_GFM_N919 ), .B(_GFM_N920 ), .Z(_GFM_n629 ) );
XOR2_X2 _GFM_U3853  ( .A(_GFM_N915 ), .B(_GFM_N917 ), .Z(_GFM_n6300 ) );
XOR2_X2 _GFM_U3852  ( .A(_GFM_N910 ), .B(_GFM_N914 ), .Z(_GFM_n6310 ) );
XOR2_X2 _GFM_U3851  ( .A(_GFM_N907 ), .B(_GFM_N909 ), .Z(_GFM_n632 ) );
XOR2_X2 _GFM_U3850  ( .A(_GFM_N903 ), .B(_GFM_N906 ), .Z(_GFM_n633 ) );
XOR2_X2 _GFM_U3849  ( .A(_GFM_N900 ), .B(_GFM_N902 ), .Z(_GFM_n634 ) );
XOR2_X2 _GFM_U3848  ( .A(_GFM_n6360 ), .B(_GFM_n6350 ), .Z(z_out[30]) );
XOR2_X2 _GFM_U3847  ( .A(_GFM_n6380 ), .B(_GFM_n637 ), .Z(_GFM_n6350 ) );
XOR2_X2 _GFM_U3846  ( .A(_GFM_n6400 ), .B(_GFM_n639 ), .Z(_GFM_n6360 ) );
XOR2_X2 _GFM_U3845  ( .A(_GFM_n642 ), .B(_GFM_n6410 ), .Z(_GFM_n637 ) );
XOR2_X2 _GFM_U3844  ( .A(_GFM_n6440 ), .B(_GFM_n643 ), .Z(_GFM_n6380 ) );
XOR2_X2 _GFM_U3843  ( .A(_GFM_n646 ), .B(_GFM_n6450 ), .Z(_GFM_n639 ) );
XOR2_X2 _GFM_U3842  ( .A(_GFM_n6480 ), .B(_GFM_n6470 ), .Z(_GFM_n6400 ) );
XOR2_X2 _GFM_U3841  ( .A(z_in[30]), .B(_GFM_n649 ), .Z(_GFM_n6410 ) );
XOR2_X2 _GFM_U3840  ( .A(_GFM_N957 ), .B(_GFM_N958 ), .Z(_GFM_n642 ) );
XOR2_X2 _GFM_U3839  ( .A(_GFM_N954 ), .B(_GFM_N955 ), .Z(_GFM_n643 ) );
XOR2_X2 _GFM_U3838  ( .A(_GFM_N950 ), .B(_GFM_N951 ), .Z(_GFM_n6440 ) );
XOR2_X2 _GFM_U3837  ( .A(_GFM_N946 ), .B(_GFM_N948 ), .Z(_GFM_n6450 ) );
XOR2_X2 _GFM_U3836  ( .A(_GFM_N941 ), .B(_GFM_N945 ), .Z(_GFM_n646 ) );
XOR2_X2 _GFM_U3835  ( .A(_GFM_N938 ), .B(_GFM_N940 ), .Z(_GFM_n6470 ) );
XOR2_X2 _GFM_U3834  ( .A(_GFM_N934 ), .B(_GFM_N937 ), .Z(_GFM_n6480 ) );
XOR2_X2 _GFM_U3833  ( .A(_GFM_N931 ), .B(_GFM_N933 ), .Z(_GFM_n649 ) );
XOR2_X2 _GFM_U3832  ( .A(_GFM_n651 ), .B(_GFM_n650 ), .Z(z_out[31]) );
XOR2_X2 _GFM_U3831  ( .A(_GFM_n653 ), .B(_GFM_n6520 ), .Z(_GFM_n650 ) );
XOR2_X2 _GFM_U3830  ( .A(_GFM_n6550 ), .B(_GFM_n6540 ), .Z(_GFM_n651 ) );
XOR2_X2 _GFM_U3829  ( .A(_GFM_n657 ), .B(_GFM_n656 ), .Z(_GFM_n6520 ) );
XOR2_X2 _GFM_U3828  ( .A(_GFM_n6590 ), .B(_GFM_n6580 ), .Z(_GFM_n653 ) );
XOR2_X2 _GFM_U3827  ( .A(_GFM_n6610 ), .B(_GFM_n660 ), .Z(_GFM_n6540 ) );
XOR2_X2 _GFM_U3826  ( .A(_GFM_n663 ), .B(_GFM_n6620 ), .Z(_GFM_n6550 ) );
XOR2_X2 _GFM_U3825  ( .A(z_in[31]), .B(_GFM_n664 ), .Z(_GFM_n656 ) );
XOR2_X2 _GFM_U3824  ( .A(_GFM_N988 ), .B(_GFM_N989 ), .Z(_GFM_n657 ) );
XOR2_X2 _GFM_U3823  ( .A(_GFM_N985 ), .B(_GFM_N986 ), .Z(_GFM_n6580 ) );
XOR2_X2 _GFM_U3822  ( .A(_GFM_N981 ), .B(_GFM_N982 ), .Z(_GFM_n6590 ) );
XOR2_X2 _GFM_U3821  ( .A(_GFM_N977 ), .B(_GFM_N979 ), .Z(_GFM_n660 ) );
XOR2_X2 _GFM_U3820  ( .A(_GFM_N972 ), .B(_GFM_N976 ), .Z(_GFM_n6610 ) );
XOR2_X2 _GFM_U3819  ( .A(_GFM_N969 ), .B(_GFM_N971 ), .Z(_GFM_n6620 ) );
XOR2_X2 _GFM_U3818  ( .A(_GFM_N965 ), .B(_GFM_N968 ), .Z(_GFM_n663 ) );
XOR2_X2 _GFM_U3817  ( .A(_GFM_N962 ), .B(_GFM_N964 ), .Z(_GFM_n664 ) );
XOR2_X2 _GFM_U3816  ( .A(_GFM_n6660 ), .B(_GFM_n665 ), .Z(z_out[32]) );
XOR2_X2 _GFM_U3815  ( .A(_GFM_n668 ), .B(_GFM_n6670 ), .Z(_GFM_n665 ) );
XOR2_X2 _GFM_U3814  ( .A(_GFM_n670 ), .B(_GFM_n6690 ), .Z(_GFM_n6660 ) );
XOR2_X2 _GFM_U3813  ( .A(_GFM_n6720 ), .B(_GFM_n6710 ), .Z(_GFM_n6670 ) );
XOR2_X2 _GFM_U3812  ( .A(_GFM_n674 ), .B(_GFM_n673 ), .Z(_GFM_n668 ) );
XOR2_X2 _GFM_U3811  ( .A(_GFM_n6760 ), .B(_GFM_n6750 ), .Z(_GFM_n6690 ) );
XOR2_X2 _GFM_U3810  ( .A(_GFM_n6780 ), .B(_GFM_n677 ), .Z(_GFM_n670 ) );
XOR2_X2 _GFM_U3809  ( .A(z_in[32]), .B(_GFM_n6790 ), .Z(_GFM_n6710 ) );
XOR2_X2 _GFM_U3808  ( .A(_GFM_N1019 ), .B(_GFM_N1020 ), .Z(_GFM_n6720 ) );
XOR2_X2 _GFM_U3807  ( .A(_GFM_N1016 ), .B(_GFM_N1017 ), .Z(_GFM_n673 ) );
XOR2_X2 _GFM_U3806  ( .A(_GFM_N1012 ), .B(_GFM_N1013 ), .Z(_GFM_n674 ) );
XOR2_X2 _GFM_U3805  ( .A(_GFM_N1008 ), .B(_GFM_N1010 ), .Z(_GFM_n6750 ) );
XOR2_X2 _GFM_U3804  ( .A(_GFM_N1003 ), .B(_GFM_N1007 ), .Z(_GFM_n6760 ) );
XOR2_X2 _GFM_U3803  ( .A(_GFM_N1000 ), .B(_GFM_N1002 ), .Z(_GFM_n677 ) );
XOR2_X2 _GFM_U3802  ( .A(_GFM_N996 ), .B(_GFM_N999 ), .Z(_GFM_n6780 ) );
XOR2_X2 _GFM_U3801  ( .A(_GFM_N993 ), .B(_GFM_N995 ), .Z(_GFM_n6790 ) );
XOR2_X2 _GFM_U3800  ( .A(_GFM_n681 ), .B(_GFM_n680 ), .Z(z_out[33]) );
XOR2_X2 _GFM_U3799  ( .A(_GFM_n6830 ), .B(_GFM_n682 ), .Z(_GFM_n680 ) );
XOR2_X2 _GFM_U3798  ( .A(_GFM_n6850 ), .B(_GFM_n684 ), .Z(_GFM_n681 ) );
XOR2_X2 _GFM_U3797  ( .A(_GFM_n687 ), .B(_GFM_n6860 ), .Z(_GFM_n682 ) );
XOR2_X2 _GFM_U3796  ( .A(_GFM_n6890 ), .B(_GFM_n688 ), .Z(_GFM_n6830 ) );
XOR2_X2 _GFM_U3795  ( .A(_GFM_n691 ), .B(_GFM_n6900 ), .Z(_GFM_n684 ) );
XOR2_X2 _GFM_U3794  ( .A(_GFM_n6930 ), .B(_GFM_n6920 ), .Z(_GFM_n6850 ) );
XOR2_X2 _GFM_U3793  ( .A(z_in[33]), .B(_GFM_n694 ), .Z(_GFM_n6860 ) );
XOR2_X2 _GFM_U3792  ( .A(_GFM_N1050 ), .B(_GFM_N1051 ), .Z(_GFM_n687 ) );
XOR2_X2 _GFM_U3791  ( .A(_GFM_N1047 ), .B(_GFM_N1048 ), .Z(_GFM_n688 ) );
XOR2_X2 _GFM_U3790  ( .A(_GFM_N1043 ), .B(_GFM_N1044 ), .Z(_GFM_n6890 ) );
XOR2_X2 _GFM_U3789  ( .A(_GFM_N1039 ), .B(_GFM_N1041 ), .Z(_GFM_n6900 ) );
XOR2_X2 _GFM_U3788  ( .A(_GFM_N1034 ), .B(_GFM_N1038 ), .Z(_GFM_n691 ) );
XOR2_X2 _GFM_U3787  ( .A(_GFM_N1031 ), .B(_GFM_N1033 ), .Z(_GFM_n6920 ) );
XOR2_X2 _GFM_U3786  ( .A(_GFM_N1027 ), .B(_GFM_N1030 ), .Z(_GFM_n6930 ) );
XOR2_X2 _GFM_U3785  ( .A(_GFM_N1024 ), .B(_GFM_N1026 ), .Z(_GFM_n694 ) );
XOR2_X2 _GFM_U3784  ( .A(_GFM_n696 ), .B(_GFM_n695 ), .Z(z_out[34]) );
XOR2_X2 _GFM_U3783  ( .A(_GFM_n6980 ), .B(_GFM_n6970 ), .Z(_GFM_n695 ) );
XOR2_X2 _GFM_U3782  ( .A(_GFM_n7000 ), .B(_GFM_n699 ), .Z(_GFM_n696 ) );
XOR2_X2 _GFM_U3781  ( .A(_GFM_n7020 ), .B(_GFM_n701 ), .Z(_GFM_n6970 ) );
XOR2_X2 _GFM_U3780  ( .A(_GFM_n704 ), .B(_GFM_n7030 ), .Z(_GFM_n6980 ) );
XOR2_X2 _GFM_U3779  ( .A(_GFM_n7060 ), .B(_GFM_n705 ), .Z(_GFM_n699 ) );
XOR2_X2 _GFM_U3778  ( .A(_GFM_n708 ), .B(_GFM_n7070 ), .Z(_GFM_n7000 ) );
XOR2_X2 _GFM_U3777  ( .A(z_in[34]), .B(_GFM_n7090 ), .Z(_GFM_n701 ) );
XOR2_X2 _GFM_U3776  ( .A(_GFM_N1081 ), .B(_GFM_N1082 ), .Z(_GFM_n7020 ) );
XOR2_X2 _GFM_U3775  ( .A(_GFM_N1078 ), .B(_GFM_N1079 ), .Z(_GFM_n7030 ) );
XOR2_X2 _GFM_U3774  ( .A(_GFM_N1074 ), .B(_GFM_N1075 ), .Z(_GFM_n704 ) );
XOR2_X2 _GFM_U3773  ( .A(_GFM_N1070 ), .B(_GFM_N1072 ), .Z(_GFM_n705 ) );
XOR2_X2 _GFM_U3772  ( .A(_GFM_N1065 ), .B(_GFM_N1069 ), .Z(_GFM_n7060 ) );
XOR2_X2 _GFM_U3771  ( .A(_GFM_N1062 ), .B(_GFM_N1064 ), .Z(_GFM_n7070 ) );
XOR2_X2 _GFM_U3770  ( .A(_GFM_N1058 ), .B(_GFM_N1061 ), .Z(_GFM_n708 ) );
XOR2_X2 _GFM_U3769  ( .A(_GFM_N1055 ), .B(_GFM_N1057 ), .Z(_GFM_n7090 ) );
XOR2_X2 _GFM_U3768  ( .A(_GFM_n711 ), .B(_GFM_n7100 ), .Z(z_out[35]) );
XOR2_X2 _GFM_U3767  ( .A(_GFM_n713 ), .B(_GFM_n712 ), .Z(_GFM_n7100 ) );
XOR2_X2 _GFM_U3766  ( .A(_GFM_n715 ), .B(_GFM_n7140 ), .Z(_GFM_n711 ) );
XOR2_X2 _GFM_U3765  ( .A(_GFM_n7170 ), .B(_GFM_n7160 ), .Z(_GFM_n712 ) );
XOR2_X2 _GFM_U3764  ( .A(_GFM_n719 ), .B(_GFM_n718 ), .Z(_GFM_n713 ) );
XOR2_X2 _GFM_U3763  ( .A(_GFM_n7210 ), .B(_GFM_n7200 ), .Z(_GFM_n7140 ) );
XOR2_X2 _GFM_U3762  ( .A(_GFM_n7230 ), .B(_GFM_n722 ), .Z(_GFM_n715 ) );
XOR2_X2 _GFM_U3761  ( .A(z_in[35]), .B(_GFM_n7240 ), .Z(_GFM_n7160 ) );
XOR2_X2 _GFM_U3760  ( .A(_GFM_N1112 ), .B(_GFM_N1113 ), .Z(_GFM_n7170 ) );
XOR2_X2 _GFM_U3759  ( .A(_GFM_N1109 ), .B(_GFM_N1110 ), .Z(_GFM_n718 ) );
XOR2_X2 _GFM_U3758  ( .A(_GFM_N1105 ), .B(_GFM_N1106 ), .Z(_GFM_n719 ) );
XOR2_X2 _GFM_U3757  ( .A(_GFM_N1101 ), .B(_GFM_N1103 ), .Z(_GFM_n7200 ) );
XOR2_X2 _GFM_U3756  ( .A(_GFM_N1096 ), .B(_GFM_N1100 ), .Z(_GFM_n7210 ) );
XOR2_X2 _GFM_U3755  ( .A(_GFM_N1093 ), .B(_GFM_N1095 ), .Z(_GFM_n722 ) );
XOR2_X2 _GFM_U3754  ( .A(_GFM_N1089 ), .B(_GFM_N1092 ), .Z(_GFM_n7230 ) );
XOR2_X2 _GFM_U3753  ( .A(_GFM_N1086 ), .B(_GFM_N1088 ), .Z(_GFM_n7240 ) );
XOR2_X2 _GFM_U3752  ( .A(_GFM_n726 ), .B(_GFM_n725 ), .Z(z_out[36]) );
XOR2_X2 _GFM_U3751  ( .A(_GFM_n7280 ), .B(_GFM_n727 ), .Z(_GFM_n725 ) );
XOR2_X2 _GFM_U3750  ( .A(_GFM_n730 ), .B(_GFM_n7290 ), .Z(_GFM_n726 ) );
XOR2_X2 _GFM_U3749  ( .A(_GFM_n732 ), .B(_GFM_n7310 ), .Z(_GFM_n727 ) );
XOR2_X2 _GFM_U3748  ( .A(_GFM_n7340 ), .B(_GFM_n7330 ), .Z(_GFM_n7280 ) );
XOR2_X2 _GFM_U3747  ( .A(_GFM_n736 ), .B(_GFM_n735 ), .Z(_GFM_n7290 ) );
XOR2_X2 _GFM_U3746  ( .A(_GFM_n7380 ), .B(_GFM_n7370 ), .Z(_GFM_n730 ) );
XOR2_X2 _GFM_U3745  ( .A(z_in[36]), .B(_GFM_n739 ), .Z(_GFM_n7310 ) );
XOR2_X2 _GFM_U3744  ( .A(_GFM_N1143 ), .B(_GFM_N1144 ), .Z(_GFM_n732 ) );
XOR2_X2 _GFM_U3743  ( .A(_GFM_N1140 ), .B(_GFM_N1141 ), .Z(_GFM_n7330 ) );
XOR2_X2 _GFM_U3742  ( .A(_GFM_N1136 ), .B(_GFM_N1137 ), .Z(_GFM_n7340 ) );
XOR2_X2 _GFM_U3741  ( .A(_GFM_N1132 ), .B(_GFM_N1134 ), .Z(_GFM_n735 ) );
XOR2_X2 _GFM_U3740  ( .A(_GFM_N1127 ), .B(_GFM_N1131 ), .Z(_GFM_n736 ) );
XOR2_X2 _GFM_U3739  ( .A(_GFM_N1124 ), .B(_GFM_N1126 ), .Z(_GFM_n7370 ) );
XOR2_X2 _GFM_U3738  ( .A(_GFM_N1120 ), .B(_GFM_N1123 ), .Z(_GFM_n7380 ) );
XOR2_X2 _GFM_U3737  ( .A(_GFM_N1117 ), .B(_GFM_N1119 ), .Z(_GFM_n739 ) );
XOR2_X2 _GFM_U3736  ( .A(_GFM_n7410 ), .B(_GFM_n7400 ), .Z(z_out[37]) );
XOR2_X2 _GFM_U3735  ( .A(_GFM_n743 ), .B(_GFM_n742 ), .Z(_GFM_n7400 ) );
XOR2_X2 _GFM_U3734  ( .A(_GFM_n7450 ), .B(_GFM_n744 ), .Z(_GFM_n7410 ) );
XOR2_X2 _GFM_U3733  ( .A(_GFM_n7470 ), .B(_GFM_n746 ), .Z(_GFM_n742 ) );
XOR2_X2 _GFM_U3732  ( .A(_GFM_n749 ), .B(_GFM_n7480 ), .Z(_GFM_n743 ) );
XOR2_X2 _GFM_U3731  ( .A(_GFM_n7510 ), .B(_GFM_n750 ), .Z(_GFM_n744 ) );
XOR2_X2 _GFM_U3730  ( .A(_GFM_n753 ), .B(_GFM_n7520 ), .Z(_GFM_n7450 ) );
XOR2_X2 _GFM_U3729  ( .A(z_in[37]), .B(_GFM_n7540 ), .Z(_GFM_n746 ) );
XOR2_X2 _GFM_U3728  ( .A(_GFM_N1174 ), .B(_GFM_N1175 ), .Z(_GFM_n7470 ) );
XOR2_X2 _GFM_U3727  ( .A(_GFM_N1171 ), .B(_GFM_N1172 ), .Z(_GFM_n7480 ) );
XOR2_X2 _GFM_U3726  ( .A(_GFM_N1167 ), .B(_GFM_N1168 ), .Z(_GFM_n749 ) );
XOR2_X2 _GFM_U3725  ( .A(_GFM_N1163 ), .B(_GFM_N1165 ), .Z(_GFM_n750 ) );
XOR2_X2 _GFM_U3724  ( .A(_GFM_N1158 ), .B(_GFM_N1162 ), .Z(_GFM_n7510 ) );
XOR2_X2 _GFM_U3723  ( .A(_GFM_N1155 ), .B(_GFM_N1157 ), .Z(_GFM_n7520 ) );
XOR2_X2 _GFM_U3722  ( .A(_GFM_N1151 ), .B(_GFM_N1154 ), .Z(_GFM_n753 ) );
XOR2_X2 _GFM_U3721  ( .A(_GFM_N1148 ), .B(_GFM_N1150 ), .Z(_GFM_n7540 ) );
XOR2_X2 _GFM_U3720  ( .A(_GFM_n756 ), .B(_GFM_n7550 ), .Z(z_out[38]) );
XOR2_X2 _GFM_U3719  ( .A(_GFM_n758 ), .B(_GFM_n757 ), .Z(_GFM_n7550 ) );
XOR2_X2 _GFM_U3718  ( .A(_GFM_n7600 ), .B(_GFM_n7590 ), .Z(_GFM_n756 ) );
XOR2_X2 _GFM_U3717  ( .A(_GFM_n7620 ), .B(_GFM_n761 ), .Z(_GFM_n757 ) );
XOR2_X2 _GFM_U3716  ( .A(_GFM_n7640 ), .B(_GFM_n763 ), .Z(_GFM_n758 ) );
XOR2_X2 _GFM_U3715  ( .A(_GFM_n766 ), .B(_GFM_n7650 ), .Z(_GFM_n7590 ) );
XOR2_X2 _GFM_U3714  ( .A(_GFM_n7680 ), .B(_GFM_n767 ), .Z(_GFM_n7600 ) );
XOR2_X2 _GFM_U3713  ( .A(z_in[38]), .B(_GFM_n7690 ), .Z(_GFM_n761 ) );
XOR2_X2 _GFM_U3712  ( .A(_GFM_N1205 ), .B(_GFM_N1206 ), .Z(_GFM_n7620 ) );
XOR2_X2 _GFM_U3711  ( .A(_GFM_N1202 ), .B(_GFM_N1203 ), .Z(_GFM_n763 ) );
XOR2_X2 _GFM_U3710  ( .A(_GFM_N1198 ), .B(_GFM_N1199 ), .Z(_GFM_n7640 ) );
XOR2_X2 _GFM_U3709  ( .A(_GFM_N1194 ), .B(_GFM_N1196 ), .Z(_GFM_n7650 ) );
XOR2_X2 _GFM_U3708  ( .A(_GFM_N1189 ), .B(_GFM_N1193 ), .Z(_GFM_n766 ) );
XOR2_X2 _GFM_U3707  ( .A(_GFM_N1186 ), .B(_GFM_N1188 ), .Z(_GFM_n767 ) );
XOR2_X2 _GFM_U3706  ( .A(_GFM_N1182 ), .B(_GFM_N1185 ), .Z(_GFM_n7680 ) );
XOR2_X2 _GFM_U3705  ( .A(_GFM_N1179 ), .B(_GFM_N1181 ), .Z(_GFM_n7690 ) );
XOR2_X2 _GFM_U3704  ( .A(_GFM_n7710 ), .B(_GFM_n770 ), .Z(z_out[39]) );
XOR2_X2 _GFM_U3703  ( .A(_GFM_n773 ), .B(_GFM_n7720 ), .Z(_GFM_n770 ) );
XOR2_X2 _GFM_U3702  ( .A(_GFM_n775 ), .B(_GFM_n774 ), .Z(_GFM_n7710 ) );
XOR2_X2 _GFM_U3701  ( .A(_GFM_n777 ), .B(_GFM_n7760 ), .Z(_GFM_n7720 ) );
XOR2_X2 _GFM_U3700  ( .A(_GFM_n7790 ), .B(_GFM_n7780 ), .Z(_GFM_n773 ) );
XOR2_X2 _GFM_U3699  ( .A(_GFM_n781 ), .B(_GFM_n780 ), .Z(_GFM_n774 ) );
XOR2_X2 _GFM_U3698  ( .A(_GFM_n7830 ), .B(_GFM_n7820 ), .Z(_GFM_n775 ) );
XOR2_X2 _GFM_U3697  ( .A(z_in[39]), .B(_GFM_n784 ), .Z(_GFM_n7760 ) );
XOR2_X2 _GFM_U3696  ( .A(_GFM_N1236 ), .B(_GFM_N1237 ), .Z(_GFM_n777 ) );
XOR2_X2 _GFM_U3695  ( .A(_GFM_N1233 ), .B(_GFM_N1234 ), .Z(_GFM_n7780 ) );
XOR2_X2 _GFM_U3694  ( .A(_GFM_N1229 ), .B(_GFM_N1230 ), .Z(_GFM_n7790 ) );
XOR2_X2 _GFM_U3693  ( .A(_GFM_N1225 ), .B(_GFM_N1227 ), .Z(_GFM_n780 ) );
XOR2_X2 _GFM_U3692  ( .A(_GFM_N1220 ), .B(_GFM_N1224 ), .Z(_GFM_n781 ) );
XOR2_X2 _GFM_U3691  ( .A(_GFM_N1217 ), .B(_GFM_N1219 ), .Z(_GFM_n7820 ) );
XOR2_X2 _GFM_U3690  ( .A(_GFM_N1213 ), .B(_GFM_N1216 ), .Z(_GFM_n7830 ) );
XOR2_X2 _GFM_U3689  ( .A(_GFM_N1210 ), .B(_GFM_N1212 ), .Z(_GFM_n784 ) );
XOR2_X2 _GFM_U3688  ( .A(_GFM_n7860 ), .B(_GFM_n7850 ), .Z(z_out[40]) );
XOR2_X2 _GFM_U3687  ( .A(_GFM_n788 ), .B(_GFM_n787 ), .Z(_GFM_n7850 ) );
XOR2_X2 _GFM_U3686  ( .A(_GFM_n7900 ), .B(_GFM_n789 ), .Z(_GFM_n7860 ) );
XOR2_X2 _GFM_U3685  ( .A(_GFM_n792 ), .B(_GFM_n7910 ), .Z(_GFM_n787 ) );
XOR2_X2 _GFM_U3684  ( .A(_GFM_n794 ), .B(_GFM_n7930 ), .Z(_GFM_n788 ) );
XOR2_X2 _GFM_U3683  ( .A(_GFM_n7960 ), .B(_GFM_n7950 ), .Z(_GFM_n789 ) );
XOR2_X2 _GFM_U3682  ( .A(_GFM_n798 ), .B(_GFM_n797 ), .Z(_GFM_n7900 ) );
XOR2_X2 _GFM_U3681  ( .A(z_in[40]), .B(_GFM_n7990 ), .Z(_GFM_n7910 ) );
XOR2_X2 _GFM_U3680  ( .A(_GFM_N1267 ), .B(_GFM_N1268 ), .Z(_GFM_n792 ) );
XOR2_X2 _GFM_U3679  ( .A(_GFM_N1264 ), .B(_GFM_N1265 ), .Z(_GFM_n7930 ) );
XOR2_X2 _GFM_U3678  ( .A(_GFM_N1260 ), .B(_GFM_N1261 ), .Z(_GFM_n794 ) );
XOR2_X2 _GFM_U3677  ( .A(_GFM_N1256 ), .B(_GFM_N1258 ), .Z(_GFM_n7950 ) );
XOR2_X2 _GFM_U3676  ( .A(_GFM_N1251 ), .B(_GFM_N1255 ), .Z(_GFM_n7960 ) );
XOR2_X2 _GFM_U3675  ( .A(_GFM_N1248 ), .B(_GFM_N1250 ), .Z(_GFM_n797 ) );
XOR2_X2 _GFM_U3674  ( .A(_GFM_N1244 ), .B(_GFM_N1247 ), .Z(_GFM_n798 ) );
XOR2_X2 _GFM_U3673  ( .A(_GFM_N1241 ), .B(_GFM_N1243 ), .Z(_GFM_n7990 ) );
XOR2_X2 _GFM_U3672  ( .A(_GFM_n801 ), .B(_GFM_n8000 ), .Z(z_out[41]) );
XOR2_X2 _GFM_U3671  ( .A(_GFM_n8030 ), .B(_GFM_n8020 ), .Z(_GFM_n8000 ) );
XOR2_X2 _GFM_U3670  ( .A(_GFM_n805 ), .B(_GFM_n804 ), .Z(_GFM_n801 ) );
XOR2_X2 _GFM_U3669  ( .A(_GFM_n8070 ), .B(_GFM_n806 ), .Z(_GFM_n8020 ) );
XOR2_X2 _GFM_U3668  ( .A(_GFM_n8090 ), .B(_GFM_n808 ), .Z(_GFM_n8030 ) );
XOR2_X2 _GFM_U3667  ( .A(_GFM_n811 ), .B(_GFM_n8100 ), .Z(_GFM_n804 ) );
XOR2_X2 _GFM_U3666  ( .A(_GFM_n8130 ), .B(_GFM_n812 ), .Z(_GFM_n805 ) );
XOR2_X2 _GFM_U3665  ( .A(z_in[41]), .B(_GFM_n8140 ), .Z(_GFM_n806 ) );
XOR2_X2 _GFM_U3664  ( .A(_GFM_N1298 ), .B(_GFM_N1299 ), .Z(_GFM_n8070 ) );
XOR2_X2 _GFM_U3663  ( .A(_GFM_N1295 ), .B(_GFM_N1296 ), .Z(_GFM_n808 ) );
XOR2_X2 _GFM_U3662  ( .A(_GFM_N1291 ), .B(_GFM_N1292 ), .Z(_GFM_n8090 ) );
XOR2_X2 _GFM_U3661  ( .A(_GFM_N1287 ), .B(_GFM_N1289 ), .Z(_GFM_n8100 ) );
XOR2_X2 _GFM_U3660  ( .A(_GFM_N1282 ), .B(_GFM_N1286 ), .Z(_GFM_n811 ) );
XOR2_X2 _GFM_U3659  ( .A(_GFM_N1279 ), .B(_GFM_N1281 ), .Z(_GFM_n812 ) );
XOR2_X2 _GFM_U3658  ( .A(_GFM_N1275 ), .B(_GFM_N1278 ), .Z(_GFM_n8130 ) );
XOR2_X2 _GFM_U3657  ( .A(_GFM_N1272 ), .B(_GFM_N1274 ), .Z(_GFM_n8140 ) );
XOR2_X2 _GFM_U3656  ( .A(_GFM_n8160 ), .B(_GFM_n815 ), .Z(z_out[42]) );
XOR2_X2 _GFM_U3655  ( .A(_GFM_n818 ), .B(_GFM_n8170 ), .Z(_GFM_n815 ) );
XOR2_X2 _GFM_U3654  ( .A(_GFM_n820 ), .B(_GFM_n819 ), .Z(_GFM_n8160 ) );
XOR2_X2 _GFM_U3653  ( .A(_GFM_n8220 ), .B(_GFM_n8210 ), .Z(_GFM_n8170 ) );
XOR2_X2 _GFM_U3652  ( .A(_GFM_n8240 ), .B(_GFM_n823 ), .Z(_GFM_n818 ) );
XOR2_X2 _GFM_U3651  ( .A(_GFM_n8260 ), .B(_GFM_n825 ), .Z(_GFM_n819 ) );
XOR2_X2 _GFM_U3650  ( .A(_GFM_n828 ), .B(_GFM_n8270 ), .Z(_GFM_n820 ) );
XOR2_X2 _GFM_U3649  ( .A(z_in[42]), .B(_GFM_n829 ), .Z(_GFM_n8210 ) );
XOR2_X2 _GFM_U3648  ( .A(_GFM_N1329 ), .B(_GFM_N1330 ), .Z(_GFM_n8220 ) );
XOR2_X2 _GFM_U3647  ( .A(_GFM_N1326 ), .B(_GFM_N1327 ), .Z(_GFM_n823 ) );
XOR2_X2 _GFM_U3646  ( .A(_GFM_N1322 ), .B(_GFM_N1323 ), .Z(_GFM_n8240 ) );
XOR2_X2 _GFM_U3645  ( .A(_GFM_N1318 ), .B(_GFM_N1320 ), .Z(_GFM_n825 ) );
XOR2_X2 _GFM_U3644  ( .A(_GFM_N1313 ), .B(_GFM_N1317 ), .Z(_GFM_n8260 ) );
XOR2_X2 _GFM_U3643  ( .A(_GFM_N1310 ), .B(_GFM_N1312 ), .Z(_GFM_n8270 ) );
XOR2_X2 _GFM_U3642  ( .A(_GFM_N1306 ), .B(_GFM_N1309 ), .Z(_GFM_n828 ) );
XOR2_X2 _GFM_U3641  ( .A(_GFM_N1303 ), .B(_GFM_N1305 ), .Z(_GFM_n829 ) );
XOR2_X2 _GFM_U3640  ( .A(_GFM_n8310 ), .B(_GFM_n8300 ), .Z(z_out[43]) );
XOR2_X2 _GFM_U3639  ( .A(_GFM_n8330 ), .B(_GFM_n832 ), .Z(_GFM_n8300 ) );
XOR2_X2 _GFM_U3638  ( .A(_GFM_n835 ), .B(_GFM_n8340 ), .Z(_GFM_n8310 ) );
XOR2_X2 _GFM_U3637  ( .A(_GFM_n837 ), .B(_GFM_n836 ), .Z(_GFM_n832 ) );
XOR2_X2 _GFM_U3636  ( .A(_GFM_n839 ), .B(_GFM_n8380 ), .Z(_GFM_n8330 ) );
XOR2_X2 _GFM_U3635  ( .A(_GFM_n8410 ), .B(_GFM_n8400 ), .Z(_GFM_n8340 ) );
XOR2_X2 _GFM_U3634  ( .A(_GFM_n843 ), .B(_GFM_n842 ), .Z(_GFM_n835 ) );
XOR2_X2 _GFM_U3633  ( .A(z_in[43]), .B(_GFM_n8440 ), .Z(_GFM_n836 ) );
XOR2_X2 _GFM_U3632  ( .A(_GFM_N1360 ), .B(_GFM_N1361 ), .Z(_GFM_n837 ) );
XOR2_X2 _GFM_U3631  ( .A(_GFM_N1357 ), .B(_GFM_N1358 ), .Z(_GFM_n8380 ) );
XOR2_X2 _GFM_U3630  ( .A(_GFM_N1353 ), .B(_GFM_N1354 ), .Z(_GFM_n839 ) );
XOR2_X2 _GFM_U3629  ( .A(_GFM_N1349 ), .B(_GFM_N1351 ), .Z(_GFM_n8400 ) );
XOR2_X2 _GFM_U3628  ( .A(_GFM_N1344 ), .B(_GFM_N1348 ), .Z(_GFM_n8410 ) );
XOR2_X2 _GFM_U3627  ( .A(_GFM_N1341 ), .B(_GFM_N1343 ), .Z(_GFM_n842 ) );
XOR2_X2 _GFM_U3626  ( .A(_GFM_N1337 ), .B(_GFM_N1340 ), .Z(_GFM_n843 ) );
XOR2_X2 _GFM_U3625  ( .A(_GFM_N1334 ), .B(_GFM_N1336 ), .Z(_GFM_n8440 ) );
XOR2_X2 _GFM_U3624  ( .A(_GFM_n846 ), .B(_GFM_n8450 ), .Z(z_out[44]) );
XOR2_X2 _GFM_U3623  ( .A(_GFM_n8480 ), .B(_GFM_n8470 ), .Z(_GFM_n8450 ) );
XOR2_X2 _GFM_U3622  ( .A(_GFM_n850 ), .B(_GFM_n849 ), .Z(_GFM_n846 ) );
XOR2_X2 _GFM_U3621  ( .A(_GFM_n8520 ), .B(_GFM_n851 ), .Z(_GFM_n8470 ) );
XOR2_X2 _GFM_U3620  ( .A(_GFM_n854 ), .B(_GFM_n8530 ), .Z(_GFM_n8480 ) );
XOR2_X2 _GFM_U3619  ( .A(_GFM_n856 ), .B(_GFM_n8550 ), .Z(_GFM_n849 ) );
XOR2_X2 _GFM_U3618  ( .A(_GFM_n8580 ), .B(_GFM_n8570 ), .Z(_GFM_n850 ) );
XOR2_X2 _GFM_U3617  ( .A(z_in[44]), .B(_GFM_n859 ), .Z(_GFM_n851 ) );
XOR2_X2 _GFM_U3616  ( .A(_GFM_N1391 ), .B(_GFM_N1392 ), .Z(_GFM_n8520 ) );
XOR2_X2 _GFM_U3615  ( .A(_GFM_N1388 ), .B(_GFM_N1389 ), .Z(_GFM_n8530 ) );
XOR2_X2 _GFM_U3614  ( .A(_GFM_N1384 ), .B(_GFM_N1385 ), .Z(_GFM_n854 ) );
XOR2_X2 _GFM_U3613  ( .A(_GFM_N1380 ), .B(_GFM_N1382 ), .Z(_GFM_n8550 ) );
XOR2_X2 _GFM_U3612  ( .A(_GFM_N1375 ), .B(_GFM_N1379 ), .Z(_GFM_n856 ) );
XOR2_X2 _GFM_U3611  ( .A(_GFM_N1372 ), .B(_GFM_N1374 ), .Z(_GFM_n8570 ) );
XOR2_X2 _GFM_U3610  ( .A(_GFM_N1368 ), .B(_GFM_N1371 ), .Z(_GFM_n8580 ) );
XOR2_X2 _GFM_U3609  ( .A(_GFM_N1365 ), .B(_GFM_N1367 ), .Z(_GFM_n859 ) );
XOR2_X2 _GFM_U3608  ( .A(_GFM_n8610 ), .B(_GFM_n860 ), .Z(z_out[45]) );
XOR2_X2 _GFM_U3607  ( .A(_GFM_n863 ), .B(_GFM_n8620 ), .Z(_GFM_n860 ) );
XOR2_X2 _GFM_U3606  ( .A(_GFM_n8650 ), .B(_GFM_n8640 ), .Z(_GFM_n8610 ) );
XOR2_X2 _GFM_U3605  ( .A(_GFM_n867 ), .B(_GFM_n866 ), .Z(_GFM_n8620 ) );
XOR2_X2 _GFM_U3604  ( .A(_GFM_n8690 ), .B(_GFM_n868 ), .Z(_GFM_n863 ) );
XOR2_X2 _GFM_U3603  ( .A(_GFM_n8710 ), .B(_GFM_n870 ), .Z(_GFM_n8640 ) );
XOR2_X2 _GFM_U3602  ( .A(_GFM_n873 ), .B(_GFM_n8720 ), .Z(_GFM_n8650 ) );
XOR2_X2 _GFM_U3601  ( .A(z_in[45]), .B(_GFM_n874 ), .Z(_GFM_n866 ) );
XOR2_X2 _GFM_U3600  ( .A(_GFM_N1422 ), .B(_GFM_N1423 ), .Z(_GFM_n867 ) );
XOR2_X2 _GFM_U3599  ( .A(_GFM_N1419 ), .B(_GFM_N1420 ), .Z(_GFM_n868 ) );
XOR2_X2 _GFM_U3598  ( .A(_GFM_N1415 ), .B(_GFM_N1416 ), .Z(_GFM_n8690 ) );
XOR2_X2 _GFM_U3597  ( .A(_GFM_N1411 ), .B(_GFM_N1413 ), .Z(_GFM_n870 ) );
XOR2_X2 _GFM_U3596  ( .A(_GFM_N1406 ), .B(_GFM_N1410 ), .Z(_GFM_n8710 ) );
XOR2_X2 _GFM_U3595  ( .A(_GFM_N1403 ), .B(_GFM_N1405 ), .Z(_GFM_n8720 ) );
XOR2_X2 _GFM_U3594  ( .A(_GFM_N1399 ), .B(_GFM_N1402 ), .Z(_GFM_n873 ) );
XOR2_X2 _GFM_U3593  ( .A(_GFM_N1396 ), .B(_GFM_N1398 ), .Z(_GFM_n874 ) );
XOR2_X2 _GFM_U3592  ( .A(_GFM_n8760 ), .B(_GFM_n8750 ), .Z(z_out[46]) );
XOR2_X2 _GFM_U3591  ( .A(_GFM_n8780 ), .B(_GFM_n877 ), .Z(_GFM_n8750 ) );
XOR2_X2 _GFM_U3590  ( .A(_GFM_n880 ), .B(_GFM_n8790 ), .Z(_GFM_n8760 ) );
XOR2_X2 _GFM_U3589  ( .A(_GFM_n882 ), .B(_GFM_n881 ), .Z(_GFM_n877 ) );
XOR2_X2 _GFM_U3588  ( .A(_GFM_n8840 ), .B(_GFM_n8830 ), .Z(_GFM_n8780 ) );
XOR2_X2 _GFM_U3587  ( .A(_GFM_n8860 ), .B(_GFM_n885 ), .Z(_GFM_n8790 ) );
XOR2_X2 _GFM_U3586  ( .A(_GFM_n8880 ), .B(_GFM_n887 ), .Z(_GFM_n880 ) );
XOR2_X2 _GFM_U3585  ( .A(z_in[46]), .B(_GFM_n8890 ), .Z(_GFM_n881 ) );
XOR2_X2 _GFM_U3584  ( .A(_GFM_N1453 ), .B(_GFM_N1454 ), .Z(_GFM_n882 ) );
XOR2_X2 _GFM_U3583  ( .A(_GFM_N1450 ), .B(_GFM_N1451 ), .Z(_GFM_n8830 ) );
XOR2_X2 _GFM_U3582  ( .A(_GFM_N1446 ), .B(_GFM_N1447 ), .Z(_GFM_n8840 ) );
XOR2_X2 _GFM_U3581  ( .A(_GFM_N1442 ), .B(_GFM_N1444 ), .Z(_GFM_n885 ) );
XOR2_X2 _GFM_U3580  ( .A(_GFM_N1437 ), .B(_GFM_N1441 ), .Z(_GFM_n8860 ) );
XOR2_X2 _GFM_U3579  ( .A(_GFM_N1434 ), .B(_GFM_N1436 ), .Z(_GFM_n887 ) );
XOR2_X2 _GFM_U3578  ( .A(_GFM_N1430 ), .B(_GFM_N1433 ), .Z(_GFM_n8880 ) );
XOR2_X2 _GFM_U3577  ( .A(_GFM_N1427 ), .B(_GFM_N1429 ), .Z(_GFM_n8890 ) );
XOR2_X2 _GFM_U3576  ( .A(_GFM_n891 ), .B(_GFM_n890 ), .Z(z_out[47]) );
XOR2_X2 _GFM_U3575  ( .A(_GFM_n8930 ), .B(_GFM_n8920 ), .Z(_GFM_n890 ) );
XOR2_X2 _GFM_U3574  ( .A(_GFM_n8950 ), .B(_GFM_n894 ), .Z(_GFM_n891 ) );
XOR2_X2 _GFM_U3573  ( .A(_GFM_n897 ), .B(_GFM_n8960 ), .Z(_GFM_n8920 ) );
XOR2_X2 _GFM_U3572  ( .A(_GFM_n899 ), .B(_GFM_n898 ), .Z(_GFM_n8930 ) );
XOR2_X2 _GFM_U3571  ( .A(_GFM_n901 ), .B(_GFM_n9000 ), .Z(_GFM_n894 ) );
XOR2_X2 _GFM_U3570  ( .A(_GFM_n9030 ), .B(_GFM_n9020 ), .Z(_GFM_n8950 ) );
XOR2_X2 _GFM_U3569  ( .A(z_in[47]), .B(_GFM_n904 ), .Z(_GFM_n8960 ) );
XOR2_X2 _GFM_U3568  ( .A(_GFM_N1484 ), .B(_GFM_N1485 ), .Z(_GFM_n897 ) );
XOR2_X2 _GFM_U3567  ( .A(_GFM_N1481 ), .B(_GFM_N1482 ), .Z(_GFM_n898 ) );
XOR2_X2 _GFM_U3566  ( .A(_GFM_N1477 ), .B(_GFM_N1478 ), .Z(_GFM_n899 ) );
XOR2_X2 _GFM_U3565  ( .A(_GFM_N1473 ), .B(_GFM_N1475 ), .Z(_GFM_n9000 ) );
XOR2_X2 _GFM_U3564  ( .A(_GFM_N1468 ), .B(_GFM_N1472 ), .Z(_GFM_n901 ) );
XOR2_X2 _GFM_U3563  ( .A(_GFM_N1465 ), .B(_GFM_N1467 ), .Z(_GFM_n9020 ) );
XOR2_X2 _GFM_U3562  ( .A(_GFM_N1461 ), .B(_GFM_N1464 ), .Z(_GFM_n9030 ) );
XOR2_X2 _GFM_U3561  ( .A(_GFM_N1458 ), .B(_GFM_N1460 ), .Z(_GFM_n904 ) );
XOR2_X2 _GFM_U3560  ( .A(_GFM_n9060 ), .B(_GFM_n905 ), .Z(z_out[48]) );
XOR2_X2 _GFM_U3559  ( .A(_GFM_n908 ), .B(_GFM_n9070 ), .Z(_GFM_n905 ) );
XOR2_X2 _GFM_U3558  ( .A(_GFM_n9100 ), .B(_GFM_n9090 ), .Z(_GFM_n9060 ) );
XOR2_X2 _GFM_U3557  ( .A(_GFM_n912 ), .B(_GFM_n911 ), .Z(_GFM_n9070 ) );
XOR2_X2 _GFM_U3556  ( .A(_GFM_n9140 ), .B(_GFM_n913 ), .Z(_GFM_n908 ) );
XOR2_X2 _GFM_U3555  ( .A(_GFM_n916 ), .B(_GFM_n9150 ), .Z(_GFM_n9090 ) );
XOR2_X2 _GFM_U3554  ( .A(_GFM_n918 ), .B(_GFM_n9170 ), .Z(_GFM_n9100 ) );
XOR2_X2 _GFM_U3553  ( .A(z_in[48]), .B(_GFM_n9190 ), .Z(_GFM_n911 ) );
XOR2_X2 _GFM_U3552  ( .A(_GFM_N1515 ), .B(_GFM_N1516 ), .Z(_GFM_n912 ) );
XOR2_X2 _GFM_U3551  ( .A(_GFM_N1512 ), .B(_GFM_N1513 ), .Z(_GFM_n913 ) );
XOR2_X2 _GFM_U3550  ( .A(_GFM_N1508 ), .B(_GFM_N1509 ), .Z(_GFM_n9140 ) );
XOR2_X2 _GFM_U3549  ( .A(_GFM_N1504 ), .B(_GFM_N1506 ), .Z(_GFM_n9150 ) );
XOR2_X2 _GFM_U3548  ( .A(_GFM_N1499 ), .B(_GFM_N1503 ), .Z(_GFM_n916 ) );
XOR2_X2 _GFM_U3547  ( .A(_GFM_N1496 ), .B(_GFM_N1498 ), .Z(_GFM_n9170 ) );
XOR2_X2 _GFM_U3546  ( .A(_GFM_N1492 ), .B(_GFM_N1495 ), .Z(_GFM_n918 ) );
XOR2_X2 _GFM_U3545  ( .A(_GFM_N1489 ), .B(_GFM_N1491 ), .Z(_GFM_n9190 ) );
XOR2_X2 _GFM_U3544  ( .A(_GFM_n921 ), .B(_GFM_n9200 ), .Z(z_out[49]) );
XOR2_X2 _GFM_U3543  ( .A(_GFM_n9230 ), .B(_GFM_n922 ), .Z(_GFM_n9200 ) );
XOR2_X2 _GFM_U3542  ( .A(_GFM_n925 ), .B(_GFM_n9240 ), .Z(_GFM_n921 ) );
XOR2_X2 _GFM_U3541  ( .A(_GFM_n9270 ), .B(_GFM_n9260 ), .Z(_GFM_n922 ) );
XOR2_X2 _GFM_U3540  ( .A(_GFM_n929 ), .B(_GFM_n928 ), .Z(_GFM_n9230 ) );
XOR2_X2 _GFM_U3539  ( .A(_GFM_n9310 ), .B(_GFM_n930 ), .Z(_GFM_n9240 ) );
XOR2_X2 _GFM_U3538  ( .A(_GFM_n9330 ), .B(_GFM_n932 ), .Z(_GFM_n925 ) );
XOR2_X2 _GFM_U3537  ( .A(z_in[49]), .B(_GFM_n9340 ), .Z(_GFM_n9260 ) );
XOR2_X2 _GFM_U3536  ( .A(_GFM_N1546 ), .B(_GFM_N1547 ), .Z(_GFM_n9270 ) );
XOR2_X2 _GFM_U3535  ( .A(_GFM_N1543 ), .B(_GFM_N1544 ), .Z(_GFM_n928 ) );
XOR2_X2 _GFM_U3534  ( .A(_GFM_N1539 ), .B(_GFM_N1540 ), .Z(_GFM_n929 ) );
XOR2_X2 _GFM_U3533  ( .A(_GFM_N1535 ), .B(_GFM_N1537 ), .Z(_GFM_n930 ) );
XOR2_X2 _GFM_U3532  ( .A(_GFM_N1530 ), .B(_GFM_N1534 ), .Z(_GFM_n9310 ) );
XOR2_X2 _GFM_U3531  ( .A(_GFM_N1527 ), .B(_GFM_N1529 ), .Z(_GFM_n932 ) );
XOR2_X2 _GFM_U3530  ( .A(_GFM_N1523 ), .B(_GFM_N1526 ), .Z(_GFM_n9330 ) );
XOR2_X2 _GFM_U3529  ( .A(_GFM_N1520 ), .B(_GFM_N1522 ), .Z(_GFM_n9340 ) );
XOR2_X2 _GFM_U3528  ( .A(_GFM_n936 ), .B(_GFM_n935 ), .Z(z_out[50]) );
XOR2_X2 _GFM_U3527  ( .A(_GFM_n9380 ), .B(_GFM_n9370 ), .Z(_GFM_n935 ) );
XOR2_X2 _GFM_U3526  ( .A(_GFM_n9400 ), .B(_GFM_n939 ), .Z(_GFM_n936 ) );
XOR2_X2 _GFM_U3525  ( .A(_GFM_n942 ), .B(_GFM_n9410 ), .Z(_GFM_n9370 ) );
XOR2_X2 _GFM_U3524  ( .A(_GFM_n944 ), .B(_GFM_n943 ), .Z(_GFM_n9380 ) );
XOR2_X2 _GFM_U3523  ( .A(_GFM_n9460 ), .B(_GFM_n9450 ), .Z(_GFM_n939 ) );
XOR2_X2 _GFM_U3522  ( .A(_GFM_n9480 ), .B(_GFM_n947 ), .Z(_GFM_n9400 ) );
XOR2_X2 _GFM_U3521  ( .A(z_in[50]), .B(_GFM_n949 ), .Z(_GFM_n9410 ) );
XOR2_X2 _GFM_U3520  ( .A(_GFM_N1577 ), .B(_GFM_N1578 ), .Z(_GFM_n942 ) );
XOR2_X2 _GFM_U3519  ( .A(_GFM_N1574 ), .B(_GFM_N1575 ), .Z(_GFM_n943 ) );
XOR2_X2 _GFM_U3518  ( .A(_GFM_N1570 ), .B(_GFM_N1571 ), .Z(_GFM_n944 ) );
XOR2_X2 _GFM_U3517  ( .A(_GFM_N1566 ), .B(_GFM_N1568 ), .Z(_GFM_n9450 ) );
XOR2_X2 _GFM_U3516  ( .A(_GFM_N1561 ), .B(_GFM_N1565 ), .Z(_GFM_n9460 ) );
XOR2_X2 _GFM_U3515  ( .A(_GFM_N1558 ), .B(_GFM_N1560 ), .Z(_GFM_n947 ) );
XOR2_X2 _GFM_U3514  ( .A(_GFM_N1554 ), .B(_GFM_N1557 ), .Z(_GFM_n9480 ) );
XOR2_X2 _GFM_U3513  ( .A(_GFM_N1551 ), .B(_GFM_N1553 ), .Z(_GFM_n949 ) );
XOR2_X2 _GFM_U3512  ( .A(_GFM_n9510 ), .B(_GFM_n9500 ), .Z(z_out[51]) );
XOR2_X2 _GFM_U3511  ( .A(_GFM_n953 ), .B(_GFM_n952 ), .Z(_GFM_n9500 ) );
XOR2_X2 _GFM_U3510  ( .A(_GFM_n9550 ), .B(_GFM_n9540 ), .Z(_GFM_n9510 ) );
XOR2_X2 _GFM_U3509  ( .A(_GFM_n9570 ), .B(_GFM_n956 ), .Z(_GFM_n952 ) );
XOR2_X2 _GFM_U3508  ( .A(_GFM_n959 ), .B(_GFM_n9580 ), .Z(_GFM_n953 ) );
XOR2_X2 _GFM_U3507  ( .A(_GFM_n961 ), .B(_GFM_n960 ), .Z(_GFM_n9540 ) );
XOR2_X2 _GFM_U3506  ( .A(_GFM_n963 ), .B(_GFM_n9620 ), .Z(_GFM_n9550 ) );
XOR2_X2 _GFM_U3505  ( .A(z_in[51]), .B(_GFM_n9640 ), .Z(_GFM_n956 ) );
XOR2_X2 _GFM_U3504  ( .A(_GFM_N1608 ), .B(_GFM_N1609 ), .Z(_GFM_n9570 ) );
XOR2_X2 _GFM_U3503  ( .A(_GFM_N1605 ), .B(_GFM_N1606 ), .Z(_GFM_n9580 ) );
XOR2_X2 _GFM_U3502  ( .A(_GFM_N1601 ), .B(_GFM_N1602 ), .Z(_GFM_n959 ) );
XOR2_X2 _GFM_U3501  ( .A(_GFM_N1597 ), .B(_GFM_N1599 ), .Z(_GFM_n960 ) );
XOR2_X2 _GFM_U3500  ( .A(_GFM_N1592 ), .B(_GFM_N1596 ), .Z(_GFM_n961 ) );
XOR2_X2 _GFM_U3499  ( .A(_GFM_N1589 ), .B(_GFM_N1591 ), .Z(_GFM_n9620 ) );
XOR2_X2 _GFM_U3498  ( .A(_GFM_N1585 ), .B(_GFM_N1588 ), .Z(_GFM_n963 ) );
XOR2_X2 _GFM_U3497  ( .A(_GFM_N1582 ), .B(_GFM_N1584 ), .Z(_GFM_n9640 ) );
XOR2_X2 _GFM_U3496  ( .A(_GFM_n966 ), .B(_GFM_n9650 ), .Z(z_out[52]) );
XOR2_X2 _GFM_U3495  ( .A(_GFM_n9680 ), .B(_GFM_n967 ), .Z(_GFM_n9650 ) );
XOR2_X2 _GFM_U3494  ( .A(_GFM_n970 ), .B(_GFM_n9690 ), .Z(_GFM_n966 ) );
XOR2_X2 _GFM_U3493  ( .A(_GFM_n9720 ), .B(_GFM_n9710 ), .Z(_GFM_n967 ) );
XOR2_X2 _GFM_U3492  ( .A(_GFM_n974 ), .B(_GFM_n973 ), .Z(_GFM_n9680 ) );
XOR2_X2 _GFM_U3491  ( .A(_GFM_n9760 ), .B(_GFM_n975 ), .Z(_GFM_n9690 ) );
XOR2_X2 _GFM_U3490  ( .A(_GFM_n978 ), .B(_GFM_n9770 ), .Z(_GFM_n970 ) );
XOR2_X2 _GFM_U3489  ( .A(z_in[52]), .B(_GFM_n9790 ), .Z(_GFM_n9710 ) );
XOR2_X2 _GFM_U3488  ( .A(_GFM_N1639 ), .B(_GFM_N1640 ), .Z(_GFM_n9720 ) );
XOR2_X2 _GFM_U3487  ( .A(_GFM_N1636 ), .B(_GFM_N1637 ), .Z(_GFM_n973 ) );
XOR2_X2 _GFM_U3486  ( .A(_GFM_N1632 ), .B(_GFM_N1633 ), .Z(_GFM_n974 ) );
XOR2_X2 _GFM_U3485  ( .A(_GFM_N1628 ), .B(_GFM_N1630 ), .Z(_GFM_n975 ) );
XOR2_X2 _GFM_U3484  ( .A(_GFM_N1623 ), .B(_GFM_N1627 ), .Z(_GFM_n9760 ) );
XOR2_X2 _GFM_U3483  ( .A(_GFM_N1620 ), .B(_GFM_N1622 ), .Z(_GFM_n9770 ) );
XOR2_X2 _GFM_U3482  ( .A(_GFM_N1616 ), .B(_GFM_N1619 ), .Z(_GFM_n978 ) );
XOR2_X2 _GFM_U3481  ( .A(_GFM_N1613 ), .B(_GFM_N1615 ), .Z(_GFM_n9790 ) );
XOR2_X2 _GFM_U3480  ( .A(_GFM_n9810 ), .B(_GFM_n980 ), .Z(z_out[53]) );
XOR2_X2 _GFM_U3479  ( .A(_GFM_n983 ), .B(_GFM_n9820 ), .Z(_GFM_n980 ) );
XOR2_X2 _GFM_U3478  ( .A(_GFM_n9850 ), .B(_GFM_n984 ), .Z(_GFM_n9810 ) );
XOR2_X2 _GFM_U3477  ( .A(_GFM_n987 ), .B(_GFM_n9860 ), .Z(_GFM_n9820 ) );
XOR2_X2 _GFM_U3476  ( .A(_GFM_n9890 ), .B(_GFM_n9880 ), .Z(_GFM_n983 ) );
XOR2_X2 _GFM_U3475  ( .A(_GFM_n991 ), .B(_GFM_n990 ), .Z(_GFM_n984 ) );
XOR2_X2 _GFM_U3474  ( .A(_GFM_n9930 ), .B(_GFM_n992 ), .Z(_GFM_n9850 ) );
XOR2_X2 _GFM_U3473  ( .A(z_in[53]), .B(_GFM_n994 ), .Z(_GFM_n9860 ) );
XOR2_X2 _GFM_U3472  ( .A(_GFM_N1670 ), .B(_GFM_N1671 ), .Z(_GFM_n987 ) );
XOR2_X2 _GFM_U3471  ( .A(_GFM_N1667 ), .B(_GFM_N1668 ), .Z(_GFM_n9880 ) );
XOR2_X2 _GFM_U3470  ( .A(_GFM_N1663 ), .B(_GFM_N1664 ), .Z(_GFM_n9890 ) );
XOR2_X2 _GFM_U3469  ( .A(_GFM_N1659 ), .B(_GFM_N1661 ), .Z(_GFM_n990 ) );
XOR2_X2 _GFM_U3468  ( .A(_GFM_N1654 ), .B(_GFM_N1658 ), .Z(_GFM_n991 ) );
XOR2_X2 _GFM_U3467  ( .A(_GFM_N1651 ), .B(_GFM_N1653 ), .Z(_GFM_n992 ) );
XOR2_X2 _GFM_U3466  ( .A(_GFM_N1647 ), .B(_GFM_N1650 ), .Z(_GFM_n9930 ) );
XOR2_X2 _GFM_U3465  ( .A(_GFM_N1644 ), .B(_GFM_N1646 ), .Z(_GFM_n994 ) );
XOR2_X2 _GFM_U3464  ( .A(_GFM_n9960 ), .B(_GFM_n9950 ), .Z(z_out[54]) );
XOR2_X2 _GFM_U3463  ( .A(_GFM_n998 ), .B(_GFM_n997 ), .Z(_GFM_n9950 ) );
XOR2_X2 _GFM_U3462  ( .A(_GFM_n10000 ), .B(_GFM_n9990 ), .Z(_GFM_n9960 ) );
XOR2_X2 _GFM_U3461  ( .A(_GFM_n10020 ), .B(_GFM_n1001 ), .Z(_GFM_n997 ) );
XOR2_X2 _GFM_U3460  ( .A(_GFM_n1004 ), .B(_GFM_n10030 ), .Z(_GFM_n998 ) );
XOR2_X2 _GFM_U3459  ( .A(_GFM_n1006 ), .B(_GFM_n1005 ), .Z(_GFM_n9990 ) );
XOR2_X2 _GFM_U3458  ( .A(_GFM_n10080 ), .B(_GFM_n10070 ), .Z(_GFM_n10000 ));
XOR2_X2 _GFM_U3457  ( .A(z_in[54]), .B(_GFM_n1009 ), .Z(_GFM_n1001 ) );
XOR2_X2 _GFM_U3456  ( .A(_GFM_N1701 ), .B(_GFM_N1702 ), .Z(_GFM_n10020 ) );
XOR2_X2 _GFM_U3455  ( .A(_GFM_N1698 ), .B(_GFM_N1699 ), .Z(_GFM_n10030 ) );
XOR2_X2 _GFM_U3454  ( .A(_GFM_N1694 ), .B(_GFM_N1695 ), .Z(_GFM_n1004 ) );
XOR2_X2 _GFM_U3453  ( .A(_GFM_N1690 ), .B(_GFM_N1692 ), .Z(_GFM_n1005 ) );
XOR2_X2 _GFM_U3452  ( .A(_GFM_N1685 ), .B(_GFM_N1689 ), .Z(_GFM_n1006 ) );
XOR2_X2 _GFM_U3451  ( .A(_GFM_N1682 ), .B(_GFM_N1684 ), .Z(_GFM_n10070 ) );
XOR2_X2 _GFM_U3450  ( .A(_GFM_N1678 ), .B(_GFM_N1681 ), .Z(_GFM_n10080 ) );
XOR2_X2 _GFM_U3449  ( .A(_GFM_N1675 ), .B(_GFM_N1677 ), .Z(_GFM_n1009 ) );
XOR2_X2 _GFM_U3448  ( .A(_GFM_n1011 ), .B(_GFM_n10100 ), .Z(z_out[55]) );
XOR2_X2 _GFM_U3447  ( .A(_GFM_n10130 ), .B(_GFM_n10120 ), .Z(_GFM_n10100 ));
XOR2_X2 _GFM_U3446  ( .A(_GFM_n1015 ), .B(_GFM_n1014 ), .Z(_GFM_n1011 ) );
XOR2_X2 _GFM_U3445  ( .A(_GFM_n10170 ), .B(_GFM_n10160 ), .Z(_GFM_n10120 ));
XOR2_X2 _GFM_U3444  ( .A(_GFM_n10190 ), .B(_GFM_n1018 ), .Z(_GFM_n10130 ) );
XOR2_X2 _GFM_U3443  ( .A(_GFM_n1021 ), .B(_GFM_n10200 ), .Z(_GFM_n1014 ) );
XOR2_X2 _GFM_U3442  ( .A(_GFM_n1023 ), .B(_GFM_n1022 ), .Z(_GFM_n1015 ) );
XOR2_X2 _GFM_U3441  ( .A(z_in[55]), .B(_GFM_n10240 ), .Z(_GFM_n10160 ) );
XOR2_X2 _GFM_U3440  ( .A(_GFM_N1732 ), .B(_GFM_N1733 ), .Z(_GFM_n10170 ) );
XOR2_X2 _GFM_U3439  ( .A(_GFM_N1729 ), .B(_GFM_N1730 ), .Z(_GFM_n1018 ) );
XOR2_X2 _GFM_U3438  ( .A(_GFM_N1725 ), .B(_GFM_N1726 ), .Z(_GFM_n10190 ) );
XOR2_X2 _GFM_U3437  ( .A(_GFM_N1721 ), .B(_GFM_N1723 ), .Z(_GFM_n10200 ) );
XOR2_X2 _GFM_U3436  ( .A(_GFM_N1716 ), .B(_GFM_N1720 ), .Z(_GFM_n1021 ) );
XOR2_X2 _GFM_U3435  ( .A(_GFM_N1713 ), .B(_GFM_N1715 ), .Z(_GFM_n1022 ) );
XOR2_X2 _GFM_U3434  ( .A(_GFM_N1709 ), .B(_GFM_N1712 ), .Z(_GFM_n1023 ) );
XOR2_X2 _GFM_U3433  ( .A(_GFM_N1706 ), .B(_GFM_N1708 ), .Z(_GFM_n10240 ) );
XOR2_X2 _GFM_U3432  ( .A(_GFM_n10260 ), .B(_GFM_n1025 ), .Z(z_out[56]) );
XOR2_X2 _GFM_U3431  ( .A(_GFM_n1028 ), .B(_GFM_n10270 ), .Z(_GFM_n1025 ) );
XOR2_X2 _GFM_U3430  ( .A(_GFM_n10300 ), .B(_GFM_n1029 ), .Z(_GFM_n10260 ) );
XOR2_X2 _GFM_U3429  ( .A(_GFM_n1032 ), .B(_GFM_n10310 ), .Z(_GFM_n10270 ) );
XOR2_X2 _GFM_U3428  ( .A(_GFM_n10340 ), .B(_GFM_n10330 ), .Z(_GFM_n1028 ) );
XOR2_X2 _GFM_U3427  ( .A(_GFM_n1036 ), .B(_GFM_n1035 ), .Z(_GFM_n1029 ) );
XOR2_X2 _GFM_U3426  ( .A(_GFM_n10380 ), .B(_GFM_n1037 ), .Z(_GFM_n10300 ) );
XOR2_X2 _GFM_U3425  ( .A(z_in[56]), .B(_GFM_n10390 ), .Z(_GFM_n10310 ) );
XOR2_X2 _GFM_U3424  ( .A(_GFM_N1763 ), .B(_GFM_N1764 ), .Z(_GFM_n1032 ) );
XOR2_X2 _GFM_U3423  ( .A(_GFM_N1760 ), .B(_GFM_N1761 ), .Z(_GFM_n10330 ) );
XOR2_X2 _GFM_U3422  ( .A(_GFM_N1756 ), .B(_GFM_N1757 ), .Z(_GFM_n10340 ) );
XOR2_X2 _GFM_U3421  ( .A(_GFM_N1752 ), .B(_GFM_N1754 ), .Z(_GFM_n1035 ) );
XOR2_X2 _GFM_U3420  ( .A(_GFM_N1747 ), .B(_GFM_N1751 ), .Z(_GFM_n1036 ) );
XOR2_X2 _GFM_U3419  ( .A(_GFM_N1744 ), .B(_GFM_N1746 ), .Z(_GFM_n1037 ) );
XOR2_X2 _GFM_U3418  ( .A(_GFM_N1740 ), .B(_GFM_N1743 ), .Z(_GFM_n10380 ) );
XOR2_X2 _GFM_U3417  ( .A(_GFM_N1737 ), .B(_GFM_N1739 ), .Z(_GFM_n10390 ) );
XOR2_X2 _GFM_U3416  ( .A(_GFM_n10410 ), .B(_GFM_n1040 ), .Z(z_out[57]) );
XOR2_X2 _GFM_U3415  ( .A(_GFM_n10430 ), .B(_GFM_n1042 ), .Z(_GFM_n1040 ) );
XOR2_X2 _GFM_U3414  ( .A(_GFM_n1045 ), .B(_GFM_n10440 ), .Z(_GFM_n10410 ) );
XOR2_X2 _GFM_U3413  ( .A(_GFM_n10470 ), .B(_GFM_n1046 ), .Z(_GFM_n1042 ) );
XOR2_X2 _GFM_U3412  ( .A(_GFM_n1049 ), .B(_GFM_n10480 ), .Z(_GFM_n10430 ) );
XOR2_X2 _GFM_U3411  ( .A(_GFM_n10510 ), .B(_GFM_n10500 ), .Z(_GFM_n10440 ));
XOR2_X2 _GFM_U3410  ( .A(_GFM_n1053 ), .B(_GFM_n1052 ), .Z(_GFM_n1045 ) );
XOR2_X2 _GFM_U3409  ( .A(z_in[57]), .B(_GFM_n1054 ), .Z(_GFM_n1046 ) );
XOR2_X2 _GFM_U3408  ( .A(_GFM_N1794 ), .B(_GFM_N1795 ), .Z(_GFM_n10470 ) );
XOR2_X2 _GFM_U3407  ( .A(_GFM_N1791 ), .B(_GFM_N1792 ), .Z(_GFM_n10480 ) );
XOR2_X2 _GFM_U3406  ( .A(_GFM_N1787 ), .B(_GFM_N1788 ), .Z(_GFM_n1049 ) );
XOR2_X2 _GFM_U3405  ( .A(_GFM_N1783 ), .B(_GFM_N1785 ), .Z(_GFM_n10500 ) );
XOR2_X2 _GFM_U3404  ( .A(_GFM_N1778 ), .B(_GFM_N1782 ), .Z(_GFM_n10510 ) );
XOR2_X2 _GFM_U3403  ( .A(_GFM_N1775 ), .B(_GFM_N1777 ), .Z(_GFM_n1052 ) );
XOR2_X2 _GFM_U3402  ( .A(_GFM_N1771 ), .B(_GFM_N1774 ), .Z(_GFM_n1053 ) );
XOR2_X2 _GFM_U3401  ( .A(_GFM_N1768 ), .B(_GFM_N1770 ), .Z(_GFM_n1054 ) );
XOR2_X2 _GFM_U3400  ( .A(_GFM_n1056 ), .B(_GFM_n10550 ), .Z(z_out[58]) );
XOR2_X2 _GFM_U3399  ( .A(_GFM_n10580 ), .B(_GFM_n10570 ), .Z(_GFM_n10550 ));
XOR2_X2 _GFM_U3398  ( .A(_GFM_n1060 ), .B(_GFM_n1059 ), .Z(_GFM_n1056 ) );
XOR2_X2 _GFM_U3397  ( .A(_GFM_n10620 ), .B(_GFM_n10610 ), .Z(_GFM_n10570 ));
XOR2_X2 _GFM_U3396  ( .A(_GFM_n10640 ), .B(_GFM_n1063 ), .Z(_GFM_n10580 ) );
XOR2_X2 _GFM_U3395  ( .A(_GFM_n1066 ), .B(_GFM_n10650 ), .Z(_GFM_n1059 ) );
XOR2_X2 _GFM_U3394  ( .A(_GFM_n1068 ), .B(_GFM_n1067 ), .Z(_GFM_n1060 ) );
XOR2_X2 _GFM_U3393  ( .A(z_in[58]), .B(_GFM_n10690 ), .Z(_GFM_n10610 ) );
XOR2_X2 _GFM_U3392  ( .A(_GFM_N1825 ), .B(_GFM_N1826 ), .Z(_GFM_n10620 ) );
XOR2_X2 _GFM_U3391  ( .A(_GFM_N1822 ), .B(_GFM_N1823 ), .Z(_GFM_n1063 ) );
XOR2_X2 _GFM_U3390  ( .A(_GFM_N1818 ), .B(_GFM_N1819 ), .Z(_GFM_n10640 ) );
XOR2_X2 _GFM_U3389  ( .A(_GFM_N1814 ), .B(_GFM_N1816 ), .Z(_GFM_n10650 ) );
XOR2_X2 _GFM_U3388  ( .A(_GFM_N1809 ), .B(_GFM_N1813 ), .Z(_GFM_n1066 ) );
XOR2_X2 _GFM_U3387  ( .A(_GFM_N1806 ), .B(_GFM_N1808 ), .Z(_GFM_n1067 ) );
XOR2_X2 _GFM_U3386  ( .A(_GFM_N1802 ), .B(_GFM_N1805 ), .Z(_GFM_n1068 ) );
XOR2_X2 _GFM_U3385  ( .A(_GFM_N1799 ), .B(_GFM_N1801 ), .Z(_GFM_n10690 ) );
XOR2_X2 _GFM_U3384  ( .A(_GFM_n1071 ), .B(_GFM_n10700 ), .Z(z_out[59]) );
XOR2_X2 _GFM_U3383  ( .A(_GFM_n1073 ), .B(_GFM_n10720 ), .Z(_GFM_n10700 ) );
XOR2_X2 _GFM_U3382  ( .A(_GFM_n10750 ), .B(_GFM_n10740 ), .Z(_GFM_n1071 ) );
XOR2_X2 _GFM_U3381  ( .A(_GFM_n1077 ), .B(_GFM_n1076 ), .Z(_GFM_n10720 ) );
XOR2_X2 _GFM_U3380  ( .A(_GFM_n10790 ), .B(_GFM_n10780 ), .Z(_GFM_n1073 ) );
XOR2_X2 _GFM_U3379  ( .A(_GFM_n10810 ), .B(_GFM_n1080 ), .Z(_GFM_n10740 ) );
XOR2_X2 _GFM_U3378  ( .A(_GFM_n1083 ), .B(_GFM_n10820 ), .Z(_GFM_n10750 ) );
XOR2_X2 _GFM_U3377  ( .A(z_in[59]), .B(_GFM_n1084 ), .Z(_GFM_n1076 ) );
XOR2_X2 _GFM_U3376  ( .A(_GFM_N1856 ), .B(_GFM_N1857 ), .Z(_GFM_n1077 ) );
XOR2_X2 _GFM_U3375  ( .A(_GFM_N1853 ), .B(_GFM_N1854 ), .Z(_GFM_n10780 ) );
XOR2_X2 _GFM_U3374  ( .A(_GFM_N1849 ), .B(_GFM_N1850 ), .Z(_GFM_n10790 ) );
XOR2_X2 _GFM_U3373  ( .A(_GFM_N1845 ), .B(_GFM_N1847 ), .Z(_GFM_n1080 ) );
XOR2_X2 _GFM_U3372  ( .A(_GFM_N1840 ), .B(_GFM_N1844 ), .Z(_GFM_n10810 ) );
XOR2_X2 _GFM_U3371  ( .A(_GFM_N1837 ), .B(_GFM_N1839 ), .Z(_GFM_n10820 ) );
XOR2_X2 _GFM_U3370  ( .A(_GFM_N1833 ), .B(_GFM_N1836 ), .Z(_GFM_n1083 ) );
XOR2_X2 _GFM_U3369  ( .A(_GFM_N1830 ), .B(_GFM_N1832 ), .Z(_GFM_n1084 ) );
XOR2_X2 _GFM_U3368  ( .A(_GFM_n10860 ), .B(_GFM_n1085 ), .Z(z_out[60]) );
XOR2_X2 _GFM_U3367  ( .A(_GFM_n10880 ), .B(_GFM_n1087 ), .Z(_GFM_n1085 ) );
XOR2_X2 _GFM_U3366  ( .A(_GFM_n1090 ), .B(_GFM_n10890 ), .Z(_GFM_n10860 ) );
XOR2_X2 _GFM_U3365  ( .A(_GFM_n10920 ), .B(_GFM_n1091 ), .Z(_GFM_n1087 ) );
XOR2_X2 _GFM_U3364  ( .A(_GFM_n1094 ), .B(_GFM_n10930 ), .Z(_GFM_n10880 ) );
XOR2_X2 _GFM_U3363  ( .A(_GFM_n10960 ), .B(_GFM_n10950 ), .Z(_GFM_n10890 ));
XOR2_X2 _GFM_U3362  ( .A(_GFM_n1098 ), .B(_GFM_n1097 ), .Z(_GFM_n1090 ) );
XOR2_X2 _GFM_U3361  ( .A(z_in[60]), .B(_GFM_n1099 ), .Z(_GFM_n1091 ) );
XOR2_X2 _GFM_U3360  ( .A(_GFM_N1887 ), .B(_GFM_N1888 ), .Z(_GFM_n10920 ) );
XOR2_X2 _GFM_U3359  ( .A(_GFM_N1884 ), .B(_GFM_N1885 ), .Z(_GFM_n10930 ) );
XOR2_X2 _GFM_U3358  ( .A(_GFM_N1880 ), .B(_GFM_N1881 ), .Z(_GFM_n1094 ) );
XOR2_X2 _GFM_U3357  ( .A(_GFM_N1876 ), .B(_GFM_N1878 ), .Z(_GFM_n10950 ) );
XOR2_X2 _GFM_U3356  ( .A(_GFM_N1871 ), .B(_GFM_N1875 ), .Z(_GFM_n10960 ) );
XOR2_X2 _GFM_U3355  ( .A(_GFM_N1868 ), .B(_GFM_N1870 ), .Z(_GFM_n1097 ) );
XOR2_X2 _GFM_U3354  ( .A(_GFM_N1864 ), .B(_GFM_N1867 ), .Z(_GFM_n1098 ) );
XOR2_X2 _GFM_U3353  ( .A(_GFM_N1861 ), .B(_GFM_N1863 ), .Z(_GFM_n1099 ) );
XOR2_X2 _GFM_U3352  ( .A(_GFM_n11010 ), .B(_GFM_n11000 ), .Z(z_out[61]) );
XOR2_X2 _GFM_U3351  ( .A(_GFM_n11030 ), .B(_GFM_n1102 ), .Z(_GFM_n11000 ) );
XOR2_X2 _GFM_U3350  ( .A(_GFM_n11050 ), .B(_GFM_n1104 ), .Z(_GFM_n11010 ) );
XOR2_X2 _GFM_U3349  ( .A(_GFM_n1107 ), .B(_GFM_n11060 ), .Z(_GFM_n1102 ) );
XOR2_X2 _GFM_U3348  ( .A(_GFM_n11090 ), .B(_GFM_n1108 ), .Z(_GFM_n11030 ) );
XOR2_X2 _GFM_U3347  ( .A(_GFM_n1111 ), .B(_GFM_n11100 ), .Z(_GFM_n1104 ) );
XOR2_X2 _GFM_U3346  ( .A(_GFM_n11130 ), .B(_GFM_n11120 ), .Z(_GFM_n11050 ));
XOR2_X2 _GFM_U3345  ( .A(z_in[61]), .B(_GFM_n1114 ), .Z(_GFM_n11060 ) );
XOR2_X2 _GFM_U3344  ( .A(_GFM_N1918 ), .B(_GFM_N1919 ), .Z(_GFM_n1107 ) );
XOR2_X2 _GFM_U3343  ( .A(_GFM_N1915 ), .B(_GFM_N1916 ), .Z(_GFM_n1108 ) );
XOR2_X2 _GFM_U3342  ( .A(_GFM_N1911 ), .B(_GFM_N1912 ), .Z(_GFM_n11090 ) );
XOR2_X2 _GFM_U3341  ( .A(_GFM_N1907 ), .B(_GFM_N1909 ), .Z(_GFM_n11100 ) );
XOR2_X2 _GFM_U3340  ( .A(_GFM_N1902 ), .B(_GFM_N1906 ), .Z(_GFM_n1111 ) );
XOR2_X2 _GFM_U3339  ( .A(_GFM_N1899 ), .B(_GFM_N1901 ), .Z(_GFM_n11120 ) );
XOR2_X2 _GFM_U3338  ( .A(_GFM_N1895 ), .B(_GFM_N1898 ), .Z(_GFM_n11130 ) );
XOR2_X2 _GFM_U3337  ( .A(_GFM_N1892 ), .B(_GFM_N1894 ), .Z(_GFM_n1114 ) );
XOR2_X2 _GFM_U3336  ( .A(_GFM_n1116 ), .B(_GFM_n1115 ), .Z(z_out[62]) );
XOR2_X2 _GFM_U3335  ( .A(_GFM_n1118 ), .B(_GFM_n11170 ), .Z(_GFM_n1115 ) );
XOR2_X2 _GFM_U3334  ( .A(_GFM_n11200 ), .B(_GFM_n11190 ), .Z(_GFM_n1116 ) );
XOR2_X2 _GFM_U3333  ( .A(_GFM_n1122 ), .B(_GFM_n1121 ), .Z(_GFM_n11170 ) );
XOR2_X2 _GFM_U3332  ( .A(_GFM_n11240 ), .B(_GFM_n11230 ), .Z(_GFM_n1118 ) );
XOR2_X2 _GFM_U3331  ( .A(_GFM_n11260 ), .B(_GFM_n1125 ), .Z(_GFM_n11190 ) );
XOR2_X2 _GFM_U3330  ( .A(_GFM_n1128 ), .B(_GFM_n11270 ), .Z(_GFM_n11200 ) );
XOR2_X2 _GFM_U3329  ( .A(z_in[62]), .B(_GFM_n1129 ), .Z(_GFM_n1121 ) );
XOR2_X2 _GFM_U3328  ( .A(_GFM_N1949 ), .B(_GFM_N1950 ), .Z(_GFM_n1122 ) );
XOR2_X2 _GFM_U3327  ( .A(_GFM_N1946 ), .B(_GFM_N1947 ), .Z(_GFM_n11230 ) );
XOR2_X2 _GFM_U3326  ( .A(_GFM_N1942 ), .B(_GFM_N1943 ), .Z(_GFM_n11240 ) );
XOR2_X2 _GFM_U3325  ( .A(_GFM_N1938 ), .B(_GFM_N1940 ), .Z(_GFM_n1125 ) );
XOR2_X2 _GFM_U3324  ( .A(_GFM_N1933 ), .B(_GFM_N1937 ), .Z(_GFM_n11260 ) );
XOR2_X2 _GFM_U3323  ( .A(_GFM_N1930 ), .B(_GFM_N1932 ), .Z(_GFM_n11270 ) );
XOR2_X2 _GFM_U3322  ( .A(_GFM_N1926 ), .B(_GFM_N1929 ), .Z(_GFM_n1128 ) );
XOR2_X2 _GFM_U3321  ( .A(_GFM_N1923 ), .B(_GFM_N1925 ), .Z(_GFM_n1129 ) );
XOR2_X2 _GFM_U3320  ( .A(_GFM_n11310 ), .B(_GFM_n1130 ), .Z(z_out[63]) );
XOR2_X2 _GFM_U3319  ( .A(_GFM_n1133 ), .B(_GFM_n11320 ), .Z(_GFM_n1130 ) );
XOR2_X2 _GFM_U3318  ( .A(_GFM_n1135 ), .B(_GFM_n11340 ), .Z(_GFM_n11310 ) );
XOR2_X2 _GFM_U3317  ( .A(_GFM_n11370 ), .B(_GFM_n11360 ), .Z(_GFM_n11320 ));
XOR2_X2 _GFM_U3316  ( .A(_GFM_n1139 ), .B(_GFM_n1138 ), .Z(_GFM_n1133 ) );
XOR2_X2 _GFM_U3315  ( .A(_GFM_n11410 ), .B(_GFM_n11400 ), .Z(_GFM_n11340 ));
XOR2_X2 _GFM_U3314  ( .A(_GFM_n11430 ), .B(_GFM_n1142 ), .Z(_GFM_n1135 ) );
XOR2_X2 _GFM_U3313  ( .A(z_in[63]), .B(_GFM_n11440 ), .Z(_GFM_n11360 ) );
XOR2_X2 _GFM_U3312  ( .A(_GFM_N1980 ), .B(_GFM_N1981 ), .Z(_GFM_n11370 ) );
XOR2_X2 _GFM_U3311  ( .A(_GFM_N1977 ), .B(_GFM_N1978 ), .Z(_GFM_n1138 ) );
XOR2_X2 _GFM_U3310  ( .A(_GFM_N1973 ), .B(_GFM_N1974 ), .Z(_GFM_n1139 ) );
XOR2_X2 _GFM_U3309  ( .A(_GFM_N1969 ), .B(_GFM_N1971 ), .Z(_GFM_n11400 ) );
XOR2_X2 _GFM_U3308  ( .A(_GFM_N1964 ), .B(_GFM_N1968 ), .Z(_GFM_n11410 ) );
XOR2_X2 _GFM_U3307  ( .A(_GFM_N1961 ), .B(_GFM_N1963 ), .Z(_GFM_n1142 ) );
XOR2_X2 _GFM_U3306  ( .A(_GFM_N1957 ), .B(_GFM_N1960 ), .Z(_GFM_n11430 ) );
XOR2_X2 _GFM_U3305  ( .A(_GFM_N1954 ), .B(_GFM_N1956 ), .Z(_GFM_n11440 ) );
XOR2_X2 _GFM_U3304  ( .A(_GFM_n1146 ), .B(_GFM_n1145 ), .Z(z_out[64]) );
XOR2_X2 _GFM_U3303  ( .A(_GFM_n11480 ), .B(_GFM_n1147 ), .Z(_GFM_n1145 ) );
XOR2_X2 _GFM_U3302  ( .A(_GFM_n11500 ), .B(_GFM_n1149 ), .Z(_GFM_n1146 ) );
XOR2_X2 _GFM_U3301  ( .A(_GFM_n1152 ), .B(_GFM_n11510 ), .Z(_GFM_n1147 ) );
XOR2_X2 _GFM_U3300  ( .A(_GFM_n11540 ), .B(_GFM_n1153 ), .Z(_GFM_n11480 ) );
XOR2_X2 _GFM_U3299  ( .A(_GFM_n1156 ), .B(_GFM_n11550 ), .Z(_GFM_n1149 ) );
XOR2_X2 _GFM_U3298  ( .A(_GFM_n11580 ), .B(_GFM_n11570 ), .Z(_GFM_n11500 ));
XOR2_X2 _GFM_U3297  ( .A(z_in[64]), .B(_GFM_n1159 ), .Z(_GFM_n11510 ) );
XOR2_X2 _GFM_U3296  ( .A(_GFM_N2011 ), .B(_GFM_N2012 ), .Z(_GFM_n1152 ) );
XOR2_X2 _GFM_U3295  ( .A(_GFM_N2008 ), .B(_GFM_N2009 ), .Z(_GFM_n1153 ) );
XOR2_X2 _GFM_U3294  ( .A(_GFM_N2004 ), .B(_GFM_N2005 ), .Z(_GFM_n11540 ) );
XOR2_X2 _GFM_U3293  ( .A(_GFM_N2000 ), .B(_GFM_N2002 ), .Z(_GFM_n11550 ) );
XOR2_X2 _GFM_U3292  ( .A(_GFM_N1995 ), .B(_GFM_N1999 ), .Z(_GFM_n1156 ) );
XOR2_X2 _GFM_U3291  ( .A(_GFM_N1992 ), .B(_GFM_N1994 ), .Z(_GFM_n11570 ) );
XOR2_X2 _GFM_U3290  ( .A(_GFM_N1988 ), .B(_GFM_N1991 ), .Z(_GFM_n11580 ) );
XOR2_X2 _GFM_U3289  ( .A(_GFM_N1985 ), .B(_GFM_N1987 ), .Z(_GFM_n1159 ) );
XOR2_X2 _GFM_U3288  ( .A(_GFM_n1161 ), .B(_GFM_n1160 ), .Z(z_out[65]) );
XOR2_X2 _GFM_U3287  ( .A(_GFM_n11630 ), .B(_GFM_n11620 ), .Z(_GFM_n1160 ) );
XOR2_X2 _GFM_U3286  ( .A(_GFM_n11650 ), .B(_GFM_n1164 ), .Z(_GFM_n1161 ) );
XOR2_X2 _GFM_U3285  ( .A(_GFM_n11670 ), .B(_GFM_n1166 ), .Z(_GFM_n11620 ) );
XOR2_X2 _GFM_U3284  ( .A(_GFM_n1169 ), .B(_GFM_n11680 ), .Z(_GFM_n11630 ) );
XOR2_X2 _GFM_U3283  ( .A(_GFM_n11710 ), .B(_GFM_n1170 ), .Z(_GFM_n1164 ) );
XOR2_X2 _GFM_U3282  ( .A(_GFM_n1173 ), .B(_GFM_n11720 ), .Z(_GFM_n11650 ) );
XOR2_X2 _GFM_U3281  ( .A(z_in[65]), .B(_GFM_n11740 ), .Z(_GFM_n1166 ) );
XOR2_X2 _GFM_U3280  ( .A(_GFM_N2042 ), .B(_GFM_N2043 ), .Z(_GFM_n11670 ) );
XOR2_X2 _GFM_U3279  ( .A(_GFM_N2039 ), .B(_GFM_N2040 ), .Z(_GFM_n11680 ) );
XOR2_X2 _GFM_U3278  ( .A(_GFM_N2035 ), .B(_GFM_N2036 ), .Z(_GFM_n1169 ) );
XOR2_X2 _GFM_U3277  ( .A(_GFM_N2031 ), .B(_GFM_N2033 ), .Z(_GFM_n1170 ) );
XOR2_X2 _GFM_U3276  ( .A(_GFM_N2026 ), .B(_GFM_N2030 ), .Z(_GFM_n11710 ) );
XOR2_X2 _GFM_U3275  ( .A(_GFM_N2023 ), .B(_GFM_N2025 ), .Z(_GFM_n11720 ) );
XOR2_X2 _GFM_U3274  ( .A(_GFM_N2019 ), .B(_GFM_N2022 ), .Z(_GFM_n1173 ) );
XOR2_X2 _GFM_U3273  ( .A(_GFM_N2016 ), .B(_GFM_N2018 ), .Z(_GFM_n11740 ) );
XOR2_X2 _GFM_U3272  ( .A(_GFM_n1176 ), .B(_GFM_n11750 ), .Z(z_out[66]) );
XOR2_X2 _GFM_U3271  ( .A(_GFM_n1178 ), .B(_GFM_n1177 ), .Z(_GFM_n11750 ) );
XOR2_X2 _GFM_U3270  ( .A(_GFM_n1180 ), .B(_GFM_n11790 ), .Z(_GFM_n1176 ) );
XOR2_X2 _GFM_U3269  ( .A(_GFM_n11820 ), .B(_GFM_n11810 ), .Z(_GFM_n1177 ) );
XOR2_X2 _GFM_U3268  ( .A(_GFM_n1184 ), .B(_GFM_n1183 ), .Z(_GFM_n1178 ) );
XOR2_X2 _GFM_U3267  ( .A(_GFM_n11860 ), .B(_GFM_n11850 ), .Z(_GFM_n11790 ));
XOR2_X2 _GFM_U3266  ( .A(_GFM_n11880 ), .B(_GFM_n1187 ), .Z(_GFM_n1180 ) );
XOR2_X2 _GFM_U3265  ( .A(z_in[66]), .B(_GFM_n11890 ), .Z(_GFM_n11810 ) );
XOR2_X2 _GFM_U3264  ( .A(_GFM_N2073 ), .B(_GFM_N2074 ), .Z(_GFM_n11820 ) );
XOR2_X2 _GFM_U3263  ( .A(_GFM_N2070 ), .B(_GFM_N2071 ), .Z(_GFM_n1183 ) );
XOR2_X2 _GFM_U3262  ( .A(_GFM_N2066 ), .B(_GFM_N2067 ), .Z(_GFM_n1184 ) );
XOR2_X2 _GFM_U3261  ( .A(_GFM_N2062 ), .B(_GFM_N2064 ), .Z(_GFM_n11850 ) );
XOR2_X2 _GFM_U3260  ( .A(_GFM_N2057 ), .B(_GFM_N2061 ), .Z(_GFM_n11860 ) );
XOR2_X2 _GFM_U3259  ( .A(_GFM_N2054 ), .B(_GFM_N2056 ), .Z(_GFM_n1187 ) );
XOR2_X2 _GFM_U3258  ( .A(_GFM_N2050 ), .B(_GFM_N2053 ), .Z(_GFM_n11880 ) );
XOR2_X2 _GFM_U3257  ( .A(_GFM_N2047 ), .B(_GFM_N2049 ), .Z(_GFM_n11890 ) );
XOR2_X2 _GFM_U3256  ( .A(_GFM_n1191 ), .B(_GFM_n1190 ), .Z(z_out[67]) );
XOR2_X2 _GFM_U3255  ( .A(_GFM_n11930 ), .B(_GFM_n1192 ), .Z(_GFM_n1190 ) );
XOR2_X2 _GFM_U3254  ( .A(_GFM_n1195 ), .B(_GFM_n11940 ), .Z(_GFM_n1191 ) );
XOR2_X2 _GFM_U3253  ( .A(_GFM_n1197 ), .B(_GFM_n11960 ), .Z(_GFM_n1192 ) );
XOR2_X2 _GFM_U3252  ( .A(_GFM_n11990 ), .B(_GFM_n11980 ), .Z(_GFM_n11930 ));
XOR2_X2 _GFM_U3251  ( .A(_GFM_n1201 ), .B(_GFM_n1200 ), .Z(_GFM_n11940 ) );
XOR2_X2 _GFM_U3250  ( .A(_GFM_n12030 ), .B(_GFM_n12020 ), .Z(_GFM_n1195 ) );
XOR2_X2 _GFM_U3249  ( .A(z_in[67]), .B(_GFM_n1204 ), .Z(_GFM_n11960 ) );
XOR2_X2 _GFM_U3248  ( .A(_GFM_N2104 ), .B(_GFM_N2105 ), .Z(_GFM_n1197 ) );
XOR2_X2 _GFM_U3247  ( .A(_GFM_N2101 ), .B(_GFM_N2102 ), .Z(_GFM_n11980 ) );
XOR2_X2 _GFM_U3246  ( .A(_GFM_N2097 ), .B(_GFM_N2098 ), .Z(_GFM_n11990 ) );
XOR2_X2 _GFM_U3245  ( .A(_GFM_N2093 ), .B(_GFM_N2095 ), .Z(_GFM_n1200 ) );
XOR2_X2 _GFM_U3244  ( .A(_GFM_N2088 ), .B(_GFM_N2092 ), .Z(_GFM_n1201 ) );
XOR2_X2 _GFM_U3243  ( .A(_GFM_N2085 ), .B(_GFM_N2087 ), .Z(_GFM_n12020 ) );
XOR2_X2 _GFM_U3242  ( .A(_GFM_N2081 ), .B(_GFM_N2084 ), .Z(_GFM_n12030 ) );
XOR2_X2 _GFM_U3241  ( .A(_GFM_N2078 ), .B(_GFM_N2080 ), .Z(_GFM_n1204 ) );
XOR2_X2 _GFM_U3240  ( .A(_GFM_n12060 ), .B(_GFM_n12050 ), .Z(z_out[68]) );
XOR2_X2 _GFM_U3239  ( .A(_GFM_n1208 ), .B(_GFM_n1207 ), .Z(_GFM_n12050 ) );
XOR2_X2 _GFM_U3238  ( .A(_GFM_n12100 ), .B(_GFM_n1209 ), .Z(_GFM_n12060 ) );
XOR2_X2 _GFM_U3237  ( .A(_GFM_n12120 ), .B(_GFM_n1211 ), .Z(_GFM_n1207 ) );
XOR2_X2 _GFM_U3236  ( .A(_GFM_n1214 ), .B(_GFM_n12130 ), .Z(_GFM_n1208 ) );
XOR2_X2 _GFM_U3235  ( .A(_GFM_n12160 ), .B(_GFM_n1215 ), .Z(_GFM_n1209 ) );
XOR2_X2 _GFM_U3234  ( .A(_GFM_n1218 ), .B(_GFM_n12170 ), .Z(_GFM_n12100 ) );
XOR2_X2 _GFM_U3233  ( .A(z_in[68]), .B(_GFM_n12190 ), .Z(_GFM_n1211 ) );
XOR2_X2 _GFM_U3232  ( .A(_GFM_N2135 ), .B(_GFM_N2136 ), .Z(_GFM_n12120 ) );
XOR2_X2 _GFM_U3231  ( .A(_GFM_N2132 ), .B(_GFM_N2133 ), .Z(_GFM_n12130 ) );
XOR2_X2 _GFM_U3230  ( .A(_GFM_N2128 ), .B(_GFM_N2129 ), .Z(_GFM_n1214 ) );
XOR2_X2 _GFM_U3229  ( .A(_GFM_N2124 ), .B(_GFM_N2126 ), .Z(_GFM_n1215 ) );
XOR2_X2 _GFM_U3228  ( .A(_GFM_N2119 ), .B(_GFM_N2123 ), .Z(_GFM_n12160 ) );
XOR2_X2 _GFM_U3227  ( .A(_GFM_N2116 ), .B(_GFM_N2118 ), .Z(_GFM_n12170 ) );
XOR2_X2 _GFM_U3226  ( .A(_GFM_N2112 ), .B(_GFM_N2115 ), .Z(_GFM_n1218 ) );
XOR2_X2 _GFM_U3225  ( .A(_GFM_N2109 ), .B(_GFM_N2111 ), .Z(_GFM_n12190 ) );
XOR2_X2 _GFM_U3224  ( .A(_GFM_n1221 ), .B(_GFM_n12200 ), .Z(z_out[69]) );
XOR2_X2 _GFM_U3223  ( .A(_GFM_n1223 ), .B(_GFM_n1222 ), .Z(_GFM_n12200 ) );
XOR2_X2 _GFM_U3222  ( .A(_GFM_n12250 ), .B(_GFM_n12240 ), .Z(_GFM_n1221 ) );
XOR2_X2 _GFM_U3221  ( .A(_GFM_n12270 ), .B(_GFM_n1226 ), .Z(_GFM_n1222 ) );
XOR2_X2 _GFM_U3220  ( .A(_GFM_n12290 ), .B(_GFM_n1228 ), .Z(_GFM_n1223 ) );
XOR2_X2 _GFM_U3219  ( .A(_GFM_n1231 ), .B(_GFM_n12300 ), .Z(_GFM_n12240 ) );
XOR2_X2 _GFM_U3218  ( .A(_GFM_n12330 ), .B(_GFM_n1232 ), .Z(_GFM_n12250 ) );
XOR2_X2 _GFM_U3217  ( .A(z_in[69]), .B(_GFM_n12340 ), .Z(_GFM_n1226 ) );
XOR2_X2 _GFM_U3216  ( .A(_GFM_N2166 ), .B(_GFM_N2167 ), .Z(_GFM_n12270 ) );
XOR2_X2 _GFM_U3215  ( .A(_GFM_N2163 ), .B(_GFM_N2164 ), .Z(_GFM_n1228 ) );
XOR2_X2 _GFM_U3214  ( .A(_GFM_N2159 ), .B(_GFM_N2160 ), .Z(_GFM_n12290 ) );
XOR2_X2 _GFM_U3213  ( .A(_GFM_N2155 ), .B(_GFM_N2157 ), .Z(_GFM_n12300 ) );
XOR2_X2 _GFM_U3212  ( .A(_GFM_N2150 ), .B(_GFM_N2154 ), .Z(_GFM_n1231 ) );
XOR2_X2 _GFM_U3211  ( .A(_GFM_N2147 ), .B(_GFM_N2149 ), .Z(_GFM_n1232 ) );
XOR2_X2 _GFM_U3210  ( .A(_GFM_N2143 ), .B(_GFM_N2146 ), .Z(_GFM_n12330 ) );
XOR2_X2 _GFM_U3209  ( .A(_GFM_N2140 ), .B(_GFM_N2142 ), .Z(_GFM_n12340 ) );
XOR2_X2 _GFM_U3208  ( .A(_GFM_n12360 ), .B(_GFM_n1235 ), .Z(z_out[70]) );
XOR2_X2 _GFM_U3207  ( .A(_GFM_n1238 ), .B(_GFM_n12370 ), .Z(_GFM_n1235 ) );
XOR2_X2 _GFM_U3206  ( .A(_GFM_n1240 ), .B(_GFM_n1239 ), .Z(_GFM_n12360 ) );
XOR2_X2 _GFM_U3205  ( .A(_GFM_n1242 ), .B(_GFM_n12410 ), .Z(_GFM_n12370 ) );
XOR2_X2 _GFM_U3204  ( .A(_GFM_n12440 ), .B(_GFM_n12430 ), .Z(_GFM_n1238 ) );
XOR2_X2 _GFM_U3203  ( .A(_GFM_n1246 ), .B(_GFM_n1245 ), .Z(_GFM_n1239 ) );
XOR2_X2 _GFM_U3202  ( .A(_GFM_n12480 ), .B(_GFM_n12470 ), .Z(_GFM_n1240 ) );
XOR2_X2 _GFM_U3201  ( .A(z_in[70]), .B(_GFM_n1249 ), .Z(_GFM_n12410 ) );
XOR2_X2 _GFM_U3200  ( .A(_GFM_N2197 ), .B(_GFM_N2198 ), .Z(_GFM_n1242 ) );
XOR2_X2 _GFM_U3199  ( .A(_GFM_N2194 ), .B(_GFM_N2195 ), .Z(_GFM_n12430 ) );
XOR2_X2 _GFM_U3198  ( .A(_GFM_N2190 ), .B(_GFM_N2191 ), .Z(_GFM_n12440 ) );
XOR2_X2 _GFM_U3197  ( .A(_GFM_N2186 ), .B(_GFM_N2188 ), .Z(_GFM_n1245 ) );
XOR2_X2 _GFM_U3196  ( .A(_GFM_N2181 ), .B(_GFM_N2185 ), .Z(_GFM_n1246 ) );
XOR2_X2 _GFM_U3195  ( .A(_GFM_N2178 ), .B(_GFM_N2180 ), .Z(_GFM_n12470 ) );
XOR2_X2 _GFM_U3194  ( .A(_GFM_N2174 ), .B(_GFM_N2177 ), .Z(_GFM_n12480 ) );
XOR2_X2 _GFM_U3193  ( .A(_GFM_N2171 ), .B(_GFM_N2173 ), .Z(_GFM_n1249 ) );
XOR2_X2 _GFM_U3192  ( .A(_GFM_n12510 ), .B(_GFM_n12500 ), .Z(z_out[71]) );
XOR2_X2 _GFM_U3191  ( .A(_GFM_n1253 ), .B(_GFM_n1252 ), .Z(_GFM_n12500 ) );
XOR2_X2 _GFM_U3190  ( .A(_GFM_n12550 ), .B(_GFM_n1254 ), .Z(_GFM_n12510 ) );
XOR2_X2 _GFM_U3189  ( .A(_GFM_n1257 ), .B(_GFM_n12560 ), .Z(_GFM_n1252 ) );
XOR2_X2 _GFM_U3188  ( .A(_GFM_n1259 ), .B(_GFM_n12580 ), .Z(_GFM_n1253 ) );
XOR2_X2 _GFM_U3187  ( .A(_GFM_n12610 ), .B(_GFM_n12600 ), .Z(_GFM_n1254 ) );
XOR2_X2 _GFM_U3186  ( .A(_GFM_n1263 ), .B(_GFM_n1262 ), .Z(_GFM_n12550 ) );
XOR2_X2 _GFM_U3185  ( .A(z_in[71]), .B(_GFM_n12640 ), .Z(_GFM_n12560 ) );
XOR2_X2 _GFM_U3184  ( .A(_GFM_N2228 ), .B(_GFM_N2229 ), .Z(_GFM_n1257 ) );
XOR2_X2 _GFM_U3183  ( .A(_GFM_N2225 ), .B(_GFM_N2226 ), .Z(_GFM_n12580 ) );
XOR2_X2 _GFM_U3182  ( .A(_GFM_N2221 ), .B(_GFM_N2222 ), .Z(_GFM_n1259 ) );
XOR2_X2 _GFM_U3181  ( .A(_GFM_N2217 ), .B(_GFM_N2219 ), .Z(_GFM_n12600 ) );
XOR2_X2 _GFM_U3180  ( .A(_GFM_N2212 ), .B(_GFM_N2216 ), .Z(_GFM_n12610 ) );
XOR2_X2 _GFM_U3179  ( .A(_GFM_N2209 ), .B(_GFM_N2211 ), .Z(_GFM_n1262 ) );
XOR2_X2 _GFM_U3178  ( .A(_GFM_N2205 ), .B(_GFM_N2208 ), .Z(_GFM_n1263 ) );
XOR2_X2 _GFM_U3177  ( .A(_GFM_N2202 ), .B(_GFM_N2204 ), .Z(_GFM_n12640 ) );
XOR2_X2 _GFM_U3176  ( .A(_GFM_n1266 ), .B(_GFM_n12650 ), .Z(z_out[72]) );
XOR2_X2 _GFM_U3175  ( .A(_GFM_n12680 ), .B(_GFM_n12670 ), .Z(_GFM_n12650 ));
XOR2_X2 _GFM_U3174  ( .A(_GFM_n1270 ), .B(_GFM_n1269 ), .Z(_GFM_n1266 ) );
XOR2_X2 _GFM_U3173  ( .A(_GFM_n12720 ), .B(_GFM_n1271 ), .Z(_GFM_n12670 ) );
XOR2_X2 _GFM_U3172  ( .A(_GFM_n12740 ), .B(_GFM_n1273 ), .Z(_GFM_n12680 ) );
XOR2_X2 _GFM_U3171  ( .A(_GFM_n1276 ), .B(_GFM_n12750 ), .Z(_GFM_n1269 ) );
XOR2_X2 _GFM_U3170  ( .A(_GFM_n12780 ), .B(_GFM_n1277 ), .Z(_GFM_n1270 ) );
XOR2_X2 _GFM_U3169  ( .A(z_in[72]), .B(_GFM_n12790 ), .Z(_GFM_n1271 ) );
XOR2_X2 _GFM_U3168  ( .A(_GFM_N2259 ), .B(_GFM_N2260 ), .Z(_GFM_n12720 ) );
XOR2_X2 _GFM_U3167  ( .A(_GFM_N2256 ), .B(_GFM_N2257 ), .Z(_GFM_n1273 ) );
XOR2_X2 _GFM_U3166  ( .A(_GFM_N2252 ), .B(_GFM_N2253 ), .Z(_GFM_n12740 ) );
XOR2_X2 _GFM_U3165  ( .A(_GFM_N2248 ), .B(_GFM_N2250 ), .Z(_GFM_n12750 ) );
XOR2_X2 _GFM_U3164  ( .A(_GFM_N2243 ), .B(_GFM_N2247 ), .Z(_GFM_n1276 ) );
XOR2_X2 _GFM_U3163  ( .A(_GFM_N2240 ), .B(_GFM_N2242 ), .Z(_GFM_n1277 ) );
XOR2_X2 _GFM_U3162  ( .A(_GFM_N2236 ), .B(_GFM_N2239 ), .Z(_GFM_n12780 ) );
XOR2_X2 _GFM_U3161  ( .A(_GFM_N2233 ), .B(_GFM_N2235 ), .Z(_GFM_n12790 ) );
XOR2_X2 _GFM_U3160  ( .A(_GFM_n12810 ), .B(_GFM_n1280 ), .Z(z_out[73]) );
XOR2_X2 _GFM_U3159  ( .A(_GFM_n1283 ), .B(_GFM_n12820 ), .Z(_GFM_n1280 ) );
XOR2_X2 _GFM_U3158  ( .A(_GFM_n1285 ), .B(_GFM_n1284 ), .Z(_GFM_n12810 ) );
XOR2_X2 _GFM_U3157  ( .A(_GFM_n12870 ), .B(_GFM_n12860 ), .Z(_GFM_n12820 ));
XOR2_X2 _GFM_U3156  ( .A(_GFM_n12890 ), .B(_GFM_n1288 ), .Z(_GFM_n1283 ) );
XOR2_X2 _GFM_U3155  ( .A(_GFM_n12910 ), .B(_GFM_n1290 ), .Z(_GFM_n1284 ) );
XOR2_X2 _GFM_U3154  ( .A(_GFM_n1293 ), .B(_GFM_n12920 ), .Z(_GFM_n1285 ) );
XOR2_X2 _GFM_U3153  ( .A(z_in[73]), .B(_GFM_n1294 ), .Z(_GFM_n12860 ) );
XOR2_X2 _GFM_U3152  ( .A(_GFM_N2290 ), .B(_GFM_N2291 ), .Z(_GFM_n12870 ) );
XOR2_X2 _GFM_U3151  ( .A(_GFM_N2287 ), .B(_GFM_N2288 ), .Z(_GFM_n1288 ) );
XOR2_X2 _GFM_U3150  ( .A(_GFM_N2283 ), .B(_GFM_N2284 ), .Z(_GFM_n12890 ) );
XOR2_X2 _GFM_U3149  ( .A(_GFM_N2279 ), .B(_GFM_N2281 ), .Z(_GFM_n1290 ) );
XOR2_X2 _GFM_U3148  ( .A(_GFM_N2274 ), .B(_GFM_N2278 ), .Z(_GFM_n12910 ) );
XOR2_X2 _GFM_U3147  ( .A(_GFM_N2271 ), .B(_GFM_N2273 ), .Z(_GFM_n12920 ) );
XOR2_X2 _GFM_U3146  ( .A(_GFM_N2267 ), .B(_GFM_N2270 ), .Z(_GFM_n1293 ) );
XOR2_X2 _GFM_U3145  ( .A(_GFM_N2264 ), .B(_GFM_N2266 ), .Z(_GFM_n1294 ) );
XOR2_X2 _GFM_U3144  ( .A(_GFM_n12960 ), .B(_GFM_n12950 ), .Z(z_out[74]) );
XOR2_X2 _GFM_U3143  ( .A(_GFM_n12980 ), .B(_GFM_n1297 ), .Z(_GFM_n12950 ) );
XOR2_X2 _GFM_U3142  ( .A(_GFM_n1300 ), .B(_GFM_n12990 ), .Z(_GFM_n12960 ) );
XOR2_X2 _GFM_U3141  ( .A(_GFM_n1302 ), .B(_GFM_n1301 ), .Z(_GFM_n1297 ) );
XOR2_X2 _GFM_U3140  ( .A(_GFM_n1304 ), .B(_GFM_n13030 ), .Z(_GFM_n12980 ) );
XOR2_X2 _GFM_U3139  ( .A(_GFM_n13060 ), .B(_GFM_n13050 ), .Z(_GFM_n12990 ));
XOR2_X2 _GFM_U3138  ( .A(_GFM_n1308 ), .B(_GFM_n1307 ), .Z(_GFM_n1300 ) );
XOR2_X2 _GFM_U3137  ( .A(z_in[74]), .B(_GFM_n13090 ), .Z(_GFM_n1301 ) );
XOR2_X2 _GFM_U3136  ( .A(_GFM_N2321 ), .B(_GFM_N2322 ), .Z(_GFM_n1302 ) );
XOR2_X2 _GFM_U3135  ( .A(_GFM_N2318 ), .B(_GFM_N2319 ), .Z(_GFM_n13030 ) );
XOR2_X2 _GFM_U3134  ( .A(_GFM_N2314 ), .B(_GFM_N2315 ), .Z(_GFM_n1304 ) );
XOR2_X2 _GFM_U3133  ( .A(_GFM_N2310 ), .B(_GFM_N2312 ), .Z(_GFM_n13050 ) );
XOR2_X2 _GFM_U3132  ( .A(_GFM_N2305 ), .B(_GFM_N2309 ), .Z(_GFM_n13060 ) );
XOR2_X2 _GFM_U3131  ( .A(_GFM_N2302 ), .B(_GFM_N2304 ), .Z(_GFM_n1307 ) );
XOR2_X2 _GFM_U3130  ( .A(_GFM_N2298 ), .B(_GFM_N2301 ), .Z(_GFM_n1308 ) );
XOR2_X2 _GFM_U3129  ( .A(_GFM_N2295 ), .B(_GFM_N2297 ), .Z(_GFM_n13090 ) );
XOR2_X2 _GFM_U3128  ( .A(_GFM_n1311 ), .B(_GFM_n13100 ), .Z(z_out[75]) );
XOR2_X2 _GFM_U3127  ( .A(_GFM_n13130 ), .B(_GFM_n13120 ), .Z(_GFM_n13100 ));
XOR2_X2 _GFM_U3126  ( .A(_GFM_n1315 ), .B(_GFM_n1314 ), .Z(_GFM_n1311 ) );
XOR2_X2 _GFM_U3125  ( .A(_GFM_n13170 ), .B(_GFM_n1316 ), .Z(_GFM_n13120 ) );
XOR2_X2 _GFM_U3124  ( .A(_GFM_n1319 ), .B(_GFM_n13180 ), .Z(_GFM_n13130 ) );
XOR2_X2 _GFM_U3123  ( .A(_GFM_n1321 ), .B(_GFM_n13200 ), .Z(_GFM_n1314 ) );
XOR2_X2 _GFM_U3122  ( .A(_GFM_n13230 ), .B(_GFM_n13220 ), .Z(_GFM_n1315 ) );
XOR2_X2 _GFM_U3121  ( .A(z_in[75]), .B(_GFM_n1324 ), .Z(_GFM_n1316 ) );
XOR2_X2 _GFM_U3120  ( .A(_GFM_N2352 ), .B(_GFM_N2353 ), .Z(_GFM_n13170 ) );
XOR2_X2 _GFM_U3119  ( .A(_GFM_N2349 ), .B(_GFM_N2350 ), .Z(_GFM_n13180 ) );
XOR2_X2 _GFM_U3118  ( .A(_GFM_N2345 ), .B(_GFM_N2346 ), .Z(_GFM_n1319 ) );
XOR2_X2 _GFM_U3117  ( .A(_GFM_N2341 ), .B(_GFM_N2343 ), .Z(_GFM_n13200 ) );
XOR2_X2 _GFM_U3116  ( .A(_GFM_N2336 ), .B(_GFM_N2340 ), .Z(_GFM_n1321 ) );
XOR2_X2 _GFM_U3115  ( .A(_GFM_N2333 ), .B(_GFM_N2335 ), .Z(_GFM_n13220 ) );
XOR2_X2 _GFM_U3114  ( .A(_GFM_N2329 ), .B(_GFM_N2332 ), .Z(_GFM_n13230 ) );
XOR2_X2 _GFM_U3113  ( .A(_GFM_N2326 ), .B(_GFM_N2328 ), .Z(_GFM_n1324 ) );
XOR2_X2 _GFM_U3112  ( .A(_GFM_n13260 ), .B(_GFM_n1325 ), .Z(z_out[76]) );
XOR2_X2 _GFM_U3111  ( .A(_GFM_n1328 ), .B(_GFM_n13270 ), .Z(_GFM_n1325 ) );
XOR2_X2 _GFM_U3110  ( .A(_GFM_n13300 ), .B(_GFM_n13290 ), .Z(_GFM_n13260 ));
XOR2_X2 _GFM_U3109  ( .A(_GFM_n1332 ), .B(_GFM_n1331 ), .Z(_GFM_n13270 ) );
XOR2_X2 _GFM_U3108  ( .A(_GFM_n13340 ), .B(_GFM_n1333 ), .Z(_GFM_n1328 ) );
XOR2_X2 _GFM_U3107  ( .A(_GFM_n13360 ), .B(_GFM_n1335 ), .Z(_GFM_n13290 ) );
XOR2_X2 _GFM_U3106  ( .A(_GFM_n1338 ), .B(_GFM_n13370 ), .Z(_GFM_n13300 ) );
XOR2_X2 _GFM_U3105  ( .A(z_in[76]), .B(_GFM_n1339 ), .Z(_GFM_n1331 ) );
XOR2_X2 _GFM_U3104  ( .A(_GFM_N2383 ), .B(_GFM_N2384 ), .Z(_GFM_n1332 ) );
XOR2_X2 _GFM_U3103  ( .A(_GFM_N2380 ), .B(_GFM_N2381 ), .Z(_GFM_n1333 ) );
XOR2_X2 _GFM_U3102  ( .A(_GFM_N2376 ), .B(_GFM_N2377 ), .Z(_GFM_n13340 ) );
XOR2_X2 _GFM_U3101  ( .A(_GFM_N2372 ), .B(_GFM_N2374 ), .Z(_GFM_n1335 ) );
XOR2_X2 _GFM_U3100  ( .A(_GFM_N2367 ), .B(_GFM_N2371 ), .Z(_GFM_n13360 ) );
XOR2_X2 _GFM_U3099  ( .A(_GFM_N2364 ), .B(_GFM_N2366 ), .Z(_GFM_n13370 ) );
XOR2_X2 _GFM_U3098  ( .A(_GFM_N2360 ), .B(_GFM_N2363 ), .Z(_GFM_n1338 ) );
XOR2_X2 _GFM_U3097  ( .A(_GFM_N2357 ), .B(_GFM_N2359 ), .Z(_GFM_n1339 ) );
XOR2_X2 _GFM_U3096  ( .A(_GFM_n13410 ), .B(_GFM_n13400 ), .Z(z_out[77]) );
XOR2_X2 _GFM_U3095  ( .A(_GFM_n13430 ), .B(_GFM_n1342 ), .Z(_GFM_n13400 ) );
XOR2_X2 _GFM_U3094  ( .A(_GFM_n1345 ), .B(_GFM_n13440 ), .Z(_GFM_n13410 ) );
XOR2_X2 _GFM_U3093  ( .A(_GFM_n1347 ), .B(_GFM_n1346 ), .Z(_GFM_n1342 ) );
XOR2_X2 _GFM_U3092  ( .A(_GFM_n13490 ), .B(_GFM_n13480 ), .Z(_GFM_n13430 ));
XOR2_X2 _GFM_U3091  ( .A(_GFM_n13510 ), .B(_GFM_n1350 ), .Z(_GFM_n13440 ) );
XOR2_X2 _GFM_U3090  ( .A(_GFM_n13530 ), .B(_GFM_n1352 ), .Z(_GFM_n1345 ) );
XOR2_X2 _GFM_U3089  ( .A(z_in[77]), .B(_GFM_n13540 ), .Z(_GFM_n1346 ) );
XOR2_X2 _GFM_U3088  ( .A(_GFM_N2414 ), .B(_GFM_N2415 ), .Z(_GFM_n1347 ) );
XOR2_X2 _GFM_U3087  ( .A(_GFM_N2411 ), .B(_GFM_N2412 ), .Z(_GFM_n13480 ) );
XOR2_X2 _GFM_U3086  ( .A(_GFM_N2407 ), .B(_GFM_N2408 ), .Z(_GFM_n13490 ) );
XOR2_X2 _GFM_U3085  ( .A(_GFM_N2403 ), .B(_GFM_N2405 ), .Z(_GFM_n1350 ) );
XOR2_X2 _GFM_U3084  ( .A(_GFM_N2398 ), .B(_GFM_N2402 ), .Z(_GFM_n13510 ) );
XOR2_X2 _GFM_U3083  ( .A(_GFM_N2395 ), .B(_GFM_N2397 ), .Z(_GFM_n1352 ) );
XOR2_X2 _GFM_U3082  ( .A(_GFM_N2391 ), .B(_GFM_N2394 ), .Z(_GFM_n13530 ) );
XOR2_X2 _GFM_U3081  ( .A(_GFM_N2388 ), .B(_GFM_N2390 ), .Z(_GFM_n13540 ) );
XOR2_X2 _GFM_U3080  ( .A(_GFM_n1356 ), .B(_GFM_n1355 ), .Z(z_out[78]) );
XOR2_X2 _GFM_U3079  ( .A(_GFM_n13580 ), .B(_GFM_n13570 ), .Z(_GFM_n1355 ) );
XOR2_X2 _GFM_U3078  ( .A(_GFM_n13600 ), .B(_GFM_n1359 ), .Z(_GFM_n1356 ) );
XOR2_X2 _GFM_U3077  ( .A(_GFM_n1362 ), .B(_GFM_n13610 ), .Z(_GFM_n13570 ) );
XOR2_X2 _GFM_U3076  ( .A(_GFM_n1364 ), .B(_GFM_n1363 ), .Z(_GFM_n13580 ) );
XOR2_X2 _GFM_U3075  ( .A(_GFM_n1366 ), .B(_GFM_n13650 ), .Z(_GFM_n1359 ) );
XOR2_X2 _GFM_U3074  ( .A(_GFM_n13680 ), .B(_GFM_n13670 ), .Z(_GFM_n13600 ));
XOR2_X2 _GFM_U3073  ( .A(z_in[78]), .B(_GFM_n1369 ), .Z(_GFM_n13610 ) );
XOR2_X2 _GFM_U3072  ( .A(_GFM_N2445 ), .B(_GFM_N2446 ), .Z(_GFM_n1362 ) );
XOR2_X2 _GFM_U3071  ( .A(_GFM_N2442 ), .B(_GFM_N2443 ), .Z(_GFM_n1363 ) );
XOR2_X2 _GFM_U3070  ( .A(_GFM_N2438 ), .B(_GFM_N2439 ), .Z(_GFM_n1364 ) );
XOR2_X2 _GFM_U3069  ( .A(_GFM_N2434 ), .B(_GFM_N2436 ), .Z(_GFM_n13650 ) );
XOR2_X2 _GFM_U3068  ( .A(_GFM_N2429 ), .B(_GFM_N2433 ), .Z(_GFM_n1366 ) );
XOR2_X2 _GFM_U3067  ( .A(_GFM_N2426 ), .B(_GFM_N2428 ), .Z(_GFM_n13670 ) );
XOR2_X2 _GFM_U3066  ( .A(_GFM_N2422 ), .B(_GFM_N2425 ), .Z(_GFM_n13680 ) );
XOR2_X2 _GFM_U3065  ( .A(_GFM_N2419 ), .B(_GFM_N2421 ), .Z(_GFM_n1369 ) );
XOR2_X2 _GFM_U3064  ( .A(_GFM_n13710 ), .B(_GFM_n1370 ), .Z(z_out[79]) );
XOR2_X2 _GFM_U3063  ( .A(_GFM_n1373 ), .B(_GFM_n13720 ), .Z(_GFM_n1370 ) );
XOR2_X2 _GFM_U3062  ( .A(_GFM_n13750 ), .B(_GFM_n13740 ), .Z(_GFM_n13710 ));
XOR2_X2 _GFM_U3061  ( .A(_GFM_n1377 ), .B(_GFM_n1376 ), .Z(_GFM_n13720 ) );
XOR2_X2 _GFM_U3060  ( .A(_GFM_n13790 ), .B(_GFM_n1378 ), .Z(_GFM_n1373 ) );
XOR2_X2 _GFM_U3059  ( .A(_GFM_n1381 ), .B(_GFM_n13800 ), .Z(_GFM_n13740 ) );
XOR2_X2 _GFM_U3058  ( .A(_GFM_n1383 ), .B(_GFM_n13820 ), .Z(_GFM_n13750 ) );
XOR2_X2 _GFM_U3057  ( .A(z_in[79]), .B(_GFM_n13840 ), .Z(_GFM_n1376 ) );
XOR2_X2 _GFM_U3056  ( .A(_GFM_N2476 ), .B(_GFM_N2477 ), .Z(_GFM_n1377 ) );
XOR2_X2 _GFM_U3055  ( .A(_GFM_N2473 ), .B(_GFM_N2474 ), .Z(_GFM_n1378 ) );
XOR2_X2 _GFM_U3054  ( .A(_GFM_N2469 ), .B(_GFM_N2470 ), .Z(_GFM_n13790 ) );
XOR2_X2 _GFM_U3053  ( .A(_GFM_N2465 ), .B(_GFM_N2467 ), .Z(_GFM_n13800 ) );
XOR2_X2 _GFM_U3052  ( .A(_GFM_N2460 ), .B(_GFM_N2464 ), .Z(_GFM_n1381 ) );
XOR2_X2 _GFM_U3051  ( .A(_GFM_N2457 ), .B(_GFM_N2459 ), .Z(_GFM_n13820 ) );
XOR2_X2 _GFM_U3050  ( .A(_GFM_N2453 ), .B(_GFM_N2456 ), .Z(_GFM_n1383 ) );
XOR2_X2 _GFM_U3049  ( .A(_GFM_N2450 ), .B(_GFM_N2452 ), .Z(_GFM_n13840 ) );
XOR2_X2 _GFM_U3048  ( .A(_GFM_n1386 ), .B(_GFM_n13850 ), .Z(z_out[80]) );
XOR2_X2 _GFM_U3047  ( .A(_GFM_n13880 ), .B(_GFM_n1387 ), .Z(_GFM_n13850 ) );
XOR2_X2 _GFM_U3046  ( .A(_GFM_n1390 ), .B(_GFM_n13890 ), .Z(_GFM_n1386 ) );
XOR2_X2 _GFM_U3045  ( .A(_GFM_n13920 ), .B(_GFM_n13910 ), .Z(_GFM_n1387 ) );
XOR2_X2 _GFM_U3044  ( .A(_GFM_n1394 ), .B(_GFM_n1393 ), .Z(_GFM_n13880 ) );
XOR2_X2 _GFM_U3043  ( .A(_GFM_n13960 ), .B(_GFM_n1395 ), .Z(_GFM_n13890 ) );
XOR2_X2 _GFM_U3042  ( .A(_GFM_n13980 ), .B(_GFM_n1397 ), .Z(_GFM_n1390 ) );
XOR2_X2 _GFM_U3041  ( .A(z_in[80]), .B(_GFM_n13990 ), .Z(_GFM_n13910 ) );
XOR2_X2 _GFM_U3040  ( .A(_GFM_N2507 ), .B(_GFM_N2508 ), .Z(_GFM_n13920 ) );
XOR2_X2 _GFM_U3039  ( .A(_GFM_N2504 ), .B(_GFM_N2505 ), .Z(_GFM_n1393 ) );
XOR2_X2 _GFM_U3038  ( .A(_GFM_N2500 ), .B(_GFM_N2501 ), .Z(_GFM_n1394 ) );
XOR2_X2 _GFM_U3037  ( .A(_GFM_N2496 ), .B(_GFM_N2498 ), .Z(_GFM_n1395 ) );
XOR2_X2 _GFM_U3036  ( .A(_GFM_N2491 ), .B(_GFM_N2495 ), .Z(_GFM_n13960 ) );
XOR2_X2 _GFM_U3035  ( .A(_GFM_N2488 ), .B(_GFM_N2490 ), .Z(_GFM_n1397 ) );
XOR2_X2 _GFM_U3034  ( .A(_GFM_N2484 ), .B(_GFM_N2487 ), .Z(_GFM_n13980 ) );
XOR2_X2 _GFM_U3033  ( .A(_GFM_N2481 ), .B(_GFM_N2483 ), .Z(_GFM_n13990 ) );
XOR2_X2 _GFM_U3032  ( .A(_GFM_n1401 ), .B(_GFM_n1400 ), .Z(z_out[81]) );
XOR2_X2 _GFM_U3031  ( .A(_GFM_n14030 ), .B(_GFM_n14020 ), .Z(_GFM_n1400 ) );
XOR2_X2 _GFM_U3030  ( .A(_GFM_n14050 ), .B(_GFM_n1404 ), .Z(_GFM_n1401 ) );
XOR2_X2 _GFM_U3029  ( .A(_GFM_n1407 ), .B(_GFM_n14060 ), .Z(_GFM_n14020 ) );
XOR2_X2 _GFM_U3028  ( .A(_GFM_n1409 ), .B(_GFM_n1408 ), .Z(_GFM_n14030 ) );
XOR2_X2 _GFM_U3027  ( .A(_GFM_n14110 ), .B(_GFM_n14100 ), .Z(_GFM_n1404 ) );
XOR2_X2 _GFM_U3026  ( .A(_GFM_n14130 ), .B(_GFM_n1412 ), .Z(_GFM_n14050 ) );
XOR2_X2 _GFM_U3025  ( .A(z_in[81]), .B(_GFM_n1414 ), .Z(_GFM_n14060 ) );
XOR2_X2 _GFM_U3024  ( .A(_GFM_N2538 ), .B(_GFM_N2539 ), .Z(_GFM_n1407 ) );
XOR2_X2 _GFM_U3023  ( .A(_GFM_N2535 ), .B(_GFM_N2536 ), .Z(_GFM_n1408 ) );
XOR2_X2 _GFM_U3022  ( .A(_GFM_N2531 ), .B(_GFM_N2532 ), .Z(_GFM_n1409 ) );
XOR2_X2 _GFM_U3021  ( .A(_GFM_N2527 ), .B(_GFM_N2529 ), .Z(_GFM_n14100 ) );
XOR2_X2 _GFM_U3020  ( .A(_GFM_N2522 ), .B(_GFM_N2526 ), .Z(_GFM_n14110 ) );
XOR2_X2 _GFM_U3019  ( .A(_GFM_N2519 ), .B(_GFM_N2521 ), .Z(_GFM_n1412 ) );
XOR2_X2 _GFM_U3018  ( .A(_GFM_N2515 ), .B(_GFM_N2518 ), .Z(_GFM_n14130 ) );
XOR2_X2 _GFM_U3017  ( .A(_GFM_N2512 ), .B(_GFM_N2514 ), .Z(_GFM_n1414 ) );
XOR2_X2 _GFM_U3016  ( .A(_GFM_n14160 ), .B(_GFM_n14150 ), .Z(z_out[82]) );
XOR2_X2 _GFM_U3015  ( .A(_GFM_n1418 ), .B(_GFM_n1417 ), .Z(_GFM_n14150 ) );
XOR2_X2 _GFM_U3014  ( .A(_GFM_n14200 ), .B(_GFM_n14190 ), .Z(_GFM_n14160 ));
XOR2_X2 _GFM_U3013  ( .A(_GFM_n14220 ), .B(_GFM_n1421 ), .Z(_GFM_n1417 ) );
XOR2_X2 _GFM_U3012  ( .A(_GFM_n1424 ), .B(_GFM_n14230 ), .Z(_GFM_n1418 ) );
XOR2_X2 _GFM_U3011  ( .A(_GFM_n1426 ), .B(_GFM_n1425 ), .Z(_GFM_n14190 ) );
XOR2_X2 _GFM_U3010  ( .A(_GFM_n1428 ), .B(_GFM_n14270 ), .Z(_GFM_n14200 ) );
XOR2_X2 _GFM_U3009  ( .A(z_in[82]), .B(_GFM_n14290 ), .Z(_GFM_n1421 ) );
XOR2_X2 _GFM_U3008  ( .A(_GFM_N2569 ), .B(_GFM_N2570 ), .Z(_GFM_n14220 ) );
XOR2_X2 _GFM_U3007  ( .A(_GFM_N2566 ), .B(_GFM_N2567 ), .Z(_GFM_n14230 ) );
XOR2_X2 _GFM_U3006  ( .A(_GFM_N2562 ), .B(_GFM_N2563 ), .Z(_GFM_n1424 ) );
XOR2_X2 _GFM_U3005  ( .A(_GFM_N2558 ), .B(_GFM_N2560 ), .Z(_GFM_n1425 ) );
XOR2_X2 _GFM_U3004  ( .A(_GFM_N2553 ), .B(_GFM_N2557 ), .Z(_GFM_n1426 ) );
XOR2_X2 _GFM_U3003  ( .A(_GFM_N2550 ), .B(_GFM_N2552 ), .Z(_GFM_n14270 ) );
XOR2_X2 _GFM_U3002  ( .A(_GFM_N2546 ), .B(_GFM_N2549 ), .Z(_GFM_n1428 ) );
XOR2_X2 _GFM_U3001  ( .A(_GFM_N2543 ), .B(_GFM_N2545 ), .Z(_GFM_n14290 ) );
XOR2_X2 _GFM_U3000  ( .A(_GFM_n1431 ), .B(_GFM_n14300 ), .Z(z_out[83]) );
XOR2_X2 _GFM_U2999  ( .A(_GFM_n14330 ), .B(_GFM_n1432 ), .Z(_GFM_n14300 ) );
XOR2_X2 _GFM_U2998  ( .A(_GFM_n1435 ), .B(_GFM_n14340 ), .Z(_GFM_n1431 ) );
XOR2_X2 _GFM_U2997  ( .A(_GFM_n14370 ), .B(_GFM_n14360 ), .Z(_GFM_n1432 ) );
XOR2_X2 _GFM_U2996  ( .A(_GFM_n1439 ), .B(_GFM_n1438 ), .Z(_GFM_n14330 ) );
XOR2_X2 _GFM_U2995  ( .A(_GFM_n14410 ), .B(_GFM_n1440 ), .Z(_GFM_n14340 ) );
XOR2_X2 _GFM_U2994  ( .A(_GFM_n1443 ), .B(_GFM_n14420 ), .Z(_GFM_n1435 ) );
XOR2_X2 _GFM_U2993  ( .A(z_in[83]), .B(_GFM_n14440 ), .Z(_GFM_n14360 ) );
XOR2_X2 _GFM_U2992  ( .A(_GFM_N2600 ), .B(_GFM_N2601 ), .Z(_GFM_n14370 ) );
XOR2_X2 _GFM_U2991  ( .A(_GFM_N2597 ), .B(_GFM_N2598 ), .Z(_GFM_n1438 ) );
XOR2_X2 _GFM_U2990  ( .A(_GFM_N2593 ), .B(_GFM_N2594 ), .Z(_GFM_n1439 ) );
XOR2_X2 _GFM_U2989  ( .A(_GFM_N2589 ), .B(_GFM_N2591 ), .Z(_GFM_n1440 ) );
XOR2_X2 _GFM_U2988  ( .A(_GFM_N2584 ), .B(_GFM_N2588 ), .Z(_GFM_n14410 ) );
XOR2_X2 _GFM_U2987  ( .A(_GFM_N2581 ), .B(_GFM_N2583 ), .Z(_GFM_n14420 ) );
XOR2_X2 _GFM_U2986  ( .A(_GFM_N2577 ), .B(_GFM_N2580 ), .Z(_GFM_n1443 ) );
XOR2_X2 _GFM_U2985  ( .A(_GFM_N2574 ), .B(_GFM_N2576 ), .Z(_GFM_n14440 ) );
XOR2_X2 _GFM_U2984  ( .A(_GFM_n14460 ), .B(_GFM_n1445 ), .Z(z_out[84]) );
XOR2_X2 _GFM_U2983  ( .A(_GFM_n1448 ), .B(_GFM_n14470 ), .Z(_GFM_n1445 ) );
XOR2_X2 _GFM_U2982  ( .A(_GFM_n14500 ), .B(_GFM_n1449 ), .Z(_GFM_n14460 ) );
XOR2_X2 _GFM_U2981  ( .A(_GFM_n1452 ), .B(_GFM_n14510 ), .Z(_GFM_n14470 ) );
XOR2_X2 _GFM_U2980  ( .A(_GFM_n14540 ), .B(_GFM_n14530 ), .Z(_GFM_n1448 ) );
XOR2_X2 _GFM_U2979  ( .A(_GFM_n1456 ), .B(_GFM_n1455 ), .Z(_GFM_n1449 ) );
XOR2_X2 _GFM_U2978  ( .A(_GFM_n14580 ), .B(_GFM_n1457 ), .Z(_GFM_n14500 ) );
XOR2_X2 _GFM_U2977  ( .A(z_in[84]), .B(_GFM_n1459 ), .Z(_GFM_n14510 ) );
XOR2_X2 _GFM_U2976  ( .A(_GFM_N2631 ), .B(_GFM_N2632 ), .Z(_GFM_n1452 ) );
XOR2_X2 _GFM_U2975  ( .A(_GFM_N2628 ), .B(_GFM_N2629 ), .Z(_GFM_n14530 ) );
XOR2_X2 _GFM_U2974  ( .A(_GFM_N2624 ), .B(_GFM_N2625 ), .Z(_GFM_n14540 ) );
XOR2_X2 _GFM_U2973  ( .A(_GFM_N2620 ), .B(_GFM_N2622 ), .Z(_GFM_n1455 ) );
XOR2_X2 _GFM_U2972  ( .A(_GFM_N2615 ), .B(_GFM_N2619 ), .Z(_GFM_n1456 ) );
XOR2_X2 _GFM_U2971  ( .A(_GFM_N2612 ), .B(_GFM_N2614 ), .Z(_GFM_n1457 ) );
XOR2_X2 _GFM_U2970  ( .A(_GFM_N2608 ), .B(_GFM_N2611 ), .Z(_GFM_n14580 ) );
XOR2_X2 _GFM_U2969  ( .A(_GFM_N2605 ), .B(_GFM_N2607 ), .Z(_GFM_n1459 ) );
XOR2_X2 _GFM_U2968  ( .A(_GFM_n14610 ), .B(_GFM_n14600 ), .Z(z_out[85]) );
XOR2_X2 _GFM_U2967  ( .A(_GFM_n1463 ), .B(_GFM_n1462 ), .Z(_GFM_n14600 ) );
XOR2_X2 _GFM_U2966  ( .A(_GFM_n14650 ), .B(_GFM_n14640 ), .Z(_GFM_n14610 ));
XOR2_X2 _GFM_U2965  ( .A(_GFM_n14670 ), .B(_GFM_n1466 ), .Z(_GFM_n1462 ) );
XOR2_X2 _GFM_U2964  ( .A(_GFM_n1469 ), .B(_GFM_n14680 ), .Z(_GFM_n1463 ) );
XOR2_X2 _GFM_U2963  ( .A(_GFM_n1471 ), .B(_GFM_n1470 ), .Z(_GFM_n14640 ) );
XOR2_X2 _GFM_U2962  ( .A(_GFM_n14730 ), .B(_GFM_n14720 ), .Z(_GFM_n14650 ));
XOR2_X2 _GFM_U2961  ( .A(z_in[85]), .B(_GFM_n1474 ), .Z(_GFM_n1466 ) );
XOR2_X2 _GFM_U2960  ( .A(_GFM_N2662 ), .B(_GFM_N2663 ), .Z(_GFM_n14670 ) );
XOR2_X2 _GFM_U2959  ( .A(_GFM_N2659 ), .B(_GFM_N2660 ), .Z(_GFM_n14680 ) );
XOR2_X2 _GFM_U2958  ( .A(_GFM_N2655 ), .B(_GFM_N2656 ), .Z(_GFM_n1469 ) );
XOR2_X2 _GFM_U2957  ( .A(_GFM_N2651 ), .B(_GFM_N2653 ), .Z(_GFM_n1470 ) );
XOR2_X2 _GFM_U2956  ( .A(_GFM_N2646 ), .B(_GFM_N2650 ), .Z(_GFM_n1471 ) );
XOR2_X2 _GFM_U2955  ( .A(_GFM_N2643 ), .B(_GFM_N2645 ), .Z(_GFM_n14720 ) );
XOR2_X2 _GFM_U2954  ( .A(_GFM_N2639 ), .B(_GFM_N2642 ), .Z(_GFM_n14730 ) );
XOR2_X2 _GFM_U2953  ( .A(_GFM_N2636 ), .B(_GFM_N2638 ), .Z(_GFM_n1474 ) );
XOR2_X2 _GFM_U2952  ( .A(_GFM_n1476 ), .B(_GFM_n14750 ), .Z(z_out[86]) );
XOR2_X2 _GFM_U2951  ( .A(_GFM_n14780 ), .B(_GFM_n14770 ), .Z(_GFM_n14750 ));
XOR2_X2 _GFM_U2950  ( .A(_GFM_n1480 ), .B(_GFM_n1479 ), .Z(_GFM_n1476 ) );
XOR2_X2 _GFM_U2949  ( .A(_GFM_n14820 ), .B(_GFM_n14810 ), .Z(_GFM_n14770 ));
XOR2_X2 _GFM_U2948  ( .A(_GFM_n14840 ), .B(_GFM_n1483 ), .Z(_GFM_n14780 ) );
XOR2_X2 _GFM_U2947  ( .A(_GFM_n1486 ), .B(_GFM_n14850 ), .Z(_GFM_n1479 ) );
XOR2_X2 _GFM_U2946  ( .A(_GFM_n1488 ), .B(_GFM_n1487 ), .Z(_GFM_n1480 ) );
XOR2_X2 _GFM_U2945  ( .A(z_in[86]), .B(_GFM_n14890 ), .Z(_GFM_n14810 ) );
XOR2_X2 _GFM_U2944  ( .A(_GFM_N2693 ), .B(_GFM_N2694 ), .Z(_GFM_n14820 ) );
XOR2_X2 _GFM_U2943  ( .A(_GFM_N2690 ), .B(_GFM_N2691 ), .Z(_GFM_n1483 ) );
XOR2_X2 _GFM_U2942  ( .A(_GFM_N2686 ), .B(_GFM_N2687 ), .Z(_GFM_n14840 ) );
XOR2_X2 _GFM_U2941  ( .A(_GFM_N2682 ), .B(_GFM_N2684 ), .Z(_GFM_n14850 ) );
XOR2_X2 _GFM_U2940  ( .A(_GFM_N2677 ), .B(_GFM_N2681 ), .Z(_GFM_n1486 ) );
XOR2_X2 _GFM_U2939  ( .A(_GFM_N2674 ), .B(_GFM_N2676 ), .Z(_GFM_n1487 ) );
XOR2_X2 _GFM_U2938  ( .A(_GFM_N2670 ), .B(_GFM_N2673 ), .Z(_GFM_n1488 ) );
XOR2_X2 _GFM_U2937  ( .A(_GFM_N2667 ), .B(_GFM_N2669 ), .Z(_GFM_n14890 ) );
XOR2_X2 _GFM_U2936  ( .A(_GFM_n14910 ), .B(_GFM_n1490 ), .Z(z_out[87]) );
XOR2_X2 _GFM_U2935  ( .A(_GFM_n1493 ), .B(_GFM_n14920 ), .Z(_GFM_n1490 ) );
XOR2_X2 _GFM_U2934  ( .A(_GFM_n14950 ), .B(_GFM_n1494 ), .Z(_GFM_n14910 ) );
XOR2_X2 _GFM_U2933  ( .A(_GFM_n1497 ), .B(_GFM_n14960 ), .Z(_GFM_n14920 ) );
XOR2_X2 _GFM_U2932  ( .A(_GFM_n14990 ), .B(_GFM_n14980 ), .Z(_GFM_n1493 ) );
XOR2_X2 _GFM_U2931  ( .A(_GFM_n1501 ), .B(_GFM_n1500 ), .Z(_GFM_n1494 ) );
XOR2_X2 _GFM_U2930  ( .A(_GFM_n15030 ), .B(_GFM_n1502 ), .Z(_GFM_n14950 ) );
XOR2_X2 _GFM_U2929  ( .A(z_in[87]), .B(_GFM_n15040 ), .Z(_GFM_n14960 ) );
XOR2_X2 _GFM_U2928  ( .A(_GFM_N2724 ), .B(_GFM_N2725 ), .Z(_GFM_n1497 ) );
XOR2_X2 _GFM_U2927  ( .A(_GFM_N2721 ), .B(_GFM_N2722 ), .Z(_GFM_n14980 ) );
XOR2_X2 _GFM_U2926  ( .A(_GFM_N2717 ), .B(_GFM_N2718 ), .Z(_GFM_n14990 ) );
XOR2_X2 _GFM_U2925  ( .A(_GFM_N2713 ), .B(_GFM_N2715 ), .Z(_GFM_n1500 ) );
XOR2_X2 _GFM_U2924  ( .A(_GFM_N2708 ), .B(_GFM_N2712 ), .Z(_GFM_n1501 ) );
XOR2_X2 _GFM_U2923  ( .A(_GFM_N2705 ), .B(_GFM_N2707 ), .Z(_GFM_n1502 ) );
XOR2_X2 _GFM_U2922  ( .A(_GFM_N2701 ), .B(_GFM_N2704 ), .Z(_GFM_n15030 ) );
XOR2_X2 _GFM_U2921  ( .A(_GFM_N2698 ), .B(_GFM_N2700 ), .Z(_GFM_n15040 ) );
XOR2_X2 _GFM_U2920  ( .A(_GFM_n15060 ), .B(_GFM_n1505 ), .Z(z_out[88]) );
XOR2_X2 _GFM_U2919  ( .A(_GFM_n15080 ), .B(_GFM_n1507 ), .Z(_GFM_n1505 ) );
XOR2_X2 _GFM_U2918  ( .A(_GFM_n1510 ), .B(_GFM_n15090 ), .Z(_GFM_n15060 ) );
XOR2_X2 _GFM_U2917  ( .A(_GFM_n15120 ), .B(_GFM_n1511 ), .Z(_GFM_n1507 ) );
XOR2_X2 _GFM_U2916  ( .A(_GFM_n1514 ), .B(_GFM_n15130 ), .Z(_GFM_n15080 ) );
XOR2_X2 _GFM_U2915  ( .A(_GFM_n15160 ), .B(_GFM_n15150 ), .Z(_GFM_n15090 ));
XOR2_X2 _GFM_U2914  ( .A(_GFM_n1518 ), .B(_GFM_n1517 ), .Z(_GFM_n1510 ) );
XOR2_X2 _GFM_U2913  ( .A(z_in[88]), .B(_GFM_n1519 ), .Z(_GFM_n1511 ) );
XOR2_X2 _GFM_U2912  ( .A(_GFM_N2755 ), .B(_GFM_N2756 ), .Z(_GFM_n15120 ) );
XOR2_X2 _GFM_U2911  ( .A(_GFM_N2752 ), .B(_GFM_N2753 ), .Z(_GFM_n15130 ) );
XOR2_X2 _GFM_U2910  ( .A(_GFM_N2748 ), .B(_GFM_N2749 ), .Z(_GFM_n1514 ) );
XOR2_X2 _GFM_U2909  ( .A(_GFM_N2744 ), .B(_GFM_N2746 ), .Z(_GFM_n15150 ) );
XOR2_X2 _GFM_U2908  ( .A(_GFM_N2739 ), .B(_GFM_N2743 ), .Z(_GFM_n15160 ) );
XOR2_X2 _GFM_U2907  ( .A(_GFM_N2736 ), .B(_GFM_N2738 ), .Z(_GFM_n1517 ) );
XOR2_X2 _GFM_U2906  ( .A(_GFM_N2732 ), .B(_GFM_N2735 ), .Z(_GFM_n1518 ) );
XOR2_X2 _GFM_U2905  ( .A(_GFM_N2729 ), .B(_GFM_N2731 ), .Z(_GFM_n1519 ) );
XOR2_X2 _GFM_U2904  ( .A(_GFM_n1521 ), .B(_GFM_n15200 ), .Z(z_out[89]) );
XOR2_X2 _GFM_U2903  ( .A(_GFM_n15230 ), .B(_GFM_n15220 ), .Z(_GFM_n15200 ));
XOR2_X2 _GFM_U2902  ( .A(_GFM_n1525 ), .B(_GFM_n1524 ), .Z(_GFM_n1521 ) );
XOR2_X2 _GFM_U2901  ( .A(_GFM_n15270 ), .B(_GFM_n15260 ), .Z(_GFM_n15220 ));
XOR2_X2 _GFM_U2900  ( .A(_GFM_n15290 ), .B(_GFM_n1528 ), .Z(_GFM_n15230 ) );
XOR2_X2 _GFM_U2899  ( .A(_GFM_n1531 ), .B(_GFM_n15300 ), .Z(_GFM_n1524 ) );
XOR2_X2 _GFM_U2898  ( .A(_GFM_n1533 ), .B(_GFM_n1532 ), .Z(_GFM_n1525 ) );
XOR2_X2 _GFM_U2897  ( .A(z_in[89]), .B(_GFM_n15340 ), .Z(_GFM_n15260 ) );
XOR2_X2 _GFM_U2896  ( .A(_GFM_N2786 ), .B(_GFM_N2787 ), .Z(_GFM_n15270 ) );
XOR2_X2 _GFM_U2895  ( .A(_GFM_N2783 ), .B(_GFM_N2784 ), .Z(_GFM_n1528 ) );
XOR2_X2 _GFM_U2894  ( .A(_GFM_N2779 ), .B(_GFM_N2780 ), .Z(_GFM_n15290 ) );
XOR2_X2 _GFM_U2893  ( .A(_GFM_N2775 ), .B(_GFM_N2777 ), .Z(_GFM_n15300 ) );
XOR2_X2 _GFM_U2892  ( .A(_GFM_N2770 ), .B(_GFM_N2774 ), .Z(_GFM_n1531 ) );
XOR2_X2 _GFM_U2891  ( .A(_GFM_N2767 ), .B(_GFM_N2769 ), .Z(_GFM_n1532 ) );
XOR2_X2 _GFM_U2890  ( .A(_GFM_N2763 ), .B(_GFM_N2766 ), .Z(_GFM_n1533 ) );
XOR2_X2 _GFM_U2889  ( .A(_GFM_N2760 ), .B(_GFM_N2762 ), .Z(_GFM_n15340 ) );
XOR2_X2 _GFM_U2888  ( .A(_GFM_n1536 ), .B(_GFM_n15350 ), .Z(z_out[90]) );
XOR2_X2 _GFM_U2887  ( .A(_GFM_n1538 ), .B(_GFM_n15370 ), .Z(_GFM_n15350 ) );
XOR2_X2 _GFM_U2886  ( .A(_GFM_n15400 ), .B(_GFM_n15390 ), .Z(_GFM_n1536 ) );
XOR2_X2 _GFM_U2885  ( .A(_GFM_n1542 ), .B(_GFM_n1541 ), .Z(_GFM_n15370 ) );
XOR2_X2 _GFM_U2884  ( .A(_GFM_n15440 ), .B(_GFM_n15430 ), .Z(_GFM_n1538 ) );
XOR2_X2 _GFM_U2883  ( .A(_GFM_n15460 ), .B(_GFM_n1545 ), .Z(_GFM_n15390 ) );
XOR2_X2 _GFM_U2882  ( .A(_GFM_n1548 ), .B(_GFM_n15470 ), .Z(_GFM_n15400 ) );
XOR2_X2 _GFM_U2881  ( .A(z_in[90]), .B(_GFM_n1549 ), .Z(_GFM_n1541 ) );
XOR2_X2 _GFM_U2880  ( .A(_GFM_N2817 ), .B(_GFM_N2818 ), .Z(_GFM_n1542 ) );
XOR2_X2 _GFM_U2879  ( .A(_GFM_N2814 ), .B(_GFM_N2815 ), .Z(_GFM_n15430 ) );
XOR2_X2 _GFM_U2878  ( .A(_GFM_N2810 ), .B(_GFM_N2811 ), .Z(_GFM_n15440 ) );
XOR2_X2 _GFM_U2877  ( .A(_GFM_N2806 ), .B(_GFM_N2808 ), .Z(_GFM_n1545 ) );
XOR2_X2 _GFM_U2876  ( .A(_GFM_N2801 ), .B(_GFM_N2805 ), .Z(_GFM_n15460 ) );
XOR2_X2 _GFM_U2875  ( .A(_GFM_N2798 ), .B(_GFM_N2800 ), .Z(_GFM_n15470 ) );
XOR2_X2 _GFM_U2874  ( .A(_GFM_N2794 ), .B(_GFM_N2797 ), .Z(_GFM_n1548 ) );
XOR2_X2 _GFM_U2873  ( .A(_GFM_N2791 ), .B(_GFM_N2793 ), .Z(_GFM_n1549 ) );
XOR2_X2 _GFM_U2872  ( .A(_GFM_n15510 ), .B(_GFM_n1550 ), .Z(z_out[91]) );
XOR2_X2 _GFM_U2871  ( .A(_GFM_n15530 ), .B(_GFM_n1552 ), .Z(_GFM_n1550 ) );
XOR2_X2 _GFM_U2870  ( .A(_GFM_n1555 ), .B(_GFM_n15540 ), .Z(_GFM_n15510 ) );
XOR2_X2 _GFM_U2869  ( .A(_GFM_n15570 ), .B(_GFM_n1556 ), .Z(_GFM_n1552 ) );
XOR2_X2 _GFM_U2868  ( .A(_GFM_n1559 ), .B(_GFM_n15580 ), .Z(_GFM_n15530 ) );
XOR2_X2 _GFM_U2867  ( .A(_GFM_n15610 ), .B(_GFM_n15600 ), .Z(_GFM_n15540 ));
XOR2_X2 _GFM_U2866  ( .A(_GFM_n1563 ), .B(_GFM_n1562 ), .Z(_GFM_n1555 ) );
XOR2_X2 _GFM_U2865  ( .A(z_in[91]), .B(_GFM_n1564 ), .Z(_GFM_n1556 ) );
XOR2_X2 _GFM_U2864  ( .A(_GFM_N2848 ), .B(_GFM_N2849 ), .Z(_GFM_n15570 ) );
XOR2_X2 _GFM_U2863  ( .A(_GFM_N2845 ), .B(_GFM_N2846 ), .Z(_GFM_n15580 ) );
XOR2_X2 _GFM_U2862  ( .A(_GFM_N2841 ), .B(_GFM_N2842 ), .Z(_GFM_n1559 ) );
XOR2_X2 _GFM_U2861  ( .A(_GFM_N2837 ), .B(_GFM_N2839 ), .Z(_GFM_n15600 ) );
XOR2_X2 _GFM_U2860  ( .A(_GFM_N2832 ), .B(_GFM_N2836 ), .Z(_GFM_n15610 ) );
XOR2_X2 _GFM_U2859  ( .A(_GFM_N2829 ), .B(_GFM_N2831 ), .Z(_GFM_n1562 ) );
XOR2_X2 _GFM_U2858  ( .A(_GFM_N2825 ), .B(_GFM_N2828 ), .Z(_GFM_n1563 ) );
XOR2_X2 _GFM_U2857  ( .A(_GFM_N2822 ), .B(_GFM_N2824 ), .Z(_GFM_n1564 ) );
XOR2_X2 _GFM_U2856  ( .A(_GFM_n15660 ), .B(_GFM_n15650 ), .Z(z_out[92]) );
XOR2_X2 _GFM_U2855  ( .A(_GFM_n15680 ), .B(_GFM_n1567 ), .Z(_GFM_n15650 ) );
XOR2_X2 _GFM_U2854  ( .A(_GFM_n15700 ), .B(_GFM_n1569 ), .Z(_GFM_n15660 ) );
XOR2_X2 _GFM_U2853  ( .A(_GFM_n1572 ), .B(_GFM_n15710 ), .Z(_GFM_n1567 ) );
XOR2_X2 _GFM_U2852  ( .A(_GFM_n15740 ), .B(_GFM_n1573 ), .Z(_GFM_n15680 ) );
XOR2_X2 _GFM_U2851  ( .A(_GFM_n1576 ), .B(_GFM_n15750 ), .Z(_GFM_n1569 ) );
XOR2_X2 _GFM_U2850  ( .A(_GFM_n15780 ), .B(_GFM_n15770 ), .Z(_GFM_n15700 ));
XOR2_X2 _GFM_U2849  ( .A(z_in[92]), .B(_GFM_n1579 ), .Z(_GFM_n15710 ) );
XOR2_X2 _GFM_U2848  ( .A(_GFM_N2879 ), .B(_GFM_N2880 ), .Z(_GFM_n1572 ) );
XOR2_X2 _GFM_U2847  ( .A(_GFM_N2876 ), .B(_GFM_N2877 ), .Z(_GFM_n1573 ) );
XOR2_X2 _GFM_U2846  ( .A(_GFM_N2872 ), .B(_GFM_N2873 ), .Z(_GFM_n15740 ) );
XOR2_X2 _GFM_U2845  ( .A(_GFM_N2868 ), .B(_GFM_N2870 ), .Z(_GFM_n15750 ) );
XOR2_X2 _GFM_U2844  ( .A(_GFM_N2863 ), .B(_GFM_N2867 ), .Z(_GFM_n1576 ) );
XOR2_X2 _GFM_U2843  ( .A(_GFM_N2860 ), .B(_GFM_N2862 ), .Z(_GFM_n15770 ) );
XOR2_X2 _GFM_U2842  ( .A(_GFM_N2856 ), .B(_GFM_N2859 ), .Z(_GFM_n15780 ) );
XOR2_X2 _GFM_U2841  ( .A(_GFM_N2853 ), .B(_GFM_N2855 ), .Z(_GFM_n1579 ) );
XOR2_X2 _GFM_U2840  ( .A(_GFM_n1581 ), .B(_GFM_n1580 ), .Z(z_out[93]) );
XOR2_X2 _GFM_U2839  ( .A(_GFM_n1583 ), .B(_GFM_n15820 ), .Z(_GFM_n1580 ) );
XOR2_X2 _GFM_U2838  ( .A(_GFM_n15850 ), .B(_GFM_n15840 ), .Z(_GFM_n1581 ) );
XOR2_X2 _GFM_U2837  ( .A(_GFM_n1587 ), .B(_GFM_n1586 ), .Z(_GFM_n15820 ) );
XOR2_X2 _GFM_U2836  ( .A(_GFM_n15890 ), .B(_GFM_n15880 ), .Z(_GFM_n1583 ) );
XOR2_X2 _GFM_U2835  ( .A(_GFM_n15910 ), .B(_GFM_n1590 ), .Z(_GFM_n15840 ) );
XOR2_X2 _GFM_U2834  ( .A(_GFM_n1593 ), .B(_GFM_n15920 ), .Z(_GFM_n15850 ) );
XOR2_X2 _GFM_U2833  ( .A(z_in[93]), .B(_GFM_n1594 ), .Z(_GFM_n1586 ) );
XOR2_X2 _GFM_U2832  ( .A(_GFM_N2910 ), .B(_GFM_N2911 ), .Z(_GFM_n1587 ) );
XOR2_X2 _GFM_U2831  ( .A(_GFM_N2907 ), .B(_GFM_N2908 ), .Z(_GFM_n15880 ) );
XOR2_X2 _GFM_U2830  ( .A(_GFM_N2903 ), .B(_GFM_N2904 ), .Z(_GFM_n15890 ) );
XOR2_X2 _GFM_U2829  ( .A(_GFM_N2899 ), .B(_GFM_N2901 ), .Z(_GFM_n1590 ) );
XOR2_X2 _GFM_U2828  ( .A(_GFM_N2894 ), .B(_GFM_N2898 ), .Z(_GFM_n15910 ) );
XOR2_X2 _GFM_U2827  ( .A(_GFM_N2891 ), .B(_GFM_N2893 ), .Z(_GFM_n15920 ) );
XOR2_X2 _GFM_U2826  ( .A(_GFM_N2887 ), .B(_GFM_N2890 ), .Z(_GFM_n1593 ) );
XOR2_X2 _GFM_U2825  ( .A(_GFM_N2884 ), .B(_GFM_N2886 ), .Z(_GFM_n1594 ) );
XOR2_X2 _GFM_U2824  ( .A(_GFM_n15960 ), .B(_GFM_n1595 ), .Z(z_out[94]) );
XOR2_X2 _GFM_U2823  ( .A(_GFM_n1598 ), .B(_GFM_n15970 ), .Z(_GFM_n1595 ) );
XOR2_X2 _GFM_U2822  ( .A(_GFM_n1600 ), .B(_GFM_n15990 ), .Z(_GFM_n15960 ) );
XOR2_X2 _GFM_U2821  ( .A(_GFM_n16020 ), .B(_GFM_n16010 ), .Z(_GFM_n15970 ));
XOR2_X2 _GFM_U2820  ( .A(_GFM_n1604 ), .B(_GFM_n1603 ), .Z(_GFM_n1598 ) );
XOR2_X2 _GFM_U2819  ( .A(_GFM_n16060 ), .B(_GFM_n16050 ), .Z(_GFM_n15990 ));
XOR2_X2 _GFM_U2818  ( .A(_GFM_n16080 ), .B(_GFM_n1607 ), .Z(_GFM_n1600 ) );
XOR2_X2 _GFM_U2817  ( .A(z_in[94]), .B(_GFM_n16090 ), .Z(_GFM_n16010 ) );
XOR2_X2 _GFM_U2816  ( .A(_GFM_N2941 ), .B(_GFM_N2942 ), .Z(_GFM_n16020 ) );
XOR2_X2 _GFM_U2815  ( .A(_GFM_N2938 ), .B(_GFM_N2939 ), .Z(_GFM_n1603 ) );
XOR2_X2 _GFM_U2814  ( .A(_GFM_N2934 ), .B(_GFM_N2935 ), .Z(_GFM_n1604 ) );
XOR2_X2 _GFM_U2813  ( .A(_GFM_N2930 ), .B(_GFM_N2932 ), .Z(_GFM_n16050 ) );
XOR2_X2 _GFM_U2812  ( .A(_GFM_N2925 ), .B(_GFM_N2929 ), .Z(_GFM_n16060 ) );
XOR2_X2 _GFM_U2811  ( .A(_GFM_N2922 ), .B(_GFM_N2924 ), .Z(_GFM_n1607 ) );
XOR2_X2 _GFM_U2810  ( .A(_GFM_N2918 ), .B(_GFM_N2921 ), .Z(_GFM_n16080 ) );
XOR2_X2 _GFM_U2809  ( .A(_GFM_N2915 ), .B(_GFM_N2917 ), .Z(_GFM_n16090 ) );
XOR2_X2 _GFM_U2808  ( .A(_GFM_n1611 ), .B(_GFM_n1610 ), .Z(z_out[95]) );
XOR2_X2 _GFM_U2807  ( .A(_GFM_n16130 ), .B(_GFM_n1612 ), .Z(_GFM_n1610 ) );
XOR2_X2 _GFM_U2806  ( .A(_GFM_n16150 ), .B(_GFM_n1614 ), .Z(_GFM_n1611 ) );
XOR2_X2 _GFM_U2805  ( .A(_GFM_n1617 ), .B(_GFM_n16160 ), .Z(_GFM_n1612 ) );
XOR2_X2 _GFM_U2804  ( .A(_GFM_n16190 ), .B(_GFM_n1618 ), .Z(_GFM_n16130 ) );
XOR2_X2 _GFM_U2803  ( .A(_GFM_n1621 ), .B(_GFM_n16200 ), .Z(_GFM_n1614 ) );
XOR2_X2 _GFM_U2802  ( .A(_GFM_n16230 ), .B(_GFM_n16220 ), .Z(_GFM_n16150 ));
XOR2_X2 _GFM_U2801  ( .A(z_in[95]), .B(_GFM_n1624 ), .Z(_GFM_n16160 ) );
XOR2_X2 _GFM_U2800  ( .A(_GFM_N2972 ), .B(_GFM_N2973 ), .Z(_GFM_n1617 ) );
XOR2_X2 _GFM_U2799  ( .A(_GFM_N2969 ), .B(_GFM_N2970 ), .Z(_GFM_n1618 ) );
XOR2_X2 _GFM_U2798  ( .A(_GFM_N2965 ), .B(_GFM_N2966 ), .Z(_GFM_n16190 ) );
XOR2_X2 _GFM_U2797  ( .A(_GFM_N2961 ), .B(_GFM_N2963 ), .Z(_GFM_n16200 ) );
XOR2_X2 _GFM_U2796  ( .A(_GFM_N2956 ), .B(_GFM_N2960 ), .Z(_GFM_n1621 ) );
XOR2_X2 _GFM_U2795  ( .A(_GFM_N2953 ), .B(_GFM_N2955 ), .Z(_GFM_n16220 ) );
XOR2_X2 _GFM_U2794  ( .A(_GFM_N2949 ), .B(_GFM_N2952 ), .Z(_GFM_n16230 ) );
XOR2_X2 _GFM_U2793  ( .A(_GFM_N2946 ), .B(_GFM_N2948 ), .Z(_GFM_n1624 ) );
XOR2_X2 _GFM_U2792  ( .A(_GFM_n1626 ), .B(_GFM_n1625 ), .Z(z_out[96]) );
XOR2_X2 _GFM_U2791  ( .A(_GFM_n16280 ), .B(_GFM_n16270 ), .Z(_GFM_n1625 ) );
XOR2_X2 _GFM_U2790  ( .A(_GFM_n16300 ), .B(_GFM_n1629 ), .Z(_GFM_n1626 ) );
XOR2_X2 _GFM_U2789  ( .A(_GFM_n16320 ), .B(_GFM_n1631 ), .Z(_GFM_n16270 ) );
XOR2_X2 _GFM_U2788  ( .A(_GFM_n1634 ), .B(_GFM_n16330 ), .Z(_GFM_n16280 ) );
XOR2_X2 _GFM_U2787  ( .A(_GFM_n16360 ), .B(_GFM_n1635 ), .Z(_GFM_n1629 ) );
XOR2_X2 _GFM_U2786  ( .A(_GFM_n1638 ), .B(_GFM_n16370 ), .Z(_GFM_n16300 ) );
XOR2_X2 _GFM_U2785  ( .A(z_in[96]), .B(_GFM_n16390 ), .Z(_GFM_n1631 ) );
XOR2_X2 _GFM_U2784  ( .A(_GFM_N3003 ), .B(_GFM_N3004 ), .Z(_GFM_n16320 ) );
XOR2_X2 _GFM_U2783  ( .A(_GFM_N3000 ), .B(_GFM_N3001 ), .Z(_GFM_n16330 ) );
XOR2_X2 _GFM_U2782  ( .A(_GFM_N2996 ), .B(_GFM_N2997 ), .Z(_GFM_n1634 ) );
XOR2_X2 _GFM_U2781  ( .A(_GFM_N2992 ), .B(_GFM_N2994 ), .Z(_GFM_n1635 ) );
XOR2_X2 _GFM_U2780  ( .A(_GFM_N2987 ), .B(_GFM_N2991 ), .Z(_GFM_n16360 ) );
XOR2_X2 _GFM_U2779  ( .A(_GFM_N2984 ), .B(_GFM_N2986 ), .Z(_GFM_n16370 ) );
XOR2_X2 _GFM_U2778  ( .A(_GFM_N2980 ), .B(_GFM_N2983 ), .Z(_GFM_n1638 ) );
XOR2_X2 _GFM_U2777  ( .A(_GFM_N2977 ), .B(_GFM_N2979 ), .Z(_GFM_n16390 ) );
XOR2_X2 _GFM_U2776  ( .A(_GFM_n1641 ), .B(_GFM_n16400 ), .Z(z_out[97]) );
XOR2_X2 _GFM_U2775  ( .A(_GFM_n1643 ), .B(_GFM_n1642 ), .Z(_GFM_n16400 ) );
XOR2_X2 _GFM_U2774  ( .A(_GFM_n1645 ), .B(_GFM_n16440 ), .Z(_GFM_n1641 ) );
XOR2_X2 _GFM_U2773  ( .A(_GFM_n16470 ), .B(_GFM_n16460 ), .Z(_GFM_n1642 ) );
XOR2_X2 _GFM_U2772  ( .A(_GFM_n1649 ), .B(_GFM_n1648 ), .Z(_GFM_n1643 ) );
XOR2_X2 _GFM_U2771  ( .A(_GFM_n16510 ), .B(_GFM_n16500 ), .Z(_GFM_n16440 ));
XOR2_X2 _GFM_U2770  ( .A(_GFM_n16530 ), .B(_GFM_n1652 ), .Z(_GFM_n1645 ) );
XOR2_X2 _GFM_U2769  ( .A(z_in[97]), .B(_GFM_n16540 ), .Z(_GFM_n16460 ) );
XOR2_X2 _GFM_U2768  ( .A(_GFM_N3034 ), .B(_GFM_N3035 ), .Z(_GFM_n16470 ) );
XOR2_X2 _GFM_U2767  ( .A(_GFM_N3031 ), .B(_GFM_N3032 ), .Z(_GFM_n1648 ) );
XOR2_X2 _GFM_U2766  ( .A(_GFM_N3027 ), .B(_GFM_N3028 ), .Z(_GFM_n1649 ) );
XOR2_X2 _GFM_U2765  ( .A(_GFM_N3023 ), .B(_GFM_N3025 ), .Z(_GFM_n16500 ) );
XOR2_X2 _GFM_U2764  ( .A(_GFM_N3018 ), .B(_GFM_N3022 ), .Z(_GFM_n16510 ) );
XOR2_X2 _GFM_U2763  ( .A(_GFM_N3015 ), .B(_GFM_N3017 ), .Z(_GFM_n1652 ) );
XOR2_X2 _GFM_U2762  ( .A(_GFM_N3011 ), .B(_GFM_N3014 ), .Z(_GFM_n16530 ) );
XOR2_X2 _GFM_U2761  ( .A(_GFM_N3008 ), .B(_GFM_N3010 ), .Z(_GFM_n16540 ) );
XOR2_X2 _GFM_U2760  ( .A(_GFM_n1656 ), .B(_GFM_n1655 ), .Z(z_out[98]) );
XOR2_X2 _GFM_U2759  ( .A(_GFM_n16580 ), .B(_GFM_n1657 ), .Z(_GFM_n1655 ) );
XOR2_X2 _GFM_U2758  ( .A(_GFM_n1660 ), .B(_GFM_n16590 ), .Z(_GFM_n1656 ) );
XOR2_X2 _GFM_U2757  ( .A(_GFM_n1662 ), .B(_GFM_n16610 ), .Z(_GFM_n1657 ) );
XOR2_X2 _GFM_U2756  ( .A(_GFM_n16640 ), .B(_GFM_n16630 ), .Z(_GFM_n16580 ));
XOR2_X2 _GFM_U2755  ( .A(_GFM_n1666 ), .B(_GFM_n1665 ), .Z(_GFM_n16590 ) );
XOR2_X2 _GFM_U2754  ( .A(_GFM_n16680 ), .B(_GFM_n16670 ), .Z(_GFM_n1660 ) );
XOR2_X2 _GFM_U2753  ( .A(z_in[98]), .B(_GFM_n1669 ), .Z(_GFM_n16610 ) );
XOR2_X2 _GFM_U2752  ( .A(_GFM_N3065 ), .B(_GFM_N3066 ), .Z(_GFM_n1662 ) );
XOR2_X2 _GFM_U2751  ( .A(_GFM_N3062 ), .B(_GFM_N3063 ), .Z(_GFM_n16630 ) );
XOR2_X2 _GFM_U2750  ( .A(_GFM_N3058 ), .B(_GFM_N3059 ), .Z(_GFM_n16640 ) );
XOR2_X2 _GFM_U2749  ( .A(_GFM_N3054 ), .B(_GFM_N3056 ), .Z(_GFM_n1665 ) );
XOR2_X2 _GFM_U2748  ( .A(_GFM_N3049 ), .B(_GFM_N3053 ), .Z(_GFM_n1666 ) );
XOR2_X2 _GFM_U2747  ( .A(_GFM_N3046 ), .B(_GFM_N3048 ), .Z(_GFM_n16670 ) );
XOR2_X2 _GFM_U2746  ( .A(_GFM_N3042 ), .B(_GFM_N3045 ), .Z(_GFM_n16680 ) );
XOR2_X2 _GFM_U2745  ( .A(_GFM_N3039 ), .B(_GFM_N3041 ), .Z(_GFM_n1669 ) );
XOR2_X2 _GFM_U2744  ( .A(_GFM_n16710 ), .B(_GFM_n16700 ), .Z(z_out[99]) );
XOR2_X2 _GFM_U2743  ( .A(_GFM_n1673 ), .B(_GFM_n1672 ), .Z(_GFM_n16700 ) );
XOR2_X2 _GFM_U2742  ( .A(_GFM_n16750 ), .B(_GFM_n1674 ), .Z(_GFM_n16710 ) );
XOR2_X2 _GFM_U2741  ( .A(_GFM_n16770 ), .B(_GFM_n1676 ), .Z(_GFM_n1672 ) );
XOR2_X2 _GFM_U2740  ( .A(_GFM_n1679 ), .B(_GFM_n16780 ), .Z(_GFM_n1673 ) );
XOR2_X2 _GFM_U2739  ( .A(_GFM_n16810 ), .B(_GFM_n1680 ), .Z(_GFM_n1674 ) );
XOR2_X2 _GFM_U2738  ( .A(_GFM_n1683 ), .B(_GFM_n16820 ), .Z(_GFM_n16750 ) );
XOR2_X2 _GFM_U2737  ( .A(z_in[99]), .B(_GFM_n16840 ), .Z(_GFM_n1676 ) );
XOR2_X2 _GFM_U2736  ( .A(_GFM_N3096 ), .B(_GFM_N3097 ), .Z(_GFM_n16770 ) );
XOR2_X2 _GFM_U2735  ( .A(_GFM_N3093 ), .B(_GFM_N3094 ), .Z(_GFM_n16780 ) );
XOR2_X2 _GFM_U2734  ( .A(_GFM_N3089 ), .B(_GFM_N3090 ), .Z(_GFM_n1679 ) );
XOR2_X2 _GFM_U2733  ( .A(_GFM_N3085 ), .B(_GFM_N3087 ), .Z(_GFM_n1680 ) );
XOR2_X2 _GFM_U2732  ( .A(_GFM_N3080 ), .B(_GFM_N3084 ), .Z(_GFM_n16810 ) );
XOR2_X2 _GFM_U2731  ( .A(_GFM_N3077 ), .B(_GFM_N3079 ), .Z(_GFM_n16820 ) );
XOR2_X2 _GFM_U2730  ( .A(_GFM_N3073 ), .B(_GFM_N3076 ), .Z(_GFM_n1683 ) );
XOR2_X2 _GFM_U2729  ( .A(_GFM_N3070 ), .B(_GFM_N3072 ), .Z(_GFM_n16840 ) );
XOR2_X2 _GFM_U2728  ( .A(_GFM_n1686 ), .B(_GFM_n16850 ), .Z(z_out[100]) );
XOR2_X2 _GFM_U2727  ( .A(_GFM_n1688 ), .B(_GFM_n1687 ), .Z(_GFM_n16850 ) );
XOR2_X2 _GFM_U2726  ( .A(_GFM_n16900 ), .B(_GFM_n16890 ), .Z(_GFM_n1686 ) );
XOR2_X2 _GFM_U2725  ( .A(_GFM_n16920 ), .B(_GFM_n1691 ), .Z(_GFM_n1687 ) );
XOR2_X2 _GFM_U2724  ( .A(_GFM_n16940 ), .B(_GFM_n1693 ), .Z(_GFM_n1688 ) );
XOR2_X2 _GFM_U2723  ( .A(_GFM_n1696 ), .B(_GFM_n16950 ), .Z(_GFM_n16890 ) );
XOR2_X2 _GFM_U2722  ( .A(_GFM_n16980 ), .B(_GFM_n1697 ), .Z(_GFM_n16900 ) );
XOR2_X2 _GFM_U2721  ( .A(z_in[100]), .B(_GFM_n16990 ), .Z(_GFM_n1691 ) );
XOR2_X2 _GFM_U2720  ( .A(_GFM_N3127 ), .B(_GFM_N3128 ), .Z(_GFM_n16920 ) );
XOR2_X2 _GFM_U2719  ( .A(_GFM_N3124 ), .B(_GFM_N3125 ), .Z(_GFM_n1693 ) );
XOR2_X2 _GFM_U2718  ( .A(_GFM_N3120 ), .B(_GFM_N3121 ), .Z(_GFM_n16940 ) );
XOR2_X2 _GFM_U2717  ( .A(_GFM_N3116 ), .B(_GFM_N3118 ), .Z(_GFM_n16950 ) );
XOR2_X2 _GFM_U2716  ( .A(_GFM_N3111 ), .B(_GFM_N3115 ), .Z(_GFM_n1696 ) );
XOR2_X2 _GFM_U2715  ( .A(_GFM_N3108 ), .B(_GFM_N3110 ), .Z(_GFM_n1697 ) );
XOR2_X2 _GFM_U2714  ( .A(_GFM_N3104 ), .B(_GFM_N3107 ), .Z(_GFM_n16980 ) );
XOR2_X2 _GFM_U2713  ( .A(_GFM_N3101 ), .B(_GFM_N3103 ), .Z(_GFM_n16990 ) );
XOR2_X2 _GFM_U2712  ( .A(_GFM_n17010 ), .B(_GFM_n1700 ), .Z(z_out[101]) );
XOR2_X2 _GFM_U2711  ( .A(_GFM_n1703 ), .B(_GFM_n17020 ), .Z(_GFM_n1700 ) );
XOR2_X2 _GFM_U2710  ( .A(_GFM_n1705 ), .B(_GFM_n1704 ), .Z(_GFM_n17010 ) );
XOR2_X2 _GFM_U2709  ( .A(_GFM_n1707 ), .B(_GFM_n17060 ), .Z(_GFM_n17020 ) );
XOR2_X2 _GFM_U2708  ( .A(_GFM_n17090 ), .B(_GFM_n17080 ), .Z(_GFM_n1703 ) );
XOR2_X2 _GFM_U2707  ( .A(_GFM_n1711 ), .B(_GFM_n1710 ), .Z(_GFM_n1704 ) );
XOR2_X2 _GFM_U2706  ( .A(_GFM_n17130 ), .B(_GFM_n17120 ), .Z(_GFM_n1705 ) );
XOR2_X2 _GFM_U2705  ( .A(z_in[101]), .B(_GFM_n1714 ), .Z(_GFM_n17060 ) );
XOR2_X2 _GFM_U2704  ( .A(_GFM_N3158 ), .B(_GFM_N3159 ), .Z(_GFM_n1707 ) );
XOR2_X2 _GFM_U2703  ( .A(_GFM_N3155 ), .B(_GFM_N3156 ), .Z(_GFM_n17080 ) );
XOR2_X2 _GFM_U2702  ( .A(_GFM_N3151 ), .B(_GFM_N3152 ), .Z(_GFM_n17090 ) );
XOR2_X2 _GFM_U2701  ( .A(_GFM_N3147 ), .B(_GFM_N3149 ), .Z(_GFM_n1710 ) );
XOR2_X2 _GFM_U2700  ( .A(_GFM_N3142 ), .B(_GFM_N3146 ), .Z(_GFM_n1711 ) );
XOR2_X2 _GFM_U2699  ( .A(_GFM_N3139 ), .B(_GFM_N3141 ), .Z(_GFM_n17120 ) );
XOR2_X2 _GFM_U2698  ( .A(_GFM_N3135 ), .B(_GFM_N3138 ), .Z(_GFM_n17130 ) );
XOR2_X2 _GFM_U2697  ( .A(_GFM_N3132 ), .B(_GFM_N3134 ), .Z(_GFM_n1714 ) );
XOR2_X2 _GFM_U2696  ( .A(_GFM_n17160 ), .B(_GFM_n17150 ), .Z(z_out[102]) );
XOR2_X2 _GFM_U2695  ( .A(_GFM_n1718 ), .B(_GFM_n1717 ), .Z(_GFM_n17150 ) );
XOR2_X2 _GFM_U2694  ( .A(_GFM_n17200 ), .B(_GFM_n1719 ), .Z(_GFM_n17160 ) );
XOR2_X2 _GFM_U2693  ( .A(_GFM_n1722 ), .B(_GFM_n17210 ), .Z(_GFM_n1717 ) );
XOR2_X2 _GFM_U2692  ( .A(_GFM_n1724 ), .B(_GFM_n17230 ), .Z(_GFM_n1718 ) );
XOR2_X2 _GFM_U2691  ( .A(_GFM_n17260 ), .B(_GFM_n17250 ), .Z(_GFM_n1719 ) );
XOR2_X2 _GFM_U2690  ( .A(_GFM_n1728 ), .B(_GFM_n1727 ), .Z(_GFM_n17200 ) );
XOR2_X2 _GFM_U2689  ( .A(z_in[102]), .B(_GFM_n17290 ), .Z(_GFM_n17210 ) );
XOR2_X2 _GFM_U2688  ( .A(_GFM_N3189 ), .B(_GFM_N3190 ), .Z(_GFM_n1722 ) );
XOR2_X2 _GFM_U2687  ( .A(_GFM_N3186 ), .B(_GFM_N3187 ), .Z(_GFM_n17230 ) );
XOR2_X2 _GFM_U2686  ( .A(_GFM_N3182 ), .B(_GFM_N3183 ), .Z(_GFM_n1724 ) );
XOR2_X2 _GFM_U2685  ( .A(_GFM_N3178 ), .B(_GFM_N3180 ), .Z(_GFM_n17250 ) );
XOR2_X2 _GFM_U2684  ( .A(_GFM_N3173 ), .B(_GFM_N3177 ), .Z(_GFM_n17260 ) );
XOR2_X2 _GFM_U2683  ( .A(_GFM_N3170 ), .B(_GFM_N3172 ), .Z(_GFM_n1727 ) );
XOR2_X2 _GFM_U2682  ( .A(_GFM_N3166 ), .B(_GFM_N3169 ), .Z(_GFM_n1728 ) );
XOR2_X2 _GFM_U2681  ( .A(_GFM_N3163 ), .B(_GFM_N3165 ), .Z(_GFM_n17290 ) );
XOR2_X2 _GFM_U2680  ( .A(_GFM_n1731 ), .B(_GFM_n17300 ), .Z(z_out[103]) );
XOR2_X2 _GFM_U2679  ( .A(_GFM_n17330 ), .B(_GFM_n17320 ), .Z(_GFM_n17300 ));
XOR2_X2 _GFM_U2678  ( .A(_GFM_n1735 ), .B(_GFM_n1734 ), .Z(_GFM_n1731 ) );
XOR2_X2 _GFM_U2677  ( .A(_GFM_n17370 ), .B(_GFM_n1736 ), .Z(_GFM_n17320 ) );
XOR2_X2 _GFM_U2676  ( .A(_GFM_n17390 ), .B(_GFM_n1738 ), .Z(_GFM_n17330 ) );
XOR2_X2 _GFM_U2675  ( .A(_GFM_n1741 ), .B(_GFM_n17400 ), .Z(_GFM_n1734 ) );
XOR2_X2 _GFM_U2674  ( .A(_GFM_n17430 ), .B(_GFM_n1742 ), .Z(_GFM_n1735 ) );
XOR2_X2 _GFM_U2673  ( .A(z_in[103]), .B(_GFM_n17440 ), .Z(_GFM_n1736 ) );
XOR2_X2 _GFM_U2672  ( .A(_GFM_N3220 ), .B(_GFM_N3221 ), .Z(_GFM_n17370 ) );
XOR2_X2 _GFM_U2671  ( .A(_GFM_N3217 ), .B(_GFM_N3218 ), .Z(_GFM_n1738 ) );
XOR2_X2 _GFM_U2670  ( .A(_GFM_N3213 ), .B(_GFM_N3214 ), .Z(_GFM_n17390 ) );
XOR2_X2 _GFM_U2669  ( .A(_GFM_N3209 ), .B(_GFM_N3211 ), .Z(_GFM_n17400 ) );
XOR2_X2 _GFM_U2668  ( .A(_GFM_N3204 ), .B(_GFM_N3208 ), .Z(_GFM_n1741 ) );
XOR2_X2 _GFM_U2667  ( .A(_GFM_N3201 ), .B(_GFM_N3203 ), .Z(_GFM_n1742 ) );
XOR2_X2 _GFM_U2666  ( .A(_GFM_N3197 ), .B(_GFM_N3200 ), .Z(_GFM_n17430 ) );
XOR2_X2 _GFM_U2665  ( .A(_GFM_N3194 ), .B(_GFM_N3196 ), .Z(_GFM_n17440 ) );
XOR2_X2 _GFM_U2664  ( .A(_GFM_n17460 ), .B(_GFM_n1745 ), .Z(z_out[104]) );
XOR2_X2 _GFM_U2663  ( .A(_GFM_n1748 ), .B(_GFM_n17470 ), .Z(_GFM_n1745 ) );
XOR2_X2 _GFM_U2662  ( .A(_GFM_n1750 ), .B(_GFM_n1749 ), .Z(_GFM_n17460 ) );
XOR2_X2 _GFM_U2661  ( .A(_GFM_n17520 ), .B(_GFM_n17510 ), .Z(_GFM_n17470 ));
XOR2_X2 _GFM_U2660  ( .A(_GFM_n17540 ), .B(_GFM_n1753 ), .Z(_GFM_n1748 ) );
XOR2_X2 _GFM_U2659  ( .A(_GFM_n17560 ), .B(_GFM_n1755 ), .Z(_GFM_n1749 ) );
XOR2_X2 _GFM_U2658  ( .A(_GFM_n1758 ), .B(_GFM_n17570 ), .Z(_GFM_n1750 ) );
XOR2_X2 _GFM_U2657  ( .A(z_in[104]), .B(_GFM_n1759 ), .Z(_GFM_n17510 ) );
XOR2_X2 _GFM_U2656  ( .A(_GFM_N3251 ), .B(_GFM_N3252 ), .Z(_GFM_n17520 ) );
XOR2_X2 _GFM_U2655  ( .A(_GFM_N3248 ), .B(_GFM_N3249 ), .Z(_GFM_n1753 ) );
XOR2_X2 _GFM_U2654  ( .A(_GFM_N3244 ), .B(_GFM_N3245 ), .Z(_GFM_n17540 ) );
XOR2_X2 _GFM_U2653  ( .A(_GFM_N3240 ), .B(_GFM_N3242 ), .Z(_GFM_n1755 ) );
XOR2_X2 _GFM_U2652  ( .A(_GFM_N3235 ), .B(_GFM_N3239 ), .Z(_GFM_n17560 ) );
XOR2_X2 _GFM_U2651  ( .A(_GFM_N3232 ), .B(_GFM_N3234 ), .Z(_GFM_n17570 ) );
XOR2_X2 _GFM_U2650  ( .A(_GFM_N3228 ), .B(_GFM_N3231 ), .Z(_GFM_n1758 ) );
XOR2_X2 _GFM_U2649  ( .A(_GFM_N3225 ), .B(_GFM_N3227 ), .Z(_GFM_n1759 ) );
XOR2_X2 _GFM_U2648  ( .A(_GFM_n17610 ), .B(_GFM_n17600 ), .Z(z_out[105]) );
XOR2_X2 _GFM_U2647  ( .A(_GFM_n17630 ), .B(_GFM_n1762 ), .Z(_GFM_n17600 ) );
XOR2_X2 _GFM_U2646  ( .A(_GFM_n1765 ), .B(_GFM_n17640 ), .Z(_GFM_n17610 ) );
XOR2_X2 _GFM_U2645  ( .A(_GFM_n1767 ), .B(_GFM_n1766 ), .Z(_GFM_n1762 ) );
XOR2_X2 _GFM_U2644  ( .A(_GFM_n1769 ), .B(_GFM_n17680 ), .Z(_GFM_n17630 ) );
XOR2_X2 _GFM_U2643  ( .A(_GFM_n17710 ), .B(_GFM_n17700 ), .Z(_GFM_n17640 ));
XOR2_X2 _GFM_U2642  ( .A(_GFM_n1773 ), .B(_GFM_n1772 ), .Z(_GFM_n1765 ) );
XOR2_X2 _GFM_U2641  ( .A(z_in[105]), .B(_GFM_n17740 ), .Z(_GFM_n1766 ) );
XOR2_X2 _GFM_U2640  ( .A(_GFM_N3282 ), .B(_GFM_N3283 ), .Z(_GFM_n1767 ) );
XOR2_X2 _GFM_U2639  ( .A(_GFM_N3279 ), .B(_GFM_N3280 ), .Z(_GFM_n17680 ) );
XOR2_X2 _GFM_U2638  ( .A(_GFM_N3275 ), .B(_GFM_N3276 ), .Z(_GFM_n1769 ) );
XOR2_X2 _GFM_U2637  ( .A(_GFM_N3271 ), .B(_GFM_N3273 ), .Z(_GFM_n17700 ) );
XOR2_X2 _GFM_U2636  ( .A(_GFM_N3266 ), .B(_GFM_N3270 ), .Z(_GFM_n17710 ) );
XOR2_X2 _GFM_U2635  ( .A(_GFM_N3263 ), .B(_GFM_N3265 ), .Z(_GFM_n1772 ) );
XOR2_X2 _GFM_U2634  ( .A(_GFM_N3259 ), .B(_GFM_N3262 ), .Z(_GFM_n1773 ) );
XOR2_X2 _GFM_U2633  ( .A(_GFM_N3256 ), .B(_GFM_N3258 ), .Z(_GFM_n17740 ) );
XOR2_X2 _GFM_U2632  ( .A(_GFM_n1776 ), .B(_GFM_n17750 ), .Z(z_out[106]) );
XOR2_X2 _GFM_U2631  ( .A(_GFM_n17780 ), .B(_GFM_n17770 ), .Z(_GFM_n17750 ));
XOR2_X2 _GFM_U2630  ( .A(_GFM_n1780 ), .B(_GFM_n1779 ), .Z(_GFM_n1776 ) );
XOR2_X2 _GFM_U2629  ( .A(_GFM_n17820 ), .B(_GFM_n1781 ), .Z(_GFM_n17770 ) );
XOR2_X2 _GFM_U2628  ( .A(_GFM_n1784 ), .B(_GFM_n17830 ), .Z(_GFM_n17780 ) );
XOR2_X2 _GFM_U2627  ( .A(_GFM_n1786 ), .B(_GFM_n17850 ), .Z(_GFM_n1779 ) );
XOR2_X2 _GFM_U2626  ( .A(_GFM_n17880 ), .B(_GFM_n17870 ), .Z(_GFM_n1780 ) );
XOR2_X2 _GFM_U2625  ( .A(z_in[106]), .B(_GFM_n1789 ), .Z(_GFM_n1781 ) );
XOR2_X2 _GFM_U2624  ( .A(_GFM_N3313 ), .B(_GFM_N3316 ), .Z(_GFM_n17820 ) );
XOR2_X2 _GFM_U2623  ( .A(_GFM_N3309 ), .B(_GFM_N3312 ), .Z(_GFM_n17830 ) );
XOR2_X2 _GFM_U2622  ( .A(_GFM_N3306 ), .B(_GFM_N3308 ), .Z(_GFM_n1784 ) );
XOR2_X2 _GFM_U2621  ( .A(_GFM_N3303 ), .B(_GFM_N3304 ), .Z(_GFM_n17850 ) );
XOR2_X2 _GFM_U2620  ( .A(_GFM_N3298 ), .B(_GFM_N3299 ), .Z(_GFM_n1786 ) );
XOR2_X2 _GFM_U2619  ( .A(_GFM_N3294 ), .B(_GFM_N3296 ), .Z(_GFM_n17870 ) );
XOR2_X2 _GFM_U2618  ( .A(_GFM_N3290 ), .B(_GFM_N3293 ), .Z(_GFM_n17880 ) );
XOR2_X2 _GFM_U2617  ( .A(_GFM_N3287 ), .B(_GFM_N3289 ), .Z(_GFM_n1789 ) );
XOR2_X2 _GFM_U2616  ( .A(_GFM_n17910 ), .B(_GFM_n1790 ), .Z(z_out[107]) );
XOR2_X2 _GFM_U2615  ( .A(_GFM_n1793 ), .B(_GFM_n17920 ), .Z(_GFM_n1790 ) );
XOR2_X2 _GFM_U2614  ( .A(_GFM_n17950 ), .B(_GFM_n17940 ), .Z(_GFM_n17910 ));
XOR2_X2 _GFM_U2613  ( .A(_GFM_n1797 ), .B(_GFM_n1796 ), .Z(_GFM_n17920 ) );
XOR2_X2 _GFM_U2612  ( .A(_GFM_n17990 ), .B(_GFM_n1798 ), .Z(_GFM_n1793 ) );
XOR2_X2 _GFM_U2611  ( .A(_GFM_n18010 ), .B(_GFM_n1800 ), .Z(_GFM_n17940 ) );
XOR2_X2 _GFM_U2610  ( .A(_GFM_n1803 ), .B(_GFM_n18020 ), .Z(_GFM_n17950 ) );
XOR2_X2 _GFM_U2609  ( .A(z_in[107]), .B(_GFM_n1804 ), .Z(_GFM_n1796 ) );
XOR2_X2 _GFM_U2608  ( .A(_GFM_N3346 ), .B(_GFM_N3349 ), .Z(_GFM_n1797 ) );
XOR2_X2 _GFM_U2607  ( .A(_GFM_N3341 ), .B(_GFM_N3345 ), .Z(_GFM_n1798 ) );
XOR2_X2 _GFM_U2606  ( .A(_GFM_N3338 ), .B(_GFM_N3340 ), .Z(_GFM_n17990 ) );
XOR2_X2 _GFM_U2605  ( .A(_GFM_N3335 ), .B(_GFM_N3336 ), .Z(_GFM_n1800 ) );
XOR2_X2 _GFM_U2604  ( .A(_GFM_N3330 ), .B(_GFM_N3331 ), .Z(_GFM_n18010 ) );
XOR2_X2 _GFM_U2603  ( .A(_GFM_N3326 ), .B(_GFM_N3328 ), .Z(_GFM_n18020 ) );
XOR2_X2 _GFM_U2602  ( .A(_GFM_N3322 ), .B(_GFM_N3325 ), .Z(_GFM_n1803 ) );
XOR2_X2 _GFM_U2601  ( .A(_GFM_N3319 ), .B(_GFM_N3321 ), .Z(_GFM_n1804 ) );
XOR2_X2 _GFM_U2600  ( .A(_GFM_n18060 ), .B(_GFM_n18050 ), .Z(z_out[108]) );
XOR2_X2 _GFM_U2599  ( .A(_GFM_n18080 ), .B(_GFM_n1807 ), .Z(_GFM_n18050 ) );
XOR2_X2 _GFM_U2598  ( .A(_GFM_n1810 ), .B(_GFM_n18090 ), .Z(_GFM_n18060 ) );
XOR2_X2 _GFM_U2597  ( .A(_GFM_n1812 ), .B(_GFM_n1811 ), .Z(_GFM_n1807 ) );
XOR2_X2 _GFM_U2596  ( .A(_GFM_n18140 ), .B(_GFM_n18130 ), .Z(_GFM_n18080 ));
XOR2_X2 _GFM_U2595  ( .A(_GFM_n18160 ), .B(_GFM_n1815 ), .Z(_GFM_n18090 ) );
XOR2_X2 _GFM_U2594  ( .A(_GFM_n18180 ), .B(_GFM_n1817 ), .Z(_GFM_n1810 ) );
XOR2_X2 _GFM_U2593  ( .A(z_in[108]), .B(_GFM_n18190 ), .Z(_GFM_n1811 ) );
XOR2_X2 _GFM_U2592  ( .A(_GFM_N3380 ), .B(_GFM_N3383 ), .Z(_GFM_n1812 ) );
XOR2_X2 _GFM_U2591  ( .A(_GFM_N3374 ), .B(_GFM_N3378 ), .Z(_GFM_n18130 ) );
XOR2_X2 _GFM_U2590  ( .A(_GFM_N3371 ), .B(_GFM_N3373 ), .Z(_GFM_n18140 ) );
XOR2_X2 _GFM_U2589  ( .A(_GFM_N3368 ), .B(_GFM_N3369 ), .Z(_GFM_n1815 ) );
XOR2_X2 _GFM_U2588  ( .A(_GFM_N3363 ), .B(_GFM_N3364 ), .Z(_GFM_n18160 ) );
XOR2_X2 _GFM_U2587  ( .A(_GFM_N3359 ), .B(_GFM_N3361 ), .Z(_GFM_n1817 ) );
XOR2_X2 _GFM_U2586  ( .A(_GFM_N3355 ), .B(_GFM_N3358 ), .Z(_GFM_n18180 ) );
XOR2_X2 _GFM_U2585  ( .A(_GFM_N3352 ), .B(_GFM_N3354 ), .Z(_GFM_n18190 ) );
XOR2_X2 _GFM_U2584  ( .A(_GFM_n1821 ), .B(_GFM_n1820 ), .Z(z_out[109]) );
XOR2_X2 _GFM_U2583  ( .A(_GFM_n18230 ), .B(_GFM_n18220 ), .Z(_GFM_n1820 ) );
XOR2_X2 _GFM_U2582  ( .A(_GFM_n18250 ), .B(_GFM_n1824 ), .Z(_GFM_n1821 ) );
XOR2_X2 _GFM_U2581  ( .A(_GFM_n1827 ), .B(_GFM_n18260 ), .Z(_GFM_n18220 ) );
XOR2_X2 _GFM_U2580  ( .A(_GFM_n1829 ), .B(_GFM_n1828 ), .Z(_GFM_n18230 ) );
XOR2_X2 _GFM_U2579  ( .A(_GFM_n1831 ), .B(_GFM_n18300 ), .Z(_GFM_n1824 ) );
XOR2_X2 _GFM_U2578  ( .A(_GFM_n18330 ), .B(_GFM_n18320 ), .Z(_GFM_n18250 ));
XOR2_X2 _GFM_U2577  ( .A(z_in[109]), .B(_GFM_n1834 ), .Z(_GFM_n18260 ) );
XOR2_X2 _GFM_U2576  ( .A(_GFM_N3415 ), .B(_GFM_N3418 ), .Z(_GFM_n1827 ) );
XOR2_X2 _GFM_U2575  ( .A(_GFM_N3409 ), .B(_GFM_N3413 ), .Z(_GFM_n1828 ) );
XOR2_X2 _GFM_U2574  ( .A(_GFM_N3406 ), .B(_GFM_N3407 ), .Z(_GFM_n1829 ) );
XOR2_X2 _GFM_U2573  ( .A(_GFM_N3402 ), .B(_GFM_N3404 ), .Z(_GFM_n18300 ) );
XOR2_X2 _GFM_U2572  ( .A(_GFM_N3397 ), .B(_GFM_N3398 ), .Z(_GFM_n1831 ) );
XOR2_X2 _GFM_U2571  ( .A(_GFM_N3393 ), .B(_GFM_N3395 ), .Z(_GFM_n18320 ) );
XOR2_X2 _GFM_U2570  ( .A(_GFM_N3389 ), .B(_GFM_N3392 ), .Z(_GFM_n18330 ) );
XOR2_X2 _GFM_U2569  ( .A(_GFM_N3386 ), .B(_GFM_N3388 ), .Z(_GFM_n1834 ) );
XOR2_X2 _GFM_U2568  ( .A(_GFM_n18360 ), .B(_GFM_n1835 ), .Z(z_out[110]) );
XOR2_X2 _GFM_U2567  ( .A(_GFM_n1838 ), .B(_GFM_n18370 ), .Z(_GFM_n1835 ) );
XOR2_X2 _GFM_U2566  ( .A(_GFM_n18400 ), .B(_GFM_n18390 ), .Z(_GFM_n18360 ));
XOR2_X2 _GFM_U2565  ( .A(_GFM_n1842 ), .B(_GFM_n1841 ), .Z(_GFM_n18370 ) );
XOR2_X2 _GFM_U2564  ( .A(_GFM_n18440 ), .B(_GFM_n1843 ), .Z(_GFM_n1838 ) );
XOR2_X2 _GFM_U2563  ( .A(_GFM_n1846 ), .B(_GFM_n18450 ), .Z(_GFM_n18390 ) );
XOR2_X2 _GFM_U2562  ( .A(_GFM_n1848 ), .B(_GFM_n18470 ), .Z(_GFM_n18400 ) );
XOR2_X2 _GFM_U2561  ( .A(z_in[110]), .B(_GFM_n18490 ), .Z(_GFM_n1841 ) );
XOR2_X2 _GFM_U2560  ( .A(_GFM_N3452 ), .B(_GFM_N3455 ), .Z(_GFM_n1842 ) );
XOR2_X2 _GFM_U2559  ( .A(_GFM_N3446 ), .B(_GFM_N3450 ), .Z(_GFM_n1843 ) );
XOR2_X2 _GFM_U2558  ( .A(_GFM_N3443 ), .B(_GFM_N3444 ), .Z(_GFM_n18440 ) );
XOR2_X2 _GFM_U2557  ( .A(_GFM_N3439 ), .B(_GFM_N3441 ), .Z(_GFM_n18450 ) );
XOR2_X2 _GFM_U2556  ( .A(_GFM_N3433 ), .B(_GFM_N3434 ), .Z(_GFM_n1846 ) );
XOR2_X2 _GFM_U2555  ( .A(_GFM_N3429 ), .B(_GFM_N3431 ), .Z(_GFM_n18470 ) );
XOR2_X2 _GFM_U2554  ( .A(_GFM_N3425 ), .B(_GFM_N3428 ), .Z(_GFM_n1848 ) );
XOR2_X2 _GFM_U2553  ( .A(_GFM_N3422 ), .B(_GFM_N3424 ), .Z(_GFM_n18490 ) );
XOR2_X2 _GFM_U2552  ( .A(_GFM_n1851 ), .B(_GFM_n18500 ), .Z(z_out[111]) );
XOR2_X2 _GFM_U2551  ( .A(_GFM_n18530 ), .B(_GFM_n1852 ), .Z(_GFM_n18500 ) );
XOR2_X2 _GFM_U2550  ( .A(_GFM_n1855 ), .B(_GFM_n18540 ), .Z(_GFM_n1851 ) );
XOR2_X2 _GFM_U2549  ( .A(_GFM_n18570 ), .B(_GFM_n18560 ), .Z(_GFM_n1852 ) );
XOR2_X2 _GFM_U2548  ( .A(_GFM_n1859 ), .B(_GFM_n1858 ), .Z(_GFM_n18530 ) );
XOR2_X2 _GFM_U2547  ( .A(_GFM_n18610 ), .B(_GFM_n1860 ), .Z(_GFM_n18540 ) );
XOR2_X2 _GFM_U2546  ( .A(_GFM_n18630 ), .B(_GFM_n1862 ), .Z(_GFM_n1855 ) );
XOR2_X2 _GFM_U2545  ( .A(z_in[111]), .B(_GFM_n18640 ), .Z(_GFM_n18560 ) );
XOR2_X2 _GFM_U2544  ( .A(_GFM_N3491 ), .B(_GFM_N3495 ), .Z(_GFM_n18570 ) );
XOR2_X2 _GFM_U2543  ( .A(_GFM_N3484 ), .B(_GFM_N3489 ), .Z(_GFM_n1858 ) );
XOR2_X2 _GFM_U2542  ( .A(_GFM_N3482 ), .B(_GFM_N3483 ), .Z(_GFM_n1859 ) );
XOR2_X2 _GFM_U2541  ( .A(_GFM_N3477 ), .B(_GFM_N3479 ), .Z(_GFM_n1860 ) );
XOR2_X2 _GFM_U2540  ( .A(_GFM_N3471 ), .B(_GFM_N3472 ), .Z(_GFM_n18610 ) );
XOR2_X2 _GFM_U2539  ( .A(_GFM_N3467 ), .B(_GFM_N3469 ), .Z(_GFM_n1862 ) );
XOR2_X2 _GFM_U2538  ( .A(_GFM_N3463 ), .B(_GFM_N3466 ), .Z(_GFM_n18630 ) );
XOR2_X2 _GFM_U2537  ( .A(_GFM_N3460 ), .B(_GFM_N3462 ), .Z(_GFM_n18640 ) );
XOR2_X2 _GFM_U2536  ( .A(_GFM_n1866 ), .B(_GFM_n1865 ), .Z(z_out[112]) );
XOR2_X2 _GFM_U2535  ( .A(_GFM_n18680 ), .B(_GFM_n18670 ), .Z(_GFM_n1865 ) );
XOR2_X2 _GFM_U2534  ( .A(_GFM_n18700 ), .B(_GFM_n1869 ), .Z(_GFM_n1866 ) );
XOR2_X2 _GFM_U2533  ( .A(_GFM_n18721 ), .B(_GFM_n18710 ), .Z(_GFM_n18670 ));
XOR2_X2 _GFM_U2532  ( .A(_GFM_n1874 ), .B(_GFM_n1873 ), .Z(_GFM_n18680 ) );
XOR2_X2 _GFM_U2531  ( .A(_GFM_n18760 ), .B(_GFM_n18750 ), .Z(_GFM_n1869 ) );
XOR2_X2 _GFM_U2530  ( .A(_GFM_n18780 ), .B(_GFM_n1877 ), .Z(_GFM_n18700 ) );
XOR2_X2 _GFM_U2529  ( .A(z_in[112]), .B(_GFM_n1879 ), .Z(_GFM_n18710 ) );
XOR2_X2 _GFM_U2528  ( .A(_GFM_N3534 ), .B(_GFM_N3538 ), .Z(_GFM_n18721 ) );
XOR2_X2 _GFM_U2527  ( .A(_GFM_N3527 ), .B(_GFM_N3529 ), .Z(_GFM_n1873 ) );
XOR2_X2 _GFM_U2526  ( .A(_GFM_N3521 ), .B(_GFM_N3524 ), .Z(_GFM_n1874 ) );
XOR2_X2 _GFM_U2525  ( .A(_GFM_N3514 ), .B(_GFM_N3519 ), .Z(_GFM_n18750 ) );
XOR2_X2 _GFM_U2524  ( .A(_GFM_N3511 ), .B(_GFM_N3513 ), .Z(_GFM_n18760 ) );
XOR2_X2 _GFM_U2523  ( .A(_GFM_N3508 ), .B(_GFM_N3509 ), .Z(_GFM_n1877 ) );
XOR2_X2 _GFM_U2522  ( .A(_GFM_N3503 ), .B(_GFM_N3505 ), .Z(_GFM_n18780 ) );
XOR2_X2 _GFM_U2521  ( .A(_GFM_N3500 ), .B(_GFM_N3502 ), .Z(_GFM_n1879 ) );
XOR2_X2 _GFM_U2520  ( .A(_GFM_n18810 ), .B(_GFM_n18800 ), .Z(z_out[113]) );
XOR2_X2 _GFM_U2519  ( .A(_GFM_n1883 ), .B(_GFM_n1882 ), .Z(_GFM_n18800 ) );
XOR2_X2 _GFM_U2518  ( .A(_GFM_n18850 ), .B(_GFM_n18840 ), .Z(_GFM_n18810 ));
XOR2_X2 _GFM_U2517  ( .A(_GFM_n18870 ), .B(_GFM_n1886 ), .Z(_GFM_n1882 ) );
XOR2_X2 _GFM_U2516  ( .A(_GFM_n1889 ), .B(_GFM_n18880 ), .Z(_GFM_n1883 ) );
XOR2_X2 _GFM_U2515  ( .A(_GFM_n1891 ), .B(_GFM_n18901 ), .Z(_GFM_n18840 ) );
XOR2_X2 _GFM_U2514  ( .A(_GFM_n1893 ), .B(_GFM_n18920 ), .Z(_GFM_n18850 ) );
XOR2_X2 _GFM_U2513  ( .A(z_in[113]), .B(_GFM_n18940 ), .Z(_GFM_n1886 ) );
XOR2_X2 _GFM_U2512  ( .A(_GFM_N3580 ), .B(_GFM_N3584 ), .Z(_GFM_n18870 ) );
XOR2_X2 _GFM_U2511  ( .A(_GFM_N3571 ), .B(_GFM_N3574 ), .Z(_GFM_n18880 ) );
XOR2_X2 _GFM_U2510  ( .A(_GFM_N3566 ), .B(_GFM_N3569 ), .Z(_GFM_n1889 ) );
XOR2_X2 _GFM_U2509  ( .A(_GFM_N3558 ), .B(_GFM_N3563 ), .Z(_GFM_n18901 ) );
XOR2_X2 _GFM_U2508  ( .A(_GFM_N3554 ), .B(_GFM_N3556 ), .Z(_GFM_n1891 ) );
XOR2_X2 _GFM_U2507  ( .A(_GFM_N3551 ), .B(_GFM_N3552 ), .Z(_GFM_n18920 ) );
XOR2_X2 _GFM_U2506  ( .A(_GFM_N3546 ), .B(_GFM_N3548 ), .Z(_GFM_n1893 ) );
XOR2_X2 _GFM_U2505  ( .A(_GFM_N3543 ), .B(_GFM_N3545 ), .Z(_GFM_n18940 ) );
XOR2_X2 _GFM_U2504  ( .A(_GFM_n1896 ), .B(_GFM_n18950 ), .Z(z_out[114]) );
XOR2_X2 _GFM_U2503  ( .A(_GFM_n18980 ), .B(_GFM_n1897 ), .Z(_GFM_n18950 ) );
XOR2_X2 _GFM_U2502  ( .A(_GFM_n19001 ), .B(_GFM_n18990 ), .Z(_GFM_n1896 ) );
XOR2_X2 _GFM_U2501  ( .A(_GFM_n19020 ), .B(_GFM_n19010 ), .Z(_GFM_n1897 ) );
XOR2_X2 _GFM_U2500  ( .A(_GFM_n1904 ), .B(_GFM_n1903 ), .Z(_GFM_n18980 ) );
XOR2_X2 _GFM_U2499  ( .A(_GFM_n19060 ), .B(_GFM_n1905 ), .Z(_GFM_n18990 ) );
XOR2_X2 _GFM_U2498  ( .A(_GFM_n1908 ), .B(_GFM_n19070 ), .Z(_GFM_n19001 ) );
XOR2_X2 _GFM_U2497  ( .A(z_in[114]), .B(_GFM_n19090 ), .Z(_GFM_n19010 ) );
XOR2_X2 _GFM_U2496  ( .A(_GFM_N3629 ), .B(_GFM_N3633 ), .Z(_GFM_n19020 ) );
XOR2_X2 _GFM_U2495  ( .A(_GFM_N3620 ), .B(_GFM_N3623 ), .Z(_GFM_n1903 ) );
XOR2_X2 _GFM_U2494  ( .A(_GFM_N3615 ), .B(_GFM_N3618 ), .Z(_GFM_n1904 ) );
XOR2_X2 _GFM_U2493  ( .A(_GFM_N3605 ), .B(_GFM_N3611 ), .Z(_GFM_n1905 ) );
XOR2_X2 _GFM_U2492  ( .A(_GFM_N3600 ), .B(_GFM_N3603 ), .Z(_GFM_n19060 ) );
XOR2_X2 _GFM_U2491  ( .A(_GFM_N3597 ), .B(_GFM_N3598 ), .Z(_GFM_n19070 ) );
XOR2_X2 _GFM_U2490  ( .A(_GFM_N3592 ), .B(_GFM_N3594 ), .Z(_GFM_n1908 ) );
XOR2_X2 _GFM_U2489  ( .A(_GFM_N3589 ), .B(_GFM_N3591 ), .Z(_GFM_n19090 ) );
XOR2_X2 _GFM_U2488  ( .A(_GFM_n19110 ), .B(_GFM_n1910 ), .Z(z_out[115]) );
XOR2_X2 _GFM_U2487  ( .A(_GFM_n1913 ), .B(_GFM_n19120 ), .Z(_GFM_n1910 ) );
XOR2_X2 _GFM_U2486  ( .A(_GFM_n19150 ), .B(_GFM_n1914 ), .Z(_GFM_n19110 ) );
XOR2_X2 _GFM_U2485  ( .A(_GFM_n1917 ), .B(_GFM_n19160 ), .Z(_GFM_n19120 ) );
XOR2_X2 _GFM_U2484  ( .A(_GFM_n19190 ), .B(_GFM_n19180 ), .Z(_GFM_n1913 ) );
XOR2_X2 _GFM_U2483  ( .A(_GFM_n1921 ), .B(_GFM_n1920 ), .Z(_GFM_n1914 ) );
XOR2_X2 _GFM_U2482  ( .A(_GFM_n19230 ), .B(_GFM_n1922 ), .Z(_GFM_n19150 ) );
XOR2_X2 _GFM_U2481  ( .A(z_in[115]), .B(_GFM_n1924 ), .Z(_GFM_n19160 ) );
XOR2_X2 _GFM_U2480  ( .A(_GFM_N3681 ), .B(_GFM_N3685 ), .Z(_GFM_n1917 ) );
XOR2_X2 _GFM_U2479  ( .A(_GFM_N3672 ), .B(_GFM_N3674 ), .Z(_GFM_n19180 ) );
XOR2_X2 _GFM_U2478  ( .A(_GFM_N3666 ), .B(_GFM_N3670 ), .Z(_GFM_n19190 ) );
XOR2_X2 _GFM_U2477  ( .A(_GFM_N3655 ), .B(_GFM_N3662 ), .Z(_GFM_n1920 ) );
XOR2_X2 _GFM_U2476  ( .A(_GFM_N3649 ), .B(_GFM_N3653 ), .Z(_GFM_n1921 ) );
XOR2_X2 _GFM_U2475  ( .A(_GFM_N3647 ), .B(_GFM_N3648 ), .Z(_GFM_n1922 ) );
XOR2_X2 _GFM_U2474  ( .A(_GFM_N3641 ), .B(_GFM_N3643 ), .Z(_GFM_n19230 ) );
XOR2_X2 _GFM_U2473  ( .A(_GFM_N3638 ), .B(_GFM_N3640 ), .Z(_GFM_n1924 ) );
XOR2_X2 _GFM_U2472  ( .A(_GFM_n19260 ), .B(_GFM_n19250 ), .Z(z_out[116]) );
XOR2_X2 _GFM_U2471  ( .A(_GFM_n1928 ), .B(_GFM_n1927 ), .Z(_GFM_n19250 ) );
XOR2_X2 _GFM_U2470  ( .A(_GFM_n19300 ), .B(_GFM_n19290 ), .Z(_GFM_n19260 ));
XOR2_X2 _GFM_U2469  ( .A(_GFM_n19320 ), .B(_GFM_n19311 ), .Z(_GFM_n1927 ) );
XOR2_X2 _GFM_U2468  ( .A(_GFM_n1934 ), .B(_GFM_n19330 ), .Z(_GFM_n1928 ) );
XOR2_X2 _GFM_U2467  ( .A(_GFM_n1936 ), .B(_GFM_n1935 ), .Z(_GFM_n19290 ) );
XOR2_X2 _GFM_U2466  ( .A(_GFM_n19380 ), .B(_GFM_n19370 ), .Z(_GFM_n19300 ));
XOR2_X2 _GFM_U2465  ( .A(z_in[116]), .B(_GFM_n1939 ), .Z(_GFM_n19311 ) );
XOR2_X2 _GFM_U2464  ( .A(_GFM_N3735 ), .B(_GFM_N3740 ), .Z(_GFM_n19320 ) );
XOR2_X2 _GFM_U2463  ( .A(_GFM_N3725 ), .B(_GFM_N3731 ), .Z(_GFM_n19330 ) );
XOR2_X2 _GFM_U2462  ( .A(_GFM_N3719 ), .B(_GFM_N3723 ), .Z(_GFM_n1934 ) );
XOR2_X2 _GFM_U2461  ( .A(_GFM_N3708 ), .B(_GFM_N3715 ), .Z(_GFM_n1935 ) );
XOR2_X2 _GFM_U2460  ( .A(_GFM_N3703 ), .B(_GFM_N3706 ), .Z(_GFM_n1936 ) );
XOR2_X2 _GFM_U2459  ( .A(_GFM_N3699 ), .B(_GFM_N3701 ), .Z(_GFM_n19370 ) );
XOR2_X2 _GFM_U2458  ( .A(_GFM_N3693 ), .B(_GFM_N3695 ), .Z(_GFM_n19380 ) );
XOR2_X2 _GFM_U2457  ( .A(_GFM_N3690 ), .B(_GFM_N3692 ), .Z(_GFM_n1939 ) );
XOR2_X2 _GFM_U2456  ( .A(_GFM_n19411 ), .B(_GFM_n19400 ), .Z(z_out[117]) );
XOR2_X2 _GFM_U2455  ( .A(_GFM_n19430 ), .B(_GFM_n19420 ), .Z(_GFM_n19400 ));
XOR2_X2 _GFM_U2454  ( .A(_GFM_n1945 ), .B(_GFM_n1944 ), .Z(_GFM_n19411 ) );
XOR2_X2 _GFM_U2453  ( .A(_GFM_n19470 ), .B(_GFM_n19460 ), .Z(_GFM_n19420 ));
XOR2_X2 _GFM_U2452  ( .A(_GFM_n19490 ), .B(_GFM_n1948 ), .Z(_GFM_n19430 ) );
XOR2_X2 _GFM_U2451  ( .A(_GFM_n1951 ), .B(_GFM_n19500 ), .Z(_GFM_n1944 ) );
XOR2_X2 _GFM_U2450  ( .A(_GFM_n1953 ), .B(_GFM_n1952 ), .Z(_GFM_n1945 ) );
XOR2_X2 _GFM_U2449  ( .A(z_in[117]), .B(_GFM_n19540 ), .Z(_GFM_n19460 ) );
XOR2_X2 _GFM_U2448  ( .A(_GFM_N3793 ), .B(_GFM_N3798 ), .Z(_GFM_n19470 ) );
XOR2_X2 _GFM_U2447  ( .A(_GFM_N3783 ), .B(_GFM_N3789 ), .Z(_GFM_n1948 ) );
XOR2_X2 _GFM_U2446  ( .A(_GFM_N3775 ), .B(_GFM_N3780 ), .Z(_GFM_n19490 ) );
XOR2_X2 _GFM_U2445  ( .A(_GFM_N3764 ), .B(_GFM_N3771 ), .Z(_GFM_n19500 ) );
XOR2_X2 _GFM_U2444  ( .A(_GFM_N3759 ), .B(_GFM_N3762 ), .Z(_GFM_n1951 ) );
XOR2_X2 _GFM_U2443  ( .A(_GFM_N3754 ), .B(_GFM_N3756 ), .Z(_GFM_n1952 ) );
XOR2_X2 _GFM_U2442  ( .A(_GFM_N3748 ), .B(_GFM_N3750 ), .Z(_GFM_n1953 ) );
XOR2_X2 _GFM_U2441  ( .A(_GFM_N3745 ), .B(_GFM_N3747 ), .Z(_GFM_n19540 ) );
XOR2_X2 _GFM_U2440  ( .A(_GFM_n19560 ), .B(_GFM_n1955 ), .Z(z_out[118]) );
XOR2_X2 _GFM_U2439  ( .A(_GFM_n1958 ), .B(_GFM_n19570 ), .Z(_GFM_n1955 ) );
XOR2_X2 _GFM_U2438  ( .A(_GFM_n19600 ), .B(_GFM_n1959 ), .Z(_GFM_n19560 ) );
XOR2_X2 _GFM_U2437  ( .A(_GFM_n19621 ), .B(_GFM_n19610 ), .Z(_GFM_n19570 ));
XOR2_X2 _GFM_U2436  ( .A(_GFM_n19640 ), .B(_GFM_n19630 ), .Z(_GFM_n1958 ) );
XOR2_X2 _GFM_U2435  ( .A(_GFM_n1966 ), .B(_GFM_n1965 ), .Z(_GFM_n1959 ) );
XOR2_X2 _GFM_U2434  ( .A(_GFM_n19680 ), .B(_GFM_n1967 ), .Z(_GFM_n19600 ) );
XOR2_X2 _GFM_U2433  ( .A(z_in[118]), .B(_GFM_n19690 ), .Z(_GFM_n19610 ) );
XOR2_X2 _GFM_U2432  ( .A(_GFM_N3854 ), .B(_GFM_N3859 ), .Z(_GFM_n19621 ) );
XOR2_X2 _GFM_U2431  ( .A(_GFM_N3844 ), .B(_GFM_N3850 ), .Z(_GFM_n19630 ) );
XOR2_X2 _GFM_U2430  ( .A(_GFM_N3835 ), .B(_GFM_N3840 ), .Z(_GFM_n19640 ) );
XOR2_X2 _GFM_U2429  ( .A(_GFM_N3825 ), .B(_GFM_N3831 ), .Z(_GFM_n1965 ) );
XOR2_X2 _GFM_U2428  ( .A(_GFM_N3818 ), .B(_GFM_N3821 ), .Z(_GFM_n1966 ) );
XOR2_X2 _GFM_U2427  ( .A(_GFM_N3812 ), .B(_GFM_N3816 ), .Z(_GFM_n1967 ) );
XOR2_X2 _GFM_U2426  ( .A(_GFM_N3808 ), .B(_GFM_N3809 ), .Z(_GFM_n19680 ) );
XOR2_X2 _GFM_U2425  ( .A(_GFM_N3803 ), .B(_GFM_N3804 ), .Z(_GFM_n19690 ) );
XOR2_X2 _GFM_U2424  ( .A(_GFM_n19710 ), .B(_GFM_n19701 ), .Z(z_out[119]) );
XOR2_X2 _GFM_U2423  ( .A(_GFM_n19730 ), .B(_GFM_n1972 ), .Z(_GFM_n19701 ) );
XOR2_X2 _GFM_U2422  ( .A(_GFM_n1975 ), .B(_GFM_n19740 ), .Z(_GFM_n19710 ) );
XOR2_X2 _GFM_U2421  ( .A(_GFM_n19770 ), .B(_GFM_n1976 ), .Z(_GFM_n1972 ) );
XOR2_X2 _GFM_U2420  ( .A(_GFM_n1979 ), .B(_GFM_n19780 ), .Z(_GFM_n19730 ) );
XOR2_X2 _GFM_U2419  ( .A(_GFM_n19810 ), .B(_GFM_n19800 ), .Z(_GFM_n19740 ));
XOR2_X2 _GFM_U2418  ( .A(_GFM_n1983 ), .B(_GFM_n1982 ), .Z(_GFM_n1975 ) );
XOR2_X2 _GFM_U2417  ( .A(z_in[119]), .B(_GFM_n1984 ), .Z(_GFM_n1976 ) );
XOR2_X2 _GFM_U2416  ( .A(_GFM_N3918 ), .B(_GFM_N3923 ), .Z(_GFM_n19770 ) );
XOR2_X2 _GFM_U2415  ( .A(_GFM_N3908 ), .B(_GFM_N3914 ), .Z(_GFM_n19780 ) );
XOR2_X2 _GFM_U2414  ( .A(_GFM_N3899 ), .B(_GFM_N3904 ), .Z(_GFM_n1979 ) );
XOR2_X2 _GFM_U2413  ( .A(_GFM_N3889 ), .B(_GFM_N3895 ), .Z(_GFM_n19800 ) );
XOR2_X2 _GFM_U2412  ( .A(_GFM_N3881 ), .B(_GFM_N3883 ), .Z(_GFM_n19810 ) );
XOR2_X2 _GFM_U2411  ( .A(_GFM_N3874 ), .B(_GFM_N3879 ), .Z(_GFM_n1982 ) );
XOR2_X2 _GFM_U2410  ( .A(_GFM_N3869 ), .B(_GFM_N3871 ), .Z(_GFM_n1983 ) );
XOR2_X2 _GFM_U2409  ( .A(_GFM_N3864 ), .B(_GFM_N3865 ), .Z(_GFM_n1984 ) );
XOR2_X2 _GFM_U2408  ( .A(_GFM_n1986 ), .B(_GFM_n19850 ), .Z(z_out[120]) );
XOR2_X2 _GFM_U2407  ( .A(_GFM_n19880 ), .B(_GFM_n19870 ), .Z(_GFM_n19850 ));
XOR2_X2 _GFM_U2406  ( .A(_GFM_n1990 ), .B(_GFM_n1989 ), .Z(_GFM_n1986 ) );
XOR2_X2 _GFM_U2405  ( .A(_GFM_n19920 ), .B(_GFM_n19910 ), .Z(_GFM_n19870 ));
XOR2_X2 _GFM_U2404  ( .A(_GFM_n19940 ), .B(_GFM_n1993 ), .Z(_GFM_n19880 ) );
XOR2_X2 _GFM_U2403  ( .A(_GFM_n1996 ), .B(_GFM_n19950 ), .Z(_GFM_n1989 ) );
XOR2_X2 _GFM_U2402  ( .A(_GFM_n1998 ), .B(_GFM_n1997 ), .Z(_GFM_n1990 ) );
XOR2_X2 _GFM_U2401  ( .A(z_in[120]), .B(_GFM_n19990 ), .Z(_GFM_n19910 ) );
XOR2_X2 _GFM_U2400  ( .A(_GFM_N3985 ), .B(_GFM_N3990 ), .Z(_GFM_n19920 ) );
XOR2_X2 _GFM_U2399  ( .A(_GFM_N3975 ), .B(_GFM_N3981 ), .Z(_GFM_n1993 ) );
XOR2_X2 _GFM_U2398  ( .A(_GFM_N3966 ), .B(_GFM_N3971 ), .Z(_GFM_n19940 ) );
XOR2_X2 _GFM_U2397  ( .A(_GFM_N3955 ), .B(_GFM_N3962 ), .Z(_GFM_n19950 ) );
XOR2_X2 _GFM_U2396  ( .A(_GFM_N3946 ), .B(_GFM_N3951 ), .Z(_GFM_n1996 ) );
XOR2_X2 _GFM_U2395  ( .A(_GFM_N3939 ), .B(_GFM_N3944 ), .Z(_GFM_n1997 ) );
XOR2_X2 _GFM_U2394  ( .A(_GFM_N3934 ), .B(_GFM_N3936 ), .Z(_GFM_n1998 ) );
XOR2_X2 _GFM_U2393  ( .A(_GFM_N3928 ), .B(_GFM_N3931 ), .Z(_GFM_n19990 ) );
XOR2_X2 _GFM_U2392  ( .A(_GFM_n2001 ), .B(_GFM_n20000 ), .Z(z_out[121]) );
XOR2_X2 _GFM_U2391  ( .A(_GFM_n2003 ), .B(_GFM_n20020 ), .Z(_GFM_n20000 ) );
XOR2_X2 _GFM_U2390  ( .A(_GFM_n20050 ), .B(_GFM_n20040 ), .Z(_GFM_n2001 ) );
XOR2_X2 _GFM_U2389  ( .A(_GFM_n2007 ), .B(_GFM_n2006 ), .Z(_GFM_n20020 ) );
XOR2_X2 _GFM_U2388  ( .A(_GFM_n20090 ), .B(_GFM_n20080 ), .Z(_GFM_n2003 ) );
XOR2_X2 _GFM_U2387  ( .A(_GFM_n20110 ), .B(_GFM_n20101 ), .Z(_GFM_n20040 ));
XOR2_X2 _GFM_U2386  ( .A(_GFM_n2013 ), .B(_GFM_n20120 ), .Z(_GFM_n20050 ) );
XOR2_X2 _GFM_U2385  ( .A(z_in[121]), .B(_GFM_n2014 ), .Z(_GFM_n2006 ) );
XOR2_X2 _GFM_U2384  ( .A(_GFM_N4039 ), .B(_GFM_N4042 ), .Z(_GFM_n2007 ) );
XOR2_X2 _GFM_U2383  ( .A(_GFM_N4032 ), .B(_GFM_N4035 ), .Z(_GFM_n20080 ) );
XOR2_X2 _GFM_U2382  ( .A(_GFM_N4024 ), .B(_GFM_N4027 ), .Z(_GFM_n20090 ) );
XOR2_X2 _GFM_U2381  ( .A(_GFM_N4017 ), .B(_GFM_N4020 ), .Z(_GFM_n20101 ) );
XOR2_X2 _GFM_U2380  ( .A(_GFM_N4007 ), .B(_GFM_N4012 ), .Z(_GFM_n20110 ) );
XOR2_X2 _GFM_U2379  ( .A(_GFM_N4004 ), .B(_GFM_N4006 ), .Z(_GFM_n20120 ) );
XOR2_X2 _GFM_U2378  ( .A(_GFM_N3997 ), .B(_GFM_N3999 ), .Z(_GFM_n2013 ) );
XOR2_X2 _GFM_U2377  ( .A(_GFM_N3994 ), .B(_GFM_N3996 ), .Z(_GFM_n2014 ) );
XOR2_X2 _GFM_U2376  ( .A(_GFM_n20160 ), .B(_GFM_n2015 ), .Z(z_out[122]) );
XOR2_X2 _GFM_U2375  ( .A(_GFM_n20180 ), .B(_GFM_n2017 ), .Z(_GFM_n2015 ) );
XOR2_X2 _GFM_U2374  ( .A(_GFM_n20201 ), .B(_GFM_n20190 ), .Z(_GFM_n20160 ));
XOR2_X2 _GFM_U2373  ( .A(_GFM_n20220 ), .B(_GFM_n2021 ), .Z(_GFM_n2017 ) );
XOR2_X2 _GFM_U2372  ( .A(_GFM_n2024 ), .B(_GFM_n20230 ), .Z(_GFM_n20180 ) );
XOR2_X2 _GFM_U2371  ( .A(_GFM_n20260 ), .B(_GFM_n20250 ), .Z(_GFM_n20190 ));
XOR2_X2 _GFM_U2370  ( .A(_GFM_n2028 ), .B(_GFM_n2027 ), .Z(_GFM_n20201 ) );
XOR2_X2 _GFM_U2369  ( .A(z_in[122]), .B(_GFM_n2029 ), .Z(_GFM_n2021 ) );
XOR2_X2 _GFM_U2368  ( .A(_GFM_N4094 ), .B(_GFM_N4097 ), .Z(_GFM_n20220 ) );
XOR2_X2 _GFM_U2367  ( .A(_GFM_N4087 ), .B(_GFM_N4090 ), .Z(_GFM_n20230 ) );
XOR2_X2 _GFM_U2366  ( .A(_GFM_N4079 ), .B(_GFM_N4082 ), .Z(_GFM_n2024 ) );
XOR2_X2 _GFM_U2365  ( .A(_GFM_N4072 ), .B(_GFM_N4075 ), .Z(_GFM_n20250 ) );
XOR2_X2 _GFM_U2364  ( .A(_GFM_N4063 ), .B(_GFM_N4066 ), .Z(_GFM_n20260 ) );
XOR2_X2 _GFM_U2363  ( .A(_GFM_N4057 ), .B(_GFM_N4059 ), .Z(_GFM_n2027 ) );
XOR2_X2 _GFM_U2362  ( .A(_GFM_N4050 ), .B(_GFM_N4052 ), .Z(_GFM_n2028 ) );
XOR2_X2 _GFM_U2361  ( .A(_GFM_N4047 ), .B(_GFM_N4049 ), .Z(_GFM_n2029 ) );
XOR2_X2 _GFM_U2360  ( .A(_GFM_n20310 ), .B(_GFM_n20300 ), .Z(z_out[123]) );
XOR2_X2 _GFM_U2359  ( .A(_GFM_n20330 ), .B(_GFM_n2032 ), .Z(_GFM_n20300 ) );
XOR2_X2 _GFM_U2358  ( .A(_GFM_n20350 ), .B(_GFM_n2034 ), .Z(_GFM_n20310 ) );
XOR2_X2 _GFM_U2357  ( .A(_GFM_n2037 ), .B(_GFM_n20360 ), .Z(_GFM_n2032 ) );
XOR2_X2 _GFM_U2356  ( .A(_GFM_n20390 ), .B(_GFM_n2038 ), .Z(_GFM_n20330 ) );
XOR2_X2 _GFM_U2355  ( .A(_GFM_n20411 ), .B(_GFM_n20400 ), .Z(_GFM_n2034 ) );
XOR2_X2 _GFM_U2354  ( .A(_GFM_n20430 ), .B(_GFM_n20420 ), .Z(_GFM_n20350 ));
XOR2_X2 _GFM_U2353  ( .A(z_in[123]), .B(_GFM_n2044 ), .Z(_GFM_n20360 ) );
XOR2_X2 _GFM_U2352  ( .A(_GFM_N4151 ), .B(_GFM_N4154 ), .Z(_GFM_n2037 ) );
XOR2_X2 _GFM_U2351  ( .A(_GFM_N4144 ), .B(_GFM_N4147 ), .Z(_GFM_n2038 ) );
XOR2_X2 _GFM_U2350  ( .A(_GFM_N4136 ), .B(_GFM_N4139 ), .Z(_GFM_n20390 ) );
XOR2_X2 _GFM_U2349  ( .A(_GFM_N4129 ), .B(_GFM_N4132 ), .Z(_GFM_n20400 ) );
XOR2_X2 _GFM_U2348  ( .A(_GFM_N4120 ), .B(_GFM_N4123 ), .Z(_GFM_n20411 ) );
XOR2_X2 _GFM_U2347  ( .A(_GFM_N4113 ), .B(_GFM_N4116 ), .Z(_GFM_n20420 ) );
XOR2_X2 _GFM_U2346  ( .A(_GFM_N4106 ), .B(_GFM_N4108 ), .Z(_GFM_n20430 ) );
XOR2_X2 _GFM_U2345  ( .A(_GFM_N4102 ), .B(_GFM_N4103 ), .Z(_GFM_n2044 ) );
XOR2_X2 _GFM_U2344  ( .A(_GFM_n2046 ), .B(_GFM_n2045 ), .Z(z_out[124]) );
XOR2_X2 _GFM_U2343  ( .A(_GFM_n2048 ), .B(_GFM_n20470 ), .Z(_GFM_n2045 ) );
XOR2_X2 _GFM_U2342  ( .A(_GFM_n20500 ), .B(_GFM_n20490 ), .Z(_GFM_n2046 ) );
XOR2_X2 _GFM_U2341  ( .A(_GFM_n2052 ), .B(_GFM_n2051 ), .Z(_GFM_n20470 ) );
XOR2_X2 _GFM_U2340  ( .A(_GFM_n20540 ), .B(_GFM_n20530 ), .Z(_GFM_n2048 ) );
XOR2_X2 _GFM_U2339  ( .A(_GFM_n20560 ), .B(_GFM_n2055 ), .Z(_GFM_n20490 ) );
XOR2_X2 _GFM_U2338  ( .A(_GFM_n2058 ), .B(_GFM_n20570 ), .Z(_GFM_n20500 ) );
XOR2_X2 _GFM_U2337  ( .A(z_in[124]), .B(_GFM_n2059 ), .Z(_GFM_n2051 ) );
XOR2_X2 _GFM_U2336  ( .A(_GFM_N4210 ), .B(_GFM_N4213 ), .Z(_GFM_n2052 ) );
XOR2_X2 _GFM_U2335  ( .A(_GFM_N4203 ), .B(_GFM_N4206 ), .Z(_GFM_n20530 ) );
XOR2_X2 _GFM_U2334  ( .A(_GFM_N4195 ), .B(_GFM_N4198 ), .Z(_GFM_n20540 ) );
XOR2_X2 _GFM_U2333  ( .A(_GFM_N4188 ), .B(_GFM_N4191 ), .Z(_GFM_n2055 ) );
XOR2_X2 _GFM_U2332  ( .A(_GFM_N4179 ), .B(_GFM_N4182 ), .Z(_GFM_n20560 ) );
XOR2_X2 _GFM_U2331  ( .A(_GFM_N4172 ), .B(_GFM_N4175 ), .Z(_GFM_n20570 ) );
XOR2_X2 _GFM_U2330  ( .A(_GFM_N4164 ), .B(_GFM_N4167 ), .Z(_GFM_n2058 ) );
XOR2_X2 _GFM_U2329  ( .A(_GFM_N4159 ), .B(_GFM_N4160 ), .Z(_GFM_n2059 ) );
XOR2_X2 _GFM_U2328  ( .A(_GFM_n20610 ), .B(_GFM_n20601 ), .Z(z_out[125]) );
XOR2_X2 _GFM_U2327  ( .A(_GFM_n2063 ), .B(_GFM_n20620 ), .Z(_GFM_n20601 ) );
XOR2_X2 _GFM_U2326  ( .A(_GFM_n2065 ), .B(_GFM_n20640 ), .Z(_GFM_n20610 ) );
XOR2_X2 _GFM_U2325  ( .A(_GFM_n20670 ), .B(_GFM_n20660 ), .Z(_GFM_n20620 ));
XOR2_X2 _GFM_U2324  ( .A(_GFM_n2069 ), .B(_GFM_n2068 ), .Z(_GFM_n2063 ) );
XOR2_X2 _GFM_U2323  ( .A(_GFM_n20710 ), .B(_GFM_n20700 ), .Z(_GFM_n20640 ));
XOR2_X2 _GFM_U2322  ( .A(_GFM_n20730 ), .B(_GFM_n20721 ), .Z(_GFM_n2065 ) );
XOR2_X2 _GFM_U2321  ( .A(z_in[125]), .B(_GFM_n20740 ), .Z(_GFM_n20660 ) );
XOR2_X2 _GFM_U2320  ( .A(_GFM_N4269 ), .B(_GFM_N4272 ), .Z(_GFM_n20670 ) );
XOR2_X2 _GFM_U2319  ( .A(_GFM_N4263 ), .B(_GFM_N4265 ), .Z(_GFM_n2068 ) );
XOR2_X2 _GFM_U2318  ( .A(_GFM_N4255 ), .B(_GFM_N4258 ), .Z(_GFM_n2069 ) );
XOR2_X2 _GFM_U2317  ( .A(_GFM_N4249 ), .B(_GFM_N4251 ), .Z(_GFM_n20700 ) );
XOR2_X2 _GFM_U2316  ( .A(_GFM_N4240 ), .B(_GFM_N4243 ), .Z(_GFM_n20710 ) );
XOR2_X2 _GFM_U2315  ( .A(_GFM_N4233 ), .B(_GFM_N4236 ), .Z(_GFM_n20721 ) );
XOR2_X2 _GFM_U2314  ( .A(_GFM_N4225 ), .B(_GFM_N4228 ), .Z(_GFM_n20730 ) );
XOR2_X2 _GFM_U2313  ( .A(_GFM_N4218 ), .B(_GFM_N4221 ), .Z(_GFM_n20740 ) );
XOR2_X2 _GFM_U2312  ( .A(_GFM_n2076 ), .B(_GFM_n2075 ), .Z(z_out[126]) );
XOR2_X2 _GFM_U2311  ( .A(_GFM_n20780 ), .B(_GFM_n2077 ), .Z(_GFM_n2075 ) );
XOR2_X2 _GFM_U2310  ( .A(_GFM_n20800 ), .B(_GFM_n2079 ), .Z(_GFM_n2076 ) );
XOR2_X2 _GFM_U2309  ( .A(_GFM_n2082 ), .B(_GFM_n20810 ), .Z(_GFM_n2077 ) );
XOR2_X2 _GFM_U2308  ( .A(_GFM_n20840 ), .B(_GFM_n2083 ), .Z(_GFM_n20780 ) );
XOR2_X2 _GFM_U2307  ( .A(_GFM_n2086 ), .B(_GFM_n20850 ), .Z(_GFM_n2079 ) );
XOR2_X2 _GFM_U2306  ( .A(_GFM_n20880 ), .B(_GFM_n20870 ), .Z(_GFM_n20800 ));
XOR2_X2 _GFM_U2305  ( .A(z_in[126]), .B(_GFM_n2089 ), .Z(_GFM_n20810 ) );
XOR2_X2 _GFM_U2304  ( .A(_GFM_N4316 ), .B(_GFM_N4318 ), .Z(_GFM_n2082 ) );
XOR2_X2 _GFM_U2303  ( .A(_GFM_N4311 ), .B(_GFM_N4313 ), .Z(_GFM_n2083 ) );
XOR2_X2 _GFM_U2302  ( .A(_GFM_N4305 ), .B(_GFM_N4307 ), .Z(_GFM_n20840 ) );
XOR2_X2 _GFM_U2301  ( .A(_GFM_N4300 ), .B(_GFM_N4302 ), .Z(_GFM_n20850 ) );
XOR2_X2 _GFM_U2300  ( .A(_GFM_N4293 ), .B(_GFM_N4295 ), .Z(_GFM_n2086 ) );
XOR2_X2 _GFM_U2299  ( .A(_GFM_N4288 ), .B(_GFM_N4290 ), .Z(_GFM_n20870 ) );
XOR2_X2 _GFM_U2298  ( .A(_GFM_N4282 ), .B(_GFM_N4284 ), .Z(_GFM_n20880 ) );
XOR2_X2 _GFM_U2297  ( .A(_GFM_N4276 ), .B(_GFM_N4279 ), .Z(_GFM_n2089 ) );
XOR2_X2 _GFM_U2296  ( .A(_GFM_n2091 ), .B(_GFM_n2090 ), .Z(z_out[127]) );
XOR2_X2 _GFM_U2295  ( .A(_GFM_n20930 ), .B(_GFM_n20920 ), .Z(_GFM_n2090 ) );
XOR2_X2 _GFM_U2294  ( .A(_GFM_n20950 ), .B(_GFM_n2094 ), .Z(_GFM_n2091 ) );
XOR2_X2 _GFM_U2293  ( .A(_GFM_n20970 ), .B(_GFM_n2096 ), .Z(_GFM_n20920 ) );
XOR2_X2 _GFM_U2292  ( .A(_GFM_n2099 ), .B(_GFM_n20980 ), .Z(_GFM_n20930 ) );
XOR2_X2 _GFM_U2291  ( .A(_GFM_n21010 ), .B(_GFM_n21001 ), .Z(_GFM_n2094 ) );
XOR2_X2 _GFM_U2290  ( .A(_GFM_n2103 ), .B(_GFM_n21020 ), .Z(_GFM_n20950 ) );
XOR2_X2 _GFM_U2289  ( .A(z_in[127]), .B(_GFM_n21040 ), .Z(_GFM_n2096 ) );
XOR2_X2 _GFM_U2288  ( .A(_GFM_N4348 ), .B(_GFM_N4349 ), .Z(_GFM_n20970 ) );
XOR2_X2 _GFM_U2287  ( .A(_GFM_N4345 ), .B(_GFM_N4346 ), .Z(_GFM_n20980 ) );
XOR2_X2 _GFM_U2286  ( .A(_GFM_N4341 ), .B(_GFM_N4342 ), .Z(_GFM_n2099 ) );
XOR2_X2 _GFM_U2285  ( .A(_GFM_N4337 ), .B(_GFM_N4339 ), .Z(_GFM_n21001 ) );
XOR2_X2 _GFM_U2284  ( .A(_GFM_N4332 ), .B(_GFM_N4336 ), .Z(_GFM_n21010 ) );
XOR2_X2 _GFM_U2283  ( .A(_GFM_N4329 ), .B(_GFM_N4331 ), .Z(_GFM_n21020 ) );
XOR2_X2 _GFM_U2282  ( .A(_GFM_N4325 ), .B(_GFM_N4328 ), .Z(_GFM_n2103 ) );
XOR2_X2 _GFM_U2281  ( .A(_GFM_N4322 ), .B(_GFM_N4324 ), .Z(_GFM_n21040 ) );
XOR2_X2 _GFM_U2280  ( .A(v_in[0]), .B(_GFM_n21050 ), .Z(v_out[110]) );
XOR2_X2 _GFM_U2279  ( .A(v_in[126]), .B(v_in[5]), .Z(_GFM_n21050 ) );
XOR2_X2 _GFM_U2278  ( .A(v_in[0]), .B(_GFM_n2106 ), .Z(_GFM_N4224 ) );
XOR2_X2 _GFM_U2277  ( .A(v_in[127]), .B(v_in[1]), .Z(_GFM_n2106 ) );
XOR2_X2 _GFM_U2276  ( .A(v_in[6]), .B(_GFM_N4224 ), .Z(v_out[111]) );
XOR2_X2 _GFM_U2275  ( .A(v_in[0]), .B(_GFM_n2107 ), .Z(_GFM_N4227 ) );
XOR2_X2 _GFM_U2274  ( .A(v_in[2]), .B(v_in[1]), .Z(_GFM_n2107 ) );
XOR2_X2 _GFM_U2273  ( .A(v_in[7]), .B(_GFM_N4227 ), .Z(v_out[112]) );
XOR2_X2 _GFM_U2272  ( .A(v_in[1]), .B(_GFM_n2108 ), .Z(_GFM_N4235 ) );
XOR2_X2 _GFM_U2271  ( .A(v_in[3]), .B(v_in[2]), .Z(_GFM_n2108 ) );
XOR2_X2 _GFM_U2270  ( .A(v_in[8]), .B(_GFM_N4235 ), .Z(v_out[113]) );
XOR2_X2 _GFM_U2269  ( .A(v_in[2]), .B(_GFM_n21090 ), .Z(_GFM_N4232 ) );
XOR2_X2 _GFM_U2268  ( .A(v_in[4]), .B(v_in[3]), .Z(_GFM_n21090 ) );
XOR2_X2 _GFM_U2267  ( .A(v_in[9]), .B(_GFM_N4232 ), .Z(v_out[114]) );
XOR2_X2 _GFM_U2266  ( .A(v_in[3]), .B(_GFM_n21101 ), .Z(_GFM_N4239 ) );
XOR2_X2 _GFM_U2265  ( .A(v_in[5]), .B(v_in[4]), .Z(_GFM_n21101 ) );
XOR2_X2 _GFM_U2264  ( .A(v_in[10]), .B(_GFM_N4239 ), .Z(v_out[115]) );
XOR2_X2 _GFM_U2263  ( .A(v_in[4]), .B(_GFM_n21110 ), .Z(_GFM_N4242 ) );
XOR2_X2 _GFM_U2262  ( .A(v_in[6]), .B(v_in[5]), .Z(_GFM_n21110 ) );
XOR2_X2 _GFM_U2261  ( .A(v_in[11]), .B(_GFM_N4242 ), .Z(v_out[116]) );
XOR2_X2 _GFM_U2260  ( .A(v_in[5]), .B(_GFM_n21120 ), .Z(_GFM_N4257 ) );
XOR2_X2 _GFM_U2259  ( .A(v_in[7]), .B(v_in[6]), .Z(_GFM_n21120 ) );
XOR2_X2 _GFM_U2258  ( .A(v_in[12]), .B(_GFM_N4257 ), .Z(v_out[117]) );
XOR2_X2 _GFM_U2257  ( .A(v_in[6]), .B(_GFM_n2113 ), .Z(_GFM_N4254 ) );
XOR2_X2 _GFM_U2256  ( .A(v_in[8]), .B(v_in[7]), .Z(_GFM_n2113 ) );
XOR2_X2 _GFM_U2255  ( .A(v_in[13]), .B(_GFM_N4254 ), .Z(v_out[118]) );
XOR2_X2 _GFM_U2254  ( .A(v_in[7]), .B(_GFM_n2114 ), .Z(_GFM_N4248 ) );
XOR2_X2 _GFM_U2253  ( .A(v_in[9]), .B(v_in[8]), .Z(_GFM_n2114 ) );
XOR2_X2 _GFM_U2252  ( .A(v_in[14]), .B(_GFM_N4248 ), .Z(v_out[119]) );
XOR2_X2 _GFM_U2251  ( .A(v_in[8]), .B(_GFM_n21150 ), .Z(_GFM_N4250 ) );
XOR2_X2 _GFM_U2250  ( .A(v_in[10]), .B(v_in[9]), .Z(_GFM_n21150 ) );
XOR2_X2 _GFM_U2249  ( .A(v_in[15]), .B(_GFM_N4250 ), .Z(v_out[120]) );
XOR2_X2 _GFM_U2248  ( .A(v_in[9]), .B(_GFM_n21160 ), .Z(v_out[121]) );
XOR2_X2 _GFM_U2247  ( .A(v_in[11]), .B(v_in[10]), .Z(_GFM_n21160 ) );
XOR2_X2 _GFM_U2246  ( .A(v_in[10]), .B(_GFM_n2117 ), .Z(v_out[122]) );
XOR2_X2 _GFM_U2245  ( .A(v_in[12]), .B(v_in[11]), .Z(_GFM_n2117 ) );
XOR2_X2 _GFM_U2244  ( .A(v_in[11]), .B(_GFM_n21180 ), .Z(v_out[123]) );
XOR2_X2 _GFM_U2243  ( .A(v_in[13]), .B(v_in[12]), .Z(_GFM_n21180 ) );
XOR2_X2 _GFM_U2242  ( .A(v_in[12]), .B(_GFM_n21190 ), .Z(v_out[124]) );
XOR2_X2 _GFM_U2241  ( .A(v_in[14]), .B(v_in[13]), .Z(_GFM_n21190 ) );
XOR2_X2 _GFM_U2240  ( .A(v_in[13]), .B(_GFM_n2120 ), .Z(v_out[125]) );
XOR2_X2 _GFM_U2239  ( .A(v_in[15]), .B(v_in[14]), .Z(_GFM_n2120 ) );
INV_X4 _AES_ENC_U1636  ( .A(rst), .ZN(_AES_ENC_n1267 ) );
INV_X4 _AES_ENC_U1635  ( .A(_AES_ENC_n17 ), .ZN(_AES_ENC_n1266 ) );
NAND3_X2 _AES_ENC_U1634  ( .A1(_AES_ENC_n15 ), .A2(_AES_ENC_n1258 ), .A3(_AES_ENC_n16 ), .ZN(_AES_ENC_n796 ) );
NOR2_X2 _AES_ENC_U1633  ( .A1(_AES_ENC_n22 ), .A2(_AES_ENC_n2 ), .ZN(_AES_ENC_n17 ) );
NOR2_X2 _AES_ENC_U1632  ( .A1(_AES_ENC_n1234 ), .A2(_AES_ENC_n1231 ), .ZN(_AES_ENC_n14 ) );
NOR2_X2 _AES_ENC_U1631  ( .A1(_AES_ENC_n1232 ), .A2(_AES_ENC_n22 ), .ZN(_AES_ENC_n11 ) );
INV_X4 _AES_ENC_U1630  ( .A(_AES_ENC_n1258 ), .ZN(_AES_ENC_n1265 ) );
INV_X4 _AES_ENC_U1629  ( .A(_AES_ENC_n1256 ), .ZN(_AES_ENC_n1250 ) );
INV_X4 _AES_ENC_U1628  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1246 ) );
INV_X4 _AES_ENC_U1627  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1247 ) );
INV_X4 _AES_ENC_U1626  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1245 ) );
INV_X4 _AES_ENC_U1625  ( .A(_AES_ENC_n1255 ), .ZN(_AES_ENC_n1248 ) );
INV_X4 _AES_ENC_U1624  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1249 ) );
INV_X4 _AES_ENC_U1623  ( .A(_AES_ENC_n1265 ), .ZN(_AES_ENC_n1259 ) );
INV_X4 _AES_ENC_U1622  ( .A(_AES_ENC_n1238 ), .ZN(_AES_ENC_n1254 ) );
INV_X4 _AES_ENC_U1621  ( .A(_AES_ENC_n1238 ), .ZN(_AES_ENC_n1253 ) );
INV_X4 _AES_ENC_U1620  ( .A(_AES_ENC_n1238 ), .ZN(_AES_ENC_n1252 ) );
INV_X4 _AES_ENC_U1619  ( .A(_AES_ENC_n1238 ), .ZN(_AES_ENC_n1256 ) );
INV_X4 _AES_ENC_U1618  ( .A(_AES_ENC_n1238 ), .ZN(_AES_ENC_n1255 ) );
INV_X4 _AES_ENC_U1617  ( .A(_AES_ENC_n1238 ), .ZN(_AES_ENC_n1251 ) );
INV_X4 _AES_ENC_U1616  ( .A(_AES_ENC_n1265 ), .ZN(_AES_ENC_n12601 ) );
INV_X4 _AES_ENC_U1615  ( .A(_AES_ENC_n1265 ), .ZN(_AES_ENC_n1261 ) );
INV_X4 _AES_ENC_U1614  ( .A(_AES_ENC_n1265 ), .ZN(_AES_ENC_n1262 ) );
INV_X4 _AES_ENC_U1613  ( .A(_AES_ENC_n1265 ), .ZN(_AES_ENC_n1263 ) );
INV_X4 _AES_ENC_U1052  ( .A(_AES_ENC_n1265 ), .ZN(_AES_ENC_n1264 ) );
INV_X4 _AES_ENC_U1051  ( .A(aes_kld), .ZN(_AES_ENC_n1258 ) );
INV_X4 _AES_ENC_U1050  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1244 ) );
INV_X4 _AES_ENC_U1049  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1241 ) );
INV_X4 _AES_ENC_U1048  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1239 ) );
INV_X4 _AES_ENC_U1047  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1242 ) );
INV_X4 _AES_ENC_U1046  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1243 ) );
INV_X4 _AES_ENC_U1045  ( .A(_AES_ENC_n793 ), .ZN(_AES_ENC_n1240 ) );
INV_X4 _AES_ENC_U876  ( .A(_AES_ENC_n1258 ), .ZN(_AES_ENC_n1257 ) );
INV_X4 _AES_ENC_U16  ( .A(_AES_ENC_n1258 ), .ZN(_AES_ENC_n1237 ) );
INV_X4 _AES_ENC_U14  ( .A(_AES_ENC_n1258 ), .ZN(_AES_ENC_n1236 ) );
INV_X4 _AES_ENC_U7  ( .A(_AES_ENC_n1258 ), .ZN(_AES_ENC_n1235 ) );
CLKBUFX1 gbuf_d_780(.A(aes_kld), .Y(ddout__780));
CLKBUFX1 gbuf_q_780(.A(qq_in780), .Y(_AES_ENC_n1238));
CLKBUFX1 gbuf_qn_780(.A(qnn_in_780), .Y(_AES_ENC_n793));
NAND2_X2 _AES_ENC_U1044  ( .A1(_AES_ENC_sa32_next[6]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n7891 ) );
XOR2_X2 _AES_ENC_U1043  ( .A(_AES_ENC_w2[6] ), .B(_AES_ENC_text_in_r[38] ),.Z(_AES_ENC_n791 ) );
NAND2_X2 _AES_ENC_U1042  ( .A1(_AES_ENC_n791 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n7901 ) );
NAND2_X2 _AES_ENC_U1041  ( .A1(_AES_ENC_n7891 ), .A2(_AES_ENC_n7901 ), .ZN(_AES_ENC_N100 ) );
NAND2_X2 _AES_ENC_U1040  ( .A1(_AES_ENC_sa32_next[7]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n658 ) );
XOR2_X2 _AES_ENC_U1039  ( .A(_AES_ENC_w2[7] ), .B(_AES_ENC_text_in_r[39] ),.Z(_AES_ENC_n6601 ) );
NAND2_X2 _AES_ENC_U1038  ( .A1(_AES_ENC_n6601 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n659 ) );
NAND2_X2 _AES_ENC_U1037  ( .A1(_AES_ENC_n658 ), .A2(_AES_ENC_n659 ), .ZN(_AES_ENC_N101 ) );
NAND2_X2 _AES_ENC_U1036  ( .A1(_AES_ENC_sa22_next[0]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n655 ) );
XOR2_X2 _AES_ENC_U1035  ( .A(_AES_ENC_w2[8] ), .B(_AES_ENC_text_in_r[40] ),.Z(_AES_ENC_n657 ) );
NAND2_X2 _AES_ENC_U1034  ( .A1(_AES_ENC_n657 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n656 ) );
NAND2_X2 _AES_ENC_U1033  ( .A1(_AES_ENC_n655 ), .A2(_AES_ENC_n656 ), .ZN(_AES_ENC_N110 ) );
NAND2_X2 _AES_ENC_U1032  ( .A1(_AES_ENC_sa22_next[1]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n652 ) );
XOR2_X2 _AES_ENC_U1031  ( .A(_AES_ENC_w2[9] ), .B(_AES_ENC_text_in_r[41] ),.Z(_AES_ENC_n654 ) );
NAND2_X2 _AES_ENC_U1030  ( .A1(_AES_ENC_n654 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n653 ) );
NAND2_X2 _AES_ENC_U1029  ( .A1(_AES_ENC_n652 ), .A2(_AES_ENC_n653 ), .ZN(_AES_ENC_N111 ) );
NAND2_X2 _AES_ENC_U1028  ( .A1(_AES_ENC_sa22_next[2]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n649 ) );
XOR2_X2 _AES_ENC_U1027  ( .A(_AES_ENC_w2[10] ), .B(_AES_ENC_text_in_r[42] ),.Z(_AES_ENC_n651 ) );
NAND2_X2 _AES_ENC_U1026  ( .A1(_AES_ENC_n651 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n6501 ) );
NAND2_X2 _AES_ENC_U1025  ( .A1(_AES_ENC_n649 ), .A2(_AES_ENC_n6501 ), .ZN(_AES_ENC_N112 ) );
NAND2_X2 _AES_ENC_U1024  ( .A1(_AES_ENC_sa22_next[3]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n646 ) );
XOR2_X2 _AES_ENC_U1023  ( .A(_AES_ENC_w2[11] ), .B(_AES_ENC_text_in_r[43] ),.Z(_AES_ENC_n648 ) );
NAND2_X2 _AES_ENC_U1022  ( .A1(_AES_ENC_n648 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n647 ) );
NAND2_X2 _AES_ENC_U1021  ( .A1(_AES_ENC_n646 ), .A2(_AES_ENC_n647 ), .ZN(_AES_ENC_N113 ) );
NAND2_X2 _AES_ENC_U1020  ( .A1(_AES_ENC_sa22_next[4]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n643 ) );
XOR2_X2 _AES_ENC_U1019  ( .A(_AES_ENC_w2[12] ), .B(_AES_ENC_text_in_r[44] ),.Z(_AES_ENC_n645 ) );
NAND2_X2 _AES_ENC_U1018  ( .A1(_AES_ENC_n645 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n644 ) );
NAND2_X2 _AES_ENC_U1017  ( .A1(_AES_ENC_n643 ), .A2(_AES_ENC_n644 ), .ZN(_AES_ENC_N114 ) );
NAND2_X2 _AES_ENC_U1016  ( .A1(_AES_ENC_sa22_next[5]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n6401 ) );
XOR2_X2 _AES_ENC_U1015  ( .A(_AES_ENC_w2[13] ), .B(_AES_ENC_text_in_r[45] ),.Z(_AES_ENC_n642 ) );
NAND2_X2 _AES_ENC_U1014  ( .A1(_AES_ENC_n642 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n641 ) );
NAND2_X2 _AES_ENC_U1013  ( .A1(_AES_ENC_n6401 ), .A2(_AES_ENC_n641 ), .ZN(_AES_ENC_N115 ) );
NAND2_X2 _AES_ENC_U1012  ( .A1(_AES_ENC_sa22_next[6]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n637 ) );
XOR2_X2 _AES_ENC_U1011  ( .A(_AES_ENC_w2[14] ), .B(_AES_ENC_text_in_r[46] ),.Z(_AES_ENC_n639 ) );
NAND2_X2 _AES_ENC_U1010  ( .A1(_AES_ENC_n639 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n638 ) );
NAND2_X2 _AES_ENC_U1009  ( .A1(_AES_ENC_n637 ), .A2(_AES_ENC_n638 ), .ZN(_AES_ENC_N116 ) );
NAND2_X2 _AES_ENC_U1008  ( .A1(_AES_ENC_sa22_next[7]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n634 ) );
XOR2_X2 _AES_ENC_U1007  ( .A(_AES_ENC_w2[15] ), .B(_AES_ENC_text_in_r[47] ),.Z(_AES_ENC_n636 ) );
NAND2_X2 _AES_ENC_U1006  ( .A1(_AES_ENC_n636 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n635 ) );
NAND2_X2 _AES_ENC_U1005  ( .A1(_AES_ENC_n634 ), .A2(_AES_ENC_n635 ), .ZN(_AES_ENC_N117 ) );
NAND2_X2 _AES_ENC_U1004  ( .A1(_AES_ENC_sa12_next[0]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n631 ) );
XOR2_X2 _AES_ENC_U1003  ( .A(_AES_ENC_w2[16] ), .B(_AES_ENC_text_in_r[48] ),.Z(_AES_ENC_n633 ) );
NAND2_X2 _AES_ENC_U1002  ( .A1(_AES_ENC_n633 ), .A2(_AES_ENC_n1239 ), .ZN(_AES_ENC_n632 ) );
NAND2_X2 _AES_ENC_U1001  ( .A1(_AES_ENC_n631 ), .A2(_AES_ENC_n632 ), .ZN(_AES_ENC_N126 ) );
NAND2_X2 _AES_ENC_U1000  ( .A1(_AES_ENC_sa12_next[1]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n628 ) );
XOR2_X2 _AES_ENC_U999  ( .A(_AES_ENC_w2[17] ), .B(_AES_ENC_text_in_r[49] ),.Z(_AES_ENC_n6301 ) );
NAND2_X2 _AES_ENC_U998  ( .A1(_AES_ENC_n6301 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n629 ) );
NAND2_X2 _AES_ENC_U997  ( .A1(_AES_ENC_n628 ), .A2(_AES_ENC_n629 ), .ZN(_AES_ENC_N127 ) );
NAND2_X2 _AES_ENC_U996  ( .A1(_AES_ENC_sa12_next[2]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n625 ) );
XOR2_X2 _AES_ENC_U995  ( .A(_AES_ENC_w2[18] ), .B(_AES_ENC_text_in_r[50] ),.Z(_AES_ENC_n627 ) );
NAND2_X2 _AES_ENC_U994  ( .A1(_AES_ENC_n627 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n626 ) );
NAND2_X2 _AES_ENC_U993  ( .A1(_AES_ENC_n625 ), .A2(_AES_ENC_n626 ), .ZN(_AES_ENC_N128 ) );
NAND2_X2 _AES_ENC_U992  ( .A1(_AES_ENC_sa12_next[3]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n622 ) );
XOR2_X2 _AES_ENC_U991  ( .A(_AES_ENC_w2[19] ), .B(_AES_ENC_text_in_r[51] ),.Z(_AES_ENC_n624 ) );
NAND2_X2 _AES_ENC_U990  ( .A1(_AES_ENC_n624 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n623 ) );
NAND2_X2 _AES_ENC_U989  ( .A1(_AES_ENC_n622 ), .A2(_AES_ENC_n623 ), .ZN(_AES_ENC_N129 ) );
NAND2_X2 _AES_ENC_U988  ( .A1(_AES_ENC_sa12_next[4]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n619 ) );
XOR2_X2 _AES_ENC_U987  ( .A(_AES_ENC_w2[20] ), .B(_AES_ENC_text_in_r[52] ),.Z(_AES_ENC_n621 ) );
NAND2_X2 _AES_ENC_U986  ( .A1(_AES_ENC_n621 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n6201 ) );
NAND2_X2 _AES_ENC_U985  ( .A1(_AES_ENC_n619 ), .A2(_AES_ENC_n6201 ), .ZN(_AES_ENC_N130 ) );
NAND2_X2 _AES_ENC_U984  ( .A1(_AES_ENC_sa12_next[5]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n616 ) );
XOR2_X2 _AES_ENC_U983  ( .A(_AES_ENC_w2[21] ), .B(_AES_ENC_text_in_r[53] ),.Z(_AES_ENC_n618 ) );
NAND2_X2 _AES_ENC_U982  ( .A1(_AES_ENC_n618 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n617 ) );
NAND2_X2 _AES_ENC_U981  ( .A1(_AES_ENC_n616 ), .A2(_AES_ENC_n617 ), .ZN(_AES_ENC_N131 ) );
NAND2_X2 _AES_ENC_U980  ( .A1(_AES_ENC_sa12_next[6]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n613 ) );
XOR2_X2 _AES_ENC_U979  ( .A(_AES_ENC_w2[22] ), .B(_AES_ENC_text_in_r[54] ),.Z(_AES_ENC_n615 ) );
NAND2_X2 _AES_ENC_U978  ( .A1(_AES_ENC_n615 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n614 ) );
NAND2_X2 _AES_ENC_U977  ( .A1(_AES_ENC_n613 ), .A2(_AES_ENC_n614 ), .ZN(_AES_ENC_N132 ) );
NAND2_X2 _AES_ENC_U976  ( .A1(_AES_ENC_sa12_next[7]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n610 ) );
XOR2_X2 _AES_ENC_U975  ( .A(_AES_ENC_w2[23] ), .B(_AES_ENC_text_in_r[55] ),.Z(_AES_ENC_n612 ) );
NAND2_X2 _AES_ENC_U974  ( .A1(_AES_ENC_n612 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n611 ) );
NAND2_X2 _AES_ENC_U973  ( .A1(_AES_ENC_n610 ), .A2(_AES_ENC_n611 ), .ZN(_AES_ENC_N133 ) );
NAND2_X2 _AES_ENC_U972  ( .A1(_AES_ENC_sa02_next[0]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n607 ) );
XOR2_X2 _AES_ENC_U971  ( .A(_AES_ENC_w2[24] ), .B(_AES_ENC_text_in_r[56] ),.Z(_AES_ENC_n609 ) );
NAND2_X2 _AES_ENC_U970  ( .A1(_AES_ENC_n609 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n608 ) );
NAND2_X2 _AES_ENC_U969  ( .A1(_AES_ENC_n607 ), .A2(_AES_ENC_n608 ), .ZN(_AES_ENC_N142 ) );
NAND2_X2 _AES_ENC_U968  ( .A1(_AES_ENC_sa02_next[1]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n604 ) );
XOR2_X2 _AES_ENC_U967  ( .A(_AES_ENC_w2[25] ), .B(_AES_ENC_text_in_r[57] ),.Z(_AES_ENC_n606 ) );
NAND2_X2 _AES_ENC_U966  ( .A1(_AES_ENC_n606 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n605 ) );
NAND2_X2 _AES_ENC_U965  ( .A1(_AES_ENC_n604 ), .A2(_AES_ENC_n605 ), .ZN(_AES_ENC_N143 ) );
NAND2_X2 _AES_ENC_U964  ( .A1(_AES_ENC_sa02_next[2]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n601 ) );
XOR2_X2 _AES_ENC_U963  ( .A(_AES_ENC_w2[26] ), .B(_AES_ENC_text_in_r[58] ),.Z(_AES_ENC_n603 ) );
NAND2_X2 _AES_ENC_U962  ( .A1(_AES_ENC_n603 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n602 ) );
NAND2_X2 _AES_ENC_U961  ( .A1(_AES_ENC_n601 ), .A2(_AES_ENC_n602 ), .ZN(_AES_ENC_N144 ) );
NAND2_X2 _AES_ENC_U960  ( .A1(_AES_ENC_sa02_next[3]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n598 ) );
XOR2_X2 _AES_ENC_U959  ( .A(_AES_ENC_w2[27] ), .B(_AES_ENC_text_in_r[59] ),.Z(_AES_ENC_n600 ) );
NAND2_X2 _AES_ENC_U958  ( .A1(_AES_ENC_n600 ), .A2(_AES_ENC_n1240 ), .ZN(_AES_ENC_n599 ) );
NAND2_X2 _AES_ENC_U957  ( .A1(_AES_ENC_n598 ), .A2(_AES_ENC_n599 ), .ZN(_AES_ENC_N145 ) );
NAND2_X2 _AES_ENC_U956  ( .A1(_AES_ENC_sa02_next[4]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n595 ) );
XOR2_X2 _AES_ENC_U955  ( .A(_AES_ENC_w2[28] ), .B(_AES_ENC_text_in_r[60] ),.Z(_AES_ENC_n597 ) );
NAND2_X2 _AES_ENC_U954  ( .A1(_AES_ENC_n597 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n596 ) );
NAND2_X2 _AES_ENC_U953  ( .A1(_AES_ENC_n595 ), .A2(_AES_ENC_n596 ), .ZN(_AES_ENC_N146 ) );
NAND2_X2 _AES_ENC_U952  ( .A1(_AES_ENC_sa02_next[5]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n592 ) );
XOR2_X2 _AES_ENC_U951  ( .A(_AES_ENC_w2[29] ), .B(_AES_ENC_text_in_r[61] ),.Z(_AES_ENC_n594 ) );
NAND2_X2 _AES_ENC_U950  ( .A1(_AES_ENC_n594 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n593 ) );
NAND2_X2 _AES_ENC_U949  ( .A1(_AES_ENC_n592 ), .A2(_AES_ENC_n593 ), .ZN(_AES_ENC_N147 ) );
NAND2_X2 _AES_ENC_U948  ( .A1(_AES_ENC_sa02_next[6]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n589 ) );
XOR2_X2 _AES_ENC_U947  ( .A(_AES_ENC_w2[30] ), .B(_AES_ENC_text_in_r[62] ),.Z(_AES_ENC_n591 ) );
NAND2_X2 _AES_ENC_U946  ( .A1(_AES_ENC_n591 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n590 ) );
NAND2_X2 _AES_ENC_U945  ( .A1(_AES_ENC_n589 ), .A2(_AES_ENC_n590 ), .ZN(_AES_ENC_N148 ) );
NAND2_X2 _AES_ENC_U944  ( .A1(_AES_ENC_sa02_next[7]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n586 ) );
XOR2_X2 _AES_ENC_U943  ( .A(_AES_ENC_w2[31] ), .B(_AES_ENC_text_in_r[63] ),.Z(_AES_ENC_n588 ) );
NAND2_X2 _AES_ENC_U942  ( .A1(_AES_ENC_n588 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n587 ) );
NAND2_X2 _AES_ENC_U941  ( .A1(_AES_ENC_n586 ), .A2(_AES_ENC_n587 ), .ZN(_AES_ENC_N149 ) );
NAND2_X2 _AES_ENC_U940  ( .A1(_AES_ENC_sa31_next[0]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n583 ) );
XOR2_X2 _AES_ENC_U939  ( .A(_AES_ENC_w1[0] ), .B(_AES_ENC_text_in_r[64] ),.Z(_AES_ENC_n585 ) );
NAND2_X2 _AES_ENC_U938  ( .A1(_AES_ENC_n585 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n584 ) );
NAND2_X2 _AES_ENC_U937  ( .A1(_AES_ENC_n583 ), .A2(_AES_ENC_n584 ), .ZN(_AES_ENC_N158 ) );
NAND2_X2 _AES_ENC_U936  ( .A1(_AES_ENC_sa31_next[1]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n580 ) );
XOR2_X2 _AES_ENC_U935  ( .A(_AES_ENC_w1[1] ), .B(_AES_ENC_text_in_r[65] ),.Z(_AES_ENC_n582 ) );
NAND2_X2 _AES_ENC_U934  ( .A1(_AES_ENC_n582 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n581 ) );
NAND2_X2 _AES_ENC_U933  ( .A1(_AES_ENC_n580 ), .A2(_AES_ENC_n581 ), .ZN(_AES_ENC_N159 ) );
NAND2_X2 _AES_ENC_U932  ( .A1(_AES_ENC_sa31_next[2]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n577 ) );
XOR2_X2 _AES_ENC_U931  ( .A(_AES_ENC_w1[2] ), .B(_AES_ENC_text_in_r[66] ),.Z(_AES_ENC_n579 ) );
NAND2_X2 _AES_ENC_U930  ( .A1(_AES_ENC_n579 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n578 ) );
NAND2_X2 _AES_ENC_U929  ( .A1(_AES_ENC_n577 ), .A2(_AES_ENC_n578 ), .ZN(_AES_ENC_N160 ) );
NAND2_X2 _AES_ENC_U928  ( .A1(_AES_ENC_sa31_next[3]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n574 ) );
XOR2_X2 _AES_ENC_U927  ( .A(_AES_ENC_w1[3] ), .B(_AES_ENC_text_in_r[67] ),.Z(_AES_ENC_n576 ) );
NAND2_X2 _AES_ENC_U926  ( .A1(_AES_ENC_n576 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n575 ) );
NAND2_X2 _AES_ENC_U925  ( .A1(_AES_ENC_n574 ), .A2(_AES_ENC_n575 ), .ZN(_AES_ENC_N161 ) );
NAND2_X2 _AES_ENC_U924  ( .A1(_AES_ENC_sa31_next[4]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n571 ) );
XOR2_X2 _AES_ENC_U923  ( .A(_AES_ENC_w1[4] ), .B(_AES_ENC_text_in_r[68] ),.Z(_AES_ENC_n573 ) );
NAND2_X2 _AES_ENC_U922  ( .A1(_AES_ENC_n573 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n572 ) );
NAND2_X2 _AES_ENC_U921  ( .A1(_AES_ENC_n571 ), .A2(_AES_ENC_n572 ), .ZN(_AES_ENC_N162 ) );
NAND2_X2 _AES_ENC_U920  ( .A1(_AES_ENC_sa31_next[5]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n568 ) );
XOR2_X2 _AES_ENC_U919  ( .A(_AES_ENC_w1[5] ), .B(_AES_ENC_text_in_r[69] ),.Z(_AES_ENC_n570 ) );
NAND2_X2 _AES_ENC_U918  ( .A1(_AES_ENC_n570 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n569 ) );
NAND2_X2 _AES_ENC_U917  ( .A1(_AES_ENC_n568 ), .A2(_AES_ENC_n569 ), .ZN(_AES_ENC_N163 ) );
NAND2_X2 _AES_ENC_U916  ( .A1(_AES_ENC_sa31_next[6]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n565 ) );
XOR2_X2 _AES_ENC_U915  ( .A(_AES_ENC_w1[6] ), .B(_AES_ENC_text_in_r[70] ),.Z(_AES_ENC_n567 ) );
NAND2_X2 _AES_ENC_U914  ( .A1(_AES_ENC_n567 ), .A2(_AES_ENC_n1241 ), .ZN(_AES_ENC_n566 ) );
NAND2_X2 _AES_ENC_U913  ( .A1(_AES_ENC_n565 ), .A2(_AES_ENC_n566 ), .ZN(_AES_ENC_N164 ) );
NAND2_X2 _AES_ENC_U912  ( .A1(_AES_ENC_sa31_next[7]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n562 ) );
XOR2_X2 _AES_ENC_U911  ( .A(_AES_ENC_w1[7] ), .B(_AES_ENC_text_in_r[71] ),.Z(_AES_ENC_n564 ) );
NAND2_X2 _AES_ENC_U910  ( .A1(_AES_ENC_n564 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n563 ) );
NAND2_X2 _AES_ENC_U909  ( .A1(_AES_ENC_n562 ), .A2(_AES_ENC_n563 ), .ZN(_AES_ENC_N165 ) );
NAND2_X2 _AES_ENC_U908  ( .A1(_AES_ENC_sa21_next[0]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n559 ) );
XOR2_X2 _AES_ENC_U907  ( .A(_AES_ENC_w1[8] ), .B(_AES_ENC_text_in_r[72] ),.Z(_AES_ENC_n561 ) );
NAND2_X2 _AES_ENC_U906  ( .A1(_AES_ENC_n561 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n560 ) );
NAND2_X2 _AES_ENC_U905  ( .A1(_AES_ENC_n559 ), .A2(_AES_ENC_n560 ), .ZN(_AES_ENC_N174 ) );
NAND2_X2 _AES_ENC_U904  ( .A1(_AES_ENC_sa21_next[1]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n556 ) );
XOR2_X2 _AES_ENC_U903  ( .A(_AES_ENC_w1[9] ), .B(_AES_ENC_text_in_r[73] ),.Z(_AES_ENC_n558 ) );
NAND2_X2 _AES_ENC_U902  ( .A1(_AES_ENC_n558 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n557 ) );
NAND2_X2 _AES_ENC_U901  ( .A1(_AES_ENC_n556 ), .A2(_AES_ENC_n557 ), .ZN(_AES_ENC_N175 ) );
NAND2_X2 _AES_ENC_U900  ( .A1(_AES_ENC_sa21_next[2]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n553 ) );
XOR2_X2 _AES_ENC_U899  ( .A(_AES_ENC_w1[10] ), .B(_AES_ENC_text_in_r[74] ),.Z(_AES_ENC_n555 ) );
NAND2_X2 _AES_ENC_U898  ( .A1(_AES_ENC_n555 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n554 ) );
NAND2_X2 _AES_ENC_U897  ( .A1(_AES_ENC_n553 ), .A2(_AES_ENC_n554 ), .ZN(_AES_ENC_N176 ) );
NAND2_X2 _AES_ENC_U896  ( .A1(_AES_ENC_sa21_next[3]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n550 ) );
XOR2_X2 _AES_ENC_U895  ( .A(_AES_ENC_w1[11] ), .B(_AES_ENC_text_in_r[75] ),.Z(_AES_ENC_n552 ) );
NAND2_X2 _AES_ENC_U894  ( .A1(_AES_ENC_n552 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n551 ) );
NAND2_X2 _AES_ENC_U893  ( .A1(_AES_ENC_n550 ), .A2(_AES_ENC_n551 ), .ZN(_AES_ENC_N177 ) );
NAND2_X2 _AES_ENC_U892  ( .A1(_AES_ENC_sa21_next[4]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n547 ) );
XOR2_X2 _AES_ENC_U891  ( .A(_AES_ENC_w1[12] ), .B(_AES_ENC_text_in_r[76] ),.Z(_AES_ENC_n549 ) );
NAND2_X2 _AES_ENC_U890  ( .A1(_AES_ENC_n549 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n548 ) );
NAND2_X2 _AES_ENC_U889  ( .A1(_AES_ENC_n547 ), .A2(_AES_ENC_n548 ), .ZN(_AES_ENC_N178 ) );
NAND2_X2 _AES_ENC_U888  ( .A1(_AES_ENC_sa21_next[5]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n544 ) );
XOR2_X2 _AES_ENC_U887  ( .A(_AES_ENC_w1[13] ), .B(_AES_ENC_text_in_r[77] ),.Z(_AES_ENC_n546 ) );
NAND2_X2 _AES_ENC_U886  ( .A1(_AES_ENC_n546 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n545 ) );
NAND2_X2 _AES_ENC_U885  ( .A1(_AES_ENC_n544 ), .A2(_AES_ENC_n545 ), .ZN(_AES_ENC_N179 ) );
NAND2_X2 _AES_ENC_U884  ( .A1(_AES_ENC_sa21_next[6]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n541 ) );
XOR2_X2 _AES_ENC_U883  ( .A(_AES_ENC_w1[14] ), .B(_AES_ENC_text_in_r[78] ),.Z(_AES_ENC_n543 ) );
NAND2_X2 _AES_ENC_U882  ( .A1(_AES_ENC_n543 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n542 ) );
NAND2_X2 _AES_ENC_U881  ( .A1(_AES_ENC_n541 ), .A2(_AES_ENC_n542 ), .ZN(_AES_ENC_N180 ) );
NAND2_X2 _AES_ENC_U880  ( .A1(_AES_ENC_sa21_next[7]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n538 ) );
XOR2_X2 _AES_ENC_U879  ( .A(_AES_ENC_w1[15] ), .B(_AES_ENC_text_in_r[79] ),.Z(_AES_ENC_n540 ) );
NAND2_X2 _AES_ENC_U878  ( .A1(_AES_ENC_n540 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n539 ) );
NAND2_X2 _AES_ENC_U877  ( .A1(_AES_ENC_n538 ), .A2(_AES_ENC_n539 ), .ZN(_AES_ENC_N181 ) );
AND4_X2 _AES_ENC_U875  ( .A1(_AES_ENC_n1232 ), .A2(_AES_ENC_n1259 ), .A3(_AES_ENC_n14 ), .A4(_AES_ENC_n792 ), .ZN(_AES_ENC_N19 ) );
NAND2_X2 _AES_ENC_U874  ( .A1(_AES_ENC_sa11_next[0]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n535 ) );
XOR2_X2 _AES_ENC_U873  ( .A(_AES_ENC_w1[16] ), .B(_AES_ENC_text_in_r[80] ),.Z(_AES_ENC_n537 ) );
NAND2_X2 _AES_ENC_U872  ( .A1(_AES_ENC_n537 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n536 ) );
NAND2_X2 _AES_ENC_U871  ( .A1(_AES_ENC_n535 ), .A2(_AES_ENC_n536 ), .ZN(_AES_ENC_N190 ) );
NAND2_X2 _AES_ENC_U870  ( .A1(_AES_ENC_sa11_next[1]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n532 ) );
XOR2_X2 _AES_ENC_U869  ( .A(_AES_ENC_w1[17] ), .B(_AES_ENC_text_in_r[81] ),.Z(_AES_ENC_n534 ) );
NAND2_X2 _AES_ENC_U868  ( .A1(_AES_ENC_n534 ), .A2(_AES_ENC_n1242 ), .ZN(_AES_ENC_n533 ) );
NAND2_X2 _AES_ENC_U867  ( .A1(_AES_ENC_n532 ), .A2(_AES_ENC_n533 ), .ZN(_AES_ENC_N191 ) );
NAND2_X2 _AES_ENC_U866  ( .A1(_AES_ENC_sa11_next[2]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n529 ) );
XOR2_X2 _AES_ENC_U865  ( .A(_AES_ENC_w1[18] ), .B(_AES_ENC_text_in_r[82] ),.Z(_AES_ENC_n531 ) );
NAND2_X2 _AES_ENC_U864  ( .A1(_AES_ENC_n531 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n5301 ) );
NAND2_X2 _AES_ENC_U863  ( .A1(_AES_ENC_n529 ), .A2(_AES_ENC_n5301 ), .ZN(_AES_ENC_N192 ) );
NAND2_X2 _AES_ENC_U862  ( .A1(_AES_ENC_sa11_next[3]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n526 ) );
XOR2_X2 _AES_ENC_U861  ( .A(_AES_ENC_w1[19] ), .B(_AES_ENC_text_in_r[83] ),.Z(_AES_ENC_n528 ) );
NAND2_X2 _AES_ENC_U860  ( .A1(_AES_ENC_n528 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n527 ) );
NAND2_X2 _AES_ENC_U859  ( .A1(_AES_ENC_n526 ), .A2(_AES_ENC_n527 ), .ZN(_AES_ENC_N193 ) );
NAND2_X2 _AES_ENC_U858  ( .A1(_AES_ENC_sa11_next[4]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n523 ) );
XOR2_X2 _AES_ENC_U857  ( .A(_AES_ENC_w1[20] ), .B(_AES_ENC_text_in_r[84] ),.Z(_AES_ENC_n525 ) );
NAND2_X2 _AES_ENC_U856  ( .A1(_AES_ENC_n525 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n524 ) );
NAND2_X2 _AES_ENC_U855  ( .A1(_AES_ENC_n523 ), .A2(_AES_ENC_n524 ), .ZN(_AES_ENC_N194 ) );
NAND2_X2 _AES_ENC_U854  ( .A1(_AES_ENC_sa11_next[5]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n5201 ) );
XOR2_X2 _AES_ENC_U853  ( .A(_AES_ENC_w1[21] ), .B(_AES_ENC_text_in_r[85] ),.Z(_AES_ENC_n522 ) );
NAND2_X2 _AES_ENC_U852  ( .A1(_AES_ENC_n522 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n521 ) );
NAND2_X2 _AES_ENC_U851  ( .A1(_AES_ENC_n5201 ), .A2(_AES_ENC_n521 ), .ZN(_AES_ENC_N195 ) );
NAND2_X2 _AES_ENC_U850  ( .A1(_AES_ENC_sa11_next[6]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n517 ) );
XOR2_X2 _AES_ENC_U849  ( .A(_AES_ENC_w1[22] ), .B(_AES_ENC_text_in_r[86] ),.Z(_AES_ENC_n519 ) );
NAND2_X2 _AES_ENC_U848  ( .A1(_AES_ENC_n519 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n518 ) );
NAND2_X2 _AES_ENC_U847  ( .A1(_AES_ENC_n517 ), .A2(_AES_ENC_n518 ), .ZN(_AES_ENC_N196 ) );
NAND2_X2 _AES_ENC_U846  ( .A1(_AES_ENC_sa11_next[7]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n514 ) );
XOR2_X2 _AES_ENC_U845  ( .A(_AES_ENC_w1[23] ), .B(_AES_ENC_text_in_r[87] ),.Z(_AES_ENC_n516 ) );
NAND2_X2 _AES_ENC_U844  ( .A1(_AES_ENC_n516 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n515 ) );
NAND2_X2 _AES_ENC_U843  ( .A1(_AES_ENC_n514 ), .A2(_AES_ENC_n515 ), .ZN(_AES_ENC_N197 ) );
NAND2_X2 _AES_ENC_U842  ( .A1(_AES_ENC_sa01_next[0]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n511 ) );
XOR2_X2 _AES_ENC_U841  ( .A(_AES_ENC_w1[24] ), .B(_AES_ENC_text_in_r[88] ),.Z(_AES_ENC_n513 ) );
NAND2_X2 _AES_ENC_U840  ( .A1(_AES_ENC_n513 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n512 ) );
NAND2_X2 _AES_ENC_U839  ( .A1(_AES_ENC_n511 ), .A2(_AES_ENC_n512 ), .ZN(_AES_ENC_N206 ) );
NAND2_X2 _AES_ENC_U838  ( .A1(_AES_ENC_sa01_next[1]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n508 ) );
XOR2_X2 _AES_ENC_U837  ( .A(_AES_ENC_w1[25] ), .B(_AES_ENC_text_in_r[89] ),.Z(_AES_ENC_n5101 ) );
NAND2_X2 _AES_ENC_U836  ( .A1(_AES_ENC_n5101 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n509 ) );
NAND2_X2 _AES_ENC_U835  ( .A1(_AES_ENC_n508 ), .A2(_AES_ENC_n509 ), .ZN(_AES_ENC_N207 ) );
NAND2_X2 _AES_ENC_U834  ( .A1(_AES_ENC_sa01_next[2]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n505 ) );
XOR2_X2 _AES_ENC_U833  ( .A(_AES_ENC_w1[26] ), .B(_AES_ENC_text_in_r[90] ),.Z(_AES_ENC_n507 ) );
NAND2_X2 _AES_ENC_U832  ( .A1(_AES_ENC_n507 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n506 ) );
NAND2_X2 _AES_ENC_U831  ( .A1(_AES_ENC_n505 ), .A2(_AES_ENC_n506 ), .ZN(_AES_ENC_N208 ) );
NAND2_X2 _AES_ENC_U830  ( .A1(_AES_ENC_sa01_next[3]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n5021 ) );
XOR2_X2 _AES_ENC_U829  ( .A(_AES_ENC_w1[27] ), .B(_AES_ENC_text_in_r[91] ),.Z(_AES_ENC_n504 ) );
NAND2_X2 _AES_ENC_U828  ( .A1(_AES_ENC_n504 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n503 ) );
NAND2_X2 _AES_ENC_U827  ( .A1(_AES_ENC_n5021 ), .A2(_AES_ENC_n503 ), .ZN(_AES_ENC_N209 ) );
NAND2_X2 _AES_ENC_U826  ( .A1(_AES_ENC_sa01_next[4]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4990 ) );
XOR2_X2 _AES_ENC_U825  ( .A(_AES_ENC_w1[28] ), .B(_AES_ENC_text_in_r[92] ),.Z(_AES_ENC_n5010 ) );
NAND2_X2 _AES_ENC_U824  ( .A1(_AES_ENC_n5010 ), .A2(_AES_ENC_n1243 ), .ZN(_AES_ENC_n5000 ) );
NAND2_X2 _AES_ENC_U823  ( .A1(_AES_ENC_n4990 ), .A2(_AES_ENC_n5000 ), .ZN(_AES_ENC_N210 ) );
NAND2_X2 _AES_ENC_U822  ( .A1(_AES_ENC_sa01_next[5]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4960 ) );
XOR2_X2 _AES_ENC_U821  ( .A(_AES_ENC_w1[29] ), .B(_AES_ENC_text_in_r[93] ),.Z(_AES_ENC_n4980 ) );
NAND2_X2 _AES_ENC_U820  ( .A1(_AES_ENC_n4980 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4970 ) );
NAND2_X2 _AES_ENC_U819  ( .A1(_AES_ENC_n4960 ), .A2(_AES_ENC_n4970 ), .ZN(_AES_ENC_N211 ) );
NAND2_X2 _AES_ENC_U818  ( .A1(_AES_ENC_sa01_next[6]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4930 ) );
XOR2_X2 _AES_ENC_U817  ( .A(_AES_ENC_w1[30] ), .B(_AES_ENC_text_in_r[94] ),.Z(_AES_ENC_n4950 ) );
NAND2_X2 _AES_ENC_U816  ( .A1(_AES_ENC_n4950 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4940 ) );
NAND2_X2 _AES_ENC_U815  ( .A1(_AES_ENC_n4930 ), .A2(_AES_ENC_n4940 ), .ZN(_AES_ENC_N212 ) );
NAND2_X2 _AES_ENC_U814  ( .A1(_AES_ENC_sa01_next[7]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4900 ) );
XOR2_X2 _AES_ENC_U813  ( .A(_AES_ENC_w1[31] ), .B(_AES_ENC_text_in_r[95] ),.Z(_AES_ENC_n4920 ) );
NAND2_X2 _AES_ENC_U812  ( .A1(_AES_ENC_n4920 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4911 ) );
NAND2_X2 _AES_ENC_U811  ( .A1(_AES_ENC_n4900 ), .A2(_AES_ENC_n4911 ), .ZN(_AES_ENC_N213 ) );
NAND2_X2 _AES_ENC_U810  ( .A1(_AES_ENC_sa30_next[0]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4870 ) );
XOR2_X2 _AES_ENC_U809  ( .A(_AES_ENC_w0[0] ), .B(_AES_ENC_text_in_r[96] ),.Z(_AES_ENC_n4890 ) );
NAND2_X2 _AES_ENC_U808  ( .A1(_AES_ENC_n4890 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4880 ) );
NAND2_X2 _AES_ENC_U807  ( .A1(_AES_ENC_n4870 ), .A2(_AES_ENC_n4880 ), .ZN(_AES_ENC_N222 ) );
NAND2_X2 _AES_ENC_U806  ( .A1(_AES_ENC_sa30_next[1]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4840 ) );
XOR2_X2 _AES_ENC_U805  ( .A(_AES_ENC_w0[1] ), .B(_AES_ENC_text_in_r[97] ),.Z(_AES_ENC_n4860 ) );
NAND2_X2 _AES_ENC_U804  ( .A1(_AES_ENC_n4860 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4850 ) );
NAND2_X2 _AES_ENC_U803  ( .A1(_AES_ENC_n4840 ), .A2(_AES_ENC_n4850 ), .ZN(_AES_ENC_N223 ) );
NAND2_X2 _AES_ENC_U802  ( .A1(_AES_ENC_sa30_next[2]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4811 ) );
XOR2_X2 _AES_ENC_U801  ( .A(_AES_ENC_w0[2] ), .B(_AES_ENC_text_in_r[98] ),.Z(_AES_ENC_n4830 ) );
NAND2_X2 _AES_ENC_U800  ( .A1(_AES_ENC_n4830 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4820 ) );
NAND2_X2 _AES_ENC_U799  ( .A1(_AES_ENC_n4811 ), .A2(_AES_ENC_n4820 ), .ZN(_AES_ENC_N224 ) );
NAND2_X2 _AES_ENC_U798  ( .A1(_AES_ENC_sa30_next[3]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4780 ) );
XOR2_X2 _AES_ENC_U797  ( .A(_AES_ENC_w0[3] ), .B(_AES_ENC_text_in_r[99] ),.Z(_AES_ENC_n4800 ) );
NAND2_X2 _AES_ENC_U796  ( .A1(_AES_ENC_n4800 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4790 ) );
NAND2_X2 _AES_ENC_U795  ( .A1(_AES_ENC_n4780 ), .A2(_AES_ENC_n4790 ), .ZN(_AES_ENC_N225 ) );
NAND2_X2 _AES_ENC_U794  ( .A1(_AES_ENC_sa30_next[4]), .A2(_AES_ENC_n1253 ),.ZN(_AES_ENC_n4750 ) );
XOR2_X2 _AES_ENC_U793  ( .A(_AES_ENC_w0[4] ), .B(_AES_ENC_text_in_r[100] ),.Z(_AES_ENC_n4770 ) );
NAND2_X2 _AES_ENC_U792  ( .A1(_AES_ENC_n4770 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4760 ) );
NAND2_X2 _AES_ENC_U791  ( .A1(_AES_ENC_n4750 ), .A2(_AES_ENC_n4760 ), .ZN(_AES_ENC_N226 ) );
NAND2_X2 _AES_ENC_U790  ( .A1(_AES_ENC_sa30_next[5]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4720 ) );
XOR2_X2 _AES_ENC_U789  ( .A(_AES_ENC_w0[5] ), .B(_AES_ENC_text_in_r[101] ),.Z(_AES_ENC_n4740 ) );
NAND2_X2 _AES_ENC_U788  ( .A1(_AES_ENC_n4740 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4730 ) );
NAND2_X2 _AES_ENC_U787  ( .A1(_AES_ENC_n4720 ), .A2(_AES_ENC_n4730 ), .ZN(_AES_ENC_N227 ) );
NAND2_X2 _AES_ENC_U786  ( .A1(_AES_ENC_sa30_next[6]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4690 ) );
XOR2_X2 _AES_ENC_U785  ( .A(_AES_ENC_w0[6] ), .B(_AES_ENC_text_in_r[102] ),.Z(_AES_ENC_n4711 ) );
NAND2_X2 _AES_ENC_U784  ( .A1(_AES_ENC_n4711 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4700 ) );
NAND2_X2 _AES_ENC_U783  ( .A1(_AES_ENC_n4690 ), .A2(_AES_ENC_n4700 ), .ZN(_AES_ENC_N228 ) );
NAND2_X2 _AES_ENC_U782  ( .A1(_AES_ENC_sa30_next[7]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4660 ) );
XOR2_X2 _AES_ENC_U781  ( .A(_AES_ENC_w0[7] ), .B(_AES_ENC_text_in_r[103] ),.Z(_AES_ENC_n4680 ) );
NAND2_X2 _AES_ENC_U780  ( .A1(_AES_ENC_n4680 ), .A2(_AES_ENC_n1244 ), .ZN(_AES_ENC_n4670 ) );
NAND2_X2 _AES_ENC_U779  ( .A1(_AES_ENC_n4660 ), .A2(_AES_ENC_n4670 ), .ZN(_AES_ENC_N229 ) );
NAND2_X2 _AES_ENC_U778  ( .A1(_AES_ENC_sa20_next[0]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4630 ) );
XOR2_X2 _AES_ENC_U777  ( .A(_AES_ENC_w0[8] ), .B(_AES_ENC_text_in_r[104] ),.Z(_AES_ENC_n4650 ) );
NAND2_X2 _AES_ENC_U776  ( .A1(_AES_ENC_n4650 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4640 ) );
NAND2_X2 _AES_ENC_U775  ( .A1(_AES_ENC_n4630 ), .A2(_AES_ENC_n4640 ), .ZN(_AES_ENC_N238 ) );
NAND2_X2 _AES_ENC_U774  ( .A1(_AES_ENC_sa20_next[1]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4600 ) );
XOR2_X2 _AES_ENC_U773  ( .A(_AES_ENC_w0[9] ), .B(_AES_ENC_text_in_r[105] ),.Z(_AES_ENC_n4620 ) );
NAND2_X2 _AES_ENC_U772  ( .A1(_AES_ENC_n4620 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4611 ) );
NAND2_X2 _AES_ENC_U771  ( .A1(_AES_ENC_n4600 ), .A2(_AES_ENC_n4611 ), .ZN(_AES_ENC_N239 ) );
NAND2_X2 _AES_ENC_U770  ( .A1(_AES_ENC_sa20_next[2]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4570 ) );
XOR2_X2 _AES_ENC_U769  ( .A(_AES_ENC_w0[10] ), .B(_AES_ENC_text_in_r[106] ),.Z(_AES_ENC_n4590 ) );
NAND2_X2 _AES_ENC_U768  ( .A1(_AES_ENC_n4590 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4580 ) );
NAND2_X2 _AES_ENC_U767  ( .A1(_AES_ENC_n4570 ), .A2(_AES_ENC_n4580 ), .ZN(_AES_ENC_N240 ) );
NAND2_X2 _AES_ENC_U766  ( .A1(_AES_ENC_sa20_next[3]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4540 ) );
XOR2_X2 _AES_ENC_U765  ( .A(_AES_ENC_w0[11] ), .B(_AES_ENC_text_in_r[107] ),.Z(_AES_ENC_n4560 ) );
NAND2_X2 _AES_ENC_U764  ( .A1(_AES_ENC_n4560 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4550 ) );
NAND2_X2 _AES_ENC_U763  ( .A1(_AES_ENC_n4540 ), .A2(_AES_ENC_n4550 ), .ZN(_AES_ENC_N241 ) );
NAND2_X2 _AES_ENC_U762  ( .A1(_AES_ENC_sa20_next[4]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4510 ) );
XOR2_X2 _AES_ENC_U761  ( .A(_AES_ENC_w0[12] ), .B(_AES_ENC_text_in_r[108] ),.Z(_AES_ENC_n4530 ) );
NAND2_X2 _AES_ENC_U760  ( .A1(_AES_ENC_n4530 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4520 ) );
NAND2_X2 _AES_ENC_U759  ( .A1(_AES_ENC_n4510 ), .A2(_AES_ENC_n4520 ), .ZN(_AES_ENC_N242 ) );
NAND2_X2 _AES_ENC_U758  ( .A1(_AES_ENC_sa20_next[5]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4480 ) );
XOR2_X2 _AES_ENC_U757  ( .A(_AES_ENC_w0[13] ), .B(_AES_ENC_text_in_r[109] ),.Z(_AES_ENC_n4500 ) );
NAND2_X2 _AES_ENC_U756  ( .A1(_AES_ENC_n4500 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4490 ) );
NAND2_X2 _AES_ENC_U755  ( .A1(_AES_ENC_n4480 ), .A2(_AES_ENC_n4490 ), .ZN(_AES_ENC_N243 ) );
NAND2_X2 _AES_ENC_U754  ( .A1(_AES_ENC_sa20_next[6]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4450 ) );
XOR2_X2 _AES_ENC_U753  ( .A(_AES_ENC_w0[14] ), .B(_AES_ENC_text_in_r[110] ),.Z(_AES_ENC_n4470 ) );
NAND2_X2 _AES_ENC_U752  ( .A1(_AES_ENC_n4470 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4460 ) );
NAND2_X2 _AES_ENC_U751  ( .A1(_AES_ENC_n4450 ), .A2(_AES_ENC_n4460 ), .ZN(_AES_ENC_N244 ) );
NAND2_X2 _AES_ENC_U750  ( .A1(_AES_ENC_sa20_next[7]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4420 ) );
XOR2_X2 _AES_ENC_U749  ( .A(_AES_ENC_w0[15] ), .B(_AES_ENC_text_in_r[111] ),.Z(_AES_ENC_n4440 ) );
NAND2_X2 _AES_ENC_U748  ( .A1(_AES_ENC_n4440 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4430 ) );
NAND2_X2 _AES_ENC_U747  ( .A1(_AES_ENC_n4420 ), .A2(_AES_ENC_n4430 ), .ZN(_AES_ENC_N245 ) );
NAND2_X2 _AES_ENC_U746  ( .A1(_AES_ENC_sa10_next[0]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4390 ) );
XOR2_X2 _AES_ENC_U745  ( .A(_AES_ENC_w0[16] ), .B(_AES_ENC_text_in_r[112] ),.Z(_AES_ENC_n4410 ) );
NAND2_X2 _AES_ENC_U744  ( .A1(_AES_ENC_n4410 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4400 ) );
NAND2_X2 _AES_ENC_U743  ( .A1(_AES_ENC_n4390 ), .A2(_AES_ENC_n4400 ), .ZN(_AES_ENC_N254 ) );
NAND2_X2 _AES_ENC_U742  ( .A1(_AES_ENC_sa10_next[1]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4360 ) );
XOR2_X2 _AES_ENC_U741  ( .A(_AES_ENC_w0[17] ), .B(_AES_ENC_text_in_r[113] ),.Z(_AES_ENC_n4380 ) );
NAND2_X2 _AES_ENC_U740  ( .A1(_AES_ENC_n4380 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4370 ) );
NAND2_X2 _AES_ENC_U739  ( .A1(_AES_ENC_n4360 ), .A2(_AES_ENC_n4370 ), .ZN(_AES_ENC_N255 ) );
NAND2_X2 _AES_ENC_U738  ( .A1(_AES_ENC_sa10_next[2]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4330 ) );
XOR2_X2 _AES_ENC_U737  ( .A(_AES_ENC_w0[18] ), .B(_AES_ENC_text_in_r[114] ),.Z(_AES_ENC_n4350 ) );
NAND2_X2 _AES_ENC_U736  ( .A1(_AES_ENC_n4350 ), .A2(_AES_ENC_n1245 ), .ZN(_AES_ENC_n4340 ) );
NAND2_X2 _AES_ENC_U735  ( .A1(_AES_ENC_n4330 ), .A2(_AES_ENC_n4340 ), .ZN(_AES_ENC_N256 ) );
NAND2_X2 _AES_ENC_U734  ( .A1(_AES_ENC_sa10_next[3]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4300 ) );
XOR2_X2 _AES_ENC_U733  ( .A(_AES_ENC_w0[19] ), .B(_AES_ENC_text_in_r[115] ),.Z(_AES_ENC_n4320 ) );
NAND2_X2 _AES_ENC_U732  ( .A1(_AES_ENC_n4320 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4310 ) );
NAND2_X2 _AES_ENC_U731  ( .A1(_AES_ENC_n4300 ), .A2(_AES_ENC_n4310 ), .ZN(_AES_ENC_N257 ) );
NAND2_X2 _AES_ENC_U730  ( .A1(_AES_ENC_sa10_next[4]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4270 ) );
XOR2_X2 _AES_ENC_U729  ( .A(_AES_ENC_w0[20] ), .B(_AES_ENC_text_in_r[116] ),.Z(_AES_ENC_n4290 ) );
NAND2_X2 _AES_ENC_U728  ( .A1(_AES_ENC_n4290 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4280 ) );
NAND2_X2 _AES_ENC_U727  ( .A1(_AES_ENC_n4270 ), .A2(_AES_ENC_n4280 ), .ZN(_AES_ENC_N258 ) );
NAND2_X2 _AES_ENC_U726  ( .A1(_AES_ENC_sa10_next[5]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4240 ) );
XOR2_X2 _AES_ENC_U725  ( .A(_AES_ENC_w0[21] ), .B(_AES_ENC_text_in_r[117] ),.Z(_AES_ENC_n4260 ) );
NAND2_X2 _AES_ENC_U724  ( .A1(_AES_ENC_n4260 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4250 ) );
NAND2_X2 _AES_ENC_U723  ( .A1(_AES_ENC_n4240 ), .A2(_AES_ENC_n4250 ), .ZN(_AES_ENC_N259 ) );
NAND2_X2 _AES_ENC_U722  ( .A1(_AES_ENC_sa10_next[6]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4210 ) );
XOR2_X2 _AES_ENC_U721  ( .A(_AES_ENC_w0[22] ), .B(_AES_ENC_text_in_r[118] ),.Z(_AES_ENC_n4230 ) );
NAND2_X2 _AES_ENC_U720  ( .A1(_AES_ENC_n4230 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4220 ) );
NAND2_X2 _AES_ENC_U719  ( .A1(_AES_ENC_n4210 ), .A2(_AES_ENC_n4220 ), .ZN(_AES_ENC_N260 ) );
NAND2_X2 _AES_ENC_U718  ( .A1(_AES_ENC_sa10_next[7]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4180 ) );
XOR2_X2 _AES_ENC_U717  ( .A(_AES_ENC_w0[23] ), .B(_AES_ENC_text_in_r[119] ),.Z(_AES_ENC_n4200 ) );
NAND2_X2 _AES_ENC_U716  ( .A1(_AES_ENC_n4200 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4190 ) );
NAND2_X2 _AES_ENC_U715  ( .A1(_AES_ENC_n4180 ), .A2(_AES_ENC_n4190 ), .ZN(_AES_ENC_N261 ) );
NAND2_X2 _AES_ENC_U714  ( .A1(_AES_ENC_sa00_next[0]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4150 ) );
XOR2_X2 _AES_ENC_U713  ( .A(_AES_ENC_w0[24] ), .B(_AES_ENC_text_in_r[120] ),.Z(_AES_ENC_n4170 ) );
NAND2_X2 _AES_ENC_U712  ( .A1(_AES_ENC_n4170 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4160 ) );
NAND2_X2 _AES_ENC_U711  ( .A1(_AES_ENC_n4150 ), .A2(_AES_ENC_n4160 ), .ZN(_AES_ENC_N270 ) );
NAND2_X2 _AES_ENC_U710  ( .A1(_AES_ENC_sa00_next[1]), .A2(_AES_ENC_n1254 ),.ZN(_AES_ENC_n4120 ) );
XOR2_X2 _AES_ENC_U709  ( .A(_AES_ENC_w0[25] ), .B(_AES_ENC_text_in_r[121] ),.Z(_AES_ENC_n4140 ) );
NAND2_X2 _AES_ENC_U708  ( .A1(_AES_ENC_n4140 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4130 ) );
NAND2_X2 _AES_ENC_U707  ( .A1(_AES_ENC_n4120 ), .A2(_AES_ENC_n4130 ), .ZN(_AES_ENC_N271 ) );
NAND2_X2 _AES_ENC_U706  ( .A1(_AES_ENC_sa00_next[2]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n4090 ) );
XOR2_X2 _AES_ENC_U705  ( .A(_AES_ENC_w0[26] ), .B(_AES_ENC_text_in_r[122] ),.Z(_AES_ENC_n4110 ) );
NAND2_X2 _AES_ENC_U704  ( .A1(_AES_ENC_n4110 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4100 ) );
NAND2_X2 _AES_ENC_U703  ( .A1(_AES_ENC_n4090 ), .A2(_AES_ENC_n4100 ), .ZN(_AES_ENC_N272 ) );
NAND2_X2 _AES_ENC_U702  ( .A1(_AES_ENC_sa00_next[3]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n4060 ) );
XOR2_X2 _AES_ENC_U701  ( .A(_AES_ENC_w0[27] ), .B(_AES_ENC_text_in_r[123] ),.Z(_AES_ENC_n4080 ) );
NAND2_X2 _AES_ENC_U700  ( .A1(_AES_ENC_n4080 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4070 ) );
NAND2_X2 _AES_ENC_U699  ( .A1(_AES_ENC_n4060 ), .A2(_AES_ENC_n4070 ), .ZN(_AES_ENC_N273 ) );
NAND2_X2 _AES_ENC_U698  ( .A1(_AES_ENC_sa00_next[4]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n4030 ) );
XOR2_X2 _AES_ENC_U697  ( .A(_AES_ENC_w0[28] ), .B(_AES_ENC_text_in_r[124] ),.Z(_AES_ENC_n4050 ) );
NAND2_X2 _AES_ENC_U696  ( .A1(_AES_ENC_n4050 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4040 ) );
NAND2_X2 _AES_ENC_U695  ( .A1(_AES_ENC_n4030 ), .A2(_AES_ENC_n4040 ), .ZN(_AES_ENC_N274 ) );
NAND2_X2 _AES_ENC_U694  ( .A1(_AES_ENC_sa00_next[5]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n4000 ) );
XOR2_X2 _AES_ENC_U693  ( .A(_AES_ENC_w0[29] ), .B(_AES_ENC_text_in_r[125] ),.Z(_AES_ENC_n4020 ) );
NAND2_X2 _AES_ENC_U692  ( .A1(_AES_ENC_n4020 ), .A2(_AES_ENC_n1246 ), .ZN(_AES_ENC_n4010 ) );
NAND2_X2 _AES_ENC_U691  ( .A1(_AES_ENC_n4000 ), .A2(_AES_ENC_n4010 ), .ZN(_AES_ENC_N275 ) );
NAND2_X2 _AES_ENC_U690  ( .A1(_AES_ENC_sa00_next[6]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3970 ) );
XOR2_X2 _AES_ENC_U689  ( .A(_AES_ENC_w0[30] ), .B(_AES_ENC_text_in_r[126] ),.Z(_AES_ENC_n3990 ) );
NAND2_X2 _AES_ENC_U688  ( .A1(_AES_ENC_n3990 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3980 ) );
NAND2_X2 _AES_ENC_U687  ( .A1(_AES_ENC_n3970 ), .A2(_AES_ENC_n3980 ), .ZN(_AES_ENC_N276 ) );
NAND2_X2 _AES_ENC_U686  ( .A1(_AES_ENC_sa00_next[7]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3940 ) );
XOR2_X2 _AES_ENC_U685  ( .A(_AES_ENC_w0[31] ), .B(_AES_ENC_text_in_r[127] ),.Z(_AES_ENC_n3960 ) );
NAND2_X2 _AES_ENC_U684  ( .A1(_AES_ENC_n3960 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3950 ) );
NAND2_X2 _AES_ENC_U683  ( .A1(_AES_ENC_n3940 ), .A2(_AES_ENC_n3950 ), .ZN(_AES_ENC_N277 ) );
NAND2_X2 _AES_ENC_U682  ( .A1(__AES_ENC_sa33_next[0]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3910 ) );
XOR2_X2 _AES_ENC_U681  ( .A(_AES_ENC_w3[0] ), .B(_AES_ENC_text_in_r[0] ),.Z(_AES_ENC_n3930 ) );
NAND2_X2 _AES_ENC_U680  ( .A1(_AES_ENC_n3930 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3920 ) );
NAND2_X2 _AES_ENC_U679  ( .A1(_AES_ENC_n3910 ), .A2(_AES_ENC_n3920 ), .ZN(_AES_ENC_N30 ) );
NAND2_X2 _AES_ENC_U678  ( .A1(__AES_ENC_sa33_next[1]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3880 ) );
XOR2_X2 _AES_ENC_U677  ( .A(_AES_ENC_w3[1] ), .B(_AES_ENC_text_in_r[1] ),.Z(_AES_ENC_n3900 ) );
NAND2_X2 _AES_ENC_U676  ( .A1(_AES_ENC_n3900 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3890 ) );
NAND2_X2 _AES_ENC_U675  ( .A1(_AES_ENC_n3880 ), .A2(_AES_ENC_n3890 ), .ZN(_AES_ENC_N31 ) );
NAND2_X2 _AES_ENC_U674  ( .A1(__AES_ENC_sa33_next[2]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3850 ) );
XOR2_X2 _AES_ENC_U673  ( .A(_AES_ENC_w3[2] ), .B(_AES_ENC_text_in_r[2] ),.Z(_AES_ENC_n3870 ) );
NAND2_X2 _AES_ENC_U672  ( .A1(_AES_ENC_n3870 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3860 ) );
NAND2_X2 _AES_ENC_U671  ( .A1(_AES_ENC_n3850 ), .A2(_AES_ENC_n3860 ), .ZN(_AES_ENC_N32 ) );
NAND2_X2 _AES_ENC_U670  ( .A1(__AES_ENC_sa33_next[3]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3820 ) );
XOR2_X2 _AES_ENC_U669  ( .A(_AES_ENC_w3[3] ), .B(_AES_ENC_text_in_r[3] ),.Z(_AES_ENC_n3840 ) );
NAND2_X2 _AES_ENC_U668  ( .A1(_AES_ENC_n3840 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3830 ) );
NAND2_X2 _AES_ENC_U667  ( .A1(_AES_ENC_n3820 ), .A2(_AES_ENC_n3830 ), .ZN(_AES_ENC_N33 ) );
NAND2_X2 _AES_ENC_U666  ( .A1(__AES_ENC_sa33_next[4]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3790 ) );
XOR2_X2 _AES_ENC_U665  ( .A(_AES_ENC_w3[4] ), .B(_AES_ENC_text_in_r[4] ),.Z(_AES_ENC_n3810 ) );
NAND2_X2 _AES_ENC_U664  ( .A1(_AES_ENC_n3810 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3800 ) );
NAND2_X2 _AES_ENC_U663  ( .A1(_AES_ENC_n3790 ), .A2(_AES_ENC_n3800 ), .ZN(_AES_ENC_N34 ) );
NAND2_X2 _AES_ENC_U662  ( .A1(__AES_ENC_sa33_next[5]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3760 ) );
XOR2_X2 _AES_ENC_U661  ( .A(_AES_ENC_w3[5] ), .B(_AES_ENC_text_in_r[5] ),.Z(_AES_ENC_n3780 ) );
NAND2_X2 _AES_ENC_U660  ( .A1(_AES_ENC_n3780 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3770 ) );
NAND2_X2 _AES_ENC_U659  ( .A1(_AES_ENC_n3760 ), .A2(_AES_ENC_n3770 ), .ZN(_AES_ENC_N35 ) );
NAND2_X2 _AES_ENC_U658  ( .A1(__AES_ENC_sa33_next[6]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n373 ) );
XOR2_X2 _AES_ENC_U657  ( .A(_AES_ENC_w3[6] ), .B(_AES_ENC_text_in_r[6] ),.Z(_AES_ENC_n3750 ) );
NAND2_X2 _AES_ENC_U656  ( .A1(_AES_ENC_n3750 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n3740 ) );
NAND2_X2 _AES_ENC_U655  ( .A1(_AES_ENC_n373 ), .A2(_AES_ENC_n3740 ), .ZN(_AES_ENC_N36 ) );
NAND2_X2 _AES_ENC_U654  ( .A1(__AES_ENC_sa33_next[7]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n3701 ) );
XOR2_X2 _AES_ENC_U653  ( .A(_AES_ENC_w3[7] ), .B(_AES_ENC_text_in_r[7] ),.Z(_AES_ENC_n372 ) );
NAND2_X2 _AES_ENC_U652  ( .A1(_AES_ENC_n372 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n371 ) );
NAND2_X2 _AES_ENC_U651  ( .A1(_AES_ENC_n3701 ), .A2(_AES_ENC_n371 ), .ZN(_AES_ENC_N37 ) );
XOR2_X2 _AES_ENC_U650  ( .A(_AES_ENC_w0[31] ), .B(_AES_ENC_sa00_sub[7] ),.Z(_AES_ENC_N374 ) );
XOR2_X2 _AES_ENC_U649  ( .A(_AES_ENC_w0[30] ), .B(_AES_ENC_sa00_sub[6] ),.Z(_AES_ENC_N375 ) );
XOR2_X2 _AES_ENC_U648  ( .A(_AES_ENC_w0[29] ), .B(_AES_ENC_sa00_sub[5] ),.Z(_AES_ENC_N376 ) );
XOR2_X2 _AES_ENC_U647  ( .A(_AES_ENC_w0[28] ), .B(_AES_ENC_sa00_sub[4] ),.Z(_AES_ENC_N377 ) );
XOR2_X2 _AES_ENC_U646  ( .A(_AES_ENC_w0[27] ), .B(_AES_ENC_sa00_sub[3] ),.Z(_AES_ENC_N378 ) );
XOR2_X2 _AES_ENC_U645  ( .A(_AES_ENC_w0[26] ), .B(_AES_ENC_sa00_sub[2] ),.Z(_AES_ENC_N379 ) );
XOR2_X2 _AES_ENC_U644  ( .A(_AES_ENC_w0[25] ), .B(_AES_ENC_sa00_sub[1] ),.Z(_AES_ENC_N380 ) );
XOR2_X2 _AES_ENC_U643  ( .A(_AES_ENC_w0[24] ), .B(_AES_ENC_sa00_sub[0] ),.Z(_AES_ENC_N381 ) );
XOR2_X2 _AES_ENC_U642  ( .A(_AES_ENC_w1[31] ), .B(_AES_ENC_sa01_sub[7] ),.Z(_AES_ENC_N382 ) );
XOR2_X2 _AES_ENC_U641  ( .A(_AES_ENC_w1[30] ), .B(_AES_ENC_sa01_sub[6] ),.Z(_AES_ENC_N383 ) );
XOR2_X2 _AES_ENC_U640  ( .A(_AES_ENC_w1[29] ), .B(_AES_ENC_sa01_sub[5] ),.Z(_AES_ENC_N384 ) );
XOR2_X2 _AES_ENC_U639  ( .A(_AES_ENC_w1[28] ), .B(_AES_ENC_sa01_sub[4] ),.Z(_AES_ENC_N385 ) );
XOR2_X2 _AES_ENC_U638  ( .A(_AES_ENC_w1[27] ), .B(_AES_ENC_sa01_sub[3] ),.Z(_AES_ENC_N386 ) );
XOR2_X2 _AES_ENC_U637  ( .A(_AES_ENC_w1[26] ), .B(_AES_ENC_sa01_sub[2] ),.Z(_AES_ENC_N387 ) );
XOR2_X2 _AES_ENC_U636  ( .A(_AES_ENC_w1[25] ), .B(_AES_ENC_sa01_sub[1] ),.Z(_AES_ENC_N388 ) );
XOR2_X2 _AES_ENC_U635  ( .A(_AES_ENC_w1[24] ), .B(_AES_ENC_sa01_sub[0] ),.Z(_AES_ENC_N389 ) );
XOR2_X2 _AES_ENC_U634  ( .A(_AES_ENC_w2[31] ), .B(_AES_ENC_sa02_sub[7] ),.Z(_AES_ENC_N390 ) );
XOR2_X2 _AES_ENC_U633  ( .A(_AES_ENC_w2[30] ), .B(_AES_ENC_sa02_sub[6] ),.Z(_AES_ENC_N391 ) );
XOR2_X2 _AES_ENC_U632  ( .A(_AES_ENC_w2[29] ), .B(_AES_ENC_sa02_sub[5] ),.Z(_AES_ENC_N392 ) );
XOR2_X2 _AES_ENC_U631  ( .A(_AES_ENC_w2[28] ), .B(_AES_ENC_sa02_sub[4] ),.Z(_AES_ENC_N393 ) );
XOR2_X2 _AES_ENC_U630  ( .A(_AES_ENC_w2[27] ), .B(_AES_ENC_sa02_sub[3] ),.Z(_AES_ENC_N394 ) );
XOR2_X2 _AES_ENC_U629  ( .A(_AES_ENC_w2[26] ), .B(_AES_ENC_sa02_sub[2] ),.Z(_AES_ENC_N395 ) );
XOR2_X2 _AES_ENC_U628  ( .A(_AES_ENC_w2[25] ), .B(_AES_ENC_sa02_sub[1] ),.Z(_AES_ENC_N396 ) );
XOR2_X2 _AES_ENC_U627  ( .A(_AES_ENC_w2[24] ), .B(_AES_ENC_sa02_sub[0] ),.Z(_AES_ENC_N397 ) );
XOR2_X2 _AES_ENC_U626  ( .A(_AES_ENC_w3[31] ), .B(_AES_ENC_sa03_sub[7] ),.Z(_AES_ENC_N398 ) );
XOR2_X2 _AES_ENC_U625  ( .A(_AES_ENC_w3[30] ), .B(_AES_ENC_sa03_sub[6] ),.Z(_AES_ENC_N399 ) );
XOR2_X2 _AES_ENC_U624  ( .A(_AES_ENC_w3[29] ), .B(_AES_ENC_sa03_sub[5] ),.Z(_AES_ENC_N400 ) );
XOR2_X2 _AES_ENC_U623  ( .A(_AES_ENC_w3[28] ), .B(_AES_ENC_sa03_sub[4] ),.Z(_AES_ENC_N401 ) );
XOR2_X2 _AES_ENC_U622  ( .A(_AES_ENC_w3[27] ), .B(_AES_ENC_sa03_sub[3] ),.Z(_AES_ENC_N402 ) );
XOR2_X2 _AES_ENC_U621  ( .A(_AES_ENC_w3[26] ), .B(_AES_ENC_sa03_sub[2] ),.Z(_AES_ENC_N403 ) );
XOR2_X2 _AES_ENC_U620  ( .A(_AES_ENC_w3[25] ), .B(_AES_ENC_sa03_sub[1] ),.Z(_AES_ENC_N404 ) );
XOR2_X2 _AES_ENC_U619  ( .A(_AES_ENC_w3[24] ), .B(_AES_ENC_sa03_sub[0] ),.Z(_AES_ENC_N405 ) );
XOR2_X2 _AES_ENC_U618  ( .A(_AES_ENC_w0[23] ), .B(_AES_ENC_sa11_sub[7] ),.Z(_AES_ENC_N406 ) );
XOR2_X2 _AES_ENC_U617  ( .A(_AES_ENC_w0[22] ), .B(_AES_ENC_sa11_sub[6] ),.Z(_AES_ENC_N407 ) );
XOR2_X2 _AES_ENC_U616  ( .A(_AES_ENC_w0[21] ), .B(_AES_ENC_sa11_sub[5] ),.Z(_AES_ENC_N408 ) );
XOR2_X2 _AES_ENC_U615  ( .A(_AES_ENC_w0[20] ), .B(_AES_ENC_sa11_sub[4] ),.Z(_AES_ENC_N409 ) );
XOR2_X2 _AES_ENC_U614  ( .A(_AES_ENC_w0[19] ), .B(_AES_ENC_sa11_sub[3] ),.Z(_AES_ENC_N410 ) );
XOR2_X2 _AES_ENC_U613  ( .A(_AES_ENC_w0[18] ), .B(_AES_ENC_sa11_sub[2] ),.Z(_AES_ENC_N411 ) );
XOR2_X2 _AES_ENC_U612  ( .A(_AES_ENC_w0[17] ), .B(_AES_ENC_sa11_sub[1] ),.Z(_AES_ENC_N412 ) );
XOR2_X2 _AES_ENC_U611  ( .A(_AES_ENC_w0[16] ), .B(_AES_ENC_sa11_sub[0] ),.Z(_AES_ENC_N413 ) );
XOR2_X2 _AES_ENC_U610  ( .A(_AES_ENC_w1[23] ), .B(_AES_ENC_sa12_sub[7] ),.Z(_AES_ENC_N414 ) );
XOR2_X2 _AES_ENC_U609  ( .A(_AES_ENC_w1[22] ), .B(_AES_ENC_sa12_sub[6] ),.Z(_AES_ENC_N415 ) );
XOR2_X2 _AES_ENC_U608  ( .A(_AES_ENC_w1[21] ), .B(_AES_ENC_sa12_sub[5] ),.Z(_AES_ENC_N416 ) );
XOR2_X2 _AES_ENC_U607  ( .A(_AES_ENC_w1[20] ), .B(_AES_ENC_sa12_sub[4] ),.Z(_AES_ENC_N417 ) );
XOR2_X2 _AES_ENC_U606  ( .A(_AES_ENC_w1[19] ), .B(_AES_ENC_sa12_sub[3] ),.Z(_AES_ENC_N418 ) );
XOR2_X2 _AES_ENC_U605  ( .A(_AES_ENC_w1[18] ), .B(_AES_ENC_sa12_sub[2] ),.Z(_AES_ENC_N419 ) );
XOR2_X2 _AES_ENC_U604  ( .A(_AES_ENC_w1[17] ), .B(_AES_ENC_sa12_sub[1] ),.Z(_AES_ENC_N420 ) );
XOR2_X2 _AES_ENC_U603  ( .A(_AES_ENC_w1[16] ), .B(_AES_ENC_sa12_sub[0] ),.Z(_AES_ENC_N421 ) );
XOR2_X2 _AES_ENC_U602  ( .A(_AES_ENC_w2[23] ), .B(_AES_ENC_sa13_sub[7] ),.Z(_AES_ENC_N422 ) );
XOR2_X2 _AES_ENC_U601  ( .A(_AES_ENC_w2[22] ), .B(_AES_ENC_sa13_sub[6] ),.Z(_AES_ENC_N423 ) );
XOR2_X2 _AES_ENC_U600  ( .A(_AES_ENC_w2[21] ), .B(_AES_ENC_sa13_sub[5] ),.Z(_AES_ENC_N424 ) );
XOR2_X2 _AES_ENC_U599  ( .A(_AES_ENC_w2[20] ), .B(_AES_ENC_sa13_sub[4] ),.Z(_AES_ENC_N425 ) );
XOR2_X2 _AES_ENC_U598  ( .A(_AES_ENC_w2[19] ), .B(_AES_ENC_sa13_sub[3] ),.Z(_AES_ENC_N426 ) );
XOR2_X2 _AES_ENC_U597  ( .A(_AES_ENC_w2[18] ), .B(_AES_ENC_sa13_sub[2] ),.Z(_AES_ENC_N427 ) );
XOR2_X2 _AES_ENC_U596  ( .A(_AES_ENC_w2[17] ), .B(_AES_ENC_sa13_sub[1] ),.Z(_AES_ENC_N428 ) );
XOR2_X2 _AES_ENC_U595  ( .A(_AES_ENC_w2[16] ), .B(_AES_ENC_sa13_sub[0] ),.Z(_AES_ENC_N429 ) );
XOR2_X2 _AES_ENC_U594  ( .A(_AES_ENC_w3[23] ), .B(_AES_ENC_sa10_sub[7] ),.Z(_AES_ENC_N430 ) );
XOR2_X2 _AES_ENC_U593  ( .A(_AES_ENC_w3[22] ), .B(_AES_ENC_sa10_sub[6] ),.Z(_AES_ENC_N431 ) );
XOR2_X2 _AES_ENC_U592  ( .A(_AES_ENC_w3[21] ), .B(_AES_ENC_sa10_sub[5] ),.Z(_AES_ENC_N432 ) );
XOR2_X2 _AES_ENC_U591  ( .A(_AES_ENC_w3[20] ), .B(_AES_ENC_sa10_sub[4] ),.Z(_AES_ENC_N433 ) );
XOR2_X2 _AES_ENC_U590  ( .A(_AES_ENC_w3[19] ), .B(_AES_ENC_sa10_sub[3] ),.Z(_AES_ENC_N434 ) );
XOR2_X2 _AES_ENC_U589  ( .A(_AES_ENC_w3[18] ), .B(_AES_ENC_sa10_sub[2] ),.Z(_AES_ENC_N435 ) );
XOR2_X2 _AES_ENC_U588  ( .A(_AES_ENC_w3[17] ), .B(_AES_ENC_sa10_sub[1] ),.Z(_AES_ENC_N436 ) );
XOR2_X2 _AES_ENC_U587  ( .A(_AES_ENC_w3[16] ), .B(_AES_ENC_sa10_sub[0] ),.Z(_AES_ENC_N437 ) );
XOR2_X2 _AES_ENC_U586  ( .A(_AES_ENC_w0[15] ), .B(_AES_ENC_sa22_sub[7] ),.Z(_AES_ENC_N438 ) );
XOR2_X2 _AES_ENC_U585  ( .A(_AES_ENC_w0[14] ), .B(_AES_ENC_sa22_sub[6] ),.Z(_AES_ENC_N439 ) );
XOR2_X2 _AES_ENC_U584  ( .A(_AES_ENC_w0[13] ), .B(_AES_ENC_sa22_sub[5] ),.Z(_AES_ENC_N440 ) );
XOR2_X2 _AES_ENC_U583  ( .A(_AES_ENC_w0[12] ), .B(_AES_ENC_sa22_sub[4] ),.Z(_AES_ENC_N441 ) );
XOR2_X2 _AES_ENC_U582  ( .A(_AES_ENC_w0[11] ), .B(_AES_ENC_sa22_sub[3] ),.Z(_AES_ENC_N442 ) );
XOR2_X2 _AES_ENC_U581  ( .A(_AES_ENC_w0[10] ), .B(_AES_ENC_sa22_sub[2] ),.Z(_AES_ENC_N443 ) );
XOR2_X2 _AES_ENC_U580  ( .A(_AES_ENC_w0[9] ), .B(_AES_ENC_sa22_sub[1] ), .Z(_AES_ENC_N444 ) );
XOR2_X2 _AES_ENC_U579  ( .A(_AES_ENC_w0[8] ), .B(_AES_ENC_sa22_sub[0] ), .Z(_AES_ENC_N445 ) );
XOR2_X2 _AES_ENC_U578  ( .A(_AES_ENC_w1[15] ), .B(_AES_ENC_sa23_sub[7] ),.Z(_AES_ENC_N446 ) );
XOR2_X2 _AES_ENC_U577  ( .A(_AES_ENC_w1[14] ), .B(_AES_ENC_sa23_sub[6] ),.Z(_AES_ENC_N447 ) );
XOR2_X2 _AES_ENC_U576  ( .A(_AES_ENC_w1[13] ), .B(_AES_ENC_sa23_sub[5] ),.Z(_AES_ENC_N448 ) );
XOR2_X2 _AES_ENC_U575  ( .A(_AES_ENC_w1[12] ), .B(_AES_ENC_sa23_sub[4] ),.Z(_AES_ENC_N449 ) );
XOR2_X2 _AES_ENC_U574  ( .A(_AES_ENC_w1[11] ), .B(_AES_ENC_sa23_sub[3] ),.Z(_AES_ENC_N450 ) );
XOR2_X2 _AES_ENC_U573  ( .A(_AES_ENC_w1[10] ), .B(_AES_ENC_sa23_sub[2] ),.Z(_AES_ENC_N451 ) );
XOR2_X2 _AES_ENC_U572  ( .A(_AES_ENC_w1[9] ), .B(_AES_ENC_sa23_sub[1] ), .Z(_AES_ENC_N452 ) );
XOR2_X2 _AES_ENC_U571  ( .A(_AES_ENC_w1[8] ), .B(_AES_ENC_sa23_sub[0] ), .Z(_AES_ENC_N453 ) );
XOR2_X2 _AES_ENC_U570  ( .A(_AES_ENC_w2[15] ), .B(_AES_ENC_sa20_sub[7] ),.Z(_AES_ENC_N454 ) );
XOR2_X2 _AES_ENC_U569  ( .A(_AES_ENC_w2[14] ), .B(_AES_ENC_sa20_sub[6] ),.Z(_AES_ENC_N455 ) );
XOR2_X2 _AES_ENC_U568  ( .A(_AES_ENC_w2[13] ), .B(_AES_ENC_sa20_sub[5] ),.Z(_AES_ENC_N456 ) );
XOR2_X2 _AES_ENC_U567  ( .A(_AES_ENC_w2[12] ), .B(_AES_ENC_sa20_sub[4] ),.Z(_AES_ENC_N457 ) );
XOR2_X2 _AES_ENC_U566  ( .A(_AES_ENC_w2[11] ), .B(_AES_ENC_sa20_sub[3] ),.Z(_AES_ENC_N458 ) );
XOR2_X2 _AES_ENC_U565  ( .A(_AES_ENC_w2[10] ), .B(_AES_ENC_sa20_sub[2] ),.Z(_AES_ENC_N459 ) );
NAND2_X2 _AES_ENC_U564  ( .A1(_AES_ENC_sa23_next[0]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n367 ) );
XOR2_X2 _AES_ENC_U563  ( .A(_AES_ENC_w3[8] ), .B(_AES_ENC_text_in_r[8] ),.Z(_AES_ENC_n369 ) );
NAND2_X2 _AES_ENC_U562  ( .A1(_AES_ENC_n369 ), .A2(_AES_ENC_n1247 ), .ZN(_AES_ENC_n368 ) );
NAND2_X2 _AES_ENC_U561  ( .A1(_AES_ENC_n367 ), .A2(_AES_ENC_n368 ), .ZN(_AES_ENC_N46 ) );
XOR2_X2 _AES_ENC_U560  ( .A(_AES_ENC_w2[9] ), .B(_AES_ENC_sa20_sub[1] ), .Z(_AES_ENC_N460 ) );
XOR2_X2 _AES_ENC_U559  ( .A(_AES_ENC_w2[8] ), .B(_AES_ENC_sa20_sub[0] ), .Z(_AES_ENC_N461 ) );
XOR2_X2 _AES_ENC_U558  ( .A(_AES_ENC_w3[15] ), .B(_AES_ENC_sa21_sub[7] ),.Z(_AES_ENC_N462 ) );
XOR2_X2 _AES_ENC_U557  ( .A(_AES_ENC_w3[14] ), .B(_AES_ENC_sa21_sub[6] ),.Z(_AES_ENC_N463 ) );
XOR2_X2 _AES_ENC_U556  ( .A(_AES_ENC_w3[13] ), .B(_AES_ENC_sa21_sub[5] ),.Z(_AES_ENC_N464 ) );
XOR2_X2 _AES_ENC_U555  ( .A(_AES_ENC_w3[12] ), .B(_AES_ENC_sa21_sub[4] ),.Z(_AES_ENC_N465 ) );
XOR2_X2 _AES_ENC_U554  ( .A(_AES_ENC_w3[11] ), .B(_AES_ENC_sa21_sub[3] ),.Z(_AES_ENC_N466 ) );
XOR2_X2 _AES_ENC_U553  ( .A(_AES_ENC_w3[10] ), .B(_AES_ENC_sa21_sub[2] ),.Z(_AES_ENC_N467 ) );
XOR2_X2 _AES_ENC_U552  ( .A(_AES_ENC_w3[9] ), .B(_AES_ENC_sa21_sub[1] ), .Z(_AES_ENC_N468 ) );
XOR2_X2 _AES_ENC_U551  ( .A(_AES_ENC_w3[8] ), .B(_AES_ENC_sa21_sub[0] ), .Z(_AES_ENC_N469 ) );
NAND2_X2 _AES_ENC_U550  ( .A1(_AES_ENC_sa23_next[1]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n364 ) );
XOR2_X2 _AES_ENC_U549  ( .A(_AES_ENC_w3[9] ), .B(_AES_ENC_text_in_r[9] ),.Z(_AES_ENC_n366 ) );
NAND2_X2 _AES_ENC_U548  ( .A1(_AES_ENC_n366 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n365 ) );
NAND2_X2 _AES_ENC_U547  ( .A1(_AES_ENC_n364 ), .A2(_AES_ENC_n365 ), .ZN(_AES_ENC_N47 ) );
XOR2_X2 _AES_ENC_U546  ( .A(_AES_ENC_w0[7] ), .B(_AES_ENC_sa33_sub[7] ), .Z(_AES_ENC_N470 ) );
XOR2_X2 _AES_ENC_U545  ( .A(_AES_ENC_w0[6] ), .B(_AES_ENC_sa33_sub[6] ), .Z(_AES_ENC_N471 ) );
XOR2_X2 _AES_ENC_U544  ( .A(_AES_ENC_w0[5] ), .B(_AES_ENC_sa33_sub[5] ), .Z(_AES_ENC_N472 ) );
XOR2_X2 _AES_ENC_U543  ( .A(_AES_ENC_w0[4] ), .B(_AES_ENC_sa33_sub[4] ), .Z(_AES_ENC_N473 ) );
XOR2_X2 _AES_ENC_U542  ( .A(_AES_ENC_w0[3] ), .B(_AES_ENC_sa33_sub[3] ), .Z(_AES_ENC_N474 ) );
XOR2_X2 _AES_ENC_U541  ( .A(_AES_ENC_w0[2] ), .B(_AES_ENC_sa33_sub[2] ), .Z(_AES_ENC_N475 ) );
XOR2_X2 _AES_ENC_U540  ( .A(_AES_ENC_w0[1] ), .B(_AES_ENC_sa33_sub[1] ), .Z(_AES_ENC_N476 ) );
XOR2_X2 _AES_ENC_U539  ( .A(_AES_ENC_w0[0] ), .B(_AES_ENC_sa33_sub[0] ), .Z(_AES_ENC_N477 ) );
XOR2_X2 _AES_ENC_U538  ( .A(_AES_ENC_w1[7] ), .B(_AES_ENC_sa30_sub[7] ), .Z(_AES_ENC_N478 ) );
XOR2_X2 _AES_ENC_U537  ( .A(_AES_ENC_w1[6] ), .B(_AES_ENC_sa30_sub[6] ), .Z(_AES_ENC_N479 ) );
NAND2_X2 _AES_ENC_U536  ( .A1(_AES_ENC_sa23_next[2]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n361 ) );
XOR2_X2 _AES_ENC_U535  ( .A(_AES_ENC_w3[10] ), .B(_AES_ENC_text_in_r[10] ),.Z(_AES_ENC_n363 ) );
NAND2_X2 _AES_ENC_U534  ( .A1(_AES_ENC_n363 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n362 ) );
NAND2_X2 _AES_ENC_U533  ( .A1(_AES_ENC_n361 ), .A2(_AES_ENC_n362 ), .ZN(_AES_ENC_N48 ) );
XOR2_X2 _AES_ENC_U532  ( .A(_AES_ENC_w1[5] ), .B(_AES_ENC_sa30_sub[5] ), .Z(_AES_ENC_N480 ) );
XOR2_X2 _AES_ENC_U531  ( .A(_AES_ENC_w1[4] ), .B(_AES_ENC_sa30_sub[4] ), .Z(_AES_ENC_N481 ) );
XOR2_X2 _AES_ENC_U530  ( .A(_AES_ENC_w1[3] ), .B(_AES_ENC_sa30_sub[3] ), .Z(_AES_ENC_N482 ) );
XOR2_X2 _AES_ENC_U529  ( .A(_AES_ENC_w1[2] ), .B(_AES_ENC_sa30_sub[2] ), .Z(_AES_ENC_N483 ) );
XOR2_X2 _AES_ENC_U528  ( .A(_AES_ENC_w1[1] ), .B(_AES_ENC_sa30_sub[1] ), .Z(_AES_ENC_N484 ) );
XOR2_X2 _AES_ENC_U527  ( .A(_AES_ENC_w1[0] ), .B(_AES_ENC_sa30_sub[0] ), .Z(_AES_ENC_N485 ) );
XOR2_X2 _AES_ENC_U526  ( .A(_AES_ENC_w2[7] ), .B(_AES_ENC_sa31_sub[7] ), .Z(_AES_ENC_N486 ) );
XOR2_X2 _AES_ENC_U525  ( .A(_AES_ENC_w2[6] ), .B(_AES_ENC_sa31_sub[6] ), .Z(_AES_ENC_N487 ) );
XOR2_X2 _AES_ENC_U524  ( .A(_AES_ENC_w2[5] ), .B(_AES_ENC_sa31_sub[5] ), .Z(_AES_ENC_N488 ) );
XOR2_X2 _AES_ENC_U523  ( .A(_AES_ENC_w2[4] ), .B(_AES_ENC_sa31_sub[4] ), .Z(_AES_ENC_N489 ) );
NAND2_X2 _AES_ENC_U522  ( .A1(_AES_ENC_sa23_next[3]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n358 ) );
XOR2_X2 _AES_ENC_U521  ( .A(_AES_ENC_w3[11] ), .B(_AES_ENC_text_in_r[11] ),.Z(_AES_ENC_n3601 ) );
NAND2_X2 _AES_ENC_U520  ( .A1(_AES_ENC_n3601 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n359 ) );
NAND2_X2 _AES_ENC_U519  ( .A1(_AES_ENC_n358 ), .A2(_AES_ENC_n359 ), .ZN(_AES_ENC_N49 ) );
XOR2_X2 _AES_ENC_U518  ( .A(_AES_ENC_w2[3] ), .B(_AES_ENC_sa31_sub[3] ), .Z(_AES_ENC_N490 ) );
XOR2_X2 _AES_ENC_U517  ( .A(_AES_ENC_w2[2] ), .B(_AES_ENC_sa31_sub[2] ), .Z(_AES_ENC_N491 ) );
XOR2_X2 _AES_ENC_U516  ( .A(_AES_ENC_w2[1] ), .B(_AES_ENC_sa31_sub[1] ), .Z(_AES_ENC_N492 ) );
XOR2_X2 _AES_ENC_U515  ( .A(_AES_ENC_w2[0] ), .B(_AES_ENC_sa31_sub[0] ), .Z(_AES_ENC_N493 ) );
XOR2_X2 _AES_ENC_U514  ( .A(_AES_ENC_w3[7] ), .B(_AES_ENC_sa32_sub[7] ), .Z(_AES_ENC_N494 ) );
XOR2_X2 _AES_ENC_U513  ( .A(_AES_ENC_w3[6] ), .B(_AES_ENC_sa32_sub[6] ), .Z(_AES_ENC_N495 ) );
XOR2_X2 _AES_ENC_U512  ( .A(_AES_ENC_w3[5] ), .B(_AES_ENC_sa32_sub[5] ), .Z(_AES_ENC_N496 ) );
XOR2_X2 _AES_ENC_U511  ( .A(_AES_ENC_w3[4] ), .B(_AES_ENC_sa32_sub[4] ), .Z(_AES_ENC_N497 ) );
XOR2_X2 _AES_ENC_U510  ( .A(_AES_ENC_w3[3] ), .B(_AES_ENC_sa32_sub[3] ), .Z(_AES_ENC_N498 ) );
XOR2_X2 _AES_ENC_U509  ( .A(_AES_ENC_w3[2] ), .B(_AES_ENC_sa32_sub[2] ), .Z(_AES_ENC_N499 ) );
NAND2_X2 _AES_ENC_U508  ( .A1(_AES_ENC_sa23_next[4]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n355 ) );
XOR2_X2 _AES_ENC_U507  ( .A(_AES_ENC_w3[12] ), .B(_AES_ENC_text_in_r[12] ),.Z(_AES_ENC_n357 ) );
NAND2_X2 _AES_ENC_U506  ( .A1(_AES_ENC_n357 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n356 ) );
NAND2_X2 _AES_ENC_U505  ( .A1(_AES_ENC_n355 ), .A2(_AES_ENC_n356 ), .ZN(_AES_ENC_N50 ) );
XOR2_X2 _AES_ENC_U504  ( .A(_AES_ENC_w3[1] ), .B(_AES_ENC_sa32_sub[1] ), .Z(_AES_ENC_N500 ) );
XOR2_X2 _AES_ENC_U503  ( .A(_AES_ENC_w3[0] ), .B(_AES_ENC_sa32_sub[0] ), .Z(_AES_ENC_N501 ) );
NAND2_X2 _AES_ENC_U502  ( .A1(_AES_ENC_sa23_next[5]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n352 ) );
XOR2_X2 _AES_ENC_U501  ( .A(_AES_ENC_w3[13] ), .B(_AES_ENC_text_in_r[13] ),.Z(_AES_ENC_n354 ) );
NAND2_X2 _AES_ENC_U500  ( .A1(_AES_ENC_n354 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n353 ) );
NAND2_X2 _AES_ENC_U499  ( .A1(_AES_ENC_n352 ), .A2(_AES_ENC_n353 ), .ZN(_AES_ENC_N51 ) );
NAND2_X2 _AES_ENC_U498  ( .A1(_AES_ENC_sa23_next[6]), .A2(_AES_ENC_n1255 ),.ZN(_AES_ENC_n349 ) );
XOR2_X2 _AES_ENC_U497  ( .A(_AES_ENC_w3[14] ), .B(_AES_ENC_text_in_r[14] ),.Z(_AES_ENC_n351 ) );
NAND2_X2 _AES_ENC_U496  ( .A1(_AES_ENC_n351 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n3501 ) );
NAND2_X2 _AES_ENC_U495  ( .A1(_AES_ENC_n349 ), .A2(_AES_ENC_n3501 ), .ZN(_AES_ENC_N52 ) );
NAND2_X2 _AES_ENC_U494  ( .A1(_AES_ENC_sa23_next[7]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n346 ) );
XOR2_X2 _AES_ENC_U493  ( .A(_AES_ENC_w3[15] ), .B(_AES_ENC_text_in_r[15] ),.Z(_AES_ENC_n348 ) );
NAND2_X2 _AES_ENC_U492  ( .A1(_AES_ENC_n348 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n347 ) );
NAND2_X2 _AES_ENC_U491  ( .A1(_AES_ENC_n346 ), .A2(_AES_ENC_n347 ), .ZN(_AES_ENC_N53 ) );
NAND2_X2 _AES_ENC_U490  ( .A1(_AES_ENC_sa13_next[0]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n343 ) );
XOR2_X2 _AES_ENC_U489  ( .A(_AES_ENC_w3[16] ), .B(_AES_ENC_text_in_r[16] ),.Z(_AES_ENC_n345 ) );
NAND2_X2 _AES_ENC_U488  ( .A1(_AES_ENC_n345 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n344 ) );
NAND2_X2 _AES_ENC_U487  ( .A1(_AES_ENC_n343 ), .A2(_AES_ENC_n344 ), .ZN(_AES_ENC_N62 ) );
NAND2_X2 _AES_ENC_U486  ( .A1(_AES_ENC_sa13_next[1]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n3401 ) );
XOR2_X2 _AES_ENC_U485  ( .A(_AES_ENC_w3[17] ), .B(_AES_ENC_text_in_r[17] ),.Z(_AES_ENC_n342 ) );
NAND2_X2 _AES_ENC_U484  ( .A1(_AES_ENC_n342 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n341 ) );
NAND2_X2 _AES_ENC_U483  ( .A1(_AES_ENC_n3401 ), .A2(_AES_ENC_n341 ), .ZN(_AES_ENC_N63 ) );
NAND2_X2 _AES_ENC_U482  ( .A1(_AES_ENC_sa13_next[2]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n337 ) );
XOR2_X2 _AES_ENC_U481  ( .A(_AES_ENC_w3[18] ), .B(_AES_ENC_text_in_r[18] ),.Z(_AES_ENC_n339 ) );
NAND2_X2 _AES_ENC_U480  ( .A1(_AES_ENC_n339 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n338 ) );
NAND2_X2 _AES_ENC_U479  ( .A1(_AES_ENC_n337 ), .A2(_AES_ENC_n338 ), .ZN(_AES_ENC_N64 ) );
NAND2_X2 _AES_ENC_U478  ( .A1(_AES_ENC_sa13_next[3]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n334 ) );
XOR2_X2 _AES_ENC_U477  ( .A(_AES_ENC_w3[19] ), .B(_AES_ENC_text_in_r[19] ),.Z(_AES_ENC_n336 ) );
NAND2_X2 _AES_ENC_U476  ( .A1(_AES_ENC_n336 ), .A2(_AES_ENC_n1248 ), .ZN(_AES_ENC_n335 ) );
NAND2_X2 _AES_ENC_U475  ( .A1(_AES_ENC_n334 ), .A2(_AES_ENC_n335 ), .ZN(_AES_ENC_N65 ) );
NAND2_X2 _AES_ENC_U474  ( .A1(_AES_ENC_sa13_next[4]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n331 ) );
XOR2_X2 _AES_ENC_U473  ( .A(_AES_ENC_w3[20] ), .B(_AES_ENC_text_in_r[20] ),.Z(_AES_ENC_n333 ) );
NAND2_X2 _AES_ENC_U472  ( .A1(_AES_ENC_n333 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n332 ) );
NAND2_X2 _AES_ENC_U471  ( .A1(_AES_ENC_n331 ), .A2(_AES_ENC_n332 ), .ZN(_AES_ENC_N66 ) );
NAND2_X2 _AES_ENC_U470  ( .A1(_AES_ENC_sa13_next[5]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n328 ) );
XOR2_X2 _AES_ENC_U469  ( .A(_AES_ENC_w3[21] ), .B(_AES_ENC_text_in_r[21] ),.Z(_AES_ENC_n3301 ) );
NAND2_X2 _AES_ENC_U468  ( .A1(_AES_ENC_n3301 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n329 ) );
NAND2_X2 _AES_ENC_U467  ( .A1(_AES_ENC_n328 ), .A2(_AES_ENC_n329 ), .ZN(_AES_ENC_N67 ) );
NAND2_X2 _AES_ENC_U466  ( .A1(_AES_ENC_sa13_next[6]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n325 ) );
XOR2_X2 _AES_ENC_U465  ( .A(_AES_ENC_w3[22] ), .B(_AES_ENC_text_in_r[22] ),.Z(_AES_ENC_n327 ) );
NAND2_X2 _AES_ENC_U464  ( .A1(_AES_ENC_n327 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n326 ) );
NAND2_X2 _AES_ENC_U463  ( .A1(_AES_ENC_n325 ), .A2(_AES_ENC_n326 ), .ZN(_AES_ENC_N68 ) );
NAND2_X2 _AES_ENC_U462  ( .A1(_AES_ENC_sa13_next[7]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n322 ) );
XOR2_X2 _AES_ENC_U461  ( .A(_AES_ENC_w3[23] ), .B(_AES_ENC_text_in_r[23] ),.Z(_AES_ENC_n324 ) );
NAND2_X2 _AES_ENC_U460  ( .A1(_AES_ENC_n324 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n323 ) );
NAND2_X2 _AES_ENC_U459  ( .A1(_AES_ENC_n322 ), .A2(_AES_ENC_n323 ), .ZN(_AES_ENC_N69 ) );
NAND2_X2 _AES_ENC_U458  ( .A1(_AES_ENC_sa03_next[0]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n319 ) );
XOR2_X2 _AES_ENC_U457  ( .A(_AES_ENC_w3[24] ), .B(_AES_ENC_text_in_r[24] ),.Z(_AES_ENC_n321 ) );
NAND2_X2 _AES_ENC_U456  ( .A1(_AES_ENC_n321 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n3201 ) );
NAND2_X2 _AES_ENC_U455  ( .A1(_AES_ENC_n319 ), .A2(_AES_ENC_n3201 ), .ZN(_AES_ENC_N78 ) );
NAND2_X2 _AES_ENC_U454  ( .A1(_AES_ENC_sa03_next[1]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n316 ) );
XOR2_X2 _AES_ENC_U453  ( .A(_AES_ENC_w3[25] ), .B(_AES_ENC_text_in_r[25] ),.Z(_AES_ENC_n318 ) );
NAND2_X2 _AES_ENC_U452  ( .A1(_AES_ENC_n318 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n317 ) );
NAND2_X2 _AES_ENC_U451  ( .A1(_AES_ENC_n316 ), .A2(_AES_ENC_n317 ), .ZN(_AES_ENC_N79 ) );
NAND2_X2 _AES_ENC_U450  ( .A1(_AES_ENC_sa03_next[2]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n313 ) );
XOR2_X2 _AES_ENC_U449  ( .A(_AES_ENC_w3[26] ), .B(_AES_ENC_text_in_r[26] ),.Z(_AES_ENC_n315 ) );
NAND2_X2 _AES_ENC_U448  ( .A1(_AES_ENC_n315 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n314 ) );
NAND2_X2 _AES_ENC_U447  ( .A1(_AES_ENC_n313 ), .A2(_AES_ENC_n314 ), .ZN(_AES_ENC_N80 ) );
NAND2_X2 _AES_ENC_U446  ( .A1(_AES_ENC_sa03_next[3]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n3101 ) );
XOR2_X2 _AES_ENC_U445  ( .A(_AES_ENC_w3[27] ), .B(_AES_ENC_text_in_r[27] ),.Z(_AES_ENC_n312 ) );
NAND2_X2 _AES_ENC_U444  ( .A1(_AES_ENC_n312 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n311 ) );
NAND2_X2 _AES_ENC_U443  ( .A1(_AES_ENC_n3101 ), .A2(_AES_ENC_n311 ), .ZN(_AES_ENC_N81 ) );
NAND2_X2 _AES_ENC_U442  ( .A1(_AES_ENC_sa03_next[4]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n307 ) );
XOR2_X2 _AES_ENC_U441  ( .A(_AES_ENC_w3[28] ), .B(_AES_ENC_text_in_r[28] ),.Z(_AES_ENC_n309 ) );
NAND2_X2 _AES_ENC_U440  ( .A1(_AES_ENC_n309 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n308 ) );
NAND2_X2 _AES_ENC_U439  ( .A1(_AES_ENC_n307 ), .A2(_AES_ENC_n308 ), .ZN(_AES_ENC_N82 ) );
NAND2_X2 _AES_ENC_U438  ( .A1(_AES_ENC_sa03_next[5]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n304 ) );
XOR2_X2 _AES_ENC_U437  ( .A(_AES_ENC_w3[29] ), .B(_AES_ENC_text_in_r[29] ),.Z(_AES_ENC_n306 ) );
NAND2_X2 _AES_ENC_U436  ( .A1(_AES_ENC_n306 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n305 ) );
NAND2_X2 _AES_ENC_U435  ( .A1(_AES_ENC_n304 ), .A2(_AES_ENC_n305 ), .ZN(_AES_ENC_N83 ) );
NAND2_X2 _AES_ENC_U434  ( .A1(_AES_ENC_sa03_next[6]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n301 ) );
XOR2_X2 _AES_ENC_U433  ( .A(_AES_ENC_w3[30] ), .B(_AES_ENC_text_in_r[30] ),.Z(_AES_ENC_n303 ) );
NAND2_X2 _AES_ENC_U432  ( .A1(_AES_ENC_n303 ), .A2(_AES_ENC_n1249 ), .ZN(_AES_ENC_n302 ) );
NAND2_X2 _AES_ENC_U431  ( .A1(_AES_ENC_n301 ), .A2(_AES_ENC_n302 ), .ZN(_AES_ENC_N84 ) );
NAND2_X2 _AES_ENC_U430  ( .A1(_AES_ENC_sa03_next[7]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n298 ) );
XOR2_X2 _AES_ENC_U429  ( .A(_AES_ENC_w3[31] ), .B(_AES_ENC_text_in_r[31] ),.Z(_AES_ENC_n3001 ) );
NAND2_X2 _AES_ENC_U428  ( .A1(_AES_ENC_n3001 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n299 ) );
NAND2_X2 _AES_ENC_U427  ( .A1(_AES_ENC_n298 ), .A2(_AES_ENC_n299 ), .ZN(_AES_ENC_N85 ) );
NAND2_X2 _AES_ENC_U426  ( .A1(_AES_ENC_sa32_next[0]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n295 ) );
XOR2_X2 _AES_ENC_U425  ( .A(_AES_ENC_w2[0] ), .B(_AES_ENC_text_in_r[32] ),.Z(_AES_ENC_n297 ) );
NAND2_X2 _AES_ENC_U424  ( .A1(_AES_ENC_n297 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n296 ) );
NAND2_X2 _AES_ENC_U423  ( .A1(_AES_ENC_n295 ), .A2(_AES_ENC_n296 ), .ZN(_AES_ENC_N94 ) );
NAND2_X2 _AES_ENC_U422  ( .A1(_AES_ENC_sa32_next[1]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n292 ) );
XOR2_X2 _AES_ENC_U421  ( .A(_AES_ENC_w2[1] ), .B(_AES_ENC_text_in_r[33] ),.Z(_AES_ENC_n294 ) );
NAND2_X2 _AES_ENC_U420  ( .A1(_AES_ENC_n294 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n293 ) );
NAND2_X2 _AES_ENC_U419  ( .A1(_AES_ENC_n292 ), .A2(_AES_ENC_n293 ), .ZN(_AES_ENC_N95 ) );
NAND2_X2 _AES_ENC_U418  ( .A1(_AES_ENC_sa32_next[2]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n289 ) );
XOR2_X2 _AES_ENC_U417  ( .A(_AES_ENC_w2[2] ), .B(_AES_ENC_text_in_r[34] ),.Z(_AES_ENC_n291 ) );
NAND2_X2 _AES_ENC_U416  ( .A1(_AES_ENC_n291 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n290 ) );
NAND2_X2 _AES_ENC_U415  ( .A1(_AES_ENC_n289 ), .A2(_AES_ENC_n290 ), .ZN(_AES_ENC_N96 ) );
NAND2_X2 _AES_ENC_U414  ( .A1(_AES_ENC_sa32_next[3]), .A2(_AES_ENC_n1256 ),.ZN(_AES_ENC_n286 ) );
XOR2_X2 _AES_ENC_U413  ( .A(_AES_ENC_w2[3] ), .B(_AES_ENC_text_in_r[35] ),.Z(_AES_ENC_n288 ) );
NAND2_X2 _AES_ENC_U412  ( .A1(_AES_ENC_n288 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n287 ) );
NAND2_X2 _AES_ENC_U411  ( .A1(_AES_ENC_n286 ), .A2(_AES_ENC_n287 ), .ZN(_AES_ENC_N97 ) );
NAND2_X2 _AES_ENC_U410  ( .A1(_AES_ENC_sa32_next[4]), .A2(_AES_ENC_n1252 ),.ZN(_AES_ENC_n283 ) );
XOR2_X2 _AES_ENC_U409  ( .A(_AES_ENC_w2[4] ), .B(_AES_ENC_text_in_r[36] ),.Z(_AES_ENC_n285 ) );
NAND2_X2 _AES_ENC_U408  ( .A1(_AES_ENC_n285 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n284 ) );
NAND2_X2 _AES_ENC_U407  ( .A1(_AES_ENC_n283 ), .A2(_AES_ENC_n284 ), .ZN(_AES_ENC_N98 ) );
NAND2_X2 _AES_ENC_U406  ( .A1(_AES_ENC_sa32_next[5]), .A2(_AES_ENC_n1251 ),.ZN(_AES_ENC_n280 ) );
XOR2_X2 _AES_ENC_U405  ( .A(_AES_ENC_w2[5] ), .B(_AES_ENC_text_in_r[37] ),.Z(_AES_ENC_n282 ) );
NAND2_X2 _AES_ENC_U404  ( .A1(_AES_ENC_n282 ), .A2(_AES_ENC_n1250 ), .ZN(_AES_ENC_n281 ) );
NAND2_X2 _AES_ENC_U403  ( .A1(_AES_ENC_n280 ), .A2(_AES_ENC_n281 ), .ZN(_AES_ENC_N99 ) );
NAND2_X2 _AES_ENC_U402  ( .A1(aes_text_in[0]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n278 ) );
NAND2_X2 _AES_ENC_U401  ( .A1(_AES_ENC_text_in_r[0] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n279 ) );
NAND2_X2 _AES_ENC_U400  ( .A1(_AES_ENC_n278 ), .A2(_AES_ENC_n279 ), .ZN(_AES_ENC_n661 ) );
NAND2_X2 _AES_ENC_U399  ( .A1(aes_text_in[1]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2760 ) );
NAND2_X2 _AES_ENC_U398  ( .A1(_AES_ENC_text_in_r[1] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2770 ) );
NAND2_X2 _AES_ENC_U397  ( .A1(_AES_ENC_n2760 ), .A2(_AES_ENC_n2770 ), .ZN(_AES_ENC_n662 ) );
NAND2_X2 _AES_ENC_U396  ( .A1(aes_text_in[2]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2740 ) );
NAND2_X2 _AES_ENC_U395  ( .A1(_AES_ENC_text_in_r[2] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2750 ) );
NAND2_X2 _AES_ENC_U394  ( .A1(_AES_ENC_n2740 ), .A2(_AES_ENC_n2750 ), .ZN(_AES_ENC_n663 ) );
NAND2_X2 _AES_ENC_U393  ( .A1(aes_text_in[3]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2720 ) );
NAND2_X2 _AES_ENC_U392  ( .A1(_AES_ENC_text_in_r[3] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2730 ) );
NAND2_X2 _AES_ENC_U391  ( .A1(_AES_ENC_n2720 ), .A2(_AES_ENC_n2730 ), .ZN(_AES_ENC_n664 ) );
NAND2_X2 _AES_ENC_U390  ( .A1(aes_text_in[4]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2700 ) );
NAND2_X2 _AES_ENC_U389  ( .A1(_AES_ENC_text_in_r[4] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2710 ) );
NAND2_X2 _AES_ENC_U388  ( .A1(_AES_ENC_n2700 ), .A2(_AES_ENC_n2710 ), .ZN(_AES_ENC_n665 ) );
NAND2_X2 _AES_ENC_U387  ( .A1(aes_text_in[5]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n268 ) );
NAND2_X2 _AES_ENC_U386  ( .A1(_AES_ENC_text_in_r[5] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n269 ) );
NAND2_X2 _AES_ENC_U385  ( .A1(_AES_ENC_n268 ), .A2(_AES_ENC_n269 ), .ZN(_AES_ENC_n666 ) );
NAND2_X2 _AES_ENC_U384  ( .A1(aes_text_in[6]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n266 ) );
NAND2_X2 _AES_ENC_U383  ( .A1(_AES_ENC_text_in_r[6] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n267 ) );
NAND2_X2 _AES_ENC_U382  ( .A1(_AES_ENC_n266 ), .A2(_AES_ENC_n267 ), .ZN(_AES_ENC_n667 ) );
NAND2_X2 _AES_ENC_U381  ( .A1(aes_text_in[7]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n264 ) );
NAND2_X2 _AES_ENC_U380  ( .A1(_AES_ENC_text_in_r[7] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n265 ) );
NAND2_X2 _AES_ENC_U379  ( .A1(_AES_ENC_n264 ), .A2(_AES_ENC_n265 ), .ZN(_AES_ENC_n668 ) );
NAND2_X2 _AES_ENC_U378  ( .A1(aes_text_in[8]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n262 ) );
NAND2_X2 _AES_ENC_U377  ( .A1(_AES_ENC_text_in_r[8] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n263 ) );
NAND2_X2 _AES_ENC_U376  ( .A1(_AES_ENC_n262 ), .A2(_AES_ENC_n263 ), .ZN(_AES_ENC_n669 ) );
NAND2_X2 _AES_ENC_U375  ( .A1(aes_text_in[9]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2600 ) );
NAND2_X2 _AES_ENC_U374  ( .A1(_AES_ENC_text_in_r[9] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2610 ) );
NAND2_X2 _AES_ENC_U373  ( .A1(_AES_ENC_n2600 ), .A2(_AES_ENC_n2610 ), .ZN(_AES_ENC_n670 ) );
NAND2_X2 _AES_ENC_U372  ( .A1(aes_text_in[10]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2580 ) );
NAND2_X2 _AES_ENC_U371  ( .A1(_AES_ENC_text_in_r[10] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2590 ) );
NAND2_X2 _AES_ENC_U370  ( .A1(_AES_ENC_n2580 ), .A2(_AES_ENC_n2590 ), .ZN(_AES_ENC_n671 ) );
NAND2_X2 _AES_ENC_U369  ( .A1(aes_text_in[11]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2560 ) );
NAND2_X2 _AES_ENC_U368  ( .A1(_AES_ENC_text_in_r[11] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2570 ) );
NAND2_X2 _AES_ENC_U367  ( .A1(_AES_ENC_n2560 ), .A2(_AES_ENC_n2570 ), .ZN(_AES_ENC_n672 ) );
NAND2_X2 _AES_ENC_U366  ( .A1(aes_text_in[12]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2540 ) );
NAND2_X2 _AES_ENC_U365  ( .A1(_AES_ENC_text_in_r[12] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2550 ) );
NAND2_X2 _AES_ENC_U364  ( .A1(_AES_ENC_n2540 ), .A2(_AES_ENC_n2550 ), .ZN(_AES_ENC_n673 ) );
NAND2_X2 _AES_ENC_U363  ( .A1(aes_text_in[13]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n252 ) );
NAND2_X2 _AES_ENC_U362  ( .A1(_AES_ENC_text_in_r[13] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n253 ) );
NAND2_X2 _AES_ENC_U361  ( .A1(_AES_ENC_n252 ), .A2(_AES_ENC_n253 ), .ZN(_AES_ENC_n674 ) );
NAND2_X2 _AES_ENC_U360  ( .A1(aes_text_in[14]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n250 ) );
NAND2_X2 _AES_ENC_U359  ( .A1(_AES_ENC_text_in_r[14] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n251 ) );
NAND2_X2 _AES_ENC_U358  ( .A1(_AES_ENC_n250 ), .A2(_AES_ENC_n251 ), .ZN(_AES_ENC_n675 ) );
NAND2_X2 _AES_ENC_U357  ( .A1(aes_text_in[15]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n248 ) );
NAND2_X2 _AES_ENC_U356  ( .A1(_AES_ENC_text_in_r[15] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n249 ) );
NAND2_X2 _AES_ENC_U355  ( .A1(_AES_ENC_n248 ), .A2(_AES_ENC_n249 ), .ZN(_AES_ENC_n676 ) );
NAND2_X2 _AES_ENC_U354  ( .A1(aes_text_in[16]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n246 ) );
NAND2_X2 _AES_ENC_U353  ( .A1(_AES_ENC_text_in_r[16] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n247 ) );
NAND2_X2 _AES_ENC_U352  ( .A1(_AES_ENC_n246 ), .A2(_AES_ENC_n247 ), .ZN(_AES_ENC_n677 ) );
NAND2_X2 _AES_ENC_U351  ( .A1(aes_text_in[17]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2440 ) );
NAND2_X2 _AES_ENC_U350  ( .A1(_AES_ENC_text_in_r[17] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2450 ) );
NAND2_X2 _AES_ENC_U349  ( .A1(_AES_ENC_n2440 ), .A2(_AES_ENC_n2450 ), .ZN(_AES_ENC_n678 ) );
NAND2_X2 _AES_ENC_U348  ( .A1(aes_text_in[18]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2420 ) );
NAND2_X2 _AES_ENC_U347  ( .A1(_AES_ENC_text_in_r[18] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2430 ) );
NAND2_X2 _AES_ENC_U346  ( .A1(_AES_ENC_n2420 ), .A2(_AES_ENC_n2430 ), .ZN(_AES_ENC_n679 ) );
NAND2_X2 _AES_ENC_U345  ( .A1(aes_text_in[19]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2400 ) );
NAND2_X2 _AES_ENC_U344  ( .A1(_AES_ENC_text_in_r[19] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2410 ) );
NAND2_X2 _AES_ENC_U343  ( .A1(_AES_ENC_n2400 ), .A2(_AES_ENC_n2410 ), .ZN(_AES_ENC_n680 ) );
NAND2_X2 _AES_ENC_U342  ( .A1(aes_text_in[20]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2380 ) );
NAND2_X2 _AES_ENC_U341  ( .A1(_AES_ENC_text_in_r[20] ), .A2(_AES_ENC_n1264 ),.ZN(_AES_ENC_n2390 ) );
NAND2_X2 _AES_ENC_U340  ( .A1(_AES_ENC_n2380 ), .A2(_AES_ENC_n2390 ), .ZN(_AES_ENC_n681 ) );
NAND2_X2 _AES_ENC_U339  ( .A1(aes_text_in[21]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n236 ) );
NAND2_X2 _AES_ENC_U338  ( .A1(_AES_ENC_text_in_r[21] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n237 ) );
NAND2_X2 _AES_ENC_U337  ( .A1(_AES_ENC_n236 ), .A2(_AES_ENC_n237 ), .ZN(_AES_ENC_n682 ) );
NAND2_X2 _AES_ENC_U336  ( .A1(aes_text_in[22]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n234 ) );
NAND2_X2 _AES_ENC_U335  ( .A1(_AES_ENC_text_in_r[22] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n235 ) );
NAND2_X2 _AES_ENC_U334  ( .A1(_AES_ENC_n234 ), .A2(_AES_ENC_n235 ), .ZN(_AES_ENC_n683 ) );
NAND2_X2 _AES_ENC_U333  ( .A1(aes_text_in[23]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n232 ) );
NAND2_X2 _AES_ENC_U332  ( .A1(_AES_ENC_text_in_r[23] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n233 ) );
NAND2_X2 _AES_ENC_U331  ( .A1(_AES_ENC_n232 ), .A2(_AES_ENC_n233 ), .ZN(_AES_ENC_n684 ) );
NAND2_X2 _AES_ENC_U330  ( .A1(aes_text_in[24]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n230 ) );
NAND2_X2 _AES_ENC_U329  ( .A1(_AES_ENC_text_in_r[24] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n231 ) );
NAND2_X2 _AES_ENC_U328  ( .A1(_AES_ENC_n230 ), .A2(_AES_ENC_n231 ), .ZN(_AES_ENC_n685 ) );
NAND2_X2 _AES_ENC_U327  ( .A1(aes_text_in[25]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2280 ) );
NAND2_X2 _AES_ENC_U326  ( .A1(_AES_ENC_text_in_r[25] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2290 ) );
NAND2_X2 _AES_ENC_U325  ( .A1(_AES_ENC_n2280 ), .A2(_AES_ENC_n2290 ), .ZN(_AES_ENC_n686 ) );
NAND2_X2 _AES_ENC_U324  ( .A1(aes_text_in[26]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2260 ) );
NAND2_X2 _AES_ENC_U323  ( .A1(_AES_ENC_text_in_r[26] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2270 ) );
NAND2_X2 _AES_ENC_U322  ( .A1(_AES_ENC_n2260 ), .A2(_AES_ENC_n2270 ), .ZN(_AES_ENC_n687 ) );
NAND2_X2 _AES_ENC_U321  ( .A1(aes_text_in[27]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2240 ) );
NAND2_X2 _AES_ENC_U320  ( .A1(_AES_ENC_text_in_r[27] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2250 ) );
NAND2_X2 _AES_ENC_U319  ( .A1(_AES_ENC_n2240 ), .A2(_AES_ENC_n2250 ), .ZN(_AES_ENC_n688 ) );
NAND2_X2 _AES_ENC_U318  ( .A1(aes_text_in[28]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2220 ) );
NAND2_X2 _AES_ENC_U317  ( .A1(_AES_ENC_text_in_r[28] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2230 ) );
NAND2_X2 _AES_ENC_U316  ( .A1(_AES_ENC_n2220 ), .A2(_AES_ENC_n2230 ), .ZN(_AES_ENC_n689 ) );
NAND2_X2 _AES_ENC_U315  ( .A1(aes_text_in[29]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n220 ) );
NAND2_X2 _AES_ENC_U314  ( .A1(_AES_ENC_text_in_r[29] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n221 ) );
NAND2_X2 _AES_ENC_U313  ( .A1(_AES_ENC_n220 ), .A2(_AES_ENC_n221 ), .ZN(_AES_ENC_n690 ) );
NAND2_X2 _AES_ENC_U312  ( .A1(aes_text_in[30]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n218 ) );
NAND2_X2 _AES_ENC_U311  ( .A1(_AES_ENC_text_in_r[30] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n219 ) );
NAND2_X2 _AES_ENC_U310  ( .A1(_AES_ENC_n218 ), .A2(_AES_ENC_n219 ), .ZN(_AES_ENC_n691 ) );
NAND2_X2 _AES_ENC_U309  ( .A1(aes_text_in[31]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n216 ) );
NAND2_X2 _AES_ENC_U308  ( .A1(_AES_ENC_text_in_r[31] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n217 ) );
NAND2_X2 _AES_ENC_U307  ( .A1(_AES_ENC_n216 ), .A2(_AES_ENC_n217 ), .ZN(_AES_ENC_n692 ) );
NAND2_X2 _AES_ENC_U306  ( .A1(aes_text_in[32]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n214 ) );
NAND2_X2 _AES_ENC_U305  ( .A1(_AES_ENC_text_in_r[32] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n215 ) );
NAND2_X2 _AES_ENC_U304  ( .A1(_AES_ENC_n214 ), .A2(_AES_ENC_n215 ), .ZN(_AES_ENC_n693 ) );
NAND2_X2 _AES_ENC_U303  ( .A1(aes_text_in[33]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2120 ) );
NAND2_X2 _AES_ENC_U302  ( .A1(_AES_ENC_text_in_r[33] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2130 ) );
NAND2_X2 _AES_ENC_U301  ( .A1(_AES_ENC_n2120 ), .A2(_AES_ENC_n2130 ), .ZN(_AES_ENC_n694 ) );
NAND2_X2 _AES_ENC_U300  ( .A1(aes_text_in[34]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2100 ) );
NAND2_X2 _AES_ENC_U299  ( .A1(_AES_ENC_text_in_r[34] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2110 ) );
NAND2_X2 _AES_ENC_U298  ( .A1(_AES_ENC_n2100 ), .A2(_AES_ENC_n2110 ), .ZN(_AES_ENC_n695 ) );
NAND2_X2 _AES_ENC_U297  ( .A1(aes_text_in[35]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2080 ) );
NAND2_X2 _AES_ENC_U296  ( .A1(_AES_ENC_text_in_r[35] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2090 ) );
NAND2_X2 _AES_ENC_U295  ( .A1(_AES_ENC_n2080 ), .A2(_AES_ENC_n2090 ), .ZN(_AES_ENC_n696 ) );
NAND2_X2 _AES_ENC_U294  ( .A1(aes_text_in[36]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n2060 ) );
NAND2_X2 _AES_ENC_U293  ( .A1(_AES_ENC_text_in_r[36] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n2070 ) );
NAND2_X2 _AES_ENC_U292  ( .A1(_AES_ENC_n2060 ), .A2(_AES_ENC_n2070 ), .ZN(_AES_ENC_n697 ) );
NAND2_X2 _AES_ENC_U291  ( .A1(aes_text_in[37]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n204 ) );
NAND2_X2 _AES_ENC_U290  ( .A1(_AES_ENC_text_in_r[37] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n205 ) );
NAND2_X2 _AES_ENC_U289  ( .A1(_AES_ENC_n204 ), .A2(_AES_ENC_n205 ), .ZN(_AES_ENC_n698 ) );
NAND2_X2 _AES_ENC_U288  ( .A1(aes_text_in[38]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n202 ) );
NAND2_X2 _AES_ENC_U287  ( .A1(_AES_ENC_text_in_r[38] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n203 ) );
NAND2_X2 _AES_ENC_U286  ( .A1(_AES_ENC_n202 ), .A2(_AES_ENC_n203 ), .ZN(_AES_ENC_n699 ) );
NAND2_X2 _AES_ENC_U285  ( .A1(aes_text_in[39]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n200 ) );
NAND2_X2 _AES_ENC_U284  ( .A1(_AES_ENC_text_in_r[39] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n201 ) );
NAND2_X2 _AES_ENC_U283  ( .A1(_AES_ENC_n200 ), .A2(_AES_ENC_n201 ), .ZN(_AES_ENC_n700 ) );
NAND2_X2 _AES_ENC_U282  ( .A1(aes_text_in[40]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1981 ) );
NAND2_X2 _AES_ENC_U281  ( .A1(_AES_ENC_text_in_r[40] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n199 ) );
NAND2_X2 _AES_ENC_U280  ( .A1(_AES_ENC_n1981 ), .A2(_AES_ENC_n199 ), .ZN(_AES_ENC_n701 ) );
NAND2_X2 _AES_ENC_U279  ( .A1(aes_text_in[41]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1960 ) );
NAND2_X2 _AES_ENC_U278  ( .A1(_AES_ENC_text_in_r[41] ), .A2(_AES_ENC_n1263 ),.ZN(_AES_ENC_n1970 ) );
NAND2_X2 _AES_ENC_U277  ( .A1(_AES_ENC_n1960 ), .A2(_AES_ENC_n1970 ), .ZN(_AES_ENC_n702 ) );
NAND2_X2 _AES_ENC_U276  ( .A1(aes_text_in[42]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1940 ) );
NAND2_X2 _AES_ENC_U275  ( .A1(_AES_ENC_text_in_r[42] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1950 ) );
NAND2_X2 _AES_ENC_U274  ( .A1(_AES_ENC_n1940 ), .A2(_AES_ENC_n1950 ), .ZN(_AES_ENC_n703 ) );
NAND2_X2 _AES_ENC_U273  ( .A1(aes_text_in[43]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1920 ) );
NAND2_X2 _AES_ENC_U272  ( .A1(_AES_ENC_text_in_r[43] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1930 ) );
NAND2_X2 _AES_ENC_U271  ( .A1(_AES_ENC_n1920 ), .A2(_AES_ENC_n1930 ), .ZN(_AES_ENC_n704 ) );
NAND2_X2 _AES_ENC_U270  ( .A1(aes_text_in[44]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1900 ) );
NAND2_X2 _AES_ENC_U269  ( .A1(_AES_ENC_text_in_r[44] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1910 ) );
NAND2_X2 _AES_ENC_U268  ( .A1(_AES_ENC_n1900 ), .A2(_AES_ENC_n1910 ), .ZN(_AES_ENC_n705 ) );
NAND2_X2 _AES_ENC_U267  ( .A1(aes_text_in[45]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n188 ) );
NAND2_X2 _AES_ENC_U266  ( .A1(_AES_ENC_text_in_r[45] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n189 ) );
NAND2_X2 _AES_ENC_U265  ( .A1(_AES_ENC_n188 ), .A2(_AES_ENC_n189 ), .ZN(_AES_ENC_n706 ) );
NAND2_X2 _AES_ENC_U264  ( .A1(aes_text_in[46]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n186 ) );
NAND2_X2 _AES_ENC_U263  ( .A1(_AES_ENC_text_in_r[46] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n187 ) );
NAND2_X2 _AES_ENC_U262  ( .A1(_AES_ENC_n186 ), .A2(_AES_ENC_n187 ), .ZN(_AES_ENC_n707 ) );
NAND2_X2 _AES_ENC_U261  ( .A1(aes_text_in[47]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n184 ) );
NAND2_X2 _AES_ENC_U260  ( .A1(_AES_ENC_text_in_r[47] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n185 ) );
NAND2_X2 _AES_ENC_U259  ( .A1(_AES_ENC_n184 ), .A2(_AES_ENC_n185 ), .ZN(_AES_ENC_n708 ) );
NAND2_X2 _AES_ENC_U258  ( .A1(aes_text_in[48]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n182 ) );
NAND2_X2 _AES_ENC_U257  ( .A1(_AES_ENC_text_in_r[48] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n183 ) );
NAND2_X2 _AES_ENC_U256  ( .A1(_AES_ENC_n182 ), .A2(_AES_ENC_n183 ), .ZN(_AES_ENC_n709 ) );
NAND2_X2 _AES_ENC_U255  ( .A1(aes_text_in[49]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1800 ) );
NAND2_X2 _AES_ENC_U254  ( .A1(_AES_ENC_text_in_r[49] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1810 ) );
NAND2_X2 _AES_ENC_U253  ( .A1(_AES_ENC_n1800 ), .A2(_AES_ENC_n1810 ), .ZN(_AES_ENC_n710 ) );
NAND2_X2 _AES_ENC_U252  ( .A1(aes_text_in[50]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1780 ) );
NAND2_X2 _AES_ENC_U251  ( .A1(_AES_ENC_text_in_r[50] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1790 ) );
NAND2_X2 _AES_ENC_U250  ( .A1(_AES_ENC_n1780 ), .A2(_AES_ENC_n1790 ), .ZN(_AES_ENC_n711 ) );
NAND2_X2 _AES_ENC_U249  ( .A1(aes_text_in[51]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1760 ) );
NAND2_X2 _AES_ENC_U248  ( .A1(_AES_ENC_text_in_r[51] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1770 ) );
NAND2_X2 _AES_ENC_U247  ( .A1(_AES_ENC_n1760 ), .A2(_AES_ENC_n1770 ), .ZN(_AES_ENC_n712 ) );
NAND2_X2 _AES_ENC_U246  ( .A1(aes_text_in[52]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n1740 ) );
NAND2_X2 _AES_ENC_U245  ( .A1(_AES_ENC_text_in_r[52] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1750 ) );
NAND2_X2 _AES_ENC_U244  ( .A1(_AES_ENC_n1740 ), .A2(_AES_ENC_n1750 ), .ZN(_AES_ENC_n713 ) );
NAND2_X2 _AES_ENC_U243  ( .A1(aes_text_in[53]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n172 ) );
NAND2_X2 _AES_ENC_U242  ( .A1(_AES_ENC_text_in_r[53] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n173 ) );
NAND2_X2 _AES_ENC_U241  ( .A1(_AES_ENC_n172 ), .A2(_AES_ENC_n173 ), .ZN(_AES_ENC_n714 ) );
NAND2_X2 _AES_ENC_U240  ( .A1(aes_text_in[54]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n170 ) );
NAND2_X2 _AES_ENC_U239  ( .A1(_AES_ENC_text_in_r[54] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n171 ) );
NAND2_X2 _AES_ENC_U238  ( .A1(_AES_ENC_n170 ), .A2(_AES_ENC_n171 ), .ZN(_AES_ENC_n715 ) );
NAND2_X2 _AES_ENC_U237  ( .A1(aes_text_in[55]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n168 ) );
NAND2_X2 _AES_ENC_U236  ( .A1(_AES_ENC_text_in_r[55] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n169 ) );
NAND2_X2 _AES_ENC_U235  ( .A1(_AES_ENC_n168 ), .A2(_AES_ENC_n169 ), .ZN(_AES_ENC_n716 ) );
NAND2_X2 _AES_ENC_U234  ( .A1(aes_text_in[56]), .A2(_AES_ENC_n1257 ), .ZN(_AES_ENC_n166 ) );
NAND2_X2 _AES_ENC_U233  ( .A1(_AES_ENC_text_in_r[56] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n167 ) );
NAND2_X2 _AES_ENC_U232  ( .A1(_AES_ENC_n166 ), .A2(_AES_ENC_n167 ), .ZN(_AES_ENC_n717 ) );
NAND2_X2 _AES_ENC_U231  ( .A1(aes_text_in[57]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n1640 ) );
NAND2_X2 _AES_ENC_U230  ( .A1(_AES_ENC_text_in_r[57] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1650 ) );
NAND2_X2 _AES_ENC_U229  ( .A1(_AES_ENC_n1640 ), .A2(_AES_ENC_n1650 ), .ZN(_AES_ENC_n718 ) );
NAND2_X2 _AES_ENC_U228  ( .A1(aes_text_in[58]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n1620 ) );
NAND2_X2 _AES_ENC_U227  ( .A1(_AES_ENC_text_in_r[58] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1630 ) );
NAND2_X2 _AES_ENC_U226  ( .A1(_AES_ENC_n1620 ), .A2(_AES_ENC_n1630 ), .ZN(_AES_ENC_n719 ) );
NAND2_X2 _AES_ENC_U225  ( .A1(aes_text_in[59]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n1600 ) );
NAND2_X2 _AES_ENC_U224  ( .A1(_AES_ENC_text_in_r[59] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1610 ) );
NAND2_X2 _AES_ENC_U223  ( .A1(_AES_ENC_n1600 ), .A2(_AES_ENC_n1610 ), .ZN(_AES_ENC_n720 ) );
NAND2_X2 _AES_ENC_U222  ( .A1(aes_text_in[60]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n1580 ) );
NAND2_X2 _AES_ENC_U221  ( .A1(_AES_ENC_text_in_r[60] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n1590 ) );
NAND2_X2 _AES_ENC_U220  ( .A1(_AES_ENC_n1580 ), .A2(_AES_ENC_n1590 ), .ZN(_AES_ENC_n721 ) );
NAND2_X2 _AES_ENC_U219  ( .A1(aes_text_in[61]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n156 ) );
NAND2_X2 _AES_ENC_U218  ( .A1(_AES_ENC_text_in_r[61] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n157 ) );
NAND2_X2 _AES_ENC_U217  ( .A1(_AES_ENC_n156 ), .A2(_AES_ENC_n157 ), .ZN(_AES_ENC_n722 ) );
NAND2_X2 _AES_ENC_U216  ( .A1(aes_text_in[62]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n154 ) );
NAND2_X2 _AES_ENC_U215  ( .A1(_AES_ENC_text_in_r[62] ), .A2(_AES_ENC_n1262 ),.ZN(_AES_ENC_n155 ) );
NAND2_X2 _AES_ENC_U214  ( .A1(_AES_ENC_n154 ), .A2(_AES_ENC_n155 ), .ZN(_AES_ENC_n723 ) );
NAND2_X2 _AES_ENC_U213  ( .A1(aes_text_in[63]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n152 ) );
NAND2_X2 _AES_ENC_U212  ( .A1(_AES_ENC_text_in_r[63] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n153 ) );
NAND2_X2 _AES_ENC_U211  ( .A1(_AES_ENC_n152 ), .A2(_AES_ENC_n153 ), .ZN(_AES_ENC_n724 ) );
NAND2_X2 _AES_ENC_U210  ( .A1(aes_text_in[64]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n150 ) );
NAND2_X2 _AES_ENC_U209  ( .A1(_AES_ENC_text_in_r[64] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n151 ) );
NAND2_X2 _AES_ENC_U208  ( .A1(_AES_ENC_n150 ), .A2(_AES_ENC_n151 ), .ZN(_AES_ENC_n725 ) );
NAND2_X2 _AES_ENC_U207  ( .A1(aes_text_in[65]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n1480 ) );
NAND2_X2 _AES_ENC_U206  ( .A1(_AES_ENC_text_in_r[65] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1490 ) );
NAND2_X2 _AES_ENC_U205  ( .A1(_AES_ENC_n1480 ), .A2(_AES_ENC_n1490 ), .ZN(_AES_ENC_n726 ) );
NAND2_X2 _AES_ENC_U204  ( .A1(aes_text_in[66]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n1460 ) );
NAND2_X2 _AES_ENC_U203  ( .A1(_AES_ENC_text_in_r[66] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1470 ) );
NAND2_X2 _AES_ENC_U202  ( .A1(_AES_ENC_n1460 ), .A2(_AES_ENC_n1470 ), .ZN(_AES_ENC_n727 ) );
NAND2_X2 _AES_ENC_U201  ( .A1(aes_text_in[67]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n1440 ) );
NAND2_X2 _AES_ENC_U200  ( .A1(_AES_ENC_text_in_r[67] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1450 ) );
NAND2_X2 _AES_ENC_U199  ( .A1(_AES_ENC_n1440 ), .A2(_AES_ENC_n1450 ), .ZN(_AES_ENC_n728 ) );
NAND2_X2 _AES_ENC_U198  ( .A1(aes_text_in[68]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n1420 ) );
NAND2_X2 _AES_ENC_U197  ( .A1(_AES_ENC_text_in_r[68] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1430 ) );
NAND2_X2 _AES_ENC_U196  ( .A1(_AES_ENC_n1420 ), .A2(_AES_ENC_n1430 ), .ZN(_AES_ENC_n729 ) );
NAND2_X2 _AES_ENC_U195  ( .A1(aes_text_in[69]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n140 ) );
NAND2_X2 _AES_ENC_U194  ( .A1(_AES_ENC_text_in_r[69] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n141 ) );
NAND2_X2 _AES_ENC_U193  ( .A1(_AES_ENC_n140 ), .A2(_AES_ENC_n141 ), .ZN(_AES_ENC_n730 ) );
NAND2_X2 _AES_ENC_U192  ( .A1(aes_text_in[70]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n138 ) );
NAND2_X2 _AES_ENC_U191  ( .A1(_AES_ENC_text_in_r[70] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n139 ) );
NAND2_X2 _AES_ENC_U190  ( .A1(_AES_ENC_n138 ), .A2(_AES_ENC_n139 ), .ZN(_AES_ENC_n731 ) );
NAND2_X2 _AES_ENC_U189  ( .A1(aes_text_in[71]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n136 ) );
NAND2_X2 _AES_ENC_U188  ( .A1(_AES_ENC_text_in_r[71] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n137 ) );
NAND2_X2 _AES_ENC_U187  ( .A1(_AES_ENC_n136 ), .A2(_AES_ENC_n137 ), .ZN(_AES_ENC_n732 ) );
NAND2_X2 _AES_ENC_U186  ( .A1(aes_text_in[72]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n134 ) );
NAND2_X2 _AES_ENC_U185  ( .A1(_AES_ENC_text_in_r[72] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n135 ) );
NAND2_X2 _AES_ENC_U184  ( .A1(_AES_ENC_n134 ), .A2(_AES_ENC_n135 ), .ZN(_AES_ENC_n733 ) );
NAND2_X2 _AES_ENC_U183  ( .A1(aes_text_in[73]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n1320 ) );
NAND2_X2 _AES_ENC_U182  ( .A1(_AES_ENC_text_in_r[73] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1330 ) );
NAND2_X2 _AES_ENC_U181  ( .A1(_AES_ENC_n1320 ), .A2(_AES_ENC_n1330 ), .ZN(_AES_ENC_n734 ) );
NAND2_X2 _AES_ENC_U180  ( .A1(aes_text_in[74]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n1300 ) );
NAND2_X2 _AES_ENC_U179  ( .A1(_AES_ENC_text_in_r[74] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1310 ) );
NAND2_X2 _AES_ENC_U178  ( .A1(_AES_ENC_n1300 ), .A2(_AES_ENC_n1310 ), .ZN(_AES_ENC_n735 ) );
NAND2_X2 _AES_ENC_U177  ( .A1(aes_text_in[75]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n1280 ) );
NAND2_X2 _AES_ENC_U176  ( .A1(_AES_ENC_text_in_r[75] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1290 ) );
NAND2_X2 _AES_ENC_U175  ( .A1(_AES_ENC_n1280 ), .A2(_AES_ENC_n1290 ), .ZN(_AES_ENC_n736 ) );
NAND2_X2 _AES_ENC_U174  ( .A1(aes_text_in[76]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n12600 ) );
NAND2_X2 _AES_ENC_U173  ( .A1(_AES_ENC_text_in_r[76] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n1270 ) );
NAND2_X2 _AES_ENC_U172  ( .A1(_AES_ENC_n12600 ), .A2(_AES_ENC_n1270 ), .ZN(_AES_ENC_n737 ) );
NAND2_X2 _AES_ENC_U171  ( .A1(aes_text_in[77]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n124 ) );
NAND2_X2 _AES_ENC_U170  ( .A1(_AES_ENC_text_in_r[77] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n125 ) );
NAND2_X2 _AES_ENC_U169  ( .A1(_AES_ENC_n124 ), .A2(_AES_ENC_n125 ), .ZN(_AES_ENC_n738 ) );
NAND2_X2 _AES_ENC_U168  ( .A1(aes_text_in[78]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n122 ) );
NAND2_X2 _AES_ENC_U167  ( .A1(_AES_ENC_text_in_r[78] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n123 ) );
NAND2_X2 _AES_ENC_U166  ( .A1(_AES_ENC_n122 ), .A2(_AES_ENC_n123 ), .ZN(_AES_ENC_n739 ) );
NAND2_X2 _AES_ENC_U165  ( .A1(aes_text_in[79]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n120 ) );
NAND2_X2 _AES_ENC_U164  ( .A1(_AES_ENC_text_in_r[79] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n121 ) );
NAND2_X2 _AES_ENC_U163  ( .A1(_AES_ENC_n120 ), .A2(_AES_ENC_n121 ), .ZN(_AES_ENC_n740 ) );
NAND2_X2 _AES_ENC_U162  ( .A1(aes_text_in[80]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n118 ) );
NAND2_X2 _AES_ENC_U161  ( .A1(_AES_ENC_text_in_r[80] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n119 ) );
NAND2_X2 _AES_ENC_U160  ( .A1(_AES_ENC_n118 ), .A2(_AES_ENC_n119 ), .ZN(_AES_ENC_n741 ) );
NAND2_X2 _AES_ENC_U159  ( .A1(aes_text_in[81]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n11610 ) );
NAND2_X2 _AES_ENC_U158  ( .A1(_AES_ENC_text_in_r[81] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n11710 ) );
NAND2_X2 _AES_ENC_U157  ( .A1(_AES_ENC_n11610 ), .A2(_AES_ENC_n11710 ), .ZN(_AES_ENC_n742 ) );
NAND2_X2 _AES_ENC_U156  ( .A1(aes_text_in[82]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n11410 ) );
NAND2_X2 _AES_ENC_U155  ( .A1(_AES_ENC_text_in_r[82] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n11510 ) );
NAND2_X2 _AES_ENC_U154  ( .A1(_AES_ENC_n11410 ), .A2(_AES_ENC_n11510 ), .ZN(_AES_ENC_n743 ) );
NAND2_X2 _AES_ENC_U153  ( .A1(aes_text_in[83]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n11210 ) );
NAND2_X2 _AES_ENC_U152  ( .A1(_AES_ENC_text_in_r[83] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n11310 ) );
NAND2_X2 _AES_ENC_U151  ( .A1(_AES_ENC_n11210 ), .A2(_AES_ENC_n11310 ), .ZN(_AES_ENC_n744 ) );
NAND2_X2 _AES_ENC_U150  ( .A1(aes_text_in[84]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n11010 ) );
NAND2_X2 _AES_ENC_U149  ( .A1(_AES_ENC_text_in_r[84] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n11110 ) );
NAND2_X2 _AES_ENC_U148  ( .A1(_AES_ENC_n11010 ), .A2(_AES_ENC_n11110 ), .ZN(_AES_ENC_n745 ) );
NAND2_X2 _AES_ENC_U147  ( .A1(aes_text_in[85]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n108 ) );
NAND2_X2 _AES_ENC_U146  ( .A1(_AES_ENC_text_in_r[85] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n109 ) );
NAND2_X2 _AES_ENC_U145  ( .A1(_AES_ENC_n108 ), .A2(_AES_ENC_n109 ), .ZN(_AES_ENC_n746 ) );
NAND2_X2 _AES_ENC_U144  ( .A1(aes_text_in[86]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n106 ) );
NAND2_X2 _AES_ENC_U143  ( .A1(_AES_ENC_text_in_r[86] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n107 ) );
NAND2_X2 _AES_ENC_U142  ( .A1(_AES_ENC_n106 ), .A2(_AES_ENC_n107 ), .ZN(_AES_ENC_n747 ) );
NAND2_X2 _AES_ENC_U141  ( .A1(aes_text_in[87]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n104 ) );
NAND2_X2 _AES_ENC_U140  ( .A1(_AES_ENC_text_in_r[87] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n105 ) );
NAND2_X2 _AES_ENC_U139  ( .A1(_AES_ENC_n104 ), .A2(_AES_ENC_n105 ), .ZN(_AES_ENC_n748 ) );
NAND2_X2 _AES_ENC_U138  ( .A1(aes_text_in[88]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n102 ) );
NAND2_X2 _AES_ENC_U137  ( .A1(_AES_ENC_text_in_r[88] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n103 ) );
NAND2_X2 _AES_ENC_U136  ( .A1(_AES_ENC_n102 ), .A2(_AES_ENC_n103 ), .ZN(_AES_ENC_n749 ) );
NAND2_X2 _AES_ENC_U135  ( .A1(aes_text_in[89]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n10010 ) );
NAND2_X2 _AES_ENC_U134  ( .A1(_AES_ENC_text_in_r[89] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n10110 ) );
NAND2_X2 _AES_ENC_U133  ( .A1(_AES_ENC_n10010 ), .A2(_AES_ENC_n10110 ), .ZN(_AES_ENC_n750 ) );
NAND2_X2 _AES_ENC_U132  ( .A1(aes_text_in[90]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n9810 ) );
NAND2_X2 _AES_ENC_U131  ( .A1(_AES_ENC_text_in_r[90] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n9910 ) );
NAND2_X2 _AES_ENC_U130  ( .A1(_AES_ENC_n9810 ), .A2(_AES_ENC_n9910 ), .ZN(_AES_ENC_n751 ) );
NAND2_X2 _AES_ENC_U129  ( .A1(aes_text_in[91]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n9610 ) );
NAND2_X2 _AES_ENC_U128  ( .A1(_AES_ENC_text_in_r[91] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n9710 ) );
NAND2_X2 _AES_ENC_U127  ( .A1(_AES_ENC_n9610 ), .A2(_AES_ENC_n9710 ), .ZN(_AES_ENC_n752 ) );
NAND2_X2 _AES_ENC_U126  ( .A1(aes_text_in[92]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n9410 ) );
NAND2_X2 _AES_ENC_U125  ( .A1(_AES_ENC_text_in_r[92] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n9510 ) );
NAND2_X2 _AES_ENC_U124  ( .A1(_AES_ENC_n9410 ), .A2(_AES_ENC_n9510 ), .ZN(_AES_ENC_n753 ) );
NAND2_X2 _AES_ENC_U123  ( .A1(aes_text_in[93]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n92 ) );
NAND2_X2 _AES_ENC_U122  ( .A1(_AES_ENC_text_in_r[93] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n93 ) );
NAND2_X2 _AES_ENC_U121  ( .A1(_AES_ENC_n92 ), .A2(_AES_ENC_n93 ), .ZN(_AES_ENC_n754 ) );
NAND2_X2 _AES_ENC_U120  ( .A1(aes_text_in[94]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n90 ) );
NAND2_X2 _AES_ENC_U119  ( .A1(_AES_ENC_text_in_r[94] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n91 ) );
NAND2_X2 _AES_ENC_U118  ( .A1(_AES_ENC_n90 ), .A2(_AES_ENC_n91 ), .ZN(_AES_ENC_n755 ) );
NAND2_X2 _AES_ENC_U117  ( .A1(aes_text_in[95]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n88 ) );
NAND2_X2 _AES_ENC_U116  ( .A1(_AES_ENC_text_in_r[95] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n89 ) );
NAND2_X2 _AES_ENC_U115  ( .A1(_AES_ENC_n88 ), .A2(_AES_ENC_n89 ), .ZN(_AES_ENC_n756 ) );
NAND2_X2 _AES_ENC_U114  ( .A1(aes_text_in[96]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n86 ) );
NAND2_X2 _AES_ENC_U113  ( .A1(_AES_ENC_text_in_r[96] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n87 ) );
NAND2_X2 _AES_ENC_U112  ( .A1(_AES_ENC_n86 ), .A2(_AES_ENC_n87 ), .ZN(_AES_ENC_n757 ) );
NAND2_X2 _AES_ENC_U111  ( .A1(aes_text_in[97]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n8410 ) );
NAND2_X2 _AES_ENC_U110  ( .A1(_AES_ENC_text_in_r[97] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n8510 ) );
NAND2_X2 _AES_ENC_U109  ( .A1(_AES_ENC_n8410 ), .A2(_AES_ENC_n8510 ), .ZN(_AES_ENC_n758 ) );
NAND2_X2 _AES_ENC_U108  ( .A1(aes_text_in[98]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n8210 ) );
NAND2_X2 _AES_ENC_U107  ( .A1(_AES_ENC_text_in_r[98] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n8310 ) );
NAND2_X2 _AES_ENC_U106  ( .A1(_AES_ENC_n8210 ), .A2(_AES_ENC_n8310 ), .ZN(_AES_ENC_n759 ) );
NAND2_X2 _AES_ENC_U105  ( .A1(aes_text_in[99]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n8010 ) );
NAND2_X2 _AES_ENC_U104  ( .A1(_AES_ENC_text_in_r[99] ), .A2(_AES_ENC_n1261 ),.ZN(_AES_ENC_n8110 ) );
NAND2_X2 _AES_ENC_U103  ( .A1(_AES_ENC_n8010 ), .A2(_AES_ENC_n8110 ), .ZN(_AES_ENC_n760 ) );
NAND2_X2 _AES_ENC_U102  ( .A1(aes_text_in[100]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n7890 ) );
NAND2_X2 _AES_ENC_U101  ( .A1(_AES_ENC_text_in_r[100] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n7900 ) );
NAND2_X2 _AES_ENC_U100  ( .A1(_AES_ENC_n7890 ), .A2(_AES_ENC_n7900 ), .ZN(_AES_ENC_n761 ) );
NAND2_X2 _AES_ENC_U99  ( .A1(aes_text_in[101]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n76 ) );
NAND2_X2 _AES_ENC_U98  ( .A1(_AES_ENC_text_in_r[101] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n77 ) );
NAND2_X2 _AES_ENC_U97  ( .A1(_AES_ENC_n76 ), .A2(_AES_ENC_n77 ), .ZN(_AES_ENC_n762 ) );
NAND2_X2 _AES_ENC_U96  ( .A1(aes_text_in[102]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n74 ) );
NAND2_X2 _AES_ENC_U95  ( .A1(_AES_ENC_text_in_r[102] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n75 ) );
NAND2_X2 _AES_ENC_U94  ( .A1(_AES_ENC_n74 ), .A2(_AES_ENC_n75 ), .ZN(_AES_ENC_n763 ) );
NAND2_X2 _AES_ENC_U93  ( .A1(aes_text_in[103]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n72 ) );
NAND2_X2 _AES_ENC_U92  ( .A1(_AES_ENC_text_in_r[103] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n73 ) );
NAND2_X2 _AES_ENC_U91  ( .A1(_AES_ENC_n72 ), .A2(_AES_ENC_n73 ), .ZN(_AES_ENC_n764 ) );
NAND2_X2 _AES_ENC_U90  ( .A1(aes_text_in[104]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n70 ) );
NAND2_X2 _AES_ENC_U89  ( .A1(_AES_ENC_text_in_r[104] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n71 ) );
NAND2_X2 _AES_ENC_U88  ( .A1(_AES_ENC_n70 ), .A2(_AES_ENC_n71 ), .ZN(_AES_ENC_n765 ) );
NAND2_X2 _AES_ENC_U87  ( .A1(aes_text_in[105]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n6810 ) );
NAND2_X2 _AES_ENC_U86  ( .A1(_AES_ENC_text_in_r[105] ), .A2(_AES_ENC_n12601 ), .ZN(_AES_ENC_n6910 ) );
NAND2_X2 _AES_ENC_U85  ( .A1(_AES_ENC_n6810 ), .A2(_AES_ENC_n6910 ), .ZN(_AES_ENC_n766 ) );
NAND2_X2 _AES_ENC_U84  ( .A1(aes_text_in[106]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n6600 ) );
NAND2_X2 _AES_ENC_U83  ( .A1(_AES_ENC_text_in_r[106] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n6710 ) );
NAND2_X2 _AES_ENC_U82  ( .A1(_AES_ENC_n6600 ), .A2(_AES_ENC_n6710 ), .ZN(_AES_ENC_n767 ) );
NAND2_X2 _AES_ENC_U81  ( .A1(aes_text_in[107]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n6400 ) );
NAND2_X2 _AES_ENC_U80  ( .A1(_AES_ENC_text_in_r[107] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n6500 ) );
NAND2_X2 _AES_ENC_U79  ( .A1(_AES_ENC_n6400 ), .A2(_AES_ENC_n6500 ), .ZN(_AES_ENC_n768 ) );
NAND2_X2 _AES_ENC_U78  ( .A1(aes_text_in[108]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n6200 ) );
NAND2_X2 _AES_ENC_U77  ( .A1(_AES_ENC_text_in_r[108] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n6300 ) );
NAND2_X2 _AES_ENC_U76  ( .A1(_AES_ENC_n6200 ), .A2(_AES_ENC_n6300 ), .ZN(_AES_ENC_n769 ) );
NAND2_X2 _AES_ENC_U75  ( .A1(aes_text_in[109]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n60 ) );
NAND2_X2 _AES_ENC_U74  ( .A1(_AES_ENC_text_in_r[109] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n61 ) );
NAND2_X2 _AES_ENC_U73  ( .A1(_AES_ENC_n60 ), .A2(_AES_ENC_n61 ), .ZN(_AES_ENC_n770 ) );
NAND2_X2 _AES_ENC_U72  ( .A1(aes_text_in[110]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n58 ) );
NAND2_X2 _AES_ENC_U71  ( .A1(_AES_ENC_text_in_r[110] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n59 ) );
NAND2_X2 _AES_ENC_U70  ( .A1(_AES_ENC_n58 ), .A2(_AES_ENC_n59 ), .ZN(_AES_ENC_n771 ) );
NAND2_X2 _AES_ENC_U69  ( .A1(aes_text_in[111]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n56 ) );
NAND2_X2 _AES_ENC_U68  ( .A1(_AES_ENC_text_in_r[111] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n57 ) );
NAND2_X2 _AES_ENC_U67  ( .A1(_AES_ENC_n56 ), .A2(_AES_ENC_n57 ), .ZN(_AES_ENC_n772 ) );
NAND2_X2 _AES_ENC_U66  ( .A1(aes_text_in[112]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n54 ) );
NAND2_X2 _AES_ENC_U65  ( .A1(_AES_ENC_text_in_r[112] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n55 ) );
NAND2_X2 _AES_ENC_U64  ( .A1(_AES_ENC_n54 ), .A2(_AES_ENC_n55 ), .ZN(_AES_ENC_n773 ) );
NAND2_X2 _AES_ENC_U63  ( .A1(aes_text_in[113]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n5200 ) );
NAND2_X2 _AES_ENC_U62  ( .A1(_AES_ENC_text_in_r[113] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n5300 ) );
NAND2_X2 _AES_ENC_U61  ( .A1(_AES_ENC_n5200 ), .A2(_AES_ENC_n5300 ), .ZN(_AES_ENC_n774 ) );
NAND2_X2 _AES_ENC_U60  ( .A1(aes_text_in[114]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n5020 ) );
NAND2_X2 _AES_ENC_U59  ( .A1(_AES_ENC_text_in_r[114] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n5100 ) );
NAND2_X2 _AES_ENC_U58  ( .A1(_AES_ENC_n5020 ), .A2(_AES_ENC_n5100 ), .ZN(_AES_ENC_n775 ) );
NAND2_X2 _AES_ENC_U57  ( .A1(aes_text_in[115]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n4810 ) );
NAND2_X2 _AES_ENC_U56  ( .A1(_AES_ENC_text_in_r[115] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n4910 ) );
NAND2_X2 _AES_ENC_U55  ( .A1(_AES_ENC_n4810 ), .A2(_AES_ENC_n4910 ), .ZN(_AES_ENC_n776 ) );
NAND2_X2 _AES_ENC_U54  ( .A1(aes_text_in[116]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n4610 ) );
NAND2_X2 _AES_ENC_U53  ( .A1(_AES_ENC_text_in_r[116] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n4710 ) );
NAND2_X2 _AES_ENC_U52  ( .A1(_AES_ENC_n4610 ), .A2(_AES_ENC_n4710 ), .ZN(_AES_ENC_n777 ) );
NAND2_X2 _AES_ENC_U51  ( .A1(aes_text_in[117]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n44 ) );
NAND2_X2 _AES_ENC_U50  ( .A1(_AES_ENC_text_in_r[117] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n45 ) );
NAND2_X2 _AES_ENC_U49  ( .A1(_AES_ENC_n44 ), .A2(_AES_ENC_n45 ), .ZN(_AES_ENC_n778 ) );
NAND2_X2 _AES_ENC_U48  ( .A1(aes_text_in[118]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n42 ) );
NAND2_X2 _AES_ENC_U47  ( .A1(_AES_ENC_text_in_r[118] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n43 ) );
NAND2_X2 _AES_ENC_U46  ( .A1(_AES_ENC_n42 ), .A2(_AES_ENC_n43 ), .ZN(_AES_ENC_n779 ) );
NAND2_X2 _AES_ENC_U45  ( .A1(aes_text_in[119]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n40 ) );
NAND2_X2 _AES_ENC_U44  ( .A1(_AES_ENC_text_in_r[119] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n41 ) );
NAND2_X2 _AES_ENC_U43  ( .A1(_AES_ENC_n40 ), .A2(_AES_ENC_n41 ), .ZN(_AES_ENC_n780 ) );
NAND2_X2 _AES_ENC_U42  ( .A1(aes_text_in[120]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n38 ) );
NAND2_X2 _AES_ENC_U41  ( .A1(_AES_ENC_text_in_r[120] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n39 ) );
NAND2_X2 _AES_ENC_U40  ( .A1(_AES_ENC_n38 ), .A2(_AES_ENC_n39 ), .ZN(_AES_ENC_n781 ) );
NAND2_X2 _AES_ENC_U39  ( .A1(aes_text_in[121]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n3600 ) );
NAND2_X2 _AES_ENC_U38  ( .A1(_AES_ENC_text_in_r[121] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n3700 ) );
NAND2_X2 _AES_ENC_U37  ( .A1(_AES_ENC_n3600 ), .A2(_AES_ENC_n3700 ), .ZN(_AES_ENC_n782 ) );
NAND2_X2 _AES_ENC_U36  ( .A1(aes_text_in[122]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n3400 ) );
NAND2_X2 _AES_ENC_U35  ( .A1(_AES_ENC_text_in_r[122] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n3500 ) );
NAND2_X2 _AES_ENC_U34  ( .A1(_AES_ENC_n3400 ), .A2(_AES_ENC_n3500 ), .ZN(_AES_ENC_n783 ) );
NAND2_X2 _AES_ENC_U33  ( .A1(aes_text_in[123]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n3200 ) );
NAND2_X2 _AES_ENC_U32  ( .A1(_AES_ENC_text_in_r[123] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n3300 ) );
NAND2_X2 _AES_ENC_U31  ( .A1(_AES_ENC_n3200 ), .A2(_AES_ENC_n3300 ), .ZN(_AES_ENC_n784 ) );
NAND2_X2 _AES_ENC_U30  ( .A1(aes_text_in[124]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n3000 ) );
NAND2_X2 _AES_ENC_U29  ( .A1(_AES_ENC_text_in_r[124] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n3100 ) );
NAND2_X2 _AES_ENC_U28  ( .A1(_AES_ENC_n3000 ), .A2(_AES_ENC_n3100 ), .ZN(_AES_ENC_n785 ) );
NAND2_X2 _AES_ENC_U27  ( .A1(aes_text_in[125]), .A2(_AES_ENC_n1235 ), .ZN(_AES_ENC_n28 ) );
NAND2_X2 _AES_ENC_U26  ( .A1(_AES_ENC_text_in_r[125] ), .A2(_AES_ENC_n1259 ),.ZN(_AES_ENC_n29 ) );
NAND2_X2 _AES_ENC_U25  ( .A1(_AES_ENC_n28 ), .A2(_AES_ENC_n29 ), .ZN(_AES_ENC_n786 ) );
NAND2_X2 _AES_ENC_U24  ( .A1(aes_text_in[126]), .A2(_AES_ENC_n1236 ), .ZN(_AES_ENC_n26 ) );
NAND2_X2 _AES_ENC_U23  ( .A1(_AES_ENC_text_in_r[126] ), .A2(_AES_ENC_n1258 ),.ZN(_AES_ENC_n27 ) );
NAND2_X2 _AES_ENC_U22  ( .A1(_AES_ENC_n26 ), .A2(_AES_ENC_n27 ), .ZN(_AES_ENC_n787 ) );
NAND2_X2 _AES_ENC_U21  ( .A1(aes_text_in[127]), .A2(_AES_ENC_n1237 ), .ZN(_AES_ENC_n24 ) );
NAND2_X2 _AES_ENC_U20  ( .A1(_AES_ENC_text_in_r[127] ), .A2(_AES_ENC_n1258 ),.ZN(_AES_ENC_n25 ) );
NAND2_X2 _AES_ENC_U19  ( .A1(_AES_ENC_n24 ), .A2(_AES_ENC_n25 ), .ZN(_AES_ENC_n788 ) );
NAND2_X2 _AES_ENC_U18  ( .A1(_AES_ENC_n792 ), .A2(_AES_ENC_n14 ), .ZN(_AES_ENC_n23 ) );
NAND2_X2 _AES_ENC_U17  ( .A1(_AES_ENC_n1258 ), .A2(_AES_ENC_n23 ), .ZN(_AES_ENC_n22 ) );
NAND2_X2 _AES_ENC_U15  ( .A1(_AES_ENC_n11 ), .A2(_AES_ENC_n14 ), .ZN(_AES_ENC_n18 ) );
NAND2_X2 _AES_ENC_U13  ( .A1(_AES_ENC_n1258 ), .A2(_AES_ENC_n1231 ), .ZN(_AES_ENC_n21 ) );
NAND2_X2 _AES_ENC_U12  ( .A1(_AES_ENC_n1266 ), .A2(_AES_ENC_n21 ), .ZN(_AES_ENC_n20 ) );
NAND2_X2 _AES_ENC_U11  ( .A1(_AES_ENC_n20 ), .A2(_AES_ENC_n1234 ), .ZN(_AES_ENC_n1980 ) );
NAND2_X2 _AES_ENC_U10  ( .A1(_AES_ENC_n18 ), .A2(_AES_ENC_n1980 ), .ZN(_AES_ENC_n795 ) );
NAND2_X2 _AES_ENC_U9  ( .A1(_AES_ENC_n17 ), .A2(_AES_ENC_n1231 ), .ZN(_AES_ENC_n15 ) );
NAND2_X2 _AES_ENC_U8  ( .A1(_AES_ENC_n11 ), .A2(_AES_ENC_n794 ), .ZN(_AES_ENC_n16 ) );
NAND2_X2 _AES_ENC_U6  ( .A1(_AES_ENC_n14 ), .A2(_AES_ENC_n1266 ), .ZN(_AES_ENC_n13 ) );
NAND2_X2 _AES_ENC_U5  ( .A1(_AES_ENC_n13 ), .A2(_AES_ENC_n1233 ), .ZN(_AES_ENC_n12 ) );
NAND2_X2 _AES_ENC_U4  ( .A1(_AES_ENC_n1258 ), .A2(_AES_ENC_n12 ), .ZN(_AES_ENC_n797 ) );
OR2_X2 _AES_ENC_U3  ( .A1(_AES_ENC_n1257 ), .A2(_AES_ENC_n11 ), .ZN(_AES_ENC_n798 ) );
CLKBUFX1 gbuf_d_781(.A(_AES_ENC_N501), .Y(ddout__781));
CLKBUFX1 gbuf_q_781(.A(qq_in781), .Y(aes_text_out[0]));
CLKBUFX1 gbuf_d_782(.A(_AES_ENC_N500), .Y(ddout__782));
CLKBUFX1 gbuf_q_782(.A(qq_in782), .Y(aes_text_out[1]));
CLKBUFX1 gbuf_d_783(.A(_AES_ENC_N499), .Y(ddout__783));
CLKBUFX1 gbuf_q_783(.A(qq_in783), .Y(aes_text_out[2]));
CLKBUFX1 gbuf_d_784(.A(_AES_ENC_N498), .Y(ddout__784));
CLKBUFX1 gbuf_q_784(.A(qq_in784), .Y(aes_text_out[3]));
CLKBUFX1 gbuf_d_785(.A(_AES_ENC_N497), .Y(ddout__785));
CLKBUFX1 gbuf_q_785(.A(qq_in785), .Y(aes_text_out[4]));
CLKBUFX1 gbuf_d_786(.A(_AES_ENC_N496), .Y(ddout__786));
CLKBUFX1 gbuf_q_786(.A(qq_in786), .Y(aes_text_out[5]));
CLKBUFX1 gbuf_d_787(.A(_AES_ENC_N495), .Y(ddout__787));
CLKBUFX1 gbuf_q_787(.A(qq_in787), .Y(aes_text_out[6]));
CLKBUFX1 gbuf_d_788(.A(_AES_ENC_N494), .Y(ddout__788));
CLKBUFX1 gbuf_q_788(.A(qq_in788), .Y(aes_text_out[7]));
CLKBUFX1 gbuf_d_789(.A(_AES_ENC_N469), .Y(ddout__789));
CLKBUFX1 gbuf_q_789(.A(qq_in789), .Y(aes_text_out[8]));
CLKBUFX1 gbuf_d_790(.A(_AES_ENC_N468), .Y(ddout__790));
CLKBUFX1 gbuf_q_790(.A(qq_in790), .Y(aes_text_out[9]));
CLKBUFX1 gbuf_d_791(.A(_AES_ENC_N467), .Y(ddout__791));
CLKBUFX1 gbuf_q_791(.A(qq_in791), .Y(aes_text_out[10]));
CLKBUFX1 gbuf_d_792(.A(_AES_ENC_N466), .Y(ddout__792));
CLKBUFX1 gbuf_q_792(.A(qq_in792), .Y(aes_text_out[11]));
CLKBUFX1 gbuf_d_793(.A(_AES_ENC_N465), .Y(ddout__793));
CLKBUFX1 gbuf_q_793(.A(qq_in793), .Y(aes_text_out[12]));
CLKBUFX1 gbuf_d_794(.A(_AES_ENC_N464), .Y(ddout__794));
CLKBUFX1 gbuf_q_794(.A(qq_in794), .Y(aes_text_out[13]));
CLKBUFX1 gbuf_d_795(.A(_AES_ENC_N463), .Y(ddout__795));
CLKBUFX1 gbuf_q_795(.A(qq_in795), .Y(aes_text_out[14]));
CLKBUFX1 gbuf_d_796(.A(_AES_ENC_N462), .Y(ddout__796));
CLKBUFX1 gbuf_q_796(.A(qq_in796), .Y(aes_text_out[15]));
CLKBUFX1 gbuf_d_797(.A(_AES_ENC_N437), .Y(ddout__797));
CLKBUFX1 gbuf_q_797(.A(qq_in797), .Y(aes_text_out[16]));
CLKBUFX1 gbuf_d_798(.A(_AES_ENC_N436), .Y(ddout__798));
CLKBUFX1 gbuf_q_798(.A(qq_in798), .Y(aes_text_out[17]));
CLKBUFX1 gbuf_d_799(.A(_AES_ENC_N435), .Y(ddout__799));
CLKBUFX1 gbuf_q_799(.A(qq_in799), .Y(aes_text_out[18]));
CLKBUFX1 gbuf_d_800(.A(_AES_ENC_N434), .Y(ddout__800));
CLKBUFX1 gbuf_q_800(.A(qq_in800), .Y(aes_text_out[19]));
CLKBUFX1 gbuf_d_801(.A(_AES_ENC_N433), .Y(ddout__801));
CLKBUFX1 gbuf_q_801(.A(qq_in801), .Y(aes_text_out[20]));
CLKBUFX1 gbuf_d_802(.A(_AES_ENC_N432), .Y(ddout__802));
CLKBUFX1 gbuf_q_802(.A(qq_in802), .Y(aes_text_out[21]));
CLKBUFX1 gbuf_d_803(.A(_AES_ENC_N431), .Y(ddout__803));
CLKBUFX1 gbuf_q_803(.A(qq_in803), .Y(aes_text_out[22]));
CLKBUFX1 gbuf_d_804(.A(_AES_ENC_N430), .Y(ddout__804));
CLKBUFX1 gbuf_q_804(.A(qq_in804), .Y(aes_text_out[23]));
CLKBUFX1 gbuf_d_805(.A(_AES_ENC_N405), .Y(ddout__805));
CLKBUFX1 gbuf_q_805(.A(qq_in805), .Y(aes_text_out[24]));
CLKBUFX1 gbuf_d_806(.A(_AES_ENC_N404), .Y(ddout__806));
CLKBUFX1 gbuf_q_806(.A(qq_in806), .Y(aes_text_out[25]));
CLKBUFX1 gbuf_d_807(.A(_AES_ENC_N403), .Y(ddout__807));
CLKBUFX1 gbuf_q_807(.A(qq_in807), .Y(aes_text_out[26]));
CLKBUFX1 gbuf_d_808(.A(_AES_ENC_N402), .Y(ddout__808));
CLKBUFX1 gbuf_q_808(.A(qq_in808), .Y(aes_text_out[27]));
CLKBUFX1 gbuf_d_809(.A(_AES_ENC_N401), .Y(ddout__809));
CLKBUFX1 gbuf_q_809(.A(qq_in809), .Y(aes_text_out[28]));
CLKBUFX1 gbuf_d_810(.A(_AES_ENC_N400), .Y(ddout__810));
CLKBUFX1 gbuf_q_810(.A(qq_in810), .Y(aes_text_out[29]));
CLKBUFX1 gbuf_d_811(.A(_AES_ENC_N399), .Y(ddout__811));
CLKBUFX1 gbuf_q_811(.A(qq_in811), .Y(aes_text_out[30]));
CLKBUFX1 gbuf_d_812(.A(_AES_ENC_N398), .Y(ddout__812));
CLKBUFX1 gbuf_q_812(.A(qq_in812), .Y(aes_text_out[31]));
CLKBUFX1 gbuf_d_813(.A(_AES_ENC_N493), .Y(ddout__813));
CLKBUFX1 gbuf_q_813(.A(qq_in813), .Y(aes_text_out[32]));
CLKBUFX1 gbuf_d_814(.A(_AES_ENC_N492), .Y(ddout__814));
CLKBUFX1 gbuf_q_814(.A(qq_in814), .Y(aes_text_out[33]));
CLKBUFX1 gbuf_d_815(.A(_AES_ENC_N491), .Y(ddout__815));
CLKBUFX1 gbuf_q_815(.A(qq_in815), .Y(aes_text_out[34]));
CLKBUFX1 gbuf_d_816(.A(_AES_ENC_N490), .Y(ddout__816));
CLKBUFX1 gbuf_q_816(.A(qq_in816), .Y(aes_text_out[35]));
CLKBUFX1 gbuf_d_817(.A(_AES_ENC_N489), .Y(ddout__817));
CLKBUFX1 gbuf_q_817(.A(qq_in817), .Y(aes_text_out[36]));
CLKBUFX1 gbuf_d_818(.A(_AES_ENC_N488), .Y(ddout__818));
CLKBUFX1 gbuf_q_818(.A(qq_in818), .Y(aes_text_out[37]));
CLKBUFX1 gbuf_d_819(.A(_AES_ENC_N487), .Y(ddout__819));
CLKBUFX1 gbuf_q_819(.A(qq_in819), .Y(aes_text_out[38]));
CLKBUFX1 gbuf_d_820(.A(_AES_ENC_N486), .Y(ddout__820));
CLKBUFX1 gbuf_q_820(.A(qq_in820), .Y(aes_text_out[39]));
CLKBUFX1 gbuf_d_821(.A(_AES_ENC_N461), .Y(ddout__821));
CLKBUFX1 gbuf_q_821(.A(qq_in821), .Y(aes_text_out[40]));
CLKBUFX1 gbuf_d_822(.A(_AES_ENC_N460), .Y(ddout__822));
CLKBUFX1 gbuf_q_822(.A(qq_in822), .Y(aes_text_out[41]));
CLKBUFX1 gbuf_d_823(.A(_AES_ENC_N459), .Y(ddout__823));
CLKBUFX1 gbuf_q_823(.A(qq_in823), .Y(aes_text_out[42]));
CLKBUFX1 gbuf_d_824(.A(_AES_ENC_N458), .Y(ddout__824));
CLKBUFX1 gbuf_q_824(.A(qq_in824), .Y(aes_text_out[43]));
CLKBUFX1 gbuf_d_825(.A(_AES_ENC_N457), .Y(ddout__825));
CLKBUFX1 gbuf_q_825(.A(qq_in825), .Y(aes_text_out[44]));
CLKBUFX1 gbuf_d_826(.A(_AES_ENC_N456), .Y(ddout__826));
CLKBUFX1 gbuf_q_826(.A(qq_in826), .Y(aes_text_out[45]));
CLKBUFX1 gbuf_d_827(.A(_AES_ENC_N455), .Y(ddout__827));
CLKBUFX1 gbuf_q_827(.A(qq_in827), .Y(aes_text_out[46]));
CLKBUFX1 gbuf_d_828(.A(_AES_ENC_N454), .Y(ddout__828));
CLKBUFX1 gbuf_q_828(.A(qq_in828), .Y(aes_text_out[47]));
CLKBUFX1 gbuf_d_829(.A(_AES_ENC_N429), .Y(ddout__829));
CLKBUFX1 gbuf_q_829(.A(qq_in829), .Y(aes_text_out[48]));
CLKBUFX1 gbuf_d_830(.A(_AES_ENC_N428), .Y(ddout__830));
CLKBUFX1 gbuf_q_830(.A(qq_in830), .Y(aes_text_out[49]));
CLKBUFX1 gbuf_d_831(.A(_AES_ENC_N427), .Y(ddout__831));
CLKBUFX1 gbuf_q_831(.A(qq_in831), .Y(aes_text_out[50]));
CLKBUFX1 gbuf_d_832(.A(_AES_ENC_N426), .Y(ddout__832));
CLKBUFX1 gbuf_q_832(.A(qq_in832), .Y(aes_text_out[51]));
CLKBUFX1 gbuf_d_833(.A(_AES_ENC_N425), .Y(ddout__833));
CLKBUFX1 gbuf_q_833(.A(qq_in833), .Y(aes_text_out[52]));
CLKBUFX1 gbuf_d_834(.A(_AES_ENC_N424), .Y(ddout__834));
CLKBUFX1 gbuf_q_834(.A(qq_in834), .Y(aes_text_out[53]));
CLKBUFX1 gbuf_d_835(.A(_AES_ENC_N423), .Y(ddout__835));
CLKBUFX1 gbuf_q_835(.A(qq_in835), .Y(aes_text_out[54]));
CLKBUFX1 gbuf_d_836(.A(_AES_ENC_N422), .Y(ddout__836));
CLKBUFX1 gbuf_q_836(.A(qq_in836), .Y(aes_text_out[55]));
CLKBUFX1 gbuf_d_837(.A(_AES_ENC_N397), .Y(ddout__837));
CLKBUFX1 gbuf_q_837(.A(qq_in837), .Y(aes_text_out[56]));
CLKBUFX1 gbuf_d_838(.A(_AES_ENC_N396), .Y(ddout__838));
CLKBUFX1 gbuf_q_838(.A(qq_in838), .Y(aes_text_out[57]));
CLKBUFX1 gbuf_d_839(.A(_AES_ENC_N395), .Y(ddout__839));
CLKBUFX1 gbuf_q_839(.A(qq_in839), .Y(aes_text_out[58]));
CLKBUFX1 gbuf_d_840(.A(_AES_ENC_N394), .Y(ddout__840));
CLKBUFX1 gbuf_q_840(.A(qq_in840), .Y(aes_text_out[59]));
CLKBUFX1 gbuf_d_841(.A(_AES_ENC_N393), .Y(ddout__841));
CLKBUFX1 gbuf_q_841(.A(qq_in841), .Y(aes_text_out[60]));
CLKBUFX1 gbuf_d_842(.A(_AES_ENC_N392), .Y(ddout__842));
CLKBUFX1 gbuf_q_842(.A(qq_in842), .Y(aes_text_out[61]));
CLKBUFX1 gbuf_d_843(.A(_AES_ENC_N391), .Y(ddout__843));
CLKBUFX1 gbuf_q_843(.A(qq_in843), .Y(aes_text_out[62]));
CLKBUFX1 gbuf_d_844(.A(_AES_ENC_N390), .Y(ddout__844));
CLKBUFX1 gbuf_q_844(.A(qq_in844), .Y(aes_text_out[63]));
CLKBUFX1 gbuf_d_845(.A(_AES_ENC_N485), .Y(ddout__845));
CLKBUFX1 gbuf_q_845(.A(qq_in845), .Y(aes_text_out[64]));
CLKBUFX1 gbuf_d_846(.A(_AES_ENC_N484), .Y(ddout__846));
CLKBUFX1 gbuf_q_846(.A(qq_in846), .Y(aes_text_out[65]));
CLKBUFX1 gbuf_d_847(.A(_AES_ENC_N483), .Y(ddout__847));
CLKBUFX1 gbuf_q_847(.A(qq_in847), .Y(aes_text_out[66]));
CLKBUFX1 gbuf_d_848(.A(_AES_ENC_N482), .Y(ddout__848));
CLKBUFX1 gbuf_q_848(.A(qq_in848), .Y(aes_text_out[67]));
CLKBUFX1 gbuf_d_849(.A(_AES_ENC_N481), .Y(ddout__849));
CLKBUFX1 gbuf_q_849(.A(qq_in849), .Y(aes_text_out[68]));
CLKBUFX1 gbuf_d_850(.A(_AES_ENC_N480), .Y(ddout__850));
CLKBUFX1 gbuf_q_850(.A(qq_in850), .Y(aes_text_out[69]));
CLKBUFX1 gbuf_d_851(.A(_AES_ENC_N479), .Y(ddout__851));
CLKBUFX1 gbuf_q_851(.A(qq_in851), .Y(aes_text_out[70]));
CLKBUFX1 gbuf_d_852(.A(_AES_ENC_N478), .Y(ddout__852));
CLKBUFX1 gbuf_q_852(.A(qq_in852), .Y(aes_text_out[71]));
CLKBUFX1 gbuf_d_853(.A(_AES_ENC_N453), .Y(ddout__853));
CLKBUFX1 gbuf_q_853(.A(qq_in853), .Y(aes_text_out[72]));
CLKBUFX1 gbuf_d_854(.A(_AES_ENC_N452), .Y(ddout__854));
CLKBUFX1 gbuf_q_854(.A(qq_in854), .Y(aes_text_out[73]));
CLKBUFX1 gbuf_d_855(.A(_AES_ENC_N451), .Y(ddout__855));
CLKBUFX1 gbuf_q_855(.A(qq_in855), .Y(aes_text_out[74]));
CLKBUFX1 gbuf_d_856(.A(_AES_ENC_N450), .Y(ddout__856));
CLKBUFX1 gbuf_q_856(.A(qq_in856), .Y(aes_text_out[75]));
CLKBUFX1 gbuf_d_857(.A(_AES_ENC_N449), .Y(ddout__857));
CLKBUFX1 gbuf_q_857(.A(qq_in857), .Y(aes_text_out[76]));
CLKBUFX1 gbuf_d_858(.A(_AES_ENC_N448), .Y(ddout__858));
CLKBUFX1 gbuf_q_858(.A(qq_in858), .Y(aes_text_out[77]));
CLKBUFX1 gbuf_d_859(.A(_AES_ENC_N447), .Y(ddout__859));
CLKBUFX1 gbuf_q_859(.A(qq_in859), .Y(aes_text_out[78]));
CLKBUFX1 gbuf_d_860(.A(_AES_ENC_N446), .Y(ddout__860));
CLKBUFX1 gbuf_q_860(.A(qq_in860), .Y(aes_text_out[79]));
CLKBUFX1 gbuf_d_861(.A(_AES_ENC_N421), .Y(ddout__861));
CLKBUFX1 gbuf_q_861(.A(qq_in861), .Y(aes_text_out[80]));
CLKBUFX1 gbuf_d_862(.A(_AES_ENC_N420), .Y(ddout__862));
CLKBUFX1 gbuf_q_862(.A(qq_in862), .Y(aes_text_out[81]));
CLKBUFX1 gbuf_d_863(.A(_AES_ENC_N419), .Y(ddout__863));
CLKBUFX1 gbuf_q_863(.A(qq_in863), .Y(aes_text_out[82]));
CLKBUFX1 gbuf_d_864(.A(_AES_ENC_N418), .Y(ddout__864));
CLKBUFX1 gbuf_q_864(.A(qq_in864), .Y(aes_text_out[83]));
CLKBUFX1 gbuf_d_865(.A(_AES_ENC_N417), .Y(ddout__865));
CLKBUFX1 gbuf_q_865(.A(qq_in865), .Y(aes_text_out[84]));
CLKBUFX1 gbuf_d_866(.A(_AES_ENC_N416), .Y(ddout__866));
CLKBUFX1 gbuf_q_866(.A(qq_in866), .Y(aes_text_out[85]));
CLKBUFX1 gbuf_d_867(.A(_AES_ENC_N415), .Y(ddout__867));
CLKBUFX1 gbuf_q_867(.A(qq_in867), .Y(aes_text_out[86]));
CLKBUFX1 gbuf_d_868(.A(_AES_ENC_N414), .Y(ddout__868));
CLKBUFX1 gbuf_q_868(.A(qq_in868), .Y(aes_text_out[87]));
CLKBUFX1 gbuf_d_869(.A(_AES_ENC_N389), .Y(ddout__869));
CLKBUFX1 gbuf_q_869(.A(qq_in869), .Y(aes_text_out[88]));
CLKBUFX1 gbuf_d_870(.A(_AES_ENC_N388), .Y(ddout__870));
CLKBUFX1 gbuf_q_870(.A(qq_in870), .Y(aes_text_out[89]));
CLKBUFX1 gbuf_d_871(.A(_AES_ENC_N387), .Y(ddout__871));
CLKBUFX1 gbuf_q_871(.A(qq_in871), .Y(aes_text_out[90]));
CLKBUFX1 gbuf_d_872(.A(_AES_ENC_N386), .Y(ddout__872));
CLKBUFX1 gbuf_q_872(.A(qq_in872), .Y(aes_text_out[91]));
CLKBUFX1 gbuf_d_873(.A(_AES_ENC_N385), .Y(ddout__873));
CLKBUFX1 gbuf_q_873(.A(qq_in873), .Y(aes_text_out[92]));
CLKBUFX1 gbuf_d_874(.A(_AES_ENC_N384), .Y(ddout__874));
CLKBUFX1 gbuf_q_874(.A(qq_in874), .Y(aes_text_out[93]));
CLKBUFX1 gbuf_d_875(.A(_AES_ENC_N383), .Y(ddout__875));
CLKBUFX1 gbuf_q_875(.A(qq_in875), .Y(aes_text_out[94]));
CLKBUFX1 gbuf_d_876(.A(_AES_ENC_N382), .Y(ddout__876));
CLKBUFX1 gbuf_q_876(.A(qq_in876), .Y(aes_text_out[95]));
CLKBUFX1 gbuf_d_877(.A(_AES_ENC_N477), .Y(ddout__877));
CLKBUFX1 gbuf_q_877(.A(qq_in877), .Y(aes_text_out[96]));
CLKBUFX1 gbuf_d_878(.A(_AES_ENC_N476), .Y(ddout__878));
CLKBUFX1 gbuf_q_878(.A(qq_in878), .Y(aes_text_out[97]));
CLKBUFX1 gbuf_d_879(.A(_AES_ENC_N475), .Y(ddout__879));
CLKBUFX1 gbuf_q_879(.A(qq_in879), .Y(aes_text_out[98]));
CLKBUFX1 gbuf_d_880(.A(_AES_ENC_N474), .Y(ddout__880));
CLKBUFX1 gbuf_q_880(.A(qq_in880), .Y(aes_text_out[99]));
CLKBUFX1 gbuf_d_881(.A(_AES_ENC_N473), .Y(ddout__881));
CLKBUFX1 gbuf_q_881(.A(qq_in881), .Y(aes_text_out[100]));
CLKBUFX1 gbuf_d_882(.A(_AES_ENC_N472), .Y(ddout__882));
CLKBUFX1 gbuf_q_882(.A(qq_in882), .Y(aes_text_out[101]));
CLKBUFX1 gbuf_d_883(.A(_AES_ENC_N471), .Y(ddout__883));
CLKBUFX1 gbuf_q_883(.A(qq_in883), .Y(aes_text_out[102]));
CLKBUFX1 gbuf_d_884(.A(_AES_ENC_N470), .Y(ddout__884));
CLKBUFX1 gbuf_q_884(.A(qq_in884), .Y(aes_text_out[103]));
CLKBUFX1 gbuf_d_885(.A(_AES_ENC_N445), .Y(ddout__885));
CLKBUFX1 gbuf_q_885(.A(qq_in885), .Y(aes_text_out[104]));
CLKBUFX1 gbuf_d_886(.A(_AES_ENC_N444), .Y(ddout__886));
CLKBUFX1 gbuf_q_886(.A(qq_in886), .Y(aes_text_out[105]));
CLKBUFX1 gbuf_d_887(.A(_AES_ENC_N443), .Y(ddout__887));
CLKBUFX1 gbuf_q_887(.A(qq_in887), .Y(aes_text_out[106]));
CLKBUFX1 gbuf_d_888(.A(_AES_ENC_N442), .Y(ddout__888));
CLKBUFX1 gbuf_q_888(.A(qq_in888), .Y(aes_text_out[107]));
CLKBUFX1 gbuf_d_889(.A(_AES_ENC_N441), .Y(ddout__889));
CLKBUFX1 gbuf_q_889(.A(qq_in889), .Y(aes_text_out[108]));
CLKBUFX1 gbuf_d_890(.A(_AES_ENC_N440), .Y(ddout__890));
CLKBUFX1 gbuf_q_890(.A(qq_in890), .Y(aes_text_out[109]));
CLKBUFX1 gbuf_d_891(.A(_AES_ENC_N439), .Y(ddout__891));
CLKBUFX1 gbuf_q_891(.A(qq_in891), .Y(aes_text_out[110]));
CLKBUFX1 gbuf_d_892(.A(_AES_ENC_N438), .Y(ddout__892));
CLKBUFX1 gbuf_q_892(.A(qq_in892), .Y(aes_text_out[111]));
CLKBUFX1 gbuf_d_893(.A(_AES_ENC_N413), .Y(ddout__893));
CLKBUFX1 gbuf_q_893(.A(qq_in893), .Y(aes_text_out[112]));
CLKBUFX1 gbuf_d_894(.A(_AES_ENC_N412), .Y(ddout__894));
CLKBUFX1 gbuf_q_894(.A(qq_in894), .Y(aes_text_out[113]));
CLKBUFX1 gbuf_d_895(.A(_AES_ENC_N411), .Y(ddout__895));
CLKBUFX1 gbuf_q_895(.A(qq_in895), .Y(aes_text_out[114]));
CLKBUFX1 gbuf_d_896(.A(_AES_ENC_N410), .Y(ddout__896));
CLKBUFX1 gbuf_q_896(.A(qq_in896), .Y(aes_text_out[115]));
CLKBUFX1 gbuf_d_897(.A(_AES_ENC_N409), .Y(ddout__897));
CLKBUFX1 gbuf_q_897(.A(qq_in897), .Y(aes_text_out[116]));
CLKBUFX1 gbuf_d_898(.A(_AES_ENC_N408), .Y(ddout__898));
CLKBUFX1 gbuf_q_898(.A(qq_in898), .Y(aes_text_out[117]));
CLKBUFX1 gbuf_d_899(.A(_AES_ENC_N407), .Y(ddout__899));
CLKBUFX1 gbuf_q_899(.A(qq_in899), .Y(aes_text_out[118]));
CLKBUFX1 gbuf_d_900(.A(_AES_ENC_N406), .Y(ddout__900));
CLKBUFX1 gbuf_q_900(.A(qq_in900), .Y(aes_text_out[119]));
CLKBUFX1 gbuf_d_901(.A(_AES_ENC_N381), .Y(ddout__901));
CLKBUFX1 gbuf_q_901(.A(qq_in901), .Y(aes_text_out[120]));
CLKBUFX1 gbuf_d_902(.A(_AES_ENC_N380), .Y(ddout__902));
CLKBUFX1 gbuf_q_902(.A(qq_in902), .Y(aes_text_out[121]));
CLKBUFX1 gbuf_d_903(.A(_AES_ENC_N379), .Y(ddout__903));
CLKBUFX1 gbuf_q_903(.A(qq_in903), .Y(aes_text_out[122]));
CLKBUFX1 gbuf_d_904(.A(_AES_ENC_N378), .Y(ddout__904));
CLKBUFX1 gbuf_q_904(.A(qq_in904), .Y(aes_text_out[123]));
CLKBUFX1 gbuf_d_905(.A(_AES_ENC_N377), .Y(ddout__905));
CLKBUFX1 gbuf_q_905(.A(qq_in905), .Y(aes_text_out[124]));
CLKBUFX1 gbuf_d_906(.A(_AES_ENC_N376), .Y(ddout__906));
CLKBUFX1 gbuf_q_906(.A(qq_in906), .Y(aes_text_out[125]));
CLKBUFX1 gbuf_d_907(.A(_AES_ENC_N375), .Y(ddout__907));
CLKBUFX1 gbuf_q_907(.A(qq_in907), .Y(aes_text_out[126]));
CLKBUFX1 gbuf_d_908(.A(_AES_ENC_N374), .Y(ddout__908));
CLKBUFX1 gbuf_q_908(.A(qq_in908), .Y(aes_text_out[127]));
CLKBUFX1 gbuf_d_909(.A(_AES_ENC_N101), .Y(ddout__909));
CLKBUFX1 gbuf_q_909(.A(qq_in909), .Y(_AES_ENC_sa32[7]));
CLKBUFX1 gbuf_d_910(.A(_AES_ENC_N229), .Y(ddout__910));
CLKBUFX1 gbuf_q_910(.A(qq_in910), .Y(_AES_ENC_sa30[7]));
CLKBUFX1 gbuf_d_911(.A(_AES_ENC_N238), .Y(ddout__911));
CLKBUFX1 gbuf_q_911(.A(qq_in911), .Y(_AES_ENC_sa20[0]));
CLKBUFX1 gbuf_d_912(.A(_AES_ENC_N239), .Y(ddout__912));
CLKBUFX1 gbuf_q_912(.A(qq_in912), .Y(_AES_ENC_sa20[1]));
CLKBUFX1 gbuf_d_913(.A(_AES_ENC_N241), .Y(ddout__913));
CLKBUFX1 gbuf_q_913(.A(qq_in913), .Y(_AES_ENC_sa20[3]));
CLKBUFX1 gbuf_d_914(.A(_AES_ENC_N242), .Y(ddout__914));
CLKBUFX1 gbuf_q_914(.A(qq_in914), .Y(_AES_ENC_sa20[4]));
CLKBUFX1 gbuf_d_915(.A(_AES_ENC_N261), .Y(ddout__915));
CLKBUFX1 gbuf_q_915(.A(qq_in915), .Y(_AES_ENC_sa10[7]));
CLKBUFX1 gbuf_d_916(.A(_AES_ENC_N277), .Y(ddout__916));
CLKBUFX1 gbuf_q_916(.A(qq_in916), .Y(_AES_ENC_sa00[7]));
CLKBUFX1 gbuf_d_917(.A(_AES_ENC_N228), .Y(ddout__917));
CLKBUFX1 gbuf_q_917(.A(qq_in917), .Y(_AES_ENC_sa30[6]));
CLKBUFX1 gbuf_d_918(.A(_AES_ENC_N260), .Y(ddout__918));
CLKBUFX1 gbuf_q_918(.A(qq_in918), .Y(_AES_ENC_sa10[6]));
CLKBUFX1 gbuf_d_919(.A(_AES_ENC_N276), .Y(ddout__919));
CLKBUFX1 gbuf_q_919(.A(qq_in919), .Y(_AES_ENC_sa00[6]));
CLKBUFX1 gbuf_d_920(.A(_AES_ENC_N227), .Y(ddout__920));
CLKBUFX1 gbuf_q_920(.A(qq_in920), .Y(_AES_ENC_sa30[5]));
CLKBUFX1 gbuf_d_921(.A(_AES_ENC_N244), .Y(ddout__921));
CLKBUFX1 gbuf_q_921(.A(qq_in921), .Y(_AES_ENC_sa20[6]));
CLKBUFX1 gbuf_d_922(.A(_AES_ENC_N259), .Y(ddout__922));
CLKBUFX1 gbuf_q_922(.A(qq_in922), .Y(_AES_ENC_sa10[5]));
CLKBUFX1 gbuf_d_923(.A(_AES_ENC_N275), .Y(ddout__923));
CLKBUFX1 gbuf_q_923(.A(qq_in923), .Y(_AES_ENC_sa00[5]));
CLKBUFX1 gbuf_d_924(.A(_AES_ENC_N226), .Y(ddout__924));
CLKBUFX1 gbuf_q_924(.A(qq_in924), .Y(_AES_ENC_sa30[4]));
CLKBUFX1 gbuf_d_925(.A(_AES_ENC_N243), .Y(ddout__925));
CLKBUFX1 gbuf_q_925(.A(qq_in925), .Y(_AES_ENC_sa20[5]));
CLKBUFX1 gbuf_d_926(.A(_AES_ENC_N258), .Y(ddout__926));
CLKBUFX1 gbuf_q_926(.A(qq_in926), .Y(_AES_ENC_sa10[4]));
CLKBUFX1 gbuf_d_927(.A(_AES_ENC_N274), .Y(ddout__927));
CLKBUFX1 gbuf_q_927(.A(qq_in927), .Y(_AES_ENC_sa00[4]));
CLKBUFX1 gbuf_d_928(.A(_AES_ENC_N225), .Y(ddout__928));
CLKBUFX1 gbuf_q_928(.A(qq_in928), .Y(_AES_ENC_sa30[3]));
CLKBUFX1 gbuf_d_929(.A(_AES_ENC_N257), .Y(ddout__929));
CLKBUFX1 gbuf_q_929(.A(qq_in929), .Y(_AES_ENC_sa10[3]));
CLKBUFX1 gbuf_d_930(.A(_AES_ENC_N273), .Y(ddout__930));
CLKBUFX1 gbuf_q_930(.A(qq_in930), .Y(_AES_ENC_sa00[3]));
CLKBUFX1 gbuf_d_931(.A(_AES_ENC_N224), .Y(ddout__931));
CLKBUFX1 gbuf_q_931(.A(qq_in931), .Y(_AES_ENC_sa30[2]));
CLKBUFX1 gbuf_d_932(.A(_AES_ENC_N256), .Y(ddout__932));
CLKBUFX1 gbuf_q_932(.A(qq_in932), .Y(_AES_ENC_sa10[2]));
CLKBUFX1 gbuf_d_933(.A(_AES_ENC_N272), .Y(ddout__933));
CLKBUFX1 gbuf_q_933(.A(qq_in933), .Y(_AES_ENC_sa00[2]));
CLKBUFX1 gbuf_d_934(.A(_AES_ENC_N223), .Y(ddout__934));
CLKBUFX1 gbuf_q_934(.A(qq_in934), .Y(_AES_ENC_sa30[1]));
CLKBUFX1 gbuf_d_935(.A(_AES_ENC_N240), .Y(ddout__935));
CLKBUFX1 gbuf_q_935(.A(qq_in935), .Y(_AES_ENC_sa20[2]));
CLKBUFX1 gbuf_d_936(.A(_AES_ENC_N255), .Y(ddout__936));
CLKBUFX1 gbuf_q_936(.A(qq_in936), .Y(_AES_ENC_sa10[1]));
CLKBUFX1 gbuf_d_937(.A(_AES_ENC_N271), .Y(ddout__937));
CLKBUFX1 gbuf_q_937(.A(qq_in937), .Y(_AES_ENC_sa00[1]));
CLKBUFX1 gbuf_d_938(.A(_AES_ENC_N117), .Y(ddout__938));
CLKBUFX1 gbuf_q_938(.A(qq_in938), .Y(_AES_ENC_sa22[7]));
CLKBUFX1 gbuf_d_939(.A(_AES_ENC_N133), .Y(ddout__939));
CLKBUFX1 gbuf_q_939(.A(qq_in939), .Y(_AES_ENC_sa12[7]));
CLKBUFX1 gbuf_d_940(.A(_AES_ENC_N132), .Y(ddout__940));
CLKBUFX1 gbuf_q_940(.A(qq_in940), .Y(_AES_ENC_sa12[6]));
CLKBUFX1 gbuf_d_941(.A(_AES_ENC_N100), .Y(ddout__941));
CLKBUFX1 gbuf_q_941(.A(qq_in941), .Y(_AES_ENC_sa32[6]));
CLKBUFX1 gbuf_d_942(.A(_AES_ENC_N116), .Y(ddout__942));
CLKBUFX1 gbuf_q_942(.A(qq_in942), .Y(_AES_ENC_sa22[6]));
CLKBUFX1 gbuf_d_943(.A(_AES_ENC_N149), .Y(ddout__943));
CLKBUFX1 gbuf_q_943(.A(qq_in943), .Y(_AES_ENC_sa02[7]));
CLKBUFX1 gbuf_d_944(.A(_AES_ENC_N131), .Y(ddout__944));
CLKBUFX1 gbuf_q_944(.A(qq_in944), .Y(_AES_ENC_sa12[5]));
CLKBUFX1 gbuf_d_945(.A(_AES_ENC_N99), .Y(ddout__945));
CLKBUFX1 gbuf_q_945(.A(qq_in945), .Y(_AES_ENC_sa32[5]));
CLKBUFX1 gbuf_d_946(.A(_AES_ENC_N115), .Y(ddout__946));
CLKBUFX1 gbuf_q_946(.A(qq_in946), .Y(_AES_ENC_sa22[5]));
CLKBUFX1 gbuf_d_947(.A(_AES_ENC_N148), .Y(ddout__947));
CLKBUFX1 gbuf_q_947(.A(qq_in947), .Y(_AES_ENC_sa02[6]));
CLKBUFX1 gbuf_d_948(.A(_AES_ENC_N130), .Y(ddout__948));
CLKBUFX1 gbuf_q_948(.A(qq_in948), .Y(_AES_ENC_sa12[4]));
CLKBUFX1 gbuf_d_949(.A(_AES_ENC_N98), .Y(ddout__949));
CLKBUFX1 gbuf_q_949(.A(qq_in949), .Y(_AES_ENC_sa32[4]));
CLKBUFX1 gbuf_d_950(.A(_AES_ENC_N114), .Y(ddout__950));
CLKBUFX1 gbuf_q_950(.A(qq_in950), .Y(_AES_ENC_sa22[4]));
CLKBUFX1 gbuf_d_951(.A(_AES_ENC_N147), .Y(ddout__951));
CLKBUFX1 gbuf_q_951(.A(qq_in951), .Y(_AES_ENC_sa02[5]));
CLKBUFX1 gbuf_d_952(.A(_AES_ENC_N129), .Y(ddout__952));
CLKBUFX1 gbuf_q_952(.A(qq_in952), .Y(_AES_ENC_sa12[3]));
CLKBUFX1 gbuf_d_953(.A(_AES_ENC_N97), .Y(ddout__953));
CLKBUFX1 gbuf_q_953(.A(qq_in953), .Y(_AES_ENC_sa32[3]));
CLKBUFX1 gbuf_d_954(.A(_AES_ENC_N113), .Y(ddout__954));
CLKBUFX1 gbuf_q_954(.A(qq_in954), .Y(_AES_ENC_sa22[3]));
CLKBUFX1 gbuf_d_955(.A(_AES_ENC_N146), .Y(ddout__955));
CLKBUFX1 gbuf_q_955(.A(qq_in955), .Y(_AES_ENC_sa02[4]));
CLKBUFX1 gbuf_d_956(.A(_AES_ENC_N128), .Y(ddout__956));
CLKBUFX1 gbuf_q_956(.A(qq_in956), .Y(_AES_ENC_sa12[2]));
CLKBUFX1 gbuf_d_957(.A(_AES_ENC_N96), .Y(ddout__957));
CLKBUFX1 gbuf_q_957(.A(qq_in957), .Y(_AES_ENC_sa32[2]));
CLKBUFX1 gbuf_d_958(.A(_AES_ENC_N112), .Y(ddout__958));
CLKBUFX1 gbuf_q_958(.A(qq_in958), .Y(_AES_ENC_sa22[2]));
CLKBUFX1 gbuf_d_959(.A(_AES_ENC_N145), .Y(ddout__959));
CLKBUFX1 gbuf_q_959(.A(qq_in959), .Y(_AES_ENC_sa02[3]));
CLKBUFX1 gbuf_d_960(.A(_AES_ENC_N127), .Y(ddout__960));
CLKBUFX1 gbuf_q_960(.A(qq_in960), .Y(_AES_ENC_sa12[1]));
CLKBUFX1 gbuf_d_961(.A(_AES_ENC_N95), .Y(ddout__961));
CLKBUFX1 gbuf_q_961(.A(qq_in961), .Y(_AES_ENC_sa32[1]));
CLKBUFX1 gbuf_d_962(.A(_AES_ENC_N111), .Y(ddout__962));
CLKBUFX1 gbuf_q_962(.A(qq_in962), .Y(_AES_ENC_sa22[1]));
CLKBUFX1 gbuf_d_963(.A(_AES_ENC_N144), .Y(ddout__963));
CLKBUFX1 gbuf_q_963(.A(qq_in963), .Y(_AES_ENC_sa02[2]));
CLKBUFX1 gbuf_d_964(.A(_AES_ENC_N110), .Y(ddout__964));
CLKBUFX1 gbuf_q_964(.A(qq_in964), .Y(_AES_ENC_sa22[0]));
CLKBUFX1 gbuf_d_965(.A(_AES_ENC_N143), .Y(ddout__965));
CLKBUFX1 gbuf_q_965(.A(qq_in965), .Y(_AES_ENC_sa02[1]));
CLKBUFX1 gbuf_d_966(.A(_AES_ENC_N142), .Y(ddout__966));
CLKBUFX1 gbuf_q_966(.A(qq_in966), .Y(_AES_ENC_sa02[0]));
CLKBUFX1 gbuf_d_967(.A(_AES_ENC_N62), .Y(ddout__967));
CLKBUFX1 gbuf_q_967(.A(qq_in967), .Y(_AES_ENC_sa13[0]));
CLKBUFX1 gbuf_d_968(.A(_AES_ENC_N63), .Y(ddout__968));
CLKBUFX1 gbuf_q_968(.A(qq_in968), .Y(_AES_ENC_sa13[1]));
CLKBUFX1 gbuf_d_969(.A(_AES_ENC_N65), .Y(ddout__969));
CLKBUFX1 gbuf_q_969(.A(qq_in969), .Y(_AES_ENC_sa13[3]));
CLKBUFX1 gbuf_d_970(.A(_AES_ENC_N66), .Y(ddout__970));
CLKBUFX1 gbuf_q_970(.A(qq_in970), .Y(_AES_ENC_sa13[4]));
CLKBUFX1 gbuf_d_971(.A(_AES_ENC_N37), .Y(ddout__971));
CLKBUFX1 gbuf_q_971(.A(qq_in971), .Y(_AES_ENC_sa33[7]));
CLKBUFX1 gbuf_d_972(.A(_AES_ENC_N165), .Y(ddout__972));
CLKBUFX1 gbuf_q_972(.A(qq_in972), .Y(_AES_ENC_sa31[7]));
CLKBUFX1 gbuf_d_973(.A(_AES_ENC_N46), .Y(ddout__973));
CLKBUFX1 gbuf_q_973(.A(qq_in973), .Y(_AES_ENC_sa23[0]));
CLKBUFX1 gbuf_d_974(.A(_AES_ENC_N47), .Y(ddout__974));
CLKBUFX1 gbuf_q_974(.A(qq_in974), .Y(_AES_ENC_sa23[1]));
CLKBUFX1 gbuf_d_975(.A(_AES_ENC_N49), .Y(ddout__975));
CLKBUFX1 gbuf_q_975(.A(qq_in975), .Y(_AES_ENC_sa23[3]));
CLKBUFX1 gbuf_d_976(.A(_AES_ENC_N50), .Y(ddout__976));
CLKBUFX1 gbuf_q_976(.A(qq_in976), .Y(_AES_ENC_sa23[4]));
CLKBUFX1 gbuf_d_977(.A(_AES_ENC_N69), .Y(ddout__977));
CLKBUFX1 gbuf_q_977(.A(qq_in977), .Y(_AES_ENC_sa13[7]));
CLKBUFX1 gbuf_d_978(.A(_AES_ENC_N68), .Y(ddout__978));
CLKBUFX1 gbuf_q_978(.A(qq_in978), .Y(_AES_ENC_sa13[6]));
CLKBUFX1 gbuf_d_979(.A(_AES_ENC_N36), .Y(ddout__979));
CLKBUFX1 gbuf_q_979(.A(qq_in979), .Y(_AES_ENC_sa33[6]));
CLKBUFX1 gbuf_d_980(.A(_AES_ENC_N52), .Y(ddout__980));
CLKBUFX1 gbuf_q_980(.A(qq_in980), .Y(_AES_ENC_sa23[6]));
CLKBUFX1 gbuf_d_981(.A(_AES_ENC_N67), .Y(ddout__981));
CLKBUFX1 gbuf_q_981(.A(qq_in981), .Y(_AES_ENC_sa13[5]));
CLKBUFX1 gbuf_d_982(.A(_AES_ENC_N35), .Y(ddout__982));
CLKBUFX1 gbuf_q_982(.A(qq_in982), .Y(_AES_ENC_sa33[5]));
CLKBUFX1 gbuf_d_983(.A(_AES_ENC_N51), .Y(ddout__983));
CLKBUFX1 gbuf_q_983(.A(qq_in983), .Y(_AES_ENC_sa23[5]));
CLKBUFX1 gbuf_d_984(.A(_AES_ENC_N84), .Y(ddout__984));
CLKBUFX1 gbuf_q_984(.A(qq_in984), .Y(_AES_ENC_sa03[6]));
CLKBUFX1 gbuf_d_985(.A(_AES_ENC_N34), .Y(ddout__985));
CLKBUFX1 gbuf_q_985(.A(qq_in985), .Y(_AES_ENC_sa33[4]));
CLKBUFX1 gbuf_d_986(.A(_AES_ENC_N83), .Y(ddout__986));
CLKBUFX1 gbuf_q_986(.A(qq_in986), .Y(_AES_ENC_sa03[5]));
CLKBUFX1 gbuf_d_987(.A(_AES_ENC_N33), .Y(ddout__987));
CLKBUFX1 gbuf_q_987(.A(qq_in987), .Y(_AES_ENC_sa33[3]));
CLKBUFX1 gbuf_d_988(.A(_AES_ENC_N82), .Y(ddout__988));
CLKBUFX1 gbuf_q_988(.A(qq_in988), .Y(_AES_ENC_sa03[4]));
CLKBUFX1 gbuf_d_989(.A(_AES_ENC_N64), .Y(ddout__989));
CLKBUFX1 gbuf_q_989(.A(qq_in989), .Y(_AES_ENC_sa13[2]));
CLKBUFX1 gbuf_d_990(.A(_AES_ENC_N32), .Y(ddout__990));
CLKBUFX1 gbuf_q_990(.A(qq_in990), .Y(_AES_ENC_sa33[2]));
CLKBUFX1 gbuf_d_991(.A(_AES_ENC_N48), .Y(ddout__991));
CLKBUFX1 gbuf_q_991(.A(qq_in991), .Y(_AES_ENC_sa23[2]));
CLKBUFX1 gbuf_d_992(.A(_AES_ENC_N81), .Y(ddout__992));
CLKBUFX1 gbuf_q_992(.A(qq_in992), .Y(_AES_ENC_sa03[3]));
CLKBUFX1 gbuf_d_993(.A(_AES_ENC_N31), .Y(ddout__993));
CLKBUFX1 gbuf_q_993(.A(qq_in993), .Y(_AES_ENC_sa33[1]));
CLKBUFX1 gbuf_d_994(.A(_AES_ENC_N80), .Y(ddout__994));
CLKBUFX1 gbuf_q_994(.A(qq_in994), .Y(_AES_ENC_sa03[2]));
CLKBUFX1 gbuf_d_995(.A(_AES_ENC_N79), .Y(ddout__995));
CLKBUFX1 gbuf_q_995(.A(qq_in995), .Y(_AES_ENC_sa03[1]));
CLKBUFX1 gbuf_d_996(.A(_AES_ENC_N85), .Y(ddout__996));
CLKBUFX1 gbuf_q_996(.A(qq_in996), .Y(_AES_ENC_sa03[7]));
CLKBUFX1 gbuf_d_997(.A(_AES_ENC_N78), .Y(ddout__997));
CLKBUFX1 gbuf_q_997(.A(qq_in997), .Y(_AES_ENC_sa03[0]));
CLKBUFX1 gbuf_d_998(.A(_AES_ENC_N174), .Y(ddout__998));
CLKBUFX1 gbuf_q_998(.A(qq_in998), .Y(_AES_ENC_sa21[0]));
CLKBUFX1 gbuf_d_999(.A(_AES_ENC_N175), .Y(ddout__999));
CLKBUFX1 gbuf_q_999(.A(qq_in999), .Y(_AES_ENC_sa21[1]));
CLKBUFX1 gbuf_d_1000(.A(_AES_ENC_N177), .Y(ddout__1000));
CLKBUFX1 gbuf_q_1000(.A(qq_in1000), .Y(_AES_ENC_sa21[3]));
CLKBUFX1 gbuf_d_1001(.A(_AES_ENC_N178), .Y(ddout__1001));
CLKBUFX1 gbuf_q_1001(.A(qq_in1001), .Y(_AES_ENC_sa21[4]));
CLKBUFX1 gbuf_d_1002(.A(_AES_ENC_N197), .Y(ddout__1002));
CLKBUFX1 gbuf_q_1002(.A(qq_in1002), .Y(_AES_ENC_sa11[7]));
CLKBUFX1 gbuf_d_1003(.A(_AES_ENC_N181), .Y(ddout__1003));
CLKBUFX1 gbuf_q_1003(.A(qq_in1003), .Y(_AES_ENC_sa21[7]));
CLKBUFX1 gbuf_d_1004(.A(_AES_ENC_N206), .Y(ddout__1004));
CLKBUFX1 gbuf_q_1004(.A(qq_in1004), .Y(_AES_ENC_sa01[0]));
CLKBUFX1 gbuf_d_1005(.A(_AES_ENC_N207), .Y(ddout__1005));
CLKBUFX1 gbuf_q_1005(.A(qq_in1005), .Y(_AES_ENC_sa01[1]));
CLKBUFX1 gbuf_d_1006(.A(_AES_ENC_N209), .Y(ddout__1006));
CLKBUFX1 gbuf_q_1006(.A(qq_in1006), .Y(_AES_ENC_sa01[3]));
CLKBUFX1 gbuf_d_1007(.A(_AES_ENC_N210), .Y(ddout__1007));
CLKBUFX1 gbuf_q_1007(.A(qq_in1007), .Y(_AES_ENC_sa01[4]));
CLKBUFX1 gbuf_d_1008(.A(_AES_ENC_N196), .Y(ddout__1008));
CLKBUFX1 gbuf_q_1008(.A(qq_in1008), .Y(_AES_ENC_sa11[6]));
CLKBUFX1 gbuf_d_1009(.A(_AES_ENC_N164), .Y(ddout__1009));
CLKBUFX1 gbuf_q_1009(.A(qq_in1009), .Y(_AES_ENC_sa31[6]));
CLKBUFX1 gbuf_d_1010(.A(_AES_ENC_N180), .Y(ddout__1010));
CLKBUFX1 gbuf_q_1010(.A(qq_in1010), .Y(_AES_ENC_sa21[6]));
CLKBUFX1 gbuf_d_1011(.A(_AES_ENC_N195), .Y(ddout__1011));
CLKBUFX1 gbuf_q_1011(.A(qq_in1011), .Y(_AES_ENC_sa11[5]));
CLKBUFX1 gbuf_d_1012(.A(_AES_ENC_N163), .Y(ddout__1012));
CLKBUFX1 gbuf_q_1012(.A(qq_in1012), .Y(_AES_ENC_sa31[5]));
CLKBUFX1 gbuf_d_1013(.A(_AES_ENC_N179), .Y(ddout__1013));
CLKBUFX1 gbuf_q_1013(.A(qq_in1013), .Y(_AES_ENC_sa21[5]));
CLKBUFX1 gbuf_d_1014(.A(_AES_ENC_N212), .Y(ddout__1014));
CLKBUFX1 gbuf_q_1014(.A(qq_in1014), .Y(_AES_ENC_sa01[6]));
CLKBUFX1 gbuf_d_1015(.A(_AES_ENC_N194), .Y(ddout__1015));
CLKBUFX1 gbuf_q_1015(.A(qq_in1015), .Y(_AES_ENC_sa11[4]));
CLKBUFX1 gbuf_d_1016(.A(_AES_ENC_N162), .Y(ddout__1016));
CLKBUFX1 gbuf_q_1016(.A(qq_in1016), .Y(_AES_ENC_sa31[4]));
CLKBUFX1 gbuf_d_1017(.A(_AES_ENC_N211), .Y(ddout__1017));
CLKBUFX1 gbuf_q_1017(.A(qq_in1017), .Y(_AES_ENC_sa01[5]));
CLKBUFX1 gbuf_d_1018(.A(_AES_ENC_N193), .Y(ddout__1018));
CLKBUFX1 gbuf_q_1018(.A(qq_in1018), .Y(_AES_ENC_sa11[3]));
CLKBUFX1 gbuf_d_1019(.A(_AES_ENC_N161), .Y(ddout__1019));
CLKBUFX1 gbuf_q_1019(.A(qq_in1019), .Y(_AES_ENC_sa31[3]));
CLKBUFX1 gbuf_d_1020(.A(_AES_ENC_N192), .Y(ddout__1020));
CLKBUFX1 gbuf_q_1020(.A(qq_in1020), .Y(_AES_ENC_sa11[2]));
CLKBUFX1 gbuf_d_1021(.A(_AES_ENC_N160), .Y(ddout__1021));
CLKBUFX1 gbuf_q_1021(.A(qq_in1021), .Y(_AES_ENC_sa31[2]));
CLKBUFX1 gbuf_d_1022(.A(_AES_ENC_N176), .Y(ddout__1022));
CLKBUFX1 gbuf_q_1022(.A(qq_in1022), .Y(_AES_ENC_sa21[2]));
CLKBUFX1 gbuf_d_1023(.A(_AES_ENC_N191), .Y(ddout__1023));
CLKBUFX1 gbuf_q_1023(.A(qq_in1023), .Y(_AES_ENC_sa11[1]));
CLKBUFX1 gbuf_d_1024(.A(_AES_ENC_N159), .Y(ddout__1024));
CLKBUFX1 gbuf_q_1024(.A(qq_in1024), .Y(_AES_ENC_sa31[1]));
CLKBUFX1 gbuf_d_1025(.A(_AES_ENC_N208), .Y(ddout__1025));
CLKBUFX1 gbuf_q_1025(.A(qq_in1025), .Y(_AES_ENC_sa01[2]));
CLKBUFX1 gbuf_d_1026(.A(_AES_ENC_N213), .Y(ddout__1026));
CLKBUFX1 gbuf_q_1026(.A(qq_in1026), .Y(_AES_ENC_sa01[7]));
CLKBUFX1 gbuf_d_1027(.A(_AES_ENC_N53), .Y(ddout__1027));
CLKBUFX1 gbuf_q_1027(.A(qq_in1027), .Y(_AES_ENC_sa23[7]));
CLKBUFX1 gbuf_d_1028(.A(_AES_ENC_N254), .Y(ddout__1028));
CLKBUFX1 gbuf_q_1028(.A(qq_in1028), .Y(_AES_ENC_sa10[0]));
CLKBUFX1 gbuf_d_1029(.A(_AES_ENC_N190), .Y(ddout__1029));
CLKBUFX1 gbuf_q_1029(.A(qq_in1029), .Y(_AES_ENC_sa11[0]));
CLKBUFX1 gbuf_d_1030(.A(_AES_ENC_N126), .Y(ddout__1030));
CLKBUFX1 gbuf_q_1030(.A(qq_in1030), .Y(_AES_ENC_sa12[0]));
CLKBUFX1 gbuf_d_1031(.A(_AES_ENC_N245), .Y(ddout__1031));
CLKBUFX1 gbuf_q_1031(.A(qq_in1031), .Y(_AES_ENC_sa20[7]));
CLKBUFX1 gbuf_d_1032(.A(_AES_ENC_N30), .Y(ddout__1032));
CLKBUFX1 gbuf_q_1032(.A(qq_in1032), .Y(_AES_ENC_sa33[0]));
CLKBUFX1 gbuf_d_1033(.A(_AES_ENC_N94), .Y(ddout__1033));
CLKBUFX1 gbuf_q_1033(.A(qq_in1033), .Y(_AES_ENC_sa32[0]));
CLKBUFX1 gbuf_d_1034(.A(_AES_ENC_N158), .Y(ddout__1034));
CLKBUFX1 gbuf_q_1034(.A(qq_in1034), .Y(_AES_ENC_sa31[0]));
CLKBUFX1 gbuf_d_1035(.A(_AES_ENC_N222), .Y(ddout__1035));
CLKBUFX1 gbuf_q_1035(.A(qq_in1035), .Y(_AES_ENC_sa30[0]));
CLKBUFX1 gbuf_d_1036(.A(_AES_ENC_N270), .Y(ddout__1036));
CLKBUFX1 gbuf_q_1036(.A(qq_in1036), .Y(_AES_ENC_sa00[0]));
CLKBUFX1 gbuf_d_1037(.A(_AES_ENC_n661), .Y(ddout__1037));
CLKBUFX1 gbuf_q_1037(.A(qq_in1037), .Y(_AES_ENC_text_in_r[0]));
CLKBUFX1 gbuf_d_1038(.A(_AES_ENC_n662), .Y(ddout__1038));
CLKBUFX1 gbuf_q_1038(.A(qq_in1038), .Y(_AES_ENC_text_in_r[1]));
CLKBUFX1 gbuf_d_1039(.A(_AES_ENC_n663), .Y(ddout__1039));
CLKBUFX1 gbuf_q_1039(.A(qq_in1039), .Y(_AES_ENC_text_in_r[2]));
CLKBUFX1 gbuf_d_1040(.A(_AES_ENC_n664), .Y(ddout__1040));
CLKBUFX1 gbuf_q_1040(.A(qq_in1040), .Y(_AES_ENC_text_in_r[3]));
CLKBUFX1 gbuf_d_1041(.A(_AES_ENC_n665), .Y(ddout__1041));
CLKBUFX1 gbuf_q_1041(.A(qq_in1041), .Y(_AES_ENC_text_in_r[4]));
CLKBUFX1 gbuf_d_1042(.A(_AES_ENC_n666), .Y(ddout__1042));
CLKBUFX1 gbuf_q_1042(.A(qq_in1042), .Y(_AES_ENC_text_in_r[5]));
CLKBUFX1 gbuf_d_1043(.A(_AES_ENC_n667), .Y(ddout__1043));
CLKBUFX1 gbuf_q_1043(.A(qq_in1043), .Y(_AES_ENC_text_in_r[6]));
CLKBUFX1 gbuf_d_1044(.A(_AES_ENC_n668), .Y(ddout__1044));
CLKBUFX1 gbuf_q_1044(.A(qq_in1044), .Y(_AES_ENC_text_in_r[7]));
CLKBUFX1 gbuf_d_1045(.A(_AES_ENC_n669), .Y(ddout__1045));
CLKBUFX1 gbuf_q_1045(.A(qq_in1045), .Y(_AES_ENC_text_in_r[8]));
CLKBUFX1 gbuf_d_1046(.A(_AES_ENC_n670), .Y(ddout__1046));
CLKBUFX1 gbuf_q_1046(.A(qq_in1046), .Y(_AES_ENC_text_in_r[9]));
CLKBUFX1 gbuf_d_1047(.A(_AES_ENC_n671), .Y(ddout__1047));
CLKBUFX1 gbuf_q_1047(.A(qq_in1047), .Y(_AES_ENC_text_in_r[10]));
CLKBUFX1 gbuf_d_1048(.A(_AES_ENC_n672), .Y(ddout__1048));
CLKBUFX1 gbuf_q_1048(.A(qq_in1048), .Y(_AES_ENC_text_in_r[11]));
CLKBUFX1 gbuf_d_1049(.A(_AES_ENC_n673), .Y(ddout__1049));
CLKBUFX1 gbuf_q_1049(.A(qq_in1049), .Y(_AES_ENC_text_in_r[12]));
CLKBUFX1 gbuf_d_1050(.A(_AES_ENC_n674), .Y(ddout__1050));
CLKBUFX1 gbuf_q_1050(.A(qq_in1050), .Y(_AES_ENC_text_in_r[13]));
CLKBUFX1 gbuf_d_1051(.A(_AES_ENC_n675), .Y(ddout__1051));
CLKBUFX1 gbuf_q_1051(.A(qq_in1051), .Y(_AES_ENC_text_in_r[14]));
CLKBUFX1 gbuf_d_1052(.A(_AES_ENC_n676), .Y(ddout__1052));
CLKBUFX1 gbuf_q_1052(.A(qq_in1052), .Y(_AES_ENC_text_in_r[15]));
CLKBUFX1 gbuf_d_1053(.A(_AES_ENC_n677), .Y(ddout__1053));
CLKBUFX1 gbuf_q_1053(.A(qq_in1053), .Y(_AES_ENC_text_in_r[16]));
CLKBUFX1 gbuf_d_1054(.A(_AES_ENC_n678), .Y(ddout__1054));
CLKBUFX1 gbuf_q_1054(.A(qq_in1054), .Y(_AES_ENC_text_in_r[17]));
CLKBUFX1 gbuf_d_1055(.A(_AES_ENC_n679), .Y(ddout__1055));
CLKBUFX1 gbuf_q_1055(.A(qq_in1055), .Y(_AES_ENC_text_in_r[18]));
CLKBUFX1 gbuf_d_1056(.A(_AES_ENC_n680), .Y(ddout__1056));
CLKBUFX1 gbuf_q_1056(.A(qq_in1056), .Y(_AES_ENC_text_in_r[19]));
CLKBUFX1 gbuf_d_1057(.A(_AES_ENC_n681), .Y(ddout__1057));
CLKBUFX1 gbuf_q_1057(.A(qq_in1057), .Y(_AES_ENC_text_in_r[20]));
CLKBUFX1 gbuf_d_1058(.A(_AES_ENC_n682), .Y(ddout__1058));
CLKBUFX1 gbuf_q_1058(.A(qq_in1058), .Y(_AES_ENC_text_in_r[21]));
CLKBUFX1 gbuf_d_1059(.A(_AES_ENC_n683), .Y(ddout__1059));
CLKBUFX1 gbuf_q_1059(.A(qq_in1059), .Y(_AES_ENC_text_in_r[22]));
CLKBUFX1 gbuf_d_1060(.A(_AES_ENC_n684), .Y(ddout__1060));
CLKBUFX1 gbuf_q_1060(.A(qq_in1060), .Y(_AES_ENC_text_in_r[23]));
CLKBUFX1 gbuf_d_1061(.A(_AES_ENC_n685), .Y(ddout__1061));
CLKBUFX1 gbuf_q_1061(.A(qq_in1061), .Y(_AES_ENC_text_in_r[24]));
CLKBUFX1 gbuf_d_1062(.A(_AES_ENC_n686), .Y(ddout__1062));
CLKBUFX1 gbuf_q_1062(.A(qq_in1062), .Y(_AES_ENC_text_in_r[25]));
CLKBUFX1 gbuf_d_1063(.A(_AES_ENC_n687), .Y(ddout__1063));
CLKBUFX1 gbuf_q_1063(.A(qq_in1063), .Y(_AES_ENC_text_in_r[26]));
CLKBUFX1 gbuf_d_1064(.A(_AES_ENC_n688), .Y(ddout__1064));
CLKBUFX1 gbuf_q_1064(.A(qq_in1064), .Y(_AES_ENC_text_in_r[27]));
CLKBUFX1 gbuf_d_1065(.A(_AES_ENC_n689), .Y(ddout__1065));
CLKBUFX1 gbuf_q_1065(.A(qq_in1065), .Y(_AES_ENC_text_in_r[28]));
CLKBUFX1 gbuf_d_1066(.A(_AES_ENC_n690), .Y(ddout__1066));
CLKBUFX1 gbuf_q_1066(.A(qq_in1066), .Y(_AES_ENC_text_in_r[29]));
CLKBUFX1 gbuf_d_1067(.A(_AES_ENC_n691), .Y(ddout__1067));
CLKBUFX1 gbuf_q_1067(.A(qq_in1067), .Y(_AES_ENC_text_in_r[30]));
CLKBUFX1 gbuf_d_1068(.A(_AES_ENC_n692), .Y(ddout__1068));
CLKBUFX1 gbuf_q_1068(.A(qq_in1068), .Y(_AES_ENC_text_in_r[31]));
CLKBUFX1 gbuf_d_1069(.A(_AES_ENC_n693), .Y(ddout__1069));
CLKBUFX1 gbuf_q_1069(.A(qq_in1069), .Y(_AES_ENC_text_in_r[32]));
CLKBUFX1 gbuf_d_1070(.A(_AES_ENC_n694), .Y(ddout__1070));
CLKBUFX1 gbuf_q_1070(.A(qq_in1070), .Y(_AES_ENC_text_in_r[33]));
CLKBUFX1 gbuf_d_1071(.A(_AES_ENC_n695), .Y(ddout__1071));
CLKBUFX1 gbuf_q_1071(.A(qq_in1071), .Y(_AES_ENC_text_in_r[34]));
CLKBUFX1 gbuf_d_1072(.A(_AES_ENC_n696), .Y(ddout__1072));
CLKBUFX1 gbuf_q_1072(.A(qq_in1072), .Y(_AES_ENC_text_in_r[35]));
CLKBUFX1 gbuf_d_1073(.A(_AES_ENC_n697), .Y(ddout__1073));
CLKBUFX1 gbuf_q_1073(.A(qq_in1073), .Y(_AES_ENC_text_in_r[36]));
CLKBUFX1 gbuf_d_1074(.A(_AES_ENC_n698), .Y(ddout__1074));
CLKBUFX1 gbuf_q_1074(.A(qq_in1074), .Y(_AES_ENC_text_in_r[37]));
CLKBUFX1 gbuf_d_1075(.A(_AES_ENC_n699), .Y(ddout__1075));
CLKBUFX1 gbuf_q_1075(.A(qq_in1075), .Y(_AES_ENC_text_in_r[38]));
CLKBUFX1 gbuf_d_1076(.A(_AES_ENC_n700), .Y(ddout__1076));
CLKBUFX1 gbuf_q_1076(.A(qq_in1076), .Y(_AES_ENC_text_in_r[39]));
CLKBUFX1 gbuf_d_1077(.A(_AES_ENC_n701), .Y(ddout__1077));
CLKBUFX1 gbuf_q_1077(.A(qq_in1077), .Y(_AES_ENC_text_in_r[40]));
CLKBUFX1 gbuf_d_1078(.A(_AES_ENC_n702), .Y(ddout__1078));
CLKBUFX1 gbuf_q_1078(.A(qq_in1078), .Y(_AES_ENC_text_in_r[41]));
CLKBUFX1 gbuf_d_1079(.A(_AES_ENC_n703), .Y(ddout__1079));
CLKBUFX1 gbuf_q_1079(.A(qq_in1079), .Y(_AES_ENC_text_in_r[42]));
CLKBUFX1 gbuf_d_1080(.A(_AES_ENC_n704), .Y(ddout__1080));
CLKBUFX1 gbuf_q_1080(.A(qq_in1080), .Y(_AES_ENC_text_in_r[43]));
CLKBUFX1 gbuf_d_1081(.A(_AES_ENC_n705), .Y(ddout__1081));
CLKBUFX1 gbuf_q_1081(.A(qq_in1081), .Y(_AES_ENC_text_in_r[44]));
CLKBUFX1 gbuf_d_1082(.A(_AES_ENC_n706), .Y(ddout__1082));
CLKBUFX1 gbuf_q_1082(.A(qq_in1082), .Y(_AES_ENC_text_in_r[45]));
CLKBUFX1 gbuf_d_1083(.A(_AES_ENC_n707), .Y(ddout__1083));
CLKBUFX1 gbuf_q_1083(.A(qq_in1083), .Y(_AES_ENC_text_in_r[46]));
CLKBUFX1 gbuf_d_1084(.A(_AES_ENC_n708), .Y(ddout__1084));
CLKBUFX1 gbuf_q_1084(.A(qq_in1084), .Y(_AES_ENC_text_in_r[47]));
CLKBUFX1 gbuf_d_1085(.A(_AES_ENC_n709), .Y(ddout__1085));
CLKBUFX1 gbuf_q_1085(.A(qq_in1085), .Y(_AES_ENC_text_in_r[48]));
CLKBUFX1 gbuf_d_1086(.A(_AES_ENC_n710), .Y(ddout__1086));
CLKBUFX1 gbuf_q_1086(.A(qq_in1086), .Y(_AES_ENC_text_in_r[49]));
CLKBUFX1 gbuf_d_1087(.A(_AES_ENC_n711), .Y(ddout__1087));
CLKBUFX1 gbuf_q_1087(.A(qq_in1087), .Y(_AES_ENC_text_in_r[50]));
CLKBUFX1 gbuf_d_1088(.A(_AES_ENC_n712), .Y(ddout__1088));
CLKBUFX1 gbuf_q_1088(.A(qq_in1088), .Y(_AES_ENC_text_in_r[51]));
CLKBUFX1 gbuf_d_1089(.A(_AES_ENC_n713), .Y(ddout__1089));
CLKBUFX1 gbuf_q_1089(.A(qq_in1089), .Y(_AES_ENC_text_in_r[52]));
CLKBUFX1 gbuf_d_1090(.A(_AES_ENC_n714), .Y(ddout__1090));
CLKBUFX1 gbuf_q_1090(.A(qq_in1090), .Y(_AES_ENC_text_in_r[53]));
CLKBUFX1 gbuf_d_1091(.A(_AES_ENC_n715), .Y(ddout__1091));
CLKBUFX1 gbuf_q_1091(.A(qq_in1091), .Y(_AES_ENC_text_in_r[54]));
CLKBUFX1 gbuf_d_1092(.A(_AES_ENC_n716), .Y(ddout__1092));
CLKBUFX1 gbuf_q_1092(.A(qq_in1092), .Y(_AES_ENC_text_in_r[55]));
CLKBUFX1 gbuf_d_1093(.A(_AES_ENC_n717), .Y(ddout__1093));
CLKBUFX1 gbuf_q_1093(.A(qq_in1093), .Y(_AES_ENC_text_in_r[56]));
CLKBUFX1 gbuf_d_1094(.A(_AES_ENC_n718), .Y(ddout__1094));
CLKBUFX1 gbuf_q_1094(.A(qq_in1094), .Y(_AES_ENC_text_in_r[57]));
CLKBUFX1 gbuf_d_1095(.A(_AES_ENC_n719), .Y(ddout__1095));
CLKBUFX1 gbuf_q_1095(.A(qq_in1095), .Y(_AES_ENC_text_in_r[58]));
CLKBUFX1 gbuf_d_1096(.A(_AES_ENC_n720), .Y(ddout__1096));
CLKBUFX1 gbuf_q_1096(.A(qq_in1096), .Y(_AES_ENC_text_in_r[59]));
CLKBUFX1 gbuf_d_1097(.A(_AES_ENC_n721), .Y(ddout__1097));
CLKBUFX1 gbuf_q_1097(.A(qq_in1097), .Y(_AES_ENC_text_in_r[60]));
CLKBUFX1 gbuf_d_1098(.A(_AES_ENC_n722), .Y(ddout__1098));
CLKBUFX1 gbuf_q_1098(.A(qq_in1098), .Y(_AES_ENC_text_in_r[61]));
CLKBUFX1 gbuf_d_1099(.A(_AES_ENC_n723), .Y(ddout__1099));
CLKBUFX1 gbuf_q_1099(.A(qq_in1099), .Y(_AES_ENC_text_in_r[62]));
CLKBUFX1 gbuf_d_1100(.A(_AES_ENC_n724), .Y(ddout__1100));
CLKBUFX1 gbuf_q_1100(.A(qq_in1100), .Y(_AES_ENC_text_in_r[63]));
CLKBUFX1 gbuf_d_1101(.A(_AES_ENC_n725), .Y(ddout__1101));
CLKBUFX1 gbuf_q_1101(.A(qq_in1101), .Y(_AES_ENC_text_in_r[64]));
CLKBUFX1 gbuf_d_1102(.A(_AES_ENC_n726), .Y(ddout__1102));
CLKBUFX1 gbuf_q_1102(.A(qq_in1102), .Y(_AES_ENC_text_in_r[65]));
CLKBUFX1 gbuf_d_1103(.A(_AES_ENC_n727), .Y(ddout__1103));
CLKBUFX1 gbuf_q_1103(.A(qq_in1103), .Y(_AES_ENC_text_in_r[66]));
CLKBUFX1 gbuf_d_1104(.A(_AES_ENC_n728), .Y(ddout__1104));
CLKBUFX1 gbuf_q_1104(.A(qq_in1104), .Y(_AES_ENC_text_in_r[67]));
CLKBUFX1 gbuf_d_1105(.A(_AES_ENC_n729), .Y(ddout__1105));
CLKBUFX1 gbuf_q_1105(.A(qq_in1105), .Y(_AES_ENC_text_in_r[68]));
CLKBUFX1 gbuf_d_1106(.A(_AES_ENC_n730), .Y(ddout__1106));
CLKBUFX1 gbuf_q_1106(.A(qq_in1106), .Y(_AES_ENC_text_in_r[69]));
CLKBUFX1 gbuf_d_1107(.A(_AES_ENC_n731), .Y(ddout__1107));
CLKBUFX1 gbuf_q_1107(.A(qq_in1107), .Y(_AES_ENC_text_in_r[70]));
CLKBUFX1 gbuf_d_1108(.A(_AES_ENC_n732), .Y(ddout__1108));
CLKBUFX1 gbuf_q_1108(.A(qq_in1108), .Y(_AES_ENC_text_in_r[71]));
CLKBUFX1 gbuf_d_1109(.A(_AES_ENC_n733), .Y(ddout__1109));
CLKBUFX1 gbuf_q_1109(.A(qq_in1109), .Y(_AES_ENC_text_in_r[72]));
CLKBUFX1 gbuf_d_1110(.A(_AES_ENC_n734), .Y(ddout__1110));
CLKBUFX1 gbuf_q_1110(.A(qq_in1110), .Y(_AES_ENC_text_in_r[73]));
CLKBUFX1 gbuf_d_1111(.A(_AES_ENC_n735), .Y(ddout__1111));
CLKBUFX1 gbuf_q_1111(.A(qq_in1111), .Y(_AES_ENC_text_in_r[74]));
CLKBUFX1 gbuf_d_1112(.A(_AES_ENC_n736), .Y(ddout__1112));
CLKBUFX1 gbuf_q_1112(.A(qq_in1112), .Y(_AES_ENC_text_in_r[75]));
CLKBUFX1 gbuf_d_1113(.A(_AES_ENC_n737), .Y(ddout__1113));
CLKBUFX1 gbuf_q_1113(.A(qq_in1113), .Y(_AES_ENC_text_in_r[76]));
CLKBUFX1 gbuf_d_1114(.A(_AES_ENC_n738), .Y(ddout__1114));
CLKBUFX1 gbuf_q_1114(.A(qq_in1114), .Y(_AES_ENC_text_in_r[77]));
CLKBUFX1 gbuf_d_1115(.A(_AES_ENC_n739), .Y(ddout__1115));
CLKBUFX1 gbuf_q_1115(.A(qq_in1115), .Y(_AES_ENC_text_in_r[78]));
CLKBUFX1 gbuf_d_1116(.A(_AES_ENC_n740), .Y(ddout__1116));
CLKBUFX1 gbuf_q_1116(.A(qq_in1116), .Y(_AES_ENC_text_in_r[79]));
CLKBUFX1 gbuf_d_1117(.A(_AES_ENC_n741), .Y(ddout__1117));
CLKBUFX1 gbuf_q_1117(.A(qq_in1117), .Y(_AES_ENC_text_in_r[80]));
CLKBUFX1 gbuf_d_1118(.A(_AES_ENC_n742), .Y(ddout__1118));
CLKBUFX1 gbuf_q_1118(.A(qq_in1118), .Y(_AES_ENC_text_in_r[81]));
CLKBUFX1 gbuf_d_1119(.A(_AES_ENC_n743), .Y(ddout__1119));
CLKBUFX1 gbuf_q_1119(.A(qq_in1119), .Y(_AES_ENC_text_in_r[82]));
CLKBUFX1 gbuf_d_1120(.A(_AES_ENC_n744), .Y(ddout__1120));
CLKBUFX1 gbuf_q_1120(.A(qq_in1120), .Y(_AES_ENC_text_in_r[83]));
CLKBUFX1 gbuf_d_1121(.A(_AES_ENC_n745), .Y(ddout__1121));
CLKBUFX1 gbuf_q_1121(.A(qq_in1121), .Y(_AES_ENC_text_in_r[84]));
CLKBUFX1 gbuf_d_1122(.A(_AES_ENC_n746), .Y(ddout__1122));
CLKBUFX1 gbuf_q_1122(.A(qq_in1122), .Y(_AES_ENC_text_in_r[85]));
CLKBUFX1 gbuf_d_1123(.A(_AES_ENC_n747), .Y(ddout__1123));
CLKBUFX1 gbuf_q_1123(.A(qq_in1123), .Y(_AES_ENC_text_in_r[86]));
CLKBUFX1 gbuf_d_1124(.A(_AES_ENC_n748), .Y(ddout__1124));
CLKBUFX1 gbuf_q_1124(.A(qq_in1124), .Y(_AES_ENC_text_in_r[87]));
CLKBUFX1 gbuf_d_1125(.A(_AES_ENC_n749), .Y(ddout__1125));
CLKBUFX1 gbuf_q_1125(.A(qq_in1125), .Y(_AES_ENC_text_in_r[88]));
CLKBUFX1 gbuf_d_1126(.A(_AES_ENC_n750), .Y(ddout__1126));
CLKBUFX1 gbuf_q_1126(.A(qq_in1126), .Y(_AES_ENC_text_in_r[89]));
CLKBUFX1 gbuf_d_1127(.A(_AES_ENC_n751), .Y(ddout__1127));
CLKBUFX1 gbuf_q_1127(.A(qq_in1127), .Y(_AES_ENC_text_in_r[90]));
CLKBUFX1 gbuf_d_1128(.A(_AES_ENC_n752), .Y(ddout__1128));
CLKBUFX1 gbuf_q_1128(.A(qq_in1128), .Y(_AES_ENC_text_in_r[91]));
CLKBUFX1 gbuf_d_1129(.A(_AES_ENC_n753), .Y(ddout__1129));
CLKBUFX1 gbuf_q_1129(.A(qq_in1129), .Y(_AES_ENC_text_in_r[92]));
CLKBUFX1 gbuf_d_1130(.A(_AES_ENC_n754), .Y(ddout__1130));
CLKBUFX1 gbuf_q_1130(.A(qq_in1130), .Y(_AES_ENC_text_in_r[93]));
CLKBUFX1 gbuf_d_1131(.A(_AES_ENC_n755), .Y(ddout__1131));
CLKBUFX1 gbuf_q_1131(.A(qq_in1131), .Y(_AES_ENC_text_in_r[94]));
CLKBUFX1 gbuf_d_1132(.A(_AES_ENC_n756), .Y(ddout__1132));
CLKBUFX1 gbuf_q_1132(.A(qq_in1132), .Y(_AES_ENC_text_in_r[95]));
CLKBUFX1 gbuf_d_1133(.A(_AES_ENC_n757), .Y(ddout__1133));
CLKBUFX1 gbuf_q_1133(.A(qq_in1133), .Y(_AES_ENC_text_in_r[96]));
CLKBUFX1 gbuf_d_1134(.A(_AES_ENC_n758), .Y(ddout__1134));
CLKBUFX1 gbuf_q_1134(.A(qq_in1134), .Y(_AES_ENC_text_in_r[97]));
CLKBUFX1 gbuf_d_1135(.A(_AES_ENC_n759), .Y(ddout__1135));
CLKBUFX1 gbuf_q_1135(.A(qq_in1135), .Y(_AES_ENC_text_in_r[98]));
CLKBUFX1 gbuf_d_1136(.A(_AES_ENC_n760), .Y(ddout__1136));
CLKBUFX1 gbuf_q_1136(.A(qq_in1136), .Y(_AES_ENC_text_in_r[99]));
CLKBUFX1 gbuf_d_1137(.A(_AES_ENC_n761), .Y(ddout__1137));
CLKBUFX1 gbuf_q_1137(.A(qq_in1137), .Y(_AES_ENC_text_in_r[100]));
CLKBUFX1 gbuf_d_1138(.A(_AES_ENC_n762), .Y(ddout__1138));
CLKBUFX1 gbuf_q_1138(.A(qq_in1138), .Y(_AES_ENC_text_in_r[101]));
CLKBUFX1 gbuf_d_1139(.A(_AES_ENC_n763), .Y(ddout__1139));
CLKBUFX1 gbuf_q_1139(.A(qq_in1139), .Y(_AES_ENC_text_in_r[102]));
CLKBUFX1 gbuf_d_1140(.A(_AES_ENC_n764), .Y(ddout__1140));
CLKBUFX1 gbuf_q_1140(.A(qq_in1140), .Y(_AES_ENC_text_in_r[103]));
CLKBUFX1 gbuf_d_1141(.A(_AES_ENC_n765), .Y(ddout__1141));
CLKBUFX1 gbuf_q_1141(.A(qq_in1141), .Y(_AES_ENC_text_in_r[104]));
CLKBUFX1 gbuf_d_1142(.A(_AES_ENC_n766), .Y(ddout__1142));
CLKBUFX1 gbuf_q_1142(.A(qq_in1142), .Y(_AES_ENC_text_in_r[105]));
CLKBUFX1 gbuf_d_1143(.A(_AES_ENC_n767), .Y(ddout__1143));
CLKBUFX1 gbuf_q_1143(.A(qq_in1143), .Y(_AES_ENC_text_in_r[106]));
CLKBUFX1 gbuf_d_1144(.A(_AES_ENC_n768), .Y(ddout__1144));
CLKBUFX1 gbuf_q_1144(.A(qq_in1144), .Y(_AES_ENC_text_in_r[107]));
CLKBUFX1 gbuf_d_1145(.A(_AES_ENC_n769), .Y(ddout__1145));
CLKBUFX1 gbuf_q_1145(.A(qq_in1145), .Y(_AES_ENC_text_in_r[108]));
CLKBUFX1 gbuf_d_1146(.A(_AES_ENC_n770), .Y(ddout__1146));
CLKBUFX1 gbuf_q_1146(.A(qq_in1146), .Y(_AES_ENC_text_in_r[109]));
CLKBUFX1 gbuf_d_1147(.A(_AES_ENC_n771), .Y(ddout__1147));
CLKBUFX1 gbuf_q_1147(.A(qq_in1147), .Y(_AES_ENC_text_in_r[110]));
CLKBUFX1 gbuf_d_1148(.A(_AES_ENC_n772), .Y(ddout__1148));
CLKBUFX1 gbuf_q_1148(.A(qq_in1148), .Y(_AES_ENC_text_in_r[111]));
CLKBUFX1 gbuf_d_1149(.A(_AES_ENC_n773), .Y(ddout__1149));
CLKBUFX1 gbuf_q_1149(.A(qq_in1149), .Y(_AES_ENC_text_in_r[112]));
CLKBUFX1 gbuf_d_1150(.A(_AES_ENC_n774), .Y(ddout__1150));
CLKBUFX1 gbuf_q_1150(.A(qq_in1150), .Y(_AES_ENC_text_in_r[113]));
CLKBUFX1 gbuf_d_1151(.A(_AES_ENC_n775), .Y(ddout__1151));
CLKBUFX1 gbuf_q_1151(.A(qq_in1151), .Y(_AES_ENC_text_in_r[114]));
CLKBUFX1 gbuf_d_1152(.A(_AES_ENC_n776), .Y(ddout__1152));
CLKBUFX1 gbuf_q_1152(.A(qq_in1152), .Y(_AES_ENC_text_in_r[115]));
CLKBUFX1 gbuf_d_1153(.A(_AES_ENC_n777), .Y(ddout__1153));
CLKBUFX1 gbuf_q_1153(.A(qq_in1153), .Y(_AES_ENC_text_in_r[116]));
CLKBUFX1 gbuf_d_1154(.A(_AES_ENC_n778), .Y(ddout__1154));
CLKBUFX1 gbuf_q_1154(.A(qq_in1154), .Y(_AES_ENC_text_in_r[117]));
CLKBUFX1 gbuf_d_1155(.A(_AES_ENC_n779), .Y(ddout__1155));
CLKBUFX1 gbuf_q_1155(.A(qq_in1155), .Y(_AES_ENC_text_in_r[118]));
CLKBUFX1 gbuf_d_1156(.A(_AES_ENC_n780), .Y(ddout__1156));
CLKBUFX1 gbuf_q_1156(.A(qq_in1156), .Y(_AES_ENC_text_in_r[119]));
CLKBUFX1 gbuf_d_1157(.A(_AES_ENC_n781), .Y(ddout__1157));
CLKBUFX1 gbuf_q_1157(.A(qq_in1157), .Y(_AES_ENC_text_in_r[120]));
CLKBUFX1 gbuf_d_1158(.A(_AES_ENC_n782), .Y(ddout__1158));
CLKBUFX1 gbuf_q_1158(.A(qq_in1158), .Y(_AES_ENC_text_in_r[121]));
CLKBUFX1 gbuf_d_1159(.A(_AES_ENC_n783), .Y(ddout__1159));
CLKBUFX1 gbuf_q_1159(.A(qq_in1159), .Y(_AES_ENC_text_in_r[122]));
CLKBUFX1 gbuf_d_1160(.A(_AES_ENC_n784), .Y(ddout__1160));
CLKBUFX1 gbuf_q_1160(.A(qq_in1160), .Y(_AES_ENC_text_in_r[123]));
CLKBUFX1 gbuf_d_1161(.A(_AES_ENC_n785), .Y(ddout__1161));
CLKBUFX1 gbuf_q_1161(.A(qq_in1161), .Y(_AES_ENC_text_in_r[124]));
CLKBUFX1 gbuf_d_1162(.A(_AES_ENC_n786), .Y(ddout__1162));
CLKBUFX1 gbuf_q_1162(.A(qq_in1162), .Y(_AES_ENC_text_in_r[125]));
CLKBUFX1 gbuf_d_1163(.A(_AES_ENC_n787), .Y(ddout__1163));
CLKBUFX1 gbuf_q_1163(.A(qq_in1163), .Y(_AES_ENC_text_in_r[126]));
CLKBUFX1 gbuf_d_1164(.A(_AES_ENC_n788), .Y(ddout__1164));
CLKBUFX1 gbuf_q_1164(.A(qq_in1164), .Y(_AES_ENC_text_in_r[127]));
CLKBUFX1 gbuf_d_1165(.A(_AES_ENC_N19), .Y(ddout__1165));
CLKBUFX1 gbuf_q_1165(.A(qq_in1165), .Y(aes_done));
XOR2_X2 _AES_ENC_U1612  ( .A(_AES_ENC_sa22_sub[7] ), .B(_AES_ENC_sa33_sub[7] ), .Z(_AES_ENC_n1167 ) );
XOR2_X2 _AES_ENC_U1611  ( .A(_AES_ENC_sa00_sub[6] ), .B(_AES_ENC_sa11_sub[6] ), .Z(_AES_ENC_n1169 ) );
XOR2_X2 _AES_ENC_U1610  ( .A(_AES_ENC_n800 ), .B(_AES_ENC_n799 ), .Z(_AES_ENC_sa00_next[7]) );
XOR2_X2 _AES_ENC_U1609  ( .A(_AES_ENC_n1167 ), .B(_AES_ENC_n1169 ), .Z(_AES_ENC_n799 ) );
XOR2_X2 _AES_ENC_U1608  ( .A(_AES_ENC_w0[31] ), .B(_AES_ENC_sa11_sub[7] ),.Z(_AES_ENC_n800 ) );
XOR2_X2 _AES_ENC_U1607  ( .A(_AES_ENC_sa00_sub[5] ), .B(_AES_ENC_sa11_sub[5] ), .Z(_AES_ENC_n1170 ) );
XOR2_X2 _AES_ENC_U1606  ( .A(_AES_ENC_sa22_sub[6] ), .B(_AES_ENC_sa33_sub[6] ), .Z(_AES_ENC_n1160 ) );
XOR2_X2 _AES_ENC_U1605  ( .A(_AES_ENC_n802 ), .B(_AES_ENC_n801 ), .Z(_AES_ENC_sa00_next[6]) );
XOR2_X2 _AES_ENC_U1604  ( .A(_AES_ENC_n1170 ), .B(_AES_ENC_n1160 ), .Z(_AES_ENC_n801 ) );
XOR2_X2 _AES_ENC_U1603  ( .A(_AES_ENC_w0[30] ), .B(_AES_ENC_sa11_sub[6] ),.Z(_AES_ENC_n802 ) );
XOR2_X2 _AES_ENC_U1602  ( .A(_AES_ENC_sa00_sub[4] ), .B(_AES_ENC_sa11_sub[4] ), .Z(_AES_ENC_n1171 ) );
XOR2_X2 _AES_ENC_U1601  ( .A(_AES_ENC_sa22_sub[5] ), .B(_AES_ENC_sa33_sub[5] ), .Z(_AES_ENC_n1161 ) );
XOR2_X2 _AES_ENC_U1600  ( .A(_AES_ENC_n804 ), .B(_AES_ENC_n803 ), .Z(_AES_ENC_sa00_next[5]) );
XOR2_X2 _AES_ENC_U1599  ( .A(_AES_ENC_n1171 ), .B(_AES_ENC_n1161 ), .Z(_AES_ENC_n803 ) );
XOR2_X2 _AES_ENC_U1598  ( .A(_AES_ENC_w0[29] ), .B(_AES_ENC_sa11_sub[5] ),.Z(_AES_ENC_n804 ) );
XOR2_X2 _AES_ENC_U1597  ( .A(_AES_ENC_sa00_sub[7] ), .B(_AES_ENC_sa11_sub[7] ), .Z(_AES_ENC_n1168 ) );
XOR2_X2 _AES_ENC_U1596  ( .A(_AES_ENC_sa00_sub[3] ), .B(_AES_ENC_sa11_sub[3] ), .Z(_AES_ENC_n1172 ) );
XOR2_X2 _AES_ENC_U1595  ( .A(_AES_ENC_sa22_sub[4] ), .B(_AES_ENC_sa33_sub[4] ), .Z(_AES_ENC_n1162 ) );
XOR2_X2 _AES_ENC_U1594  ( .A(_AES_ENC_n806 ), .B(_AES_ENC_n805 ), .Z(_AES_ENC_sa00_next[4]) );
XOR2_X2 _AES_ENC_U1593  ( .A(_AES_ENC_n1162 ), .B(_AES_ENC_n807 ), .Z(_AES_ENC_n805 ) );
XOR2_X2 _AES_ENC_U1592  ( .A(_AES_ENC_n1168 ), .B(_AES_ENC_n1172 ), .Z(_AES_ENC_n806 ) );
XOR2_X2 _AES_ENC_U1591  ( .A(_AES_ENC_w0[28] ), .B(_AES_ENC_sa11_sub[4] ),.Z(_AES_ENC_n807 ) );
XOR2_X2 _AES_ENC_U1590  ( .A(_AES_ENC_sa00_sub[2] ), .B(_AES_ENC_sa11_sub[2] ), .Z(_AES_ENC_n1173 ) );
XOR2_X2 _AES_ENC_U1589  ( .A(_AES_ENC_sa22_sub[3] ), .B(_AES_ENC_sa33_sub[3] ), .Z(_AES_ENC_n1163 ) );
XOR2_X2 _AES_ENC_U1588  ( .A(_AES_ENC_n809 ), .B(_AES_ENC_n808 ), .Z(_AES_ENC_sa00_next[3]) );
XOR2_X2 _AES_ENC_U1587  ( .A(_AES_ENC_n1163 ), .B(_AES_ENC_n810 ), .Z(_AES_ENC_n808 ) );
XOR2_X2 _AES_ENC_U1586  ( .A(_AES_ENC_n1168 ), .B(_AES_ENC_n1173 ), .Z(_AES_ENC_n809 ) );
XOR2_X2 _AES_ENC_U1585  ( .A(_AES_ENC_w0[27] ), .B(_AES_ENC_sa11_sub[3] ),.Z(_AES_ENC_n810 ) );
XOR2_X2 _AES_ENC_U1584  ( .A(_AES_ENC_sa00_sub[1] ), .B(_AES_ENC_sa11_sub[1] ), .Z(_AES_ENC_n1174 ) );
XOR2_X2 _AES_ENC_U1583  ( .A(_AES_ENC_sa22_sub[2] ), .B(_AES_ENC_sa33_sub[2] ), .Z(_AES_ENC_n1164 ) );
XOR2_X2 _AES_ENC_U1582  ( .A(_AES_ENC_n812 ), .B(_AES_ENC_n811 ), .Z(_AES_ENC_sa00_next[2]) );
XOR2_X2 _AES_ENC_U1581  ( .A(_AES_ENC_n1174 ), .B(_AES_ENC_n1164 ), .Z(_AES_ENC_n811 ) );
XOR2_X2 _AES_ENC_U1580  ( .A(_AES_ENC_w0[26] ), .B(_AES_ENC_sa11_sub[2] ),.Z(_AES_ENC_n812 ) );
XOR2_X2 _AES_ENC_U1579  ( .A(_AES_ENC_sa00_sub[0] ), .B(_AES_ENC_sa11_sub[0] ), .Z(_AES_ENC_n1175 ) );
XOR2_X2 _AES_ENC_U1578  ( .A(_AES_ENC_sa22_sub[1] ), .B(_AES_ENC_sa33_sub[1] ), .Z(_AES_ENC_n1165 ) );
XOR2_X2 _AES_ENC_U1577  ( .A(_AES_ENC_n814 ), .B(_AES_ENC_n813 ), .Z(_AES_ENC_sa00_next[1]) );
XOR2_X2 _AES_ENC_U1576  ( .A(_AES_ENC_n1165 ), .B(_AES_ENC_n815 ), .Z(_AES_ENC_n813 ) );
XOR2_X2 _AES_ENC_U1575  ( .A(_AES_ENC_n1168 ), .B(_AES_ENC_n1175 ), .Z(_AES_ENC_n814 ) );
XOR2_X2 _AES_ENC_U1574  ( .A(_AES_ENC_w0[25] ), .B(_AES_ENC_sa11_sub[1] ),.Z(_AES_ENC_n815 ) );
XOR2_X2 _AES_ENC_U1573  ( .A(_AES_ENC_sa22_sub[0] ), .B(_AES_ENC_sa33_sub[0] ), .Z(_AES_ENC_n1166 ) );
XOR2_X2 _AES_ENC_U1572  ( .A(_AES_ENC_n817 ), .B(_AES_ENC_n816 ), .Z(_AES_ENC_sa00_next[0]) );
XOR2_X2 _AES_ENC_U1571  ( .A(_AES_ENC_n1168 ), .B(_AES_ENC_n1166 ), .Z(_AES_ENC_n816 ) );
XOR2_X2 _AES_ENC_U1570  ( .A(_AES_ENC_w0[24] ), .B(_AES_ENC_sa11_sub[0] ),.Z(_AES_ENC_n817 ) );
XOR2_X2 _AES_ENC_U1569  ( .A(_AES_ENC_n819 ), .B(_AES_ENC_n818 ), .Z(_AES_ENC_sa10_next[7]) );
XOR2_X2 _AES_ENC_U1568  ( .A(_AES_ENC_n1167 ), .B(_AES_ENC_n820 ), .Z(_AES_ENC_n818 ) );
XOR2_X2 _AES_ENC_U1567  ( .A(_AES_ENC_sa11_sub[6] ), .B(_AES_ENC_sa22_sub[6] ), .Z(_AES_ENC_n819 ) );
XOR2_X2 _AES_ENC_U1566  ( .A(_AES_ENC_w0[23] ), .B(_AES_ENC_sa00_sub[7] ),.Z(_AES_ENC_n820 ) );
XOR2_X2 _AES_ENC_U1565  ( .A(_AES_ENC_n822 ), .B(_AES_ENC_n821 ), .Z(_AES_ENC_sa10_next[6]) );
XOR2_X2 _AES_ENC_U1564  ( .A(_AES_ENC_n1160 ), .B(_AES_ENC_n823 ), .Z(_AES_ENC_n821 ) );
XOR2_X2 _AES_ENC_U1563  ( .A(_AES_ENC_sa11_sub[5] ), .B(_AES_ENC_sa22_sub[5] ), .Z(_AES_ENC_n822 ) );
XOR2_X2 _AES_ENC_U1562  ( .A(_AES_ENC_w0[22] ), .B(_AES_ENC_sa00_sub[6] ),.Z(_AES_ENC_n823 ) );
XOR2_X2 _AES_ENC_U1561  ( .A(_AES_ENC_n825 ), .B(_AES_ENC_n824 ), .Z(_AES_ENC_sa10_next[5]) );
XOR2_X2 _AES_ENC_U1560  ( .A(_AES_ENC_n1161 ), .B(_AES_ENC_n826 ), .Z(_AES_ENC_n824 ) );
XOR2_X2 _AES_ENC_U1559  ( .A(_AES_ENC_sa11_sub[4] ), .B(_AES_ENC_sa22_sub[4] ), .Z(_AES_ENC_n825 ) );
XOR2_X2 _AES_ENC_U1558  ( .A(_AES_ENC_w0[21] ), .B(_AES_ENC_sa00_sub[5] ),.Z(_AES_ENC_n826 ) );
XOR2_X2 _AES_ENC_U1557  ( .A(_AES_ENC_sa11_sub[7] ), .B(_AES_ENC_sa22_sub[7] ), .Z(_AES_ENC_n1159 ) );
XOR2_X2 _AES_ENC_U1556  ( .A(_AES_ENC_n828 ), .B(_AES_ENC_n827 ), .Z(_AES_ENC_sa10_next[4]) );
XOR2_X2 _AES_ENC_U1555  ( .A(_AES_ENC_n830 ), .B(_AES_ENC_n829 ), .Z(_AES_ENC_n827 ) );
XOR2_X2 _AES_ENC_U1554  ( .A(_AES_ENC_n1159 ), .B(_AES_ENC_n1162 ), .Z(_AES_ENC_n828 ) );
XOR2_X2 _AES_ENC_U1553  ( .A(_AES_ENC_sa11_sub[3] ), .B(_AES_ENC_sa22_sub[3] ), .Z(_AES_ENC_n829 ) );
XOR2_X2 _AES_ENC_U1552  ( .A(_AES_ENC_w0[20] ), .B(_AES_ENC_sa00_sub[4] ),.Z(_AES_ENC_n830 ) );
XOR2_X2 _AES_ENC_U1551  ( .A(_AES_ENC_n832 ), .B(_AES_ENC_n831 ), .Z(_AES_ENC_sa10_next[3]) );
XOR2_X2 _AES_ENC_U1550  ( .A(_AES_ENC_n834 ), .B(_AES_ENC_n833 ), .Z(_AES_ENC_n831 ) );
XOR2_X2 _AES_ENC_U1549  ( .A(_AES_ENC_n1159 ), .B(_AES_ENC_n1163 ), .Z(_AES_ENC_n832 ) );
XOR2_X2 _AES_ENC_U1548  ( .A(_AES_ENC_sa11_sub[2] ), .B(_AES_ENC_sa22_sub[2] ), .Z(_AES_ENC_n833 ) );
XOR2_X2 _AES_ENC_U1547  ( .A(_AES_ENC_w0[19] ), .B(_AES_ENC_sa00_sub[3] ),.Z(_AES_ENC_n834 ) );
XOR2_X2 _AES_ENC_U1546  ( .A(_AES_ENC_n836 ), .B(_AES_ENC_n835 ), .Z(_AES_ENC_sa10_next[2]) );
XOR2_X2 _AES_ENC_U1545  ( .A(_AES_ENC_n1164 ), .B(_AES_ENC_n837 ), .Z(_AES_ENC_n835 ) );
XOR2_X2 _AES_ENC_U1544  ( .A(_AES_ENC_sa11_sub[1] ), .B(_AES_ENC_sa22_sub[1] ), .Z(_AES_ENC_n836 ) );
XOR2_X2 _AES_ENC_U1543  ( .A(_AES_ENC_w0[18] ), .B(_AES_ENC_sa00_sub[2] ),.Z(_AES_ENC_n837 ) );
XOR2_X2 _AES_ENC_U1542  ( .A(_AES_ENC_n839 ), .B(_AES_ENC_n838 ), .Z(_AES_ENC_sa10_next[1]) );
XOR2_X2 _AES_ENC_U1541  ( .A(_AES_ENC_n841 ), .B(_AES_ENC_n840 ), .Z(_AES_ENC_n838 ) );
XOR2_X2 _AES_ENC_U1540  ( .A(_AES_ENC_n1159 ), .B(_AES_ENC_n1165 ), .Z(_AES_ENC_n839 ) );
XOR2_X2 _AES_ENC_U1539  ( .A(_AES_ENC_sa11_sub[0] ), .B(_AES_ENC_sa22_sub[0] ), .Z(_AES_ENC_n840 ) );
XOR2_X2 _AES_ENC_U1538  ( .A(_AES_ENC_w0[17] ), .B(_AES_ENC_sa00_sub[1] ),.Z(_AES_ENC_n841 ) );
XOR2_X2 _AES_ENC_U1537  ( .A(_AES_ENC_n843 ), .B(_AES_ENC_n842 ), .Z(_AES_ENC_sa10_next[0]) );
XOR2_X2 _AES_ENC_U1536  ( .A(_AES_ENC_n1159 ), .B(_AES_ENC_n1166 ), .Z(_AES_ENC_n842 ) );
XOR2_X2 _AES_ENC_U1535  ( .A(_AES_ENC_w0[16] ), .B(_AES_ENC_sa00_sub[0] ),.Z(_AES_ENC_n843 ) );
XOR2_X2 _AES_ENC_U1534  ( .A(_AES_ENC_n845 ), .B(_AES_ENC_n844 ), .Z(_AES_ENC_sa20_next[7]) );
XOR2_X2 _AES_ENC_U1533  ( .A(_AES_ENC_n1168 ), .B(_AES_ENC_n1160 ), .Z(_AES_ENC_n844 ) );
XOR2_X2 _AES_ENC_U1532  ( .A(_AES_ENC_w0[15] ), .B(_AES_ENC_sa33_sub[7] ),.Z(_AES_ENC_n845 ) );
XOR2_X2 _AES_ENC_U1531  ( .A(_AES_ENC_n847 ), .B(_AES_ENC_n846 ), .Z(_AES_ENC_sa20_next[6]) );
XOR2_X2 _AES_ENC_U1530  ( .A(_AES_ENC_n1169 ), .B(_AES_ENC_n1161 ), .Z(_AES_ENC_n846 ) );
XOR2_X2 _AES_ENC_U1529  ( .A(_AES_ENC_w0[14] ), .B(_AES_ENC_sa33_sub[6] ),.Z(_AES_ENC_n847 ) );
XOR2_X2 _AES_ENC_U1528  ( .A(_AES_ENC_n849 ), .B(_AES_ENC_n848 ), .Z(_AES_ENC_sa20_next[5]) );
XOR2_X2 _AES_ENC_U1527  ( .A(_AES_ENC_n1170 ), .B(_AES_ENC_n1162 ), .Z(_AES_ENC_n848 ) );
XOR2_X2 _AES_ENC_U1526  ( .A(_AES_ENC_w0[13] ), .B(_AES_ENC_sa33_sub[5] ),.Z(_AES_ENC_n849 ) );
XOR2_X2 _AES_ENC_U1525  ( .A(_AES_ENC_n851 ), .B(_AES_ENC_n850 ), .Z(_AES_ENC_sa20_next[4]) );
XOR2_X2 _AES_ENC_U1524  ( .A(_AES_ENC_n1163 ), .B(_AES_ENC_n852 ), .Z(_AES_ENC_n850 ) );
XOR2_X2 _AES_ENC_U1523  ( .A(_AES_ENC_n1167 ), .B(_AES_ENC_n1171 ), .Z(_AES_ENC_n851 ) );
XOR2_X2 _AES_ENC_U1522  ( .A(_AES_ENC_w0[12] ), .B(_AES_ENC_sa33_sub[4] ),.Z(_AES_ENC_n852 ) );
XOR2_X2 _AES_ENC_U1521  ( .A(_AES_ENC_n854 ), .B(_AES_ENC_n853 ), .Z(_AES_ENC_sa20_next[3]) );
XOR2_X2 _AES_ENC_U1520  ( .A(_AES_ENC_n1164 ), .B(_AES_ENC_n855 ), .Z(_AES_ENC_n853 ) );
XOR2_X2 _AES_ENC_U1519  ( .A(_AES_ENC_n1167 ), .B(_AES_ENC_n1172 ), .Z(_AES_ENC_n854 ) );
XOR2_X2 _AES_ENC_U1518  ( .A(_AES_ENC_w0[11] ), .B(_AES_ENC_sa33_sub[3] ),.Z(_AES_ENC_n855 ) );
XOR2_X2 _AES_ENC_U1517  ( .A(_AES_ENC_n857 ), .B(_AES_ENC_n856 ), .Z(_AES_ENC_sa20_next[2]) );
XOR2_X2 _AES_ENC_U1516  ( .A(_AES_ENC_n1173 ), .B(_AES_ENC_n1165 ), .Z(_AES_ENC_n856 ) );
XOR2_X2 _AES_ENC_U1515  ( .A(_AES_ENC_w0[10] ), .B(_AES_ENC_sa33_sub[2] ),.Z(_AES_ENC_n857 ) );
XOR2_X2 _AES_ENC_U1514  ( .A(_AES_ENC_n859 ), .B(_AES_ENC_n858 ), .Z(_AES_ENC_sa20_next[1]) );
XOR2_X2 _AES_ENC_U1513  ( .A(_AES_ENC_n1166 ), .B(_AES_ENC_n860 ), .Z(_AES_ENC_n858 ) );
XOR2_X2 _AES_ENC_U1512  ( .A(_AES_ENC_n1167 ), .B(_AES_ENC_n1174 ), .Z(_AES_ENC_n859 ) );
XOR2_X2 _AES_ENC_U1511  ( .A(_AES_ENC_w0[9] ), .B(_AES_ENC_sa33_sub[1] ),.Z(_AES_ENC_n860 ) );
XOR2_X2 _AES_ENC_U1510  ( .A(_AES_ENC_n862 ), .B(_AES_ENC_n861 ), .Z(_AES_ENC_sa20_next[0]) );
XOR2_X2 _AES_ENC_U1509  ( .A(_AES_ENC_n1167 ), .B(_AES_ENC_n1175 ), .Z(_AES_ENC_n861 ) );
XOR2_X2 _AES_ENC_U1508  ( .A(_AES_ENC_w0[8] ), .B(_AES_ENC_sa33_sub[0] ),.Z(_AES_ENC_n862 ) );
XOR2_X2 _AES_ENC_U1507  ( .A(_AES_ENC_n864 ), .B(_AES_ENC_n863 ), .Z(_AES_ENC_sa30_next[7]) );
XOR2_X2 _AES_ENC_U1506  ( .A(_AES_ENC_n1168 ), .B(_AES_ENC_n865 ), .Z(_AES_ENC_n863 ) );
XOR2_X2 _AES_ENC_U1505  ( .A(_AES_ENC_sa22_sub[7] ), .B(_AES_ENC_sa33_sub[6] ), .Z(_AES_ENC_n864 ) );
XOR2_X2 _AES_ENC_U1504  ( .A(_AES_ENC_w0[7] ), .B(_AES_ENC_sa00_sub[6] ),.Z(_AES_ENC_n865 ) );
XOR2_X2 _AES_ENC_U1503  ( .A(_AES_ENC_n867 ), .B(_AES_ENC_n866 ), .Z(_AES_ENC_sa30_next[6]) );
XOR2_X2 _AES_ENC_U1502  ( .A(_AES_ENC_n1169 ), .B(_AES_ENC_n868 ), .Z(_AES_ENC_n866 ) );
XOR2_X2 _AES_ENC_U1501  ( .A(_AES_ENC_sa22_sub[6] ), .B(_AES_ENC_sa33_sub[5] ), .Z(_AES_ENC_n867 ) );
XOR2_X2 _AES_ENC_U1500  ( .A(_AES_ENC_w0[6] ), .B(_AES_ENC_sa00_sub[5] ),.Z(_AES_ENC_n868 ) );
XOR2_X2 _AES_ENC_U1499  ( .A(_AES_ENC_n870 ), .B(_AES_ENC_n869 ), .Z(_AES_ENC_sa30_next[5]) );
XOR2_X2 _AES_ENC_U1498  ( .A(_AES_ENC_n1170 ), .B(_AES_ENC_n871 ), .Z(_AES_ENC_n869 ) );
XOR2_X2 _AES_ENC_U1497  ( .A(_AES_ENC_sa22_sub[5] ), .B(_AES_ENC_sa33_sub[4] ), .Z(_AES_ENC_n870 ) );
XOR2_X2 _AES_ENC_U1496  ( .A(_AES_ENC_w0[5] ), .B(_AES_ENC_sa00_sub[4] ),.Z(_AES_ENC_n871 ) );
XOR2_X2 _AES_ENC_U1495  ( .A(_AES_ENC_sa00_sub[7] ), .B(_AES_ENC_sa33_sub[7] ), .Z(_AES_ENC_n1176 ) );
XOR2_X2 _AES_ENC_U1494  ( .A(_AES_ENC_n873 ), .B(_AES_ENC_n872 ), .Z(_AES_ENC_sa30_next[4]) );
XOR2_X2 _AES_ENC_U1493  ( .A(_AES_ENC_n875 ), .B(_AES_ENC_n874 ), .Z(_AES_ENC_n872 ) );
XOR2_X2 _AES_ENC_U1492  ( .A(_AES_ENC_n1176 ), .B(_AES_ENC_n1171 ), .Z(_AES_ENC_n873 ) );
XOR2_X2 _AES_ENC_U1491  ( .A(_AES_ENC_sa22_sub[4] ), .B(_AES_ENC_sa33_sub[3] ), .Z(_AES_ENC_n874 ) );
XOR2_X2 _AES_ENC_U1490  ( .A(_AES_ENC_w0[4] ), .B(_AES_ENC_sa00_sub[3] ),.Z(_AES_ENC_n875 ) );
XOR2_X2 _AES_ENC_U1489  ( .A(_AES_ENC_n877 ), .B(_AES_ENC_n876 ), .Z(_AES_ENC_sa30_next[3]) );
XOR2_X2 _AES_ENC_U1488  ( .A(_AES_ENC_n879 ), .B(_AES_ENC_n878 ), .Z(_AES_ENC_n876 ) );
XOR2_X2 _AES_ENC_U1487  ( .A(_AES_ENC_n1176 ), .B(_AES_ENC_n1172 ), .Z(_AES_ENC_n877 ) );
XOR2_X2 _AES_ENC_U1486  ( .A(_AES_ENC_sa22_sub[3] ), .B(_AES_ENC_sa33_sub[2] ), .Z(_AES_ENC_n878 ) );
XOR2_X2 _AES_ENC_U1485  ( .A(_AES_ENC_w0[3] ), .B(_AES_ENC_sa00_sub[2] ),.Z(_AES_ENC_n879 ) );
XOR2_X2 _AES_ENC_U1484  ( .A(_AES_ENC_n881 ), .B(_AES_ENC_n880 ), .Z(_AES_ENC_sa30_next[2]) );
XOR2_X2 _AES_ENC_U1483  ( .A(_AES_ENC_n1173 ), .B(_AES_ENC_n882 ), .Z(_AES_ENC_n880 ) );
XOR2_X2 _AES_ENC_U1482  ( .A(_AES_ENC_sa22_sub[2] ), .B(_AES_ENC_sa33_sub[1] ), .Z(_AES_ENC_n881 ) );
XOR2_X2 _AES_ENC_U1481  ( .A(_AES_ENC_w0[2] ), .B(_AES_ENC_sa00_sub[1] ),.Z(_AES_ENC_n882 ) );
XOR2_X2 _AES_ENC_U1480  ( .A(_AES_ENC_n884 ), .B(_AES_ENC_n883 ), .Z(_AES_ENC_sa30_next[1]) );
XOR2_X2 _AES_ENC_U1479  ( .A(_AES_ENC_n886 ), .B(_AES_ENC_n885 ), .Z(_AES_ENC_n883 ) );
XOR2_X2 _AES_ENC_U1478  ( .A(_AES_ENC_n1176 ), .B(_AES_ENC_n1174 ), .Z(_AES_ENC_n884 ) );
XOR2_X2 _AES_ENC_U1477  ( .A(_AES_ENC_sa22_sub[1] ), .B(_AES_ENC_sa33_sub[0] ), .Z(_AES_ENC_n885 ) );
XOR2_X2 _AES_ENC_U1476  ( .A(_AES_ENC_w0[1] ), .B(_AES_ENC_sa00_sub[0] ),.Z(_AES_ENC_n886 ) );
XOR2_X2 _AES_ENC_U1475  ( .A(_AES_ENC_n888 ), .B(_AES_ENC_n887 ), .Z(_AES_ENC_sa30_next[0]) );
XOR2_X2 _AES_ENC_U1474  ( .A(_AES_ENC_n1176 ), .B(_AES_ENC_n1175 ), .Z(_AES_ENC_n887 ) );
XOR2_X2 _AES_ENC_U1473  ( .A(_AES_ENC_w0[0] ), .B(_AES_ENC_sa22_sub[0] ),.Z(_AES_ENC_n888 ) );
XOR2_X2 _AES_ENC_U1472  ( .A(_AES_ENC_sa23_sub[7] ), .B(_AES_ENC_sa30_sub[7] ), .Z(_AES_ENC_n1185 ) );
XOR2_X2 _AES_ENC_U1471  ( .A(_AES_ENC_sa01_sub[6] ), .B(_AES_ENC_sa12_sub[6] ), .Z(_AES_ENC_n1187 ) );
XOR2_X2 _AES_ENC_U1470  ( .A(_AES_ENC_n890 ), .B(_AES_ENC_n889 ), .Z(_AES_ENC_sa01_next[7]) );
XOR2_X2 _AES_ENC_U1469  ( .A(_AES_ENC_n1185 ), .B(_AES_ENC_n1187 ), .Z(_AES_ENC_n889 ) );
XOR2_X2 _AES_ENC_U1468  ( .A(_AES_ENC_w1[31] ), .B(_AES_ENC_sa12_sub[7] ),.Z(_AES_ENC_n890 ) );
XOR2_X2 _AES_ENC_U1467  ( .A(_AES_ENC_sa01_sub[5] ), .B(_AES_ENC_sa12_sub[5] ), .Z(_AES_ENC_n1188 ) );
XOR2_X2 _AES_ENC_U1466  ( .A(_AES_ENC_sa23_sub[6] ), .B(_AES_ENC_sa30_sub[6] ), .Z(_AES_ENC_n1178 ) );
XOR2_X2 _AES_ENC_U1465  ( .A(_AES_ENC_n892 ), .B(_AES_ENC_n891 ), .Z(_AES_ENC_sa01_next[6]) );
XOR2_X2 _AES_ENC_U1464  ( .A(_AES_ENC_n1188 ), .B(_AES_ENC_n1178 ), .Z(_AES_ENC_n891 ) );
XOR2_X2 _AES_ENC_U1463  ( .A(_AES_ENC_w1[30] ), .B(_AES_ENC_sa12_sub[6] ),.Z(_AES_ENC_n892 ) );
XOR2_X2 _AES_ENC_U1462  ( .A(_AES_ENC_sa01_sub[4] ), .B(_AES_ENC_sa12_sub[4] ), .Z(_AES_ENC_n1189 ) );
XOR2_X2 _AES_ENC_U1461  ( .A(_AES_ENC_sa23_sub[5] ), .B(_AES_ENC_sa30_sub[5] ), .Z(_AES_ENC_n1179 ) );
XOR2_X2 _AES_ENC_U1460  ( .A(_AES_ENC_n894 ), .B(_AES_ENC_n893 ), .Z(_AES_ENC_sa01_next[5]) );
XOR2_X2 _AES_ENC_U1459  ( .A(_AES_ENC_n1189 ), .B(_AES_ENC_n1179 ), .Z(_AES_ENC_n893 ) );
XOR2_X2 _AES_ENC_U1458  ( .A(_AES_ENC_w1[29] ), .B(_AES_ENC_sa12_sub[5] ),.Z(_AES_ENC_n894 ) );
XOR2_X2 _AES_ENC_U1457  ( .A(_AES_ENC_sa01_sub[7] ), .B(_AES_ENC_sa12_sub[7] ), .Z(_AES_ENC_n1186 ) );
XOR2_X2 _AES_ENC_U1456  ( .A(_AES_ENC_sa01_sub[3] ), .B(_AES_ENC_sa12_sub[3] ), .Z(_AES_ENC_n1190 ) );
XOR2_X2 _AES_ENC_U1455  ( .A(_AES_ENC_sa23_sub[4] ), .B(_AES_ENC_sa30_sub[4] ), .Z(_AES_ENC_n1180 ) );
XOR2_X2 _AES_ENC_U1454  ( .A(_AES_ENC_n896 ), .B(_AES_ENC_n895 ), .Z(_AES_ENC_sa01_next[4]) );
XOR2_X2 _AES_ENC_U1453  ( .A(_AES_ENC_n1180 ), .B(_AES_ENC_n897 ), .Z(_AES_ENC_n895 ) );
XOR2_X2 _AES_ENC_U1452  ( .A(_AES_ENC_n1186 ), .B(_AES_ENC_n1190 ), .Z(_AES_ENC_n896 ) );
XOR2_X2 _AES_ENC_U1451  ( .A(_AES_ENC_w1[28] ), .B(_AES_ENC_sa12_sub[4] ),.Z(_AES_ENC_n897 ) );
XOR2_X2 _AES_ENC_U1450  ( .A(_AES_ENC_sa01_sub[2] ), .B(_AES_ENC_sa12_sub[2] ), .Z(_AES_ENC_n1191 ) );
XOR2_X2 _AES_ENC_U1449  ( .A(_AES_ENC_sa23_sub[3] ), .B(_AES_ENC_sa30_sub[3] ), .Z(_AES_ENC_n1181 ) );
XOR2_X2 _AES_ENC_U1448  ( .A(_AES_ENC_n899 ), .B(_AES_ENC_n898 ), .Z(_AES_ENC_sa01_next[3]) );
XOR2_X2 _AES_ENC_U1447  ( .A(_AES_ENC_n1181 ), .B(_AES_ENC_n900 ), .Z(_AES_ENC_n898 ) );
XOR2_X2 _AES_ENC_U1446  ( .A(_AES_ENC_n1186 ), .B(_AES_ENC_n1191 ), .Z(_AES_ENC_n899 ) );
XOR2_X2 _AES_ENC_U1445  ( .A(_AES_ENC_w1[27] ), .B(_AES_ENC_sa12_sub[3] ),.Z(_AES_ENC_n900 ) );
XOR2_X2 _AES_ENC_U1444  ( .A(_AES_ENC_sa01_sub[1] ), .B(_AES_ENC_sa12_sub[1] ), .Z(_AES_ENC_n1192 ) );
XOR2_X2 _AES_ENC_U1443  ( .A(_AES_ENC_sa23_sub[2] ), .B(_AES_ENC_sa30_sub[2] ), .Z(_AES_ENC_n1182 ) );
XOR2_X2 _AES_ENC_U1442  ( .A(_AES_ENC_n902 ), .B(_AES_ENC_n901 ), .Z(_AES_ENC_sa01_next[2]) );
XOR2_X2 _AES_ENC_U1441  ( .A(_AES_ENC_n1192 ), .B(_AES_ENC_n1182 ), .Z(_AES_ENC_n901 ) );
XOR2_X2 _AES_ENC_U1440  ( .A(_AES_ENC_w1[26] ), .B(_AES_ENC_sa12_sub[2] ),.Z(_AES_ENC_n902 ) );
XOR2_X2 _AES_ENC_U1439  ( .A(_AES_ENC_sa01_sub[0] ), .B(_AES_ENC_sa12_sub[0] ), .Z(_AES_ENC_n1193 ) );
XOR2_X2 _AES_ENC_U1438  ( .A(_AES_ENC_sa23_sub[1] ), .B(_AES_ENC_sa30_sub[1] ), .Z(_AES_ENC_n1183 ) );
XOR2_X2 _AES_ENC_U1437  ( .A(_AES_ENC_n904 ), .B(_AES_ENC_n903 ), .Z(_AES_ENC_sa01_next[1]) );
XOR2_X2 _AES_ENC_U1436  ( .A(_AES_ENC_n1183 ), .B(_AES_ENC_n905 ), .Z(_AES_ENC_n903 ) );
XOR2_X2 _AES_ENC_U1435  ( .A(_AES_ENC_n1186 ), .B(_AES_ENC_n1193 ), .Z(_AES_ENC_n904 ) );
XOR2_X2 _AES_ENC_U1434  ( .A(_AES_ENC_w1[25] ), .B(_AES_ENC_sa12_sub[1] ),.Z(_AES_ENC_n905 ) );
XOR2_X2 _AES_ENC_U1433  ( .A(_AES_ENC_sa23_sub[0] ), .B(_AES_ENC_sa30_sub[0] ), .Z(_AES_ENC_n1184 ) );
XOR2_X2 _AES_ENC_U1432  ( .A(_AES_ENC_n907 ), .B(_AES_ENC_n906 ), .Z(_AES_ENC_sa01_next[0]) );
XOR2_X2 _AES_ENC_U1431  ( .A(_AES_ENC_n1186 ), .B(_AES_ENC_n1184 ), .Z(_AES_ENC_n906 ) );
XOR2_X2 _AES_ENC_U1430  ( .A(_AES_ENC_w1[24] ), .B(_AES_ENC_sa12_sub[0] ),.Z(_AES_ENC_n907 ) );
XOR2_X2 _AES_ENC_U1429  ( .A(_AES_ENC_n909 ), .B(_AES_ENC_n908 ), .Z(_AES_ENC_sa11_next[7]) );
XOR2_X2 _AES_ENC_U1428  ( .A(_AES_ENC_n1185 ), .B(_AES_ENC_n910 ), .Z(_AES_ENC_n908 ) );
XOR2_X2 _AES_ENC_U1427  ( .A(_AES_ENC_sa12_sub[6] ), .B(_AES_ENC_sa23_sub[6] ), .Z(_AES_ENC_n909 ) );
XOR2_X2 _AES_ENC_U1426  ( .A(_AES_ENC_w1[23] ), .B(_AES_ENC_sa01_sub[7] ),.Z(_AES_ENC_n910 ) );
XOR2_X2 _AES_ENC_U1425  ( .A(_AES_ENC_n912 ), .B(_AES_ENC_n911 ), .Z(_AES_ENC_sa11_next[6]) );
XOR2_X2 _AES_ENC_U1424  ( .A(_AES_ENC_n1178 ), .B(_AES_ENC_n913 ), .Z(_AES_ENC_n911 ) );
XOR2_X2 _AES_ENC_U1423  ( .A(_AES_ENC_sa12_sub[5] ), .B(_AES_ENC_sa23_sub[5] ), .Z(_AES_ENC_n912 ) );
XOR2_X2 _AES_ENC_U1422  ( .A(_AES_ENC_w1[22] ), .B(_AES_ENC_sa01_sub[6] ),.Z(_AES_ENC_n913 ) );
XOR2_X2 _AES_ENC_U1421  ( .A(_AES_ENC_n915 ), .B(_AES_ENC_n914 ), .Z(_AES_ENC_sa11_next[5]) );
XOR2_X2 _AES_ENC_U1420  ( .A(_AES_ENC_n1179 ), .B(_AES_ENC_n916 ), .Z(_AES_ENC_n914 ) );
XOR2_X2 _AES_ENC_U1419  ( .A(_AES_ENC_sa12_sub[4] ), .B(_AES_ENC_sa23_sub[4] ), .Z(_AES_ENC_n915 ) );
XOR2_X2 _AES_ENC_U1418  ( .A(_AES_ENC_w1[21] ), .B(_AES_ENC_sa01_sub[5] ),.Z(_AES_ENC_n916 ) );
XOR2_X2 _AES_ENC_U1417  ( .A(_AES_ENC_sa12_sub[7] ), .B(_AES_ENC_sa23_sub[7] ), .Z(_AES_ENC_n1177 ) );
XOR2_X2 _AES_ENC_U1416  ( .A(_AES_ENC_n918 ), .B(_AES_ENC_n917 ), .Z(_AES_ENC_sa11_next[4]) );
XOR2_X2 _AES_ENC_U1415  ( .A(_AES_ENC_n920 ), .B(_AES_ENC_n919 ), .Z(_AES_ENC_n917 ) );
XOR2_X2 _AES_ENC_U1414  ( .A(_AES_ENC_n1177 ), .B(_AES_ENC_n1180 ), .Z(_AES_ENC_n918 ) );
XOR2_X2 _AES_ENC_U1413  ( .A(_AES_ENC_sa12_sub[3] ), .B(_AES_ENC_sa23_sub[3] ), .Z(_AES_ENC_n919 ) );
XOR2_X2 _AES_ENC_U1412  ( .A(_AES_ENC_w1[20] ), .B(_AES_ENC_sa01_sub[4] ),.Z(_AES_ENC_n920 ) );
XOR2_X2 _AES_ENC_U1411  ( .A(_AES_ENC_n922 ), .B(_AES_ENC_n921 ), .Z(_AES_ENC_sa11_next[3]) );
XOR2_X2 _AES_ENC_U1410  ( .A(_AES_ENC_n924 ), .B(_AES_ENC_n923 ), .Z(_AES_ENC_n921 ) );
XOR2_X2 _AES_ENC_U1409  ( .A(_AES_ENC_n1177 ), .B(_AES_ENC_n1181 ), .Z(_AES_ENC_n922 ) );
XOR2_X2 _AES_ENC_U1408  ( .A(_AES_ENC_sa12_sub[2] ), .B(_AES_ENC_sa23_sub[2] ), .Z(_AES_ENC_n923 ) );
XOR2_X2 _AES_ENC_U1407  ( .A(_AES_ENC_w1[19] ), .B(_AES_ENC_sa01_sub[3] ),.Z(_AES_ENC_n924 ) );
XOR2_X2 _AES_ENC_U1406  ( .A(_AES_ENC_n926 ), .B(_AES_ENC_n925 ), .Z(_AES_ENC_sa11_next[2]) );
XOR2_X2 _AES_ENC_U1405  ( .A(_AES_ENC_n1182 ), .B(_AES_ENC_n927 ), .Z(_AES_ENC_n925 ) );
XOR2_X2 _AES_ENC_U1404  ( .A(_AES_ENC_sa12_sub[1] ), .B(_AES_ENC_sa23_sub[1] ), .Z(_AES_ENC_n926 ) );
XOR2_X2 _AES_ENC_U1403  ( .A(_AES_ENC_w1[18] ), .B(_AES_ENC_sa01_sub[2] ),.Z(_AES_ENC_n927 ) );
XOR2_X2 _AES_ENC_U1402  ( .A(_AES_ENC_n929 ), .B(_AES_ENC_n928 ), .Z(_AES_ENC_sa11_next[1]) );
XOR2_X2 _AES_ENC_U1401  ( .A(_AES_ENC_n931 ), .B(_AES_ENC_n930 ), .Z(_AES_ENC_n928 ) );
XOR2_X2 _AES_ENC_U1400  ( .A(_AES_ENC_n1177 ), .B(_AES_ENC_n1183 ), .Z(_AES_ENC_n929 ) );
XOR2_X2 _AES_ENC_U1399  ( .A(_AES_ENC_sa12_sub[0] ), .B(_AES_ENC_sa23_sub[0] ), .Z(_AES_ENC_n930 ) );
XOR2_X2 _AES_ENC_U1398  ( .A(_AES_ENC_w1[17] ), .B(_AES_ENC_sa01_sub[1] ),.Z(_AES_ENC_n931 ) );
XOR2_X2 _AES_ENC_U1397  ( .A(_AES_ENC_n933 ), .B(_AES_ENC_n932 ), .Z(_AES_ENC_sa11_next[0]) );
XOR2_X2 _AES_ENC_U1396  ( .A(_AES_ENC_n1177 ), .B(_AES_ENC_n1184 ), .Z(_AES_ENC_n932 ) );
XOR2_X2 _AES_ENC_U1395  ( .A(_AES_ENC_w1[16] ), .B(_AES_ENC_sa01_sub[0] ),.Z(_AES_ENC_n933 ) );
XOR2_X2 _AES_ENC_U1394  ( .A(_AES_ENC_n935 ), .B(_AES_ENC_n934 ), .Z(_AES_ENC_sa21_next[7]) );
XOR2_X2 _AES_ENC_U1393  ( .A(_AES_ENC_n1186 ), .B(_AES_ENC_n1178 ), .Z(_AES_ENC_n934 ) );
XOR2_X2 _AES_ENC_U1392  ( .A(_AES_ENC_w1[15] ), .B(_AES_ENC_sa30_sub[7] ),.Z(_AES_ENC_n935 ) );
XOR2_X2 _AES_ENC_U1391  ( .A(_AES_ENC_n937 ), .B(_AES_ENC_n936 ), .Z(_AES_ENC_sa21_next[6]) );
XOR2_X2 _AES_ENC_U1390  ( .A(_AES_ENC_n1187 ), .B(_AES_ENC_n1179 ), .Z(_AES_ENC_n936 ) );
XOR2_X2 _AES_ENC_U1389  ( .A(_AES_ENC_w1[14] ), .B(_AES_ENC_sa30_sub[6] ),.Z(_AES_ENC_n937 ) );
XOR2_X2 _AES_ENC_U1388  ( .A(_AES_ENC_n939 ), .B(_AES_ENC_n938 ), .Z(_AES_ENC_sa21_next[5]) );
XOR2_X2 _AES_ENC_U1387  ( .A(_AES_ENC_n1188 ), .B(_AES_ENC_n1180 ), .Z(_AES_ENC_n938 ) );
XOR2_X2 _AES_ENC_U1386  ( .A(_AES_ENC_w1[13] ), .B(_AES_ENC_sa30_sub[5] ),.Z(_AES_ENC_n939 ) );
XOR2_X2 _AES_ENC_U1385  ( .A(_AES_ENC_n941 ), .B(_AES_ENC_n940 ), .Z(_AES_ENC_sa21_next[4]) );
XOR2_X2 _AES_ENC_U1384  ( .A(_AES_ENC_n1181 ), .B(_AES_ENC_n942 ), .Z(_AES_ENC_n940 ) );
XOR2_X2 _AES_ENC_U1383  ( .A(_AES_ENC_n1185 ), .B(_AES_ENC_n1189 ), .Z(_AES_ENC_n941 ) );
XOR2_X2 _AES_ENC_U1382  ( .A(_AES_ENC_w1[12] ), .B(_AES_ENC_sa30_sub[4] ),.Z(_AES_ENC_n942 ) );
XOR2_X2 _AES_ENC_U1381  ( .A(_AES_ENC_n944 ), .B(_AES_ENC_n943 ), .Z(_AES_ENC_sa21_next[3]) );
XOR2_X2 _AES_ENC_U1380  ( .A(_AES_ENC_n1182 ), .B(_AES_ENC_n945 ), .Z(_AES_ENC_n943 ) );
XOR2_X2 _AES_ENC_U1379  ( .A(_AES_ENC_n1185 ), .B(_AES_ENC_n1190 ), .Z(_AES_ENC_n944 ) );
XOR2_X2 _AES_ENC_U1378  ( .A(_AES_ENC_w1[11] ), .B(_AES_ENC_sa30_sub[3] ),.Z(_AES_ENC_n945 ) );
XOR2_X2 _AES_ENC_U1377  ( .A(_AES_ENC_n947 ), .B(_AES_ENC_n946 ), .Z(_AES_ENC_sa21_next[2]) );
XOR2_X2 _AES_ENC_U1376  ( .A(_AES_ENC_n1191 ), .B(_AES_ENC_n1183 ), .Z(_AES_ENC_n946 ) );
XOR2_X2 _AES_ENC_U1375  ( .A(_AES_ENC_w1[10] ), .B(_AES_ENC_sa30_sub[2] ),.Z(_AES_ENC_n947 ) );
XOR2_X2 _AES_ENC_U1374  ( .A(_AES_ENC_n949 ), .B(_AES_ENC_n948 ), .Z(_AES_ENC_sa21_next[1]) );
XOR2_X2 _AES_ENC_U1373  ( .A(_AES_ENC_n1184 ), .B(_AES_ENC_n950 ), .Z(_AES_ENC_n948 ) );
XOR2_X2 _AES_ENC_U1372  ( .A(_AES_ENC_n1185 ), .B(_AES_ENC_n1192 ), .Z(_AES_ENC_n949 ) );
XOR2_X2 _AES_ENC_U1371  ( .A(_AES_ENC_w1[9] ), .B(_AES_ENC_sa30_sub[1] ),.Z(_AES_ENC_n950 ) );
XOR2_X2 _AES_ENC_U1370  ( .A(_AES_ENC_n952 ), .B(_AES_ENC_n951 ), .Z(_AES_ENC_sa21_next[0]) );
XOR2_X2 _AES_ENC_U1369  ( .A(_AES_ENC_n1185 ), .B(_AES_ENC_n1193 ), .Z(_AES_ENC_n951 ) );
XOR2_X2 _AES_ENC_U1368  ( .A(_AES_ENC_w1[8] ), .B(_AES_ENC_sa30_sub[0] ),.Z(_AES_ENC_n952 ) );
XOR2_X2 _AES_ENC_U1367  ( .A(_AES_ENC_n954 ), .B(_AES_ENC_n953 ), .Z(_AES_ENC_sa31_next[7]) );
XOR2_X2 _AES_ENC_U1366  ( .A(_AES_ENC_n1186 ), .B(_AES_ENC_n955 ), .Z(_AES_ENC_n953 ) );
XOR2_X2 _AES_ENC_U1365  ( .A(_AES_ENC_sa23_sub[7] ), .B(_AES_ENC_sa30_sub[6] ), .Z(_AES_ENC_n954 ) );
XOR2_X2 _AES_ENC_U1364  ( .A(_AES_ENC_w1[7] ), .B(_AES_ENC_sa01_sub[6] ),.Z(_AES_ENC_n955 ) );
XOR2_X2 _AES_ENC_U1363  ( .A(_AES_ENC_n957 ), .B(_AES_ENC_n956 ), .Z(_AES_ENC_sa31_next[6]) );
XOR2_X2 _AES_ENC_U1362  ( .A(_AES_ENC_n1187 ), .B(_AES_ENC_n958 ), .Z(_AES_ENC_n956 ) );
XOR2_X2 _AES_ENC_U1361  ( .A(_AES_ENC_sa23_sub[6] ), .B(_AES_ENC_sa30_sub[5] ), .Z(_AES_ENC_n957 ) );
XOR2_X2 _AES_ENC_U1360  ( .A(_AES_ENC_w1[6] ), .B(_AES_ENC_sa01_sub[5] ),.Z(_AES_ENC_n958 ) );
XOR2_X2 _AES_ENC_U1359  ( .A(_AES_ENC_n960 ), .B(_AES_ENC_n959 ), .Z(_AES_ENC_sa31_next[5]) );
XOR2_X2 _AES_ENC_U1358  ( .A(_AES_ENC_n1188 ), .B(_AES_ENC_n961 ), .Z(_AES_ENC_n959 ) );
XOR2_X2 _AES_ENC_U1357  ( .A(_AES_ENC_sa23_sub[5] ), .B(_AES_ENC_sa30_sub[4] ), .Z(_AES_ENC_n960 ) );
XOR2_X2 _AES_ENC_U1356  ( .A(_AES_ENC_w1[5] ), .B(_AES_ENC_sa01_sub[4] ),.Z(_AES_ENC_n961 ) );
XOR2_X2 _AES_ENC_U1355  ( .A(_AES_ENC_sa01_sub[7] ), .B(_AES_ENC_sa30_sub[7] ), .Z(_AES_ENC_n1194 ) );
XOR2_X2 _AES_ENC_U1354  ( .A(_AES_ENC_n963 ), .B(_AES_ENC_n962 ), .Z(_AES_ENC_sa31_next[4]) );
XOR2_X2 _AES_ENC_U1353  ( .A(_AES_ENC_n965 ), .B(_AES_ENC_n964 ), .Z(_AES_ENC_n962 ) );
XOR2_X2 _AES_ENC_U1352  ( .A(_AES_ENC_n1194 ), .B(_AES_ENC_n1189 ), .Z(_AES_ENC_n963 ) );
XOR2_X2 _AES_ENC_U1351  ( .A(_AES_ENC_sa23_sub[4] ), .B(_AES_ENC_sa30_sub[3] ), .Z(_AES_ENC_n964 ) );
XOR2_X2 _AES_ENC_U1350  ( .A(_AES_ENC_w1[4] ), .B(_AES_ENC_sa01_sub[3] ),.Z(_AES_ENC_n965 ) );
XOR2_X2 _AES_ENC_U1349  ( .A(_AES_ENC_n967 ), .B(_AES_ENC_n966 ), .Z(_AES_ENC_sa31_next[3]) );
XOR2_X2 _AES_ENC_U1348  ( .A(_AES_ENC_n969 ), .B(_AES_ENC_n968 ), .Z(_AES_ENC_n966 ) );
XOR2_X2 _AES_ENC_U1347  ( .A(_AES_ENC_n1194 ), .B(_AES_ENC_n1190 ), .Z(_AES_ENC_n967 ) );
XOR2_X2 _AES_ENC_U1346  ( .A(_AES_ENC_sa23_sub[3] ), .B(_AES_ENC_sa30_sub[2] ), .Z(_AES_ENC_n968 ) );
XOR2_X2 _AES_ENC_U1345  ( .A(_AES_ENC_w1[3] ), .B(_AES_ENC_sa01_sub[2] ),.Z(_AES_ENC_n969 ) );
XOR2_X2 _AES_ENC_U1344  ( .A(_AES_ENC_n971 ), .B(_AES_ENC_n970 ), .Z(_AES_ENC_sa31_next[2]) );
XOR2_X2 _AES_ENC_U1343  ( .A(_AES_ENC_n1191 ), .B(_AES_ENC_n972 ), .Z(_AES_ENC_n970 ) );
XOR2_X2 _AES_ENC_U1342  ( .A(_AES_ENC_sa23_sub[2] ), .B(_AES_ENC_sa30_sub[1] ), .Z(_AES_ENC_n971 ) );
XOR2_X2 _AES_ENC_U1341  ( .A(_AES_ENC_w1[2] ), .B(_AES_ENC_sa01_sub[1] ),.Z(_AES_ENC_n972 ) );
XOR2_X2 _AES_ENC_U1340  ( .A(_AES_ENC_n974 ), .B(_AES_ENC_n973 ), .Z(_AES_ENC_sa31_next[1]) );
XOR2_X2 _AES_ENC_U1339  ( .A(_AES_ENC_n976 ), .B(_AES_ENC_n975 ), .Z(_AES_ENC_n973 ) );
XOR2_X2 _AES_ENC_U1338  ( .A(_AES_ENC_n1194 ), .B(_AES_ENC_n1192 ), .Z(_AES_ENC_n974 ) );
XOR2_X2 _AES_ENC_U1337  ( .A(_AES_ENC_sa23_sub[1] ), .B(_AES_ENC_sa30_sub[0] ), .Z(_AES_ENC_n975 ) );
XOR2_X2 _AES_ENC_U1336  ( .A(_AES_ENC_w1[1] ), .B(_AES_ENC_sa01_sub[0] ),.Z(_AES_ENC_n976 ) );
XOR2_X2 _AES_ENC_U1335  ( .A(_AES_ENC_n978 ), .B(_AES_ENC_n977 ), .Z(_AES_ENC_sa31_next[0]) );
XOR2_X2 _AES_ENC_U1334  ( .A(_AES_ENC_n1194 ), .B(_AES_ENC_n1193 ), .Z(_AES_ENC_n977 ) );
XOR2_X2 _AES_ENC_U1333  ( .A(_AES_ENC_w1[0] ), .B(_AES_ENC_sa23_sub[0] ),.Z(_AES_ENC_n978 ) );
XOR2_X2 _AES_ENC_U1332  ( .A(_AES_ENC_sa20_sub[7] ), .B(_AES_ENC_sa31_sub[7] ), .Z(_AES_ENC_n1203 ) );
XOR2_X2 _AES_ENC_U1331  ( .A(_AES_ENC_sa02_sub[6] ), .B(_AES_ENC_sa13_sub[6] ), .Z(_AES_ENC_n1205 ) );
XOR2_X2 _AES_ENC_U1330  ( .A(_AES_ENC_n980 ), .B(_AES_ENC_n979 ), .Z(_AES_ENC_sa02_next[7]) );
XOR2_X2 _AES_ENC_U1329  ( .A(_AES_ENC_n1203 ), .B(_AES_ENC_n1205 ), .Z(_AES_ENC_n979 ) );
XOR2_X2 _AES_ENC_U1328  ( .A(_AES_ENC_w2[31] ), .B(_AES_ENC_sa13_sub[7] ),.Z(_AES_ENC_n980 ) );
XOR2_X2 _AES_ENC_U1327  ( .A(_AES_ENC_sa02_sub[5] ), .B(_AES_ENC_sa13_sub[5] ), .Z(_AES_ENC_n1206 ) );
XOR2_X2 _AES_ENC_U1326  ( .A(_AES_ENC_sa20_sub[6] ), .B(_AES_ENC_sa31_sub[6] ), .Z(_AES_ENC_n1196 ) );
XOR2_X2 _AES_ENC_U1325  ( .A(_AES_ENC_n982 ), .B(_AES_ENC_n981 ), .Z(_AES_ENC_sa02_next[6]) );
XOR2_X2 _AES_ENC_U1324  ( .A(_AES_ENC_n1206 ), .B(_AES_ENC_n1196 ), .Z(_AES_ENC_n981 ) );
XOR2_X2 _AES_ENC_U1323  ( .A(_AES_ENC_w2[30] ), .B(_AES_ENC_sa13_sub[6] ),.Z(_AES_ENC_n982 ) );
XOR2_X2 _AES_ENC_U1322  ( .A(_AES_ENC_sa02_sub[4] ), .B(_AES_ENC_sa13_sub[4] ), .Z(_AES_ENC_n1207 ) );
XOR2_X2 _AES_ENC_U1321  ( .A(_AES_ENC_sa20_sub[5] ), .B(_AES_ENC_sa31_sub[5] ), .Z(_AES_ENC_n1197 ) );
XOR2_X2 _AES_ENC_U1320  ( .A(_AES_ENC_n984 ), .B(_AES_ENC_n983 ), .Z(_AES_ENC_sa02_next[5]) );
XOR2_X2 _AES_ENC_U1319  ( .A(_AES_ENC_n1207 ), .B(_AES_ENC_n1197 ), .Z(_AES_ENC_n983 ) );
XOR2_X2 _AES_ENC_U1318  ( .A(_AES_ENC_w2[29] ), .B(_AES_ENC_sa13_sub[5] ),.Z(_AES_ENC_n984 ) );
XOR2_X2 _AES_ENC_U1317  ( .A(_AES_ENC_sa02_sub[7] ), .B(_AES_ENC_sa13_sub[7] ), .Z(_AES_ENC_n1204 ) );
XOR2_X2 _AES_ENC_U1316  ( .A(_AES_ENC_sa02_sub[3] ), .B(_AES_ENC_sa13_sub[3] ), .Z(_AES_ENC_n1208 ) );
XOR2_X2 _AES_ENC_U1315  ( .A(_AES_ENC_sa20_sub[4] ), .B(_AES_ENC_sa31_sub[4] ), .Z(_AES_ENC_n1198 ) );
XOR2_X2 _AES_ENC_U1314  ( .A(_AES_ENC_n986 ), .B(_AES_ENC_n985 ), .Z(_AES_ENC_sa02_next[4]) );
XOR2_X2 _AES_ENC_U1313  ( .A(_AES_ENC_n1198 ), .B(_AES_ENC_n987 ), .Z(_AES_ENC_n985 ) );
XOR2_X2 _AES_ENC_U1312  ( .A(_AES_ENC_n1204 ), .B(_AES_ENC_n1208 ), .Z(_AES_ENC_n986 ) );
XOR2_X2 _AES_ENC_U1311  ( .A(_AES_ENC_w2[28] ), .B(_AES_ENC_sa13_sub[4] ),.Z(_AES_ENC_n987 ) );
XOR2_X2 _AES_ENC_U1310  ( .A(_AES_ENC_sa02_sub[2] ), .B(_AES_ENC_sa13_sub[2] ), .Z(_AES_ENC_n1209 ) );
XOR2_X2 _AES_ENC_U1309  ( .A(_AES_ENC_sa20_sub[3] ), .B(_AES_ENC_sa31_sub[3] ), .Z(_AES_ENC_n1199 ) );
XOR2_X2 _AES_ENC_U1308  ( .A(_AES_ENC_n989 ), .B(_AES_ENC_n988 ), .Z(_AES_ENC_sa02_next[3]) );
XOR2_X2 _AES_ENC_U1307  ( .A(_AES_ENC_n1199 ), .B(_AES_ENC_n990 ), .Z(_AES_ENC_n988 ) );
XOR2_X2 _AES_ENC_U1306  ( .A(_AES_ENC_n1204 ), .B(_AES_ENC_n1209 ), .Z(_AES_ENC_n989 ) );
XOR2_X2 _AES_ENC_U1305  ( .A(_AES_ENC_w2[27] ), .B(_AES_ENC_sa13_sub[3] ),.Z(_AES_ENC_n990 ) );
XOR2_X2 _AES_ENC_U1304  ( .A(_AES_ENC_sa02_sub[1] ), .B(_AES_ENC_sa13_sub[1] ), .Z(_AES_ENC_n1210 ) );
XOR2_X2 _AES_ENC_U1303  ( .A(_AES_ENC_sa20_sub[2] ), .B(_AES_ENC_sa31_sub[2] ), .Z(_AES_ENC_n1200 ) );
XOR2_X2 _AES_ENC_U1302  ( .A(_AES_ENC_n992 ), .B(_AES_ENC_n991 ), .Z(_AES_ENC_sa02_next[2]) );
XOR2_X2 _AES_ENC_U1301  ( .A(_AES_ENC_n1210 ), .B(_AES_ENC_n1200 ), .Z(_AES_ENC_n991 ) );
XOR2_X2 _AES_ENC_U1300  ( .A(_AES_ENC_w2[26] ), .B(_AES_ENC_sa13_sub[2] ),.Z(_AES_ENC_n992 ) );
XOR2_X2 _AES_ENC_U1299  ( .A(_AES_ENC_sa02_sub[0] ), .B(_AES_ENC_sa13_sub[0] ), .Z(_AES_ENC_n1211 ) );
XOR2_X2 _AES_ENC_U1298  ( .A(_AES_ENC_sa20_sub[1] ), .B(_AES_ENC_sa31_sub[1] ), .Z(_AES_ENC_n1201 ) );
XOR2_X2 _AES_ENC_U1297  ( .A(_AES_ENC_n994 ), .B(_AES_ENC_n993 ), .Z(_AES_ENC_sa02_next[1]) );
XOR2_X2 _AES_ENC_U1296  ( .A(_AES_ENC_n1201 ), .B(_AES_ENC_n995 ), .Z(_AES_ENC_n993 ) );
XOR2_X2 _AES_ENC_U1295  ( .A(_AES_ENC_n1204 ), .B(_AES_ENC_n1211 ), .Z(_AES_ENC_n994 ) );
XOR2_X2 _AES_ENC_U1294  ( .A(_AES_ENC_w2[25] ), .B(_AES_ENC_sa13_sub[1] ),.Z(_AES_ENC_n995 ) );
XOR2_X2 _AES_ENC_U1293  ( .A(_AES_ENC_sa20_sub[0] ), .B(_AES_ENC_sa31_sub[0] ), .Z(_AES_ENC_n1202 ) );
XOR2_X2 _AES_ENC_U1292  ( .A(_AES_ENC_n997 ), .B(_AES_ENC_n996 ), .Z(_AES_ENC_sa02_next[0]) );
XOR2_X2 _AES_ENC_U1291  ( .A(_AES_ENC_n1204 ), .B(_AES_ENC_n1202 ), .Z(_AES_ENC_n996 ) );
XOR2_X2 _AES_ENC_U1290  ( .A(_AES_ENC_w2[24] ), .B(_AES_ENC_sa13_sub[0] ),.Z(_AES_ENC_n997 ) );
XOR2_X2 _AES_ENC_U1289  ( .A(_AES_ENC_n999 ), .B(_AES_ENC_n998 ), .Z(_AES_ENC_sa12_next[7]) );
XOR2_X2 _AES_ENC_U1288  ( .A(_AES_ENC_n1203 ), .B(_AES_ENC_n1000 ), .Z(_AES_ENC_n998 ) );
XOR2_X2 _AES_ENC_U1287  ( .A(_AES_ENC_sa13_sub[6] ), .B(_AES_ENC_sa20_sub[6] ), .Z(_AES_ENC_n999 ) );
XOR2_X2 _AES_ENC_U1286  ( .A(_AES_ENC_w2[23] ), .B(_AES_ENC_sa02_sub[7] ),.Z(_AES_ENC_n1000 ) );
XOR2_X2 _AES_ENC_U1285  ( .A(_AES_ENC_n1002 ), .B(_AES_ENC_n1001 ), .Z(_AES_ENC_sa12_next[6]) );
XOR2_X2 _AES_ENC_U1284  ( .A(_AES_ENC_n1196 ), .B(_AES_ENC_n1003 ), .Z(_AES_ENC_n1001 ) );
XOR2_X2 _AES_ENC_U1283  ( .A(_AES_ENC_sa13_sub[5] ), .B(_AES_ENC_sa20_sub[5] ), .Z(_AES_ENC_n1002 ) );
XOR2_X2 _AES_ENC_U1282  ( .A(_AES_ENC_w2[22] ), .B(_AES_ENC_sa02_sub[6] ),.Z(_AES_ENC_n1003 ) );
XOR2_X2 _AES_ENC_U1281  ( .A(_AES_ENC_n1005 ), .B(_AES_ENC_n1004 ), .Z(_AES_ENC_sa12_next[5]) );
XOR2_X2 _AES_ENC_U1280  ( .A(_AES_ENC_n1197 ), .B(_AES_ENC_n1006 ), .Z(_AES_ENC_n1004 ) );
XOR2_X2 _AES_ENC_U1279  ( .A(_AES_ENC_sa13_sub[4] ), .B(_AES_ENC_sa20_sub[4] ), .Z(_AES_ENC_n1005 ) );
XOR2_X2 _AES_ENC_U1278  ( .A(_AES_ENC_w2[21] ), .B(_AES_ENC_sa02_sub[5] ),.Z(_AES_ENC_n1006 ) );
XOR2_X2 _AES_ENC_U1277  ( .A(_AES_ENC_sa13_sub[7] ), .B(_AES_ENC_sa20_sub[7] ), .Z(_AES_ENC_n1195 ) );
XOR2_X2 _AES_ENC_U1276  ( .A(_AES_ENC_n1008 ), .B(_AES_ENC_n1007 ), .Z(_AES_ENC_sa12_next[4]) );
XOR2_X2 _AES_ENC_U1275  ( .A(_AES_ENC_n1010 ), .B(_AES_ENC_n1009 ), .Z(_AES_ENC_n1007 ) );
XOR2_X2 _AES_ENC_U1274  ( .A(_AES_ENC_n1195 ), .B(_AES_ENC_n1198 ), .Z(_AES_ENC_n1008 ) );
XOR2_X2 _AES_ENC_U1273  ( .A(_AES_ENC_sa13_sub[3] ), .B(_AES_ENC_sa20_sub[3] ), .Z(_AES_ENC_n1009 ) );
XOR2_X2 _AES_ENC_U1272  ( .A(_AES_ENC_w2[20] ), .B(_AES_ENC_sa02_sub[4] ),.Z(_AES_ENC_n1010 ) );
XOR2_X2 _AES_ENC_U1271  ( .A(_AES_ENC_n1012 ), .B(_AES_ENC_n1011 ), .Z(_AES_ENC_sa12_next[3]) );
XOR2_X2 _AES_ENC_U1270  ( .A(_AES_ENC_n1014 ), .B(_AES_ENC_n1013 ), .Z(_AES_ENC_n1011 ) );
XOR2_X2 _AES_ENC_U1269  ( .A(_AES_ENC_n1195 ), .B(_AES_ENC_n1199 ), .Z(_AES_ENC_n1012 ) );
XOR2_X2 _AES_ENC_U1268  ( .A(_AES_ENC_sa13_sub[2] ), .B(_AES_ENC_sa20_sub[2] ), .Z(_AES_ENC_n1013 ) );
XOR2_X2 _AES_ENC_U1267  ( .A(_AES_ENC_w2[19] ), .B(_AES_ENC_sa02_sub[3] ),.Z(_AES_ENC_n1014 ) );
XOR2_X2 _AES_ENC_U1266  ( .A(_AES_ENC_n1016 ), .B(_AES_ENC_n1015 ), .Z(_AES_ENC_sa12_next[2]) );
XOR2_X2 _AES_ENC_U1265  ( .A(_AES_ENC_n1200 ), .B(_AES_ENC_n1017 ), .Z(_AES_ENC_n1015 ) );
XOR2_X2 _AES_ENC_U1264  ( .A(_AES_ENC_sa13_sub[1] ), .B(_AES_ENC_sa20_sub[1] ), .Z(_AES_ENC_n1016 ) );
XOR2_X2 _AES_ENC_U1263  ( .A(_AES_ENC_w2[18] ), .B(_AES_ENC_sa02_sub[2] ),.Z(_AES_ENC_n1017 ) );
XOR2_X2 _AES_ENC_U1262  ( .A(_AES_ENC_n1019 ), .B(_AES_ENC_n1018 ), .Z(_AES_ENC_sa12_next[1]) );
XOR2_X2 _AES_ENC_U1261  ( .A(_AES_ENC_n1021 ), .B(_AES_ENC_n1020 ), .Z(_AES_ENC_n1018 ) );
XOR2_X2 _AES_ENC_U1260  ( .A(_AES_ENC_n1195 ), .B(_AES_ENC_n1201 ), .Z(_AES_ENC_n1019 ) );
XOR2_X2 _AES_ENC_U1259  ( .A(_AES_ENC_sa13_sub[0] ), .B(_AES_ENC_sa20_sub[0] ), .Z(_AES_ENC_n1020 ) );
XOR2_X2 _AES_ENC_U1258  ( .A(_AES_ENC_w2[17] ), .B(_AES_ENC_sa02_sub[1] ),.Z(_AES_ENC_n1021 ) );
XOR2_X2 _AES_ENC_U1257  ( .A(_AES_ENC_n1023 ), .B(_AES_ENC_n1022 ), .Z(_AES_ENC_sa12_next[0]) );
XOR2_X2 _AES_ENC_U1256  ( .A(_AES_ENC_n1195 ), .B(_AES_ENC_n1202 ), .Z(_AES_ENC_n1022 ) );
XOR2_X2 _AES_ENC_U1255  ( .A(_AES_ENC_w2[16] ), .B(_AES_ENC_sa02_sub[0] ),.Z(_AES_ENC_n1023 ) );
XOR2_X2 _AES_ENC_U1254  ( .A(_AES_ENC_n1025 ), .B(_AES_ENC_n1024 ), .Z(_AES_ENC_sa22_next[7]) );
XOR2_X2 _AES_ENC_U1253  ( .A(_AES_ENC_n1204 ), .B(_AES_ENC_n1196 ), .Z(_AES_ENC_n1024 ) );
XOR2_X2 _AES_ENC_U1252  ( .A(_AES_ENC_w2[15] ), .B(_AES_ENC_sa31_sub[7] ),.Z(_AES_ENC_n1025 ) );
XOR2_X2 _AES_ENC_U1251  ( .A(_AES_ENC_n1027 ), .B(_AES_ENC_n1026 ), .Z(_AES_ENC_sa22_next[6]) );
XOR2_X2 _AES_ENC_U1250  ( .A(_AES_ENC_n1205 ), .B(_AES_ENC_n1197 ), .Z(_AES_ENC_n1026 ) );
XOR2_X2 _AES_ENC_U1249  ( .A(_AES_ENC_w2[14] ), .B(_AES_ENC_sa31_sub[6] ),.Z(_AES_ENC_n1027 ) );
XOR2_X2 _AES_ENC_U1248  ( .A(_AES_ENC_n1029 ), .B(_AES_ENC_n1028 ), .Z(_AES_ENC_sa22_next[5]) );
XOR2_X2 _AES_ENC_U1247  ( .A(_AES_ENC_n1206 ), .B(_AES_ENC_n1198 ), .Z(_AES_ENC_n1028 ) );
XOR2_X2 _AES_ENC_U1246  ( .A(_AES_ENC_w2[13] ), .B(_AES_ENC_sa31_sub[5] ),.Z(_AES_ENC_n1029 ) );
XOR2_X2 _AES_ENC_U1245  ( .A(_AES_ENC_n1031 ), .B(_AES_ENC_n1030 ), .Z(_AES_ENC_sa22_next[4]) );
XOR2_X2 _AES_ENC_U1244  ( .A(_AES_ENC_n1199 ), .B(_AES_ENC_n1032 ), .Z(_AES_ENC_n1030 ) );
XOR2_X2 _AES_ENC_U1243  ( .A(_AES_ENC_n1203 ), .B(_AES_ENC_n1207 ), .Z(_AES_ENC_n1031 ) );
XOR2_X2 _AES_ENC_U1242  ( .A(_AES_ENC_w2[12] ), .B(_AES_ENC_sa31_sub[4] ),.Z(_AES_ENC_n1032 ) );
XOR2_X2 _AES_ENC_U1241  ( .A(_AES_ENC_n1034 ), .B(_AES_ENC_n1033 ), .Z(_AES_ENC_sa22_next[3]) );
XOR2_X2 _AES_ENC_U1240  ( .A(_AES_ENC_n1200 ), .B(_AES_ENC_n1035 ), .Z(_AES_ENC_n1033 ) );
XOR2_X2 _AES_ENC_U1239  ( .A(_AES_ENC_n1203 ), .B(_AES_ENC_n1208 ), .Z(_AES_ENC_n1034 ) );
XOR2_X2 _AES_ENC_U1238  ( .A(_AES_ENC_w2[11] ), .B(_AES_ENC_sa31_sub[3] ),.Z(_AES_ENC_n1035 ) );
XOR2_X2 _AES_ENC_U1237  ( .A(_AES_ENC_n1037 ), .B(_AES_ENC_n1036 ), .Z(_AES_ENC_sa22_next[2]) );
XOR2_X2 _AES_ENC_U1236  ( .A(_AES_ENC_n1209 ), .B(_AES_ENC_n1201 ), .Z(_AES_ENC_n1036 ) );
XOR2_X2 _AES_ENC_U1235  ( .A(_AES_ENC_w2[10] ), .B(_AES_ENC_sa31_sub[2] ),.Z(_AES_ENC_n1037 ) );
XOR2_X2 _AES_ENC_U1234  ( .A(_AES_ENC_n1039 ), .B(_AES_ENC_n1038 ), .Z(_AES_ENC_sa22_next[1]) );
XOR2_X2 _AES_ENC_U1233  ( .A(_AES_ENC_n1202 ), .B(_AES_ENC_n1040 ), .Z(_AES_ENC_n1038 ) );
XOR2_X2 _AES_ENC_U1232  ( .A(_AES_ENC_n1203 ), .B(_AES_ENC_n1210 ), .Z(_AES_ENC_n1039 ) );
XOR2_X2 _AES_ENC_U1231  ( .A(_AES_ENC_w2[9] ), .B(_AES_ENC_sa31_sub[1] ),.Z(_AES_ENC_n1040 ) );
XOR2_X2 _AES_ENC_U1230  ( .A(_AES_ENC_n1042 ), .B(_AES_ENC_n1041 ), .Z(_AES_ENC_sa22_next[0]) );
XOR2_X2 _AES_ENC_U1229  ( .A(_AES_ENC_n1203 ), .B(_AES_ENC_n1211 ), .Z(_AES_ENC_n1041 ) );
XOR2_X2 _AES_ENC_U1228  ( .A(_AES_ENC_w2[8] ), .B(_AES_ENC_sa31_sub[0] ),.Z(_AES_ENC_n1042 ) );
XOR2_X2 _AES_ENC_U1227  ( .A(_AES_ENC_n1044 ), .B(_AES_ENC_n1043 ), .Z(_AES_ENC_sa32_next[7]) );
XOR2_X2 _AES_ENC_U1226  ( .A(_AES_ENC_n1204 ), .B(_AES_ENC_n1045 ), .Z(_AES_ENC_n1043 ) );
XOR2_X2 _AES_ENC_U1225  ( .A(_AES_ENC_sa20_sub[7] ), .B(_AES_ENC_sa31_sub[6] ), .Z(_AES_ENC_n1044 ) );
XOR2_X2 _AES_ENC_U1224  ( .A(_AES_ENC_w2[7] ), .B(_AES_ENC_sa02_sub[6] ),.Z(_AES_ENC_n1045 ) );
XOR2_X2 _AES_ENC_U1223  ( .A(_AES_ENC_n1047 ), .B(_AES_ENC_n1046 ), .Z(_AES_ENC_sa32_next[6]) );
XOR2_X2 _AES_ENC_U1222  ( .A(_AES_ENC_n1205 ), .B(_AES_ENC_n1048 ), .Z(_AES_ENC_n1046 ) );
XOR2_X2 _AES_ENC_U1221  ( .A(_AES_ENC_sa20_sub[6] ), .B(_AES_ENC_sa31_sub[5] ), .Z(_AES_ENC_n1047 ) );
XOR2_X2 _AES_ENC_U1220  ( .A(_AES_ENC_w2[6] ), .B(_AES_ENC_sa02_sub[5] ),.Z(_AES_ENC_n1048 ) );
XOR2_X2 _AES_ENC_U1219  ( .A(_AES_ENC_n1050 ), .B(_AES_ENC_n1049 ), .Z(_AES_ENC_sa32_next[5]) );
XOR2_X2 _AES_ENC_U1218  ( .A(_AES_ENC_n1206 ), .B(_AES_ENC_n1051 ), .Z(_AES_ENC_n1049 ) );
XOR2_X2 _AES_ENC_U1217  ( .A(_AES_ENC_sa20_sub[5] ), .B(_AES_ENC_sa31_sub[4] ), .Z(_AES_ENC_n1050 ) );
XOR2_X2 _AES_ENC_U1216  ( .A(_AES_ENC_w2[5] ), .B(_AES_ENC_sa02_sub[4] ),.Z(_AES_ENC_n1051 ) );
XOR2_X2 _AES_ENC_U1215  ( .A(_AES_ENC_sa02_sub[7] ), .B(_AES_ENC_sa31_sub[7] ), .Z(_AES_ENC_n1212 ) );
XOR2_X2 _AES_ENC_U1214  ( .A(_AES_ENC_n1053 ), .B(_AES_ENC_n1052 ), .Z(_AES_ENC_sa32_next[4]) );
XOR2_X2 _AES_ENC_U1213  ( .A(_AES_ENC_n1055 ), .B(_AES_ENC_n1054 ), .Z(_AES_ENC_n1052 ) );
XOR2_X2 _AES_ENC_U1212  ( .A(_AES_ENC_n1212 ), .B(_AES_ENC_n1207 ), .Z(_AES_ENC_n1053 ) );
XOR2_X2 _AES_ENC_U1211  ( .A(_AES_ENC_sa20_sub[4] ), .B(_AES_ENC_sa31_sub[3] ), .Z(_AES_ENC_n1054 ) );
XOR2_X2 _AES_ENC_U1210  ( .A(_AES_ENC_w2[4] ), .B(_AES_ENC_sa02_sub[3] ),.Z(_AES_ENC_n1055 ) );
XOR2_X2 _AES_ENC_U1209  ( .A(_AES_ENC_n1057 ), .B(_AES_ENC_n1056 ), .Z(_AES_ENC_sa32_next[3]) );
XOR2_X2 _AES_ENC_U1208  ( .A(_AES_ENC_n1059 ), .B(_AES_ENC_n1058 ), .Z(_AES_ENC_n1056 ) );
XOR2_X2 _AES_ENC_U1207  ( .A(_AES_ENC_n1212 ), .B(_AES_ENC_n1208 ), .Z(_AES_ENC_n1057 ) );
XOR2_X2 _AES_ENC_U1206  ( .A(_AES_ENC_sa20_sub[3] ), .B(_AES_ENC_sa31_sub[2] ), .Z(_AES_ENC_n1058 ) );
XOR2_X2 _AES_ENC_U1205  ( .A(_AES_ENC_w2[3] ), .B(_AES_ENC_sa02_sub[2] ),.Z(_AES_ENC_n1059 ) );
XOR2_X2 _AES_ENC_U1204  ( .A(_AES_ENC_n1061 ), .B(_AES_ENC_n1060 ), .Z(_AES_ENC_sa32_next[2]) );
XOR2_X2 _AES_ENC_U1203  ( .A(_AES_ENC_n1209 ), .B(_AES_ENC_n1062 ), .Z(_AES_ENC_n1060 ) );
XOR2_X2 _AES_ENC_U1202  ( .A(_AES_ENC_sa20_sub[2] ), .B(_AES_ENC_sa31_sub[1] ), .Z(_AES_ENC_n1061 ) );
XOR2_X2 _AES_ENC_U1201  ( .A(_AES_ENC_w2[2] ), .B(_AES_ENC_sa02_sub[1] ),.Z(_AES_ENC_n1062 ) );
XOR2_X2 _AES_ENC_U1200  ( .A(_AES_ENC_n1064 ), .B(_AES_ENC_n1063 ), .Z(_AES_ENC_sa32_next[1]) );
XOR2_X2 _AES_ENC_U1199  ( .A(_AES_ENC_n1066 ), .B(_AES_ENC_n1065 ), .Z(_AES_ENC_n1063 ) );
XOR2_X2 _AES_ENC_U1198  ( .A(_AES_ENC_n1212 ), .B(_AES_ENC_n1210 ), .Z(_AES_ENC_n1064 ) );
XOR2_X2 _AES_ENC_U1197  ( .A(_AES_ENC_sa20_sub[1] ), .B(_AES_ENC_sa31_sub[0] ), .Z(_AES_ENC_n1065 ) );
XOR2_X2 _AES_ENC_U1196  ( .A(_AES_ENC_w2[1] ), .B(_AES_ENC_sa02_sub[0] ),.Z(_AES_ENC_n1066 ) );
XOR2_X2 _AES_ENC_U1195  ( .A(_AES_ENC_n1068 ), .B(_AES_ENC_n1067 ), .Z(_AES_ENC_sa32_next[0]) );
XOR2_X2 _AES_ENC_U1194  ( .A(_AES_ENC_n1212 ), .B(_AES_ENC_n1211 ), .Z(_AES_ENC_n1067 ) );
XOR2_X2 _AES_ENC_U1193  ( .A(_AES_ENC_w2[0] ), .B(_AES_ENC_sa20_sub[0] ),.Z(_AES_ENC_n1068 ) );
XOR2_X2 _AES_ENC_U1192  ( .A(_AES_ENC_sa21_sub[7] ), .B(_AES_ENC_sa32_sub[7] ), .Z(_AES_ENC_n1221 ) );
XOR2_X2 _AES_ENC_U1191  ( .A(_AES_ENC_sa03_sub[6] ), .B(_AES_ENC_sa10_sub[6] ), .Z(_AES_ENC_n1223 ) );
XOR2_X2 _AES_ENC_U1190  ( .A(_AES_ENC_n1070 ), .B(_AES_ENC_n1069 ), .Z(_AES_ENC_sa03_next[7]) );
XOR2_X2 _AES_ENC_U1189  ( .A(_AES_ENC_n1221 ), .B(_AES_ENC_n1223 ), .Z(_AES_ENC_n1069 ) );
XOR2_X2 _AES_ENC_U1188  ( .A(_AES_ENC_w3[31] ), .B(_AES_ENC_sa10_sub[7] ),.Z(_AES_ENC_n1070 ) );
XOR2_X2 _AES_ENC_U1187  ( .A(_AES_ENC_sa03_sub[5] ), .B(_AES_ENC_sa10_sub[5] ), .Z(_AES_ENC_n1224 ) );
XOR2_X2 _AES_ENC_U1186  ( .A(_AES_ENC_sa21_sub[6] ), .B(_AES_ENC_sa32_sub[6] ), .Z(_AES_ENC_n1214 ) );
XOR2_X2 _AES_ENC_U1185  ( .A(_AES_ENC_n1072 ), .B(_AES_ENC_n1071 ), .Z(_AES_ENC_sa03_next[6]) );
XOR2_X2 _AES_ENC_U1184  ( .A(_AES_ENC_n1224 ), .B(_AES_ENC_n1214 ), .Z(_AES_ENC_n1071 ) );
XOR2_X2 _AES_ENC_U1183  ( .A(_AES_ENC_w3[30] ), .B(_AES_ENC_sa10_sub[6] ),.Z(_AES_ENC_n1072 ) );
XOR2_X2 _AES_ENC_U1182  ( .A(_AES_ENC_sa03_sub[4] ), .B(_AES_ENC_sa10_sub[4] ), .Z(_AES_ENC_n1225 ) );
XOR2_X2 _AES_ENC_U1181  ( .A(_AES_ENC_sa21_sub[5] ), .B(_AES_ENC_sa32_sub[5] ), .Z(_AES_ENC_n1215 ) );
XOR2_X2 _AES_ENC_U1180  ( .A(_AES_ENC_n1074 ), .B(_AES_ENC_n1073 ), .Z(_AES_ENC_sa03_next[5]) );
XOR2_X2 _AES_ENC_U1179  ( .A(_AES_ENC_n1225 ), .B(_AES_ENC_n1215 ), .Z(_AES_ENC_n1073 ) );
XOR2_X2 _AES_ENC_U1178  ( .A(_AES_ENC_w3[29] ), .B(_AES_ENC_sa10_sub[5] ),.Z(_AES_ENC_n1074 ) );
XOR2_X2 _AES_ENC_U1177  ( .A(_AES_ENC_sa03_sub[7] ), .B(_AES_ENC_sa10_sub[7] ), .Z(_AES_ENC_n1222 ) );
XOR2_X2 _AES_ENC_U1176  ( .A(_AES_ENC_sa03_sub[3] ), .B(_AES_ENC_sa10_sub[3] ), .Z(_AES_ENC_n1226 ) );
XOR2_X2 _AES_ENC_U1175  ( .A(_AES_ENC_sa21_sub[4] ), .B(_AES_ENC_sa32_sub[4] ), .Z(_AES_ENC_n1216 ) );
XOR2_X2 _AES_ENC_U1174  ( .A(_AES_ENC_n1076 ), .B(_AES_ENC_n1075 ), .Z(_AES_ENC_sa03_next[4]) );
XOR2_X2 _AES_ENC_U1173  ( .A(_AES_ENC_n1216 ), .B(_AES_ENC_n1077 ), .Z(_AES_ENC_n1075 ) );
XOR2_X2 _AES_ENC_U1172  ( .A(_AES_ENC_n1222 ), .B(_AES_ENC_n1226 ), .Z(_AES_ENC_n1076 ) );
XOR2_X2 _AES_ENC_U1171  ( .A(_AES_ENC_w3[28] ), .B(_AES_ENC_sa10_sub[4] ),.Z(_AES_ENC_n1077 ) );
XOR2_X2 _AES_ENC_U1170  ( .A(_AES_ENC_sa03_sub[2] ), .B(_AES_ENC_sa10_sub[2] ), .Z(_AES_ENC_n1227 ) );
XOR2_X2 _AES_ENC_U1169  ( .A(_AES_ENC_sa21_sub[3] ), .B(_AES_ENC_sa32_sub[3] ), .Z(_AES_ENC_n1217 ) );
XOR2_X2 _AES_ENC_U1168  ( .A(_AES_ENC_n1079 ), .B(_AES_ENC_n1078 ), .Z(_AES_ENC_sa03_next[3]) );
XOR2_X2 _AES_ENC_U1167  ( .A(_AES_ENC_n1217 ), .B(_AES_ENC_n1080 ), .Z(_AES_ENC_n1078 ) );
XOR2_X2 _AES_ENC_U1166  ( .A(_AES_ENC_n1222 ), .B(_AES_ENC_n1227 ), .Z(_AES_ENC_n1079 ) );
XOR2_X2 _AES_ENC_U1165  ( .A(_AES_ENC_w3[27] ), .B(_AES_ENC_sa10_sub[3] ),.Z(_AES_ENC_n1080 ) );
XOR2_X2 _AES_ENC_U1164  ( .A(_AES_ENC_sa03_sub[1] ), .B(_AES_ENC_sa10_sub[1] ), .Z(_AES_ENC_n1228 ) );
XOR2_X2 _AES_ENC_U1163  ( .A(_AES_ENC_sa21_sub[2] ), .B(_AES_ENC_sa32_sub[2] ), .Z(_AES_ENC_n1218 ) );
XOR2_X2 _AES_ENC_U1162  ( .A(_AES_ENC_n1082 ), .B(_AES_ENC_n1081 ), .Z(_AES_ENC_sa03_next[2]) );
XOR2_X2 _AES_ENC_U1161  ( .A(_AES_ENC_n1228 ), .B(_AES_ENC_n1218 ), .Z(_AES_ENC_n1081 ) );
XOR2_X2 _AES_ENC_U1160  ( .A(_AES_ENC_w3[26] ), .B(_AES_ENC_sa10_sub[2] ),.Z(_AES_ENC_n1082 ) );
XOR2_X2 _AES_ENC_U1159  ( .A(_AES_ENC_sa03_sub[0] ), .B(_AES_ENC_sa10_sub[0] ), .Z(_AES_ENC_n1229 ) );
XOR2_X2 _AES_ENC_U1158  ( .A(_AES_ENC_sa21_sub[1] ), .B(_AES_ENC_sa32_sub[1] ), .Z(_AES_ENC_n1219 ) );
XOR2_X2 _AES_ENC_U1157  ( .A(_AES_ENC_n1084 ), .B(_AES_ENC_n1083 ), .Z(_AES_ENC_sa03_next[1]) );
XOR2_X2 _AES_ENC_U1156  ( .A(_AES_ENC_n1219 ), .B(_AES_ENC_n1085 ), .Z(_AES_ENC_n1083 ) );
XOR2_X2 _AES_ENC_U1155  ( .A(_AES_ENC_n1222 ), .B(_AES_ENC_n1229 ), .Z(_AES_ENC_n1084 ) );
XOR2_X2 _AES_ENC_U1154  ( .A(_AES_ENC_w3[25] ), .B(_AES_ENC_sa10_sub[1] ),.Z(_AES_ENC_n1085 ) );
XOR2_X2 _AES_ENC_U1153  ( .A(_AES_ENC_sa21_sub[0] ), .B(_AES_ENC_sa32_sub[0] ), .Z(_AES_ENC_n1220 ) );
XOR2_X2 _AES_ENC_U1152  ( .A(_AES_ENC_n1087 ), .B(_AES_ENC_n1086 ), .Z(_AES_ENC_sa03_next[0]) );
XOR2_X2 _AES_ENC_U1151  ( .A(_AES_ENC_n1222 ), .B(_AES_ENC_n1220 ), .Z(_AES_ENC_n1086 ) );
XOR2_X2 _AES_ENC_U1150  ( .A(_AES_ENC_w3[24] ), .B(_AES_ENC_sa10_sub[0] ),.Z(_AES_ENC_n1087 ) );
XOR2_X2 _AES_ENC_U1149  ( .A(_AES_ENC_n1089 ), .B(_AES_ENC_n1088 ), .Z(_AES_ENC_sa13_next[7]) );
XOR2_X2 _AES_ENC_U1148  ( .A(_AES_ENC_n1221 ), .B(_AES_ENC_n1090 ), .Z(_AES_ENC_n1088 ) );
XOR2_X2 _AES_ENC_U1147  ( .A(_AES_ENC_sa10_sub[6] ), .B(_AES_ENC_sa21_sub[6] ), .Z(_AES_ENC_n1089 ) );
XOR2_X2 _AES_ENC_U1146  ( .A(_AES_ENC_w3[23] ), .B(_AES_ENC_sa03_sub[7] ),.Z(_AES_ENC_n1090 ) );
XOR2_X2 _AES_ENC_U1145  ( .A(_AES_ENC_n1092 ), .B(_AES_ENC_n1091 ), .Z(_AES_ENC_sa13_next[6]) );
XOR2_X2 _AES_ENC_U1144  ( .A(_AES_ENC_n1214 ), .B(_AES_ENC_n1093 ), .Z(_AES_ENC_n1091 ) );
XOR2_X2 _AES_ENC_U1143  ( .A(_AES_ENC_sa10_sub[5] ), .B(_AES_ENC_sa21_sub[5] ), .Z(_AES_ENC_n1092 ) );
XOR2_X2 _AES_ENC_U1142  ( .A(_AES_ENC_w3[22] ), .B(_AES_ENC_sa03_sub[6] ),.Z(_AES_ENC_n1093 ) );
XOR2_X2 _AES_ENC_U1141  ( .A(_AES_ENC_n1095 ), .B(_AES_ENC_n1094 ), .Z(_AES_ENC_sa13_next[5]) );
XOR2_X2 _AES_ENC_U1140  ( .A(_AES_ENC_n1215 ), .B(_AES_ENC_n1096 ), .Z(_AES_ENC_n1094 ) );
XOR2_X2 _AES_ENC_U1139  ( .A(_AES_ENC_sa10_sub[4] ), .B(_AES_ENC_sa21_sub[4] ), .Z(_AES_ENC_n1095 ) );
XOR2_X2 _AES_ENC_U1138  ( .A(_AES_ENC_w3[21] ), .B(_AES_ENC_sa03_sub[5] ),.Z(_AES_ENC_n1096 ) );
XOR2_X2 _AES_ENC_U1137  ( .A(_AES_ENC_sa10_sub[7] ), .B(_AES_ENC_sa21_sub[7] ), .Z(_AES_ENC_n1213 ) );
XOR2_X2 _AES_ENC_U1136  ( .A(_AES_ENC_n1098 ), .B(_AES_ENC_n1097 ), .Z(_AES_ENC_sa13_next[4]) );
XOR2_X2 _AES_ENC_U1135  ( .A(_AES_ENC_n1100 ), .B(_AES_ENC_n1099 ), .Z(_AES_ENC_n1097 ) );
XOR2_X2 _AES_ENC_U1134  ( .A(_AES_ENC_n1213 ), .B(_AES_ENC_n1216 ), .Z(_AES_ENC_n1098 ) );
XOR2_X2 _AES_ENC_U1133  ( .A(_AES_ENC_sa10_sub[3] ), .B(_AES_ENC_sa21_sub[3] ), .Z(_AES_ENC_n1099 ) );
XOR2_X2 _AES_ENC_U1132  ( .A(_AES_ENC_w3[20] ), .B(_AES_ENC_sa03_sub[4] ),.Z(_AES_ENC_n1100 ) );
XOR2_X2 _AES_ENC_U1131  ( .A(_AES_ENC_n1102 ), .B(_AES_ENC_n1101 ), .Z(_AES_ENC_sa13_next[3]) );
XOR2_X2 _AES_ENC_U1130  ( .A(_AES_ENC_n1104 ), .B(_AES_ENC_n1103 ), .Z(_AES_ENC_n1101 ) );
XOR2_X2 _AES_ENC_U1129  ( .A(_AES_ENC_n1213 ), .B(_AES_ENC_n1217 ), .Z(_AES_ENC_n1102 ) );
XOR2_X2 _AES_ENC_U1128  ( .A(_AES_ENC_sa10_sub[2] ), .B(_AES_ENC_sa21_sub[2] ), .Z(_AES_ENC_n1103 ) );
XOR2_X2 _AES_ENC_U1127  ( .A(_AES_ENC_w3[19] ), .B(_AES_ENC_sa03_sub[3] ),.Z(_AES_ENC_n1104 ) );
XOR2_X2 _AES_ENC_U1126  ( .A(_AES_ENC_n1106 ), .B(_AES_ENC_n1105 ), .Z(_AES_ENC_sa13_next[2]) );
XOR2_X2 _AES_ENC_U1125  ( .A(_AES_ENC_n1218 ), .B(_AES_ENC_n1107 ), .Z(_AES_ENC_n1105 ) );
XOR2_X2 _AES_ENC_U1124  ( .A(_AES_ENC_sa10_sub[1] ), .B(_AES_ENC_sa21_sub[1] ), .Z(_AES_ENC_n1106 ) );
XOR2_X2 _AES_ENC_U1123  ( .A(_AES_ENC_w3[18] ), .B(_AES_ENC_sa03_sub[2] ),.Z(_AES_ENC_n1107 ) );
XOR2_X2 _AES_ENC_U1122  ( .A(_AES_ENC_n1109 ), .B(_AES_ENC_n1108 ), .Z(_AES_ENC_sa13_next[1]) );
XOR2_X2 _AES_ENC_U1121  ( .A(_AES_ENC_n1111 ), .B(_AES_ENC_n1110 ), .Z(_AES_ENC_n1108 ) );
XOR2_X2 _AES_ENC_U1120  ( .A(_AES_ENC_n1213 ), .B(_AES_ENC_n1219 ), .Z(_AES_ENC_n1109 ) );
XOR2_X2 _AES_ENC_U1119  ( .A(_AES_ENC_sa10_sub[0] ), .B(_AES_ENC_sa21_sub[0] ), .Z(_AES_ENC_n1110 ) );
XOR2_X2 _AES_ENC_U1118  ( .A(_AES_ENC_w3[17] ), .B(_AES_ENC_sa03_sub[1] ),.Z(_AES_ENC_n1111 ) );
XOR2_X2 _AES_ENC_U1117  ( .A(_AES_ENC_n1113 ), .B(_AES_ENC_n1112 ), .Z(_AES_ENC_sa13_next[0]) );
XOR2_X2 _AES_ENC_U1116  ( .A(_AES_ENC_n1213 ), .B(_AES_ENC_n1220 ), .Z(_AES_ENC_n1112 ) );
XOR2_X2 _AES_ENC_U1115  ( .A(_AES_ENC_w3[16] ), .B(_AES_ENC_sa03_sub[0] ),.Z(_AES_ENC_n1113 ) );
XOR2_X2 _AES_ENC_U1114  ( .A(_AES_ENC_n1115 ), .B(_AES_ENC_n1114 ), .Z(_AES_ENC_sa23_next[7]) );
XOR2_X2 _AES_ENC_U1113  ( .A(_AES_ENC_n1222 ), .B(_AES_ENC_n1214 ), .Z(_AES_ENC_n1114 ) );
XOR2_X2 _AES_ENC_U1112  ( .A(_AES_ENC_w3[15] ), .B(_AES_ENC_sa32_sub[7] ),.Z(_AES_ENC_n1115 ) );
XOR2_X2 _AES_ENC_U1111  ( .A(_AES_ENC_n1117 ), .B(_AES_ENC_n1116 ), .Z(_AES_ENC_sa23_next[6]) );
XOR2_X2 _AES_ENC_U1110  ( .A(_AES_ENC_n1223 ), .B(_AES_ENC_n1215 ), .Z(_AES_ENC_n1116 ) );
XOR2_X2 _AES_ENC_U1109  ( .A(_AES_ENC_w3[14] ), .B(_AES_ENC_sa32_sub[6] ),.Z(_AES_ENC_n1117 ) );
XOR2_X2 _AES_ENC_U1108  ( .A(_AES_ENC_n1119 ), .B(_AES_ENC_n1118 ), .Z(_AES_ENC_sa23_next[5]) );
XOR2_X2 _AES_ENC_U1107  ( .A(_AES_ENC_n1224 ), .B(_AES_ENC_n1216 ), .Z(_AES_ENC_n1118 ) );
XOR2_X2 _AES_ENC_U1106  ( .A(_AES_ENC_w3[13] ), .B(_AES_ENC_sa32_sub[5] ),.Z(_AES_ENC_n1119 ) );
XOR2_X2 _AES_ENC_U1105  ( .A(_AES_ENC_n1121 ), .B(_AES_ENC_n1120 ), .Z(_AES_ENC_sa23_next[4]) );
XOR2_X2 _AES_ENC_U1104  ( .A(_AES_ENC_n1217 ), .B(_AES_ENC_n1122 ), .Z(_AES_ENC_n1120 ) );
XOR2_X2 _AES_ENC_U1103  ( .A(_AES_ENC_n1221 ), .B(_AES_ENC_n1225 ), .Z(_AES_ENC_n1121 ) );
XOR2_X2 _AES_ENC_U1102  ( .A(_AES_ENC_w3[12] ), .B(_AES_ENC_sa32_sub[4] ),.Z(_AES_ENC_n1122 ) );
XOR2_X2 _AES_ENC_U1101  ( .A(_AES_ENC_n1124 ), .B(_AES_ENC_n1123 ), .Z(_AES_ENC_sa23_next[3]) );
XOR2_X2 _AES_ENC_U1100  ( .A(_AES_ENC_n1218 ), .B(_AES_ENC_n1125 ), .Z(_AES_ENC_n1123 ) );
XOR2_X2 _AES_ENC_U1099  ( .A(_AES_ENC_n1221 ), .B(_AES_ENC_n1226 ), .Z(_AES_ENC_n1124 ) );
XOR2_X2 _AES_ENC_U1098  ( .A(_AES_ENC_w3[11] ), .B(_AES_ENC_sa32_sub[3] ),.Z(_AES_ENC_n1125 ) );
XOR2_X2 _AES_ENC_U1097  ( .A(_AES_ENC_n1127 ), .B(_AES_ENC_n1126 ), .Z(_AES_ENC_sa23_next[2]) );
XOR2_X2 _AES_ENC_U1096  ( .A(_AES_ENC_n1227 ), .B(_AES_ENC_n1219 ), .Z(_AES_ENC_n1126 ) );
XOR2_X2 _AES_ENC_U1095  ( .A(_AES_ENC_w3[10] ), .B(_AES_ENC_sa32_sub[2] ),.Z(_AES_ENC_n1127 ) );
XOR2_X2 _AES_ENC_U1094  ( .A(_AES_ENC_n1129 ), .B(_AES_ENC_n1128 ), .Z(_AES_ENC_sa23_next[1]) );
XOR2_X2 _AES_ENC_U1093  ( .A(_AES_ENC_n1220 ), .B(_AES_ENC_n1130 ), .Z(_AES_ENC_n1128 ) );
XOR2_X2 _AES_ENC_U1092  ( .A(_AES_ENC_n1221 ), .B(_AES_ENC_n1228 ), .Z(_AES_ENC_n1129 ) );
XOR2_X2 _AES_ENC_U1091  ( .A(_AES_ENC_w3[9] ), .B(_AES_ENC_sa32_sub[1] ),.Z(_AES_ENC_n1130 ) );
XOR2_X2 _AES_ENC_U1090  ( .A(_AES_ENC_n1132 ), .B(_AES_ENC_n1131 ), .Z(_AES_ENC_sa23_next[0]) );
XOR2_X2 _AES_ENC_U1089  ( .A(_AES_ENC_n1221 ), .B(_AES_ENC_n1229 ), .Z(_AES_ENC_n1131 ) );
XOR2_X2 _AES_ENC_U1088  ( .A(_AES_ENC_w3[8] ), .B(_AES_ENC_sa32_sub[0] ),.Z(_AES_ENC_n1132 ) );
XOR2_X2 _AES_ENC_U1087  ( .A(_AES_ENC_n1134 ), .B(_AES_ENC_n1133 ), .Z(__AES_ENC_sa33_next[7]) );
XOR2_X2 _AES_ENC_U1086  ( .A(_AES_ENC_n1222 ), .B(_AES_ENC_n1135 ), .Z(_AES_ENC_n1133 ) );
XOR2_X2 _AES_ENC_U1085  ( .A(_AES_ENC_sa21_sub[7] ), .B(_AES_ENC_sa32_sub[6] ), .Z(_AES_ENC_n1134 ) );
XOR2_X2 _AES_ENC_U1084  ( .A(_AES_ENC_w3[7] ), .B(_AES_ENC_sa03_sub[6] ),.Z(_AES_ENC_n1135 ) );
XOR2_X2 _AES_ENC_U1083  ( .A(_AES_ENC_n1137 ), .B(_AES_ENC_n1136 ), .Z(__AES_ENC_sa33_next[6]) );
XOR2_X2 _AES_ENC_U1082  ( .A(_AES_ENC_n1223 ), .B(_AES_ENC_n1138 ), .Z(_AES_ENC_n1136 ) );
XOR2_X2 _AES_ENC_U1081  ( .A(_AES_ENC_sa21_sub[6] ), .B(_AES_ENC_sa32_sub[5] ), .Z(_AES_ENC_n1137 ) );
XOR2_X2 _AES_ENC_U1080  ( .A(_AES_ENC_w3[6] ), .B(_AES_ENC_sa03_sub[5] ),.Z(_AES_ENC_n1138 ) );
XOR2_X2 _AES_ENC_U1079  ( .A(_AES_ENC_n1140 ), .B(_AES_ENC_n1139 ), .Z(__AES_ENC_sa33_next[5]) );
XOR2_X2 _AES_ENC_U1078  ( .A(_AES_ENC_n1224 ), .B(_AES_ENC_n1141 ), .Z(_AES_ENC_n1139 ) );
XOR2_X2 _AES_ENC_U1077  ( .A(_AES_ENC_sa21_sub[5] ), .B(_AES_ENC_sa32_sub[4] ), .Z(_AES_ENC_n1140 ) );
XOR2_X2 _AES_ENC_U1076  ( .A(_AES_ENC_w3[5] ), .B(_AES_ENC_sa03_sub[4] ),.Z(_AES_ENC_n1141 ) );
XOR2_X2 _AES_ENC_U1075  ( .A(_AES_ENC_sa03_sub[7] ), .B(_AES_ENC_sa32_sub[7] ), .Z(_AES_ENC_n1230 ) );
XOR2_X2 _AES_ENC_U1074  ( .A(_AES_ENC_n1143 ), .B(_AES_ENC_n1142 ), .Z(__AES_ENC_sa33_next[4]) );
XOR2_X2 _AES_ENC_U1073  ( .A(_AES_ENC_n1145 ), .B(_AES_ENC_n1144 ), .Z(_AES_ENC_n1142 ) );
XOR2_X2 _AES_ENC_U1072  ( .A(_AES_ENC_n1230 ), .B(_AES_ENC_n1225 ), .Z(_AES_ENC_n1143 ) );
XOR2_X2 _AES_ENC_U1071  ( .A(_AES_ENC_sa21_sub[4] ), .B(_AES_ENC_sa32_sub[3] ), .Z(_AES_ENC_n1144 ) );
XOR2_X2 _AES_ENC_U1070  ( .A(_AES_ENC_w3[4] ), .B(_AES_ENC_sa03_sub[3] ),.Z(_AES_ENC_n1145 ) );
XOR2_X2 _AES_ENC_U1069  ( .A(_AES_ENC_n1147 ), .B(_AES_ENC_n1146 ), .Z(__AES_ENC_sa33_next[3]) );
XOR2_X2 _AES_ENC_U1068  ( .A(_AES_ENC_n1149 ), .B(_AES_ENC_n1148 ), .Z(_AES_ENC_n1146 ) );
XOR2_X2 _AES_ENC_U1067  ( .A(_AES_ENC_n1230 ), .B(_AES_ENC_n1226 ), .Z(_AES_ENC_n1147 ) );
XOR2_X2 _AES_ENC_U1066  ( .A(_AES_ENC_sa21_sub[3] ), .B(_AES_ENC_sa32_sub[2] ), .Z(_AES_ENC_n1148 ) );
XOR2_X2 _AES_ENC_U1065  ( .A(_AES_ENC_w3[3] ), .B(_AES_ENC_sa03_sub[2] ),.Z(_AES_ENC_n1149 ) );
XOR2_X2 _AES_ENC_U1064  ( .A(_AES_ENC_n1151 ), .B(_AES_ENC_n1150 ), .Z(__AES_ENC_sa33_next[2]) );
XOR2_X2 _AES_ENC_U1063  ( .A(_AES_ENC_n1227 ), .B(_AES_ENC_n1152 ), .Z(_AES_ENC_n1150 ) );
XOR2_X2 _AES_ENC_U1062  ( .A(_AES_ENC_sa21_sub[2] ), .B(_AES_ENC_sa32_sub[1] ), .Z(_AES_ENC_n1151 ) );
XOR2_X2 _AES_ENC_U1061  ( .A(_AES_ENC_w3[2] ), .B(_AES_ENC_sa03_sub[1] ),.Z(_AES_ENC_n1152 ) );
XOR2_X2 _AES_ENC_U1060  ( .A(_AES_ENC_n1154 ), .B(_AES_ENC_n1153 ), .Z(__AES_ENC_sa33_next[1]) );
XOR2_X2 _AES_ENC_U1059  ( .A(_AES_ENC_n1156 ), .B(_AES_ENC_n1155 ), .Z(_AES_ENC_n1153 ) );
XOR2_X2 _AES_ENC_U1058  ( .A(_AES_ENC_n1230 ), .B(_AES_ENC_n1228 ), .Z(_AES_ENC_n1154 ) );
XOR2_X2 _AES_ENC_U1057  ( .A(_AES_ENC_sa21_sub[1] ), .B(_AES_ENC_sa32_sub[0] ), .Z(_AES_ENC_n1155 ) );
XOR2_X2 _AES_ENC_U1056  ( .A(_AES_ENC_w3[1] ), .B(_AES_ENC_sa03_sub[0] ),.Z(_AES_ENC_n1156 ) );
XOR2_X2 _AES_ENC_U1055  ( .A(_AES_ENC_n1158 ), .B(_AES_ENC_n1157 ), .Z(__AES_ENC_sa33_next[0]) );
XOR2_X2 _AES_ENC_U1054  ( .A(_AES_ENC_n1230 ), .B(_AES_ENC_n1229 ), .Z(_AES_ENC_n1157 ) );
XOR2_X2 _AES_ENC_U1053  ( .A(_AES_ENC_w3[0] ), .B(_AES_ENC_sa21_sub[0] ),.Z(_AES_ENC_n1158 ) );
CLKBUFX1 gbuf_d_395(.A(_AES_ENC_n795), .Y(d_out_395));
CLKBUFX1 gbuf_q_395(.A(q_in_395), .Y(_AES_ENC_n1234));
CLKBUFX1 gbuf_d_396(.A(_AES_ENC_n796), .Y(d_out_396));
CLKBUFX1 gbuf_q_396(.A(q_in_396), .Y(_AES_ENC_n1231));
CLKBUFX1 gbuf_qn_396(.A(qn_in_396), .Y(_AES_ENC_n794));
CLKBUFX1 gbuf_d_397(.A(_AES_ENC_n797), .Y(d_out_397));
CLKBUFX1 gbuf_q_397(.A(q_in_397), .Y(_AES_ENC_n1233));
CLKBUFX1 gbuf_qn_397(.A(qn_in_397), .Y(_AES_ENC_n792));
CLKBUFX1 gbuf_d_398(.A(_AES_ENC_n798), .Y(d_out_398));
CLKBUFX1 gbuf_q_398(.A(q_in_398), .Y(_AES_ENC_n1232));
CLKBUFX1 gbuf_qn_398(.A(qn_in_398), .Y(_AES_ENC_n2));
INV_X4 _AES_ENC_u0_U558  ( .A(_AES_ENC_n1235 ), .ZN(_AES_ENC_u0_n319 ) );
INV_X4 _AES_ENC_u0_U557  ( .A(_AES_ENC_n1235 ), .ZN(_AES_ENC_u0_n325 ) );
INV_X4 _AES_ENC_u0_U556  ( .A(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n324 ) );
INV_X4 _AES_ENC_u0_U555  ( .A(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n322 ) );
INV_X4 _AES_ENC_u0_U554  ( .A(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n323 ) );
INV_X4 _AES_ENC_u0_U553  ( .A(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n321 ) );
INV_X4 _AES_ENC_u0_U552  ( .A(_AES_ENC_n1235 ), .ZN(_AES_ENC_u0_n320 ) );
INV_X4 _AES_ENC_u0_U551  ( .A(_AES_ENC_u0_n319 ), .ZN(_AES_ENC_u0_n318 ) );
INV_X4 _AES_ENC_u0_U550  ( .A(_AES_ENC_u0_n320 ), .ZN(_AES_ENC_u0_n317 ) );
INV_X4 _AES_ENC_u0_U549  ( .A(_AES_ENC_u0_n319 ), .ZN(_AES_ENC_u0_n316 ) );
INV_X4 _AES_ENC_u0_U548  ( .A(_AES_ENC_u0_n319 ), .ZN(_AES_ENC_u0_n315 ) );
NAND2_X1 _AES_ENC_u0_U411  ( .A1(n17502), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n870 ) );
NAND2_X1 _AES_ENC_u0_U410  ( .A1(n17501), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1520 ) );
NAND2_X1 _AES_ENC_u0_U407  ( .A1(n17500), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n630 ) );
NAND2_X1 _AES_ENC_u0_U404  ( .A1(n17499), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1360 ) );
NAND2_X1 _AES_ENC_u0_U401  ( .A1(n17498), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2000 ) );
NAND2_X1 _AES_ENC_u0_U398  ( .A1(n17497), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2640 ) );
NAND2_X1 _AES_ENC_u0_U395  ( .A1(n17496), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n600 ) );
NAND2_X1 _AES_ENC_u0_U392  ( .A1(n17495), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1340 ) );
NAND2_X1 _AES_ENC_u0_U389  ( .A1(n17494), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1980 ) );
NAND2_X1 _AES_ENC_u0_U386  ( .A1(n17493), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2620 ) );
NAND2_X1 _AES_ENC_u0_U383  ( .A1(n17492), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n570 ) );
NAND2_X1 _AES_ENC_u0_U380  ( .A1(n17491), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1320 ) );
NAND2_X1 _AES_ENC_u0_U377  ( .A1(n17490), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1960 ) );
NAND2_X1 _AES_ENC_u0_U374  ( .A1(n17489), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2600 ) );
NAND2_X1 _AES_ENC_u0_U371  ( .A1(n17488), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n540 ) );
NAND2_X1 _AES_ENC_u0_U368  ( .A1(n17487), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1300 ) );
NAND2_X1 _AES_ENC_u0_U365  ( .A1(n17486), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1940 ) );
NAND2_X1 _AES_ENC_u0_U362  ( .A1(n17485), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2580 ) );
NAND2_X1 _AES_ENC_u0_U359  ( .A1(n17484), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n510 ) );
NAND2_X1 _AES_ENC_u0_U356  ( .A1(n17483), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1280 ) );
NAND2_X1 _AES_ENC_u0_U353  ( .A1(n17482), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1920 ) );
NAND2_X1 _AES_ENC_u0_U350  ( .A1(n17481), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2560 ) );
NAND2_X1 _AES_ENC_u0_U347  ( .A1(n17480), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n480 ) );
NAND2_X1 _AES_ENC_u0_U344  ( .A1(n17479), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1260 ) );
NAND2_X1 _AES_ENC_u0_U341  ( .A1(n17478), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1900 ) );
NAND2_X1 _AES_ENC_u0_U338  ( .A1(n17477), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2540 ) );
NAND2_X1 _AES_ENC_u0_U335  ( .A1(n17476), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n450 ) );
NAND2_X1 _AES_ENC_u0_U332  ( .A1(n17475), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1240 ) );
NAND2_X1 _AES_ENC_u0_U329  ( .A1(n17474), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1880 ) );
NAND2_X1 _AES_ENC_u0_U326  ( .A1(n17473), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2520 ) );
NAND2_X1 _AES_ENC_u0_U323  ( .A1(n17472), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n420 ) );
NAND2_X1 _AES_ENC_u0_U320  ( .A1(n17471), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1220 ) );
NAND2_X1 _AES_ENC_u0_U317  ( .A1(n17470), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n39 ) );
NAND2_X1 _AES_ENC_u0_U314  ( .A1(n17469), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1200 ) );
NAND2_X1 _AES_ENC_u0_U311  ( .A1(n17468), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1840 ) );
NAND2_X1 _AES_ENC_u0_U308  ( .A1(n17467), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2480 ) );
NAND2_X1 _AES_ENC_u0_U305  ( .A1(n17466), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n36 ) );
NAND2_X1 _AES_ENC_u0_U30200  ( .A1(n17465), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1180 ) );
NAND2_X1 _AES_ENC_u0_U299  ( .A1(n17464), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1820 ) );
NAND2_X1 _AES_ENC_u0_U296  ( .A1(n17463), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2460 ) );
NAND2_X1 _AES_ENC_u0_U293  ( .A1(n17462), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n33 ) );
NAND2_X1 _AES_ENC_u0_U290  ( .A1(n17461), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1160 ) );
NAND2_X1 _AES_ENC_u0_U287  ( .A1(n17460), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1800 ) );
NAND2_X1 _AES_ENC_u0_U284  ( .A1(n17459), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2440 ) );
NAND2_X1 _AES_ENC_u0_U281  ( .A1(n17458), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n30 ) );
NAND2_X1 _AES_ENC_u0_U278  ( .A1(n17457), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1140 ) );
NAND2_X1 _AES_ENC_u0_U275  ( .A1(n17456), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1780 ) );
NAND2_X1 _AES_ENC_u0_U272  ( .A1(n17455), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2420 ) );
NAND2_X1 _AES_ENC_u0_U269  ( .A1(n17454), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n27 ) );
NAND2_X1 _AES_ENC_u0_U266  ( .A1(n17453), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1120 ) );
NAND2_X1 _AES_ENC_u0_U263  ( .A1(n17452), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1760 ) );
NAND2_X1 _AES_ENC_u0_U260  ( .A1(n17451), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2400 ) );
NAND2_X1 _AES_ENC_u0_U257  ( .A1(n17450), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n24 ) );
NAND2_X1 _AES_ENC_u0_U254  ( .A1(n17449), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1100 ) );
NAND2_X1 _AES_ENC_u0_U251  ( .A1(n17448), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1740 ) );
NAND2_X1 _AES_ENC_u0_U248  ( .A1(n17447), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2380 ) );
NAND2_X1 _AES_ENC_u0_U245  ( .A1(n17446), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n21 ) );
NAND2_X1 _AES_ENC_u0_U242  ( .A1(n17445), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1080 ) );
NAND2_X1 _AES_ENC_u0_U239  ( .A1(n17444), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1720 ) );
NAND2_X1 _AES_ENC_u0_U236  ( .A1(n17443), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2360 ) );
NAND2_X1 _AES_ENC_u0_U233  ( .A1(n17442), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n18 ) );
NAND2_X1 _AES_ENC_u0_U230  ( .A1(n17441), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1060 ) );
NAND2_X1 _AES_ENC_u0_U227  ( .A1(n17440), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1040 ) );
NAND2_X1 _AES_ENC_u0_U224  ( .A1(n17439), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1680 ) );
NAND2_X1 _AES_ENC_u0_U221  ( .A1(n17438), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2320 ) );
NAND2_X1 _AES_ENC_u0_U218  ( .A1(n17437), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1610 ) );
NAND2_X1 _AES_ENC_u0_U215  ( .A1(n17436), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1020 ) );
NAND2_X1 _AES_ENC_u0_U212  ( .A1(n17435), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1660 ) );
NAND2_X1 _AES_ENC_u0_U209  ( .A1(n17434), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2300 ) );
NAND2_X1 _AES_ENC_u0_U206  ( .A1(n17433), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n1400 ) );
NAND2_X1 _AES_ENC_u0_U203  ( .A1(n17432), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1000 ) );
NAND2_X1 _AES_ENC_u0_U200  ( .A1(n17431), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1640 ) );
NAND2_X1 _AES_ENC_u0_U197  ( .A1(n17430), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2280 ) );
NAND2_X1 _AES_ENC_u0_U194  ( .A1(n17429), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1210 ) );
NAND2_X1 _AES_ENC_u0_U191  ( .A1(n17428), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n980 ) );
NAND2_X1 _AES_ENC_u0_U188  ( .A1(n17427), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1620 ) );
NAND2_X1 _AES_ENC_u0_U185  ( .A1(n17426), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2260 ) );
NAND2_X1 _AES_ENC_u0_U182  ( .A1(n17425), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1010 ) );
NAND2_X1 _AES_ENC_u0_U179  ( .A1(n17424), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n960 ) );
NAND2_X1 _AES_ENC_u0_U176  ( .A1(n17423), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1600 ) );
NAND2_X1 _AES_ENC_u0_U173  ( .A1(n17422), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2240 ) );
NAND2_X1 _AES_ENC_u0_U170  ( .A1(n17421), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n8 ) );
NAND2_X1 _AES_ENC_u0_U167  ( .A1(n17420), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n940 ) );
NAND2_X1 _AES_ENC_u0_U164  ( .A1(n17419), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1580 ) );
NAND2_X1 _AES_ENC_u0_U161  ( .A1(n17418), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2220 ) );
NAND2_X1 _AES_ENC_u0_U158  ( .A1(n17417), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n6 ) );
NAND2_X1 _AES_ENC_u0_U155  ( .A1(n17416), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n920 ) );
NAND2_X1 _AES_ENC_u0_U152  ( .A1(n17415), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1560 ) );
NAND2_X1 _AES_ENC_u0_U149  ( .A1(n17414), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2200 ) );
NAND2_X1 _AES_ENC_u0_U146  ( .A1(n17413), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n4 ) );
NAND2_X1 _AES_ENC_u0_U143  ( .A1(n17412), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n900 ) );
NAND2_X1 _AES_ENC_u0_U140  ( .A1(n17411), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n840 ) );
NAND2_X1 _AES_ENC_u0_U137  ( .A1(n17410), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1500 ) );
NAND2_X1 _AES_ENC_u0_U134  ( .A1(n17409), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2140 ) );
NAND2_X1 _AES_ENC_u0_U131  ( .A1(n17408), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n278 ) );
NAND2_X1 _AES_ENC_u0_U128  ( .A1(n17407), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n810 ) );
NAND2_X1 _AES_ENC_u0_U125  ( .A1(n17406), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1480 ) );
NAND2_X1 _AES_ENC_u0_U122  ( .A1(n17405), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2120 ) );
NAND2_X1 _AES_ENC_u0_U118  ( .A1(n17404), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n276 ) );
NAND2_X1 _AES_ENC_u0_U114  ( .A1(n17403), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n780 ) );
NAND2_X1 _AES_ENC_u0_U110  ( .A1(n17402), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1460 ) );
NAND2_X1 _AES_ENC_u0_U106  ( .A1(n17401), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2100 ) );
NAND2_X1 _AES_ENC_u0_U102  ( .A1(n17400), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n274 ) );
NAND2_X1 _AES_ENC_u0_U98  ( .A1(n17399), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n75 ) );
NAND2_X1 _AES_ENC_u0_U94  ( .A1(n17398), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1440 ) );
NAND2_X1 _AES_ENC_u0_U90  ( .A1(n17397), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2080 ) );
NAND2_X1 _AES_ENC_u0_U86  ( .A1(n17396), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n272 ) );
NAND2_X1 _AES_ENC_u0_U82  ( .A1(n17395), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n720 ) );
NAND2_X1 _AES_ENC_u0_U78  ( .A1(n17394), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1420 ) );
NAND2_X1 _AES_ENC_u0_U74  ( .A1(n17393), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n206 ) );
NAND2_X1 _AES_ENC_u0_U70  ( .A1(n17392), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2700 ) );
NAND2_X1 _AES_ENC_u0_U66  ( .A1(n17391), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n690 ) );
NAND2_X1 _AES_ENC_u0_U62  ( .A1(n17390), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1401 ) );
NAND2_X1 _AES_ENC_u0_U58  ( .A1(n17389), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2040 ) );
NAND2_X1 _AES_ENC_u0_U54  ( .A1(n17388), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2680 ) );
NAND2_X1 _AES_ENC_u0_U50  ( .A1(n17387), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n660 ) );
NAND2_X1 _AES_ENC_u0_U46  ( .A1(n17386), .A2(_AES_ENC_u0_n317 ), .ZN(_AES_ENC_u0_n1380 ) );
NAND2_X1 _AES_ENC_u0_U42  ( .A1(n17385), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2020 ) );
NAND2_X1 _AES_ENC_u0_U38  ( .A1(n17384), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2660 ) );
NAND2_X1 _AES_ENC_u0_U34  ( .A1(n17383), .A2(_AES_ENC_u0_n316 ), .ZN(_AES_ENC_u0_n1540 ) );
NAND2_X1 _AES_ENC_u0_U3020  ( .A1(n17382), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2180 ) );
NAND2_X1 _AES_ENC_u0_U26  ( .A1(_AES_ENC_u0_n316 ), .A2(cii_K[127]), .ZN(_AES_ENC_u0_n2 ) );
NAND2_X1 _AES_ENC_u0_U23  ( .A1(_AES_ENC_u0_n2 ), .A2(_AES_ENC_u0_n3 ), .ZN(_AES_ENC_u0_N73 ) );
BUF_X32 _AES_ENC_u0_U20  ( .A(_AES_ENC_u0_N73 ), .Z(_AES_ENC_u0_n314 ) );
NAND2_X1 _AES_ENC_u0_U17  ( .A1(n17381), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1700 ) );
NAND2_X1 _AES_ENC_u0_U14  ( .A1(n17380), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2340 ) );
NAND2_X1 _AES_ENC_u0_U11  ( .A1(n17379), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n1860 ) );
NAND2_X1 _AES_ENC_u0_U8  ( .A1(n17378), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2500 ) );
NAND2_X1 _AES_ENC_u0_U5  ( .A1(n17377), .A2(_AES_ENC_u0_n318 ), .ZN(_AES_ENC_u0_n2160 ) );
NAND2_X1 _AES_ENC_u0_U3010  ( .A1(n17376), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_n280 ) );
NAND2_X2 _AES_ENC_u0_U409  ( .A1(_AES_ENC_u0_N107 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n281 ) );
NAND2_X2 _AES_ENC_u0_U408  ( .A1(_AES_ENC_u0_n280 ), .A2(_AES_ENC_u0_n281 ),.ZN(_AES_ENC_u0_N108 ) );
NAND2_X2 _AES_ENC_u0_U406  ( .A1(_AES_ENC_u0_N106 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n279 ) );
NAND2_X2 _AES_ENC_u0_U405  ( .A1(_AES_ENC_u0_n278 ), .A2(_AES_ENC_u0_n279 ),.ZN(_AES_ENC_u0_N109 ) );
NAND2_X2 _AES_ENC_u0_U403  ( .A1(_AES_ENC_u0_N105 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n277 ) );
NAND2_X2 _AES_ENC_u0_U402  ( .A1(_AES_ENC_u0_n276 ), .A2(_AES_ENC_u0_n277 ),.ZN(_AES_ENC_u0_N110 ) );
NAND2_X2 _AES_ENC_u0_U400  ( .A1(_AES_ENC_u0_N104 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n275 ) );
NAND2_X2 _AES_ENC_u0_U399  ( .A1(_AES_ENC_u0_n274 ), .A2(_AES_ENC_u0_n275 ),.ZN(_AES_ENC_u0_N111 ) );
NAND2_X2 _AES_ENC_u0_U397  ( .A1(_AES_ENC_u0_N103 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n273 ) );
NAND2_X2 _AES_ENC_u0_U396  ( .A1(_AES_ENC_u0_n272 ), .A2(_AES_ENC_u0_n273 ),.ZN(_AES_ENC_u0_N112 ) );
NAND2_X2 _AES_ENC_u0_U394  ( .A1(_AES_ENC_u0_N102 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n2710 ) );
NAND2_X2 _AES_ENC_u0_U393  ( .A1(_AES_ENC_u0_n2700 ), .A2(_AES_ENC_u0_n2710 ), .ZN(_AES_ENC_u0_N113 ) );
NAND2_X2 _AES_ENC_u0_U391  ( .A1(_AES_ENC_u0_N101 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n2690 ) );
NAND2_X2 _AES_ENC_u0_U390  ( .A1(_AES_ENC_u0_n2680 ), .A2(_AES_ENC_u0_n2690 ), .ZN(_AES_ENC_u0_N114 ) );
NAND2_X2 _AES_ENC_u0_U388  ( .A1(_AES_ENC_u0_N100 ), .A2(_AES_ENC_u0_n319 ),.ZN(_AES_ENC_u0_n2670 ) );
NAND2_X2 _AES_ENC_u0_U387  ( .A1(_AES_ENC_u0_n2660 ), .A2(_AES_ENC_u0_n2670 ), .ZN(_AES_ENC_u0_N115 ) );
NAND2_X2 _AES_ENC_u0_U385  ( .A1(_AES_ENC_u0_N99 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2650 ) );
NAND2_X2 _AES_ENC_u0_U384  ( .A1(_AES_ENC_u0_n2640 ), .A2(_AES_ENC_u0_n2650 ), .ZN(_AES_ENC_u0_N116 ) );
NAND2_X2 _AES_ENC_u0_U382  ( .A1(_AES_ENC_u0_N98 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2630 ) );
NAND2_X2 _AES_ENC_u0_U381  ( .A1(_AES_ENC_u0_n2620 ), .A2(_AES_ENC_u0_n2630 ), .ZN(_AES_ENC_u0_N117 ) );
NAND2_X2 _AES_ENC_u0_U379  ( .A1(_AES_ENC_u0_N97 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2610 ) );
NAND2_X2 _AES_ENC_u0_U378  ( .A1(_AES_ENC_u0_n2600 ), .A2(_AES_ENC_u0_n2610 ), .ZN(_AES_ENC_u0_N118 ) );
NAND2_X2 _AES_ENC_u0_U376  ( .A1(_AES_ENC_u0_N96 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2590 ) );
NAND2_X2 _AES_ENC_u0_U375  ( .A1(_AES_ENC_u0_n2580 ), .A2(_AES_ENC_u0_n2590 ), .ZN(_AES_ENC_u0_N119 ) );
NAND2_X2 _AES_ENC_u0_U373  ( .A1(_AES_ENC_u0_N95 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2570 ) );
NAND2_X2 _AES_ENC_u0_U372  ( .A1(_AES_ENC_u0_n2560 ), .A2(_AES_ENC_u0_n2570 ), .ZN(_AES_ENC_u0_N120 ) );
NAND2_X2 _AES_ENC_u0_U370  ( .A1(_AES_ENC_u0_N94 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2550 ) );
NAND2_X2 _AES_ENC_u0_U369  ( .A1(_AES_ENC_u0_n2540 ), .A2(_AES_ENC_u0_n2550 ), .ZN(_AES_ENC_u0_N121 ) );
NAND2_X2 _AES_ENC_u0_U367  ( .A1(_AES_ENC_u0_N93 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2530 ) );
NAND2_X2 _AES_ENC_u0_U366  ( .A1(_AES_ENC_u0_n2520 ), .A2(_AES_ENC_u0_n2530 ), .ZN(_AES_ENC_u0_N122 ) );
NAND2_X2 _AES_ENC_u0_U364  ( .A1(_AES_ENC_u0_N92 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2510 ) );
NAND2_X2 _AES_ENC_u0_U363  ( .A1(_AES_ENC_u0_n2500 ), .A2(_AES_ENC_u0_n2510 ), .ZN(_AES_ENC_u0_N123 ) );
NAND2_X2 _AES_ENC_u0_U361  ( .A1(_AES_ENC_u0_N91 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2490 ) );
NAND2_X2 _AES_ENC_u0_U360  ( .A1(_AES_ENC_u0_n2480 ), .A2(_AES_ENC_u0_n2490 ), .ZN(_AES_ENC_u0_N124 ) );
NAND2_X2 _AES_ENC_u0_U358  ( .A1(_AES_ENC_u0_N90 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2470 ) );
NAND2_X2 _AES_ENC_u0_U357  ( .A1(_AES_ENC_u0_n2460 ), .A2(_AES_ENC_u0_n2470 ), .ZN(_AES_ENC_u0_N125 ) );
NAND2_X2 _AES_ENC_u0_U355  ( .A1(_AES_ENC_u0_N89 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2450 ) );
NAND2_X2 _AES_ENC_u0_U354  ( .A1(_AES_ENC_u0_n2440 ), .A2(_AES_ENC_u0_n2450 ), .ZN(_AES_ENC_u0_N126 ) );
NAND2_X2 _AES_ENC_u0_U352  ( .A1(_AES_ENC_u0_N88 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2430 ) );
NAND2_X2 _AES_ENC_u0_U351  ( .A1(_AES_ENC_u0_n2420 ), .A2(_AES_ENC_u0_n2430 ), .ZN(_AES_ENC_u0_N127 ) );
NAND2_X2 _AES_ENC_u0_U349  ( .A1(_AES_ENC_u0_N87 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2410 ) );
NAND2_X2 _AES_ENC_u0_U348  ( .A1(_AES_ENC_u0_n2400 ), .A2(_AES_ENC_u0_n2410 ), .ZN(_AES_ENC_u0_N128 ) );
NAND2_X2 _AES_ENC_u0_U346  ( .A1(_AES_ENC_u0_N86 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2390 ) );
NAND2_X2 _AES_ENC_u0_U345  ( .A1(_AES_ENC_u0_n2380 ), .A2(_AES_ENC_u0_n2390 ), .ZN(_AES_ENC_u0_N129 ) );
NAND2_X2 _AES_ENC_u0_U343  ( .A1(_AES_ENC_u0_N85 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2370 ) );
NAND2_X2 _AES_ENC_u0_U342  ( .A1(_AES_ENC_u0_n2360 ), .A2(_AES_ENC_u0_n2370 ), .ZN(_AES_ENC_u0_N130 ) );
NAND2_X2 _AES_ENC_u0_U340  ( .A1(_AES_ENC_u0_N84 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2350 ) );
NAND2_X2 _AES_ENC_u0_U339  ( .A1(_AES_ENC_u0_n2340 ), .A2(_AES_ENC_u0_n2350 ), .ZN(_AES_ENC_u0_N131 ) );
NAND2_X2 _AES_ENC_u0_U337  ( .A1(_AES_ENC_u0_N83 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2330 ) );
NAND2_X2 _AES_ENC_u0_U336  ( .A1(_AES_ENC_u0_n2320 ), .A2(_AES_ENC_u0_n2330 ), .ZN(_AES_ENC_u0_N132 ) );
NAND2_X2 _AES_ENC_u0_U334  ( .A1(_AES_ENC_u0_N82 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2310 ) );
NAND2_X2 _AES_ENC_u0_U333  ( .A1(_AES_ENC_u0_n2300 ), .A2(_AES_ENC_u0_n2310 ), .ZN(_AES_ENC_u0_N133 ) );
NAND2_X2 _AES_ENC_u0_U331  ( .A1(_AES_ENC_u0_N81 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2290 ) );
NAND2_X2 _AES_ENC_u0_U330  ( .A1(_AES_ENC_u0_n2280 ), .A2(_AES_ENC_u0_n2290 ), .ZN(_AES_ENC_u0_N134 ) );
NAND2_X2 _AES_ENC_u0_U328  ( .A1(_AES_ENC_u0_N80 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2270 ) );
NAND2_X2 _AES_ENC_u0_U327  ( .A1(_AES_ENC_u0_n2260 ), .A2(_AES_ENC_u0_n2270 ), .ZN(_AES_ENC_u0_N135 ) );
NAND2_X2 _AES_ENC_u0_U325  ( .A1(_AES_ENC_u0_N79 ), .A2(_AES_ENC_u0_n320 ),.ZN(_AES_ENC_u0_n2250 ) );
NAND2_X2 _AES_ENC_u0_U324  ( .A1(_AES_ENC_u0_n2240 ), .A2(_AES_ENC_u0_n2250 ), .ZN(_AES_ENC_u0_N136 ) );
NAND2_X2 _AES_ENC_u0_U322  ( .A1(_AES_ENC_u0_N78 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2230 ) );
NAND2_X2 _AES_ENC_u0_U321  ( .A1(_AES_ENC_u0_n2220 ), .A2(_AES_ENC_u0_n2230 ), .ZN(_AES_ENC_u0_N137 ) );
NAND2_X2 _AES_ENC_u0_U319  ( .A1(_AES_ENC_u0_N77 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2210 ) );
NAND2_X2 _AES_ENC_u0_U318  ( .A1(_AES_ENC_u0_n2200 ), .A2(_AES_ENC_u0_n2210 ), .ZN(_AES_ENC_u0_N138 ) );
NAND2_X2 _AES_ENC_u0_U316  ( .A1(_AES_ENC_u0_N76 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2190 ) );
NAND2_X2 _AES_ENC_u0_U315  ( .A1(_AES_ENC_u0_n2180 ), .A2(_AES_ENC_u0_n2190 ), .ZN(_AES_ENC_u0_N139 ) );
NAND2_X2 _AES_ENC_u0_U313  ( .A1(_AES_ENC_u0_N173 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2170 ) );
NAND2_X2 _AES_ENC_u0_U312  ( .A1(_AES_ENC_u0_n2160 ), .A2(_AES_ENC_u0_n2170 ), .ZN(_AES_ENC_u0_N174 ) );
NAND2_X2 _AES_ENC_u0_U310  ( .A1(_AES_ENC_u0_N172 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2150 ) );
NAND2_X2 _AES_ENC_u0_U309  ( .A1(_AES_ENC_u0_n2140 ), .A2(_AES_ENC_u0_n2150 ), .ZN(_AES_ENC_u0_N175 ) );
NAND2_X2 _AES_ENC_u0_U307  ( .A1(_AES_ENC_u0_N171 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2130 ) );
NAND2_X2 _AES_ENC_u0_U306  ( .A1(_AES_ENC_u0_n2120 ), .A2(_AES_ENC_u0_n2130 ), .ZN(_AES_ENC_u0_N176 ) );
NAND2_X2 _AES_ENC_u0_U304  ( .A1(_AES_ENC_u0_N170 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2110 ) );
NAND2_X2 _AES_ENC_u0_U303  ( .A1(_AES_ENC_u0_n2100 ), .A2(_AES_ENC_u0_n2110 ), .ZN(_AES_ENC_u0_N177 ) );
NAND2_X2 _AES_ENC_u0_U301  ( .A1(_AES_ENC_u0_N169 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2090 ) );
NAND2_X2 _AES_ENC_u0_U300  ( .A1(_AES_ENC_u0_n2080 ), .A2(_AES_ENC_u0_n2090 ), .ZN(_AES_ENC_u0_N178 ) );
NAND2_X2 _AES_ENC_u0_U298  ( .A1(_AES_ENC_u0_N168 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n207 ) );
NAND2_X2 _AES_ENC_u0_U297  ( .A1(_AES_ENC_u0_n206 ), .A2(_AES_ENC_u0_n207 ),.ZN(_AES_ENC_u0_N179 ) );
NAND2_X2 _AES_ENC_u0_U295  ( .A1(_AES_ENC_u0_N167 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2050 ) );
NAND2_X2 _AES_ENC_u0_U294  ( .A1(_AES_ENC_u0_n2040 ), .A2(_AES_ENC_u0_n2050 ), .ZN(_AES_ENC_u0_N180 ) );
NAND2_X2 _AES_ENC_u0_U292  ( .A1(_AES_ENC_u0_N166 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2030 ) );
NAND2_X2 _AES_ENC_u0_U291  ( .A1(_AES_ENC_u0_n2020 ), .A2(_AES_ENC_u0_n2030 ), .ZN(_AES_ENC_u0_N181 ) );
NAND2_X2 _AES_ENC_u0_U289  ( .A1(_AES_ENC_u0_N165 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n2010 ) );
NAND2_X2 _AES_ENC_u0_U288  ( .A1(_AES_ENC_u0_n2000 ), .A2(_AES_ENC_u0_n2010 ), .ZN(_AES_ENC_u0_N182 ) );
NAND2_X2 _AES_ENC_u0_U286  ( .A1(_AES_ENC_u0_N164 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1990 ) );
NAND2_X2 _AES_ENC_u0_U285  ( .A1(_AES_ENC_u0_n1980 ), .A2(_AES_ENC_u0_n1990 ), .ZN(_AES_ENC_u0_N183 ) );
NAND2_X2 _AES_ENC_u0_U283  ( .A1(_AES_ENC_u0_N163 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1970 ) );
NAND2_X2 _AES_ENC_u0_U282  ( .A1(_AES_ENC_u0_n1960 ), .A2(_AES_ENC_u0_n1970 ), .ZN(_AES_ENC_u0_N184 ) );
NAND2_X2 _AES_ENC_u0_U280  ( .A1(_AES_ENC_u0_N162 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1950 ) );
NAND2_X2 _AES_ENC_u0_U279  ( .A1(_AES_ENC_u0_n1940 ), .A2(_AES_ENC_u0_n1950 ), .ZN(_AES_ENC_u0_N185 ) );
NAND2_X2 _AES_ENC_u0_U277  ( .A1(_AES_ENC_u0_N161 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1930 ) );
NAND2_X2 _AES_ENC_u0_U276  ( .A1(_AES_ENC_u0_n1920 ), .A2(_AES_ENC_u0_n1930 ), .ZN(_AES_ENC_u0_N186 ) );
NAND2_X2 _AES_ENC_u0_U274  ( .A1(_AES_ENC_u0_N160 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1910 ) );
NAND2_X2 _AES_ENC_u0_U273  ( .A1(_AES_ENC_u0_n1900 ), .A2(_AES_ENC_u0_n1910 ), .ZN(_AES_ENC_u0_N187 ) );
NAND2_X2 _AES_ENC_u0_U271  ( .A1(_AES_ENC_u0_N159 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1890 ) );
NAND2_X2 _AES_ENC_u0_U270  ( .A1(_AES_ENC_u0_n1880 ), .A2(_AES_ENC_u0_n1890 ), .ZN(_AES_ENC_u0_N188 ) );
NAND2_X2 _AES_ENC_u0_U268  ( .A1(_AES_ENC_u0_N158 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1870 ) );
NAND2_X2 _AES_ENC_u0_U267  ( .A1(_AES_ENC_u0_n1860 ), .A2(_AES_ENC_u0_n1870 ), .ZN(_AES_ENC_u0_N189 ) );
NAND2_X2 _AES_ENC_u0_U265  ( .A1(_AES_ENC_u0_N157 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1850 ) );
NAND2_X2 _AES_ENC_u0_U264  ( .A1(_AES_ENC_u0_n1840 ), .A2(_AES_ENC_u0_n1850 ), .ZN(_AES_ENC_u0_N190 ) );
NAND2_X2 _AES_ENC_u0_U262  ( .A1(_AES_ENC_u0_N156 ), .A2(_AES_ENC_u0_n321 ),.ZN(_AES_ENC_u0_n1830 ) );
NAND2_X2 _AES_ENC_u0_U261  ( .A1(_AES_ENC_u0_n1820 ), .A2(_AES_ENC_u0_n1830 ), .ZN(_AES_ENC_u0_N191 ) );
NAND2_X2 _AES_ENC_u0_U259  ( .A1(_AES_ENC_u0_N155 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1810 ) );
NAND2_X2 _AES_ENC_u0_U258  ( .A1(_AES_ENC_u0_n1800 ), .A2(_AES_ENC_u0_n1810 ), .ZN(_AES_ENC_u0_N192 ) );
NAND2_X2 _AES_ENC_u0_U256  ( .A1(_AES_ENC_u0_N154 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1790 ) );
NAND2_X2 _AES_ENC_u0_U255  ( .A1(_AES_ENC_u0_n1780 ), .A2(_AES_ENC_u0_n1790 ), .ZN(_AES_ENC_u0_N193 ) );
NAND2_X2 _AES_ENC_u0_U253  ( .A1(_AES_ENC_u0_N153 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1770 ) );
NAND2_X2 _AES_ENC_u0_U252  ( .A1(_AES_ENC_u0_n1760 ), .A2(_AES_ENC_u0_n1770 ), .ZN(_AES_ENC_u0_N194 ) );
NAND2_X2 _AES_ENC_u0_U250  ( .A1(_AES_ENC_u0_N152 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1750 ) );
NAND2_X2 _AES_ENC_u0_U249  ( .A1(_AES_ENC_u0_n1740 ), .A2(_AES_ENC_u0_n1750 ), .ZN(_AES_ENC_u0_N195 ) );
NAND2_X2 _AES_ENC_u0_U247  ( .A1(_AES_ENC_u0_N151 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1730 ) );
NAND2_X2 _AES_ENC_u0_U246  ( .A1(_AES_ENC_u0_n1720 ), .A2(_AES_ENC_u0_n1730 ), .ZN(_AES_ENC_u0_N196 ) );
NAND2_X2 _AES_ENC_u0_U244  ( .A1(_AES_ENC_u0_N150 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1711 ) );
NAND2_X2 _AES_ENC_u0_U243  ( .A1(_AES_ENC_u0_n1700 ), .A2(_AES_ENC_u0_n1711 ), .ZN(_AES_ENC_u0_N197 ) );
NAND2_X2 _AES_ENC_u0_U241  ( .A1(_AES_ENC_u0_N149 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1690 ) );
NAND2_X2 _AES_ENC_u0_U240  ( .A1(_AES_ENC_u0_n1680 ), .A2(_AES_ENC_u0_n1690 ), .ZN(_AES_ENC_u0_N198 ) );
NAND2_X2 _AES_ENC_u0_U238  ( .A1(_AES_ENC_u0_N148 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1670 ) );
NAND2_X2 _AES_ENC_u0_U237  ( .A1(_AES_ENC_u0_n1660 ), .A2(_AES_ENC_u0_n1670 ), .ZN(_AES_ENC_u0_N199 ) );
NAND2_X2 _AES_ENC_u0_U235  ( .A1(_AES_ENC_u0_N147 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1650 ) );
NAND2_X2 _AES_ENC_u0_U234  ( .A1(_AES_ENC_u0_n1640 ), .A2(_AES_ENC_u0_n1650 ), .ZN(_AES_ENC_u0_N200 ) );
NAND2_X2 _AES_ENC_u0_U232  ( .A1(_AES_ENC_u0_N146 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1630 ) );
NAND2_X2 _AES_ENC_u0_U231  ( .A1(_AES_ENC_u0_n1620 ), .A2(_AES_ENC_u0_n1630 ), .ZN(_AES_ENC_u0_N201 ) );
NAND2_X2 _AES_ENC_u0_U229  ( .A1(_AES_ENC_u0_N145 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1611 ) );
NAND2_X2 _AES_ENC_u0_U228  ( .A1(_AES_ENC_u0_n1600 ), .A2(_AES_ENC_u0_n1611 ), .ZN(_AES_ENC_u0_N202 ) );
NAND2_X2 _AES_ENC_u0_U226  ( .A1(_AES_ENC_u0_N144 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1590 ) );
NAND2_X2 _AES_ENC_u0_U225  ( .A1(_AES_ENC_u0_n1580 ), .A2(_AES_ENC_u0_n1590 ), .ZN(_AES_ENC_u0_N203 ) );
NAND2_X2 _AES_ENC_u0_U223  ( .A1(_AES_ENC_u0_N143 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1570 ) );
NAND2_X2 _AES_ENC_u0_U222  ( .A1(_AES_ENC_u0_n1560 ), .A2(_AES_ENC_u0_n1570 ), .ZN(_AES_ENC_u0_N204 ) );
NAND2_X2 _AES_ENC_u0_U220  ( .A1(_AES_ENC_u0_N142 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1550 ) );
NAND2_X2 _AES_ENC_u0_U219  ( .A1(_AES_ENC_u0_n1540 ), .A2(_AES_ENC_u0_n1550 ), .ZN(_AES_ENC_u0_N205 ) );
NAND2_X2 _AES_ENC_u0_U217  ( .A1(_AES_ENC_u0_N239 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1530 ) );
NAND2_X2 _AES_ENC_u0_U216  ( .A1(_AES_ENC_u0_n1520 ), .A2(_AES_ENC_u0_n1530 ), .ZN(_AES_ENC_u0_N240 ) );
NAND2_X2 _AES_ENC_u0_U214  ( .A1(_AES_ENC_u0_N238 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1511 ) );
NAND2_X2 _AES_ENC_u0_U213  ( .A1(_AES_ENC_u0_n1500 ), .A2(_AES_ENC_u0_n1511 ), .ZN(_AES_ENC_u0_N241 ) );
NAND2_X2 _AES_ENC_u0_U211  ( .A1(_AES_ENC_u0_N237 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1490 ) );
NAND2_X2 _AES_ENC_u0_U210  ( .A1(_AES_ENC_u0_n1480 ), .A2(_AES_ENC_u0_n1490 ), .ZN(_AES_ENC_u0_N242 ) );
NAND2_X2 _AES_ENC_u0_U208  ( .A1(_AES_ENC_u0_N236 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1470 ) );
NAND2_X2 _AES_ENC_u0_U207  ( .A1(_AES_ENC_u0_n1460 ), .A2(_AES_ENC_u0_n1470 ), .ZN(_AES_ENC_u0_N243 ) );
NAND2_X2 _AES_ENC_u0_U205  ( .A1(_AES_ENC_u0_N235 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1450 ) );
NAND2_X2 _AES_ENC_u0_U204  ( .A1(_AES_ENC_u0_n1440 ), .A2(_AES_ENC_u0_n1450 ), .ZN(_AES_ENC_u0_N244 ) );
NAND2_X2 _AES_ENC_u0_U202  ( .A1(_AES_ENC_u0_N234 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n1430 ) );
NAND2_X2 _AES_ENC_u0_U201  ( .A1(_AES_ENC_u0_n1420 ), .A2(_AES_ENC_u0_n1430 ), .ZN(_AES_ENC_u0_N245 ) );
NAND2_X2 _AES_ENC_u0_U199  ( .A1(_AES_ENC_u0_N233 ), .A2(_AES_ENC_u0_n322 ),.ZN(_AES_ENC_u0_n141 ) );
NAND2_X2 _AES_ENC_u0_U198  ( .A1(_AES_ENC_u0_n1401 ), .A2(_AES_ENC_u0_n141 ),.ZN(_AES_ENC_u0_N246 ) );
NAND2_X2 _AES_ENC_u0_U196  ( .A1(_AES_ENC_u0_N232 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1390 ) );
NAND2_X2 _AES_ENC_u0_U195  ( .A1(_AES_ENC_u0_n1380 ), .A2(_AES_ENC_u0_n1390 ), .ZN(_AES_ENC_u0_N247 ) );
NAND2_X2 _AES_ENC_u0_U193  ( .A1(_AES_ENC_u0_N231 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1370 ) );
NAND2_X2 _AES_ENC_u0_U192  ( .A1(_AES_ENC_u0_n1360 ), .A2(_AES_ENC_u0_n1370 ), .ZN(_AES_ENC_u0_N248 ) );
NAND2_X2 _AES_ENC_u0_U190  ( .A1(_AES_ENC_u0_N230 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1350 ) );
NAND2_X2 _AES_ENC_u0_U189  ( .A1(_AES_ENC_u0_n1340 ), .A2(_AES_ENC_u0_n1350 ), .ZN(_AES_ENC_u0_N249 ) );
NAND2_X2 _AES_ENC_u0_U187  ( .A1(_AES_ENC_u0_N229 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1330 ) );
NAND2_X2 _AES_ENC_u0_U186  ( .A1(_AES_ENC_u0_n1320 ), .A2(_AES_ENC_u0_n1330 ), .ZN(_AES_ENC_u0_N250 ) );
NAND2_X2 _AES_ENC_u0_U184  ( .A1(_AES_ENC_u0_N228 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1311 ) );
NAND2_X2 _AES_ENC_u0_U183  ( .A1(_AES_ENC_u0_n1300 ), .A2(_AES_ENC_u0_n1311 ), .ZN(_AES_ENC_u0_N251 ) );
NAND2_X2 _AES_ENC_u0_U181  ( .A1(_AES_ENC_u0_N227 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1290 ) );
NAND2_X2 _AES_ENC_u0_U180  ( .A1(_AES_ENC_u0_n1280 ), .A2(_AES_ENC_u0_n1290 ), .ZN(_AES_ENC_u0_N252 ) );
NAND2_X2 _AES_ENC_u0_U178  ( .A1(_AES_ENC_u0_N226 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1270 ) );
NAND2_X2 _AES_ENC_u0_U177  ( .A1(_AES_ENC_u0_n1260 ), .A2(_AES_ENC_u0_n1270 ), .ZN(_AES_ENC_u0_N253 ) );
NAND2_X2 _AES_ENC_u0_U175  ( .A1(_AES_ENC_u0_N225 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1250 ) );
NAND2_X2 _AES_ENC_u0_U174  ( .A1(_AES_ENC_u0_n1240 ), .A2(_AES_ENC_u0_n1250 ), .ZN(_AES_ENC_u0_N254 ) );
NAND2_X2 _AES_ENC_u0_U172  ( .A1(_AES_ENC_u0_N224 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1230 ) );
NAND2_X2 _AES_ENC_u0_U171  ( .A1(_AES_ENC_u0_n1220 ), .A2(_AES_ENC_u0_n1230 ), .ZN(_AES_ENC_u0_N255 ) );
NAND2_X2 _AES_ENC_u0_U169  ( .A1(_AES_ENC_u0_N223 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1211 ) );
NAND2_X2 _AES_ENC_u0_U168  ( .A1(_AES_ENC_u0_n1200 ), .A2(_AES_ENC_u0_n1211 ), .ZN(_AES_ENC_u0_N256 ) );
NAND2_X2 _AES_ENC_u0_U166  ( .A1(_AES_ENC_u0_N222 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1190 ) );
NAND2_X2 _AES_ENC_u0_U165  ( .A1(_AES_ENC_u0_n1180 ), .A2(_AES_ENC_u0_n1190 ), .ZN(_AES_ENC_u0_N257 ) );
NAND2_X2 _AES_ENC_u0_U163  ( .A1(_AES_ENC_u0_N221 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1170 ) );
NAND2_X2 _AES_ENC_u0_U162  ( .A1(_AES_ENC_u0_n1160 ), .A2(_AES_ENC_u0_n1170 ), .ZN(_AES_ENC_u0_N258 ) );
NAND2_X2 _AES_ENC_u0_U160  ( .A1(_AES_ENC_u0_N220 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1150 ) );
NAND2_X2 _AES_ENC_u0_U159  ( .A1(_AES_ENC_u0_n1140 ), .A2(_AES_ENC_u0_n1150 ), .ZN(_AES_ENC_u0_N259 ) );
NAND2_X2 _AES_ENC_u0_U157  ( .A1(_AES_ENC_u0_N219 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1130 ) );
NAND2_X2 _AES_ENC_u0_U156  ( .A1(_AES_ENC_u0_n1120 ), .A2(_AES_ENC_u0_n1130 ), .ZN(_AES_ENC_u0_N260 ) );
NAND2_X2 _AES_ENC_u0_U154  ( .A1(_AES_ENC_u0_N218 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1111 ) );
NAND2_X2 _AES_ENC_u0_U153  ( .A1(_AES_ENC_u0_n1100 ), .A2(_AES_ENC_u0_n1111 ), .ZN(_AES_ENC_u0_N261 ) );
NAND2_X2 _AES_ENC_u0_U151  ( .A1(_AES_ENC_u0_N217 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1090 ) );
NAND2_X2 _AES_ENC_u0_U150  ( .A1(_AES_ENC_u0_n1080 ), .A2(_AES_ENC_u0_n1090 ), .ZN(_AES_ENC_u0_N262 ) );
NAND2_X2 _AES_ENC_u0_U148  ( .A1(_AES_ENC_u0_N216 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1070 ) );
NAND2_X2 _AES_ENC_u0_U147  ( .A1(_AES_ENC_u0_n1060 ), .A2(_AES_ENC_u0_n1070 ), .ZN(_AES_ENC_u0_N263 ) );
NAND2_X2 _AES_ENC_u0_U145  ( .A1(_AES_ENC_u0_N215 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1050 ) );
NAND2_X2 _AES_ENC_u0_U144  ( .A1(_AES_ENC_u0_n1040 ), .A2(_AES_ENC_u0_n1050 ), .ZN(_AES_ENC_u0_N264 ) );
NAND2_X2 _AES_ENC_u0_U142  ( .A1(_AES_ENC_u0_N214 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1030 ) );
NAND2_X2 _AES_ENC_u0_U141  ( .A1(_AES_ENC_u0_n1020 ), .A2(_AES_ENC_u0_n1030 ), .ZN(_AES_ENC_u0_N265 ) );
NAND2_X2 _AES_ENC_u0_U139  ( .A1(_AES_ENC_u0_N213 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n1011 ) );
NAND2_X2 _AES_ENC_u0_U138  ( .A1(_AES_ENC_u0_n1000 ), .A2(_AES_ENC_u0_n1011 ), .ZN(_AES_ENC_u0_N266 ) );
NAND2_X2 _AES_ENC_u0_U136  ( .A1(_AES_ENC_u0_N212 ), .A2(_AES_ENC_u0_n323 ),.ZN(_AES_ENC_u0_n990 ) );
NAND2_X2 _AES_ENC_u0_U135  ( .A1(_AES_ENC_u0_n980 ), .A2(_AES_ENC_u0_n990 ),.ZN(_AES_ENC_u0_N267 ) );
NAND2_X2 _AES_ENC_u0_U133  ( .A1(_AES_ENC_u0_N211 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n970 ) );
NAND2_X2 _AES_ENC_u0_U132  ( .A1(_AES_ENC_u0_n960 ), .A2(_AES_ENC_u0_n970 ),.ZN(_AES_ENC_u0_N268 ) );
NAND2_X2 _AES_ENC_u0_U130  ( .A1(_AES_ENC_u0_N210 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n950 ) );
NAND2_X2 _AES_ENC_u0_U129  ( .A1(_AES_ENC_u0_n940 ), .A2(_AES_ENC_u0_n950 ),.ZN(_AES_ENC_u0_N269 ) );
NAND2_X2 _AES_ENC_u0_U127  ( .A1(_AES_ENC_u0_N209 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n930 ) );
NAND2_X2 _AES_ENC_u0_U126  ( .A1(_AES_ENC_u0_n920 ), .A2(_AES_ENC_u0_n930 ),.ZN(_AES_ENC_u0_N270 ) );
NAND2_X2 _AES_ENC_u0_U124  ( .A1(_AES_ENC_u0_N208 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n910 ) );
NAND2_X2 _AES_ENC_u0_U123  ( .A1(_AES_ENC_u0_n900 ), .A2(_AES_ENC_u0_n910 ),.ZN(_AES_ENC_u0_N271 ) );
XOR2_X2 _AES_ENC_u0_U121  ( .A(_AES_ENC_w0[0] ), .B(_AES_ENC_u0_subword[0] ),.Z(_AES_ENC_u0_n890 ) );
NAND2_X2 _AES_ENC_u0_U120  ( .A1(_AES_ENC_u0_n890 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n880 ) );
NAND2_X2 _AES_ENC_u0_U119  ( .A1(_AES_ENC_u0_n870 ), .A2(_AES_ENC_u0_n880 ),.ZN(_AES_ENC_u0_N42 ) );
XOR2_X2 _AES_ENC_u0_U117  ( .A(_AES_ENC_w0[1] ), .B(_AES_ENC_u0_subword[1] ),.Z(_AES_ENC_u0_n860 ) );
NAND2_X2 _AES_ENC_u0_U116  ( .A1(_AES_ENC_u0_n860 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n850 ) );
NAND2_X2 _AES_ENC_u0_U115  ( .A1(_AES_ENC_u0_n840 ), .A2(_AES_ENC_u0_n850 ),.ZN(_AES_ENC_u0_N43 ) );
XOR2_X2 _AES_ENC_u0_U113  ( .A(_AES_ENC_w0[2] ), .B(_AES_ENC_u0_subword[2] ),.Z(_AES_ENC_u0_n830 ) );
NAND2_X2 _AES_ENC_u0_U112  ( .A1(_AES_ENC_u0_n830 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n820 ) );
NAND2_X2 _AES_ENC_u0_U111  ( .A1(_AES_ENC_u0_n810 ), .A2(_AES_ENC_u0_n820 ),.ZN(_AES_ENC_u0_N44 ) );
XOR2_X2 _AES_ENC_u0_U109  ( .A(_AES_ENC_w0[3] ), .B(_AES_ENC_u0_subword[3] ),.Z(_AES_ENC_u0_n800 ) );
NAND2_X2 _AES_ENC_u0_U108  ( .A1(_AES_ENC_u0_n800 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n790 ) );
NAND2_X2 _AES_ENC_u0_U107  ( .A1(_AES_ENC_u0_n780 ), .A2(_AES_ENC_u0_n790 ),.ZN(_AES_ENC_u0_N45 ) );
XOR2_X2 _AES_ENC_u0_U105  ( .A(_AES_ENC_w0[4] ), .B(_AES_ENC_u0_subword[4] ),.Z(_AES_ENC_u0_n770 ) );
NAND2_X2 _AES_ENC_u0_U104  ( .A1(_AES_ENC_u0_n770 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n760 ) );
NAND2_X2 _AES_ENC_u0_U103  ( .A1(_AES_ENC_u0_n75 ), .A2(_AES_ENC_u0_n760 ),.ZN(_AES_ENC_u0_N46 ) );
XOR2_X2 _AES_ENC_u0_U101  ( .A(_AES_ENC_w0[5] ), .B(_AES_ENC_u0_subword[5] ),.Z(_AES_ENC_u0_n74 ) );
NAND2_X2 _AES_ENC_u0_U100  ( .A1(_AES_ENC_u0_n74 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n730 ) );
NAND2_X2 _AES_ENC_u0_U99  ( .A1(_AES_ENC_u0_n720 ), .A2(_AES_ENC_u0_n730 ),.ZN(_AES_ENC_u0_N47 ) );
XOR2_X2 _AES_ENC_u0_U97  ( .A(_AES_ENC_w0[6] ), .B(_AES_ENC_u0_subword[6] ),.Z(_AES_ENC_u0_n710 ) );
NAND2_X2 _AES_ENC_u0_U96  ( .A1(_AES_ENC_u0_n710 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n700 ) );
NAND2_X2 _AES_ENC_u0_U95  ( .A1(_AES_ENC_u0_n690 ), .A2(_AES_ENC_u0_n700 ),.ZN(_AES_ENC_u0_N48 ) );
XOR2_X2 _AES_ENC_u0_U93  ( .A(_AES_ENC_w0[7] ), .B(_AES_ENC_u0_subword[7] ),.Z(_AES_ENC_u0_n680 ) );
NAND2_X2 _AES_ENC_u0_U92  ( .A1(_AES_ENC_u0_n680 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n670 ) );
NAND2_X2 _AES_ENC_u0_U91  ( .A1(_AES_ENC_u0_n660 ), .A2(_AES_ENC_u0_n670 ),.ZN(_AES_ENC_u0_N49 ) );
XOR2_X2 _AES_ENC_u0_U89  ( .A(_AES_ENC_w0[8] ), .B(_AES_ENC_u0_subword[8] ),.Z(_AES_ENC_u0_n650 ) );
NAND2_X2 _AES_ENC_u0_U88  ( .A1(_AES_ENC_u0_n650 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n640 ) );
NAND2_X2 _AES_ENC_u0_U87  ( .A1(_AES_ENC_u0_n630 ), .A2(_AES_ENC_u0_n640 ),.ZN(_AES_ENC_u0_N50 ) );
XOR2_X2 _AES_ENC_u0_U85  ( .A(_AES_ENC_w0[9] ), .B(_AES_ENC_u0_subword[9] ),.Z(_AES_ENC_u0_n620 ) );
NAND2_X2 _AES_ENC_u0_U84  ( .A1(_AES_ENC_u0_n620 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n610 ) );
NAND2_X2 _AES_ENC_u0_U83  ( .A1(_AES_ENC_u0_n600 ), .A2(_AES_ENC_u0_n610 ),.ZN(_AES_ENC_u0_N51 ) );
XOR2_X2 _AES_ENC_u0_U81  ( .A(_AES_ENC_w0[10] ), .B(_AES_ENC_u0_subword[10] ), .Z(_AES_ENC_u0_n590 ) );
NAND2_X2 _AES_ENC_u0_U80  ( .A1(_AES_ENC_u0_n590 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n580 ) );
NAND2_X2 _AES_ENC_u0_U79  ( .A1(_AES_ENC_u0_n570 ), .A2(_AES_ENC_u0_n580 ),.ZN(_AES_ENC_u0_N52 ) );
XOR2_X2 _AES_ENC_u0_U77  ( .A(_AES_ENC_w0[11] ), .B(_AES_ENC_u0_subword[11] ), .Z(_AES_ENC_u0_n560 ) );
NAND2_X2 _AES_ENC_u0_U76  ( .A1(_AES_ENC_u0_n560 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n550 ) );
NAND2_X2 _AES_ENC_u0_U75  ( .A1(_AES_ENC_u0_n540 ), .A2(_AES_ENC_u0_n550 ),.ZN(_AES_ENC_u0_N53 ) );
XOR2_X2 _AES_ENC_u0_U73  ( .A(_AES_ENC_w0[12] ), .B(_AES_ENC_u0_subword[12] ), .Z(_AES_ENC_u0_n530 ) );
NAND2_X2 _AES_ENC_u0_U72  ( .A1(_AES_ENC_u0_n530 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n520 ) );
NAND2_X2 _AES_ENC_u0_U71  ( .A1(_AES_ENC_u0_n510 ), .A2(_AES_ENC_u0_n520 ),.ZN(_AES_ENC_u0_N54 ) );
XOR2_X2 _AES_ENC_u0_U69  ( .A(_AES_ENC_w0[13] ), .B(_AES_ENC_u0_subword[13] ), .Z(_AES_ENC_u0_n500 ) );
NAND2_X2 _AES_ENC_u0_U68  ( .A1(_AES_ENC_u0_n500 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n490 ) );
NAND2_X2 _AES_ENC_u0_U67  ( .A1(_AES_ENC_u0_n480 ), .A2(_AES_ENC_u0_n490 ),.ZN(_AES_ENC_u0_N55 ) );
XOR2_X2 _AES_ENC_u0_U65  ( .A(_AES_ENC_w0[14] ), .B(_AES_ENC_u0_subword[14] ), .Z(_AES_ENC_u0_n470 ) );
NAND2_X2 _AES_ENC_u0_U64  ( .A1(_AES_ENC_u0_n470 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n460 ) );
NAND2_X2 _AES_ENC_u0_U63  ( .A1(_AES_ENC_u0_n450 ), .A2(_AES_ENC_u0_n460 ),.ZN(_AES_ENC_u0_N56 ) );
XOR2_X2 _AES_ENC_u0_U61  ( .A(_AES_ENC_w0[15] ), .B(_AES_ENC_u0_subword[15] ), .Z(_AES_ENC_u0_n440 ) );
NAND2_X2 _AES_ENC_u0_U60  ( .A1(_AES_ENC_u0_n440 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n430 ) );
NAND2_X2 _AES_ENC_u0_U59  ( .A1(_AES_ENC_u0_n420 ), .A2(_AES_ENC_u0_n430 ),.ZN(_AES_ENC_u0_N57 ) );
XOR2_X2 _AES_ENC_u0_U57  ( .A(_AES_ENC_w0[16] ), .B(_AES_ENC_u0_subword[16] ), .Z(_AES_ENC_u0_n41 ) );
NAND2_X2 _AES_ENC_u0_U56  ( .A1(_AES_ENC_u0_n41 ), .A2(_AES_ENC_u0_n324 ),.ZN(_AES_ENC_u0_n40 ) );
NAND2_X2 _AES_ENC_u0_U55  ( .A1(_AES_ENC_u0_n39 ), .A2(_AES_ENC_u0_n40 ),.ZN(_AES_ENC_u0_N58 ) );
XOR2_X2 _AES_ENC_u0_U53  ( .A(_AES_ENC_w0[17] ), .B(_AES_ENC_u0_subword[17] ), .Z(_AES_ENC_u0_n38 ) );
NAND2_X2 _AES_ENC_u0_U52  ( .A1(_AES_ENC_u0_n38 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n37 ) );
NAND2_X2 _AES_ENC_u0_U51  ( .A1(_AES_ENC_u0_n36 ), .A2(_AES_ENC_u0_n37 ),.ZN(_AES_ENC_u0_N59 ) );
XOR2_X2 _AES_ENC_u0_U49  ( .A(_AES_ENC_w0[18] ), .B(_AES_ENC_u0_subword[18] ), .Z(_AES_ENC_u0_n35 ) );
NAND2_X2 _AES_ENC_u0_U48  ( .A1(_AES_ENC_u0_n35 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n34 ) );
NAND2_X2 _AES_ENC_u0_U47  ( .A1(_AES_ENC_u0_n33 ), .A2(_AES_ENC_u0_n34 ),.ZN(_AES_ENC_u0_N60 ) );
XOR2_X2 _AES_ENC_u0_U45  ( .A(_AES_ENC_w0[19] ), .B(_AES_ENC_u0_subword[19] ), .Z(_AES_ENC_u0_n32 ) );
NAND2_X2 _AES_ENC_u0_U44  ( .A1(_AES_ENC_u0_n32 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n31 ) );
NAND2_X2 _AES_ENC_u0_U43  ( .A1(_AES_ENC_u0_n30 ), .A2(_AES_ENC_u0_n31 ),.ZN(_AES_ENC_u0_N61 ) );
XOR2_X2 _AES_ENC_u0_U41  ( .A(_AES_ENC_w0[20] ), .B(_AES_ENC_u0_subword[20] ), .Z(_AES_ENC_u0_n29 ) );
NAND2_X2 _AES_ENC_u0_U40  ( .A1(_AES_ENC_u0_n29 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n28 ) );
NAND2_X2 _AES_ENC_u0_U39  ( .A1(_AES_ENC_u0_n27 ), .A2(_AES_ENC_u0_n28 ),.ZN(_AES_ENC_u0_N62 ) );
XOR2_X2 _AES_ENC_u0_U37  ( .A(_AES_ENC_w0[21] ), .B(_AES_ENC_u0_subword[21] ), .Z(_AES_ENC_u0_n26 ) );
NAND2_X2 _AES_ENC_u0_U36  ( .A1(_AES_ENC_u0_n26 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n25 ) );
NAND2_X2 _AES_ENC_u0_U35  ( .A1(_AES_ENC_u0_n24 ), .A2(_AES_ENC_u0_n25 ),.ZN(_AES_ENC_u0_N63 ) );
XOR2_X2 _AES_ENC_u0_U33  ( .A(_AES_ENC_w0[22] ), .B(_AES_ENC_u0_subword[22] ), .Z(_AES_ENC_u0_n23 ) );
NAND2_X2 _AES_ENC_u0_U32  ( .A1(_AES_ENC_u0_n23 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n22 ) );
NAND2_X2 _AES_ENC_u0_U31  ( .A1(_AES_ENC_u0_n21 ), .A2(_AES_ENC_u0_n22 ),.ZN(_AES_ENC_u0_N64 ) );
XOR2_X2 _AES_ENC_u0_U29  ( .A(_AES_ENC_w0[23] ), .B(_AES_ENC_u0_subword[23] ), .Z(_AES_ENC_u0_n20 ) );
NAND2_X2 _AES_ENC_u0_U28  ( .A1(_AES_ENC_u0_n20 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n19 ) );
NAND2_X2 _AES_ENC_u0_U27  ( .A1(_AES_ENC_u0_n18 ), .A2(_AES_ENC_u0_n19 ),.ZN(_AES_ENC_u0_N65 ) );
NAND2_X2 _AES_ENC_u0_U25  ( .A1(_AES_ENC_u0_N17 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n1710 ) );
NAND2_X2 _AES_ENC_u0_U24  ( .A1(_AES_ENC_u0_n1610 ), .A2(_AES_ENC_u0_n1710 ),.ZN(_AES_ENC_u0_N66 ) );
NAND2_X2 _AES_ENC_u0_U22  ( .A1(_AES_ENC_u0_N16 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n1510 ) );
NAND2_X2 _AES_ENC_u0_U21  ( .A1(_AES_ENC_u0_n1400 ), .A2(_AES_ENC_u0_n1510 ),.ZN(_AES_ENC_u0_N67 ) );
NAND2_X2 _AES_ENC_u0_U19  ( .A1(_AES_ENC_u0_N15 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n1310 ) );
NAND2_X2 _AES_ENC_u0_U18  ( .A1(_AES_ENC_u0_n1210 ), .A2(_AES_ENC_u0_n1310 ),.ZN(_AES_ENC_u0_N68 ) );
NAND2_X2 _AES_ENC_u0_U16  ( .A1(_AES_ENC_u0_N14 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n1110 ) );
NAND2_X2 _AES_ENC_u0_U15  ( .A1(_AES_ENC_u0_n1010 ), .A2(_AES_ENC_u0_n1110 ),.ZN(_AES_ENC_u0_N69 ) );
NAND2_X2 _AES_ENC_u0_U13  ( .A1(_AES_ENC_u0_N13 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n9 ) );
NAND2_X2 _AES_ENC_u0_U12  ( .A1(_AES_ENC_u0_n8 ), .A2(_AES_ENC_u0_n9 ), .ZN(_AES_ENC_u0_N70 ) );
NAND2_X2 _AES_ENC_u0_U10  ( .A1(_AES_ENC_u0_N12 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n7 ) );
NAND2_X2 _AES_ENC_u0_U9  ( .A1(_AES_ENC_u0_n6 ), .A2(_AES_ENC_u0_n7 ), .ZN(_AES_ENC_u0_N71 ) );
NAND2_X2 _AES_ENC_u0_U7  ( .A1(_AES_ENC_u0_N11 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n5 ) );
NAND2_X2 _AES_ENC_u0_U6  ( .A1(_AES_ENC_u0_n4 ), .A2(_AES_ENC_u0_n5 ), .ZN(_AES_ENC_u0_N72 ) );
NAND2_X2 _AES_ENC_u0_U4  ( .A1(_AES_ENC_u0_N10 ), .A2(_AES_ENC_u0_n325 ),.ZN(_AES_ENC_u0_n3 ) );
CLKBUFX1 gbuf_d_1166(.A(_AES_ENC_u0_N108), .Y(ddout__1166));
CLKBUFX1 gbuf_q_1166(.A(qq_in1166), .Y(_AES_ENC_w1[0]));
CLKBUFX1 gbuf_d_1167(.A(_AES_ENC_u0_N174), .Y(ddout__1167));
CLKBUFX1 gbuf_q_1167(.A(qq_in1167), .Y(_AES_ENC_w2[0]));
CLKBUFX1 gbuf_d_1168(.A(_AES_ENC_u0_N123), .Y(ddout__1168));
CLKBUFX1 gbuf_q_1168(.A(qq_in1168), .Y(_AES_ENC_w1[15]));
CLKBUFX1 gbuf_d_1169(.A(_AES_ENC_u0_N189), .Y(ddout__1169));
CLKBUFX1 gbuf_q_1169(.A(qq_in1169), .Y(_AES_ENC_w2[15]));
CLKBUFX1 gbuf_d_1170(.A(_AES_ENC_u0_N131), .Y(ddout__1170));
CLKBUFX1 gbuf_q_1170(.A(qq_in1170), .Y(_AES_ENC_w1[23]));
CLKBUFX1 gbuf_d_1171(.A(_AES_ENC_u0_N197), .Y(ddout__1171));
CLKBUFX1 gbuf_q_1171(.A(qq_in1171), .Y(_AES_ENC_w2[23]));
CLKBUFX1 gbuf_d_1172(.A(_AES_ENC_u0_n314), .Y(ddout__1172));
CLKBUFX1 gbuf_q_1172(.A(qq_in1172), .Y(_AES_ENC_w0[31]));
CLKBUFX1 gbuf_d_1173(.A(_AES_ENC_u0_N139), .Y(ddout__1173));
CLKBUFX1 gbuf_q_1173(.A(qq_in1173), .Y(_AES_ENC_w1[31]));
CLKBUFX1 gbuf_d_1174(.A(_AES_ENC_u0_N205), .Y(ddout__1174));
CLKBUFX1 gbuf_q_1174(.A(qq_in1174), .Y(_AES_ENC_w2[31]));
CLKBUFX1 gbuf_d_1175(.A(_AES_ENC_u0_N115), .Y(ddout__1175));
CLKBUFX1 gbuf_q_1175(.A(qq_in1175), .Y(_AES_ENC_w1[7]));
CLKBUFX1 gbuf_d_1176(.A(_AES_ENC_u0_N181), .Y(ddout__1176));
CLKBUFX1 gbuf_q_1176(.A(qq_in1176), .Y(_AES_ENC_w2[7]));
CLKBUFX1 gbuf_d_1177(.A(_AES_ENC_u0_N247), .Y(ddout__1177));
CLKBUFX1 gbuf_q_1177(.A(qq_in1177), .Y(_AES_ENC_w3[7]));
CLKBUFX1 gbuf_d_1178(.A(_AES_ENC_u0_N49), .Y(ddout__1178));
CLKBUFX1 gbuf_q_1178(.A(qq_in1178), .Y(_AES_ENC_w0[7]));
CLKBUFX1 gbuf_d_1179(.A(_AES_ENC_u0_N114), .Y(ddout__1179));
CLKBUFX1 gbuf_q_1179(.A(qq_in1179), .Y(_AES_ENC_w1[6]));
CLKBUFX1 gbuf_d_1180(.A(_AES_ENC_u0_N180), .Y(ddout__1180));
CLKBUFX1 gbuf_q_1180(.A(qq_in1180), .Y(_AES_ENC_w2[6]));
CLKBUFX1 gbuf_d_1181(.A(_AES_ENC_u0_N246), .Y(ddout__1181));
CLKBUFX1 gbuf_q_1181(.A(qq_in1181), .Y(_AES_ENC_w3[6]));
CLKBUFX1 gbuf_d_1182(.A(_AES_ENC_u0_N48), .Y(ddout__1182));
CLKBUFX1 gbuf_q_1182(.A(qq_in1182), .Y(_AES_ENC_w0[6]));
CLKBUFX1 gbuf_d_1183(.A(_AES_ENC_u0_N113), .Y(ddout__1183));
CLKBUFX1 gbuf_q_1183(.A(qq_in1183), .Y(_AES_ENC_w1[5]));
CLKBUFX1 gbuf_d_1184(.A(_AES_ENC_u0_N179), .Y(ddout__1184));
CLKBUFX1 gbuf_q_1184(.A(qq_in1184), .Y(_AES_ENC_w2[5]));
CLKBUFX1 gbuf_d_1185(.A(_AES_ENC_u0_N245), .Y(ddout__1185));
CLKBUFX1 gbuf_q_1185(.A(qq_in1185), .Y(_AES_ENC_w3[5]));
CLKBUFX1 gbuf_d_1186(.A(_AES_ENC_u0_N47), .Y(ddout__1186));
CLKBUFX1 gbuf_q_1186(.A(qq_in1186), .Y(_AES_ENC_w0[5]));
CLKBUFX1 gbuf_d_1187(.A(_AES_ENC_u0_N112), .Y(ddout__1187));
CLKBUFX1 gbuf_q_1187(.A(qq_in1187), .Y(_AES_ENC_w1[4]));
CLKBUFX1 gbuf_d_1188(.A(_AES_ENC_u0_N178), .Y(ddout__1188));
CLKBUFX1 gbuf_q_1188(.A(qq_in1188), .Y(_AES_ENC_w2[4]));
CLKBUFX1 gbuf_d_1189(.A(_AES_ENC_u0_N244), .Y(ddout__1189));
CLKBUFX1 gbuf_q_1189(.A(qq_in1189), .Y(_AES_ENC_w3[4]));
CLKBUFX1 gbuf_d_1190(.A(_AES_ENC_u0_N46), .Y(ddout__1190));
CLKBUFX1 gbuf_q_1190(.A(qq_in1190), .Y(_AES_ENC_w0[4]));
CLKBUFX1 gbuf_d_1191(.A(_AES_ENC_u0_N111), .Y(ddout__1191));
CLKBUFX1 gbuf_q_1191(.A(qq_in1191), .Y(_AES_ENC_w1[3]));
CLKBUFX1 gbuf_d_1192(.A(_AES_ENC_u0_N177), .Y(ddout__1192));
CLKBUFX1 gbuf_q_1192(.A(qq_in1192), .Y(_AES_ENC_w2[3]));
CLKBUFX1 gbuf_d_1193(.A(_AES_ENC_u0_N243), .Y(ddout__1193));
CLKBUFX1 gbuf_q_1193(.A(qq_in1193), .Y(_AES_ENC_w3[3]));
CLKBUFX1 gbuf_d_1194(.A(_AES_ENC_u0_N45), .Y(ddout__1194));
CLKBUFX1 gbuf_q_1194(.A(qq_in1194), .Y(_AES_ENC_w0[3]));
CLKBUFX1 gbuf_d_1195(.A(_AES_ENC_u0_N110), .Y(ddout__1195));
CLKBUFX1 gbuf_q_1195(.A(qq_in1195), .Y(_AES_ENC_w1[2]));
CLKBUFX1 gbuf_d_1196(.A(_AES_ENC_u0_N176), .Y(ddout__1196));
CLKBUFX1 gbuf_q_1196(.A(qq_in1196), .Y(_AES_ENC_w2[2]));
CLKBUFX1 gbuf_d_1197(.A(_AES_ENC_u0_N242), .Y(ddout__1197));
CLKBUFX1 gbuf_q_1197(.A(qq_in1197), .Y(_AES_ENC_w3[2]));
CLKBUFX1 gbuf_d_1198(.A(_AES_ENC_u0_N44), .Y(ddout__1198));
CLKBUFX1 gbuf_q_1198(.A(qq_in1198), .Y(_AES_ENC_w0[2]));
CLKBUFX1 gbuf_d_1199(.A(_AES_ENC_u0_N109), .Y(ddout__1199));
CLKBUFX1 gbuf_q_1199(.A(qq_in1199), .Y(_AES_ENC_w1[1]));
CLKBUFX1 gbuf_d_1200(.A(_AES_ENC_u0_N175), .Y(ddout__1200));
CLKBUFX1 gbuf_q_1200(.A(qq_in1200), .Y(_AES_ENC_w2[1]));
CLKBUFX1 gbuf_d_1201(.A(_AES_ENC_u0_N241), .Y(ddout__1201));
CLKBUFX1 gbuf_q_1201(.A(qq_in1201), .Y(_AES_ENC_w3[1]));
CLKBUFX1 gbuf_d_1202(.A(_AES_ENC_u0_N43), .Y(ddout__1202));
CLKBUFX1 gbuf_q_1202(.A(qq_in1202), .Y(_AES_ENC_w0[1]));
CLKBUFX1 gbuf_d_1203(.A(_AES_ENC_u0_N271), .Y(ddout__1203));
CLKBUFX1 gbuf_q_1203(.A(qq_in1203), .Y(_AES_ENC_w3[31]));
CLKBUFX1 gbuf_d_1204(.A(_AES_ENC_u0_N72), .Y(ddout__1204));
CLKBUFX1 gbuf_q_1204(.A(qq_in1204), .Y(_AES_ENC_w0[30]));
CLKBUFX1 gbuf_d_1205(.A(_AES_ENC_u0_N138), .Y(ddout__1205));
CLKBUFX1 gbuf_q_1205(.A(qq_in1205), .Y(_AES_ENC_w1[30]));
CLKBUFX1 gbuf_d_1206(.A(_AES_ENC_u0_N204), .Y(ddout__1206));
CLKBUFX1 gbuf_q_1206(.A(qq_in1206), .Y(_AES_ENC_w2[30]));
CLKBUFX1 gbuf_d_1207(.A(_AES_ENC_u0_N270), .Y(ddout__1207));
CLKBUFX1 gbuf_q_1207(.A(qq_in1207), .Y(_AES_ENC_w3[30]));
CLKBUFX1 gbuf_d_1208(.A(_AES_ENC_u0_N71), .Y(ddout__1208));
CLKBUFX1 gbuf_q_1208(.A(qq_in1208), .Y(_AES_ENC_w0[29]));
CLKBUFX1 gbuf_d_1209(.A(_AES_ENC_u0_N137), .Y(ddout__1209));
CLKBUFX1 gbuf_q_1209(.A(qq_in1209), .Y(_AES_ENC_w1[29]));
CLKBUFX1 gbuf_d_1210(.A(_AES_ENC_u0_N203), .Y(ddout__1210));
CLKBUFX1 gbuf_q_1210(.A(qq_in1210), .Y(_AES_ENC_w2[29]));
CLKBUFX1 gbuf_d_1211(.A(_AES_ENC_u0_N269), .Y(ddout__1211));
CLKBUFX1 gbuf_q_1211(.A(qq_in1211), .Y(_AES_ENC_w3[29]));
CLKBUFX1 gbuf_d_1212(.A(_AES_ENC_u0_N70), .Y(ddout__1212));
CLKBUFX1 gbuf_q_1212(.A(qq_in1212), .Y(_AES_ENC_w0[28]));
CLKBUFX1 gbuf_d_1213(.A(_AES_ENC_u0_N136), .Y(ddout__1213));
CLKBUFX1 gbuf_q_1213(.A(qq_in1213), .Y(_AES_ENC_w1[28]));
CLKBUFX1 gbuf_d_1214(.A(_AES_ENC_u0_N202), .Y(ddout__1214));
CLKBUFX1 gbuf_q_1214(.A(qq_in1214), .Y(_AES_ENC_w2[28]));
CLKBUFX1 gbuf_d_1215(.A(_AES_ENC_u0_N268), .Y(ddout__1215));
CLKBUFX1 gbuf_q_1215(.A(qq_in1215), .Y(_AES_ENC_w3[28]));
CLKBUFX1 gbuf_d_1216(.A(_AES_ENC_u0_N69), .Y(ddout__1216));
CLKBUFX1 gbuf_q_1216(.A(qq_in1216), .Y(_AES_ENC_w0[27]));
CLKBUFX1 gbuf_d_1217(.A(_AES_ENC_u0_N135), .Y(ddout__1217));
CLKBUFX1 gbuf_q_1217(.A(qq_in1217), .Y(_AES_ENC_w1[27]));
CLKBUFX1 gbuf_d_1218(.A(_AES_ENC_u0_N201), .Y(ddout__1218));
CLKBUFX1 gbuf_q_1218(.A(qq_in1218), .Y(_AES_ENC_w2[27]));
CLKBUFX1 gbuf_d_1219(.A(_AES_ENC_u0_N267), .Y(ddout__1219));
CLKBUFX1 gbuf_q_1219(.A(qq_in1219), .Y(_AES_ENC_w3[27]));
CLKBUFX1 gbuf_d_1220(.A(_AES_ENC_u0_N68), .Y(ddout__1220));
CLKBUFX1 gbuf_q_1220(.A(qq_in1220), .Y(_AES_ENC_w0[26]));
CLKBUFX1 gbuf_d_1221(.A(_AES_ENC_u0_N134), .Y(ddout__1221));
CLKBUFX1 gbuf_q_1221(.A(qq_in1221), .Y(_AES_ENC_w1[26]));
CLKBUFX1 gbuf_d_1222(.A(_AES_ENC_u0_N200), .Y(ddout__1222));
CLKBUFX1 gbuf_q_1222(.A(qq_in1222), .Y(_AES_ENC_w2[26]));
CLKBUFX1 gbuf_d_1223(.A(_AES_ENC_u0_N266), .Y(ddout__1223));
CLKBUFX1 gbuf_q_1223(.A(qq_in1223), .Y(_AES_ENC_w3[26]));
CLKBUFX1 gbuf_d_1224(.A(_AES_ENC_u0_N67), .Y(ddout__1224));
CLKBUFX1 gbuf_q_1224(.A(qq_in1224), .Y(_AES_ENC_w0[25]));
CLKBUFX1 gbuf_d_1225(.A(_AES_ENC_u0_N133), .Y(ddout__1225));
CLKBUFX1 gbuf_q_1225(.A(qq_in1225), .Y(_AES_ENC_w1[25]));
CLKBUFX1 gbuf_d_1226(.A(_AES_ENC_u0_N199), .Y(ddout__1226));
CLKBUFX1 gbuf_q_1226(.A(qq_in1226), .Y(_AES_ENC_w2[25]));
CLKBUFX1 gbuf_d_1227(.A(_AES_ENC_u0_N265), .Y(ddout__1227));
CLKBUFX1 gbuf_q_1227(.A(qq_in1227), .Y(_AES_ENC_w3[25]));
CLKBUFX1 gbuf_d_1228(.A(_AES_ENC_u0_N66), .Y(ddout__1228));
CLKBUFX1 gbuf_q_1228(.A(qq_in1228), .Y(_AES_ENC_w0[24]));
CLKBUFX1 gbuf_d_1229(.A(_AES_ENC_u0_N132), .Y(ddout__1229));
CLKBUFX1 gbuf_q_1229(.A(qq_in1229), .Y(_AES_ENC_w1[24]));
CLKBUFX1 gbuf_d_1230(.A(_AES_ENC_u0_N198), .Y(ddout__1230));
CLKBUFX1 gbuf_q_1230(.A(qq_in1230), .Y(_AES_ENC_w2[24]));
CLKBUFX1 gbuf_d_1231(.A(_AES_ENC_u0_N264), .Y(ddout__1231));
CLKBUFX1 gbuf_q_1231(.A(qq_in1231), .Y(_AES_ENC_w3[24]));
CLKBUFX1 gbuf_d_1232(.A(_AES_ENC_u0_N263), .Y(ddout__1232));
CLKBUFX1 gbuf_q_1232(.A(qq_in1232), .Y(_AES_ENC_w3[23]));
CLKBUFX1 gbuf_d_1233(.A(_AES_ENC_u0_N65), .Y(ddout__1233));
CLKBUFX1 gbuf_q_1233(.A(qq_in1233), .Y(_AES_ENC_w0[23]));
CLKBUFX1 gbuf_d_1234(.A(_AES_ENC_u0_N130), .Y(ddout__1234));
CLKBUFX1 gbuf_q_1234(.A(qq_in1234), .Y(_AES_ENC_w1[22]));
CLKBUFX1 gbuf_d_1235(.A(_AES_ENC_u0_N196), .Y(ddout__1235));
CLKBUFX1 gbuf_q_1235(.A(qq_in1235), .Y(_AES_ENC_w2[22]));
CLKBUFX1 gbuf_d_1236(.A(_AES_ENC_u0_N262), .Y(ddout__1236));
CLKBUFX1 gbuf_q_1236(.A(qq_in1236), .Y(_AES_ENC_w3[22]));
CLKBUFX1 gbuf_d_1237(.A(_AES_ENC_u0_N64), .Y(ddout__1237));
CLKBUFX1 gbuf_q_1237(.A(qq_in1237), .Y(_AES_ENC_w0[22]));
CLKBUFX1 gbuf_d_1238(.A(_AES_ENC_u0_N129), .Y(ddout__1238));
CLKBUFX1 gbuf_q_1238(.A(qq_in1238), .Y(_AES_ENC_w1[21]));
CLKBUFX1 gbuf_d_1239(.A(_AES_ENC_u0_N195), .Y(ddout__1239));
CLKBUFX1 gbuf_q_1239(.A(qq_in1239), .Y(_AES_ENC_w2[21]));
CLKBUFX1 gbuf_d_1240(.A(_AES_ENC_u0_N261), .Y(ddout__1240));
CLKBUFX1 gbuf_q_1240(.A(qq_in1240), .Y(_AES_ENC_w3[21]));
CLKBUFX1 gbuf_d_1241(.A(_AES_ENC_u0_N63), .Y(ddout__1241));
CLKBUFX1 gbuf_q_1241(.A(qq_in1241), .Y(_AES_ENC_w0[21]));
CLKBUFX1 gbuf_d_1242(.A(_AES_ENC_u0_N128), .Y(ddout__1242));
CLKBUFX1 gbuf_q_1242(.A(qq_in1242), .Y(_AES_ENC_w1[20]));
CLKBUFX1 gbuf_d_1243(.A(_AES_ENC_u0_N194), .Y(ddout__1243));
CLKBUFX1 gbuf_q_1243(.A(qq_in1243), .Y(_AES_ENC_w2[20]));
CLKBUFX1 gbuf_d_1244(.A(_AES_ENC_u0_N260), .Y(ddout__1244));
CLKBUFX1 gbuf_q_1244(.A(qq_in1244), .Y(_AES_ENC_w3[20]));
CLKBUFX1 gbuf_d_1245(.A(_AES_ENC_u0_N62), .Y(ddout__1245));
CLKBUFX1 gbuf_q_1245(.A(qq_in1245), .Y(_AES_ENC_w0[20]));
CLKBUFX1 gbuf_d_1246(.A(_AES_ENC_u0_N127), .Y(ddout__1246));
CLKBUFX1 gbuf_q_1246(.A(qq_in1246), .Y(_AES_ENC_w1[19]));
CLKBUFX1 gbuf_d_1247(.A(_AES_ENC_u0_N193), .Y(ddout__1247));
CLKBUFX1 gbuf_q_1247(.A(qq_in1247), .Y(_AES_ENC_w2[19]));
CLKBUFX1 gbuf_d_1248(.A(_AES_ENC_u0_N259), .Y(ddout__1248));
CLKBUFX1 gbuf_q_1248(.A(qq_in1248), .Y(_AES_ENC_w3[19]));
CLKBUFX1 gbuf_d_1249(.A(_AES_ENC_u0_N61), .Y(ddout__1249));
CLKBUFX1 gbuf_q_1249(.A(qq_in1249), .Y(_AES_ENC_w0[19]));
CLKBUFX1 gbuf_d_1250(.A(_AES_ENC_u0_N126), .Y(ddout__1250));
CLKBUFX1 gbuf_q_1250(.A(qq_in1250), .Y(_AES_ENC_w1[18]));
CLKBUFX1 gbuf_d_1251(.A(_AES_ENC_u0_N192), .Y(ddout__1251));
CLKBUFX1 gbuf_q_1251(.A(qq_in1251), .Y(_AES_ENC_w2[18]));
CLKBUFX1 gbuf_d_1252(.A(_AES_ENC_u0_N258), .Y(ddout__1252));
CLKBUFX1 gbuf_q_1252(.A(qq_in1252), .Y(_AES_ENC_w3[18]));
CLKBUFX1 gbuf_d_1253(.A(_AES_ENC_u0_N60), .Y(ddout__1253));
CLKBUFX1 gbuf_q_1253(.A(qq_in1253), .Y(_AES_ENC_w0[18]));
CLKBUFX1 gbuf_d_1254(.A(_AES_ENC_u0_N125), .Y(ddout__1254));
CLKBUFX1 gbuf_q_1254(.A(qq_in1254), .Y(_AES_ENC_w1[17]));
CLKBUFX1 gbuf_d_1255(.A(_AES_ENC_u0_N191), .Y(ddout__1255));
CLKBUFX1 gbuf_q_1255(.A(qq_in1255), .Y(_AES_ENC_w2[17]));
CLKBUFX1 gbuf_d_1256(.A(_AES_ENC_u0_N257), .Y(ddout__1256));
CLKBUFX1 gbuf_q_1256(.A(qq_in1256), .Y(_AES_ENC_w3[17]));
CLKBUFX1 gbuf_d_1257(.A(_AES_ENC_u0_N59), .Y(ddout__1257));
CLKBUFX1 gbuf_q_1257(.A(qq_in1257), .Y(_AES_ENC_w0[17]));
CLKBUFX1 gbuf_d_1258(.A(_AES_ENC_u0_N124), .Y(ddout__1258));
CLKBUFX1 gbuf_q_1258(.A(qq_in1258), .Y(_AES_ENC_w1[16]));
CLKBUFX1 gbuf_d_1259(.A(_AES_ENC_u0_N190), .Y(ddout__1259));
CLKBUFX1 gbuf_q_1259(.A(qq_in1259), .Y(_AES_ENC_w2[16]));
CLKBUFX1 gbuf_d_1260(.A(_AES_ENC_u0_N256), .Y(ddout__1260));
CLKBUFX1 gbuf_q_1260(.A(qq_in1260), .Y(_AES_ENC_w3[16]));
CLKBUFX1 gbuf_d_1261(.A(_AES_ENC_u0_N58), .Y(ddout__1261));
CLKBUFX1 gbuf_q_1261(.A(qq_in1261), .Y(_AES_ENC_w0[16]));
CLKBUFX1 gbuf_d_1262(.A(_AES_ENC_u0_N255), .Y(ddout__1262));
CLKBUFX1 gbuf_q_1262(.A(qq_in1262), .Y(_AES_ENC_w3[15]));
CLKBUFX1 gbuf_d_1263(.A(_AES_ENC_u0_N57), .Y(ddout__1263));
CLKBUFX1 gbuf_q_1263(.A(qq_in1263), .Y(_AES_ENC_w0[15]));
CLKBUFX1 gbuf_d_1264(.A(_AES_ENC_u0_N122), .Y(ddout__1264));
CLKBUFX1 gbuf_q_1264(.A(qq_in1264), .Y(_AES_ENC_w1[14]));
CLKBUFX1 gbuf_d_1265(.A(_AES_ENC_u0_N188), .Y(ddout__1265));
CLKBUFX1 gbuf_q_1265(.A(qq_in1265), .Y(_AES_ENC_w2[14]));
CLKBUFX1 gbuf_d_1266(.A(_AES_ENC_u0_N254), .Y(ddout__1266));
CLKBUFX1 gbuf_q_1266(.A(qq_in1266), .Y(_AES_ENC_w3[14]));
CLKBUFX1 gbuf_d_1267(.A(_AES_ENC_u0_N56), .Y(ddout__1267));
CLKBUFX1 gbuf_q_1267(.A(qq_in1267), .Y(_AES_ENC_w0[14]));
CLKBUFX1 gbuf_d_1268(.A(_AES_ENC_u0_N121), .Y(ddout__1268));
CLKBUFX1 gbuf_q_1268(.A(qq_in1268), .Y(_AES_ENC_w1[13]));
CLKBUFX1 gbuf_d_1269(.A(_AES_ENC_u0_N187), .Y(ddout__1269));
CLKBUFX1 gbuf_q_1269(.A(qq_in1269), .Y(_AES_ENC_w2[13]));
CLKBUFX1 gbuf_d_1270(.A(_AES_ENC_u0_N253), .Y(ddout__1270));
CLKBUFX1 gbuf_q_1270(.A(qq_in1270), .Y(_AES_ENC_w3[13]));
CLKBUFX1 gbuf_d_1271(.A(_AES_ENC_u0_N55), .Y(ddout__1271));
CLKBUFX1 gbuf_q_1271(.A(qq_in1271), .Y(_AES_ENC_w0[13]));
CLKBUFX1 gbuf_d_1272(.A(_AES_ENC_u0_N120), .Y(ddout__1272));
CLKBUFX1 gbuf_q_1272(.A(qq_in1272), .Y(_AES_ENC_w1[12]));
CLKBUFX1 gbuf_d_1273(.A(_AES_ENC_u0_N186), .Y(ddout__1273));
CLKBUFX1 gbuf_q_1273(.A(qq_in1273), .Y(_AES_ENC_w2[12]));
CLKBUFX1 gbuf_d_1274(.A(_AES_ENC_u0_N252), .Y(ddout__1274));
CLKBUFX1 gbuf_q_1274(.A(qq_in1274), .Y(_AES_ENC_w3[12]));
CLKBUFX1 gbuf_d_1275(.A(_AES_ENC_u0_N54), .Y(ddout__1275));
CLKBUFX1 gbuf_q_1275(.A(qq_in1275), .Y(_AES_ENC_w0[12]));
CLKBUFX1 gbuf_d_1276(.A(_AES_ENC_u0_N119), .Y(ddout__1276));
CLKBUFX1 gbuf_q_1276(.A(qq_in1276), .Y(_AES_ENC_w1[11]));
CLKBUFX1 gbuf_d_1277(.A(_AES_ENC_u0_N185), .Y(ddout__1277));
CLKBUFX1 gbuf_q_1277(.A(qq_in1277), .Y(_AES_ENC_w2[11]));
CLKBUFX1 gbuf_d_1278(.A(_AES_ENC_u0_N251), .Y(ddout__1278));
CLKBUFX1 gbuf_q_1278(.A(qq_in1278), .Y(_AES_ENC_w3[11]));
CLKBUFX1 gbuf_d_1279(.A(_AES_ENC_u0_N53), .Y(ddout__1279));
CLKBUFX1 gbuf_q_1279(.A(qq_in1279), .Y(_AES_ENC_w0[11]));
CLKBUFX1 gbuf_d_1280(.A(_AES_ENC_u0_N118), .Y(ddout__1280));
CLKBUFX1 gbuf_q_1280(.A(qq_in1280), .Y(_AES_ENC_w1[10]));
CLKBUFX1 gbuf_d_1281(.A(_AES_ENC_u0_N184), .Y(ddout__1281));
CLKBUFX1 gbuf_q_1281(.A(qq_in1281), .Y(_AES_ENC_w2[10]));
CLKBUFX1 gbuf_d_1282(.A(_AES_ENC_u0_N250), .Y(ddout__1282));
CLKBUFX1 gbuf_q_1282(.A(qq_in1282), .Y(_AES_ENC_w3[10]));
CLKBUFX1 gbuf_d_1283(.A(_AES_ENC_u0_N52), .Y(ddout__1283));
CLKBUFX1 gbuf_q_1283(.A(qq_in1283), .Y(_AES_ENC_w0[10]));
CLKBUFX1 gbuf_d_1284(.A(_AES_ENC_u0_N117), .Y(ddout__1284));
CLKBUFX1 gbuf_q_1284(.A(qq_in1284), .Y(_AES_ENC_w1[9]));
CLKBUFX1 gbuf_d_1285(.A(_AES_ENC_u0_N183), .Y(ddout__1285));
CLKBUFX1 gbuf_q_1285(.A(qq_in1285), .Y(_AES_ENC_w2[9]));
CLKBUFX1 gbuf_d_1286(.A(_AES_ENC_u0_N249), .Y(ddout__1286));
CLKBUFX1 gbuf_q_1286(.A(qq_in1286), .Y(_AES_ENC_w3[9]));
CLKBUFX1 gbuf_d_1287(.A(_AES_ENC_u0_N51), .Y(ddout__1287));
CLKBUFX1 gbuf_q_1287(.A(qq_in1287), .Y(_AES_ENC_w0[9]));
CLKBUFX1 gbuf_d_1288(.A(_AES_ENC_u0_N116), .Y(ddout__1288));
CLKBUFX1 gbuf_q_1288(.A(qq_in1288), .Y(_AES_ENC_w1[8]));
CLKBUFX1 gbuf_d_1289(.A(_AES_ENC_u0_N182), .Y(ddout__1289));
CLKBUFX1 gbuf_q_1289(.A(qq_in1289), .Y(_AES_ENC_w2[8]));
CLKBUFX1 gbuf_d_1290(.A(_AES_ENC_u0_N248), .Y(ddout__1290));
CLKBUFX1 gbuf_q_1290(.A(qq_in1290), .Y(_AES_ENC_w3[8]));
CLKBUFX1 gbuf_d_1291(.A(_AES_ENC_u0_N50), .Y(ddout__1291));
CLKBUFX1 gbuf_q_1291(.A(qq_in1291), .Y(_AES_ENC_w0[8]));
CLKBUFX1 gbuf_d_1292(.A(_AES_ENC_u0_N240), .Y(ddout__1292));
CLKBUFX1 gbuf_q_1292(.A(qq_in1292), .Y(_AES_ENC_w3[0]));
CLKBUFX1 gbuf_d_1293(.A(_AES_ENC_u0_N42), .Y(ddout__1293));
CLKBUFX1 gbuf_q_1293(.A(qq_in1293), .Y(_AES_ENC_w0[0]));
XOR2_X2 _AES_ENC_u0_U547  ( .A(_AES_ENC_u0_rcon[31]), .B(_AES_ENC_u0_n282 ),.Z(_AES_ENC_u0_N10 ) );
XOR2_X2 _AES_ENC_u0_U546  ( .A(_AES_ENC_w0[31] ), .B(_AES_ENC_u0_subword[31] ), .Z(_AES_ENC_u0_n282 ) );
XOR2_X2 _AES_ENC_u0_U545  ( .A(_AES_ENC_w1[31] ), .B(_AES_ENC_u0_N10 ), .Z(_AES_ENC_u0_N76 ) );
XOR2_X2 _AES_ENC_u0_U544  ( .A(_AES_ENC_w2[31] ), .B(_AES_ENC_u0_N76 ), .Z(_AES_ENC_u0_N142 ) );
XOR2_X2 _AES_ENC_u0_U543  ( .A(_AES_ENC_w3[31] ), .B(_AES_ENC_u0_N142 ), .Z(_AES_ENC_u0_N208 ) );
XOR2_X2 _AES_ENC_u0_U542  ( .A(_AES_ENC_u0_rcon[30]), .B(_AES_ENC_u0_n283 ),.Z(_AES_ENC_u0_N11 ) );
XOR2_X2 _AES_ENC_u0_U541  ( .A(_AES_ENC_w0[30] ), .B(_AES_ENC_u0_subword[30] ), .Z(_AES_ENC_u0_n283 ) );
XOR2_X2 _AES_ENC_u0_U540  ( .A(_AES_ENC_w1[30] ), .B(_AES_ENC_u0_N11 ), .Z(_AES_ENC_u0_N77 ) );
XOR2_X2 _AES_ENC_u0_U539  ( .A(_AES_ENC_w2[30] ), .B(_AES_ENC_u0_N77 ), .Z(_AES_ENC_u0_N143 ) );
XOR2_X2 _AES_ENC_u0_U538  ( .A(_AES_ENC_w3[30] ), .B(_AES_ENC_u0_N143 ), .Z(_AES_ENC_u0_N209 ) );
XOR2_X2 _AES_ENC_u0_U537  ( .A(_AES_ENC_u0_rcon[29]), .B(_AES_ENC_u0_n284 ),.Z(_AES_ENC_u0_N12 ) );
XOR2_X2 _AES_ENC_u0_U536  ( .A(_AES_ENC_w0[29] ), .B(_AES_ENC_u0_subword[29] ), .Z(_AES_ENC_u0_n284 ) );
XOR2_X2 _AES_ENC_u0_U535  ( .A(_AES_ENC_w1[29] ), .B(_AES_ENC_u0_N12 ), .Z(_AES_ENC_u0_N78 ) );
XOR2_X2 _AES_ENC_u0_U534  ( .A(_AES_ENC_w2[29] ), .B(_AES_ENC_u0_N78 ), .Z(_AES_ENC_u0_N144 ) );
XOR2_X2 _AES_ENC_u0_U533  ( .A(_AES_ENC_w3[29] ), .B(_AES_ENC_u0_N144 ), .Z(_AES_ENC_u0_N210 ) );
XOR2_X2 _AES_ENC_u0_U532  ( .A(_AES_ENC_u0_rcon[28]), .B(_AES_ENC_u0_n285 ),.Z(_AES_ENC_u0_N13 ) );
XOR2_X2 _AES_ENC_u0_U531  ( .A(_AES_ENC_w0[28] ), .B(_AES_ENC_u0_subword[28] ), .Z(_AES_ENC_u0_n285 ) );
XOR2_X2 _AES_ENC_u0_U530  ( .A(_AES_ENC_w1[28] ), .B(_AES_ENC_u0_N13 ), .Z(_AES_ENC_u0_N79 ) );
XOR2_X2 _AES_ENC_u0_U529  ( .A(_AES_ENC_w2[28] ), .B(_AES_ENC_u0_N79 ), .Z(_AES_ENC_u0_N145 ) );
XOR2_X2 _AES_ENC_u0_U528  ( .A(_AES_ENC_w3[28] ), .B(_AES_ENC_u0_N145 ), .Z(_AES_ENC_u0_N211 ) );
XOR2_X2 _AES_ENC_u0_U527  ( .A(_AES_ENC_u0_rcon[27]), .B(_AES_ENC_u0_n286 ),.Z(_AES_ENC_u0_N14 ) );
XOR2_X2 _AES_ENC_u0_U526  ( .A(_AES_ENC_w0[27] ), .B(_AES_ENC_u0_subword[27] ), .Z(_AES_ENC_u0_n286 ) );
XOR2_X2 _AES_ENC_u0_U525  ( .A(_AES_ENC_w1[27] ), .B(_AES_ENC_u0_N14 ), .Z(_AES_ENC_u0_N80 ) );
XOR2_X2 _AES_ENC_u0_U524  ( .A(_AES_ENC_w2[27] ), .B(_AES_ENC_u0_N80 ), .Z(_AES_ENC_u0_N146 ) );
XOR2_X2 _AES_ENC_u0_U523  ( .A(_AES_ENC_w3[27] ), .B(_AES_ENC_u0_N146 ), .Z(_AES_ENC_u0_N212 ) );
XOR2_X2 _AES_ENC_u0_U522  ( .A(_AES_ENC_u0_rcon[26]), .B(_AES_ENC_u0_n287 ),.Z(_AES_ENC_u0_N15 ) );
XOR2_X2 _AES_ENC_u0_U521  ( .A(_AES_ENC_w0[26] ), .B(_AES_ENC_u0_subword[26] ), .Z(_AES_ENC_u0_n287 ) );
XOR2_X2 _AES_ENC_u0_U520  ( .A(_AES_ENC_w1[26] ), .B(_AES_ENC_u0_N15 ), .Z(_AES_ENC_u0_N81 ) );
XOR2_X2 _AES_ENC_u0_U519  ( .A(_AES_ENC_w2[26] ), .B(_AES_ENC_u0_N81 ), .Z(_AES_ENC_u0_N147 ) );
XOR2_X2 _AES_ENC_u0_U518  ( .A(_AES_ENC_w3[26] ), .B(_AES_ENC_u0_N147 ), .Z(_AES_ENC_u0_N213 ) );
XOR2_X2 _AES_ENC_u0_U517  ( .A(_AES_ENC_u0_rcon[25]), .B(_AES_ENC_u0_n288 ),.Z(_AES_ENC_u0_N16 ) );
XOR2_X2 _AES_ENC_u0_U516  ( .A(_AES_ENC_w0[25] ), .B(_AES_ENC_u0_subword[25] ), .Z(_AES_ENC_u0_n288 ) );
XOR2_X2 _AES_ENC_u0_U515  ( .A(_AES_ENC_w1[25] ), .B(_AES_ENC_u0_N16 ), .Z(_AES_ENC_u0_N82 ) );
XOR2_X2 _AES_ENC_u0_U514  ( .A(_AES_ENC_w2[25] ), .B(_AES_ENC_u0_N82 ), .Z(_AES_ENC_u0_N148 ) );
XOR2_X2 _AES_ENC_u0_U513  ( .A(_AES_ENC_w3[25] ), .B(_AES_ENC_u0_N148 ), .Z(_AES_ENC_u0_N214 ) );
XOR2_X2 _AES_ENC_u0_U512  ( .A(_AES_ENC_u0_rcon[24]), .B(_AES_ENC_u0_n289 ),.Z(_AES_ENC_u0_N17 ) );
XOR2_X2 _AES_ENC_u0_U511  ( .A(_AES_ENC_w0[24] ), .B(_AES_ENC_u0_subword[24] ), .Z(_AES_ENC_u0_n289 ) );
XOR2_X2 _AES_ENC_u0_U510  ( .A(_AES_ENC_w1[24] ), .B(_AES_ENC_u0_N17 ), .Z(_AES_ENC_u0_N83 ) );
XOR2_X2 _AES_ENC_u0_U509  ( .A(_AES_ENC_w2[24] ), .B(_AES_ENC_u0_N83 ), .Z(_AES_ENC_u0_N149 ) );
XOR2_X2 _AES_ENC_u0_U508  ( .A(_AES_ENC_w3[24] ), .B(_AES_ENC_u0_N149 ), .Z(_AES_ENC_u0_N215 ) );
XOR2_X2 _AES_ENC_u0_U507  ( .A(_AES_ENC_u0_subword[23] ), .B(_AES_ENC_u0_n290 ), .Z(_AES_ENC_u0_N84 ) );
XOR2_X2 _AES_ENC_u0_U506  ( .A(_AES_ENC_w1[23] ), .B(_AES_ENC_w0[23] ), .Z(_AES_ENC_u0_n290 ) );
XOR2_X2 _AES_ENC_u0_U505  ( .A(_AES_ENC_w2[23] ), .B(_AES_ENC_u0_N84 ), .Z(_AES_ENC_u0_N150 ) );
XOR2_X2 _AES_ENC_u0_U504  ( .A(_AES_ENC_w3[23] ), .B(_AES_ENC_u0_N150 ), .Z(_AES_ENC_u0_N216 ) );
XOR2_X2 _AES_ENC_u0_U503  ( .A(_AES_ENC_u0_subword[22] ), .B(_AES_ENC_u0_n291 ), .Z(_AES_ENC_u0_N85 ) );
XOR2_X2 _AES_ENC_u0_U502  ( .A(_AES_ENC_w1[22] ), .B(_AES_ENC_w0[22] ), .Z(_AES_ENC_u0_n291 ) );
XOR2_X2 _AES_ENC_u0_U501  ( .A(_AES_ENC_w2[22] ), .B(_AES_ENC_u0_N85 ), .Z(_AES_ENC_u0_N151 ) );
XOR2_X2 _AES_ENC_u0_U500  ( .A(_AES_ENC_w3[22] ), .B(_AES_ENC_u0_N151 ), .Z(_AES_ENC_u0_N217 ) );
XOR2_X2 _AES_ENC_u0_U499  ( .A(_AES_ENC_u0_subword[21] ), .B(_AES_ENC_u0_n292 ), .Z(_AES_ENC_u0_N86 ) );
XOR2_X2 _AES_ENC_u0_U498  ( .A(_AES_ENC_w1[21] ), .B(_AES_ENC_w0[21] ), .Z(_AES_ENC_u0_n292 ) );
XOR2_X2 _AES_ENC_u0_U497  ( .A(_AES_ENC_w2[21] ), .B(_AES_ENC_u0_N86 ), .Z(_AES_ENC_u0_N152 ) );
XOR2_X2 _AES_ENC_u0_U496  ( .A(_AES_ENC_w3[21] ), .B(_AES_ENC_u0_N152 ), .Z(_AES_ENC_u0_N218 ) );
XOR2_X2 _AES_ENC_u0_U495  ( .A(_AES_ENC_u0_subword[20] ), .B(_AES_ENC_u0_n293 ), .Z(_AES_ENC_u0_N87 ) );
XOR2_X2 _AES_ENC_u0_U494  ( .A(_AES_ENC_w1[20] ), .B(_AES_ENC_w0[20] ), .Z(_AES_ENC_u0_n293 ) );
XOR2_X2 _AES_ENC_u0_U493  ( .A(_AES_ENC_w2[20] ), .B(_AES_ENC_u0_N87 ), .Z(_AES_ENC_u0_N153 ) );
XOR2_X2 _AES_ENC_u0_U492  ( .A(_AES_ENC_w3[20] ), .B(_AES_ENC_u0_N153 ), .Z(_AES_ENC_u0_N219 ) );
XOR2_X2 _AES_ENC_u0_U491  ( .A(_AES_ENC_u0_subword[19] ), .B(_AES_ENC_u0_n294 ), .Z(_AES_ENC_u0_N88 ) );
XOR2_X2 _AES_ENC_u0_U490  ( .A(_AES_ENC_w1[19] ), .B(_AES_ENC_w0[19] ), .Z(_AES_ENC_u0_n294 ) );
XOR2_X2 _AES_ENC_u0_U489  ( .A(_AES_ENC_w2[19] ), .B(_AES_ENC_u0_N88 ), .Z(_AES_ENC_u0_N154 ) );
XOR2_X2 _AES_ENC_u0_U488  ( .A(_AES_ENC_w3[19] ), .B(_AES_ENC_u0_N154 ), .Z(_AES_ENC_u0_N220 ) );
XOR2_X2 _AES_ENC_u0_U487  ( .A(_AES_ENC_u0_subword[18] ), .B(_AES_ENC_u0_n295 ), .Z(_AES_ENC_u0_N89 ) );
XOR2_X2 _AES_ENC_u0_U486  ( .A(_AES_ENC_w1[18] ), .B(_AES_ENC_w0[18] ), .Z(_AES_ENC_u0_n295 ) );
XOR2_X2 _AES_ENC_u0_U485  ( .A(_AES_ENC_w2[18] ), .B(_AES_ENC_u0_N89 ), .Z(_AES_ENC_u0_N155 ) );
XOR2_X2 _AES_ENC_u0_U484  ( .A(_AES_ENC_w3[18] ), .B(_AES_ENC_u0_N155 ), .Z(_AES_ENC_u0_N221 ) );
XOR2_X2 _AES_ENC_u0_U483  ( .A(_AES_ENC_u0_subword[17] ), .B(_AES_ENC_u0_n296 ), .Z(_AES_ENC_u0_N90 ) );
XOR2_X2 _AES_ENC_u0_U482  ( .A(_AES_ENC_w1[17] ), .B(_AES_ENC_w0[17] ), .Z(_AES_ENC_u0_n296 ) );
XOR2_X2 _AES_ENC_u0_U481  ( .A(_AES_ENC_w2[17] ), .B(_AES_ENC_u0_N90 ), .Z(_AES_ENC_u0_N156 ) );
XOR2_X2 _AES_ENC_u0_U480  ( .A(_AES_ENC_w3[17] ), .B(_AES_ENC_u0_N156 ), .Z(_AES_ENC_u0_N222 ) );
XOR2_X2 _AES_ENC_u0_U479  ( .A(_AES_ENC_u0_subword[16] ), .B(_AES_ENC_u0_n297 ), .Z(_AES_ENC_u0_N91 ) );
XOR2_X2 _AES_ENC_u0_U478  ( .A(_AES_ENC_w1[16] ), .B(_AES_ENC_w0[16] ), .Z(_AES_ENC_u0_n297 ) );
XOR2_X2 _AES_ENC_u0_U477  ( .A(_AES_ENC_w2[16] ), .B(_AES_ENC_u0_N91 ), .Z(_AES_ENC_u0_N157 ) );
XOR2_X2 _AES_ENC_u0_U476  ( .A(_AES_ENC_w3[16] ), .B(_AES_ENC_u0_N157 ), .Z(_AES_ENC_u0_N223 ) );
XOR2_X2 _AES_ENC_u0_U475  ( .A(_AES_ENC_u0_subword[15] ), .B(_AES_ENC_u0_n298 ), .Z(_AES_ENC_u0_N92 ) );
XOR2_X2 _AES_ENC_u0_U474  ( .A(_AES_ENC_w1[15] ), .B(_AES_ENC_w0[15] ), .Z(_AES_ENC_u0_n298 ) );
XOR2_X2 _AES_ENC_u0_U473  ( .A(_AES_ENC_w2[15] ), .B(_AES_ENC_u0_N92 ), .Z(_AES_ENC_u0_N158 ) );
XOR2_X2 _AES_ENC_u0_U472  ( .A(_AES_ENC_w3[15] ), .B(_AES_ENC_u0_N158 ), .Z(_AES_ENC_u0_N224 ) );
XOR2_X2 _AES_ENC_u0_U471  ( .A(_AES_ENC_u0_subword[14] ), .B(_AES_ENC_u0_n299 ), .Z(_AES_ENC_u0_N93 ) );
XOR2_X2 _AES_ENC_u0_U470  ( .A(_AES_ENC_w1[14] ), .B(_AES_ENC_w0[14] ), .Z(_AES_ENC_u0_n299 ) );
XOR2_X2 _AES_ENC_u0_U469  ( .A(_AES_ENC_w2[14] ), .B(_AES_ENC_u0_N93 ), .Z(_AES_ENC_u0_N159 ) );
XOR2_X2 _AES_ENC_u0_U468  ( .A(_AES_ENC_w3[14] ), .B(_AES_ENC_u0_N159 ), .Z(_AES_ENC_u0_N225 ) );
XOR2_X2 _AES_ENC_u0_U467  ( .A(_AES_ENC_u0_subword[13] ), .B(_AES_ENC_u0_n300 ), .Z(_AES_ENC_u0_N94 ) );
XOR2_X2 _AES_ENC_u0_U466  ( .A(_AES_ENC_w1[13] ), .B(_AES_ENC_w0[13] ), .Z(_AES_ENC_u0_n300 ) );
XOR2_X2 _AES_ENC_u0_U465  ( .A(_AES_ENC_w2[13] ), .B(_AES_ENC_u0_N94 ), .Z(_AES_ENC_u0_N160 ) );
XOR2_X2 _AES_ENC_u0_U464  ( .A(_AES_ENC_w3[13] ), .B(_AES_ENC_u0_N160 ), .Z(_AES_ENC_u0_N226 ) );
XOR2_X2 _AES_ENC_u0_U463  ( .A(_AES_ENC_u0_subword[12] ), .B(_AES_ENC_u0_n301 ), .Z(_AES_ENC_u0_N95 ) );
XOR2_X2 _AES_ENC_u0_U462  ( .A(_AES_ENC_w1[12] ), .B(_AES_ENC_w0[12] ), .Z(_AES_ENC_u0_n301 ) );
XOR2_X2 _AES_ENC_u0_U461  ( .A(_AES_ENC_w2[12] ), .B(_AES_ENC_u0_N95 ), .Z(_AES_ENC_u0_N161 ) );
XOR2_X2 _AES_ENC_u0_U460  ( .A(_AES_ENC_w3[12] ), .B(_AES_ENC_u0_N161 ), .Z(_AES_ENC_u0_N227 ) );
XOR2_X2 _AES_ENC_u0_U459  ( .A(_AES_ENC_u0_subword[11] ), .B(_AES_ENC_u0_n302 ), .Z(_AES_ENC_u0_N96 ) );
XOR2_X2 _AES_ENC_u0_U458  ( .A(_AES_ENC_w1[11] ), .B(_AES_ENC_w0[11] ), .Z(_AES_ENC_u0_n302 ) );
XOR2_X2 _AES_ENC_u0_U457  ( .A(_AES_ENC_w2[11] ), .B(_AES_ENC_u0_N96 ), .Z(_AES_ENC_u0_N162 ) );
XOR2_X2 _AES_ENC_u0_U456  ( .A(_AES_ENC_w3[11] ), .B(_AES_ENC_u0_N162 ), .Z(_AES_ENC_u0_N228 ) );
XOR2_X2 _AES_ENC_u0_U455  ( .A(_AES_ENC_u0_subword[10] ), .B(_AES_ENC_u0_n303 ), .Z(_AES_ENC_u0_N97 ) );
XOR2_X2 _AES_ENC_u0_U454  ( .A(_AES_ENC_w1[10] ), .B(_AES_ENC_w0[10] ), .Z(_AES_ENC_u0_n303 ) );
XOR2_X2 _AES_ENC_u0_U453  ( .A(_AES_ENC_w2[10] ), .B(_AES_ENC_u0_N97 ), .Z(_AES_ENC_u0_N163 ) );
XOR2_X2 _AES_ENC_u0_U452  ( .A(_AES_ENC_w3[10] ), .B(_AES_ENC_u0_N163 ), .Z(_AES_ENC_u0_N229 ) );
XOR2_X2 _AES_ENC_u0_U451  ( .A(_AES_ENC_u0_subword[9] ), .B(_AES_ENC_u0_n304 ), .Z(_AES_ENC_u0_N98 ) );
XOR2_X2 _AES_ENC_u0_U450  ( .A(_AES_ENC_w1[9] ), .B(_AES_ENC_w0[9] ), .Z(_AES_ENC_u0_n304 ) );
XOR2_X2 _AES_ENC_u0_U449  ( .A(_AES_ENC_w2[9] ), .B(_AES_ENC_u0_N98 ), .Z(_AES_ENC_u0_N164 ) );
XOR2_X2 _AES_ENC_u0_U448  ( .A(_AES_ENC_w3[9] ), .B(_AES_ENC_u0_N164 ), .Z(_AES_ENC_u0_N230 ) );
XOR2_X2 _AES_ENC_u0_U447  ( .A(_AES_ENC_u0_subword[8] ), .B(_AES_ENC_u0_n305 ), .Z(_AES_ENC_u0_N99 ) );
XOR2_X2 _AES_ENC_u0_U446  ( .A(_AES_ENC_w1[8] ), .B(_AES_ENC_w0[8] ), .Z(_AES_ENC_u0_n305 ) );
XOR2_X2 _AES_ENC_u0_U445  ( .A(_AES_ENC_w2[8] ), .B(_AES_ENC_u0_N99 ), .Z(_AES_ENC_u0_N165 ) );
XOR2_X2 _AES_ENC_u0_U444  ( .A(_AES_ENC_w3[8] ), .B(_AES_ENC_u0_N165 ), .Z(_AES_ENC_u0_N231 ) );
XOR2_X2 _AES_ENC_u0_U443  ( .A(_AES_ENC_u0_subword[7] ), .B(_AES_ENC_u0_n306 ), .Z(_AES_ENC_u0_N100 ) );
XOR2_X2 _AES_ENC_u0_U442  ( .A(_AES_ENC_w1[7] ), .B(_AES_ENC_w0[7] ), .Z(_AES_ENC_u0_n306 ) );
XOR2_X2 _AES_ENC_u0_U441  ( .A(_AES_ENC_w2[7] ), .B(_AES_ENC_u0_N100 ), .Z(_AES_ENC_u0_N166 ) );
XOR2_X2 _AES_ENC_u0_U440  ( .A(_AES_ENC_w3[7] ), .B(_AES_ENC_u0_N166 ), .Z(_AES_ENC_u0_N232 ) );
XOR2_X2 _AES_ENC_u0_U439  ( .A(_AES_ENC_u0_subword[6] ), .B(_AES_ENC_u0_n307 ), .Z(_AES_ENC_u0_N101 ) );
XOR2_X2 _AES_ENC_u0_U438  ( .A(_AES_ENC_w1[6] ), .B(_AES_ENC_w0[6] ), .Z(_AES_ENC_u0_n307 ) );
XOR2_X2 _AES_ENC_u0_U437  ( .A(_AES_ENC_w2[6] ), .B(_AES_ENC_u0_N101 ), .Z(_AES_ENC_u0_N167 ) );
XOR2_X2 _AES_ENC_u0_U436  ( .A(_AES_ENC_w3[6] ), .B(_AES_ENC_u0_N167 ), .Z(_AES_ENC_u0_N233 ) );
XOR2_X2 _AES_ENC_u0_U435  ( .A(_AES_ENC_u0_subword[5] ), .B(_AES_ENC_u0_n308 ), .Z(_AES_ENC_u0_N102 ) );
XOR2_X2 _AES_ENC_u0_U434  ( .A(_AES_ENC_w1[5] ), .B(_AES_ENC_w0[5] ), .Z(_AES_ENC_u0_n308 ) );
XOR2_X2 _AES_ENC_u0_U433  ( .A(_AES_ENC_w2[5] ), .B(_AES_ENC_u0_N102 ), .Z(_AES_ENC_u0_N168 ) );
XOR2_X2 _AES_ENC_u0_U432  ( .A(_AES_ENC_w3[5] ), .B(_AES_ENC_u0_N168 ), .Z(_AES_ENC_u0_N234 ) );
XOR2_X2 _AES_ENC_u0_U431  ( .A(_AES_ENC_u0_subword[4] ), .B(_AES_ENC_u0_n309 ), .Z(_AES_ENC_u0_N103 ) );
XOR2_X2 _AES_ENC_u0_U430  ( .A(_AES_ENC_w1[4] ), .B(_AES_ENC_w0[4] ), .Z(_AES_ENC_u0_n309 ) );
XOR2_X2 _AES_ENC_u0_U429  ( .A(_AES_ENC_w2[4] ), .B(_AES_ENC_u0_N103 ), .Z(_AES_ENC_u0_N169 ) );
XOR2_X2 _AES_ENC_u0_U428  ( .A(_AES_ENC_w3[4] ), .B(_AES_ENC_u0_N169 ), .Z(_AES_ENC_u0_N235 ) );
XOR2_X2 _AES_ENC_u0_U427  ( .A(_AES_ENC_u0_subword[3] ), .B(_AES_ENC_u0_n310 ), .Z(_AES_ENC_u0_N104 ) );
XOR2_X2 _AES_ENC_u0_U426  ( .A(_AES_ENC_w1[3] ), .B(_AES_ENC_w0[3] ), .Z(_AES_ENC_u0_n310 ) );
XOR2_X2 _AES_ENC_u0_U425  ( .A(_AES_ENC_w2[3] ), .B(_AES_ENC_u0_N104 ), .Z(_AES_ENC_u0_N170 ) );
XOR2_X2 _AES_ENC_u0_U424  ( .A(_AES_ENC_w3[3] ), .B(_AES_ENC_u0_N170 ), .Z(_AES_ENC_u0_N236 ) );
XOR2_X2 _AES_ENC_u0_U423  ( .A(_AES_ENC_u0_subword[2] ), .B(_AES_ENC_u0_n311 ), .Z(_AES_ENC_u0_N105 ) );
XOR2_X2 _AES_ENC_u0_U422  ( .A(_AES_ENC_w1[2] ), .B(_AES_ENC_w0[2] ), .Z(_AES_ENC_u0_n311 ) );
XOR2_X2 _AES_ENC_u0_U421  ( .A(_AES_ENC_w2[2] ), .B(_AES_ENC_u0_N105 ), .Z(_AES_ENC_u0_N171 ) );
XOR2_X2 _AES_ENC_u0_U420  ( .A(_AES_ENC_w3[2] ), .B(_AES_ENC_u0_N171 ), .Z(_AES_ENC_u0_N237 ) );
XOR2_X2 _AES_ENC_u0_U419  ( .A(_AES_ENC_u0_subword[1] ), .B(_AES_ENC_u0_n312 ), .Z(_AES_ENC_u0_N106 ) );
XOR2_X2 _AES_ENC_u0_U418  ( .A(_AES_ENC_w1[1] ), .B(_AES_ENC_w0[1] ), .Z(_AES_ENC_u0_n312 ) );
XOR2_X2 _AES_ENC_u0_U417  ( .A(_AES_ENC_w2[1] ), .B(_AES_ENC_u0_N106 ), .Z(_AES_ENC_u0_N172 ) );
XOR2_X2 _AES_ENC_u0_U416  ( .A(_AES_ENC_w3[1] ), .B(_AES_ENC_u0_N172 ), .Z(_AES_ENC_u0_N238 ) );
XOR2_X2 _AES_ENC_u0_U415  ( .A(_AES_ENC_u0_subword[0] ), .B(_AES_ENC_u0_n313 ), .Z(_AES_ENC_u0_N107 ) );
XOR2_X2 _AES_ENC_u0_U414  ( .A(_AES_ENC_w1[0] ), .B(_AES_ENC_w0[0] ), .Z(_AES_ENC_u0_n313 ) );
XOR2_X2 _AES_ENC_u0_U413  ( .A(_AES_ENC_w2[0] ), .B(_AES_ENC_u0_N107 ), .Z(_AES_ENC_u0_N173 ) );
XOR2_X2 _AES_ENC_u0_U412  ( .A(_AES_ENC_w3[0] ), .B(_AES_ENC_u0_N173 ), .Z(_AES_ENC_u0_N239 ) );
INV_X4 _AES_ENC_u0_u0_U575  ( .A(_AES_ENC_w3[23] ), .ZN(_AES_ENC_u0_u0_n627 ) );
INV_X4 _AES_ENC_u0_u0_U574  ( .A(_AES_ENC_u0_u0_n1114 ), .ZN(_AES_ENC_u0_u0_n625 ) );
INV_X4 _AES_ENC_u0_u0_U573  ( .A(_AES_ENC_w3[20] ), .ZN(_AES_ENC_u0_u0_n624 ) );
INV_X4 _AES_ENC_u0_u0_U572  ( .A(_AES_ENC_u0_u0_n1025 ), .ZN(_AES_ENC_u0_u0_n622 ) );
INV_X4 _AES_ENC_u0_u0_U571  ( .A(_AES_ENC_u0_u0_n1120 ), .ZN(_AES_ENC_u0_u0_n620 ) );
INV_X4 _AES_ENC_u0_u0_U570  ( .A(_AES_ENC_u0_u0_n1121 ), .ZN(_AES_ENC_u0_u0_n619 ) );
INV_X4 _AES_ENC_u0_u0_U569  ( .A(_AES_ENC_u0_u0_n1048 ), .ZN(_AES_ENC_u0_u0_n618 ) );
INV_X4 _AES_ENC_u0_u0_U568  ( .A(_AES_ENC_u0_u0_n974 ), .ZN(_AES_ENC_u0_u0_n616 ) );
INV_X4 _AES_ENC_u0_u0_U567  ( .A(_AES_ENC_u0_u0_n794 ), .ZN(_AES_ENC_u0_u0_n614 ) );
INV_X4 _AES_ENC_u0_u0_U566  ( .A(_AES_ENC_w3[18] ), .ZN(_AES_ENC_u0_u0_n611 ) );
INV_X4 _AES_ENC_u0_u0_U565  ( .A(_AES_ENC_u0_u0_n800 ), .ZN(_AES_ENC_u0_u0_n610 ) );
INV_X4 _AES_ENC_u0_u0_U564  ( .A(_AES_ENC_u0_u0_n925 ), .ZN(_AES_ENC_u0_u0_n609 ) );
INV_X4 _AES_ENC_u0_u0_U563  ( .A(_AES_ENC_u0_u0_n779 ), .ZN(_AES_ENC_u0_u0_n607 ) );
INV_X4 _AES_ENC_u0_u0_U562  ( .A(_AES_ENC_u0_u0_n1022 ), .ZN(_AES_ENC_u0_u0_n603 ) );
INV_X4 _AES_ENC_u0_u0_U561  ( .A(_AES_ENC_u0_u0_n1102 ), .ZN(_AES_ENC_u0_u0_n602 ) );
INV_X4 _AES_ENC_u0_u0_U560  ( .A(_AES_ENC_u0_u0_n929 ), .ZN(_AES_ENC_u0_u0_n601 ) );
INV_X4 _AES_ENC_u0_u0_U559  ( .A(_AES_ENC_u0_u0_n1056 ), .ZN(_AES_ENC_u0_u0_n600 ) );
INV_X4 _AES_ENC_u0_u0_U558  ( .A(_AES_ENC_u0_u0_n1054 ), .ZN(_AES_ENC_u0_u0_n599 ) );
INV_X4 _AES_ENC_u0_u0_U557  ( .A(_AES_ENC_u0_u0_n881 ), .ZN(_AES_ENC_u0_u0_n598 ) );
INV_X4 _AES_ENC_u0_u0_U556  ( .A(_AES_ENC_u0_u0_n926 ), .ZN(_AES_ENC_u0_u0_n597 ) );
INV_X4 _AES_ENC_u0_u0_U555  ( .A(_AES_ENC_u0_u0_n977 ), .ZN(_AES_ENC_u0_u0_n595 ) );
INV_X4 _AES_ENC_u0_u0_U554  ( .A(_AES_ENC_u0_u0_n1031 ), .ZN(_AES_ENC_u0_u0_n594 ) );
INV_X4 _AES_ENC_u0_u0_U553  ( .A(_AES_ENC_u0_u0_n1103 ), .ZN(_AES_ENC_u0_u0_n593 ) );
INV_X4 _AES_ENC_u0_u0_U552  ( .A(_AES_ENC_u0_u0_n1009 ), .ZN(_AES_ENC_u0_u0_n592 ) );
INV_X4 _AES_ENC_u0_u0_U551  ( .A(_AES_ENC_u0_u0_n990 ), .ZN(_AES_ENC_u0_u0_n591 ) );
INV_X4 _AES_ENC_u0_u0_U550  ( .A(_AES_ENC_u0_u0_n1058 ), .ZN(_AES_ENC_u0_u0_n590 ) );
INV_X4 _AES_ENC_u0_u0_U549  ( .A(_AES_ENC_u0_u0_n1074 ), .ZN(_AES_ENC_u0_u0_n589 ) );
INV_X4 _AES_ENC_u0_u0_U548  ( .A(_AES_ENC_u0_u0_n1053 ), .ZN(_AES_ENC_u0_u0_n588 ) );
INV_X4 _AES_ENC_u0_u0_U547  ( .A(_AES_ENC_u0_u0_n826 ), .ZN(_AES_ENC_u0_u0_n587 ) );
INV_X4 _AES_ENC_u0_u0_U546  ( .A(_AES_ENC_u0_u0_n992 ), .ZN(_AES_ENC_u0_u0_n586 ) );
INV_X4 _AES_ENC_u0_u0_U545  ( .A(_AES_ENC_u0_u0_n821 ), .ZN(_AES_ENC_u0_u0_n585 ) );
INV_X4 _AES_ENC_u0_u0_U544  ( .A(_AES_ENC_u0_u0_n910 ), .ZN(_AES_ENC_u0_u0_n584 ) );
INV_X4 _AES_ENC_u0_u0_U543  ( .A(_AES_ENC_u0_u0_n906 ), .ZN(_AES_ENC_u0_u0_n583 ) );
INV_X4 _AES_ENC_u0_u0_U542  ( .A(_AES_ENC_u0_u0_n880 ), .ZN(_AES_ENC_u0_u0_n581 ) );
INV_X4 _AES_ENC_u0_u0_U541  ( .A(_AES_ENC_u0_u0_n1013 ), .ZN(_AES_ENC_u0_u0_n580 ) );
INV_X4 _AES_ENC_u0_u0_U540  ( .A(_AES_ENC_u0_u0_n1092 ), .ZN(_AES_ENC_u0_u0_n579 ) );
INV_X4 _AES_ENC_u0_u0_U539  ( .A(_AES_ENC_u0_u0_n824 ), .ZN(_AES_ENC_u0_u0_n578 ) );
INV_X4 _AES_ENC_u0_u0_U538  ( .A(_AES_ENC_u0_u0_n1091 ), .ZN(_AES_ENC_u0_u0_n577 ) );
INV_X4 _AES_ENC_u0_u0_U537  ( .A(_AES_ENC_u0_u0_n1080 ), .ZN(_AES_ENC_u0_u0_n576 ) );
INV_X4 _AES_ENC_u0_u0_U536  ( .A(_AES_ENC_u0_u0_n959 ), .ZN(_AES_ENC_u0_u0_n575 ) );
INV_X4 _AES_ENC_u0_u0_U535  ( .A(_AES_ENC_w3[16] ), .ZN(_AES_ENC_u0_u0_n574 ) );
NOR2_X2 _AES_ENC_u0_u0_U534  ( .A1(_AES_ENC_w3[20] ), .A2(_AES_ENC_w3[19] ),.ZN(_AES_ENC_u0_u0_n1025 ) );
INV_X4 _AES_ENC_u0_u0_U533  ( .A(_AES_ENC_u0_u0_n569 ), .ZN(_AES_ENC_u0_u0_n572 ) );
NOR2_X2 _AES_ENC_u0_u0_U532  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n765 ) );
NOR2_X2 _AES_ENC_u0_u0_U531  ( .A1(_AES_ENC_w3[20] ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n764 ) );
NOR2_X2 _AES_ENC_u0_u0_U530  ( .A1(_AES_ENC_u0_u0_n765 ), .A2(_AES_ENC_u0_u0_n764 ), .ZN(_AES_ENC_u0_u0_n766 ) );
NOR2_X2 _AES_ENC_u0_u0_U529  ( .A1(_AES_ENC_u0_u0_n766 ), .A2(_AES_ENC_u0_u0_n575 ), .ZN(_AES_ENC_u0_u0_n767 ) );
NOR2_X2 _AES_ENC_u0_u0_U528  ( .A1(_AES_ENC_u0_u0_n1117 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n707 ) );
NOR3_X2 _AES_ENC_u0_u0_U527  ( .A1(_AES_ENC_u0_u0_n627 ), .A2(_AES_ENC_w3[21] ), .A3(_AES_ENC_u0_u0_n704 ), .ZN(_AES_ENC_u0_u0_n706 ) );
NOR2_X2 _AES_ENC_u0_u0_U526  ( .A1(_AES_ENC_w3[20] ), .A2(_AES_ENC_u0_u0_n579 ), .ZN(_AES_ENC_u0_u0_n705 ) );
NOR3_X2 _AES_ENC_u0_u0_U525  ( .A1(_AES_ENC_u0_u0_n707 ), .A2(_AES_ENC_u0_u0_n706 ), .A3(_AES_ENC_u0_u0_n705 ), .ZN(_AES_ENC_u0_u0_n713 ) );
NOR4_X2 _AES_ENC_u0_u0_U524  ( .A1(_AES_ENC_u0_u0_n633 ), .A2(_AES_ENC_u0_u0_n632 ), .A3(_AES_ENC_u0_u0_n631 ), .A4(_AES_ENC_u0_u0_n630 ), .ZN(_AES_ENC_u0_u0_n634 ) );
NOR2_X2 _AES_ENC_u0_u0_U523  ( .A1(_AES_ENC_u0_u0_n629 ), .A2(_AES_ENC_u0_u0_n628 ), .ZN(_AES_ENC_u0_u0_n635 ) );
NAND3_X2 _AES_ENC_u0_u0_U522  ( .A1(_AES_ENC_w3[18] ), .A2(_AES_ENC_w3[23] ),.A3(_AES_ENC_u0_u0_n1059 ), .ZN(_AES_ENC_u0_u0_n636 ) );
INV_X4 _AES_ENC_u0_u0_U521  ( .A(_AES_ENC_w3[19] ), .ZN(_AES_ENC_u0_u0_n621 ) );
NOR2_X2 _AES_ENC_u0_u0_U520  ( .A1(_AES_ENC_w3[21] ), .A2(_AES_ENC_w3[18] ),.ZN(_AES_ENC_u0_u0_n974 ) );
NAND3_X2 _AES_ENC_u0_u0_U519  ( .A1(_AES_ENC_u0_u0_n652 ), .A2(_AES_ENC_u0_u0_n626 ), .A3(_AES_ENC_w3[23] ), .ZN(_AES_ENC_u0_u0_n653 ) );
NOR2_X2 _AES_ENC_u0_u0_U518  ( .A1(_AES_ENC_u0_u0_n611 ), .A2(_AES_ENC_w3[21] ), .ZN(_AES_ENC_u0_u0_n925 ) );
NOR2_X2 _AES_ENC_u0_u0_U517  ( .A1(_AES_ENC_u0_u0_n626 ), .A2(_AES_ENC_w3[18] ), .ZN(_AES_ENC_u0_u0_n1048 ) );
INV_X4 _AES_ENC_u0_u0_U516  ( .A(_AES_ENC_w3[21] ), .ZN(_AES_ENC_u0_u0_n626 ) );
NOR2_X2 _AES_ENC_u0_u0_U515  ( .A1(_AES_ENC_u0_u0_n611 ), .A2(_AES_ENC_w3[23] ), .ZN(_AES_ENC_u0_u0_n779 ) );
NOR2_X2 _AES_ENC_u0_u0_U512  ( .A1(_AES_ENC_w3[23] ), .A2(_AES_ENC_w3[18] ),.ZN(_AES_ENC_u0_u0_n794 ) );
NAND3_X2 _AES_ENC_u0_u0_U510  ( .A1(_AES_ENC_u0_u0_n679 ), .A2(_AES_ENC_u0_u0_n678 ), .A3(_AES_ENC_u0_u0_n677 ), .ZN(_AES_ENC_u0_subword[24] ) );
NOR2_X2 _AES_ENC_u0_u0_U509  ( .A1(_AES_ENC_u0_u0_n574 ), .A2(_AES_ENC_w3[22] ), .ZN(_AES_ENC_u0_u0_n1070 ) );
NOR2_X2 _AES_ENC_u0_u0_U508  ( .A1(_AES_ENC_w3[16] ), .A2(_AES_ENC_w3[22] ),.ZN(_AES_ENC_u0_u0_n1090 ) );
NOR2_X2 _AES_ENC_u0_u0_U507  ( .A1(_AES_ENC_w3[20] ), .A2(_AES_ENC_w3[17] ),.ZN(_AES_ENC_u0_u0_n1102 ) );
NOR2_X2 _AES_ENC_u0_u0_U506  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_w3[19] ), .ZN(_AES_ENC_u0_u0_n1053 ) );
NOR2_X2 _AES_ENC_u0_u0_U505  ( .A1(_AES_ENC_u0_u0_n607 ), .A2(_AES_ENC_w3[21] ), .ZN(_AES_ENC_u0_u0_n1024 ) );
NOR2_X2 _AES_ENC_u0_u0_U504  ( .A1(_AES_ENC_u0_u0_n625 ), .A2(_AES_ENC_w3[18] ), .ZN(_AES_ENC_u0_u0_n1093 ) );
NOR2_X2 _AES_ENC_u0_u0_U503  ( .A1(_AES_ENC_u0_u0_n614 ), .A2(_AES_ENC_w3[21] ), .ZN(_AES_ENC_u0_u0_n1094 ) );
NOR2_X2 _AES_ENC_u0_u0_U502  ( .A1(_AES_ENC_u0_u0_n624 ), .A2(_AES_ENC_w3[19] ), .ZN(_AES_ENC_u0_u0_n931 ) );
INV_X4 _AES_ENC_u0_u0_U501  ( .A(_AES_ENC_u0_u0_n570 ), .ZN(_AES_ENC_u0_u0_n573 ) );
NOR2_X2 _AES_ENC_u0_u0_U500  ( .A1(_AES_ENC_u0_u0_n622 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n1059 ) );
NOR4_X2 _AES_ENC_u0_u0_U499  ( .A1(_AES_ENC_u0_u0_n1125 ), .A2(_AES_ENC_u0_u0_n1124 ), .A3(_AES_ENC_u0_u0_n1123 ), .A4(_AES_ENC_u0_u0_n1122 ), .ZN(_AES_ENC_u0_u0_n1126 ) );
NOR2_X2 _AES_ENC_u0_u0_U498  ( .A1(_AES_ENC_u0_u0_n826 ), .A2(_AES_ENC_u0_u0_n572 ), .ZN(_AES_ENC_u0_u0_n827 ) );
NOR3_X2 _AES_ENC_u0_u0_U497  ( .A1(_AES_ENC_u0_u0_n769 ), .A2(_AES_ENC_u0_u0_n768 ), .A3(_AES_ENC_u0_u0_n767 ), .ZN(_AES_ENC_u0_u0_n775 ) );
NOR2_X2 _AES_ENC_u0_u0_U496  ( .A1(_AES_ENC_u0_u0_n946 ), .A2(_AES_ENC_u0_u0_n945 ), .ZN(_AES_ENC_u0_u0_n952 ) );
NOR2_X2 _AES_ENC_u0_u0_U495  ( .A1(_AES_ENC_w3[17] ), .A2(_AES_ENC_u0_u0_n623 ), .ZN(_AES_ENC_u0_u0_n913 ) );
NOR2_X2 _AES_ENC_u0_u0_U494  ( .A1(_AES_ENC_u0_u0_n913 ), .A2(_AES_ENC_u0_u0_n1091 ), .ZN(_AES_ENC_u0_u0_n914 ) );
NOR2_X2 _AES_ENC_u0_u0_U492  ( .A1(_AES_ENC_u0_u0_n1056 ), .A2(_AES_ENC_u0_u0_n1053 ), .ZN(_AES_ENC_u0_u0_n749 ) );
NOR2_X2 _AES_ENC_u0_u0_U491  ( .A1(_AES_ENC_u0_u0_n749 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n752 ) );
NOR4_X2 _AES_ENC_u0_u0_U490  ( .A1(_AES_ENC_u0_u0_n983 ), .A2(_AES_ENC_u0_u0_n698 ), .A3(_AES_ENC_u0_u0_n697 ), .A4(_AES_ENC_u0_u0_n696 ), .ZN(_AES_ENC_u0_u0_n699 ) );
NOR3_X2 _AES_ENC_u0_u0_U489  ( .A1(_AES_ENC_u0_u0_n695 ), .A2(_AES_ENC_u0_u0_n694 ), .A3(_AES_ENC_u0_u0_n693 ), .ZN(_AES_ENC_u0_u0_n700 ) );
NOR4_X2 _AES_ENC_u0_u0_U488  ( .A1(_AES_ENC_u0_u0_n757 ), .A2(_AES_ENC_u0_u0_n756 ), .A3(_AES_ENC_u0_u0_n755 ), .A4(_AES_ENC_u0_u0_n754 ), .ZN(_AES_ENC_u0_u0_n758 ) );
NOR2_X2 _AES_ENC_u0_u0_U487  ( .A1(_AES_ENC_u0_u0_n752 ), .A2(_AES_ENC_u0_u0_n751 ), .ZN(_AES_ENC_u0_u0_n759 ) );
NOR4_X2 _AES_ENC_u0_u0_U486  ( .A1(_AES_ENC_u0_u0_n870 ), .A2(_AES_ENC_u0_u0_n869 ), .A3(_AES_ENC_u0_u0_n868 ), .A4(_AES_ENC_u0_u0_n867 ), .ZN(_AES_ENC_u0_u0_n871 ) );
NOR3_X2 _AES_ENC_u0_u0_U483  ( .A1(_AES_ENC_u0_u0_n995 ), .A2(_AES_ENC_u0_u0_n586 ), .A3(_AES_ENC_u0_u0_n994 ), .ZN(_AES_ENC_u0_u0_n1002 ) );
NOR2_X2 _AES_ENC_u0_u0_U482  ( .A1(_AES_ENC_u0_u0_n1076 ), .A2(_AES_ENC_u0_u0_n1075 ), .ZN(_AES_ENC_u0_u0_n1086 ) );
NOR2_X2 _AES_ENC_u0_u0_U480  ( .A1(_AES_ENC_u0_u0_n1053 ), .A2(_AES_ENC_u0_u0_n1095 ), .ZN(_AES_ENC_u0_u0_n639 ) );
NOR2_X2 _AES_ENC_u0_u0_U479  ( .A1(_AES_ENC_u0_u0_n639 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n640 ) );
NOR2_X2 _AES_ENC_u0_u0_U478  ( .A1(_AES_ENC_u0_u0_n909 ), .A2(_AES_ENC_u0_u0_n908 ), .ZN(_AES_ENC_u0_u0_n920 ) );
INV_X4 _AES_ENC_u0_u0_U477  ( .A(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n596 ) );
NOR2_X2 _AES_ENC_u0_u0_U474  ( .A1(_AES_ENC_u0_u0_n932 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n933 ) );
NOR2_X2 _AES_ENC_u0_u0_U473  ( .A1(_AES_ENC_u0_u0_n929 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n935 ) );
NOR2_X2 _AES_ENC_u0_u0_U472  ( .A1(_AES_ENC_u0_u0_n931 ), .A2(_AES_ENC_u0_u0_n930 ), .ZN(_AES_ENC_u0_u0_n934 ) );
NOR3_X2 _AES_ENC_u0_u0_U471  ( .A1(_AES_ENC_u0_u0_n935 ), .A2(_AES_ENC_u0_u0_n934 ), .A3(_AES_ENC_u0_u0_n933 ), .ZN(_AES_ENC_u0_u0_n936 ) );
OR2_X4 _AES_ENC_u0_u0_U470  ( .A1(_AES_ENC_u0_u0_n1094 ), .A2(_AES_ENC_u0_u0_n1093 ), .ZN(_AES_ENC_u0_u0_n571 ) );
AND2_X2 _AES_ENC_u0_u0_U469  ( .A1(_AES_ENC_u0_u0_n571 ), .A2(_AES_ENC_u0_u0_n1095 ), .ZN(_AES_ENC_u0_u0_n1101 ) );
NOR2_X2 _AES_ENC_u0_u0_U468  ( .A1(_AES_ENC_u0_u0_n1074 ), .A2(_AES_ENC_u0_u0_n931 ), .ZN(_AES_ENC_u0_u0_n796 ) );
NOR2_X2 _AES_ENC_u0_u0_U467  ( .A1(_AES_ENC_u0_u0_n796 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n797 ) );
NOR2_X2 _AES_ENC_u0_u0_U466  ( .A1(_AES_ENC_u0_u0_n1054 ), .A2(_AES_ENC_u0_u0_n1053 ), .ZN(_AES_ENC_u0_u0_n1055 ) );
NOR2_X2 _AES_ENC_u0_u0_U465  ( .A1(_AES_ENC_u0_u0_n1049 ), .A2(_AES_ENC_u0_u0_n618 ), .ZN(_AES_ENC_u0_u0_n1051 ) );
NOR2_X2 _AES_ENC_u0_u0_U464  ( .A1(_AES_ENC_u0_u0_n1051 ), .A2(_AES_ENC_u0_u0_n1050 ), .ZN(_AES_ENC_u0_u0_n1052 ) );
NOR2_X2 _AES_ENC_u0_u0_U463  ( .A1(_AES_ENC_u0_u0_n1052 ), .A2(_AES_ENC_u0_u0_n592 ), .ZN(_AES_ENC_u0_u0_n1064 ) );
NOR2_X2 _AES_ENC_u0_u0_U462  ( .A1(_AES_ENC_w3[17] ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n631 ) );
NOR2_X2 _AES_ENC_u0_u0_U461  ( .A1(_AES_ENC_u0_u0_n1025 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n980 ) );
NOR2_X2 _AES_ENC_u0_u0_U460  ( .A1(_AES_ENC_u0_u0_n1073 ), .A2(_AES_ENC_u0_u0_n1094 ), .ZN(_AES_ENC_u0_u0_n795 ) );
NOR2_X2 _AES_ENC_u0_u0_U459  ( .A1(_AES_ENC_u0_u0_n795 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n799 ) );
NOR2_X2 _AES_ENC_u0_u0_U458  ( .A1(_AES_ENC_u0_u0_n624 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n1075 ) );
NOR2_X2 _AES_ENC_u0_u0_U455  ( .A1(_AES_ENC_u0_u0_n624 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n822 ) );
NOR2_X2 _AES_ENC_u0_u0_U448  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n823 ) );
NOR2_X2 _AES_ENC_u0_u0_U447  ( .A1(_AES_ENC_u0_u0_n823 ), .A2(_AES_ENC_u0_u0_n822 ), .ZN(_AES_ENC_u0_u0_n825 ) );
NOR2_X2 _AES_ENC_u0_u0_U442  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n981 ) );
NOR2_X2 _AES_ENC_u0_u0_U441  ( .A1(_AES_ENC_u0_u0_n1074 ), .A2(_AES_ENC_u0_u0_n1025 ), .ZN(_AES_ENC_u0_u0_n891 ) );
NOR2_X2 _AES_ENC_u0_u0_U438  ( .A1(_AES_ENC_u0_u0_n1102 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n643 ) );
NOR2_X2 _AES_ENC_u0_u0_U435  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n621 ), .ZN(_AES_ENC_u0_u0_n642 ) );
NOR2_X2 _AES_ENC_u0_u0_U434  ( .A1(_AES_ENC_u0_u0_n911 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n644 ) );
NOR4_X2 _AES_ENC_u0_u0_U433  ( .A1(_AES_ENC_u0_u0_n644 ), .A2(_AES_ENC_u0_u0_n643 ), .A3(_AES_ENC_u0_u0_n804 ), .A4(_AES_ENC_u0_u0_n642 ), .ZN(_AES_ENC_u0_u0_n645 ) );
NOR2_X2 _AES_ENC_u0_u0_U428  ( .A1(_AES_ENC_u0_u0_n1102 ), .A2(_AES_ENC_u0_u0_n910 ), .ZN(_AES_ENC_u0_u0_n932 ) );
NOR3_X2 _AES_ENC_u0_u0_U427  ( .A1(_AES_ENC_u0_u0_n623 ), .A2(_AES_ENC_w3[17] ), .A3(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n683 ) );
NOR2_X2 _AES_ENC_u0_u0_U421  ( .A1(_AES_ENC_u0_u0_n1102 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n755 ) );
INV_X4 _AES_ENC_u0_u0_U420  ( .A(_AES_ENC_u0_u0_n931 ), .ZN(_AES_ENC_u0_u0_n623 ) );
NOR2_X2 _AES_ENC_u0_u0_U419  ( .A1(_AES_ENC_u0_u0_n996 ), .A2(_AES_ENC_u0_u0_n931 ), .ZN(_AES_ENC_u0_u0_n704 ) );
NOR2_X2 _AES_ENC_u0_u0_U418  ( .A1(_AES_ENC_u0_u0_n1029 ), .A2(_AES_ENC_u0_u0_n1025 ), .ZN(_AES_ENC_u0_u0_n1079 ) );
NOR3_X2 _AES_ENC_u0_u0_U417  ( .A1(_AES_ENC_u0_u0_n589 ), .A2(_AES_ENC_u0_u0_n1025 ), .A3(_AES_ENC_u0_u0_n616 ), .ZN(_AES_ENC_u0_u0_n945 ) );
NOR2_X2 _AES_ENC_u0_u0_U416  ( .A1(_AES_ENC_u0_u0_n1072 ), .A2(_AES_ENC_u0_u0_n1094 ), .ZN(_AES_ENC_u0_u0_n930 ) );
NOR2_X2 _AES_ENC_u0_u0_U415  ( .A1(_AES_ENC_u0_u0_n931 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n743 ) );
NOR2_X2 _AES_ENC_u0_u0_U414  ( .A1(_AES_ENC_u0_u0_n931 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n685 ) );
NOR3_X2 _AES_ENC_u0_u0_U413  ( .A1(_AES_ENC_u0_u0_n610 ), .A2(_AES_ENC_u0_u0_n572 ), .A3(_AES_ENC_u0_u0_n575 ), .ZN(_AES_ENC_u0_u0_n962 ) );
NOR2_X2 _AES_ENC_u0_u0_U410  ( .A1(_AES_ENC_u0_u0_n626 ), .A2(_AES_ENC_u0_u0_n611 ), .ZN(_AES_ENC_u0_u0_n800 ) );
NOR3_X2 _AES_ENC_u0_u0_U409  ( .A1(_AES_ENC_u0_u0_n590 ), .A2(_AES_ENC_u0_u0_n627 ), .A3(_AES_ENC_u0_u0_n611 ), .ZN(_AES_ENC_u0_u0_n798 ) );
NOR3_X2 _AES_ENC_u0_u0_U406  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n572 ), .A3(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n694 ) );
NOR4_X2 _AES_ENC_u0_u0_U405  ( .A1(_AES_ENC_u0_u0_n946 ), .A2(_AES_ENC_u0_u0_n1046 ), .A3(_AES_ENC_u0_u0_n671 ), .A4(_AES_ENC_u0_u0_n670 ), .ZN(_AES_ENC_u0_u0_n672 ) );
NOR4_X2 _AES_ENC_u0_u0_U404  ( .A1(_AES_ENC_u0_u0_n806 ), .A2(_AES_ENC_u0_u0_n805 ), .A3(_AES_ENC_u0_u0_n804 ), .A4(_AES_ENC_u0_u0_n803 ), .ZN(_AES_ENC_u0_u0_n807 ) );
NOR3_X2 _AES_ENC_u0_u0_U403  ( .A1(_AES_ENC_u0_u0_n799 ), .A2(_AES_ENC_u0_u0_n798 ), .A3(_AES_ENC_u0_u0_n797 ), .ZN(_AES_ENC_u0_u0_n808 ) );
NOR3_X2 _AES_ENC_u0_u0_U401  ( .A1(_AES_ENC_u0_u0_n1101 ), .A2(_AES_ENC_u0_u0_n1100 ), .A3(_AES_ENC_u0_u0_n1099 ), .ZN(_AES_ENC_u0_u0_n1109 ) );
NOR2_X2 _AES_ENC_u0_u0_U400  ( .A1(_AES_ENC_u0_u0_n641 ), .A2(_AES_ENC_u0_u0_n640 ), .ZN(_AES_ENC_u0_u0_n646 ) );
NOR3_X2 _AES_ENC_u0_u0_U399  ( .A1(_AES_ENC_u0_u0_n743 ), .A2(_AES_ENC_u0_u0_n742 ), .A3(_AES_ENC_u0_u0_n741 ), .ZN(_AES_ENC_u0_u0_n744 ) );
NOR2_X2 _AES_ENC_u0_u0_U398  ( .A1(_AES_ENC_u0_u0_n697 ), .A2(_AES_ENC_u0_u0_n658 ), .ZN(_AES_ENC_u0_u0_n659 ) );
NOR3_X2 _AES_ENC_u0_u0_U397  ( .A1(_AES_ENC_u0_u0_n959 ), .A2(_AES_ENC_u0_u0_n572 ), .A3(_AES_ENC_u0_u0_n609 ), .ZN(_AES_ENC_u0_u0_n768 ) );
NOR2_X2 _AES_ENC_u0_u0_U396  ( .A1(_AES_ENC_u0_u0_n891 ), .A2(_AES_ENC_u0_u0_n609 ), .ZN(_AES_ENC_u0_u0_n894 ) );
NOR3_X2 _AES_ENC_u0_u0_U393  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n572 ), .A3(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n895 ) );
NOR3_X2 _AES_ENC_u0_u0_U390  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n1056 ), .A3(_AES_ENC_u0_u0_n990 ), .ZN(_AES_ENC_u0_u0_n896 ) );
NOR4_X2 _AES_ENC_u0_u0_U389  ( .A1(_AES_ENC_u0_u0_n896 ), .A2(_AES_ENC_u0_u0_n895 ), .A3(_AES_ENC_u0_u0_n894 ), .A4(_AES_ENC_u0_u0_n893 ), .ZN(_AES_ENC_u0_u0_n897 ) );
NOR2_X2 _AES_ENC_u0_u0_U388  ( .A1(_AES_ENC_u0_u0_n598 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n885 ) );
NOR2_X2 _AES_ENC_u0_u0_U387  ( .A1(_AES_ENC_u0_u0_n623 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n882 ) );
NOR2_X2 _AES_ENC_u0_u0_U386  ( .A1(_AES_ENC_u0_u0_n1053 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n884 ) );
NOR4_X2 _AES_ENC_u0_u0_U385  ( .A1(_AES_ENC_u0_u0_n885 ), .A2(_AES_ENC_u0_u0_n884 ), .A3(_AES_ENC_u0_u0_n883 ), .A4(_AES_ENC_u0_u0_n882 ), .ZN(_AES_ENC_u0_u0_n886 ) );
NOR2_X2 _AES_ENC_u0_u0_U384  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n569 ), .ZN(_AES_ENC_u0_u0_n947 ) );
NOR2_X2 _AES_ENC_u0_u0_U383  ( .A1(_AES_ENC_u0_u0_n572 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n949 ) );
NOR2_X2 _AES_ENC_u0_u0_U382  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n602 ), .ZN(_AES_ENC_u0_u0_n950 ) );
NOR4_X2 _AES_ENC_u0_u0_U374  ( .A1(_AES_ENC_u0_u0_n950 ), .A2(_AES_ENC_u0_u0_n949 ), .A3(_AES_ENC_u0_u0_n948 ), .A4(_AES_ENC_u0_u0_n947 ), .ZN(_AES_ENC_u0_u0_n951 ) );
NOR2_X2 _AES_ENC_u0_u0_U373  ( .A1(_AES_ENC_u0_u0_n1078 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n1033 ) );
NOR2_X2 _AES_ENC_u0_u0_U372  ( .A1(_AES_ENC_u0_u0_n1031 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n1032 ) );
NOR3_X2 _AES_ENC_u0_u0_U370  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n1025 ), .A3(_AES_ENC_u0_u0_n1074 ), .ZN(_AES_ENC_u0_u0_n1035 ) );
NOR4_X2 _AES_ENC_u0_u0_U369  ( .A1(_AES_ENC_u0_u0_n1035 ), .A2(_AES_ENC_u0_u0_n1034 ), .A3(_AES_ENC_u0_u0_n1033 ), .A4(_AES_ENC_u0_u0_n1032 ), .ZN(_AES_ENC_u0_u0_n1036 ) );
NOR2_X2 _AES_ENC_u0_u0_U368  ( .A1(_AES_ENC_u0_u0_n825 ), .A2(_AES_ENC_u0_u0_n578 ), .ZN(_AES_ENC_u0_u0_n830 ) );
NOR2_X2 _AES_ENC_u0_u0_U367  ( .A1(_AES_ENC_u0_u0_n827 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n829 ) );
NOR2_X2 _AES_ENC_u0_u0_U366  ( .A1(_AES_ENC_u0_u0_n572 ), .A2(_AES_ENC_u0_u0_n579 ), .ZN(_AES_ENC_u0_u0_n828 ) );
NOR4_X2 _AES_ENC_u0_u0_U365  ( .A1(_AES_ENC_u0_u0_n831 ), .A2(_AES_ENC_u0_u0_n830 ), .A3(_AES_ENC_u0_u0_n829 ), .A4(_AES_ENC_u0_u0_n828 ), .ZN(_AES_ENC_u0_u0_n832 ) );
NOR2_X2 _AES_ENC_u0_u0_U364  ( .A1(_AES_ENC_u0_u0_n598 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n1107 ) );
NOR2_X2 _AES_ENC_u0_u0_U363  ( .A1(_AES_ENC_u0_u0_n1102 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n1106 ) );
NOR2_X2 _AES_ENC_u0_u0_U354  ( .A1(_AES_ENC_u0_u0_n1103 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n1105 ) );
NOR4_X2 _AES_ENC_u0_u0_U353  ( .A1(_AES_ENC_u0_u0_n1107 ), .A2(_AES_ENC_u0_u0_n1106 ), .A3(_AES_ENC_u0_u0_n1105 ), .A4(_AES_ENC_u0_u0_n1104 ), .ZN(_AES_ENC_u0_u0_n1108 ) );
NOR3_X2 _AES_ENC_u0_u0_U352  ( .A1(_AES_ENC_u0_u0_n959 ), .A2(_AES_ENC_u0_u0_n621 ), .A3(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n963 ) );
NOR2_X2 _AES_ENC_u0_u0_U351  ( .A1(_AES_ENC_u0_u0_n626 ), .A2(_AES_ENC_u0_u0_n627 ), .ZN(_AES_ENC_u0_u0_n1114 ) );
NOR3_X2 _AES_ENC_u0_u0_U350  ( .A1(_AES_ENC_u0_u0_n910 ), .A2(_AES_ENC_u0_u0_n1059 ), .A3(_AES_ENC_u0_u0_n611 ), .ZN(_AES_ENC_u0_u0_n1115 ) );
INV_X4 _AES_ENC_u0_u0_U349  ( .A(_AES_ENC_u0_u0_n1024 ), .ZN(_AES_ENC_u0_u0_n606 ) );
INV_X4 _AES_ENC_u0_u0_U348  ( .A(_AES_ENC_u0_u0_n1094 ), .ZN(_AES_ENC_u0_u0_n613 ) );
NOR2_X2 _AES_ENC_u0_u0_U347  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n931 ), .ZN(_AES_ENC_u0_u0_n1100 ) );
NOR2_X2 _AES_ENC_u0_u0_U346  ( .A1(_AES_ENC_u0_u0_n569 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n929 ) );
NOR2_X2 _AES_ENC_u0_u0_U345  ( .A1(_AES_ENC_u0_u0_n620 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n926 ) );
INV_X4 _AES_ENC_u0_u0_U338  ( .A(_AES_ENC_u0_u0_n1093 ), .ZN(_AES_ENC_u0_u0_n617 ) );
NOR2_X2 _AES_ENC_u0_u0_U335  ( .A1(_AES_ENC_u0_u0_n572 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n1095 ) );
NOR2_X2 _AES_ENC_u0_u0_U329  ( .A1(_AES_ENC_u0_u0_n609 ), .A2(_AES_ENC_u0_u0_n627 ), .ZN(_AES_ENC_u0_u0_n1010 ) );
NOR2_X2 _AES_ENC_u0_u0_U328  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n1103 ) );
NOR2_X2 _AES_ENC_u0_u0_U327  ( .A1(_AES_ENC_w3[17] ), .A2(_AES_ENC_u0_u0_n1120 ), .ZN(_AES_ENC_u0_u0_n1022 ) );
NOR2_X2 _AES_ENC_u0_u0_U325  ( .A1(_AES_ENC_u0_u0_n619 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n911 ) );
NOR2_X2 _AES_ENC_u0_u0_U324  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_u0_u0_n1025 ), .ZN(_AES_ENC_u0_u0_n826 ) );
NOR2_X2 _AES_ENC_u0_u0_U319  ( .A1(_AES_ENC_u0_u0_n626 ), .A2(_AES_ENC_u0_u0_n607 ), .ZN(_AES_ENC_u0_u0_n1072 ) );
NOR2_X2 _AES_ENC_u0_u0_U318  ( .A1(_AES_ENC_u0_u0_n627 ), .A2(_AES_ENC_u0_u0_n616 ), .ZN(_AES_ENC_u0_u0_n956 ) );
NOR2_X2 _AES_ENC_u0_u0_U317  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_u0_u0_n624 ), .ZN(_AES_ENC_u0_u0_n1121 ) );
NOR2_X2 _AES_ENC_u0_u0_U316  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_u0_u0_n624 ), .ZN(_AES_ENC_u0_u0_n1058 ) );
NOR2_X2 _AES_ENC_u0_u0_U315  ( .A1(_AES_ENC_u0_u0_n625 ), .A2(_AES_ENC_u0_u0_n611 ), .ZN(_AES_ENC_u0_u0_n1073 ) );
NOR2_X2 _AES_ENC_u0_u0_U314  ( .A1(_AES_ENC_w3[17] ), .A2(_AES_ENC_u0_u0_n1025 ), .ZN(_AES_ENC_u0_u0_n1054 ) );
NOR2_X2 _AES_ENC_u0_u0_U312  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_u0_u0_n931 ), .ZN(_AES_ENC_u0_u0_n1029 ) );
NOR2_X2 _AES_ENC_u0_u0_U311  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n1056 ) );
NOR2_X2 _AES_ENC_u0_u0_U310  ( .A1(_AES_ENC_u0_u0_n614 ), .A2(_AES_ENC_u0_u0_n626 ), .ZN(_AES_ENC_u0_u0_n1050 ) );
NOR2_X2 _AES_ENC_u0_u0_U309  ( .A1(_AES_ENC_u0_u0_n1121 ), .A2(_AES_ENC_u0_u0_n1025 ), .ZN(_AES_ENC_u0_u0_n1120 ) );
NOR2_X2 _AES_ENC_u0_u0_U303  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_u0_u0_n572 ), .ZN(_AES_ENC_u0_u0_n1074 ) );
NOR2_X2 _AES_ENC_u0_u0_U302  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n584 ), .ZN(_AES_ENC_u0_u0_n838 ) );
NOR2_X2 _AES_ENC_u0_u0_U300  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n602 ), .ZN(_AES_ENC_u0_u0_n837 ) );
NOR2_X2 _AES_ENC_u0_u0_U299  ( .A1(_AES_ENC_u0_u0_n838 ), .A2(_AES_ENC_u0_u0_n837 ), .ZN(_AES_ENC_u0_u0_n845 ) );
NOR2_X2 _AES_ENC_u0_u0_U298  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n1071 ), .ZN(_AES_ENC_u0_u0_n669 ) );
NOR2_X2 _AES_ENC_u0_u0_U297  ( .A1(_AES_ENC_u0_u0_n1095 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n668 ) );
NOR2_X2 _AES_ENC_u0_u0_U296  ( .A1(_AES_ENC_u0_u0_n669 ), .A2(_AES_ENC_u0_u0_n668 ), .ZN(_AES_ENC_u0_u0_n673 ) );
NOR2_X2 _AES_ENC_u0_u0_U295  ( .A1(_AES_ENC_u0_u0_n1058 ), .A2(_AES_ENC_u0_u0_n1054 ), .ZN(_AES_ENC_u0_u0_n878 ) );
NOR2_X2 _AES_ENC_u0_u0_U294  ( .A1(_AES_ENC_u0_u0_n878 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n879 ) );
NOR2_X2 _AES_ENC_u0_u0_U293  ( .A1(_AES_ENC_u0_u0_n880 ), .A2(_AES_ENC_u0_u0_n879 ), .ZN(_AES_ENC_u0_u0_n887 ) );
NOR3_X2 _AES_ENC_u0_u0_U292  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n1091 ), .A3(_AES_ENC_u0_u0_n1022 ), .ZN(_AES_ENC_u0_u0_n720 ) );
NOR3_X2 _AES_ENC_u0_u0_U291  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n1054 ), .A3(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n719 ) );
NOR2_X2 _AES_ENC_u0_u0_U290  ( .A1(_AES_ENC_u0_u0_n720 ), .A2(_AES_ENC_u0_u0_n719 ), .ZN(_AES_ENC_u0_u0_n726 ) );
NOR2_X2 _AES_ENC_u0_u0_U284  ( .A1(_AES_ENC_u0_u0_n576 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n866 ) );
NOR2_X2 _AES_ENC_u0_u0_U283  ( .A1(_AES_ENC_u0_u0_n614 ), .A2(_AES_ENC_u0_u0_n591 ), .ZN(_AES_ENC_u0_u0_n865 ) );
NOR2_X2 _AES_ENC_u0_u0_U282  ( .A1(_AES_ENC_u0_u0_n866 ), .A2(_AES_ENC_u0_u0_n865 ), .ZN(_AES_ENC_u0_u0_n872 ) );
NOR2_X2 _AES_ENC_u0_u0_U281  ( .A1(_AES_ENC_u0_u0_n1059 ), .A2(_AES_ENC_u0_u0_n1058 ), .ZN(_AES_ENC_u0_u0_n1060 ) );
NOR2_X2 _AES_ENC_u0_u0_U280  ( .A1(_AES_ENC_u0_u0_n911 ), .A2(_AES_ENC_u0_u0_n910 ), .ZN(_AES_ENC_u0_u0_n912 ) );
NOR2_X2 _AES_ENC_u0_u0_U279  ( .A1(_AES_ENC_u0_u0_n912 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n916 ) );
NOR2_X2 _AES_ENC_u0_u0_U273  ( .A1(_AES_ENC_u0_u0_n826 ), .A2(_AES_ENC_u0_u0_n573 ), .ZN(_AES_ENC_u0_u0_n750 ) );
NOR2_X2 _AES_ENC_u0_u0_U272  ( .A1(_AES_ENC_u0_u0_n750 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n751 ) );
NOR2_X2 _AES_ENC_u0_u0_U271  ( .A1(_AES_ENC_u0_u0_n907 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n908 ) );
NOR2_X2 _AES_ENC_u0_u0_U270  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n588 ), .ZN(_AES_ENC_u0_u0_n957 ) );
NOR2_X2 _AES_ENC_u0_u0_U269  ( .A1(_AES_ENC_u0_u0_n990 ), .A2(_AES_ENC_u0_u0_n926 ), .ZN(_AES_ENC_u0_u0_n780 ) );
NOR2_X2 _AES_ENC_u0_u0_U268  ( .A1(_AES_ENC_u0_u0_n1022 ), .A2(_AES_ENC_u0_u0_n1058 ), .ZN(_AES_ENC_u0_u0_n740 ) );
NOR2_X2 _AES_ENC_u0_u0_U267  ( .A1(_AES_ENC_u0_u0_n740 ), .A2(_AES_ENC_u0_u0_n616 ), .ZN(_AES_ENC_u0_u0_n742 ) );
NOR2_X2 _AES_ENC_u0_u0_U263  ( .A1(_AES_ENC_u0_u0_n1098 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n1099 ) );
NOR2_X2 _AES_ENC_u0_u0_U262  ( .A1(_AES_ENC_u0_u0_n1120 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n993 ) );
NOR2_X2 _AES_ENC_u0_u0_U258  ( .A1(_AES_ENC_u0_u0_n993 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n994 ) );
NOR2_X2 _AES_ENC_u0_u0_U255  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n620 ), .ZN(_AES_ENC_u0_u0_n1026 ) );
NOR2_X2 _AES_ENC_u0_u0_U254  ( .A1(_AES_ENC_u0_u0_n573 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n1027 ) );
NOR2_X2 _AES_ENC_u0_u0_U253  ( .A1(_AES_ENC_u0_u0_n1027 ), .A2(_AES_ENC_u0_u0_n1026 ), .ZN(_AES_ENC_u0_u0_n1028 ) );
NOR2_X2 _AES_ENC_u0_u0_U252  ( .A1(_AES_ENC_u0_u0_n1029 ), .A2(_AES_ENC_u0_u0_n1028 ), .ZN(_AES_ENC_u0_u0_n1034 ) );
NOR2_X2 _AES_ENC_u0_u0_U251  ( .A1(_AES_ENC_u0_u0_n1056 ), .A2(_AES_ENC_u0_u0_n990 ), .ZN(_AES_ENC_u0_u0_n991 ) );
NOR2_X2 _AES_ENC_u0_u0_U250  ( .A1(_AES_ENC_u0_u0_n991 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n995 ) );
NOR2_X2 _AES_ENC_u0_u0_U243  ( .A1(_AES_ENC_u0_u0_n603 ), .A2(_AES_ENC_u0_u0_n610 ), .ZN(_AES_ENC_u0_u0_n1006 ) );
NOR2_X2 _AES_ENC_u0_u0_U242  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n577 ), .ZN(_AES_ENC_u0_u0_n1007 ) );
NOR2_X2 _AES_ENC_u0_u0_U241  ( .A1(_AES_ENC_u0_u0_n607 ), .A2(_AES_ENC_u0_u0_n590 ), .ZN(_AES_ENC_u0_u0_n1008 ) );
NOR3_X2 _AES_ENC_u0_u0_U240  ( .A1(_AES_ENC_u0_u0_n1008 ), .A2(_AES_ENC_u0_u0_n1007 ), .A3(_AES_ENC_u0_u0_n1006 ), .ZN(_AES_ENC_u0_u0_n1018 ) );
NOR2_X2 _AES_ENC_u0_u0_U239  ( .A1(_AES_ENC_u0_u0_n606 ), .A2(_AES_ENC_u0_u0_n906 ), .ZN(_AES_ENC_u0_u0_n741 ) );
NOR2_X2 _AES_ENC_u0_u0_U238  ( .A1(_AES_ENC_u0_u0_n1054 ), .A2(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n763 ) );
NOR2_X2 _AES_ENC_u0_u0_U237  ( .A1(_AES_ENC_u0_u0_n763 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n769 ) );
NOR2_X2 _AES_ENC_u0_u0_U236  ( .A1(_AES_ENC_u0_u0_n839 ), .A2(_AES_ENC_u0_u0_n582 ), .ZN(_AES_ENC_u0_u0_n693 ) );
NOR2_X2 _AES_ENC_u0_u0_U235  ( .A1(_AES_ENC_u0_u0_n609 ), .A2(_AES_ENC_u0_u0_n580 ), .ZN(_AES_ENC_u0_u0_n1123 ) );
NOR2_X2 _AES_ENC_u0_u0_U234  ( .A1(_AES_ENC_u0_u0_n780 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n784 ) );
NOR2_X2 _AES_ENC_u0_u0_U229  ( .A1(_AES_ENC_u0_u0_n1117 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n782 ) );
NOR2_X2 _AES_ENC_u0_u0_U228  ( .A1(_AES_ENC_u0_u0_n781 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n783 ) );
NOR4_X2 _AES_ENC_u0_u0_U227  ( .A1(_AES_ENC_u0_u0_n880 ), .A2(_AES_ENC_u0_u0_n784 ), .A3(_AES_ENC_u0_u0_n783 ), .A4(_AES_ENC_u0_u0_n782 ), .ZN(_AES_ENC_u0_u0_n785 ) );
INV_X4 _AES_ENC_u0_u0_U226  ( .A(_AES_ENC_u0_u0_n1029 ), .ZN(_AES_ENC_u0_u0_n582 ) );
NOR2_X2 _AES_ENC_u0_u0_U225  ( .A1(_AES_ENC_u0_u0_n593 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n1125 ) );
NOR2_X2 _AES_ENC_u0_u0_U223  ( .A1(_AES_ENC_u0_u0_n616 ), .A2(_AES_ENC_u0_u0_n580 ), .ZN(_AES_ENC_u0_u0_n771 ) );
NOR2_X2 _AES_ENC_u0_u0_U222  ( .A1(_AES_ENC_u0_u0_n616 ), .A2(_AES_ENC_u0_u0_n597 ), .ZN(_AES_ENC_u0_u0_n883 ) );
NOR2_X2 _AES_ENC_u0_u0_U221  ( .A1(_AES_ENC_u0_u0_n990 ), .A2(_AES_ENC_u0_u0_n929 ), .ZN(_AES_ENC_u0_u0_n892 ) );
NOR2_X2 _AES_ENC_u0_u0_U217  ( .A1(_AES_ENC_u0_u0_n892 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n893 ) );
NOR2_X2 _AES_ENC_u0_u0_U213  ( .A1(_AES_ENC_u0_u0_n910 ), .A2(_AES_ENC_u0_u0_n1056 ), .ZN(_AES_ENC_u0_u0_n941 ) );
NOR2_X2 _AES_ENC_u0_u0_U212  ( .A1(_AES_ENC_u0_u0_n623 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n630 ) );
NOR2_X2 _AES_ENC_u0_u0_U211  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n602 ), .ZN(_AES_ENC_u0_u0_n806 ) );
NOR2_X2 _AES_ENC_u0_u0_U210  ( .A1(_AES_ENC_u0_u0_n623 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n948 ) );
NOR2_X2 _AES_ENC_u0_u0_U209  ( .A1(_AES_ENC_u0_u0_n606 ), .A2(_AES_ENC_u0_u0_n582 ), .ZN(_AES_ENC_u0_u0_n1104 ) );
NOR2_X2 _AES_ENC_u0_u0_U208  ( .A1(_AES_ENC_u0_u0_n1121 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n1122 ) );
NOR2_X2 _AES_ENC_u0_u0_U207  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n1023 ), .ZN(_AES_ENC_u0_u0_n756 ) );
NOR2_X2 _AES_ENC_u0_u0_U201  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n602 ), .ZN(_AES_ENC_u0_u0_n870 ) );
NOR2_X2 _AES_ENC_u0_u0_U200  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n589 ), .ZN(_AES_ENC_u0_u0_n868 ) );
NOR2_X2 _AES_ENC_u0_u0_U199  ( .A1(_AES_ENC_u0_u0_n1120 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n1124 ) );
NOR2_X2 _AES_ENC_u0_u0_U198  ( .A1(_AES_ENC_u0_u0_n1120 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n696 ) );
NOR2_X2 _AES_ENC_u0_u0_U197  ( .A1(_AES_ENC_u0_u0_n1074 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n1076 ) );
NOR2_X2 _AES_ENC_u0_u0_U196  ( .A1(_AES_ENC_u0_u0_n1074 ), .A2(_AES_ENC_u0_u0_n620 ), .ZN(_AES_ENC_u0_u0_n781 ) );
NOR3_X2 _AES_ENC_u0_u0_U195  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n1056 ), .A3(_AES_ENC_u0_u0_n990 ), .ZN(_AES_ENC_u0_u0_n979 ) );
NOR3_X2 _AES_ENC_u0_u0_U194  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n1058 ), .A3(_AES_ENC_u0_u0_n1059 ), .ZN(_AES_ENC_u0_u0_n854 ) );
NOR2_X2 _AES_ENC_u0_u0_U187  ( .A1(_AES_ENC_u0_u0_n996 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n869 ) );
NOR2_X2 _AES_ENC_u0_u0_U186  ( .A1(_AES_ENC_u0_u0_n1056 ), .A2(_AES_ENC_u0_u0_n1074 ), .ZN(_AES_ENC_u0_u0_n1057 ) );
NOR3_X2 _AES_ENC_u0_u0_U185  ( .A1(_AES_ENC_u0_u0_n607 ), .A2(_AES_ENC_u0_u0_n1120 ), .A3(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n978 ) );
NOR2_X2 _AES_ENC_u0_u0_U184  ( .A1(_AES_ENC_u0_u0_n996 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n998 ) );
NOR2_X2 _AES_ENC_u0_u0_U183  ( .A1(_AES_ENC_u0_u0_n996 ), .A2(_AES_ENC_u0_u0_n911 ), .ZN(_AES_ENC_u0_u0_n1116 ) );
NOR2_X2 _AES_ENC_u0_u0_U182  ( .A1(_AES_ENC_u0_u0_n1074 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n754 ) );
NOR2_X2 _AES_ENC_u0_u0_U181  ( .A1(_AES_ENC_u0_u0_n926 ), .A2(_AES_ENC_u0_u0_n1103 ), .ZN(_AES_ENC_u0_u0_n977 ) );
NOR2_X2 _AES_ENC_u0_u0_U180  ( .A1(_AES_ENC_u0_u0_n839 ), .A2(_AES_ENC_u0_u0_n824 ), .ZN(_AES_ENC_u0_u0_n1092 ) );
NOR2_X2 _AES_ENC_u0_u0_U174  ( .A1(_AES_ENC_u0_u0_n573 ), .A2(_AES_ENC_u0_u0_n1074 ), .ZN(_AES_ENC_u0_u0_n684 ) );
NOR2_X2 _AES_ENC_u0_u0_U173  ( .A1(_AES_ENC_u0_u0_n826 ), .A2(_AES_ENC_u0_u0_n1059 ), .ZN(_AES_ENC_u0_u0_n907 ) );
NOR3_X2 _AES_ENC_u0_u0_U172  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n573 ), .A3(_AES_ENC_u0_u0_n1074 ), .ZN(_AES_ENC_u0_u0_n641 ) );
NOR3_X2 _AES_ENC_u0_u0_U171  ( .A1(_AES_ENC_u0_u0_n625 ), .A2(_AES_ENC_u0_u0_n1115 ), .A3(_AES_ENC_u0_u0_n585 ), .ZN(_AES_ENC_u0_u0_n831 ) );
NOR3_X2 _AES_ENC_u0_u0_U170  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n573 ), .A3(_AES_ENC_u0_u0_n1013 ), .ZN(_AES_ENC_u0_u0_n670 ) );
NOR2_X2 _AES_ENC_u0_u0_U169  ( .A1(_AES_ENC_u0_u0_n1029 ), .A2(_AES_ENC_u0_u0_n1095 ), .ZN(_AES_ENC_u0_u0_n735 ) );
NOR2_X2 _AES_ENC_u0_u0_U168  ( .A1(_AES_ENC_u0_u0_n1100 ), .A2(_AES_ENC_u0_u0_n854 ), .ZN(_AES_ENC_u0_u0_n860 ) );
NAND3_X2 _AES_ENC_u0_u0_U162  ( .A1(_AES_ENC_u0_u0_n569 ), .A2(_AES_ENC_u0_u0_n582 ), .A3(_AES_ENC_u0_u0_n681 ), .ZN(_AES_ENC_u0_u0_n691 ) );
NOR2_X2 _AES_ENC_u0_u0_U161  ( .A1(_AES_ENC_u0_u0_n683 ), .A2(_AES_ENC_u0_u0_n682 ), .ZN(_AES_ENC_u0_u0_n690 ) );
NOR4_X2 _AES_ENC_u0_u0_U160  ( .A1(_AES_ENC_u0_u0_n963 ), .A2(_AES_ENC_u0_u0_n962 ), .A3(_AES_ENC_u0_u0_n961 ), .A4(_AES_ENC_u0_u0_n960 ), .ZN(_AES_ENC_u0_u0_n964 ) );
NOR2_X2 _AES_ENC_u0_u0_U159  ( .A1(_AES_ENC_u0_u0_n958 ), .A2(_AES_ENC_u0_u0_n957 ), .ZN(_AES_ENC_u0_u0_n965 ) );
NOR4_X2 _AES_ENC_u0_u0_U158  ( .A1(_AES_ENC_u0_u0_n983 ), .A2(_AES_ENC_u0_u0_n982 ), .A3(_AES_ENC_u0_u0_n981 ), .A4(_AES_ENC_u0_u0_n980 ), .ZN(_AES_ENC_u0_u0_n984 ) );
NOR2_X2 _AES_ENC_u0_u0_U157  ( .A1(_AES_ENC_u0_u0_n979 ), .A2(_AES_ENC_u0_u0_n978 ), .ZN(_AES_ENC_u0_u0_n985 ) );
NOR3_X2 _AES_ENC_u0_u0_U156  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n1054 ), .A3(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n961 ) );
NOR3_X2 _AES_ENC_u0_u0_U155  ( .A1(_AES_ENC_u0_u0_n620 ), .A2(_AES_ENC_u0_u0_n1074 ), .A3(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n671 ) );
NOR2_X2 _AES_ENC_u0_u0_U154  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n1077 ), .ZN(_AES_ENC_u0_u0_n1084 ) );
NOR2_X2 _AES_ENC_u0_u0_U153  ( .A1(_AES_ENC_u0_u0_n1079 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n1082 ) );
NOR2_X2 _AES_ENC_u0_u0_U152  ( .A1(_AES_ENC_u0_u0_n1078 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n1083 ) );
NOR4_X2 _AES_ENC_u0_u0_U143  ( .A1(_AES_ENC_u0_u0_n1084 ), .A2(_AES_ENC_u0_u0_n1083 ), .A3(_AES_ENC_u0_u0_n1082 ), .A4(_AES_ENC_u0_u0_n1081 ), .ZN(_AES_ENC_u0_u0_n1085 ) );
NOR2_X2 _AES_ENC_u0_u0_U142  ( .A1(_AES_ENC_u0_u0_n1057 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n1062 ) );
NOR2_X2 _AES_ENC_u0_u0_U141  ( .A1(_AES_ENC_u0_u0_n1060 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n1061 ) );
NOR2_X2 _AES_ENC_u0_u0_U140  ( .A1(_AES_ENC_u0_u0_n1055 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n1063 ) );
NOR4_X2 _AES_ENC_u0_u0_U132  ( .A1(_AES_ENC_u0_u0_n1064 ), .A2(_AES_ENC_u0_u0_n1063 ), .A3(_AES_ENC_u0_u0_n1062 ), .A4(_AES_ENC_u0_u0_n1061 ), .ZN(_AES_ENC_u0_u0_n1065 ) );
NOR2_X2 _AES_ENC_u0_u0_U131  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n582 ), .ZN(_AES_ENC_u0_u0_n770 ) );
NOR2_X2 _AES_ENC_u0_u0_U130  ( .A1(_AES_ENC_u0_u0_n1103 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n772 ) );
NOR2_X2 _AES_ENC_u0_u0_U129  ( .A1(_AES_ENC_u0_u0_n610 ), .A2(_AES_ENC_u0_u0_n599 ), .ZN(_AES_ENC_u0_u0_n773 ) );
NOR4_X2 _AES_ENC_u0_u0_U128  ( .A1(_AES_ENC_u0_u0_n773 ), .A2(_AES_ENC_u0_u0_n772 ), .A3(_AES_ENC_u0_u0_n771 ), .A4(_AES_ENC_u0_u0_n770 ), .ZN(_AES_ENC_u0_u0_n774 ) );
NOR3_X2 _AES_ENC_u0_u0_U127  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n1091 ), .A3(_AES_ENC_u0_u0_n1022 ), .ZN(_AES_ENC_u0_u0_n843 ) );
NOR2_X2 _AES_ENC_u0_u0_U126  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n1077 ), .ZN(_AES_ENC_u0_u0_n841 ) );
NOR2_X2 _AES_ENC_u0_u0_U121  ( .A1(_AES_ENC_u0_u0_n1120 ), .A2(_AES_ENC_u0_u0_n839 ), .ZN(_AES_ENC_u0_u0_n842 ) );
NOR4_X2 _AES_ENC_u0_u0_U120  ( .A1(_AES_ENC_u0_u0_n843 ), .A2(_AES_ENC_u0_u0_n842 ), .A3(_AES_ENC_u0_u0_n841 ), .A4(_AES_ENC_u0_u0_n840 ), .ZN(_AES_ENC_u0_u0_n844 ) );
NOR2_X2 _AES_ENC_u0_u0_U119  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n595 ), .ZN(_AES_ENC_u0_u0_n858 ) );
NOR2_X2 _AES_ENC_u0_u0_U118  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n855 ), .ZN(_AES_ENC_u0_u0_n857 ) );
NOR2_X2 _AES_ENC_u0_u0_U117  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n587 ), .ZN(_AES_ENC_u0_u0_n856 ) );
NOR4_X2 _AES_ENC_u0_u0_U116  ( .A1(_AES_ENC_u0_u0_n858 ), .A2(_AES_ENC_u0_u0_n857 ), .A3(_AES_ENC_u0_u0_n856 ), .A4(_AES_ENC_u0_u0_n958 ), .ZN(_AES_ENC_u0_u0_n859 ) );
NOR3_X2 _AES_ENC_u0_u0_U115  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n1120 ), .A3(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n918 ) );
NOR2_X2 _AES_ENC_u0_u0_U106  ( .A1(_AES_ENC_u0_u0_n914 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n915 ) );
NOR3_X2 _AES_ENC_u0_u0_U105  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n573 ), .A3(_AES_ENC_u0_u0_n1013 ), .ZN(_AES_ENC_u0_u0_n917 ) );
NOR4_X2 _AES_ENC_u0_u0_U104  ( .A1(_AES_ENC_u0_u0_n918 ), .A2(_AES_ENC_u0_u0_n917 ), .A3(_AES_ENC_u0_u0_n916 ), .A4(_AES_ENC_u0_u0_n915 ), .ZN(_AES_ENC_u0_u0_n919 ) );
NOR2_X2 _AES_ENC_u0_u0_U103  ( .A1(_AES_ENC_u0_u0_n735 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n687 ) );
NOR2_X2 _AES_ENC_u0_u0_U102  ( .A1(_AES_ENC_u0_u0_n684 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n688 ) );
NOR2_X2 _AES_ENC_u0_u0_U101  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n600 ), .ZN(_AES_ENC_u0_u0_n686 ) );
NOR4_X2 _AES_ENC_u0_u0_U100  ( .A1(_AES_ENC_u0_u0_n688 ), .A2(_AES_ENC_u0_u0_n687 ), .A3(_AES_ENC_u0_u0_n686 ), .A4(_AES_ENC_u0_u0_n685 ), .ZN(_AES_ENC_u0_u0_n689 ) );
NOR2_X2 _AES_ENC_u0_u0_U95  ( .A1(_AES_ENC_u0_u0_n583 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n814 ) );
NOR3_X2 _AES_ENC_u0_u0_U94  ( .A1(_AES_ENC_u0_u0_n606 ), .A2(_AES_ENC_u0_u0_n1058 ), .A3(_AES_ENC_u0_u0_n1059 ), .ZN(_AES_ENC_u0_u0_n815 ) );
NOR2_X2 _AES_ENC_u0_u0_U93  ( .A1(_AES_ENC_u0_u0_n907 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n813 ) );
NOR4_X2 _AES_ENC_u0_u0_U92  ( .A1(_AES_ENC_u0_u0_n815 ), .A2(_AES_ENC_u0_u0_n814 ), .A3(_AES_ENC_u0_u0_n813 ), .A4(_AES_ENC_u0_u0_n812 ), .ZN(_AES_ENC_u0_u0_n816 ) );
NOR2_X2 _AES_ENC_u0_u0_U91  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n881 ), .ZN(_AES_ENC_u0_u0_n711 ) );
NOR2_X2 _AES_ENC_u0_u0_U90  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n855 ), .ZN(_AES_ENC_u0_u0_n709 ) );
NOR2_X2 _AES_ENC_u0_u0_U89  ( .A1(_AES_ENC_u0_u0_n609 ), .A2(_AES_ENC_u0_u0_n590 ), .ZN(_AES_ENC_u0_u0_n710 ) );
NOR4_X2 _AES_ENC_u0_u0_U88  ( .A1(_AES_ENC_u0_u0_n711 ), .A2(_AES_ENC_u0_u0_n710 ), .A3(_AES_ENC_u0_u0_n709 ), .A4(_AES_ENC_u0_u0_n708 ), .ZN(_AES_ENC_u0_u0_n712 ) );
NOR2_X2 _AES_ENC_u0_u0_U87  ( .A1(_AES_ENC_u0_u0_n617 ), .A2(_AES_ENC_u0_u0_n569 ), .ZN(_AES_ENC_u0_u0_n721 ) );
NOR2_X2 _AES_ENC_u0_u0_U86  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n1096 ), .ZN(_AES_ENC_u0_u0_n722 ) );
NOR2_X2 _AES_ENC_u0_u0_U81  ( .A1(_AES_ENC_u0_u0_n1031 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n723 ) );
NOR4_X2 _AES_ENC_u0_u0_U80  ( .A1(_AES_ENC_u0_u0_n724 ), .A2(_AES_ENC_u0_u0_n723 ), .A3(_AES_ENC_u0_u0_n722 ), .A4(_AES_ENC_u0_u0_n721 ), .ZN(_AES_ENC_u0_u0_n725 ) );
NOR2_X2 _AES_ENC_u0_u0_U79  ( .A1(_AES_ENC_u0_u0_n911 ), .A2(_AES_ENC_u0_u0_n990 ), .ZN(_AES_ENC_u0_u0_n1009 ) );
NOR2_X2 _AES_ENC_u0_u0_U78  ( .A1(_AES_ENC_u0_u0_n1013 ), .A2(_AES_ENC_u0_u0_n573 ), .ZN(_AES_ENC_u0_u0_n1014 ) );
NOR2_X2 _AES_ENC_u0_u0_U74  ( .A1(_AES_ENC_u0_u0_n1014 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n1015 ) );
NOR4_X2 _AES_ENC_u0_u0_U73  ( .A1(_AES_ENC_u0_u0_n1016 ), .A2(_AES_ENC_u0_u0_n1015 ), .A3(_AES_ENC_u0_u0_n1119 ), .A4(_AES_ENC_u0_u0_n1046 ), .ZN(_AES_ENC_u0_u0_n1017 ) );
NOR2_X2 _AES_ENC_u0_u0_U72  ( .A1(_AES_ENC_u0_u0_n606 ), .A2(_AES_ENC_u0_u0_n589 ), .ZN(_AES_ENC_u0_u0_n997 ) );
NOR2_X2 _AES_ENC_u0_u0_U71  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n577 ), .ZN(_AES_ENC_u0_u0_n1000 ) );
NOR2_X2 _AES_ENC_u0_u0_U65  ( .A1(_AES_ENC_u0_u0_n616 ), .A2(_AES_ENC_u0_u0_n1096 ), .ZN(_AES_ENC_u0_u0_n999 ) );
NOR4_X2 _AES_ENC_u0_u0_U64  ( .A1(_AES_ENC_u0_u0_n1000 ), .A2(_AES_ENC_u0_u0_n999 ), .A3(_AES_ENC_u0_u0_n998 ), .A4(_AES_ENC_u0_u0_n997 ), .ZN(_AES_ENC_u0_u0_n1001 ) );
NOR2_X2 _AES_ENC_u0_u0_U63  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n1096 ), .ZN(_AES_ENC_u0_u0_n697 ) );
NOR2_X2 _AES_ENC_u0_u0_U62  ( .A1(_AES_ENC_u0_u0_n620 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n958 ) );
NOR2_X2 _AES_ENC_u0_u0_U61  ( .A1(_AES_ENC_u0_u0_n911 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n983 ) );
NOR2_X2 _AES_ENC_u0_u0_U59  ( .A1(_AES_ENC_u0_u0_n1054 ), .A2(_AES_ENC_u0_u0_n1103 ), .ZN(_AES_ENC_u0_u0_n1031 ) );
INV_X4 _AES_ENC_u0_u0_U58  ( .A(_AES_ENC_u0_u0_n1050 ), .ZN(_AES_ENC_u0_u0_n612 ) );
INV_X4 _AES_ENC_u0_u0_U57  ( .A(_AES_ENC_u0_u0_n1072 ), .ZN(_AES_ENC_u0_u0_n605 ) );
INV_X4 _AES_ENC_u0_u0_U50  ( .A(_AES_ENC_u0_u0_n1073 ), .ZN(_AES_ENC_u0_u0_n604 ) );
NOR2_X2 _AES_ENC_u0_u0_U49  ( .A1(_AES_ENC_u0_u0_n582 ), .A2(_AES_ENC_u0_u0_n613 ), .ZN(_AES_ENC_u0_u0_n880 ) );
NOR3_X2 _AES_ENC_u0_u0_U48  ( .A1(_AES_ENC_u0_u0_n826 ), .A2(_AES_ENC_u0_u0_n1121 ), .A3(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n946 ) );
INV_X4 _AES_ENC_u0_u0_U47  ( .A(_AES_ENC_u0_u0_n1010 ), .ZN(_AES_ENC_u0_u0_n608 ) );
NOR3_X2 _AES_ENC_u0_u0_U46  ( .A1(_AES_ENC_u0_u0_n573 ), .A2(_AES_ENC_u0_u0_n1029 ), .A3(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n1119 ) );
INV_X4 _AES_ENC_u0_u0_U45  ( .A(_AES_ENC_u0_u0_n956 ), .ZN(_AES_ENC_u0_u0_n615 ) );
NOR2_X2 _AES_ENC_u0_u0_U44  ( .A1(_AES_ENC_u0_u0_n623 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n1013 ) );
NOR2_X2 _AES_ENC_u0_u0_U43  ( .A1(_AES_ENC_u0_u0_n620 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n910 ) );
NOR2_X2 _AES_ENC_u0_u0_U42  ( .A1(_AES_ENC_u0_u0_n569 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n1091 ) );
NOR2_X2 _AES_ENC_u0_u0_U41  ( .A1(_AES_ENC_u0_u0_n622 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n990 ) );
NOR2_X2 _AES_ENC_u0_u0_U36  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_u0_u0_n1121 ), .ZN(_AES_ENC_u0_u0_n996 ) );
NOR2_X2 _AES_ENC_u0_u0_U35  ( .A1(_AES_ENC_u0_u0_n610 ), .A2(_AES_ENC_u0_u0_n600 ), .ZN(_AES_ENC_u0_u0_n628 ) );
NOR2_X2 _AES_ENC_u0_u0_U34  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n1117 ), .ZN(_AES_ENC_u0_u0_n1118 ) );
NOR2_X2 _AES_ENC_u0_u0_U33  ( .A1(_AES_ENC_u0_u0_n1119 ), .A2(_AES_ENC_u0_u0_n1118 ), .ZN(_AES_ENC_u0_u0_n1127 ) );
NOR2_X2 _AES_ENC_u0_u0_U32  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n594 ), .ZN(_AES_ENC_u0_u0_n629 ) );
NOR2_X2 _AES_ENC_u0_u0_U31  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n906 ), .ZN(_AES_ENC_u0_u0_n909 ) );
NOR2_X2 _AES_ENC_u0_u0_U30  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n597 ), .ZN(_AES_ENC_u0_u0_n658 ) );
NOR2_X2 _AES_ENC_u0_u0_U29  ( .A1(_AES_ENC_u0_u0_n1116 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n695 ) );
NOR2_X2 _AES_ENC_u0_u0_U24  ( .A1(_AES_ENC_u0_u0_n941 ), .A2(_AES_ENC_u0_u0_n608 ), .ZN(_AES_ENC_u0_u0_n724 ) );
NOR2_X2 _AES_ENC_u0_u0_U23  ( .A1(_AES_ENC_u0_u0_n576 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n840 ) );
NOR2_X2 _AES_ENC_u0_u0_U21  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n593 ), .ZN(_AES_ENC_u0_u0_n633 ) );
NOR2_X2 _AES_ENC_u0_u0_U20  ( .A1(_AES_ENC_u0_u0_n1009 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n960 ) );
NOR2_X2 _AES_ENC_u0_u0_U19  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n1045 ), .ZN(_AES_ENC_u0_u0_n812 ) );
NOR2_X2 _AES_ENC_u0_u0_U18  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n1080 ), .ZN(_AES_ENC_u0_u0_n1081 ) );
NOR2_X2 _AES_ENC_u0_u0_U17  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n601 ), .ZN(_AES_ENC_u0_u0_n982 ) );
NOR2_X2 _AES_ENC_u0_u0_U16  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n594 ), .ZN(_AES_ENC_u0_u0_n757 ) );
NOR2_X2 _AES_ENC_u0_u0_U15  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n590 ), .ZN(_AES_ENC_u0_u0_n698 ) );
NOR2_X2 _AES_ENC_u0_u0_U10  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n619 ), .ZN(_AES_ENC_u0_u0_n708 ) );
NOR2_X2 _AES_ENC_u0_u0_U9  ( .A1(_AES_ENC_u0_u0_n619 ), .A2(_AES_ENC_u0_u0_n604 ), .ZN(_AES_ENC_u0_u0_n803 ) );
NOR2_X2 _AES_ENC_u0_u0_U8  ( .A1(_AES_ENC_u0_u0_n615 ), .A2(_AES_ENC_u0_u0_n582 ), .ZN(_AES_ENC_u0_u0_n867 ) );
NOR2_X2 _AES_ENC_u0_u0_U7  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n599 ), .ZN(_AES_ENC_u0_u0_n804 ) );
NOR2_X2 _AES_ENC_u0_u0_U6  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n620 ), .ZN(_AES_ENC_u0_u0_n1046 ) );
OR2_X4 _AES_ENC_u0_u0_U5  ( .A1(_AES_ENC_u0_u0_n624 ), .A2(_AES_ENC_w3[17] ),.ZN(_AES_ENC_u0_u0_n570 ) );
OR2_X4 _AES_ENC_u0_u0_U4  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_w3[20] ),.ZN(_AES_ENC_u0_u0_n569 ) );
NAND2_X2 _AES_ENC_u0_u0_U514  ( .A1(_AES_ENC_u0_u0_n1121 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n1030 ) );
AND2_X2 _AES_ENC_u0_u0_U513  ( .A1(_AES_ENC_u0_u0_n597 ), .A2(_AES_ENC_u0_u0_n1030 ), .ZN(_AES_ENC_u0_u0_n1049 ) );
NAND2_X2 _AES_ENC_u0_u0_U511  ( .A1(_AES_ENC_u0_u0_n1049 ), .A2(_AES_ENC_u0_u0_n794 ), .ZN(_AES_ENC_u0_u0_n637 ) );
AND2_X2 _AES_ENC_u0_u0_U493  ( .A1(_AES_ENC_u0_u0_n779 ), .A2(_AES_ENC_u0_u0_n996 ), .ZN(_AES_ENC_u0_u0_n632 ) );
NAND4_X2 _AES_ENC_u0_u0_U485  ( .A1(_AES_ENC_u0_u0_n637 ), .A2(_AES_ENC_u0_u0_n636 ), .A3(_AES_ENC_u0_u0_n635 ), .A4(_AES_ENC_u0_u0_n634 ), .ZN(_AES_ENC_u0_u0_n638 ) );
NAND2_X2 _AES_ENC_u0_u0_U484  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n638 ), .ZN(_AES_ENC_u0_u0_n679 ) );
NAND2_X2 _AES_ENC_u0_u0_U481  ( .A1(_AES_ENC_u0_u0_n1094 ), .A2(_AES_ENC_u0_u0_n591 ), .ZN(_AES_ENC_u0_u0_n648 ) );
NAND2_X2 _AES_ENC_u0_u0_U476  ( .A1(_AES_ENC_u0_u0_n601 ), .A2(_AES_ENC_u0_u0_n590 ), .ZN(_AES_ENC_u0_u0_n762 ) );
NAND2_X2 _AES_ENC_u0_u0_U475  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n762 ), .ZN(_AES_ENC_u0_u0_n647 ) );
NAND4_X2 _AES_ENC_u0_u0_U457  ( .A1(_AES_ENC_u0_u0_n648 ), .A2(_AES_ENC_u0_u0_n647 ), .A3(_AES_ENC_u0_u0_n646 ), .A4(_AES_ENC_u0_u0_n645 ), .ZN(_AES_ENC_u0_u0_n649 ) );
NAND2_X2 _AES_ENC_u0_u0_U456  ( .A1(_AES_ENC_w3[16] ), .A2(_AES_ENC_u0_u0_n649 ), .ZN(_AES_ENC_u0_u0_n665 ) );
NAND2_X2 _AES_ENC_u0_u0_U454  ( .A1(_AES_ENC_u0_u0_n596 ), .A2(_AES_ENC_u0_u0_n623 ), .ZN(_AES_ENC_u0_u0_n855 ) );
NAND2_X2 _AES_ENC_u0_u0_U453  ( .A1(_AES_ENC_u0_u0_n587 ), .A2(_AES_ENC_u0_u0_n855 ), .ZN(_AES_ENC_u0_u0_n821 ) );
NAND2_X2 _AES_ENC_u0_u0_U452  ( .A1(_AES_ENC_u0_u0_n1093 ), .A2(_AES_ENC_u0_u0_n821 ), .ZN(_AES_ENC_u0_u0_n662 ) );
NAND2_X2 _AES_ENC_u0_u0_U451  ( .A1(_AES_ENC_u0_u0_n619 ), .A2(_AES_ENC_u0_u0_n589 ), .ZN(_AES_ENC_u0_u0_n650 ) );
NAND2_X2 _AES_ENC_u0_u0_U450  ( .A1(_AES_ENC_u0_u0_n956 ), .A2(_AES_ENC_u0_u0_n650 ), .ZN(_AES_ENC_u0_u0_n661 ) );
NAND2_X2 _AES_ENC_u0_u0_U449  ( .A1(_AES_ENC_u0_u0_n626 ), .A2(_AES_ENC_u0_u0_n627 ), .ZN(_AES_ENC_u0_u0_n839 ) );
OR2_X2 _AES_ENC_u0_u0_U446  ( .A1(_AES_ENC_u0_u0_n839 ), .A2(_AES_ENC_u0_u0_n932 ), .ZN(_AES_ENC_u0_u0_n656 ) );
NAND2_X2 _AES_ENC_u0_u0_U445  ( .A1(_AES_ENC_u0_u0_n621 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n1096 ) );
NAND2_X2 _AES_ENC_u0_u0_U444  ( .A1(_AES_ENC_u0_u0_n1030 ), .A2(_AES_ENC_u0_u0_n1096 ), .ZN(_AES_ENC_u0_u0_n651 ) );
NAND2_X2 _AES_ENC_u0_u0_U443  ( .A1(_AES_ENC_u0_u0_n1114 ), .A2(_AES_ENC_u0_u0_n651 ), .ZN(_AES_ENC_u0_u0_n655 ) );
OR3_X2 _AES_ENC_u0_u0_U440  ( .A1(_AES_ENC_u0_u0_n1079 ), .A2(_AES_ENC_w3[23] ), .A3(_AES_ENC_u0_u0_n626 ), .ZN(_AES_ENC_u0_u0_n654 ) );
NAND2_X2 _AES_ENC_u0_u0_U439  ( .A1(_AES_ENC_u0_u0_n593 ), .A2(_AES_ENC_u0_u0_n601 ), .ZN(_AES_ENC_u0_u0_n652 ) );
NAND4_X2 _AES_ENC_u0_u0_U437  ( .A1(_AES_ENC_u0_u0_n656 ), .A2(_AES_ENC_u0_u0_n655 ), .A3(_AES_ENC_u0_u0_n654 ), .A4(_AES_ENC_u0_u0_n653 ), .ZN(_AES_ENC_u0_u0_n657 ) );
NAND2_X2 _AES_ENC_u0_u0_U436  ( .A1(_AES_ENC_w3[18] ), .A2(_AES_ENC_u0_u0_n657 ), .ZN(_AES_ENC_u0_u0_n660 ) );
NAND4_X2 _AES_ENC_u0_u0_U432  ( .A1(_AES_ENC_u0_u0_n662 ), .A2(_AES_ENC_u0_u0_n661 ), .A3(_AES_ENC_u0_u0_n660 ), .A4(_AES_ENC_u0_u0_n659 ), .ZN(_AES_ENC_u0_u0_n663 ) );
NAND2_X2 _AES_ENC_u0_u0_U431  ( .A1(_AES_ENC_u0_u0_n663 ), .A2(_AES_ENC_u0_u0_n574 ), .ZN(_AES_ENC_u0_u0_n664 ) );
NAND2_X2 _AES_ENC_u0_u0_U430  ( .A1(_AES_ENC_u0_u0_n665 ), .A2(_AES_ENC_u0_u0_n664 ), .ZN(_AES_ENC_u0_u0_n666 ) );
NAND2_X2 _AES_ENC_u0_u0_U429  ( .A1(_AES_ENC_w3[22] ), .A2(_AES_ENC_u0_u0_n666 ), .ZN(_AES_ENC_u0_u0_n678 ) );
NAND2_X2 _AES_ENC_u0_u0_U426  ( .A1(_AES_ENC_u0_u0_n735 ), .A2(_AES_ENC_u0_u0_n1093 ), .ZN(_AES_ENC_u0_u0_n675 ) );
NAND2_X2 _AES_ENC_u0_u0_U425  ( .A1(_AES_ENC_u0_u0_n588 ), .A2(_AES_ENC_u0_u0_n597 ), .ZN(_AES_ENC_u0_u0_n1045 ) );
OR2_X2 _AES_ENC_u0_u0_U424  ( .A1(_AES_ENC_u0_u0_n1045 ), .A2(_AES_ENC_u0_u0_n605 ), .ZN(_AES_ENC_u0_u0_n674 ) );
NAND2_X2 _AES_ENC_u0_u0_U423  ( .A1(_AES_ENC_w3[17] ), .A2(_AES_ENC_u0_u0_n620 ), .ZN(_AES_ENC_u0_u0_n667 ) );
NAND2_X2 _AES_ENC_u0_u0_U422  ( .A1(_AES_ENC_u0_u0_n619 ), .A2(_AES_ENC_u0_u0_n667 ), .ZN(_AES_ENC_u0_u0_n1071 ) );
NAND4_X2 _AES_ENC_u0_u0_U412  ( .A1(_AES_ENC_u0_u0_n675 ), .A2(_AES_ENC_u0_u0_n674 ), .A3(_AES_ENC_u0_u0_n673 ), .A4(_AES_ENC_u0_u0_n672 ), .ZN(_AES_ENC_u0_u0_n676 ) );
NAND2_X2 _AES_ENC_u0_u0_U411  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n676 ), .ZN(_AES_ENC_u0_u0_n677 ) );
NAND2_X2 _AES_ENC_u0_u0_U408  ( .A1(_AES_ENC_u0_u0_n800 ), .A2(_AES_ENC_u0_u0_n1022 ), .ZN(_AES_ENC_u0_u0_n680 ) );
NAND2_X2 _AES_ENC_u0_u0_U407  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n680 ), .ZN(_AES_ENC_u0_u0_n681 ) );
AND2_X2 _AES_ENC_u0_u0_U402  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n684 ), .ZN(_AES_ENC_u0_u0_n682 ) );
NAND4_X2 _AES_ENC_u0_u0_U395  ( .A1(_AES_ENC_u0_u0_n691 ), .A2(_AES_ENC_u0_u0_n581 ), .A3(_AES_ENC_u0_u0_n690 ), .A4(_AES_ENC_u0_u0_n689 ), .ZN(_AES_ENC_u0_u0_n692 ) );
NAND2_X2 _AES_ENC_u0_u0_U394  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n692 ), .ZN(_AES_ENC_u0_u0_n733 ) );
NAND2_X2 _AES_ENC_u0_u0_U392  ( .A1(_AES_ENC_u0_u0_n977 ), .A2(_AES_ENC_u0_u0_n1050 ), .ZN(_AES_ENC_u0_u0_n702 ) );
NAND2_X2 _AES_ENC_u0_u0_U391  ( .A1(_AES_ENC_u0_u0_n1093 ), .A2(_AES_ENC_u0_u0_n1045 ), .ZN(_AES_ENC_u0_u0_n701 ) );
NAND4_X2 _AES_ENC_u0_u0_U381  ( .A1(_AES_ENC_u0_u0_n702 ), .A2(_AES_ENC_u0_u0_n701 ), .A3(_AES_ENC_u0_u0_n700 ), .A4(_AES_ENC_u0_u0_n699 ), .ZN(_AES_ENC_u0_u0_n703 ) );
NAND2_X2 _AES_ENC_u0_u0_U380  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n703 ), .ZN(_AES_ENC_u0_u0_n732 ) );
AND2_X2 _AES_ENC_u0_u0_U379  ( .A1(_AES_ENC_w3[16] ), .A2(_AES_ENC_w3[22] ),.ZN(_AES_ENC_u0_u0_n1113 ) );
NAND2_X2 _AES_ENC_u0_u0_U378  ( .A1(_AES_ENC_u0_u0_n601 ), .A2(_AES_ENC_u0_u0_n1030 ), .ZN(_AES_ENC_u0_u0_n881 ) );
NAND2_X2 _AES_ENC_u0_u0_U377  ( .A1(_AES_ENC_u0_u0_n1093 ), .A2(_AES_ENC_u0_u0_n881 ), .ZN(_AES_ENC_u0_u0_n715 ) );
NAND2_X2 _AES_ENC_u0_u0_U376  ( .A1(_AES_ENC_u0_u0_n1010 ), .A2(_AES_ENC_u0_u0_n600 ), .ZN(_AES_ENC_u0_u0_n714 ) );
NAND2_X2 _AES_ENC_u0_u0_U375  ( .A1(_AES_ENC_u0_u0_n855 ), .A2(_AES_ENC_u0_u0_n588 ), .ZN(_AES_ENC_u0_u0_n1117 ) );
XNOR2_X2 _AES_ENC_u0_u0_U371  ( .A(_AES_ENC_u0_u0_n611 ), .B(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n824 ) );
NAND4_X2 _AES_ENC_u0_u0_U362  ( .A1(_AES_ENC_u0_u0_n715 ), .A2(_AES_ENC_u0_u0_n714 ), .A3(_AES_ENC_u0_u0_n713 ), .A4(_AES_ENC_u0_u0_n712 ), .ZN(_AES_ENC_u0_u0_n716 ) );
NAND2_X2 _AES_ENC_u0_u0_U361  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n716 ), .ZN(_AES_ENC_u0_u0_n731 ) );
AND2_X2 _AES_ENC_u0_u0_U360  ( .A1(_AES_ENC_w3[22] ), .A2(_AES_ENC_u0_u0_n574 ), .ZN(_AES_ENC_u0_u0_n1131 ) );
NAND2_X2 _AES_ENC_u0_u0_U359  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n717 ) );
NAND2_X2 _AES_ENC_u0_u0_U358  ( .A1(_AES_ENC_u0_u0_n1029 ), .A2(_AES_ENC_u0_u0_n717 ), .ZN(_AES_ENC_u0_u0_n728 ) );
NAND2_X2 _AES_ENC_u0_u0_U357  ( .A1(_AES_ENC_w3[17] ), .A2(_AES_ENC_u0_u0_n624 ), .ZN(_AES_ENC_u0_u0_n1097 ) );
NAND2_X2 _AES_ENC_u0_u0_U356  ( .A1(_AES_ENC_u0_u0_n603 ), .A2(_AES_ENC_u0_u0_n1097 ), .ZN(_AES_ENC_u0_u0_n718 ) );
NAND2_X2 _AES_ENC_u0_u0_U355  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n718 ), .ZN(_AES_ENC_u0_u0_n727 ) );
NAND4_X2 _AES_ENC_u0_u0_U344  ( .A1(_AES_ENC_u0_u0_n728 ), .A2(_AES_ENC_u0_u0_n727 ), .A3(_AES_ENC_u0_u0_n726 ), .A4(_AES_ENC_u0_u0_n725 ), .ZN(_AES_ENC_u0_u0_n729 ) );
NAND2_X2 _AES_ENC_u0_u0_U343  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n729 ), .ZN(_AES_ENC_u0_u0_n730 ) );
NAND4_X2 _AES_ENC_u0_u0_U342  ( .A1(_AES_ENC_u0_u0_n733 ), .A2(_AES_ENC_u0_u0_n732 ), .A3(_AES_ENC_u0_u0_n731 ), .A4(_AES_ENC_u0_u0_n730 ), .ZN(_AES_ENC_u0_subword[25] ) );
NAND2_X2 _AES_ENC_u0_u0_U341  ( .A1(_AES_ENC_w3[23] ), .A2(_AES_ENC_u0_u0_n611 ), .ZN(_AES_ENC_u0_u0_n734 ) );
NAND2_X2 _AES_ENC_u0_u0_U340  ( .A1(_AES_ENC_u0_u0_n734 ), .A2(_AES_ENC_u0_u0_n607 ), .ZN(_AES_ENC_u0_u0_n738 ) );
OR4_X2 _AES_ENC_u0_u0_U339  ( .A1(_AES_ENC_u0_u0_n738 ), .A2(_AES_ENC_u0_u0_n626 ), .A3(_AES_ENC_u0_u0_n826 ), .A4(_AES_ENC_u0_u0_n1121 ), .ZN(_AES_ENC_u0_u0_n746 ) );
NAND2_X2 _AES_ENC_u0_u0_U337  ( .A1(_AES_ENC_u0_u0_n1100 ), .A2(_AES_ENC_u0_u0_n587 ), .ZN(_AES_ENC_u0_u0_n992 ) );
OR2_X2 _AES_ENC_u0_u0_U336  ( .A1(_AES_ENC_u0_u0_n610 ), .A2(_AES_ENC_u0_u0_n735 ), .ZN(_AES_ENC_u0_u0_n737 ) );
NAND2_X2 _AES_ENC_u0_u0_U334  ( .A1(_AES_ENC_u0_u0_n619 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n753 ) );
NAND2_X2 _AES_ENC_u0_u0_U333  ( .A1(_AES_ENC_u0_u0_n582 ), .A2(_AES_ENC_u0_u0_n753 ), .ZN(_AES_ENC_u0_u0_n1080 ) );
NAND2_X2 _AES_ENC_u0_u0_U332  ( .A1(_AES_ENC_u0_u0_n1048 ), .A2(_AES_ENC_u0_u0_n576 ), .ZN(_AES_ENC_u0_u0_n736 ) );
NAND2_X2 _AES_ENC_u0_u0_U331  ( .A1(_AES_ENC_u0_u0_n737 ), .A2(_AES_ENC_u0_u0_n736 ), .ZN(_AES_ENC_u0_u0_n739 ) );
NAND2_X2 _AES_ENC_u0_u0_U330  ( .A1(_AES_ENC_u0_u0_n739 ), .A2(_AES_ENC_u0_u0_n738 ), .ZN(_AES_ENC_u0_u0_n745 ) );
NAND2_X2 _AES_ENC_u0_u0_U326  ( .A1(_AES_ENC_u0_u0_n1096 ), .A2(_AES_ENC_u0_u0_n590 ), .ZN(_AES_ENC_u0_u0_n906 ) );
NAND4_X2 _AES_ENC_u0_u0_U323  ( .A1(_AES_ENC_u0_u0_n746 ), .A2(_AES_ENC_u0_u0_n992 ), .A3(_AES_ENC_u0_u0_n745 ), .A4(_AES_ENC_u0_u0_n744 ), .ZN(_AES_ENC_u0_u0_n747 ) );
NAND2_X2 _AES_ENC_u0_u0_U322  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n747 ), .ZN(_AES_ENC_u0_u0_n793 ) );
NAND2_X2 _AES_ENC_u0_u0_U321  ( .A1(_AES_ENC_u0_u0_n584 ), .A2(_AES_ENC_u0_u0_n855 ), .ZN(_AES_ENC_u0_u0_n748 ) );
NAND2_X2 _AES_ENC_u0_u0_U320  ( .A1(_AES_ENC_u0_u0_n956 ), .A2(_AES_ENC_u0_u0_n748 ), .ZN(_AES_ENC_u0_u0_n760 ) );
NAND2_X2 _AES_ENC_u0_u0_U313  ( .A1(_AES_ENC_u0_u0_n590 ), .A2(_AES_ENC_u0_u0_n753 ), .ZN(_AES_ENC_u0_u0_n1023 ) );
NAND4_X2 _AES_ENC_u0_u0_U308  ( .A1(_AES_ENC_u0_u0_n760 ), .A2(_AES_ENC_u0_u0_n992 ), .A3(_AES_ENC_u0_u0_n759 ), .A4(_AES_ENC_u0_u0_n758 ), .ZN(_AES_ENC_u0_u0_n761 ) );
NAND2_X2 _AES_ENC_u0_u0_U307  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n761 ), .ZN(_AES_ENC_u0_u0_n792 ) );
NAND2_X2 _AES_ENC_u0_u0_U306  ( .A1(_AES_ENC_u0_u0_n584 ), .A2(_AES_ENC_u0_u0_n603 ), .ZN(_AES_ENC_u0_u0_n989 ) );
NAND2_X2 _AES_ENC_u0_u0_U305  ( .A1(_AES_ENC_u0_u0_n1050 ), .A2(_AES_ENC_u0_u0_n989 ), .ZN(_AES_ENC_u0_u0_n777 ) );
NAND2_X2 _AES_ENC_u0_u0_U304  ( .A1(_AES_ENC_u0_u0_n1093 ), .A2(_AES_ENC_u0_u0_n762 ), .ZN(_AES_ENC_u0_u0_n776 ) );
XNOR2_X2 _AES_ENC_u0_u0_U301  ( .A(_AES_ENC_w3[23] ), .B(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n959 ) );
NAND4_X2 _AES_ENC_u0_u0_U289  ( .A1(_AES_ENC_u0_u0_n777 ), .A2(_AES_ENC_u0_u0_n776 ), .A3(_AES_ENC_u0_u0_n775 ), .A4(_AES_ENC_u0_u0_n774 ), .ZN(_AES_ENC_u0_u0_n778 ) );
NAND2_X2 _AES_ENC_u0_u0_U288  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n778 ), .ZN(_AES_ENC_u0_u0_n791 ) );
NAND2_X2 _AES_ENC_u0_u0_U287  ( .A1(_AES_ENC_u0_u0_n1056 ), .A2(_AES_ENC_u0_u0_n1050 ), .ZN(_AES_ENC_u0_u0_n788 ) );
NAND2_X2 _AES_ENC_u0_u0_U286  ( .A1(_AES_ENC_u0_u0_n1091 ), .A2(_AES_ENC_u0_u0_n779 ), .ZN(_AES_ENC_u0_u0_n787 ) );
NAND2_X2 _AES_ENC_u0_u0_U285  ( .A1(_AES_ENC_u0_u0_n956 ), .A2(_AES_ENC_w3[17] ), .ZN(_AES_ENC_u0_u0_n786 ) );
NAND4_X2 _AES_ENC_u0_u0_U278  ( .A1(_AES_ENC_u0_u0_n788 ), .A2(_AES_ENC_u0_u0_n787 ), .A3(_AES_ENC_u0_u0_n786 ), .A4(_AES_ENC_u0_u0_n785 ), .ZN(_AES_ENC_u0_u0_n789 ) );
NAND2_X2 _AES_ENC_u0_u0_U277  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n789 ), .ZN(_AES_ENC_u0_u0_n790 ) );
NAND4_X2 _AES_ENC_u0_u0_U276  ( .A1(_AES_ENC_u0_u0_n793 ), .A2(_AES_ENC_u0_u0_n792 ), .A3(_AES_ENC_u0_u0_n791 ), .A4(_AES_ENC_u0_u0_n790 ), .ZN(_AES_ENC_u0_subword[26] ) );
NAND2_X2 _AES_ENC_u0_u0_U275  ( .A1(_AES_ENC_u0_u0_n1059 ), .A2(_AES_ENC_u0_u0_n794 ), .ZN(_AES_ENC_u0_u0_n810 ) );
NAND2_X2 _AES_ENC_u0_u0_U274  ( .A1(_AES_ENC_u0_u0_n1049 ), .A2(_AES_ENC_u0_u0_n956 ), .ZN(_AES_ENC_u0_u0_n809 ) );
OR2_X2 _AES_ENC_u0_u0_U266  ( .A1(_AES_ENC_u0_u0_n1096 ), .A2(_AES_ENC_u0_u0_n606 ), .ZN(_AES_ENC_u0_u0_n802 ) );
NAND2_X2 _AES_ENC_u0_u0_U265  ( .A1(_AES_ENC_u0_u0_n1053 ), .A2(_AES_ENC_u0_u0_n800 ), .ZN(_AES_ENC_u0_u0_n801 ) );
NAND2_X2 _AES_ENC_u0_u0_U264  ( .A1(_AES_ENC_u0_u0_n802 ), .A2(_AES_ENC_u0_u0_n801 ), .ZN(_AES_ENC_u0_u0_n805 ) );
NAND4_X2 _AES_ENC_u0_u0_U261  ( .A1(_AES_ENC_u0_u0_n810 ), .A2(_AES_ENC_u0_u0_n809 ), .A3(_AES_ENC_u0_u0_n808 ), .A4(_AES_ENC_u0_u0_n807 ), .ZN(_AES_ENC_u0_u0_n811 ) );
NAND2_X2 _AES_ENC_u0_u0_U260  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n811 ), .ZN(_AES_ENC_u0_u0_n852 ) );
OR2_X2 _AES_ENC_u0_u0_U259  ( .A1(_AES_ENC_u0_u0_n1023 ), .A2(_AES_ENC_u0_u0_n617 ), .ZN(_AES_ENC_u0_u0_n819 ) );
OR2_X2 _AES_ENC_u0_u0_U257  ( .A1(_AES_ENC_u0_u0_n570 ), .A2(_AES_ENC_u0_u0_n930 ), .ZN(_AES_ENC_u0_u0_n818 ) );
NAND2_X2 _AES_ENC_u0_u0_U256  ( .A1(_AES_ENC_u0_u0_n1013 ), .A2(_AES_ENC_u0_u0_n1094 ), .ZN(_AES_ENC_u0_u0_n817 ) );
NAND4_X2 _AES_ENC_u0_u0_U249  ( .A1(_AES_ENC_u0_u0_n819 ), .A2(_AES_ENC_u0_u0_n818 ), .A3(_AES_ENC_u0_u0_n817 ), .A4(_AES_ENC_u0_u0_n816 ), .ZN(_AES_ENC_u0_u0_n820 ) );
NAND2_X2 _AES_ENC_u0_u0_U248  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n820 ), .ZN(_AES_ENC_u0_u0_n851 ) );
NAND2_X2 _AES_ENC_u0_u0_U247  ( .A1(_AES_ENC_u0_u0_n956 ), .A2(_AES_ENC_u0_u0_n1080 ), .ZN(_AES_ENC_u0_u0_n835 ) );
NAND2_X2 _AES_ENC_u0_u0_U246  ( .A1(_AES_ENC_u0_u0_n570 ), .A2(_AES_ENC_u0_u0_n1030 ), .ZN(_AES_ENC_u0_u0_n1047 ) );
OR2_X2 _AES_ENC_u0_u0_U245  ( .A1(_AES_ENC_u0_u0_n1047 ), .A2(_AES_ENC_u0_u0_n612 ), .ZN(_AES_ENC_u0_u0_n834 ) );
NAND2_X2 _AES_ENC_u0_u0_U244  ( .A1(_AES_ENC_u0_u0_n1072 ), .A2(_AES_ENC_u0_u0_n589 ), .ZN(_AES_ENC_u0_u0_n833 ) );
NAND4_X2 _AES_ENC_u0_u0_U233  ( .A1(_AES_ENC_u0_u0_n835 ), .A2(_AES_ENC_u0_u0_n834 ), .A3(_AES_ENC_u0_u0_n833 ), .A4(_AES_ENC_u0_u0_n832 ), .ZN(_AES_ENC_u0_u0_n836 ) );
NAND2_X2 _AES_ENC_u0_u0_U232  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n836 ), .ZN(_AES_ENC_u0_u0_n850 ) );
NAND2_X2 _AES_ENC_u0_u0_U231  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n623 ), .ZN(_AES_ENC_u0_u0_n847 ) );
NAND2_X2 _AES_ENC_u0_u0_U230  ( .A1(_AES_ENC_u0_u0_n1050 ), .A2(_AES_ENC_u0_u0_n1071 ), .ZN(_AES_ENC_u0_u0_n846 ) );
OR2_X2 _AES_ENC_u0_u0_U224  ( .A1(_AES_ENC_u0_u0_n1053 ), .A2(_AES_ENC_u0_u0_n911 ), .ZN(_AES_ENC_u0_u0_n1077 ) );
NAND4_X2 _AES_ENC_u0_u0_U220  ( .A1(_AES_ENC_u0_u0_n847 ), .A2(_AES_ENC_u0_u0_n846 ), .A3(_AES_ENC_u0_u0_n845 ), .A4(_AES_ENC_u0_u0_n844 ), .ZN(_AES_ENC_u0_u0_n848 ) );
NAND2_X2 _AES_ENC_u0_u0_U219  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n848 ), .ZN(_AES_ENC_u0_u0_n849 ) );
NAND4_X2 _AES_ENC_u0_u0_U218  ( .A1(_AES_ENC_u0_u0_n852 ), .A2(_AES_ENC_u0_u0_n851 ), .A3(_AES_ENC_u0_u0_n850 ), .A4(_AES_ENC_u0_u0_n849 ), .ZN(_AES_ENC_u0_subword[27] ) );
NAND2_X2 _AES_ENC_u0_u0_U216  ( .A1(_AES_ENC_u0_u0_n1009 ), .A2(_AES_ENC_u0_u0_n1072 ), .ZN(_AES_ENC_u0_u0_n862 ) );
NAND2_X2 _AES_ENC_u0_u0_U215  ( .A1(_AES_ENC_u0_u0_n603 ), .A2(_AES_ENC_u0_u0_n577 ), .ZN(_AES_ENC_u0_u0_n853 ) );
NAND2_X2 _AES_ENC_u0_u0_U214  ( .A1(_AES_ENC_u0_u0_n1050 ), .A2(_AES_ENC_u0_u0_n853 ), .ZN(_AES_ENC_u0_u0_n861 ) );
NAND4_X2 _AES_ENC_u0_u0_U206  ( .A1(_AES_ENC_u0_u0_n862 ), .A2(_AES_ENC_u0_u0_n861 ), .A3(_AES_ENC_u0_u0_n860 ), .A4(_AES_ENC_u0_u0_n859 ), .ZN(_AES_ENC_u0_u0_n863 ) );
NAND2_X2 _AES_ENC_u0_u0_U205  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n863 ), .ZN(_AES_ENC_u0_u0_n905 ) );
NAND2_X2 _AES_ENC_u0_u0_U204  ( .A1(_AES_ENC_u0_u0_n1010 ), .A2(_AES_ENC_u0_u0_n989 ), .ZN(_AES_ENC_u0_u0_n874 ) );
NAND2_X2 _AES_ENC_u0_u0_U203  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n610 ), .ZN(_AES_ENC_u0_u0_n864 ) );
NAND2_X2 _AES_ENC_u0_u0_U202  ( .A1(_AES_ENC_u0_u0_n929 ), .A2(_AES_ENC_u0_u0_n864 ), .ZN(_AES_ENC_u0_u0_n873 ) );
NAND4_X2 _AES_ENC_u0_u0_U193  ( .A1(_AES_ENC_u0_u0_n874 ), .A2(_AES_ENC_u0_u0_n873 ), .A3(_AES_ENC_u0_u0_n872 ), .A4(_AES_ENC_u0_u0_n871 ), .ZN(_AES_ENC_u0_u0_n875 ) );
NAND2_X2 _AES_ENC_u0_u0_U192  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n875 ), .ZN(_AES_ENC_u0_u0_n904 ) );
NAND2_X2 _AES_ENC_u0_u0_U191  ( .A1(_AES_ENC_u0_u0_n583 ), .A2(_AES_ENC_u0_u0_n1050 ), .ZN(_AES_ENC_u0_u0_n889 ) );
NAND2_X2 _AES_ENC_u0_u0_U190  ( .A1(_AES_ENC_u0_u0_n1093 ), .A2(_AES_ENC_u0_u0_n587 ), .ZN(_AES_ENC_u0_u0_n876 ) );
NAND2_X2 _AES_ENC_u0_u0_U189  ( .A1(_AES_ENC_u0_u0_n604 ), .A2(_AES_ENC_u0_u0_n876 ), .ZN(_AES_ENC_u0_u0_n877 ) );
NAND2_X2 _AES_ENC_u0_u0_U188  ( .A1(_AES_ENC_u0_u0_n877 ), .A2(_AES_ENC_u0_u0_n623 ), .ZN(_AES_ENC_u0_u0_n888 ) );
NAND4_X2 _AES_ENC_u0_u0_U179  ( .A1(_AES_ENC_u0_u0_n889 ), .A2(_AES_ENC_u0_u0_n888 ), .A3(_AES_ENC_u0_u0_n887 ), .A4(_AES_ENC_u0_u0_n886 ), .ZN(_AES_ENC_u0_u0_n890 ) );
NAND2_X2 _AES_ENC_u0_u0_U178  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n890 ), .ZN(_AES_ENC_u0_u0_n903 ) );
OR2_X2 _AES_ENC_u0_u0_U177  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n1059 ), .ZN(_AES_ENC_u0_u0_n900 ) );
NAND2_X2 _AES_ENC_u0_u0_U176  ( .A1(_AES_ENC_u0_u0_n1073 ), .A2(_AES_ENC_u0_u0_n1047 ), .ZN(_AES_ENC_u0_u0_n899 ) );
NAND2_X2 _AES_ENC_u0_u0_U175  ( .A1(_AES_ENC_u0_u0_n1094 ), .A2(_AES_ENC_u0_u0_n595 ), .ZN(_AES_ENC_u0_u0_n898 ) );
NAND4_X2 _AES_ENC_u0_u0_U167  ( .A1(_AES_ENC_u0_u0_n900 ), .A2(_AES_ENC_u0_u0_n899 ), .A3(_AES_ENC_u0_u0_n898 ), .A4(_AES_ENC_u0_u0_n897 ), .ZN(_AES_ENC_u0_u0_n901 ) );
NAND2_X2 _AES_ENC_u0_u0_U166  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n901 ), .ZN(_AES_ENC_u0_u0_n902 ) );
NAND4_X2 _AES_ENC_u0_u0_U165  ( .A1(_AES_ENC_u0_u0_n905 ), .A2(_AES_ENC_u0_u0_n904 ), .A3(_AES_ENC_u0_u0_n903 ), .A4(_AES_ENC_u0_u0_n902 ), .ZN(_AES_ENC_u0_subword[28] ) );
NAND2_X2 _AES_ENC_u0_u0_U164  ( .A1(_AES_ENC_u0_u0_n1094 ), .A2(_AES_ENC_u0_u0_n599 ), .ZN(_AES_ENC_u0_u0_n922 ) );
NAND2_X2 _AES_ENC_u0_u0_U163  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n989 ), .ZN(_AES_ENC_u0_u0_n921 ) );
NAND4_X2 _AES_ENC_u0_u0_U151  ( .A1(_AES_ENC_u0_u0_n922 ), .A2(_AES_ENC_u0_u0_n921 ), .A3(_AES_ENC_u0_u0_n920 ), .A4(_AES_ENC_u0_u0_n919 ), .ZN(_AES_ENC_u0_u0_n923 ) );
NAND2_X2 _AES_ENC_u0_u0_U150  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n923 ), .ZN(_AES_ENC_u0_u0_n972 ) );
NAND2_X2 _AES_ENC_u0_u0_U149  ( .A1(_AES_ENC_u0_u0_n582 ), .A2(_AES_ENC_u0_u0_n619 ), .ZN(_AES_ENC_u0_u0_n924 ) );
NAND2_X2 _AES_ENC_u0_u0_U148  ( .A1(_AES_ENC_u0_u0_n1073 ), .A2(_AES_ENC_u0_u0_n924 ), .ZN(_AES_ENC_u0_u0_n939 ) );
NAND2_X2 _AES_ENC_u0_u0_U147  ( .A1(_AES_ENC_u0_u0_n926 ), .A2(_AES_ENC_u0_u0_n925 ), .ZN(_AES_ENC_u0_u0_n927 ) );
NAND2_X2 _AES_ENC_u0_u0_U146  ( .A1(_AES_ENC_u0_u0_n606 ), .A2(_AES_ENC_u0_u0_n927 ), .ZN(_AES_ENC_u0_u0_n928 ) );
NAND2_X2 _AES_ENC_u0_u0_U145  ( .A1(_AES_ENC_u0_u0_n928 ), .A2(_AES_ENC_u0_u0_n1080 ), .ZN(_AES_ENC_u0_u0_n938 ) );
OR2_X2 _AES_ENC_u0_u0_U144  ( .A1(_AES_ENC_u0_u0_n1117 ), .A2(_AES_ENC_u0_u0_n615 ), .ZN(_AES_ENC_u0_u0_n937 ) );
NAND4_X2 _AES_ENC_u0_u0_U139  ( .A1(_AES_ENC_u0_u0_n939 ), .A2(_AES_ENC_u0_u0_n938 ), .A3(_AES_ENC_u0_u0_n937 ), .A4(_AES_ENC_u0_u0_n936 ), .ZN(_AES_ENC_u0_u0_n940 ) );
NAND2_X2 _AES_ENC_u0_u0_U138  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n940 ), .ZN(_AES_ENC_u0_u0_n971 ) );
OR2_X2 _AES_ENC_u0_u0_U137  ( .A1(_AES_ENC_u0_u0_n605 ), .A2(_AES_ENC_u0_u0_n941 ), .ZN(_AES_ENC_u0_u0_n954 ) );
NAND2_X2 _AES_ENC_u0_u0_U136  ( .A1(_AES_ENC_u0_u0_n1096 ), .A2(_AES_ENC_u0_u0_n577 ), .ZN(_AES_ENC_u0_u0_n942 ) );
NAND2_X2 _AES_ENC_u0_u0_U135  ( .A1(_AES_ENC_u0_u0_n1048 ), .A2(_AES_ENC_u0_u0_n942 ), .ZN(_AES_ENC_u0_u0_n943 ) );
NAND2_X2 _AES_ENC_u0_u0_U134  ( .A1(_AES_ENC_u0_u0_n612 ), .A2(_AES_ENC_u0_u0_n943 ), .ZN(_AES_ENC_u0_u0_n944 ) );
NAND2_X2 _AES_ENC_u0_u0_U133  ( .A1(_AES_ENC_u0_u0_n944 ), .A2(_AES_ENC_u0_u0_n580 ), .ZN(_AES_ENC_u0_u0_n953 ) );
NAND4_X2 _AES_ENC_u0_u0_U125  ( .A1(_AES_ENC_u0_u0_n954 ), .A2(_AES_ENC_u0_u0_n953 ), .A3(_AES_ENC_u0_u0_n952 ), .A4(_AES_ENC_u0_u0_n951 ), .ZN(_AES_ENC_u0_u0_n955 ) );
NAND2_X2 _AES_ENC_u0_u0_U124  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n955 ), .ZN(_AES_ENC_u0_u0_n970 ) );
NAND2_X2 _AES_ENC_u0_u0_U123  ( .A1(_AES_ENC_u0_u0_n1094 ), .A2(_AES_ENC_u0_u0_n1071 ), .ZN(_AES_ENC_u0_u0_n967 ) );
NAND2_X2 _AES_ENC_u0_u0_U122  ( .A1(_AES_ENC_u0_u0_n956 ), .A2(_AES_ENC_u0_u0_n1030 ), .ZN(_AES_ENC_u0_u0_n966 ) );
NAND4_X2 _AES_ENC_u0_u0_U114  ( .A1(_AES_ENC_u0_u0_n967 ), .A2(_AES_ENC_u0_u0_n966 ), .A3(_AES_ENC_u0_u0_n965 ), .A4(_AES_ENC_u0_u0_n964 ), .ZN(_AES_ENC_u0_u0_n968 ) );
NAND2_X2 _AES_ENC_u0_u0_U113  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n968 ), .ZN(_AES_ENC_u0_u0_n969 ) );
NAND4_X2 _AES_ENC_u0_u0_U112  ( .A1(_AES_ENC_u0_u0_n972 ), .A2(_AES_ENC_u0_u0_n971 ), .A3(_AES_ENC_u0_u0_n970 ), .A4(_AES_ENC_u0_u0_n969 ), .ZN(_AES_ENC_u0_subword[29] ) );
NAND2_X2 _AES_ENC_u0_u0_U111  ( .A1(_AES_ENC_u0_u0_n570 ), .A2(_AES_ENC_u0_u0_n1097 ), .ZN(_AES_ENC_u0_u0_n973 ) );
NAND2_X2 _AES_ENC_u0_u0_U110  ( .A1(_AES_ENC_u0_u0_n1073 ), .A2(_AES_ENC_u0_u0_n973 ), .ZN(_AES_ENC_u0_u0_n987 ) );
NAND2_X2 _AES_ENC_u0_u0_U109  ( .A1(_AES_ENC_u0_u0_n974 ), .A2(_AES_ENC_u0_u0_n1077 ), .ZN(_AES_ENC_u0_u0_n975 ) );
NAND2_X2 _AES_ENC_u0_u0_U108  ( .A1(_AES_ENC_u0_u0_n613 ), .A2(_AES_ENC_u0_u0_n975 ), .ZN(_AES_ENC_u0_u0_n976 ) );
NAND2_X2 _AES_ENC_u0_u0_U107  ( .A1(_AES_ENC_u0_u0_n977 ), .A2(_AES_ENC_u0_u0_n976 ), .ZN(_AES_ENC_u0_u0_n986 ) );
NAND4_X2 _AES_ENC_u0_u0_U99  ( .A1(_AES_ENC_u0_u0_n987 ), .A2(_AES_ENC_u0_u0_n986 ), .A3(_AES_ENC_u0_u0_n985 ), .A4(_AES_ENC_u0_u0_n984 ), .ZN(_AES_ENC_u0_u0_n988 ) );
NAND2_X2 _AES_ENC_u0_u0_U98  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n988 ), .ZN(_AES_ENC_u0_u0_n1044 ) );
NAND2_X2 _AES_ENC_u0_u0_U97  ( .A1(_AES_ENC_u0_u0_n1073 ), .A2(_AES_ENC_u0_u0_n989 ), .ZN(_AES_ENC_u0_u0_n1004 ) );
NAND2_X2 _AES_ENC_u0_u0_U96  ( .A1(_AES_ENC_u0_u0_n1092 ), .A2(_AES_ENC_u0_u0_n619 ), .ZN(_AES_ENC_u0_u0_n1003 ) );
NAND4_X2 _AES_ENC_u0_u0_U85  ( .A1(_AES_ENC_u0_u0_n1004 ), .A2(_AES_ENC_u0_u0_n1003 ), .A3(_AES_ENC_u0_u0_n1002 ), .A4(_AES_ENC_u0_u0_n1001 ), .ZN(_AES_ENC_u0_u0_n1005 ) );
NAND2_X2 _AES_ENC_u0_u0_U84  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n1005 ), .ZN(_AES_ENC_u0_u0_n1043 ) );
NAND2_X2 _AES_ENC_u0_u0_U83  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n596 ), .ZN(_AES_ENC_u0_u0_n1020 ) );
NAND2_X2 _AES_ENC_u0_u0_U82  ( .A1(_AES_ENC_u0_u0_n1050 ), .A2(_AES_ENC_u0_u0_n624 ), .ZN(_AES_ENC_u0_u0_n1019 ) );
NAND2_X2 _AES_ENC_u0_u0_U77  ( .A1(_AES_ENC_u0_u0_n1059 ), .A2(_AES_ENC_u0_u0_n1114 ), .ZN(_AES_ENC_u0_u0_n1012 ) );
NAND2_X2 _AES_ENC_u0_u0_U76  ( .A1(_AES_ENC_u0_u0_n1010 ), .A2(_AES_ENC_u0_u0_n592 ), .ZN(_AES_ENC_u0_u0_n1011 ) );
NAND2_X2 _AES_ENC_u0_u0_U75  ( .A1(_AES_ENC_u0_u0_n1012 ), .A2(_AES_ENC_u0_u0_n1011 ), .ZN(_AES_ENC_u0_u0_n1016 ) );
NAND4_X2 _AES_ENC_u0_u0_U70  ( .A1(_AES_ENC_u0_u0_n1020 ), .A2(_AES_ENC_u0_u0_n1019 ), .A3(_AES_ENC_u0_u0_n1018 ), .A4(_AES_ENC_u0_u0_n1017 ), .ZN(_AES_ENC_u0_u0_n1021 ) );
NAND2_X2 _AES_ENC_u0_u0_U69  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n1021 ), .ZN(_AES_ENC_u0_u0_n1042 ) );
NAND2_X2 _AES_ENC_u0_u0_U68  ( .A1(_AES_ENC_u0_u0_n1022 ), .A2(_AES_ENC_u0_u0_n1093 ), .ZN(_AES_ENC_u0_u0_n1039 ) );
NAND2_X2 _AES_ENC_u0_u0_U67  ( .A1(_AES_ENC_u0_u0_n1050 ), .A2(_AES_ENC_u0_u0_n1023 ), .ZN(_AES_ENC_u0_u0_n1038 ) );
NAND2_X2 _AES_ENC_u0_u0_U66  ( .A1(_AES_ENC_u0_u0_n1024 ), .A2(_AES_ENC_u0_u0_n1071 ), .ZN(_AES_ENC_u0_u0_n1037 ) );
AND2_X2 _AES_ENC_u0_u0_U60  ( .A1(_AES_ENC_u0_u0_n1030 ), .A2(_AES_ENC_u0_u0_n602 ), .ZN(_AES_ENC_u0_u0_n1078 ) );
NAND4_X2 _AES_ENC_u0_u0_U56  ( .A1(_AES_ENC_u0_u0_n1039 ), .A2(_AES_ENC_u0_u0_n1038 ), .A3(_AES_ENC_u0_u0_n1037 ), .A4(_AES_ENC_u0_u0_n1036 ), .ZN(_AES_ENC_u0_u0_n1040 ) );
NAND2_X2 _AES_ENC_u0_u0_U55  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n1040 ), .ZN(_AES_ENC_u0_u0_n1041 ) );
NAND4_X2 _AES_ENC_u0_u0_U54  ( .A1(_AES_ENC_u0_u0_n1044 ), .A2(_AES_ENC_u0_u0_n1043 ), .A3(_AES_ENC_u0_u0_n1042 ), .A4(_AES_ENC_u0_u0_n1041 ), .ZN(_AES_ENC_u0_subword[30] ) );
NAND2_X2 _AES_ENC_u0_u0_U53  ( .A1(_AES_ENC_u0_u0_n1072 ), .A2(_AES_ENC_u0_u0_n1045 ), .ZN(_AES_ENC_u0_u0_n1068 ) );
NAND2_X2 _AES_ENC_u0_u0_U52  ( .A1(_AES_ENC_u0_u0_n1046 ), .A2(_AES_ENC_u0_u0_n582 ), .ZN(_AES_ENC_u0_u0_n1067 ) );
NAND2_X2 _AES_ENC_u0_u0_U51  ( .A1(_AES_ENC_u0_u0_n1094 ), .A2(_AES_ENC_u0_u0_n1047 ), .ZN(_AES_ENC_u0_u0_n1066 ) );
NAND4_X2 _AES_ENC_u0_u0_U40  ( .A1(_AES_ENC_u0_u0_n1068 ), .A2(_AES_ENC_u0_u0_n1067 ), .A3(_AES_ENC_u0_u0_n1066 ), .A4(_AES_ENC_u0_u0_n1065 ), .ZN(_AES_ENC_u0_u0_n1069 ) );
NAND2_X2 _AES_ENC_u0_u0_U39  ( .A1(_AES_ENC_u0_u0_n1070 ), .A2(_AES_ENC_u0_u0_n1069 ), .ZN(_AES_ENC_u0_u0_n1135 ) );
NAND2_X2 _AES_ENC_u0_u0_U38  ( .A1(_AES_ENC_u0_u0_n1072 ), .A2(_AES_ENC_u0_u0_n1071 ), .ZN(_AES_ENC_u0_u0_n1088 ) );
NAND2_X2 _AES_ENC_u0_u0_U37  ( .A1(_AES_ENC_u0_u0_n1073 ), .A2(_AES_ENC_u0_u0_n595 ), .ZN(_AES_ENC_u0_u0_n1087 ) );
NAND4_X2 _AES_ENC_u0_u0_U28  ( .A1(_AES_ENC_u0_u0_n1088 ), .A2(_AES_ENC_u0_u0_n1087 ), .A3(_AES_ENC_u0_u0_n1086 ), .A4(_AES_ENC_u0_u0_n1085 ), .ZN(_AES_ENC_u0_u0_n1089 ) );
NAND2_X2 _AES_ENC_u0_u0_U27  ( .A1(_AES_ENC_u0_u0_n1090 ), .A2(_AES_ENC_u0_u0_n1089 ), .ZN(_AES_ENC_u0_u0_n1134 ) );
NAND2_X2 _AES_ENC_u0_u0_U26  ( .A1(_AES_ENC_u0_u0_n1091 ), .A2(_AES_ENC_u0_u0_n1093 ), .ZN(_AES_ENC_u0_u0_n1111 ) );
NAND2_X2 _AES_ENC_u0_u0_U25  ( .A1(_AES_ENC_u0_u0_n1092 ), .A2(_AES_ENC_u0_u0_n1120 ), .ZN(_AES_ENC_u0_u0_n1110 ) );
AND2_X2 _AES_ENC_u0_u0_U22  ( .A1(_AES_ENC_u0_u0_n1097 ), .A2(_AES_ENC_u0_u0_n1096 ), .ZN(_AES_ENC_u0_u0_n1098 ) );
NAND4_X2 _AES_ENC_u0_u0_U14  ( .A1(_AES_ENC_u0_u0_n1111 ), .A2(_AES_ENC_u0_u0_n1110 ), .A3(_AES_ENC_u0_u0_n1109 ), .A4(_AES_ENC_u0_u0_n1108 ), .ZN(_AES_ENC_u0_u0_n1112 ) );
NAND2_X2 _AES_ENC_u0_u0_U13  ( .A1(_AES_ENC_u0_u0_n1113 ), .A2(_AES_ENC_u0_u0_n1112 ), .ZN(_AES_ENC_u0_u0_n1133 ) );
NAND2_X2 _AES_ENC_u0_u0_U12  ( .A1(_AES_ENC_u0_u0_n1115 ), .A2(_AES_ENC_u0_u0_n1114 ), .ZN(_AES_ENC_u0_u0_n1129 ) );
OR2_X2 _AES_ENC_u0_u0_U11  ( .A1(_AES_ENC_u0_u0_n608 ), .A2(_AES_ENC_u0_u0_n1116 ), .ZN(_AES_ENC_u0_u0_n1128 ) );
NAND4_X2 _AES_ENC_u0_u0_U3  ( .A1(_AES_ENC_u0_u0_n1129 ), .A2(_AES_ENC_u0_u0_n1128 ), .A3(_AES_ENC_u0_u0_n1127 ), .A4(_AES_ENC_u0_u0_n1126 ), .ZN(_AES_ENC_u0_u0_n1130 ) );
NAND2_X2 _AES_ENC_u0_u0_U2  ( .A1(_AES_ENC_u0_u0_n1131 ), .A2(_AES_ENC_u0_u0_n1130 ), .ZN(_AES_ENC_u0_u0_n1132 ) );
NAND4_X2 _AES_ENC_u0_u0_U1  ( .A1(_AES_ENC_u0_u0_n1135 ), .A2(_AES_ENC_u0_u0_n1134 ), .A3(_AES_ENC_u0_u0_n1133 ), .A4(_AES_ENC_u0_u0_n1132 ), .ZN(_AES_ENC_u0_subword[31] ) );
INV_X4 _AES_ENC_u0_u1_U575  ( .A(_AES_ENC_w3[15] ), .ZN(_AES_ENC_u0_u1_n627 ) );
INV_X4 _AES_ENC_u0_u1_U574  ( .A(_AES_ENC_u0_u1_n1114 ), .ZN(_AES_ENC_u0_u1_n625 ) );
INV_X4 _AES_ENC_u0_u1_U573  ( .A(_AES_ENC_w3[12] ), .ZN(_AES_ENC_u0_u1_n624 ) );
INV_X4 _AES_ENC_u0_u1_U572  ( .A(_AES_ENC_u0_u1_n1025 ), .ZN(_AES_ENC_u0_u1_n622 ) );
INV_X4 _AES_ENC_u0_u1_U571  ( .A(_AES_ENC_u0_u1_n1120 ), .ZN(_AES_ENC_u0_u1_n620 ) );
INV_X4 _AES_ENC_u0_u1_U570  ( .A(_AES_ENC_u0_u1_n1121 ), .ZN(_AES_ENC_u0_u1_n619 ) );
INV_X4 _AES_ENC_u0_u1_U569  ( .A(_AES_ENC_u0_u1_n1048 ), .ZN(_AES_ENC_u0_u1_n618 ) );
INV_X4 _AES_ENC_u0_u1_U568  ( .A(_AES_ENC_u0_u1_n974 ), .ZN(_AES_ENC_u0_u1_n616 ) );
INV_X4 _AES_ENC_u0_u1_U567  ( .A(_AES_ENC_u0_u1_n794 ), .ZN(_AES_ENC_u0_u1_n614 ) );
INV_X4 _AES_ENC_u0_u1_U566  ( .A(_AES_ENC_w3[10] ), .ZN(_AES_ENC_u0_u1_n611 ) );
INV_X4 _AES_ENC_u0_u1_U565  ( .A(_AES_ENC_u0_u1_n800 ), .ZN(_AES_ENC_u0_u1_n610 ) );
INV_X4 _AES_ENC_u0_u1_U564  ( .A(_AES_ENC_u0_u1_n925 ), .ZN(_AES_ENC_u0_u1_n609 ) );
INV_X4 _AES_ENC_u0_u1_U563  ( .A(_AES_ENC_u0_u1_n779 ), .ZN(_AES_ENC_u0_u1_n607 ) );
INV_X4 _AES_ENC_u0_u1_U562  ( .A(_AES_ENC_u0_u1_n1022 ), .ZN(_AES_ENC_u0_u1_n603 ) );
INV_X4 _AES_ENC_u0_u1_U561  ( .A(_AES_ENC_u0_u1_n1102 ), .ZN(_AES_ENC_u0_u1_n602 ) );
INV_X4 _AES_ENC_u0_u1_U560  ( .A(_AES_ENC_u0_u1_n929 ), .ZN(_AES_ENC_u0_u1_n601 ) );
INV_X4 _AES_ENC_u0_u1_U559  ( .A(_AES_ENC_u0_u1_n1056 ), .ZN(_AES_ENC_u0_u1_n600 ) );
INV_X4 _AES_ENC_u0_u1_U558  ( .A(_AES_ENC_u0_u1_n1054 ), .ZN(_AES_ENC_u0_u1_n599 ) );
INV_X4 _AES_ENC_u0_u1_U557  ( .A(_AES_ENC_u0_u1_n881 ), .ZN(_AES_ENC_u0_u1_n598 ) );
INV_X4 _AES_ENC_u0_u1_U556  ( .A(_AES_ENC_u0_u1_n926 ), .ZN(_AES_ENC_u0_u1_n597 ) );
INV_X4 _AES_ENC_u0_u1_U555  ( .A(_AES_ENC_u0_u1_n977 ), .ZN(_AES_ENC_u0_u1_n595 ) );
INV_X4 _AES_ENC_u0_u1_U554  ( .A(_AES_ENC_u0_u1_n1031 ), .ZN(_AES_ENC_u0_u1_n594 ) );
INV_X4 _AES_ENC_u0_u1_U553  ( .A(_AES_ENC_u0_u1_n1103 ), .ZN(_AES_ENC_u0_u1_n593 ) );
INV_X4 _AES_ENC_u0_u1_U552  ( .A(_AES_ENC_u0_u1_n1009 ), .ZN(_AES_ENC_u0_u1_n592 ) );
INV_X4 _AES_ENC_u0_u1_U551  ( .A(_AES_ENC_u0_u1_n990 ), .ZN(_AES_ENC_u0_u1_n591 ) );
INV_X4 _AES_ENC_u0_u1_U550  ( .A(_AES_ENC_u0_u1_n1058 ), .ZN(_AES_ENC_u0_u1_n590 ) );
INV_X4 _AES_ENC_u0_u1_U549  ( .A(_AES_ENC_u0_u1_n1074 ), .ZN(_AES_ENC_u0_u1_n589 ) );
INV_X4 _AES_ENC_u0_u1_U548  ( .A(_AES_ENC_u0_u1_n1053 ), .ZN(_AES_ENC_u0_u1_n588 ) );
INV_X4 _AES_ENC_u0_u1_U547  ( .A(_AES_ENC_u0_u1_n826 ), .ZN(_AES_ENC_u0_u1_n587 ) );
INV_X4 _AES_ENC_u0_u1_U546  ( .A(_AES_ENC_u0_u1_n992 ), .ZN(_AES_ENC_u0_u1_n586 ) );
INV_X4 _AES_ENC_u0_u1_U545  ( .A(_AES_ENC_u0_u1_n821 ), .ZN(_AES_ENC_u0_u1_n585 ) );
INV_X4 _AES_ENC_u0_u1_U544  ( .A(_AES_ENC_u0_u1_n910 ), .ZN(_AES_ENC_u0_u1_n584 ) );
INV_X4 _AES_ENC_u0_u1_U543  ( .A(_AES_ENC_u0_u1_n906 ), .ZN(_AES_ENC_u0_u1_n583 ) );
INV_X4 _AES_ENC_u0_u1_U542  ( .A(_AES_ENC_u0_u1_n880 ), .ZN(_AES_ENC_u0_u1_n581 ) );
INV_X4 _AES_ENC_u0_u1_U541  ( .A(_AES_ENC_u0_u1_n1013 ), .ZN(_AES_ENC_u0_u1_n580 ) );
INV_X4 _AES_ENC_u0_u1_U540  ( .A(_AES_ENC_u0_u1_n1092 ), .ZN(_AES_ENC_u0_u1_n579 ) );
INV_X4 _AES_ENC_u0_u1_U539  ( .A(_AES_ENC_u0_u1_n824 ), .ZN(_AES_ENC_u0_u1_n578 ) );
INV_X4 _AES_ENC_u0_u1_U538  ( .A(_AES_ENC_u0_u1_n1091 ), .ZN(_AES_ENC_u0_u1_n577 ) );
INV_X4 _AES_ENC_u0_u1_U537  ( .A(_AES_ENC_u0_u1_n1080 ), .ZN(_AES_ENC_u0_u1_n576 ) );
INV_X4 _AES_ENC_u0_u1_U536  ( .A(_AES_ENC_u0_u1_n959 ), .ZN(_AES_ENC_u0_u1_n575 ) );
INV_X4 _AES_ENC_u0_u1_U535  ( .A(_AES_ENC_w3[8] ), .ZN(_AES_ENC_u0_u1_n574 ));
NOR2_X2 _AES_ENC_u0_u1_U534  ( .A1(_AES_ENC_u0_u1_n574 ), .A2(_AES_ENC_w3[14] ), .ZN(_AES_ENC_u0_u1_n1070 ) );
NOR2_X2 _AES_ENC_u0_u1_U533  ( .A1(_AES_ENC_w3[8] ), .A2(_AES_ENC_w3[14] ),.ZN(_AES_ENC_u0_u1_n1090 ) );
NOR2_X2 _AES_ENC_u0_u1_U532  ( .A1(_AES_ENC_w3[12] ), .A2(_AES_ENC_w3[11] ),.ZN(_AES_ENC_u0_u1_n1025 ) );
NAND3_X2 _AES_ENC_u0_u1_U531  ( .A1(_AES_ENC_u0_u1_n679 ), .A2(_AES_ENC_u0_u1_n678 ), .A3(_AES_ENC_u0_u1_n677 ), .ZN(_AES_ENC_u0_subword[16] ) );
NOR2_X2 _AES_ENC_u0_u1_U530  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n765 ) );
NOR2_X2 _AES_ENC_u0_u1_U529  ( .A1(_AES_ENC_w3[12] ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n764 ) );
NOR2_X2 _AES_ENC_u0_u1_U528  ( .A1(_AES_ENC_u0_u1_n765 ), .A2(_AES_ENC_u0_u1_n764 ), .ZN(_AES_ENC_u0_u1_n766 ) );
NOR2_X2 _AES_ENC_u0_u1_U527  ( .A1(_AES_ENC_u0_u1_n766 ), .A2(_AES_ENC_u0_u1_n575 ), .ZN(_AES_ENC_u0_u1_n767 ) );
NOR2_X2 _AES_ENC_u0_u1_U526  ( .A1(_AES_ENC_u0_u1_n1117 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n707 ) );
NOR3_X2 _AES_ENC_u0_u1_U525  ( .A1(_AES_ENC_u0_u1_n627 ), .A2(_AES_ENC_w3[13] ), .A3(_AES_ENC_u0_u1_n704 ), .ZN(_AES_ENC_u0_u1_n706 ) );
NOR2_X2 _AES_ENC_u0_u1_U524  ( .A1(_AES_ENC_w3[12] ), .A2(_AES_ENC_u0_u1_n579 ), .ZN(_AES_ENC_u0_u1_n705 ) );
NOR3_X2 _AES_ENC_u0_u1_U523  ( .A1(_AES_ENC_u0_u1_n707 ), .A2(_AES_ENC_u0_u1_n706 ), .A3(_AES_ENC_u0_u1_n705 ), .ZN(_AES_ENC_u0_u1_n713 ) );
NOR4_X2 _AES_ENC_u0_u1_U522  ( .A1(_AES_ENC_u0_u1_n633 ), .A2(_AES_ENC_u0_u1_n632 ), .A3(_AES_ENC_u0_u1_n631 ), .A4(_AES_ENC_u0_u1_n630 ), .ZN(_AES_ENC_u0_u1_n634 ) );
NOR2_X2 _AES_ENC_u0_u1_U521  ( .A1(_AES_ENC_u0_u1_n629 ), .A2(_AES_ENC_u0_u1_n628 ), .ZN(_AES_ENC_u0_u1_n635 ) );
NAND3_X2 _AES_ENC_u0_u1_U520  ( .A1(_AES_ENC_w3[10] ), .A2(_AES_ENC_w3[15] ),.A3(_AES_ENC_u0_u1_n1059 ), .ZN(_AES_ENC_u0_u1_n636 ) );
INV_X4 _AES_ENC_u0_u1_U519  ( .A(_AES_ENC_w3[11] ), .ZN(_AES_ENC_u0_u1_n621 ) );
NOR2_X2 _AES_ENC_u0_u1_U518  ( .A1(_AES_ENC_w3[13] ), .A2(_AES_ENC_w3[10] ),.ZN(_AES_ENC_u0_u1_n974 ) );
NAND3_X2 _AES_ENC_u0_u1_U517  ( .A1(_AES_ENC_u0_u1_n652 ), .A2(_AES_ENC_u0_u1_n626 ), .A3(_AES_ENC_w3[15] ), .ZN(_AES_ENC_u0_u1_n653 ) );
NOR2_X2 _AES_ENC_u0_u1_U516  ( .A1(_AES_ENC_u0_u1_n611 ), .A2(_AES_ENC_w3[13] ), .ZN(_AES_ENC_u0_u1_n925 ) );
NOR2_X2 _AES_ENC_u0_u1_U515  ( .A1(_AES_ENC_u0_u1_n626 ), .A2(_AES_ENC_w3[10] ), .ZN(_AES_ENC_u0_u1_n1048 ) );
INV_X4 _AES_ENC_u0_u1_U512  ( .A(_AES_ENC_w3[13] ), .ZN(_AES_ENC_u0_u1_n626 ) );
NOR2_X2 _AES_ENC_u0_u1_U510  ( .A1(_AES_ENC_u0_u1_n611 ), .A2(_AES_ENC_w3[15] ), .ZN(_AES_ENC_u0_u1_n779 ) );
NOR2_X2 _AES_ENC_u0_u1_U509  ( .A1(_AES_ENC_w3[15] ), .A2(_AES_ENC_w3[10] ),.ZN(_AES_ENC_u0_u1_n794 ) );
NOR2_X2 _AES_ENC_u0_u1_U508  ( .A1(_AES_ENC_w3[12] ), .A2(_AES_ENC_w3[9] ),.ZN(_AES_ENC_u0_u1_n1102 ) );
INV_X4 _AES_ENC_u0_u1_U507  ( .A(_AES_ENC_u0_u1_n569 ), .ZN(_AES_ENC_u0_u1_n572 ) );
NOR2_X2 _AES_ENC_u0_u1_U506  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_w3[11] ), .ZN(_AES_ENC_u0_u1_n1053 ) );
NOR2_X2 _AES_ENC_u0_u1_U505  ( .A1(_AES_ENC_u0_u1_n607 ), .A2(_AES_ENC_w3[13] ), .ZN(_AES_ENC_u0_u1_n1024 ) );
NOR2_X2 _AES_ENC_u0_u1_U504  ( .A1(_AES_ENC_u0_u1_n625 ), .A2(_AES_ENC_w3[10] ), .ZN(_AES_ENC_u0_u1_n1093 ) );
NOR2_X2 _AES_ENC_u0_u1_U503  ( .A1(_AES_ENC_u0_u1_n614 ), .A2(_AES_ENC_w3[13] ), .ZN(_AES_ENC_u0_u1_n1094 ) );
NOR2_X2 _AES_ENC_u0_u1_U502  ( .A1(_AES_ENC_u0_u1_n624 ), .A2(_AES_ENC_w3[11] ), .ZN(_AES_ENC_u0_u1_n931 ) );
INV_X4 _AES_ENC_u0_u1_U501  ( .A(_AES_ENC_u0_u1_n570 ), .ZN(_AES_ENC_u0_u1_n573 ) );
NOR2_X2 _AES_ENC_u0_u1_U500  ( .A1(_AES_ENC_u0_u1_n622 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n1059 ) );
NOR2_X2 _AES_ENC_u0_u1_U499  ( .A1(_AES_ENC_u0_u1_n1053 ), .A2(_AES_ENC_u0_u1_n1095 ), .ZN(_AES_ENC_u0_u1_n639 ) );
NOR3_X2 _AES_ENC_u0_u1_U498  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n573 ), .A3(_AES_ENC_u0_u1_n1074 ), .ZN(_AES_ENC_u0_u1_n641 ) );
NOR2_X2 _AES_ENC_u0_u1_U497  ( .A1(_AES_ENC_u0_u1_n639 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n640 ) );
NOR2_X2 _AES_ENC_u0_u1_U496  ( .A1(_AES_ENC_u0_u1_n641 ), .A2(_AES_ENC_u0_u1_n640 ), .ZN(_AES_ENC_u0_u1_n646 ) );
NOR2_X2 _AES_ENC_u0_u1_U495  ( .A1(_AES_ENC_u0_u1_n826 ), .A2(_AES_ENC_u0_u1_n572 ), .ZN(_AES_ENC_u0_u1_n827 ) );
NOR3_X2 _AES_ENC_u0_u1_U494  ( .A1(_AES_ENC_u0_u1_n769 ), .A2(_AES_ENC_u0_u1_n768 ), .A3(_AES_ENC_u0_u1_n767 ), .ZN(_AES_ENC_u0_u1_n775 ) );
NOR2_X2 _AES_ENC_u0_u1_U492  ( .A1(_AES_ENC_w3[9] ), .A2(_AES_ENC_u0_u1_n623 ), .ZN(_AES_ENC_u0_u1_n913 ) );
NOR2_X2 _AES_ENC_u0_u1_U491  ( .A1(_AES_ENC_u0_u1_n913 ), .A2(_AES_ENC_u0_u1_n1091 ), .ZN(_AES_ENC_u0_u1_n914 ) );
NOR2_X2 _AES_ENC_u0_u1_U490  ( .A1(_AES_ENC_u0_u1_n1056 ), .A2(_AES_ENC_u0_u1_n1053 ), .ZN(_AES_ENC_u0_u1_n749 ) );
NOR2_X2 _AES_ENC_u0_u1_U489  ( .A1(_AES_ENC_u0_u1_n749 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n752 ) );
NOR3_X2 _AES_ENC_u0_u1_U488  ( .A1(_AES_ENC_u0_u1_n995 ), .A2(_AES_ENC_u0_u1_n586 ), .A3(_AES_ENC_u0_u1_n994 ), .ZN(_AES_ENC_u0_u1_n1002 ) );
NOR2_X2 _AES_ENC_u0_u1_U487  ( .A1(_AES_ENC_u0_u1_n909 ), .A2(_AES_ENC_u0_u1_n908 ), .ZN(_AES_ENC_u0_u1_n920 ) );
INV_X4 _AES_ENC_u0_u1_U486  ( .A(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n596 ));
NOR2_X2 _AES_ENC_u0_u1_U483  ( .A1(_AES_ENC_u0_u1_n932 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n933 ) );
NOR2_X2 _AES_ENC_u0_u1_U482  ( .A1(_AES_ENC_u0_u1_n929 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n935 ) );
NOR2_X2 _AES_ENC_u0_u1_U480  ( .A1(_AES_ENC_u0_u1_n931 ), .A2(_AES_ENC_u0_u1_n930 ), .ZN(_AES_ENC_u0_u1_n934 ) );
NOR3_X2 _AES_ENC_u0_u1_U479  ( .A1(_AES_ENC_u0_u1_n935 ), .A2(_AES_ENC_u0_u1_n934 ), .A3(_AES_ENC_u0_u1_n933 ), .ZN(_AES_ENC_u0_u1_n936 ) );
OR2_X4 _AES_ENC_u0_u1_U478  ( .A1(_AES_ENC_u0_u1_n1094 ), .A2(_AES_ENC_u0_u1_n1093 ), .ZN(_AES_ENC_u0_u1_n571 ) );
AND2_X2 _AES_ENC_u0_u1_U477  ( .A1(_AES_ENC_u0_u1_n571 ), .A2(_AES_ENC_u0_u1_n1095 ), .ZN(_AES_ENC_u0_u1_n1101 ) );
NOR2_X2 _AES_ENC_u0_u1_U474  ( .A1(_AES_ENC_u0_u1_n1074 ), .A2(_AES_ENC_u0_u1_n931 ), .ZN(_AES_ENC_u0_u1_n796 ) );
NOR2_X2 _AES_ENC_u0_u1_U473  ( .A1(_AES_ENC_u0_u1_n796 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n797 ) );
NOR2_X2 _AES_ENC_u0_u1_U472  ( .A1(_AES_ENC_u0_u1_n1054 ), .A2(_AES_ENC_u0_u1_n1053 ), .ZN(_AES_ENC_u0_u1_n1055 ) );
NOR2_X2 _AES_ENC_u0_u1_U471  ( .A1(_AES_ENC_u0_u1_n572 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n949 ) );
NOR2_X2 _AES_ENC_u0_u1_U470  ( .A1(_AES_ENC_u0_u1_n1049 ), .A2(_AES_ENC_u0_u1_n618 ), .ZN(_AES_ENC_u0_u1_n1051 ) );
NOR2_X2 _AES_ENC_u0_u1_U469  ( .A1(_AES_ENC_u0_u1_n1051 ), .A2(_AES_ENC_u0_u1_n1050 ), .ZN(_AES_ENC_u0_u1_n1052 ) );
NOR2_X2 _AES_ENC_u0_u1_U468  ( .A1(_AES_ENC_u0_u1_n1052 ), .A2(_AES_ENC_u0_u1_n592 ), .ZN(_AES_ENC_u0_u1_n1064 ) );
NOR2_X2 _AES_ENC_u0_u1_U467  ( .A1(_AES_ENC_w3[9] ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n631 ) );
NOR2_X2 _AES_ENC_u0_u1_U466  ( .A1(_AES_ENC_u0_u1_n1025 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n980 ) );
NOR2_X2 _AES_ENC_u0_u1_U465  ( .A1(_AES_ENC_u0_u1_n1074 ), .A2(_AES_ENC_u0_u1_n1025 ), .ZN(_AES_ENC_u0_u1_n891 ) );
NOR2_X2 _AES_ENC_u0_u1_U464  ( .A1(_AES_ENC_u0_u1_n891 ), .A2(_AES_ENC_u0_u1_n609 ), .ZN(_AES_ENC_u0_u1_n894 ) );
NOR2_X2 _AES_ENC_u0_u1_U463  ( .A1(_AES_ENC_u0_u1_n1073 ), .A2(_AES_ENC_u0_u1_n1094 ), .ZN(_AES_ENC_u0_u1_n795 ) );
NOR2_X2 _AES_ENC_u0_u1_U462  ( .A1(_AES_ENC_u0_u1_n795 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n799 ) );
NOR2_X2 _AES_ENC_u0_u1_U461  ( .A1(_AES_ENC_u0_u1_n624 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n1075 ) );
NOR2_X2 _AES_ENC_u0_u1_U460  ( .A1(_AES_ENC_u0_u1_n624 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n822 ) );
NOR2_X2 _AES_ENC_u0_u1_U459  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n823 ) );
NOR2_X2 _AES_ENC_u0_u1_U458  ( .A1(_AES_ENC_u0_u1_n823 ), .A2(_AES_ENC_u0_u1_n822 ), .ZN(_AES_ENC_u0_u1_n825 ) );
NOR2_X2 _AES_ENC_u0_u1_U455  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n981 ) );
NOR2_X2 _AES_ENC_u0_u1_U448  ( .A1(_AES_ENC_u0_u1_n1102 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n643 ) );
NOR2_X2 _AES_ENC_u0_u1_U447  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n621 ), .ZN(_AES_ENC_u0_u1_n642 ) );
NOR2_X2 _AES_ENC_u0_u1_U442  ( .A1(_AES_ENC_u0_u1_n911 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n644 ) );
NOR4_X2 _AES_ENC_u0_u1_U441  ( .A1(_AES_ENC_u0_u1_n644 ), .A2(_AES_ENC_u0_u1_n643 ), .A3(_AES_ENC_u0_u1_n804 ), .A4(_AES_ENC_u0_u1_n642 ), .ZN(_AES_ENC_u0_u1_n645 ) );
NOR2_X2 _AES_ENC_u0_u1_U438  ( .A1(_AES_ENC_u0_u1_n1102 ), .A2(_AES_ENC_u0_u1_n910 ), .ZN(_AES_ENC_u0_u1_n932 ) );
NOR3_X2 _AES_ENC_u0_u1_U435  ( .A1(_AES_ENC_u0_u1_n623 ), .A2(_AES_ENC_w3[9] ), .A3(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n683 ));
NOR2_X2 _AES_ENC_u0_u1_U434  ( .A1(_AES_ENC_u0_u1_n1102 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n755 ) );
INV_X4 _AES_ENC_u0_u1_U433  ( .A(_AES_ENC_u0_u1_n931 ), .ZN(_AES_ENC_u0_u1_n623 ) );
NOR2_X2 _AES_ENC_u0_u1_U428  ( .A1(_AES_ENC_u0_u1_n996 ), .A2(_AES_ENC_u0_u1_n931 ), .ZN(_AES_ENC_u0_u1_n704 ) );
NOR2_X2 _AES_ENC_u0_u1_U427  ( .A1(_AES_ENC_u0_u1_n1029 ), .A2(_AES_ENC_u0_u1_n1025 ), .ZN(_AES_ENC_u0_u1_n1079 ) );
NOR3_X2 _AES_ENC_u0_u1_U421  ( .A1(_AES_ENC_u0_u1_n589 ), .A2(_AES_ENC_u0_u1_n1025 ), .A3(_AES_ENC_u0_u1_n616 ), .ZN(_AES_ENC_u0_u1_n945 ) );
NOR2_X2 _AES_ENC_u0_u1_U420  ( .A1(_AES_ENC_u0_u1_n1072 ), .A2(_AES_ENC_u0_u1_n1094 ), .ZN(_AES_ENC_u0_u1_n930 ) );
NOR2_X2 _AES_ENC_u0_u1_U419  ( .A1(_AES_ENC_u0_u1_n931 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n743 ) );
NOR2_X2 _AES_ENC_u0_u1_U418  ( .A1(_AES_ENC_u0_u1_n931 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n685 ) );
NOR3_X2 _AES_ENC_u0_u1_U417  ( .A1(_AES_ENC_u0_u1_n610 ), .A2(_AES_ENC_u0_u1_n572 ), .A3(_AES_ENC_u0_u1_n575 ), .ZN(_AES_ENC_u0_u1_n962 ) );
NOR2_X2 _AES_ENC_u0_u1_U416  ( .A1(_AES_ENC_u0_u1_n626 ), .A2(_AES_ENC_u0_u1_n611 ), .ZN(_AES_ENC_u0_u1_n800 ) );
NOR3_X2 _AES_ENC_u0_u1_U415  ( .A1(_AES_ENC_u0_u1_n590 ), .A2(_AES_ENC_u0_u1_n627 ), .A3(_AES_ENC_u0_u1_n611 ), .ZN(_AES_ENC_u0_u1_n798 ) );
NOR3_X2 _AES_ENC_u0_u1_U414  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n572 ), .A3(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n694 ) );
NOR3_X2 _AES_ENC_u0_u1_U413  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n572 ), .A3(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n895 ) );
NOR3_X2 _AES_ENC_u0_u1_U410  ( .A1(_AES_ENC_u0_u1_n1008 ), .A2(_AES_ENC_u0_u1_n1007 ), .A3(_AES_ENC_u0_u1_n1006 ), .ZN(_AES_ENC_u0_u1_n1018 ) );
NOR2_X2 _AES_ENC_u0_u1_U409  ( .A1(_AES_ENC_u0_u1_n669 ), .A2(_AES_ENC_u0_u1_n668 ), .ZN(_AES_ENC_u0_u1_n673 ) );
NOR4_X2 _AES_ENC_u0_u1_U406  ( .A1(_AES_ENC_u0_u1_n946 ), .A2(_AES_ENC_u0_u1_n1046 ), .A3(_AES_ENC_u0_u1_n671 ), .A4(_AES_ENC_u0_u1_n670 ), .ZN(_AES_ENC_u0_u1_n672 ) );
NOR4_X2 _AES_ENC_u0_u1_U405  ( .A1(_AES_ENC_u0_u1_n711 ), .A2(_AES_ENC_u0_u1_n710 ), .A3(_AES_ENC_u0_u1_n709 ), .A4(_AES_ENC_u0_u1_n708 ), .ZN(_AES_ENC_u0_u1_n712 ) );
NOR4_X2 _AES_ENC_u0_u1_U404  ( .A1(_AES_ENC_u0_u1_n806 ), .A2(_AES_ENC_u0_u1_n805 ), .A3(_AES_ENC_u0_u1_n804 ), .A4(_AES_ENC_u0_u1_n803 ), .ZN(_AES_ENC_u0_u1_n807 ) );
NOR3_X2 _AES_ENC_u0_u1_U403  ( .A1(_AES_ENC_u0_u1_n799 ), .A2(_AES_ENC_u0_u1_n798 ), .A3(_AES_ENC_u0_u1_n797 ), .ZN(_AES_ENC_u0_u1_n808 ) );
NOR4_X2 _AES_ENC_u0_u1_U401  ( .A1(_AES_ENC_u0_u1_n843 ), .A2(_AES_ENC_u0_u1_n842 ), .A3(_AES_ENC_u0_u1_n841 ), .A4(_AES_ENC_u0_u1_n840 ), .ZN(_AES_ENC_u0_u1_n844 ) );
NOR3_X2 _AES_ENC_u0_u1_U400  ( .A1(_AES_ENC_u0_u1_n1101 ), .A2(_AES_ENC_u0_u1_n1100 ), .A3(_AES_ENC_u0_u1_n1099 ), .ZN(_AES_ENC_u0_u1_n1109 ) );
NOR3_X2 _AES_ENC_u0_u1_U399  ( .A1(_AES_ENC_u0_u1_n743 ), .A2(_AES_ENC_u0_u1_n742 ), .A3(_AES_ENC_u0_u1_n741 ), .ZN(_AES_ENC_u0_u1_n744 ) );
NOR2_X2 _AES_ENC_u0_u1_U398  ( .A1(_AES_ENC_u0_u1_n697 ), .A2(_AES_ENC_u0_u1_n658 ), .ZN(_AES_ENC_u0_u1_n659 ) );
NOR3_X2 _AES_ENC_u0_u1_U397  ( .A1(_AES_ENC_u0_u1_n959 ), .A2(_AES_ENC_u0_u1_n572 ), .A3(_AES_ENC_u0_u1_n609 ), .ZN(_AES_ENC_u0_u1_n768 ) );
NOR2_X2 _AES_ENC_u0_u1_U396  ( .A1(_AES_ENC_u0_u1_n598 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n885 ) );
NOR2_X2 _AES_ENC_u0_u1_U393  ( .A1(_AES_ENC_u0_u1_n623 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n882 ) );
NOR2_X2 _AES_ENC_u0_u1_U390  ( .A1(_AES_ENC_u0_u1_n1053 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n884 ) );
NOR4_X2 _AES_ENC_u0_u1_U389  ( .A1(_AES_ENC_u0_u1_n885 ), .A2(_AES_ENC_u0_u1_n884 ), .A3(_AES_ENC_u0_u1_n883 ), .A4(_AES_ENC_u0_u1_n882 ), .ZN(_AES_ENC_u0_u1_n886 ) );
NOR2_X2 _AES_ENC_u0_u1_U388  ( .A1(_AES_ENC_u0_u1_n1078 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n1033 ) );
NOR2_X2 _AES_ENC_u0_u1_U387  ( .A1(_AES_ENC_u0_u1_n1031 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n1032 ) );
NOR3_X2 _AES_ENC_u0_u1_U386  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n1025 ), .A3(_AES_ENC_u0_u1_n1074 ), .ZN(_AES_ENC_u0_u1_n1035 ) );
NOR4_X2 _AES_ENC_u0_u1_U385  ( .A1(_AES_ENC_u0_u1_n1035 ), .A2(_AES_ENC_u0_u1_n1034 ), .A3(_AES_ENC_u0_u1_n1033 ), .A4(_AES_ENC_u0_u1_n1032 ), .ZN(_AES_ENC_u0_u1_n1036 ) );
NOR2_X2 _AES_ENC_u0_u1_U384  ( .A1(_AES_ENC_u0_u1_n825 ), .A2(_AES_ENC_u0_u1_n578 ), .ZN(_AES_ENC_u0_u1_n830 ) );
NOR2_X2 _AES_ENC_u0_u1_U383  ( .A1(_AES_ENC_u0_u1_n827 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n829 ) );
NOR2_X2 _AES_ENC_u0_u1_U382  ( .A1(_AES_ENC_u0_u1_n572 ), .A2(_AES_ENC_u0_u1_n579 ), .ZN(_AES_ENC_u0_u1_n828 ) );
NOR4_X2 _AES_ENC_u0_u1_U374  ( .A1(_AES_ENC_u0_u1_n831 ), .A2(_AES_ENC_u0_u1_n830 ), .A3(_AES_ENC_u0_u1_n829 ), .A4(_AES_ENC_u0_u1_n828 ), .ZN(_AES_ENC_u0_u1_n832 ) );
NOR2_X2 _AES_ENC_u0_u1_U373  ( .A1(_AES_ENC_u0_u1_n598 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n1107 ) );
NOR2_X2 _AES_ENC_u0_u1_U372  ( .A1(_AES_ENC_u0_u1_n1102 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n1106 ) );
NOR2_X2 _AES_ENC_u0_u1_U370  ( .A1(_AES_ENC_u0_u1_n1103 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n1105 ) );
NOR4_X2 _AES_ENC_u0_u1_U369  ( .A1(_AES_ENC_u0_u1_n1107 ), .A2(_AES_ENC_u0_u1_n1106 ), .A3(_AES_ENC_u0_u1_n1105 ), .A4(_AES_ENC_u0_u1_n1104 ), .ZN(_AES_ENC_u0_u1_n1108 ) );
NOR3_X2 _AES_ENC_u0_u1_U368  ( .A1(_AES_ENC_u0_u1_n959 ), .A2(_AES_ENC_u0_u1_n621 ), .A3(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n963 ) );
NOR2_X2 _AES_ENC_u0_u1_U367  ( .A1(_AES_ENC_u0_u1_n626 ), .A2(_AES_ENC_u0_u1_n627 ), .ZN(_AES_ENC_u0_u1_n1114 ) );
NOR3_X2 _AES_ENC_u0_u1_U366  ( .A1(_AES_ENC_u0_u1_n910 ), .A2(_AES_ENC_u0_u1_n1059 ), .A3(_AES_ENC_u0_u1_n611 ), .ZN(_AES_ENC_u0_u1_n1115 ) );
INV_X4 _AES_ENC_u0_u1_U365  ( .A(_AES_ENC_u0_u1_n1024 ), .ZN(_AES_ENC_u0_u1_n606 ) );
INV_X4 _AES_ENC_u0_u1_U364  ( .A(_AES_ENC_u0_u1_n1094 ), .ZN(_AES_ENC_u0_u1_n613 ) );
NOR2_X2 _AES_ENC_u0_u1_U363  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n931 ), .ZN(_AES_ENC_u0_u1_n1100 ) );
NOR2_X2 _AES_ENC_u0_u1_U354  ( .A1(_AES_ENC_u0_u1_n569 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n929 ) );
NOR2_X2 _AES_ENC_u0_u1_U353  ( .A1(_AES_ENC_u0_u1_n620 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n926 ) );
INV_X4 _AES_ENC_u0_u1_U352  ( .A(_AES_ENC_u0_u1_n1093 ), .ZN(_AES_ENC_u0_u1_n617 ) );
NOR2_X2 _AES_ENC_u0_u1_U351  ( .A1(_AES_ENC_u0_u1_n572 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n1095 ) );
NOR2_X2 _AES_ENC_u0_u1_U350  ( .A1(_AES_ENC_u0_u1_n609 ), .A2(_AES_ENC_u0_u1_n627 ), .ZN(_AES_ENC_u0_u1_n1010 ) );
NOR2_X2 _AES_ENC_u0_u1_U349  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n1103 ) );
NOR2_X2 _AES_ENC_u0_u1_U348  ( .A1(_AES_ENC_w3[9] ), .A2(_AES_ENC_u0_u1_n1120 ), .ZN(_AES_ENC_u0_u1_n1022 ) );
NOR2_X2 _AES_ENC_u0_u1_U347  ( .A1(_AES_ENC_u0_u1_n619 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n911 ) );
NOR2_X2 _AES_ENC_u0_u1_U346  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_u0_u1_n1025 ), .ZN(_AES_ENC_u0_u1_n826 ) );
NOR2_X2 _AES_ENC_u0_u1_U345  ( .A1(_AES_ENC_u0_u1_n626 ), .A2(_AES_ENC_u0_u1_n607 ), .ZN(_AES_ENC_u0_u1_n1072 ) );
NOR2_X2 _AES_ENC_u0_u1_U338  ( .A1(_AES_ENC_u0_u1_n627 ), .A2(_AES_ENC_u0_u1_n616 ), .ZN(_AES_ENC_u0_u1_n956 ) );
NOR2_X2 _AES_ENC_u0_u1_U335  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_u0_u1_n624 ), .ZN(_AES_ENC_u0_u1_n1121 ) );
NOR2_X2 _AES_ENC_u0_u1_U329  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_u0_u1_n624 ), .ZN(_AES_ENC_u0_u1_n1058 ) );
NOR2_X2 _AES_ENC_u0_u1_U328  ( .A1(_AES_ENC_u0_u1_n625 ), .A2(_AES_ENC_u0_u1_n611 ), .ZN(_AES_ENC_u0_u1_n1073 ) );
NOR2_X2 _AES_ENC_u0_u1_U327  ( .A1(_AES_ENC_w3[9] ), .A2(_AES_ENC_u0_u1_n1025 ), .ZN(_AES_ENC_u0_u1_n1054 ) );
NOR2_X2 _AES_ENC_u0_u1_U325  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_u0_u1_n931 ), .ZN(_AES_ENC_u0_u1_n1029 ) );
NOR2_X2 _AES_ENC_u0_u1_U324  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n1056 ) );
NOR2_X2 _AES_ENC_u0_u1_U319  ( .A1(_AES_ENC_u0_u1_n614 ), .A2(_AES_ENC_u0_u1_n626 ), .ZN(_AES_ENC_u0_u1_n1050 ) );
NOR2_X2 _AES_ENC_u0_u1_U318  ( .A1(_AES_ENC_u0_u1_n1121 ), .A2(_AES_ENC_u0_u1_n1025 ), .ZN(_AES_ENC_u0_u1_n1120 ) );
NOR2_X2 _AES_ENC_u0_u1_U317  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_u0_u1_n572 ), .ZN(_AES_ENC_u0_u1_n1074 ) );
NOR2_X2 _AES_ENC_u0_u1_U316  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n584 ), .ZN(_AES_ENC_u0_u1_n838 ) );
NOR2_X2 _AES_ENC_u0_u1_U315  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n602 ), .ZN(_AES_ENC_u0_u1_n837 ) );
NOR2_X2 _AES_ENC_u0_u1_U314  ( .A1(_AES_ENC_u0_u1_n838 ), .A2(_AES_ENC_u0_u1_n837 ), .ZN(_AES_ENC_u0_u1_n845 ) );
NOR2_X2 _AES_ENC_u0_u1_U312  ( .A1(_AES_ENC_u0_u1_n1058 ), .A2(_AES_ENC_u0_u1_n1054 ), .ZN(_AES_ENC_u0_u1_n878 ) );
NOR2_X2 _AES_ENC_u0_u1_U311  ( .A1(_AES_ENC_u0_u1_n878 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n879 ) );
NOR2_X2 _AES_ENC_u0_u1_U310  ( .A1(_AES_ENC_u0_u1_n880 ), .A2(_AES_ENC_u0_u1_n879 ), .ZN(_AES_ENC_u0_u1_n887 ) );
NOR3_X2 _AES_ENC_u0_u1_U309  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n1091 ), .A3(_AES_ENC_u0_u1_n1022 ), .ZN(_AES_ENC_u0_u1_n720 ) );
NOR3_X2 _AES_ENC_u0_u1_U303  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n1054 ), .A3(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n719 ) );
NOR2_X2 _AES_ENC_u0_u1_U302  ( .A1(_AES_ENC_u0_u1_n720 ), .A2(_AES_ENC_u0_u1_n719 ), .ZN(_AES_ENC_u0_u1_n726 ) );
NOR2_X2 _AES_ENC_u0_u1_U300  ( .A1(_AES_ENC_u0_u1_n614 ), .A2(_AES_ENC_u0_u1_n591 ), .ZN(_AES_ENC_u0_u1_n865 ) );
NOR2_X2 _AES_ENC_u0_u1_U299  ( .A1(_AES_ENC_u0_u1_n1059 ), .A2(_AES_ENC_u0_u1_n1058 ), .ZN(_AES_ENC_u0_u1_n1060 ) );
NOR2_X2 _AES_ENC_u0_u1_U298  ( .A1(_AES_ENC_u0_u1_n1095 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n668 ) );
NOR2_X2 _AES_ENC_u0_u1_U297  ( .A1(_AES_ENC_u0_u1_n826 ), .A2(_AES_ENC_u0_u1_n573 ), .ZN(_AES_ENC_u0_u1_n750 ) );
NOR2_X2 _AES_ENC_u0_u1_U296  ( .A1(_AES_ENC_u0_u1_n750 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n751 ) );
NOR2_X2 _AES_ENC_u0_u1_U295  ( .A1(_AES_ENC_u0_u1_n907 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n908 ) );
NOR2_X2 _AES_ENC_u0_u1_U294  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n588 ), .ZN(_AES_ENC_u0_u1_n957 ) );
NOR2_X2 _AES_ENC_u0_u1_U293  ( .A1(_AES_ENC_u0_u1_n990 ), .A2(_AES_ENC_u0_u1_n926 ), .ZN(_AES_ENC_u0_u1_n780 ) );
NOR2_X2 _AES_ENC_u0_u1_U292  ( .A1(_AES_ENC_u0_u1_n1022 ), .A2(_AES_ENC_u0_u1_n1058 ), .ZN(_AES_ENC_u0_u1_n740 ) );
NOR2_X2 _AES_ENC_u0_u1_U291  ( .A1(_AES_ENC_u0_u1_n740 ), .A2(_AES_ENC_u0_u1_n616 ), .ZN(_AES_ENC_u0_u1_n742 ) );
NOR2_X2 _AES_ENC_u0_u1_U290  ( .A1(_AES_ENC_u0_u1_n1098 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n1099 ) );
NOR2_X2 _AES_ENC_u0_u1_U284  ( .A1(_AES_ENC_u0_u1_n1120 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n993 ) );
NOR2_X2 _AES_ENC_u0_u1_U283  ( .A1(_AES_ENC_u0_u1_n993 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n994 ) );
NOR2_X2 _AES_ENC_u0_u1_U282  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n620 ), .ZN(_AES_ENC_u0_u1_n1026 ) );
NOR2_X2 _AES_ENC_u0_u1_U281  ( .A1(_AES_ENC_u0_u1_n573 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n1027 ) );
NOR2_X2 _AES_ENC_u0_u1_U280  ( .A1(_AES_ENC_u0_u1_n1027 ), .A2(_AES_ENC_u0_u1_n1026 ), .ZN(_AES_ENC_u0_u1_n1028 ) );
NOR2_X2 _AES_ENC_u0_u1_U279  ( .A1(_AES_ENC_u0_u1_n1029 ), .A2(_AES_ENC_u0_u1_n1028 ), .ZN(_AES_ENC_u0_u1_n1034 ) );
NOR2_X2 _AES_ENC_u0_u1_U273  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n1071 ), .ZN(_AES_ENC_u0_u1_n669 ) );
NOR2_X2 _AES_ENC_u0_u1_U272  ( .A1(_AES_ENC_u0_u1_n1056 ), .A2(_AES_ENC_u0_u1_n990 ), .ZN(_AES_ENC_u0_u1_n991 ) );
NOR2_X2 _AES_ENC_u0_u1_U271  ( .A1(_AES_ENC_u0_u1_n991 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n995 ) );
NOR4_X2 _AES_ENC_u0_u1_U270  ( .A1(_AES_ENC_u0_u1_n757 ), .A2(_AES_ENC_u0_u1_n756 ), .A3(_AES_ENC_u0_u1_n755 ), .A4(_AES_ENC_u0_u1_n754 ), .ZN(_AES_ENC_u0_u1_n758 ) );
NOR2_X2 _AES_ENC_u0_u1_U269  ( .A1(_AES_ENC_u0_u1_n752 ), .A2(_AES_ENC_u0_u1_n751 ), .ZN(_AES_ENC_u0_u1_n759 ) );
NOR2_X2 _AES_ENC_u0_u1_U268  ( .A1(_AES_ENC_u0_u1_n607 ), .A2(_AES_ENC_u0_u1_n590 ), .ZN(_AES_ENC_u0_u1_n1008 ) );
NOR2_X2 _AES_ENC_u0_u1_U267  ( .A1(_AES_ENC_u0_u1_n606 ), .A2(_AES_ENC_u0_u1_n906 ), .ZN(_AES_ENC_u0_u1_n741 ) );
NOR2_X2 _AES_ENC_u0_u1_U263  ( .A1(_AES_ENC_u0_u1_n1054 ), .A2(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n763 ) );
NOR2_X2 _AES_ENC_u0_u1_U262  ( .A1(_AES_ENC_u0_u1_n763 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n769 ) );
NOR2_X2 _AES_ENC_u0_u1_U258  ( .A1(_AES_ENC_u0_u1_n839 ), .A2(_AES_ENC_u0_u1_n582 ), .ZN(_AES_ENC_u0_u1_n693 ) );
NOR2_X2 _AES_ENC_u0_u1_U255  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n577 ), .ZN(_AES_ENC_u0_u1_n1007 ) );
NOR2_X2 _AES_ENC_u0_u1_U254  ( .A1(_AES_ENC_u0_u1_n609 ), .A2(_AES_ENC_u0_u1_n580 ), .ZN(_AES_ENC_u0_u1_n1123 ) );
NOR2_X2 _AES_ENC_u0_u1_U253  ( .A1(_AES_ENC_u0_u1_n780 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n784 ) );
NOR2_X2 _AES_ENC_u0_u1_U252  ( .A1(_AES_ENC_u0_u1_n1117 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n782 ) );
NOR2_X2 _AES_ENC_u0_u1_U251  ( .A1(_AES_ENC_u0_u1_n781 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n783 ) );
NOR4_X2 _AES_ENC_u0_u1_U250  ( .A1(_AES_ENC_u0_u1_n880 ), .A2(_AES_ENC_u0_u1_n784 ), .A3(_AES_ENC_u0_u1_n783 ), .A4(_AES_ENC_u0_u1_n782 ), .ZN(_AES_ENC_u0_u1_n785 ) );
NOR2_X2 _AES_ENC_u0_u1_U243  ( .A1(_AES_ENC_u0_u1_n609 ), .A2(_AES_ENC_u0_u1_n590 ), .ZN(_AES_ENC_u0_u1_n710 ) );
INV_X4 _AES_ENC_u0_u1_U242  ( .A(_AES_ENC_u0_u1_n1029 ), .ZN(_AES_ENC_u0_u1_n582 ) );
NOR2_X2 _AES_ENC_u0_u1_U241  ( .A1(_AES_ENC_u0_u1_n593 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n1125 ) );
NOR2_X2 _AES_ENC_u0_u1_U240  ( .A1(_AES_ENC_u0_u1_n616 ), .A2(_AES_ENC_u0_u1_n580 ), .ZN(_AES_ENC_u0_u1_n771 ) );
NOR2_X2 _AES_ENC_u0_u1_U239  ( .A1(_AES_ENC_u0_u1_n616 ), .A2(_AES_ENC_u0_u1_n597 ), .ZN(_AES_ENC_u0_u1_n883 ) );
NOR2_X2 _AES_ENC_u0_u1_U238  ( .A1(_AES_ENC_u0_u1_n911 ), .A2(_AES_ENC_u0_u1_n910 ), .ZN(_AES_ENC_u0_u1_n912 ) );
NOR2_X2 _AES_ENC_u0_u1_U237  ( .A1(_AES_ENC_u0_u1_n912 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n916 ) );
NOR2_X2 _AES_ENC_u0_u1_U236  ( .A1(_AES_ENC_u0_u1_n990 ), .A2(_AES_ENC_u0_u1_n929 ), .ZN(_AES_ENC_u0_u1_n892 ) );
NOR2_X2 _AES_ENC_u0_u1_U235  ( .A1(_AES_ENC_u0_u1_n892 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n893 ) );
NOR2_X2 _AES_ENC_u0_u1_U234  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n602 ), .ZN(_AES_ENC_u0_u1_n950 ) );
NOR2_X2 _AES_ENC_u0_u1_U229  ( .A1(_AES_ENC_u0_u1_n1079 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n1082 ) );
NOR2_X2 _AES_ENC_u0_u1_U228  ( .A1(_AES_ENC_u0_u1_n910 ), .A2(_AES_ENC_u0_u1_n1056 ), .ZN(_AES_ENC_u0_u1_n941 ) );
NOR2_X2 _AES_ENC_u0_u1_U227  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n1077 ), .ZN(_AES_ENC_u0_u1_n841 ) );
NOR2_X2 _AES_ENC_u0_u1_U226  ( .A1(_AES_ENC_u0_u1_n623 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n630 ) );
NOR2_X2 _AES_ENC_u0_u1_U225  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n602 ), .ZN(_AES_ENC_u0_u1_n806 ) );
NOR2_X2 _AES_ENC_u0_u1_U223  ( .A1(_AES_ENC_u0_u1_n623 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n948 ) );
NOR2_X2 _AES_ENC_u0_u1_U222  ( .A1(_AES_ENC_u0_u1_n606 ), .A2(_AES_ENC_u0_u1_n582 ), .ZN(_AES_ENC_u0_u1_n1104 ) );
NOR2_X2 _AES_ENC_u0_u1_U221  ( .A1(_AES_ENC_u0_u1_n1121 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n1122 ) );
NOR2_X2 _AES_ENC_u0_u1_U217  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n1023 ), .ZN(_AES_ENC_u0_u1_n756 ) );
NOR2_X2 _AES_ENC_u0_u1_U213  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n602 ), .ZN(_AES_ENC_u0_u1_n870 ) );
NOR2_X2 _AES_ENC_u0_u1_U212  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n569 ), .ZN(_AES_ENC_u0_u1_n947 ) );
NOR2_X2 _AES_ENC_u0_u1_U211  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n1077 ), .ZN(_AES_ENC_u0_u1_n1084 ) );
NOR2_X2 _AES_ENC_u0_u1_U210  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n855 ), .ZN(_AES_ENC_u0_u1_n709 ) );
NOR2_X2 _AES_ENC_u0_u1_U209  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n589 ), .ZN(_AES_ENC_u0_u1_n868 ) );
NOR2_X2 _AES_ENC_u0_u1_U208  ( .A1(_AES_ENC_u0_u1_n1120 ), .A2(_AES_ENC_u0_u1_n839 ), .ZN(_AES_ENC_u0_u1_n842 ) );
NOR2_X2 _AES_ENC_u0_u1_U207  ( .A1(_AES_ENC_u0_u1_n1120 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n1124 ) );
NOR2_X2 _AES_ENC_u0_u1_U201  ( .A1(_AES_ENC_u0_u1_n1120 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n696 ) );
NOR2_X2 _AES_ENC_u0_u1_U200  ( .A1(_AES_ENC_u0_u1_n1074 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n1076 ) );
NOR2_X2 _AES_ENC_u0_u1_U199  ( .A1(_AES_ENC_u0_u1_n1074 ), .A2(_AES_ENC_u0_u1_n620 ), .ZN(_AES_ENC_u0_u1_n781 ) );
NOR3_X2 _AES_ENC_u0_u1_U198  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n1056 ), .A3(_AES_ENC_u0_u1_n990 ), .ZN(_AES_ENC_u0_u1_n979 ) );
NOR3_X2 _AES_ENC_u0_u1_U197  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n1058 ), .A3(_AES_ENC_u0_u1_n1059 ), .ZN(_AES_ENC_u0_u1_n854 ) );
NOR2_X2 _AES_ENC_u0_u1_U196  ( .A1(_AES_ENC_u0_u1_n996 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n869 ) );
NOR2_X2 _AES_ENC_u0_u1_U195  ( .A1(_AES_ENC_u0_u1_n1056 ), .A2(_AES_ENC_u0_u1_n1074 ), .ZN(_AES_ENC_u0_u1_n1057 ) );
NOR3_X2 _AES_ENC_u0_u1_U194  ( .A1(_AES_ENC_u0_u1_n607 ), .A2(_AES_ENC_u0_u1_n1120 ), .A3(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n978 ) );
NOR2_X2 _AES_ENC_u0_u1_U187  ( .A1(_AES_ENC_u0_u1_n996 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n998 ) );
NOR2_X2 _AES_ENC_u0_u1_U186  ( .A1(_AES_ENC_u0_u1_n996 ), .A2(_AES_ENC_u0_u1_n911 ), .ZN(_AES_ENC_u0_u1_n1116 ) );
NOR2_X2 _AES_ENC_u0_u1_U185  ( .A1(_AES_ENC_u0_u1_n1074 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n754 ) );
NOR2_X2 _AES_ENC_u0_u1_U184  ( .A1(_AES_ENC_u0_u1_n926 ), .A2(_AES_ENC_u0_u1_n1103 ), .ZN(_AES_ENC_u0_u1_n977 ) );
NOR2_X2 _AES_ENC_u0_u1_U183  ( .A1(_AES_ENC_u0_u1_n839 ), .A2(_AES_ENC_u0_u1_n824 ), .ZN(_AES_ENC_u0_u1_n1092 ) );
NOR2_X2 _AES_ENC_u0_u1_U182  ( .A1(_AES_ENC_u0_u1_n573 ), .A2(_AES_ENC_u0_u1_n1074 ), .ZN(_AES_ENC_u0_u1_n684 ) );
NOR2_X2 _AES_ENC_u0_u1_U181  ( .A1(_AES_ENC_u0_u1_n826 ), .A2(_AES_ENC_u0_u1_n1059 ), .ZN(_AES_ENC_u0_u1_n907 ) );
NOR3_X2 _AES_ENC_u0_u1_U180  ( .A1(_AES_ENC_u0_u1_n625 ), .A2(_AES_ENC_u0_u1_n1115 ), .A3(_AES_ENC_u0_u1_n585 ), .ZN(_AES_ENC_u0_u1_n831 ) );
NOR3_X2 _AES_ENC_u0_u1_U174  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n1056 ), .A3(_AES_ENC_u0_u1_n990 ), .ZN(_AES_ENC_u0_u1_n896 ) );
NOR3_X2 _AES_ENC_u0_u1_U173  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n573 ), .A3(_AES_ENC_u0_u1_n1013 ), .ZN(_AES_ENC_u0_u1_n670 ) );
NOR3_X2 _AES_ENC_u0_u1_U172  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n1091 ), .A3(_AES_ENC_u0_u1_n1022 ), .ZN(_AES_ENC_u0_u1_n843 ) );
NOR2_X2 _AES_ENC_u0_u1_U171  ( .A1(_AES_ENC_u0_u1_n1029 ), .A2(_AES_ENC_u0_u1_n1095 ), .ZN(_AES_ENC_u0_u1_n735 ) );
NAND3_X2 _AES_ENC_u0_u1_U170  ( .A1(_AES_ENC_u0_u1_n569 ), .A2(_AES_ENC_u0_u1_n582 ), .A3(_AES_ENC_u0_u1_n681 ), .ZN(_AES_ENC_u0_u1_n691 ) );
NOR2_X2 _AES_ENC_u0_u1_U169  ( .A1(_AES_ENC_u0_u1_n683 ), .A2(_AES_ENC_u0_u1_n682 ), .ZN(_AES_ENC_u0_u1_n690 ) );
NOR4_X2 _AES_ENC_u0_u1_U168  ( .A1(_AES_ENC_u0_u1_n983 ), .A2(_AES_ENC_u0_u1_n698 ), .A3(_AES_ENC_u0_u1_n697 ), .A4(_AES_ENC_u0_u1_n696 ), .ZN(_AES_ENC_u0_u1_n699 ) );
NOR3_X2 _AES_ENC_u0_u1_U162  ( .A1(_AES_ENC_u0_u1_n695 ), .A2(_AES_ENC_u0_u1_n694 ), .A3(_AES_ENC_u0_u1_n693 ), .ZN(_AES_ENC_u0_u1_n700 ) );
NOR2_X2 _AES_ENC_u0_u1_U161  ( .A1(_AES_ENC_u0_u1_n1100 ), .A2(_AES_ENC_u0_u1_n854 ), .ZN(_AES_ENC_u0_u1_n860 ) );
NOR4_X2 _AES_ENC_u0_u1_U160  ( .A1(_AES_ENC_u0_u1_n896 ), .A2(_AES_ENC_u0_u1_n895 ), .A3(_AES_ENC_u0_u1_n894 ), .A4(_AES_ENC_u0_u1_n893 ), .ZN(_AES_ENC_u0_u1_n897 ) );
NOR2_X2 _AES_ENC_u0_u1_U159  ( .A1(_AES_ENC_u0_u1_n866 ), .A2(_AES_ENC_u0_u1_n865 ), .ZN(_AES_ENC_u0_u1_n872 ) );
NOR4_X2 _AES_ENC_u0_u1_U158  ( .A1(_AES_ENC_u0_u1_n870 ), .A2(_AES_ENC_u0_u1_n869 ), .A3(_AES_ENC_u0_u1_n868 ), .A4(_AES_ENC_u0_u1_n867 ), .ZN(_AES_ENC_u0_u1_n871 ) );
NOR4_X2 _AES_ENC_u0_u1_U157  ( .A1(_AES_ENC_u0_u1_n963 ), .A2(_AES_ENC_u0_u1_n962 ), .A3(_AES_ENC_u0_u1_n961 ), .A4(_AES_ENC_u0_u1_n960 ), .ZN(_AES_ENC_u0_u1_n964 ) );
NOR2_X2 _AES_ENC_u0_u1_U156  ( .A1(_AES_ENC_u0_u1_n958 ), .A2(_AES_ENC_u0_u1_n957 ), .ZN(_AES_ENC_u0_u1_n965 ) );
NOR4_X2 _AES_ENC_u0_u1_U155  ( .A1(_AES_ENC_u0_u1_n950 ), .A2(_AES_ENC_u0_u1_n949 ), .A3(_AES_ENC_u0_u1_n948 ), .A4(_AES_ENC_u0_u1_n947 ), .ZN(_AES_ENC_u0_u1_n951 ) );
NOR2_X2 _AES_ENC_u0_u1_U154  ( .A1(_AES_ENC_u0_u1_n946 ), .A2(_AES_ENC_u0_u1_n945 ), .ZN(_AES_ENC_u0_u1_n952 ) );
NOR4_X2 _AES_ENC_u0_u1_U153  ( .A1(_AES_ENC_u0_u1_n983 ), .A2(_AES_ENC_u0_u1_n982 ), .A3(_AES_ENC_u0_u1_n981 ), .A4(_AES_ENC_u0_u1_n980 ), .ZN(_AES_ENC_u0_u1_n984 ) );
NOR2_X2 _AES_ENC_u0_u1_U152  ( .A1(_AES_ENC_u0_u1_n979 ), .A2(_AES_ENC_u0_u1_n978 ), .ZN(_AES_ENC_u0_u1_n985 ) );
NOR4_X2 _AES_ENC_u0_u1_U143  ( .A1(_AES_ENC_u0_u1_n1125 ), .A2(_AES_ENC_u0_u1_n1124 ), .A3(_AES_ENC_u0_u1_n1123 ), .A4(_AES_ENC_u0_u1_n1122 ), .ZN(_AES_ENC_u0_u1_n1126 ) );
NOR4_X2 _AES_ENC_u0_u1_U142  ( .A1(_AES_ENC_u0_u1_n1084 ), .A2(_AES_ENC_u0_u1_n1083 ), .A3(_AES_ENC_u0_u1_n1082 ), .A4(_AES_ENC_u0_u1_n1081 ), .ZN(_AES_ENC_u0_u1_n1085 ) );
NOR2_X2 _AES_ENC_u0_u1_U141  ( .A1(_AES_ENC_u0_u1_n1076 ), .A2(_AES_ENC_u0_u1_n1075 ), .ZN(_AES_ENC_u0_u1_n1086 ) );
NOR3_X2 _AES_ENC_u0_u1_U140  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n1054 ), .A3(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n961 ) );
NOR3_X2 _AES_ENC_u0_u1_U132  ( .A1(_AES_ENC_u0_u1_n620 ), .A2(_AES_ENC_u0_u1_n1074 ), .A3(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n671 ) );
NOR2_X2 _AES_ENC_u0_u1_U131  ( .A1(_AES_ENC_u0_u1_n1057 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n1062 ) );
NOR2_X2 _AES_ENC_u0_u1_U130  ( .A1(_AES_ENC_u0_u1_n1060 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n1061 ) );
NOR2_X2 _AES_ENC_u0_u1_U129  ( .A1(_AES_ENC_u0_u1_n1055 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n1063 ) );
NOR4_X2 _AES_ENC_u0_u1_U128  ( .A1(_AES_ENC_u0_u1_n1064 ), .A2(_AES_ENC_u0_u1_n1063 ), .A3(_AES_ENC_u0_u1_n1062 ), .A4(_AES_ENC_u0_u1_n1061 ), .ZN(_AES_ENC_u0_u1_n1065 ) );
NOR3_X2 _AES_ENC_u0_u1_U127  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n1120 ), .A3(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n918 ) );
NOR2_X2 _AES_ENC_u0_u1_U126  ( .A1(_AES_ENC_u0_u1_n914 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n915 ) );
NOR3_X2 _AES_ENC_u0_u1_U121  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n573 ), .A3(_AES_ENC_u0_u1_n1013 ), .ZN(_AES_ENC_u0_u1_n917 ) );
NOR4_X2 _AES_ENC_u0_u1_U120  ( .A1(_AES_ENC_u0_u1_n918 ), .A2(_AES_ENC_u0_u1_n917 ), .A3(_AES_ENC_u0_u1_n916 ), .A4(_AES_ENC_u0_u1_n915 ), .ZN(_AES_ENC_u0_u1_n919 ) );
NOR2_X2 _AES_ENC_u0_u1_U119  ( .A1(_AES_ENC_u0_u1_n735 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n687 ) );
NOR2_X2 _AES_ENC_u0_u1_U118  ( .A1(_AES_ENC_u0_u1_n684 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n688 ) );
NOR2_X2 _AES_ENC_u0_u1_U117  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n600 ), .ZN(_AES_ENC_u0_u1_n686 ) );
NOR4_X2 _AES_ENC_u0_u1_U116  ( .A1(_AES_ENC_u0_u1_n688 ), .A2(_AES_ENC_u0_u1_n687 ), .A3(_AES_ENC_u0_u1_n686 ), .A4(_AES_ENC_u0_u1_n685 ), .ZN(_AES_ENC_u0_u1_n689 ) );
NOR2_X2 _AES_ENC_u0_u1_U115  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n582 ), .ZN(_AES_ENC_u0_u1_n770 ) );
NOR2_X2 _AES_ENC_u0_u1_U106  ( .A1(_AES_ENC_u0_u1_n1103 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n772 ) );
NOR2_X2 _AES_ENC_u0_u1_U105  ( .A1(_AES_ENC_u0_u1_n610 ), .A2(_AES_ENC_u0_u1_n599 ), .ZN(_AES_ENC_u0_u1_n773 ) );
NOR4_X2 _AES_ENC_u0_u1_U104  ( .A1(_AES_ENC_u0_u1_n773 ), .A2(_AES_ENC_u0_u1_n772 ), .A3(_AES_ENC_u0_u1_n771 ), .A4(_AES_ENC_u0_u1_n770 ), .ZN(_AES_ENC_u0_u1_n774 ) );
NOR2_X2 _AES_ENC_u0_u1_U103  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n595 ), .ZN(_AES_ENC_u0_u1_n858 ) );
NOR2_X2 _AES_ENC_u0_u1_U102  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n855 ), .ZN(_AES_ENC_u0_u1_n857 ) );
NOR2_X2 _AES_ENC_u0_u1_U101  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n587 ), .ZN(_AES_ENC_u0_u1_n856 ) );
NOR4_X2 _AES_ENC_u0_u1_U100  ( .A1(_AES_ENC_u0_u1_n858 ), .A2(_AES_ENC_u0_u1_n857 ), .A3(_AES_ENC_u0_u1_n856 ), .A4(_AES_ENC_u0_u1_n958 ), .ZN(_AES_ENC_u0_u1_n859 ) );
NOR2_X2 _AES_ENC_u0_u1_U95  ( .A1(_AES_ENC_u0_u1_n583 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n814 ) );
NOR3_X2 _AES_ENC_u0_u1_U94  ( .A1(_AES_ENC_u0_u1_n606 ), .A2(_AES_ENC_u0_u1_n1058 ), .A3(_AES_ENC_u0_u1_n1059 ), .ZN(_AES_ENC_u0_u1_n815 ) );
NOR2_X2 _AES_ENC_u0_u1_U93  ( .A1(_AES_ENC_u0_u1_n907 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n813 ) );
NOR4_X2 _AES_ENC_u0_u1_U92  ( .A1(_AES_ENC_u0_u1_n815 ), .A2(_AES_ENC_u0_u1_n814 ), .A3(_AES_ENC_u0_u1_n813 ), .A4(_AES_ENC_u0_u1_n812 ), .ZN(_AES_ENC_u0_u1_n816 ) );
NOR2_X2 _AES_ENC_u0_u1_U91  ( .A1(_AES_ENC_u0_u1_n617 ), .A2(_AES_ENC_u0_u1_n569 ), .ZN(_AES_ENC_u0_u1_n721 ) );
NOR2_X2 _AES_ENC_u0_u1_U90  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n1096 ), .ZN(_AES_ENC_u0_u1_n722 ) );
NOR2_X2 _AES_ENC_u0_u1_U89  ( .A1(_AES_ENC_u0_u1_n1031 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n723 ) );
NOR4_X2 _AES_ENC_u0_u1_U88  ( .A1(_AES_ENC_u0_u1_n724 ), .A2(_AES_ENC_u0_u1_n723 ), .A3(_AES_ENC_u0_u1_n722 ), .A4(_AES_ENC_u0_u1_n721 ), .ZN(_AES_ENC_u0_u1_n725 ) );
NOR2_X2 _AES_ENC_u0_u1_U87  ( .A1(_AES_ENC_u0_u1_n911 ), .A2(_AES_ENC_u0_u1_n990 ), .ZN(_AES_ENC_u0_u1_n1009 ) );
NOR2_X2 _AES_ENC_u0_u1_U86  ( .A1(_AES_ENC_u0_u1_n1013 ), .A2(_AES_ENC_u0_u1_n573 ), .ZN(_AES_ENC_u0_u1_n1014 ) );
NOR2_X2 _AES_ENC_u0_u1_U81  ( .A1(_AES_ENC_u0_u1_n1014 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n1015 ) );
NOR4_X2 _AES_ENC_u0_u1_U80  ( .A1(_AES_ENC_u0_u1_n1016 ), .A2(_AES_ENC_u0_u1_n1015 ), .A3(_AES_ENC_u0_u1_n1119 ), .A4(_AES_ENC_u0_u1_n1046 ), .ZN(_AES_ENC_u0_u1_n1017 ) );
NOR2_X2 _AES_ENC_u0_u1_U79  ( .A1(_AES_ENC_u0_u1_n606 ), .A2(_AES_ENC_u0_u1_n589 ), .ZN(_AES_ENC_u0_u1_n997 ) );
NOR2_X2 _AES_ENC_u0_u1_U78  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n577 ), .ZN(_AES_ENC_u0_u1_n1000 ) );
NOR2_X2 _AES_ENC_u0_u1_U74  ( .A1(_AES_ENC_u0_u1_n616 ), .A2(_AES_ENC_u0_u1_n1096 ), .ZN(_AES_ENC_u0_u1_n999 ) );
NOR4_X2 _AES_ENC_u0_u1_U73  ( .A1(_AES_ENC_u0_u1_n1000 ), .A2(_AES_ENC_u0_u1_n999 ), .A3(_AES_ENC_u0_u1_n998 ), .A4(_AES_ENC_u0_u1_n997 ), .ZN(_AES_ENC_u0_u1_n1001 ) );
NOR2_X2 _AES_ENC_u0_u1_U72  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n1096 ), .ZN(_AES_ENC_u0_u1_n697 ) );
NOR2_X2 _AES_ENC_u0_u1_U71  ( .A1(_AES_ENC_u0_u1_n620 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n958 ) );
NOR2_X2 _AES_ENC_u0_u1_U65  ( .A1(_AES_ENC_u0_u1_n911 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n983 ) );
NOR2_X2 _AES_ENC_u0_u1_U64  ( .A1(_AES_ENC_u0_u1_n1054 ), .A2(_AES_ENC_u0_u1_n1103 ), .ZN(_AES_ENC_u0_u1_n1031 ) );
INV_X4 _AES_ENC_u0_u1_U63  ( .A(_AES_ENC_u0_u1_n1050 ), .ZN(_AES_ENC_u0_u1_n612 ) );
INV_X4 _AES_ENC_u0_u1_U62  ( .A(_AES_ENC_u0_u1_n1072 ), .ZN(_AES_ENC_u0_u1_n605 ) );
INV_X4 _AES_ENC_u0_u1_U61  ( .A(_AES_ENC_u0_u1_n1073 ), .ZN(_AES_ENC_u0_u1_n604 ) );
NOR2_X2 _AES_ENC_u0_u1_U59  ( .A1(_AES_ENC_u0_u1_n582 ), .A2(_AES_ENC_u0_u1_n613 ), .ZN(_AES_ENC_u0_u1_n880 ) );
NOR3_X2 _AES_ENC_u0_u1_U58  ( .A1(_AES_ENC_u0_u1_n826 ), .A2(_AES_ENC_u0_u1_n1121 ), .A3(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n946 ) );
INV_X4 _AES_ENC_u0_u1_U57  ( .A(_AES_ENC_u0_u1_n1010 ), .ZN(_AES_ENC_u0_u1_n608 ) );
NOR3_X2 _AES_ENC_u0_u1_U50  ( .A1(_AES_ENC_u0_u1_n573 ), .A2(_AES_ENC_u0_u1_n1029 ), .A3(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n1119 ) );
INV_X4 _AES_ENC_u0_u1_U49  ( .A(_AES_ENC_u0_u1_n956 ), .ZN(_AES_ENC_u0_u1_n615 ) );
NOR2_X2 _AES_ENC_u0_u1_U48  ( .A1(_AES_ENC_u0_u1_n623 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n1013 ) );
NOR2_X2 _AES_ENC_u0_u1_U47  ( .A1(_AES_ENC_u0_u1_n620 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n910 ) );
NOR2_X2 _AES_ENC_u0_u1_U46  ( .A1(_AES_ENC_u0_u1_n569 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n1091 ) );
NOR2_X2 _AES_ENC_u0_u1_U45  ( .A1(_AES_ENC_u0_u1_n622 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n990 ) );
NOR2_X2 _AES_ENC_u0_u1_U44  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_u0_u1_n1121 ), .ZN(_AES_ENC_u0_u1_n996 ) );
NOR2_X2 _AES_ENC_u0_u1_U43  ( .A1(_AES_ENC_u0_u1_n610 ), .A2(_AES_ENC_u0_u1_n600 ), .ZN(_AES_ENC_u0_u1_n628 ) );
NOR2_X2 _AES_ENC_u0_u1_U42  ( .A1(_AES_ENC_u0_u1_n576 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n866 ) );
NOR2_X2 _AES_ENC_u0_u1_U41  ( .A1(_AES_ENC_u0_u1_n603 ), .A2(_AES_ENC_u0_u1_n610 ), .ZN(_AES_ENC_u0_u1_n1006 ) );
NOR2_X2 _AES_ENC_u0_u1_U36  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n1117 ), .ZN(_AES_ENC_u0_u1_n1118 ) );
NOR2_X2 _AES_ENC_u0_u1_U35  ( .A1(_AES_ENC_u0_u1_n1119 ), .A2(_AES_ENC_u0_u1_n1118 ), .ZN(_AES_ENC_u0_u1_n1127 ) );
NOR2_X2 _AES_ENC_u0_u1_U34  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n594 ), .ZN(_AES_ENC_u0_u1_n629 ) );
NOR2_X2 _AES_ENC_u0_u1_U33  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n906 ), .ZN(_AES_ENC_u0_u1_n909 ) );
NOR2_X2 _AES_ENC_u0_u1_U32  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n597 ), .ZN(_AES_ENC_u0_u1_n658 ) );
NOR2_X2 _AES_ENC_u0_u1_U31  ( .A1(_AES_ENC_u0_u1_n1116 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n695 ) );
NOR2_X2 _AES_ENC_u0_u1_U30  ( .A1(_AES_ENC_u0_u1_n1078 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n1083 ) );
NOR2_X2 _AES_ENC_u0_u1_U29  ( .A1(_AES_ENC_u0_u1_n941 ), .A2(_AES_ENC_u0_u1_n608 ), .ZN(_AES_ENC_u0_u1_n724 ) );
NOR2_X2 _AES_ENC_u0_u1_U24  ( .A1(_AES_ENC_u0_u1_n576 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n840 ) );
NOR2_X2 _AES_ENC_u0_u1_U23  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n593 ), .ZN(_AES_ENC_u0_u1_n633 ) );
NOR2_X2 _AES_ENC_u0_u1_U21  ( .A1(_AES_ENC_u0_u1_n1009 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n960 ) );
NOR2_X2 _AES_ENC_u0_u1_U20  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n1045 ), .ZN(_AES_ENC_u0_u1_n812 ) );
NOR2_X2 _AES_ENC_u0_u1_U19  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n1080 ), .ZN(_AES_ENC_u0_u1_n1081 ) );
NOR2_X2 _AES_ENC_u0_u1_U18  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n601 ), .ZN(_AES_ENC_u0_u1_n982 ) );
NOR2_X2 _AES_ENC_u0_u1_U17  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n594 ), .ZN(_AES_ENC_u0_u1_n757 ) );
NOR2_X2 _AES_ENC_u0_u1_U16  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n590 ), .ZN(_AES_ENC_u0_u1_n698 ) );
NOR2_X2 _AES_ENC_u0_u1_U15  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n619 ), .ZN(_AES_ENC_u0_u1_n708 ) );
NOR2_X2 _AES_ENC_u0_u1_U10  ( .A1(_AES_ENC_u0_u1_n619 ), .A2(_AES_ENC_u0_u1_n604 ), .ZN(_AES_ENC_u0_u1_n803 ) );
NOR2_X2 _AES_ENC_u0_u1_U9  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n881 ), .ZN(_AES_ENC_u0_u1_n711 ) );
NOR2_X2 _AES_ENC_u0_u1_U8  ( .A1(_AES_ENC_u0_u1_n615 ), .A2(_AES_ENC_u0_u1_n582 ), .ZN(_AES_ENC_u0_u1_n867 ) );
NOR2_X2 _AES_ENC_u0_u1_U7  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n599 ), .ZN(_AES_ENC_u0_u1_n804 ) );
NOR2_X2 _AES_ENC_u0_u1_U6  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n620 ), .ZN(_AES_ENC_u0_u1_n1046 ) );
OR2_X4 _AES_ENC_u0_u1_U5  ( .A1(_AES_ENC_u0_u1_n624 ), .A2(_AES_ENC_w3[9] ),.ZN(_AES_ENC_u0_u1_n570 ) );
OR2_X4 _AES_ENC_u0_u1_U4  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_w3[12] ),.ZN(_AES_ENC_u0_u1_n569 ) );
NAND2_X2 _AES_ENC_u0_u1_U514  ( .A1(_AES_ENC_u0_u1_n1121 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n1030 ) );
AND2_X2 _AES_ENC_u0_u1_U513  ( .A1(_AES_ENC_u0_u1_n597 ), .A2(_AES_ENC_u0_u1_n1030 ), .ZN(_AES_ENC_u0_u1_n1049 ) );
NAND2_X2 _AES_ENC_u0_u1_U511  ( .A1(_AES_ENC_u0_u1_n1049 ), .A2(_AES_ENC_u0_u1_n794 ), .ZN(_AES_ENC_u0_u1_n637 ) );
AND2_X2 _AES_ENC_u0_u1_U493  ( .A1(_AES_ENC_u0_u1_n779 ), .A2(_AES_ENC_u0_u1_n996 ), .ZN(_AES_ENC_u0_u1_n632 ) );
NAND4_X2 _AES_ENC_u0_u1_U485  ( .A1(_AES_ENC_u0_u1_n637 ), .A2(_AES_ENC_u0_u1_n636 ), .A3(_AES_ENC_u0_u1_n635 ), .A4(_AES_ENC_u0_u1_n634 ), .ZN(_AES_ENC_u0_u1_n638 ) );
NAND2_X2 _AES_ENC_u0_u1_U484  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n638 ), .ZN(_AES_ENC_u0_u1_n679 ) );
NAND2_X2 _AES_ENC_u0_u1_U481  ( .A1(_AES_ENC_u0_u1_n1094 ), .A2(_AES_ENC_u0_u1_n591 ), .ZN(_AES_ENC_u0_u1_n648 ) );
NAND2_X2 _AES_ENC_u0_u1_U476  ( .A1(_AES_ENC_u0_u1_n601 ), .A2(_AES_ENC_u0_u1_n590 ), .ZN(_AES_ENC_u0_u1_n762 ) );
NAND2_X2 _AES_ENC_u0_u1_U475  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n762 ), .ZN(_AES_ENC_u0_u1_n647 ) );
NAND4_X2 _AES_ENC_u0_u1_U457  ( .A1(_AES_ENC_u0_u1_n648 ), .A2(_AES_ENC_u0_u1_n647 ), .A3(_AES_ENC_u0_u1_n646 ), .A4(_AES_ENC_u0_u1_n645 ), .ZN(_AES_ENC_u0_u1_n649 ) );
NAND2_X2 _AES_ENC_u0_u1_U456  ( .A1(_AES_ENC_w3[8] ), .A2(_AES_ENC_u0_u1_n649 ), .ZN(_AES_ENC_u0_u1_n665 ) );
NAND2_X2 _AES_ENC_u0_u1_U454  ( .A1(_AES_ENC_u0_u1_n596 ), .A2(_AES_ENC_u0_u1_n623 ), .ZN(_AES_ENC_u0_u1_n855 ) );
NAND2_X2 _AES_ENC_u0_u1_U453  ( .A1(_AES_ENC_u0_u1_n587 ), .A2(_AES_ENC_u0_u1_n855 ), .ZN(_AES_ENC_u0_u1_n821 ) );
NAND2_X2 _AES_ENC_u0_u1_U452  ( .A1(_AES_ENC_u0_u1_n1093 ), .A2(_AES_ENC_u0_u1_n821 ), .ZN(_AES_ENC_u0_u1_n662 ) );
NAND2_X2 _AES_ENC_u0_u1_U451  ( .A1(_AES_ENC_u0_u1_n619 ), .A2(_AES_ENC_u0_u1_n589 ), .ZN(_AES_ENC_u0_u1_n650 ) );
NAND2_X2 _AES_ENC_u0_u1_U450  ( .A1(_AES_ENC_u0_u1_n956 ), .A2(_AES_ENC_u0_u1_n650 ), .ZN(_AES_ENC_u0_u1_n661 ) );
NAND2_X2 _AES_ENC_u0_u1_U449  ( .A1(_AES_ENC_u0_u1_n626 ), .A2(_AES_ENC_u0_u1_n627 ), .ZN(_AES_ENC_u0_u1_n839 ) );
OR2_X2 _AES_ENC_u0_u1_U446  ( .A1(_AES_ENC_u0_u1_n839 ), .A2(_AES_ENC_u0_u1_n932 ), .ZN(_AES_ENC_u0_u1_n656 ) );
NAND2_X2 _AES_ENC_u0_u1_U445  ( .A1(_AES_ENC_u0_u1_n621 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n1096 ) );
NAND2_X2 _AES_ENC_u0_u1_U444  ( .A1(_AES_ENC_u0_u1_n1030 ), .A2(_AES_ENC_u0_u1_n1096 ), .ZN(_AES_ENC_u0_u1_n651 ) );
NAND2_X2 _AES_ENC_u0_u1_U443  ( .A1(_AES_ENC_u0_u1_n1114 ), .A2(_AES_ENC_u0_u1_n651 ), .ZN(_AES_ENC_u0_u1_n655 ) );
OR3_X2 _AES_ENC_u0_u1_U440  ( .A1(_AES_ENC_u0_u1_n1079 ), .A2(_AES_ENC_w3[15] ), .A3(_AES_ENC_u0_u1_n626 ), .ZN(_AES_ENC_u0_u1_n654 ) );
NAND2_X2 _AES_ENC_u0_u1_U439  ( .A1(_AES_ENC_u0_u1_n593 ), .A2(_AES_ENC_u0_u1_n601 ), .ZN(_AES_ENC_u0_u1_n652 ) );
NAND4_X2 _AES_ENC_u0_u1_U437  ( .A1(_AES_ENC_u0_u1_n656 ), .A2(_AES_ENC_u0_u1_n655 ), .A3(_AES_ENC_u0_u1_n654 ), .A4(_AES_ENC_u0_u1_n653 ), .ZN(_AES_ENC_u0_u1_n657 ) );
NAND2_X2 _AES_ENC_u0_u1_U436  ( .A1(_AES_ENC_w3[10] ), .A2(_AES_ENC_u0_u1_n657 ), .ZN(_AES_ENC_u0_u1_n660 ) );
NAND4_X2 _AES_ENC_u0_u1_U432  ( .A1(_AES_ENC_u0_u1_n662 ), .A2(_AES_ENC_u0_u1_n661 ), .A3(_AES_ENC_u0_u1_n660 ), .A4(_AES_ENC_u0_u1_n659 ), .ZN(_AES_ENC_u0_u1_n663 ) );
NAND2_X2 _AES_ENC_u0_u1_U431  ( .A1(_AES_ENC_u0_u1_n663 ), .A2(_AES_ENC_u0_u1_n574 ), .ZN(_AES_ENC_u0_u1_n664 ) );
NAND2_X2 _AES_ENC_u0_u1_U430  ( .A1(_AES_ENC_u0_u1_n665 ), .A2(_AES_ENC_u0_u1_n664 ), .ZN(_AES_ENC_u0_u1_n666 ) );
NAND2_X2 _AES_ENC_u0_u1_U429  ( .A1(_AES_ENC_w3[14] ), .A2(_AES_ENC_u0_u1_n666 ), .ZN(_AES_ENC_u0_u1_n678 ) );
NAND2_X2 _AES_ENC_u0_u1_U426  ( .A1(_AES_ENC_u0_u1_n735 ), .A2(_AES_ENC_u0_u1_n1093 ), .ZN(_AES_ENC_u0_u1_n675 ) );
NAND2_X2 _AES_ENC_u0_u1_U425  ( .A1(_AES_ENC_u0_u1_n588 ), .A2(_AES_ENC_u0_u1_n597 ), .ZN(_AES_ENC_u0_u1_n1045 ) );
OR2_X2 _AES_ENC_u0_u1_U424  ( .A1(_AES_ENC_u0_u1_n1045 ), .A2(_AES_ENC_u0_u1_n605 ), .ZN(_AES_ENC_u0_u1_n674 ) );
NAND2_X2 _AES_ENC_u0_u1_U423  ( .A1(_AES_ENC_w3[9] ), .A2(_AES_ENC_u0_u1_n620 ), .ZN(_AES_ENC_u0_u1_n667 ) );
NAND2_X2 _AES_ENC_u0_u1_U422  ( .A1(_AES_ENC_u0_u1_n619 ), .A2(_AES_ENC_u0_u1_n667 ), .ZN(_AES_ENC_u0_u1_n1071 ) );
NAND4_X2 _AES_ENC_u0_u1_U412  ( .A1(_AES_ENC_u0_u1_n675 ), .A2(_AES_ENC_u0_u1_n674 ), .A3(_AES_ENC_u0_u1_n673 ), .A4(_AES_ENC_u0_u1_n672 ), .ZN(_AES_ENC_u0_u1_n676 ) );
NAND2_X2 _AES_ENC_u0_u1_U411  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n676 ), .ZN(_AES_ENC_u0_u1_n677 ) );
NAND2_X2 _AES_ENC_u0_u1_U408  ( .A1(_AES_ENC_u0_u1_n800 ), .A2(_AES_ENC_u0_u1_n1022 ), .ZN(_AES_ENC_u0_u1_n680 ) );
NAND2_X2 _AES_ENC_u0_u1_U407  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n680 ), .ZN(_AES_ENC_u0_u1_n681 ) );
AND2_X2 _AES_ENC_u0_u1_U402  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n684 ), .ZN(_AES_ENC_u0_u1_n682 ) );
NAND4_X2 _AES_ENC_u0_u1_U395  ( .A1(_AES_ENC_u0_u1_n691 ), .A2(_AES_ENC_u0_u1_n581 ), .A3(_AES_ENC_u0_u1_n690 ), .A4(_AES_ENC_u0_u1_n689 ), .ZN(_AES_ENC_u0_u1_n692 ) );
NAND2_X2 _AES_ENC_u0_u1_U394  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n692 ), .ZN(_AES_ENC_u0_u1_n733 ) );
NAND2_X2 _AES_ENC_u0_u1_U392  ( .A1(_AES_ENC_u0_u1_n977 ), .A2(_AES_ENC_u0_u1_n1050 ), .ZN(_AES_ENC_u0_u1_n702 ) );
NAND2_X2 _AES_ENC_u0_u1_U391  ( .A1(_AES_ENC_u0_u1_n1093 ), .A2(_AES_ENC_u0_u1_n1045 ), .ZN(_AES_ENC_u0_u1_n701 ) );
NAND4_X2 _AES_ENC_u0_u1_U381  ( .A1(_AES_ENC_u0_u1_n702 ), .A2(_AES_ENC_u0_u1_n701 ), .A3(_AES_ENC_u0_u1_n700 ), .A4(_AES_ENC_u0_u1_n699 ), .ZN(_AES_ENC_u0_u1_n703 ) );
NAND2_X2 _AES_ENC_u0_u1_U380  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n703 ), .ZN(_AES_ENC_u0_u1_n732 ) );
AND2_X2 _AES_ENC_u0_u1_U379  ( .A1(_AES_ENC_w3[8] ), .A2(_AES_ENC_w3[14] ),.ZN(_AES_ENC_u0_u1_n1113 ) );
NAND2_X2 _AES_ENC_u0_u1_U378  ( .A1(_AES_ENC_u0_u1_n601 ), .A2(_AES_ENC_u0_u1_n1030 ), .ZN(_AES_ENC_u0_u1_n881 ) );
NAND2_X2 _AES_ENC_u0_u1_U377  ( .A1(_AES_ENC_u0_u1_n1093 ), .A2(_AES_ENC_u0_u1_n881 ), .ZN(_AES_ENC_u0_u1_n715 ) );
NAND2_X2 _AES_ENC_u0_u1_U376  ( .A1(_AES_ENC_u0_u1_n1010 ), .A2(_AES_ENC_u0_u1_n600 ), .ZN(_AES_ENC_u0_u1_n714 ) );
NAND2_X2 _AES_ENC_u0_u1_U375  ( .A1(_AES_ENC_u0_u1_n855 ), .A2(_AES_ENC_u0_u1_n588 ), .ZN(_AES_ENC_u0_u1_n1117 ) );
XNOR2_X2 _AES_ENC_u0_u1_U371  ( .A(_AES_ENC_u0_u1_n611 ), .B(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n824 ) );
NAND4_X2 _AES_ENC_u0_u1_U362  ( .A1(_AES_ENC_u0_u1_n715 ), .A2(_AES_ENC_u0_u1_n714 ), .A3(_AES_ENC_u0_u1_n713 ), .A4(_AES_ENC_u0_u1_n712 ), .ZN(_AES_ENC_u0_u1_n716 ) );
NAND2_X2 _AES_ENC_u0_u1_U361  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n716 ), .ZN(_AES_ENC_u0_u1_n731 ) );
AND2_X2 _AES_ENC_u0_u1_U360  ( .A1(_AES_ENC_w3[14] ), .A2(_AES_ENC_u0_u1_n574 ), .ZN(_AES_ENC_u0_u1_n1131 ) );
NAND2_X2 _AES_ENC_u0_u1_U359  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n717 ) );
NAND2_X2 _AES_ENC_u0_u1_U358  ( .A1(_AES_ENC_u0_u1_n1029 ), .A2(_AES_ENC_u0_u1_n717 ), .ZN(_AES_ENC_u0_u1_n728 ) );
NAND2_X2 _AES_ENC_u0_u1_U357  ( .A1(_AES_ENC_w3[9] ), .A2(_AES_ENC_u0_u1_n624 ), .ZN(_AES_ENC_u0_u1_n1097 ) );
NAND2_X2 _AES_ENC_u0_u1_U356  ( .A1(_AES_ENC_u0_u1_n603 ), .A2(_AES_ENC_u0_u1_n1097 ), .ZN(_AES_ENC_u0_u1_n718 ) );
NAND2_X2 _AES_ENC_u0_u1_U355  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n718 ), .ZN(_AES_ENC_u0_u1_n727 ) );
NAND4_X2 _AES_ENC_u0_u1_U344  ( .A1(_AES_ENC_u0_u1_n728 ), .A2(_AES_ENC_u0_u1_n727 ), .A3(_AES_ENC_u0_u1_n726 ), .A4(_AES_ENC_u0_u1_n725 ), .ZN(_AES_ENC_u0_u1_n729 ) );
NAND2_X2 _AES_ENC_u0_u1_U343  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n729 ), .ZN(_AES_ENC_u0_u1_n730 ) );
NAND4_X2 _AES_ENC_u0_u1_U342  ( .A1(_AES_ENC_u0_u1_n733 ), .A2(_AES_ENC_u0_u1_n732 ), .A3(_AES_ENC_u0_u1_n731 ), .A4(_AES_ENC_u0_u1_n730 ), .ZN(_AES_ENC_u0_subword[17] ) );
NAND2_X2 _AES_ENC_u0_u1_U341  ( .A1(_AES_ENC_w3[15] ), .A2(_AES_ENC_u0_u1_n611 ), .ZN(_AES_ENC_u0_u1_n734 ) );
NAND2_X2 _AES_ENC_u0_u1_U340  ( .A1(_AES_ENC_u0_u1_n734 ), .A2(_AES_ENC_u0_u1_n607 ), .ZN(_AES_ENC_u0_u1_n738 ) );
OR4_X2 _AES_ENC_u0_u1_U339  ( .A1(_AES_ENC_u0_u1_n738 ), .A2(_AES_ENC_u0_u1_n626 ), .A3(_AES_ENC_u0_u1_n826 ), .A4(_AES_ENC_u0_u1_n1121 ), .ZN(_AES_ENC_u0_u1_n746 ) );
NAND2_X2 _AES_ENC_u0_u1_U337  ( .A1(_AES_ENC_u0_u1_n1100 ), .A2(_AES_ENC_u0_u1_n587 ), .ZN(_AES_ENC_u0_u1_n992 ) );
OR2_X2 _AES_ENC_u0_u1_U336  ( .A1(_AES_ENC_u0_u1_n610 ), .A2(_AES_ENC_u0_u1_n735 ), .ZN(_AES_ENC_u0_u1_n737 ) );
NAND2_X2 _AES_ENC_u0_u1_U334  ( .A1(_AES_ENC_u0_u1_n619 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n753 ) );
NAND2_X2 _AES_ENC_u0_u1_U333  ( .A1(_AES_ENC_u0_u1_n582 ), .A2(_AES_ENC_u0_u1_n753 ), .ZN(_AES_ENC_u0_u1_n1080 ) );
NAND2_X2 _AES_ENC_u0_u1_U332  ( .A1(_AES_ENC_u0_u1_n1048 ), .A2(_AES_ENC_u0_u1_n576 ), .ZN(_AES_ENC_u0_u1_n736 ) );
NAND2_X2 _AES_ENC_u0_u1_U331  ( .A1(_AES_ENC_u0_u1_n737 ), .A2(_AES_ENC_u0_u1_n736 ), .ZN(_AES_ENC_u0_u1_n739 ) );
NAND2_X2 _AES_ENC_u0_u1_U330  ( .A1(_AES_ENC_u0_u1_n739 ), .A2(_AES_ENC_u0_u1_n738 ), .ZN(_AES_ENC_u0_u1_n745 ) );
NAND2_X2 _AES_ENC_u0_u1_U326  ( .A1(_AES_ENC_u0_u1_n1096 ), .A2(_AES_ENC_u0_u1_n590 ), .ZN(_AES_ENC_u0_u1_n906 ) );
NAND4_X2 _AES_ENC_u0_u1_U323  ( .A1(_AES_ENC_u0_u1_n746 ), .A2(_AES_ENC_u0_u1_n992 ), .A3(_AES_ENC_u0_u1_n745 ), .A4(_AES_ENC_u0_u1_n744 ), .ZN(_AES_ENC_u0_u1_n747 ) );
NAND2_X2 _AES_ENC_u0_u1_U322  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n747 ), .ZN(_AES_ENC_u0_u1_n793 ) );
NAND2_X2 _AES_ENC_u0_u1_U321  ( .A1(_AES_ENC_u0_u1_n584 ), .A2(_AES_ENC_u0_u1_n855 ), .ZN(_AES_ENC_u0_u1_n748 ) );
NAND2_X2 _AES_ENC_u0_u1_U320  ( .A1(_AES_ENC_u0_u1_n956 ), .A2(_AES_ENC_u0_u1_n748 ), .ZN(_AES_ENC_u0_u1_n760 ) );
NAND2_X2 _AES_ENC_u0_u1_U313  ( .A1(_AES_ENC_u0_u1_n590 ), .A2(_AES_ENC_u0_u1_n753 ), .ZN(_AES_ENC_u0_u1_n1023 ) );
NAND4_X2 _AES_ENC_u0_u1_U308  ( .A1(_AES_ENC_u0_u1_n760 ), .A2(_AES_ENC_u0_u1_n992 ), .A3(_AES_ENC_u0_u1_n759 ), .A4(_AES_ENC_u0_u1_n758 ), .ZN(_AES_ENC_u0_u1_n761 ) );
NAND2_X2 _AES_ENC_u0_u1_U307  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n761 ), .ZN(_AES_ENC_u0_u1_n792 ) );
NAND2_X2 _AES_ENC_u0_u1_U306  ( .A1(_AES_ENC_u0_u1_n584 ), .A2(_AES_ENC_u0_u1_n603 ), .ZN(_AES_ENC_u0_u1_n989 ) );
NAND2_X2 _AES_ENC_u0_u1_U305  ( .A1(_AES_ENC_u0_u1_n1050 ), .A2(_AES_ENC_u0_u1_n989 ), .ZN(_AES_ENC_u0_u1_n777 ) );
NAND2_X2 _AES_ENC_u0_u1_U304  ( .A1(_AES_ENC_u0_u1_n1093 ), .A2(_AES_ENC_u0_u1_n762 ), .ZN(_AES_ENC_u0_u1_n776 ) );
XNOR2_X2 _AES_ENC_u0_u1_U301  ( .A(_AES_ENC_w3[15] ), .B(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n959 ) );
NAND4_X2 _AES_ENC_u0_u1_U289  ( .A1(_AES_ENC_u0_u1_n777 ), .A2(_AES_ENC_u0_u1_n776 ), .A3(_AES_ENC_u0_u1_n775 ), .A4(_AES_ENC_u0_u1_n774 ), .ZN(_AES_ENC_u0_u1_n778 ) );
NAND2_X2 _AES_ENC_u0_u1_U288  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n778 ), .ZN(_AES_ENC_u0_u1_n791 ) );
NAND2_X2 _AES_ENC_u0_u1_U287  ( .A1(_AES_ENC_u0_u1_n1056 ), .A2(_AES_ENC_u0_u1_n1050 ), .ZN(_AES_ENC_u0_u1_n788 ) );
NAND2_X2 _AES_ENC_u0_u1_U286  ( .A1(_AES_ENC_u0_u1_n1091 ), .A2(_AES_ENC_u0_u1_n779 ), .ZN(_AES_ENC_u0_u1_n787 ) );
NAND2_X2 _AES_ENC_u0_u1_U285  ( .A1(_AES_ENC_u0_u1_n956 ), .A2(_AES_ENC_w3[9] ), .ZN(_AES_ENC_u0_u1_n786 ) );
NAND4_X2 _AES_ENC_u0_u1_U278  ( .A1(_AES_ENC_u0_u1_n788 ), .A2(_AES_ENC_u0_u1_n787 ), .A3(_AES_ENC_u0_u1_n786 ), .A4(_AES_ENC_u0_u1_n785 ), .ZN(_AES_ENC_u0_u1_n789 ) );
NAND2_X2 _AES_ENC_u0_u1_U277  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n789 ), .ZN(_AES_ENC_u0_u1_n790 ) );
NAND4_X2 _AES_ENC_u0_u1_U276  ( .A1(_AES_ENC_u0_u1_n793 ), .A2(_AES_ENC_u0_u1_n792 ), .A3(_AES_ENC_u0_u1_n791 ), .A4(_AES_ENC_u0_u1_n790 ), .ZN(_AES_ENC_u0_subword[18] ) );
NAND2_X2 _AES_ENC_u0_u1_U275  ( .A1(_AES_ENC_u0_u1_n1059 ), .A2(_AES_ENC_u0_u1_n794 ), .ZN(_AES_ENC_u0_u1_n810 ) );
NAND2_X2 _AES_ENC_u0_u1_U274  ( .A1(_AES_ENC_u0_u1_n1049 ), .A2(_AES_ENC_u0_u1_n956 ), .ZN(_AES_ENC_u0_u1_n809 ) );
OR2_X2 _AES_ENC_u0_u1_U266  ( .A1(_AES_ENC_u0_u1_n1096 ), .A2(_AES_ENC_u0_u1_n606 ), .ZN(_AES_ENC_u0_u1_n802 ) );
NAND2_X2 _AES_ENC_u0_u1_U265  ( .A1(_AES_ENC_u0_u1_n1053 ), .A2(_AES_ENC_u0_u1_n800 ), .ZN(_AES_ENC_u0_u1_n801 ) );
NAND2_X2 _AES_ENC_u0_u1_U264  ( .A1(_AES_ENC_u0_u1_n802 ), .A2(_AES_ENC_u0_u1_n801 ), .ZN(_AES_ENC_u0_u1_n805 ) );
NAND4_X2 _AES_ENC_u0_u1_U261  ( .A1(_AES_ENC_u0_u1_n810 ), .A2(_AES_ENC_u0_u1_n809 ), .A3(_AES_ENC_u0_u1_n808 ), .A4(_AES_ENC_u0_u1_n807 ), .ZN(_AES_ENC_u0_u1_n811 ) );
NAND2_X2 _AES_ENC_u0_u1_U260  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n811 ), .ZN(_AES_ENC_u0_u1_n852 ) );
OR2_X2 _AES_ENC_u0_u1_U259  ( .A1(_AES_ENC_u0_u1_n1023 ), .A2(_AES_ENC_u0_u1_n617 ), .ZN(_AES_ENC_u0_u1_n819 ) );
OR2_X2 _AES_ENC_u0_u1_U257  ( .A1(_AES_ENC_u0_u1_n570 ), .A2(_AES_ENC_u0_u1_n930 ), .ZN(_AES_ENC_u0_u1_n818 ) );
NAND2_X2 _AES_ENC_u0_u1_U256  ( .A1(_AES_ENC_u0_u1_n1013 ), .A2(_AES_ENC_u0_u1_n1094 ), .ZN(_AES_ENC_u0_u1_n817 ) );
NAND4_X2 _AES_ENC_u0_u1_U249  ( .A1(_AES_ENC_u0_u1_n819 ), .A2(_AES_ENC_u0_u1_n818 ), .A3(_AES_ENC_u0_u1_n817 ), .A4(_AES_ENC_u0_u1_n816 ), .ZN(_AES_ENC_u0_u1_n820 ) );
NAND2_X2 _AES_ENC_u0_u1_U248  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n820 ), .ZN(_AES_ENC_u0_u1_n851 ) );
NAND2_X2 _AES_ENC_u0_u1_U247  ( .A1(_AES_ENC_u0_u1_n956 ), .A2(_AES_ENC_u0_u1_n1080 ), .ZN(_AES_ENC_u0_u1_n835 ) );
NAND2_X2 _AES_ENC_u0_u1_U246  ( .A1(_AES_ENC_u0_u1_n570 ), .A2(_AES_ENC_u0_u1_n1030 ), .ZN(_AES_ENC_u0_u1_n1047 ) );
OR2_X2 _AES_ENC_u0_u1_U245  ( .A1(_AES_ENC_u0_u1_n1047 ), .A2(_AES_ENC_u0_u1_n612 ), .ZN(_AES_ENC_u0_u1_n834 ) );
NAND2_X2 _AES_ENC_u0_u1_U244  ( .A1(_AES_ENC_u0_u1_n1072 ), .A2(_AES_ENC_u0_u1_n589 ), .ZN(_AES_ENC_u0_u1_n833 ) );
NAND4_X2 _AES_ENC_u0_u1_U233  ( .A1(_AES_ENC_u0_u1_n835 ), .A2(_AES_ENC_u0_u1_n834 ), .A3(_AES_ENC_u0_u1_n833 ), .A4(_AES_ENC_u0_u1_n832 ), .ZN(_AES_ENC_u0_u1_n836 ) );
NAND2_X2 _AES_ENC_u0_u1_U232  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n836 ), .ZN(_AES_ENC_u0_u1_n850 ) );
NAND2_X2 _AES_ENC_u0_u1_U231  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n623 ), .ZN(_AES_ENC_u0_u1_n847 ) );
NAND2_X2 _AES_ENC_u0_u1_U230  ( .A1(_AES_ENC_u0_u1_n1050 ), .A2(_AES_ENC_u0_u1_n1071 ), .ZN(_AES_ENC_u0_u1_n846 ) );
OR2_X2 _AES_ENC_u0_u1_U224  ( .A1(_AES_ENC_u0_u1_n1053 ), .A2(_AES_ENC_u0_u1_n911 ), .ZN(_AES_ENC_u0_u1_n1077 ) );
NAND4_X2 _AES_ENC_u0_u1_U220  ( .A1(_AES_ENC_u0_u1_n847 ), .A2(_AES_ENC_u0_u1_n846 ), .A3(_AES_ENC_u0_u1_n845 ), .A4(_AES_ENC_u0_u1_n844 ), .ZN(_AES_ENC_u0_u1_n848 ) );
NAND2_X2 _AES_ENC_u0_u1_U219  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n848 ), .ZN(_AES_ENC_u0_u1_n849 ) );
NAND4_X2 _AES_ENC_u0_u1_U218  ( .A1(_AES_ENC_u0_u1_n852 ), .A2(_AES_ENC_u0_u1_n851 ), .A3(_AES_ENC_u0_u1_n850 ), .A4(_AES_ENC_u0_u1_n849 ), .ZN(_AES_ENC_u0_subword[19] ) );
NAND2_X2 _AES_ENC_u0_u1_U216  ( .A1(_AES_ENC_u0_u1_n1009 ), .A2(_AES_ENC_u0_u1_n1072 ), .ZN(_AES_ENC_u0_u1_n862 ) );
NAND2_X2 _AES_ENC_u0_u1_U215  ( .A1(_AES_ENC_u0_u1_n603 ), .A2(_AES_ENC_u0_u1_n577 ), .ZN(_AES_ENC_u0_u1_n853 ) );
NAND2_X2 _AES_ENC_u0_u1_U214  ( .A1(_AES_ENC_u0_u1_n1050 ), .A2(_AES_ENC_u0_u1_n853 ), .ZN(_AES_ENC_u0_u1_n861 ) );
NAND4_X2 _AES_ENC_u0_u1_U206  ( .A1(_AES_ENC_u0_u1_n862 ), .A2(_AES_ENC_u0_u1_n861 ), .A3(_AES_ENC_u0_u1_n860 ), .A4(_AES_ENC_u0_u1_n859 ), .ZN(_AES_ENC_u0_u1_n863 ) );
NAND2_X2 _AES_ENC_u0_u1_U205  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n863 ), .ZN(_AES_ENC_u0_u1_n905 ) );
NAND2_X2 _AES_ENC_u0_u1_U204  ( .A1(_AES_ENC_u0_u1_n1010 ), .A2(_AES_ENC_u0_u1_n989 ), .ZN(_AES_ENC_u0_u1_n874 ) );
NAND2_X2 _AES_ENC_u0_u1_U203  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n610 ), .ZN(_AES_ENC_u0_u1_n864 ) );
NAND2_X2 _AES_ENC_u0_u1_U202  ( .A1(_AES_ENC_u0_u1_n929 ), .A2(_AES_ENC_u0_u1_n864 ), .ZN(_AES_ENC_u0_u1_n873 ) );
NAND4_X2 _AES_ENC_u0_u1_U193  ( .A1(_AES_ENC_u0_u1_n874 ), .A2(_AES_ENC_u0_u1_n873 ), .A3(_AES_ENC_u0_u1_n872 ), .A4(_AES_ENC_u0_u1_n871 ), .ZN(_AES_ENC_u0_u1_n875 ) );
NAND2_X2 _AES_ENC_u0_u1_U192  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n875 ), .ZN(_AES_ENC_u0_u1_n904 ) );
NAND2_X2 _AES_ENC_u0_u1_U191  ( .A1(_AES_ENC_u0_u1_n583 ), .A2(_AES_ENC_u0_u1_n1050 ), .ZN(_AES_ENC_u0_u1_n889 ) );
NAND2_X2 _AES_ENC_u0_u1_U190  ( .A1(_AES_ENC_u0_u1_n1093 ), .A2(_AES_ENC_u0_u1_n587 ), .ZN(_AES_ENC_u0_u1_n876 ) );
NAND2_X2 _AES_ENC_u0_u1_U189  ( .A1(_AES_ENC_u0_u1_n604 ), .A2(_AES_ENC_u0_u1_n876 ), .ZN(_AES_ENC_u0_u1_n877 ) );
NAND2_X2 _AES_ENC_u0_u1_U188  ( .A1(_AES_ENC_u0_u1_n877 ), .A2(_AES_ENC_u0_u1_n623 ), .ZN(_AES_ENC_u0_u1_n888 ) );
NAND4_X2 _AES_ENC_u0_u1_U179  ( .A1(_AES_ENC_u0_u1_n889 ), .A2(_AES_ENC_u0_u1_n888 ), .A3(_AES_ENC_u0_u1_n887 ), .A4(_AES_ENC_u0_u1_n886 ), .ZN(_AES_ENC_u0_u1_n890 ) );
NAND2_X2 _AES_ENC_u0_u1_U178  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n890 ), .ZN(_AES_ENC_u0_u1_n903 ) );
OR2_X2 _AES_ENC_u0_u1_U177  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n1059 ), .ZN(_AES_ENC_u0_u1_n900 ) );
NAND2_X2 _AES_ENC_u0_u1_U176  ( .A1(_AES_ENC_u0_u1_n1073 ), .A2(_AES_ENC_u0_u1_n1047 ), .ZN(_AES_ENC_u0_u1_n899 ) );
NAND2_X2 _AES_ENC_u0_u1_U175  ( .A1(_AES_ENC_u0_u1_n1094 ), .A2(_AES_ENC_u0_u1_n595 ), .ZN(_AES_ENC_u0_u1_n898 ) );
NAND4_X2 _AES_ENC_u0_u1_U167  ( .A1(_AES_ENC_u0_u1_n900 ), .A2(_AES_ENC_u0_u1_n899 ), .A3(_AES_ENC_u0_u1_n898 ), .A4(_AES_ENC_u0_u1_n897 ), .ZN(_AES_ENC_u0_u1_n901 ) );
NAND2_X2 _AES_ENC_u0_u1_U166  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n901 ), .ZN(_AES_ENC_u0_u1_n902 ) );
NAND4_X2 _AES_ENC_u0_u1_U165  ( .A1(_AES_ENC_u0_u1_n905 ), .A2(_AES_ENC_u0_u1_n904 ), .A3(_AES_ENC_u0_u1_n903 ), .A4(_AES_ENC_u0_u1_n902 ), .ZN(_AES_ENC_u0_subword[20] ) );
NAND2_X2 _AES_ENC_u0_u1_U164  ( .A1(_AES_ENC_u0_u1_n1094 ), .A2(_AES_ENC_u0_u1_n599 ), .ZN(_AES_ENC_u0_u1_n922 ) );
NAND2_X2 _AES_ENC_u0_u1_U163  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n989 ), .ZN(_AES_ENC_u0_u1_n921 ) );
NAND4_X2 _AES_ENC_u0_u1_U151  ( .A1(_AES_ENC_u0_u1_n922 ), .A2(_AES_ENC_u0_u1_n921 ), .A3(_AES_ENC_u0_u1_n920 ), .A4(_AES_ENC_u0_u1_n919 ), .ZN(_AES_ENC_u0_u1_n923 ) );
NAND2_X2 _AES_ENC_u0_u1_U150  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n923 ), .ZN(_AES_ENC_u0_u1_n972 ) );
NAND2_X2 _AES_ENC_u0_u1_U149  ( .A1(_AES_ENC_u0_u1_n582 ), .A2(_AES_ENC_u0_u1_n619 ), .ZN(_AES_ENC_u0_u1_n924 ) );
NAND2_X2 _AES_ENC_u0_u1_U148  ( .A1(_AES_ENC_u0_u1_n1073 ), .A2(_AES_ENC_u0_u1_n924 ), .ZN(_AES_ENC_u0_u1_n939 ) );
NAND2_X2 _AES_ENC_u0_u1_U147  ( .A1(_AES_ENC_u0_u1_n926 ), .A2(_AES_ENC_u0_u1_n925 ), .ZN(_AES_ENC_u0_u1_n927 ) );
NAND2_X2 _AES_ENC_u0_u1_U146  ( .A1(_AES_ENC_u0_u1_n606 ), .A2(_AES_ENC_u0_u1_n927 ), .ZN(_AES_ENC_u0_u1_n928 ) );
NAND2_X2 _AES_ENC_u0_u1_U145  ( .A1(_AES_ENC_u0_u1_n928 ), .A2(_AES_ENC_u0_u1_n1080 ), .ZN(_AES_ENC_u0_u1_n938 ) );
OR2_X2 _AES_ENC_u0_u1_U144  ( .A1(_AES_ENC_u0_u1_n1117 ), .A2(_AES_ENC_u0_u1_n615 ), .ZN(_AES_ENC_u0_u1_n937 ) );
NAND4_X2 _AES_ENC_u0_u1_U139  ( .A1(_AES_ENC_u0_u1_n939 ), .A2(_AES_ENC_u0_u1_n938 ), .A3(_AES_ENC_u0_u1_n937 ), .A4(_AES_ENC_u0_u1_n936 ), .ZN(_AES_ENC_u0_u1_n940 ) );
NAND2_X2 _AES_ENC_u0_u1_U138  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n940 ), .ZN(_AES_ENC_u0_u1_n971 ) );
OR2_X2 _AES_ENC_u0_u1_U137  ( .A1(_AES_ENC_u0_u1_n605 ), .A2(_AES_ENC_u0_u1_n941 ), .ZN(_AES_ENC_u0_u1_n954 ) );
NAND2_X2 _AES_ENC_u0_u1_U136  ( .A1(_AES_ENC_u0_u1_n1096 ), .A2(_AES_ENC_u0_u1_n577 ), .ZN(_AES_ENC_u0_u1_n942 ) );
NAND2_X2 _AES_ENC_u0_u1_U135  ( .A1(_AES_ENC_u0_u1_n1048 ), .A2(_AES_ENC_u0_u1_n942 ), .ZN(_AES_ENC_u0_u1_n943 ) );
NAND2_X2 _AES_ENC_u0_u1_U134  ( .A1(_AES_ENC_u0_u1_n612 ), .A2(_AES_ENC_u0_u1_n943 ), .ZN(_AES_ENC_u0_u1_n944 ) );
NAND2_X2 _AES_ENC_u0_u1_U133  ( .A1(_AES_ENC_u0_u1_n944 ), .A2(_AES_ENC_u0_u1_n580 ), .ZN(_AES_ENC_u0_u1_n953 ) );
NAND4_X2 _AES_ENC_u0_u1_U125  ( .A1(_AES_ENC_u0_u1_n954 ), .A2(_AES_ENC_u0_u1_n953 ), .A3(_AES_ENC_u0_u1_n952 ), .A4(_AES_ENC_u0_u1_n951 ), .ZN(_AES_ENC_u0_u1_n955 ) );
NAND2_X2 _AES_ENC_u0_u1_U124  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n955 ), .ZN(_AES_ENC_u0_u1_n970 ) );
NAND2_X2 _AES_ENC_u0_u1_U123  ( .A1(_AES_ENC_u0_u1_n1094 ), .A2(_AES_ENC_u0_u1_n1071 ), .ZN(_AES_ENC_u0_u1_n967 ) );
NAND2_X2 _AES_ENC_u0_u1_U122  ( .A1(_AES_ENC_u0_u1_n956 ), .A2(_AES_ENC_u0_u1_n1030 ), .ZN(_AES_ENC_u0_u1_n966 ) );
NAND4_X2 _AES_ENC_u0_u1_U114  ( .A1(_AES_ENC_u0_u1_n967 ), .A2(_AES_ENC_u0_u1_n966 ), .A3(_AES_ENC_u0_u1_n965 ), .A4(_AES_ENC_u0_u1_n964 ), .ZN(_AES_ENC_u0_u1_n968 ) );
NAND2_X2 _AES_ENC_u0_u1_U113  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n968 ), .ZN(_AES_ENC_u0_u1_n969 ) );
NAND4_X2 _AES_ENC_u0_u1_U112  ( .A1(_AES_ENC_u0_u1_n972 ), .A2(_AES_ENC_u0_u1_n971 ), .A3(_AES_ENC_u0_u1_n970 ), .A4(_AES_ENC_u0_u1_n969 ), .ZN(_AES_ENC_u0_subword[21] ) );
NAND2_X2 _AES_ENC_u0_u1_U111  ( .A1(_AES_ENC_u0_u1_n570 ), .A2(_AES_ENC_u0_u1_n1097 ), .ZN(_AES_ENC_u0_u1_n973 ) );
NAND2_X2 _AES_ENC_u0_u1_U110  ( .A1(_AES_ENC_u0_u1_n1073 ), .A2(_AES_ENC_u0_u1_n973 ), .ZN(_AES_ENC_u0_u1_n987 ) );
NAND2_X2 _AES_ENC_u0_u1_U109  ( .A1(_AES_ENC_u0_u1_n974 ), .A2(_AES_ENC_u0_u1_n1077 ), .ZN(_AES_ENC_u0_u1_n975 ) );
NAND2_X2 _AES_ENC_u0_u1_U108  ( .A1(_AES_ENC_u0_u1_n613 ), .A2(_AES_ENC_u0_u1_n975 ), .ZN(_AES_ENC_u0_u1_n976 ) );
NAND2_X2 _AES_ENC_u0_u1_U107  ( .A1(_AES_ENC_u0_u1_n977 ), .A2(_AES_ENC_u0_u1_n976 ), .ZN(_AES_ENC_u0_u1_n986 ) );
NAND4_X2 _AES_ENC_u0_u1_U99  ( .A1(_AES_ENC_u0_u1_n987 ), .A2(_AES_ENC_u0_u1_n986 ), .A3(_AES_ENC_u0_u1_n985 ), .A4(_AES_ENC_u0_u1_n984 ), .ZN(_AES_ENC_u0_u1_n988 ) );
NAND2_X2 _AES_ENC_u0_u1_U98  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n988 ), .ZN(_AES_ENC_u0_u1_n1044 ) );
NAND2_X2 _AES_ENC_u0_u1_U97  ( .A1(_AES_ENC_u0_u1_n1073 ), .A2(_AES_ENC_u0_u1_n989 ), .ZN(_AES_ENC_u0_u1_n1004 ) );
NAND2_X2 _AES_ENC_u0_u1_U96  ( .A1(_AES_ENC_u0_u1_n1092 ), .A2(_AES_ENC_u0_u1_n619 ), .ZN(_AES_ENC_u0_u1_n1003 ) );
NAND4_X2 _AES_ENC_u0_u1_U85  ( .A1(_AES_ENC_u0_u1_n1004 ), .A2(_AES_ENC_u0_u1_n1003 ), .A3(_AES_ENC_u0_u1_n1002 ), .A4(_AES_ENC_u0_u1_n1001 ), .ZN(_AES_ENC_u0_u1_n1005 ) );
NAND2_X2 _AES_ENC_u0_u1_U84  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n1005 ), .ZN(_AES_ENC_u0_u1_n1043 ) );
NAND2_X2 _AES_ENC_u0_u1_U83  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n596 ), .ZN(_AES_ENC_u0_u1_n1020 ) );
NAND2_X2 _AES_ENC_u0_u1_U82  ( .A1(_AES_ENC_u0_u1_n1050 ), .A2(_AES_ENC_u0_u1_n624 ), .ZN(_AES_ENC_u0_u1_n1019 ) );
NAND2_X2 _AES_ENC_u0_u1_U77  ( .A1(_AES_ENC_u0_u1_n1059 ), .A2(_AES_ENC_u0_u1_n1114 ), .ZN(_AES_ENC_u0_u1_n1012 ) );
NAND2_X2 _AES_ENC_u0_u1_U76  ( .A1(_AES_ENC_u0_u1_n1010 ), .A2(_AES_ENC_u0_u1_n592 ), .ZN(_AES_ENC_u0_u1_n1011 ) );
NAND2_X2 _AES_ENC_u0_u1_U75  ( .A1(_AES_ENC_u0_u1_n1012 ), .A2(_AES_ENC_u0_u1_n1011 ), .ZN(_AES_ENC_u0_u1_n1016 ) );
NAND4_X2 _AES_ENC_u0_u1_U70  ( .A1(_AES_ENC_u0_u1_n1020 ), .A2(_AES_ENC_u0_u1_n1019 ), .A3(_AES_ENC_u0_u1_n1018 ), .A4(_AES_ENC_u0_u1_n1017 ), .ZN(_AES_ENC_u0_u1_n1021 ) );
NAND2_X2 _AES_ENC_u0_u1_U69  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n1021 ), .ZN(_AES_ENC_u0_u1_n1042 ) );
NAND2_X2 _AES_ENC_u0_u1_U68  ( .A1(_AES_ENC_u0_u1_n1022 ), .A2(_AES_ENC_u0_u1_n1093 ), .ZN(_AES_ENC_u0_u1_n1039 ) );
NAND2_X2 _AES_ENC_u0_u1_U67  ( .A1(_AES_ENC_u0_u1_n1050 ), .A2(_AES_ENC_u0_u1_n1023 ), .ZN(_AES_ENC_u0_u1_n1038 ) );
NAND2_X2 _AES_ENC_u0_u1_U66  ( .A1(_AES_ENC_u0_u1_n1024 ), .A2(_AES_ENC_u0_u1_n1071 ), .ZN(_AES_ENC_u0_u1_n1037 ) );
AND2_X2 _AES_ENC_u0_u1_U60  ( .A1(_AES_ENC_u0_u1_n1030 ), .A2(_AES_ENC_u0_u1_n602 ), .ZN(_AES_ENC_u0_u1_n1078 ) );
NAND4_X2 _AES_ENC_u0_u1_U56  ( .A1(_AES_ENC_u0_u1_n1039 ), .A2(_AES_ENC_u0_u1_n1038 ), .A3(_AES_ENC_u0_u1_n1037 ), .A4(_AES_ENC_u0_u1_n1036 ), .ZN(_AES_ENC_u0_u1_n1040 ) );
NAND2_X2 _AES_ENC_u0_u1_U55  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n1040 ), .ZN(_AES_ENC_u0_u1_n1041 ) );
NAND4_X2 _AES_ENC_u0_u1_U54  ( .A1(_AES_ENC_u0_u1_n1044 ), .A2(_AES_ENC_u0_u1_n1043 ), .A3(_AES_ENC_u0_u1_n1042 ), .A4(_AES_ENC_u0_u1_n1041 ), .ZN(_AES_ENC_u0_subword[22] ) );
NAND2_X2 _AES_ENC_u0_u1_U53  ( .A1(_AES_ENC_u0_u1_n1072 ), .A2(_AES_ENC_u0_u1_n1045 ), .ZN(_AES_ENC_u0_u1_n1068 ) );
NAND2_X2 _AES_ENC_u0_u1_U52  ( .A1(_AES_ENC_u0_u1_n1046 ), .A2(_AES_ENC_u0_u1_n582 ), .ZN(_AES_ENC_u0_u1_n1067 ) );
NAND2_X2 _AES_ENC_u0_u1_U51  ( .A1(_AES_ENC_u0_u1_n1094 ), .A2(_AES_ENC_u0_u1_n1047 ), .ZN(_AES_ENC_u0_u1_n1066 ) );
NAND4_X2 _AES_ENC_u0_u1_U40  ( .A1(_AES_ENC_u0_u1_n1068 ), .A2(_AES_ENC_u0_u1_n1067 ), .A3(_AES_ENC_u0_u1_n1066 ), .A4(_AES_ENC_u0_u1_n1065 ), .ZN(_AES_ENC_u0_u1_n1069 ) );
NAND2_X2 _AES_ENC_u0_u1_U39  ( .A1(_AES_ENC_u0_u1_n1070 ), .A2(_AES_ENC_u0_u1_n1069 ), .ZN(_AES_ENC_u0_u1_n1135 ) );
NAND2_X2 _AES_ENC_u0_u1_U38  ( .A1(_AES_ENC_u0_u1_n1072 ), .A2(_AES_ENC_u0_u1_n1071 ), .ZN(_AES_ENC_u0_u1_n1088 ) );
NAND2_X2 _AES_ENC_u0_u1_U37  ( .A1(_AES_ENC_u0_u1_n1073 ), .A2(_AES_ENC_u0_u1_n595 ), .ZN(_AES_ENC_u0_u1_n1087 ) );
NAND4_X2 _AES_ENC_u0_u1_U28  ( .A1(_AES_ENC_u0_u1_n1088 ), .A2(_AES_ENC_u0_u1_n1087 ), .A3(_AES_ENC_u0_u1_n1086 ), .A4(_AES_ENC_u0_u1_n1085 ), .ZN(_AES_ENC_u0_u1_n1089 ) );
NAND2_X2 _AES_ENC_u0_u1_U27  ( .A1(_AES_ENC_u0_u1_n1090 ), .A2(_AES_ENC_u0_u1_n1089 ), .ZN(_AES_ENC_u0_u1_n1134 ) );
NAND2_X2 _AES_ENC_u0_u1_U26  ( .A1(_AES_ENC_u0_u1_n1091 ), .A2(_AES_ENC_u0_u1_n1093 ), .ZN(_AES_ENC_u0_u1_n1111 ) );
NAND2_X2 _AES_ENC_u0_u1_U25  ( .A1(_AES_ENC_u0_u1_n1092 ), .A2(_AES_ENC_u0_u1_n1120 ), .ZN(_AES_ENC_u0_u1_n1110 ) );
AND2_X2 _AES_ENC_u0_u1_U22  ( .A1(_AES_ENC_u0_u1_n1097 ), .A2(_AES_ENC_u0_u1_n1096 ), .ZN(_AES_ENC_u0_u1_n1098 ) );
NAND4_X2 _AES_ENC_u0_u1_U14  ( .A1(_AES_ENC_u0_u1_n1111 ), .A2(_AES_ENC_u0_u1_n1110 ), .A3(_AES_ENC_u0_u1_n1109 ), .A4(_AES_ENC_u0_u1_n1108 ), .ZN(_AES_ENC_u0_u1_n1112 ) );
NAND2_X2 _AES_ENC_u0_u1_U13  ( .A1(_AES_ENC_u0_u1_n1113 ), .A2(_AES_ENC_u0_u1_n1112 ), .ZN(_AES_ENC_u0_u1_n1133 ) );
NAND2_X2 _AES_ENC_u0_u1_U12  ( .A1(_AES_ENC_u0_u1_n1115 ), .A2(_AES_ENC_u0_u1_n1114 ), .ZN(_AES_ENC_u0_u1_n1129 ) );
OR2_X2 _AES_ENC_u0_u1_U11  ( .A1(_AES_ENC_u0_u1_n608 ), .A2(_AES_ENC_u0_u1_n1116 ), .ZN(_AES_ENC_u0_u1_n1128 ) );
NAND4_X2 _AES_ENC_u0_u1_U3  ( .A1(_AES_ENC_u0_u1_n1129 ), .A2(_AES_ENC_u0_u1_n1128 ), .A3(_AES_ENC_u0_u1_n1127 ), .A4(_AES_ENC_u0_u1_n1126 ), .ZN(_AES_ENC_u0_u1_n1130 ) );
NAND2_X2 _AES_ENC_u0_u1_U2  ( .A1(_AES_ENC_u0_u1_n1131 ), .A2(_AES_ENC_u0_u1_n1130 ), .ZN(_AES_ENC_u0_u1_n1132 ) );
NAND4_X2 _AES_ENC_u0_u1_U1  ( .A1(_AES_ENC_u0_u1_n1135 ), .A2(_AES_ENC_u0_u1_n1134 ), .A3(_AES_ENC_u0_u1_n1133 ), .A4(_AES_ENC_u0_u1_n1132 ), .ZN(_AES_ENC_u0_subword[23] ) );
INV_X4 _AES_ENC_u0_u2_U575  ( .A(_AES_ENC_w3[7] ), .ZN(_AES_ENC_u0_u2_n627 ));
INV_X4 _AES_ENC_u0_u2_U574  ( .A(_AES_ENC_u0_u2_n1114 ), .ZN(_AES_ENC_u0_u2_n625 ) );
INV_X4 _AES_ENC_u0_u2_U573  ( .A(_AES_ENC_w3[4] ), .ZN(_AES_ENC_u0_u2_n624 ));
INV_X4 _AES_ENC_u0_u2_U572  ( .A(_AES_ENC_u0_u2_n1025 ), .ZN(_AES_ENC_u0_u2_n622 ) );
INV_X4 _AES_ENC_u0_u2_U571  ( .A(_AES_ENC_u0_u2_n1120 ), .ZN(_AES_ENC_u0_u2_n620 ) );
INV_X4 _AES_ENC_u0_u2_U570  ( .A(_AES_ENC_u0_u2_n1121 ), .ZN(_AES_ENC_u0_u2_n619 ) );
INV_X4 _AES_ENC_u0_u2_U569  ( .A(_AES_ENC_u0_u2_n1048 ), .ZN(_AES_ENC_u0_u2_n618 ) );
INV_X4 _AES_ENC_u0_u2_U568  ( .A(_AES_ENC_u0_u2_n974 ), .ZN(_AES_ENC_u0_u2_n616 ) );
INV_X4 _AES_ENC_u0_u2_U567  ( .A(_AES_ENC_u0_u2_n794 ), .ZN(_AES_ENC_u0_u2_n614 ) );
INV_X4 _AES_ENC_u0_u2_U566  ( .A(_AES_ENC_w3[2] ), .ZN(_AES_ENC_u0_u2_n611 ));
INV_X4 _AES_ENC_u0_u2_U565  ( .A(_AES_ENC_u0_u2_n800 ), .ZN(_AES_ENC_u0_u2_n610 ) );
INV_X4 _AES_ENC_u0_u2_U564  ( .A(_AES_ENC_u0_u2_n925 ), .ZN(_AES_ENC_u0_u2_n609 ) );
INV_X4 _AES_ENC_u0_u2_U563  ( .A(_AES_ENC_u0_u2_n779 ), .ZN(_AES_ENC_u0_u2_n607 ) );
INV_X4 _AES_ENC_u0_u2_U562  ( .A(_AES_ENC_u0_u2_n1022 ), .ZN(_AES_ENC_u0_u2_n603 ) );
INV_X4 _AES_ENC_u0_u2_U561  ( .A(_AES_ENC_u0_u2_n1102 ), .ZN(_AES_ENC_u0_u2_n602 ) );
INV_X4 _AES_ENC_u0_u2_U560  ( .A(_AES_ENC_u0_u2_n929 ), .ZN(_AES_ENC_u0_u2_n601 ) );
INV_X4 _AES_ENC_u0_u2_U559  ( .A(_AES_ENC_u0_u2_n1056 ), .ZN(_AES_ENC_u0_u2_n600 ) );
INV_X4 _AES_ENC_u0_u2_U558  ( .A(_AES_ENC_u0_u2_n1054 ), .ZN(_AES_ENC_u0_u2_n599 ) );
INV_X4 _AES_ENC_u0_u2_U557  ( .A(_AES_ENC_u0_u2_n881 ), .ZN(_AES_ENC_u0_u2_n598 ) );
INV_X4 _AES_ENC_u0_u2_U556  ( .A(_AES_ENC_u0_u2_n926 ), .ZN(_AES_ENC_u0_u2_n597 ) );
INV_X4 _AES_ENC_u0_u2_U555  ( .A(_AES_ENC_u0_u2_n977 ), .ZN(_AES_ENC_u0_u2_n595 ) );
INV_X4 _AES_ENC_u0_u2_U554  ( .A(_AES_ENC_u0_u2_n1031 ), .ZN(_AES_ENC_u0_u2_n594 ) );
INV_X4 _AES_ENC_u0_u2_U553  ( .A(_AES_ENC_u0_u2_n1103 ), .ZN(_AES_ENC_u0_u2_n593 ) );
INV_X4 _AES_ENC_u0_u2_U552  ( .A(_AES_ENC_u0_u2_n1009 ), .ZN(_AES_ENC_u0_u2_n592 ) );
INV_X4 _AES_ENC_u0_u2_U551  ( .A(_AES_ENC_u0_u2_n990 ), .ZN(_AES_ENC_u0_u2_n591 ) );
INV_X4 _AES_ENC_u0_u2_U550  ( .A(_AES_ENC_u0_u2_n1058 ), .ZN(_AES_ENC_u0_u2_n590 ) );
INV_X4 _AES_ENC_u0_u2_U549  ( .A(_AES_ENC_u0_u2_n1074 ), .ZN(_AES_ENC_u0_u2_n589 ) );
INV_X4 _AES_ENC_u0_u2_U548  ( .A(_AES_ENC_u0_u2_n1053 ), .ZN(_AES_ENC_u0_u2_n588 ) );
INV_X4 _AES_ENC_u0_u2_U547  ( .A(_AES_ENC_u0_u2_n826 ), .ZN(_AES_ENC_u0_u2_n587 ) );
INV_X4 _AES_ENC_u0_u2_U546  ( .A(_AES_ENC_u0_u2_n992 ), .ZN(_AES_ENC_u0_u2_n586 ) );
INV_X4 _AES_ENC_u0_u2_U545  ( .A(_AES_ENC_u0_u2_n821 ), .ZN(_AES_ENC_u0_u2_n585 ) );
INV_X4 _AES_ENC_u0_u2_U544  ( .A(_AES_ENC_u0_u2_n910 ), .ZN(_AES_ENC_u0_u2_n584 ) );
INV_X4 _AES_ENC_u0_u2_U543  ( .A(_AES_ENC_u0_u2_n906 ), .ZN(_AES_ENC_u0_u2_n583 ) );
INV_X4 _AES_ENC_u0_u2_U542  ( .A(_AES_ENC_u0_u2_n880 ), .ZN(_AES_ENC_u0_u2_n581 ) );
INV_X4 _AES_ENC_u0_u2_U541  ( .A(_AES_ENC_u0_u2_n1013 ), .ZN(_AES_ENC_u0_u2_n580 ) );
INV_X4 _AES_ENC_u0_u2_U540  ( .A(_AES_ENC_u0_u2_n1092 ), .ZN(_AES_ENC_u0_u2_n579 ) );
INV_X4 _AES_ENC_u0_u2_U539  ( .A(_AES_ENC_u0_u2_n824 ), .ZN(_AES_ENC_u0_u2_n578 ) );
INV_X4 _AES_ENC_u0_u2_U538  ( .A(_AES_ENC_u0_u2_n1091 ), .ZN(_AES_ENC_u0_u2_n577 ) );
INV_X4 _AES_ENC_u0_u2_U537  ( .A(_AES_ENC_u0_u2_n1080 ), .ZN(_AES_ENC_u0_u2_n576 ) );
INV_X4 _AES_ENC_u0_u2_U536  ( .A(_AES_ENC_u0_u2_n959 ), .ZN(_AES_ENC_u0_u2_n575 ) );
INV_X4 _AES_ENC_u0_u2_U535  ( .A(_AES_ENC_w3[0] ), .ZN(_AES_ENC_u0_u2_n574 ));
NOR2_X2 _AES_ENC_u0_u2_U534  ( .A1(_AES_ENC_u0_u2_n574 ), .A2(_AES_ENC_w3[6] ), .ZN(_AES_ENC_u0_u2_n1070 ) );
NOR2_X2 _AES_ENC_u0_u2_U533  ( .A1(_AES_ENC_w3[0] ), .A2(_AES_ENC_w3[6] ),.ZN(_AES_ENC_u0_u2_n1090 ) );
NOR2_X2 _AES_ENC_u0_u2_U532  ( .A1(_AES_ENC_w3[4] ), .A2(_AES_ENC_w3[3] ),.ZN(_AES_ENC_u0_u2_n1025 ) );
NAND3_X2 _AES_ENC_u0_u2_U531  ( .A1(_AES_ENC_u0_u2_n679 ), .A2(_AES_ENC_u0_u2_n678 ), .A3(_AES_ENC_u0_u2_n677 ), .ZN(_AES_ENC_u0_subword[8] ) );
NOR2_X2 _AES_ENC_u0_u2_U530  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n765 ) );
NOR2_X2 _AES_ENC_u0_u2_U529  ( .A1(_AES_ENC_w3[4] ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n764 ) );
NOR2_X2 _AES_ENC_u0_u2_U528  ( .A1(_AES_ENC_u0_u2_n765 ), .A2(_AES_ENC_u0_u2_n764 ), .ZN(_AES_ENC_u0_u2_n766 ) );
NOR2_X2 _AES_ENC_u0_u2_U527  ( .A1(_AES_ENC_u0_u2_n766 ), .A2(_AES_ENC_u0_u2_n575 ), .ZN(_AES_ENC_u0_u2_n767 ) );
NOR2_X2 _AES_ENC_u0_u2_U526  ( .A1(_AES_ENC_u0_u2_n1117 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n707 ) );
NOR3_X2 _AES_ENC_u0_u2_U525  ( .A1(_AES_ENC_u0_u2_n627 ), .A2(_AES_ENC_w3[5] ), .A3(_AES_ENC_u0_u2_n704 ), .ZN(_AES_ENC_u0_u2_n706 ));
NOR2_X2 _AES_ENC_u0_u2_U524  ( .A1(_AES_ENC_w3[4] ), .A2(_AES_ENC_u0_u2_n579 ), .ZN(_AES_ENC_u0_u2_n705 ) );
NOR3_X2 _AES_ENC_u0_u2_U523  ( .A1(_AES_ENC_u0_u2_n707 ), .A2(_AES_ENC_u0_u2_n706 ), .A3(_AES_ENC_u0_u2_n705 ), .ZN(_AES_ENC_u0_u2_n713 ) );
NOR4_X2 _AES_ENC_u0_u2_U522  ( .A1(_AES_ENC_u0_u2_n633 ), .A2(_AES_ENC_u0_u2_n632 ), .A3(_AES_ENC_u0_u2_n631 ), .A4(_AES_ENC_u0_u2_n630 ), .ZN(_AES_ENC_u0_u2_n634 ) );
NOR2_X2 _AES_ENC_u0_u2_U521  ( .A1(_AES_ENC_u0_u2_n629 ), .A2(_AES_ENC_u0_u2_n628 ), .ZN(_AES_ENC_u0_u2_n635 ) );
NAND3_X2 _AES_ENC_u0_u2_U520  ( .A1(_AES_ENC_w3[2] ), .A2(_AES_ENC_w3[7] ),.A3(_AES_ENC_u0_u2_n1059 ), .ZN(_AES_ENC_u0_u2_n636 ) );
INV_X4 _AES_ENC_u0_u2_U519  ( .A(_AES_ENC_w3[3] ), .ZN(_AES_ENC_u0_u2_n621 ));
NOR2_X2 _AES_ENC_u0_u2_U518  ( .A1(_AES_ENC_w3[5] ), .A2(_AES_ENC_w3[2] ),.ZN(_AES_ENC_u0_u2_n974 ) );
NAND3_X2 _AES_ENC_u0_u2_U517  ( .A1(_AES_ENC_u0_u2_n652 ), .A2(_AES_ENC_u0_u2_n626 ), .A3(_AES_ENC_w3[7] ), .ZN(_AES_ENC_u0_u2_n653 ));
NOR2_X2 _AES_ENC_u0_u2_U516  ( .A1(_AES_ENC_u0_u2_n611 ), .A2(_AES_ENC_w3[5] ), .ZN(_AES_ENC_u0_u2_n925 ) );
NOR2_X2 _AES_ENC_u0_u2_U515  ( .A1(_AES_ENC_u0_u2_n626 ), .A2(_AES_ENC_w3[2] ), .ZN(_AES_ENC_u0_u2_n1048 ) );
INV_X4 _AES_ENC_u0_u2_U512  ( .A(_AES_ENC_w3[5] ), .ZN(_AES_ENC_u0_u2_n626 ));
NOR2_X2 _AES_ENC_u0_u2_U510  ( .A1(_AES_ENC_u0_u2_n611 ), .A2(_AES_ENC_w3[7] ), .ZN(_AES_ENC_u0_u2_n779 ) );
NOR2_X2 _AES_ENC_u0_u2_U509  ( .A1(_AES_ENC_w3[7] ), .A2(_AES_ENC_w3[2] ),.ZN(_AES_ENC_u0_u2_n794 ) );
NOR2_X2 _AES_ENC_u0_u2_U508  ( .A1(_AES_ENC_w3[4] ), .A2(_AES_ENC_w3[1] ),.ZN(_AES_ENC_u0_u2_n1102 ) );
INV_X4 _AES_ENC_u0_u2_U507  ( .A(_AES_ENC_u0_u2_n569 ), .ZN(_AES_ENC_u0_u2_n572 ) );
NOR2_X2 _AES_ENC_u0_u2_U506  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_w3[3] ), .ZN(_AES_ENC_u0_u2_n1053 ) );
NOR2_X2 _AES_ENC_u0_u2_U505  ( .A1(_AES_ENC_u0_u2_n607 ), .A2(_AES_ENC_w3[5] ), .ZN(_AES_ENC_u0_u2_n1024 ) );
NOR2_X2 _AES_ENC_u0_u2_U504  ( .A1(_AES_ENC_u0_u2_n625 ), .A2(_AES_ENC_w3[2] ), .ZN(_AES_ENC_u0_u2_n1093 ) );
NOR2_X2 _AES_ENC_u0_u2_U503  ( .A1(_AES_ENC_u0_u2_n614 ), .A2(_AES_ENC_w3[5] ), .ZN(_AES_ENC_u0_u2_n1094 ) );
NOR2_X2 _AES_ENC_u0_u2_U502  ( .A1(_AES_ENC_u0_u2_n624 ), .A2(_AES_ENC_w3[3] ), .ZN(_AES_ENC_u0_u2_n931 ) );
INV_X4 _AES_ENC_u0_u2_U501  ( .A(_AES_ENC_u0_u2_n570 ), .ZN(_AES_ENC_u0_u2_n573 ) );
NOR2_X2 _AES_ENC_u0_u2_U500  ( .A1(_AES_ENC_u0_u2_n622 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n1059 ) );
NOR2_X2 _AES_ENC_u0_u2_U499  ( .A1(_AES_ENC_u0_u2_n1053 ), .A2(_AES_ENC_u0_u2_n1095 ), .ZN(_AES_ENC_u0_u2_n639 ) );
NOR3_X2 _AES_ENC_u0_u2_U498  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n573 ), .A3(_AES_ENC_u0_u2_n1074 ), .ZN(_AES_ENC_u0_u2_n641 ) );
NOR2_X2 _AES_ENC_u0_u2_U497  ( .A1(_AES_ENC_u0_u2_n639 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n640 ) );
NOR2_X2 _AES_ENC_u0_u2_U496  ( .A1(_AES_ENC_u0_u2_n641 ), .A2(_AES_ENC_u0_u2_n640 ), .ZN(_AES_ENC_u0_u2_n646 ) );
NOR2_X2 _AES_ENC_u0_u2_U495  ( .A1(_AES_ENC_u0_u2_n826 ), .A2(_AES_ENC_u0_u2_n572 ), .ZN(_AES_ENC_u0_u2_n827 ) );
NOR3_X2 _AES_ENC_u0_u2_U494  ( .A1(_AES_ENC_u0_u2_n769 ), .A2(_AES_ENC_u0_u2_n768 ), .A3(_AES_ENC_u0_u2_n767 ), .ZN(_AES_ENC_u0_u2_n775 ) );
NOR2_X2 _AES_ENC_u0_u2_U492  ( .A1(_AES_ENC_w3[1] ), .A2(_AES_ENC_u0_u2_n623 ), .ZN(_AES_ENC_u0_u2_n913 ) );
NOR2_X2 _AES_ENC_u0_u2_U491  ( .A1(_AES_ENC_u0_u2_n913 ), .A2(_AES_ENC_u0_u2_n1091 ), .ZN(_AES_ENC_u0_u2_n914 ) );
NOR2_X2 _AES_ENC_u0_u2_U490  ( .A1(_AES_ENC_u0_u2_n1056 ), .A2(_AES_ENC_u0_u2_n1053 ), .ZN(_AES_ENC_u0_u2_n749 ) );
NOR2_X2 _AES_ENC_u0_u2_U489  ( .A1(_AES_ENC_u0_u2_n749 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n752 ) );
NOR3_X2 _AES_ENC_u0_u2_U488  ( .A1(_AES_ENC_u0_u2_n995 ), .A2(_AES_ENC_u0_u2_n586 ), .A3(_AES_ENC_u0_u2_n994 ), .ZN(_AES_ENC_u0_u2_n1002 ) );
NOR2_X2 _AES_ENC_u0_u2_U487  ( .A1(_AES_ENC_u0_u2_n909 ), .A2(_AES_ENC_u0_u2_n908 ), .ZN(_AES_ENC_u0_u2_n920 ) );
INV_X4 _AES_ENC_u0_u2_U486  ( .A(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n596 ));
NOR2_X2 _AES_ENC_u0_u2_U483  ( .A1(_AES_ENC_u0_u2_n932 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n933 ) );
NOR2_X2 _AES_ENC_u0_u2_U482  ( .A1(_AES_ENC_u0_u2_n929 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n935 ) );
NOR2_X2 _AES_ENC_u0_u2_U480  ( .A1(_AES_ENC_u0_u2_n931 ), .A2(_AES_ENC_u0_u2_n930 ), .ZN(_AES_ENC_u0_u2_n934 ) );
NOR3_X2 _AES_ENC_u0_u2_U479  ( .A1(_AES_ENC_u0_u2_n935 ), .A2(_AES_ENC_u0_u2_n934 ), .A3(_AES_ENC_u0_u2_n933 ), .ZN(_AES_ENC_u0_u2_n936 ) );
OR2_X4 _AES_ENC_u0_u2_U478  ( .A1(_AES_ENC_u0_u2_n1094 ), .A2(_AES_ENC_u0_u2_n1093 ), .ZN(_AES_ENC_u0_u2_n571 ) );
AND2_X2 _AES_ENC_u0_u2_U477  ( .A1(_AES_ENC_u0_u2_n571 ), .A2(_AES_ENC_u0_u2_n1095 ), .ZN(_AES_ENC_u0_u2_n1101 ) );
NOR2_X2 _AES_ENC_u0_u2_U474  ( .A1(_AES_ENC_u0_u2_n1074 ), .A2(_AES_ENC_u0_u2_n931 ), .ZN(_AES_ENC_u0_u2_n796 ) );
NOR2_X2 _AES_ENC_u0_u2_U473  ( .A1(_AES_ENC_u0_u2_n796 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n797 ) );
NOR2_X2 _AES_ENC_u0_u2_U472  ( .A1(_AES_ENC_u0_u2_n1054 ), .A2(_AES_ENC_u0_u2_n1053 ), .ZN(_AES_ENC_u0_u2_n1055 ) );
NOR2_X2 _AES_ENC_u0_u2_U471  ( .A1(_AES_ENC_u0_u2_n572 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n949 ) );
NOR2_X2 _AES_ENC_u0_u2_U470  ( .A1(_AES_ENC_u0_u2_n1049 ), .A2(_AES_ENC_u0_u2_n618 ), .ZN(_AES_ENC_u0_u2_n1051 ) );
NOR2_X2 _AES_ENC_u0_u2_U469  ( .A1(_AES_ENC_u0_u2_n1051 ), .A2(_AES_ENC_u0_u2_n1050 ), .ZN(_AES_ENC_u0_u2_n1052 ) );
NOR2_X2 _AES_ENC_u0_u2_U468  ( .A1(_AES_ENC_u0_u2_n1052 ), .A2(_AES_ENC_u0_u2_n592 ), .ZN(_AES_ENC_u0_u2_n1064 ) );
NOR2_X2 _AES_ENC_u0_u2_U467  ( .A1(_AES_ENC_w3[1] ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n631 ) );
NOR2_X2 _AES_ENC_u0_u2_U466  ( .A1(_AES_ENC_u0_u2_n1025 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n980 ) );
NOR2_X2 _AES_ENC_u0_u2_U465  ( .A1(_AES_ENC_u0_u2_n1074 ), .A2(_AES_ENC_u0_u2_n1025 ), .ZN(_AES_ENC_u0_u2_n891 ) );
NOR2_X2 _AES_ENC_u0_u2_U464  ( .A1(_AES_ENC_u0_u2_n891 ), .A2(_AES_ENC_u0_u2_n609 ), .ZN(_AES_ENC_u0_u2_n894 ) );
NOR2_X2 _AES_ENC_u0_u2_U463  ( .A1(_AES_ENC_u0_u2_n1073 ), .A2(_AES_ENC_u0_u2_n1094 ), .ZN(_AES_ENC_u0_u2_n795 ) );
NOR2_X2 _AES_ENC_u0_u2_U462  ( .A1(_AES_ENC_u0_u2_n795 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n799 ) );
NOR2_X2 _AES_ENC_u0_u2_U461  ( .A1(_AES_ENC_u0_u2_n624 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n1075 ) );
NOR2_X2 _AES_ENC_u0_u2_U460  ( .A1(_AES_ENC_u0_u2_n624 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n822 ) );
NOR2_X2 _AES_ENC_u0_u2_U459  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n823 ) );
NOR2_X2 _AES_ENC_u0_u2_U458  ( .A1(_AES_ENC_u0_u2_n823 ), .A2(_AES_ENC_u0_u2_n822 ), .ZN(_AES_ENC_u0_u2_n825 ) );
NOR2_X2 _AES_ENC_u0_u2_U455  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n981 ) );
NOR2_X2 _AES_ENC_u0_u2_U448  ( .A1(_AES_ENC_u0_u2_n1102 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n643 ) );
NOR2_X2 _AES_ENC_u0_u2_U447  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n621 ), .ZN(_AES_ENC_u0_u2_n642 ) );
NOR2_X2 _AES_ENC_u0_u2_U442  ( .A1(_AES_ENC_u0_u2_n911 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n644 ) );
NOR4_X2 _AES_ENC_u0_u2_U441  ( .A1(_AES_ENC_u0_u2_n644 ), .A2(_AES_ENC_u0_u2_n643 ), .A3(_AES_ENC_u0_u2_n804 ), .A4(_AES_ENC_u0_u2_n642 ), .ZN(_AES_ENC_u0_u2_n645 ) );
NOR2_X2 _AES_ENC_u0_u2_U438  ( .A1(_AES_ENC_u0_u2_n1102 ), .A2(_AES_ENC_u0_u2_n910 ), .ZN(_AES_ENC_u0_u2_n932 ) );
NOR3_X2 _AES_ENC_u0_u2_U435  ( .A1(_AES_ENC_u0_u2_n623 ), .A2(_AES_ENC_w3[1] ), .A3(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n683 ));
NOR2_X2 _AES_ENC_u0_u2_U434  ( .A1(_AES_ENC_u0_u2_n1102 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n755 ) );
INV_X4 _AES_ENC_u0_u2_U433  ( .A(_AES_ENC_u0_u2_n931 ), .ZN(_AES_ENC_u0_u2_n623 ) );
NOR2_X2 _AES_ENC_u0_u2_U428  ( .A1(_AES_ENC_u0_u2_n996 ), .A2(_AES_ENC_u0_u2_n931 ), .ZN(_AES_ENC_u0_u2_n704 ) );
NOR2_X2 _AES_ENC_u0_u2_U427  ( .A1(_AES_ENC_u0_u2_n1029 ), .A2(_AES_ENC_u0_u2_n1025 ), .ZN(_AES_ENC_u0_u2_n1079 ) );
NOR3_X2 _AES_ENC_u0_u2_U421  ( .A1(_AES_ENC_u0_u2_n589 ), .A2(_AES_ENC_u0_u2_n1025 ), .A3(_AES_ENC_u0_u2_n616 ), .ZN(_AES_ENC_u0_u2_n945 ) );
NOR2_X2 _AES_ENC_u0_u2_U420  ( .A1(_AES_ENC_u0_u2_n1072 ), .A2(_AES_ENC_u0_u2_n1094 ), .ZN(_AES_ENC_u0_u2_n930 ) );
NOR2_X2 _AES_ENC_u0_u2_U419  ( .A1(_AES_ENC_u0_u2_n931 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n743 ) );
NOR2_X2 _AES_ENC_u0_u2_U418  ( .A1(_AES_ENC_u0_u2_n931 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n685 ) );
NOR3_X2 _AES_ENC_u0_u2_U417  ( .A1(_AES_ENC_u0_u2_n610 ), .A2(_AES_ENC_u0_u2_n572 ), .A3(_AES_ENC_u0_u2_n575 ), .ZN(_AES_ENC_u0_u2_n962 ) );
NOR2_X2 _AES_ENC_u0_u2_U416  ( .A1(_AES_ENC_u0_u2_n626 ), .A2(_AES_ENC_u0_u2_n611 ), .ZN(_AES_ENC_u0_u2_n800 ) );
NOR3_X2 _AES_ENC_u0_u2_U415  ( .A1(_AES_ENC_u0_u2_n590 ), .A2(_AES_ENC_u0_u2_n627 ), .A3(_AES_ENC_u0_u2_n611 ), .ZN(_AES_ENC_u0_u2_n798 ) );
NOR3_X2 _AES_ENC_u0_u2_U414  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n572 ), .A3(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n694 ) );
NOR3_X2 _AES_ENC_u0_u2_U413  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n572 ), .A3(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n895 ) );
NOR3_X2 _AES_ENC_u0_u2_U410  ( .A1(_AES_ENC_u0_u2_n1008 ), .A2(_AES_ENC_u0_u2_n1007 ), .A3(_AES_ENC_u0_u2_n1006 ), .ZN(_AES_ENC_u0_u2_n1018 ) );
NOR4_X2 _AES_ENC_u0_u2_U409  ( .A1(_AES_ENC_u0_u2_n806 ), .A2(_AES_ENC_u0_u2_n805 ), .A3(_AES_ENC_u0_u2_n804 ), .A4(_AES_ENC_u0_u2_n803 ), .ZN(_AES_ENC_u0_u2_n807 ) );
NOR3_X2 _AES_ENC_u0_u2_U406  ( .A1(_AES_ENC_u0_u2_n799 ), .A2(_AES_ENC_u0_u2_n798 ), .A3(_AES_ENC_u0_u2_n797 ), .ZN(_AES_ENC_u0_u2_n808 ) );
NOR2_X2 _AES_ENC_u0_u2_U405  ( .A1(_AES_ENC_u0_u2_n669 ), .A2(_AES_ENC_u0_u2_n668 ), .ZN(_AES_ENC_u0_u2_n673 ) );
NOR4_X2 _AES_ENC_u0_u2_U404  ( .A1(_AES_ENC_u0_u2_n946 ), .A2(_AES_ENC_u0_u2_n1046 ), .A3(_AES_ENC_u0_u2_n671 ), .A4(_AES_ENC_u0_u2_n670 ), .ZN(_AES_ENC_u0_u2_n672 ) );
NOR4_X2 _AES_ENC_u0_u2_U403  ( .A1(_AES_ENC_u0_u2_n711 ), .A2(_AES_ENC_u0_u2_n710 ), .A3(_AES_ENC_u0_u2_n709 ), .A4(_AES_ENC_u0_u2_n708 ), .ZN(_AES_ENC_u0_u2_n712 ) );
NOR4_X2 _AES_ENC_u0_u2_U401  ( .A1(_AES_ENC_u0_u2_n843 ), .A2(_AES_ENC_u0_u2_n842 ), .A3(_AES_ENC_u0_u2_n841 ), .A4(_AES_ENC_u0_u2_n840 ), .ZN(_AES_ENC_u0_u2_n844 ) );
NOR3_X2 _AES_ENC_u0_u2_U400  ( .A1(_AES_ENC_u0_u2_n1101 ), .A2(_AES_ENC_u0_u2_n1100 ), .A3(_AES_ENC_u0_u2_n1099 ), .ZN(_AES_ENC_u0_u2_n1109 ) );
NOR3_X2 _AES_ENC_u0_u2_U399  ( .A1(_AES_ENC_u0_u2_n743 ), .A2(_AES_ENC_u0_u2_n742 ), .A3(_AES_ENC_u0_u2_n741 ), .ZN(_AES_ENC_u0_u2_n744 ) );
NOR2_X2 _AES_ENC_u0_u2_U398  ( .A1(_AES_ENC_u0_u2_n697 ), .A2(_AES_ENC_u0_u2_n658 ), .ZN(_AES_ENC_u0_u2_n659 ) );
NOR3_X2 _AES_ENC_u0_u2_U397  ( .A1(_AES_ENC_u0_u2_n959 ), .A2(_AES_ENC_u0_u2_n572 ), .A3(_AES_ENC_u0_u2_n609 ), .ZN(_AES_ENC_u0_u2_n768 ) );
NOR2_X2 _AES_ENC_u0_u2_U396  ( .A1(_AES_ENC_u0_u2_n1078 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n1033 ) );
NOR2_X2 _AES_ENC_u0_u2_U393  ( .A1(_AES_ENC_u0_u2_n1031 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n1032 ) );
NOR3_X2 _AES_ENC_u0_u2_U390  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n1025 ), .A3(_AES_ENC_u0_u2_n1074 ), .ZN(_AES_ENC_u0_u2_n1035 ) );
NOR4_X2 _AES_ENC_u0_u2_U389  ( .A1(_AES_ENC_u0_u2_n1035 ), .A2(_AES_ENC_u0_u2_n1034 ), .A3(_AES_ENC_u0_u2_n1033 ), .A4(_AES_ENC_u0_u2_n1032 ), .ZN(_AES_ENC_u0_u2_n1036 ) );
NOR2_X2 _AES_ENC_u0_u2_U388  ( .A1(_AES_ENC_u0_u2_n598 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n885 ) );
NOR2_X2 _AES_ENC_u0_u2_U387  ( .A1(_AES_ENC_u0_u2_n623 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n882 ) );
NOR2_X2 _AES_ENC_u0_u2_U386  ( .A1(_AES_ENC_u0_u2_n1053 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n884 ) );
NOR4_X2 _AES_ENC_u0_u2_U385  ( .A1(_AES_ENC_u0_u2_n885 ), .A2(_AES_ENC_u0_u2_n884 ), .A3(_AES_ENC_u0_u2_n883 ), .A4(_AES_ENC_u0_u2_n882 ), .ZN(_AES_ENC_u0_u2_n886 ) );
NOR2_X2 _AES_ENC_u0_u2_U384  ( .A1(_AES_ENC_u0_u2_n825 ), .A2(_AES_ENC_u0_u2_n578 ), .ZN(_AES_ENC_u0_u2_n830 ) );
NOR2_X2 _AES_ENC_u0_u2_U383  ( .A1(_AES_ENC_u0_u2_n827 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n829 ) );
NOR2_X2 _AES_ENC_u0_u2_U382  ( .A1(_AES_ENC_u0_u2_n572 ), .A2(_AES_ENC_u0_u2_n579 ), .ZN(_AES_ENC_u0_u2_n828 ) );
NOR4_X2 _AES_ENC_u0_u2_U374  ( .A1(_AES_ENC_u0_u2_n831 ), .A2(_AES_ENC_u0_u2_n830 ), .A3(_AES_ENC_u0_u2_n829 ), .A4(_AES_ENC_u0_u2_n828 ), .ZN(_AES_ENC_u0_u2_n832 ) );
NOR2_X2 _AES_ENC_u0_u2_U373  ( .A1(_AES_ENC_u0_u2_n598 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n1107 ) );
NOR2_X2 _AES_ENC_u0_u2_U372  ( .A1(_AES_ENC_u0_u2_n1102 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n1106 ) );
NOR2_X2 _AES_ENC_u0_u2_U370  ( .A1(_AES_ENC_u0_u2_n1103 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n1105 ) );
NOR4_X2 _AES_ENC_u0_u2_U369  ( .A1(_AES_ENC_u0_u2_n1107 ), .A2(_AES_ENC_u0_u2_n1106 ), .A3(_AES_ENC_u0_u2_n1105 ), .A4(_AES_ENC_u0_u2_n1104 ), .ZN(_AES_ENC_u0_u2_n1108 ) );
NOR3_X2 _AES_ENC_u0_u2_U368  ( .A1(_AES_ENC_u0_u2_n959 ), .A2(_AES_ENC_u0_u2_n621 ), .A3(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n963 ) );
NOR2_X2 _AES_ENC_u0_u2_U367  ( .A1(_AES_ENC_u0_u2_n626 ), .A2(_AES_ENC_u0_u2_n627 ), .ZN(_AES_ENC_u0_u2_n1114 ) );
NOR3_X2 _AES_ENC_u0_u2_U366  ( .A1(_AES_ENC_u0_u2_n910 ), .A2(_AES_ENC_u0_u2_n1059 ), .A3(_AES_ENC_u0_u2_n611 ), .ZN(_AES_ENC_u0_u2_n1115 ) );
INV_X4 _AES_ENC_u0_u2_U365  ( .A(_AES_ENC_u0_u2_n1024 ), .ZN(_AES_ENC_u0_u2_n606 ) );
INV_X4 _AES_ENC_u0_u2_U364  ( .A(_AES_ENC_u0_u2_n1094 ), .ZN(_AES_ENC_u0_u2_n613 ) );
NOR2_X2 _AES_ENC_u0_u2_U363  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n931 ), .ZN(_AES_ENC_u0_u2_n1100 ) );
NOR2_X2 _AES_ENC_u0_u2_U354  ( .A1(_AES_ENC_u0_u2_n569 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n929 ) );
NOR2_X2 _AES_ENC_u0_u2_U353  ( .A1(_AES_ENC_u0_u2_n620 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n926 ) );
INV_X4 _AES_ENC_u0_u2_U352  ( .A(_AES_ENC_u0_u2_n1093 ), .ZN(_AES_ENC_u0_u2_n617 ) );
NOR2_X2 _AES_ENC_u0_u2_U351  ( .A1(_AES_ENC_u0_u2_n572 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n1095 ) );
NOR2_X2 _AES_ENC_u0_u2_U350  ( .A1(_AES_ENC_u0_u2_n609 ), .A2(_AES_ENC_u0_u2_n627 ), .ZN(_AES_ENC_u0_u2_n1010 ) );
NOR2_X2 _AES_ENC_u0_u2_U349  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n1103 ) );
NOR2_X2 _AES_ENC_u0_u2_U348  ( .A1(_AES_ENC_w3[1] ), .A2(_AES_ENC_u0_u2_n1120 ), .ZN(_AES_ENC_u0_u2_n1022 ) );
NOR2_X2 _AES_ENC_u0_u2_U347  ( .A1(_AES_ENC_u0_u2_n619 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n911 ) );
NOR2_X2 _AES_ENC_u0_u2_U346  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_u0_u2_n1025 ), .ZN(_AES_ENC_u0_u2_n826 ) );
NOR2_X2 _AES_ENC_u0_u2_U345  ( .A1(_AES_ENC_u0_u2_n626 ), .A2(_AES_ENC_u0_u2_n607 ), .ZN(_AES_ENC_u0_u2_n1072 ) );
NOR2_X2 _AES_ENC_u0_u2_U338  ( .A1(_AES_ENC_u0_u2_n627 ), .A2(_AES_ENC_u0_u2_n616 ), .ZN(_AES_ENC_u0_u2_n956 ) );
NOR2_X2 _AES_ENC_u0_u2_U335  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_u0_u2_n624 ), .ZN(_AES_ENC_u0_u2_n1121 ) );
NOR2_X2 _AES_ENC_u0_u2_U329  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_u0_u2_n624 ), .ZN(_AES_ENC_u0_u2_n1058 ) );
NOR2_X2 _AES_ENC_u0_u2_U328  ( .A1(_AES_ENC_u0_u2_n625 ), .A2(_AES_ENC_u0_u2_n611 ), .ZN(_AES_ENC_u0_u2_n1073 ) );
NOR2_X2 _AES_ENC_u0_u2_U327  ( .A1(_AES_ENC_w3[1] ), .A2(_AES_ENC_u0_u2_n1025 ), .ZN(_AES_ENC_u0_u2_n1054 ) );
NOR2_X2 _AES_ENC_u0_u2_U325  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_u0_u2_n931 ), .ZN(_AES_ENC_u0_u2_n1029 ) );
NOR2_X2 _AES_ENC_u0_u2_U324  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n1056 ) );
NOR2_X2 _AES_ENC_u0_u2_U319  ( .A1(_AES_ENC_u0_u2_n614 ), .A2(_AES_ENC_u0_u2_n626 ), .ZN(_AES_ENC_u0_u2_n1050 ) );
NOR2_X2 _AES_ENC_u0_u2_U318  ( .A1(_AES_ENC_u0_u2_n1121 ), .A2(_AES_ENC_u0_u2_n1025 ), .ZN(_AES_ENC_u0_u2_n1120 ) );
NOR2_X2 _AES_ENC_u0_u2_U317  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_u0_u2_n572 ), .ZN(_AES_ENC_u0_u2_n1074 ) );
NOR2_X2 _AES_ENC_u0_u2_U316  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n584 ), .ZN(_AES_ENC_u0_u2_n838 ) );
NOR2_X2 _AES_ENC_u0_u2_U315  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n602 ), .ZN(_AES_ENC_u0_u2_n837 ) );
NOR2_X2 _AES_ENC_u0_u2_U314  ( .A1(_AES_ENC_u0_u2_n838 ), .A2(_AES_ENC_u0_u2_n837 ), .ZN(_AES_ENC_u0_u2_n845 ) );
NOR2_X2 _AES_ENC_u0_u2_U312  ( .A1(_AES_ENC_u0_u2_n1058 ), .A2(_AES_ENC_u0_u2_n1054 ), .ZN(_AES_ENC_u0_u2_n878 ) );
NOR2_X2 _AES_ENC_u0_u2_U311  ( .A1(_AES_ENC_u0_u2_n878 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n879 ) );
NOR2_X2 _AES_ENC_u0_u2_U310  ( .A1(_AES_ENC_u0_u2_n880 ), .A2(_AES_ENC_u0_u2_n879 ), .ZN(_AES_ENC_u0_u2_n887 ) );
NOR3_X2 _AES_ENC_u0_u2_U309  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n1091 ), .A3(_AES_ENC_u0_u2_n1022 ), .ZN(_AES_ENC_u0_u2_n720 ) );
NOR3_X2 _AES_ENC_u0_u2_U303  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n1054 ), .A3(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n719 ) );
NOR2_X2 _AES_ENC_u0_u2_U302  ( .A1(_AES_ENC_u0_u2_n720 ), .A2(_AES_ENC_u0_u2_n719 ), .ZN(_AES_ENC_u0_u2_n726 ) );
NOR2_X2 _AES_ENC_u0_u2_U300  ( .A1(_AES_ENC_u0_u2_n614 ), .A2(_AES_ENC_u0_u2_n591 ), .ZN(_AES_ENC_u0_u2_n865 ) );
NOR2_X2 _AES_ENC_u0_u2_U299  ( .A1(_AES_ENC_u0_u2_n1059 ), .A2(_AES_ENC_u0_u2_n1058 ), .ZN(_AES_ENC_u0_u2_n1060 ) );
NOR2_X2 _AES_ENC_u0_u2_U298  ( .A1(_AES_ENC_u0_u2_n1095 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n668 ) );
NOR2_X2 _AES_ENC_u0_u2_U297  ( .A1(_AES_ENC_u0_u2_n826 ), .A2(_AES_ENC_u0_u2_n573 ), .ZN(_AES_ENC_u0_u2_n750 ) );
NOR2_X2 _AES_ENC_u0_u2_U296  ( .A1(_AES_ENC_u0_u2_n750 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n751 ) );
NOR2_X2 _AES_ENC_u0_u2_U295  ( .A1(_AES_ENC_u0_u2_n907 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n908 ) );
NOR2_X2 _AES_ENC_u0_u2_U294  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n588 ), .ZN(_AES_ENC_u0_u2_n957 ) );
NOR2_X2 _AES_ENC_u0_u2_U293  ( .A1(_AES_ENC_u0_u2_n990 ), .A2(_AES_ENC_u0_u2_n926 ), .ZN(_AES_ENC_u0_u2_n780 ) );
NOR2_X2 _AES_ENC_u0_u2_U292  ( .A1(_AES_ENC_u0_u2_n1022 ), .A2(_AES_ENC_u0_u2_n1058 ), .ZN(_AES_ENC_u0_u2_n740 ) );
NOR2_X2 _AES_ENC_u0_u2_U291  ( .A1(_AES_ENC_u0_u2_n740 ), .A2(_AES_ENC_u0_u2_n616 ), .ZN(_AES_ENC_u0_u2_n742 ) );
NOR2_X2 _AES_ENC_u0_u2_U290  ( .A1(_AES_ENC_u0_u2_n1098 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n1099 ) );
NOR2_X2 _AES_ENC_u0_u2_U284  ( .A1(_AES_ENC_u0_u2_n1120 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n993 ) );
NOR2_X2 _AES_ENC_u0_u2_U283  ( .A1(_AES_ENC_u0_u2_n993 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n994 ) );
NOR2_X2 _AES_ENC_u0_u2_U282  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n620 ), .ZN(_AES_ENC_u0_u2_n1026 ) );
NOR2_X2 _AES_ENC_u0_u2_U281  ( .A1(_AES_ENC_u0_u2_n573 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n1027 ) );
NOR2_X2 _AES_ENC_u0_u2_U280  ( .A1(_AES_ENC_u0_u2_n1027 ), .A2(_AES_ENC_u0_u2_n1026 ), .ZN(_AES_ENC_u0_u2_n1028 ) );
NOR2_X2 _AES_ENC_u0_u2_U279  ( .A1(_AES_ENC_u0_u2_n1029 ), .A2(_AES_ENC_u0_u2_n1028 ), .ZN(_AES_ENC_u0_u2_n1034 ) );
NOR2_X2 _AES_ENC_u0_u2_U273  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n1071 ), .ZN(_AES_ENC_u0_u2_n669 ) );
NOR2_X2 _AES_ENC_u0_u2_U272  ( .A1(_AES_ENC_u0_u2_n1056 ), .A2(_AES_ENC_u0_u2_n990 ), .ZN(_AES_ENC_u0_u2_n991 ) );
NOR2_X2 _AES_ENC_u0_u2_U271  ( .A1(_AES_ENC_u0_u2_n991 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n995 ) );
NOR4_X2 _AES_ENC_u0_u2_U270  ( .A1(_AES_ENC_u0_u2_n757 ), .A2(_AES_ENC_u0_u2_n756 ), .A3(_AES_ENC_u0_u2_n755 ), .A4(_AES_ENC_u0_u2_n754 ), .ZN(_AES_ENC_u0_u2_n758 ) );
NOR2_X2 _AES_ENC_u0_u2_U269  ( .A1(_AES_ENC_u0_u2_n752 ), .A2(_AES_ENC_u0_u2_n751 ), .ZN(_AES_ENC_u0_u2_n759 ) );
NOR2_X2 _AES_ENC_u0_u2_U268  ( .A1(_AES_ENC_u0_u2_n607 ), .A2(_AES_ENC_u0_u2_n590 ), .ZN(_AES_ENC_u0_u2_n1008 ) );
NOR2_X2 _AES_ENC_u0_u2_U267  ( .A1(_AES_ENC_u0_u2_n606 ), .A2(_AES_ENC_u0_u2_n906 ), .ZN(_AES_ENC_u0_u2_n741 ) );
NOR2_X2 _AES_ENC_u0_u2_U263  ( .A1(_AES_ENC_u0_u2_n1054 ), .A2(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n763 ) );
NOR2_X2 _AES_ENC_u0_u2_U262  ( .A1(_AES_ENC_u0_u2_n763 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n769 ) );
NOR2_X2 _AES_ENC_u0_u2_U258  ( .A1(_AES_ENC_u0_u2_n839 ), .A2(_AES_ENC_u0_u2_n582 ), .ZN(_AES_ENC_u0_u2_n693 ) );
NOR2_X2 _AES_ENC_u0_u2_U255  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n577 ), .ZN(_AES_ENC_u0_u2_n1007 ) );
NOR2_X2 _AES_ENC_u0_u2_U254  ( .A1(_AES_ENC_u0_u2_n609 ), .A2(_AES_ENC_u0_u2_n580 ), .ZN(_AES_ENC_u0_u2_n1123 ) );
NOR2_X2 _AES_ENC_u0_u2_U253  ( .A1(_AES_ENC_u0_u2_n780 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n784 ) );
NOR2_X2 _AES_ENC_u0_u2_U252  ( .A1(_AES_ENC_u0_u2_n1117 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n782 ) );
NOR2_X2 _AES_ENC_u0_u2_U251  ( .A1(_AES_ENC_u0_u2_n781 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n783 ) );
NOR4_X2 _AES_ENC_u0_u2_U250  ( .A1(_AES_ENC_u0_u2_n880 ), .A2(_AES_ENC_u0_u2_n784 ), .A3(_AES_ENC_u0_u2_n783 ), .A4(_AES_ENC_u0_u2_n782 ), .ZN(_AES_ENC_u0_u2_n785 ) );
NOR2_X2 _AES_ENC_u0_u2_U243  ( .A1(_AES_ENC_u0_u2_n609 ), .A2(_AES_ENC_u0_u2_n590 ), .ZN(_AES_ENC_u0_u2_n710 ) );
INV_X4 _AES_ENC_u0_u2_U242  ( .A(_AES_ENC_u0_u2_n1029 ), .ZN(_AES_ENC_u0_u2_n582 ) );
NOR2_X2 _AES_ENC_u0_u2_U241  ( .A1(_AES_ENC_u0_u2_n593 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n1125 ) );
NOR2_X2 _AES_ENC_u0_u2_U240  ( .A1(_AES_ENC_u0_u2_n616 ), .A2(_AES_ENC_u0_u2_n580 ), .ZN(_AES_ENC_u0_u2_n771 ) );
NOR2_X2 _AES_ENC_u0_u2_U239  ( .A1(_AES_ENC_u0_u2_n616 ), .A2(_AES_ENC_u0_u2_n597 ), .ZN(_AES_ENC_u0_u2_n883 ) );
NOR2_X2 _AES_ENC_u0_u2_U238  ( .A1(_AES_ENC_u0_u2_n911 ), .A2(_AES_ENC_u0_u2_n910 ), .ZN(_AES_ENC_u0_u2_n912 ) );
NOR2_X2 _AES_ENC_u0_u2_U237  ( .A1(_AES_ENC_u0_u2_n912 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n916 ) );
NOR2_X2 _AES_ENC_u0_u2_U236  ( .A1(_AES_ENC_u0_u2_n990 ), .A2(_AES_ENC_u0_u2_n929 ), .ZN(_AES_ENC_u0_u2_n892 ) );
NOR2_X2 _AES_ENC_u0_u2_U235  ( .A1(_AES_ENC_u0_u2_n892 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n893 ) );
NOR2_X2 _AES_ENC_u0_u2_U234  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n602 ), .ZN(_AES_ENC_u0_u2_n950 ) );
NOR2_X2 _AES_ENC_u0_u2_U229  ( .A1(_AES_ENC_u0_u2_n1079 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n1082 ) );
NOR2_X2 _AES_ENC_u0_u2_U228  ( .A1(_AES_ENC_u0_u2_n910 ), .A2(_AES_ENC_u0_u2_n1056 ), .ZN(_AES_ENC_u0_u2_n941 ) );
NOR2_X2 _AES_ENC_u0_u2_U227  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n1077 ), .ZN(_AES_ENC_u0_u2_n841 ) );
NOR2_X2 _AES_ENC_u0_u2_U226  ( .A1(_AES_ENC_u0_u2_n623 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n630 ) );
NOR2_X2 _AES_ENC_u0_u2_U225  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n602 ), .ZN(_AES_ENC_u0_u2_n806 ) );
NOR2_X2 _AES_ENC_u0_u2_U223  ( .A1(_AES_ENC_u0_u2_n623 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n948 ) );
NOR2_X2 _AES_ENC_u0_u2_U222  ( .A1(_AES_ENC_u0_u2_n606 ), .A2(_AES_ENC_u0_u2_n582 ), .ZN(_AES_ENC_u0_u2_n1104 ) );
NOR2_X2 _AES_ENC_u0_u2_U221  ( .A1(_AES_ENC_u0_u2_n1121 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n1122 ) );
NOR2_X2 _AES_ENC_u0_u2_U217  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n1023 ), .ZN(_AES_ENC_u0_u2_n756 ) );
NOR2_X2 _AES_ENC_u0_u2_U213  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n602 ), .ZN(_AES_ENC_u0_u2_n870 ) );
NOR2_X2 _AES_ENC_u0_u2_U212  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n569 ), .ZN(_AES_ENC_u0_u2_n947 ) );
NOR2_X2 _AES_ENC_u0_u2_U211  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n1077 ), .ZN(_AES_ENC_u0_u2_n1084 ) );
NOR2_X2 _AES_ENC_u0_u2_U210  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n855 ), .ZN(_AES_ENC_u0_u2_n709 ) );
NOR2_X2 _AES_ENC_u0_u2_U209  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n589 ), .ZN(_AES_ENC_u0_u2_n868 ) );
NOR2_X2 _AES_ENC_u0_u2_U208  ( .A1(_AES_ENC_u0_u2_n1120 ), .A2(_AES_ENC_u0_u2_n839 ), .ZN(_AES_ENC_u0_u2_n842 ) );
NOR2_X2 _AES_ENC_u0_u2_U207  ( .A1(_AES_ENC_u0_u2_n1120 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n1124 ) );
NOR2_X2 _AES_ENC_u0_u2_U201  ( .A1(_AES_ENC_u0_u2_n1120 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n696 ) );
NOR2_X2 _AES_ENC_u0_u2_U200  ( .A1(_AES_ENC_u0_u2_n1074 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n1076 ) );
NOR2_X2 _AES_ENC_u0_u2_U199  ( .A1(_AES_ENC_u0_u2_n1074 ), .A2(_AES_ENC_u0_u2_n620 ), .ZN(_AES_ENC_u0_u2_n781 ) );
NOR3_X2 _AES_ENC_u0_u2_U198  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n1056 ), .A3(_AES_ENC_u0_u2_n990 ), .ZN(_AES_ENC_u0_u2_n979 ) );
NOR3_X2 _AES_ENC_u0_u2_U197  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n1058 ), .A3(_AES_ENC_u0_u2_n1059 ), .ZN(_AES_ENC_u0_u2_n854 ) );
NOR2_X2 _AES_ENC_u0_u2_U196  ( .A1(_AES_ENC_u0_u2_n996 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n869 ) );
NOR2_X2 _AES_ENC_u0_u2_U195  ( .A1(_AES_ENC_u0_u2_n1056 ), .A2(_AES_ENC_u0_u2_n1074 ), .ZN(_AES_ENC_u0_u2_n1057 ) );
NOR3_X2 _AES_ENC_u0_u2_U194  ( .A1(_AES_ENC_u0_u2_n607 ), .A2(_AES_ENC_u0_u2_n1120 ), .A3(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n978 ) );
NOR2_X2 _AES_ENC_u0_u2_U187  ( .A1(_AES_ENC_u0_u2_n996 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n998 ) );
NOR2_X2 _AES_ENC_u0_u2_U186  ( .A1(_AES_ENC_u0_u2_n996 ), .A2(_AES_ENC_u0_u2_n911 ), .ZN(_AES_ENC_u0_u2_n1116 ) );
NOR2_X2 _AES_ENC_u0_u2_U185  ( .A1(_AES_ENC_u0_u2_n1074 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n754 ) );
NOR2_X2 _AES_ENC_u0_u2_U184  ( .A1(_AES_ENC_u0_u2_n926 ), .A2(_AES_ENC_u0_u2_n1103 ), .ZN(_AES_ENC_u0_u2_n977 ) );
NOR2_X2 _AES_ENC_u0_u2_U183  ( .A1(_AES_ENC_u0_u2_n839 ), .A2(_AES_ENC_u0_u2_n824 ), .ZN(_AES_ENC_u0_u2_n1092 ) );
NOR2_X2 _AES_ENC_u0_u2_U182  ( .A1(_AES_ENC_u0_u2_n573 ), .A2(_AES_ENC_u0_u2_n1074 ), .ZN(_AES_ENC_u0_u2_n684 ) );
NOR2_X2 _AES_ENC_u0_u2_U181  ( .A1(_AES_ENC_u0_u2_n826 ), .A2(_AES_ENC_u0_u2_n1059 ), .ZN(_AES_ENC_u0_u2_n907 ) );
NOR3_X2 _AES_ENC_u0_u2_U180  ( .A1(_AES_ENC_u0_u2_n625 ), .A2(_AES_ENC_u0_u2_n1115 ), .A3(_AES_ENC_u0_u2_n585 ), .ZN(_AES_ENC_u0_u2_n831 ) );
NOR3_X2 _AES_ENC_u0_u2_U174  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n1056 ), .A3(_AES_ENC_u0_u2_n990 ), .ZN(_AES_ENC_u0_u2_n896 ) );
NOR3_X2 _AES_ENC_u0_u2_U173  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n573 ), .A3(_AES_ENC_u0_u2_n1013 ), .ZN(_AES_ENC_u0_u2_n670 ) );
NOR3_X2 _AES_ENC_u0_u2_U172  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n1091 ), .A3(_AES_ENC_u0_u2_n1022 ), .ZN(_AES_ENC_u0_u2_n843 ) );
NOR2_X2 _AES_ENC_u0_u2_U171  ( .A1(_AES_ENC_u0_u2_n1029 ), .A2(_AES_ENC_u0_u2_n1095 ), .ZN(_AES_ENC_u0_u2_n735 ) );
NOR2_X2 _AES_ENC_u0_u2_U170  ( .A1(_AES_ENC_u0_u2_n1100 ), .A2(_AES_ENC_u0_u2_n854 ), .ZN(_AES_ENC_u0_u2_n860 ) );
NOR4_X2 _AES_ENC_u0_u2_U169  ( .A1(_AES_ENC_u0_u2_n1125 ), .A2(_AES_ENC_u0_u2_n1124 ), .A3(_AES_ENC_u0_u2_n1123 ), .A4(_AES_ENC_u0_u2_n1122 ), .ZN(_AES_ENC_u0_u2_n1126 ) );
NOR4_X2 _AES_ENC_u0_u2_U168  ( .A1(_AES_ENC_u0_u2_n1084 ), .A2(_AES_ENC_u0_u2_n1083 ), .A3(_AES_ENC_u0_u2_n1082 ), .A4(_AES_ENC_u0_u2_n1081 ), .ZN(_AES_ENC_u0_u2_n1085 ) );
NOR2_X2 _AES_ENC_u0_u2_U162  ( .A1(_AES_ENC_u0_u2_n1076 ), .A2(_AES_ENC_u0_u2_n1075 ), .ZN(_AES_ENC_u0_u2_n1086 ) );
NAND3_X2 _AES_ENC_u0_u2_U161  ( .A1(_AES_ENC_u0_u2_n569 ), .A2(_AES_ENC_u0_u2_n582 ), .A3(_AES_ENC_u0_u2_n681 ), .ZN(_AES_ENC_u0_u2_n691 ) );
NOR2_X2 _AES_ENC_u0_u2_U160  ( .A1(_AES_ENC_u0_u2_n683 ), .A2(_AES_ENC_u0_u2_n682 ), .ZN(_AES_ENC_u0_u2_n690 ) );
NOR4_X2 _AES_ENC_u0_u2_U159  ( .A1(_AES_ENC_u0_u2_n983 ), .A2(_AES_ENC_u0_u2_n698 ), .A3(_AES_ENC_u0_u2_n697 ), .A4(_AES_ENC_u0_u2_n696 ), .ZN(_AES_ENC_u0_u2_n699 ) );
NOR3_X2 _AES_ENC_u0_u2_U158  ( .A1(_AES_ENC_u0_u2_n695 ), .A2(_AES_ENC_u0_u2_n694 ), .A3(_AES_ENC_u0_u2_n693 ), .ZN(_AES_ENC_u0_u2_n700 ) );
NOR4_X2 _AES_ENC_u0_u2_U157  ( .A1(_AES_ENC_u0_u2_n896 ), .A2(_AES_ENC_u0_u2_n895 ), .A3(_AES_ENC_u0_u2_n894 ), .A4(_AES_ENC_u0_u2_n893 ), .ZN(_AES_ENC_u0_u2_n897 ) );
NOR2_X2 _AES_ENC_u0_u2_U156  ( .A1(_AES_ENC_u0_u2_n866 ), .A2(_AES_ENC_u0_u2_n865 ), .ZN(_AES_ENC_u0_u2_n872 ) );
NOR4_X2 _AES_ENC_u0_u2_U155  ( .A1(_AES_ENC_u0_u2_n870 ), .A2(_AES_ENC_u0_u2_n869 ), .A3(_AES_ENC_u0_u2_n868 ), .A4(_AES_ENC_u0_u2_n867 ), .ZN(_AES_ENC_u0_u2_n871 ) );
NOR4_X2 _AES_ENC_u0_u2_U154  ( .A1(_AES_ENC_u0_u2_n963 ), .A2(_AES_ENC_u0_u2_n962 ), .A3(_AES_ENC_u0_u2_n961 ), .A4(_AES_ENC_u0_u2_n960 ), .ZN(_AES_ENC_u0_u2_n964 ) );
NOR2_X2 _AES_ENC_u0_u2_U153  ( .A1(_AES_ENC_u0_u2_n958 ), .A2(_AES_ENC_u0_u2_n957 ), .ZN(_AES_ENC_u0_u2_n965 ) );
NOR4_X2 _AES_ENC_u0_u2_U152  ( .A1(_AES_ENC_u0_u2_n950 ), .A2(_AES_ENC_u0_u2_n949 ), .A3(_AES_ENC_u0_u2_n948 ), .A4(_AES_ENC_u0_u2_n947 ), .ZN(_AES_ENC_u0_u2_n951 ) );
NOR2_X2 _AES_ENC_u0_u2_U143  ( .A1(_AES_ENC_u0_u2_n946 ), .A2(_AES_ENC_u0_u2_n945 ), .ZN(_AES_ENC_u0_u2_n952 ) );
NOR4_X2 _AES_ENC_u0_u2_U142  ( .A1(_AES_ENC_u0_u2_n983 ), .A2(_AES_ENC_u0_u2_n982 ), .A3(_AES_ENC_u0_u2_n981 ), .A4(_AES_ENC_u0_u2_n980 ), .ZN(_AES_ENC_u0_u2_n984 ) );
NOR2_X2 _AES_ENC_u0_u2_U141  ( .A1(_AES_ENC_u0_u2_n979 ), .A2(_AES_ENC_u0_u2_n978 ), .ZN(_AES_ENC_u0_u2_n985 ) );
NOR3_X2 _AES_ENC_u0_u2_U140  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n1054 ), .A3(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n961 ) );
NOR3_X2 _AES_ENC_u0_u2_U132  ( .A1(_AES_ENC_u0_u2_n620 ), .A2(_AES_ENC_u0_u2_n1074 ), .A3(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n671 ) );
NOR2_X2 _AES_ENC_u0_u2_U131  ( .A1(_AES_ENC_u0_u2_n1057 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n1062 ) );
NOR2_X2 _AES_ENC_u0_u2_U130  ( .A1(_AES_ENC_u0_u2_n1060 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n1061 ) );
NOR2_X2 _AES_ENC_u0_u2_U129  ( .A1(_AES_ENC_u0_u2_n1055 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n1063 ) );
NOR4_X2 _AES_ENC_u0_u2_U128  ( .A1(_AES_ENC_u0_u2_n1064 ), .A2(_AES_ENC_u0_u2_n1063 ), .A3(_AES_ENC_u0_u2_n1062 ), .A4(_AES_ENC_u0_u2_n1061 ), .ZN(_AES_ENC_u0_u2_n1065 ) );
NOR3_X2 _AES_ENC_u0_u2_U127  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n1120 ), .A3(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n918 ) );
NOR2_X2 _AES_ENC_u0_u2_U126  ( .A1(_AES_ENC_u0_u2_n914 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n915 ) );
NOR3_X2 _AES_ENC_u0_u2_U121  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n573 ), .A3(_AES_ENC_u0_u2_n1013 ), .ZN(_AES_ENC_u0_u2_n917 ) );
NOR4_X2 _AES_ENC_u0_u2_U120  ( .A1(_AES_ENC_u0_u2_n918 ), .A2(_AES_ENC_u0_u2_n917 ), .A3(_AES_ENC_u0_u2_n916 ), .A4(_AES_ENC_u0_u2_n915 ), .ZN(_AES_ENC_u0_u2_n919 ) );
NOR2_X2 _AES_ENC_u0_u2_U119  ( .A1(_AES_ENC_u0_u2_n735 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n687 ) );
NOR2_X2 _AES_ENC_u0_u2_U118  ( .A1(_AES_ENC_u0_u2_n684 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n688 ) );
NOR2_X2 _AES_ENC_u0_u2_U117  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n600 ), .ZN(_AES_ENC_u0_u2_n686 ) );
NOR4_X2 _AES_ENC_u0_u2_U116  ( .A1(_AES_ENC_u0_u2_n688 ), .A2(_AES_ENC_u0_u2_n687 ), .A3(_AES_ENC_u0_u2_n686 ), .A4(_AES_ENC_u0_u2_n685 ), .ZN(_AES_ENC_u0_u2_n689 ) );
NOR2_X2 _AES_ENC_u0_u2_U115  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n582 ), .ZN(_AES_ENC_u0_u2_n770 ) );
NOR2_X2 _AES_ENC_u0_u2_U106  ( .A1(_AES_ENC_u0_u2_n1103 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n772 ) );
NOR2_X2 _AES_ENC_u0_u2_U105  ( .A1(_AES_ENC_u0_u2_n610 ), .A2(_AES_ENC_u0_u2_n599 ), .ZN(_AES_ENC_u0_u2_n773 ) );
NOR4_X2 _AES_ENC_u0_u2_U104  ( .A1(_AES_ENC_u0_u2_n773 ), .A2(_AES_ENC_u0_u2_n772 ), .A3(_AES_ENC_u0_u2_n771 ), .A4(_AES_ENC_u0_u2_n770 ), .ZN(_AES_ENC_u0_u2_n774 ) );
NOR2_X2 _AES_ENC_u0_u2_U103  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n595 ), .ZN(_AES_ENC_u0_u2_n858 ) );
NOR2_X2 _AES_ENC_u0_u2_U102  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n855 ), .ZN(_AES_ENC_u0_u2_n857 ) );
NOR2_X2 _AES_ENC_u0_u2_U101  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n587 ), .ZN(_AES_ENC_u0_u2_n856 ) );
NOR4_X2 _AES_ENC_u0_u2_U100  ( .A1(_AES_ENC_u0_u2_n858 ), .A2(_AES_ENC_u0_u2_n857 ), .A3(_AES_ENC_u0_u2_n856 ), .A4(_AES_ENC_u0_u2_n958 ), .ZN(_AES_ENC_u0_u2_n859 ) );
NOR2_X2 _AES_ENC_u0_u2_U95  ( .A1(_AES_ENC_u0_u2_n583 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n814 ) );
NOR3_X2 _AES_ENC_u0_u2_U94  ( .A1(_AES_ENC_u0_u2_n606 ), .A2(_AES_ENC_u0_u2_n1058 ), .A3(_AES_ENC_u0_u2_n1059 ), .ZN(_AES_ENC_u0_u2_n815 ) );
NOR2_X2 _AES_ENC_u0_u2_U93  ( .A1(_AES_ENC_u0_u2_n907 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n813 ) );
NOR4_X2 _AES_ENC_u0_u2_U92  ( .A1(_AES_ENC_u0_u2_n815 ), .A2(_AES_ENC_u0_u2_n814 ), .A3(_AES_ENC_u0_u2_n813 ), .A4(_AES_ENC_u0_u2_n812 ), .ZN(_AES_ENC_u0_u2_n816 ) );
NOR2_X2 _AES_ENC_u0_u2_U91  ( .A1(_AES_ENC_u0_u2_n617 ), .A2(_AES_ENC_u0_u2_n569 ), .ZN(_AES_ENC_u0_u2_n721 ) );
NOR2_X2 _AES_ENC_u0_u2_U90  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n1096 ), .ZN(_AES_ENC_u0_u2_n722 ) );
NOR2_X2 _AES_ENC_u0_u2_U89  ( .A1(_AES_ENC_u0_u2_n1031 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n723 ) );
NOR4_X2 _AES_ENC_u0_u2_U88  ( .A1(_AES_ENC_u0_u2_n724 ), .A2(_AES_ENC_u0_u2_n723 ), .A3(_AES_ENC_u0_u2_n722 ), .A4(_AES_ENC_u0_u2_n721 ), .ZN(_AES_ENC_u0_u2_n725 ) );
NOR2_X2 _AES_ENC_u0_u2_U87  ( .A1(_AES_ENC_u0_u2_n911 ), .A2(_AES_ENC_u0_u2_n990 ), .ZN(_AES_ENC_u0_u2_n1009 ) );
NOR2_X2 _AES_ENC_u0_u2_U86  ( .A1(_AES_ENC_u0_u2_n1013 ), .A2(_AES_ENC_u0_u2_n573 ), .ZN(_AES_ENC_u0_u2_n1014 ) );
NOR2_X2 _AES_ENC_u0_u2_U81  ( .A1(_AES_ENC_u0_u2_n1014 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n1015 ) );
NOR4_X2 _AES_ENC_u0_u2_U80  ( .A1(_AES_ENC_u0_u2_n1016 ), .A2(_AES_ENC_u0_u2_n1015 ), .A3(_AES_ENC_u0_u2_n1119 ), .A4(_AES_ENC_u0_u2_n1046 ), .ZN(_AES_ENC_u0_u2_n1017 ) );
NOR2_X2 _AES_ENC_u0_u2_U79  ( .A1(_AES_ENC_u0_u2_n606 ), .A2(_AES_ENC_u0_u2_n589 ), .ZN(_AES_ENC_u0_u2_n997 ) );
NOR2_X2 _AES_ENC_u0_u2_U78  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n577 ), .ZN(_AES_ENC_u0_u2_n1000 ) );
NOR2_X2 _AES_ENC_u0_u2_U74  ( .A1(_AES_ENC_u0_u2_n616 ), .A2(_AES_ENC_u0_u2_n1096 ), .ZN(_AES_ENC_u0_u2_n999 ) );
NOR4_X2 _AES_ENC_u0_u2_U73  ( .A1(_AES_ENC_u0_u2_n1000 ), .A2(_AES_ENC_u0_u2_n999 ), .A3(_AES_ENC_u0_u2_n998 ), .A4(_AES_ENC_u0_u2_n997 ), .ZN(_AES_ENC_u0_u2_n1001 ) );
NOR2_X2 _AES_ENC_u0_u2_U72  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n1096 ), .ZN(_AES_ENC_u0_u2_n697 ) );
NOR2_X2 _AES_ENC_u0_u2_U71  ( .A1(_AES_ENC_u0_u2_n620 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n958 ) );
NOR2_X2 _AES_ENC_u0_u2_U65  ( .A1(_AES_ENC_u0_u2_n911 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n983 ) );
NOR2_X2 _AES_ENC_u0_u2_U64  ( .A1(_AES_ENC_u0_u2_n1054 ), .A2(_AES_ENC_u0_u2_n1103 ), .ZN(_AES_ENC_u0_u2_n1031 ) );
INV_X4 _AES_ENC_u0_u2_U63  ( .A(_AES_ENC_u0_u2_n1050 ), .ZN(_AES_ENC_u0_u2_n612 ) );
INV_X4 _AES_ENC_u0_u2_U62  ( .A(_AES_ENC_u0_u2_n1072 ), .ZN(_AES_ENC_u0_u2_n605 ) );
INV_X4 _AES_ENC_u0_u2_U61  ( .A(_AES_ENC_u0_u2_n1073 ), .ZN(_AES_ENC_u0_u2_n604 ) );
NOR2_X2 _AES_ENC_u0_u2_U59  ( .A1(_AES_ENC_u0_u2_n582 ), .A2(_AES_ENC_u0_u2_n613 ), .ZN(_AES_ENC_u0_u2_n880 ) );
NOR3_X2 _AES_ENC_u0_u2_U58  ( .A1(_AES_ENC_u0_u2_n826 ), .A2(_AES_ENC_u0_u2_n1121 ), .A3(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n946 ) );
INV_X4 _AES_ENC_u0_u2_U57  ( .A(_AES_ENC_u0_u2_n1010 ), .ZN(_AES_ENC_u0_u2_n608 ) );
NOR3_X2 _AES_ENC_u0_u2_U50  ( .A1(_AES_ENC_u0_u2_n573 ), .A2(_AES_ENC_u0_u2_n1029 ), .A3(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n1119 ) );
INV_X4 _AES_ENC_u0_u2_U49  ( .A(_AES_ENC_u0_u2_n956 ), .ZN(_AES_ENC_u0_u2_n615 ) );
NOR2_X2 _AES_ENC_u0_u2_U48  ( .A1(_AES_ENC_u0_u2_n623 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n1013 ) );
NOR2_X2 _AES_ENC_u0_u2_U47  ( .A1(_AES_ENC_u0_u2_n620 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n910 ) );
NOR2_X2 _AES_ENC_u0_u2_U46  ( .A1(_AES_ENC_u0_u2_n569 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n1091 ) );
NOR2_X2 _AES_ENC_u0_u2_U45  ( .A1(_AES_ENC_u0_u2_n622 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n990 ) );
NOR2_X2 _AES_ENC_u0_u2_U44  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_u0_u2_n1121 ), .ZN(_AES_ENC_u0_u2_n996 ) );
NOR2_X2 _AES_ENC_u0_u2_U43  ( .A1(_AES_ENC_u0_u2_n610 ), .A2(_AES_ENC_u0_u2_n600 ), .ZN(_AES_ENC_u0_u2_n628 ) );
NOR2_X2 _AES_ENC_u0_u2_U42  ( .A1(_AES_ENC_u0_u2_n576 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n866 ) );
NOR2_X2 _AES_ENC_u0_u2_U41  ( .A1(_AES_ENC_u0_u2_n603 ), .A2(_AES_ENC_u0_u2_n610 ), .ZN(_AES_ENC_u0_u2_n1006 ) );
NOR2_X2 _AES_ENC_u0_u2_U36  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n1117 ), .ZN(_AES_ENC_u0_u2_n1118 ) );
NOR2_X2 _AES_ENC_u0_u2_U35  ( .A1(_AES_ENC_u0_u2_n1119 ), .A2(_AES_ENC_u0_u2_n1118 ), .ZN(_AES_ENC_u0_u2_n1127 ) );
NOR2_X2 _AES_ENC_u0_u2_U34  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n594 ), .ZN(_AES_ENC_u0_u2_n629 ) );
NOR2_X2 _AES_ENC_u0_u2_U33  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n906 ), .ZN(_AES_ENC_u0_u2_n909 ) );
NOR2_X2 _AES_ENC_u0_u2_U32  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n597 ), .ZN(_AES_ENC_u0_u2_n658 ) );
NOR2_X2 _AES_ENC_u0_u2_U31  ( .A1(_AES_ENC_u0_u2_n1116 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n695 ) );
NOR2_X2 _AES_ENC_u0_u2_U30  ( .A1(_AES_ENC_u0_u2_n1078 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n1083 ) );
NOR2_X2 _AES_ENC_u0_u2_U29  ( .A1(_AES_ENC_u0_u2_n941 ), .A2(_AES_ENC_u0_u2_n608 ), .ZN(_AES_ENC_u0_u2_n724 ) );
NOR2_X2 _AES_ENC_u0_u2_U24  ( .A1(_AES_ENC_u0_u2_n576 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n840 ) );
NOR2_X2 _AES_ENC_u0_u2_U23  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n593 ), .ZN(_AES_ENC_u0_u2_n633 ) );
NOR2_X2 _AES_ENC_u0_u2_U21  ( .A1(_AES_ENC_u0_u2_n1009 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n960 ) );
NOR2_X2 _AES_ENC_u0_u2_U20  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n1045 ), .ZN(_AES_ENC_u0_u2_n812 ) );
NOR2_X2 _AES_ENC_u0_u2_U19  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n1080 ), .ZN(_AES_ENC_u0_u2_n1081 ) );
NOR2_X2 _AES_ENC_u0_u2_U18  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n601 ), .ZN(_AES_ENC_u0_u2_n982 ) );
NOR2_X2 _AES_ENC_u0_u2_U17  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n594 ), .ZN(_AES_ENC_u0_u2_n757 ) );
NOR2_X2 _AES_ENC_u0_u2_U16  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n590 ), .ZN(_AES_ENC_u0_u2_n698 ) );
NOR2_X2 _AES_ENC_u0_u2_U15  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n619 ), .ZN(_AES_ENC_u0_u2_n708 ) );
NOR2_X2 _AES_ENC_u0_u2_U10  ( .A1(_AES_ENC_u0_u2_n619 ), .A2(_AES_ENC_u0_u2_n604 ), .ZN(_AES_ENC_u0_u2_n803 ) );
NOR2_X2 _AES_ENC_u0_u2_U9  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n881 ), .ZN(_AES_ENC_u0_u2_n711 ) );
NOR2_X2 _AES_ENC_u0_u2_U8  ( .A1(_AES_ENC_u0_u2_n615 ), .A2(_AES_ENC_u0_u2_n582 ), .ZN(_AES_ENC_u0_u2_n867 ) );
NOR2_X2 _AES_ENC_u0_u2_U7  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n599 ), .ZN(_AES_ENC_u0_u2_n804 ) );
NOR2_X2 _AES_ENC_u0_u2_U6  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n620 ), .ZN(_AES_ENC_u0_u2_n1046 ) );
OR2_X4 _AES_ENC_u0_u2_U5  ( .A1(_AES_ENC_u0_u2_n624 ), .A2(_AES_ENC_w3[1] ),.ZN(_AES_ENC_u0_u2_n570 ) );
OR2_X4 _AES_ENC_u0_u2_U4  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_w3[4] ),.ZN(_AES_ENC_u0_u2_n569 ) );
NAND2_X2 _AES_ENC_u0_u2_U514  ( .A1(_AES_ENC_u0_u2_n1121 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n1030 ) );
AND2_X2 _AES_ENC_u0_u2_U513  ( .A1(_AES_ENC_u0_u2_n597 ), .A2(_AES_ENC_u0_u2_n1030 ), .ZN(_AES_ENC_u0_u2_n1049 ) );
NAND2_X2 _AES_ENC_u0_u2_U511  ( .A1(_AES_ENC_u0_u2_n1049 ), .A2(_AES_ENC_u0_u2_n794 ), .ZN(_AES_ENC_u0_u2_n637 ) );
AND2_X2 _AES_ENC_u0_u2_U493  ( .A1(_AES_ENC_u0_u2_n779 ), .A2(_AES_ENC_u0_u2_n996 ), .ZN(_AES_ENC_u0_u2_n632 ) );
NAND4_X2 _AES_ENC_u0_u2_U485  ( .A1(_AES_ENC_u0_u2_n637 ), .A2(_AES_ENC_u0_u2_n636 ), .A3(_AES_ENC_u0_u2_n635 ), .A4(_AES_ENC_u0_u2_n634 ), .ZN(_AES_ENC_u0_u2_n638 ) );
NAND2_X2 _AES_ENC_u0_u2_U484  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n638 ), .ZN(_AES_ENC_u0_u2_n679 ) );
NAND2_X2 _AES_ENC_u0_u2_U481  ( .A1(_AES_ENC_u0_u2_n1094 ), .A2(_AES_ENC_u0_u2_n591 ), .ZN(_AES_ENC_u0_u2_n648 ) );
NAND2_X2 _AES_ENC_u0_u2_U476  ( .A1(_AES_ENC_u0_u2_n601 ), .A2(_AES_ENC_u0_u2_n590 ), .ZN(_AES_ENC_u0_u2_n762 ) );
NAND2_X2 _AES_ENC_u0_u2_U475  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n762 ), .ZN(_AES_ENC_u0_u2_n647 ) );
NAND4_X2 _AES_ENC_u0_u2_U457  ( .A1(_AES_ENC_u0_u2_n648 ), .A2(_AES_ENC_u0_u2_n647 ), .A3(_AES_ENC_u0_u2_n646 ), .A4(_AES_ENC_u0_u2_n645 ), .ZN(_AES_ENC_u0_u2_n649 ) );
NAND2_X2 _AES_ENC_u0_u2_U456  ( .A1(_AES_ENC_w3[0] ), .A2(_AES_ENC_u0_u2_n649 ), .ZN(_AES_ENC_u0_u2_n665 ) );
NAND2_X2 _AES_ENC_u0_u2_U454  ( .A1(_AES_ENC_u0_u2_n596 ), .A2(_AES_ENC_u0_u2_n623 ), .ZN(_AES_ENC_u0_u2_n855 ) );
NAND2_X2 _AES_ENC_u0_u2_U453  ( .A1(_AES_ENC_u0_u2_n587 ), .A2(_AES_ENC_u0_u2_n855 ), .ZN(_AES_ENC_u0_u2_n821 ) );
NAND2_X2 _AES_ENC_u0_u2_U452  ( .A1(_AES_ENC_u0_u2_n1093 ), .A2(_AES_ENC_u0_u2_n821 ), .ZN(_AES_ENC_u0_u2_n662 ) );
NAND2_X2 _AES_ENC_u0_u2_U451  ( .A1(_AES_ENC_u0_u2_n619 ), .A2(_AES_ENC_u0_u2_n589 ), .ZN(_AES_ENC_u0_u2_n650 ) );
NAND2_X2 _AES_ENC_u0_u2_U450  ( .A1(_AES_ENC_u0_u2_n956 ), .A2(_AES_ENC_u0_u2_n650 ), .ZN(_AES_ENC_u0_u2_n661 ) );
NAND2_X2 _AES_ENC_u0_u2_U449  ( .A1(_AES_ENC_u0_u2_n626 ), .A2(_AES_ENC_u0_u2_n627 ), .ZN(_AES_ENC_u0_u2_n839 ) );
OR2_X2 _AES_ENC_u0_u2_U446  ( .A1(_AES_ENC_u0_u2_n839 ), .A2(_AES_ENC_u0_u2_n932 ), .ZN(_AES_ENC_u0_u2_n656 ) );
NAND2_X2 _AES_ENC_u0_u2_U445  ( .A1(_AES_ENC_u0_u2_n621 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n1096 ) );
NAND2_X2 _AES_ENC_u0_u2_U444  ( .A1(_AES_ENC_u0_u2_n1030 ), .A2(_AES_ENC_u0_u2_n1096 ), .ZN(_AES_ENC_u0_u2_n651 ) );
NAND2_X2 _AES_ENC_u0_u2_U443  ( .A1(_AES_ENC_u0_u2_n1114 ), .A2(_AES_ENC_u0_u2_n651 ), .ZN(_AES_ENC_u0_u2_n655 ) );
OR3_X2 _AES_ENC_u0_u2_U440  ( .A1(_AES_ENC_u0_u2_n1079 ), .A2(_AES_ENC_w3[7] ), .A3(_AES_ENC_u0_u2_n626 ), .ZN(_AES_ENC_u0_u2_n654 ));
NAND2_X2 _AES_ENC_u0_u2_U439  ( .A1(_AES_ENC_u0_u2_n593 ), .A2(_AES_ENC_u0_u2_n601 ), .ZN(_AES_ENC_u0_u2_n652 ) );
NAND4_X2 _AES_ENC_u0_u2_U437  ( .A1(_AES_ENC_u0_u2_n656 ), .A2(_AES_ENC_u0_u2_n655 ), .A3(_AES_ENC_u0_u2_n654 ), .A4(_AES_ENC_u0_u2_n653 ), .ZN(_AES_ENC_u0_u2_n657 ) );
NAND2_X2 _AES_ENC_u0_u2_U436  ( .A1(_AES_ENC_w3[2] ), .A2(_AES_ENC_u0_u2_n657 ), .ZN(_AES_ENC_u0_u2_n660 ) );
NAND4_X2 _AES_ENC_u0_u2_U432  ( .A1(_AES_ENC_u0_u2_n662 ), .A2(_AES_ENC_u0_u2_n661 ), .A3(_AES_ENC_u0_u2_n660 ), .A4(_AES_ENC_u0_u2_n659 ), .ZN(_AES_ENC_u0_u2_n663 ) );
NAND2_X2 _AES_ENC_u0_u2_U431  ( .A1(_AES_ENC_u0_u2_n663 ), .A2(_AES_ENC_u0_u2_n574 ), .ZN(_AES_ENC_u0_u2_n664 ) );
NAND2_X2 _AES_ENC_u0_u2_U430  ( .A1(_AES_ENC_u0_u2_n665 ), .A2(_AES_ENC_u0_u2_n664 ), .ZN(_AES_ENC_u0_u2_n666 ) );
NAND2_X2 _AES_ENC_u0_u2_U429  ( .A1(_AES_ENC_w3[6] ), .A2(_AES_ENC_u0_u2_n666 ), .ZN(_AES_ENC_u0_u2_n678 ) );
NAND2_X2 _AES_ENC_u0_u2_U426  ( .A1(_AES_ENC_u0_u2_n735 ), .A2(_AES_ENC_u0_u2_n1093 ), .ZN(_AES_ENC_u0_u2_n675 ) );
NAND2_X2 _AES_ENC_u0_u2_U425  ( .A1(_AES_ENC_u0_u2_n588 ), .A2(_AES_ENC_u0_u2_n597 ), .ZN(_AES_ENC_u0_u2_n1045 ) );
OR2_X2 _AES_ENC_u0_u2_U424  ( .A1(_AES_ENC_u0_u2_n1045 ), .A2(_AES_ENC_u0_u2_n605 ), .ZN(_AES_ENC_u0_u2_n674 ) );
NAND2_X2 _AES_ENC_u0_u2_U423  ( .A1(_AES_ENC_w3[1] ), .A2(_AES_ENC_u0_u2_n620 ), .ZN(_AES_ENC_u0_u2_n667 ) );
NAND2_X2 _AES_ENC_u0_u2_U422  ( .A1(_AES_ENC_u0_u2_n619 ), .A2(_AES_ENC_u0_u2_n667 ), .ZN(_AES_ENC_u0_u2_n1071 ) );
NAND4_X2 _AES_ENC_u0_u2_U412  ( .A1(_AES_ENC_u0_u2_n675 ), .A2(_AES_ENC_u0_u2_n674 ), .A3(_AES_ENC_u0_u2_n673 ), .A4(_AES_ENC_u0_u2_n672 ), .ZN(_AES_ENC_u0_u2_n676 ) );
NAND2_X2 _AES_ENC_u0_u2_U411  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n676 ), .ZN(_AES_ENC_u0_u2_n677 ) );
NAND2_X2 _AES_ENC_u0_u2_U408  ( .A1(_AES_ENC_u0_u2_n800 ), .A2(_AES_ENC_u0_u2_n1022 ), .ZN(_AES_ENC_u0_u2_n680 ) );
NAND2_X2 _AES_ENC_u0_u2_U407  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n680 ), .ZN(_AES_ENC_u0_u2_n681 ) );
AND2_X2 _AES_ENC_u0_u2_U402  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n684 ), .ZN(_AES_ENC_u0_u2_n682 ) );
NAND4_X2 _AES_ENC_u0_u2_U395  ( .A1(_AES_ENC_u0_u2_n691 ), .A2(_AES_ENC_u0_u2_n581 ), .A3(_AES_ENC_u0_u2_n690 ), .A4(_AES_ENC_u0_u2_n689 ), .ZN(_AES_ENC_u0_u2_n692 ) );
NAND2_X2 _AES_ENC_u0_u2_U394  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n692 ), .ZN(_AES_ENC_u0_u2_n733 ) );
NAND2_X2 _AES_ENC_u0_u2_U392  ( .A1(_AES_ENC_u0_u2_n977 ), .A2(_AES_ENC_u0_u2_n1050 ), .ZN(_AES_ENC_u0_u2_n702 ) );
NAND2_X2 _AES_ENC_u0_u2_U391  ( .A1(_AES_ENC_u0_u2_n1093 ), .A2(_AES_ENC_u0_u2_n1045 ), .ZN(_AES_ENC_u0_u2_n701 ) );
NAND4_X2 _AES_ENC_u0_u2_U381  ( .A1(_AES_ENC_u0_u2_n702 ), .A2(_AES_ENC_u0_u2_n701 ), .A3(_AES_ENC_u0_u2_n700 ), .A4(_AES_ENC_u0_u2_n699 ), .ZN(_AES_ENC_u0_u2_n703 ) );
NAND2_X2 _AES_ENC_u0_u2_U380  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n703 ), .ZN(_AES_ENC_u0_u2_n732 ) );
AND2_X2 _AES_ENC_u0_u2_U379  ( .A1(_AES_ENC_w3[0] ), .A2(_AES_ENC_w3[6] ),.ZN(_AES_ENC_u0_u2_n1113 ) );
NAND2_X2 _AES_ENC_u0_u2_U378  ( .A1(_AES_ENC_u0_u2_n601 ), .A2(_AES_ENC_u0_u2_n1030 ), .ZN(_AES_ENC_u0_u2_n881 ) );
NAND2_X2 _AES_ENC_u0_u2_U377  ( .A1(_AES_ENC_u0_u2_n1093 ), .A2(_AES_ENC_u0_u2_n881 ), .ZN(_AES_ENC_u0_u2_n715 ) );
NAND2_X2 _AES_ENC_u0_u2_U376  ( .A1(_AES_ENC_u0_u2_n1010 ), .A2(_AES_ENC_u0_u2_n600 ), .ZN(_AES_ENC_u0_u2_n714 ) );
NAND2_X2 _AES_ENC_u0_u2_U375  ( .A1(_AES_ENC_u0_u2_n855 ), .A2(_AES_ENC_u0_u2_n588 ), .ZN(_AES_ENC_u0_u2_n1117 ) );
XNOR2_X2 _AES_ENC_u0_u2_U371  ( .A(_AES_ENC_u0_u2_n611 ), .B(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n824 ) );
NAND4_X2 _AES_ENC_u0_u2_U362  ( .A1(_AES_ENC_u0_u2_n715 ), .A2(_AES_ENC_u0_u2_n714 ), .A3(_AES_ENC_u0_u2_n713 ), .A4(_AES_ENC_u0_u2_n712 ), .ZN(_AES_ENC_u0_u2_n716 ) );
NAND2_X2 _AES_ENC_u0_u2_U361  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n716 ), .ZN(_AES_ENC_u0_u2_n731 ) );
AND2_X2 _AES_ENC_u0_u2_U360  ( .A1(_AES_ENC_w3[6] ), .A2(_AES_ENC_u0_u2_n574 ), .ZN(_AES_ENC_u0_u2_n1131 ) );
NAND2_X2 _AES_ENC_u0_u2_U359  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n717 ) );
NAND2_X2 _AES_ENC_u0_u2_U358  ( .A1(_AES_ENC_u0_u2_n1029 ), .A2(_AES_ENC_u0_u2_n717 ), .ZN(_AES_ENC_u0_u2_n728 ) );
NAND2_X2 _AES_ENC_u0_u2_U357  ( .A1(_AES_ENC_w3[1] ), .A2(_AES_ENC_u0_u2_n624 ), .ZN(_AES_ENC_u0_u2_n1097 ) );
NAND2_X2 _AES_ENC_u0_u2_U356  ( .A1(_AES_ENC_u0_u2_n603 ), .A2(_AES_ENC_u0_u2_n1097 ), .ZN(_AES_ENC_u0_u2_n718 ) );
NAND2_X2 _AES_ENC_u0_u2_U355  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n718 ), .ZN(_AES_ENC_u0_u2_n727 ) );
NAND4_X2 _AES_ENC_u0_u2_U344  ( .A1(_AES_ENC_u0_u2_n728 ), .A2(_AES_ENC_u0_u2_n727 ), .A3(_AES_ENC_u0_u2_n726 ), .A4(_AES_ENC_u0_u2_n725 ), .ZN(_AES_ENC_u0_u2_n729 ) );
NAND2_X2 _AES_ENC_u0_u2_U343  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n729 ), .ZN(_AES_ENC_u0_u2_n730 ) );
NAND4_X2 _AES_ENC_u0_u2_U342  ( .A1(_AES_ENC_u0_u2_n733 ), .A2(_AES_ENC_u0_u2_n732 ), .A3(_AES_ENC_u0_u2_n731 ), .A4(_AES_ENC_u0_u2_n730 ), .ZN(_AES_ENC_u0_subword[9] ) );
NAND2_X2 _AES_ENC_u0_u2_U341  ( .A1(_AES_ENC_w3[7] ), .A2(_AES_ENC_u0_u2_n611 ), .ZN(_AES_ENC_u0_u2_n734 ) );
NAND2_X2 _AES_ENC_u0_u2_U340  ( .A1(_AES_ENC_u0_u2_n734 ), .A2(_AES_ENC_u0_u2_n607 ), .ZN(_AES_ENC_u0_u2_n738 ) );
OR4_X2 _AES_ENC_u0_u2_U339  ( .A1(_AES_ENC_u0_u2_n738 ), .A2(_AES_ENC_u0_u2_n626 ), .A3(_AES_ENC_u0_u2_n826 ), .A4(_AES_ENC_u0_u2_n1121 ), .ZN(_AES_ENC_u0_u2_n746 ) );
NAND2_X2 _AES_ENC_u0_u2_U337  ( .A1(_AES_ENC_u0_u2_n1100 ), .A2(_AES_ENC_u0_u2_n587 ), .ZN(_AES_ENC_u0_u2_n992 ) );
OR2_X2 _AES_ENC_u0_u2_U336  ( .A1(_AES_ENC_u0_u2_n610 ), .A2(_AES_ENC_u0_u2_n735 ), .ZN(_AES_ENC_u0_u2_n737 ) );
NAND2_X2 _AES_ENC_u0_u2_U334  ( .A1(_AES_ENC_u0_u2_n619 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n753 ) );
NAND2_X2 _AES_ENC_u0_u2_U333  ( .A1(_AES_ENC_u0_u2_n582 ), .A2(_AES_ENC_u0_u2_n753 ), .ZN(_AES_ENC_u0_u2_n1080 ) );
NAND2_X2 _AES_ENC_u0_u2_U332  ( .A1(_AES_ENC_u0_u2_n1048 ), .A2(_AES_ENC_u0_u2_n576 ), .ZN(_AES_ENC_u0_u2_n736 ) );
NAND2_X2 _AES_ENC_u0_u2_U331  ( .A1(_AES_ENC_u0_u2_n737 ), .A2(_AES_ENC_u0_u2_n736 ), .ZN(_AES_ENC_u0_u2_n739 ) );
NAND2_X2 _AES_ENC_u0_u2_U330  ( .A1(_AES_ENC_u0_u2_n739 ), .A2(_AES_ENC_u0_u2_n738 ), .ZN(_AES_ENC_u0_u2_n745 ) );
NAND2_X2 _AES_ENC_u0_u2_U326  ( .A1(_AES_ENC_u0_u2_n1096 ), .A2(_AES_ENC_u0_u2_n590 ), .ZN(_AES_ENC_u0_u2_n906 ) );
NAND4_X2 _AES_ENC_u0_u2_U323  ( .A1(_AES_ENC_u0_u2_n746 ), .A2(_AES_ENC_u0_u2_n992 ), .A3(_AES_ENC_u0_u2_n745 ), .A4(_AES_ENC_u0_u2_n744 ), .ZN(_AES_ENC_u0_u2_n747 ) );
NAND2_X2 _AES_ENC_u0_u2_U322  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n747 ), .ZN(_AES_ENC_u0_u2_n793 ) );
NAND2_X2 _AES_ENC_u0_u2_U321  ( .A1(_AES_ENC_u0_u2_n584 ), .A2(_AES_ENC_u0_u2_n855 ), .ZN(_AES_ENC_u0_u2_n748 ) );
NAND2_X2 _AES_ENC_u0_u2_U320  ( .A1(_AES_ENC_u0_u2_n956 ), .A2(_AES_ENC_u0_u2_n748 ), .ZN(_AES_ENC_u0_u2_n760 ) );
NAND2_X2 _AES_ENC_u0_u2_U313  ( .A1(_AES_ENC_u0_u2_n590 ), .A2(_AES_ENC_u0_u2_n753 ), .ZN(_AES_ENC_u0_u2_n1023 ) );
NAND4_X2 _AES_ENC_u0_u2_U308  ( .A1(_AES_ENC_u0_u2_n760 ), .A2(_AES_ENC_u0_u2_n992 ), .A3(_AES_ENC_u0_u2_n759 ), .A4(_AES_ENC_u0_u2_n758 ), .ZN(_AES_ENC_u0_u2_n761 ) );
NAND2_X2 _AES_ENC_u0_u2_U307  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n761 ), .ZN(_AES_ENC_u0_u2_n792 ) );
NAND2_X2 _AES_ENC_u0_u2_U306  ( .A1(_AES_ENC_u0_u2_n584 ), .A2(_AES_ENC_u0_u2_n603 ), .ZN(_AES_ENC_u0_u2_n989 ) );
NAND2_X2 _AES_ENC_u0_u2_U305  ( .A1(_AES_ENC_u0_u2_n1050 ), .A2(_AES_ENC_u0_u2_n989 ), .ZN(_AES_ENC_u0_u2_n777 ) );
NAND2_X2 _AES_ENC_u0_u2_U304  ( .A1(_AES_ENC_u0_u2_n1093 ), .A2(_AES_ENC_u0_u2_n762 ), .ZN(_AES_ENC_u0_u2_n776 ) );
XNOR2_X2 _AES_ENC_u0_u2_U301  ( .A(_AES_ENC_w3[7] ), .B(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n959 ) );
NAND4_X2 _AES_ENC_u0_u2_U289  ( .A1(_AES_ENC_u0_u2_n777 ), .A2(_AES_ENC_u0_u2_n776 ), .A3(_AES_ENC_u0_u2_n775 ), .A4(_AES_ENC_u0_u2_n774 ), .ZN(_AES_ENC_u0_u2_n778 ) );
NAND2_X2 _AES_ENC_u0_u2_U288  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n778 ), .ZN(_AES_ENC_u0_u2_n791 ) );
NAND2_X2 _AES_ENC_u0_u2_U287  ( .A1(_AES_ENC_u0_u2_n1056 ), .A2(_AES_ENC_u0_u2_n1050 ), .ZN(_AES_ENC_u0_u2_n788 ) );
NAND2_X2 _AES_ENC_u0_u2_U286  ( .A1(_AES_ENC_u0_u2_n1091 ), .A2(_AES_ENC_u0_u2_n779 ), .ZN(_AES_ENC_u0_u2_n787 ) );
NAND2_X2 _AES_ENC_u0_u2_U285  ( .A1(_AES_ENC_u0_u2_n956 ), .A2(_AES_ENC_w3[1] ), .ZN(_AES_ENC_u0_u2_n786 ) );
NAND4_X2 _AES_ENC_u0_u2_U278  ( .A1(_AES_ENC_u0_u2_n788 ), .A2(_AES_ENC_u0_u2_n787 ), .A3(_AES_ENC_u0_u2_n786 ), .A4(_AES_ENC_u0_u2_n785 ), .ZN(_AES_ENC_u0_u2_n789 ) );
NAND2_X2 _AES_ENC_u0_u2_U277  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n789 ), .ZN(_AES_ENC_u0_u2_n790 ) );
NAND4_X2 _AES_ENC_u0_u2_U276  ( .A1(_AES_ENC_u0_u2_n793 ), .A2(_AES_ENC_u0_u2_n792 ), .A3(_AES_ENC_u0_u2_n791 ), .A4(_AES_ENC_u0_u2_n790 ), .ZN(_AES_ENC_u0_subword[10] ) );
NAND2_X2 _AES_ENC_u0_u2_U275  ( .A1(_AES_ENC_u0_u2_n1059 ), .A2(_AES_ENC_u0_u2_n794 ), .ZN(_AES_ENC_u0_u2_n810 ) );
NAND2_X2 _AES_ENC_u0_u2_U274  ( .A1(_AES_ENC_u0_u2_n1049 ), .A2(_AES_ENC_u0_u2_n956 ), .ZN(_AES_ENC_u0_u2_n809 ) );
OR2_X2 _AES_ENC_u0_u2_U266  ( .A1(_AES_ENC_u0_u2_n1096 ), .A2(_AES_ENC_u0_u2_n606 ), .ZN(_AES_ENC_u0_u2_n802 ) );
NAND2_X2 _AES_ENC_u0_u2_U265  ( .A1(_AES_ENC_u0_u2_n1053 ), .A2(_AES_ENC_u0_u2_n800 ), .ZN(_AES_ENC_u0_u2_n801 ) );
NAND2_X2 _AES_ENC_u0_u2_U264  ( .A1(_AES_ENC_u0_u2_n802 ), .A2(_AES_ENC_u0_u2_n801 ), .ZN(_AES_ENC_u0_u2_n805 ) );
NAND4_X2 _AES_ENC_u0_u2_U261  ( .A1(_AES_ENC_u0_u2_n810 ), .A2(_AES_ENC_u0_u2_n809 ), .A3(_AES_ENC_u0_u2_n808 ), .A4(_AES_ENC_u0_u2_n807 ), .ZN(_AES_ENC_u0_u2_n811 ) );
NAND2_X2 _AES_ENC_u0_u2_U260  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n811 ), .ZN(_AES_ENC_u0_u2_n852 ) );
OR2_X2 _AES_ENC_u0_u2_U259  ( .A1(_AES_ENC_u0_u2_n1023 ), .A2(_AES_ENC_u0_u2_n617 ), .ZN(_AES_ENC_u0_u2_n819 ) );
OR2_X2 _AES_ENC_u0_u2_U257  ( .A1(_AES_ENC_u0_u2_n570 ), .A2(_AES_ENC_u0_u2_n930 ), .ZN(_AES_ENC_u0_u2_n818 ) );
NAND2_X2 _AES_ENC_u0_u2_U256  ( .A1(_AES_ENC_u0_u2_n1013 ), .A2(_AES_ENC_u0_u2_n1094 ), .ZN(_AES_ENC_u0_u2_n817 ) );
NAND4_X2 _AES_ENC_u0_u2_U249  ( .A1(_AES_ENC_u0_u2_n819 ), .A2(_AES_ENC_u0_u2_n818 ), .A3(_AES_ENC_u0_u2_n817 ), .A4(_AES_ENC_u0_u2_n816 ), .ZN(_AES_ENC_u0_u2_n820 ) );
NAND2_X2 _AES_ENC_u0_u2_U248  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n820 ), .ZN(_AES_ENC_u0_u2_n851 ) );
NAND2_X2 _AES_ENC_u0_u2_U247  ( .A1(_AES_ENC_u0_u2_n956 ), .A2(_AES_ENC_u0_u2_n1080 ), .ZN(_AES_ENC_u0_u2_n835 ) );
NAND2_X2 _AES_ENC_u0_u2_U246  ( .A1(_AES_ENC_u0_u2_n570 ), .A2(_AES_ENC_u0_u2_n1030 ), .ZN(_AES_ENC_u0_u2_n1047 ) );
OR2_X2 _AES_ENC_u0_u2_U245  ( .A1(_AES_ENC_u0_u2_n1047 ), .A2(_AES_ENC_u0_u2_n612 ), .ZN(_AES_ENC_u0_u2_n834 ) );
NAND2_X2 _AES_ENC_u0_u2_U244  ( .A1(_AES_ENC_u0_u2_n1072 ), .A2(_AES_ENC_u0_u2_n589 ), .ZN(_AES_ENC_u0_u2_n833 ) );
NAND4_X2 _AES_ENC_u0_u2_U233  ( .A1(_AES_ENC_u0_u2_n835 ), .A2(_AES_ENC_u0_u2_n834 ), .A3(_AES_ENC_u0_u2_n833 ), .A4(_AES_ENC_u0_u2_n832 ), .ZN(_AES_ENC_u0_u2_n836 ) );
NAND2_X2 _AES_ENC_u0_u2_U232  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n836 ), .ZN(_AES_ENC_u0_u2_n850 ) );
NAND2_X2 _AES_ENC_u0_u2_U231  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n623 ), .ZN(_AES_ENC_u0_u2_n847 ) );
NAND2_X2 _AES_ENC_u0_u2_U230  ( .A1(_AES_ENC_u0_u2_n1050 ), .A2(_AES_ENC_u0_u2_n1071 ), .ZN(_AES_ENC_u0_u2_n846 ) );
OR2_X2 _AES_ENC_u0_u2_U224  ( .A1(_AES_ENC_u0_u2_n1053 ), .A2(_AES_ENC_u0_u2_n911 ), .ZN(_AES_ENC_u0_u2_n1077 ) );
NAND4_X2 _AES_ENC_u0_u2_U220  ( .A1(_AES_ENC_u0_u2_n847 ), .A2(_AES_ENC_u0_u2_n846 ), .A3(_AES_ENC_u0_u2_n845 ), .A4(_AES_ENC_u0_u2_n844 ), .ZN(_AES_ENC_u0_u2_n848 ) );
NAND2_X2 _AES_ENC_u0_u2_U219  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n848 ), .ZN(_AES_ENC_u0_u2_n849 ) );
NAND4_X2 _AES_ENC_u0_u2_U218  ( .A1(_AES_ENC_u0_u2_n852 ), .A2(_AES_ENC_u0_u2_n851 ), .A3(_AES_ENC_u0_u2_n850 ), .A4(_AES_ENC_u0_u2_n849 ), .ZN(_AES_ENC_u0_subword[11] ) );
NAND2_X2 _AES_ENC_u0_u2_U216  ( .A1(_AES_ENC_u0_u2_n1009 ), .A2(_AES_ENC_u0_u2_n1072 ), .ZN(_AES_ENC_u0_u2_n862 ) );
NAND2_X2 _AES_ENC_u0_u2_U215  ( .A1(_AES_ENC_u0_u2_n603 ), .A2(_AES_ENC_u0_u2_n577 ), .ZN(_AES_ENC_u0_u2_n853 ) );
NAND2_X2 _AES_ENC_u0_u2_U214  ( .A1(_AES_ENC_u0_u2_n1050 ), .A2(_AES_ENC_u0_u2_n853 ), .ZN(_AES_ENC_u0_u2_n861 ) );
NAND4_X2 _AES_ENC_u0_u2_U206  ( .A1(_AES_ENC_u0_u2_n862 ), .A2(_AES_ENC_u0_u2_n861 ), .A3(_AES_ENC_u0_u2_n860 ), .A4(_AES_ENC_u0_u2_n859 ), .ZN(_AES_ENC_u0_u2_n863 ) );
NAND2_X2 _AES_ENC_u0_u2_U205  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n863 ), .ZN(_AES_ENC_u0_u2_n905 ) );
NAND2_X2 _AES_ENC_u0_u2_U204  ( .A1(_AES_ENC_u0_u2_n1010 ), .A2(_AES_ENC_u0_u2_n989 ), .ZN(_AES_ENC_u0_u2_n874 ) );
NAND2_X2 _AES_ENC_u0_u2_U203  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n610 ), .ZN(_AES_ENC_u0_u2_n864 ) );
NAND2_X2 _AES_ENC_u0_u2_U202  ( .A1(_AES_ENC_u0_u2_n929 ), .A2(_AES_ENC_u0_u2_n864 ), .ZN(_AES_ENC_u0_u2_n873 ) );
NAND4_X2 _AES_ENC_u0_u2_U193  ( .A1(_AES_ENC_u0_u2_n874 ), .A2(_AES_ENC_u0_u2_n873 ), .A3(_AES_ENC_u0_u2_n872 ), .A4(_AES_ENC_u0_u2_n871 ), .ZN(_AES_ENC_u0_u2_n875 ) );
NAND2_X2 _AES_ENC_u0_u2_U192  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n875 ), .ZN(_AES_ENC_u0_u2_n904 ) );
NAND2_X2 _AES_ENC_u0_u2_U191  ( .A1(_AES_ENC_u0_u2_n583 ), .A2(_AES_ENC_u0_u2_n1050 ), .ZN(_AES_ENC_u0_u2_n889 ) );
NAND2_X2 _AES_ENC_u0_u2_U190  ( .A1(_AES_ENC_u0_u2_n1093 ), .A2(_AES_ENC_u0_u2_n587 ), .ZN(_AES_ENC_u0_u2_n876 ) );
NAND2_X2 _AES_ENC_u0_u2_U189  ( .A1(_AES_ENC_u0_u2_n604 ), .A2(_AES_ENC_u0_u2_n876 ), .ZN(_AES_ENC_u0_u2_n877 ) );
NAND2_X2 _AES_ENC_u0_u2_U188  ( .A1(_AES_ENC_u0_u2_n877 ), .A2(_AES_ENC_u0_u2_n623 ), .ZN(_AES_ENC_u0_u2_n888 ) );
NAND4_X2 _AES_ENC_u0_u2_U179  ( .A1(_AES_ENC_u0_u2_n889 ), .A2(_AES_ENC_u0_u2_n888 ), .A3(_AES_ENC_u0_u2_n887 ), .A4(_AES_ENC_u0_u2_n886 ), .ZN(_AES_ENC_u0_u2_n890 ) );
NAND2_X2 _AES_ENC_u0_u2_U178  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n890 ), .ZN(_AES_ENC_u0_u2_n903 ) );
OR2_X2 _AES_ENC_u0_u2_U177  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n1059 ), .ZN(_AES_ENC_u0_u2_n900 ) );
NAND2_X2 _AES_ENC_u0_u2_U176  ( .A1(_AES_ENC_u0_u2_n1073 ), .A2(_AES_ENC_u0_u2_n1047 ), .ZN(_AES_ENC_u0_u2_n899 ) );
NAND2_X2 _AES_ENC_u0_u2_U175  ( .A1(_AES_ENC_u0_u2_n1094 ), .A2(_AES_ENC_u0_u2_n595 ), .ZN(_AES_ENC_u0_u2_n898 ) );
NAND4_X2 _AES_ENC_u0_u2_U167  ( .A1(_AES_ENC_u0_u2_n900 ), .A2(_AES_ENC_u0_u2_n899 ), .A3(_AES_ENC_u0_u2_n898 ), .A4(_AES_ENC_u0_u2_n897 ), .ZN(_AES_ENC_u0_u2_n901 ) );
NAND2_X2 _AES_ENC_u0_u2_U166  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n901 ), .ZN(_AES_ENC_u0_u2_n902 ) );
NAND4_X2 _AES_ENC_u0_u2_U165  ( .A1(_AES_ENC_u0_u2_n905 ), .A2(_AES_ENC_u0_u2_n904 ), .A3(_AES_ENC_u0_u2_n903 ), .A4(_AES_ENC_u0_u2_n902 ), .ZN(_AES_ENC_u0_subword[12] ) );
NAND2_X2 _AES_ENC_u0_u2_U164  ( .A1(_AES_ENC_u0_u2_n1094 ), .A2(_AES_ENC_u0_u2_n599 ), .ZN(_AES_ENC_u0_u2_n922 ) );
NAND2_X2 _AES_ENC_u0_u2_U163  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n989 ), .ZN(_AES_ENC_u0_u2_n921 ) );
NAND4_X2 _AES_ENC_u0_u2_U151  ( .A1(_AES_ENC_u0_u2_n922 ), .A2(_AES_ENC_u0_u2_n921 ), .A3(_AES_ENC_u0_u2_n920 ), .A4(_AES_ENC_u0_u2_n919 ), .ZN(_AES_ENC_u0_u2_n923 ) );
NAND2_X2 _AES_ENC_u0_u2_U150  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n923 ), .ZN(_AES_ENC_u0_u2_n972 ) );
NAND2_X2 _AES_ENC_u0_u2_U149  ( .A1(_AES_ENC_u0_u2_n582 ), .A2(_AES_ENC_u0_u2_n619 ), .ZN(_AES_ENC_u0_u2_n924 ) );
NAND2_X2 _AES_ENC_u0_u2_U148  ( .A1(_AES_ENC_u0_u2_n1073 ), .A2(_AES_ENC_u0_u2_n924 ), .ZN(_AES_ENC_u0_u2_n939 ) );
NAND2_X2 _AES_ENC_u0_u2_U147  ( .A1(_AES_ENC_u0_u2_n926 ), .A2(_AES_ENC_u0_u2_n925 ), .ZN(_AES_ENC_u0_u2_n927 ) );
NAND2_X2 _AES_ENC_u0_u2_U146  ( .A1(_AES_ENC_u0_u2_n606 ), .A2(_AES_ENC_u0_u2_n927 ), .ZN(_AES_ENC_u0_u2_n928 ) );
NAND2_X2 _AES_ENC_u0_u2_U145  ( .A1(_AES_ENC_u0_u2_n928 ), .A2(_AES_ENC_u0_u2_n1080 ), .ZN(_AES_ENC_u0_u2_n938 ) );
OR2_X2 _AES_ENC_u0_u2_U144  ( .A1(_AES_ENC_u0_u2_n1117 ), .A2(_AES_ENC_u0_u2_n615 ), .ZN(_AES_ENC_u0_u2_n937 ) );
NAND4_X2 _AES_ENC_u0_u2_U139  ( .A1(_AES_ENC_u0_u2_n939 ), .A2(_AES_ENC_u0_u2_n938 ), .A3(_AES_ENC_u0_u2_n937 ), .A4(_AES_ENC_u0_u2_n936 ), .ZN(_AES_ENC_u0_u2_n940 ) );
NAND2_X2 _AES_ENC_u0_u2_U138  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n940 ), .ZN(_AES_ENC_u0_u2_n971 ) );
OR2_X2 _AES_ENC_u0_u2_U137  ( .A1(_AES_ENC_u0_u2_n605 ), .A2(_AES_ENC_u0_u2_n941 ), .ZN(_AES_ENC_u0_u2_n954 ) );
NAND2_X2 _AES_ENC_u0_u2_U136  ( .A1(_AES_ENC_u0_u2_n1096 ), .A2(_AES_ENC_u0_u2_n577 ), .ZN(_AES_ENC_u0_u2_n942 ) );
NAND2_X2 _AES_ENC_u0_u2_U135  ( .A1(_AES_ENC_u0_u2_n1048 ), .A2(_AES_ENC_u0_u2_n942 ), .ZN(_AES_ENC_u0_u2_n943 ) );
NAND2_X2 _AES_ENC_u0_u2_U134  ( .A1(_AES_ENC_u0_u2_n612 ), .A2(_AES_ENC_u0_u2_n943 ), .ZN(_AES_ENC_u0_u2_n944 ) );
NAND2_X2 _AES_ENC_u0_u2_U133  ( .A1(_AES_ENC_u0_u2_n944 ), .A2(_AES_ENC_u0_u2_n580 ), .ZN(_AES_ENC_u0_u2_n953 ) );
NAND4_X2 _AES_ENC_u0_u2_U125  ( .A1(_AES_ENC_u0_u2_n954 ), .A2(_AES_ENC_u0_u2_n953 ), .A3(_AES_ENC_u0_u2_n952 ), .A4(_AES_ENC_u0_u2_n951 ), .ZN(_AES_ENC_u0_u2_n955 ) );
NAND2_X2 _AES_ENC_u0_u2_U124  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n955 ), .ZN(_AES_ENC_u0_u2_n970 ) );
NAND2_X2 _AES_ENC_u0_u2_U123  ( .A1(_AES_ENC_u0_u2_n1094 ), .A2(_AES_ENC_u0_u2_n1071 ), .ZN(_AES_ENC_u0_u2_n967 ) );
NAND2_X2 _AES_ENC_u0_u2_U122  ( .A1(_AES_ENC_u0_u2_n956 ), .A2(_AES_ENC_u0_u2_n1030 ), .ZN(_AES_ENC_u0_u2_n966 ) );
NAND4_X2 _AES_ENC_u0_u2_U114  ( .A1(_AES_ENC_u0_u2_n967 ), .A2(_AES_ENC_u0_u2_n966 ), .A3(_AES_ENC_u0_u2_n965 ), .A4(_AES_ENC_u0_u2_n964 ), .ZN(_AES_ENC_u0_u2_n968 ) );
NAND2_X2 _AES_ENC_u0_u2_U113  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n968 ), .ZN(_AES_ENC_u0_u2_n969 ) );
NAND4_X2 _AES_ENC_u0_u2_U112  ( .A1(_AES_ENC_u0_u2_n972 ), .A2(_AES_ENC_u0_u2_n971 ), .A3(_AES_ENC_u0_u2_n970 ), .A4(_AES_ENC_u0_u2_n969 ), .ZN(_AES_ENC_u0_subword[13] ) );
NAND2_X2 _AES_ENC_u0_u2_U111  ( .A1(_AES_ENC_u0_u2_n570 ), .A2(_AES_ENC_u0_u2_n1097 ), .ZN(_AES_ENC_u0_u2_n973 ) );
NAND2_X2 _AES_ENC_u0_u2_U110  ( .A1(_AES_ENC_u0_u2_n1073 ), .A2(_AES_ENC_u0_u2_n973 ), .ZN(_AES_ENC_u0_u2_n987 ) );
NAND2_X2 _AES_ENC_u0_u2_U109  ( .A1(_AES_ENC_u0_u2_n974 ), .A2(_AES_ENC_u0_u2_n1077 ), .ZN(_AES_ENC_u0_u2_n975 ) );
NAND2_X2 _AES_ENC_u0_u2_U108  ( .A1(_AES_ENC_u0_u2_n613 ), .A2(_AES_ENC_u0_u2_n975 ), .ZN(_AES_ENC_u0_u2_n976 ) );
NAND2_X2 _AES_ENC_u0_u2_U107  ( .A1(_AES_ENC_u0_u2_n977 ), .A2(_AES_ENC_u0_u2_n976 ), .ZN(_AES_ENC_u0_u2_n986 ) );
NAND4_X2 _AES_ENC_u0_u2_U99  ( .A1(_AES_ENC_u0_u2_n987 ), .A2(_AES_ENC_u0_u2_n986 ), .A3(_AES_ENC_u0_u2_n985 ), .A4(_AES_ENC_u0_u2_n984 ), .ZN(_AES_ENC_u0_u2_n988 ) );
NAND2_X2 _AES_ENC_u0_u2_U98  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n988 ), .ZN(_AES_ENC_u0_u2_n1044 ) );
NAND2_X2 _AES_ENC_u0_u2_U97  ( .A1(_AES_ENC_u0_u2_n1073 ), .A2(_AES_ENC_u0_u2_n989 ), .ZN(_AES_ENC_u0_u2_n1004 ) );
NAND2_X2 _AES_ENC_u0_u2_U96  ( .A1(_AES_ENC_u0_u2_n1092 ), .A2(_AES_ENC_u0_u2_n619 ), .ZN(_AES_ENC_u0_u2_n1003 ) );
NAND4_X2 _AES_ENC_u0_u2_U85  ( .A1(_AES_ENC_u0_u2_n1004 ), .A2(_AES_ENC_u0_u2_n1003 ), .A3(_AES_ENC_u0_u2_n1002 ), .A4(_AES_ENC_u0_u2_n1001 ), .ZN(_AES_ENC_u0_u2_n1005 ) );
NAND2_X2 _AES_ENC_u0_u2_U84  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n1005 ), .ZN(_AES_ENC_u0_u2_n1043 ) );
NAND2_X2 _AES_ENC_u0_u2_U83  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n596 ), .ZN(_AES_ENC_u0_u2_n1020 ) );
NAND2_X2 _AES_ENC_u0_u2_U82  ( .A1(_AES_ENC_u0_u2_n1050 ), .A2(_AES_ENC_u0_u2_n624 ), .ZN(_AES_ENC_u0_u2_n1019 ) );
NAND2_X2 _AES_ENC_u0_u2_U77  ( .A1(_AES_ENC_u0_u2_n1059 ), .A2(_AES_ENC_u0_u2_n1114 ), .ZN(_AES_ENC_u0_u2_n1012 ) );
NAND2_X2 _AES_ENC_u0_u2_U76  ( .A1(_AES_ENC_u0_u2_n1010 ), .A2(_AES_ENC_u0_u2_n592 ), .ZN(_AES_ENC_u0_u2_n1011 ) );
NAND2_X2 _AES_ENC_u0_u2_U75  ( .A1(_AES_ENC_u0_u2_n1012 ), .A2(_AES_ENC_u0_u2_n1011 ), .ZN(_AES_ENC_u0_u2_n1016 ) );
NAND4_X2 _AES_ENC_u0_u2_U70  ( .A1(_AES_ENC_u0_u2_n1020 ), .A2(_AES_ENC_u0_u2_n1019 ), .A3(_AES_ENC_u0_u2_n1018 ), .A4(_AES_ENC_u0_u2_n1017 ), .ZN(_AES_ENC_u0_u2_n1021 ) );
NAND2_X2 _AES_ENC_u0_u2_U69  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n1021 ), .ZN(_AES_ENC_u0_u2_n1042 ) );
NAND2_X2 _AES_ENC_u0_u2_U68  ( .A1(_AES_ENC_u0_u2_n1022 ), .A2(_AES_ENC_u0_u2_n1093 ), .ZN(_AES_ENC_u0_u2_n1039 ) );
NAND2_X2 _AES_ENC_u0_u2_U67  ( .A1(_AES_ENC_u0_u2_n1050 ), .A2(_AES_ENC_u0_u2_n1023 ), .ZN(_AES_ENC_u0_u2_n1038 ) );
NAND2_X2 _AES_ENC_u0_u2_U66  ( .A1(_AES_ENC_u0_u2_n1024 ), .A2(_AES_ENC_u0_u2_n1071 ), .ZN(_AES_ENC_u0_u2_n1037 ) );
AND2_X2 _AES_ENC_u0_u2_U60  ( .A1(_AES_ENC_u0_u2_n1030 ), .A2(_AES_ENC_u0_u2_n602 ), .ZN(_AES_ENC_u0_u2_n1078 ) );
NAND4_X2 _AES_ENC_u0_u2_U56  ( .A1(_AES_ENC_u0_u2_n1039 ), .A2(_AES_ENC_u0_u2_n1038 ), .A3(_AES_ENC_u0_u2_n1037 ), .A4(_AES_ENC_u0_u2_n1036 ), .ZN(_AES_ENC_u0_u2_n1040 ) );
NAND2_X2 _AES_ENC_u0_u2_U55  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n1040 ), .ZN(_AES_ENC_u0_u2_n1041 ) );
NAND4_X2 _AES_ENC_u0_u2_U54  ( .A1(_AES_ENC_u0_u2_n1044 ), .A2(_AES_ENC_u0_u2_n1043 ), .A3(_AES_ENC_u0_u2_n1042 ), .A4(_AES_ENC_u0_u2_n1041 ), .ZN(_AES_ENC_u0_subword[14] ) );
NAND2_X2 _AES_ENC_u0_u2_U53  ( .A1(_AES_ENC_u0_u2_n1072 ), .A2(_AES_ENC_u0_u2_n1045 ), .ZN(_AES_ENC_u0_u2_n1068 ) );
NAND2_X2 _AES_ENC_u0_u2_U52  ( .A1(_AES_ENC_u0_u2_n1046 ), .A2(_AES_ENC_u0_u2_n582 ), .ZN(_AES_ENC_u0_u2_n1067 ) );
NAND2_X2 _AES_ENC_u0_u2_U51  ( .A1(_AES_ENC_u0_u2_n1094 ), .A2(_AES_ENC_u0_u2_n1047 ), .ZN(_AES_ENC_u0_u2_n1066 ) );
NAND4_X2 _AES_ENC_u0_u2_U40  ( .A1(_AES_ENC_u0_u2_n1068 ), .A2(_AES_ENC_u0_u2_n1067 ), .A3(_AES_ENC_u0_u2_n1066 ), .A4(_AES_ENC_u0_u2_n1065 ), .ZN(_AES_ENC_u0_u2_n1069 ) );
NAND2_X2 _AES_ENC_u0_u2_U39  ( .A1(_AES_ENC_u0_u2_n1070 ), .A2(_AES_ENC_u0_u2_n1069 ), .ZN(_AES_ENC_u0_u2_n1135 ) );
NAND2_X2 _AES_ENC_u0_u2_U38  ( .A1(_AES_ENC_u0_u2_n1072 ), .A2(_AES_ENC_u0_u2_n1071 ), .ZN(_AES_ENC_u0_u2_n1088 ) );
NAND2_X2 _AES_ENC_u0_u2_U37  ( .A1(_AES_ENC_u0_u2_n1073 ), .A2(_AES_ENC_u0_u2_n595 ), .ZN(_AES_ENC_u0_u2_n1087 ) );
NAND4_X2 _AES_ENC_u0_u2_U28  ( .A1(_AES_ENC_u0_u2_n1088 ), .A2(_AES_ENC_u0_u2_n1087 ), .A3(_AES_ENC_u0_u2_n1086 ), .A4(_AES_ENC_u0_u2_n1085 ), .ZN(_AES_ENC_u0_u2_n1089 ) );
NAND2_X2 _AES_ENC_u0_u2_U27  ( .A1(_AES_ENC_u0_u2_n1090 ), .A2(_AES_ENC_u0_u2_n1089 ), .ZN(_AES_ENC_u0_u2_n1134 ) );
NAND2_X2 _AES_ENC_u0_u2_U26  ( .A1(_AES_ENC_u0_u2_n1091 ), .A2(_AES_ENC_u0_u2_n1093 ), .ZN(_AES_ENC_u0_u2_n1111 ) );
NAND2_X2 _AES_ENC_u0_u2_U25  ( .A1(_AES_ENC_u0_u2_n1092 ), .A2(_AES_ENC_u0_u2_n1120 ), .ZN(_AES_ENC_u0_u2_n1110 ) );
AND2_X2 _AES_ENC_u0_u2_U22  ( .A1(_AES_ENC_u0_u2_n1097 ), .A2(_AES_ENC_u0_u2_n1096 ), .ZN(_AES_ENC_u0_u2_n1098 ) );
NAND4_X2 _AES_ENC_u0_u2_U14  ( .A1(_AES_ENC_u0_u2_n1111 ), .A2(_AES_ENC_u0_u2_n1110 ), .A3(_AES_ENC_u0_u2_n1109 ), .A4(_AES_ENC_u0_u2_n1108 ), .ZN(_AES_ENC_u0_u2_n1112 ) );
NAND2_X2 _AES_ENC_u0_u2_U13  ( .A1(_AES_ENC_u0_u2_n1113 ), .A2(_AES_ENC_u0_u2_n1112 ), .ZN(_AES_ENC_u0_u2_n1133 ) );
NAND2_X2 _AES_ENC_u0_u2_U12  ( .A1(_AES_ENC_u0_u2_n1115 ), .A2(_AES_ENC_u0_u2_n1114 ), .ZN(_AES_ENC_u0_u2_n1129 ) );
OR2_X2 _AES_ENC_u0_u2_U11  ( .A1(_AES_ENC_u0_u2_n608 ), .A2(_AES_ENC_u0_u2_n1116 ), .ZN(_AES_ENC_u0_u2_n1128 ) );
NAND4_X2 _AES_ENC_u0_u2_U3  ( .A1(_AES_ENC_u0_u2_n1129 ), .A2(_AES_ENC_u0_u2_n1128 ), .A3(_AES_ENC_u0_u2_n1127 ), .A4(_AES_ENC_u0_u2_n1126 ), .ZN(_AES_ENC_u0_u2_n1130 ) );
NAND2_X2 _AES_ENC_u0_u2_U2  ( .A1(_AES_ENC_u0_u2_n1131 ), .A2(_AES_ENC_u0_u2_n1130 ), .ZN(_AES_ENC_u0_u2_n1132 ) );
NAND4_X2 _AES_ENC_u0_u2_U1  ( .A1(_AES_ENC_u0_u2_n1135 ), .A2(_AES_ENC_u0_u2_n1134 ), .A3(_AES_ENC_u0_u2_n1133 ), .A4(_AES_ENC_u0_u2_n1132 ), .ZN(_AES_ENC_u0_subword[15] ) );
INV_X4 _AES_ENC_u0_u3_U575  ( .A(_AES_ENC_w3[31] ), .ZN(_AES_ENC_u0_u3_n627 ) );
INV_X4 _AES_ENC_u0_u3_U574  ( .A(_AES_ENC_u0_u3_n1114 ), .ZN(_AES_ENC_u0_u3_n625 ) );
INV_X4 _AES_ENC_u0_u3_U573  ( .A(_AES_ENC_w3[28] ), .ZN(_AES_ENC_u0_u3_n624 ) );
INV_X4 _AES_ENC_u0_u3_U572  ( .A(_AES_ENC_u0_u3_n1025 ), .ZN(_AES_ENC_u0_u3_n622 ) );
INV_X4 _AES_ENC_u0_u3_U571  ( .A(_AES_ENC_u0_u3_n1120 ), .ZN(_AES_ENC_u0_u3_n620 ) );
INV_X4 _AES_ENC_u0_u3_U570  ( .A(_AES_ENC_u0_u3_n1121 ), .ZN(_AES_ENC_u0_u3_n619 ) );
INV_X4 _AES_ENC_u0_u3_U569  ( .A(_AES_ENC_u0_u3_n1048 ), .ZN(_AES_ENC_u0_u3_n618 ) );
INV_X4 _AES_ENC_u0_u3_U568  ( .A(_AES_ENC_u0_u3_n974 ), .ZN(_AES_ENC_u0_u3_n616 ) );
INV_X4 _AES_ENC_u0_u3_U567  ( .A(_AES_ENC_u0_u3_n794 ), .ZN(_AES_ENC_u0_u3_n614 ) );
INV_X4 _AES_ENC_u0_u3_U566  ( .A(_AES_ENC_w3[26] ), .ZN(_AES_ENC_u0_u3_n611 ) );
INV_X4 _AES_ENC_u0_u3_U565  ( .A(_AES_ENC_u0_u3_n800 ), .ZN(_AES_ENC_u0_u3_n610 ) );
INV_X4 _AES_ENC_u0_u3_U564  ( .A(_AES_ENC_u0_u3_n925 ), .ZN(_AES_ENC_u0_u3_n609 ) );
INV_X4 _AES_ENC_u0_u3_U563  ( .A(_AES_ENC_u0_u3_n779 ), .ZN(_AES_ENC_u0_u3_n607 ) );
INV_X4 _AES_ENC_u0_u3_U562  ( .A(_AES_ENC_u0_u3_n1022 ), .ZN(_AES_ENC_u0_u3_n603 ) );
INV_X4 _AES_ENC_u0_u3_U561  ( .A(_AES_ENC_u0_u3_n1102 ), .ZN(_AES_ENC_u0_u3_n602 ) );
INV_X4 _AES_ENC_u0_u3_U560  ( .A(_AES_ENC_u0_u3_n929 ), .ZN(_AES_ENC_u0_u3_n601 ) );
INV_X4 _AES_ENC_u0_u3_U559  ( .A(_AES_ENC_u0_u3_n1056 ), .ZN(_AES_ENC_u0_u3_n600 ) );
INV_X4 _AES_ENC_u0_u3_U558  ( .A(_AES_ENC_u0_u3_n1054 ), .ZN(_AES_ENC_u0_u3_n599 ) );
INV_X4 _AES_ENC_u0_u3_U557  ( .A(_AES_ENC_u0_u3_n881 ), .ZN(_AES_ENC_u0_u3_n598 ) );
INV_X4 _AES_ENC_u0_u3_U556  ( .A(_AES_ENC_u0_u3_n926 ), .ZN(_AES_ENC_u0_u3_n597 ) );
INV_X4 _AES_ENC_u0_u3_U555  ( .A(_AES_ENC_u0_u3_n977 ), .ZN(_AES_ENC_u0_u3_n595 ) );
INV_X4 _AES_ENC_u0_u3_U554  ( .A(_AES_ENC_u0_u3_n1031 ), .ZN(_AES_ENC_u0_u3_n594 ) );
INV_X4 _AES_ENC_u0_u3_U553  ( .A(_AES_ENC_u0_u3_n1103 ), .ZN(_AES_ENC_u0_u3_n593 ) );
INV_X4 _AES_ENC_u0_u3_U552  ( .A(_AES_ENC_u0_u3_n1009 ), .ZN(_AES_ENC_u0_u3_n592 ) );
INV_X4 _AES_ENC_u0_u3_U551  ( .A(_AES_ENC_u0_u3_n990 ), .ZN(_AES_ENC_u0_u3_n591 ) );
INV_X4 _AES_ENC_u0_u3_U550  ( .A(_AES_ENC_u0_u3_n1058 ), .ZN(_AES_ENC_u0_u3_n590 ) );
INV_X4 _AES_ENC_u0_u3_U549  ( .A(_AES_ENC_u0_u3_n1074 ), .ZN(_AES_ENC_u0_u3_n589 ) );
INV_X4 _AES_ENC_u0_u3_U548  ( .A(_AES_ENC_u0_u3_n1053 ), .ZN(_AES_ENC_u0_u3_n588 ) );
INV_X4 _AES_ENC_u0_u3_U547  ( .A(_AES_ENC_u0_u3_n826 ), .ZN(_AES_ENC_u0_u3_n587 ) );
INV_X4 _AES_ENC_u0_u3_U546  ( .A(_AES_ENC_u0_u3_n992 ), .ZN(_AES_ENC_u0_u3_n586 ) );
INV_X4 _AES_ENC_u0_u3_U545  ( .A(_AES_ENC_u0_u3_n821 ), .ZN(_AES_ENC_u0_u3_n585 ) );
INV_X4 _AES_ENC_u0_u3_U544  ( .A(_AES_ENC_u0_u3_n910 ), .ZN(_AES_ENC_u0_u3_n584 ) );
INV_X4 _AES_ENC_u0_u3_U543  ( .A(_AES_ENC_u0_u3_n906 ), .ZN(_AES_ENC_u0_u3_n583 ) );
INV_X4 _AES_ENC_u0_u3_U542  ( .A(_AES_ENC_u0_u3_n880 ), .ZN(_AES_ENC_u0_u3_n581 ) );
INV_X4 _AES_ENC_u0_u3_U541  ( .A(_AES_ENC_u0_u3_n1013 ), .ZN(_AES_ENC_u0_u3_n580 ) );
INV_X4 _AES_ENC_u0_u3_U540  ( .A(_AES_ENC_u0_u3_n1092 ), .ZN(_AES_ENC_u0_u3_n579 ) );
INV_X4 _AES_ENC_u0_u3_U539  ( .A(_AES_ENC_u0_u3_n824 ), .ZN(_AES_ENC_u0_u3_n578 ) );
INV_X4 _AES_ENC_u0_u3_U538  ( .A(_AES_ENC_u0_u3_n1091 ), .ZN(_AES_ENC_u0_u3_n577 ) );
INV_X4 _AES_ENC_u0_u3_U537  ( .A(_AES_ENC_u0_u3_n1080 ), .ZN(_AES_ENC_u0_u3_n576 ) );
INV_X4 _AES_ENC_u0_u3_U536  ( .A(_AES_ENC_u0_u3_n959 ), .ZN(_AES_ENC_u0_u3_n575 ) );
INV_X4 _AES_ENC_u0_u3_U535  ( .A(_AES_ENC_w3[24] ), .ZN(_AES_ENC_u0_u3_n574 ) );
NOR2_X2 _AES_ENC_u0_u3_U534  ( .A1(_AES_ENC_u0_u3_n574 ), .A2(_AES_ENC_w3[30] ), .ZN(_AES_ENC_u0_u3_n1070 ) );
NOR2_X2 _AES_ENC_u0_u3_U533  ( .A1(_AES_ENC_w3[24] ), .A2(_AES_ENC_w3[30] ),.ZN(_AES_ENC_u0_u3_n1090 ) );
NOR2_X2 _AES_ENC_u0_u3_U532  ( .A1(_AES_ENC_w3[28] ), .A2(_AES_ENC_w3[27] ),.ZN(_AES_ENC_u0_u3_n1025 ) );
NAND3_X2 _AES_ENC_u0_u3_U531  ( .A1(_AES_ENC_u0_u3_n679 ), .A2(_AES_ENC_u0_u3_n678 ), .A3(_AES_ENC_u0_u3_n677 ), .ZN(_AES_ENC_u0_subword[0] ) );
NOR2_X2 _AES_ENC_u0_u3_U530  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n765 ) );
NOR2_X2 _AES_ENC_u0_u3_U529  ( .A1(_AES_ENC_w3[28] ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n764 ) );
NOR2_X2 _AES_ENC_u0_u3_U528  ( .A1(_AES_ENC_u0_u3_n765 ), .A2(_AES_ENC_u0_u3_n764 ), .ZN(_AES_ENC_u0_u3_n766 ) );
NOR2_X2 _AES_ENC_u0_u3_U527  ( .A1(_AES_ENC_u0_u3_n766 ), .A2(_AES_ENC_u0_u3_n575 ), .ZN(_AES_ENC_u0_u3_n767 ) );
NOR2_X2 _AES_ENC_u0_u3_U526  ( .A1(_AES_ENC_u0_u3_n1117 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n707 ) );
NOR3_X2 _AES_ENC_u0_u3_U525  ( .A1(_AES_ENC_u0_u3_n627 ), .A2(_AES_ENC_w3[29] ), .A3(_AES_ENC_u0_u3_n704 ), .ZN(_AES_ENC_u0_u3_n706 ) );
NOR2_X2 _AES_ENC_u0_u3_U524  ( .A1(_AES_ENC_w3[28] ), .A2(_AES_ENC_u0_u3_n579 ), .ZN(_AES_ENC_u0_u3_n705 ) );
NOR3_X2 _AES_ENC_u0_u3_U523  ( .A1(_AES_ENC_u0_u3_n707 ), .A2(_AES_ENC_u0_u3_n706 ), .A3(_AES_ENC_u0_u3_n705 ), .ZN(_AES_ENC_u0_u3_n713 ) );
NOR4_X2 _AES_ENC_u0_u3_U522  ( .A1(_AES_ENC_u0_u3_n633 ), .A2(_AES_ENC_u0_u3_n632 ), .A3(_AES_ENC_u0_u3_n631 ), .A4(_AES_ENC_u0_u3_n630 ), .ZN(_AES_ENC_u0_u3_n634 ) );
NOR2_X2 _AES_ENC_u0_u3_U521  ( .A1(_AES_ENC_u0_u3_n629 ), .A2(_AES_ENC_u0_u3_n628 ), .ZN(_AES_ENC_u0_u3_n635 ) );
NAND3_X2 _AES_ENC_u0_u3_U520  ( .A1(_AES_ENC_w3[26] ), .A2(_AES_ENC_w3[31] ),.A3(_AES_ENC_u0_u3_n1059 ), .ZN(_AES_ENC_u0_u3_n636 ) );
INV_X4 _AES_ENC_u0_u3_U519  ( .A(_AES_ENC_w3[27] ), .ZN(_AES_ENC_u0_u3_n621 ) );
NOR2_X2 _AES_ENC_u0_u3_U518  ( .A1(_AES_ENC_w3[29] ), .A2(_AES_ENC_w3[26] ),.ZN(_AES_ENC_u0_u3_n974 ) );
NAND3_X2 _AES_ENC_u0_u3_U517  ( .A1(_AES_ENC_u0_u3_n652 ), .A2(_AES_ENC_u0_u3_n626 ), .A3(_AES_ENC_w3[31] ), .ZN(_AES_ENC_u0_u3_n653 ) );
NOR2_X2 _AES_ENC_u0_u3_U516  ( .A1(_AES_ENC_u0_u3_n611 ), .A2(_AES_ENC_w3[29] ), .ZN(_AES_ENC_u0_u3_n925 ) );
NOR2_X2 _AES_ENC_u0_u3_U515  ( .A1(_AES_ENC_u0_u3_n626 ), .A2(_AES_ENC_w3[26] ), .ZN(_AES_ENC_u0_u3_n1048 ) );
INV_X4 _AES_ENC_u0_u3_U512  ( .A(_AES_ENC_w3[29] ), .ZN(_AES_ENC_u0_u3_n626 ) );
NOR2_X2 _AES_ENC_u0_u3_U510  ( .A1(_AES_ENC_u0_u3_n611 ), .A2(_AES_ENC_w3[31] ), .ZN(_AES_ENC_u0_u3_n779 ) );
NOR2_X2 _AES_ENC_u0_u3_U509  ( .A1(_AES_ENC_w3[31] ), .A2(_AES_ENC_w3[26] ),.ZN(_AES_ENC_u0_u3_n794 ) );
NOR2_X2 _AES_ENC_u0_u3_U508  ( .A1(_AES_ENC_w3[28] ), .A2(_AES_ENC_w3[25] ),.ZN(_AES_ENC_u0_u3_n1102 ) );
INV_X4 _AES_ENC_u0_u3_U507  ( .A(_AES_ENC_u0_u3_n569 ), .ZN(_AES_ENC_u0_u3_n572 ) );
NOR2_X2 _AES_ENC_u0_u3_U506  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_w3[27] ), .ZN(_AES_ENC_u0_u3_n1053 ) );
NOR2_X2 _AES_ENC_u0_u3_U505  ( .A1(_AES_ENC_u0_u3_n607 ), .A2(_AES_ENC_w3[29] ), .ZN(_AES_ENC_u0_u3_n1024 ) );
NOR2_X2 _AES_ENC_u0_u3_U504  ( .A1(_AES_ENC_u0_u3_n625 ), .A2(_AES_ENC_w3[26] ), .ZN(_AES_ENC_u0_u3_n1093 ) );
NOR2_X2 _AES_ENC_u0_u3_U503  ( .A1(_AES_ENC_u0_u3_n614 ), .A2(_AES_ENC_w3[29] ), .ZN(_AES_ENC_u0_u3_n1094 ) );
NOR2_X2 _AES_ENC_u0_u3_U502  ( .A1(_AES_ENC_u0_u3_n624 ), .A2(_AES_ENC_w3[27] ), .ZN(_AES_ENC_u0_u3_n931 ) );
INV_X4 _AES_ENC_u0_u3_U501  ( .A(_AES_ENC_u0_u3_n570 ), .ZN(_AES_ENC_u0_u3_n573 ) );
NOR2_X2 _AES_ENC_u0_u3_U500  ( .A1(_AES_ENC_u0_u3_n622 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n1059 ) );
NOR2_X2 _AES_ENC_u0_u3_U499  ( .A1(_AES_ENC_u0_u3_n1053 ), .A2(_AES_ENC_u0_u3_n1095 ), .ZN(_AES_ENC_u0_u3_n639 ) );
NOR3_X2 _AES_ENC_u0_u3_U498  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n573 ), .A3(_AES_ENC_u0_u3_n1074 ), .ZN(_AES_ENC_u0_u3_n641 ) );
NOR2_X2 _AES_ENC_u0_u3_U497  ( .A1(_AES_ENC_u0_u3_n639 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n640 ) );
NOR2_X2 _AES_ENC_u0_u3_U496  ( .A1(_AES_ENC_u0_u3_n641 ), .A2(_AES_ENC_u0_u3_n640 ), .ZN(_AES_ENC_u0_u3_n646 ) );
NOR2_X2 _AES_ENC_u0_u3_U495  ( .A1(_AES_ENC_u0_u3_n826 ), .A2(_AES_ENC_u0_u3_n572 ), .ZN(_AES_ENC_u0_u3_n827 ) );
NOR3_X2 _AES_ENC_u0_u3_U494  ( .A1(_AES_ENC_u0_u3_n769 ), .A2(_AES_ENC_u0_u3_n768 ), .A3(_AES_ENC_u0_u3_n767 ), .ZN(_AES_ENC_u0_u3_n775 ) );
NOR2_X2 _AES_ENC_u0_u3_U492  ( .A1(_AES_ENC_w3[25] ), .A2(_AES_ENC_u0_u3_n623 ), .ZN(_AES_ENC_u0_u3_n913 ) );
NOR2_X2 _AES_ENC_u0_u3_U491  ( .A1(_AES_ENC_u0_u3_n913 ), .A2(_AES_ENC_u0_u3_n1091 ), .ZN(_AES_ENC_u0_u3_n914 ) );
NOR2_X2 _AES_ENC_u0_u3_U490  ( .A1(_AES_ENC_u0_u3_n1056 ), .A2(_AES_ENC_u0_u3_n1053 ), .ZN(_AES_ENC_u0_u3_n749 ) );
NOR2_X2 _AES_ENC_u0_u3_U489  ( .A1(_AES_ENC_u0_u3_n749 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n752 ) );
NOR3_X2 _AES_ENC_u0_u3_U488  ( .A1(_AES_ENC_u0_u3_n995 ), .A2(_AES_ENC_u0_u3_n586 ), .A3(_AES_ENC_u0_u3_n994 ), .ZN(_AES_ENC_u0_u3_n1002 ) );
NOR2_X2 _AES_ENC_u0_u3_U487  ( .A1(_AES_ENC_u0_u3_n909 ), .A2(_AES_ENC_u0_u3_n908 ), .ZN(_AES_ENC_u0_u3_n920 ) );
INV_X4 _AES_ENC_u0_u3_U486  ( .A(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n596 ) );
NOR2_X2 _AES_ENC_u0_u3_U483  ( .A1(_AES_ENC_u0_u3_n932 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n933 ) );
NOR2_X2 _AES_ENC_u0_u3_U482  ( .A1(_AES_ENC_u0_u3_n929 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n935 ) );
NOR2_X2 _AES_ENC_u0_u3_U480  ( .A1(_AES_ENC_u0_u3_n931 ), .A2(_AES_ENC_u0_u3_n930 ), .ZN(_AES_ENC_u0_u3_n934 ) );
NOR3_X2 _AES_ENC_u0_u3_U479  ( .A1(_AES_ENC_u0_u3_n935 ), .A2(_AES_ENC_u0_u3_n934 ), .A3(_AES_ENC_u0_u3_n933 ), .ZN(_AES_ENC_u0_u3_n936 ) );
OR2_X4 _AES_ENC_u0_u3_U478  ( .A1(_AES_ENC_u0_u3_n1094 ), .A2(_AES_ENC_u0_u3_n1093 ), .ZN(_AES_ENC_u0_u3_n571 ) );
AND2_X2 _AES_ENC_u0_u3_U477  ( .A1(_AES_ENC_u0_u3_n571 ), .A2(_AES_ENC_u0_u3_n1095 ), .ZN(_AES_ENC_u0_u3_n1101 ) );
NOR2_X2 _AES_ENC_u0_u3_U474  ( .A1(_AES_ENC_u0_u3_n1074 ), .A2(_AES_ENC_u0_u3_n931 ), .ZN(_AES_ENC_u0_u3_n796 ) );
NOR2_X2 _AES_ENC_u0_u3_U473  ( .A1(_AES_ENC_u0_u3_n796 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n797 ) );
NOR2_X2 _AES_ENC_u0_u3_U472  ( .A1(_AES_ENC_u0_u3_n1054 ), .A2(_AES_ENC_u0_u3_n1053 ), .ZN(_AES_ENC_u0_u3_n1055 ) );
NOR2_X2 _AES_ENC_u0_u3_U471  ( .A1(_AES_ENC_u0_u3_n572 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n949 ) );
NOR2_X2 _AES_ENC_u0_u3_U470  ( .A1(_AES_ENC_u0_u3_n1049 ), .A2(_AES_ENC_u0_u3_n618 ), .ZN(_AES_ENC_u0_u3_n1051 ) );
NOR2_X2 _AES_ENC_u0_u3_U469  ( .A1(_AES_ENC_u0_u3_n1051 ), .A2(_AES_ENC_u0_u3_n1050 ), .ZN(_AES_ENC_u0_u3_n1052 ) );
NOR2_X2 _AES_ENC_u0_u3_U468  ( .A1(_AES_ENC_u0_u3_n1052 ), .A2(_AES_ENC_u0_u3_n592 ), .ZN(_AES_ENC_u0_u3_n1064 ) );
NOR2_X2 _AES_ENC_u0_u3_U467  ( .A1(_AES_ENC_w3[25] ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n631 ) );
NOR2_X2 _AES_ENC_u0_u3_U466  ( .A1(_AES_ENC_u0_u3_n1025 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n980 ) );
NOR2_X2 _AES_ENC_u0_u3_U465  ( .A1(_AES_ENC_u0_u3_n1074 ), .A2(_AES_ENC_u0_u3_n1025 ), .ZN(_AES_ENC_u0_u3_n891 ) );
NOR2_X2 _AES_ENC_u0_u3_U464  ( .A1(_AES_ENC_u0_u3_n891 ), .A2(_AES_ENC_u0_u3_n609 ), .ZN(_AES_ENC_u0_u3_n894 ) );
NOR2_X2 _AES_ENC_u0_u3_U463  ( .A1(_AES_ENC_u0_u3_n1073 ), .A2(_AES_ENC_u0_u3_n1094 ), .ZN(_AES_ENC_u0_u3_n795 ) );
NOR2_X2 _AES_ENC_u0_u3_U462  ( .A1(_AES_ENC_u0_u3_n795 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n799 ) );
NOR2_X2 _AES_ENC_u0_u3_U461  ( .A1(_AES_ENC_u0_u3_n624 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n1075 ) );
NOR2_X2 _AES_ENC_u0_u3_U460  ( .A1(_AES_ENC_u0_u3_n624 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n822 ) );
NOR2_X2 _AES_ENC_u0_u3_U459  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n823 ) );
NOR2_X2 _AES_ENC_u0_u3_U458  ( .A1(_AES_ENC_u0_u3_n823 ), .A2(_AES_ENC_u0_u3_n822 ), .ZN(_AES_ENC_u0_u3_n825 ) );
NOR2_X2 _AES_ENC_u0_u3_U455  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n981 ) );
NOR2_X2 _AES_ENC_u0_u3_U448  ( .A1(_AES_ENC_u0_u3_n1102 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n643 ) );
NOR2_X2 _AES_ENC_u0_u3_U447  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n621 ), .ZN(_AES_ENC_u0_u3_n642 ) );
NOR2_X2 _AES_ENC_u0_u3_U442  ( .A1(_AES_ENC_u0_u3_n911 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n644 ) );
NOR4_X2 _AES_ENC_u0_u3_U441  ( .A1(_AES_ENC_u0_u3_n644 ), .A2(_AES_ENC_u0_u3_n643 ), .A3(_AES_ENC_u0_u3_n804 ), .A4(_AES_ENC_u0_u3_n642 ), .ZN(_AES_ENC_u0_u3_n645 ) );
NOR2_X2 _AES_ENC_u0_u3_U438  ( .A1(_AES_ENC_u0_u3_n1102 ), .A2(_AES_ENC_u0_u3_n910 ), .ZN(_AES_ENC_u0_u3_n932 ) );
NOR3_X2 _AES_ENC_u0_u3_U435  ( .A1(_AES_ENC_u0_u3_n623 ), .A2(_AES_ENC_w3[25] ), .A3(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n683 ) );
NOR2_X2 _AES_ENC_u0_u3_U434  ( .A1(_AES_ENC_u0_u3_n1102 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n755 ) );
INV_X4 _AES_ENC_u0_u3_U433  ( .A(_AES_ENC_u0_u3_n931 ), .ZN(_AES_ENC_u0_u3_n623 ) );
NOR2_X2 _AES_ENC_u0_u3_U428  ( .A1(_AES_ENC_u0_u3_n996 ), .A2(_AES_ENC_u0_u3_n931 ), .ZN(_AES_ENC_u0_u3_n704 ) );
NOR2_X2 _AES_ENC_u0_u3_U427  ( .A1(_AES_ENC_u0_u3_n1029 ), .A2(_AES_ENC_u0_u3_n1025 ), .ZN(_AES_ENC_u0_u3_n1079 ) );
NOR3_X2 _AES_ENC_u0_u3_U421  ( .A1(_AES_ENC_u0_u3_n589 ), .A2(_AES_ENC_u0_u3_n1025 ), .A3(_AES_ENC_u0_u3_n616 ), .ZN(_AES_ENC_u0_u3_n945 ) );
NOR2_X2 _AES_ENC_u0_u3_U420  ( .A1(_AES_ENC_u0_u3_n1072 ), .A2(_AES_ENC_u0_u3_n1094 ), .ZN(_AES_ENC_u0_u3_n930 ) );
NOR2_X2 _AES_ENC_u0_u3_U419  ( .A1(_AES_ENC_u0_u3_n931 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n743 ) );
NOR2_X2 _AES_ENC_u0_u3_U418  ( .A1(_AES_ENC_u0_u3_n931 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n685 ) );
NOR3_X2 _AES_ENC_u0_u3_U417  ( .A1(_AES_ENC_u0_u3_n610 ), .A2(_AES_ENC_u0_u3_n572 ), .A3(_AES_ENC_u0_u3_n575 ), .ZN(_AES_ENC_u0_u3_n962 ) );
NOR2_X2 _AES_ENC_u0_u3_U416  ( .A1(_AES_ENC_u0_u3_n626 ), .A2(_AES_ENC_u0_u3_n611 ), .ZN(_AES_ENC_u0_u3_n800 ) );
NOR3_X2 _AES_ENC_u0_u3_U415  ( .A1(_AES_ENC_u0_u3_n590 ), .A2(_AES_ENC_u0_u3_n627 ), .A3(_AES_ENC_u0_u3_n611 ), .ZN(_AES_ENC_u0_u3_n798 ) );
NOR3_X2 _AES_ENC_u0_u3_U414  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n572 ), .A3(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n694 ) );
NOR3_X2 _AES_ENC_u0_u3_U413  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n572 ), .A3(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n895 ) );
NOR3_X2 _AES_ENC_u0_u3_U410  ( .A1(_AES_ENC_u0_u3_n1008 ), .A2(_AES_ENC_u0_u3_n1007 ), .A3(_AES_ENC_u0_u3_n1006 ), .ZN(_AES_ENC_u0_u3_n1018 ) );
NOR4_X2 _AES_ENC_u0_u3_U409  ( .A1(_AES_ENC_u0_u3_n711 ), .A2(_AES_ENC_u0_u3_n710 ), .A3(_AES_ENC_u0_u3_n709 ), .A4(_AES_ENC_u0_u3_n708 ), .ZN(_AES_ENC_u0_u3_n712 ) );
NOR4_X2 _AES_ENC_u0_u3_U406  ( .A1(_AES_ENC_u0_u3_n806 ), .A2(_AES_ENC_u0_u3_n805 ), .A3(_AES_ENC_u0_u3_n804 ), .A4(_AES_ENC_u0_u3_n803 ), .ZN(_AES_ENC_u0_u3_n807 ) );
NOR3_X2 _AES_ENC_u0_u3_U405  ( .A1(_AES_ENC_u0_u3_n799 ), .A2(_AES_ENC_u0_u3_n798 ), .A3(_AES_ENC_u0_u3_n797 ), .ZN(_AES_ENC_u0_u3_n808 ) );
NOR2_X2 _AES_ENC_u0_u3_U404  ( .A1(_AES_ENC_u0_u3_n669 ), .A2(_AES_ENC_u0_u3_n668 ), .ZN(_AES_ENC_u0_u3_n673 ) );
NOR4_X2 _AES_ENC_u0_u3_U403  ( .A1(_AES_ENC_u0_u3_n946 ), .A2(_AES_ENC_u0_u3_n1046 ), .A3(_AES_ENC_u0_u3_n671 ), .A4(_AES_ENC_u0_u3_n670 ), .ZN(_AES_ENC_u0_u3_n672 ) );
NOR4_X2 _AES_ENC_u0_u3_U401  ( .A1(_AES_ENC_u0_u3_n843 ), .A2(_AES_ENC_u0_u3_n842 ), .A3(_AES_ENC_u0_u3_n841 ), .A4(_AES_ENC_u0_u3_n840 ), .ZN(_AES_ENC_u0_u3_n844 ) );
NOR3_X2 _AES_ENC_u0_u3_U400  ( .A1(_AES_ENC_u0_u3_n1101 ), .A2(_AES_ENC_u0_u3_n1100 ), .A3(_AES_ENC_u0_u3_n1099 ), .ZN(_AES_ENC_u0_u3_n1109 ) );
NOR3_X2 _AES_ENC_u0_u3_U399  ( .A1(_AES_ENC_u0_u3_n743 ), .A2(_AES_ENC_u0_u3_n742 ), .A3(_AES_ENC_u0_u3_n741 ), .ZN(_AES_ENC_u0_u3_n744 ) );
NOR2_X2 _AES_ENC_u0_u3_U398  ( .A1(_AES_ENC_u0_u3_n697 ), .A2(_AES_ENC_u0_u3_n658 ), .ZN(_AES_ENC_u0_u3_n659 ) );
NOR3_X2 _AES_ENC_u0_u3_U397  ( .A1(_AES_ENC_u0_u3_n959 ), .A2(_AES_ENC_u0_u3_n572 ), .A3(_AES_ENC_u0_u3_n609 ), .ZN(_AES_ENC_u0_u3_n768 ) );
NOR2_X2 _AES_ENC_u0_u3_U396  ( .A1(_AES_ENC_u0_u3_n1078 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n1033 ) );
NOR2_X2 _AES_ENC_u0_u3_U393  ( .A1(_AES_ENC_u0_u3_n1031 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n1032 ) );
NOR3_X2 _AES_ENC_u0_u3_U390  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n1025 ), .A3(_AES_ENC_u0_u3_n1074 ), .ZN(_AES_ENC_u0_u3_n1035 ) );
NOR4_X2 _AES_ENC_u0_u3_U389  ( .A1(_AES_ENC_u0_u3_n1035 ), .A2(_AES_ENC_u0_u3_n1034 ), .A3(_AES_ENC_u0_u3_n1033 ), .A4(_AES_ENC_u0_u3_n1032 ), .ZN(_AES_ENC_u0_u3_n1036 ) );
NOR2_X2 _AES_ENC_u0_u3_U388  ( .A1(_AES_ENC_u0_u3_n598 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n885 ) );
NOR2_X2 _AES_ENC_u0_u3_U387  ( .A1(_AES_ENC_u0_u3_n623 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n882 ) );
NOR2_X2 _AES_ENC_u0_u3_U386  ( .A1(_AES_ENC_u0_u3_n1053 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n884 ) );
NOR4_X2 _AES_ENC_u0_u3_U385  ( .A1(_AES_ENC_u0_u3_n885 ), .A2(_AES_ENC_u0_u3_n884 ), .A3(_AES_ENC_u0_u3_n883 ), .A4(_AES_ENC_u0_u3_n882 ), .ZN(_AES_ENC_u0_u3_n886 ) );
NOR2_X2 _AES_ENC_u0_u3_U384  ( .A1(_AES_ENC_u0_u3_n825 ), .A2(_AES_ENC_u0_u3_n578 ), .ZN(_AES_ENC_u0_u3_n830 ) );
NOR2_X2 _AES_ENC_u0_u3_U383  ( .A1(_AES_ENC_u0_u3_n827 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n829 ) );
NOR2_X2 _AES_ENC_u0_u3_U382  ( .A1(_AES_ENC_u0_u3_n572 ), .A2(_AES_ENC_u0_u3_n579 ), .ZN(_AES_ENC_u0_u3_n828 ) );
NOR4_X2 _AES_ENC_u0_u3_U374  ( .A1(_AES_ENC_u0_u3_n831 ), .A2(_AES_ENC_u0_u3_n830 ), .A3(_AES_ENC_u0_u3_n829 ), .A4(_AES_ENC_u0_u3_n828 ), .ZN(_AES_ENC_u0_u3_n832 ) );
NOR2_X2 _AES_ENC_u0_u3_U373  ( .A1(_AES_ENC_u0_u3_n598 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n1107 ) );
NOR2_X2 _AES_ENC_u0_u3_U372  ( .A1(_AES_ENC_u0_u3_n1102 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n1106 ) );
NOR2_X2 _AES_ENC_u0_u3_U370  ( .A1(_AES_ENC_u0_u3_n1103 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n1105 ) );
NOR4_X2 _AES_ENC_u0_u3_U369  ( .A1(_AES_ENC_u0_u3_n1107 ), .A2(_AES_ENC_u0_u3_n1106 ), .A3(_AES_ENC_u0_u3_n1105 ), .A4(_AES_ENC_u0_u3_n1104 ), .ZN(_AES_ENC_u0_u3_n1108 ) );
NOR3_X2 _AES_ENC_u0_u3_U368  ( .A1(_AES_ENC_u0_u3_n959 ), .A2(_AES_ENC_u0_u3_n621 ), .A3(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n963 ) );
NOR2_X2 _AES_ENC_u0_u3_U367  ( .A1(_AES_ENC_u0_u3_n626 ), .A2(_AES_ENC_u0_u3_n627 ), .ZN(_AES_ENC_u0_u3_n1114 ) );
NOR3_X2 _AES_ENC_u0_u3_U366  ( .A1(_AES_ENC_u0_u3_n910 ), .A2(_AES_ENC_u0_u3_n1059 ), .A3(_AES_ENC_u0_u3_n611 ), .ZN(_AES_ENC_u0_u3_n1115 ) );
INV_X4 _AES_ENC_u0_u3_U365  ( .A(_AES_ENC_u0_u3_n1024 ), .ZN(_AES_ENC_u0_u3_n606 ) );
INV_X4 _AES_ENC_u0_u3_U364  ( .A(_AES_ENC_u0_u3_n1094 ), .ZN(_AES_ENC_u0_u3_n613 ) );
NOR2_X2 _AES_ENC_u0_u3_U363  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n931 ), .ZN(_AES_ENC_u0_u3_n1100 ) );
NOR2_X2 _AES_ENC_u0_u3_U354  ( .A1(_AES_ENC_u0_u3_n569 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n929 ) );
NOR2_X2 _AES_ENC_u0_u3_U353  ( .A1(_AES_ENC_u0_u3_n620 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n926 ) );
INV_X4 _AES_ENC_u0_u3_U352  ( .A(_AES_ENC_u0_u3_n1093 ), .ZN(_AES_ENC_u0_u3_n617 ) );
NOR2_X2 _AES_ENC_u0_u3_U351  ( .A1(_AES_ENC_u0_u3_n572 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n1095 ) );
NOR2_X2 _AES_ENC_u0_u3_U350  ( .A1(_AES_ENC_u0_u3_n609 ), .A2(_AES_ENC_u0_u3_n627 ), .ZN(_AES_ENC_u0_u3_n1010 ) );
NOR2_X2 _AES_ENC_u0_u3_U349  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n1103 ) );
NOR2_X2 _AES_ENC_u0_u3_U348  ( .A1(_AES_ENC_w3[25] ), .A2(_AES_ENC_u0_u3_n1120 ), .ZN(_AES_ENC_u0_u3_n1022 ) );
NOR2_X2 _AES_ENC_u0_u3_U347  ( .A1(_AES_ENC_u0_u3_n619 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n911 ) );
NOR2_X2 _AES_ENC_u0_u3_U346  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_u0_u3_n1025 ), .ZN(_AES_ENC_u0_u3_n826 ) );
NOR2_X2 _AES_ENC_u0_u3_U345  ( .A1(_AES_ENC_u0_u3_n626 ), .A2(_AES_ENC_u0_u3_n607 ), .ZN(_AES_ENC_u0_u3_n1072 ) );
NOR2_X2 _AES_ENC_u0_u3_U338  ( .A1(_AES_ENC_u0_u3_n627 ), .A2(_AES_ENC_u0_u3_n616 ), .ZN(_AES_ENC_u0_u3_n956 ) );
NOR2_X2 _AES_ENC_u0_u3_U335  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_u0_u3_n624 ), .ZN(_AES_ENC_u0_u3_n1121 ) );
NOR2_X2 _AES_ENC_u0_u3_U329  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_u0_u3_n624 ), .ZN(_AES_ENC_u0_u3_n1058 ) );
NOR2_X2 _AES_ENC_u0_u3_U328  ( .A1(_AES_ENC_u0_u3_n625 ), .A2(_AES_ENC_u0_u3_n611 ), .ZN(_AES_ENC_u0_u3_n1073 ) );
NOR2_X2 _AES_ENC_u0_u3_U327  ( .A1(_AES_ENC_w3[25] ), .A2(_AES_ENC_u0_u3_n1025 ), .ZN(_AES_ENC_u0_u3_n1054 ) );
NOR2_X2 _AES_ENC_u0_u3_U325  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_u0_u3_n931 ), .ZN(_AES_ENC_u0_u3_n1029 ) );
NOR2_X2 _AES_ENC_u0_u3_U324  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n1056 ) );
NOR2_X2 _AES_ENC_u0_u3_U319  ( .A1(_AES_ENC_u0_u3_n614 ), .A2(_AES_ENC_u0_u3_n626 ), .ZN(_AES_ENC_u0_u3_n1050 ) );
NOR2_X2 _AES_ENC_u0_u3_U318  ( .A1(_AES_ENC_u0_u3_n1121 ), .A2(_AES_ENC_u0_u3_n1025 ), .ZN(_AES_ENC_u0_u3_n1120 ) );
NOR2_X2 _AES_ENC_u0_u3_U317  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_u0_u3_n572 ), .ZN(_AES_ENC_u0_u3_n1074 ) );
NOR2_X2 _AES_ENC_u0_u3_U316  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n584 ), .ZN(_AES_ENC_u0_u3_n838 ) );
NOR2_X2 _AES_ENC_u0_u3_U315  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n602 ), .ZN(_AES_ENC_u0_u3_n837 ) );
NOR2_X2 _AES_ENC_u0_u3_U314  ( .A1(_AES_ENC_u0_u3_n838 ), .A2(_AES_ENC_u0_u3_n837 ), .ZN(_AES_ENC_u0_u3_n845 ) );
NOR2_X2 _AES_ENC_u0_u3_U312  ( .A1(_AES_ENC_u0_u3_n1058 ), .A2(_AES_ENC_u0_u3_n1054 ), .ZN(_AES_ENC_u0_u3_n878 ) );
NOR2_X2 _AES_ENC_u0_u3_U311  ( .A1(_AES_ENC_u0_u3_n878 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n879 ) );
NOR2_X2 _AES_ENC_u0_u3_U310  ( .A1(_AES_ENC_u0_u3_n880 ), .A2(_AES_ENC_u0_u3_n879 ), .ZN(_AES_ENC_u0_u3_n887 ) );
NOR3_X2 _AES_ENC_u0_u3_U309  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n1091 ), .A3(_AES_ENC_u0_u3_n1022 ), .ZN(_AES_ENC_u0_u3_n720 ) );
NOR3_X2 _AES_ENC_u0_u3_U303  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n1054 ), .A3(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n719 ) );
NOR2_X2 _AES_ENC_u0_u3_U302  ( .A1(_AES_ENC_u0_u3_n720 ), .A2(_AES_ENC_u0_u3_n719 ), .ZN(_AES_ENC_u0_u3_n726 ) );
NOR2_X2 _AES_ENC_u0_u3_U300  ( .A1(_AES_ENC_u0_u3_n614 ), .A2(_AES_ENC_u0_u3_n591 ), .ZN(_AES_ENC_u0_u3_n865 ) );
NOR2_X2 _AES_ENC_u0_u3_U299  ( .A1(_AES_ENC_u0_u3_n1059 ), .A2(_AES_ENC_u0_u3_n1058 ), .ZN(_AES_ENC_u0_u3_n1060 ) );
NOR2_X2 _AES_ENC_u0_u3_U298  ( .A1(_AES_ENC_u0_u3_n1095 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n668 ) );
NOR2_X2 _AES_ENC_u0_u3_U297  ( .A1(_AES_ENC_u0_u3_n826 ), .A2(_AES_ENC_u0_u3_n573 ), .ZN(_AES_ENC_u0_u3_n750 ) );
NOR2_X2 _AES_ENC_u0_u3_U296  ( .A1(_AES_ENC_u0_u3_n750 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n751 ) );
NOR2_X2 _AES_ENC_u0_u3_U295  ( .A1(_AES_ENC_u0_u3_n907 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n908 ) );
NOR2_X2 _AES_ENC_u0_u3_U294  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n588 ), .ZN(_AES_ENC_u0_u3_n957 ) );
NOR2_X2 _AES_ENC_u0_u3_U293  ( .A1(_AES_ENC_u0_u3_n990 ), .A2(_AES_ENC_u0_u3_n926 ), .ZN(_AES_ENC_u0_u3_n780 ) );
NOR2_X2 _AES_ENC_u0_u3_U292  ( .A1(_AES_ENC_u0_u3_n1022 ), .A2(_AES_ENC_u0_u3_n1058 ), .ZN(_AES_ENC_u0_u3_n740 ) );
NOR2_X2 _AES_ENC_u0_u3_U291  ( .A1(_AES_ENC_u0_u3_n740 ), .A2(_AES_ENC_u0_u3_n616 ), .ZN(_AES_ENC_u0_u3_n742 ) );
NOR2_X2 _AES_ENC_u0_u3_U290  ( .A1(_AES_ENC_u0_u3_n1098 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n1099 ) );
NOR2_X2 _AES_ENC_u0_u3_U284  ( .A1(_AES_ENC_u0_u3_n1120 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n993 ) );
NOR2_X2 _AES_ENC_u0_u3_U283  ( .A1(_AES_ENC_u0_u3_n993 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n994 ) );
NOR2_X2 _AES_ENC_u0_u3_U282  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n620 ), .ZN(_AES_ENC_u0_u3_n1026 ) );
NOR2_X2 _AES_ENC_u0_u3_U281  ( .A1(_AES_ENC_u0_u3_n573 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n1027 ) );
NOR2_X2 _AES_ENC_u0_u3_U280  ( .A1(_AES_ENC_u0_u3_n1027 ), .A2(_AES_ENC_u0_u3_n1026 ), .ZN(_AES_ENC_u0_u3_n1028 ) );
NOR2_X2 _AES_ENC_u0_u3_U279  ( .A1(_AES_ENC_u0_u3_n1029 ), .A2(_AES_ENC_u0_u3_n1028 ), .ZN(_AES_ENC_u0_u3_n1034 ) );
NOR2_X2 _AES_ENC_u0_u3_U273  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n1071 ), .ZN(_AES_ENC_u0_u3_n669 ) );
NOR2_X2 _AES_ENC_u0_u3_U272  ( .A1(_AES_ENC_u0_u3_n1056 ), .A2(_AES_ENC_u0_u3_n990 ), .ZN(_AES_ENC_u0_u3_n991 ) );
NOR2_X2 _AES_ENC_u0_u3_U271  ( .A1(_AES_ENC_u0_u3_n991 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n995 ) );
NOR4_X2 _AES_ENC_u0_u3_U270  ( .A1(_AES_ENC_u0_u3_n757 ), .A2(_AES_ENC_u0_u3_n756 ), .A3(_AES_ENC_u0_u3_n755 ), .A4(_AES_ENC_u0_u3_n754 ), .ZN(_AES_ENC_u0_u3_n758 ) );
NOR2_X2 _AES_ENC_u0_u3_U269  ( .A1(_AES_ENC_u0_u3_n752 ), .A2(_AES_ENC_u0_u3_n751 ), .ZN(_AES_ENC_u0_u3_n759 ) );
NOR2_X2 _AES_ENC_u0_u3_U268  ( .A1(_AES_ENC_u0_u3_n607 ), .A2(_AES_ENC_u0_u3_n590 ), .ZN(_AES_ENC_u0_u3_n1008 ) );
NOR2_X2 _AES_ENC_u0_u3_U267  ( .A1(_AES_ENC_u0_u3_n606 ), .A2(_AES_ENC_u0_u3_n906 ), .ZN(_AES_ENC_u0_u3_n741 ) );
NOR2_X2 _AES_ENC_u0_u3_U263  ( .A1(_AES_ENC_u0_u3_n1054 ), .A2(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n763 ) );
NOR2_X2 _AES_ENC_u0_u3_U262  ( .A1(_AES_ENC_u0_u3_n763 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n769 ) );
NOR2_X2 _AES_ENC_u0_u3_U258  ( .A1(_AES_ENC_u0_u3_n839 ), .A2(_AES_ENC_u0_u3_n582 ), .ZN(_AES_ENC_u0_u3_n693 ) );
NOR2_X2 _AES_ENC_u0_u3_U255  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n577 ), .ZN(_AES_ENC_u0_u3_n1007 ) );
NOR2_X2 _AES_ENC_u0_u3_U254  ( .A1(_AES_ENC_u0_u3_n609 ), .A2(_AES_ENC_u0_u3_n580 ), .ZN(_AES_ENC_u0_u3_n1123 ) );
NOR2_X2 _AES_ENC_u0_u3_U253  ( .A1(_AES_ENC_u0_u3_n780 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n784 ) );
NOR2_X2 _AES_ENC_u0_u3_U252  ( .A1(_AES_ENC_u0_u3_n1117 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n782 ) );
NOR2_X2 _AES_ENC_u0_u3_U251  ( .A1(_AES_ENC_u0_u3_n781 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n783 ) );
NOR4_X2 _AES_ENC_u0_u3_U250  ( .A1(_AES_ENC_u0_u3_n880 ), .A2(_AES_ENC_u0_u3_n784 ), .A3(_AES_ENC_u0_u3_n783 ), .A4(_AES_ENC_u0_u3_n782 ), .ZN(_AES_ENC_u0_u3_n785 ) );
NOR2_X2 _AES_ENC_u0_u3_U243  ( .A1(_AES_ENC_u0_u3_n609 ), .A2(_AES_ENC_u0_u3_n590 ), .ZN(_AES_ENC_u0_u3_n710 ) );
INV_X4 _AES_ENC_u0_u3_U242  ( .A(_AES_ENC_u0_u3_n1029 ), .ZN(_AES_ENC_u0_u3_n582 ) );
NOR2_X2 _AES_ENC_u0_u3_U241  ( .A1(_AES_ENC_u0_u3_n593 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n1125 ) );
NOR2_X2 _AES_ENC_u0_u3_U240  ( .A1(_AES_ENC_u0_u3_n616 ), .A2(_AES_ENC_u0_u3_n580 ), .ZN(_AES_ENC_u0_u3_n771 ) );
NOR2_X2 _AES_ENC_u0_u3_U239  ( .A1(_AES_ENC_u0_u3_n616 ), .A2(_AES_ENC_u0_u3_n597 ), .ZN(_AES_ENC_u0_u3_n883 ) );
NOR2_X2 _AES_ENC_u0_u3_U238  ( .A1(_AES_ENC_u0_u3_n911 ), .A2(_AES_ENC_u0_u3_n910 ), .ZN(_AES_ENC_u0_u3_n912 ) );
NOR2_X2 _AES_ENC_u0_u3_U237  ( .A1(_AES_ENC_u0_u3_n912 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n916 ) );
NOR2_X2 _AES_ENC_u0_u3_U236  ( .A1(_AES_ENC_u0_u3_n990 ), .A2(_AES_ENC_u0_u3_n929 ), .ZN(_AES_ENC_u0_u3_n892 ) );
NOR2_X2 _AES_ENC_u0_u3_U235  ( .A1(_AES_ENC_u0_u3_n892 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n893 ) );
NOR2_X2 _AES_ENC_u0_u3_U234  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n602 ), .ZN(_AES_ENC_u0_u3_n950 ) );
NOR2_X2 _AES_ENC_u0_u3_U229  ( .A1(_AES_ENC_u0_u3_n1079 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n1082 ) );
NOR2_X2 _AES_ENC_u0_u3_U228  ( .A1(_AES_ENC_u0_u3_n910 ), .A2(_AES_ENC_u0_u3_n1056 ), .ZN(_AES_ENC_u0_u3_n941 ) );
NOR2_X2 _AES_ENC_u0_u3_U227  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n1077 ), .ZN(_AES_ENC_u0_u3_n841 ) );
NOR2_X2 _AES_ENC_u0_u3_U226  ( .A1(_AES_ENC_u0_u3_n623 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n630 ) );
NOR2_X2 _AES_ENC_u0_u3_U225  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n602 ), .ZN(_AES_ENC_u0_u3_n806 ) );
NOR2_X2 _AES_ENC_u0_u3_U223  ( .A1(_AES_ENC_u0_u3_n623 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n948 ) );
NOR2_X2 _AES_ENC_u0_u3_U222  ( .A1(_AES_ENC_u0_u3_n606 ), .A2(_AES_ENC_u0_u3_n582 ), .ZN(_AES_ENC_u0_u3_n1104 ) );
NOR2_X2 _AES_ENC_u0_u3_U221  ( .A1(_AES_ENC_u0_u3_n1121 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n1122 ) );
NOR2_X2 _AES_ENC_u0_u3_U217  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n1023 ), .ZN(_AES_ENC_u0_u3_n756 ) );
NOR2_X2 _AES_ENC_u0_u3_U213  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n602 ), .ZN(_AES_ENC_u0_u3_n870 ) );
NOR2_X2 _AES_ENC_u0_u3_U212  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n569 ), .ZN(_AES_ENC_u0_u3_n947 ) );
NOR2_X2 _AES_ENC_u0_u3_U211  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n1077 ), .ZN(_AES_ENC_u0_u3_n1084 ) );
NOR2_X2 _AES_ENC_u0_u3_U210  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n855 ), .ZN(_AES_ENC_u0_u3_n709 ) );
NOR2_X2 _AES_ENC_u0_u3_U209  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n589 ), .ZN(_AES_ENC_u0_u3_n868 ) );
NOR2_X2 _AES_ENC_u0_u3_U208  ( .A1(_AES_ENC_u0_u3_n1120 ), .A2(_AES_ENC_u0_u3_n839 ), .ZN(_AES_ENC_u0_u3_n842 ) );
NOR2_X2 _AES_ENC_u0_u3_U207  ( .A1(_AES_ENC_u0_u3_n1120 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n1124 ) );
NOR2_X2 _AES_ENC_u0_u3_U201  ( .A1(_AES_ENC_u0_u3_n1120 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n696 ) );
NOR2_X2 _AES_ENC_u0_u3_U200  ( .A1(_AES_ENC_u0_u3_n1074 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n1076 ) );
NOR2_X2 _AES_ENC_u0_u3_U199  ( .A1(_AES_ENC_u0_u3_n1074 ), .A2(_AES_ENC_u0_u3_n620 ), .ZN(_AES_ENC_u0_u3_n781 ) );
NOR3_X2 _AES_ENC_u0_u3_U198  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n1056 ), .A3(_AES_ENC_u0_u3_n990 ), .ZN(_AES_ENC_u0_u3_n979 ) );
NOR3_X2 _AES_ENC_u0_u3_U197  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n1058 ), .A3(_AES_ENC_u0_u3_n1059 ), .ZN(_AES_ENC_u0_u3_n854 ) );
NOR2_X2 _AES_ENC_u0_u3_U196  ( .A1(_AES_ENC_u0_u3_n996 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n869 ) );
NOR2_X2 _AES_ENC_u0_u3_U195  ( .A1(_AES_ENC_u0_u3_n1056 ), .A2(_AES_ENC_u0_u3_n1074 ), .ZN(_AES_ENC_u0_u3_n1057 ) );
NOR3_X2 _AES_ENC_u0_u3_U194  ( .A1(_AES_ENC_u0_u3_n607 ), .A2(_AES_ENC_u0_u3_n1120 ), .A3(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n978 ) );
NOR2_X2 _AES_ENC_u0_u3_U187  ( .A1(_AES_ENC_u0_u3_n996 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n998 ) );
NOR2_X2 _AES_ENC_u0_u3_U186  ( .A1(_AES_ENC_u0_u3_n996 ), .A2(_AES_ENC_u0_u3_n911 ), .ZN(_AES_ENC_u0_u3_n1116 ) );
NOR2_X2 _AES_ENC_u0_u3_U185  ( .A1(_AES_ENC_u0_u3_n1074 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n754 ) );
NOR2_X2 _AES_ENC_u0_u3_U184  ( .A1(_AES_ENC_u0_u3_n926 ), .A2(_AES_ENC_u0_u3_n1103 ), .ZN(_AES_ENC_u0_u3_n977 ) );
NOR2_X2 _AES_ENC_u0_u3_U183  ( .A1(_AES_ENC_u0_u3_n839 ), .A2(_AES_ENC_u0_u3_n824 ), .ZN(_AES_ENC_u0_u3_n1092 ) );
NOR2_X2 _AES_ENC_u0_u3_U182  ( .A1(_AES_ENC_u0_u3_n573 ), .A2(_AES_ENC_u0_u3_n1074 ), .ZN(_AES_ENC_u0_u3_n684 ) );
NOR2_X2 _AES_ENC_u0_u3_U181  ( .A1(_AES_ENC_u0_u3_n826 ), .A2(_AES_ENC_u0_u3_n1059 ), .ZN(_AES_ENC_u0_u3_n907 ) );
NOR3_X2 _AES_ENC_u0_u3_U180  ( .A1(_AES_ENC_u0_u3_n625 ), .A2(_AES_ENC_u0_u3_n1115 ), .A3(_AES_ENC_u0_u3_n585 ), .ZN(_AES_ENC_u0_u3_n831 ) );
NOR3_X2 _AES_ENC_u0_u3_U174  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n1056 ), .A3(_AES_ENC_u0_u3_n990 ), .ZN(_AES_ENC_u0_u3_n896 ) );
NOR3_X2 _AES_ENC_u0_u3_U173  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n573 ), .A3(_AES_ENC_u0_u3_n1013 ), .ZN(_AES_ENC_u0_u3_n670 ) );
NOR3_X2 _AES_ENC_u0_u3_U172  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n1091 ), .A3(_AES_ENC_u0_u3_n1022 ), .ZN(_AES_ENC_u0_u3_n843 ) );
NOR2_X2 _AES_ENC_u0_u3_U171  ( .A1(_AES_ENC_u0_u3_n1029 ), .A2(_AES_ENC_u0_u3_n1095 ), .ZN(_AES_ENC_u0_u3_n735 ) );
NOR4_X2 _AES_ENC_u0_u3_U170  ( .A1(_AES_ENC_u0_u3_n983 ), .A2(_AES_ENC_u0_u3_n698 ), .A3(_AES_ENC_u0_u3_n697 ), .A4(_AES_ENC_u0_u3_n696 ), .ZN(_AES_ENC_u0_u3_n699 ) );
NOR3_X2 _AES_ENC_u0_u3_U169  ( .A1(_AES_ENC_u0_u3_n695 ), .A2(_AES_ENC_u0_u3_n694 ), .A3(_AES_ENC_u0_u3_n693 ), .ZN(_AES_ENC_u0_u3_n700 ) );
NOR2_X2 _AES_ENC_u0_u3_U168  ( .A1(_AES_ENC_u0_u3_n1100 ), .A2(_AES_ENC_u0_u3_n854 ), .ZN(_AES_ENC_u0_u3_n860 ) );
NAND3_X2 _AES_ENC_u0_u3_U162  ( .A1(_AES_ENC_u0_u3_n569 ), .A2(_AES_ENC_u0_u3_n582 ), .A3(_AES_ENC_u0_u3_n681 ), .ZN(_AES_ENC_u0_u3_n691 ) );
NOR2_X2 _AES_ENC_u0_u3_U161  ( .A1(_AES_ENC_u0_u3_n683 ), .A2(_AES_ENC_u0_u3_n682 ), .ZN(_AES_ENC_u0_u3_n690 ) );
NOR4_X2 _AES_ENC_u0_u3_U160  ( .A1(_AES_ENC_u0_u3_n896 ), .A2(_AES_ENC_u0_u3_n895 ), .A3(_AES_ENC_u0_u3_n894 ), .A4(_AES_ENC_u0_u3_n893 ), .ZN(_AES_ENC_u0_u3_n897 ) );
NOR2_X2 _AES_ENC_u0_u3_U159  ( .A1(_AES_ENC_u0_u3_n866 ), .A2(_AES_ENC_u0_u3_n865 ), .ZN(_AES_ENC_u0_u3_n872 ) );
NOR4_X2 _AES_ENC_u0_u3_U158  ( .A1(_AES_ENC_u0_u3_n870 ), .A2(_AES_ENC_u0_u3_n869 ), .A3(_AES_ENC_u0_u3_n868 ), .A4(_AES_ENC_u0_u3_n867 ), .ZN(_AES_ENC_u0_u3_n871 ) );
NOR4_X2 _AES_ENC_u0_u3_U157  ( .A1(_AES_ENC_u0_u3_n963 ), .A2(_AES_ENC_u0_u3_n962 ), .A3(_AES_ENC_u0_u3_n961 ), .A4(_AES_ENC_u0_u3_n960 ), .ZN(_AES_ENC_u0_u3_n964 ) );
NOR2_X2 _AES_ENC_u0_u3_U156  ( .A1(_AES_ENC_u0_u3_n958 ), .A2(_AES_ENC_u0_u3_n957 ), .ZN(_AES_ENC_u0_u3_n965 ) );
NOR4_X2 _AES_ENC_u0_u3_U155  ( .A1(_AES_ENC_u0_u3_n950 ), .A2(_AES_ENC_u0_u3_n949 ), .A3(_AES_ENC_u0_u3_n948 ), .A4(_AES_ENC_u0_u3_n947 ), .ZN(_AES_ENC_u0_u3_n951 ) );
NOR2_X2 _AES_ENC_u0_u3_U154  ( .A1(_AES_ENC_u0_u3_n946 ), .A2(_AES_ENC_u0_u3_n945 ), .ZN(_AES_ENC_u0_u3_n952 ) );
NOR4_X2 _AES_ENC_u0_u3_U153  ( .A1(_AES_ENC_u0_u3_n983 ), .A2(_AES_ENC_u0_u3_n982 ), .A3(_AES_ENC_u0_u3_n981 ), .A4(_AES_ENC_u0_u3_n980 ), .ZN(_AES_ENC_u0_u3_n984 ) );
NOR2_X2 _AES_ENC_u0_u3_U152  ( .A1(_AES_ENC_u0_u3_n979 ), .A2(_AES_ENC_u0_u3_n978 ), .ZN(_AES_ENC_u0_u3_n985 ) );
NOR4_X2 _AES_ENC_u0_u3_U143  ( .A1(_AES_ENC_u0_u3_n1125 ), .A2(_AES_ENC_u0_u3_n1124 ), .A3(_AES_ENC_u0_u3_n1123 ), .A4(_AES_ENC_u0_u3_n1122 ), .ZN(_AES_ENC_u0_u3_n1126 ) );
NOR4_X2 _AES_ENC_u0_u3_U142  ( .A1(_AES_ENC_u0_u3_n1084 ), .A2(_AES_ENC_u0_u3_n1083 ), .A3(_AES_ENC_u0_u3_n1082 ), .A4(_AES_ENC_u0_u3_n1081 ), .ZN(_AES_ENC_u0_u3_n1085 ) );
NOR2_X2 _AES_ENC_u0_u3_U141  ( .A1(_AES_ENC_u0_u3_n1076 ), .A2(_AES_ENC_u0_u3_n1075 ), .ZN(_AES_ENC_u0_u3_n1086 ) );
NOR3_X2 _AES_ENC_u0_u3_U140  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n1054 ), .A3(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n961 ) );
NOR3_X2 _AES_ENC_u0_u3_U132  ( .A1(_AES_ENC_u0_u3_n620 ), .A2(_AES_ENC_u0_u3_n1074 ), .A3(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n671 ) );
NOR2_X2 _AES_ENC_u0_u3_U131  ( .A1(_AES_ENC_u0_u3_n1057 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n1062 ) );
NOR2_X2 _AES_ENC_u0_u3_U130  ( .A1(_AES_ENC_u0_u3_n1060 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n1061 ) );
NOR2_X2 _AES_ENC_u0_u3_U129  ( .A1(_AES_ENC_u0_u3_n1055 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n1063 ) );
NOR4_X2 _AES_ENC_u0_u3_U128  ( .A1(_AES_ENC_u0_u3_n1064 ), .A2(_AES_ENC_u0_u3_n1063 ), .A3(_AES_ENC_u0_u3_n1062 ), .A4(_AES_ENC_u0_u3_n1061 ), .ZN(_AES_ENC_u0_u3_n1065 ) );
NOR3_X2 _AES_ENC_u0_u3_U127  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n1120 ), .A3(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n918 ) );
NOR2_X2 _AES_ENC_u0_u3_U126  ( .A1(_AES_ENC_u0_u3_n914 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n915 ) );
NOR3_X2 _AES_ENC_u0_u3_U121  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n573 ), .A3(_AES_ENC_u0_u3_n1013 ), .ZN(_AES_ENC_u0_u3_n917 ) );
NOR4_X2 _AES_ENC_u0_u3_U120  ( .A1(_AES_ENC_u0_u3_n918 ), .A2(_AES_ENC_u0_u3_n917 ), .A3(_AES_ENC_u0_u3_n916 ), .A4(_AES_ENC_u0_u3_n915 ), .ZN(_AES_ENC_u0_u3_n919 ) );
NOR2_X2 _AES_ENC_u0_u3_U119  ( .A1(_AES_ENC_u0_u3_n735 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n687 ) );
NOR2_X2 _AES_ENC_u0_u3_U118  ( .A1(_AES_ENC_u0_u3_n684 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n688 ) );
NOR2_X2 _AES_ENC_u0_u3_U117  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n600 ), .ZN(_AES_ENC_u0_u3_n686 ) );
NOR4_X2 _AES_ENC_u0_u3_U116  ( .A1(_AES_ENC_u0_u3_n688 ), .A2(_AES_ENC_u0_u3_n687 ), .A3(_AES_ENC_u0_u3_n686 ), .A4(_AES_ENC_u0_u3_n685 ), .ZN(_AES_ENC_u0_u3_n689 ) );
NOR2_X2 _AES_ENC_u0_u3_U115  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n582 ), .ZN(_AES_ENC_u0_u3_n770 ) );
NOR2_X2 _AES_ENC_u0_u3_U106  ( .A1(_AES_ENC_u0_u3_n1103 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n772 ) );
NOR2_X2 _AES_ENC_u0_u3_U105  ( .A1(_AES_ENC_u0_u3_n610 ), .A2(_AES_ENC_u0_u3_n599 ), .ZN(_AES_ENC_u0_u3_n773 ) );
NOR4_X2 _AES_ENC_u0_u3_U104  ( .A1(_AES_ENC_u0_u3_n773 ), .A2(_AES_ENC_u0_u3_n772 ), .A3(_AES_ENC_u0_u3_n771 ), .A4(_AES_ENC_u0_u3_n770 ), .ZN(_AES_ENC_u0_u3_n774 ) );
NOR2_X2 _AES_ENC_u0_u3_U103  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n595 ), .ZN(_AES_ENC_u0_u3_n858 ) );
NOR2_X2 _AES_ENC_u0_u3_U102  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n855 ), .ZN(_AES_ENC_u0_u3_n857 ) );
NOR2_X2 _AES_ENC_u0_u3_U101  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n587 ), .ZN(_AES_ENC_u0_u3_n856 ) );
NOR4_X2 _AES_ENC_u0_u3_U100  ( .A1(_AES_ENC_u0_u3_n858 ), .A2(_AES_ENC_u0_u3_n857 ), .A3(_AES_ENC_u0_u3_n856 ), .A4(_AES_ENC_u0_u3_n958 ), .ZN(_AES_ENC_u0_u3_n859 ) );
NOR2_X2 _AES_ENC_u0_u3_U95  ( .A1(_AES_ENC_u0_u3_n583 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n814 ) );
NOR3_X2 _AES_ENC_u0_u3_U94  ( .A1(_AES_ENC_u0_u3_n606 ), .A2(_AES_ENC_u0_u3_n1058 ), .A3(_AES_ENC_u0_u3_n1059 ), .ZN(_AES_ENC_u0_u3_n815 ) );
NOR2_X2 _AES_ENC_u0_u3_U93  ( .A1(_AES_ENC_u0_u3_n907 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n813 ) );
NOR4_X2 _AES_ENC_u0_u3_U92  ( .A1(_AES_ENC_u0_u3_n815 ), .A2(_AES_ENC_u0_u3_n814 ), .A3(_AES_ENC_u0_u3_n813 ), .A4(_AES_ENC_u0_u3_n812 ), .ZN(_AES_ENC_u0_u3_n816 ) );
NOR2_X2 _AES_ENC_u0_u3_U91  ( .A1(_AES_ENC_u0_u3_n617 ), .A2(_AES_ENC_u0_u3_n569 ), .ZN(_AES_ENC_u0_u3_n721 ) );
NOR2_X2 _AES_ENC_u0_u3_U90  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n1096 ), .ZN(_AES_ENC_u0_u3_n722 ) );
NOR2_X2 _AES_ENC_u0_u3_U89  ( .A1(_AES_ENC_u0_u3_n1031 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n723 ) );
NOR4_X2 _AES_ENC_u0_u3_U88  ( .A1(_AES_ENC_u0_u3_n724 ), .A2(_AES_ENC_u0_u3_n723 ), .A3(_AES_ENC_u0_u3_n722 ), .A4(_AES_ENC_u0_u3_n721 ), .ZN(_AES_ENC_u0_u3_n725 ) );
NOR2_X2 _AES_ENC_u0_u3_U87  ( .A1(_AES_ENC_u0_u3_n911 ), .A2(_AES_ENC_u0_u3_n990 ), .ZN(_AES_ENC_u0_u3_n1009 ) );
NOR2_X2 _AES_ENC_u0_u3_U86  ( .A1(_AES_ENC_u0_u3_n1013 ), .A2(_AES_ENC_u0_u3_n573 ), .ZN(_AES_ENC_u0_u3_n1014 ) );
NOR2_X2 _AES_ENC_u0_u3_U81  ( .A1(_AES_ENC_u0_u3_n1014 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n1015 ) );
NOR4_X2 _AES_ENC_u0_u3_U80  ( .A1(_AES_ENC_u0_u3_n1016 ), .A2(_AES_ENC_u0_u3_n1015 ), .A3(_AES_ENC_u0_u3_n1119 ), .A4(_AES_ENC_u0_u3_n1046 ), .ZN(_AES_ENC_u0_u3_n1017 ) );
NOR2_X2 _AES_ENC_u0_u3_U79  ( .A1(_AES_ENC_u0_u3_n606 ), .A2(_AES_ENC_u0_u3_n589 ), .ZN(_AES_ENC_u0_u3_n997 ) );
NOR2_X2 _AES_ENC_u0_u3_U78  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n577 ), .ZN(_AES_ENC_u0_u3_n1000 ) );
NOR2_X2 _AES_ENC_u0_u3_U74  ( .A1(_AES_ENC_u0_u3_n616 ), .A2(_AES_ENC_u0_u3_n1096 ), .ZN(_AES_ENC_u0_u3_n999 ) );
NOR4_X2 _AES_ENC_u0_u3_U73  ( .A1(_AES_ENC_u0_u3_n1000 ), .A2(_AES_ENC_u0_u3_n999 ), .A3(_AES_ENC_u0_u3_n998 ), .A4(_AES_ENC_u0_u3_n997 ), .ZN(_AES_ENC_u0_u3_n1001 ) );
NOR2_X2 _AES_ENC_u0_u3_U72  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n1096 ), .ZN(_AES_ENC_u0_u3_n697 ) );
NOR2_X2 _AES_ENC_u0_u3_U71  ( .A1(_AES_ENC_u0_u3_n620 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n958 ) );
NOR2_X2 _AES_ENC_u0_u3_U65  ( .A1(_AES_ENC_u0_u3_n911 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n983 ) );
NOR2_X2 _AES_ENC_u0_u3_U64  ( .A1(_AES_ENC_u0_u3_n1054 ), .A2(_AES_ENC_u0_u3_n1103 ), .ZN(_AES_ENC_u0_u3_n1031 ) );
INV_X4 _AES_ENC_u0_u3_U63  ( .A(_AES_ENC_u0_u3_n1050 ), .ZN(_AES_ENC_u0_u3_n612 ) );
INV_X4 _AES_ENC_u0_u3_U62  ( .A(_AES_ENC_u0_u3_n1072 ), .ZN(_AES_ENC_u0_u3_n605 ) );
INV_X4 _AES_ENC_u0_u3_U61  ( .A(_AES_ENC_u0_u3_n1073 ), .ZN(_AES_ENC_u0_u3_n604 ) );
NOR2_X2 _AES_ENC_u0_u3_U59  ( .A1(_AES_ENC_u0_u3_n582 ), .A2(_AES_ENC_u0_u3_n613 ), .ZN(_AES_ENC_u0_u3_n880 ) );
NOR3_X2 _AES_ENC_u0_u3_U58  ( .A1(_AES_ENC_u0_u3_n826 ), .A2(_AES_ENC_u0_u3_n1121 ), .A3(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n946 ) );
INV_X4 _AES_ENC_u0_u3_U57  ( .A(_AES_ENC_u0_u3_n1010 ), .ZN(_AES_ENC_u0_u3_n608 ) );
NOR3_X2 _AES_ENC_u0_u3_U50  ( .A1(_AES_ENC_u0_u3_n573 ), .A2(_AES_ENC_u0_u3_n1029 ), .A3(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n1119 ) );
INV_X4 _AES_ENC_u0_u3_U49  ( .A(_AES_ENC_u0_u3_n956 ), .ZN(_AES_ENC_u0_u3_n615 ) );
NOR2_X2 _AES_ENC_u0_u3_U48  ( .A1(_AES_ENC_u0_u3_n623 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n1013 ) );
NOR2_X2 _AES_ENC_u0_u3_U47  ( .A1(_AES_ENC_u0_u3_n620 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n910 ) );
NOR2_X2 _AES_ENC_u0_u3_U46  ( .A1(_AES_ENC_u0_u3_n569 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n1091 ) );
NOR2_X2 _AES_ENC_u0_u3_U45  ( .A1(_AES_ENC_u0_u3_n622 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n990 ) );
NOR2_X2 _AES_ENC_u0_u3_U44  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_u0_u3_n1121 ), .ZN(_AES_ENC_u0_u3_n996 ) );
NOR2_X2 _AES_ENC_u0_u3_U43  ( .A1(_AES_ENC_u0_u3_n610 ), .A2(_AES_ENC_u0_u3_n600 ), .ZN(_AES_ENC_u0_u3_n628 ) );
NOR2_X2 _AES_ENC_u0_u3_U42  ( .A1(_AES_ENC_u0_u3_n576 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n866 ) );
NOR2_X2 _AES_ENC_u0_u3_U41  ( .A1(_AES_ENC_u0_u3_n603 ), .A2(_AES_ENC_u0_u3_n610 ), .ZN(_AES_ENC_u0_u3_n1006 ) );
NOR2_X2 _AES_ENC_u0_u3_U36  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n1117 ), .ZN(_AES_ENC_u0_u3_n1118 ) );
NOR2_X2 _AES_ENC_u0_u3_U35  ( .A1(_AES_ENC_u0_u3_n1119 ), .A2(_AES_ENC_u0_u3_n1118 ), .ZN(_AES_ENC_u0_u3_n1127 ) );
NOR2_X2 _AES_ENC_u0_u3_U34  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n594 ), .ZN(_AES_ENC_u0_u3_n629 ) );
NOR2_X2 _AES_ENC_u0_u3_U33  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n906 ), .ZN(_AES_ENC_u0_u3_n909 ) );
NOR2_X2 _AES_ENC_u0_u3_U32  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n597 ), .ZN(_AES_ENC_u0_u3_n658 ) );
NOR2_X2 _AES_ENC_u0_u3_U31  ( .A1(_AES_ENC_u0_u3_n1116 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n695 ) );
NOR2_X2 _AES_ENC_u0_u3_U30  ( .A1(_AES_ENC_u0_u3_n1078 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n1083 ) );
NOR2_X2 _AES_ENC_u0_u3_U29  ( .A1(_AES_ENC_u0_u3_n941 ), .A2(_AES_ENC_u0_u3_n608 ), .ZN(_AES_ENC_u0_u3_n724 ) );
NOR2_X2 _AES_ENC_u0_u3_U24  ( .A1(_AES_ENC_u0_u3_n576 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n840 ) );
NOR2_X2 _AES_ENC_u0_u3_U23  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n593 ), .ZN(_AES_ENC_u0_u3_n633 ) );
NOR2_X2 _AES_ENC_u0_u3_U21  ( .A1(_AES_ENC_u0_u3_n1009 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n960 ) );
NOR2_X2 _AES_ENC_u0_u3_U20  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n1045 ), .ZN(_AES_ENC_u0_u3_n812 ) );
NOR2_X2 _AES_ENC_u0_u3_U19  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n1080 ), .ZN(_AES_ENC_u0_u3_n1081 ) );
NOR2_X2 _AES_ENC_u0_u3_U18  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n601 ), .ZN(_AES_ENC_u0_u3_n982 ) );
NOR2_X2 _AES_ENC_u0_u3_U17  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n594 ), .ZN(_AES_ENC_u0_u3_n757 ) );
NOR2_X2 _AES_ENC_u0_u3_U16  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n590 ), .ZN(_AES_ENC_u0_u3_n698 ) );
NOR2_X2 _AES_ENC_u0_u3_U15  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n619 ), .ZN(_AES_ENC_u0_u3_n708 ) );
NOR2_X2 _AES_ENC_u0_u3_U10  ( .A1(_AES_ENC_u0_u3_n619 ), .A2(_AES_ENC_u0_u3_n604 ), .ZN(_AES_ENC_u0_u3_n803 ) );
NOR2_X2 _AES_ENC_u0_u3_U9  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n881 ), .ZN(_AES_ENC_u0_u3_n711 ) );
NOR2_X2 _AES_ENC_u0_u3_U8  ( .A1(_AES_ENC_u0_u3_n615 ), .A2(_AES_ENC_u0_u3_n582 ), .ZN(_AES_ENC_u0_u3_n867 ) );
NOR2_X2 _AES_ENC_u0_u3_U7  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n599 ), .ZN(_AES_ENC_u0_u3_n804 ) );
NOR2_X2 _AES_ENC_u0_u3_U6  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n620 ), .ZN(_AES_ENC_u0_u3_n1046 ) );
OR2_X4 _AES_ENC_u0_u3_U5  ( .A1(_AES_ENC_u0_u3_n624 ), .A2(_AES_ENC_w3[25] ),.ZN(_AES_ENC_u0_u3_n570 ) );
OR2_X4 _AES_ENC_u0_u3_U4  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_w3[28] ),.ZN(_AES_ENC_u0_u3_n569 ) );
NAND2_X2 _AES_ENC_u0_u3_U514  ( .A1(_AES_ENC_u0_u3_n1121 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n1030 ) );
AND2_X2 _AES_ENC_u0_u3_U513  ( .A1(_AES_ENC_u0_u3_n597 ), .A2(_AES_ENC_u0_u3_n1030 ), .ZN(_AES_ENC_u0_u3_n1049 ) );
NAND2_X2 _AES_ENC_u0_u3_U511  ( .A1(_AES_ENC_u0_u3_n1049 ), .A2(_AES_ENC_u0_u3_n794 ), .ZN(_AES_ENC_u0_u3_n637 ) );
AND2_X2 _AES_ENC_u0_u3_U493  ( .A1(_AES_ENC_u0_u3_n779 ), .A2(_AES_ENC_u0_u3_n996 ), .ZN(_AES_ENC_u0_u3_n632 ) );
NAND4_X2 _AES_ENC_u0_u3_U485  ( .A1(_AES_ENC_u0_u3_n637 ), .A2(_AES_ENC_u0_u3_n636 ), .A3(_AES_ENC_u0_u3_n635 ), .A4(_AES_ENC_u0_u3_n634 ), .ZN(_AES_ENC_u0_u3_n638 ) );
NAND2_X2 _AES_ENC_u0_u3_U484  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n638 ), .ZN(_AES_ENC_u0_u3_n679 ) );
NAND2_X2 _AES_ENC_u0_u3_U481  ( .A1(_AES_ENC_u0_u3_n1094 ), .A2(_AES_ENC_u0_u3_n591 ), .ZN(_AES_ENC_u0_u3_n648 ) );
NAND2_X2 _AES_ENC_u0_u3_U476  ( .A1(_AES_ENC_u0_u3_n601 ), .A2(_AES_ENC_u0_u3_n590 ), .ZN(_AES_ENC_u0_u3_n762 ) );
NAND2_X2 _AES_ENC_u0_u3_U475  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n762 ), .ZN(_AES_ENC_u0_u3_n647 ) );
NAND4_X2 _AES_ENC_u0_u3_U457  ( .A1(_AES_ENC_u0_u3_n648 ), .A2(_AES_ENC_u0_u3_n647 ), .A3(_AES_ENC_u0_u3_n646 ), .A4(_AES_ENC_u0_u3_n645 ), .ZN(_AES_ENC_u0_u3_n649 ) );
NAND2_X2 _AES_ENC_u0_u3_U456  ( .A1(_AES_ENC_w3[24] ), .A2(_AES_ENC_u0_u3_n649 ), .ZN(_AES_ENC_u0_u3_n665 ) );
NAND2_X2 _AES_ENC_u0_u3_U454  ( .A1(_AES_ENC_u0_u3_n596 ), .A2(_AES_ENC_u0_u3_n623 ), .ZN(_AES_ENC_u0_u3_n855 ) );
NAND2_X2 _AES_ENC_u0_u3_U453  ( .A1(_AES_ENC_u0_u3_n587 ), .A2(_AES_ENC_u0_u3_n855 ), .ZN(_AES_ENC_u0_u3_n821 ) );
NAND2_X2 _AES_ENC_u0_u3_U452  ( .A1(_AES_ENC_u0_u3_n1093 ), .A2(_AES_ENC_u0_u3_n821 ), .ZN(_AES_ENC_u0_u3_n662 ) );
NAND2_X2 _AES_ENC_u0_u3_U451  ( .A1(_AES_ENC_u0_u3_n619 ), .A2(_AES_ENC_u0_u3_n589 ), .ZN(_AES_ENC_u0_u3_n650 ) );
NAND2_X2 _AES_ENC_u0_u3_U450  ( .A1(_AES_ENC_u0_u3_n956 ), .A2(_AES_ENC_u0_u3_n650 ), .ZN(_AES_ENC_u0_u3_n661 ) );
NAND2_X2 _AES_ENC_u0_u3_U449  ( .A1(_AES_ENC_u0_u3_n626 ), .A2(_AES_ENC_u0_u3_n627 ), .ZN(_AES_ENC_u0_u3_n839 ) );
OR2_X2 _AES_ENC_u0_u3_U446  ( .A1(_AES_ENC_u0_u3_n839 ), .A2(_AES_ENC_u0_u3_n932 ), .ZN(_AES_ENC_u0_u3_n656 ) );
NAND2_X2 _AES_ENC_u0_u3_U445  ( .A1(_AES_ENC_u0_u3_n621 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n1096 ) );
NAND2_X2 _AES_ENC_u0_u3_U444  ( .A1(_AES_ENC_u0_u3_n1030 ), .A2(_AES_ENC_u0_u3_n1096 ), .ZN(_AES_ENC_u0_u3_n651 ) );
NAND2_X2 _AES_ENC_u0_u3_U443  ( .A1(_AES_ENC_u0_u3_n1114 ), .A2(_AES_ENC_u0_u3_n651 ), .ZN(_AES_ENC_u0_u3_n655 ) );
OR3_X2 _AES_ENC_u0_u3_U440  ( .A1(_AES_ENC_u0_u3_n1079 ), .A2(_AES_ENC_w3[31] ), .A3(_AES_ENC_u0_u3_n626 ), .ZN(_AES_ENC_u0_u3_n654 ) );
NAND2_X2 _AES_ENC_u0_u3_U439  ( .A1(_AES_ENC_u0_u3_n593 ), .A2(_AES_ENC_u0_u3_n601 ), .ZN(_AES_ENC_u0_u3_n652 ) );
NAND4_X2 _AES_ENC_u0_u3_U437  ( .A1(_AES_ENC_u0_u3_n656 ), .A2(_AES_ENC_u0_u3_n655 ), .A3(_AES_ENC_u0_u3_n654 ), .A4(_AES_ENC_u0_u3_n653 ), .ZN(_AES_ENC_u0_u3_n657 ) );
NAND2_X2 _AES_ENC_u0_u3_U436  ( .A1(_AES_ENC_w3[26] ), .A2(_AES_ENC_u0_u3_n657 ), .ZN(_AES_ENC_u0_u3_n660 ) );
NAND4_X2 _AES_ENC_u0_u3_U432  ( .A1(_AES_ENC_u0_u3_n662 ), .A2(_AES_ENC_u0_u3_n661 ), .A3(_AES_ENC_u0_u3_n660 ), .A4(_AES_ENC_u0_u3_n659 ), .ZN(_AES_ENC_u0_u3_n663 ) );
NAND2_X2 _AES_ENC_u0_u3_U431  ( .A1(_AES_ENC_u0_u3_n663 ), .A2(_AES_ENC_u0_u3_n574 ), .ZN(_AES_ENC_u0_u3_n664 ) );
NAND2_X2 _AES_ENC_u0_u3_U430  ( .A1(_AES_ENC_u0_u3_n665 ), .A2(_AES_ENC_u0_u3_n664 ), .ZN(_AES_ENC_u0_u3_n666 ) );
NAND2_X2 _AES_ENC_u0_u3_U429  ( .A1(_AES_ENC_w3[30] ), .A2(_AES_ENC_u0_u3_n666 ), .ZN(_AES_ENC_u0_u3_n678 ) );
NAND2_X2 _AES_ENC_u0_u3_U426  ( .A1(_AES_ENC_u0_u3_n735 ), .A2(_AES_ENC_u0_u3_n1093 ), .ZN(_AES_ENC_u0_u3_n675 ) );
NAND2_X2 _AES_ENC_u0_u3_U425  ( .A1(_AES_ENC_u0_u3_n588 ), .A2(_AES_ENC_u0_u3_n597 ), .ZN(_AES_ENC_u0_u3_n1045 ) );
OR2_X2 _AES_ENC_u0_u3_U424  ( .A1(_AES_ENC_u0_u3_n1045 ), .A2(_AES_ENC_u0_u3_n605 ), .ZN(_AES_ENC_u0_u3_n674 ) );
NAND2_X2 _AES_ENC_u0_u3_U423  ( .A1(_AES_ENC_w3[25] ), .A2(_AES_ENC_u0_u3_n620 ), .ZN(_AES_ENC_u0_u3_n667 ) );
NAND2_X2 _AES_ENC_u0_u3_U422  ( .A1(_AES_ENC_u0_u3_n619 ), .A2(_AES_ENC_u0_u3_n667 ), .ZN(_AES_ENC_u0_u3_n1071 ) );
NAND4_X2 _AES_ENC_u0_u3_U412  ( .A1(_AES_ENC_u0_u3_n675 ), .A2(_AES_ENC_u0_u3_n674 ), .A3(_AES_ENC_u0_u3_n673 ), .A4(_AES_ENC_u0_u3_n672 ), .ZN(_AES_ENC_u0_u3_n676 ) );
NAND2_X2 _AES_ENC_u0_u3_U411  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n676 ), .ZN(_AES_ENC_u0_u3_n677 ) );
NAND2_X2 _AES_ENC_u0_u3_U408  ( .A1(_AES_ENC_u0_u3_n800 ), .A2(_AES_ENC_u0_u3_n1022 ), .ZN(_AES_ENC_u0_u3_n680 ) );
NAND2_X2 _AES_ENC_u0_u3_U407  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n680 ), .ZN(_AES_ENC_u0_u3_n681 ) );
AND2_X2 _AES_ENC_u0_u3_U402  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n684 ), .ZN(_AES_ENC_u0_u3_n682 ) );
NAND4_X2 _AES_ENC_u0_u3_U395  ( .A1(_AES_ENC_u0_u3_n691 ), .A2(_AES_ENC_u0_u3_n581 ), .A3(_AES_ENC_u0_u3_n690 ), .A4(_AES_ENC_u0_u3_n689 ), .ZN(_AES_ENC_u0_u3_n692 ) );
NAND2_X2 _AES_ENC_u0_u3_U394  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n692 ), .ZN(_AES_ENC_u0_u3_n733 ) );
NAND2_X2 _AES_ENC_u0_u3_U392  ( .A1(_AES_ENC_u0_u3_n977 ), .A2(_AES_ENC_u0_u3_n1050 ), .ZN(_AES_ENC_u0_u3_n702 ) );
NAND2_X2 _AES_ENC_u0_u3_U391  ( .A1(_AES_ENC_u0_u3_n1093 ), .A2(_AES_ENC_u0_u3_n1045 ), .ZN(_AES_ENC_u0_u3_n701 ) );
NAND4_X2 _AES_ENC_u0_u3_U381  ( .A1(_AES_ENC_u0_u3_n702 ), .A2(_AES_ENC_u0_u3_n701 ), .A3(_AES_ENC_u0_u3_n700 ), .A4(_AES_ENC_u0_u3_n699 ), .ZN(_AES_ENC_u0_u3_n703 ) );
NAND2_X2 _AES_ENC_u0_u3_U380  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n703 ), .ZN(_AES_ENC_u0_u3_n732 ) );
AND2_X2 _AES_ENC_u0_u3_U379  ( .A1(_AES_ENC_w3[24] ), .A2(_AES_ENC_w3[30] ),.ZN(_AES_ENC_u0_u3_n1113 ) );
NAND2_X2 _AES_ENC_u0_u3_U378  ( .A1(_AES_ENC_u0_u3_n601 ), .A2(_AES_ENC_u0_u3_n1030 ), .ZN(_AES_ENC_u0_u3_n881 ) );
NAND2_X2 _AES_ENC_u0_u3_U377  ( .A1(_AES_ENC_u0_u3_n1093 ), .A2(_AES_ENC_u0_u3_n881 ), .ZN(_AES_ENC_u0_u3_n715 ) );
NAND2_X2 _AES_ENC_u0_u3_U376  ( .A1(_AES_ENC_u0_u3_n1010 ), .A2(_AES_ENC_u0_u3_n600 ), .ZN(_AES_ENC_u0_u3_n714 ) );
NAND2_X2 _AES_ENC_u0_u3_U375  ( .A1(_AES_ENC_u0_u3_n855 ), .A2(_AES_ENC_u0_u3_n588 ), .ZN(_AES_ENC_u0_u3_n1117 ) );
XNOR2_X2 _AES_ENC_u0_u3_U371  ( .A(_AES_ENC_u0_u3_n611 ), .B(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n824 ) );
NAND4_X2 _AES_ENC_u0_u3_U362  ( .A1(_AES_ENC_u0_u3_n715 ), .A2(_AES_ENC_u0_u3_n714 ), .A3(_AES_ENC_u0_u3_n713 ), .A4(_AES_ENC_u0_u3_n712 ), .ZN(_AES_ENC_u0_u3_n716 ) );
NAND2_X2 _AES_ENC_u0_u3_U361  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n716 ), .ZN(_AES_ENC_u0_u3_n731 ) );
AND2_X2 _AES_ENC_u0_u3_U360  ( .A1(_AES_ENC_w3[30] ), .A2(_AES_ENC_u0_u3_n574 ), .ZN(_AES_ENC_u0_u3_n1131 ) );
NAND2_X2 _AES_ENC_u0_u3_U359  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n717 ) );
NAND2_X2 _AES_ENC_u0_u3_U358  ( .A1(_AES_ENC_u0_u3_n1029 ), .A2(_AES_ENC_u0_u3_n717 ), .ZN(_AES_ENC_u0_u3_n728 ) );
NAND2_X2 _AES_ENC_u0_u3_U357  ( .A1(_AES_ENC_w3[25] ), .A2(_AES_ENC_u0_u3_n624 ), .ZN(_AES_ENC_u0_u3_n1097 ) );
NAND2_X2 _AES_ENC_u0_u3_U356  ( .A1(_AES_ENC_u0_u3_n603 ), .A2(_AES_ENC_u0_u3_n1097 ), .ZN(_AES_ENC_u0_u3_n718 ) );
NAND2_X2 _AES_ENC_u0_u3_U355  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n718 ), .ZN(_AES_ENC_u0_u3_n727 ) );
NAND4_X2 _AES_ENC_u0_u3_U344  ( .A1(_AES_ENC_u0_u3_n728 ), .A2(_AES_ENC_u0_u3_n727 ), .A3(_AES_ENC_u0_u3_n726 ), .A4(_AES_ENC_u0_u3_n725 ), .ZN(_AES_ENC_u0_u3_n729 ) );
NAND2_X2 _AES_ENC_u0_u3_U343  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n729 ), .ZN(_AES_ENC_u0_u3_n730 ) );
NAND4_X2 _AES_ENC_u0_u3_U342  ( .A1(_AES_ENC_u0_u3_n733 ), .A2(_AES_ENC_u0_u3_n732 ), .A3(_AES_ENC_u0_u3_n731 ), .A4(_AES_ENC_u0_u3_n730 ), .ZN(_AES_ENC_u0_subword[1] ) );
NAND2_X2 _AES_ENC_u0_u3_U341  ( .A1(_AES_ENC_w3[31] ), .A2(_AES_ENC_u0_u3_n611 ), .ZN(_AES_ENC_u0_u3_n734 ) );
NAND2_X2 _AES_ENC_u0_u3_U340  ( .A1(_AES_ENC_u0_u3_n734 ), .A2(_AES_ENC_u0_u3_n607 ), .ZN(_AES_ENC_u0_u3_n738 ) );
OR4_X2 _AES_ENC_u0_u3_U339  ( .A1(_AES_ENC_u0_u3_n738 ), .A2(_AES_ENC_u0_u3_n626 ), .A3(_AES_ENC_u0_u3_n826 ), .A4(_AES_ENC_u0_u3_n1121 ), .ZN(_AES_ENC_u0_u3_n746 ) );
NAND2_X2 _AES_ENC_u0_u3_U337  ( .A1(_AES_ENC_u0_u3_n1100 ), .A2(_AES_ENC_u0_u3_n587 ), .ZN(_AES_ENC_u0_u3_n992 ) );
OR2_X2 _AES_ENC_u0_u3_U336  ( .A1(_AES_ENC_u0_u3_n610 ), .A2(_AES_ENC_u0_u3_n735 ), .ZN(_AES_ENC_u0_u3_n737 ) );
NAND2_X2 _AES_ENC_u0_u3_U334  ( .A1(_AES_ENC_u0_u3_n619 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n753 ) );
NAND2_X2 _AES_ENC_u0_u3_U333  ( .A1(_AES_ENC_u0_u3_n582 ), .A2(_AES_ENC_u0_u3_n753 ), .ZN(_AES_ENC_u0_u3_n1080 ) );
NAND2_X2 _AES_ENC_u0_u3_U332  ( .A1(_AES_ENC_u0_u3_n1048 ), .A2(_AES_ENC_u0_u3_n576 ), .ZN(_AES_ENC_u0_u3_n736 ) );
NAND2_X2 _AES_ENC_u0_u3_U331  ( .A1(_AES_ENC_u0_u3_n737 ), .A2(_AES_ENC_u0_u3_n736 ), .ZN(_AES_ENC_u0_u3_n739 ) );
NAND2_X2 _AES_ENC_u0_u3_U330  ( .A1(_AES_ENC_u0_u3_n739 ), .A2(_AES_ENC_u0_u3_n738 ), .ZN(_AES_ENC_u0_u3_n745 ) );
NAND2_X2 _AES_ENC_u0_u3_U326  ( .A1(_AES_ENC_u0_u3_n1096 ), .A2(_AES_ENC_u0_u3_n590 ), .ZN(_AES_ENC_u0_u3_n906 ) );
NAND4_X2 _AES_ENC_u0_u3_U323  ( .A1(_AES_ENC_u0_u3_n746 ), .A2(_AES_ENC_u0_u3_n992 ), .A3(_AES_ENC_u0_u3_n745 ), .A4(_AES_ENC_u0_u3_n744 ), .ZN(_AES_ENC_u0_u3_n747 ) );
NAND2_X2 _AES_ENC_u0_u3_U322  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n747 ), .ZN(_AES_ENC_u0_u3_n793 ) );
NAND2_X2 _AES_ENC_u0_u3_U321  ( .A1(_AES_ENC_u0_u3_n584 ), .A2(_AES_ENC_u0_u3_n855 ), .ZN(_AES_ENC_u0_u3_n748 ) );
NAND2_X2 _AES_ENC_u0_u3_U320  ( .A1(_AES_ENC_u0_u3_n956 ), .A2(_AES_ENC_u0_u3_n748 ), .ZN(_AES_ENC_u0_u3_n760 ) );
NAND2_X2 _AES_ENC_u0_u3_U313  ( .A1(_AES_ENC_u0_u3_n590 ), .A2(_AES_ENC_u0_u3_n753 ), .ZN(_AES_ENC_u0_u3_n1023 ) );
NAND4_X2 _AES_ENC_u0_u3_U308  ( .A1(_AES_ENC_u0_u3_n760 ), .A2(_AES_ENC_u0_u3_n992 ), .A3(_AES_ENC_u0_u3_n759 ), .A4(_AES_ENC_u0_u3_n758 ), .ZN(_AES_ENC_u0_u3_n761 ) );
NAND2_X2 _AES_ENC_u0_u3_U307  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n761 ), .ZN(_AES_ENC_u0_u3_n792 ) );
NAND2_X2 _AES_ENC_u0_u3_U306  ( .A1(_AES_ENC_u0_u3_n584 ), .A2(_AES_ENC_u0_u3_n603 ), .ZN(_AES_ENC_u0_u3_n989 ) );
NAND2_X2 _AES_ENC_u0_u3_U305  ( .A1(_AES_ENC_u0_u3_n1050 ), .A2(_AES_ENC_u0_u3_n989 ), .ZN(_AES_ENC_u0_u3_n777 ) );
NAND2_X2 _AES_ENC_u0_u3_U304  ( .A1(_AES_ENC_u0_u3_n1093 ), .A2(_AES_ENC_u0_u3_n762 ), .ZN(_AES_ENC_u0_u3_n776 ) );
XNOR2_X2 _AES_ENC_u0_u3_U301  ( .A(_AES_ENC_w3[31] ), .B(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n959 ) );
NAND4_X2 _AES_ENC_u0_u3_U289  ( .A1(_AES_ENC_u0_u3_n777 ), .A2(_AES_ENC_u0_u3_n776 ), .A3(_AES_ENC_u0_u3_n775 ), .A4(_AES_ENC_u0_u3_n774 ), .ZN(_AES_ENC_u0_u3_n778 ) );
NAND2_X2 _AES_ENC_u0_u3_U288  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n778 ), .ZN(_AES_ENC_u0_u3_n791 ) );
NAND2_X2 _AES_ENC_u0_u3_U287  ( .A1(_AES_ENC_u0_u3_n1056 ), .A2(_AES_ENC_u0_u3_n1050 ), .ZN(_AES_ENC_u0_u3_n788 ) );
NAND2_X2 _AES_ENC_u0_u3_U286  ( .A1(_AES_ENC_u0_u3_n1091 ), .A2(_AES_ENC_u0_u3_n779 ), .ZN(_AES_ENC_u0_u3_n787 ) );
NAND2_X2 _AES_ENC_u0_u3_U285  ( .A1(_AES_ENC_u0_u3_n956 ), .A2(_AES_ENC_w3[25] ), .ZN(_AES_ENC_u0_u3_n786 ) );
NAND4_X2 _AES_ENC_u0_u3_U278  ( .A1(_AES_ENC_u0_u3_n788 ), .A2(_AES_ENC_u0_u3_n787 ), .A3(_AES_ENC_u0_u3_n786 ), .A4(_AES_ENC_u0_u3_n785 ), .ZN(_AES_ENC_u0_u3_n789 ) );
NAND2_X2 _AES_ENC_u0_u3_U277  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n789 ), .ZN(_AES_ENC_u0_u3_n790 ) );
NAND4_X2 _AES_ENC_u0_u3_U276  ( .A1(_AES_ENC_u0_u3_n793 ), .A2(_AES_ENC_u0_u3_n792 ), .A3(_AES_ENC_u0_u3_n791 ), .A4(_AES_ENC_u0_u3_n790 ), .ZN(_AES_ENC_u0_subword[2] ) );
NAND2_X2 _AES_ENC_u0_u3_U275  ( .A1(_AES_ENC_u0_u3_n1059 ), .A2(_AES_ENC_u0_u3_n794 ), .ZN(_AES_ENC_u0_u3_n810 ) );
NAND2_X2 _AES_ENC_u0_u3_U274  ( .A1(_AES_ENC_u0_u3_n1049 ), .A2(_AES_ENC_u0_u3_n956 ), .ZN(_AES_ENC_u0_u3_n809 ) );
OR2_X2 _AES_ENC_u0_u3_U266  ( .A1(_AES_ENC_u0_u3_n1096 ), .A2(_AES_ENC_u0_u3_n606 ), .ZN(_AES_ENC_u0_u3_n802 ) );
NAND2_X2 _AES_ENC_u0_u3_U265  ( .A1(_AES_ENC_u0_u3_n1053 ), .A2(_AES_ENC_u0_u3_n800 ), .ZN(_AES_ENC_u0_u3_n801 ) );
NAND2_X2 _AES_ENC_u0_u3_U264  ( .A1(_AES_ENC_u0_u3_n802 ), .A2(_AES_ENC_u0_u3_n801 ), .ZN(_AES_ENC_u0_u3_n805 ) );
NAND4_X2 _AES_ENC_u0_u3_U261  ( .A1(_AES_ENC_u0_u3_n810 ), .A2(_AES_ENC_u0_u3_n809 ), .A3(_AES_ENC_u0_u3_n808 ), .A4(_AES_ENC_u0_u3_n807 ), .ZN(_AES_ENC_u0_u3_n811 ) );
NAND2_X2 _AES_ENC_u0_u3_U260  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n811 ), .ZN(_AES_ENC_u0_u3_n852 ) );
OR2_X2 _AES_ENC_u0_u3_U259  ( .A1(_AES_ENC_u0_u3_n1023 ), .A2(_AES_ENC_u0_u3_n617 ), .ZN(_AES_ENC_u0_u3_n819 ) );
OR2_X2 _AES_ENC_u0_u3_U257  ( .A1(_AES_ENC_u0_u3_n570 ), .A2(_AES_ENC_u0_u3_n930 ), .ZN(_AES_ENC_u0_u3_n818 ) );
NAND2_X2 _AES_ENC_u0_u3_U256  ( .A1(_AES_ENC_u0_u3_n1013 ), .A2(_AES_ENC_u0_u3_n1094 ), .ZN(_AES_ENC_u0_u3_n817 ) );
NAND4_X2 _AES_ENC_u0_u3_U249  ( .A1(_AES_ENC_u0_u3_n819 ), .A2(_AES_ENC_u0_u3_n818 ), .A3(_AES_ENC_u0_u3_n817 ), .A4(_AES_ENC_u0_u3_n816 ), .ZN(_AES_ENC_u0_u3_n820 ) );
NAND2_X2 _AES_ENC_u0_u3_U248  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n820 ), .ZN(_AES_ENC_u0_u3_n851 ) );
NAND2_X2 _AES_ENC_u0_u3_U247  ( .A1(_AES_ENC_u0_u3_n956 ), .A2(_AES_ENC_u0_u3_n1080 ), .ZN(_AES_ENC_u0_u3_n835 ) );
NAND2_X2 _AES_ENC_u0_u3_U246  ( .A1(_AES_ENC_u0_u3_n570 ), .A2(_AES_ENC_u0_u3_n1030 ), .ZN(_AES_ENC_u0_u3_n1047 ) );
OR2_X2 _AES_ENC_u0_u3_U245  ( .A1(_AES_ENC_u0_u3_n1047 ), .A2(_AES_ENC_u0_u3_n612 ), .ZN(_AES_ENC_u0_u3_n834 ) );
NAND2_X2 _AES_ENC_u0_u3_U244  ( .A1(_AES_ENC_u0_u3_n1072 ), .A2(_AES_ENC_u0_u3_n589 ), .ZN(_AES_ENC_u0_u3_n833 ) );
NAND4_X2 _AES_ENC_u0_u3_U233  ( .A1(_AES_ENC_u0_u3_n835 ), .A2(_AES_ENC_u0_u3_n834 ), .A3(_AES_ENC_u0_u3_n833 ), .A4(_AES_ENC_u0_u3_n832 ), .ZN(_AES_ENC_u0_u3_n836 ) );
NAND2_X2 _AES_ENC_u0_u3_U232  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n836 ), .ZN(_AES_ENC_u0_u3_n850 ) );
NAND2_X2 _AES_ENC_u0_u3_U231  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n623 ), .ZN(_AES_ENC_u0_u3_n847 ) );
NAND2_X2 _AES_ENC_u0_u3_U230  ( .A1(_AES_ENC_u0_u3_n1050 ), .A2(_AES_ENC_u0_u3_n1071 ), .ZN(_AES_ENC_u0_u3_n846 ) );
OR2_X2 _AES_ENC_u0_u3_U224  ( .A1(_AES_ENC_u0_u3_n1053 ), .A2(_AES_ENC_u0_u3_n911 ), .ZN(_AES_ENC_u0_u3_n1077 ) );
NAND4_X2 _AES_ENC_u0_u3_U220  ( .A1(_AES_ENC_u0_u3_n847 ), .A2(_AES_ENC_u0_u3_n846 ), .A3(_AES_ENC_u0_u3_n845 ), .A4(_AES_ENC_u0_u3_n844 ), .ZN(_AES_ENC_u0_u3_n848 ) );
NAND2_X2 _AES_ENC_u0_u3_U219  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n848 ), .ZN(_AES_ENC_u0_u3_n849 ) );
NAND4_X2 _AES_ENC_u0_u3_U218  ( .A1(_AES_ENC_u0_u3_n852 ), .A2(_AES_ENC_u0_u3_n851 ), .A3(_AES_ENC_u0_u3_n850 ), .A4(_AES_ENC_u0_u3_n849 ), .ZN(_AES_ENC_u0_subword[3] ) );
NAND2_X2 _AES_ENC_u0_u3_U216  ( .A1(_AES_ENC_u0_u3_n1009 ), .A2(_AES_ENC_u0_u3_n1072 ), .ZN(_AES_ENC_u0_u3_n862 ) );
NAND2_X2 _AES_ENC_u0_u3_U215  ( .A1(_AES_ENC_u0_u3_n603 ), .A2(_AES_ENC_u0_u3_n577 ), .ZN(_AES_ENC_u0_u3_n853 ) );
NAND2_X2 _AES_ENC_u0_u3_U214  ( .A1(_AES_ENC_u0_u3_n1050 ), .A2(_AES_ENC_u0_u3_n853 ), .ZN(_AES_ENC_u0_u3_n861 ) );
NAND4_X2 _AES_ENC_u0_u3_U206  ( .A1(_AES_ENC_u0_u3_n862 ), .A2(_AES_ENC_u0_u3_n861 ), .A3(_AES_ENC_u0_u3_n860 ), .A4(_AES_ENC_u0_u3_n859 ), .ZN(_AES_ENC_u0_u3_n863 ) );
NAND2_X2 _AES_ENC_u0_u3_U205  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n863 ), .ZN(_AES_ENC_u0_u3_n905 ) );
NAND2_X2 _AES_ENC_u0_u3_U204  ( .A1(_AES_ENC_u0_u3_n1010 ), .A2(_AES_ENC_u0_u3_n989 ), .ZN(_AES_ENC_u0_u3_n874 ) );
NAND2_X2 _AES_ENC_u0_u3_U203  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n610 ), .ZN(_AES_ENC_u0_u3_n864 ) );
NAND2_X2 _AES_ENC_u0_u3_U202  ( .A1(_AES_ENC_u0_u3_n929 ), .A2(_AES_ENC_u0_u3_n864 ), .ZN(_AES_ENC_u0_u3_n873 ) );
NAND4_X2 _AES_ENC_u0_u3_U193  ( .A1(_AES_ENC_u0_u3_n874 ), .A2(_AES_ENC_u0_u3_n873 ), .A3(_AES_ENC_u0_u3_n872 ), .A4(_AES_ENC_u0_u3_n871 ), .ZN(_AES_ENC_u0_u3_n875 ) );
NAND2_X2 _AES_ENC_u0_u3_U192  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n875 ), .ZN(_AES_ENC_u0_u3_n904 ) );
NAND2_X2 _AES_ENC_u0_u3_U191  ( .A1(_AES_ENC_u0_u3_n583 ), .A2(_AES_ENC_u0_u3_n1050 ), .ZN(_AES_ENC_u0_u3_n889 ) );
NAND2_X2 _AES_ENC_u0_u3_U190  ( .A1(_AES_ENC_u0_u3_n1093 ), .A2(_AES_ENC_u0_u3_n587 ), .ZN(_AES_ENC_u0_u3_n876 ) );
NAND2_X2 _AES_ENC_u0_u3_U189  ( .A1(_AES_ENC_u0_u3_n604 ), .A2(_AES_ENC_u0_u3_n876 ), .ZN(_AES_ENC_u0_u3_n877 ) );
NAND2_X2 _AES_ENC_u0_u3_U188  ( .A1(_AES_ENC_u0_u3_n877 ), .A2(_AES_ENC_u0_u3_n623 ), .ZN(_AES_ENC_u0_u3_n888 ) );
NAND4_X2 _AES_ENC_u0_u3_U179  ( .A1(_AES_ENC_u0_u3_n889 ), .A2(_AES_ENC_u0_u3_n888 ), .A3(_AES_ENC_u0_u3_n887 ), .A4(_AES_ENC_u0_u3_n886 ), .ZN(_AES_ENC_u0_u3_n890 ) );
NAND2_X2 _AES_ENC_u0_u3_U178  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n890 ), .ZN(_AES_ENC_u0_u3_n903 ) );
OR2_X2 _AES_ENC_u0_u3_U177  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n1059 ), .ZN(_AES_ENC_u0_u3_n900 ) );
NAND2_X2 _AES_ENC_u0_u3_U176  ( .A1(_AES_ENC_u0_u3_n1073 ), .A2(_AES_ENC_u0_u3_n1047 ), .ZN(_AES_ENC_u0_u3_n899 ) );
NAND2_X2 _AES_ENC_u0_u3_U175  ( .A1(_AES_ENC_u0_u3_n1094 ), .A2(_AES_ENC_u0_u3_n595 ), .ZN(_AES_ENC_u0_u3_n898 ) );
NAND4_X2 _AES_ENC_u0_u3_U167  ( .A1(_AES_ENC_u0_u3_n900 ), .A2(_AES_ENC_u0_u3_n899 ), .A3(_AES_ENC_u0_u3_n898 ), .A4(_AES_ENC_u0_u3_n897 ), .ZN(_AES_ENC_u0_u3_n901 ) );
NAND2_X2 _AES_ENC_u0_u3_U166  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n901 ), .ZN(_AES_ENC_u0_u3_n902 ) );
NAND4_X2 _AES_ENC_u0_u3_U165  ( .A1(_AES_ENC_u0_u3_n905 ), .A2(_AES_ENC_u0_u3_n904 ), .A3(_AES_ENC_u0_u3_n903 ), .A4(_AES_ENC_u0_u3_n902 ), .ZN(_AES_ENC_u0_subword[4] ) );
NAND2_X2 _AES_ENC_u0_u3_U164  ( .A1(_AES_ENC_u0_u3_n1094 ), .A2(_AES_ENC_u0_u3_n599 ), .ZN(_AES_ENC_u0_u3_n922 ) );
NAND2_X2 _AES_ENC_u0_u3_U163  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n989 ), .ZN(_AES_ENC_u0_u3_n921 ) );
NAND4_X2 _AES_ENC_u0_u3_U151  ( .A1(_AES_ENC_u0_u3_n922 ), .A2(_AES_ENC_u0_u3_n921 ), .A3(_AES_ENC_u0_u3_n920 ), .A4(_AES_ENC_u0_u3_n919 ), .ZN(_AES_ENC_u0_u3_n923 ) );
NAND2_X2 _AES_ENC_u0_u3_U150  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n923 ), .ZN(_AES_ENC_u0_u3_n972 ) );
NAND2_X2 _AES_ENC_u0_u3_U149  ( .A1(_AES_ENC_u0_u3_n582 ), .A2(_AES_ENC_u0_u3_n619 ), .ZN(_AES_ENC_u0_u3_n924 ) );
NAND2_X2 _AES_ENC_u0_u3_U148  ( .A1(_AES_ENC_u0_u3_n1073 ), .A2(_AES_ENC_u0_u3_n924 ), .ZN(_AES_ENC_u0_u3_n939 ) );
NAND2_X2 _AES_ENC_u0_u3_U147  ( .A1(_AES_ENC_u0_u3_n926 ), .A2(_AES_ENC_u0_u3_n925 ), .ZN(_AES_ENC_u0_u3_n927 ) );
NAND2_X2 _AES_ENC_u0_u3_U146  ( .A1(_AES_ENC_u0_u3_n606 ), .A2(_AES_ENC_u0_u3_n927 ), .ZN(_AES_ENC_u0_u3_n928 ) );
NAND2_X2 _AES_ENC_u0_u3_U145  ( .A1(_AES_ENC_u0_u3_n928 ), .A2(_AES_ENC_u0_u3_n1080 ), .ZN(_AES_ENC_u0_u3_n938 ) );
OR2_X2 _AES_ENC_u0_u3_U144  ( .A1(_AES_ENC_u0_u3_n1117 ), .A2(_AES_ENC_u0_u3_n615 ), .ZN(_AES_ENC_u0_u3_n937 ) );
NAND4_X2 _AES_ENC_u0_u3_U139  ( .A1(_AES_ENC_u0_u3_n939 ), .A2(_AES_ENC_u0_u3_n938 ), .A3(_AES_ENC_u0_u3_n937 ), .A4(_AES_ENC_u0_u3_n936 ), .ZN(_AES_ENC_u0_u3_n940 ) );
NAND2_X2 _AES_ENC_u0_u3_U138  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n940 ), .ZN(_AES_ENC_u0_u3_n971 ) );
OR2_X2 _AES_ENC_u0_u3_U137  ( .A1(_AES_ENC_u0_u3_n605 ), .A2(_AES_ENC_u0_u3_n941 ), .ZN(_AES_ENC_u0_u3_n954 ) );
NAND2_X2 _AES_ENC_u0_u3_U136  ( .A1(_AES_ENC_u0_u3_n1096 ), .A2(_AES_ENC_u0_u3_n577 ), .ZN(_AES_ENC_u0_u3_n942 ) );
NAND2_X2 _AES_ENC_u0_u3_U135  ( .A1(_AES_ENC_u0_u3_n1048 ), .A2(_AES_ENC_u0_u3_n942 ), .ZN(_AES_ENC_u0_u3_n943 ) );
NAND2_X2 _AES_ENC_u0_u3_U134  ( .A1(_AES_ENC_u0_u3_n612 ), .A2(_AES_ENC_u0_u3_n943 ), .ZN(_AES_ENC_u0_u3_n944 ) );
NAND2_X2 _AES_ENC_u0_u3_U133  ( .A1(_AES_ENC_u0_u3_n944 ), .A2(_AES_ENC_u0_u3_n580 ), .ZN(_AES_ENC_u0_u3_n953 ) );
NAND4_X2 _AES_ENC_u0_u3_U125  ( .A1(_AES_ENC_u0_u3_n954 ), .A2(_AES_ENC_u0_u3_n953 ), .A3(_AES_ENC_u0_u3_n952 ), .A4(_AES_ENC_u0_u3_n951 ), .ZN(_AES_ENC_u0_u3_n955 ) );
NAND2_X2 _AES_ENC_u0_u3_U124  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n955 ), .ZN(_AES_ENC_u0_u3_n970 ) );
NAND2_X2 _AES_ENC_u0_u3_U123  ( .A1(_AES_ENC_u0_u3_n1094 ), .A2(_AES_ENC_u0_u3_n1071 ), .ZN(_AES_ENC_u0_u3_n967 ) );
NAND2_X2 _AES_ENC_u0_u3_U122  ( .A1(_AES_ENC_u0_u3_n956 ), .A2(_AES_ENC_u0_u3_n1030 ), .ZN(_AES_ENC_u0_u3_n966 ) );
NAND4_X2 _AES_ENC_u0_u3_U114  ( .A1(_AES_ENC_u0_u3_n967 ), .A2(_AES_ENC_u0_u3_n966 ), .A3(_AES_ENC_u0_u3_n965 ), .A4(_AES_ENC_u0_u3_n964 ), .ZN(_AES_ENC_u0_u3_n968 ) );
NAND2_X2 _AES_ENC_u0_u3_U113  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n968 ), .ZN(_AES_ENC_u0_u3_n969 ) );
NAND4_X2 _AES_ENC_u0_u3_U112  ( .A1(_AES_ENC_u0_u3_n972 ), .A2(_AES_ENC_u0_u3_n971 ), .A3(_AES_ENC_u0_u3_n970 ), .A4(_AES_ENC_u0_u3_n969 ), .ZN(_AES_ENC_u0_subword[5] ) );
NAND2_X2 _AES_ENC_u0_u3_U111  ( .A1(_AES_ENC_u0_u3_n570 ), .A2(_AES_ENC_u0_u3_n1097 ), .ZN(_AES_ENC_u0_u3_n973 ) );
NAND2_X2 _AES_ENC_u0_u3_U110  ( .A1(_AES_ENC_u0_u3_n1073 ), .A2(_AES_ENC_u0_u3_n973 ), .ZN(_AES_ENC_u0_u3_n987 ) );
NAND2_X2 _AES_ENC_u0_u3_U109  ( .A1(_AES_ENC_u0_u3_n974 ), .A2(_AES_ENC_u0_u3_n1077 ), .ZN(_AES_ENC_u0_u3_n975 ) );
NAND2_X2 _AES_ENC_u0_u3_U108  ( .A1(_AES_ENC_u0_u3_n613 ), .A2(_AES_ENC_u0_u3_n975 ), .ZN(_AES_ENC_u0_u3_n976 ) );
NAND2_X2 _AES_ENC_u0_u3_U107  ( .A1(_AES_ENC_u0_u3_n977 ), .A2(_AES_ENC_u0_u3_n976 ), .ZN(_AES_ENC_u0_u3_n986 ) );
NAND4_X2 _AES_ENC_u0_u3_U99  ( .A1(_AES_ENC_u0_u3_n987 ), .A2(_AES_ENC_u0_u3_n986 ), .A3(_AES_ENC_u0_u3_n985 ), .A4(_AES_ENC_u0_u3_n984 ), .ZN(_AES_ENC_u0_u3_n988 ) );
NAND2_X2 _AES_ENC_u0_u3_U98  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n988 ), .ZN(_AES_ENC_u0_u3_n1044 ) );
NAND2_X2 _AES_ENC_u0_u3_U97  ( .A1(_AES_ENC_u0_u3_n1073 ), .A2(_AES_ENC_u0_u3_n989 ), .ZN(_AES_ENC_u0_u3_n1004 ) );
NAND2_X2 _AES_ENC_u0_u3_U96  ( .A1(_AES_ENC_u0_u3_n1092 ), .A2(_AES_ENC_u0_u3_n619 ), .ZN(_AES_ENC_u0_u3_n1003 ) );
NAND4_X2 _AES_ENC_u0_u3_U85  ( .A1(_AES_ENC_u0_u3_n1004 ), .A2(_AES_ENC_u0_u3_n1003 ), .A3(_AES_ENC_u0_u3_n1002 ), .A4(_AES_ENC_u0_u3_n1001 ), .ZN(_AES_ENC_u0_u3_n1005 ) );
NAND2_X2 _AES_ENC_u0_u3_U84  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n1005 ), .ZN(_AES_ENC_u0_u3_n1043 ) );
NAND2_X2 _AES_ENC_u0_u3_U83  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n596 ), .ZN(_AES_ENC_u0_u3_n1020 ) );
NAND2_X2 _AES_ENC_u0_u3_U82  ( .A1(_AES_ENC_u0_u3_n1050 ), .A2(_AES_ENC_u0_u3_n624 ), .ZN(_AES_ENC_u0_u3_n1019 ) );
NAND2_X2 _AES_ENC_u0_u3_U77  ( .A1(_AES_ENC_u0_u3_n1059 ), .A2(_AES_ENC_u0_u3_n1114 ), .ZN(_AES_ENC_u0_u3_n1012 ) );
NAND2_X2 _AES_ENC_u0_u3_U76  ( .A1(_AES_ENC_u0_u3_n1010 ), .A2(_AES_ENC_u0_u3_n592 ), .ZN(_AES_ENC_u0_u3_n1011 ) );
NAND2_X2 _AES_ENC_u0_u3_U75  ( .A1(_AES_ENC_u0_u3_n1012 ), .A2(_AES_ENC_u0_u3_n1011 ), .ZN(_AES_ENC_u0_u3_n1016 ) );
NAND4_X2 _AES_ENC_u0_u3_U70  ( .A1(_AES_ENC_u0_u3_n1020 ), .A2(_AES_ENC_u0_u3_n1019 ), .A3(_AES_ENC_u0_u3_n1018 ), .A4(_AES_ENC_u0_u3_n1017 ), .ZN(_AES_ENC_u0_u3_n1021 ) );
NAND2_X2 _AES_ENC_u0_u3_U69  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n1021 ), .ZN(_AES_ENC_u0_u3_n1042 ) );
NAND2_X2 _AES_ENC_u0_u3_U68  ( .A1(_AES_ENC_u0_u3_n1022 ), .A2(_AES_ENC_u0_u3_n1093 ), .ZN(_AES_ENC_u0_u3_n1039 ) );
NAND2_X2 _AES_ENC_u0_u3_U67  ( .A1(_AES_ENC_u0_u3_n1050 ), .A2(_AES_ENC_u0_u3_n1023 ), .ZN(_AES_ENC_u0_u3_n1038 ) );
NAND2_X2 _AES_ENC_u0_u3_U66  ( .A1(_AES_ENC_u0_u3_n1024 ), .A2(_AES_ENC_u0_u3_n1071 ), .ZN(_AES_ENC_u0_u3_n1037 ) );
AND2_X2 _AES_ENC_u0_u3_U60  ( .A1(_AES_ENC_u0_u3_n1030 ), .A2(_AES_ENC_u0_u3_n602 ), .ZN(_AES_ENC_u0_u3_n1078 ) );
NAND4_X2 _AES_ENC_u0_u3_U56  ( .A1(_AES_ENC_u0_u3_n1039 ), .A2(_AES_ENC_u0_u3_n1038 ), .A3(_AES_ENC_u0_u3_n1037 ), .A4(_AES_ENC_u0_u3_n1036 ), .ZN(_AES_ENC_u0_u3_n1040 ) );
NAND2_X2 _AES_ENC_u0_u3_U55  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n1040 ), .ZN(_AES_ENC_u0_u3_n1041 ) );
NAND4_X2 _AES_ENC_u0_u3_U54  ( .A1(_AES_ENC_u0_u3_n1044 ), .A2(_AES_ENC_u0_u3_n1043 ), .A3(_AES_ENC_u0_u3_n1042 ), .A4(_AES_ENC_u0_u3_n1041 ), .ZN(_AES_ENC_u0_subword[6] ) );
NAND2_X2 _AES_ENC_u0_u3_U53  ( .A1(_AES_ENC_u0_u3_n1072 ), .A2(_AES_ENC_u0_u3_n1045 ), .ZN(_AES_ENC_u0_u3_n1068 ) );
NAND2_X2 _AES_ENC_u0_u3_U52  ( .A1(_AES_ENC_u0_u3_n1046 ), .A2(_AES_ENC_u0_u3_n582 ), .ZN(_AES_ENC_u0_u3_n1067 ) );
NAND2_X2 _AES_ENC_u0_u3_U51  ( .A1(_AES_ENC_u0_u3_n1094 ), .A2(_AES_ENC_u0_u3_n1047 ), .ZN(_AES_ENC_u0_u3_n1066 ) );
NAND4_X2 _AES_ENC_u0_u3_U40  ( .A1(_AES_ENC_u0_u3_n1068 ), .A2(_AES_ENC_u0_u3_n1067 ), .A3(_AES_ENC_u0_u3_n1066 ), .A4(_AES_ENC_u0_u3_n1065 ), .ZN(_AES_ENC_u0_u3_n1069 ) );
NAND2_X2 _AES_ENC_u0_u3_U39  ( .A1(_AES_ENC_u0_u3_n1070 ), .A2(_AES_ENC_u0_u3_n1069 ), .ZN(_AES_ENC_u0_u3_n1135 ) );
NAND2_X2 _AES_ENC_u0_u3_U38  ( .A1(_AES_ENC_u0_u3_n1072 ), .A2(_AES_ENC_u0_u3_n1071 ), .ZN(_AES_ENC_u0_u3_n1088 ) );
NAND2_X2 _AES_ENC_u0_u3_U37  ( .A1(_AES_ENC_u0_u3_n1073 ), .A2(_AES_ENC_u0_u3_n595 ), .ZN(_AES_ENC_u0_u3_n1087 ) );
NAND4_X2 _AES_ENC_u0_u3_U28  ( .A1(_AES_ENC_u0_u3_n1088 ), .A2(_AES_ENC_u0_u3_n1087 ), .A3(_AES_ENC_u0_u3_n1086 ), .A4(_AES_ENC_u0_u3_n1085 ), .ZN(_AES_ENC_u0_u3_n1089 ) );
NAND2_X2 _AES_ENC_u0_u3_U27  ( .A1(_AES_ENC_u0_u3_n1090 ), .A2(_AES_ENC_u0_u3_n1089 ), .ZN(_AES_ENC_u0_u3_n1134 ) );
NAND2_X2 _AES_ENC_u0_u3_U26  ( .A1(_AES_ENC_u0_u3_n1091 ), .A2(_AES_ENC_u0_u3_n1093 ), .ZN(_AES_ENC_u0_u3_n1111 ) );
NAND2_X2 _AES_ENC_u0_u3_U25  ( .A1(_AES_ENC_u0_u3_n1092 ), .A2(_AES_ENC_u0_u3_n1120 ), .ZN(_AES_ENC_u0_u3_n1110 ) );
AND2_X2 _AES_ENC_u0_u3_U22  ( .A1(_AES_ENC_u0_u3_n1097 ), .A2(_AES_ENC_u0_u3_n1096 ), .ZN(_AES_ENC_u0_u3_n1098 ) );
NAND4_X2 _AES_ENC_u0_u3_U14  ( .A1(_AES_ENC_u0_u3_n1111 ), .A2(_AES_ENC_u0_u3_n1110 ), .A3(_AES_ENC_u0_u3_n1109 ), .A4(_AES_ENC_u0_u3_n1108 ), .ZN(_AES_ENC_u0_u3_n1112 ) );
NAND2_X2 _AES_ENC_u0_u3_U13  ( .A1(_AES_ENC_u0_u3_n1113 ), .A2(_AES_ENC_u0_u3_n1112 ), .ZN(_AES_ENC_u0_u3_n1133 ) );
NAND2_X2 _AES_ENC_u0_u3_U12  ( .A1(_AES_ENC_u0_u3_n1115 ), .A2(_AES_ENC_u0_u3_n1114 ), .ZN(_AES_ENC_u0_u3_n1129 ) );
OR2_X2 _AES_ENC_u0_u3_U11  ( .A1(_AES_ENC_u0_u3_n608 ), .A2(_AES_ENC_u0_u3_n1116 ), .ZN(_AES_ENC_u0_u3_n1128 ) );
NAND4_X2 _AES_ENC_u0_u3_U3  ( .A1(_AES_ENC_u0_u3_n1129 ), .A2(_AES_ENC_u0_u3_n1128 ), .A3(_AES_ENC_u0_u3_n1127 ), .A4(_AES_ENC_u0_u3_n1126 ), .ZN(_AES_ENC_u0_u3_n1130 ) );
NAND2_X2 _AES_ENC_u0_u3_U2  ( .A1(_AES_ENC_u0_u3_n1131 ), .A2(_AES_ENC_u0_u3_n1130 ), .ZN(_AES_ENC_u0_u3_n1132 ) );
NAND4_X2 _AES_ENC_u0_u3_U1  ( .A1(_AES_ENC_u0_u3_n1135 ), .A2(_AES_ENC_u0_u3_n1134 ), .A3(_AES_ENC_u0_u3_n1133 ), .A4(_AES_ENC_u0_u3_n1132 ), .ZN(_AES_ENC_u0_subword[7] ) );
INV_X4 _AES_ENC_u0_r0_U41  ( .A(_AES_ENC_u0_r0_n32 ), .ZN(_AES_ENC_u0_r0_n38 ) );
INV_X4 _AES_ENC_u0_r0_U40  ( .A(_AES_ENC_u0_r0_n9 ), .ZN(_AES_ENC_u0_r0_n37 ) );
INV_X4 _AES_ENC_u0_r0_U39  ( .A(_AES_ENC_u0_r0_n11 ), .ZN(_AES_ENC_u0_r0_n36 ) );
NAND3_X2 _AES_ENC_u0_r0_U38  ( .A1(_AES_ENC_u0_r0_rcnt[0] ), .A2(_AES_ENC_u0_r0_n35 ), .A3(_AES_ENC_u0_r0_n17 ), .ZN(_AES_ENC_u0_r0_n19 ) );
NOR3_X2 _AES_ENC_u0_r0_U27  ( .A1(_AES_ENC_u0_r0_n38 ), .A2(_AES_ENC_u0_r0_n13 ), .A3(_AES_ENC_u0_r0_n36 ), .ZN(_AES_ENC_u0_r0_N49 ) );
NAND3_X2 _AES_ENC_u0_r0_U24  ( .A1(_AES_ENC_u0_r0_n16 ), .A2(_AES_ENC_u0_r0_rcnt[0] ), .A3(_AES_ENC_u0_r0_N54 ), .ZN(_AES_ENC_u0_r0_n12 ) );
NOR2_X2 _AES_ENC_u0_r0_U23  ( .A1(_AES_ENC_u0_n315 ), .A2(_AES_ENC_u0_r0_rcnt[0] ), .ZN(_AES_ENC_u0_r0_n32 ) );
NOR2_X2 _AES_ENC_u0_r0_U22  ( .A1(_AES_ENC_u0_r0_n24 ), .A2(_AES_ENC_u0_r0_n34 ), .ZN(_AES_ENC_u0_r0_n22 ) );
NOR2_X2 _AES_ENC_u0_r0_U20  ( .A1(_AES_ENC_u0_r0_n22 ), .A2(_AES_ENC_u0_r0_n23 ), .ZN(_AES_ENC_u0_r0_n9 ) );
NOR2_X2 _AES_ENC_u0_r0_U15  ( .A1(_AES_ENC_u0_r0_n11 ), .A2(_AES_ENC_u0_r0_n12 ), .ZN(_AES_ENC_u0_r0_N50 ) );
NOR2_X2 _AES_ENC_u0_r0_U12  ( .A1(_AES_ENC_u0_r0_n11 ), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_r0_N53 ) );
NOR3_X2 _AES_ENC_u0_r0_U11  ( .A1(_AES_ENC_u0_r0_n16 ), .A2(_AES_ENC_u0_r0_n9 ), .A3(_AES_ENC_u0_r0_n36 ), .ZN(_AES_ENC_u0_r0_n17 ) );
NOR2_X2 _AES_ENC_u0_r0_U7  ( .A1(_AES_ENC_u0_r0_n37 ), .A2(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_r0_N54 ) );
INV_X4 _AES_ENC_u0_r0_U6  ( .A(_AES_ENC_u0_n315 ), .ZN(_AES_ENC_u0_r0_n35 ));
XNOR2_X2 _AES_ENC_u0_r0_U37  ( .A(_AES_ENC_u0_r0_rcnt[1] ), .B(_AES_ENC_u0_r0_rcnt[0] ), .ZN(_AES_ENC_u0_r0_n11 ) );
XOR2_X2 _AES_ENC_u0_r0_U36  ( .A(_AES_ENC_u0_r0_n34 ), .B(_AES_ENC_u0_r0_n11 ), .Z(_AES_ENC_u0_r0_n26 ) );
NAND2_X2 _AES_ENC_u0_r0_U35  ( .A1(_AES_ENC_u0_r0_rcnt[0] ), .A2(_AES_ENC_u0_r0_rcnt[1] ), .ZN(_AES_ENC_u0_r0_n24 ) );
NAND2_X2 _AES_ENC_u0_r0_U34  ( .A1(_AES_ENC_u0_r0_rcnt[2] ), .A2(_AES_ENC_u0_r0_n36 ), .ZN(_AES_ENC_u0_r0_n29 ) );
NAND2_X2 _AES_ENC_u0_r0_U33  ( .A1(_AES_ENC_u0_r0_n24 ), .A2(_AES_ENC_u0_r0_n29 ), .ZN(_AES_ENC_u0_r0_n27 ) );
NAND2_X2 _AES_ENC_u0_r0_U32  ( .A1(_AES_ENC_u0_r0_n26 ), .A2(_AES_ENC_u0_r0_n27 ), .ZN(_AES_ENC_u0_r0_n28 ) );
NAND2_X2 _AES_ENC_u0_r0_U31  ( .A1(_AES_ENC_u0_r0_n35 ), .A2(_AES_ENC_u0_r0_n28 ), .ZN(_AES_ENC_u0_r0_N44 ) );
NAND4_X2 _AES_ENC_u0_r0_U30  ( .A1(_AES_ENC_u0_r0_n26 ), .A2(_AES_ENC_u0_r0_n27 ), .A3(_AES_ENC_u0_r0_n35 ), .A4(_AES_ENC_u0_r0_n33 ), .ZN(_AES_ENC_u0_r0_n7 ) );
OR3_X2 _AES_ENC_u0_r0_U29  ( .A1(_AES_ENC_u0_r0_n26 ), .A2(_AES_ENC_u0_n315 ), .A3(_AES_ENC_u0_r0_n27 ), .ZN(_AES_ENC_u0_r0_n25 ) );
NAND2_X2 _AES_ENC_u0_r0_U28  ( .A1(_AES_ENC_u0_r0_n7 ), .A2(_AES_ENC_u0_r0_n25 ), .ZN(_AES_ENC_u0_r0_N45 ) );
XOR2_X2 _AES_ENC_u0_r0_U26  ( .A(_AES_ENC_u0_r0_n33 ), .B(_AES_ENC_u0_r0_n22 ), .Z(_AES_ENC_u0_r0_n16 ) );
AND2_X2 _AES_ENC_u0_r0_U25  ( .A1(_AES_ENC_u0_r0_n24 ), .A2(_AES_ENC_u0_r0_n34 ), .ZN(_AES_ENC_u0_r0_n23 ) );
NAND2_X2 _AES_ENC_u0_r0_U21  ( .A1(_AES_ENC_u0_r0_n17 ), .A2(_AES_ENC_u0_r0_n32 ), .ZN(_AES_ENC_u0_r0_n20 ) );
NAND4_X2 _AES_ENC_u0_r0_U19  ( .A1(_AES_ENC_u0_r0_n16 ), .A2(_AES_ENC_u0_r0_N53 ), .A3(_AES_ENC_u0_r0_rcnt[0] ), .A4(_AES_ENC_u0_r0_n37 ), .ZN(_AES_ENC_u0_r0_n21 ) );
NAND2_X2 _AES_ENC_u0_r0_U18  ( .A1(_AES_ENC_u0_r0_n20 ), .A2(_AES_ENC_u0_r0_n21 ), .ZN(_AES_ENC_u0_r0_N46 ) );
AND3_X2 _AES_ENC_u0_r0_U17  ( .A1(_AES_ENC_u0_r0_n16 ), .A2(_AES_ENC_u0_r0_n36 ), .A3(_AES_ENC_u0_r0_n32 ), .ZN(_AES_ENC_u0_r0_n10 ) );
NAND2_X2 _AES_ENC_u0_r0_U16  ( .A1(_AES_ENC_u0_r0_n10 ), .A2(_AES_ENC_u0_r0_n37 ), .ZN(_AES_ENC_u0_r0_n18 ) );
NAND2_X2 _AES_ENC_u0_r0_U14  ( .A1(_AES_ENC_u0_r0_n18 ), .A2(_AES_ENC_u0_r0_n19 ), .ZN(_AES_ENC_u0_r0_N47 ) );
NAND2_X2 _AES_ENC_u0_r0_U13  ( .A1(_AES_ENC_u0_r0_n17 ), .A2(_AES_ENC_u0_r0_n35 ), .ZN(_AES_ENC_u0_r0_n14 ) );
OR2_X2 _AES_ENC_u0_r0_U10  ( .A1(_AES_ENC_u0_r0_n12 ), .A2(_AES_ENC_u0_r0_n36 ), .ZN(_AES_ENC_u0_r0_n15 ) );
NAND2_X2 _AES_ENC_u0_r0_U9  ( .A1(_AES_ENC_u0_r0_n14 ), .A2(_AES_ENC_u0_r0_n15 ), .ZN(_AES_ENC_u0_r0_N48 ) );
XOR2_X2 _AES_ENC_u0_r0_U8  ( .A(_AES_ENC_u0_r0_n33 ), .B(_AES_ENC_u0_r0_rcnt[2] ), .Z(_AES_ENC_u0_r0_n13 ) );
AND2_X2 _AES_ENC_u0_r0_U5  ( .A1(_AES_ENC_u0_r0_n9 ), .A2(_AES_ENC_u0_r0_n10 ), .ZN(_AES_ENC_u0_r0_N51 ) );
OR2_X2 _AES_ENC_u0_r0_U4  ( .A1(_AES_ENC_u0_r0_n33 ), .A2(_AES_ENC_u0_r0_N44 ), .ZN(_AES_ENC_u0_r0_n8 ) );
NAND2_X2 _AES_ENC_u0_r0_U3  ( .A1(_AES_ENC_u0_r0_n7 ), .A2(_AES_ENC_u0_r0_n8 ), .ZN(_AES_ENC_u0_r0_N55 ) );
CLKBUFX1 gbuf_d_1294(.A(_AES_ENC_u0_r0_N45), .Y(ddout__1294));
CLKBUFX1 gbuf_q_1294(.A(qq_in1294), .Y(_AES_ENC_u0_rcon[25]));
CLKBUFX1 gbuf_d_1295(.A(_AES_ENC_u0_r0_N46), .Y(ddout__1295));
CLKBUFX1 gbuf_q_1295(.A(qq_in1295), .Y(_AES_ENC_u0_rcon[26]));
CLKBUFX1 gbuf_d_1296(.A(_AES_ENC_u0_r0_N47), .Y(ddout__1296));
CLKBUFX1 gbuf_q_1296(.A(qq_in1296), .Y(_AES_ENC_u0_rcon[27]));
CLKBUFX1 gbuf_d_1297(.A(_AES_ENC_u0_r0_N48), .Y(ddout__1297));
CLKBUFX1 gbuf_q_1297(.A(qq_in1297), .Y(_AES_ENC_u0_rcon[28]));
CLKBUFX1 gbuf_d_1298(.A(_AES_ENC_u0_r0_N50), .Y(ddout__1298));
CLKBUFX1 gbuf_q_1298(.A(qq_in1298), .Y(_AES_ENC_u0_rcon[30]));
CLKBUFX1 gbuf_d_1299(.A(_AES_ENC_u0_r0_N49), .Y(ddout__1299));
CLKBUFX1 gbuf_q_1299(.A(qq_in1299), .Y(_AES_ENC_u0_rcon[29]));
CLKBUFX1 gbuf_d_1300(.A(_AES_ENC_u0_r0_N51), .Y(ddout__1300));
CLKBUFX1 gbuf_q_1300(.A(qq_in1300), .Y(_AES_ENC_u0_rcon[31]));
CLKBUFX1 gbuf_d_1301(.A(_AES_ENC_u0_r0_N55), .Y(ddout__1301));
CLKBUFX1 gbuf_qn_1301(.A(qnn_in_1301), .Y(_AES_ENC_u0_r0_n33));
CLKBUFX1 gbuf_d_1302(.A(_AES_ENC_u0_r0_N44), .Y(ddout__1302));
CLKBUFX1 gbuf_q_1302(.A(qq_in1302), .Y(_AES_ENC_u0_rcon[24]));
CLKBUFX1 gbuf_d_1303(.A(_AES_ENC_u0_r0_N54), .Y(ddout__1303));
CLKBUFX1 gbuf_q_1303(.A(qq_in1303), .Y(_AES_ENC_u0_r0_rcnt[2]));
CLKBUFX1 gbuf_qn_1303(.A(qnn_in_1303), .Y(_AES_ENC_u0_r0_n34));
CLKBUFX1 gbuf_d_1304(.A(_AES_ENC_u0_r0_N53), .Y(ddout__1304));
CLKBUFX1 gbuf_q_1304(.A(qq_in1304), .Y(_AES_ENC_u0_r0_rcnt[1]));
CLKBUFX1 gbuf_d_1305(.A(_AES_ENC_u0_r0_n32), .Y(ddout__1305));
CLKBUFX1 gbuf_q_1305(.A(qq_in1305), .Y(_AES_ENC_u0_r0_rcnt[0]));
INV_X4 _AES_ENC_us00_U575  ( .A(_AES_ENC_sa00[7]), .ZN(_AES_ENC_us00_n627 ));
INV_X4 _AES_ENC_us00_U574  ( .A(_AES_ENC_us00_n79 ), .ZN(_AES_ENC_us00_n625 ) );
INV_X4 _AES_ENC_us00_U573  ( .A(_AES_ENC_sa00[4]), .ZN(_AES_ENC_us00_n624 ));
INV_X4 _AES_ENC_us00_U572  ( .A(_AES_ENC_us00_n170 ), .ZN(_AES_ENC_us00_n622 ) );
INV_X4 _AES_ENC_us00_U571  ( .A(_AES_ENC_us00_n73 ), .ZN(_AES_ENC_us00_n620 ) );
INV_X4 _AES_ENC_us00_U570  ( .A(_AES_ENC_us00_n72 ), .ZN(_AES_ENC_us00_n619 ) );
INV_X4 _AES_ENC_us00_U569  ( .A(_AES_ENC_us00_n146 ), .ZN(_AES_ENC_us00_n618 ) );
INV_X4 _AES_ENC_us00_U568  ( .A(_AES_ENC_us00_n221 ), .ZN(_AES_ENC_us00_n616 ) );
INV_X4 _AES_ENC_us00_U567  ( .A(_AES_ENC_us00_n402 ), .ZN(_AES_ENC_us00_n614 ) );
INV_X4 _AES_ENC_us00_U566  ( .A(_AES_ENC_sa00[2]), .ZN(_AES_ENC_us00_n611 ));
INV_X4 _AES_ENC_us00_U565  ( .A(_AES_ENC_us00_n396 ), .ZN(_AES_ENC_us00_n610 ) );
INV_X4 _AES_ENC_us00_U564  ( .A(_AES_ENC_us00_n271 ), .ZN(_AES_ENC_us00_n609 ) );
INV_X4 _AES_ENC_us00_U563  ( .A(_AES_ENC_us00_n417 ), .ZN(_AES_ENC_us00_n607 ) );
INV_X4 _AES_ENC_us00_U562  ( .A(_AES_ENC_us00_n173 ), .ZN(_AES_ENC_us00_n603 ) );
INV_X4 _AES_ENC_us00_U561  ( .A(_AES_ENC_us00_n91 ), .ZN(_AES_ENC_us00_n602 ) );
INV_X4 _AES_ENC_us00_U560  ( .A(_AES_ENC_us00_n267 ), .ZN(_AES_ENC_us00_n601 ) );
INV_X4 _AES_ENC_us00_U559  ( .A(_AES_ENC_us00_n138 ), .ZN(_AES_ENC_us00_n600 ) );
INV_X4 _AES_ENC_us00_U558  ( .A(_AES_ENC_us00_n140 ), .ZN(_AES_ENC_us00_n599 ) );
INV_X4 _AES_ENC_us00_U557  ( .A(_AES_ENC_us00_n315 ), .ZN(_AES_ENC_us00_n598 ) );
INV_X4 _AES_ENC_us00_U556  ( .A(_AES_ENC_us00_n270 ), .ZN(_AES_ENC_us00_n597 ) );
INV_X4 _AES_ENC_us00_U555  ( .A(_AES_ENC_us00_n218 ), .ZN(_AES_ENC_us00_n595 ) );
INV_X4 _AES_ENC_us00_U554  ( .A(_AES_ENC_us00_n163 ), .ZN(_AES_ENC_us00_n594 ) );
INV_X4 _AES_ENC_us00_U553  ( .A(_AES_ENC_us00_n90 ), .ZN(_AES_ENC_us00_n593 ) );
INV_X4 _AES_ENC_us00_U552  ( .A(_AES_ENC_us00_n186 ), .ZN(_AES_ENC_us00_n592 ) );
INV_X4 _AES_ENC_us00_U551  ( .A(_AES_ENC_us00_n205 ), .ZN(_AES_ENC_us00_n591 ) );
INV_X4 _AES_ENC_us00_U550  ( .A(_AES_ENC_us00_n136 ), .ZN(_AES_ENC_us00_n590 ) );
INV_X4 _AES_ENC_us00_U549  ( .A(_AES_ENC_us00_n120 ), .ZN(_AES_ENC_us00_n589 ) );
INV_X4 _AES_ENC_us00_U548  ( .A(_AES_ENC_us00_n141 ), .ZN(_AES_ENC_us00_n588 ) );
INV_X4 _AES_ENC_us00_U547  ( .A(_AES_ENC_us00_n370 ), .ZN(_AES_ENC_us00_n587 ) );
INV_X4 _AES_ENC_us00_U546  ( .A(_AES_ENC_us00_n203 ), .ZN(_AES_ENC_us00_n586 ) );
INV_X4 _AES_ENC_us00_U545  ( .A(_AES_ENC_us00_n375 ), .ZN(_AES_ENC_us00_n585 ) );
INV_X4 _AES_ENC_us00_U544  ( .A(_AES_ENC_us00_n286 ), .ZN(_AES_ENC_us00_n584 ) );
INV_X4 _AES_ENC_us00_U543  ( .A(_AES_ENC_us00_n290 ), .ZN(_AES_ENC_us00_n583 ) );
INV_X4 _AES_ENC_us00_U542  ( .A(_AES_ENC_us00_n316 ), .ZN(_AES_ENC_us00_n581 ) );
INV_X4 _AES_ENC_us00_U541  ( .A(_AES_ENC_us00_n182 ), .ZN(_AES_ENC_us00_n580 ) );
INV_X4 _AES_ENC_us00_U540  ( .A(_AES_ENC_us00_n102 ), .ZN(_AES_ENC_us00_n579 ) );
INV_X4 _AES_ENC_us00_U539  ( .A(_AES_ENC_us00_n372 ), .ZN(_AES_ENC_us00_n578 ) );
INV_X4 _AES_ENC_us00_U538  ( .A(_AES_ENC_us00_n103 ), .ZN(_AES_ENC_us00_n577 ) );
INV_X4 _AES_ENC_us00_U537  ( .A(_AES_ENC_us00_n114 ), .ZN(_AES_ENC_us00_n576 ) );
INV_X4 _AES_ENC_us00_U536  ( .A(_AES_ENC_us00_n237 ), .ZN(_AES_ENC_us00_n575 ) );
INV_X4 _AES_ENC_us00_U535  ( .A(_AES_ENC_sa00[0]), .ZN(_AES_ENC_us00_n574 ));
NOR2_X2 _AES_ENC_us00_U534  ( .A1(_AES_ENC_sa00[0]), .A2(_AES_ENC_sa00[6]),.ZN(_AES_ENC_us00_n104 ) );
NOR2_X2 _AES_ENC_us00_U533  ( .A1(_AES_ENC_us00_n574 ), .A2(_AES_ENC_sa00[6]), .ZN(_AES_ENC_us00_n124 ) );
NOR2_X2 _AES_ENC_us00_U532  ( .A1(_AES_ENC_sa00[4]), .A2(_AES_ENC_sa00[3]),.ZN(_AES_ENC_us00_n170 ) );
INV_X4 _AES_ENC_us00_U531  ( .A(_AES_ENC_us00_n569 ), .ZN(_AES_ENC_us00_n572 ) );
NOR2_X2 _AES_ENC_us00_U530  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n431 ) );
NOR2_X2 _AES_ENC_us00_U529  ( .A1(_AES_ENC_sa00[4]), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n432 ) );
NOR2_X2 _AES_ENC_us00_U528  ( .A1(_AES_ENC_us00_n431 ), .A2(_AES_ENC_us00_n432 ), .ZN(_AES_ENC_us00_n430 ) );
NOR2_X2 _AES_ENC_us00_U527  ( .A1(_AES_ENC_us00_n430 ), .A2(_AES_ENC_us00_n575 ), .ZN(_AES_ENC_us00_n429 ) );
NOR3_X2 _AES_ENC_us00_U526  ( .A1(_AES_ENC_us00_n627 ), .A2(_AES_ENC_sa00[5]), .A3(_AES_ENC_us00_n492 ), .ZN(_AES_ENC_us00_n490 ));
NOR2_X2 _AES_ENC_us00_U525  ( .A1(_AES_ENC_us00_n76 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n489 ) );
NOR2_X2 _AES_ENC_us00_U524  ( .A1(_AES_ENC_sa00[4]), .A2(_AES_ENC_us00_n579 ), .ZN(_AES_ENC_us00_n491 ) );
NOR3_X2 _AES_ENC_us00_U523  ( .A1(_AES_ENC_us00_n489 ), .A2(_AES_ENC_us00_n490 ), .A3(_AES_ENC_us00_n491 ), .ZN(_AES_ENC_us00_n483 ) );
INV_X4 _AES_ENC_us00_U522  ( .A(_AES_ENC_sa00[3]), .ZN(_AES_ENC_us00_n621 ));
NAND3_X2 _AES_ENC_us00_U521  ( .A1(_AES_ENC_us00_n544 ), .A2(_AES_ENC_us00_n626 ), .A3(_AES_ENC_sa00[7]), .ZN(_AES_ENC_us00_n543 ));
NOR2_X2 _AES_ENC_us00_U520  ( .A1(_AES_ENC_us00_n611 ), .A2(_AES_ENC_sa00[5]), .ZN(_AES_ENC_us00_n271 ) );
NOR2_X2 _AES_ENC_us00_U519  ( .A1(_AES_ENC_sa00[5]), .A2(_AES_ENC_sa00[2]),.ZN(_AES_ENC_us00_n221 ) );
INV_X4 _AES_ENC_us00_U518  ( .A(_AES_ENC_sa00[5]), .ZN(_AES_ENC_us00_n626 ));
NOR2_X2 _AES_ENC_us00_U517  ( .A1(_AES_ENC_us00_n611 ), .A2(_AES_ENC_sa00[7]), .ZN(_AES_ENC_us00_n417 ) );
NAND3_X2 _AES_ENC_us00_U516  ( .A1(_AES_ENC_us00_n517 ), .A2(_AES_ENC_us00_n518 ), .A3(_AES_ENC_us00_n519 ), .ZN(_AES_ENC_sa00_sub[0] ) );
NOR2_X2 _AES_ENC_us00_U515  ( .A1(_AES_ENC_us00_n626 ), .A2(_AES_ENC_sa00[2]), .ZN(_AES_ENC_us00_n146 ) );
NOR4_X2 _AES_ENC_us00_U512  ( .A1(_AES_ENC_us00_n563 ), .A2(_AES_ENC_us00_n564 ), .A3(_AES_ENC_us00_n565 ), .A4(_AES_ENC_us00_n566 ), .ZN(_AES_ENC_us00_n562 ) );
NOR2_X2 _AES_ENC_us00_U510  ( .A1(_AES_ENC_us00_n567 ), .A2(_AES_ENC_us00_n568 ), .ZN(_AES_ENC_us00_n561 ) );
NAND3_X2 _AES_ENC_us00_U509  ( .A1(_AES_ENC_sa00[2]), .A2(_AES_ENC_sa00[7]), .A3(_AES_ENC_us00_n135 ), .ZN(_AES_ENC_us00_n560 ) );
NOR2_X2 _AES_ENC_us00_U508  ( .A1(_AES_ENC_sa00[7]), .A2(_AES_ENC_sa00[2]),.ZN(_AES_ENC_us00_n402 ) );
NOR2_X2 _AES_ENC_us00_U507  ( .A1(_AES_ENC_sa00[4]), .A2(_AES_ENC_sa00[1]),.ZN(_AES_ENC_us00_n91 ) );
NOR2_X2 _AES_ENC_us00_U506  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_sa00[3]), .ZN(_AES_ENC_us00_n141 ) );
NOR2_X2 _AES_ENC_us00_U505  ( .A1(_AES_ENC_us00_n607 ), .A2(_AES_ENC_sa00[5]), .ZN(_AES_ENC_us00_n171 ) );
NOR2_X2 _AES_ENC_us00_U504  ( .A1(_AES_ENC_us00_n625 ), .A2(_AES_ENC_sa00[2]), .ZN(_AES_ENC_us00_n101 ) );
NOR2_X2 _AES_ENC_us00_U503  ( .A1(_AES_ENC_us00_n614 ), .A2(_AES_ENC_sa00[5]), .ZN(_AES_ENC_us00_n100 ) );
NOR2_X2 _AES_ENC_us00_U502  ( .A1(_AES_ENC_us00_n624 ), .A2(_AES_ENC_sa00[3]), .ZN(_AES_ENC_us00_n265 ) );
INV_X4 _AES_ENC_us00_U501  ( .A(_AES_ENC_us00_n570 ), .ZN(_AES_ENC_us00_n573 ) );
NOR2_X2 _AES_ENC_us00_U500  ( .A1(_AES_ENC_us00_n141 ), .A2(_AES_ENC_us00_n99 ), .ZN(_AES_ENC_us00_n557 ) );
NOR3_X2 _AES_ENC_us00_U499  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n573 ), .A3(_AES_ENC_us00_n120 ), .ZN(_AES_ENC_us00_n555 ) );
NOR2_X2 _AES_ENC_us00_U498  ( .A1(_AES_ENC_us00_n557 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n556 ) );
NOR2_X2 _AES_ENC_us00_U497  ( .A1(_AES_ENC_us00_n555 ), .A2(_AES_ENC_us00_n556 ), .ZN(_AES_ENC_us00_n550 ) );
NOR3_X2 _AES_ENC_us00_U496  ( .A1(_AES_ENC_us00_n200 ), .A2(_AES_ENC_us00_n586 ), .A3(_AES_ENC_us00_n201 ), .ZN(_AES_ENC_us00_n193 ) );
NOR2_X2 _AES_ENC_us00_U495  ( .A1(_AES_ENC_us00_n287 ), .A2(_AES_ENC_us00_n288 ), .ZN(_AES_ENC_us00_n276 ) );
NOR2_X2 _AES_ENC_us00_U494  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n373 ) );
NOR2_X2 _AES_ENC_us00_U492  ( .A1(_AES_ENC_us00_n624 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n374 ) );
NOR2_X2 _AES_ENC_us00_U491  ( .A1(_AES_ENC_us00_n373 ), .A2(_AES_ENC_us00_n374 ), .ZN(_AES_ENC_us00_n371 ) );
NOR2_X2 _AES_ENC_us00_U490  ( .A1(_AES_ENC_sa00[1]), .A2(_AES_ENC_us00_n623 ), .ZN(_AES_ENC_us00_n283 ) );
NOR2_X2 _AES_ENC_us00_U489  ( .A1(_AES_ENC_us00_n283 ), .A2(_AES_ENC_us00_n103 ), .ZN(_AES_ENC_us00_n282 ) );
NOR2_X2 _AES_ENC_us00_U488  ( .A1(_AES_ENC_us00_n370 ), .A2(_AES_ENC_us00_n572 ), .ZN(_AES_ENC_us00_n369 ) );
NOR3_X2 _AES_ENC_us00_U487  ( .A1(_AES_ENC_us00_n427 ), .A2(_AES_ENC_us00_n428 ), .A3(_AES_ENC_us00_n429 ), .ZN(_AES_ENC_us00_n421 ) );
NOR2_X2 _AES_ENC_us00_U486  ( .A1(_AES_ENC_us00_n138 ), .A2(_AES_ENC_us00_n141 ), .ZN(_AES_ENC_us00_n447 ) );
NOR2_X2 _AES_ENC_us00_U483  ( .A1(_AES_ENC_us00_n447 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n444 ) );
INV_X4 _AES_ENC_us00_U482  ( .A(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n596 ));
NOR2_X2 _AES_ENC_us00_U480  ( .A1(_AES_ENC_us00_n140 ), .A2(_AES_ENC_us00_n141 ), .ZN(_AES_ENC_us00_n139 ) );
OR2_X4 _AES_ENC_us00_U479  ( .A1(_AES_ENC_us00_n100 ), .A2(_AES_ENC_us00_n101 ), .ZN(_AES_ENC_us00_n571 ) );
AND2_X2 _AES_ENC_us00_U478  ( .A1(_AES_ENC_us00_n571 ), .A2(_AES_ENC_us00_n99 ), .ZN(_AES_ENC_us00_n92 ) );
NOR2_X2 _AES_ENC_us00_U477  ( .A1(_AES_ENC_us00_n120 ), .A2(_AES_ENC_us00_n265 ), .ZN(_AES_ENC_us00_n400 ) );
NOR2_X2 _AES_ENC_us00_U474  ( .A1(_AES_ENC_us00_n400 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n399 ) );
NOR2_X2 _AES_ENC_us00_U473  ( .A1(_AES_ENC_us00_n264 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n263 ) );
NOR2_X2 _AES_ENC_us00_U472  ( .A1(_AES_ENC_us00_n267 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n261 ) );
NOR2_X2 _AES_ENC_us00_U471  ( .A1(_AES_ENC_us00_n265 ), .A2(_AES_ENC_us00_n266 ), .ZN(_AES_ENC_us00_n262 ) );
NOR3_X2 _AES_ENC_us00_U470  ( .A1(_AES_ENC_us00_n261 ), .A2(_AES_ENC_us00_n262 ), .A3(_AES_ENC_us00_n263 ), .ZN(_AES_ENC_us00_n260 ) );
NOR2_X2 _AES_ENC_us00_U469  ( .A1(_AES_ENC_us00_n624 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n119 ) );
NOR2_X2 _AES_ENC_us00_U468  ( .A1(_AES_ENC_us00_n572 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n247 ) );
NOR2_X2 _AES_ENC_us00_U467  ( .A1(_AES_ENC_us00_n145 ), .A2(_AES_ENC_us00_n618 ), .ZN(_AES_ENC_us00_n143 ) );
NOR2_X2 _AES_ENC_us00_U466  ( .A1(_AES_ENC_us00_n143 ), .A2(_AES_ENC_us00_n144 ), .ZN(_AES_ENC_us00_n142 ) );
NOR2_X2 _AES_ENC_us00_U465  ( .A1(_AES_ENC_us00_n142 ), .A2(_AES_ENC_us00_n592 ), .ZN(_AES_ENC_us00_n130 ) );
NOR2_X2 _AES_ENC_us00_U464  ( .A1(_AES_ENC_sa00[1]), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n565 ) );
NOR2_X2 _AES_ENC_us00_U463  ( .A1(_AES_ENC_us00_n170 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n215 ) );
NOR2_X2 _AES_ENC_us00_U462  ( .A1(_AES_ENC_us00_n121 ), .A2(_AES_ENC_us00_n100 ), .ZN(_AES_ENC_us00_n401 ) );
NOR2_X2 _AES_ENC_us00_U461  ( .A1(_AES_ENC_us00_n401 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n397 ) );
NOR2_X2 _AES_ENC_us00_U460  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n214 ) );
NOR2_X2 _AES_ENC_us00_U459  ( .A1(_AES_ENC_us00_n91 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n553 ) );
NOR2_X2 _AES_ENC_us00_U458  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n621 ), .ZN(_AES_ENC_us00_n554 ) );
NOR2_X2 _AES_ENC_us00_U455  ( .A1(_AES_ENC_us00_n285 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n552 ) );
NOR4_X2 _AES_ENC_us00_U448  ( .A1(_AES_ENC_us00_n552 ), .A2(_AES_ENC_us00_n553 ), .A3(_AES_ENC_us00_n392 ), .A4(_AES_ENC_us00_n554 ), .ZN(_AES_ENC_us00_n551 ) );
NOR2_X2 _AES_ENC_us00_U447  ( .A1(_AES_ENC_us00_n91 ), .A2(_AES_ENC_us00_n286 ), .ZN(_AES_ENC_us00_n264 ) );
NOR2_X2 _AES_ENC_us00_U442  ( .A1(_AES_ENC_us00_n91 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n441 ) );
NOR2_X2 _AES_ENC_us00_U441  ( .A1(_AES_ENC_us00_n265 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n453 ) );
NOR2_X2 _AES_ENC_us00_U438  ( .A1(_AES_ENC_us00_n122 ), .A2(_AES_ENC_us00_n100 ), .ZN(_AES_ENC_us00_n266 ) );
NOR2_X2 _AES_ENC_us00_U435  ( .A1(_AES_ENC_us00_n120 ), .A2(_AES_ENC_us00_n170 ), .ZN(_AES_ENC_us00_n305 ) );
NOR2_X2 _AES_ENC_us00_U434  ( .A1(_AES_ENC_us00_n305 ), .A2(_AES_ENC_us00_n609 ), .ZN(_AES_ENC_us00_n302 ) );
NOR3_X2 _AES_ENC_us00_U433  ( .A1(_AES_ENC_us00_n623 ), .A2(_AES_ENC_sa00[1]), .A3(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n513 ));
INV_X4 _AES_ENC_us00_U428  ( .A(_AES_ENC_us00_n265 ), .ZN(_AES_ENC_us00_n623 ) );
NOR2_X2 _AES_ENC_us00_U427  ( .A1(_AES_ENC_us00_n199 ), .A2(_AES_ENC_us00_n265 ), .ZN(_AES_ENC_us00_n492 ) );
NOR2_X2 _AES_ENC_us00_U421  ( .A1(_AES_ENC_us00_n265 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n511 ) );
NOR2_X2 _AES_ENC_us00_U420  ( .A1(_AES_ENC_us00_n165 ), .A2(_AES_ENC_us00_n170 ), .ZN(_AES_ENC_us00_n115 ) );
NOR3_X2 _AES_ENC_us00_U419  ( .A1(_AES_ENC_us00_n589 ), .A2(_AES_ENC_us00_n170 ), .A3(_AES_ENC_us00_n616 ), .ZN(_AES_ENC_us00_n251 ) );
NOR2_X2 _AES_ENC_us00_U418  ( .A1(_AES_ENC_us00_n626 ), .A2(_AES_ENC_us00_n611 ), .ZN(_AES_ENC_us00_n396 ) );
NOR3_X2 _AES_ENC_us00_U417  ( .A1(_AES_ENC_us00_n590 ), .A2(_AES_ENC_us00_n627 ), .A3(_AES_ENC_us00_n611 ), .ZN(_AES_ENC_us00_n398 ) );
NOR3_X2 _AES_ENC_us00_U416  ( .A1(_AES_ENC_us00_n610 ), .A2(_AES_ENC_us00_n572 ), .A3(_AES_ENC_us00_n575 ), .ZN(_AES_ENC_us00_n233 ) );
NOR3_X2 _AES_ENC_us00_U415  ( .A1(_AES_ENC_us00_n237 ), .A2(_AES_ENC_us00_n572 ), .A3(_AES_ENC_us00_n609 ), .ZN(_AES_ENC_us00_n428 ) );
NOR3_X2 _AES_ENC_us00_U414  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n572 ), .A3(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n502 ) );
NOR3_X2 _AES_ENC_us00_U413  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n572 ), .A3(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n301 ) );
NOR3_X2 _AES_ENC_us00_U410  ( .A1(_AES_ENC_us00_n187 ), .A2(_AES_ENC_us00_n188 ), .A3(_AES_ENC_us00_n189 ), .ZN(_AES_ENC_us00_n177 ) );
NOR4_X2 _AES_ENC_us00_U409  ( .A1(_AES_ENC_us00_n390 ), .A2(_AES_ENC_us00_n391 ), .A3(_AES_ENC_us00_n392 ), .A4(_AES_ENC_us00_n393 ), .ZN(_AES_ENC_us00_n389 ) );
NOR3_X2 _AES_ENC_us00_U406  ( .A1(_AES_ENC_us00_n397 ), .A2(_AES_ENC_us00_n398 ), .A3(_AES_ENC_us00_n399 ), .ZN(_AES_ENC_us00_n388 ) );
NOR2_X2 _AES_ENC_us00_U405  ( .A1(_AES_ENC_us00_n527 ), .A2(_AES_ENC_us00_n528 ), .ZN(_AES_ENC_us00_n523 ) );
NOR4_X2 _AES_ENC_us00_U404  ( .A1(_AES_ENC_us00_n250 ), .A2(_AES_ENC_us00_n148 ), .A3(_AES_ENC_us00_n525 ), .A4(_AES_ENC_us00_n526 ), .ZN(_AES_ENC_us00_n524 ) );
NOR3_X2 _AES_ENC_us00_U403  ( .A1(_AES_ENC_us00_n92 ), .A2(_AES_ENC_us00_n93 ), .A3(_AES_ENC_us00_n94 ), .ZN(_AES_ENC_us00_n84 ));
NOR4_X2 _AES_ENC_us00_U401  ( .A1(_AES_ENC_us00_n485 ), .A2(_AES_ENC_us00_n486 ), .A3(_AES_ENC_us00_n487 ), .A4(_AES_ENC_us00_n488 ), .ZN(_AES_ENC_us00_n484 ) );
NOR4_X2 _AES_ENC_us00_U400  ( .A1(_AES_ENC_us00_n353 ), .A2(_AES_ENC_us00_n354 ), .A3(_AES_ENC_us00_n355 ), .A4(_AES_ENC_us00_n356 ), .ZN(_AES_ENC_us00_n352 ) );
NOR4_X2 _AES_ENC_us00_U399  ( .A1(_AES_ENC_us00_n232 ), .A2(_AES_ENC_us00_n233 ), .A3(_AES_ENC_us00_n234 ), .A4(_AES_ENC_us00_n235 ), .ZN(_AES_ENC_us00_n231 ) );
NOR3_X2 _AES_ENC_us00_U398  ( .A1(_AES_ENC_us00_n453 ), .A2(_AES_ENC_us00_n454 ), .A3(_AES_ENC_us00_n455 ), .ZN(_AES_ENC_us00_n452 ) );
NOR2_X2 _AES_ENC_us00_U397  ( .A1(_AES_ENC_us00_n499 ), .A2(_AES_ENC_us00_n538 ), .ZN(_AES_ENC_us00_n537 ) );
NOR2_X2 _AES_ENC_us00_U396  ( .A1(_AES_ENC_us00_n598 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n311 ) );
NOR2_X2 _AES_ENC_us00_U393  ( .A1(_AES_ENC_us00_n623 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n314 ) );
NOR2_X2 _AES_ENC_us00_U390  ( .A1(_AES_ENC_us00_n141 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n312 ) );
NOR4_X2 _AES_ENC_us00_U389  ( .A1(_AES_ENC_us00_n311 ), .A2(_AES_ENC_us00_n312 ), .A3(_AES_ENC_us00_n313 ), .A4(_AES_ENC_us00_n314 ), .ZN(_AES_ENC_us00_n310 ) );
NOR2_X2 _AES_ENC_us00_U388  ( .A1(_AES_ENC_us00_n116 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n161 ) );
NOR2_X2 _AES_ENC_us00_U387  ( .A1(_AES_ENC_us00_n163 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n162 ) );
NOR3_X2 _AES_ENC_us00_U386  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n170 ), .A3(_AES_ENC_us00_n120 ), .ZN(_AES_ENC_us00_n159 ) );
NOR4_X2 _AES_ENC_us00_U385  ( .A1(_AES_ENC_us00_n159 ), .A2(_AES_ENC_us00_n160 ), .A3(_AES_ENC_us00_n161 ), .A4(_AES_ENC_us00_n162 ), .ZN(_AES_ENC_us00_n158 ) );
NOR2_X2 _AES_ENC_us00_U384  ( .A1(_AES_ENC_us00_n371 ), .A2(_AES_ENC_us00_n578 ), .ZN(_AES_ENC_us00_n366 ) );
NOR2_X2 _AES_ENC_us00_U383  ( .A1(_AES_ENC_us00_n369 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n367 ) );
NOR2_X2 _AES_ENC_us00_U382  ( .A1(_AES_ENC_us00_n572 ), .A2(_AES_ENC_us00_n579 ), .ZN(_AES_ENC_us00_n368 ) );
NOR4_X2 _AES_ENC_us00_U374  ( .A1(_AES_ENC_us00_n365 ), .A2(_AES_ENC_us00_n366 ), .A3(_AES_ENC_us00_n367 ), .A4(_AES_ENC_us00_n368 ), .ZN(_AES_ENC_us00_n364 ) );
NOR2_X2 _AES_ENC_us00_U373  ( .A1(_AES_ENC_us00_n606 ), .A2(_AES_ENC_us00_n582 ), .ZN(_AES_ENC_us00_n89 ) );
NOR2_X2 _AES_ENC_us00_U372  ( .A1(_AES_ENC_us00_n91 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n87 ) );
NOR2_X2 _AES_ENC_us00_U370  ( .A1(_AES_ENC_us00_n90 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n88 ) );
NOR4_X2 _AES_ENC_us00_U369  ( .A1(_AES_ENC_us00_n86 ), .A2(_AES_ENC_us00_n87 ), .A3(_AES_ENC_us00_n88 ), .A4(_AES_ENC_us00_n89 ),.ZN(_AES_ENC_us00_n85 ) );
NOR3_X2 _AES_ENC_us00_U368  ( .A1(_AES_ENC_us00_n237 ), .A2(_AES_ENC_us00_n621 ), .A3(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n232 ) );
NOR2_X2 _AES_ENC_us00_U367  ( .A1(_AES_ENC_us00_n626 ), .A2(_AES_ENC_us00_n627 ), .ZN(_AES_ENC_us00_n79 ) );
INV_X4 _AES_ENC_us00_U366  ( .A(_AES_ENC_us00_n171 ), .ZN(_AES_ENC_us00_n606 ) );
NOR3_X2 _AES_ENC_us00_U365  ( .A1(_AES_ENC_us00_n286 ), .A2(_AES_ENC_us00_n135 ), .A3(_AES_ENC_us00_n611 ), .ZN(_AES_ENC_us00_n78 ) );
INV_X4 _AES_ENC_us00_U364  ( .A(_AES_ENC_us00_n100 ), .ZN(_AES_ENC_us00_n613 ) );
NOR2_X2 _AES_ENC_us00_U363  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n265 ), .ZN(_AES_ENC_us00_n93 ) );
INV_X4 _AES_ENC_us00_U354  ( .A(_AES_ENC_us00_n101 ), .ZN(_AES_ENC_us00_n617 ) );
NOR2_X2 _AES_ENC_us00_U353  ( .A1(_AES_ENC_us00_n569 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n267 ) );
NOR2_X2 _AES_ENC_us00_U352  ( .A1(_AES_ENC_us00_n620 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n270 ) );
NOR2_X2 _AES_ENC_us00_U351  ( .A1(_AES_ENC_us00_n572 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n99 ) );
NOR2_X2 _AES_ENC_us00_U350  ( .A1(_AES_ENC_us00_n609 ), .A2(_AES_ENC_us00_n627 ), .ZN(_AES_ENC_us00_n185 ) );
NOR2_X2 _AES_ENC_us00_U349  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n90 ) );
NOR2_X2 _AES_ENC_us00_U348  ( .A1(_AES_ENC_us00_n622 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n135 ) );
NOR2_X2 _AES_ENC_us00_U347  ( .A1(_AES_ENC_sa00[1]), .A2(_AES_ENC_us00_n73 ), .ZN(_AES_ENC_us00_n173 ) );
NOR2_X2 _AES_ENC_us00_U346  ( .A1(_AES_ENC_us00_n619 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n285 ) );
NOR2_X2 _AES_ENC_us00_U345  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_us00_n170 ), .ZN(_AES_ENC_us00_n370 ) );
NOR2_X2 _AES_ENC_us00_U338  ( .A1(_AES_ENC_us00_n626 ), .A2(_AES_ENC_us00_n607 ), .ZN(_AES_ENC_us00_n122 ) );
NOR2_X2 _AES_ENC_us00_U335  ( .A1(_AES_ENC_us00_n627 ), .A2(_AES_ENC_us00_n616 ), .ZN(_AES_ENC_us00_n240 ) );
NOR2_X2 _AES_ENC_us00_U329  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_us00_n624 ), .ZN(_AES_ENC_us00_n72 ) );
NOR2_X2 _AES_ENC_us00_U328  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_us00_n624 ), .ZN(_AES_ENC_us00_n136 ) );
NOR2_X2 _AES_ENC_us00_U327  ( .A1(_AES_ENC_us00_n625 ), .A2(_AES_ENC_us00_n611 ), .ZN(_AES_ENC_us00_n121 ) );
NOR2_X2 _AES_ENC_us00_U325  ( .A1(_AES_ENC_sa00[1]), .A2(_AES_ENC_us00_n170 ), .ZN(_AES_ENC_us00_n140 ) );
NOR2_X2 _AES_ENC_us00_U324  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_us00_n265 ), .ZN(_AES_ENC_us00_n165 ) );
NOR2_X2 _AES_ENC_us00_U319  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n138 ) );
NOR2_X2 _AES_ENC_us00_U318  ( .A1(_AES_ENC_us00_n614 ), .A2(_AES_ENC_us00_n626 ), .ZN(_AES_ENC_us00_n144 ) );
NOR2_X2 _AES_ENC_us00_U317  ( .A1(_AES_ENC_us00_n72 ), .A2(_AES_ENC_us00_n170 ), .ZN(_AES_ENC_us00_n73 ) );
NOR2_X2 _AES_ENC_us00_U316  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_us00_n572 ), .ZN(_AES_ENC_us00_n120 ) );
NOR2_X2 _AES_ENC_us00_U315  ( .A1(_AES_ENC_us00_n136 ), .A2(_AES_ENC_us00_n140 ), .ZN(_AES_ENC_us00_n318 ) );
NOR2_X2 _AES_ENC_us00_U314  ( .A1(_AES_ENC_us00_n318 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n317 ) );
NOR2_X2 _AES_ENC_us00_U312  ( .A1(_AES_ENC_us00_n316 ), .A2(_AES_ENC_us00_n317 ), .ZN(_AES_ENC_us00_n309 ) );
NOR2_X2 _AES_ENC_us00_U311  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n588 ), .ZN(_AES_ENC_us00_n239 ) );
NOR2_X2 _AES_ENC_us00_U310  ( .A1(_AES_ENC_us00_n238 ), .A2(_AES_ENC_us00_n239 ), .ZN(_AES_ENC_us00_n230 ) );
NOR3_X2 _AES_ENC_us00_U309  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n103 ), .A3(_AES_ENC_us00_n173 ), .ZN(_AES_ENC_us00_n476 ) );
NOR3_X2 _AES_ENC_us00_U303  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n140 ), .A3(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n477 ) );
NOR2_X2 _AES_ENC_us00_U302  ( .A1(_AES_ENC_us00_n476 ), .A2(_AES_ENC_us00_n477 ), .ZN(_AES_ENC_us00_n470 ) );
NOR2_X2 _AES_ENC_us00_U300  ( .A1(_AES_ENC_us00_n614 ), .A2(_AES_ENC_us00_n591 ), .ZN(_AES_ENC_us00_n331 ) );
NOR2_X2 _AES_ENC_us00_U299  ( .A1(_AES_ENC_us00_n135 ), .A2(_AES_ENC_us00_n136 ), .ZN(_AES_ENC_us00_n134 ) );
NOR2_X2 _AES_ENC_us00_U298  ( .A1(_AES_ENC_us00_n99 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n528 ) );
NOR2_X2 _AES_ENC_us00_U297  ( .A1(_AES_ENC_us00_n285 ), .A2(_AES_ENC_us00_n286 ), .ZN(_AES_ENC_us00_n284 ) );
NOR2_X2 _AES_ENC_us00_U296  ( .A1(_AES_ENC_us00_n284 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n280 ) );
NOR2_X2 _AES_ENC_us00_U295  ( .A1(_AES_ENC_us00_n370 ), .A2(_AES_ENC_us00_n573 ), .ZN(_AES_ENC_us00_n446 ) );
NOR2_X2 _AES_ENC_us00_U294  ( .A1(_AES_ENC_us00_n446 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n445 ) );
NOR2_X2 _AES_ENC_us00_U293  ( .A1(_AES_ENC_us00_n289 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n288 ) );
NOR2_X2 _AES_ENC_us00_U292  ( .A1(_AES_ENC_us00_n205 ), .A2(_AES_ENC_us00_n270 ), .ZN(_AES_ENC_us00_n416 ) );
NOR2_X2 _AES_ENC_us00_U291  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n584 ), .ZN(_AES_ENC_us00_n358 ) );
NOR2_X2 _AES_ENC_us00_U290  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n602 ), .ZN(_AES_ENC_us00_n359 ) );
NOR2_X2 _AES_ENC_us00_U284  ( .A1(_AES_ENC_us00_n358 ), .A2(_AES_ENC_us00_n359 ), .ZN(_AES_ENC_us00_n351 ) );
NOR2_X2 _AES_ENC_us00_U283  ( .A1(_AES_ENC_us00_n173 ), .A2(_AES_ENC_us00_n136 ), .ZN(_AES_ENC_us00_n456 ) );
NOR2_X2 _AES_ENC_us00_U282  ( .A1(_AES_ENC_us00_n456 ), .A2(_AES_ENC_us00_n616 ), .ZN(_AES_ENC_us00_n454 ) );
NOR2_X2 _AES_ENC_us00_U281  ( .A1(_AES_ENC_us00_n95 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n94 ) );
NOR2_X2 _AES_ENC_us00_U280  ( .A1(_AES_ENC_us00_n73 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n202 ) );
NOR2_X2 _AES_ENC_us00_U279  ( .A1(_AES_ENC_us00_n202 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n201 ) );
NOR2_X2 _AES_ENC_us00_U273  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n620 ), .ZN(_AES_ENC_us00_n168 ) );
NOR2_X2 _AES_ENC_us00_U272  ( .A1(_AES_ENC_us00_n573 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n167 ) );
NOR2_X2 _AES_ENC_us00_U271  ( .A1(_AES_ENC_us00_n167 ), .A2(_AES_ENC_us00_n168 ), .ZN(_AES_ENC_us00_n166 ) );
NOR2_X2 _AES_ENC_us00_U270  ( .A1(_AES_ENC_us00_n165 ), .A2(_AES_ENC_us00_n166 ), .ZN(_AES_ENC_us00_n160 ) );
NOR4_X2 _AES_ENC_us00_U269  ( .A1(_AES_ENC_us00_n439 ), .A2(_AES_ENC_us00_n440 ), .A3(_AES_ENC_us00_n441 ), .A4(_AES_ENC_us00_n442 ), .ZN(_AES_ENC_us00_n438 ) );
NOR2_X2 _AES_ENC_us00_U268  ( .A1(_AES_ENC_us00_n444 ), .A2(_AES_ENC_us00_n445 ), .ZN(_AES_ENC_us00_n437 ) );
NOR2_X2 _AES_ENC_us00_U267  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n123 ), .ZN(_AES_ENC_us00_n527 ) );
NOR2_X2 _AES_ENC_us00_U263  ( .A1(_AES_ENC_us00_n138 ), .A2(_AES_ENC_us00_n205 ), .ZN(_AES_ENC_us00_n204 ) );
NOR2_X2 _AES_ENC_us00_U262  ( .A1(_AES_ENC_us00_n204 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n200 ) );
NOR2_X2 _AES_ENC_us00_U258  ( .A1(_AES_ENC_us00_n607 ), .A2(_AES_ENC_us00_n590 ), .ZN(_AES_ENC_us00_n187 ) );
NOR2_X2 _AES_ENC_us00_U255  ( .A1(_AES_ENC_us00_n357 ), .A2(_AES_ENC_us00_n582 ), .ZN(_AES_ENC_us00_n503 ) );
NOR2_X2 _AES_ENC_us00_U254  ( .A1(_AES_ENC_us00_n606 ), .A2(_AES_ENC_us00_n290 ), .ZN(_AES_ENC_us00_n455 ) );
NOR2_X2 _AES_ENC_us00_U253  ( .A1(_AES_ENC_us00_n140 ), .A2(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n433 ) );
NOR2_X2 _AES_ENC_us00_U252  ( .A1(_AES_ENC_us00_n433 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n427 ) );
NOR2_X2 _AES_ENC_us00_U251  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n577 ), .ZN(_AES_ENC_us00_n188 ) );
NOR2_X2 _AES_ENC_us00_U250  ( .A1(_AES_ENC_us00_n609 ), .A2(_AES_ENC_us00_n580 ), .ZN(_AES_ENC_us00_n70 ) );
NOR2_X2 _AES_ENC_us00_U243  ( .A1(_AES_ENC_us00_n609 ), .A2(_AES_ENC_us00_n590 ), .ZN(_AES_ENC_us00_n486 ) );
INV_X4 _AES_ENC_us00_U242  ( .A(_AES_ENC_us00_n165 ), .ZN(_AES_ENC_us00_n582 ) );
NOR2_X2 _AES_ENC_us00_U241  ( .A1(_AES_ENC_us00_n616 ), .A2(_AES_ENC_us00_n597 ), .ZN(_AES_ENC_us00_n313 ) );
NOR2_X2 _AES_ENC_us00_U240  ( .A1(_AES_ENC_us00_n593 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n68 ) );
NOR2_X2 _AES_ENC_us00_U239  ( .A1(_AES_ENC_us00_n205 ), .A2(_AES_ENC_us00_n267 ), .ZN(_AES_ENC_us00_n304 ) );
NOR2_X2 _AES_ENC_us00_U238  ( .A1(_AES_ENC_us00_n304 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n303 ) );
NOR2_X2 _AES_ENC_us00_U237  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n602 ), .ZN(_AES_ENC_us00_n246 ) );
NOR2_X2 _AES_ENC_us00_U236  ( .A1(_AES_ENC_us00_n115 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n112 ) );
NOR2_X2 _AES_ENC_us00_U235  ( .A1(_AES_ENC_us00_n286 ), .A2(_AES_ENC_us00_n138 ), .ZN(_AES_ENC_us00_n255 ) );
NOR2_X2 _AES_ENC_us00_U234  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n117 ), .ZN(_AES_ENC_us00_n355 ) );
NOR2_X2 _AES_ENC_us00_U229  ( .A1(_AES_ENC_us00_n623 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n566 ) );
NOR2_X2 _AES_ENC_us00_U228  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n602 ), .ZN(_AES_ENC_us00_n390 ) );
NOR2_X2 _AES_ENC_us00_U227  ( .A1(_AES_ENC_us00_n623 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n248 ) );
NOR2_X2 _AES_ENC_us00_U226  ( .A1(_AES_ENC_us00_n606 ), .A2(_AES_ENC_us00_n589 ), .ZN(_AES_ENC_us00_n198 ) );
NOR2_X2 _AES_ENC_us00_U225  ( .A1(_AES_ENC_us00_n72 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n71 ) );
NOR2_X2 _AES_ENC_us00_U223  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n172 ), .ZN(_AES_ENC_us00_n440 ) );
NOR2_X2 _AES_ENC_us00_U222  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n602 ), .ZN(_AES_ENC_us00_n326 ) );
NOR2_X2 _AES_ENC_us00_U221  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n569 ), .ZN(_AES_ENC_us00_n249 ) );
NOR2_X2 _AES_ENC_us00_U217  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n117 ), .ZN(_AES_ENC_us00_n110 ) );
NOR2_X2 _AES_ENC_us00_U213  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n341 ), .ZN(_AES_ENC_us00_n487 ) );
NOR2_X2 _AES_ENC_us00_U212  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n589 ), .ZN(_AES_ENC_us00_n328 ) );
NOR2_X2 _AES_ENC_us00_U211  ( .A1(_AES_ENC_us00_n73 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n69 ) );
NOR2_X2 _AES_ENC_us00_U210  ( .A1(_AES_ENC_us00_n73 ), .A2(_AES_ENC_us00_n357 ), .ZN(_AES_ENC_us00_n354 ) );
NOR2_X2 _AES_ENC_us00_U209  ( .A1(_AES_ENC_us00_n73 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n500 ) );
NOR2_X2 _AES_ENC_us00_U208  ( .A1(_AES_ENC_us00_n120 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n118 ) );
NOR2_X2 _AES_ENC_us00_U207  ( .A1(_AES_ENC_us00_n120 ), .A2(_AES_ENC_us00_n620 ), .ZN(_AES_ENC_us00_n415 ) );
NOR3_X2 _AES_ENC_us00_U201  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n138 ), .A3(_AES_ENC_us00_n205 ), .ZN(_AES_ENC_us00_n216 ) );
NOR3_X2 _AES_ENC_us00_U200  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n136 ), .A3(_AES_ENC_us00_n135 ), .ZN(_AES_ENC_us00_n342 ) );
NOR2_X2 _AES_ENC_us00_U199  ( .A1(_AES_ENC_us00_n199 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n327 ) );
NOR2_X2 _AES_ENC_us00_U198  ( .A1(_AES_ENC_us00_n138 ), .A2(_AES_ENC_us00_n120 ), .ZN(_AES_ENC_us00_n137 ) );
NOR3_X2 _AES_ENC_us00_U197  ( .A1(_AES_ENC_us00_n607 ), .A2(_AES_ENC_us00_n73 ), .A3(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n217 ) );
NOR2_X2 _AES_ENC_us00_U196  ( .A1(_AES_ENC_us00_n199 ), .A2(_AES_ENC_us00_n285 ), .ZN(_AES_ENC_us00_n77 ) );
NOR2_X2 _AES_ENC_us00_U195  ( .A1(_AES_ENC_us00_n120 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n442 ) );
NOR2_X2 _AES_ENC_us00_U194  ( .A1(_AES_ENC_us00_n270 ), .A2(_AES_ENC_us00_n90 ), .ZN(_AES_ENC_us00_n218 ) );
NOR2_X2 _AES_ENC_us00_U187  ( .A1(_AES_ENC_us00_n357 ), .A2(_AES_ENC_us00_n372 ), .ZN(_AES_ENC_us00_n102 ) );
NOR2_X2 _AES_ENC_us00_U186  ( .A1(_AES_ENC_us00_n573 ), .A2(_AES_ENC_us00_n120 ), .ZN(_AES_ENC_us00_n512 ) );
NOR2_X2 _AES_ENC_us00_U185  ( .A1(_AES_ENC_us00_n370 ), .A2(_AES_ENC_us00_n135 ), .ZN(_AES_ENC_us00_n289 ) );
NOR3_X2 _AES_ENC_us00_U184  ( .A1(_AES_ENC_us00_n625 ), .A2(_AES_ENC_us00_n78 ), .A3(_AES_ENC_us00_n585 ), .ZN(_AES_ENC_us00_n365 ) );
NOR3_X2 _AES_ENC_us00_U183  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n138 ), .A3(_AES_ENC_us00_n205 ), .ZN(_AES_ENC_us00_n300 ) );
NOR3_X2 _AES_ENC_us00_U182  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n573 ), .A3(_AES_ENC_us00_n182 ), .ZN(_AES_ENC_us00_n526 ) );
NOR3_X2 _AES_ENC_us00_U181  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n103 ), .A3(_AES_ENC_us00_n173 ), .ZN(_AES_ENC_us00_n353 ) );
NOR2_X2 _AES_ENC_us00_U180  ( .A1(_AES_ENC_us00_n165 ), .A2(_AES_ENC_us00_n99 ), .ZN(_AES_ENC_us00_n461 ) );
NOR2_X2 _AES_ENC_us00_U174  ( .A1(_AES_ENC_us00_n93 ), .A2(_AES_ENC_us00_n342 ), .ZN(_AES_ENC_us00_n336 ) );
NOR4_X2 _AES_ENC_us00_U173  ( .A1(_AES_ENC_us00_n68 ), .A2(_AES_ENC_us00_n69 ), .A3(_AES_ENC_us00_n70 ), .A4(_AES_ENC_us00_n71 ),.ZN(_AES_ENC_us00_n67 ) );
NOR4_X2 _AES_ENC_us00_U172  ( .A1(_AES_ENC_us00_n110 ), .A2(_AES_ENC_us00_n111 ), .A3(_AES_ENC_us00_n112 ), .A4(_AES_ENC_us00_n113 ), .ZN(_AES_ENC_us00_n109 ) );
NOR2_X2 _AES_ENC_us00_U171  ( .A1(_AES_ENC_us00_n118 ), .A2(_AES_ENC_us00_n119 ), .ZN(_AES_ENC_us00_n108 ) );
NAND3_X2 _AES_ENC_us00_U170  ( .A1(_AES_ENC_us00_n569 ), .A2(_AES_ENC_us00_n582 ), .A3(_AES_ENC_us00_n515 ), .ZN(_AES_ENC_us00_n505 ) );
NOR2_X2 _AES_ENC_us00_U169  ( .A1(_AES_ENC_us00_n513 ), .A2(_AES_ENC_us00_n514 ), .ZN(_AES_ENC_us00_n506 ) );
NOR3_X2 _AES_ENC_us00_U168  ( .A1(_AES_ENC_us00_n501 ), .A2(_AES_ENC_us00_n502 ), .A3(_AES_ENC_us00_n503 ), .ZN(_AES_ENC_us00_n496 ) );
NOR4_X2 _AES_ENC_us00_U162  ( .A1(_AES_ENC_us00_n212 ), .A2(_AES_ENC_us00_n498 ), .A3(_AES_ENC_us00_n499 ), .A4(_AES_ENC_us00_n500 ), .ZN(_AES_ENC_us00_n497 ) );
NOR4_X2 _AES_ENC_us00_U161  ( .A1(_AES_ENC_us00_n300 ), .A2(_AES_ENC_us00_n301 ), .A3(_AES_ENC_us00_n302 ), .A4(_AES_ENC_us00_n303 ), .ZN(_AES_ENC_us00_n299 ) );
NOR2_X2 _AES_ENC_us00_U160  ( .A1(_AES_ENC_us00_n330 ), .A2(_AES_ENC_us00_n331 ), .ZN(_AES_ENC_us00_n324 ) );
NOR4_X2 _AES_ENC_us00_U159  ( .A1(_AES_ENC_us00_n326 ), .A2(_AES_ENC_us00_n327 ), .A3(_AES_ENC_us00_n328 ), .A4(_AES_ENC_us00_n329 ), .ZN(_AES_ENC_us00_n325 ) );
NOR2_X2 _AES_ENC_us00_U158  ( .A1(_AES_ENC_us00_n250 ), .A2(_AES_ENC_us00_n251 ), .ZN(_AES_ENC_us00_n244 ) );
NOR4_X2 _AES_ENC_us00_U157  ( .A1(_AES_ENC_us00_n246 ), .A2(_AES_ENC_us00_n247 ), .A3(_AES_ENC_us00_n248 ), .A4(_AES_ENC_us00_n249 ), .ZN(_AES_ENC_us00_n245 ) );
NOR4_X2 _AES_ENC_us00_U156  ( .A1(_AES_ENC_us00_n212 ), .A2(_AES_ENC_us00_n213 ), .A3(_AES_ENC_us00_n214 ), .A4(_AES_ENC_us00_n215 ), .ZN(_AES_ENC_us00_n211 ) );
NOR2_X2 _AES_ENC_us00_U155  ( .A1(_AES_ENC_us00_n216 ), .A2(_AES_ENC_us00_n217 ), .ZN(_AES_ENC_us00_n210 ) );
NOR3_X2 _AES_ENC_us00_U154  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n140 ), .A3(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n234 ) );
NOR3_X2 _AES_ENC_us00_U153  ( .A1(_AES_ENC_us00_n620 ), .A2(_AES_ENC_us00_n120 ), .A3(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n525 ) );
NOR2_X2 _AES_ENC_us00_U152  ( .A1(_AES_ENC_us00_n137 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n132 ) );
NOR2_X2 _AES_ENC_us00_U143  ( .A1(_AES_ENC_us00_n139 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n131 ) );
NOR2_X2 _AES_ENC_us00_U142  ( .A1(_AES_ENC_us00_n134 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n133 ) );
NOR4_X2 _AES_ENC_us00_U141  ( .A1(_AES_ENC_us00_n130 ), .A2(_AES_ENC_us00_n131 ), .A3(_AES_ENC_us00_n132 ), .A4(_AES_ENC_us00_n133 ), .ZN(_AES_ENC_us00_n129 ) );
NOR2_X2 _AES_ENC_us00_U140  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n595 ), .ZN(_AES_ENC_us00_n338 ) );
NOR2_X2 _AES_ENC_us00_U132  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n341 ), .ZN(_AES_ENC_us00_n339 ) );
NOR2_X2 _AES_ENC_us00_U131  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n587 ), .ZN(_AES_ENC_us00_n340 ) );
NOR4_X2 _AES_ENC_us00_U130  ( .A1(_AES_ENC_us00_n338 ), .A2(_AES_ENC_us00_n339 ), .A3(_AES_ENC_us00_n340 ), .A4(_AES_ENC_us00_n238 ), .ZN(_AES_ENC_us00_n337 ) );
NOR3_X2 _AES_ENC_us00_U129  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n73 ), .A3(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n278 ) );
NOR3_X2 _AES_ENC_us00_U128  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n573 ), .A3(_AES_ENC_us00_n182 ), .ZN(_AES_ENC_us00_n279 ) );
NOR2_X2 _AES_ENC_us00_U127  ( .A1(_AES_ENC_us00_n282 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n281 ) );
NOR4_X2 _AES_ENC_us00_U126  ( .A1(_AES_ENC_us00_n278 ), .A2(_AES_ENC_us00_n279 ), .A3(_AES_ENC_us00_n280 ), .A4(_AES_ENC_us00_n281 ), .ZN(_AES_ENC_us00_n277 ) );
NOR2_X2 _AES_ENC_us00_U121  ( .A1(_AES_ENC_us00_n461 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n509 ) );
NOR2_X2 _AES_ENC_us00_U120  ( .A1(_AES_ENC_us00_n512 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n508 ) );
NOR2_X2 _AES_ENC_us00_U119  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n600 ), .ZN(_AES_ENC_us00_n510 ) );
NOR4_X2 _AES_ENC_us00_U118  ( .A1(_AES_ENC_us00_n508 ), .A2(_AES_ENC_us00_n509 ), .A3(_AES_ENC_us00_n510 ), .A4(_AES_ENC_us00_n511 ), .ZN(_AES_ENC_us00_n507 ) );
NOR2_X2 _AES_ENC_us00_U117  ( .A1(_AES_ENC_us00_n616 ), .A2(_AES_ENC_us00_n580 ), .ZN(_AES_ENC_us00_n425 ) );
NOR2_X2 _AES_ENC_us00_U116  ( .A1(_AES_ENC_us00_n90 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n424 ) );
NOR2_X2 _AES_ENC_us00_U115  ( .A1(_AES_ENC_us00_n610 ), .A2(_AES_ENC_us00_n599 ), .ZN(_AES_ENC_us00_n423 ) );
NOR4_X2 _AES_ENC_us00_U106  ( .A1(_AES_ENC_us00_n423 ), .A2(_AES_ENC_us00_n424 ), .A3(_AES_ENC_us00_n425 ), .A4(_AES_ENC_us00_n426 ), .ZN(_AES_ENC_us00_n422 ) );
NOR2_X2 _AES_ENC_us00_U105  ( .A1(_AES_ENC_us00_n416 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n412 ) );
NOR2_X2 _AES_ENC_us00_U104  ( .A1(_AES_ENC_us00_n76 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n414 ) );
NOR2_X2 _AES_ENC_us00_U103  ( .A1(_AES_ENC_us00_n415 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n413 ) );
NOR4_X2 _AES_ENC_us00_U102  ( .A1(_AES_ENC_us00_n316 ), .A2(_AES_ENC_us00_n412 ), .A3(_AES_ENC_us00_n413 ), .A4(_AES_ENC_us00_n414 ), .ZN(_AES_ENC_us00_n411 ) );
NOR2_X2 _AES_ENC_us00_U101  ( .A1(_AES_ENC_us00_n583 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n382 ) );
NOR2_X2 _AES_ENC_us00_U100  ( .A1(_AES_ENC_us00_n289 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n383 ) );
NOR3_X2 _AES_ENC_us00_U95  ( .A1(_AES_ENC_us00_n606 ), .A2(_AES_ENC_us00_n136 ), .A3(_AES_ENC_us00_n135 ), .ZN(_AES_ENC_us00_n381 ) );
NOR4_X2 _AES_ENC_us00_U94  ( .A1(_AES_ENC_us00_n381 ), .A2(_AES_ENC_us00_n382 ), .A3(_AES_ENC_us00_n383 ), .A4(_AES_ENC_us00_n384 ), .ZN(_AES_ENC_us00_n380 ) );
NOR2_X2 _AES_ENC_us00_U93  ( .A1(_AES_ENC_us00_n617 ), .A2(_AES_ENC_us00_n569 ), .ZN(_AES_ENC_us00_n475 ) );
NOR2_X2 _AES_ENC_us00_U92  ( .A1(_AES_ENC_us00_n163 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n473 ) );
NOR2_X2 _AES_ENC_us00_U91  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n97 ), .ZN(_AES_ENC_us00_n474 ) );
NOR4_X2 _AES_ENC_us00_U90  ( .A1(_AES_ENC_us00_n472 ), .A2(_AES_ENC_us00_n473 ), .A3(_AES_ENC_us00_n474 ), .A4(_AES_ENC_us00_n475 ), .ZN(_AES_ENC_us00_n471 ) );
NOR2_X2 _AES_ENC_us00_U89  ( .A1(_AES_ENC_us00_n285 ), .A2(_AES_ENC_us00_n205 ), .ZN(_AES_ENC_us00_n186 ) );
NOR2_X2 _AES_ENC_us00_U88  ( .A1(_AES_ENC_us00_n182 ), .A2(_AES_ENC_us00_n573 ), .ZN(_AES_ENC_us00_n181 ) );
NOR2_X2 _AES_ENC_us00_U87  ( .A1(_AES_ENC_us00_n181 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n180 ) );
NOR4_X2 _AES_ENC_us00_U86  ( .A1(_AES_ENC_us00_n179 ), .A2(_AES_ENC_us00_n180 ), .A3(_AES_ENC_us00_n74 ), .A4(_AES_ENC_us00_n148 ), .ZN(_AES_ENC_us00_n178 ) );
NOR2_X2 _AES_ENC_us00_U81  ( .A1(_AES_ENC_us00_n199 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n197 ) );
NOR2_X2 _AES_ENC_us00_U80  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n577 ), .ZN(_AES_ENC_us00_n195 ) );
NOR2_X2 _AES_ENC_us00_U79  ( .A1(_AES_ENC_us00_n616 ), .A2(_AES_ENC_us00_n97 ), .ZN(_AES_ENC_us00_n196 ) );
NOR4_X2 _AES_ENC_us00_U78  ( .A1(_AES_ENC_us00_n195 ), .A2(_AES_ENC_us00_n196 ), .A3(_AES_ENC_us00_n197 ), .A4(_AES_ENC_us00_n198 ), .ZN(_AES_ENC_us00_n194 ) );
NOR2_X2 _AES_ENC_us00_U74  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n97 ), .ZN(_AES_ENC_us00_n499 ) );
NOR2_X2 _AES_ENC_us00_U73  ( .A1(_AES_ENC_us00_n620 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n238 ) );
NOR2_X2 _AES_ENC_us00_U72  ( .A1(_AES_ENC_us00_n285 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n212 ) );
NOR2_X2 _AES_ENC_us00_U71  ( .A1(_AES_ENC_us00_n140 ), .A2(_AES_ENC_us00_n90 ), .ZN(_AES_ENC_us00_n163 ) );
INV_X4 _AES_ENC_us00_U65  ( .A(_AES_ENC_us00_n144 ), .ZN(_AES_ENC_us00_n612 ) );
INV_X4 _AES_ENC_us00_U64  ( .A(_AES_ENC_us00_n122 ), .ZN(_AES_ENC_us00_n605 ) );
INV_X4 _AES_ENC_us00_U63  ( .A(_AES_ENC_us00_n121 ), .ZN(_AES_ENC_us00_n604 ) );
NOR2_X2 _AES_ENC_us00_U62  ( .A1(_AES_ENC_us00_n582 ), .A2(_AES_ENC_us00_n613 ), .ZN(_AES_ENC_us00_n316 ) );
NOR3_X2 _AES_ENC_us00_U61  ( .A1(_AES_ENC_us00_n370 ), .A2(_AES_ENC_us00_n72 ), .A3(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n250 ) );
INV_X4 _AES_ENC_us00_U59  ( .A(_AES_ENC_us00_n185 ), .ZN(_AES_ENC_us00_n608 ) );
NOR3_X2 _AES_ENC_us00_U58  ( .A1(_AES_ENC_us00_n573 ), .A2(_AES_ENC_us00_n165 ), .A3(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n74 ) );
INV_X4 _AES_ENC_us00_U57  ( .A(_AES_ENC_us00_n240 ), .ZN(_AES_ENC_us00_n615 ) );
NOR2_X2 _AES_ENC_us00_U50  ( .A1(_AES_ENC_us00_n623 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n182 ) );
NOR2_X2 _AES_ENC_us00_U49  ( .A1(_AES_ENC_us00_n620 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n286 ) );
NOR2_X2 _AES_ENC_us00_U48  ( .A1(_AES_ENC_us00_n569 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n103 ) );
NOR2_X2 _AES_ENC_us00_U47  ( .A1(_AES_ENC_us00_n622 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n205 ) );
NOR2_X2 _AES_ENC_us00_U46  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_us00_n72 ), .ZN(_AES_ENC_us00_n199 ) );
NOR2_X2 _AES_ENC_us00_U45  ( .A1(_AES_ENC_us00_n610 ), .A2(_AES_ENC_us00_n600 ), .ZN(_AES_ENC_us00_n568 ) );
NOR2_X2 _AES_ENC_us00_U44  ( .A1(_AES_ENC_us00_n576 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n330 ) );
NOR2_X2 _AES_ENC_us00_U43  ( .A1(_AES_ENC_us00_n603 ), .A2(_AES_ENC_us00_n610 ), .ZN(_AES_ENC_us00_n189 ) );
NOR2_X2 _AES_ENC_us00_U42  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n76 ), .ZN(_AES_ENC_us00_n75 ) );
NOR2_X2 _AES_ENC_us00_U41  ( .A1(_AES_ENC_us00_n74 ), .A2(_AES_ENC_us00_n75 ), .ZN(_AES_ENC_us00_n66 ) );
NOR2_X2 _AES_ENC_us00_U36  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n594 ), .ZN(_AES_ENC_us00_n567 ) );
NOR2_X2 _AES_ENC_us00_U35  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n290 ), .ZN(_AES_ENC_us00_n287 ) );
NOR2_X2 _AES_ENC_us00_U34  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n597 ), .ZN(_AES_ENC_us00_n538 ) );
NOR2_X2 _AES_ENC_us00_U33  ( .A1(_AES_ENC_us00_n77 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n501 ) );
NOR2_X2 _AES_ENC_us00_U32  ( .A1(_AES_ENC_us00_n116 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n111 ) );
NOR2_X2 _AES_ENC_us00_U31  ( .A1(_AES_ENC_us00_n255 ), .A2(_AES_ENC_us00_n608 ), .ZN(_AES_ENC_us00_n472 ) );
NOR2_X2 _AES_ENC_us00_U30  ( .A1(_AES_ENC_us00_n598 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n86 ) );
NOR2_X2 _AES_ENC_us00_U29  ( .A1(_AES_ENC_us00_n576 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n356 ) );
NOR2_X2 _AES_ENC_us00_U24  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n593 ), .ZN(_AES_ENC_us00_n563 ) );
NOR2_X2 _AES_ENC_us00_U23  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n114 ), .ZN(_AES_ENC_us00_n113 ) );
NOR2_X2 _AES_ENC_us00_U21  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n149 ), .ZN(_AES_ENC_us00_n384 ) );
NOR2_X2 _AES_ENC_us00_U20  ( .A1(_AES_ENC_us00_n186 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n235 ) );
NOR2_X2 _AES_ENC_us00_U19  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n601 ), .ZN(_AES_ENC_us00_n213 ) );
NOR2_X2 _AES_ENC_us00_U18  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n594 ), .ZN(_AES_ENC_us00_n439 ) );
NOR2_X2 _AES_ENC_us00_U17  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n590 ), .ZN(_AES_ENC_us00_n498 ) );
NOR2_X2 _AES_ENC_us00_U16  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n619 ), .ZN(_AES_ENC_us00_n488 ) );
NOR2_X2 _AES_ENC_us00_U15  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n582 ), .ZN(_AES_ENC_us00_n426 ) );
NOR2_X2 _AES_ENC_us00_U10  ( .A1(_AES_ENC_us00_n619 ), .A2(_AES_ENC_us00_n604 ), .ZN(_AES_ENC_us00_n393 ) );
NOR2_X2 _AES_ENC_us00_U9  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n315 ), .ZN(_AES_ENC_us00_n485 ) );
NOR2_X2 _AES_ENC_us00_U8  ( .A1(_AES_ENC_us00_n615 ), .A2(_AES_ENC_us00_n582 ), .ZN(_AES_ENC_us00_n329 ) );
NOR2_X2 _AES_ENC_us00_U7  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n599 ), .ZN(_AES_ENC_us00_n392 ) );
NOR2_X2 _AES_ENC_us00_U6  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n620 ), .ZN(_AES_ENC_us00_n148 ) );
OR2_X4 _AES_ENC_us00_U5  ( .A1(_AES_ENC_us00_n624 ), .A2(_AES_ENC_sa00[1]),.ZN(_AES_ENC_us00_n570 ) );
OR2_X4 _AES_ENC_us00_U4  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_sa00[4]),.ZN(_AES_ENC_us00_n569 ) );
NAND2_X2 _AES_ENC_us00_U514  ( .A1(_AES_ENC_us00_n72 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n164 ) );
AND2_X2 _AES_ENC_us00_U513  ( .A1(_AES_ENC_us00_n597 ), .A2(_AES_ENC_us00_n164 ), .ZN(_AES_ENC_us00_n145 ) );
NAND2_X2 _AES_ENC_us00_U511  ( .A1(_AES_ENC_us00_n145 ), .A2(_AES_ENC_us00_n402 ), .ZN(_AES_ENC_us00_n559 ) );
AND2_X2 _AES_ENC_us00_U493  ( .A1(_AES_ENC_us00_n417 ), .A2(_AES_ENC_us00_n199 ), .ZN(_AES_ENC_us00_n564 ) );
NAND4_X2 _AES_ENC_us00_U485  ( .A1(_AES_ENC_us00_n559 ), .A2(_AES_ENC_us00_n560 ), .A3(_AES_ENC_us00_n561 ), .A4(_AES_ENC_us00_n562 ), .ZN(_AES_ENC_us00_n558 ) );
NAND2_X2 _AES_ENC_us00_U484  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n558 ), .ZN(_AES_ENC_us00_n517 ) );
NAND2_X2 _AES_ENC_us00_U481  ( .A1(_AES_ENC_us00_n100 ), .A2(_AES_ENC_us00_n591 ), .ZN(_AES_ENC_us00_n548 ) );
NAND2_X2 _AES_ENC_us00_U476  ( .A1(_AES_ENC_us00_n601 ), .A2(_AES_ENC_us00_n590 ), .ZN(_AES_ENC_us00_n434 ) );
NAND2_X2 _AES_ENC_us00_U475  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n434 ), .ZN(_AES_ENC_us00_n549 ) );
NAND4_X2 _AES_ENC_us00_U457  ( .A1(_AES_ENC_us00_n548 ), .A2(_AES_ENC_us00_n549 ), .A3(_AES_ENC_us00_n550 ), .A4(_AES_ENC_us00_n551 ), .ZN(_AES_ENC_us00_n547 ) );
NAND2_X2 _AES_ENC_us00_U456  ( .A1(_AES_ENC_sa00[0]), .A2(_AES_ENC_us00_n547 ), .ZN(_AES_ENC_us00_n531 ) );
NAND2_X2 _AES_ENC_us00_U454  ( .A1(_AES_ENC_us00_n596 ), .A2(_AES_ENC_us00_n623 ), .ZN(_AES_ENC_us00_n341 ) );
NAND2_X2 _AES_ENC_us00_U453  ( .A1(_AES_ENC_us00_n587 ), .A2(_AES_ENC_us00_n341 ), .ZN(_AES_ENC_us00_n375 ) );
NAND2_X2 _AES_ENC_us00_U452  ( .A1(_AES_ENC_us00_n101 ), .A2(_AES_ENC_us00_n375 ), .ZN(_AES_ENC_us00_n534 ) );
NAND2_X2 _AES_ENC_us00_U451  ( .A1(_AES_ENC_us00_n619 ), .A2(_AES_ENC_us00_n589 ), .ZN(_AES_ENC_us00_n546 ) );
NAND2_X2 _AES_ENC_us00_U450  ( .A1(_AES_ENC_us00_n240 ), .A2(_AES_ENC_us00_n546 ), .ZN(_AES_ENC_us00_n535 ) );
NAND2_X2 _AES_ENC_us00_U449  ( .A1(_AES_ENC_us00_n626 ), .A2(_AES_ENC_us00_n627 ), .ZN(_AES_ENC_us00_n357 ) );
OR2_X2 _AES_ENC_us00_U446  ( .A1(_AES_ENC_us00_n357 ), .A2(_AES_ENC_us00_n264 ), .ZN(_AES_ENC_us00_n540 ) );
NAND2_X2 _AES_ENC_us00_U445  ( .A1(_AES_ENC_us00_n621 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n97 ) );
NAND2_X2 _AES_ENC_us00_U444  ( .A1(_AES_ENC_us00_n164 ), .A2(_AES_ENC_us00_n97 ), .ZN(_AES_ENC_us00_n545 ) );
NAND2_X2 _AES_ENC_us00_U443  ( .A1(_AES_ENC_us00_n79 ), .A2(_AES_ENC_us00_n545 ), .ZN(_AES_ENC_us00_n541 ) );
OR3_X2 _AES_ENC_us00_U440  ( .A1(_AES_ENC_us00_n115 ), .A2(_AES_ENC_sa00[7]), .A3(_AES_ENC_us00_n626 ), .ZN(_AES_ENC_us00_n542 ) );
NAND2_X2 _AES_ENC_us00_U439  ( .A1(_AES_ENC_us00_n593 ), .A2(_AES_ENC_us00_n601 ), .ZN(_AES_ENC_us00_n544 ) );
NAND4_X2 _AES_ENC_us00_U437  ( .A1(_AES_ENC_us00_n540 ), .A2(_AES_ENC_us00_n541 ), .A3(_AES_ENC_us00_n542 ), .A4(_AES_ENC_us00_n543 ), .ZN(_AES_ENC_us00_n539 ) );
NAND2_X2 _AES_ENC_us00_U436  ( .A1(_AES_ENC_sa00[2]), .A2(_AES_ENC_us00_n539 ), .ZN(_AES_ENC_us00_n536 ) );
NAND4_X2 _AES_ENC_us00_U432  ( .A1(_AES_ENC_us00_n534 ), .A2(_AES_ENC_us00_n535 ), .A3(_AES_ENC_us00_n536 ), .A4(_AES_ENC_us00_n537 ), .ZN(_AES_ENC_us00_n533 ) );
NAND2_X2 _AES_ENC_us00_U431  ( .A1(_AES_ENC_us00_n533 ), .A2(_AES_ENC_us00_n574 ), .ZN(_AES_ENC_us00_n532 ) );
NAND2_X2 _AES_ENC_us00_U430  ( .A1(_AES_ENC_us00_n531 ), .A2(_AES_ENC_us00_n532 ), .ZN(_AES_ENC_us00_n530 ) );
NAND2_X2 _AES_ENC_us00_U429  ( .A1(_AES_ENC_sa00[6]), .A2(_AES_ENC_us00_n530 ), .ZN(_AES_ENC_us00_n518 ) );
NAND2_X2 _AES_ENC_us00_U426  ( .A1(_AES_ENC_us00_n461 ), .A2(_AES_ENC_us00_n101 ), .ZN(_AES_ENC_us00_n521 ) );
NAND2_X2 _AES_ENC_us00_U425  ( .A1(_AES_ENC_us00_n588 ), .A2(_AES_ENC_us00_n597 ), .ZN(_AES_ENC_us00_n149 ) );
OR2_X2 _AES_ENC_us00_U424  ( .A1(_AES_ENC_us00_n149 ), .A2(_AES_ENC_us00_n605 ), .ZN(_AES_ENC_us00_n522 ) );
NAND2_X2 _AES_ENC_us00_U423  ( .A1(_AES_ENC_sa00[1]), .A2(_AES_ENC_us00_n620 ), .ZN(_AES_ENC_us00_n529 ) );
NAND2_X2 _AES_ENC_us00_U422  ( .A1(_AES_ENC_us00_n619 ), .A2(_AES_ENC_us00_n529 ), .ZN(_AES_ENC_us00_n123 ) );
NAND4_X2 _AES_ENC_us00_U412  ( .A1(_AES_ENC_us00_n521 ), .A2(_AES_ENC_us00_n522 ), .A3(_AES_ENC_us00_n523 ), .A4(_AES_ENC_us00_n524 ), .ZN(_AES_ENC_us00_n520 ) );
NAND2_X2 _AES_ENC_us00_U411  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n520 ), .ZN(_AES_ENC_us00_n519 ) );
NAND2_X2 _AES_ENC_us00_U408  ( .A1(_AES_ENC_us00_n396 ), .A2(_AES_ENC_us00_n173 ), .ZN(_AES_ENC_us00_n516 ) );
NAND2_X2 _AES_ENC_us00_U407  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n516 ), .ZN(_AES_ENC_us00_n515 ) );
AND2_X2 _AES_ENC_us00_U402  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n512 ), .ZN(_AES_ENC_us00_n514 ) );
NAND4_X2 _AES_ENC_us00_U395  ( .A1(_AES_ENC_us00_n505 ), .A2(_AES_ENC_us00_n581 ), .A3(_AES_ENC_us00_n506 ), .A4(_AES_ENC_us00_n507 ), .ZN(_AES_ENC_us00_n504 ) );
NAND2_X2 _AES_ENC_us00_U394  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n504 ), .ZN(_AES_ENC_us00_n463 ) );
NAND2_X2 _AES_ENC_us00_U392  ( .A1(_AES_ENC_us00_n218 ), .A2(_AES_ENC_us00_n144 ), .ZN(_AES_ENC_us00_n494 ) );
NAND2_X2 _AES_ENC_us00_U391  ( .A1(_AES_ENC_us00_n101 ), .A2(_AES_ENC_us00_n149 ), .ZN(_AES_ENC_us00_n495 ) );
NAND4_X2 _AES_ENC_us00_U381  ( .A1(_AES_ENC_us00_n494 ), .A2(_AES_ENC_us00_n495 ), .A3(_AES_ENC_us00_n496 ), .A4(_AES_ENC_us00_n497 ), .ZN(_AES_ENC_us00_n493 ) );
NAND2_X2 _AES_ENC_us00_U380  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n493 ), .ZN(_AES_ENC_us00_n464 ) );
AND2_X2 _AES_ENC_us00_U379  ( .A1(_AES_ENC_sa00[0]), .A2(_AES_ENC_sa00[6]),.ZN(_AES_ENC_us00_n80 ) );
NAND2_X2 _AES_ENC_us00_U378  ( .A1(_AES_ENC_us00_n601 ), .A2(_AES_ENC_us00_n164 ), .ZN(_AES_ENC_us00_n315 ) );
NAND2_X2 _AES_ENC_us00_U377  ( .A1(_AES_ENC_us00_n101 ), .A2(_AES_ENC_us00_n315 ), .ZN(_AES_ENC_us00_n481 ) );
NAND2_X2 _AES_ENC_us00_U376  ( .A1(_AES_ENC_us00_n185 ), .A2(_AES_ENC_us00_n600 ), .ZN(_AES_ENC_us00_n482 ) );
NAND2_X2 _AES_ENC_us00_U375  ( .A1(_AES_ENC_us00_n341 ), .A2(_AES_ENC_us00_n588 ), .ZN(_AES_ENC_us00_n76 ) );
XNOR2_X2 _AES_ENC_us00_U371  ( .A(_AES_ENC_us00_n611 ), .B(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n372 ) );
NAND4_X2 _AES_ENC_us00_U362  ( .A1(_AES_ENC_us00_n481 ), .A2(_AES_ENC_us00_n482 ), .A3(_AES_ENC_us00_n483 ), .A4(_AES_ENC_us00_n484 ), .ZN(_AES_ENC_us00_n480 ) );
NAND2_X2 _AES_ENC_us00_U361  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n480 ), .ZN(_AES_ENC_us00_n465 ) );
AND2_X2 _AES_ENC_us00_U360  ( .A1(_AES_ENC_sa00[6]), .A2(_AES_ENC_us00_n574 ), .ZN(_AES_ENC_us00_n62 ) );
NAND2_X2 _AES_ENC_us00_U359  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n479 ) );
NAND2_X2 _AES_ENC_us00_U358  ( .A1(_AES_ENC_us00_n165 ), .A2(_AES_ENC_us00_n479 ), .ZN(_AES_ENC_us00_n468 ) );
NAND2_X2 _AES_ENC_us00_U357  ( .A1(_AES_ENC_sa00[1]), .A2(_AES_ENC_us00_n624 ), .ZN(_AES_ENC_us00_n96 ) );
NAND2_X2 _AES_ENC_us00_U356  ( .A1(_AES_ENC_us00_n603 ), .A2(_AES_ENC_us00_n96 ), .ZN(_AES_ENC_us00_n478 ) );
NAND2_X2 _AES_ENC_us00_U355  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n478 ), .ZN(_AES_ENC_us00_n469 ) );
NAND4_X2 _AES_ENC_us00_U344  ( .A1(_AES_ENC_us00_n468 ), .A2(_AES_ENC_us00_n469 ), .A3(_AES_ENC_us00_n470 ), .A4(_AES_ENC_us00_n471 ), .ZN(_AES_ENC_us00_n467 ) );
NAND2_X2 _AES_ENC_us00_U343  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n467 ), .ZN(_AES_ENC_us00_n466 ) );
NAND4_X2 _AES_ENC_us00_U342  ( .A1(_AES_ENC_us00_n463 ), .A2(_AES_ENC_us00_n464 ), .A3(_AES_ENC_us00_n465 ), .A4(_AES_ENC_us00_n466 ), .ZN(_AES_ENC_sa00_sub[1] ) );
NAND2_X2 _AES_ENC_us00_U341  ( .A1(_AES_ENC_sa00[7]), .A2(_AES_ENC_us00_n611 ), .ZN(_AES_ENC_us00_n462 ) );
NAND2_X2 _AES_ENC_us00_U340  ( .A1(_AES_ENC_us00_n462 ), .A2(_AES_ENC_us00_n607 ), .ZN(_AES_ENC_us00_n458 ) );
OR4_X2 _AES_ENC_us00_U339  ( .A1(_AES_ENC_us00_n458 ), .A2(_AES_ENC_us00_n626 ), .A3(_AES_ENC_us00_n370 ), .A4(_AES_ENC_us00_n72 ), .ZN(_AES_ENC_us00_n450 ) );
NAND2_X2 _AES_ENC_us00_U337  ( .A1(_AES_ENC_us00_n93 ), .A2(_AES_ENC_us00_n587 ), .ZN(_AES_ENC_us00_n203 ) );
OR2_X2 _AES_ENC_us00_U336  ( .A1(_AES_ENC_us00_n610 ), .A2(_AES_ENC_us00_n461 ), .ZN(_AES_ENC_us00_n459 ) );
NAND2_X2 _AES_ENC_us00_U334  ( .A1(_AES_ENC_us00_n619 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n443 ) );
NAND2_X2 _AES_ENC_us00_U333  ( .A1(_AES_ENC_us00_n582 ), .A2(_AES_ENC_us00_n443 ), .ZN(_AES_ENC_us00_n114 ) );
NAND2_X2 _AES_ENC_us00_U332  ( .A1(_AES_ENC_us00_n146 ), .A2(_AES_ENC_us00_n576 ), .ZN(_AES_ENC_us00_n460 ) );
NAND2_X2 _AES_ENC_us00_U331  ( .A1(_AES_ENC_us00_n459 ), .A2(_AES_ENC_us00_n460 ), .ZN(_AES_ENC_us00_n457 ) );
NAND2_X2 _AES_ENC_us00_U330  ( .A1(_AES_ENC_us00_n457 ), .A2(_AES_ENC_us00_n458 ), .ZN(_AES_ENC_us00_n451 ) );
NAND2_X2 _AES_ENC_us00_U326  ( .A1(_AES_ENC_us00_n97 ), .A2(_AES_ENC_us00_n590 ), .ZN(_AES_ENC_us00_n290 ) );
NAND4_X2 _AES_ENC_us00_U323  ( .A1(_AES_ENC_us00_n450 ), .A2(_AES_ENC_us00_n203 ), .A3(_AES_ENC_us00_n451 ), .A4(_AES_ENC_us00_n452 ), .ZN(_AES_ENC_us00_n449 ) );
NAND2_X2 _AES_ENC_us00_U322  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n449 ), .ZN(_AES_ENC_us00_n403 ) );
NAND2_X2 _AES_ENC_us00_U321  ( .A1(_AES_ENC_us00_n584 ), .A2(_AES_ENC_us00_n341 ), .ZN(_AES_ENC_us00_n448 ) );
NAND2_X2 _AES_ENC_us00_U320  ( .A1(_AES_ENC_us00_n240 ), .A2(_AES_ENC_us00_n448 ), .ZN(_AES_ENC_us00_n436 ) );
NAND2_X2 _AES_ENC_us00_U313  ( .A1(_AES_ENC_us00_n590 ), .A2(_AES_ENC_us00_n443 ), .ZN(_AES_ENC_us00_n172 ) );
NAND4_X2 _AES_ENC_us00_U308  ( .A1(_AES_ENC_us00_n436 ), .A2(_AES_ENC_us00_n203 ), .A3(_AES_ENC_us00_n437 ), .A4(_AES_ENC_us00_n438 ), .ZN(_AES_ENC_us00_n435 ) );
NAND2_X2 _AES_ENC_us00_U307  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n435 ), .ZN(_AES_ENC_us00_n404 ) );
NAND2_X2 _AES_ENC_us00_U306  ( .A1(_AES_ENC_us00_n584 ), .A2(_AES_ENC_us00_n603 ), .ZN(_AES_ENC_us00_n206 ) );
NAND2_X2 _AES_ENC_us00_U305  ( .A1(_AES_ENC_us00_n144 ), .A2(_AES_ENC_us00_n206 ), .ZN(_AES_ENC_us00_n419 ) );
NAND2_X2 _AES_ENC_us00_U304  ( .A1(_AES_ENC_us00_n101 ), .A2(_AES_ENC_us00_n434 ), .ZN(_AES_ENC_us00_n420 ) );
XNOR2_X2 _AES_ENC_us00_U301  ( .A(_AES_ENC_sa00[7]), .B(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n237 ) );
NAND4_X2 _AES_ENC_us00_U289  ( .A1(_AES_ENC_us00_n419 ), .A2(_AES_ENC_us00_n420 ), .A3(_AES_ENC_us00_n421 ), .A4(_AES_ENC_us00_n422 ), .ZN(_AES_ENC_us00_n418 ) );
NAND2_X2 _AES_ENC_us00_U288  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n418 ), .ZN(_AES_ENC_us00_n405 ) );
NAND2_X2 _AES_ENC_us00_U287  ( .A1(_AES_ENC_us00_n138 ), .A2(_AES_ENC_us00_n144 ), .ZN(_AES_ENC_us00_n408 ) );
NAND2_X2 _AES_ENC_us00_U286  ( .A1(_AES_ENC_us00_n103 ), .A2(_AES_ENC_us00_n417 ), .ZN(_AES_ENC_us00_n409 ) );
NAND2_X2 _AES_ENC_us00_U285  ( .A1(_AES_ENC_us00_n240 ), .A2(_AES_ENC_sa00[1]), .ZN(_AES_ENC_us00_n410 ) );
NAND4_X2 _AES_ENC_us00_U278  ( .A1(_AES_ENC_us00_n408 ), .A2(_AES_ENC_us00_n409 ), .A3(_AES_ENC_us00_n410 ), .A4(_AES_ENC_us00_n411 ), .ZN(_AES_ENC_us00_n407 ) );
NAND2_X2 _AES_ENC_us00_U277  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n407 ), .ZN(_AES_ENC_us00_n406 ) );
NAND4_X2 _AES_ENC_us00_U276  ( .A1(_AES_ENC_us00_n403 ), .A2(_AES_ENC_us00_n404 ), .A3(_AES_ENC_us00_n405 ), .A4(_AES_ENC_us00_n406 ), .ZN(_AES_ENC_sa00_sub[2] ) );
NAND2_X2 _AES_ENC_us00_U275  ( .A1(_AES_ENC_us00_n135 ), .A2(_AES_ENC_us00_n402 ), .ZN(_AES_ENC_us00_n386 ) );
NAND2_X2 _AES_ENC_us00_U274  ( .A1(_AES_ENC_us00_n145 ), .A2(_AES_ENC_us00_n240 ), .ZN(_AES_ENC_us00_n387 ) );
OR2_X2 _AES_ENC_us00_U266  ( .A1(_AES_ENC_us00_n97 ), .A2(_AES_ENC_us00_n606 ), .ZN(_AES_ENC_us00_n394 ) );
NAND2_X2 _AES_ENC_us00_U265  ( .A1(_AES_ENC_us00_n141 ), .A2(_AES_ENC_us00_n396 ), .ZN(_AES_ENC_us00_n395 ) );
NAND2_X2 _AES_ENC_us00_U264  ( .A1(_AES_ENC_us00_n394 ), .A2(_AES_ENC_us00_n395 ), .ZN(_AES_ENC_us00_n391 ) );
NAND4_X2 _AES_ENC_us00_U261  ( .A1(_AES_ENC_us00_n386 ), .A2(_AES_ENC_us00_n387 ), .A3(_AES_ENC_us00_n388 ), .A4(_AES_ENC_us00_n389 ), .ZN(_AES_ENC_us00_n385 ) );
NAND2_X2 _AES_ENC_us00_U260  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n385 ), .ZN(_AES_ENC_us00_n344 ) );
OR2_X2 _AES_ENC_us00_U259  ( .A1(_AES_ENC_us00_n172 ), .A2(_AES_ENC_us00_n617 ), .ZN(_AES_ENC_us00_n377 ) );
OR2_X2 _AES_ENC_us00_U257  ( .A1(_AES_ENC_us00_n570 ), .A2(_AES_ENC_us00_n266 ), .ZN(_AES_ENC_us00_n378 ) );
NAND2_X2 _AES_ENC_us00_U256  ( .A1(_AES_ENC_us00_n182 ), .A2(_AES_ENC_us00_n100 ), .ZN(_AES_ENC_us00_n379 ) );
NAND4_X2 _AES_ENC_us00_U249  ( .A1(_AES_ENC_us00_n377 ), .A2(_AES_ENC_us00_n378 ), .A3(_AES_ENC_us00_n379 ), .A4(_AES_ENC_us00_n380 ), .ZN(_AES_ENC_us00_n376 ) );
NAND2_X2 _AES_ENC_us00_U248  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n376 ), .ZN(_AES_ENC_us00_n345 ) );
NAND2_X2 _AES_ENC_us00_U247  ( .A1(_AES_ENC_us00_n240 ), .A2(_AES_ENC_us00_n114 ), .ZN(_AES_ENC_us00_n361 ) );
NAND2_X2 _AES_ENC_us00_U246  ( .A1(_AES_ENC_us00_n570 ), .A2(_AES_ENC_us00_n164 ), .ZN(_AES_ENC_us00_n147 ) );
OR2_X2 _AES_ENC_us00_U245  ( .A1(_AES_ENC_us00_n147 ), .A2(_AES_ENC_us00_n612 ), .ZN(_AES_ENC_us00_n362 ) );
NAND2_X2 _AES_ENC_us00_U244  ( .A1(_AES_ENC_us00_n122 ), .A2(_AES_ENC_us00_n589 ), .ZN(_AES_ENC_us00_n363 ) );
NAND4_X2 _AES_ENC_us00_U233  ( .A1(_AES_ENC_us00_n361 ), .A2(_AES_ENC_us00_n362 ), .A3(_AES_ENC_us00_n363 ), .A4(_AES_ENC_us00_n364 ), .ZN(_AES_ENC_us00_n360 ) );
NAND2_X2 _AES_ENC_us00_U232  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n360 ), .ZN(_AES_ENC_us00_n346 ) );
NAND2_X2 _AES_ENC_us00_U231  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n623 ), .ZN(_AES_ENC_us00_n349 ) );
NAND2_X2 _AES_ENC_us00_U230  ( .A1(_AES_ENC_us00_n144 ), .A2(_AES_ENC_us00_n123 ), .ZN(_AES_ENC_us00_n350 ) );
OR2_X2 _AES_ENC_us00_U224  ( .A1(_AES_ENC_us00_n141 ), .A2(_AES_ENC_us00_n285 ), .ZN(_AES_ENC_us00_n117 ) );
NAND4_X2 _AES_ENC_us00_U220  ( .A1(_AES_ENC_us00_n349 ), .A2(_AES_ENC_us00_n350 ), .A3(_AES_ENC_us00_n351 ), .A4(_AES_ENC_us00_n352 ), .ZN(_AES_ENC_us00_n348 ) );
NAND2_X2 _AES_ENC_us00_U219  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n348 ), .ZN(_AES_ENC_us00_n347 ) );
NAND4_X2 _AES_ENC_us00_U218  ( .A1(_AES_ENC_us00_n344 ), .A2(_AES_ENC_us00_n345 ), .A3(_AES_ENC_us00_n346 ), .A4(_AES_ENC_us00_n347 ), .ZN(_AES_ENC_sa00_sub[3] ) );
NAND2_X2 _AES_ENC_us00_U216  ( .A1(_AES_ENC_us00_n186 ), .A2(_AES_ENC_us00_n122 ), .ZN(_AES_ENC_us00_n334 ) );
NAND2_X2 _AES_ENC_us00_U215  ( .A1(_AES_ENC_us00_n603 ), .A2(_AES_ENC_us00_n577 ), .ZN(_AES_ENC_us00_n343 ) );
NAND2_X2 _AES_ENC_us00_U214  ( .A1(_AES_ENC_us00_n144 ), .A2(_AES_ENC_us00_n343 ), .ZN(_AES_ENC_us00_n335 ) );
NAND4_X2 _AES_ENC_us00_U206  ( .A1(_AES_ENC_us00_n334 ), .A2(_AES_ENC_us00_n335 ), .A3(_AES_ENC_us00_n336 ), .A4(_AES_ENC_us00_n337 ), .ZN(_AES_ENC_us00_n333 ) );
NAND2_X2 _AES_ENC_us00_U205  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n333 ), .ZN(_AES_ENC_us00_n291 ) );
NAND2_X2 _AES_ENC_us00_U204  ( .A1(_AES_ENC_us00_n185 ), .A2(_AES_ENC_us00_n206 ), .ZN(_AES_ENC_us00_n322 ) );
NAND2_X2 _AES_ENC_us00_U203  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n610 ), .ZN(_AES_ENC_us00_n332 ) );
NAND2_X2 _AES_ENC_us00_U202  ( .A1(_AES_ENC_us00_n267 ), .A2(_AES_ENC_us00_n332 ), .ZN(_AES_ENC_us00_n323 ) );
NAND4_X2 _AES_ENC_us00_U193  ( .A1(_AES_ENC_us00_n322 ), .A2(_AES_ENC_us00_n323 ), .A3(_AES_ENC_us00_n324 ), .A4(_AES_ENC_us00_n325 ), .ZN(_AES_ENC_us00_n321 ) );
NAND2_X2 _AES_ENC_us00_U192  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n321 ), .ZN(_AES_ENC_us00_n292 ) );
NAND2_X2 _AES_ENC_us00_U191  ( .A1(_AES_ENC_us00_n583 ), .A2(_AES_ENC_us00_n144 ), .ZN(_AES_ENC_us00_n307 ) );
NAND2_X2 _AES_ENC_us00_U190  ( .A1(_AES_ENC_us00_n101 ), .A2(_AES_ENC_us00_n587 ), .ZN(_AES_ENC_us00_n320 ) );
NAND2_X2 _AES_ENC_us00_U189  ( .A1(_AES_ENC_us00_n604 ), .A2(_AES_ENC_us00_n320 ), .ZN(_AES_ENC_us00_n319 ) );
NAND2_X2 _AES_ENC_us00_U188  ( .A1(_AES_ENC_us00_n319 ), .A2(_AES_ENC_us00_n623 ), .ZN(_AES_ENC_us00_n308 ) );
NAND4_X2 _AES_ENC_us00_U179  ( .A1(_AES_ENC_us00_n307 ), .A2(_AES_ENC_us00_n308 ), .A3(_AES_ENC_us00_n309 ), .A4(_AES_ENC_us00_n310 ), .ZN(_AES_ENC_us00_n306 ) );
NAND2_X2 _AES_ENC_us00_U178  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n306 ), .ZN(_AES_ENC_us00_n293 ) );
OR2_X2 _AES_ENC_us00_U177  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n135 ), .ZN(_AES_ENC_us00_n296 ) );
NAND2_X2 _AES_ENC_us00_U176  ( .A1(_AES_ENC_us00_n121 ), .A2(_AES_ENC_us00_n147 ), .ZN(_AES_ENC_us00_n297 ) );
NAND2_X2 _AES_ENC_us00_U175  ( .A1(_AES_ENC_us00_n100 ), .A2(_AES_ENC_us00_n595 ), .ZN(_AES_ENC_us00_n298 ) );
NAND4_X2 _AES_ENC_us00_U167  ( .A1(_AES_ENC_us00_n296 ), .A2(_AES_ENC_us00_n297 ), .A3(_AES_ENC_us00_n298 ), .A4(_AES_ENC_us00_n299 ), .ZN(_AES_ENC_us00_n295 ) );
NAND2_X2 _AES_ENC_us00_U166  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n295 ), .ZN(_AES_ENC_us00_n294 ) );
NAND4_X2 _AES_ENC_us00_U165  ( .A1(_AES_ENC_us00_n291 ), .A2(_AES_ENC_us00_n292 ), .A3(_AES_ENC_us00_n293 ), .A4(_AES_ENC_us00_n294 ), .ZN(_AES_ENC_sa00_sub[4] ) );
NAND2_X2 _AES_ENC_us00_U164  ( .A1(_AES_ENC_us00_n100 ), .A2(_AES_ENC_us00_n599 ), .ZN(_AES_ENC_us00_n274 ) );
NAND2_X2 _AES_ENC_us00_U163  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n206 ), .ZN(_AES_ENC_us00_n275 ) );
NAND4_X2 _AES_ENC_us00_U151  ( .A1(_AES_ENC_us00_n274 ), .A2(_AES_ENC_us00_n275 ), .A3(_AES_ENC_us00_n276 ), .A4(_AES_ENC_us00_n277 ), .ZN(_AES_ENC_us00_n273 ) );
NAND2_X2 _AES_ENC_us00_U150  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n273 ), .ZN(_AES_ENC_us00_n223 ) );
NAND2_X2 _AES_ENC_us00_U149  ( .A1(_AES_ENC_us00_n582 ), .A2(_AES_ENC_us00_n619 ), .ZN(_AES_ENC_us00_n272 ) );
NAND2_X2 _AES_ENC_us00_U148  ( .A1(_AES_ENC_us00_n121 ), .A2(_AES_ENC_us00_n272 ), .ZN(_AES_ENC_us00_n257 ) );
NAND2_X2 _AES_ENC_us00_U147  ( .A1(_AES_ENC_us00_n270 ), .A2(_AES_ENC_us00_n271 ), .ZN(_AES_ENC_us00_n269 ) );
NAND2_X2 _AES_ENC_us00_U146  ( .A1(_AES_ENC_us00_n606 ), .A2(_AES_ENC_us00_n269 ), .ZN(_AES_ENC_us00_n268 ) );
NAND2_X2 _AES_ENC_us00_U145  ( .A1(_AES_ENC_us00_n268 ), .A2(_AES_ENC_us00_n114 ), .ZN(_AES_ENC_us00_n258 ) );
OR2_X2 _AES_ENC_us00_U144  ( .A1(_AES_ENC_us00_n76 ), .A2(_AES_ENC_us00_n615 ), .ZN(_AES_ENC_us00_n259 ) );
NAND4_X2 _AES_ENC_us00_U139  ( .A1(_AES_ENC_us00_n257 ), .A2(_AES_ENC_us00_n258 ), .A3(_AES_ENC_us00_n259 ), .A4(_AES_ENC_us00_n260 ), .ZN(_AES_ENC_us00_n256 ) );
NAND2_X2 _AES_ENC_us00_U138  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n256 ), .ZN(_AES_ENC_us00_n224 ) );
OR2_X2 _AES_ENC_us00_U137  ( .A1(_AES_ENC_us00_n605 ), .A2(_AES_ENC_us00_n255 ), .ZN(_AES_ENC_us00_n242 ) );
NAND2_X2 _AES_ENC_us00_U136  ( .A1(_AES_ENC_us00_n97 ), .A2(_AES_ENC_us00_n577 ), .ZN(_AES_ENC_us00_n254 ) );
NAND2_X2 _AES_ENC_us00_U135  ( .A1(_AES_ENC_us00_n146 ), .A2(_AES_ENC_us00_n254 ), .ZN(_AES_ENC_us00_n253 ) );
NAND2_X2 _AES_ENC_us00_U134  ( .A1(_AES_ENC_us00_n612 ), .A2(_AES_ENC_us00_n253 ), .ZN(_AES_ENC_us00_n252 ) );
NAND2_X2 _AES_ENC_us00_U133  ( .A1(_AES_ENC_us00_n252 ), .A2(_AES_ENC_us00_n580 ), .ZN(_AES_ENC_us00_n243 ) );
NAND4_X2 _AES_ENC_us00_U125  ( .A1(_AES_ENC_us00_n242 ), .A2(_AES_ENC_us00_n243 ), .A3(_AES_ENC_us00_n244 ), .A4(_AES_ENC_us00_n245 ), .ZN(_AES_ENC_us00_n241 ) );
NAND2_X2 _AES_ENC_us00_U124  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n241 ), .ZN(_AES_ENC_us00_n225 ) );
NAND2_X2 _AES_ENC_us00_U123  ( .A1(_AES_ENC_us00_n100 ), .A2(_AES_ENC_us00_n123 ), .ZN(_AES_ENC_us00_n228 ) );
NAND2_X2 _AES_ENC_us00_U122  ( .A1(_AES_ENC_us00_n240 ), .A2(_AES_ENC_us00_n164 ), .ZN(_AES_ENC_us00_n229 ) );
NAND4_X2 _AES_ENC_us00_U114  ( .A1(_AES_ENC_us00_n228 ), .A2(_AES_ENC_us00_n229 ), .A3(_AES_ENC_us00_n230 ), .A4(_AES_ENC_us00_n231 ), .ZN(_AES_ENC_us00_n227 ) );
NAND2_X2 _AES_ENC_us00_U113  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n227 ), .ZN(_AES_ENC_us00_n226 ) );
NAND4_X2 _AES_ENC_us00_U112  ( .A1(_AES_ENC_us00_n223 ), .A2(_AES_ENC_us00_n224 ), .A3(_AES_ENC_us00_n225 ), .A4(_AES_ENC_us00_n226 ), .ZN(_AES_ENC_sa00_sub[5] ) );
NAND2_X2 _AES_ENC_us00_U111  ( .A1(_AES_ENC_us00_n570 ), .A2(_AES_ENC_us00_n96 ), .ZN(_AES_ENC_us00_n222 ) );
NAND2_X2 _AES_ENC_us00_U110  ( .A1(_AES_ENC_us00_n121 ), .A2(_AES_ENC_us00_n222 ), .ZN(_AES_ENC_us00_n208 ) );
NAND2_X2 _AES_ENC_us00_U109  ( .A1(_AES_ENC_us00_n221 ), .A2(_AES_ENC_us00_n117 ), .ZN(_AES_ENC_us00_n220 ) );
NAND2_X2 _AES_ENC_us00_U108  ( .A1(_AES_ENC_us00_n613 ), .A2(_AES_ENC_us00_n220 ), .ZN(_AES_ENC_us00_n219 ) );
NAND2_X2 _AES_ENC_us00_U107  ( .A1(_AES_ENC_us00_n218 ), .A2(_AES_ENC_us00_n219 ), .ZN(_AES_ENC_us00_n209 ) );
NAND4_X2 _AES_ENC_us00_U99  ( .A1(_AES_ENC_us00_n208 ), .A2(_AES_ENC_us00_n209 ), .A3(_AES_ENC_us00_n210 ), .A4(_AES_ENC_us00_n211 ), .ZN(_AES_ENC_us00_n207 ) );
NAND2_X2 _AES_ENC_us00_U98  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n207 ), .ZN(_AES_ENC_us00_n150 ) );
NAND2_X2 _AES_ENC_us00_U97  ( .A1(_AES_ENC_us00_n121 ), .A2(_AES_ENC_us00_n206 ), .ZN(_AES_ENC_us00_n191 ) );
NAND2_X2 _AES_ENC_us00_U96  ( .A1(_AES_ENC_us00_n102 ), .A2(_AES_ENC_us00_n619 ), .ZN(_AES_ENC_us00_n192 ) );
NAND4_X2 _AES_ENC_us00_U85  ( .A1(_AES_ENC_us00_n191 ), .A2(_AES_ENC_us00_n192 ), .A3(_AES_ENC_us00_n193 ), .A4(_AES_ENC_us00_n194 ), .ZN(_AES_ENC_us00_n190 ) );
NAND2_X2 _AES_ENC_us00_U84  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n190 ), .ZN(_AES_ENC_us00_n151 ) );
NAND2_X2 _AES_ENC_us00_U83  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n596 ), .ZN(_AES_ENC_us00_n175 ) );
NAND2_X2 _AES_ENC_us00_U82  ( .A1(_AES_ENC_us00_n144 ), .A2(_AES_ENC_us00_n624 ), .ZN(_AES_ENC_us00_n176 ) );
NAND2_X2 _AES_ENC_us00_U77  ( .A1(_AES_ENC_us00_n135 ), .A2(_AES_ENC_us00_n79 ), .ZN(_AES_ENC_us00_n183 ) );
NAND2_X2 _AES_ENC_us00_U76  ( .A1(_AES_ENC_us00_n185 ), .A2(_AES_ENC_us00_n592 ), .ZN(_AES_ENC_us00_n184 ) );
NAND2_X2 _AES_ENC_us00_U75  ( .A1(_AES_ENC_us00_n183 ), .A2(_AES_ENC_us00_n184 ), .ZN(_AES_ENC_us00_n179 ) );
NAND4_X2 _AES_ENC_us00_U70  ( .A1(_AES_ENC_us00_n175 ), .A2(_AES_ENC_us00_n176 ), .A3(_AES_ENC_us00_n177 ), .A4(_AES_ENC_us00_n178 ), .ZN(_AES_ENC_us00_n174 ) );
NAND2_X2 _AES_ENC_us00_U69  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n174 ), .ZN(_AES_ENC_us00_n152 ) );
NAND2_X2 _AES_ENC_us00_U68  ( .A1(_AES_ENC_us00_n173 ), .A2(_AES_ENC_us00_n101 ), .ZN(_AES_ENC_us00_n155 ) );
NAND2_X2 _AES_ENC_us00_U67  ( .A1(_AES_ENC_us00_n144 ), .A2(_AES_ENC_us00_n172 ), .ZN(_AES_ENC_us00_n156 ) );
NAND2_X2 _AES_ENC_us00_U66  ( .A1(_AES_ENC_us00_n171 ), .A2(_AES_ENC_us00_n123 ), .ZN(_AES_ENC_us00_n157 ) );
AND2_X2 _AES_ENC_us00_U60  ( .A1(_AES_ENC_us00_n164 ), .A2(_AES_ENC_us00_n602 ), .ZN(_AES_ENC_us00_n116 ) );
NAND4_X2 _AES_ENC_us00_U56  ( .A1(_AES_ENC_us00_n155 ), .A2(_AES_ENC_us00_n156 ), .A3(_AES_ENC_us00_n157 ), .A4(_AES_ENC_us00_n158 ), .ZN(_AES_ENC_us00_n154 ) );
NAND2_X2 _AES_ENC_us00_U55  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n154 ), .ZN(_AES_ENC_us00_n153 ) );
NAND4_X2 _AES_ENC_us00_U54  ( .A1(_AES_ENC_us00_n150 ), .A2(_AES_ENC_us00_n151 ), .A3(_AES_ENC_us00_n152 ), .A4(_AES_ENC_us00_n153 ), .ZN(_AES_ENC_sa00_sub[6] ) );
NAND2_X2 _AES_ENC_us00_U53  ( .A1(_AES_ENC_us00_n122 ), .A2(_AES_ENC_us00_n149 ), .ZN(_AES_ENC_us00_n126 ) );
NAND2_X2 _AES_ENC_us00_U52  ( .A1(_AES_ENC_us00_n148 ), .A2(_AES_ENC_us00_n582 ), .ZN(_AES_ENC_us00_n127 ) );
NAND2_X2 _AES_ENC_us00_U51  ( .A1(_AES_ENC_us00_n100 ), .A2(_AES_ENC_us00_n147 ), .ZN(_AES_ENC_us00_n128 ) );
NAND4_X2 _AES_ENC_us00_U40  ( .A1(_AES_ENC_us00_n126 ), .A2(_AES_ENC_us00_n127 ), .A3(_AES_ENC_us00_n128 ), .A4(_AES_ENC_us00_n129 ), .ZN(_AES_ENC_us00_n125 ) );
NAND2_X2 _AES_ENC_us00_U39  ( .A1(_AES_ENC_us00_n124 ), .A2(_AES_ENC_us00_n125 ), .ZN(_AES_ENC_us00_n58 ) );
NAND2_X2 _AES_ENC_us00_U38  ( .A1(_AES_ENC_us00_n122 ), .A2(_AES_ENC_us00_n123 ), .ZN(_AES_ENC_us00_n106 ) );
NAND2_X2 _AES_ENC_us00_U37  ( .A1(_AES_ENC_us00_n121 ), .A2(_AES_ENC_us00_n595 ), .ZN(_AES_ENC_us00_n107 ) );
NAND4_X2 _AES_ENC_us00_U28  ( .A1(_AES_ENC_us00_n106 ), .A2(_AES_ENC_us00_n107 ), .A3(_AES_ENC_us00_n108 ), .A4(_AES_ENC_us00_n109 ), .ZN(_AES_ENC_us00_n105 ) );
NAND2_X2 _AES_ENC_us00_U27  ( .A1(_AES_ENC_us00_n104 ), .A2(_AES_ENC_us00_n105 ), .ZN(_AES_ENC_us00_n59 ) );
NAND2_X2 _AES_ENC_us00_U26  ( .A1(_AES_ENC_us00_n103 ), .A2(_AES_ENC_us00_n101 ), .ZN(_AES_ENC_us00_n82 ) );
NAND2_X2 _AES_ENC_us00_U25  ( .A1(_AES_ENC_us00_n102 ), .A2(_AES_ENC_us00_n73 ), .ZN(_AES_ENC_us00_n83 ) );
AND2_X2 _AES_ENC_us00_U22  ( .A1(_AES_ENC_us00_n96 ), .A2(_AES_ENC_us00_n97 ), .ZN(_AES_ENC_us00_n95 ) );
NAND4_X2 _AES_ENC_us00_U14  ( .A1(_AES_ENC_us00_n82 ), .A2(_AES_ENC_us00_n83 ), .A3(_AES_ENC_us00_n84 ), .A4(_AES_ENC_us00_n85 ),.ZN(_AES_ENC_us00_n81 ) );
NAND2_X2 _AES_ENC_us00_U13  ( .A1(_AES_ENC_us00_n80 ), .A2(_AES_ENC_us00_n81 ), .ZN(_AES_ENC_us00_n60 ) );
NAND2_X2 _AES_ENC_us00_U12  ( .A1(_AES_ENC_us00_n78 ), .A2(_AES_ENC_us00_n79 ), .ZN(_AES_ENC_us00_n64 ) );
OR2_X2 _AES_ENC_us00_U11  ( .A1(_AES_ENC_us00_n608 ), .A2(_AES_ENC_us00_n77 ), .ZN(_AES_ENC_us00_n65 ) );
NAND4_X2 _AES_ENC_us00_U3  ( .A1(_AES_ENC_us00_n64 ), .A2(_AES_ENC_us00_n65 ), .A3(_AES_ENC_us00_n66 ), .A4(_AES_ENC_us00_n67 ), .ZN(_AES_ENC_us00_n63 ) );
NAND2_X2 _AES_ENC_us00_U2  ( .A1(_AES_ENC_us00_n62 ), .A2(_AES_ENC_us00_n63 ), .ZN(_AES_ENC_us00_n61 ) );
NAND4_X2 _AES_ENC_us00_U1  ( .A1(_AES_ENC_us00_n58 ), .A2(_AES_ENC_us00_n59 ), .A3(_AES_ENC_us00_n60 ), .A4(_AES_ENC_us00_n61 ), .ZN(_AES_ENC_sa00_sub[7] ));
INV_X4 _AES_ENC_us01_U575  ( .A(_AES_ENC_sa01[0]), .ZN(_AES_ENC_us01_n627 ));
INV_X4 _AES_ENC_us01_U574  ( .A(_AES_ENC_us01_n1053 ), .ZN(_AES_ENC_us01_n625 ) );
INV_X4 _AES_ENC_us01_U573  ( .A(_AES_ENC_us01_n1103 ), .ZN(_AES_ENC_us01_n623 ) );
INV_X4 _AES_ENC_us01_U572  ( .A(_AES_ENC_us01_n1056 ), .ZN(_AES_ENC_us01_n622 ) );
INV_X4 _AES_ENC_us01_U571  ( .A(_AES_ENC_us01_n1102 ), .ZN(_AES_ENC_us01_n621 ) );
INV_X4 _AES_ENC_us01_U570  ( .A(_AES_ENC_us01_n1074 ), .ZN(_AES_ENC_us01_n620 ) );
INV_X4 _AES_ENC_us01_U569  ( .A(_AES_ENC_us01_n929 ), .ZN(_AES_ENC_us01_n619 ) );
INV_X4 _AES_ENC_us01_U568  ( .A(_AES_ENC_us01_n1091 ), .ZN(_AES_ENC_us01_n618 ) );
INV_X4 _AES_ENC_us01_U567  ( .A(_AES_ENC_us01_n826 ), .ZN(_AES_ENC_us01_n617 ) );
INV_X4 _AES_ENC_us01_U566  ( .A(_AES_ENC_us01_n1031 ), .ZN(_AES_ENC_us01_n616 ) );
INV_X4 _AES_ENC_us01_U565  ( .A(_AES_ENC_us01_n1054 ), .ZN(_AES_ENC_us01_n615 ) );
INV_X4 _AES_ENC_us01_U564  ( .A(_AES_ENC_us01_n1025 ), .ZN(_AES_ENC_us01_n614 ) );
INV_X4 _AES_ENC_us01_U563  ( .A(_AES_ENC_us01_n990 ), .ZN(_AES_ENC_us01_n613 ) );
INV_X4 _AES_ENC_us01_U562  ( .A(_AES_ENC_sa01[4]), .ZN(_AES_ENC_us01_n612 ));
INV_X4 _AES_ENC_us01_U561  ( .A(_AES_ENC_us01_n881 ), .ZN(_AES_ENC_us01_n611 ) );
INV_X4 _AES_ENC_us01_U560  ( .A(_AES_ENC_us01_n1022 ), .ZN(_AES_ENC_us01_n610 ) );
INV_X4 _AES_ENC_us01_U559  ( .A(_AES_ENC_us01_n1120 ), .ZN(_AES_ENC_us01_n609 ) );
INV_X4 _AES_ENC_us01_U558  ( .A(_AES_ENC_us01_n977 ), .ZN(_AES_ENC_us01_n608 ) );
INV_X4 _AES_ENC_us01_U557  ( .A(_AES_ENC_us01_n926 ), .ZN(_AES_ENC_us01_n607 ) );
INV_X4 _AES_ENC_us01_U556  ( .A(_AES_ENC_us01_n910 ), .ZN(_AES_ENC_us01_n606 ) );
INV_X4 _AES_ENC_us01_U555  ( .A(_AES_ENC_us01_n1121 ), .ZN(_AES_ENC_us01_n605 ) );
INV_X4 _AES_ENC_us01_U554  ( .A(_AES_ENC_us01_n1009 ), .ZN(_AES_ENC_us01_n604 ) );
INV_X4 _AES_ENC_us01_U553  ( .A(_AES_ENC_us01_n1080 ), .ZN(_AES_ENC_us01_n602 ) );
INV_X4 _AES_ENC_us01_U552  ( .A(_AES_ENC_us01_n821 ), .ZN(_AES_ENC_us01_n600 ) );
INV_X4 _AES_ENC_us01_U551  ( .A(_AES_ENC_us01_n1013 ), .ZN(_AES_ENC_us01_n599 ) );
INV_X4 _AES_ENC_us01_U550  ( .A(_AES_ENC_us01_n1058 ), .ZN(_AES_ENC_us01_n598 ) );
INV_X4 _AES_ENC_us01_U549  ( .A(_AES_ENC_us01_n906 ), .ZN(_AES_ENC_us01_n597 ) );
INV_X4 _AES_ENC_us01_U548  ( .A(_AES_ENC_us01_n1048 ), .ZN(_AES_ENC_us01_n595 ) );
INV_X4 _AES_ENC_us01_U547  ( .A(_AES_ENC_us01_n974 ), .ZN(_AES_ENC_us01_n594 ) );
INV_X4 _AES_ENC_us01_U546  ( .A(_AES_ENC_sa01[2]), .ZN(_AES_ENC_us01_n593 ));
INV_X4 _AES_ENC_us01_U545  ( .A(_AES_ENC_us01_n800 ), .ZN(_AES_ENC_us01_n592 ) );
INV_X4 _AES_ENC_us01_U544  ( .A(_AES_ENC_us01_n925 ), .ZN(_AES_ENC_us01_n591 ) );
INV_X4 _AES_ENC_us01_U543  ( .A(_AES_ENC_us01_n824 ), .ZN(_AES_ENC_us01_n590 ) );
INV_X4 _AES_ENC_us01_U542  ( .A(_AES_ENC_us01_n959 ), .ZN(_AES_ENC_us01_n589 ) );
INV_X4 _AES_ENC_us01_U541  ( .A(_AES_ENC_us01_n779 ), .ZN(_AES_ENC_us01_n588 ) );
INV_X4 _AES_ENC_us01_U540  ( .A(_AES_ENC_us01_n794 ), .ZN(_AES_ENC_us01_n585 ) );
INV_X4 _AES_ENC_us01_U539  ( .A(_AES_ENC_us01_n880 ), .ZN(_AES_ENC_us01_n583 ) );
INV_X4 _AES_ENC_us01_U538  ( .A(_AES_ENC_sa01[7]), .ZN(_AES_ENC_us01_n581 ));
INV_X4 _AES_ENC_us01_U537  ( .A(_AES_ENC_us01_n992 ), .ZN(_AES_ENC_us01_n578 ) );
INV_X4 _AES_ENC_us01_U536  ( .A(_AES_ENC_us01_n1114 ), .ZN(_AES_ENC_us01_n577 ) );
INV_X4 _AES_ENC_us01_U535  ( .A(_AES_ENC_us01_n1092 ), .ZN(_AES_ENC_us01_n574 ) );
NOR2_X2 _AES_ENC_us01_U534  ( .A1(_AES_ENC_sa01[0]), .A2(_AES_ENC_sa01[6]),.ZN(_AES_ENC_us01_n1090 ) );
NOR2_X2 _AES_ENC_us01_U533  ( .A1(_AES_ENC_us01_n627 ), .A2(_AES_ENC_sa01[6]), .ZN(_AES_ENC_us01_n1070 ) );
NOR2_X2 _AES_ENC_us01_U532  ( .A1(_AES_ENC_sa01[4]), .A2(_AES_ENC_sa01[3]),.ZN(_AES_ENC_us01_n1025 ) );
INV_X4 _AES_ENC_us01_U531  ( .A(_AES_ENC_us01_n569 ), .ZN(_AES_ENC_us01_n572 ) );
NOR2_X2 _AES_ENC_us01_U530  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n765 ) );
NOR2_X2 _AES_ENC_us01_U529  ( .A1(_AES_ENC_sa01[4]), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n764 ) );
NOR2_X2 _AES_ENC_us01_U528  ( .A1(_AES_ENC_us01_n765 ), .A2(_AES_ENC_us01_n764 ), .ZN(_AES_ENC_us01_n766 ) );
NOR2_X2 _AES_ENC_us01_U527  ( .A1(_AES_ENC_us01_n766 ), .A2(_AES_ENC_us01_n589 ), .ZN(_AES_ENC_us01_n767 ) );
NOR3_X2 _AES_ENC_us01_U526  ( .A1(_AES_ENC_us01_n581 ), .A2(_AES_ENC_sa01[5]), .A3(_AES_ENC_us01_n704 ), .ZN(_AES_ENC_us01_n706 ));
NOR2_X2 _AES_ENC_us01_U525  ( .A1(_AES_ENC_us01_n1117 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n707 ) );
NOR2_X2 _AES_ENC_us01_U524  ( .A1(_AES_ENC_sa01[4]), .A2(_AES_ENC_us01_n574 ), .ZN(_AES_ENC_us01_n705 ) );
NOR3_X2 _AES_ENC_us01_U523  ( .A1(_AES_ENC_us01_n707 ), .A2(_AES_ENC_us01_n706 ), .A3(_AES_ENC_us01_n705 ), .ZN(_AES_ENC_us01_n713 ) );
INV_X4 _AES_ENC_us01_U522  ( .A(_AES_ENC_sa01[3]), .ZN(_AES_ENC_us01_n624 ));
NAND3_X2 _AES_ENC_us01_U521  ( .A1(_AES_ENC_us01_n652 ), .A2(_AES_ENC_us01_n596 ), .A3(_AES_ENC_sa01[7]), .ZN(_AES_ENC_us01_n653 ));
NOR2_X2 _AES_ENC_us01_U520  ( .A1(_AES_ENC_us01_n593 ), .A2(_AES_ENC_sa01[5]), .ZN(_AES_ENC_us01_n925 ) );
NOR2_X2 _AES_ENC_us01_U519  ( .A1(_AES_ENC_sa01[5]), .A2(_AES_ENC_sa01[2]),.ZN(_AES_ENC_us01_n974 ) );
INV_X4 _AES_ENC_us01_U518  ( .A(_AES_ENC_sa01[5]), .ZN(_AES_ENC_us01_n596 ));
NOR2_X2 _AES_ENC_us01_U517  ( .A1(_AES_ENC_us01_n593 ), .A2(_AES_ENC_sa01[7]), .ZN(_AES_ENC_us01_n779 ) );
NAND3_X2 _AES_ENC_us01_U516  ( .A1(_AES_ENC_us01_n679 ), .A2(_AES_ENC_us01_n678 ), .A3(_AES_ENC_us01_n677 ), .ZN(_AES_ENC_sa01_sub[0] ) );
NOR2_X2 _AES_ENC_us01_U515  ( .A1(_AES_ENC_us01_n596 ), .A2(_AES_ENC_sa01[2]), .ZN(_AES_ENC_us01_n1048 ) );
NOR4_X2 _AES_ENC_us01_U512  ( .A1(_AES_ENC_us01_n633 ), .A2(_AES_ENC_us01_n632 ), .A3(_AES_ENC_us01_n631 ), .A4(_AES_ENC_us01_n630 ), .ZN(_AES_ENC_us01_n634 ) );
NOR2_X2 _AES_ENC_us01_U510  ( .A1(_AES_ENC_us01_n629 ), .A2(_AES_ENC_us01_n628 ), .ZN(_AES_ENC_us01_n635 ) );
NAND3_X2 _AES_ENC_us01_U509  ( .A1(_AES_ENC_sa01[2]), .A2(_AES_ENC_sa01[7]), .A3(_AES_ENC_us01_n1059 ), .ZN(_AES_ENC_us01_n636 ) );
NOR2_X2 _AES_ENC_us01_U508  ( .A1(_AES_ENC_sa01[7]), .A2(_AES_ENC_sa01[2]),.ZN(_AES_ENC_us01_n794 ) );
NOR2_X2 _AES_ENC_us01_U507  ( .A1(_AES_ENC_sa01[4]), .A2(_AES_ENC_sa01[1]),.ZN(_AES_ENC_us01_n1102 ) );
NOR2_X2 _AES_ENC_us01_U506  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_sa01[3]), .ZN(_AES_ENC_us01_n1053 ) );
NOR2_X2 _AES_ENC_us01_U505  ( .A1(_AES_ENC_us01_n588 ), .A2(_AES_ENC_sa01[5]), .ZN(_AES_ENC_us01_n1024 ) );
NOR2_X2 _AES_ENC_us01_U504  ( .A1(_AES_ENC_us01_n577 ), .A2(_AES_ENC_sa01[2]), .ZN(_AES_ENC_us01_n1093 ) );
NOR2_X2 _AES_ENC_us01_U503  ( .A1(_AES_ENC_us01_n585 ), .A2(_AES_ENC_sa01[5]), .ZN(_AES_ENC_us01_n1094 ) );
NOR2_X2 _AES_ENC_us01_U502  ( .A1(_AES_ENC_us01_n612 ), .A2(_AES_ENC_sa01[3]), .ZN(_AES_ENC_us01_n931 ) );
INV_X4 _AES_ENC_us01_U501  ( .A(_AES_ENC_us01_n570 ), .ZN(_AES_ENC_us01_n573 ) );
NOR2_X2 _AES_ENC_us01_U500  ( .A1(_AES_ENC_us01_n1053 ), .A2(_AES_ENC_us01_n1095 ), .ZN(_AES_ENC_us01_n639 ) );
NOR3_X2 _AES_ENC_us01_U499  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n573 ), .A3(_AES_ENC_us01_n1074 ), .ZN(_AES_ENC_us01_n641 ) );
NOR2_X2 _AES_ENC_us01_U498  ( .A1(_AES_ENC_us01_n639 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n640 ) );
NOR2_X2 _AES_ENC_us01_U497  ( .A1(_AES_ENC_us01_n641 ), .A2(_AES_ENC_us01_n640 ), .ZN(_AES_ENC_us01_n646 ) );
NOR3_X2 _AES_ENC_us01_U496  ( .A1(_AES_ENC_us01_n995 ), .A2(_AES_ENC_us01_n578 ), .A3(_AES_ENC_us01_n994 ), .ZN(_AES_ENC_us01_n1002 ) );
NOR2_X2 _AES_ENC_us01_U495  ( .A1(_AES_ENC_us01_n909 ), .A2(_AES_ENC_us01_n908 ), .ZN(_AES_ENC_us01_n920 ) );
NOR2_X2 _AES_ENC_us01_U494  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n823 ) );
NOR2_X2 _AES_ENC_us01_U492  ( .A1(_AES_ENC_us01_n612 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n822 ) );
NOR2_X2 _AES_ENC_us01_U491  ( .A1(_AES_ENC_us01_n823 ), .A2(_AES_ENC_us01_n822 ), .ZN(_AES_ENC_us01_n825 ) );
NOR2_X2 _AES_ENC_us01_U490  ( .A1(_AES_ENC_sa01[1]), .A2(_AES_ENC_us01_n601 ), .ZN(_AES_ENC_us01_n913 ) );
NOR2_X2 _AES_ENC_us01_U489  ( .A1(_AES_ENC_us01_n913 ), .A2(_AES_ENC_us01_n1091 ), .ZN(_AES_ENC_us01_n914 ) );
NOR2_X2 _AES_ENC_us01_U488  ( .A1(_AES_ENC_us01_n826 ), .A2(_AES_ENC_us01_n572 ), .ZN(_AES_ENC_us01_n827 ) );
NOR3_X2 _AES_ENC_us01_U487  ( .A1(_AES_ENC_us01_n769 ), .A2(_AES_ENC_us01_n768 ), .A3(_AES_ENC_us01_n767 ), .ZN(_AES_ENC_us01_n775 ) );
NOR2_X2 _AES_ENC_us01_U486  ( .A1(_AES_ENC_us01_n1056 ), .A2(_AES_ENC_us01_n1053 ), .ZN(_AES_ENC_us01_n749 ) );
NOR2_X2 _AES_ENC_us01_U483  ( .A1(_AES_ENC_us01_n749 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n752 ) );
INV_X4 _AES_ENC_us01_U482  ( .A(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n626 ));
NOR2_X2 _AES_ENC_us01_U480  ( .A1(_AES_ENC_us01_n1054 ), .A2(_AES_ENC_us01_n1053 ), .ZN(_AES_ENC_us01_n1055 ) );
OR2_X4 _AES_ENC_us01_U479  ( .A1(_AES_ENC_us01_n1094 ), .A2(_AES_ENC_us01_n1093 ), .ZN(_AES_ENC_us01_n571 ) );
AND2_X2 _AES_ENC_us01_U478  ( .A1(_AES_ENC_us01_n571 ), .A2(_AES_ENC_us01_n1095 ), .ZN(_AES_ENC_us01_n1101 ) );
NOR2_X2 _AES_ENC_us01_U477  ( .A1(_AES_ENC_us01_n1074 ), .A2(_AES_ENC_us01_n931 ), .ZN(_AES_ENC_us01_n796 ) );
NOR2_X2 _AES_ENC_us01_U474  ( .A1(_AES_ENC_us01_n796 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n797 ) );
NOR2_X2 _AES_ENC_us01_U473  ( .A1(_AES_ENC_us01_n932 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n933 ) );
NOR2_X2 _AES_ENC_us01_U472  ( .A1(_AES_ENC_us01_n929 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n935 ) );
NOR2_X2 _AES_ENC_us01_U471  ( .A1(_AES_ENC_us01_n931 ), .A2(_AES_ENC_us01_n930 ), .ZN(_AES_ENC_us01_n934 ) );
NOR3_X2 _AES_ENC_us01_U470  ( .A1(_AES_ENC_us01_n935 ), .A2(_AES_ENC_us01_n934 ), .A3(_AES_ENC_us01_n933 ), .ZN(_AES_ENC_us01_n936 ) );
NOR2_X2 _AES_ENC_us01_U469  ( .A1(_AES_ENC_us01_n612 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n1075 ) );
NOR2_X2 _AES_ENC_us01_U468  ( .A1(_AES_ENC_us01_n572 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n949 ) );
NOR2_X2 _AES_ENC_us01_U467  ( .A1(_AES_ENC_us01_n1049 ), .A2(_AES_ENC_us01_n595 ), .ZN(_AES_ENC_us01_n1051 ) );
NOR2_X2 _AES_ENC_us01_U466  ( .A1(_AES_ENC_us01_n1051 ), .A2(_AES_ENC_us01_n1050 ), .ZN(_AES_ENC_us01_n1052 ) );
NOR2_X2 _AES_ENC_us01_U465  ( .A1(_AES_ENC_us01_n1052 ), .A2(_AES_ENC_us01_n604 ), .ZN(_AES_ENC_us01_n1064 ) );
NOR2_X2 _AES_ENC_us01_U464  ( .A1(_AES_ENC_sa01[1]), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n631 ) );
NOR2_X2 _AES_ENC_us01_U463  ( .A1(_AES_ENC_us01_n1025 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n980 ) );
NOR2_X2 _AES_ENC_us01_U462  ( .A1(_AES_ENC_us01_n1073 ), .A2(_AES_ENC_us01_n1094 ), .ZN(_AES_ENC_us01_n795 ) );
NOR2_X2 _AES_ENC_us01_U461  ( .A1(_AES_ENC_us01_n795 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n799 ) );
NOR2_X2 _AES_ENC_us01_U460  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n981 ) );
NOR2_X2 _AES_ENC_us01_U459  ( .A1(_AES_ENC_us01_n1102 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n643 ) );
NOR2_X2 _AES_ENC_us01_U458  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n624 ), .ZN(_AES_ENC_us01_n642 ) );
NOR2_X2 _AES_ENC_us01_U455  ( .A1(_AES_ENC_us01_n911 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n644 ) );
NOR4_X2 _AES_ENC_us01_U448  ( .A1(_AES_ENC_us01_n644 ), .A2(_AES_ENC_us01_n643 ), .A3(_AES_ENC_us01_n804 ), .A4(_AES_ENC_us01_n642 ), .ZN(_AES_ENC_us01_n645 ) );
NOR2_X2 _AES_ENC_us01_U447  ( .A1(_AES_ENC_us01_n1102 ), .A2(_AES_ENC_us01_n910 ), .ZN(_AES_ENC_us01_n932 ) );
NOR2_X2 _AES_ENC_us01_U442  ( .A1(_AES_ENC_us01_n1102 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n755 ) );
NOR2_X2 _AES_ENC_us01_U441  ( .A1(_AES_ENC_us01_n931 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n743 ) );
NOR2_X2 _AES_ENC_us01_U438  ( .A1(_AES_ENC_us01_n1072 ), .A2(_AES_ENC_us01_n1094 ), .ZN(_AES_ENC_us01_n930 ) );
NOR2_X2 _AES_ENC_us01_U435  ( .A1(_AES_ENC_us01_n1074 ), .A2(_AES_ENC_us01_n1025 ), .ZN(_AES_ENC_us01_n891 ) );
NOR2_X2 _AES_ENC_us01_U434  ( .A1(_AES_ENC_us01_n891 ), .A2(_AES_ENC_us01_n591 ), .ZN(_AES_ENC_us01_n894 ) );
NOR3_X2 _AES_ENC_us01_U433  ( .A1(_AES_ENC_us01_n601 ), .A2(_AES_ENC_sa01[1]), .A3(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n683 ));
INV_X4 _AES_ENC_us01_U428  ( .A(_AES_ENC_us01_n931 ), .ZN(_AES_ENC_us01_n601 ) );
NOR2_X2 _AES_ENC_us01_U427  ( .A1(_AES_ENC_us01_n996 ), .A2(_AES_ENC_us01_n931 ), .ZN(_AES_ENC_us01_n704 ) );
NOR2_X2 _AES_ENC_us01_U421  ( .A1(_AES_ENC_us01_n931 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n685 ) );
NOR2_X2 _AES_ENC_us01_U420  ( .A1(_AES_ENC_us01_n1029 ), .A2(_AES_ENC_us01_n1025 ), .ZN(_AES_ENC_us01_n1079 ) );
NOR3_X2 _AES_ENC_us01_U419  ( .A1(_AES_ENC_us01_n620 ), .A2(_AES_ENC_us01_n1025 ), .A3(_AES_ENC_us01_n594 ), .ZN(_AES_ENC_us01_n945 ) );
NOR2_X2 _AES_ENC_us01_U418  ( .A1(_AES_ENC_us01_n596 ), .A2(_AES_ENC_us01_n593 ), .ZN(_AES_ENC_us01_n800 ) );
NOR3_X2 _AES_ENC_us01_U417  ( .A1(_AES_ENC_us01_n598 ), .A2(_AES_ENC_us01_n581 ), .A3(_AES_ENC_us01_n593 ), .ZN(_AES_ENC_us01_n798 ) );
NOR3_X2 _AES_ENC_us01_U416  ( .A1(_AES_ENC_us01_n592 ), .A2(_AES_ENC_us01_n572 ), .A3(_AES_ENC_us01_n589 ), .ZN(_AES_ENC_us01_n962 ) );
NOR3_X2 _AES_ENC_us01_U415  ( .A1(_AES_ENC_us01_n959 ), .A2(_AES_ENC_us01_n572 ), .A3(_AES_ENC_us01_n591 ), .ZN(_AES_ENC_us01_n768 ) );
NOR3_X2 _AES_ENC_us01_U414  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n572 ), .A3(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n694 ) );
NOR3_X2 _AES_ENC_us01_U413  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n572 ), .A3(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n895 ) );
NOR3_X2 _AES_ENC_us01_U410  ( .A1(_AES_ENC_us01_n1008 ), .A2(_AES_ENC_us01_n1007 ), .A3(_AES_ENC_us01_n1006 ), .ZN(_AES_ENC_us01_n1018 ) );
NOR4_X2 _AES_ENC_us01_U409  ( .A1(_AES_ENC_us01_n806 ), .A2(_AES_ENC_us01_n805 ), .A3(_AES_ENC_us01_n804 ), .A4(_AES_ENC_us01_n803 ), .ZN(_AES_ENC_us01_n807 ) );
NOR3_X2 _AES_ENC_us01_U406  ( .A1(_AES_ENC_us01_n799 ), .A2(_AES_ENC_us01_n798 ), .A3(_AES_ENC_us01_n797 ), .ZN(_AES_ENC_us01_n808 ) );
NOR4_X2 _AES_ENC_us01_U405  ( .A1(_AES_ENC_us01_n843 ), .A2(_AES_ENC_us01_n842 ), .A3(_AES_ENC_us01_n841 ), .A4(_AES_ENC_us01_n840 ), .ZN(_AES_ENC_us01_n844 ) );
NOR2_X2 _AES_ENC_us01_U404  ( .A1(_AES_ENC_us01_n669 ), .A2(_AES_ENC_us01_n668 ), .ZN(_AES_ENC_us01_n673 ) );
NOR4_X2 _AES_ENC_us01_U403  ( .A1(_AES_ENC_us01_n946 ), .A2(_AES_ENC_us01_n1046 ), .A3(_AES_ENC_us01_n671 ), .A4(_AES_ENC_us01_n670 ), .ZN(_AES_ENC_us01_n672 ) );
NOR3_X2 _AES_ENC_us01_U401  ( .A1(_AES_ENC_us01_n1101 ), .A2(_AES_ENC_us01_n1100 ), .A3(_AES_ENC_us01_n1099 ), .ZN(_AES_ENC_us01_n1109 ) );
NOR4_X2 _AES_ENC_us01_U400  ( .A1(_AES_ENC_us01_n711 ), .A2(_AES_ENC_us01_n710 ), .A3(_AES_ENC_us01_n709 ), .A4(_AES_ENC_us01_n708 ), .ZN(_AES_ENC_us01_n712 ) );
NOR4_X2 _AES_ENC_us01_U399  ( .A1(_AES_ENC_us01_n963 ), .A2(_AES_ENC_us01_n962 ), .A3(_AES_ENC_us01_n961 ), .A4(_AES_ENC_us01_n960 ), .ZN(_AES_ENC_us01_n964 ) );
NOR3_X2 _AES_ENC_us01_U398  ( .A1(_AES_ENC_us01_n743 ), .A2(_AES_ENC_us01_n742 ), .A3(_AES_ENC_us01_n741 ), .ZN(_AES_ENC_us01_n744 ) );
NOR2_X2 _AES_ENC_us01_U397  ( .A1(_AES_ENC_us01_n697 ), .A2(_AES_ENC_us01_n658 ), .ZN(_AES_ENC_us01_n659 ) );
NOR2_X2 _AES_ENC_us01_U396  ( .A1(_AES_ENC_us01_n1078 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n1033 ) );
NOR2_X2 _AES_ENC_us01_U393  ( .A1(_AES_ENC_us01_n1031 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n1032 ) );
NOR3_X2 _AES_ENC_us01_U390  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n1025 ), .A3(_AES_ENC_us01_n1074 ), .ZN(_AES_ENC_us01_n1035 ) );
NOR4_X2 _AES_ENC_us01_U389  ( .A1(_AES_ENC_us01_n1035 ), .A2(_AES_ENC_us01_n1034 ), .A3(_AES_ENC_us01_n1033 ), .A4(_AES_ENC_us01_n1032 ), .ZN(_AES_ENC_us01_n1036 ) );
NOR2_X2 _AES_ENC_us01_U388  ( .A1(_AES_ENC_us01_n611 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n885 ) );
NOR2_X2 _AES_ENC_us01_U387  ( .A1(_AES_ENC_us01_n601 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n882 ) );
NOR2_X2 _AES_ENC_us01_U386  ( .A1(_AES_ENC_us01_n1053 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n884 ) );
NOR4_X2 _AES_ENC_us01_U385  ( .A1(_AES_ENC_us01_n885 ), .A2(_AES_ENC_us01_n884 ), .A3(_AES_ENC_us01_n883 ), .A4(_AES_ENC_us01_n882 ), .ZN(_AES_ENC_us01_n886 ) );
NOR2_X2 _AES_ENC_us01_U384  ( .A1(_AES_ENC_us01_n825 ), .A2(_AES_ENC_us01_n590 ), .ZN(_AES_ENC_us01_n830 ) );
NOR2_X2 _AES_ENC_us01_U383  ( .A1(_AES_ENC_us01_n827 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n829 ) );
NOR2_X2 _AES_ENC_us01_U382  ( .A1(_AES_ENC_us01_n572 ), .A2(_AES_ENC_us01_n574 ), .ZN(_AES_ENC_us01_n828 ) );
NOR4_X2 _AES_ENC_us01_U374  ( .A1(_AES_ENC_us01_n831 ), .A2(_AES_ENC_us01_n830 ), .A3(_AES_ENC_us01_n829 ), .A4(_AES_ENC_us01_n828 ), .ZN(_AES_ENC_us01_n832 ) );
NOR2_X2 _AES_ENC_us01_U373  ( .A1(_AES_ENC_us01_n587 ), .A2(_AES_ENC_us01_n603 ), .ZN(_AES_ENC_us01_n1104 ) );
NOR2_X2 _AES_ENC_us01_U372  ( .A1(_AES_ENC_us01_n1102 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n1106 ) );
NOR2_X2 _AES_ENC_us01_U370  ( .A1(_AES_ENC_us01_n1103 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n1105 ) );
NOR4_X2 _AES_ENC_us01_U369  ( .A1(_AES_ENC_us01_n1107 ), .A2(_AES_ENC_us01_n1106 ), .A3(_AES_ENC_us01_n1105 ), .A4(_AES_ENC_us01_n1104 ), .ZN(_AES_ENC_us01_n1108 ) );
NOR3_X2 _AES_ENC_us01_U368  ( .A1(_AES_ENC_us01_n959 ), .A2(_AES_ENC_us01_n624 ), .A3(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n963 ) );
NOR2_X2 _AES_ENC_us01_U367  ( .A1(_AES_ENC_us01_n596 ), .A2(_AES_ENC_us01_n581 ), .ZN(_AES_ENC_us01_n1114 ) );
INV_X4 _AES_ENC_us01_U366  ( .A(_AES_ENC_us01_n1024 ), .ZN(_AES_ENC_us01_n587 ) );
NOR3_X2 _AES_ENC_us01_U365  ( .A1(_AES_ENC_us01_n910 ), .A2(_AES_ENC_us01_n1059 ), .A3(_AES_ENC_us01_n593 ), .ZN(_AES_ENC_us01_n1115 ) );
INV_X4 _AES_ENC_us01_U364  ( .A(_AES_ENC_us01_n1094 ), .ZN(_AES_ENC_us01_n584 ) );
NOR2_X2 _AES_ENC_us01_U363  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n931 ), .ZN(_AES_ENC_us01_n1100 ) );
INV_X4 _AES_ENC_us01_U354  ( .A(_AES_ENC_us01_n1093 ), .ZN(_AES_ENC_us01_n575 ) );
NOR2_X2 _AES_ENC_us01_U353  ( .A1(_AES_ENC_us01_n569 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n929 ) );
NOR2_X2 _AES_ENC_us01_U352  ( .A1(_AES_ENC_us01_n609 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n926 ) );
NOR2_X2 _AES_ENC_us01_U351  ( .A1(_AES_ENC_us01_n572 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n1095 ) );
NOR2_X2 _AES_ENC_us01_U350  ( .A1(_AES_ENC_us01_n591 ), .A2(_AES_ENC_us01_n581 ), .ZN(_AES_ENC_us01_n1010 ) );
NOR2_X2 _AES_ENC_us01_U349  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n1103 ) );
NOR2_X2 _AES_ENC_us01_U348  ( .A1(_AES_ENC_us01_n614 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n1059 ) );
NOR2_X2 _AES_ENC_us01_U347  ( .A1(_AES_ENC_sa01[1]), .A2(_AES_ENC_us01_n1120 ), .ZN(_AES_ENC_us01_n1022 ) );
NOR2_X2 _AES_ENC_us01_U346  ( .A1(_AES_ENC_us01_n605 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n911 ) );
NOR2_X2 _AES_ENC_us01_U345  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_us01_n1025 ), .ZN(_AES_ENC_us01_n826 ) );
NOR2_X2 _AES_ENC_us01_U338  ( .A1(_AES_ENC_us01_n596 ), .A2(_AES_ENC_us01_n588 ), .ZN(_AES_ENC_us01_n1072 ) );
NOR2_X2 _AES_ENC_us01_U335  ( .A1(_AES_ENC_us01_n581 ), .A2(_AES_ENC_us01_n594 ), .ZN(_AES_ENC_us01_n956 ) );
NOR2_X2 _AES_ENC_us01_U329  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_us01_n612 ), .ZN(_AES_ENC_us01_n1121 ) );
NOR2_X2 _AES_ENC_us01_U328  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_us01_n612 ), .ZN(_AES_ENC_us01_n1058 ) );
NOR2_X2 _AES_ENC_us01_U327  ( .A1(_AES_ENC_us01_n577 ), .A2(_AES_ENC_us01_n593 ), .ZN(_AES_ENC_us01_n1073 ) );
NOR2_X2 _AES_ENC_us01_U325  ( .A1(_AES_ENC_sa01[1]), .A2(_AES_ENC_us01_n1025 ), .ZN(_AES_ENC_us01_n1054 ) );
NOR2_X2 _AES_ENC_us01_U324  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_us01_n931 ), .ZN(_AES_ENC_us01_n1029 ) );
NOR2_X2 _AES_ENC_us01_U319  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n1056 ) );
NOR2_X2 _AES_ENC_us01_U318  ( .A1(_AES_ENC_us01_n585 ), .A2(_AES_ENC_us01_n596 ), .ZN(_AES_ENC_us01_n1050 ) );
NOR2_X2 _AES_ENC_us01_U317  ( .A1(_AES_ENC_us01_n1121 ), .A2(_AES_ENC_us01_n1025 ), .ZN(_AES_ENC_us01_n1120 ) );
NOR2_X2 _AES_ENC_us01_U316  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_us01_n572 ), .ZN(_AES_ENC_us01_n1074 ) );
NOR2_X2 _AES_ENC_us01_U315  ( .A1(_AES_ENC_us01_n1058 ), .A2(_AES_ENC_us01_n1054 ), .ZN(_AES_ENC_us01_n878 ) );
NOR2_X2 _AES_ENC_us01_U314  ( .A1(_AES_ENC_us01_n878 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n879 ) );
NOR2_X2 _AES_ENC_us01_U312  ( .A1(_AES_ENC_us01_n880 ), .A2(_AES_ENC_us01_n879 ), .ZN(_AES_ENC_us01_n887 ) );
NOR2_X2 _AES_ENC_us01_U311  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n625 ), .ZN(_AES_ENC_us01_n957 ) );
NOR2_X2 _AES_ENC_us01_U310  ( .A1(_AES_ENC_us01_n958 ), .A2(_AES_ENC_us01_n957 ), .ZN(_AES_ENC_us01_n965 ) );
NOR3_X2 _AES_ENC_us01_U309  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n1091 ), .A3(_AES_ENC_us01_n1022 ), .ZN(_AES_ENC_us01_n720 ) );
NOR3_X2 _AES_ENC_us01_U303  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n1054 ), .A3(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n719 ) );
NOR2_X2 _AES_ENC_us01_U302  ( .A1(_AES_ENC_us01_n720 ), .A2(_AES_ENC_us01_n719 ), .ZN(_AES_ENC_us01_n726 ) );
NOR2_X2 _AES_ENC_us01_U300  ( .A1(_AES_ENC_us01_n585 ), .A2(_AES_ENC_us01_n613 ), .ZN(_AES_ENC_us01_n865 ) );
NOR2_X2 _AES_ENC_us01_U299  ( .A1(_AES_ENC_us01_n1059 ), .A2(_AES_ENC_us01_n1058 ), .ZN(_AES_ENC_us01_n1060 ) );
NOR2_X2 _AES_ENC_us01_U298  ( .A1(_AES_ENC_us01_n1095 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n668 ) );
NOR2_X2 _AES_ENC_us01_U297  ( .A1(_AES_ENC_us01_n911 ), .A2(_AES_ENC_us01_n910 ), .ZN(_AES_ENC_us01_n912 ) );
NOR2_X2 _AES_ENC_us01_U296  ( .A1(_AES_ENC_us01_n912 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n916 ) );
NOR2_X2 _AES_ENC_us01_U295  ( .A1(_AES_ENC_us01_n826 ), .A2(_AES_ENC_us01_n573 ), .ZN(_AES_ENC_us01_n750 ) );
NOR2_X2 _AES_ENC_us01_U294  ( .A1(_AES_ENC_us01_n750 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n751 ) );
NOR2_X2 _AES_ENC_us01_U293  ( .A1(_AES_ENC_us01_n907 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n908 ) );
NOR2_X2 _AES_ENC_us01_U292  ( .A1(_AES_ENC_us01_n990 ), .A2(_AES_ENC_us01_n926 ), .ZN(_AES_ENC_us01_n780 ) );
NOR2_X2 _AES_ENC_us01_U291  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n606 ), .ZN(_AES_ENC_us01_n838 ) );
NOR2_X2 _AES_ENC_us01_U290  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n621 ), .ZN(_AES_ENC_us01_n837 ) );
NOR2_X2 _AES_ENC_us01_U284  ( .A1(_AES_ENC_us01_n838 ), .A2(_AES_ENC_us01_n837 ), .ZN(_AES_ENC_us01_n845 ) );
NOR2_X2 _AES_ENC_us01_U283  ( .A1(_AES_ENC_us01_n1022 ), .A2(_AES_ENC_us01_n1058 ), .ZN(_AES_ENC_us01_n740 ) );
NOR2_X2 _AES_ENC_us01_U282  ( .A1(_AES_ENC_us01_n740 ), .A2(_AES_ENC_us01_n594 ), .ZN(_AES_ENC_us01_n742 ) );
NOR2_X2 _AES_ENC_us01_U281  ( .A1(_AES_ENC_us01_n1098 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n1099 ) );
NOR2_X2 _AES_ENC_us01_U280  ( .A1(_AES_ENC_us01_n1120 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n993 ) );
NOR2_X2 _AES_ENC_us01_U279  ( .A1(_AES_ENC_us01_n993 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n994 ) );
NOR2_X2 _AES_ENC_us01_U273  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n609 ), .ZN(_AES_ENC_us01_n1026 ) );
NOR2_X2 _AES_ENC_us01_U272  ( .A1(_AES_ENC_us01_n573 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n1027 ) );
NOR2_X2 _AES_ENC_us01_U271  ( .A1(_AES_ENC_us01_n1027 ), .A2(_AES_ENC_us01_n1026 ), .ZN(_AES_ENC_us01_n1028 ) );
NOR2_X2 _AES_ENC_us01_U270  ( .A1(_AES_ENC_us01_n1029 ), .A2(_AES_ENC_us01_n1028 ), .ZN(_AES_ENC_us01_n1034 ) );
NOR4_X2 _AES_ENC_us01_U269  ( .A1(_AES_ENC_us01_n757 ), .A2(_AES_ENC_us01_n756 ), .A3(_AES_ENC_us01_n755 ), .A4(_AES_ENC_us01_n754 ), .ZN(_AES_ENC_us01_n758 ) );
NOR2_X2 _AES_ENC_us01_U268  ( .A1(_AES_ENC_us01_n752 ), .A2(_AES_ENC_us01_n751 ), .ZN(_AES_ENC_us01_n759 ) );
NOR2_X2 _AES_ENC_us01_U267  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n1071 ), .ZN(_AES_ENC_us01_n669 ) );
NOR2_X2 _AES_ENC_us01_U263  ( .A1(_AES_ENC_us01_n1056 ), .A2(_AES_ENC_us01_n990 ), .ZN(_AES_ENC_us01_n991 ) );
NOR2_X2 _AES_ENC_us01_U262  ( .A1(_AES_ENC_us01_n991 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n995 ) );
NOR2_X2 _AES_ENC_us01_U258  ( .A1(_AES_ENC_us01_n588 ), .A2(_AES_ENC_us01_n598 ), .ZN(_AES_ENC_us01_n1008 ) );
NOR2_X2 _AES_ENC_us01_U255  ( .A1(_AES_ENC_us01_n839 ), .A2(_AES_ENC_us01_n603 ), .ZN(_AES_ENC_us01_n693 ) );
NOR2_X2 _AES_ENC_us01_U254  ( .A1(_AES_ENC_us01_n587 ), .A2(_AES_ENC_us01_n906 ), .ZN(_AES_ENC_us01_n741 ) );
NOR2_X2 _AES_ENC_us01_U253  ( .A1(_AES_ENC_us01_n1054 ), .A2(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n763 ) );
NOR2_X2 _AES_ENC_us01_U252  ( .A1(_AES_ENC_us01_n763 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n769 ) );
NOR2_X2 _AES_ENC_us01_U251  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n618 ), .ZN(_AES_ENC_us01_n1007 ) );
NOR2_X2 _AES_ENC_us01_U250  ( .A1(_AES_ENC_us01_n591 ), .A2(_AES_ENC_us01_n599 ), .ZN(_AES_ENC_us01_n1123 ) );
NOR2_X2 _AES_ENC_us01_U243  ( .A1(_AES_ENC_us01_n591 ), .A2(_AES_ENC_us01_n598 ), .ZN(_AES_ENC_us01_n710 ) );
INV_X4 _AES_ENC_us01_U242  ( .A(_AES_ENC_us01_n1029 ), .ZN(_AES_ENC_us01_n603 ) );
NOR2_X2 _AES_ENC_us01_U241  ( .A1(_AES_ENC_us01_n594 ), .A2(_AES_ENC_us01_n607 ), .ZN(_AES_ENC_us01_n883 ) );
NOR2_X2 _AES_ENC_us01_U240  ( .A1(_AES_ENC_us01_n623 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n1125 ) );
NOR2_X2 _AES_ENC_us01_U239  ( .A1(_AES_ENC_us01_n990 ), .A2(_AES_ENC_us01_n929 ), .ZN(_AES_ENC_us01_n892 ) );
NOR2_X2 _AES_ENC_us01_U238  ( .A1(_AES_ENC_us01_n892 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n893 ) );
NOR2_X2 _AES_ENC_us01_U237  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n621 ), .ZN(_AES_ENC_us01_n950 ) );
NOR2_X2 _AES_ENC_us01_U236  ( .A1(_AES_ENC_us01_n1079 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n1082 ) );
NOR2_X2 _AES_ENC_us01_U235  ( .A1(_AES_ENC_us01_n910 ), .A2(_AES_ENC_us01_n1056 ), .ZN(_AES_ENC_us01_n941 ) );
NOR2_X2 _AES_ENC_us01_U234  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n1077 ), .ZN(_AES_ENC_us01_n841 ) );
NOR2_X2 _AES_ENC_us01_U229  ( .A1(_AES_ENC_us01_n601 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n630 ) );
NOR2_X2 _AES_ENC_us01_U228  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n621 ), .ZN(_AES_ENC_us01_n806 ) );
NOR2_X2 _AES_ENC_us01_U227  ( .A1(_AES_ENC_us01_n601 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n948 ) );
NOR2_X2 _AES_ENC_us01_U226  ( .A1(_AES_ENC_us01_n587 ), .A2(_AES_ENC_us01_n620 ), .ZN(_AES_ENC_us01_n997 ) );
NOR2_X2 _AES_ENC_us01_U225  ( .A1(_AES_ENC_us01_n1121 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n1122 ) );
NOR2_X2 _AES_ENC_us01_U223  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n1023 ), .ZN(_AES_ENC_us01_n756 ) );
NOR2_X2 _AES_ENC_us01_U222  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n621 ), .ZN(_AES_ENC_us01_n870 ) );
NOR2_X2 _AES_ENC_us01_U221  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n569 ), .ZN(_AES_ENC_us01_n947 ) );
NOR2_X2 _AES_ENC_us01_U217  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n1077 ), .ZN(_AES_ENC_us01_n1084 ) );
NOR2_X2 _AES_ENC_us01_U213  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n855 ), .ZN(_AES_ENC_us01_n709 ) );
NOR2_X2 _AES_ENC_us01_U212  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n620 ), .ZN(_AES_ENC_us01_n868 ) );
NOR2_X2 _AES_ENC_us01_U211  ( .A1(_AES_ENC_us01_n1120 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n1124 ) );
NOR2_X2 _AES_ENC_us01_U210  ( .A1(_AES_ENC_us01_n1120 ), .A2(_AES_ENC_us01_n839 ), .ZN(_AES_ENC_us01_n842 ) );
NOR2_X2 _AES_ENC_us01_U209  ( .A1(_AES_ENC_us01_n1120 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n696 ) );
NOR2_X2 _AES_ENC_us01_U208  ( .A1(_AES_ENC_us01_n1074 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n1076 ) );
NOR2_X2 _AES_ENC_us01_U207  ( .A1(_AES_ENC_us01_n1074 ), .A2(_AES_ENC_us01_n609 ), .ZN(_AES_ENC_us01_n781 ) );
NOR3_X2 _AES_ENC_us01_U201  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n1056 ), .A3(_AES_ENC_us01_n990 ), .ZN(_AES_ENC_us01_n979 ) );
NOR3_X2 _AES_ENC_us01_U200  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n1058 ), .A3(_AES_ENC_us01_n1059 ), .ZN(_AES_ENC_us01_n854 ) );
NOR2_X2 _AES_ENC_us01_U199  ( .A1(_AES_ENC_us01_n996 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n869 ) );
NOR2_X2 _AES_ENC_us01_U198  ( .A1(_AES_ENC_us01_n1056 ), .A2(_AES_ENC_us01_n1074 ), .ZN(_AES_ENC_us01_n1057 ) );
NOR3_X2 _AES_ENC_us01_U197  ( .A1(_AES_ENC_us01_n588 ), .A2(_AES_ENC_us01_n1120 ), .A3(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n978 ) );
NOR2_X2 _AES_ENC_us01_U196  ( .A1(_AES_ENC_us01_n996 ), .A2(_AES_ENC_us01_n911 ), .ZN(_AES_ENC_us01_n1116 ) );
NOR2_X2 _AES_ENC_us01_U195  ( .A1(_AES_ENC_us01_n1074 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n754 ) );
NOR2_X2 _AES_ENC_us01_U194  ( .A1(_AES_ENC_us01_n926 ), .A2(_AES_ENC_us01_n1103 ), .ZN(_AES_ENC_us01_n977 ) );
NOR2_X2 _AES_ENC_us01_U187  ( .A1(_AES_ENC_us01_n839 ), .A2(_AES_ENC_us01_n824 ), .ZN(_AES_ENC_us01_n1092 ) );
NOR2_X2 _AES_ENC_us01_U186  ( .A1(_AES_ENC_us01_n573 ), .A2(_AES_ENC_us01_n1074 ), .ZN(_AES_ENC_us01_n684 ) );
NOR2_X2 _AES_ENC_us01_U185  ( .A1(_AES_ENC_us01_n826 ), .A2(_AES_ENC_us01_n1059 ), .ZN(_AES_ENC_us01_n907 ) );
NOR3_X2 _AES_ENC_us01_U184  ( .A1(_AES_ENC_us01_n577 ), .A2(_AES_ENC_us01_n1115 ), .A3(_AES_ENC_us01_n600 ), .ZN(_AES_ENC_us01_n831 ) );
NOR3_X2 _AES_ENC_us01_U183  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n1056 ), .A3(_AES_ENC_us01_n990 ), .ZN(_AES_ENC_us01_n896 ) );
NOR3_X2 _AES_ENC_us01_U182  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n573 ), .A3(_AES_ENC_us01_n1013 ), .ZN(_AES_ENC_us01_n670 ) );
NOR3_X2 _AES_ENC_us01_U181  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n1091 ), .A3(_AES_ENC_us01_n1022 ), .ZN(_AES_ENC_us01_n843 ) );
NOR2_X2 _AES_ENC_us01_U180  ( .A1(_AES_ENC_us01_n1029 ), .A2(_AES_ENC_us01_n1095 ), .ZN(_AES_ENC_us01_n735 ) );
NOR2_X2 _AES_ENC_us01_U174  ( .A1(_AES_ENC_us01_n1100 ), .A2(_AES_ENC_us01_n854 ), .ZN(_AES_ENC_us01_n860 ) );
NOR4_X2 _AES_ENC_us01_U173  ( .A1(_AES_ENC_us01_n1125 ), .A2(_AES_ENC_us01_n1124 ), .A3(_AES_ENC_us01_n1123 ), .A4(_AES_ENC_us01_n1122 ), .ZN(_AES_ENC_us01_n1126 ) );
NOR4_X2 _AES_ENC_us01_U172  ( .A1(_AES_ENC_us01_n1084 ), .A2(_AES_ENC_us01_n1083 ), .A3(_AES_ENC_us01_n1082 ), .A4(_AES_ENC_us01_n1081 ), .ZN(_AES_ENC_us01_n1085 ) );
NOR2_X2 _AES_ENC_us01_U171  ( .A1(_AES_ENC_us01_n1076 ), .A2(_AES_ENC_us01_n1075 ), .ZN(_AES_ENC_us01_n1086 ) );
NOR4_X2 _AES_ENC_us01_U170  ( .A1(_AES_ENC_us01_n983 ), .A2(_AES_ENC_us01_n982 ), .A3(_AES_ENC_us01_n981 ), .A4(_AES_ENC_us01_n980 ), .ZN(_AES_ENC_us01_n984 ) );
NOR2_X2 _AES_ENC_us01_U169  ( .A1(_AES_ENC_us01_n979 ), .A2(_AES_ENC_us01_n978 ), .ZN(_AES_ENC_us01_n985 ) );
NAND3_X2 _AES_ENC_us01_U168  ( .A1(_AES_ENC_us01_n569 ), .A2(_AES_ENC_us01_n603 ), .A3(_AES_ENC_us01_n681 ), .ZN(_AES_ENC_us01_n691 ) );
NOR2_X2 _AES_ENC_us01_U162  ( .A1(_AES_ENC_us01_n683 ), .A2(_AES_ENC_us01_n682 ), .ZN(_AES_ENC_us01_n690 ) );
NOR3_X2 _AES_ENC_us01_U161  ( .A1(_AES_ENC_us01_n695 ), .A2(_AES_ENC_us01_n694 ), .A3(_AES_ENC_us01_n693 ), .ZN(_AES_ENC_us01_n700 ) );
NOR4_X2 _AES_ENC_us01_U160  ( .A1(_AES_ENC_us01_n983 ), .A2(_AES_ENC_us01_n698 ), .A3(_AES_ENC_us01_n697 ), .A4(_AES_ENC_us01_n696 ), .ZN(_AES_ENC_us01_n699 ) );
NOR4_X2 _AES_ENC_us01_U159  ( .A1(_AES_ENC_us01_n896 ), .A2(_AES_ENC_us01_n895 ), .A3(_AES_ENC_us01_n894 ), .A4(_AES_ENC_us01_n893 ), .ZN(_AES_ENC_us01_n897 ) );
NOR2_X2 _AES_ENC_us01_U158  ( .A1(_AES_ENC_us01_n866 ), .A2(_AES_ENC_us01_n865 ), .ZN(_AES_ENC_us01_n872 ) );
NOR4_X2 _AES_ENC_us01_U157  ( .A1(_AES_ENC_us01_n870 ), .A2(_AES_ENC_us01_n869 ), .A3(_AES_ENC_us01_n868 ), .A4(_AES_ENC_us01_n867 ), .ZN(_AES_ENC_us01_n871 ) );
NOR2_X2 _AES_ENC_us01_U156  ( .A1(_AES_ENC_us01_n946 ), .A2(_AES_ENC_us01_n945 ), .ZN(_AES_ENC_us01_n952 ) );
NOR4_X2 _AES_ENC_us01_U155  ( .A1(_AES_ENC_us01_n950 ), .A2(_AES_ENC_us01_n949 ), .A3(_AES_ENC_us01_n948 ), .A4(_AES_ENC_us01_n947 ), .ZN(_AES_ENC_us01_n951 ) );
NOR3_X2 _AES_ENC_us01_U154  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n1054 ), .A3(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n961 ) );
NOR3_X2 _AES_ENC_us01_U153  ( .A1(_AES_ENC_us01_n609 ), .A2(_AES_ENC_us01_n1074 ), .A3(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n671 ) );
NOR2_X2 _AES_ENC_us01_U152  ( .A1(_AES_ENC_us01_n1057 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n1062 ) );
NOR2_X2 _AES_ENC_us01_U143  ( .A1(_AES_ENC_us01_n1055 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n1063 ) );
NOR2_X2 _AES_ENC_us01_U142  ( .A1(_AES_ENC_us01_n1060 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n1061 ) );
NOR4_X2 _AES_ENC_us01_U141  ( .A1(_AES_ENC_us01_n1064 ), .A2(_AES_ENC_us01_n1063 ), .A3(_AES_ENC_us01_n1062 ), .A4(_AES_ENC_us01_n1061 ), .ZN(_AES_ENC_us01_n1065 ) );
NOR2_X2 _AES_ENC_us01_U140  ( .A1(_AES_ENC_us01_n735 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n687 ) );
NOR2_X2 _AES_ENC_us01_U132  ( .A1(_AES_ENC_us01_n684 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n688 ) );
NOR2_X2 _AES_ENC_us01_U131  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n622 ), .ZN(_AES_ENC_us01_n686 ) );
NOR4_X2 _AES_ENC_us01_U130  ( .A1(_AES_ENC_us01_n688 ), .A2(_AES_ENC_us01_n687 ), .A3(_AES_ENC_us01_n686 ), .A4(_AES_ENC_us01_n685 ), .ZN(_AES_ENC_us01_n689 ) );
NOR2_X2 _AES_ENC_us01_U129  ( .A1(_AES_ENC_us01_n594 ), .A2(_AES_ENC_us01_n599 ), .ZN(_AES_ENC_us01_n771 ) );
NOR2_X2 _AES_ENC_us01_U128  ( .A1(_AES_ENC_us01_n1103 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n772 ) );
NOR2_X2 _AES_ENC_us01_U127  ( .A1(_AES_ENC_us01_n592 ), .A2(_AES_ENC_us01_n615 ), .ZN(_AES_ENC_us01_n773 ) );
NOR4_X2 _AES_ENC_us01_U126  ( .A1(_AES_ENC_us01_n773 ), .A2(_AES_ENC_us01_n772 ), .A3(_AES_ENC_us01_n771 ), .A4(_AES_ENC_us01_n770 ), .ZN(_AES_ENC_us01_n774 ) );
NOR2_X2 _AES_ENC_us01_U121  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n608 ), .ZN(_AES_ENC_us01_n858 ) );
NOR2_X2 _AES_ENC_us01_U120  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n855 ), .ZN(_AES_ENC_us01_n857 ) );
NOR2_X2 _AES_ENC_us01_U119  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n617 ), .ZN(_AES_ENC_us01_n856 ) );
NOR4_X2 _AES_ENC_us01_U118  ( .A1(_AES_ENC_us01_n858 ), .A2(_AES_ENC_us01_n857 ), .A3(_AES_ENC_us01_n856 ), .A4(_AES_ENC_us01_n958 ), .ZN(_AES_ENC_us01_n859 ) );
NOR3_X2 _AES_ENC_us01_U117  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n1120 ), .A3(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n918 ) );
NOR3_X2 _AES_ENC_us01_U116  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n573 ), .A3(_AES_ENC_us01_n1013 ), .ZN(_AES_ENC_us01_n917 ) );
NOR2_X2 _AES_ENC_us01_U115  ( .A1(_AES_ENC_us01_n914 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n915 ) );
NOR4_X2 _AES_ENC_us01_U106  ( .A1(_AES_ENC_us01_n918 ), .A2(_AES_ENC_us01_n917 ), .A3(_AES_ENC_us01_n916 ), .A4(_AES_ENC_us01_n915 ), .ZN(_AES_ENC_us01_n919 ) );
NOR2_X2 _AES_ENC_us01_U105  ( .A1(_AES_ENC_us01_n780 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n784 ) );
NOR2_X2 _AES_ENC_us01_U104  ( .A1(_AES_ENC_us01_n1117 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n782 ) );
NOR2_X2 _AES_ENC_us01_U103  ( .A1(_AES_ENC_us01_n781 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n783 ) );
NOR4_X2 _AES_ENC_us01_U102  ( .A1(_AES_ENC_us01_n880 ), .A2(_AES_ENC_us01_n784 ), .A3(_AES_ENC_us01_n783 ), .A4(_AES_ENC_us01_n782 ), .ZN(_AES_ENC_us01_n785 ) );
NOR2_X2 _AES_ENC_us01_U101  ( .A1(_AES_ENC_us01_n597 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n814 ) );
NOR2_X2 _AES_ENC_us01_U100  ( .A1(_AES_ENC_us01_n907 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n813 ) );
NOR3_X2 _AES_ENC_us01_U95  ( .A1(_AES_ENC_us01_n587 ), .A2(_AES_ENC_us01_n1058 ), .A3(_AES_ENC_us01_n1059 ), .ZN(_AES_ENC_us01_n815 ) );
NOR4_X2 _AES_ENC_us01_U94  ( .A1(_AES_ENC_us01_n815 ), .A2(_AES_ENC_us01_n814 ), .A3(_AES_ENC_us01_n813 ), .A4(_AES_ENC_us01_n812 ), .ZN(_AES_ENC_us01_n816 ) );
NOR2_X2 _AES_ENC_us01_U93  ( .A1(_AES_ENC_us01_n575 ), .A2(_AES_ENC_us01_n569 ), .ZN(_AES_ENC_us01_n721 ) );
NOR2_X2 _AES_ENC_us01_U92  ( .A1(_AES_ENC_us01_n1031 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n723 ) );
NOR2_X2 _AES_ENC_us01_U91  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n1096 ), .ZN(_AES_ENC_us01_n722 ) );
NOR4_X2 _AES_ENC_us01_U90  ( .A1(_AES_ENC_us01_n724 ), .A2(_AES_ENC_us01_n723 ), .A3(_AES_ENC_us01_n722 ), .A4(_AES_ENC_us01_n721 ), .ZN(_AES_ENC_us01_n725 ) );
NOR2_X2 _AES_ENC_us01_U89  ( .A1(_AES_ENC_us01_n911 ), .A2(_AES_ENC_us01_n990 ), .ZN(_AES_ENC_us01_n1009 ) );
NOR2_X2 _AES_ENC_us01_U88  ( .A1(_AES_ENC_us01_n1013 ), .A2(_AES_ENC_us01_n573 ), .ZN(_AES_ENC_us01_n1014 ) );
NOR2_X2 _AES_ENC_us01_U87  ( .A1(_AES_ENC_us01_n1014 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n1015 ) );
NOR4_X2 _AES_ENC_us01_U86  ( .A1(_AES_ENC_us01_n1016 ), .A2(_AES_ENC_us01_n1015 ), .A3(_AES_ENC_us01_n1119 ), .A4(_AES_ENC_us01_n1046 ), .ZN(_AES_ENC_us01_n1017 ) );
NOR2_X2 _AES_ENC_us01_U81  ( .A1(_AES_ENC_us01_n996 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n998 ) );
NOR2_X2 _AES_ENC_us01_U80  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n618 ), .ZN(_AES_ENC_us01_n1000 ) );
NOR2_X2 _AES_ENC_us01_U79  ( .A1(_AES_ENC_us01_n594 ), .A2(_AES_ENC_us01_n1096 ), .ZN(_AES_ENC_us01_n999 ) );
NOR4_X2 _AES_ENC_us01_U78  ( .A1(_AES_ENC_us01_n1000 ), .A2(_AES_ENC_us01_n999 ), .A3(_AES_ENC_us01_n998 ), .A4(_AES_ENC_us01_n997 ), .ZN(_AES_ENC_us01_n1001 ) );
NOR2_X2 _AES_ENC_us01_U74  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n1096 ), .ZN(_AES_ENC_us01_n697 ) );
NOR2_X2 _AES_ENC_us01_U73  ( .A1(_AES_ENC_us01_n609 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n958 ) );
NOR2_X2 _AES_ENC_us01_U72  ( .A1(_AES_ENC_us01_n911 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n983 ) );
NOR2_X2 _AES_ENC_us01_U71  ( .A1(_AES_ENC_us01_n1054 ), .A2(_AES_ENC_us01_n1103 ), .ZN(_AES_ENC_us01_n1031 ) );
INV_X4 _AES_ENC_us01_U65  ( .A(_AES_ENC_us01_n1050 ), .ZN(_AES_ENC_us01_n582 ) );
INV_X4 _AES_ENC_us01_U64  ( .A(_AES_ENC_us01_n1072 ), .ZN(_AES_ENC_us01_n586 ) );
INV_X4 _AES_ENC_us01_U63  ( .A(_AES_ENC_us01_n1073 ), .ZN(_AES_ENC_us01_n576 ) );
NOR2_X2 _AES_ENC_us01_U62  ( .A1(_AES_ENC_us01_n603 ), .A2(_AES_ENC_us01_n584 ), .ZN(_AES_ENC_us01_n880 ) );
NOR3_X2 _AES_ENC_us01_U61  ( .A1(_AES_ENC_us01_n826 ), .A2(_AES_ENC_us01_n1121 ), .A3(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n946 ) );
INV_X4 _AES_ENC_us01_U59  ( .A(_AES_ENC_us01_n1010 ), .ZN(_AES_ENC_us01_n579 ) );
NOR3_X2 _AES_ENC_us01_U58  ( .A1(_AES_ENC_us01_n573 ), .A2(_AES_ENC_us01_n1029 ), .A3(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n1119 ) );
INV_X4 _AES_ENC_us01_U57  ( .A(_AES_ENC_us01_n956 ), .ZN(_AES_ENC_us01_n580 ) );
NOR2_X2 _AES_ENC_us01_U50  ( .A1(_AES_ENC_us01_n601 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n1013 ) );
NOR2_X2 _AES_ENC_us01_U49  ( .A1(_AES_ENC_us01_n609 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n910 ) );
NOR2_X2 _AES_ENC_us01_U48  ( .A1(_AES_ENC_us01_n569 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n1091 ) );
NOR2_X2 _AES_ENC_us01_U47  ( .A1(_AES_ENC_us01_n614 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n990 ) );
NOR2_X2 _AES_ENC_us01_U46  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_us01_n1121 ), .ZN(_AES_ENC_us01_n996 ) );
NOR2_X2 _AES_ENC_us01_U45  ( .A1(_AES_ENC_us01_n592 ), .A2(_AES_ENC_us01_n622 ), .ZN(_AES_ENC_us01_n628 ) );
NOR2_X2 _AES_ENC_us01_U44  ( .A1(_AES_ENC_us01_n602 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n866 ) );
NOR2_X2 _AES_ENC_us01_U43  ( .A1(_AES_ENC_us01_n610 ), .A2(_AES_ENC_us01_n592 ), .ZN(_AES_ENC_us01_n1006 ) );
NOR2_X2 _AES_ENC_us01_U42  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n1117 ), .ZN(_AES_ENC_us01_n1118 ) );
NOR2_X2 _AES_ENC_us01_U41  ( .A1(_AES_ENC_us01_n1119 ), .A2(_AES_ENC_us01_n1118 ), .ZN(_AES_ENC_us01_n1127 ) );
NOR2_X2 _AES_ENC_us01_U36  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n616 ), .ZN(_AES_ENC_us01_n629 ) );
NOR2_X2 _AES_ENC_us01_U35  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n906 ), .ZN(_AES_ENC_us01_n909 ) );
NOR2_X2 _AES_ENC_us01_U34  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n607 ), .ZN(_AES_ENC_us01_n658 ) );
NOR2_X2 _AES_ENC_us01_U33  ( .A1(_AES_ENC_us01_n1116 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n695 ) );
NOR2_X2 _AES_ENC_us01_U32  ( .A1(_AES_ENC_us01_n1078 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n1083 ) );
NOR2_X2 _AES_ENC_us01_U31  ( .A1(_AES_ENC_us01_n941 ), .A2(_AES_ENC_us01_n579 ), .ZN(_AES_ENC_us01_n724 ) );
NOR2_X2 _AES_ENC_us01_U30  ( .A1(_AES_ENC_us01_n611 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n1107 ) );
NOR2_X2 _AES_ENC_us01_U29  ( .A1(_AES_ENC_us01_n602 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n840 ) );
NOR2_X2 _AES_ENC_us01_U24  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n623 ), .ZN(_AES_ENC_us01_n633 ) );
NOR2_X2 _AES_ENC_us01_U23  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n1080 ), .ZN(_AES_ENC_us01_n1081 ) );
NOR2_X2 _AES_ENC_us01_U21  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n1045 ), .ZN(_AES_ENC_us01_n812 ) );
NOR2_X2 _AES_ENC_us01_U20  ( .A1(_AES_ENC_us01_n1009 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n960 ) );
NOR2_X2 _AES_ENC_us01_U19  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n619 ), .ZN(_AES_ENC_us01_n982 ) );
NOR2_X2 _AES_ENC_us01_U18  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n616 ), .ZN(_AES_ENC_us01_n757 ) );
NOR2_X2 _AES_ENC_us01_U17  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n598 ), .ZN(_AES_ENC_us01_n698 ) );
NOR2_X2 _AES_ENC_us01_U16  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n605 ), .ZN(_AES_ENC_us01_n708 ) );
NOR2_X2 _AES_ENC_us01_U15  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n603 ), .ZN(_AES_ENC_us01_n770 ) );
NOR2_X2 _AES_ENC_us01_U10  ( .A1(_AES_ENC_us01_n605 ), .A2(_AES_ENC_us01_n576 ), .ZN(_AES_ENC_us01_n803 ) );
NOR2_X2 _AES_ENC_us01_U9  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n881 ), .ZN(_AES_ENC_us01_n711 ) );
NOR2_X2 _AES_ENC_us01_U8  ( .A1(_AES_ENC_us01_n580 ), .A2(_AES_ENC_us01_n603 ), .ZN(_AES_ENC_us01_n867 ) );
NOR2_X2 _AES_ENC_us01_U7  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n615 ), .ZN(_AES_ENC_us01_n804 ) );
NOR2_X2 _AES_ENC_us01_U6  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n609 ), .ZN(_AES_ENC_us01_n1046 ) );
OR2_X4 _AES_ENC_us01_U5  ( .A1(_AES_ENC_us01_n612 ), .A2(_AES_ENC_sa01[1]),.ZN(_AES_ENC_us01_n570 ) );
OR2_X4 _AES_ENC_us01_U4  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_sa01[4]),.ZN(_AES_ENC_us01_n569 ) );
NAND2_X2 _AES_ENC_us01_U514  ( .A1(_AES_ENC_us01_n1121 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n1030 ) );
AND2_X2 _AES_ENC_us01_U513  ( .A1(_AES_ENC_us01_n607 ), .A2(_AES_ENC_us01_n1030 ), .ZN(_AES_ENC_us01_n1049 ) );
NAND2_X2 _AES_ENC_us01_U511  ( .A1(_AES_ENC_us01_n1049 ), .A2(_AES_ENC_us01_n794 ), .ZN(_AES_ENC_us01_n637 ) );
AND2_X2 _AES_ENC_us01_U493  ( .A1(_AES_ENC_us01_n779 ), .A2(_AES_ENC_us01_n996 ), .ZN(_AES_ENC_us01_n632 ) );
NAND4_X2 _AES_ENC_us01_U485  ( .A1(_AES_ENC_us01_n637 ), .A2(_AES_ENC_us01_n636 ), .A3(_AES_ENC_us01_n635 ), .A4(_AES_ENC_us01_n634 ), .ZN(_AES_ENC_us01_n638 ) );
NAND2_X2 _AES_ENC_us01_U484  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n638 ), .ZN(_AES_ENC_us01_n679 ) );
NAND2_X2 _AES_ENC_us01_U481  ( .A1(_AES_ENC_us01_n1094 ), .A2(_AES_ENC_us01_n613 ), .ZN(_AES_ENC_us01_n648 ) );
NAND2_X2 _AES_ENC_us01_U476  ( .A1(_AES_ENC_us01_n619 ), .A2(_AES_ENC_us01_n598 ), .ZN(_AES_ENC_us01_n762 ) );
NAND2_X2 _AES_ENC_us01_U475  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n762 ), .ZN(_AES_ENC_us01_n647 ) );
NAND4_X2 _AES_ENC_us01_U457  ( .A1(_AES_ENC_us01_n648 ), .A2(_AES_ENC_us01_n647 ), .A3(_AES_ENC_us01_n646 ), .A4(_AES_ENC_us01_n645 ), .ZN(_AES_ENC_us01_n649 ) );
NAND2_X2 _AES_ENC_us01_U456  ( .A1(_AES_ENC_sa01[0]), .A2(_AES_ENC_us01_n649 ), .ZN(_AES_ENC_us01_n665 ) );
NAND2_X2 _AES_ENC_us01_U454  ( .A1(_AES_ENC_us01_n626 ), .A2(_AES_ENC_us01_n601 ), .ZN(_AES_ENC_us01_n855 ) );
NAND2_X2 _AES_ENC_us01_U453  ( .A1(_AES_ENC_us01_n617 ), .A2(_AES_ENC_us01_n855 ), .ZN(_AES_ENC_us01_n821 ) );
NAND2_X2 _AES_ENC_us01_U452  ( .A1(_AES_ENC_us01_n1093 ), .A2(_AES_ENC_us01_n821 ), .ZN(_AES_ENC_us01_n662 ) );
NAND2_X2 _AES_ENC_us01_U451  ( .A1(_AES_ENC_us01_n605 ), .A2(_AES_ENC_us01_n620 ), .ZN(_AES_ENC_us01_n650 ) );
NAND2_X2 _AES_ENC_us01_U450  ( .A1(_AES_ENC_us01_n956 ), .A2(_AES_ENC_us01_n650 ), .ZN(_AES_ENC_us01_n661 ) );
NAND2_X2 _AES_ENC_us01_U449  ( .A1(_AES_ENC_us01_n596 ), .A2(_AES_ENC_us01_n581 ), .ZN(_AES_ENC_us01_n839 ) );
OR2_X2 _AES_ENC_us01_U446  ( .A1(_AES_ENC_us01_n839 ), .A2(_AES_ENC_us01_n932 ), .ZN(_AES_ENC_us01_n656 ) );
NAND2_X2 _AES_ENC_us01_U445  ( .A1(_AES_ENC_us01_n624 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n1096 ) );
NAND2_X2 _AES_ENC_us01_U444  ( .A1(_AES_ENC_us01_n1030 ), .A2(_AES_ENC_us01_n1096 ), .ZN(_AES_ENC_us01_n651 ) );
NAND2_X2 _AES_ENC_us01_U443  ( .A1(_AES_ENC_us01_n1114 ), .A2(_AES_ENC_us01_n651 ), .ZN(_AES_ENC_us01_n655 ) );
OR3_X2 _AES_ENC_us01_U440  ( .A1(_AES_ENC_us01_n1079 ), .A2(_AES_ENC_sa01[7]), .A3(_AES_ENC_us01_n596 ), .ZN(_AES_ENC_us01_n654 ));
NAND2_X2 _AES_ENC_us01_U439  ( .A1(_AES_ENC_us01_n623 ), .A2(_AES_ENC_us01_n619 ), .ZN(_AES_ENC_us01_n652 ) );
NAND4_X2 _AES_ENC_us01_U437  ( .A1(_AES_ENC_us01_n656 ), .A2(_AES_ENC_us01_n655 ), .A3(_AES_ENC_us01_n654 ), .A4(_AES_ENC_us01_n653 ), .ZN(_AES_ENC_us01_n657 ) );
NAND2_X2 _AES_ENC_us01_U436  ( .A1(_AES_ENC_sa01[2]), .A2(_AES_ENC_us01_n657 ), .ZN(_AES_ENC_us01_n660 ) );
NAND4_X2 _AES_ENC_us01_U432  ( .A1(_AES_ENC_us01_n662 ), .A2(_AES_ENC_us01_n661 ), .A3(_AES_ENC_us01_n660 ), .A4(_AES_ENC_us01_n659 ), .ZN(_AES_ENC_us01_n663 ) );
NAND2_X2 _AES_ENC_us01_U431  ( .A1(_AES_ENC_us01_n663 ), .A2(_AES_ENC_us01_n627 ), .ZN(_AES_ENC_us01_n664 ) );
NAND2_X2 _AES_ENC_us01_U430  ( .A1(_AES_ENC_us01_n665 ), .A2(_AES_ENC_us01_n664 ), .ZN(_AES_ENC_us01_n666 ) );
NAND2_X2 _AES_ENC_us01_U429  ( .A1(_AES_ENC_sa01[6]), .A2(_AES_ENC_us01_n666 ), .ZN(_AES_ENC_us01_n678 ) );
NAND2_X2 _AES_ENC_us01_U426  ( .A1(_AES_ENC_us01_n735 ), .A2(_AES_ENC_us01_n1093 ), .ZN(_AES_ENC_us01_n675 ) );
NAND2_X2 _AES_ENC_us01_U425  ( .A1(_AES_ENC_us01_n625 ), .A2(_AES_ENC_us01_n607 ), .ZN(_AES_ENC_us01_n1045 ) );
OR2_X2 _AES_ENC_us01_U424  ( .A1(_AES_ENC_us01_n1045 ), .A2(_AES_ENC_us01_n586 ), .ZN(_AES_ENC_us01_n674 ) );
NAND2_X2 _AES_ENC_us01_U423  ( .A1(_AES_ENC_sa01[1]), .A2(_AES_ENC_us01_n609 ), .ZN(_AES_ENC_us01_n667 ) );
NAND2_X2 _AES_ENC_us01_U422  ( .A1(_AES_ENC_us01_n605 ), .A2(_AES_ENC_us01_n667 ), .ZN(_AES_ENC_us01_n1071 ) );
NAND4_X2 _AES_ENC_us01_U412  ( .A1(_AES_ENC_us01_n675 ), .A2(_AES_ENC_us01_n674 ), .A3(_AES_ENC_us01_n673 ), .A4(_AES_ENC_us01_n672 ), .ZN(_AES_ENC_us01_n676 ) );
NAND2_X2 _AES_ENC_us01_U411  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n676 ), .ZN(_AES_ENC_us01_n677 ) );
NAND2_X2 _AES_ENC_us01_U408  ( .A1(_AES_ENC_us01_n800 ), .A2(_AES_ENC_us01_n1022 ), .ZN(_AES_ENC_us01_n680 ) );
NAND2_X2 _AES_ENC_us01_U407  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n680 ), .ZN(_AES_ENC_us01_n681 ) );
AND2_X2 _AES_ENC_us01_U402  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n684 ), .ZN(_AES_ENC_us01_n682 ) );
NAND4_X2 _AES_ENC_us01_U395  ( .A1(_AES_ENC_us01_n691 ), .A2(_AES_ENC_us01_n583 ), .A3(_AES_ENC_us01_n690 ), .A4(_AES_ENC_us01_n689 ), .ZN(_AES_ENC_us01_n692 ) );
NAND2_X2 _AES_ENC_us01_U394  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n692 ), .ZN(_AES_ENC_us01_n733 ) );
NAND2_X2 _AES_ENC_us01_U392  ( .A1(_AES_ENC_us01_n977 ), .A2(_AES_ENC_us01_n1050 ), .ZN(_AES_ENC_us01_n702 ) );
NAND2_X2 _AES_ENC_us01_U391  ( .A1(_AES_ENC_us01_n1093 ), .A2(_AES_ENC_us01_n1045 ), .ZN(_AES_ENC_us01_n701 ) );
NAND4_X2 _AES_ENC_us01_U381  ( .A1(_AES_ENC_us01_n702 ), .A2(_AES_ENC_us01_n701 ), .A3(_AES_ENC_us01_n700 ), .A4(_AES_ENC_us01_n699 ), .ZN(_AES_ENC_us01_n703 ) );
NAND2_X2 _AES_ENC_us01_U380  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n703 ), .ZN(_AES_ENC_us01_n732 ) );
AND2_X2 _AES_ENC_us01_U379  ( .A1(_AES_ENC_sa01[0]), .A2(_AES_ENC_sa01[6]),.ZN(_AES_ENC_us01_n1113 ) );
NAND2_X2 _AES_ENC_us01_U378  ( .A1(_AES_ENC_us01_n619 ), .A2(_AES_ENC_us01_n1030 ), .ZN(_AES_ENC_us01_n881 ) );
NAND2_X2 _AES_ENC_us01_U377  ( .A1(_AES_ENC_us01_n1093 ), .A2(_AES_ENC_us01_n881 ), .ZN(_AES_ENC_us01_n715 ) );
NAND2_X2 _AES_ENC_us01_U376  ( .A1(_AES_ENC_us01_n1010 ), .A2(_AES_ENC_us01_n622 ), .ZN(_AES_ENC_us01_n714 ) );
NAND2_X2 _AES_ENC_us01_U375  ( .A1(_AES_ENC_us01_n855 ), .A2(_AES_ENC_us01_n625 ), .ZN(_AES_ENC_us01_n1117 ) );
XNOR2_X2 _AES_ENC_us01_U371  ( .A(_AES_ENC_us01_n593 ), .B(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n824 ) );
NAND4_X2 _AES_ENC_us01_U362  ( .A1(_AES_ENC_us01_n715 ), .A2(_AES_ENC_us01_n714 ), .A3(_AES_ENC_us01_n713 ), .A4(_AES_ENC_us01_n712 ), .ZN(_AES_ENC_us01_n716 ) );
NAND2_X2 _AES_ENC_us01_U361  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n716 ), .ZN(_AES_ENC_us01_n731 ) );
AND2_X2 _AES_ENC_us01_U360  ( .A1(_AES_ENC_sa01[6]), .A2(_AES_ENC_us01_n627 ), .ZN(_AES_ENC_us01_n1131 ) );
NAND2_X2 _AES_ENC_us01_U359  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n717 ) );
NAND2_X2 _AES_ENC_us01_U358  ( .A1(_AES_ENC_us01_n1029 ), .A2(_AES_ENC_us01_n717 ), .ZN(_AES_ENC_us01_n728 ) );
NAND2_X2 _AES_ENC_us01_U357  ( .A1(_AES_ENC_sa01[1]), .A2(_AES_ENC_us01_n612 ), .ZN(_AES_ENC_us01_n1097 ) );
NAND2_X2 _AES_ENC_us01_U356  ( .A1(_AES_ENC_us01_n610 ), .A2(_AES_ENC_us01_n1097 ), .ZN(_AES_ENC_us01_n718 ) );
NAND2_X2 _AES_ENC_us01_U355  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n718 ), .ZN(_AES_ENC_us01_n727 ) );
NAND4_X2 _AES_ENC_us01_U344  ( .A1(_AES_ENC_us01_n728 ), .A2(_AES_ENC_us01_n727 ), .A3(_AES_ENC_us01_n726 ), .A4(_AES_ENC_us01_n725 ), .ZN(_AES_ENC_us01_n729 ) );
NAND2_X2 _AES_ENC_us01_U343  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n729 ), .ZN(_AES_ENC_us01_n730 ) );
NAND4_X2 _AES_ENC_us01_U342  ( .A1(_AES_ENC_us01_n733 ), .A2(_AES_ENC_us01_n732 ), .A3(_AES_ENC_us01_n731 ), .A4(_AES_ENC_us01_n730 ), .ZN(_AES_ENC_sa01_sub[1] ) );
NAND2_X2 _AES_ENC_us01_U341  ( .A1(_AES_ENC_sa01[7]), .A2(_AES_ENC_us01_n593 ), .ZN(_AES_ENC_us01_n734 ) );
NAND2_X2 _AES_ENC_us01_U340  ( .A1(_AES_ENC_us01_n734 ), .A2(_AES_ENC_us01_n588 ), .ZN(_AES_ENC_us01_n738 ) );
OR4_X2 _AES_ENC_us01_U339  ( .A1(_AES_ENC_us01_n738 ), .A2(_AES_ENC_us01_n596 ), .A3(_AES_ENC_us01_n826 ), .A4(_AES_ENC_us01_n1121 ), .ZN(_AES_ENC_us01_n746 ) );
NAND2_X2 _AES_ENC_us01_U337  ( .A1(_AES_ENC_us01_n1100 ), .A2(_AES_ENC_us01_n617 ), .ZN(_AES_ENC_us01_n992 ) );
OR2_X2 _AES_ENC_us01_U336  ( .A1(_AES_ENC_us01_n592 ), .A2(_AES_ENC_us01_n735 ), .ZN(_AES_ENC_us01_n737 ) );
NAND2_X2 _AES_ENC_us01_U334  ( .A1(_AES_ENC_us01_n605 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n753 ) );
NAND2_X2 _AES_ENC_us01_U333  ( .A1(_AES_ENC_us01_n603 ), .A2(_AES_ENC_us01_n753 ), .ZN(_AES_ENC_us01_n1080 ) );
NAND2_X2 _AES_ENC_us01_U332  ( .A1(_AES_ENC_us01_n1048 ), .A2(_AES_ENC_us01_n602 ), .ZN(_AES_ENC_us01_n736 ) );
NAND2_X2 _AES_ENC_us01_U331  ( .A1(_AES_ENC_us01_n737 ), .A2(_AES_ENC_us01_n736 ), .ZN(_AES_ENC_us01_n739 ) );
NAND2_X2 _AES_ENC_us01_U330  ( .A1(_AES_ENC_us01_n739 ), .A2(_AES_ENC_us01_n738 ), .ZN(_AES_ENC_us01_n745 ) );
NAND2_X2 _AES_ENC_us01_U326  ( .A1(_AES_ENC_us01_n1096 ), .A2(_AES_ENC_us01_n598 ), .ZN(_AES_ENC_us01_n906 ) );
NAND4_X2 _AES_ENC_us01_U323  ( .A1(_AES_ENC_us01_n746 ), .A2(_AES_ENC_us01_n992 ), .A3(_AES_ENC_us01_n745 ), .A4(_AES_ENC_us01_n744 ), .ZN(_AES_ENC_us01_n747 ) );
NAND2_X2 _AES_ENC_us01_U322  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n747 ), .ZN(_AES_ENC_us01_n793 ) );
NAND2_X2 _AES_ENC_us01_U321  ( .A1(_AES_ENC_us01_n606 ), .A2(_AES_ENC_us01_n855 ), .ZN(_AES_ENC_us01_n748 ) );
NAND2_X2 _AES_ENC_us01_U320  ( .A1(_AES_ENC_us01_n956 ), .A2(_AES_ENC_us01_n748 ), .ZN(_AES_ENC_us01_n760 ) );
NAND2_X2 _AES_ENC_us01_U313  ( .A1(_AES_ENC_us01_n598 ), .A2(_AES_ENC_us01_n753 ), .ZN(_AES_ENC_us01_n1023 ) );
NAND4_X2 _AES_ENC_us01_U308  ( .A1(_AES_ENC_us01_n760 ), .A2(_AES_ENC_us01_n992 ), .A3(_AES_ENC_us01_n759 ), .A4(_AES_ENC_us01_n758 ), .ZN(_AES_ENC_us01_n761 ) );
NAND2_X2 _AES_ENC_us01_U307  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n761 ), .ZN(_AES_ENC_us01_n792 ) );
NAND2_X2 _AES_ENC_us01_U306  ( .A1(_AES_ENC_us01_n606 ), .A2(_AES_ENC_us01_n610 ), .ZN(_AES_ENC_us01_n989 ) );
NAND2_X2 _AES_ENC_us01_U305  ( .A1(_AES_ENC_us01_n1050 ), .A2(_AES_ENC_us01_n989 ), .ZN(_AES_ENC_us01_n777 ) );
NAND2_X2 _AES_ENC_us01_U304  ( .A1(_AES_ENC_us01_n1093 ), .A2(_AES_ENC_us01_n762 ), .ZN(_AES_ENC_us01_n776 ) );
XNOR2_X2 _AES_ENC_us01_U301  ( .A(_AES_ENC_sa01[7]), .B(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n959 ) );
NAND4_X2 _AES_ENC_us01_U289  ( .A1(_AES_ENC_us01_n777 ), .A2(_AES_ENC_us01_n776 ), .A3(_AES_ENC_us01_n775 ), .A4(_AES_ENC_us01_n774 ), .ZN(_AES_ENC_us01_n778 ) );
NAND2_X2 _AES_ENC_us01_U288  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n778 ), .ZN(_AES_ENC_us01_n791 ) );
NAND2_X2 _AES_ENC_us01_U287  ( .A1(_AES_ENC_us01_n1056 ), .A2(_AES_ENC_us01_n1050 ), .ZN(_AES_ENC_us01_n788 ) );
NAND2_X2 _AES_ENC_us01_U286  ( .A1(_AES_ENC_us01_n1091 ), .A2(_AES_ENC_us01_n779 ), .ZN(_AES_ENC_us01_n787 ) );
NAND2_X2 _AES_ENC_us01_U285  ( .A1(_AES_ENC_us01_n956 ), .A2(_AES_ENC_sa01[1]), .ZN(_AES_ENC_us01_n786 ) );
NAND4_X2 _AES_ENC_us01_U278  ( .A1(_AES_ENC_us01_n788 ), .A2(_AES_ENC_us01_n787 ), .A3(_AES_ENC_us01_n786 ), .A4(_AES_ENC_us01_n785 ), .ZN(_AES_ENC_us01_n789 ) );
NAND2_X2 _AES_ENC_us01_U277  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n789 ), .ZN(_AES_ENC_us01_n790 ) );
NAND4_X2 _AES_ENC_us01_U276  ( .A1(_AES_ENC_us01_n793 ), .A2(_AES_ENC_us01_n792 ), .A3(_AES_ENC_us01_n791 ), .A4(_AES_ENC_us01_n790 ), .ZN(_AES_ENC_sa01_sub[2] ) );
NAND2_X2 _AES_ENC_us01_U275  ( .A1(_AES_ENC_us01_n1059 ), .A2(_AES_ENC_us01_n794 ), .ZN(_AES_ENC_us01_n810 ) );
NAND2_X2 _AES_ENC_us01_U274  ( .A1(_AES_ENC_us01_n1049 ), .A2(_AES_ENC_us01_n956 ), .ZN(_AES_ENC_us01_n809 ) );
OR2_X2 _AES_ENC_us01_U266  ( .A1(_AES_ENC_us01_n1096 ), .A2(_AES_ENC_us01_n587 ), .ZN(_AES_ENC_us01_n802 ) );
NAND2_X2 _AES_ENC_us01_U265  ( .A1(_AES_ENC_us01_n1053 ), .A2(_AES_ENC_us01_n800 ), .ZN(_AES_ENC_us01_n801 ) );
NAND2_X2 _AES_ENC_us01_U264  ( .A1(_AES_ENC_us01_n802 ), .A2(_AES_ENC_us01_n801 ), .ZN(_AES_ENC_us01_n805 ) );
NAND4_X2 _AES_ENC_us01_U261  ( .A1(_AES_ENC_us01_n810 ), .A2(_AES_ENC_us01_n809 ), .A3(_AES_ENC_us01_n808 ), .A4(_AES_ENC_us01_n807 ), .ZN(_AES_ENC_us01_n811 ) );
NAND2_X2 _AES_ENC_us01_U260  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n811 ), .ZN(_AES_ENC_us01_n852 ) );
OR2_X2 _AES_ENC_us01_U259  ( .A1(_AES_ENC_us01_n1023 ), .A2(_AES_ENC_us01_n575 ), .ZN(_AES_ENC_us01_n819 ) );
OR2_X2 _AES_ENC_us01_U257  ( .A1(_AES_ENC_us01_n570 ), .A2(_AES_ENC_us01_n930 ), .ZN(_AES_ENC_us01_n818 ) );
NAND2_X2 _AES_ENC_us01_U256  ( .A1(_AES_ENC_us01_n1013 ), .A2(_AES_ENC_us01_n1094 ), .ZN(_AES_ENC_us01_n817 ) );
NAND4_X2 _AES_ENC_us01_U249  ( .A1(_AES_ENC_us01_n819 ), .A2(_AES_ENC_us01_n818 ), .A3(_AES_ENC_us01_n817 ), .A4(_AES_ENC_us01_n816 ), .ZN(_AES_ENC_us01_n820 ) );
NAND2_X2 _AES_ENC_us01_U248  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n820 ), .ZN(_AES_ENC_us01_n851 ) );
NAND2_X2 _AES_ENC_us01_U247  ( .A1(_AES_ENC_us01_n956 ), .A2(_AES_ENC_us01_n1080 ), .ZN(_AES_ENC_us01_n835 ) );
NAND2_X2 _AES_ENC_us01_U246  ( .A1(_AES_ENC_us01_n570 ), .A2(_AES_ENC_us01_n1030 ), .ZN(_AES_ENC_us01_n1047 ) );
OR2_X2 _AES_ENC_us01_U245  ( .A1(_AES_ENC_us01_n1047 ), .A2(_AES_ENC_us01_n582 ), .ZN(_AES_ENC_us01_n834 ) );
NAND2_X2 _AES_ENC_us01_U244  ( .A1(_AES_ENC_us01_n1072 ), .A2(_AES_ENC_us01_n620 ), .ZN(_AES_ENC_us01_n833 ) );
NAND4_X2 _AES_ENC_us01_U233  ( .A1(_AES_ENC_us01_n835 ), .A2(_AES_ENC_us01_n834 ), .A3(_AES_ENC_us01_n833 ), .A4(_AES_ENC_us01_n832 ), .ZN(_AES_ENC_us01_n836 ) );
NAND2_X2 _AES_ENC_us01_U232  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n836 ), .ZN(_AES_ENC_us01_n850 ) );
NAND2_X2 _AES_ENC_us01_U231  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n601 ), .ZN(_AES_ENC_us01_n847 ) );
NAND2_X2 _AES_ENC_us01_U230  ( .A1(_AES_ENC_us01_n1050 ), .A2(_AES_ENC_us01_n1071 ), .ZN(_AES_ENC_us01_n846 ) );
OR2_X2 _AES_ENC_us01_U224  ( .A1(_AES_ENC_us01_n1053 ), .A2(_AES_ENC_us01_n911 ), .ZN(_AES_ENC_us01_n1077 ) );
NAND4_X2 _AES_ENC_us01_U220  ( .A1(_AES_ENC_us01_n847 ), .A2(_AES_ENC_us01_n846 ), .A3(_AES_ENC_us01_n845 ), .A4(_AES_ENC_us01_n844 ), .ZN(_AES_ENC_us01_n848 ) );
NAND2_X2 _AES_ENC_us01_U219  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n848 ), .ZN(_AES_ENC_us01_n849 ) );
NAND4_X2 _AES_ENC_us01_U218  ( .A1(_AES_ENC_us01_n852 ), .A2(_AES_ENC_us01_n851 ), .A3(_AES_ENC_us01_n850 ), .A4(_AES_ENC_us01_n849 ), .ZN(_AES_ENC_sa01_sub[3] ) );
NAND2_X2 _AES_ENC_us01_U216  ( .A1(_AES_ENC_us01_n1009 ), .A2(_AES_ENC_us01_n1072 ), .ZN(_AES_ENC_us01_n862 ) );
NAND2_X2 _AES_ENC_us01_U215  ( .A1(_AES_ENC_us01_n610 ), .A2(_AES_ENC_us01_n618 ), .ZN(_AES_ENC_us01_n853 ) );
NAND2_X2 _AES_ENC_us01_U214  ( .A1(_AES_ENC_us01_n1050 ), .A2(_AES_ENC_us01_n853 ), .ZN(_AES_ENC_us01_n861 ) );
NAND4_X2 _AES_ENC_us01_U206  ( .A1(_AES_ENC_us01_n862 ), .A2(_AES_ENC_us01_n861 ), .A3(_AES_ENC_us01_n860 ), .A4(_AES_ENC_us01_n859 ), .ZN(_AES_ENC_us01_n863 ) );
NAND2_X2 _AES_ENC_us01_U205  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n863 ), .ZN(_AES_ENC_us01_n905 ) );
NAND2_X2 _AES_ENC_us01_U204  ( .A1(_AES_ENC_us01_n1010 ), .A2(_AES_ENC_us01_n989 ), .ZN(_AES_ENC_us01_n874 ) );
NAND2_X2 _AES_ENC_us01_U203  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n592 ), .ZN(_AES_ENC_us01_n864 ) );
NAND2_X2 _AES_ENC_us01_U202  ( .A1(_AES_ENC_us01_n929 ), .A2(_AES_ENC_us01_n864 ), .ZN(_AES_ENC_us01_n873 ) );
NAND4_X2 _AES_ENC_us01_U193  ( .A1(_AES_ENC_us01_n874 ), .A2(_AES_ENC_us01_n873 ), .A3(_AES_ENC_us01_n872 ), .A4(_AES_ENC_us01_n871 ), .ZN(_AES_ENC_us01_n875 ) );
NAND2_X2 _AES_ENC_us01_U192  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n875 ), .ZN(_AES_ENC_us01_n904 ) );
NAND2_X2 _AES_ENC_us01_U191  ( .A1(_AES_ENC_us01_n597 ), .A2(_AES_ENC_us01_n1050 ), .ZN(_AES_ENC_us01_n889 ) );
NAND2_X2 _AES_ENC_us01_U190  ( .A1(_AES_ENC_us01_n1093 ), .A2(_AES_ENC_us01_n617 ), .ZN(_AES_ENC_us01_n876 ) );
NAND2_X2 _AES_ENC_us01_U189  ( .A1(_AES_ENC_us01_n576 ), .A2(_AES_ENC_us01_n876 ), .ZN(_AES_ENC_us01_n877 ) );
NAND2_X2 _AES_ENC_us01_U188  ( .A1(_AES_ENC_us01_n877 ), .A2(_AES_ENC_us01_n601 ), .ZN(_AES_ENC_us01_n888 ) );
NAND4_X2 _AES_ENC_us01_U179  ( .A1(_AES_ENC_us01_n889 ), .A2(_AES_ENC_us01_n888 ), .A3(_AES_ENC_us01_n887 ), .A4(_AES_ENC_us01_n886 ), .ZN(_AES_ENC_us01_n890 ) );
NAND2_X2 _AES_ENC_us01_U178  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n890 ), .ZN(_AES_ENC_us01_n903 ) );
OR2_X2 _AES_ENC_us01_U177  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n1059 ), .ZN(_AES_ENC_us01_n900 ) );
NAND2_X2 _AES_ENC_us01_U176  ( .A1(_AES_ENC_us01_n1073 ), .A2(_AES_ENC_us01_n1047 ), .ZN(_AES_ENC_us01_n899 ) );
NAND2_X2 _AES_ENC_us01_U175  ( .A1(_AES_ENC_us01_n1094 ), .A2(_AES_ENC_us01_n608 ), .ZN(_AES_ENC_us01_n898 ) );
NAND4_X2 _AES_ENC_us01_U167  ( .A1(_AES_ENC_us01_n900 ), .A2(_AES_ENC_us01_n899 ), .A3(_AES_ENC_us01_n898 ), .A4(_AES_ENC_us01_n897 ), .ZN(_AES_ENC_us01_n901 ) );
NAND2_X2 _AES_ENC_us01_U166  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n901 ), .ZN(_AES_ENC_us01_n902 ) );
NAND4_X2 _AES_ENC_us01_U165  ( .A1(_AES_ENC_us01_n905 ), .A2(_AES_ENC_us01_n904 ), .A3(_AES_ENC_us01_n903 ), .A4(_AES_ENC_us01_n902 ), .ZN(_AES_ENC_sa01_sub[4] ) );
NAND2_X2 _AES_ENC_us01_U164  ( .A1(_AES_ENC_us01_n1094 ), .A2(_AES_ENC_us01_n615 ), .ZN(_AES_ENC_us01_n922 ) );
NAND2_X2 _AES_ENC_us01_U163  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n989 ), .ZN(_AES_ENC_us01_n921 ) );
NAND4_X2 _AES_ENC_us01_U151  ( .A1(_AES_ENC_us01_n922 ), .A2(_AES_ENC_us01_n921 ), .A3(_AES_ENC_us01_n920 ), .A4(_AES_ENC_us01_n919 ), .ZN(_AES_ENC_us01_n923 ) );
NAND2_X2 _AES_ENC_us01_U150  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n923 ), .ZN(_AES_ENC_us01_n972 ) );
NAND2_X2 _AES_ENC_us01_U149  ( .A1(_AES_ENC_us01_n603 ), .A2(_AES_ENC_us01_n605 ), .ZN(_AES_ENC_us01_n924 ) );
NAND2_X2 _AES_ENC_us01_U148  ( .A1(_AES_ENC_us01_n1073 ), .A2(_AES_ENC_us01_n924 ), .ZN(_AES_ENC_us01_n939 ) );
NAND2_X2 _AES_ENC_us01_U147  ( .A1(_AES_ENC_us01_n926 ), .A2(_AES_ENC_us01_n925 ), .ZN(_AES_ENC_us01_n927 ) );
NAND2_X2 _AES_ENC_us01_U146  ( .A1(_AES_ENC_us01_n587 ), .A2(_AES_ENC_us01_n927 ), .ZN(_AES_ENC_us01_n928 ) );
NAND2_X2 _AES_ENC_us01_U145  ( .A1(_AES_ENC_us01_n928 ), .A2(_AES_ENC_us01_n1080 ), .ZN(_AES_ENC_us01_n938 ) );
OR2_X2 _AES_ENC_us01_U144  ( .A1(_AES_ENC_us01_n1117 ), .A2(_AES_ENC_us01_n580 ), .ZN(_AES_ENC_us01_n937 ) );
NAND4_X2 _AES_ENC_us01_U139  ( .A1(_AES_ENC_us01_n939 ), .A2(_AES_ENC_us01_n938 ), .A3(_AES_ENC_us01_n937 ), .A4(_AES_ENC_us01_n936 ), .ZN(_AES_ENC_us01_n940 ) );
NAND2_X2 _AES_ENC_us01_U138  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n940 ), .ZN(_AES_ENC_us01_n971 ) );
OR2_X2 _AES_ENC_us01_U137  ( .A1(_AES_ENC_us01_n586 ), .A2(_AES_ENC_us01_n941 ), .ZN(_AES_ENC_us01_n954 ) );
NAND2_X2 _AES_ENC_us01_U136  ( .A1(_AES_ENC_us01_n1096 ), .A2(_AES_ENC_us01_n618 ), .ZN(_AES_ENC_us01_n942 ) );
NAND2_X2 _AES_ENC_us01_U135  ( .A1(_AES_ENC_us01_n1048 ), .A2(_AES_ENC_us01_n942 ), .ZN(_AES_ENC_us01_n943 ) );
NAND2_X2 _AES_ENC_us01_U134  ( .A1(_AES_ENC_us01_n582 ), .A2(_AES_ENC_us01_n943 ), .ZN(_AES_ENC_us01_n944 ) );
NAND2_X2 _AES_ENC_us01_U133  ( .A1(_AES_ENC_us01_n944 ), .A2(_AES_ENC_us01_n599 ), .ZN(_AES_ENC_us01_n953 ) );
NAND4_X2 _AES_ENC_us01_U125  ( .A1(_AES_ENC_us01_n954 ), .A2(_AES_ENC_us01_n953 ), .A3(_AES_ENC_us01_n952 ), .A4(_AES_ENC_us01_n951 ), .ZN(_AES_ENC_us01_n955 ) );
NAND2_X2 _AES_ENC_us01_U124  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n955 ), .ZN(_AES_ENC_us01_n970 ) );
NAND2_X2 _AES_ENC_us01_U123  ( .A1(_AES_ENC_us01_n1094 ), .A2(_AES_ENC_us01_n1071 ), .ZN(_AES_ENC_us01_n967 ) );
NAND2_X2 _AES_ENC_us01_U122  ( .A1(_AES_ENC_us01_n956 ), .A2(_AES_ENC_us01_n1030 ), .ZN(_AES_ENC_us01_n966 ) );
NAND4_X2 _AES_ENC_us01_U114  ( .A1(_AES_ENC_us01_n967 ), .A2(_AES_ENC_us01_n966 ), .A3(_AES_ENC_us01_n965 ), .A4(_AES_ENC_us01_n964 ), .ZN(_AES_ENC_us01_n968 ) );
NAND2_X2 _AES_ENC_us01_U113  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n968 ), .ZN(_AES_ENC_us01_n969 ) );
NAND4_X2 _AES_ENC_us01_U112  ( .A1(_AES_ENC_us01_n972 ), .A2(_AES_ENC_us01_n971 ), .A3(_AES_ENC_us01_n970 ), .A4(_AES_ENC_us01_n969 ), .ZN(_AES_ENC_sa01_sub[5] ) );
NAND2_X2 _AES_ENC_us01_U111  ( .A1(_AES_ENC_us01_n570 ), .A2(_AES_ENC_us01_n1097 ), .ZN(_AES_ENC_us01_n973 ) );
NAND2_X2 _AES_ENC_us01_U110  ( .A1(_AES_ENC_us01_n1073 ), .A2(_AES_ENC_us01_n973 ), .ZN(_AES_ENC_us01_n987 ) );
NAND2_X2 _AES_ENC_us01_U109  ( .A1(_AES_ENC_us01_n974 ), .A2(_AES_ENC_us01_n1077 ), .ZN(_AES_ENC_us01_n975 ) );
NAND2_X2 _AES_ENC_us01_U108  ( .A1(_AES_ENC_us01_n584 ), .A2(_AES_ENC_us01_n975 ), .ZN(_AES_ENC_us01_n976 ) );
NAND2_X2 _AES_ENC_us01_U107  ( .A1(_AES_ENC_us01_n977 ), .A2(_AES_ENC_us01_n976 ), .ZN(_AES_ENC_us01_n986 ) );
NAND4_X2 _AES_ENC_us01_U99  ( .A1(_AES_ENC_us01_n987 ), .A2(_AES_ENC_us01_n986 ), .A3(_AES_ENC_us01_n985 ), .A4(_AES_ENC_us01_n984 ), .ZN(_AES_ENC_us01_n988 ) );
NAND2_X2 _AES_ENC_us01_U98  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n988 ), .ZN(_AES_ENC_us01_n1044 ) );
NAND2_X2 _AES_ENC_us01_U97  ( .A1(_AES_ENC_us01_n1073 ), .A2(_AES_ENC_us01_n989 ), .ZN(_AES_ENC_us01_n1004 ) );
NAND2_X2 _AES_ENC_us01_U96  ( .A1(_AES_ENC_us01_n1092 ), .A2(_AES_ENC_us01_n605 ), .ZN(_AES_ENC_us01_n1003 ) );
NAND4_X2 _AES_ENC_us01_U85  ( .A1(_AES_ENC_us01_n1004 ), .A2(_AES_ENC_us01_n1003 ), .A3(_AES_ENC_us01_n1002 ), .A4(_AES_ENC_us01_n1001 ), .ZN(_AES_ENC_us01_n1005 ) );
NAND2_X2 _AES_ENC_us01_U84  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n1005 ), .ZN(_AES_ENC_us01_n1043 ) );
NAND2_X2 _AES_ENC_us01_U83  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n626 ), .ZN(_AES_ENC_us01_n1020 ) );
NAND2_X2 _AES_ENC_us01_U82  ( .A1(_AES_ENC_us01_n1050 ), .A2(_AES_ENC_us01_n612 ), .ZN(_AES_ENC_us01_n1019 ) );
NAND2_X2 _AES_ENC_us01_U77  ( .A1(_AES_ENC_us01_n1059 ), .A2(_AES_ENC_us01_n1114 ), .ZN(_AES_ENC_us01_n1012 ) );
NAND2_X2 _AES_ENC_us01_U76  ( .A1(_AES_ENC_us01_n1010 ), .A2(_AES_ENC_us01_n604 ), .ZN(_AES_ENC_us01_n1011 ) );
NAND2_X2 _AES_ENC_us01_U75  ( .A1(_AES_ENC_us01_n1012 ), .A2(_AES_ENC_us01_n1011 ), .ZN(_AES_ENC_us01_n1016 ) );
NAND4_X2 _AES_ENC_us01_U70  ( .A1(_AES_ENC_us01_n1020 ), .A2(_AES_ENC_us01_n1019 ), .A3(_AES_ENC_us01_n1018 ), .A4(_AES_ENC_us01_n1017 ), .ZN(_AES_ENC_us01_n1021 ) );
NAND2_X2 _AES_ENC_us01_U69  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n1021 ), .ZN(_AES_ENC_us01_n1042 ) );
NAND2_X2 _AES_ENC_us01_U68  ( .A1(_AES_ENC_us01_n1022 ), .A2(_AES_ENC_us01_n1093 ), .ZN(_AES_ENC_us01_n1039 ) );
NAND2_X2 _AES_ENC_us01_U67  ( .A1(_AES_ENC_us01_n1050 ), .A2(_AES_ENC_us01_n1023 ), .ZN(_AES_ENC_us01_n1038 ) );
NAND2_X2 _AES_ENC_us01_U66  ( .A1(_AES_ENC_us01_n1024 ), .A2(_AES_ENC_us01_n1071 ), .ZN(_AES_ENC_us01_n1037 ) );
AND2_X2 _AES_ENC_us01_U60  ( .A1(_AES_ENC_us01_n1030 ), .A2(_AES_ENC_us01_n621 ), .ZN(_AES_ENC_us01_n1078 ) );
NAND4_X2 _AES_ENC_us01_U56  ( .A1(_AES_ENC_us01_n1039 ), .A2(_AES_ENC_us01_n1038 ), .A3(_AES_ENC_us01_n1037 ), .A4(_AES_ENC_us01_n1036 ), .ZN(_AES_ENC_us01_n1040 ) );
NAND2_X2 _AES_ENC_us01_U55  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n1040 ), .ZN(_AES_ENC_us01_n1041 ) );
NAND4_X2 _AES_ENC_us01_U54  ( .A1(_AES_ENC_us01_n1044 ), .A2(_AES_ENC_us01_n1043 ), .A3(_AES_ENC_us01_n1042 ), .A4(_AES_ENC_us01_n1041 ), .ZN(_AES_ENC_sa01_sub[6] ) );
NAND2_X2 _AES_ENC_us01_U53  ( .A1(_AES_ENC_us01_n1072 ), .A2(_AES_ENC_us01_n1045 ), .ZN(_AES_ENC_us01_n1068 ) );
NAND2_X2 _AES_ENC_us01_U52  ( .A1(_AES_ENC_us01_n1046 ), .A2(_AES_ENC_us01_n603 ), .ZN(_AES_ENC_us01_n1067 ) );
NAND2_X2 _AES_ENC_us01_U51  ( .A1(_AES_ENC_us01_n1094 ), .A2(_AES_ENC_us01_n1047 ), .ZN(_AES_ENC_us01_n1066 ) );
NAND4_X2 _AES_ENC_us01_U40  ( .A1(_AES_ENC_us01_n1068 ), .A2(_AES_ENC_us01_n1067 ), .A3(_AES_ENC_us01_n1066 ), .A4(_AES_ENC_us01_n1065 ), .ZN(_AES_ENC_us01_n1069 ) );
NAND2_X2 _AES_ENC_us01_U39  ( .A1(_AES_ENC_us01_n1070 ), .A2(_AES_ENC_us01_n1069 ), .ZN(_AES_ENC_us01_n1135 ) );
NAND2_X2 _AES_ENC_us01_U38  ( .A1(_AES_ENC_us01_n1072 ), .A2(_AES_ENC_us01_n1071 ), .ZN(_AES_ENC_us01_n1088 ) );
NAND2_X2 _AES_ENC_us01_U37  ( .A1(_AES_ENC_us01_n1073 ), .A2(_AES_ENC_us01_n608 ), .ZN(_AES_ENC_us01_n1087 ) );
NAND4_X2 _AES_ENC_us01_U28  ( .A1(_AES_ENC_us01_n1088 ), .A2(_AES_ENC_us01_n1087 ), .A3(_AES_ENC_us01_n1086 ), .A4(_AES_ENC_us01_n1085 ), .ZN(_AES_ENC_us01_n1089 ) );
NAND2_X2 _AES_ENC_us01_U27  ( .A1(_AES_ENC_us01_n1090 ), .A2(_AES_ENC_us01_n1089 ), .ZN(_AES_ENC_us01_n1134 ) );
NAND2_X2 _AES_ENC_us01_U26  ( .A1(_AES_ENC_us01_n1091 ), .A2(_AES_ENC_us01_n1093 ), .ZN(_AES_ENC_us01_n1111 ) );
NAND2_X2 _AES_ENC_us01_U25  ( .A1(_AES_ENC_us01_n1092 ), .A2(_AES_ENC_us01_n1120 ), .ZN(_AES_ENC_us01_n1110 ) );
AND2_X2 _AES_ENC_us01_U22  ( .A1(_AES_ENC_us01_n1097 ), .A2(_AES_ENC_us01_n1096 ), .ZN(_AES_ENC_us01_n1098 ) );
NAND4_X2 _AES_ENC_us01_U14  ( .A1(_AES_ENC_us01_n1111 ), .A2(_AES_ENC_us01_n1110 ), .A3(_AES_ENC_us01_n1109 ), .A4(_AES_ENC_us01_n1108 ), .ZN(_AES_ENC_us01_n1112 ) );
NAND2_X2 _AES_ENC_us01_U13  ( .A1(_AES_ENC_us01_n1113 ), .A2(_AES_ENC_us01_n1112 ), .ZN(_AES_ENC_us01_n1133 ) );
NAND2_X2 _AES_ENC_us01_U12  ( .A1(_AES_ENC_us01_n1115 ), .A2(_AES_ENC_us01_n1114 ), .ZN(_AES_ENC_us01_n1129 ) );
OR2_X2 _AES_ENC_us01_U11  ( .A1(_AES_ENC_us01_n579 ), .A2(_AES_ENC_us01_n1116 ), .ZN(_AES_ENC_us01_n1128 ) );
NAND4_X2 _AES_ENC_us01_U3  ( .A1(_AES_ENC_us01_n1129 ), .A2(_AES_ENC_us01_n1128 ), .A3(_AES_ENC_us01_n1127 ), .A4(_AES_ENC_us01_n1126 ), .ZN(_AES_ENC_us01_n1130 ) );
NAND2_X2 _AES_ENC_us01_U2  ( .A1(_AES_ENC_us01_n1131 ), .A2(_AES_ENC_us01_n1130 ), .ZN(_AES_ENC_us01_n1132 ) );
NAND4_X2 _AES_ENC_us01_U1  ( .A1(_AES_ENC_us01_n1135 ), .A2(_AES_ENC_us01_n1134 ), .A3(_AES_ENC_us01_n1133 ), .A4(_AES_ENC_us01_n1132 ), .ZN(_AES_ENC_sa01_sub[7] ) );
INV_X4 _AES_ENC_us02_U575  ( .A(_AES_ENC_sa02[7]), .ZN(_AES_ENC_us02_n627 ));
INV_X4 _AES_ENC_us02_U574  ( .A(_AES_ENC_us02_n1114 ), .ZN(_AES_ENC_us02_n625 ) );
INV_X4 _AES_ENC_us02_U573  ( .A(_AES_ENC_sa02[4]), .ZN(_AES_ENC_us02_n624 ));
INV_X4 _AES_ENC_us02_U572  ( .A(_AES_ENC_us02_n1025 ), .ZN(_AES_ENC_us02_n622 ) );
INV_X4 _AES_ENC_us02_U571  ( .A(_AES_ENC_us02_n1120 ), .ZN(_AES_ENC_us02_n620 ) );
INV_X4 _AES_ENC_us02_U570  ( .A(_AES_ENC_us02_n1121 ), .ZN(_AES_ENC_us02_n619 ) );
INV_X4 _AES_ENC_us02_U569  ( .A(_AES_ENC_us02_n1048 ), .ZN(_AES_ENC_us02_n618 ) );
INV_X4 _AES_ENC_us02_U568  ( .A(_AES_ENC_us02_n974 ), .ZN(_AES_ENC_us02_n616 ) );
INV_X4 _AES_ENC_us02_U567  ( .A(_AES_ENC_us02_n794 ), .ZN(_AES_ENC_us02_n614 ) );
INV_X4 _AES_ENC_us02_U566  ( .A(_AES_ENC_sa02[2]), .ZN(_AES_ENC_us02_n611 ));
INV_X4 _AES_ENC_us02_U565  ( .A(_AES_ENC_us02_n800 ), .ZN(_AES_ENC_us02_n610 ) );
INV_X4 _AES_ENC_us02_U564  ( .A(_AES_ENC_us02_n925 ), .ZN(_AES_ENC_us02_n609 ) );
INV_X4 _AES_ENC_us02_U563  ( .A(_AES_ENC_us02_n779 ), .ZN(_AES_ENC_us02_n607 ) );
INV_X4 _AES_ENC_us02_U562  ( .A(_AES_ENC_us02_n1022 ), .ZN(_AES_ENC_us02_n603 ) );
INV_X4 _AES_ENC_us02_U561  ( .A(_AES_ENC_us02_n1102 ), .ZN(_AES_ENC_us02_n602 ) );
INV_X4 _AES_ENC_us02_U560  ( .A(_AES_ENC_us02_n929 ), .ZN(_AES_ENC_us02_n601 ) );
INV_X4 _AES_ENC_us02_U559  ( .A(_AES_ENC_us02_n1056 ), .ZN(_AES_ENC_us02_n600 ) );
INV_X4 _AES_ENC_us02_U558  ( .A(_AES_ENC_us02_n1054 ), .ZN(_AES_ENC_us02_n599 ) );
INV_X4 _AES_ENC_us02_U557  ( .A(_AES_ENC_us02_n881 ), .ZN(_AES_ENC_us02_n598 ) );
INV_X4 _AES_ENC_us02_U556  ( .A(_AES_ENC_us02_n926 ), .ZN(_AES_ENC_us02_n597 ) );
INV_X4 _AES_ENC_us02_U555  ( .A(_AES_ENC_us02_n977 ), .ZN(_AES_ENC_us02_n595 ) );
INV_X4 _AES_ENC_us02_U554  ( .A(_AES_ENC_us02_n1031 ), .ZN(_AES_ENC_us02_n594 ) );
INV_X4 _AES_ENC_us02_U553  ( .A(_AES_ENC_us02_n1103 ), .ZN(_AES_ENC_us02_n593 ) );
INV_X4 _AES_ENC_us02_U552  ( .A(_AES_ENC_us02_n1009 ), .ZN(_AES_ENC_us02_n592 ) );
INV_X4 _AES_ENC_us02_U551  ( .A(_AES_ENC_us02_n990 ), .ZN(_AES_ENC_us02_n591 ) );
INV_X4 _AES_ENC_us02_U550  ( .A(_AES_ENC_us02_n1058 ), .ZN(_AES_ENC_us02_n590 ) );
INV_X4 _AES_ENC_us02_U549  ( .A(_AES_ENC_us02_n1074 ), .ZN(_AES_ENC_us02_n589 ) );
INV_X4 _AES_ENC_us02_U548  ( .A(_AES_ENC_us02_n1053 ), .ZN(_AES_ENC_us02_n588 ) );
INV_X4 _AES_ENC_us02_U547  ( .A(_AES_ENC_us02_n826 ), .ZN(_AES_ENC_us02_n587 ) );
INV_X4 _AES_ENC_us02_U546  ( .A(_AES_ENC_us02_n992 ), .ZN(_AES_ENC_us02_n586 ) );
INV_X4 _AES_ENC_us02_U545  ( .A(_AES_ENC_us02_n821 ), .ZN(_AES_ENC_us02_n585 ) );
INV_X4 _AES_ENC_us02_U544  ( .A(_AES_ENC_us02_n910 ), .ZN(_AES_ENC_us02_n584 ) );
INV_X4 _AES_ENC_us02_U543  ( .A(_AES_ENC_us02_n906 ), .ZN(_AES_ENC_us02_n583 ) );
INV_X4 _AES_ENC_us02_U542  ( .A(_AES_ENC_us02_n880 ), .ZN(_AES_ENC_us02_n581 ) );
INV_X4 _AES_ENC_us02_U541  ( .A(_AES_ENC_us02_n1013 ), .ZN(_AES_ENC_us02_n580 ) );
INV_X4 _AES_ENC_us02_U540  ( .A(_AES_ENC_us02_n1092 ), .ZN(_AES_ENC_us02_n579 ) );
INV_X4 _AES_ENC_us02_U539  ( .A(_AES_ENC_us02_n824 ), .ZN(_AES_ENC_us02_n578 ) );
INV_X4 _AES_ENC_us02_U538  ( .A(_AES_ENC_us02_n1091 ), .ZN(_AES_ENC_us02_n577 ) );
INV_X4 _AES_ENC_us02_U537  ( .A(_AES_ENC_us02_n1080 ), .ZN(_AES_ENC_us02_n576 ) );
INV_X4 _AES_ENC_us02_U536  ( .A(_AES_ENC_us02_n959 ), .ZN(_AES_ENC_us02_n575 ) );
INV_X4 _AES_ENC_us02_U535  ( .A(_AES_ENC_sa02[0]), .ZN(_AES_ENC_us02_n574 ));
NOR2_X2 _AES_ENC_us02_U534  ( .A1(_AES_ENC_sa02[0]), .A2(_AES_ENC_sa02[6]),.ZN(_AES_ENC_us02_n1090 ) );
NOR2_X2 _AES_ENC_us02_U533  ( .A1(_AES_ENC_us02_n574 ), .A2(_AES_ENC_sa02[6]), .ZN(_AES_ENC_us02_n1070 ) );
NOR2_X2 _AES_ENC_us02_U532  ( .A1(_AES_ENC_sa02[4]), .A2(_AES_ENC_sa02[3]),.ZN(_AES_ENC_us02_n1025 ) );
INV_X4 _AES_ENC_us02_U531  ( .A(_AES_ENC_us02_n569 ), .ZN(_AES_ENC_us02_n572 ) );
NOR2_X2 _AES_ENC_us02_U530  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n765 ) );
NOR2_X2 _AES_ENC_us02_U529  ( .A1(_AES_ENC_sa02[4]), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n764 ) );
NOR2_X2 _AES_ENC_us02_U528  ( .A1(_AES_ENC_us02_n765 ), .A2(_AES_ENC_us02_n764 ), .ZN(_AES_ENC_us02_n766 ) );
NOR2_X2 _AES_ENC_us02_U527  ( .A1(_AES_ENC_us02_n766 ), .A2(_AES_ENC_us02_n575 ), .ZN(_AES_ENC_us02_n767 ) );
NOR3_X2 _AES_ENC_us02_U526  ( .A1(_AES_ENC_us02_n627 ), .A2(_AES_ENC_sa02[5]), .A3(_AES_ENC_us02_n704 ), .ZN(_AES_ENC_us02_n706 ));
NOR2_X2 _AES_ENC_us02_U525  ( .A1(_AES_ENC_us02_n1117 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n707 ) );
NOR2_X2 _AES_ENC_us02_U524  ( .A1(_AES_ENC_sa02[4]), .A2(_AES_ENC_us02_n579 ), .ZN(_AES_ENC_us02_n705 ) );
NOR3_X2 _AES_ENC_us02_U523  ( .A1(_AES_ENC_us02_n707 ), .A2(_AES_ENC_us02_n706 ), .A3(_AES_ENC_us02_n705 ), .ZN(_AES_ENC_us02_n713 ) );
INV_X4 _AES_ENC_us02_U522  ( .A(_AES_ENC_sa02[3]), .ZN(_AES_ENC_us02_n621 ));
NAND3_X2 _AES_ENC_us02_U521  ( .A1(_AES_ENC_us02_n652 ), .A2(_AES_ENC_us02_n626 ), .A3(_AES_ENC_sa02[7]), .ZN(_AES_ENC_us02_n653 ));
NOR2_X2 _AES_ENC_us02_U520  ( .A1(_AES_ENC_us02_n611 ), .A2(_AES_ENC_sa02[5]), .ZN(_AES_ENC_us02_n925 ) );
NOR2_X2 _AES_ENC_us02_U519  ( .A1(_AES_ENC_sa02[5]), .A2(_AES_ENC_sa02[2]),.ZN(_AES_ENC_us02_n974 ) );
INV_X4 _AES_ENC_us02_U518  ( .A(_AES_ENC_sa02[5]), .ZN(_AES_ENC_us02_n626 ));
NOR2_X2 _AES_ENC_us02_U517  ( .A1(_AES_ENC_us02_n611 ), .A2(_AES_ENC_sa02[7]), .ZN(_AES_ENC_us02_n779 ) );
NAND3_X2 _AES_ENC_us02_U516  ( .A1(_AES_ENC_us02_n679 ), .A2(_AES_ENC_us02_n678 ), .A3(_AES_ENC_us02_n677 ), .ZN(_AES_ENC_sa02_sub[0] ) );
NOR2_X2 _AES_ENC_us02_U515  ( .A1(_AES_ENC_us02_n626 ), .A2(_AES_ENC_sa02[2]), .ZN(_AES_ENC_us02_n1048 ) );
NOR4_X2 _AES_ENC_us02_U512  ( .A1(_AES_ENC_us02_n633 ), .A2(_AES_ENC_us02_n632 ), .A3(_AES_ENC_us02_n631 ), .A4(_AES_ENC_us02_n630 ), .ZN(_AES_ENC_us02_n634 ) );
NOR2_X2 _AES_ENC_us02_U510  ( .A1(_AES_ENC_us02_n629 ), .A2(_AES_ENC_us02_n628 ), .ZN(_AES_ENC_us02_n635 ) );
NAND3_X2 _AES_ENC_us02_U509  ( .A1(_AES_ENC_sa02[2]), .A2(_AES_ENC_sa02[7]), .A3(_AES_ENC_us02_n1059 ), .ZN(_AES_ENC_us02_n636 ) );
NOR2_X2 _AES_ENC_us02_U508  ( .A1(_AES_ENC_sa02[7]), .A2(_AES_ENC_sa02[2]),.ZN(_AES_ENC_us02_n794 ) );
NOR2_X2 _AES_ENC_us02_U507  ( .A1(_AES_ENC_sa02[4]), .A2(_AES_ENC_sa02[1]),.ZN(_AES_ENC_us02_n1102 ) );
NOR2_X2 _AES_ENC_us02_U506  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_sa02[3]), .ZN(_AES_ENC_us02_n1053 ) );
NOR2_X2 _AES_ENC_us02_U505  ( .A1(_AES_ENC_us02_n607 ), .A2(_AES_ENC_sa02[5]), .ZN(_AES_ENC_us02_n1024 ) );
NOR2_X2 _AES_ENC_us02_U504  ( .A1(_AES_ENC_us02_n625 ), .A2(_AES_ENC_sa02[2]), .ZN(_AES_ENC_us02_n1093 ) );
NOR2_X2 _AES_ENC_us02_U503  ( .A1(_AES_ENC_us02_n614 ), .A2(_AES_ENC_sa02[5]), .ZN(_AES_ENC_us02_n1094 ) );
NOR2_X2 _AES_ENC_us02_U502  ( .A1(_AES_ENC_us02_n624 ), .A2(_AES_ENC_sa02[3]), .ZN(_AES_ENC_us02_n931 ) );
INV_X4 _AES_ENC_us02_U501  ( .A(_AES_ENC_us02_n570 ), .ZN(_AES_ENC_us02_n573 ) );
NOR2_X2 _AES_ENC_us02_U500  ( .A1(_AES_ENC_us02_n1053 ), .A2(_AES_ENC_us02_n1095 ), .ZN(_AES_ENC_us02_n639 ) );
NOR3_X2 _AES_ENC_us02_U499  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n573 ), .A3(_AES_ENC_us02_n1074 ), .ZN(_AES_ENC_us02_n641 ) );
NOR2_X2 _AES_ENC_us02_U498  ( .A1(_AES_ENC_us02_n639 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n640 ) );
NOR2_X2 _AES_ENC_us02_U497  ( .A1(_AES_ENC_us02_n641 ), .A2(_AES_ENC_us02_n640 ), .ZN(_AES_ENC_us02_n646 ) );
NOR3_X2 _AES_ENC_us02_U496  ( .A1(_AES_ENC_us02_n995 ), .A2(_AES_ENC_us02_n586 ), .A3(_AES_ENC_us02_n994 ), .ZN(_AES_ENC_us02_n1002 ) );
NOR2_X2 _AES_ENC_us02_U495  ( .A1(_AES_ENC_us02_n909 ), .A2(_AES_ENC_us02_n908 ), .ZN(_AES_ENC_us02_n920 ) );
NOR2_X2 _AES_ENC_us02_U494  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n823 ) );
NOR2_X2 _AES_ENC_us02_U492  ( .A1(_AES_ENC_us02_n624 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n822 ) );
NOR2_X2 _AES_ENC_us02_U491  ( .A1(_AES_ENC_us02_n823 ), .A2(_AES_ENC_us02_n822 ), .ZN(_AES_ENC_us02_n825 ) );
NOR2_X2 _AES_ENC_us02_U490  ( .A1(_AES_ENC_sa02[1]), .A2(_AES_ENC_us02_n623 ), .ZN(_AES_ENC_us02_n913 ) );
NOR2_X2 _AES_ENC_us02_U489  ( .A1(_AES_ENC_us02_n913 ), .A2(_AES_ENC_us02_n1091 ), .ZN(_AES_ENC_us02_n914 ) );
NOR2_X2 _AES_ENC_us02_U488  ( .A1(_AES_ENC_us02_n826 ), .A2(_AES_ENC_us02_n572 ), .ZN(_AES_ENC_us02_n827 ) );
NOR3_X2 _AES_ENC_us02_U487  ( .A1(_AES_ENC_us02_n769 ), .A2(_AES_ENC_us02_n768 ), .A3(_AES_ENC_us02_n767 ), .ZN(_AES_ENC_us02_n775 ) );
NOR2_X2 _AES_ENC_us02_U486  ( .A1(_AES_ENC_us02_n1056 ), .A2(_AES_ENC_us02_n1053 ), .ZN(_AES_ENC_us02_n749 ) );
NOR2_X2 _AES_ENC_us02_U483  ( .A1(_AES_ENC_us02_n749 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n752 ) );
INV_X4 _AES_ENC_us02_U482  ( .A(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n596 ));
NOR2_X2 _AES_ENC_us02_U480  ( .A1(_AES_ENC_us02_n1054 ), .A2(_AES_ENC_us02_n1053 ), .ZN(_AES_ENC_us02_n1055 ) );
OR2_X4 _AES_ENC_us02_U479  ( .A1(_AES_ENC_us02_n1094 ), .A2(_AES_ENC_us02_n1093 ), .ZN(_AES_ENC_us02_n571 ) );
AND2_X2 _AES_ENC_us02_U478  ( .A1(_AES_ENC_us02_n571 ), .A2(_AES_ENC_us02_n1095 ), .ZN(_AES_ENC_us02_n1101 ) );
NOR2_X2 _AES_ENC_us02_U477  ( .A1(_AES_ENC_us02_n1074 ), .A2(_AES_ENC_us02_n931 ), .ZN(_AES_ENC_us02_n796 ) );
NOR2_X2 _AES_ENC_us02_U474  ( .A1(_AES_ENC_us02_n796 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n797 ) );
NOR2_X2 _AES_ENC_us02_U473  ( .A1(_AES_ENC_us02_n932 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n933 ) );
NOR2_X2 _AES_ENC_us02_U472  ( .A1(_AES_ENC_us02_n929 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n935 ) );
NOR2_X2 _AES_ENC_us02_U471  ( .A1(_AES_ENC_us02_n931 ), .A2(_AES_ENC_us02_n930 ), .ZN(_AES_ENC_us02_n934 ) );
NOR3_X2 _AES_ENC_us02_U470  ( .A1(_AES_ENC_us02_n935 ), .A2(_AES_ENC_us02_n934 ), .A3(_AES_ENC_us02_n933 ), .ZN(_AES_ENC_us02_n936 ) );
NOR2_X2 _AES_ENC_us02_U469  ( .A1(_AES_ENC_us02_n624 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n1075 ) );
NOR2_X2 _AES_ENC_us02_U468  ( .A1(_AES_ENC_us02_n572 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n949 ) );
NOR2_X2 _AES_ENC_us02_U467  ( .A1(_AES_ENC_us02_n1049 ), .A2(_AES_ENC_us02_n618 ), .ZN(_AES_ENC_us02_n1051 ) );
NOR2_X2 _AES_ENC_us02_U466  ( .A1(_AES_ENC_us02_n1051 ), .A2(_AES_ENC_us02_n1050 ), .ZN(_AES_ENC_us02_n1052 ) );
NOR2_X2 _AES_ENC_us02_U465  ( .A1(_AES_ENC_us02_n1052 ), .A2(_AES_ENC_us02_n592 ), .ZN(_AES_ENC_us02_n1064 ) );
NOR2_X2 _AES_ENC_us02_U464  ( .A1(_AES_ENC_sa02[1]), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n631 ) );
NOR2_X2 _AES_ENC_us02_U463  ( .A1(_AES_ENC_us02_n1025 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n980 ) );
NOR2_X2 _AES_ENC_us02_U462  ( .A1(_AES_ENC_us02_n1073 ), .A2(_AES_ENC_us02_n1094 ), .ZN(_AES_ENC_us02_n795 ) );
NOR2_X2 _AES_ENC_us02_U461  ( .A1(_AES_ENC_us02_n795 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n799 ) );
NOR2_X2 _AES_ENC_us02_U460  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n981 ) );
NOR2_X2 _AES_ENC_us02_U459  ( .A1(_AES_ENC_us02_n1102 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n643 ) );
NOR2_X2 _AES_ENC_us02_U458  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n621 ), .ZN(_AES_ENC_us02_n642 ) );
NOR2_X2 _AES_ENC_us02_U455  ( .A1(_AES_ENC_us02_n911 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n644 ) );
NOR4_X2 _AES_ENC_us02_U448  ( .A1(_AES_ENC_us02_n644 ), .A2(_AES_ENC_us02_n643 ), .A3(_AES_ENC_us02_n804 ), .A4(_AES_ENC_us02_n642 ), .ZN(_AES_ENC_us02_n645 ) );
NOR2_X2 _AES_ENC_us02_U447  ( .A1(_AES_ENC_us02_n1102 ), .A2(_AES_ENC_us02_n910 ), .ZN(_AES_ENC_us02_n932 ) );
NOR2_X2 _AES_ENC_us02_U442  ( .A1(_AES_ENC_us02_n1102 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n755 ) );
NOR2_X2 _AES_ENC_us02_U441  ( .A1(_AES_ENC_us02_n931 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n743 ) );
NOR2_X2 _AES_ENC_us02_U438  ( .A1(_AES_ENC_us02_n1072 ), .A2(_AES_ENC_us02_n1094 ), .ZN(_AES_ENC_us02_n930 ) );
NOR2_X2 _AES_ENC_us02_U435  ( .A1(_AES_ENC_us02_n1074 ), .A2(_AES_ENC_us02_n1025 ), .ZN(_AES_ENC_us02_n891 ) );
NOR2_X2 _AES_ENC_us02_U434  ( .A1(_AES_ENC_us02_n891 ), .A2(_AES_ENC_us02_n609 ), .ZN(_AES_ENC_us02_n894 ) );
NOR3_X2 _AES_ENC_us02_U433  ( .A1(_AES_ENC_us02_n623 ), .A2(_AES_ENC_sa02[1]), .A3(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n683 ));
INV_X4 _AES_ENC_us02_U428  ( .A(_AES_ENC_us02_n931 ), .ZN(_AES_ENC_us02_n623 ) );
NOR2_X2 _AES_ENC_us02_U427  ( .A1(_AES_ENC_us02_n996 ), .A2(_AES_ENC_us02_n931 ), .ZN(_AES_ENC_us02_n704 ) );
NOR2_X2 _AES_ENC_us02_U421  ( .A1(_AES_ENC_us02_n931 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n685 ) );
NOR2_X2 _AES_ENC_us02_U420  ( .A1(_AES_ENC_us02_n1029 ), .A2(_AES_ENC_us02_n1025 ), .ZN(_AES_ENC_us02_n1079 ) );
NOR3_X2 _AES_ENC_us02_U419  ( .A1(_AES_ENC_us02_n589 ), .A2(_AES_ENC_us02_n1025 ), .A3(_AES_ENC_us02_n616 ), .ZN(_AES_ENC_us02_n945 ) );
NOR2_X2 _AES_ENC_us02_U418  ( .A1(_AES_ENC_us02_n626 ), .A2(_AES_ENC_us02_n611 ), .ZN(_AES_ENC_us02_n800 ) );
NOR3_X2 _AES_ENC_us02_U417  ( .A1(_AES_ENC_us02_n590 ), .A2(_AES_ENC_us02_n627 ), .A3(_AES_ENC_us02_n611 ), .ZN(_AES_ENC_us02_n798 ) );
NOR3_X2 _AES_ENC_us02_U416  ( .A1(_AES_ENC_us02_n610 ), .A2(_AES_ENC_us02_n572 ), .A3(_AES_ENC_us02_n575 ), .ZN(_AES_ENC_us02_n962 ) );
NOR3_X2 _AES_ENC_us02_U415  ( .A1(_AES_ENC_us02_n959 ), .A2(_AES_ENC_us02_n572 ), .A3(_AES_ENC_us02_n609 ), .ZN(_AES_ENC_us02_n768 ) );
NOR3_X2 _AES_ENC_us02_U414  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n572 ), .A3(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n694 ) );
NOR3_X2 _AES_ENC_us02_U413  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n572 ), .A3(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n895 ) );
NOR3_X2 _AES_ENC_us02_U410  ( .A1(_AES_ENC_us02_n1008 ), .A2(_AES_ENC_us02_n1007 ), .A3(_AES_ENC_us02_n1006 ), .ZN(_AES_ENC_us02_n1018 ) );
NOR4_X2 _AES_ENC_us02_U409  ( .A1(_AES_ENC_us02_n711 ), .A2(_AES_ENC_us02_n710 ), .A3(_AES_ENC_us02_n709 ), .A4(_AES_ENC_us02_n708 ), .ZN(_AES_ENC_us02_n712 ) );
NOR4_X2 _AES_ENC_us02_U406  ( .A1(_AES_ENC_us02_n806 ), .A2(_AES_ENC_us02_n805 ), .A3(_AES_ENC_us02_n804 ), .A4(_AES_ENC_us02_n803 ), .ZN(_AES_ENC_us02_n807 ) );
NOR3_X2 _AES_ENC_us02_U405  ( .A1(_AES_ENC_us02_n799 ), .A2(_AES_ENC_us02_n798 ), .A3(_AES_ENC_us02_n797 ), .ZN(_AES_ENC_us02_n808 ) );
NOR2_X2 _AES_ENC_us02_U404  ( .A1(_AES_ENC_us02_n669 ), .A2(_AES_ENC_us02_n668 ), .ZN(_AES_ENC_us02_n673 ) );
NOR4_X2 _AES_ENC_us02_U403  ( .A1(_AES_ENC_us02_n946 ), .A2(_AES_ENC_us02_n1046 ), .A3(_AES_ENC_us02_n671 ), .A4(_AES_ENC_us02_n670 ), .ZN(_AES_ENC_us02_n672 ) );
NOR3_X2 _AES_ENC_us02_U401  ( .A1(_AES_ENC_us02_n1101 ), .A2(_AES_ENC_us02_n1100 ), .A3(_AES_ENC_us02_n1099 ), .ZN(_AES_ENC_us02_n1109 ) );
NOR4_X2 _AES_ENC_us02_U400  ( .A1(_AES_ENC_us02_n843 ), .A2(_AES_ENC_us02_n842 ), .A3(_AES_ENC_us02_n841 ), .A4(_AES_ENC_us02_n840 ), .ZN(_AES_ENC_us02_n844 ) );
NOR4_X2 _AES_ENC_us02_U399  ( .A1(_AES_ENC_us02_n963 ), .A2(_AES_ENC_us02_n962 ), .A3(_AES_ENC_us02_n961 ), .A4(_AES_ENC_us02_n960 ), .ZN(_AES_ENC_us02_n964 ) );
NOR3_X2 _AES_ENC_us02_U398  ( .A1(_AES_ENC_us02_n743 ), .A2(_AES_ENC_us02_n742 ), .A3(_AES_ENC_us02_n741 ), .ZN(_AES_ENC_us02_n744 ) );
NOR2_X2 _AES_ENC_us02_U397  ( .A1(_AES_ENC_us02_n697 ), .A2(_AES_ENC_us02_n658 ), .ZN(_AES_ENC_us02_n659 ) );
NOR2_X2 _AES_ENC_us02_U396  ( .A1(_AES_ENC_us02_n598 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n885 ) );
NOR2_X2 _AES_ENC_us02_U393  ( .A1(_AES_ENC_us02_n623 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n882 ) );
NOR2_X2 _AES_ENC_us02_U390  ( .A1(_AES_ENC_us02_n1053 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n884 ) );
NOR4_X2 _AES_ENC_us02_U389  ( .A1(_AES_ENC_us02_n885 ), .A2(_AES_ENC_us02_n884 ), .A3(_AES_ENC_us02_n883 ), .A4(_AES_ENC_us02_n882 ), .ZN(_AES_ENC_us02_n886 ) );
NOR2_X2 _AES_ENC_us02_U388  ( .A1(_AES_ENC_us02_n1078 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n1033 ) );
NOR2_X2 _AES_ENC_us02_U387  ( .A1(_AES_ENC_us02_n1031 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n1032 ) );
NOR3_X2 _AES_ENC_us02_U386  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n1025 ), .A3(_AES_ENC_us02_n1074 ), .ZN(_AES_ENC_us02_n1035 ) );
NOR4_X2 _AES_ENC_us02_U385  ( .A1(_AES_ENC_us02_n1035 ), .A2(_AES_ENC_us02_n1034 ), .A3(_AES_ENC_us02_n1033 ), .A4(_AES_ENC_us02_n1032 ), .ZN(_AES_ENC_us02_n1036 ) );
NOR2_X2 _AES_ENC_us02_U384  ( .A1(_AES_ENC_us02_n825 ), .A2(_AES_ENC_us02_n578 ), .ZN(_AES_ENC_us02_n830 ) );
NOR2_X2 _AES_ENC_us02_U383  ( .A1(_AES_ENC_us02_n827 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n829 ) );
NOR2_X2 _AES_ENC_us02_U382  ( .A1(_AES_ENC_us02_n572 ), .A2(_AES_ENC_us02_n579 ), .ZN(_AES_ENC_us02_n828 ) );
NOR4_X2 _AES_ENC_us02_U374  ( .A1(_AES_ENC_us02_n831 ), .A2(_AES_ENC_us02_n830 ), .A3(_AES_ENC_us02_n829 ), .A4(_AES_ENC_us02_n828 ), .ZN(_AES_ENC_us02_n832 ) );
NOR2_X2 _AES_ENC_us02_U373  ( .A1(_AES_ENC_us02_n606 ), .A2(_AES_ENC_us02_n582 ), .ZN(_AES_ENC_us02_n1104 ) );
NOR2_X2 _AES_ENC_us02_U372  ( .A1(_AES_ENC_us02_n1102 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n1106 ) );
NOR2_X2 _AES_ENC_us02_U370  ( .A1(_AES_ENC_us02_n1103 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n1105 ) );
NOR4_X2 _AES_ENC_us02_U369  ( .A1(_AES_ENC_us02_n1107 ), .A2(_AES_ENC_us02_n1106 ), .A3(_AES_ENC_us02_n1105 ), .A4(_AES_ENC_us02_n1104 ), .ZN(_AES_ENC_us02_n1108 ) );
NOR3_X2 _AES_ENC_us02_U368  ( .A1(_AES_ENC_us02_n959 ), .A2(_AES_ENC_us02_n621 ), .A3(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n963 ) );
NOR2_X2 _AES_ENC_us02_U367  ( .A1(_AES_ENC_us02_n626 ), .A2(_AES_ENC_us02_n627 ), .ZN(_AES_ENC_us02_n1114 ) );
INV_X4 _AES_ENC_us02_U366  ( .A(_AES_ENC_us02_n1024 ), .ZN(_AES_ENC_us02_n606 ) );
NOR3_X2 _AES_ENC_us02_U365  ( .A1(_AES_ENC_us02_n910 ), .A2(_AES_ENC_us02_n1059 ), .A3(_AES_ENC_us02_n611 ), .ZN(_AES_ENC_us02_n1115 ) );
INV_X4 _AES_ENC_us02_U364  ( .A(_AES_ENC_us02_n1094 ), .ZN(_AES_ENC_us02_n613 ) );
NOR2_X2 _AES_ENC_us02_U363  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n931 ), .ZN(_AES_ENC_us02_n1100 ) );
INV_X4 _AES_ENC_us02_U354  ( .A(_AES_ENC_us02_n1093 ), .ZN(_AES_ENC_us02_n617 ) );
NOR2_X2 _AES_ENC_us02_U353  ( .A1(_AES_ENC_us02_n569 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n929 ) );
NOR2_X2 _AES_ENC_us02_U352  ( .A1(_AES_ENC_us02_n620 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n926 ) );
NOR2_X2 _AES_ENC_us02_U351  ( .A1(_AES_ENC_us02_n572 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n1095 ) );
NOR2_X2 _AES_ENC_us02_U350  ( .A1(_AES_ENC_us02_n609 ), .A2(_AES_ENC_us02_n627 ), .ZN(_AES_ENC_us02_n1010 ) );
NOR2_X2 _AES_ENC_us02_U349  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n1103 ) );
NOR2_X2 _AES_ENC_us02_U348  ( .A1(_AES_ENC_us02_n622 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n1059 ) );
NOR2_X2 _AES_ENC_us02_U347  ( .A1(_AES_ENC_sa02[1]), .A2(_AES_ENC_us02_n1120 ), .ZN(_AES_ENC_us02_n1022 ) );
NOR2_X2 _AES_ENC_us02_U346  ( .A1(_AES_ENC_us02_n619 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n911 ) );
NOR2_X2 _AES_ENC_us02_U345  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_us02_n1025 ), .ZN(_AES_ENC_us02_n826 ) );
NOR2_X2 _AES_ENC_us02_U338  ( .A1(_AES_ENC_us02_n626 ), .A2(_AES_ENC_us02_n607 ), .ZN(_AES_ENC_us02_n1072 ) );
NOR2_X2 _AES_ENC_us02_U335  ( .A1(_AES_ENC_us02_n627 ), .A2(_AES_ENC_us02_n616 ), .ZN(_AES_ENC_us02_n956 ) );
NOR2_X2 _AES_ENC_us02_U329  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_us02_n624 ), .ZN(_AES_ENC_us02_n1121 ) );
NOR2_X2 _AES_ENC_us02_U328  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_us02_n624 ), .ZN(_AES_ENC_us02_n1058 ) );
NOR2_X2 _AES_ENC_us02_U327  ( .A1(_AES_ENC_us02_n625 ), .A2(_AES_ENC_us02_n611 ), .ZN(_AES_ENC_us02_n1073 ) );
NOR2_X2 _AES_ENC_us02_U325  ( .A1(_AES_ENC_sa02[1]), .A2(_AES_ENC_us02_n1025 ), .ZN(_AES_ENC_us02_n1054 ) );
NOR2_X2 _AES_ENC_us02_U324  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_us02_n931 ), .ZN(_AES_ENC_us02_n1029 ) );
NOR2_X2 _AES_ENC_us02_U319  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n1056 ) );
NOR2_X2 _AES_ENC_us02_U318  ( .A1(_AES_ENC_us02_n614 ), .A2(_AES_ENC_us02_n626 ), .ZN(_AES_ENC_us02_n1050 ) );
NOR2_X2 _AES_ENC_us02_U317  ( .A1(_AES_ENC_us02_n1121 ), .A2(_AES_ENC_us02_n1025 ), .ZN(_AES_ENC_us02_n1120 ) );
NOR2_X2 _AES_ENC_us02_U316  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_us02_n572 ), .ZN(_AES_ENC_us02_n1074 ) );
NOR2_X2 _AES_ENC_us02_U315  ( .A1(_AES_ENC_us02_n1058 ), .A2(_AES_ENC_us02_n1054 ), .ZN(_AES_ENC_us02_n878 ) );
NOR2_X2 _AES_ENC_us02_U314  ( .A1(_AES_ENC_us02_n878 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n879 ) );
NOR2_X2 _AES_ENC_us02_U312  ( .A1(_AES_ENC_us02_n880 ), .A2(_AES_ENC_us02_n879 ), .ZN(_AES_ENC_us02_n887 ) );
NOR2_X2 _AES_ENC_us02_U311  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n588 ), .ZN(_AES_ENC_us02_n957 ) );
NOR2_X2 _AES_ENC_us02_U310  ( .A1(_AES_ENC_us02_n958 ), .A2(_AES_ENC_us02_n957 ), .ZN(_AES_ENC_us02_n965 ) );
NOR3_X2 _AES_ENC_us02_U309  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n1091 ), .A3(_AES_ENC_us02_n1022 ), .ZN(_AES_ENC_us02_n720 ) );
NOR3_X2 _AES_ENC_us02_U303  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n1054 ), .A3(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n719 ) );
NOR2_X2 _AES_ENC_us02_U302  ( .A1(_AES_ENC_us02_n720 ), .A2(_AES_ENC_us02_n719 ), .ZN(_AES_ENC_us02_n726 ) );
NOR2_X2 _AES_ENC_us02_U300  ( .A1(_AES_ENC_us02_n614 ), .A2(_AES_ENC_us02_n591 ), .ZN(_AES_ENC_us02_n865 ) );
NOR2_X2 _AES_ENC_us02_U299  ( .A1(_AES_ENC_us02_n1059 ), .A2(_AES_ENC_us02_n1058 ), .ZN(_AES_ENC_us02_n1060 ) );
NOR2_X2 _AES_ENC_us02_U298  ( .A1(_AES_ENC_us02_n1095 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n668 ) );
NOR2_X2 _AES_ENC_us02_U297  ( .A1(_AES_ENC_us02_n911 ), .A2(_AES_ENC_us02_n910 ), .ZN(_AES_ENC_us02_n912 ) );
NOR2_X2 _AES_ENC_us02_U296  ( .A1(_AES_ENC_us02_n912 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n916 ) );
NOR2_X2 _AES_ENC_us02_U295  ( .A1(_AES_ENC_us02_n826 ), .A2(_AES_ENC_us02_n573 ), .ZN(_AES_ENC_us02_n750 ) );
NOR2_X2 _AES_ENC_us02_U294  ( .A1(_AES_ENC_us02_n750 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n751 ) );
NOR2_X2 _AES_ENC_us02_U293  ( .A1(_AES_ENC_us02_n907 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n908 ) );
NOR2_X2 _AES_ENC_us02_U292  ( .A1(_AES_ENC_us02_n990 ), .A2(_AES_ENC_us02_n926 ), .ZN(_AES_ENC_us02_n780 ) );
NOR2_X2 _AES_ENC_us02_U291  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n584 ), .ZN(_AES_ENC_us02_n838 ) );
NOR2_X2 _AES_ENC_us02_U290  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n602 ), .ZN(_AES_ENC_us02_n837 ) );
NOR2_X2 _AES_ENC_us02_U284  ( .A1(_AES_ENC_us02_n838 ), .A2(_AES_ENC_us02_n837 ), .ZN(_AES_ENC_us02_n845 ) );
NOR2_X2 _AES_ENC_us02_U283  ( .A1(_AES_ENC_us02_n1022 ), .A2(_AES_ENC_us02_n1058 ), .ZN(_AES_ENC_us02_n740 ) );
NOR2_X2 _AES_ENC_us02_U282  ( .A1(_AES_ENC_us02_n740 ), .A2(_AES_ENC_us02_n616 ), .ZN(_AES_ENC_us02_n742 ) );
NOR2_X2 _AES_ENC_us02_U281  ( .A1(_AES_ENC_us02_n1098 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n1099 ) );
NOR2_X2 _AES_ENC_us02_U280  ( .A1(_AES_ENC_us02_n1120 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n993 ) );
NOR2_X2 _AES_ENC_us02_U279  ( .A1(_AES_ENC_us02_n993 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n994 ) );
NOR2_X2 _AES_ENC_us02_U273  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n620 ), .ZN(_AES_ENC_us02_n1026 ) );
NOR2_X2 _AES_ENC_us02_U272  ( .A1(_AES_ENC_us02_n573 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n1027 ) );
NOR2_X2 _AES_ENC_us02_U271  ( .A1(_AES_ENC_us02_n1027 ), .A2(_AES_ENC_us02_n1026 ), .ZN(_AES_ENC_us02_n1028 ) );
NOR2_X2 _AES_ENC_us02_U270  ( .A1(_AES_ENC_us02_n1029 ), .A2(_AES_ENC_us02_n1028 ), .ZN(_AES_ENC_us02_n1034 ) );
NOR4_X2 _AES_ENC_us02_U269  ( .A1(_AES_ENC_us02_n757 ), .A2(_AES_ENC_us02_n756 ), .A3(_AES_ENC_us02_n755 ), .A4(_AES_ENC_us02_n754 ), .ZN(_AES_ENC_us02_n758 ) );
NOR2_X2 _AES_ENC_us02_U268  ( .A1(_AES_ENC_us02_n752 ), .A2(_AES_ENC_us02_n751 ), .ZN(_AES_ENC_us02_n759 ) );
NOR2_X2 _AES_ENC_us02_U267  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n1071 ), .ZN(_AES_ENC_us02_n669 ) );
NOR2_X2 _AES_ENC_us02_U263  ( .A1(_AES_ENC_us02_n1056 ), .A2(_AES_ENC_us02_n990 ), .ZN(_AES_ENC_us02_n991 ) );
NOR2_X2 _AES_ENC_us02_U262  ( .A1(_AES_ENC_us02_n991 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n995 ) );
NOR2_X2 _AES_ENC_us02_U258  ( .A1(_AES_ENC_us02_n607 ), .A2(_AES_ENC_us02_n590 ), .ZN(_AES_ENC_us02_n1008 ) );
NOR2_X2 _AES_ENC_us02_U255  ( .A1(_AES_ENC_us02_n839 ), .A2(_AES_ENC_us02_n582 ), .ZN(_AES_ENC_us02_n693 ) );
NOR2_X2 _AES_ENC_us02_U254  ( .A1(_AES_ENC_us02_n606 ), .A2(_AES_ENC_us02_n906 ), .ZN(_AES_ENC_us02_n741 ) );
NOR2_X2 _AES_ENC_us02_U253  ( .A1(_AES_ENC_us02_n1054 ), .A2(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n763 ) );
NOR2_X2 _AES_ENC_us02_U252  ( .A1(_AES_ENC_us02_n763 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n769 ) );
NOR2_X2 _AES_ENC_us02_U251  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n577 ), .ZN(_AES_ENC_us02_n1007 ) );
NOR2_X2 _AES_ENC_us02_U250  ( .A1(_AES_ENC_us02_n609 ), .A2(_AES_ENC_us02_n580 ), .ZN(_AES_ENC_us02_n1123 ) );
NOR2_X2 _AES_ENC_us02_U243  ( .A1(_AES_ENC_us02_n609 ), .A2(_AES_ENC_us02_n590 ), .ZN(_AES_ENC_us02_n710 ) );
INV_X4 _AES_ENC_us02_U242  ( .A(_AES_ENC_us02_n1029 ), .ZN(_AES_ENC_us02_n582 ) );
NOR2_X2 _AES_ENC_us02_U241  ( .A1(_AES_ENC_us02_n616 ), .A2(_AES_ENC_us02_n597 ), .ZN(_AES_ENC_us02_n883 ) );
NOR2_X2 _AES_ENC_us02_U240  ( .A1(_AES_ENC_us02_n593 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n1125 ) );
NOR2_X2 _AES_ENC_us02_U239  ( .A1(_AES_ENC_us02_n990 ), .A2(_AES_ENC_us02_n929 ), .ZN(_AES_ENC_us02_n892 ) );
NOR2_X2 _AES_ENC_us02_U238  ( .A1(_AES_ENC_us02_n892 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n893 ) );
NOR2_X2 _AES_ENC_us02_U237  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n602 ), .ZN(_AES_ENC_us02_n950 ) );
NOR2_X2 _AES_ENC_us02_U236  ( .A1(_AES_ENC_us02_n1079 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n1082 ) );
NOR2_X2 _AES_ENC_us02_U235  ( .A1(_AES_ENC_us02_n910 ), .A2(_AES_ENC_us02_n1056 ), .ZN(_AES_ENC_us02_n941 ) );
NOR2_X2 _AES_ENC_us02_U234  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n1077 ), .ZN(_AES_ENC_us02_n841 ) );
NOR2_X2 _AES_ENC_us02_U229  ( .A1(_AES_ENC_us02_n623 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n630 ) );
NOR2_X2 _AES_ENC_us02_U228  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n602 ), .ZN(_AES_ENC_us02_n806 ) );
NOR2_X2 _AES_ENC_us02_U227  ( .A1(_AES_ENC_us02_n623 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n948 ) );
NOR2_X2 _AES_ENC_us02_U226  ( .A1(_AES_ENC_us02_n606 ), .A2(_AES_ENC_us02_n589 ), .ZN(_AES_ENC_us02_n997 ) );
NOR2_X2 _AES_ENC_us02_U225  ( .A1(_AES_ENC_us02_n1121 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n1122 ) );
NOR2_X2 _AES_ENC_us02_U223  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n1023 ), .ZN(_AES_ENC_us02_n756 ) );
NOR2_X2 _AES_ENC_us02_U222  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n602 ), .ZN(_AES_ENC_us02_n870 ) );
NOR2_X2 _AES_ENC_us02_U221  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n569 ), .ZN(_AES_ENC_us02_n947 ) );
NOR2_X2 _AES_ENC_us02_U217  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n1077 ), .ZN(_AES_ENC_us02_n1084 ) );
NOR2_X2 _AES_ENC_us02_U213  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n855 ), .ZN(_AES_ENC_us02_n709 ) );
NOR2_X2 _AES_ENC_us02_U212  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n589 ), .ZN(_AES_ENC_us02_n868 ) );
NOR2_X2 _AES_ENC_us02_U211  ( .A1(_AES_ENC_us02_n1120 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n1124 ) );
NOR2_X2 _AES_ENC_us02_U210  ( .A1(_AES_ENC_us02_n1120 ), .A2(_AES_ENC_us02_n839 ), .ZN(_AES_ENC_us02_n842 ) );
NOR2_X2 _AES_ENC_us02_U209  ( .A1(_AES_ENC_us02_n1120 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n696 ) );
NOR2_X2 _AES_ENC_us02_U208  ( .A1(_AES_ENC_us02_n1074 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n1076 ) );
NOR2_X2 _AES_ENC_us02_U207  ( .A1(_AES_ENC_us02_n1074 ), .A2(_AES_ENC_us02_n620 ), .ZN(_AES_ENC_us02_n781 ) );
NOR3_X2 _AES_ENC_us02_U201  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n1056 ), .A3(_AES_ENC_us02_n990 ), .ZN(_AES_ENC_us02_n979 ) );
NOR3_X2 _AES_ENC_us02_U200  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n1058 ), .A3(_AES_ENC_us02_n1059 ), .ZN(_AES_ENC_us02_n854 ) );
NOR2_X2 _AES_ENC_us02_U199  ( .A1(_AES_ENC_us02_n996 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n869 ) );
NOR2_X2 _AES_ENC_us02_U198  ( .A1(_AES_ENC_us02_n1056 ), .A2(_AES_ENC_us02_n1074 ), .ZN(_AES_ENC_us02_n1057 ) );
NOR3_X2 _AES_ENC_us02_U197  ( .A1(_AES_ENC_us02_n607 ), .A2(_AES_ENC_us02_n1120 ), .A3(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n978 ) );
NOR2_X2 _AES_ENC_us02_U196  ( .A1(_AES_ENC_us02_n996 ), .A2(_AES_ENC_us02_n911 ), .ZN(_AES_ENC_us02_n1116 ) );
NOR2_X2 _AES_ENC_us02_U195  ( .A1(_AES_ENC_us02_n1074 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n754 ) );
NOR2_X2 _AES_ENC_us02_U194  ( .A1(_AES_ENC_us02_n926 ), .A2(_AES_ENC_us02_n1103 ), .ZN(_AES_ENC_us02_n977 ) );
NOR2_X2 _AES_ENC_us02_U187  ( .A1(_AES_ENC_us02_n839 ), .A2(_AES_ENC_us02_n824 ), .ZN(_AES_ENC_us02_n1092 ) );
NOR2_X2 _AES_ENC_us02_U186  ( .A1(_AES_ENC_us02_n573 ), .A2(_AES_ENC_us02_n1074 ), .ZN(_AES_ENC_us02_n684 ) );
NOR2_X2 _AES_ENC_us02_U185  ( .A1(_AES_ENC_us02_n826 ), .A2(_AES_ENC_us02_n1059 ), .ZN(_AES_ENC_us02_n907 ) );
NOR3_X2 _AES_ENC_us02_U184  ( .A1(_AES_ENC_us02_n625 ), .A2(_AES_ENC_us02_n1115 ), .A3(_AES_ENC_us02_n585 ), .ZN(_AES_ENC_us02_n831 ) );
NOR3_X2 _AES_ENC_us02_U183  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n1056 ), .A3(_AES_ENC_us02_n990 ), .ZN(_AES_ENC_us02_n896 ) );
NOR3_X2 _AES_ENC_us02_U182  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n573 ), .A3(_AES_ENC_us02_n1013 ), .ZN(_AES_ENC_us02_n670 ) );
NOR3_X2 _AES_ENC_us02_U181  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n1091 ), .A3(_AES_ENC_us02_n1022 ), .ZN(_AES_ENC_us02_n843 ) );
NOR2_X2 _AES_ENC_us02_U180  ( .A1(_AES_ENC_us02_n1029 ), .A2(_AES_ENC_us02_n1095 ), .ZN(_AES_ENC_us02_n735 ) );
NAND3_X2 _AES_ENC_us02_U174  ( .A1(_AES_ENC_us02_n569 ), .A2(_AES_ENC_us02_n582 ), .A3(_AES_ENC_us02_n681 ), .ZN(_AES_ENC_us02_n691 ) );
NOR2_X2 _AES_ENC_us02_U173  ( .A1(_AES_ENC_us02_n683 ), .A2(_AES_ENC_us02_n682 ), .ZN(_AES_ENC_us02_n690 ) );
NOR3_X2 _AES_ENC_us02_U172  ( .A1(_AES_ENC_us02_n695 ), .A2(_AES_ENC_us02_n694 ), .A3(_AES_ENC_us02_n693 ), .ZN(_AES_ENC_us02_n700 ) );
NOR4_X2 _AES_ENC_us02_U171  ( .A1(_AES_ENC_us02_n983 ), .A2(_AES_ENC_us02_n698 ), .A3(_AES_ENC_us02_n697 ), .A4(_AES_ENC_us02_n696 ), .ZN(_AES_ENC_us02_n699 ) );
NOR2_X2 _AES_ENC_us02_U170  ( .A1(_AES_ENC_us02_n1100 ), .A2(_AES_ENC_us02_n854 ), .ZN(_AES_ENC_us02_n860 ) );
NOR4_X2 _AES_ENC_us02_U169  ( .A1(_AES_ENC_us02_n1125 ), .A2(_AES_ENC_us02_n1124 ), .A3(_AES_ENC_us02_n1123 ), .A4(_AES_ENC_us02_n1122 ), .ZN(_AES_ENC_us02_n1126 ) );
NOR4_X2 _AES_ENC_us02_U168  ( .A1(_AES_ENC_us02_n1084 ), .A2(_AES_ENC_us02_n1083 ), .A3(_AES_ENC_us02_n1082 ), .A4(_AES_ENC_us02_n1081 ), .ZN(_AES_ENC_us02_n1085 ) );
NOR2_X2 _AES_ENC_us02_U162  ( .A1(_AES_ENC_us02_n1076 ), .A2(_AES_ENC_us02_n1075 ), .ZN(_AES_ENC_us02_n1086 ) );
NOR4_X2 _AES_ENC_us02_U161  ( .A1(_AES_ENC_us02_n896 ), .A2(_AES_ENC_us02_n895 ), .A3(_AES_ENC_us02_n894 ), .A4(_AES_ENC_us02_n893 ), .ZN(_AES_ENC_us02_n897 ) );
NOR2_X2 _AES_ENC_us02_U160  ( .A1(_AES_ENC_us02_n866 ), .A2(_AES_ENC_us02_n865 ), .ZN(_AES_ENC_us02_n872 ) );
NOR4_X2 _AES_ENC_us02_U159  ( .A1(_AES_ENC_us02_n870 ), .A2(_AES_ENC_us02_n869 ), .A3(_AES_ENC_us02_n868 ), .A4(_AES_ENC_us02_n867 ), .ZN(_AES_ENC_us02_n871 ) );
NOR2_X2 _AES_ENC_us02_U158  ( .A1(_AES_ENC_us02_n946 ), .A2(_AES_ENC_us02_n945 ), .ZN(_AES_ENC_us02_n952 ) );
NOR4_X2 _AES_ENC_us02_U157  ( .A1(_AES_ENC_us02_n950 ), .A2(_AES_ENC_us02_n949 ), .A3(_AES_ENC_us02_n948 ), .A4(_AES_ENC_us02_n947 ), .ZN(_AES_ENC_us02_n951 ) );
NOR4_X2 _AES_ENC_us02_U156  ( .A1(_AES_ENC_us02_n983 ), .A2(_AES_ENC_us02_n982 ), .A3(_AES_ENC_us02_n981 ), .A4(_AES_ENC_us02_n980 ), .ZN(_AES_ENC_us02_n984 ) );
NOR2_X2 _AES_ENC_us02_U155  ( .A1(_AES_ENC_us02_n979 ), .A2(_AES_ENC_us02_n978 ), .ZN(_AES_ENC_us02_n985 ) );
NOR3_X2 _AES_ENC_us02_U154  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n1054 ), .A3(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n961 ) );
NOR3_X2 _AES_ENC_us02_U153  ( .A1(_AES_ENC_us02_n620 ), .A2(_AES_ENC_us02_n1074 ), .A3(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n671 ) );
NOR2_X2 _AES_ENC_us02_U152  ( .A1(_AES_ENC_us02_n1057 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n1062 ) );
NOR2_X2 _AES_ENC_us02_U143  ( .A1(_AES_ENC_us02_n1055 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n1063 ) );
NOR2_X2 _AES_ENC_us02_U142  ( .A1(_AES_ENC_us02_n1060 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n1061 ) );
NOR4_X2 _AES_ENC_us02_U141  ( .A1(_AES_ENC_us02_n1064 ), .A2(_AES_ENC_us02_n1063 ), .A3(_AES_ENC_us02_n1062 ), .A4(_AES_ENC_us02_n1061 ), .ZN(_AES_ENC_us02_n1065 ) );
NOR2_X2 _AES_ENC_us02_U140  ( .A1(_AES_ENC_us02_n735 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n687 ) );
NOR2_X2 _AES_ENC_us02_U132  ( .A1(_AES_ENC_us02_n684 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n688 ) );
NOR2_X2 _AES_ENC_us02_U131  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n600 ), .ZN(_AES_ENC_us02_n686 ) );
NOR4_X2 _AES_ENC_us02_U130  ( .A1(_AES_ENC_us02_n688 ), .A2(_AES_ENC_us02_n687 ), .A3(_AES_ENC_us02_n686 ), .A4(_AES_ENC_us02_n685 ), .ZN(_AES_ENC_us02_n689 ) );
NOR2_X2 _AES_ENC_us02_U129  ( .A1(_AES_ENC_us02_n616 ), .A2(_AES_ENC_us02_n580 ), .ZN(_AES_ENC_us02_n771 ) );
NOR2_X2 _AES_ENC_us02_U128  ( .A1(_AES_ENC_us02_n1103 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n772 ) );
NOR2_X2 _AES_ENC_us02_U127  ( .A1(_AES_ENC_us02_n610 ), .A2(_AES_ENC_us02_n599 ), .ZN(_AES_ENC_us02_n773 ) );
NOR4_X2 _AES_ENC_us02_U126  ( .A1(_AES_ENC_us02_n773 ), .A2(_AES_ENC_us02_n772 ), .A3(_AES_ENC_us02_n771 ), .A4(_AES_ENC_us02_n770 ), .ZN(_AES_ENC_us02_n774 ) );
NOR2_X2 _AES_ENC_us02_U121  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n595 ), .ZN(_AES_ENC_us02_n858 ) );
NOR2_X2 _AES_ENC_us02_U120  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n855 ), .ZN(_AES_ENC_us02_n857 ) );
NOR2_X2 _AES_ENC_us02_U119  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n587 ), .ZN(_AES_ENC_us02_n856 ) );
NOR4_X2 _AES_ENC_us02_U118  ( .A1(_AES_ENC_us02_n858 ), .A2(_AES_ENC_us02_n857 ), .A3(_AES_ENC_us02_n856 ), .A4(_AES_ENC_us02_n958 ), .ZN(_AES_ENC_us02_n859 ) );
NOR3_X2 _AES_ENC_us02_U117  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n1120 ), .A3(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n918 ) );
NOR3_X2 _AES_ENC_us02_U116  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n573 ), .A3(_AES_ENC_us02_n1013 ), .ZN(_AES_ENC_us02_n917 ) );
NOR2_X2 _AES_ENC_us02_U115  ( .A1(_AES_ENC_us02_n914 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n915 ) );
NOR4_X2 _AES_ENC_us02_U106  ( .A1(_AES_ENC_us02_n918 ), .A2(_AES_ENC_us02_n917 ), .A3(_AES_ENC_us02_n916 ), .A4(_AES_ENC_us02_n915 ), .ZN(_AES_ENC_us02_n919 ) );
NOR2_X2 _AES_ENC_us02_U105  ( .A1(_AES_ENC_us02_n780 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n784 ) );
NOR2_X2 _AES_ENC_us02_U104  ( .A1(_AES_ENC_us02_n1117 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n782 ) );
NOR2_X2 _AES_ENC_us02_U103  ( .A1(_AES_ENC_us02_n781 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n783 ) );
NOR4_X2 _AES_ENC_us02_U102  ( .A1(_AES_ENC_us02_n880 ), .A2(_AES_ENC_us02_n784 ), .A3(_AES_ENC_us02_n783 ), .A4(_AES_ENC_us02_n782 ), .ZN(_AES_ENC_us02_n785 ) );
NOR2_X2 _AES_ENC_us02_U101  ( .A1(_AES_ENC_us02_n583 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n814 ) );
NOR2_X2 _AES_ENC_us02_U100  ( .A1(_AES_ENC_us02_n907 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n813 ) );
NOR3_X2 _AES_ENC_us02_U95  ( .A1(_AES_ENC_us02_n606 ), .A2(_AES_ENC_us02_n1058 ), .A3(_AES_ENC_us02_n1059 ), .ZN(_AES_ENC_us02_n815 ) );
NOR4_X2 _AES_ENC_us02_U94  ( .A1(_AES_ENC_us02_n815 ), .A2(_AES_ENC_us02_n814 ), .A3(_AES_ENC_us02_n813 ), .A4(_AES_ENC_us02_n812 ), .ZN(_AES_ENC_us02_n816 ) );
NOR2_X2 _AES_ENC_us02_U93  ( .A1(_AES_ENC_us02_n617 ), .A2(_AES_ENC_us02_n569 ), .ZN(_AES_ENC_us02_n721 ) );
NOR2_X2 _AES_ENC_us02_U92  ( .A1(_AES_ENC_us02_n1031 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n723 ) );
NOR2_X2 _AES_ENC_us02_U91  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n1096 ), .ZN(_AES_ENC_us02_n722 ) );
NOR4_X2 _AES_ENC_us02_U90  ( .A1(_AES_ENC_us02_n724 ), .A2(_AES_ENC_us02_n723 ), .A3(_AES_ENC_us02_n722 ), .A4(_AES_ENC_us02_n721 ), .ZN(_AES_ENC_us02_n725 ) );
NOR2_X2 _AES_ENC_us02_U89  ( .A1(_AES_ENC_us02_n911 ), .A2(_AES_ENC_us02_n990 ), .ZN(_AES_ENC_us02_n1009 ) );
NOR2_X2 _AES_ENC_us02_U88  ( .A1(_AES_ENC_us02_n1013 ), .A2(_AES_ENC_us02_n573 ), .ZN(_AES_ENC_us02_n1014 ) );
NOR2_X2 _AES_ENC_us02_U87  ( .A1(_AES_ENC_us02_n1014 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n1015 ) );
NOR4_X2 _AES_ENC_us02_U86  ( .A1(_AES_ENC_us02_n1016 ), .A2(_AES_ENC_us02_n1015 ), .A3(_AES_ENC_us02_n1119 ), .A4(_AES_ENC_us02_n1046 ), .ZN(_AES_ENC_us02_n1017 ) );
NOR2_X2 _AES_ENC_us02_U81  ( .A1(_AES_ENC_us02_n996 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n998 ) );
NOR2_X2 _AES_ENC_us02_U80  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n577 ), .ZN(_AES_ENC_us02_n1000 ) );
NOR2_X2 _AES_ENC_us02_U79  ( .A1(_AES_ENC_us02_n616 ), .A2(_AES_ENC_us02_n1096 ), .ZN(_AES_ENC_us02_n999 ) );
NOR4_X2 _AES_ENC_us02_U78  ( .A1(_AES_ENC_us02_n1000 ), .A2(_AES_ENC_us02_n999 ), .A3(_AES_ENC_us02_n998 ), .A4(_AES_ENC_us02_n997 ), .ZN(_AES_ENC_us02_n1001 ) );
NOR2_X2 _AES_ENC_us02_U74  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n1096 ), .ZN(_AES_ENC_us02_n697 ) );
NOR2_X2 _AES_ENC_us02_U73  ( .A1(_AES_ENC_us02_n620 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n958 ) );
NOR2_X2 _AES_ENC_us02_U72  ( .A1(_AES_ENC_us02_n911 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n983 ) );
NOR2_X2 _AES_ENC_us02_U71  ( .A1(_AES_ENC_us02_n1054 ), .A2(_AES_ENC_us02_n1103 ), .ZN(_AES_ENC_us02_n1031 ) );
INV_X4 _AES_ENC_us02_U65  ( .A(_AES_ENC_us02_n1050 ), .ZN(_AES_ENC_us02_n612 ) );
INV_X4 _AES_ENC_us02_U64  ( .A(_AES_ENC_us02_n1072 ), .ZN(_AES_ENC_us02_n605 ) );
INV_X4 _AES_ENC_us02_U63  ( .A(_AES_ENC_us02_n1073 ), .ZN(_AES_ENC_us02_n604 ) );
NOR2_X2 _AES_ENC_us02_U62  ( .A1(_AES_ENC_us02_n582 ), .A2(_AES_ENC_us02_n613 ), .ZN(_AES_ENC_us02_n880 ) );
NOR3_X2 _AES_ENC_us02_U61  ( .A1(_AES_ENC_us02_n826 ), .A2(_AES_ENC_us02_n1121 ), .A3(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n946 ) );
INV_X4 _AES_ENC_us02_U59  ( .A(_AES_ENC_us02_n1010 ), .ZN(_AES_ENC_us02_n608 ) );
NOR3_X2 _AES_ENC_us02_U58  ( .A1(_AES_ENC_us02_n573 ), .A2(_AES_ENC_us02_n1029 ), .A3(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n1119 ) );
INV_X4 _AES_ENC_us02_U57  ( .A(_AES_ENC_us02_n956 ), .ZN(_AES_ENC_us02_n615 ) );
NOR2_X2 _AES_ENC_us02_U50  ( .A1(_AES_ENC_us02_n623 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n1013 ) );
NOR2_X2 _AES_ENC_us02_U49  ( .A1(_AES_ENC_us02_n620 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n910 ) );
NOR2_X2 _AES_ENC_us02_U48  ( .A1(_AES_ENC_us02_n569 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n1091 ) );
NOR2_X2 _AES_ENC_us02_U47  ( .A1(_AES_ENC_us02_n622 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n990 ) );
NOR2_X2 _AES_ENC_us02_U46  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_us02_n1121 ), .ZN(_AES_ENC_us02_n996 ) );
NOR2_X2 _AES_ENC_us02_U45  ( .A1(_AES_ENC_us02_n610 ), .A2(_AES_ENC_us02_n600 ), .ZN(_AES_ENC_us02_n628 ) );
NOR2_X2 _AES_ENC_us02_U44  ( .A1(_AES_ENC_us02_n576 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n866 ) );
NOR2_X2 _AES_ENC_us02_U43  ( .A1(_AES_ENC_us02_n603 ), .A2(_AES_ENC_us02_n610 ), .ZN(_AES_ENC_us02_n1006 ) );
NOR2_X2 _AES_ENC_us02_U42  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n1117 ), .ZN(_AES_ENC_us02_n1118 ) );
NOR2_X2 _AES_ENC_us02_U41  ( .A1(_AES_ENC_us02_n1119 ), .A2(_AES_ENC_us02_n1118 ), .ZN(_AES_ENC_us02_n1127 ) );
NOR2_X2 _AES_ENC_us02_U36  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n594 ), .ZN(_AES_ENC_us02_n629 ) );
NOR2_X2 _AES_ENC_us02_U35  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n906 ), .ZN(_AES_ENC_us02_n909 ) );
NOR2_X2 _AES_ENC_us02_U34  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n597 ), .ZN(_AES_ENC_us02_n658 ) );
NOR2_X2 _AES_ENC_us02_U33  ( .A1(_AES_ENC_us02_n1116 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n695 ) );
NOR2_X2 _AES_ENC_us02_U32  ( .A1(_AES_ENC_us02_n1078 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n1083 ) );
NOR2_X2 _AES_ENC_us02_U31  ( .A1(_AES_ENC_us02_n941 ), .A2(_AES_ENC_us02_n608 ), .ZN(_AES_ENC_us02_n724 ) );
NOR2_X2 _AES_ENC_us02_U30  ( .A1(_AES_ENC_us02_n598 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n1107 ) );
NOR2_X2 _AES_ENC_us02_U29  ( .A1(_AES_ENC_us02_n576 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n840 ) );
NOR2_X2 _AES_ENC_us02_U24  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n593 ), .ZN(_AES_ENC_us02_n633 ) );
NOR2_X2 _AES_ENC_us02_U23  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n1080 ), .ZN(_AES_ENC_us02_n1081 ) );
NOR2_X2 _AES_ENC_us02_U21  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n1045 ), .ZN(_AES_ENC_us02_n812 ) );
NOR2_X2 _AES_ENC_us02_U20  ( .A1(_AES_ENC_us02_n1009 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n960 ) );
NOR2_X2 _AES_ENC_us02_U19  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n601 ), .ZN(_AES_ENC_us02_n982 ) );
NOR2_X2 _AES_ENC_us02_U18  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n594 ), .ZN(_AES_ENC_us02_n757 ) );
NOR2_X2 _AES_ENC_us02_U17  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n590 ), .ZN(_AES_ENC_us02_n698 ) );
NOR2_X2 _AES_ENC_us02_U16  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n619 ), .ZN(_AES_ENC_us02_n708 ) );
NOR2_X2 _AES_ENC_us02_U15  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n582 ), .ZN(_AES_ENC_us02_n770 ) );
NOR2_X2 _AES_ENC_us02_U10  ( .A1(_AES_ENC_us02_n619 ), .A2(_AES_ENC_us02_n604 ), .ZN(_AES_ENC_us02_n803 ) );
NOR2_X2 _AES_ENC_us02_U9  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n881 ), .ZN(_AES_ENC_us02_n711 ) );
NOR2_X2 _AES_ENC_us02_U8  ( .A1(_AES_ENC_us02_n615 ), .A2(_AES_ENC_us02_n582 ), .ZN(_AES_ENC_us02_n867 ) );
NOR2_X2 _AES_ENC_us02_U7  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n599 ), .ZN(_AES_ENC_us02_n804 ) );
NOR2_X2 _AES_ENC_us02_U6  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n620 ), .ZN(_AES_ENC_us02_n1046 ) );
OR2_X4 _AES_ENC_us02_U5  ( .A1(_AES_ENC_us02_n624 ), .A2(_AES_ENC_sa02[1]),.ZN(_AES_ENC_us02_n570 ) );
OR2_X4 _AES_ENC_us02_U4  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_sa02[4]),.ZN(_AES_ENC_us02_n569 ) );
NAND2_X2 _AES_ENC_us02_U514  ( .A1(_AES_ENC_us02_n1121 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n1030 ) );
AND2_X2 _AES_ENC_us02_U513  ( .A1(_AES_ENC_us02_n597 ), .A2(_AES_ENC_us02_n1030 ), .ZN(_AES_ENC_us02_n1049 ) );
NAND2_X2 _AES_ENC_us02_U511  ( .A1(_AES_ENC_us02_n1049 ), .A2(_AES_ENC_us02_n794 ), .ZN(_AES_ENC_us02_n637 ) );
AND2_X2 _AES_ENC_us02_U493  ( .A1(_AES_ENC_us02_n779 ), .A2(_AES_ENC_us02_n996 ), .ZN(_AES_ENC_us02_n632 ) );
NAND4_X2 _AES_ENC_us02_U485  ( .A1(_AES_ENC_us02_n637 ), .A2(_AES_ENC_us02_n636 ), .A3(_AES_ENC_us02_n635 ), .A4(_AES_ENC_us02_n634 ), .ZN(_AES_ENC_us02_n638 ) );
NAND2_X2 _AES_ENC_us02_U484  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n638 ), .ZN(_AES_ENC_us02_n679 ) );
NAND2_X2 _AES_ENC_us02_U481  ( .A1(_AES_ENC_us02_n1094 ), .A2(_AES_ENC_us02_n591 ), .ZN(_AES_ENC_us02_n648 ) );
NAND2_X2 _AES_ENC_us02_U476  ( .A1(_AES_ENC_us02_n601 ), .A2(_AES_ENC_us02_n590 ), .ZN(_AES_ENC_us02_n762 ) );
NAND2_X2 _AES_ENC_us02_U475  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n762 ), .ZN(_AES_ENC_us02_n647 ) );
NAND4_X2 _AES_ENC_us02_U457  ( .A1(_AES_ENC_us02_n648 ), .A2(_AES_ENC_us02_n647 ), .A3(_AES_ENC_us02_n646 ), .A4(_AES_ENC_us02_n645 ), .ZN(_AES_ENC_us02_n649 ) );
NAND2_X2 _AES_ENC_us02_U456  ( .A1(_AES_ENC_sa02[0]), .A2(_AES_ENC_us02_n649 ), .ZN(_AES_ENC_us02_n665 ) );
NAND2_X2 _AES_ENC_us02_U454  ( .A1(_AES_ENC_us02_n596 ), .A2(_AES_ENC_us02_n623 ), .ZN(_AES_ENC_us02_n855 ) );
NAND2_X2 _AES_ENC_us02_U453  ( .A1(_AES_ENC_us02_n587 ), .A2(_AES_ENC_us02_n855 ), .ZN(_AES_ENC_us02_n821 ) );
NAND2_X2 _AES_ENC_us02_U452  ( .A1(_AES_ENC_us02_n1093 ), .A2(_AES_ENC_us02_n821 ), .ZN(_AES_ENC_us02_n662 ) );
NAND2_X2 _AES_ENC_us02_U451  ( .A1(_AES_ENC_us02_n619 ), .A2(_AES_ENC_us02_n589 ), .ZN(_AES_ENC_us02_n650 ) );
NAND2_X2 _AES_ENC_us02_U450  ( .A1(_AES_ENC_us02_n956 ), .A2(_AES_ENC_us02_n650 ), .ZN(_AES_ENC_us02_n661 ) );
NAND2_X2 _AES_ENC_us02_U449  ( .A1(_AES_ENC_us02_n626 ), .A2(_AES_ENC_us02_n627 ), .ZN(_AES_ENC_us02_n839 ) );
OR2_X2 _AES_ENC_us02_U446  ( .A1(_AES_ENC_us02_n839 ), .A2(_AES_ENC_us02_n932 ), .ZN(_AES_ENC_us02_n656 ) );
NAND2_X2 _AES_ENC_us02_U445  ( .A1(_AES_ENC_us02_n621 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n1096 ) );
NAND2_X2 _AES_ENC_us02_U444  ( .A1(_AES_ENC_us02_n1030 ), .A2(_AES_ENC_us02_n1096 ), .ZN(_AES_ENC_us02_n651 ) );
NAND2_X2 _AES_ENC_us02_U443  ( .A1(_AES_ENC_us02_n1114 ), .A2(_AES_ENC_us02_n651 ), .ZN(_AES_ENC_us02_n655 ) );
OR3_X2 _AES_ENC_us02_U440  ( .A1(_AES_ENC_us02_n1079 ), .A2(_AES_ENC_sa02[7]), .A3(_AES_ENC_us02_n626 ), .ZN(_AES_ENC_us02_n654 ));
NAND2_X2 _AES_ENC_us02_U439  ( .A1(_AES_ENC_us02_n593 ), .A2(_AES_ENC_us02_n601 ), .ZN(_AES_ENC_us02_n652 ) );
NAND4_X2 _AES_ENC_us02_U437  ( .A1(_AES_ENC_us02_n656 ), .A2(_AES_ENC_us02_n655 ), .A3(_AES_ENC_us02_n654 ), .A4(_AES_ENC_us02_n653 ), .ZN(_AES_ENC_us02_n657 ) );
NAND2_X2 _AES_ENC_us02_U436  ( .A1(_AES_ENC_sa02[2]), .A2(_AES_ENC_us02_n657 ), .ZN(_AES_ENC_us02_n660 ) );
NAND4_X2 _AES_ENC_us02_U432  ( .A1(_AES_ENC_us02_n662 ), .A2(_AES_ENC_us02_n661 ), .A3(_AES_ENC_us02_n660 ), .A4(_AES_ENC_us02_n659 ), .ZN(_AES_ENC_us02_n663 ) );
NAND2_X2 _AES_ENC_us02_U431  ( .A1(_AES_ENC_us02_n663 ), .A2(_AES_ENC_us02_n574 ), .ZN(_AES_ENC_us02_n664 ) );
NAND2_X2 _AES_ENC_us02_U430  ( .A1(_AES_ENC_us02_n665 ), .A2(_AES_ENC_us02_n664 ), .ZN(_AES_ENC_us02_n666 ) );
NAND2_X2 _AES_ENC_us02_U429  ( .A1(_AES_ENC_sa02[6]), .A2(_AES_ENC_us02_n666 ), .ZN(_AES_ENC_us02_n678 ) );
NAND2_X2 _AES_ENC_us02_U426  ( .A1(_AES_ENC_us02_n735 ), .A2(_AES_ENC_us02_n1093 ), .ZN(_AES_ENC_us02_n675 ) );
NAND2_X2 _AES_ENC_us02_U425  ( .A1(_AES_ENC_us02_n588 ), .A2(_AES_ENC_us02_n597 ), .ZN(_AES_ENC_us02_n1045 ) );
OR2_X2 _AES_ENC_us02_U424  ( .A1(_AES_ENC_us02_n1045 ), .A2(_AES_ENC_us02_n605 ), .ZN(_AES_ENC_us02_n674 ) );
NAND2_X2 _AES_ENC_us02_U423  ( .A1(_AES_ENC_sa02[1]), .A2(_AES_ENC_us02_n620 ), .ZN(_AES_ENC_us02_n667 ) );
NAND2_X2 _AES_ENC_us02_U422  ( .A1(_AES_ENC_us02_n619 ), .A2(_AES_ENC_us02_n667 ), .ZN(_AES_ENC_us02_n1071 ) );
NAND4_X2 _AES_ENC_us02_U412  ( .A1(_AES_ENC_us02_n675 ), .A2(_AES_ENC_us02_n674 ), .A3(_AES_ENC_us02_n673 ), .A4(_AES_ENC_us02_n672 ), .ZN(_AES_ENC_us02_n676 ) );
NAND2_X2 _AES_ENC_us02_U411  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n676 ), .ZN(_AES_ENC_us02_n677 ) );
NAND2_X2 _AES_ENC_us02_U408  ( .A1(_AES_ENC_us02_n800 ), .A2(_AES_ENC_us02_n1022 ), .ZN(_AES_ENC_us02_n680 ) );
NAND2_X2 _AES_ENC_us02_U407  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n680 ), .ZN(_AES_ENC_us02_n681 ) );
AND2_X2 _AES_ENC_us02_U402  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n684 ), .ZN(_AES_ENC_us02_n682 ) );
NAND4_X2 _AES_ENC_us02_U395  ( .A1(_AES_ENC_us02_n691 ), .A2(_AES_ENC_us02_n581 ), .A3(_AES_ENC_us02_n690 ), .A4(_AES_ENC_us02_n689 ), .ZN(_AES_ENC_us02_n692 ) );
NAND2_X2 _AES_ENC_us02_U394  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n692 ), .ZN(_AES_ENC_us02_n733 ) );
NAND2_X2 _AES_ENC_us02_U392  ( .A1(_AES_ENC_us02_n977 ), .A2(_AES_ENC_us02_n1050 ), .ZN(_AES_ENC_us02_n702 ) );
NAND2_X2 _AES_ENC_us02_U391  ( .A1(_AES_ENC_us02_n1093 ), .A2(_AES_ENC_us02_n1045 ), .ZN(_AES_ENC_us02_n701 ) );
NAND4_X2 _AES_ENC_us02_U381  ( .A1(_AES_ENC_us02_n702 ), .A2(_AES_ENC_us02_n701 ), .A3(_AES_ENC_us02_n700 ), .A4(_AES_ENC_us02_n699 ), .ZN(_AES_ENC_us02_n703 ) );
NAND2_X2 _AES_ENC_us02_U380  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n703 ), .ZN(_AES_ENC_us02_n732 ) );
AND2_X2 _AES_ENC_us02_U379  ( .A1(_AES_ENC_sa02[0]), .A2(_AES_ENC_sa02[6]),.ZN(_AES_ENC_us02_n1113 ) );
NAND2_X2 _AES_ENC_us02_U378  ( .A1(_AES_ENC_us02_n601 ), .A2(_AES_ENC_us02_n1030 ), .ZN(_AES_ENC_us02_n881 ) );
NAND2_X2 _AES_ENC_us02_U377  ( .A1(_AES_ENC_us02_n1093 ), .A2(_AES_ENC_us02_n881 ), .ZN(_AES_ENC_us02_n715 ) );
NAND2_X2 _AES_ENC_us02_U376  ( .A1(_AES_ENC_us02_n1010 ), .A2(_AES_ENC_us02_n600 ), .ZN(_AES_ENC_us02_n714 ) );
NAND2_X2 _AES_ENC_us02_U375  ( .A1(_AES_ENC_us02_n855 ), .A2(_AES_ENC_us02_n588 ), .ZN(_AES_ENC_us02_n1117 ) );
XNOR2_X2 _AES_ENC_us02_U371  ( .A(_AES_ENC_us02_n611 ), .B(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n824 ) );
NAND4_X2 _AES_ENC_us02_U362  ( .A1(_AES_ENC_us02_n715 ), .A2(_AES_ENC_us02_n714 ), .A3(_AES_ENC_us02_n713 ), .A4(_AES_ENC_us02_n712 ), .ZN(_AES_ENC_us02_n716 ) );
NAND2_X2 _AES_ENC_us02_U361  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n716 ), .ZN(_AES_ENC_us02_n731 ) );
AND2_X2 _AES_ENC_us02_U360  ( .A1(_AES_ENC_sa02[6]), .A2(_AES_ENC_us02_n574 ), .ZN(_AES_ENC_us02_n1131 ) );
NAND2_X2 _AES_ENC_us02_U359  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n717 ) );
NAND2_X2 _AES_ENC_us02_U358  ( .A1(_AES_ENC_us02_n1029 ), .A2(_AES_ENC_us02_n717 ), .ZN(_AES_ENC_us02_n728 ) );
NAND2_X2 _AES_ENC_us02_U357  ( .A1(_AES_ENC_sa02[1]), .A2(_AES_ENC_us02_n624 ), .ZN(_AES_ENC_us02_n1097 ) );
NAND2_X2 _AES_ENC_us02_U356  ( .A1(_AES_ENC_us02_n603 ), .A2(_AES_ENC_us02_n1097 ), .ZN(_AES_ENC_us02_n718 ) );
NAND2_X2 _AES_ENC_us02_U355  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n718 ), .ZN(_AES_ENC_us02_n727 ) );
NAND4_X2 _AES_ENC_us02_U344  ( .A1(_AES_ENC_us02_n728 ), .A2(_AES_ENC_us02_n727 ), .A3(_AES_ENC_us02_n726 ), .A4(_AES_ENC_us02_n725 ), .ZN(_AES_ENC_us02_n729 ) );
NAND2_X2 _AES_ENC_us02_U343  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n729 ), .ZN(_AES_ENC_us02_n730 ) );
NAND4_X2 _AES_ENC_us02_U342  ( .A1(_AES_ENC_us02_n733 ), .A2(_AES_ENC_us02_n732 ), .A3(_AES_ENC_us02_n731 ), .A4(_AES_ENC_us02_n730 ), .ZN(_AES_ENC_sa02_sub[1] ) );
NAND2_X2 _AES_ENC_us02_U341  ( .A1(_AES_ENC_sa02[7]), .A2(_AES_ENC_us02_n611 ), .ZN(_AES_ENC_us02_n734 ) );
NAND2_X2 _AES_ENC_us02_U340  ( .A1(_AES_ENC_us02_n734 ), .A2(_AES_ENC_us02_n607 ), .ZN(_AES_ENC_us02_n738 ) );
OR4_X2 _AES_ENC_us02_U339  ( .A1(_AES_ENC_us02_n738 ), .A2(_AES_ENC_us02_n626 ), .A3(_AES_ENC_us02_n826 ), .A4(_AES_ENC_us02_n1121 ), .ZN(_AES_ENC_us02_n746 ) );
NAND2_X2 _AES_ENC_us02_U337  ( .A1(_AES_ENC_us02_n1100 ), .A2(_AES_ENC_us02_n587 ), .ZN(_AES_ENC_us02_n992 ) );
OR2_X2 _AES_ENC_us02_U336  ( .A1(_AES_ENC_us02_n610 ), .A2(_AES_ENC_us02_n735 ), .ZN(_AES_ENC_us02_n737 ) );
NAND2_X2 _AES_ENC_us02_U334  ( .A1(_AES_ENC_us02_n619 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n753 ) );
NAND2_X2 _AES_ENC_us02_U333  ( .A1(_AES_ENC_us02_n582 ), .A2(_AES_ENC_us02_n753 ), .ZN(_AES_ENC_us02_n1080 ) );
NAND2_X2 _AES_ENC_us02_U332  ( .A1(_AES_ENC_us02_n1048 ), .A2(_AES_ENC_us02_n576 ), .ZN(_AES_ENC_us02_n736 ) );
NAND2_X2 _AES_ENC_us02_U331  ( .A1(_AES_ENC_us02_n737 ), .A2(_AES_ENC_us02_n736 ), .ZN(_AES_ENC_us02_n739 ) );
NAND2_X2 _AES_ENC_us02_U330  ( .A1(_AES_ENC_us02_n739 ), .A2(_AES_ENC_us02_n738 ), .ZN(_AES_ENC_us02_n745 ) );
NAND2_X2 _AES_ENC_us02_U326  ( .A1(_AES_ENC_us02_n1096 ), .A2(_AES_ENC_us02_n590 ), .ZN(_AES_ENC_us02_n906 ) );
NAND4_X2 _AES_ENC_us02_U323  ( .A1(_AES_ENC_us02_n746 ), .A2(_AES_ENC_us02_n992 ), .A3(_AES_ENC_us02_n745 ), .A4(_AES_ENC_us02_n744 ), .ZN(_AES_ENC_us02_n747 ) );
NAND2_X2 _AES_ENC_us02_U322  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n747 ), .ZN(_AES_ENC_us02_n793 ) );
NAND2_X2 _AES_ENC_us02_U321  ( .A1(_AES_ENC_us02_n584 ), .A2(_AES_ENC_us02_n855 ), .ZN(_AES_ENC_us02_n748 ) );
NAND2_X2 _AES_ENC_us02_U320  ( .A1(_AES_ENC_us02_n956 ), .A2(_AES_ENC_us02_n748 ), .ZN(_AES_ENC_us02_n760 ) );
NAND2_X2 _AES_ENC_us02_U313  ( .A1(_AES_ENC_us02_n590 ), .A2(_AES_ENC_us02_n753 ), .ZN(_AES_ENC_us02_n1023 ) );
NAND4_X2 _AES_ENC_us02_U308  ( .A1(_AES_ENC_us02_n760 ), .A2(_AES_ENC_us02_n992 ), .A3(_AES_ENC_us02_n759 ), .A4(_AES_ENC_us02_n758 ), .ZN(_AES_ENC_us02_n761 ) );
NAND2_X2 _AES_ENC_us02_U307  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n761 ), .ZN(_AES_ENC_us02_n792 ) );
NAND2_X2 _AES_ENC_us02_U306  ( .A1(_AES_ENC_us02_n584 ), .A2(_AES_ENC_us02_n603 ), .ZN(_AES_ENC_us02_n989 ) );
NAND2_X2 _AES_ENC_us02_U305  ( .A1(_AES_ENC_us02_n1050 ), .A2(_AES_ENC_us02_n989 ), .ZN(_AES_ENC_us02_n777 ) );
NAND2_X2 _AES_ENC_us02_U304  ( .A1(_AES_ENC_us02_n1093 ), .A2(_AES_ENC_us02_n762 ), .ZN(_AES_ENC_us02_n776 ) );
XNOR2_X2 _AES_ENC_us02_U301  ( .A(_AES_ENC_sa02[7]), .B(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n959 ) );
NAND4_X2 _AES_ENC_us02_U289  ( .A1(_AES_ENC_us02_n777 ), .A2(_AES_ENC_us02_n776 ), .A3(_AES_ENC_us02_n775 ), .A4(_AES_ENC_us02_n774 ), .ZN(_AES_ENC_us02_n778 ) );
NAND2_X2 _AES_ENC_us02_U288  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n778 ), .ZN(_AES_ENC_us02_n791 ) );
NAND2_X2 _AES_ENC_us02_U287  ( .A1(_AES_ENC_us02_n1056 ), .A2(_AES_ENC_us02_n1050 ), .ZN(_AES_ENC_us02_n788 ) );
NAND2_X2 _AES_ENC_us02_U286  ( .A1(_AES_ENC_us02_n1091 ), .A2(_AES_ENC_us02_n779 ), .ZN(_AES_ENC_us02_n787 ) );
NAND2_X2 _AES_ENC_us02_U285  ( .A1(_AES_ENC_us02_n956 ), .A2(_AES_ENC_sa02[1]), .ZN(_AES_ENC_us02_n786 ) );
NAND4_X2 _AES_ENC_us02_U278  ( .A1(_AES_ENC_us02_n788 ), .A2(_AES_ENC_us02_n787 ), .A3(_AES_ENC_us02_n786 ), .A4(_AES_ENC_us02_n785 ), .ZN(_AES_ENC_us02_n789 ) );
NAND2_X2 _AES_ENC_us02_U277  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n789 ), .ZN(_AES_ENC_us02_n790 ) );
NAND4_X2 _AES_ENC_us02_U276  ( .A1(_AES_ENC_us02_n793 ), .A2(_AES_ENC_us02_n792 ), .A3(_AES_ENC_us02_n791 ), .A4(_AES_ENC_us02_n790 ), .ZN(_AES_ENC_sa02_sub[2] ) );
NAND2_X2 _AES_ENC_us02_U275  ( .A1(_AES_ENC_us02_n1059 ), .A2(_AES_ENC_us02_n794 ), .ZN(_AES_ENC_us02_n810 ) );
NAND2_X2 _AES_ENC_us02_U274  ( .A1(_AES_ENC_us02_n1049 ), .A2(_AES_ENC_us02_n956 ), .ZN(_AES_ENC_us02_n809 ) );
OR2_X2 _AES_ENC_us02_U266  ( .A1(_AES_ENC_us02_n1096 ), .A2(_AES_ENC_us02_n606 ), .ZN(_AES_ENC_us02_n802 ) );
NAND2_X2 _AES_ENC_us02_U265  ( .A1(_AES_ENC_us02_n1053 ), .A2(_AES_ENC_us02_n800 ), .ZN(_AES_ENC_us02_n801 ) );
NAND2_X2 _AES_ENC_us02_U264  ( .A1(_AES_ENC_us02_n802 ), .A2(_AES_ENC_us02_n801 ), .ZN(_AES_ENC_us02_n805 ) );
NAND4_X2 _AES_ENC_us02_U261  ( .A1(_AES_ENC_us02_n810 ), .A2(_AES_ENC_us02_n809 ), .A3(_AES_ENC_us02_n808 ), .A4(_AES_ENC_us02_n807 ), .ZN(_AES_ENC_us02_n811 ) );
NAND2_X2 _AES_ENC_us02_U260  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n811 ), .ZN(_AES_ENC_us02_n852 ) );
OR2_X2 _AES_ENC_us02_U259  ( .A1(_AES_ENC_us02_n1023 ), .A2(_AES_ENC_us02_n617 ), .ZN(_AES_ENC_us02_n819 ) );
OR2_X2 _AES_ENC_us02_U257  ( .A1(_AES_ENC_us02_n570 ), .A2(_AES_ENC_us02_n930 ), .ZN(_AES_ENC_us02_n818 ) );
NAND2_X2 _AES_ENC_us02_U256  ( .A1(_AES_ENC_us02_n1013 ), .A2(_AES_ENC_us02_n1094 ), .ZN(_AES_ENC_us02_n817 ) );
NAND4_X2 _AES_ENC_us02_U249  ( .A1(_AES_ENC_us02_n819 ), .A2(_AES_ENC_us02_n818 ), .A3(_AES_ENC_us02_n817 ), .A4(_AES_ENC_us02_n816 ), .ZN(_AES_ENC_us02_n820 ) );
NAND2_X2 _AES_ENC_us02_U248  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n820 ), .ZN(_AES_ENC_us02_n851 ) );
NAND2_X2 _AES_ENC_us02_U247  ( .A1(_AES_ENC_us02_n956 ), .A2(_AES_ENC_us02_n1080 ), .ZN(_AES_ENC_us02_n835 ) );
NAND2_X2 _AES_ENC_us02_U246  ( .A1(_AES_ENC_us02_n570 ), .A2(_AES_ENC_us02_n1030 ), .ZN(_AES_ENC_us02_n1047 ) );
OR2_X2 _AES_ENC_us02_U245  ( .A1(_AES_ENC_us02_n1047 ), .A2(_AES_ENC_us02_n612 ), .ZN(_AES_ENC_us02_n834 ) );
NAND2_X2 _AES_ENC_us02_U244  ( .A1(_AES_ENC_us02_n1072 ), .A2(_AES_ENC_us02_n589 ), .ZN(_AES_ENC_us02_n833 ) );
NAND4_X2 _AES_ENC_us02_U233  ( .A1(_AES_ENC_us02_n835 ), .A2(_AES_ENC_us02_n834 ), .A3(_AES_ENC_us02_n833 ), .A4(_AES_ENC_us02_n832 ), .ZN(_AES_ENC_us02_n836 ) );
NAND2_X2 _AES_ENC_us02_U232  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n836 ), .ZN(_AES_ENC_us02_n850 ) );
NAND2_X2 _AES_ENC_us02_U231  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n623 ), .ZN(_AES_ENC_us02_n847 ) );
NAND2_X2 _AES_ENC_us02_U230  ( .A1(_AES_ENC_us02_n1050 ), .A2(_AES_ENC_us02_n1071 ), .ZN(_AES_ENC_us02_n846 ) );
OR2_X2 _AES_ENC_us02_U224  ( .A1(_AES_ENC_us02_n1053 ), .A2(_AES_ENC_us02_n911 ), .ZN(_AES_ENC_us02_n1077 ) );
NAND4_X2 _AES_ENC_us02_U220  ( .A1(_AES_ENC_us02_n847 ), .A2(_AES_ENC_us02_n846 ), .A3(_AES_ENC_us02_n845 ), .A4(_AES_ENC_us02_n844 ), .ZN(_AES_ENC_us02_n848 ) );
NAND2_X2 _AES_ENC_us02_U219  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n848 ), .ZN(_AES_ENC_us02_n849 ) );
NAND4_X2 _AES_ENC_us02_U218  ( .A1(_AES_ENC_us02_n852 ), .A2(_AES_ENC_us02_n851 ), .A3(_AES_ENC_us02_n850 ), .A4(_AES_ENC_us02_n849 ), .ZN(_AES_ENC_sa02_sub[3] ) );
NAND2_X2 _AES_ENC_us02_U216  ( .A1(_AES_ENC_us02_n1009 ), .A2(_AES_ENC_us02_n1072 ), .ZN(_AES_ENC_us02_n862 ) );
NAND2_X2 _AES_ENC_us02_U215  ( .A1(_AES_ENC_us02_n603 ), .A2(_AES_ENC_us02_n577 ), .ZN(_AES_ENC_us02_n853 ) );
NAND2_X2 _AES_ENC_us02_U214  ( .A1(_AES_ENC_us02_n1050 ), .A2(_AES_ENC_us02_n853 ), .ZN(_AES_ENC_us02_n861 ) );
NAND4_X2 _AES_ENC_us02_U206  ( .A1(_AES_ENC_us02_n862 ), .A2(_AES_ENC_us02_n861 ), .A3(_AES_ENC_us02_n860 ), .A4(_AES_ENC_us02_n859 ), .ZN(_AES_ENC_us02_n863 ) );
NAND2_X2 _AES_ENC_us02_U205  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n863 ), .ZN(_AES_ENC_us02_n905 ) );
NAND2_X2 _AES_ENC_us02_U204  ( .A1(_AES_ENC_us02_n1010 ), .A2(_AES_ENC_us02_n989 ), .ZN(_AES_ENC_us02_n874 ) );
NAND2_X2 _AES_ENC_us02_U203  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n610 ), .ZN(_AES_ENC_us02_n864 ) );
NAND2_X2 _AES_ENC_us02_U202  ( .A1(_AES_ENC_us02_n929 ), .A2(_AES_ENC_us02_n864 ), .ZN(_AES_ENC_us02_n873 ) );
NAND4_X2 _AES_ENC_us02_U193  ( .A1(_AES_ENC_us02_n874 ), .A2(_AES_ENC_us02_n873 ), .A3(_AES_ENC_us02_n872 ), .A4(_AES_ENC_us02_n871 ), .ZN(_AES_ENC_us02_n875 ) );
NAND2_X2 _AES_ENC_us02_U192  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n875 ), .ZN(_AES_ENC_us02_n904 ) );
NAND2_X2 _AES_ENC_us02_U191  ( .A1(_AES_ENC_us02_n583 ), .A2(_AES_ENC_us02_n1050 ), .ZN(_AES_ENC_us02_n889 ) );
NAND2_X2 _AES_ENC_us02_U190  ( .A1(_AES_ENC_us02_n1093 ), .A2(_AES_ENC_us02_n587 ), .ZN(_AES_ENC_us02_n876 ) );
NAND2_X2 _AES_ENC_us02_U189  ( .A1(_AES_ENC_us02_n604 ), .A2(_AES_ENC_us02_n876 ), .ZN(_AES_ENC_us02_n877 ) );
NAND2_X2 _AES_ENC_us02_U188  ( .A1(_AES_ENC_us02_n877 ), .A2(_AES_ENC_us02_n623 ), .ZN(_AES_ENC_us02_n888 ) );
NAND4_X2 _AES_ENC_us02_U179  ( .A1(_AES_ENC_us02_n889 ), .A2(_AES_ENC_us02_n888 ), .A3(_AES_ENC_us02_n887 ), .A4(_AES_ENC_us02_n886 ), .ZN(_AES_ENC_us02_n890 ) );
NAND2_X2 _AES_ENC_us02_U178  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n890 ), .ZN(_AES_ENC_us02_n903 ) );
OR2_X2 _AES_ENC_us02_U177  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n1059 ), .ZN(_AES_ENC_us02_n900 ) );
NAND2_X2 _AES_ENC_us02_U176  ( .A1(_AES_ENC_us02_n1073 ), .A2(_AES_ENC_us02_n1047 ), .ZN(_AES_ENC_us02_n899 ) );
NAND2_X2 _AES_ENC_us02_U175  ( .A1(_AES_ENC_us02_n1094 ), .A2(_AES_ENC_us02_n595 ), .ZN(_AES_ENC_us02_n898 ) );
NAND4_X2 _AES_ENC_us02_U167  ( .A1(_AES_ENC_us02_n900 ), .A2(_AES_ENC_us02_n899 ), .A3(_AES_ENC_us02_n898 ), .A4(_AES_ENC_us02_n897 ), .ZN(_AES_ENC_us02_n901 ) );
NAND2_X2 _AES_ENC_us02_U166  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n901 ), .ZN(_AES_ENC_us02_n902 ) );
NAND4_X2 _AES_ENC_us02_U165  ( .A1(_AES_ENC_us02_n905 ), .A2(_AES_ENC_us02_n904 ), .A3(_AES_ENC_us02_n903 ), .A4(_AES_ENC_us02_n902 ), .ZN(_AES_ENC_sa02_sub[4] ) );
NAND2_X2 _AES_ENC_us02_U164  ( .A1(_AES_ENC_us02_n1094 ), .A2(_AES_ENC_us02_n599 ), .ZN(_AES_ENC_us02_n922 ) );
NAND2_X2 _AES_ENC_us02_U163  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n989 ), .ZN(_AES_ENC_us02_n921 ) );
NAND4_X2 _AES_ENC_us02_U151  ( .A1(_AES_ENC_us02_n922 ), .A2(_AES_ENC_us02_n921 ), .A3(_AES_ENC_us02_n920 ), .A4(_AES_ENC_us02_n919 ), .ZN(_AES_ENC_us02_n923 ) );
NAND2_X2 _AES_ENC_us02_U150  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n923 ), .ZN(_AES_ENC_us02_n972 ) );
NAND2_X2 _AES_ENC_us02_U149  ( .A1(_AES_ENC_us02_n582 ), .A2(_AES_ENC_us02_n619 ), .ZN(_AES_ENC_us02_n924 ) );
NAND2_X2 _AES_ENC_us02_U148  ( .A1(_AES_ENC_us02_n1073 ), .A2(_AES_ENC_us02_n924 ), .ZN(_AES_ENC_us02_n939 ) );
NAND2_X2 _AES_ENC_us02_U147  ( .A1(_AES_ENC_us02_n926 ), .A2(_AES_ENC_us02_n925 ), .ZN(_AES_ENC_us02_n927 ) );
NAND2_X2 _AES_ENC_us02_U146  ( .A1(_AES_ENC_us02_n606 ), .A2(_AES_ENC_us02_n927 ), .ZN(_AES_ENC_us02_n928 ) );
NAND2_X2 _AES_ENC_us02_U145  ( .A1(_AES_ENC_us02_n928 ), .A2(_AES_ENC_us02_n1080 ), .ZN(_AES_ENC_us02_n938 ) );
OR2_X2 _AES_ENC_us02_U144  ( .A1(_AES_ENC_us02_n1117 ), .A2(_AES_ENC_us02_n615 ), .ZN(_AES_ENC_us02_n937 ) );
NAND4_X2 _AES_ENC_us02_U139  ( .A1(_AES_ENC_us02_n939 ), .A2(_AES_ENC_us02_n938 ), .A3(_AES_ENC_us02_n937 ), .A4(_AES_ENC_us02_n936 ), .ZN(_AES_ENC_us02_n940 ) );
NAND2_X2 _AES_ENC_us02_U138  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n940 ), .ZN(_AES_ENC_us02_n971 ) );
OR2_X2 _AES_ENC_us02_U137  ( .A1(_AES_ENC_us02_n605 ), .A2(_AES_ENC_us02_n941 ), .ZN(_AES_ENC_us02_n954 ) );
NAND2_X2 _AES_ENC_us02_U136  ( .A1(_AES_ENC_us02_n1096 ), .A2(_AES_ENC_us02_n577 ), .ZN(_AES_ENC_us02_n942 ) );
NAND2_X2 _AES_ENC_us02_U135  ( .A1(_AES_ENC_us02_n1048 ), .A2(_AES_ENC_us02_n942 ), .ZN(_AES_ENC_us02_n943 ) );
NAND2_X2 _AES_ENC_us02_U134  ( .A1(_AES_ENC_us02_n612 ), .A2(_AES_ENC_us02_n943 ), .ZN(_AES_ENC_us02_n944 ) );
NAND2_X2 _AES_ENC_us02_U133  ( .A1(_AES_ENC_us02_n944 ), .A2(_AES_ENC_us02_n580 ), .ZN(_AES_ENC_us02_n953 ) );
NAND4_X2 _AES_ENC_us02_U125  ( .A1(_AES_ENC_us02_n954 ), .A2(_AES_ENC_us02_n953 ), .A3(_AES_ENC_us02_n952 ), .A4(_AES_ENC_us02_n951 ), .ZN(_AES_ENC_us02_n955 ) );
NAND2_X2 _AES_ENC_us02_U124  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n955 ), .ZN(_AES_ENC_us02_n970 ) );
NAND2_X2 _AES_ENC_us02_U123  ( .A1(_AES_ENC_us02_n1094 ), .A2(_AES_ENC_us02_n1071 ), .ZN(_AES_ENC_us02_n967 ) );
NAND2_X2 _AES_ENC_us02_U122  ( .A1(_AES_ENC_us02_n956 ), .A2(_AES_ENC_us02_n1030 ), .ZN(_AES_ENC_us02_n966 ) );
NAND4_X2 _AES_ENC_us02_U114  ( .A1(_AES_ENC_us02_n967 ), .A2(_AES_ENC_us02_n966 ), .A3(_AES_ENC_us02_n965 ), .A4(_AES_ENC_us02_n964 ), .ZN(_AES_ENC_us02_n968 ) );
NAND2_X2 _AES_ENC_us02_U113  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n968 ), .ZN(_AES_ENC_us02_n969 ) );
NAND4_X2 _AES_ENC_us02_U112  ( .A1(_AES_ENC_us02_n972 ), .A2(_AES_ENC_us02_n971 ), .A3(_AES_ENC_us02_n970 ), .A4(_AES_ENC_us02_n969 ), .ZN(_AES_ENC_sa02_sub[5] ) );
NAND2_X2 _AES_ENC_us02_U111  ( .A1(_AES_ENC_us02_n570 ), .A2(_AES_ENC_us02_n1097 ), .ZN(_AES_ENC_us02_n973 ) );
NAND2_X2 _AES_ENC_us02_U110  ( .A1(_AES_ENC_us02_n1073 ), .A2(_AES_ENC_us02_n973 ), .ZN(_AES_ENC_us02_n987 ) );
NAND2_X2 _AES_ENC_us02_U109  ( .A1(_AES_ENC_us02_n974 ), .A2(_AES_ENC_us02_n1077 ), .ZN(_AES_ENC_us02_n975 ) );
NAND2_X2 _AES_ENC_us02_U108  ( .A1(_AES_ENC_us02_n613 ), .A2(_AES_ENC_us02_n975 ), .ZN(_AES_ENC_us02_n976 ) );
NAND2_X2 _AES_ENC_us02_U107  ( .A1(_AES_ENC_us02_n977 ), .A2(_AES_ENC_us02_n976 ), .ZN(_AES_ENC_us02_n986 ) );
NAND4_X2 _AES_ENC_us02_U99  ( .A1(_AES_ENC_us02_n987 ), .A2(_AES_ENC_us02_n986 ), .A3(_AES_ENC_us02_n985 ), .A4(_AES_ENC_us02_n984 ), .ZN(_AES_ENC_us02_n988 ) );
NAND2_X2 _AES_ENC_us02_U98  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n988 ), .ZN(_AES_ENC_us02_n1044 ) );
NAND2_X2 _AES_ENC_us02_U97  ( .A1(_AES_ENC_us02_n1073 ), .A2(_AES_ENC_us02_n989 ), .ZN(_AES_ENC_us02_n1004 ) );
NAND2_X2 _AES_ENC_us02_U96  ( .A1(_AES_ENC_us02_n1092 ), .A2(_AES_ENC_us02_n619 ), .ZN(_AES_ENC_us02_n1003 ) );
NAND4_X2 _AES_ENC_us02_U85  ( .A1(_AES_ENC_us02_n1004 ), .A2(_AES_ENC_us02_n1003 ), .A3(_AES_ENC_us02_n1002 ), .A4(_AES_ENC_us02_n1001 ), .ZN(_AES_ENC_us02_n1005 ) );
NAND2_X2 _AES_ENC_us02_U84  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n1005 ), .ZN(_AES_ENC_us02_n1043 ) );
NAND2_X2 _AES_ENC_us02_U83  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n596 ), .ZN(_AES_ENC_us02_n1020 ) );
NAND2_X2 _AES_ENC_us02_U82  ( .A1(_AES_ENC_us02_n1050 ), .A2(_AES_ENC_us02_n624 ), .ZN(_AES_ENC_us02_n1019 ) );
NAND2_X2 _AES_ENC_us02_U77  ( .A1(_AES_ENC_us02_n1059 ), .A2(_AES_ENC_us02_n1114 ), .ZN(_AES_ENC_us02_n1012 ) );
NAND2_X2 _AES_ENC_us02_U76  ( .A1(_AES_ENC_us02_n1010 ), .A2(_AES_ENC_us02_n592 ), .ZN(_AES_ENC_us02_n1011 ) );
NAND2_X2 _AES_ENC_us02_U75  ( .A1(_AES_ENC_us02_n1012 ), .A2(_AES_ENC_us02_n1011 ), .ZN(_AES_ENC_us02_n1016 ) );
NAND4_X2 _AES_ENC_us02_U70  ( .A1(_AES_ENC_us02_n1020 ), .A2(_AES_ENC_us02_n1019 ), .A3(_AES_ENC_us02_n1018 ), .A4(_AES_ENC_us02_n1017 ), .ZN(_AES_ENC_us02_n1021 ) );
NAND2_X2 _AES_ENC_us02_U69  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n1021 ), .ZN(_AES_ENC_us02_n1042 ) );
NAND2_X2 _AES_ENC_us02_U68  ( .A1(_AES_ENC_us02_n1022 ), .A2(_AES_ENC_us02_n1093 ), .ZN(_AES_ENC_us02_n1039 ) );
NAND2_X2 _AES_ENC_us02_U67  ( .A1(_AES_ENC_us02_n1050 ), .A2(_AES_ENC_us02_n1023 ), .ZN(_AES_ENC_us02_n1038 ) );
NAND2_X2 _AES_ENC_us02_U66  ( .A1(_AES_ENC_us02_n1024 ), .A2(_AES_ENC_us02_n1071 ), .ZN(_AES_ENC_us02_n1037 ) );
AND2_X2 _AES_ENC_us02_U60  ( .A1(_AES_ENC_us02_n1030 ), .A2(_AES_ENC_us02_n602 ), .ZN(_AES_ENC_us02_n1078 ) );
NAND4_X2 _AES_ENC_us02_U56  ( .A1(_AES_ENC_us02_n1039 ), .A2(_AES_ENC_us02_n1038 ), .A3(_AES_ENC_us02_n1037 ), .A4(_AES_ENC_us02_n1036 ), .ZN(_AES_ENC_us02_n1040 ) );
NAND2_X2 _AES_ENC_us02_U55  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n1040 ), .ZN(_AES_ENC_us02_n1041 ) );
NAND4_X2 _AES_ENC_us02_U54  ( .A1(_AES_ENC_us02_n1044 ), .A2(_AES_ENC_us02_n1043 ), .A3(_AES_ENC_us02_n1042 ), .A4(_AES_ENC_us02_n1041 ), .ZN(_AES_ENC_sa02_sub[6] ) );
NAND2_X2 _AES_ENC_us02_U53  ( .A1(_AES_ENC_us02_n1072 ), .A2(_AES_ENC_us02_n1045 ), .ZN(_AES_ENC_us02_n1068 ) );
NAND2_X2 _AES_ENC_us02_U52  ( .A1(_AES_ENC_us02_n1046 ), .A2(_AES_ENC_us02_n582 ), .ZN(_AES_ENC_us02_n1067 ) );
NAND2_X2 _AES_ENC_us02_U51  ( .A1(_AES_ENC_us02_n1094 ), .A2(_AES_ENC_us02_n1047 ), .ZN(_AES_ENC_us02_n1066 ) );
NAND4_X2 _AES_ENC_us02_U40  ( .A1(_AES_ENC_us02_n1068 ), .A2(_AES_ENC_us02_n1067 ), .A3(_AES_ENC_us02_n1066 ), .A4(_AES_ENC_us02_n1065 ), .ZN(_AES_ENC_us02_n1069 ) );
NAND2_X2 _AES_ENC_us02_U39  ( .A1(_AES_ENC_us02_n1070 ), .A2(_AES_ENC_us02_n1069 ), .ZN(_AES_ENC_us02_n1135 ) );
NAND2_X2 _AES_ENC_us02_U38  ( .A1(_AES_ENC_us02_n1072 ), .A2(_AES_ENC_us02_n1071 ), .ZN(_AES_ENC_us02_n1088 ) );
NAND2_X2 _AES_ENC_us02_U37  ( .A1(_AES_ENC_us02_n1073 ), .A2(_AES_ENC_us02_n595 ), .ZN(_AES_ENC_us02_n1087 ) );
NAND4_X2 _AES_ENC_us02_U28  ( .A1(_AES_ENC_us02_n1088 ), .A2(_AES_ENC_us02_n1087 ), .A3(_AES_ENC_us02_n1086 ), .A4(_AES_ENC_us02_n1085 ), .ZN(_AES_ENC_us02_n1089 ) );
NAND2_X2 _AES_ENC_us02_U27  ( .A1(_AES_ENC_us02_n1090 ), .A2(_AES_ENC_us02_n1089 ), .ZN(_AES_ENC_us02_n1134 ) );
NAND2_X2 _AES_ENC_us02_U26  ( .A1(_AES_ENC_us02_n1091 ), .A2(_AES_ENC_us02_n1093 ), .ZN(_AES_ENC_us02_n1111 ) );
NAND2_X2 _AES_ENC_us02_U25  ( .A1(_AES_ENC_us02_n1092 ), .A2(_AES_ENC_us02_n1120 ), .ZN(_AES_ENC_us02_n1110 ) );
AND2_X2 _AES_ENC_us02_U22  ( .A1(_AES_ENC_us02_n1097 ), .A2(_AES_ENC_us02_n1096 ), .ZN(_AES_ENC_us02_n1098 ) );
NAND4_X2 _AES_ENC_us02_U14  ( .A1(_AES_ENC_us02_n1111 ), .A2(_AES_ENC_us02_n1110 ), .A3(_AES_ENC_us02_n1109 ), .A4(_AES_ENC_us02_n1108 ), .ZN(_AES_ENC_us02_n1112 ) );
NAND2_X2 _AES_ENC_us02_U13  ( .A1(_AES_ENC_us02_n1113 ), .A2(_AES_ENC_us02_n1112 ), .ZN(_AES_ENC_us02_n1133 ) );
NAND2_X2 _AES_ENC_us02_U12  ( .A1(_AES_ENC_us02_n1115 ), .A2(_AES_ENC_us02_n1114 ), .ZN(_AES_ENC_us02_n1129 ) );
OR2_X2 _AES_ENC_us02_U11  ( .A1(_AES_ENC_us02_n608 ), .A2(_AES_ENC_us02_n1116 ), .ZN(_AES_ENC_us02_n1128 ) );
NAND4_X2 _AES_ENC_us02_U3  ( .A1(_AES_ENC_us02_n1129 ), .A2(_AES_ENC_us02_n1128 ), .A3(_AES_ENC_us02_n1127 ), .A4(_AES_ENC_us02_n1126 ), .ZN(_AES_ENC_us02_n1130 ) );
NAND2_X2 _AES_ENC_us02_U2  ( .A1(_AES_ENC_us02_n1131 ), .A2(_AES_ENC_us02_n1130 ), .ZN(_AES_ENC_us02_n1132 ) );
NAND4_X2 _AES_ENC_us02_U1  ( .A1(_AES_ENC_us02_n1135 ), .A2(_AES_ENC_us02_n1134 ), .A3(_AES_ENC_us02_n1133 ), .A4(_AES_ENC_us02_n1132 ), .ZN(_AES_ENC_sa02_sub[7] ) );
INV_X4 _AES_ENC_us03_U575  ( .A(_AES_ENC_sa03[4]), .ZN(_AES_ENC_us03_n626 ));
INV_X4 _AES_ENC_us03_U574  ( .A(_AES_ENC_us03_n1025 ), .ZN(_AES_ENC_us03_n624 ) );
INV_X4 _AES_ENC_us03_U573  ( .A(_AES_ENC_us03_n1120 ), .ZN(_AES_ENC_us03_n622 ) );
INV_X4 _AES_ENC_us03_U572  ( .A(_AES_ENC_us03_n1121 ), .ZN(_AES_ENC_us03_n621 ) );
INV_X4 _AES_ENC_us03_U571  ( .A(_AES_ENC_us03_n1048 ), .ZN(_AES_ENC_us03_n620 ) );
INV_X4 _AES_ENC_us03_U570  ( .A(_AES_ENC_us03_n974 ), .ZN(_AES_ENC_us03_n619 ) );
INV_X4 _AES_ENC_us03_U569  ( .A(_AES_ENC_sa03[2]), .ZN(_AES_ENC_us03_n618 ));
INV_X4 _AES_ENC_us03_U568  ( .A(_AES_ENC_us03_n800 ), .ZN(_AES_ENC_us03_n617 ) );
INV_X4 _AES_ENC_us03_U567  ( .A(_AES_ENC_us03_n925 ), .ZN(_AES_ENC_us03_n616 ) );
INV_X4 _AES_ENC_us03_U566  ( .A(_AES_ENC_us03_n1022 ), .ZN(_AES_ENC_us03_n615 ) );
INV_X4 _AES_ENC_us03_U565  ( .A(_AES_ENC_us03_n1102 ), .ZN(_AES_ENC_us03_n614 ) );
INV_X4 _AES_ENC_us03_U564  ( .A(_AES_ENC_us03_n929 ), .ZN(_AES_ENC_us03_n613 ) );
INV_X4 _AES_ENC_us03_U563  ( .A(_AES_ENC_us03_n1056 ), .ZN(_AES_ENC_us03_n612 ) );
INV_X4 _AES_ENC_us03_U562  ( .A(_AES_ENC_us03_n1054 ), .ZN(_AES_ENC_us03_n611 ) );
INV_X4 _AES_ENC_us03_U561  ( .A(_AES_ENC_us03_n881 ), .ZN(_AES_ENC_us03_n610 ) );
INV_X4 _AES_ENC_us03_U560  ( .A(_AES_ENC_us03_n926 ), .ZN(_AES_ENC_us03_n609 ) );
INV_X4 _AES_ENC_us03_U559  ( .A(_AES_ENC_us03_n977 ), .ZN(_AES_ENC_us03_n607 ) );
INV_X4 _AES_ENC_us03_U558  ( .A(_AES_ENC_us03_n1031 ), .ZN(_AES_ENC_us03_n606 ) );
INV_X4 _AES_ENC_us03_U557  ( .A(_AES_ENC_us03_n1103 ), .ZN(_AES_ENC_us03_n605 ) );
INV_X4 _AES_ENC_us03_U556  ( .A(_AES_ENC_us03_n1009 ), .ZN(_AES_ENC_us03_n604 ) );
INV_X4 _AES_ENC_us03_U555  ( .A(_AES_ENC_us03_n990 ), .ZN(_AES_ENC_us03_n603 ) );
INV_X4 _AES_ENC_us03_U554  ( .A(_AES_ENC_us03_n1058 ), .ZN(_AES_ENC_us03_n602 ) );
INV_X4 _AES_ENC_us03_U553  ( .A(_AES_ENC_us03_n1074 ), .ZN(_AES_ENC_us03_n601 ) );
INV_X4 _AES_ENC_us03_U552  ( .A(_AES_ENC_us03_n1053 ), .ZN(_AES_ENC_us03_n600 ) );
INV_X4 _AES_ENC_us03_U551  ( .A(_AES_ENC_us03_n826 ), .ZN(_AES_ENC_us03_n599 ) );
INV_X4 _AES_ENC_us03_U550  ( .A(_AES_ENC_us03_n821 ), .ZN(_AES_ENC_us03_n598 ) );
INV_X4 _AES_ENC_us03_U549  ( .A(_AES_ENC_us03_n910 ), .ZN(_AES_ENC_us03_n597 ) );
INV_X4 _AES_ENC_us03_U548  ( .A(_AES_ENC_us03_n906 ), .ZN(_AES_ENC_us03_n596 ) );
INV_X4 _AES_ENC_us03_U547  ( .A(_AES_ENC_us03_n1013 ), .ZN(_AES_ENC_us03_n594 ) );
INV_X4 _AES_ENC_us03_U546  ( .A(_AES_ENC_us03_n824 ), .ZN(_AES_ENC_us03_n593 ) );
INV_X4 _AES_ENC_us03_U545  ( .A(_AES_ENC_us03_n1091 ), .ZN(_AES_ENC_us03_n592 ) );
INV_X4 _AES_ENC_us03_U544  ( .A(_AES_ENC_us03_n1080 ), .ZN(_AES_ENC_us03_n591 ) );
INV_X4 _AES_ENC_us03_U543  ( .A(_AES_ENC_us03_n959 ), .ZN(_AES_ENC_us03_n590 ) );
INV_X4 _AES_ENC_us03_U542  ( .A(_AES_ENC_us03_n779 ), .ZN(_AES_ENC_us03_n589 ) );
INV_X4 _AES_ENC_us03_U541  ( .A(_AES_ENC_us03_n794 ), .ZN(_AES_ENC_us03_n586 ) );
INV_X4 _AES_ENC_us03_U540  ( .A(_AES_ENC_us03_n880 ), .ZN(_AES_ENC_us03_n584 ) );
INV_X4 _AES_ENC_us03_U539  ( .A(_AES_ENC_sa03[7]), .ZN(_AES_ENC_us03_n582 ));
INV_X4 _AES_ENC_us03_U538  ( .A(_AES_ENC_us03_n992 ), .ZN(_AES_ENC_us03_n579 ) );
INV_X4 _AES_ENC_us03_U537  ( .A(_AES_ENC_us03_n1114 ), .ZN(_AES_ENC_us03_n578 ) );
INV_X4 _AES_ENC_us03_U536  ( .A(_AES_ENC_us03_n1092 ), .ZN(_AES_ENC_us03_n575 ) );
INV_X4 _AES_ENC_us03_U535  ( .A(_AES_ENC_sa03[0]), .ZN(_AES_ENC_us03_n574 ));
NOR2_X2 _AES_ENC_us03_U534  ( .A1(_AES_ENC_sa03[0]), .A2(_AES_ENC_sa03[6]),.ZN(_AES_ENC_us03_n1090 ) );
NOR2_X2 _AES_ENC_us03_U533  ( .A1(_AES_ENC_us03_n574 ), .A2(_AES_ENC_sa03[6]), .ZN(_AES_ENC_us03_n1070 ) );
NOR2_X2 _AES_ENC_us03_U532  ( .A1(_AES_ENC_sa03[4]), .A2(_AES_ENC_sa03[3]),.ZN(_AES_ENC_us03_n1025 ) );
INV_X4 _AES_ENC_us03_U531  ( .A(_AES_ENC_us03_n569 ), .ZN(_AES_ENC_us03_n572 ) );
NOR2_X2 _AES_ENC_us03_U530  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n765 ) );
NOR2_X2 _AES_ENC_us03_U529  ( .A1(_AES_ENC_sa03[4]), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n764 ) );
NOR2_X2 _AES_ENC_us03_U528  ( .A1(_AES_ENC_us03_n765 ), .A2(_AES_ENC_us03_n764 ), .ZN(_AES_ENC_us03_n766 ) );
NOR2_X2 _AES_ENC_us03_U527  ( .A1(_AES_ENC_us03_n766 ), .A2(_AES_ENC_us03_n590 ), .ZN(_AES_ENC_us03_n767 ) );
NOR3_X2 _AES_ENC_us03_U526  ( .A1(_AES_ENC_us03_n582 ), .A2(_AES_ENC_sa03[5]), .A3(_AES_ENC_us03_n704 ), .ZN(_AES_ENC_us03_n706 ));
NOR2_X2 _AES_ENC_us03_U525  ( .A1(_AES_ENC_us03_n1117 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n707 ) );
NOR2_X2 _AES_ENC_us03_U524  ( .A1(_AES_ENC_sa03[4]), .A2(_AES_ENC_us03_n575 ), .ZN(_AES_ENC_us03_n705 ) );
NOR3_X2 _AES_ENC_us03_U523  ( .A1(_AES_ENC_us03_n707 ), .A2(_AES_ENC_us03_n706 ), .A3(_AES_ENC_us03_n705 ), .ZN(_AES_ENC_us03_n713 ) );
INV_X4 _AES_ENC_us03_U522  ( .A(_AES_ENC_sa03[3]), .ZN(_AES_ENC_us03_n623 ));
NAND3_X2 _AES_ENC_us03_U521  ( .A1(_AES_ENC_us03_n652 ), .A2(_AES_ENC_us03_n627 ), .A3(_AES_ENC_sa03[7]), .ZN(_AES_ENC_us03_n653 ));
NOR2_X2 _AES_ENC_us03_U520  ( .A1(_AES_ENC_us03_n618 ), .A2(_AES_ENC_sa03[5]), .ZN(_AES_ENC_us03_n925 ) );
NOR2_X2 _AES_ENC_us03_U519  ( .A1(_AES_ENC_sa03[5]), .A2(_AES_ENC_sa03[2]),.ZN(_AES_ENC_us03_n974 ) );
INV_X4 _AES_ENC_us03_U518  ( .A(_AES_ENC_sa03[5]), .ZN(_AES_ENC_us03_n627 ));
NOR2_X2 _AES_ENC_us03_U517  ( .A1(_AES_ENC_us03_n618 ), .A2(_AES_ENC_sa03[7]), .ZN(_AES_ENC_us03_n779 ) );
NAND3_X2 _AES_ENC_us03_U516  ( .A1(_AES_ENC_us03_n679 ), .A2(_AES_ENC_us03_n678 ), .A3(_AES_ENC_us03_n677 ), .ZN(_AES_ENC_sa03_sub[0] ) );
NOR2_X2 _AES_ENC_us03_U515  ( .A1(_AES_ENC_us03_n627 ), .A2(_AES_ENC_sa03[2]), .ZN(_AES_ENC_us03_n1048 ) );
NOR4_X2 _AES_ENC_us03_U512  ( .A1(_AES_ENC_us03_n633 ), .A2(_AES_ENC_us03_n632 ), .A3(_AES_ENC_us03_n631 ), .A4(_AES_ENC_us03_n630 ), .ZN(_AES_ENC_us03_n634 ) );
NOR2_X2 _AES_ENC_us03_U510  ( .A1(_AES_ENC_us03_n629 ), .A2(_AES_ENC_us03_n628 ), .ZN(_AES_ENC_us03_n635 ) );
NAND3_X2 _AES_ENC_us03_U509  ( .A1(_AES_ENC_sa03[2]), .A2(_AES_ENC_sa03[7]), .A3(_AES_ENC_us03_n1059 ), .ZN(_AES_ENC_us03_n636 ) );
NOR2_X2 _AES_ENC_us03_U508  ( .A1(_AES_ENC_sa03[7]), .A2(_AES_ENC_sa03[2]),.ZN(_AES_ENC_us03_n794 ) );
NOR2_X2 _AES_ENC_us03_U507  ( .A1(_AES_ENC_sa03[4]), .A2(_AES_ENC_sa03[1]),.ZN(_AES_ENC_us03_n1102 ) );
NOR2_X2 _AES_ENC_us03_U506  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_sa03[3]), .ZN(_AES_ENC_us03_n1053 ) );
NOR2_X2 _AES_ENC_us03_U505  ( .A1(_AES_ENC_us03_n589 ), .A2(_AES_ENC_sa03[5]), .ZN(_AES_ENC_us03_n1024 ) );
NOR2_X2 _AES_ENC_us03_U504  ( .A1(_AES_ENC_us03_n578 ), .A2(_AES_ENC_sa03[2]), .ZN(_AES_ENC_us03_n1093 ) );
NOR2_X2 _AES_ENC_us03_U503  ( .A1(_AES_ENC_us03_n586 ), .A2(_AES_ENC_sa03[5]), .ZN(_AES_ENC_us03_n1094 ) );
NOR2_X2 _AES_ENC_us03_U502  ( .A1(_AES_ENC_us03_n626 ), .A2(_AES_ENC_sa03[3]), .ZN(_AES_ENC_us03_n931 ) );
INV_X4 _AES_ENC_us03_U501  ( .A(_AES_ENC_us03_n570 ), .ZN(_AES_ENC_us03_n573 ) );
NOR2_X2 _AES_ENC_us03_U500  ( .A1(_AES_ENC_us03_n1053 ), .A2(_AES_ENC_us03_n1095 ), .ZN(_AES_ENC_us03_n639 ) );
NOR3_X2 _AES_ENC_us03_U499  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n573 ), .A3(_AES_ENC_us03_n1074 ), .ZN(_AES_ENC_us03_n641 ) );
NOR2_X2 _AES_ENC_us03_U498  ( .A1(_AES_ENC_us03_n639 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n640 ) );
NOR2_X2 _AES_ENC_us03_U497  ( .A1(_AES_ENC_us03_n641 ), .A2(_AES_ENC_us03_n640 ), .ZN(_AES_ENC_us03_n646 ) );
NOR3_X2 _AES_ENC_us03_U496  ( .A1(_AES_ENC_us03_n995 ), .A2(_AES_ENC_us03_n579 ), .A3(_AES_ENC_us03_n994 ), .ZN(_AES_ENC_us03_n1002 ) );
NOR2_X2 _AES_ENC_us03_U495  ( .A1(_AES_ENC_us03_n909 ), .A2(_AES_ENC_us03_n908 ), .ZN(_AES_ENC_us03_n920 ) );
NOR2_X2 _AES_ENC_us03_U494  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n823 ) );
NOR2_X2 _AES_ENC_us03_U492  ( .A1(_AES_ENC_us03_n626 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n822 ) );
NOR2_X2 _AES_ENC_us03_U491  ( .A1(_AES_ENC_us03_n823 ), .A2(_AES_ENC_us03_n822 ), .ZN(_AES_ENC_us03_n825 ) );
NOR2_X2 _AES_ENC_us03_U490  ( .A1(_AES_ENC_sa03[1]), .A2(_AES_ENC_us03_n625 ), .ZN(_AES_ENC_us03_n913 ) );
NOR2_X2 _AES_ENC_us03_U489  ( .A1(_AES_ENC_us03_n913 ), .A2(_AES_ENC_us03_n1091 ), .ZN(_AES_ENC_us03_n914 ) );
NOR2_X2 _AES_ENC_us03_U488  ( .A1(_AES_ENC_us03_n826 ), .A2(_AES_ENC_us03_n572 ), .ZN(_AES_ENC_us03_n827 ) );
NOR3_X2 _AES_ENC_us03_U487  ( .A1(_AES_ENC_us03_n769 ), .A2(_AES_ENC_us03_n768 ), .A3(_AES_ENC_us03_n767 ), .ZN(_AES_ENC_us03_n775 ) );
NOR2_X2 _AES_ENC_us03_U486  ( .A1(_AES_ENC_us03_n1056 ), .A2(_AES_ENC_us03_n1053 ), .ZN(_AES_ENC_us03_n749 ) );
NOR2_X2 _AES_ENC_us03_U483  ( .A1(_AES_ENC_us03_n749 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n752 ) );
INV_X4 _AES_ENC_us03_U482  ( .A(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n608 ));
NOR2_X2 _AES_ENC_us03_U480  ( .A1(_AES_ENC_us03_n1054 ), .A2(_AES_ENC_us03_n1053 ), .ZN(_AES_ENC_us03_n1055 ) );
OR2_X4 _AES_ENC_us03_U479  ( .A1(_AES_ENC_us03_n1094 ), .A2(_AES_ENC_us03_n1093 ), .ZN(_AES_ENC_us03_n571 ) );
AND2_X2 _AES_ENC_us03_U478  ( .A1(_AES_ENC_us03_n571 ), .A2(_AES_ENC_us03_n1095 ), .ZN(_AES_ENC_us03_n1101 ) );
NOR2_X2 _AES_ENC_us03_U477  ( .A1(_AES_ENC_us03_n1074 ), .A2(_AES_ENC_us03_n931 ), .ZN(_AES_ENC_us03_n796 ) );
NOR2_X2 _AES_ENC_us03_U474  ( .A1(_AES_ENC_us03_n796 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n797 ) );
NOR2_X2 _AES_ENC_us03_U473  ( .A1(_AES_ENC_us03_n932 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n933 ) );
NOR2_X2 _AES_ENC_us03_U472  ( .A1(_AES_ENC_us03_n929 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n935 ) );
NOR2_X2 _AES_ENC_us03_U471  ( .A1(_AES_ENC_us03_n931 ), .A2(_AES_ENC_us03_n930 ), .ZN(_AES_ENC_us03_n934 ) );
NOR3_X2 _AES_ENC_us03_U470  ( .A1(_AES_ENC_us03_n935 ), .A2(_AES_ENC_us03_n934 ), .A3(_AES_ENC_us03_n933 ), .ZN(_AES_ENC_us03_n936 ) );
NOR2_X2 _AES_ENC_us03_U469  ( .A1(_AES_ENC_us03_n626 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n1075 ) );
NOR2_X2 _AES_ENC_us03_U468  ( .A1(_AES_ENC_us03_n572 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n949 ) );
NOR2_X2 _AES_ENC_us03_U467  ( .A1(_AES_ENC_us03_n1049 ), .A2(_AES_ENC_us03_n620 ), .ZN(_AES_ENC_us03_n1051 ) );
NOR2_X2 _AES_ENC_us03_U466  ( .A1(_AES_ENC_us03_n1051 ), .A2(_AES_ENC_us03_n1050 ), .ZN(_AES_ENC_us03_n1052 ) );
NOR2_X2 _AES_ENC_us03_U465  ( .A1(_AES_ENC_us03_n1052 ), .A2(_AES_ENC_us03_n604 ), .ZN(_AES_ENC_us03_n1064 ) );
NOR2_X2 _AES_ENC_us03_U464  ( .A1(_AES_ENC_sa03[1]), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n631 ) );
NOR2_X2 _AES_ENC_us03_U463  ( .A1(_AES_ENC_us03_n1025 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n980 ) );
NOR2_X2 _AES_ENC_us03_U462  ( .A1(_AES_ENC_us03_n1073 ), .A2(_AES_ENC_us03_n1094 ), .ZN(_AES_ENC_us03_n795 ) );
NOR2_X2 _AES_ENC_us03_U461  ( .A1(_AES_ENC_us03_n795 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n799 ) );
NOR2_X2 _AES_ENC_us03_U460  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n981 ) );
NOR2_X2 _AES_ENC_us03_U459  ( .A1(_AES_ENC_us03_n1102 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n643 ) );
NOR2_X2 _AES_ENC_us03_U458  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n623 ), .ZN(_AES_ENC_us03_n642 ) );
NOR2_X2 _AES_ENC_us03_U455  ( .A1(_AES_ENC_us03_n911 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n644 ) );
NOR4_X2 _AES_ENC_us03_U448  ( .A1(_AES_ENC_us03_n644 ), .A2(_AES_ENC_us03_n643 ), .A3(_AES_ENC_us03_n804 ), .A4(_AES_ENC_us03_n642 ), .ZN(_AES_ENC_us03_n645 ) );
NOR2_X2 _AES_ENC_us03_U447  ( .A1(_AES_ENC_us03_n1102 ), .A2(_AES_ENC_us03_n910 ), .ZN(_AES_ENC_us03_n932 ) );
NOR2_X2 _AES_ENC_us03_U442  ( .A1(_AES_ENC_us03_n1102 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n755 ) );
NOR2_X2 _AES_ENC_us03_U441  ( .A1(_AES_ENC_us03_n931 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n743 ) );
NOR2_X2 _AES_ENC_us03_U438  ( .A1(_AES_ENC_us03_n1072 ), .A2(_AES_ENC_us03_n1094 ), .ZN(_AES_ENC_us03_n930 ) );
NOR2_X2 _AES_ENC_us03_U435  ( .A1(_AES_ENC_us03_n1074 ), .A2(_AES_ENC_us03_n1025 ), .ZN(_AES_ENC_us03_n891 ) );
NOR2_X2 _AES_ENC_us03_U434  ( .A1(_AES_ENC_us03_n891 ), .A2(_AES_ENC_us03_n616 ), .ZN(_AES_ENC_us03_n894 ) );
NOR3_X2 _AES_ENC_us03_U433  ( .A1(_AES_ENC_us03_n625 ), .A2(_AES_ENC_sa03[1]), .A3(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n683 ));
INV_X4 _AES_ENC_us03_U428  ( .A(_AES_ENC_us03_n931 ), .ZN(_AES_ENC_us03_n625 ) );
NOR2_X2 _AES_ENC_us03_U427  ( .A1(_AES_ENC_us03_n996 ), .A2(_AES_ENC_us03_n931 ), .ZN(_AES_ENC_us03_n704 ) );
NOR2_X2 _AES_ENC_us03_U421  ( .A1(_AES_ENC_us03_n931 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n685 ) );
NOR2_X2 _AES_ENC_us03_U420  ( .A1(_AES_ENC_us03_n1029 ), .A2(_AES_ENC_us03_n1025 ), .ZN(_AES_ENC_us03_n1079 ) );
NOR3_X2 _AES_ENC_us03_U419  ( .A1(_AES_ENC_us03_n601 ), .A2(_AES_ENC_us03_n1025 ), .A3(_AES_ENC_us03_n619 ), .ZN(_AES_ENC_us03_n945 ) );
NOR2_X2 _AES_ENC_us03_U418  ( .A1(_AES_ENC_us03_n627 ), .A2(_AES_ENC_us03_n618 ), .ZN(_AES_ENC_us03_n800 ) );
NOR3_X2 _AES_ENC_us03_U417  ( .A1(_AES_ENC_us03_n602 ), .A2(_AES_ENC_us03_n582 ), .A3(_AES_ENC_us03_n618 ), .ZN(_AES_ENC_us03_n798 ) );
NOR3_X2 _AES_ENC_us03_U416  ( .A1(_AES_ENC_us03_n617 ), .A2(_AES_ENC_us03_n572 ), .A3(_AES_ENC_us03_n590 ), .ZN(_AES_ENC_us03_n962 ) );
NOR3_X2 _AES_ENC_us03_U415  ( .A1(_AES_ENC_us03_n959 ), .A2(_AES_ENC_us03_n572 ), .A3(_AES_ENC_us03_n616 ), .ZN(_AES_ENC_us03_n768 ) );
NOR3_X2 _AES_ENC_us03_U414  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n572 ), .A3(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n694 ) );
NOR3_X2 _AES_ENC_us03_U413  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n572 ), .A3(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n895 ) );
NOR3_X2 _AES_ENC_us03_U410  ( .A1(_AES_ENC_us03_n1008 ), .A2(_AES_ENC_us03_n1007 ), .A3(_AES_ENC_us03_n1006 ), .ZN(_AES_ENC_us03_n1018 ) );
NOR4_X2 _AES_ENC_us03_U409  ( .A1(_AES_ENC_us03_n711 ), .A2(_AES_ENC_us03_n710 ), .A3(_AES_ENC_us03_n709 ), .A4(_AES_ENC_us03_n708 ), .ZN(_AES_ENC_us03_n712 ) );
NOR4_X2 _AES_ENC_us03_U406  ( .A1(_AES_ENC_us03_n806 ), .A2(_AES_ENC_us03_n805 ), .A3(_AES_ENC_us03_n804 ), .A4(_AES_ENC_us03_n803 ), .ZN(_AES_ENC_us03_n807 ) );
NOR3_X2 _AES_ENC_us03_U405  ( .A1(_AES_ENC_us03_n799 ), .A2(_AES_ENC_us03_n798 ), .A3(_AES_ENC_us03_n797 ), .ZN(_AES_ENC_us03_n808 ) );
NOR2_X2 _AES_ENC_us03_U404  ( .A1(_AES_ENC_us03_n669 ), .A2(_AES_ENC_us03_n668 ), .ZN(_AES_ENC_us03_n673 ) );
NOR4_X2 _AES_ENC_us03_U403  ( .A1(_AES_ENC_us03_n946 ), .A2(_AES_ENC_us03_n1046 ), .A3(_AES_ENC_us03_n671 ), .A4(_AES_ENC_us03_n670 ), .ZN(_AES_ENC_us03_n672 ) );
NOR3_X2 _AES_ENC_us03_U401  ( .A1(_AES_ENC_us03_n1101 ), .A2(_AES_ENC_us03_n1100 ), .A3(_AES_ENC_us03_n1099 ), .ZN(_AES_ENC_us03_n1109 ) );
NOR4_X2 _AES_ENC_us03_U400  ( .A1(_AES_ENC_us03_n843 ), .A2(_AES_ENC_us03_n842 ), .A3(_AES_ENC_us03_n841 ), .A4(_AES_ENC_us03_n840 ), .ZN(_AES_ENC_us03_n844 ) );
NOR4_X2 _AES_ENC_us03_U399  ( .A1(_AES_ENC_us03_n963 ), .A2(_AES_ENC_us03_n962 ), .A3(_AES_ENC_us03_n961 ), .A4(_AES_ENC_us03_n960 ), .ZN(_AES_ENC_us03_n964 ) );
NOR3_X2 _AES_ENC_us03_U398  ( .A1(_AES_ENC_us03_n743 ), .A2(_AES_ENC_us03_n742 ), .A3(_AES_ENC_us03_n741 ), .ZN(_AES_ENC_us03_n744 ) );
NOR2_X2 _AES_ENC_us03_U397  ( .A1(_AES_ENC_us03_n697 ), .A2(_AES_ENC_us03_n658 ), .ZN(_AES_ENC_us03_n659 ) );
NOR2_X2 _AES_ENC_us03_U396  ( .A1(_AES_ENC_us03_n1078 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n1033 ) );
NOR2_X2 _AES_ENC_us03_U393  ( .A1(_AES_ENC_us03_n1031 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n1032 ) );
NOR3_X2 _AES_ENC_us03_U390  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n1025 ), .A3(_AES_ENC_us03_n1074 ), .ZN(_AES_ENC_us03_n1035 ) );
NOR4_X2 _AES_ENC_us03_U389  ( .A1(_AES_ENC_us03_n1035 ), .A2(_AES_ENC_us03_n1034 ), .A3(_AES_ENC_us03_n1033 ), .A4(_AES_ENC_us03_n1032 ), .ZN(_AES_ENC_us03_n1036 ) );
NOR2_X2 _AES_ENC_us03_U388  ( .A1(_AES_ENC_us03_n610 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n885 ) );
NOR2_X2 _AES_ENC_us03_U387  ( .A1(_AES_ENC_us03_n625 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n882 ) );
NOR2_X2 _AES_ENC_us03_U386  ( .A1(_AES_ENC_us03_n1053 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n884 ) );
NOR4_X2 _AES_ENC_us03_U385  ( .A1(_AES_ENC_us03_n885 ), .A2(_AES_ENC_us03_n884 ), .A3(_AES_ENC_us03_n883 ), .A4(_AES_ENC_us03_n882 ), .ZN(_AES_ENC_us03_n886 ) );
NOR2_X2 _AES_ENC_us03_U384  ( .A1(_AES_ENC_us03_n825 ), .A2(_AES_ENC_us03_n593 ), .ZN(_AES_ENC_us03_n830 ) );
NOR2_X2 _AES_ENC_us03_U383  ( .A1(_AES_ENC_us03_n827 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n829 ) );
NOR2_X2 _AES_ENC_us03_U382  ( .A1(_AES_ENC_us03_n572 ), .A2(_AES_ENC_us03_n575 ), .ZN(_AES_ENC_us03_n828 ) );
NOR4_X2 _AES_ENC_us03_U374  ( .A1(_AES_ENC_us03_n831 ), .A2(_AES_ENC_us03_n830 ), .A3(_AES_ENC_us03_n829 ), .A4(_AES_ENC_us03_n828 ), .ZN(_AES_ENC_us03_n832 ) );
NOR2_X2 _AES_ENC_us03_U373  ( .A1(_AES_ENC_us03_n588 ), .A2(_AES_ENC_us03_n595 ), .ZN(_AES_ENC_us03_n1104 ) );
NOR2_X2 _AES_ENC_us03_U372  ( .A1(_AES_ENC_us03_n1102 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n1106 ) );
NOR2_X2 _AES_ENC_us03_U370  ( .A1(_AES_ENC_us03_n1103 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n1105 ) );
NOR4_X2 _AES_ENC_us03_U369  ( .A1(_AES_ENC_us03_n1107 ), .A2(_AES_ENC_us03_n1106 ), .A3(_AES_ENC_us03_n1105 ), .A4(_AES_ENC_us03_n1104 ), .ZN(_AES_ENC_us03_n1108 ) );
NOR3_X2 _AES_ENC_us03_U368  ( .A1(_AES_ENC_us03_n959 ), .A2(_AES_ENC_us03_n623 ), .A3(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n963 ) );
NOR2_X2 _AES_ENC_us03_U367  ( .A1(_AES_ENC_us03_n627 ), .A2(_AES_ENC_us03_n582 ), .ZN(_AES_ENC_us03_n1114 ) );
INV_X4 _AES_ENC_us03_U366  ( .A(_AES_ENC_us03_n1024 ), .ZN(_AES_ENC_us03_n588 ) );
NOR3_X2 _AES_ENC_us03_U365  ( .A1(_AES_ENC_us03_n910 ), .A2(_AES_ENC_us03_n1059 ), .A3(_AES_ENC_us03_n618 ), .ZN(_AES_ENC_us03_n1115 ) );
INV_X4 _AES_ENC_us03_U364  ( .A(_AES_ENC_us03_n1094 ), .ZN(_AES_ENC_us03_n585 ) );
NOR2_X2 _AES_ENC_us03_U363  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n931 ), .ZN(_AES_ENC_us03_n1100 ) );
INV_X4 _AES_ENC_us03_U354  ( .A(_AES_ENC_us03_n1093 ), .ZN(_AES_ENC_us03_n576 ) );
NOR2_X2 _AES_ENC_us03_U353  ( .A1(_AES_ENC_us03_n569 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n929 ) );
NOR2_X2 _AES_ENC_us03_U352  ( .A1(_AES_ENC_us03_n622 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n926 ) );
NOR2_X2 _AES_ENC_us03_U351  ( .A1(_AES_ENC_us03_n572 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n1095 ) );
NOR2_X2 _AES_ENC_us03_U350  ( .A1(_AES_ENC_us03_n616 ), .A2(_AES_ENC_us03_n582 ), .ZN(_AES_ENC_us03_n1010 ) );
NOR2_X2 _AES_ENC_us03_U349  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n1103 ) );
NOR2_X2 _AES_ENC_us03_U348  ( .A1(_AES_ENC_us03_n624 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n1059 ) );
NOR2_X2 _AES_ENC_us03_U347  ( .A1(_AES_ENC_sa03[1]), .A2(_AES_ENC_us03_n1120 ), .ZN(_AES_ENC_us03_n1022 ) );
NOR2_X2 _AES_ENC_us03_U346  ( .A1(_AES_ENC_us03_n621 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n911 ) );
NOR2_X2 _AES_ENC_us03_U345  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_us03_n1025 ), .ZN(_AES_ENC_us03_n826 ) );
NOR2_X2 _AES_ENC_us03_U338  ( .A1(_AES_ENC_us03_n627 ), .A2(_AES_ENC_us03_n589 ), .ZN(_AES_ENC_us03_n1072 ) );
NOR2_X2 _AES_ENC_us03_U335  ( .A1(_AES_ENC_us03_n582 ), .A2(_AES_ENC_us03_n619 ), .ZN(_AES_ENC_us03_n956 ) );
NOR2_X2 _AES_ENC_us03_U329  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_us03_n626 ), .ZN(_AES_ENC_us03_n1121 ) );
NOR2_X2 _AES_ENC_us03_U328  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_us03_n626 ), .ZN(_AES_ENC_us03_n1058 ) );
NOR2_X2 _AES_ENC_us03_U327  ( .A1(_AES_ENC_us03_n578 ), .A2(_AES_ENC_us03_n618 ), .ZN(_AES_ENC_us03_n1073 ) );
NOR2_X2 _AES_ENC_us03_U325  ( .A1(_AES_ENC_sa03[1]), .A2(_AES_ENC_us03_n1025 ), .ZN(_AES_ENC_us03_n1054 ) );
NOR2_X2 _AES_ENC_us03_U324  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_us03_n931 ), .ZN(_AES_ENC_us03_n1029 ) );
NOR2_X2 _AES_ENC_us03_U319  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n1056 ) );
NOR2_X2 _AES_ENC_us03_U318  ( .A1(_AES_ENC_us03_n586 ), .A2(_AES_ENC_us03_n627 ), .ZN(_AES_ENC_us03_n1050 ) );
NOR2_X2 _AES_ENC_us03_U317  ( .A1(_AES_ENC_us03_n1121 ), .A2(_AES_ENC_us03_n1025 ), .ZN(_AES_ENC_us03_n1120 ) );
NOR2_X2 _AES_ENC_us03_U316  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_us03_n572 ), .ZN(_AES_ENC_us03_n1074 ) );
NOR2_X2 _AES_ENC_us03_U315  ( .A1(_AES_ENC_us03_n1058 ), .A2(_AES_ENC_us03_n1054 ), .ZN(_AES_ENC_us03_n878 ) );
NOR2_X2 _AES_ENC_us03_U314  ( .A1(_AES_ENC_us03_n878 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n879 ) );
NOR2_X2 _AES_ENC_us03_U312  ( .A1(_AES_ENC_us03_n880 ), .A2(_AES_ENC_us03_n879 ), .ZN(_AES_ENC_us03_n887 ) );
NOR2_X2 _AES_ENC_us03_U311  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n600 ), .ZN(_AES_ENC_us03_n957 ) );
NOR2_X2 _AES_ENC_us03_U310  ( .A1(_AES_ENC_us03_n958 ), .A2(_AES_ENC_us03_n957 ), .ZN(_AES_ENC_us03_n965 ) );
NOR3_X2 _AES_ENC_us03_U309  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n1091 ), .A3(_AES_ENC_us03_n1022 ), .ZN(_AES_ENC_us03_n720 ) );
NOR3_X2 _AES_ENC_us03_U303  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n1054 ), .A3(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n719 ) );
NOR2_X2 _AES_ENC_us03_U302  ( .A1(_AES_ENC_us03_n720 ), .A2(_AES_ENC_us03_n719 ), .ZN(_AES_ENC_us03_n726 ) );
NOR2_X2 _AES_ENC_us03_U300  ( .A1(_AES_ENC_us03_n586 ), .A2(_AES_ENC_us03_n603 ), .ZN(_AES_ENC_us03_n865 ) );
NOR2_X2 _AES_ENC_us03_U299  ( .A1(_AES_ENC_us03_n1059 ), .A2(_AES_ENC_us03_n1058 ), .ZN(_AES_ENC_us03_n1060 ) );
NOR2_X2 _AES_ENC_us03_U298  ( .A1(_AES_ENC_us03_n1095 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n668 ) );
NOR2_X2 _AES_ENC_us03_U297  ( .A1(_AES_ENC_us03_n911 ), .A2(_AES_ENC_us03_n910 ), .ZN(_AES_ENC_us03_n912 ) );
NOR2_X2 _AES_ENC_us03_U296  ( .A1(_AES_ENC_us03_n912 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n916 ) );
NOR2_X2 _AES_ENC_us03_U295  ( .A1(_AES_ENC_us03_n826 ), .A2(_AES_ENC_us03_n573 ), .ZN(_AES_ENC_us03_n750 ) );
NOR2_X2 _AES_ENC_us03_U294  ( .A1(_AES_ENC_us03_n750 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n751 ) );
NOR2_X2 _AES_ENC_us03_U293  ( .A1(_AES_ENC_us03_n907 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n908 ) );
NOR2_X2 _AES_ENC_us03_U292  ( .A1(_AES_ENC_us03_n990 ), .A2(_AES_ENC_us03_n926 ), .ZN(_AES_ENC_us03_n780 ) );
NOR2_X2 _AES_ENC_us03_U291  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n597 ), .ZN(_AES_ENC_us03_n838 ) );
NOR2_X2 _AES_ENC_us03_U290  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n614 ), .ZN(_AES_ENC_us03_n837 ) );
NOR2_X2 _AES_ENC_us03_U284  ( .A1(_AES_ENC_us03_n838 ), .A2(_AES_ENC_us03_n837 ), .ZN(_AES_ENC_us03_n845 ) );
NOR2_X2 _AES_ENC_us03_U283  ( .A1(_AES_ENC_us03_n1022 ), .A2(_AES_ENC_us03_n1058 ), .ZN(_AES_ENC_us03_n740 ) );
NOR2_X2 _AES_ENC_us03_U282  ( .A1(_AES_ENC_us03_n740 ), .A2(_AES_ENC_us03_n619 ), .ZN(_AES_ENC_us03_n742 ) );
NOR2_X2 _AES_ENC_us03_U281  ( .A1(_AES_ENC_us03_n1098 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n1099 ) );
NOR2_X2 _AES_ENC_us03_U280  ( .A1(_AES_ENC_us03_n1120 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n993 ) );
NOR2_X2 _AES_ENC_us03_U279  ( .A1(_AES_ENC_us03_n993 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n994 ) );
NOR2_X2 _AES_ENC_us03_U273  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n622 ), .ZN(_AES_ENC_us03_n1026 ) );
NOR2_X2 _AES_ENC_us03_U272  ( .A1(_AES_ENC_us03_n573 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n1027 ) );
NOR2_X2 _AES_ENC_us03_U271  ( .A1(_AES_ENC_us03_n1027 ), .A2(_AES_ENC_us03_n1026 ), .ZN(_AES_ENC_us03_n1028 ) );
NOR2_X2 _AES_ENC_us03_U270  ( .A1(_AES_ENC_us03_n1029 ), .A2(_AES_ENC_us03_n1028 ), .ZN(_AES_ENC_us03_n1034 ) );
NOR4_X2 _AES_ENC_us03_U269  ( .A1(_AES_ENC_us03_n757 ), .A2(_AES_ENC_us03_n756 ), .A3(_AES_ENC_us03_n755 ), .A4(_AES_ENC_us03_n754 ), .ZN(_AES_ENC_us03_n758 ) );
NOR2_X2 _AES_ENC_us03_U268  ( .A1(_AES_ENC_us03_n752 ), .A2(_AES_ENC_us03_n751 ), .ZN(_AES_ENC_us03_n759 ) );
NOR2_X2 _AES_ENC_us03_U267  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n1071 ), .ZN(_AES_ENC_us03_n669 ) );
NOR2_X2 _AES_ENC_us03_U263  ( .A1(_AES_ENC_us03_n1056 ), .A2(_AES_ENC_us03_n990 ), .ZN(_AES_ENC_us03_n991 ) );
NOR2_X2 _AES_ENC_us03_U262  ( .A1(_AES_ENC_us03_n991 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n995 ) );
NOR2_X2 _AES_ENC_us03_U258  ( .A1(_AES_ENC_us03_n589 ), .A2(_AES_ENC_us03_n602 ), .ZN(_AES_ENC_us03_n1008 ) );
NOR2_X2 _AES_ENC_us03_U255  ( .A1(_AES_ENC_us03_n839 ), .A2(_AES_ENC_us03_n595 ), .ZN(_AES_ENC_us03_n693 ) );
NOR2_X2 _AES_ENC_us03_U254  ( .A1(_AES_ENC_us03_n588 ), .A2(_AES_ENC_us03_n906 ), .ZN(_AES_ENC_us03_n741 ) );
NOR2_X2 _AES_ENC_us03_U253  ( .A1(_AES_ENC_us03_n1054 ), .A2(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n763 ) );
NOR2_X2 _AES_ENC_us03_U252  ( .A1(_AES_ENC_us03_n763 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n769 ) );
NOR2_X2 _AES_ENC_us03_U251  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n592 ), .ZN(_AES_ENC_us03_n1007 ) );
NOR2_X2 _AES_ENC_us03_U250  ( .A1(_AES_ENC_us03_n616 ), .A2(_AES_ENC_us03_n594 ), .ZN(_AES_ENC_us03_n1123 ) );
NOR2_X2 _AES_ENC_us03_U243  ( .A1(_AES_ENC_us03_n616 ), .A2(_AES_ENC_us03_n602 ), .ZN(_AES_ENC_us03_n710 ) );
INV_X4 _AES_ENC_us03_U242  ( .A(_AES_ENC_us03_n1029 ), .ZN(_AES_ENC_us03_n595 ) );
NOR2_X2 _AES_ENC_us03_U241  ( .A1(_AES_ENC_us03_n619 ), .A2(_AES_ENC_us03_n609 ), .ZN(_AES_ENC_us03_n883 ) );
NOR2_X2 _AES_ENC_us03_U240  ( .A1(_AES_ENC_us03_n605 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n1125 ) );
NOR2_X2 _AES_ENC_us03_U239  ( .A1(_AES_ENC_us03_n990 ), .A2(_AES_ENC_us03_n929 ), .ZN(_AES_ENC_us03_n892 ) );
NOR2_X2 _AES_ENC_us03_U238  ( .A1(_AES_ENC_us03_n892 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n893 ) );
NOR2_X2 _AES_ENC_us03_U237  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n614 ), .ZN(_AES_ENC_us03_n950 ) );
NOR2_X2 _AES_ENC_us03_U236  ( .A1(_AES_ENC_us03_n1079 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n1082 ) );
NOR2_X2 _AES_ENC_us03_U235  ( .A1(_AES_ENC_us03_n910 ), .A2(_AES_ENC_us03_n1056 ), .ZN(_AES_ENC_us03_n941 ) );
NOR2_X2 _AES_ENC_us03_U234  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n1077 ), .ZN(_AES_ENC_us03_n841 ) );
NOR2_X2 _AES_ENC_us03_U229  ( .A1(_AES_ENC_us03_n625 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n630 ) );
NOR2_X2 _AES_ENC_us03_U228  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n614 ), .ZN(_AES_ENC_us03_n806 ) );
NOR2_X2 _AES_ENC_us03_U227  ( .A1(_AES_ENC_us03_n625 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n948 ) );
NOR2_X2 _AES_ENC_us03_U226  ( .A1(_AES_ENC_us03_n588 ), .A2(_AES_ENC_us03_n601 ), .ZN(_AES_ENC_us03_n997 ) );
NOR2_X2 _AES_ENC_us03_U225  ( .A1(_AES_ENC_us03_n1121 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n1122 ) );
NOR2_X2 _AES_ENC_us03_U223  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n1023 ), .ZN(_AES_ENC_us03_n756 ) );
NOR2_X2 _AES_ENC_us03_U222  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n614 ), .ZN(_AES_ENC_us03_n870 ) );
NOR2_X2 _AES_ENC_us03_U221  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n569 ), .ZN(_AES_ENC_us03_n947 ) );
NOR2_X2 _AES_ENC_us03_U217  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n1077 ), .ZN(_AES_ENC_us03_n1084 ) );
NOR2_X2 _AES_ENC_us03_U213  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n855 ), .ZN(_AES_ENC_us03_n709 ) );
NOR2_X2 _AES_ENC_us03_U212  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n601 ), .ZN(_AES_ENC_us03_n868 ) );
NOR2_X2 _AES_ENC_us03_U211  ( .A1(_AES_ENC_us03_n1120 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n1124 ) );
NOR2_X2 _AES_ENC_us03_U210  ( .A1(_AES_ENC_us03_n1120 ), .A2(_AES_ENC_us03_n839 ), .ZN(_AES_ENC_us03_n842 ) );
NOR2_X2 _AES_ENC_us03_U209  ( .A1(_AES_ENC_us03_n1120 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n696 ) );
NOR2_X2 _AES_ENC_us03_U208  ( .A1(_AES_ENC_us03_n1074 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n1076 ) );
NOR2_X2 _AES_ENC_us03_U207  ( .A1(_AES_ENC_us03_n1074 ), .A2(_AES_ENC_us03_n622 ), .ZN(_AES_ENC_us03_n781 ) );
NOR3_X2 _AES_ENC_us03_U201  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n1056 ), .A3(_AES_ENC_us03_n990 ), .ZN(_AES_ENC_us03_n979 ) );
NOR3_X2 _AES_ENC_us03_U200  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n1058 ), .A3(_AES_ENC_us03_n1059 ), .ZN(_AES_ENC_us03_n854 ) );
NOR2_X2 _AES_ENC_us03_U199  ( .A1(_AES_ENC_us03_n996 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n869 ) );
NOR2_X2 _AES_ENC_us03_U198  ( .A1(_AES_ENC_us03_n1056 ), .A2(_AES_ENC_us03_n1074 ), .ZN(_AES_ENC_us03_n1057 ) );
NOR3_X2 _AES_ENC_us03_U197  ( .A1(_AES_ENC_us03_n589 ), .A2(_AES_ENC_us03_n1120 ), .A3(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n978 ) );
NOR2_X2 _AES_ENC_us03_U196  ( .A1(_AES_ENC_us03_n996 ), .A2(_AES_ENC_us03_n911 ), .ZN(_AES_ENC_us03_n1116 ) );
NOR2_X2 _AES_ENC_us03_U195  ( .A1(_AES_ENC_us03_n1074 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n754 ) );
NOR2_X2 _AES_ENC_us03_U194  ( .A1(_AES_ENC_us03_n926 ), .A2(_AES_ENC_us03_n1103 ), .ZN(_AES_ENC_us03_n977 ) );
NOR2_X2 _AES_ENC_us03_U187  ( .A1(_AES_ENC_us03_n839 ), .A2(_AES_ENC_us03_n824 ), .ZN(_AES_ENC_us03_n1092 ) );
NOR2_X2 _AES_ENC_us03_U186  ( .A1(_AES_ENC_us03_n573 ), .A2(_AES_ENC_us03_n1074 ), .ZN(_AES_ENC_us03_n684 ) );
NOR2_X2 _AES_ENC_us03_U185  ( .A1(_AES_ENC_us03_n826 ), .A2(_AES_ENC_us03_n1059 ), .ZN(_AES_ENC_us03_n907 ) );
NOR3_X2 _AES_ENC_us03_U184  ( .A1(_AES_ENC_us03_n578 ), .A2(_AES_ENC_us03_n1115 ), .A3(_AES_ENC_us03_n598 ), .ZN(_AES_ENC_us03_n831 ) );
NOR3_X2 _AES_ENC_us03_U183  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n1056 ), .A3(_AES_ENC_us03_n990 ), .ZN(_AES_ENC_us03_n896 ) );
NOR3_X2 _AES_ENC_us03_U182  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n573 ), .A3(_AES_ENC_us03_n1013 ), .ZN(_AES_ENC_us03_n670 ) );
NOR3_X2 _AES_ENC_us03_U181  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n1091 ), .A3(_AES_ENC_us03_n1022 ), .ZN(_AES_ENC_us03_n843 ) );
NOR2_X2 _AES_ENC_us03_U180  ( .A1(_AES_ENC_us03_n1029 ), .A2(_AES_ENC_us03_n1095 ), .ZN(_AES_ENC_us03_n735 ) );
NOR4_X2 _AES_ENC_us03_U174  ( .A1(_AES_ENC_us03_n983 ), .A2(_AES_ENC_us03_n982 ), .A3(_AES_ENC_us03_n981 ), .A4(_AES_ENC_us03_n980 ), .ZN(_AES_ENC_us03_n984 ) );
NOR2_X2 _AES_ENC_us03_U173  ( .A1(_AES_ENC_us03_n979 ), .A2(_AES_ENC_us03_n978 ), .ZN(_AES_ENC_us03_n985 ) );
NAND3_X2 _AES_ENC_us03_U172  ( .A1(_AES_ENC_us03_n569 ), .A2(_AES_ENC_us03_n595 ), .A3(_AES_ENC_us03_n681 ), .ZN(_AES_ENC_us03_n691 ) );
NOR2_X2 _AES_ENC_us03_U171  ( .A1(_AES_ENC_us03_n683 ), .A2(_AES_ENC_us03_n682 ), .ZN(_AES_ENC_us03_n690 ) );
NOR3_X2 _AES_ENC_us03_U170  ( .A1(_AES_ENC_us03_n695 ), .A2(_AES_ENC_us03_n694 ), .A3(_AES_ENC_us03_n693 ), .ZN(_AES_ENC_us03_n700 ) );
NOR4_X2 _AES_ENC_us03_U169  ( .A1(_AES_ENC_us03_n983 ), .A2(_AES_ENC_us03_n698 ), .A3(_AES_ENC_us03_n697 ), .A4(_AES_ENC_us03_n696 ), .ZN(_AES_ENC_us03_n699 ) );
NOR2_X2 _AES_ENC_us03_U168  ( .A1(_AES_ENC_us03_n1100 ), .A2(_AES_ENC_us03_n854 ), .ZN(_AES_ENC_us03_n860 ) );
NOR4_X2 _AES_ENC_us03_U162  ( .A1(_AES_ENC_us03_n1125 ), .A2(_AES_ENC_us03_n1124 ), .A3(_AES_ENC_us03_n1123 ), .A4(_AES_ENC_us03_n1122 ), .ZN(_AES_ENC_us03_n1126 ) );
NOR4_X2 _AES_ENC_us03_U161  ( .A1(_AES_ENC_us03_n1084 ), .A2(_AES_ENC_us03_n1083 ), .A3(_AES_ENC_us03_n1082 ), .A4(_AES_ENC_us03_n1081 ), .ZN(_AES_ENC_us03_n1085 ) );
NOR2_X2 _AES_ENC_us03_U160  ( .A1(_AES_ENC_us03_n1076 ), .A2(_AES_ENC_us03_n1075 ), .ZN(_AES_ENC_us03_n1086 ) );
NOR4_X2 _AES_ENC_us03_U159  ( .A1(_AES_ENC_us03_n896 ), .A2(_AES_ENC_us03_n895 ), .A3(_AES_ENC_us03_n894 ), .A4(_AES_ENC_us03_n893 ), .ZN(_AES_ENC_us03_n897 ) );
NOR2_X2 _AES_ENC_us03_U158  ( .A1(_AES_ENC_us03_n866 ), .A2(_AES_ENC_us03_n865 ), .ZN(_AES_ENC_us03_n872 ) );
NOR4_X2 _AES_ENC_us03_U157  ( .A1(_AES_ENC_us03_n870 ), .A2(_AES_ENC_us03_n869 ), .A3(_AES_ENC_us03_n868 ), .A4(_AES_ENC_us03_n867 ), .ZN(_AES_ENC_us03_n871 ) );
NOR2_X2 _AES_ENC_us03_U156  ( .A1(_AES_ENC_us03_n946 ), .A2(_AES_ENC_us03_n945 ), .ZN(_AES_ENC_us03_n952 ) );
NOR4_X2 _AES_ENC_us03_U155  ( .A1(_AES_ENC_us03_n950 ), .A2(_AES_ENC_us03_n949 ), .A3(_AES_ENC_us03_n948 ), .A4(_AES_ENC_us03_n947 ), .ZN(_AES_ENC_us03_n951 ) );
NOR3_X2 _AES_ENC_us03_U154  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n1054 ), .A3(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n961 ) );
NOR3_X2 _AES_ENC_us03_U153  ( .A1(_AES_ENC_us03_n622 ), .A2(_AES_ENC_us03_n1074 ), .A3(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n671 ) );
NOR2_X2 _AES_ENC_us03_U152  ( .A1(_AES_ENC_us03_n1057 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n1062 ) );
NOR2_X2 _AES_ENC_us03_U143  ( .A1(_AES_ENC_us03_n1055 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n1063 ) );
NOR2_X2 _AES_ENC_us03_U142  ( .A1(_AES_ENC_us03_n1060 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n1061 ) );
NOR4_X2 _AES_ENC_us03_U141  ( .A1(_AES_ENC_us03_n1064 ), .A2(_AES_ENC_us03_n1063 ), .A3(_AES_ENC_us03_n1062 ), .A4(_AES_ENC_us03_n1061 ), .ZN(_AES_ENC_us03_n1065 ) );
NOR2_X2 _AES_ENC_us03_U140  ( .A1(_AES_ENC_us03_n735 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n687 ) );
NOR2_X2 _AES_ENC_us03_U132  ( .A1(_AES_ENC_us03_n684 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n688 ) );
NOR2_X2 _AES_ENC_us03_U131  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n612 ), .ZN(_AES_ENC_us03_n686 ) );
NOR4_X2 _AES_ENC_us03_U130  ( .A1(_AES_ENC_us03_n688 ), .A2(_AES_ENC_us03_n687 ), .A3(_AES_ENC_us03_n686 ), .A4(_AES_ENC_us03_n685 ), .ZN(_AES_ENC_us03_n689 ) );
NOR2_X2 _AES_ENC_us03_U129  ( .A1(_AES_ENC_us03_n619 ), .A2(_AES_ENC_us03_n594 ), .ZN(_AES_ENC_us03_n771 ) );
NOR2_X2 _AES_ENC_us03_U128  ( .A1(_AES_ENC_us03_n1103 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n772 ) );
NOR2_X2 _AES_ENC_us03_U127  ( .A1(_AES_ENC_us03_n617 ), .A2(_AES_ENC_us03_n611 ), .ZN(_AES_ENC_us03_n773 ) );
NOR4_X2 _AES_ENC_us03_U126  ( .A1(_AES_ENC_us03_n773 ), .A2(_AES_ENC_us03_n772 ), .A3(_AES_ENC_us03_n771 ), .A4(_AES_ENC_us03_n770 ), .ZN(_AES_ENC_us03_n774 ) );
NOR2_X2 _AES_ENC_us03_U121  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n607 ), .ZN(_AES_ENC_us03_n858 ) );
NOR2_X2 _AES_ENC_us03_U120  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n855 ), .ZN(_AES_ENC_us03_n857 ) );
NOR2_X2 _AES_ENC_us03_U119  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n599 ), .ZN(_AES_ENC_us03_n856 ) );
NOR4_X2 _AES_ENC_us03_U118  ( .A1(_AES_ENC_us03_n858 ), .A2(_AES_ENC_us03_n857 ), .A3(_AES_ENC_us03_n856 ), .A4(_AES_ENC_us03_n958 ), .ZN(_AES_ENC_us03_n859 ) );
NOR3_X2 _AES_ENC_us03_U117  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n1120 ), .A3(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n918 ) );
NOR3_X2 _AES_ENC_us03_U116  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n573 ), .A3(_AES_ENC_us03_n1013 ), .ZN(_AES_ENC_us03_n917 ) );
NOR2_X2 _AES_ENC_us03_U115  ( .A1(_AES_ENC_us03_n914 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n915 ) );
NOR4_X2 _AES_ENC_us03_U106  ( .A1(_AES_ENC_us03_n918 ), .A2(_AES_ENC_us03_n917 ), .A3(_AES_ENC_us03_n916 ), .A4(_AES_ENC_us03_n915 ), .ZN(_AES_ENC_us03_n919 ) );
NOR2_X2 _AES_ENC_us03_U105  ( .A1(_AES_ENC_us03_n780 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n784 ) );
NOR2_X2 _AES_ENC_us03_U104  ( .A1(_AES_ENC_us03_n1117 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n782 ) );
NOR2_X2 _AES_ENC_us03_U103  ( .A1(_AES_ENC_us03_n781 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n783 ) );
NOR4_X2 _AES_ENC_us03_U102  ( .A1(_AES_ENC_us03_n880 ), .A2(_AES_ENC_us03_n784 ), .A3(_AES_ENC_us03_n783 ), .A4(_AES_ENC_us03_n782 ), .ZN(_AES_ENC_us03_n785 ) );
NOR2_X2 _AES_ENC_us03_U101  ( .A1(_AES_ENC_us03_n596 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n814 ) );
NOR2_X2 _AES_ENC_us03_U100  ( .A1(_AES_ENC_us03_n907 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n813 ) );
NOR3_X2 _AES_ENC_us03_U95  ( .A1(_AES_ENC_us03_n588 ), .A2(_AES_ENC_us03_n1058 ), .A3(_AES_ENC_us03_n1059 ), .ZN(_AES_ENC_us03_n815 ) );
NOR4_X2 _AES_ENC_us03_U94  ( .A1(_AES_ENC_us03_n815 ), .A2(_AES_ENC_us03_n814 ), .A3(_AES_ENC_us03_n813 ), .A4(_AES_ENC_us03_n812 ), .ZN(_AES_ENC_us03_n816 ) );
NOR2_X2 _AES_ENC_us03_U93  ( .A1(_AES_ENC_us03_n576 ), .A2(_AES_ENC_us03_n569 ), .ZN(_AES_ENC_us03_n721 ) );
NOR2_X2 _AES_ENC_us03_U92  ( .A1(_AES_ENC_us03_n1031 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n723 ) );
NOR2_X2 _AES_ENC_us03_U91  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n1096 ), .ZN(_AES_ENC_us03_n722 ) );
NOR4_X2 _AES_ENC_us03_U90  ( .A1(_AES_ENC_us03_n724 ), .A2(_AES_ENC_us03_n723 ), .A3(_AES_ENC_us03_n722 ), .A4(_AES_ENC_us03_n721 ), .ZN(_AES_ENC_us03_n725 ) );
NOR2_X2 _AES_ENC_us03_U89  ( .A1(_AES_ENC_us03_n911 ), .A2(_AES_ENC_us03_n990 ), .ZN(_AES_ENC_us03_n1009 ) );
NOR2_X2 _AES_ENC_us03_U88  ( .A1(_AES_ENC_us03_n1013 ), .A2(_AES_ENC_us03_n573 ), .ZN(_AES_ENC_us03_n1014 ) );
NOR2_X2 _AES_ENC_us03_U87  ( .A1(_AES_ENC_us03_n1014 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n1015 ) );
NOR4_X2 _AES_ENC_us03_U86  ( .A1(_AES_ENC_us03_n1016 ), .A2(_AES_ENC_us03_n1015 ), .A3(_AES_ENC_us03_n1119 ), .A4(_AES_ENC_us03_n1046 ), .ZN(_AES_ENC_us03_n1017 ) );
NOR2_X2 _AES_ENC_us03_U81  ( .A1(_AES_ENC_us03_n996 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n998 ) );
NOR2_X2 _AES_ENC_us03_U80  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n592 ), .ZN(_AES_ENC_us03_n1000 ) );
NOR2_X2 _AES_ENC_us03_U79  ( .A1(_AES_ENC_us03_n619 ), .A2(_AES_ENC_us03_n1096 ), .ZN(_AES_ENC_us03_n999 ) );
NOR4_X2 _AES_ENC_us03_U78  ( .A1(_AES_ENC_us03_n1000 ), .A2(_AES_ENC_us03_n999 ), .A3(_AES_ENC_us03_n998 ), .A4(_AES_ENC_us03_n997 ), .ZN(_AES_ENC_us03_n1001 ) );
NOR2_X2 _AES_ENC_us03_U74  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n1096 ), .ZN(_AES_ENC_us03_n697 ) );
NOR2_X2 _AES_ENC_us03_U73  ( .A1(_AES_ENC_us03_n622 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n958 ) );
NOR2_X2 _AES_ENC_us03_U72  ( .A1(_AES_ENC_us03_n911 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n983 ) );
NOR2_X2 _AES_ENC_us03_U71  ( .A1(_AES_ENC_us03_n1054 ), .A2(_AES_ENC_us03_n1103 ), .ZN(_AES_ENC_us03_n1031 ) );
INV_X4 _AES_ENC_us03_U65  ( .A(_AES_ENC_us03_n1050 ), .ZN(_AES_ENC_us03_n583 ) );
INV_X4 _AES_ENC_us03_U64  ( .A(_AES_ENC_us03_n1072 ), .ZN(_AES_ENC_us03_n587 ) );
INV_X4 _AES_ENC_us03_U63  ( .A(_AES_ENC_us03_n1073 ), .ZN(_AES_ENC_us03_n577 ) );
NOR2_X2 _AES_ENC_us03_U62  ( .A1(_AES_ENC_us03_n595 ), .A2(_AES_ENC_us03_n585 ), .ZN(_AES_ENC_us03_n880 ) );
NOR3_X2 _AES_ENC_us03_U61  ( .A1(_AES_ENC_us03_n826 ), .A2(_AES_ENC_us03_n1121 ), .A3(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n946 ) );
INV_X4 _AES_ENC_us03_U59  ( .A(_AES_ENC_us03_n1010 ), .ZN(_AES_ENC_us03_n580 ) );
NOR3_X2 _AES_ENC_us03_U58  ( .A1(_AES_ENC_us03_n573 ), .A2(_AES_ENC_us03_n1029 ), .A3(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n1119 ) );
INV_X4 _AES_ENC_us03_U57  ( .A(_AES_ENC_us03_n956 ), .ZN(_AES_ENC_us03_n581 ) );
NOR2_X2 _AES_ENC_us03_U50  ( .A1(_AES_ENC_us03_n625 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n1013 ) );
NOR2_X2 _AES_ENC_us03_U49  ( .A1(_AES_ENC_us03_n622 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n910 ) );
NOR2_X2 _AES_ENC_us03_U48  ( .A1(_AES_ENC_us03_n569 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n1091 ) );
NOR2_X2 _AES_ENC_us03_U47  ( .A1(_AES_ENC_us03_n624 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n990 ) );
NOR2_X2 _AES_ENC_us03_U46  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_us03_n1121 ), .ZN(_AES_ENC_us03_n996 ) );
NOR2_X2 _AES_ENC_us03_U45  ( .A1(_AES_ENC_us03_n617 ), .A2(_AES_ENC_us03_n612 ), .ZN(_AES_ENC_us03_n628 ) );
NOR2_X2 _AES_ENC_us03_U44  ( .A1(_AES_ENC_us03_n591 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n866 ) );
NOR2_X2 _AES_ENC_us03_U43  ( .A1(_AES_ENC_us03_n615 ), .A2(_AES_ENC_us03_n617 ), .ZN(_AES_ENC_us03_n1006 ) );
NOR2_X2 _AES_ENC_us03_U42  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n1117 ), .ZN(_AES_ENC_us03_n1118 ) );
NOR2_X2 _AES_ENC_us03_U41  ( .A1(_AES_ENC_us03_n1119 ), .A2(_AES_ENC_us03_n1118 ), .ZN(_AES_ENC_us03_n1127 ) );
NOR2_X2 _AES_ENC_us03_U36  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n606 ), .ZN(_AES_ENC_us03_n629 ) );
NOR2_X2 _AES_ENC_us03_U35  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n906 ), .ZN(_AES_ENC_us03_n909 ) );
NOR2_X2 _AES_ENC_us03_U34  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n609 ), .ZN(_AES_ENC_us03_n658 ) );
NOR2_X2 _AES_ENC_us03_U33  ( .A1(_AES_ENC_us03_n1116 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n695 ) );
NOR2_X2 _AES_ENC_us03_U32  ( .A1(_AES_ENC_us03_n1078 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n1083 ) );
NOR2_X2 _AES_ENC_us03_U31  ( .A1(_AES_ENC_us03_n941 ), .A2(_AES_ENC_us03_n580 ), .ZN(_AES_ENC_us03_n724 ) );
NOR2_X2 _AES_ENC_us03_U30  ( .A1(_AES_ENC_us03_n610 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n1107 ) );
NOR2_X2 _AES_ENC_us03_U29  ( .A1(_AES_ENC_us03_n591 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n840 ) );
NOR2_X2 _AES_ENC_us03_U24  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n605 ), .ZN(_AES_ENC_us03_n633 ) );
NOR2_X2 _AES_ENC_us03_U23  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n1080 ), .ZN(_AES_ENC_us03_n1081 ) );
NOR2_X2 _AES_ENC_us03_U21  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n1045 ), .ZN(_AES_ENC_us03_n812 ) );
NOR2_X2 _AES_ENC_us03_U20  ( .A1(_AES_ENC_us03_n1009 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n960 ) );
NOR2_X2 _AES_ENC_us03_U19  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n613 ), .ZN(_AES_ENC_us03_n982 ) );
NOR2_X2 _AES_ENC_us03_U18  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n606 ), .ZN(_AES_ENC_us03_n757 ) );
NOR2_X2 _AES_ENC_us03_U17  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n602 ), .ZN(_AES_ENC_us03_n698 ) );
NOR2_X2 _AES_ENC_us03_U16  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n621 ), .ZN(_AES_ENC_us03_n708 ) );
NOR2_X2 _AES_ENC_us03_U15  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n595 ), .ZN(_AES_ENC_us03_n770 ) );
NOR2_X2 _AES_ENC_us03_U10  ( .A1(_AES_ENC_us03_n621 ), .A2(_AES_ENC_us03_n577 ), .ZN(_AES_ENC_us03_n803 ) );
NOR2_X2 _AES_ENC_us03_U9  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n881 ), .ZN(_AES_ENC_us03_n711 ) );
NOR2_X2 _AES_ENC_us03_U8  ( .A1(_AES_ENC_us03_n581 ), .A2(_AES_ENC_us03_n595 ), .ZN(_AES_ENC_us03_n867 ) );
NOR2_X2 _AES_ENC_us03_U7  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n611 ), .ZN(_AES_ENC_us03_n804 ) );
NOR2_X2 _AES_ENC_us03_U6  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n622 ), .ZN(_AES_ENC_us03_n1046 ) );
OR2_X4 _AES_ENC_us03_U5  ( .A1(_AES_ENC_us03_n626 ), .A2(_AES_ENC_sa03[1]),.ZN(_AES_ENC_us03_n570 ) );
OR2_X4 _AES_ENC_us03_U4  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_sa03[4]),.ZN(_AES_ENC_us03_n569 ) );
NAND2_X2 _AES_ENC_us03_U514  ( .A1(_AES_ENC_us03_n1121 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n1030 ) );
AND2_X2 _AES_ENC_us03_U513  ( .A1(_AES_ENC_us03_n609 ), .A2(_AES_ENC_us03_n1030 ), .ZN(_AES_ENC_us03_n1049 ) );
NAND2_X2 _AES_ENC_us03_U511  ( .A1(_AES_ENC_us03_n1049 ), .A2(_AES_ENC_us03_n794 ), .ZN(_AES_ENC_us03_n637 ) );
AND2_X2 _AES_ENC_us03_U493  ( .A1(_AES_ENC_us03_n779 ), .A2(_AES_ENC_us03_n996 ), .ZN(_AES_ENC_us03_n632 ) );
NAND4_X2 _AES_ENC_us03_U485  ( .A1(_AES_ENC_us03_n637 ), .A2(_AES_ENC_us03_n636 ), .A3(_AES_ENC_us03_n635 ), .A4(_AES_ENC_us03_n634 ), .ZN(_AES_ENC_us03_n638 ) );
NAND2_X2 _AES_ENC_us03_U484  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n638 ), .ZN(_AES_ENC_us03_n679 ) );
NAND2_X2 _AES_ENC_us03_U481  ( .A1(_AES_ENC_us03_n1094 ), .A2(_AES_ENC_us03_n603 ), .ZN(_AES_ENC_us03_n648 ) );
NAND2_X2 _AES_ENC_us03_U476  ( .A1(_AES_ENC_us03_n613 ), .A2(_AES_ENC_us03_n602 ), .ZN(_AES_ENC_us03_n762 ) );
NAND2_X2 _AES_ENC_us03_U475  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n762 ), .ZN(_AES_ENC_us03_n647 ) );
NAND4_X2 _AES_ENC_us03_U457  ( .A1(_AES_ENC_us03_n648 ), .A2(_AES_ENC_us03_n647 ), .A3(_AES_ENC_us03_n646 ), .A4(_AES_ENC_us03_n645 ), .ZN(_AES_ENC_us03_n649 ) );
NAND2_X2 _AES_ENC_us03_U456  ( .A1(_AES_ENC_sa03[0]), .A2(_AES_ENC_us03_n649 ), .ZN(_AES_ENC_us03_n665 ) );
NAND2_X2 _AES_ENC_us03_U454  ( .A1(_AES_ENC_us03_n608 ), .A2(_AES_ENC_us03_n625 ), .ZN(_AES_ENC_us03_n855 ) );
NAND2_X2 _AES_ENC_us03_U453  ( .A1(_AES_ENC_us03_n599 ), .A2(_AES_ENC_us03_n855 ), .ZN(_AES_ENC_us03_n821 ) );
NAND2_X2 _AES_ENC_us03_U452  ( .A1(_AES_ENC_us03_n1093 ), .A2(_AES_ENC_us03_n821 ), .ZN(_AES_ENC_us03_n662 ) );
NAND2_X2 _AES_ENC_us03_U451  ( .A1(_AES_ENC_us03_n621 ), .A2(_AES_ENC_us03_n601 ), .ZN(_AES_ENC_us03_n650 ) );
NAND2_X2 _AES_ENC_us03_U450  ( .A1(_AES_ENC_us03_n956 ), .A2(_AES_ENC_us03_n650 ), .ZN(_AES_ENC_us03_n661 ) );
NAND2_X2 _AES_ENC_us03_U449  ( .A1(_AES_ENC_us03_n627 ), .A2(_AES_ENC_us03_n582 ), .ZN(_AES_ENC_us03_n839 ) );
OR2_X2 _AES_ENC_us03_U446  ( .A1(_AES_ENC_us03_n839 ), .A2(_AES_ENC_us03_n932 ), .ZN(_AES_ENC_us03_n656 ) );
NAND2_X2 _AES_ENC_us03_U445  ( .A1(_AES_ENC_us03_n623 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n1096 ) );
NAND2_X2 _AES_ENC_us03_U444  ( .A1(_AES_ENC_us03_n1030 ), .A2(_AES_ENC_us03_n1096 ), .ZN(_AES_ENC_us03_n651 ) );
NAND2_X2 _AES_ENC_us03_U443  ( .A1(_AES_ENC_us03_n1114 ), .A2(_AES_ENC_us03_n651 ), .ZN(_AES_ENC_us03_n655 ) );
OR3_X2 _AES_ENC_us03_U440  ( .A1(_AES_ENC_us03_n1079 ), .A2(_AES_ENC_sa03[7]), .A3(_AES_ENC_us03_n627 ), .ZN(_AES_ENC_us03_n654 ));
NAND2_X2 _AES_ENC_us03_U439  ( .A1(_AES_ENC_us03_n605 ), .A2(_AES_ENC_us03_n613 ), .ZN(_AES_ENC_us03_n652 ) );
NAND4_X2 _AES_ENC_us03_U437  ( .A1(_AES_ENC_us03_n656 ), .A2(_AES_ENC_us03_n655 ), .A3(_AES_ENC_us03_n654 ), .A4(_AES_ENC_us03_n653 ), .ZN(_AES_ENC_us03_n657 ) );
NAND2_X2 _AES_ENC_us03_U436  ( .A1(_AES_ENC_sa03[2]), .A2(_AES_ENC_us03_n657 ), .ZN(_AES_ENC_us03_n660 ) );
NAND4_X2 _AES_ENC_us03_U432  ( .A1(_AES_ENC_us03_n662 ), .A2(_AES_ENC_us03_n661 ), .A3(_AES_ENC_us03_n660 ), .A4(_AES_ENC_us03_n659 ), .ZN(_AES_ENC_us03_n663 ) );
NAND2_X2 _AES_ENC_us03_U431  ( .A1(_AES_ENC_us03_n663 ), .A2(_AES_ENC_us03_n574 ), .ZN(_AES_ENC_us03_n664 ) );
NAND2_X2 _AES_ENC_us03_U430  ( .A1(_AES_ENC_us03_n665 ), .A2(_AES_ENC_us03_n664 ), .ZN(_AES_ENC_us03_n666 ) );
NAND2_X2 _AES_ENC_us03_U429  ( .A1(_AES_ENC_sa03[6]), .A2(_AES_ENC_us03_n666 ), .ZN(_AES_ENC_us03_n678 ) );
NAND2_X2 _AES_ENC_us03_U426  ( .A1(_AES_ENC_us03_n735 ), .A2(_AES_ENC_us03_n1093 ), .ZN(_AES_ENC_us03_n675 ) );
NAND2_X2 _AES_ENC_us03_U425  ( .A1(_AES_ENC_us03_n600 ), .A2(_AES_ENC_us03_n609 ), .ZN(_AES_ENC_us03_n1045 ) );
OR2_X2 _AES_ENC_us03_U424  ( .A1(_AES_ENC_us03_n1045 ), .A2(_AES_ENC_us03_n587 ), .ZN(_AES_ENC_us03_n674 ) );
NAND2_X2 _AES_ENC_us03_U423  ( .A1(_AES_ENC_sa03[1]), .A2(_AES_ENC_us03_n622 ), .ZN(_AES_ENC_us03_n667 ) );
NAND2_X2 _AES_ENC_us03_U422  ( .A1(_AES_ENC_us03_n621 ), .A2(_AES_ENC_us03_n667 ), .ZN(_AES_ENC_us03_n1071 ) );
NAND4_X2 _AES_ENC_us03_U412  ( .A1(_AES_ENC_us03_n675 ), .A2(_AES_ENC_us03_n674 ), .A3(_AES_ENC_us03_n673 ), .A4(_AES_ENC_us03_n672 ), .ZN(_AES_ENC_us03_n676 ) );
NAND2_X2 _AES_ENC_us03_U411  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n676 ), .ZN(_AES_ENC_us03_n677 ) );
NAND2_X2 _AES_ENC_us03_U408  ( .A1(_AES_ENC_us03_n800 ), .A2(_AES_ENC_us03_n1022 ), .ZN(_AES_ENC_us03_n680 ) );
NAND2_X2 _AES_ENC_us03_U407  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n680 ), .ZN(_AES_ENC_us03_n681 ) );
AND2_X2 _AES_ENC_us03_U402  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n684 ), .ZN(_AES_ENC_us03_n682 ) );
NAND4_X2 _AES_ENC_us03_U395  ( .A1(_AES_ENC_us03_n691 ), .A2(_AES_ENC_us03_n584 ), .A3(_AES_ENC_us03_n690 ), .A4(_AES_ENC_us03_n689 ), .ZN(_AES_ENC_us03_n692 ) );
NAND2_X2 _AES_ENC_us03_U394  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n692 ), .ZN(_AES_ENC_us03_n733 ) );
NAND2_X2 _AES_ENC_us03_U392  ( .A1(_AES_ENC_us03_n977 ), .A2(_AES_ENC_us03_n1050 ), .ZN(_AES_ENC_us03_n702 ) );
NAND2_X2 _AES_ENC_us03_U391  ( .A1(_AES_ENC_us03_n1093 ), .A2(_AES_ENC_us03_n1045 ), .ZN(_AES_ENC_us03_n701 ) );
NAND4_X2 _AES_ENC_us03_U381  ( .A1(_AES_ENC_us03_n702 ), .A2(_AES_ENC_us03_n701 ), .A3(_AES_ENC_us03_n700 ), .A4(_AES_ENC_us03_n699 ), .ZN(_AES_ENC_us03_n703 ) );
NAND2_X2 _AES_ENC_us03_U380  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n703 ), .ZN(_AES_ENC_us03_n732 ) );
AND2_X2 _AES_ENC_us03_U379  ( .A1(_AES_ENC_sa03[0]), .A2(_AES_ENC_sa03[6]),.ZN(_AES_ENC_us03_n1113 ) );
NAND2_X2 _AES_ENC_us03_U378  ( .A1(_AES_ENC_us03_n613 ), .A2(_AES_ENC_us03_n1030 ), .ZN(_AES_ENC_us03_n881 ) );
NAND2_X2 _AES_ENC_us03_U377  ( .A1(_AES_ENC_us03_n1093 ), .A2(_AES_ENC_us03_n881 ), .ZN(_AES_ENC_us03_n715 ) );
NAND2_X2 _AES_ENC_us03_U376  ( .A1(_AES_ENC_us03_n1010 ), .A2(_AES_ENC_us03_n612 ), .ZN(_AES_ENC_us03_n714 ) );
NAND2_X2 _AES_ENC_us03_U375  ( .A1(_AES_ENC_us03_n855 ), .A2(_AES_ENC_us03_n600 ), .ZN(_AES_ENC_us03_n1117 ) );
XNOR2_X2 _AES_ENC_us03_U371  ( .A(_AES_ENC_us03_n618 ), .B(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n824 ) );
NAND4_X2 _AES_ENC_us03_U362  ( .A1(_AES_ENC_us03_n715 ), .A2(_AES_ENC_us03_n714 ), .A3(_AES_ENC_us03_n713 ), .A4(_AES_ENC_us03_n712 ), .ZN(_AES_ENC_us03_n716 ) );
NAND2_X2 _AES_ENC_us03_U361  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n716 ), .ZN(_AES_ENC_us03_n731 ) );
AND2_X2 _AES_ENC_us03_U360  ( .A1(_AES_ENC_sa03[6]), .A2(_AES_ENC_us03_n574 ), .ZN(_AES_ENC_us03_n1131 ) );
NAND2_X2 _AES_ENC_us03_U359  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n717 ) );
NAND2_X2 _AES_ENC_us03_U358  ( .A1(_AES_ENC_us03_n1029 ), .A2(_AES_ENC_us03_n717 ), .ZN(_AES_ENC_us03_n728 ) );
NAND2_X2 _AES_ENC_us03_U357  ( .A1(_AES_ENC_sa03[1]), .A2(_AES_ENC_us03_n626 ), .ZN(_AES_ENC_us03_n1097 ) );
NAND2_X2 _AES_ENC_us03_U356  ( .A1(_AES_ENC_us03_n615 ), .A2(_AES_ENC_us03_n1097 ), .ZN(_AES_ENC_us03_n718 ) );
NAND2_X2 _AES_ENC_us03_U355  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n718 ), .ZN(_AES_ENC_us03_n727 ) );
NAND4_X2 _AES_ENC_us03_U344  ( .A1(_AES_ENC_us03_n728 ), .A2(_AES_ENC_us03_n727 ), .A3(_AES_ENC_us03_n726 ), .A4(_AES_ENC_us03_n725 ), .ZN(_AES_ENC_us03_n729 ) );
NAND2_X2 _AES_ENC_us03_U343  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n729 ), .ZN(_AES_ENC_us03_n730 ) );
NAND4_X2 _AES_ENC_us03_U342  ( .A1(_AES_ENC_us03_n733 ), .A2(_AES_ENC_us03_n732 ), .A3(_AES_ENC_us03_n731 ), .A4(_AES_ENC_us03_n730 ), .ZN(_AES_ENC_sa03_sub[1] ) );
NAND2_X2 _AES_ENC_us03_U341  ( .A1(_AES_ENC_sa03[7]), .A2(_AES_ENC_us03_n618 ), .ZN(_AES_ENC_us03_n734 ) );
NAND2_X2 _AES_ENC_us03_U340  ( .A1(_AES_ENC_us03_n734 ), .A2(_AES_ENC_us03_n589 ), .ZN(_AES_ENC_us03_n738 ) );
OR4_X2 _AES_ENC_us03_U339  ( .A1(_AES_ENC_us03_n738 ), .A2(_AES_ENC_us03_n627 ), .A3(_AES_ENC_us03_n826 ), .A4(_AES_ENC_us03_n1121 ), .ZN(_AES_ENC_us03_n746 ) );
NAND2_X2 _AES_ENC_us03_U337  ( .A1(_AES_ENC_us03_n1100 ), .A2(_AES_ENC_us03_n599 ), .ZN(_AES_ENC_us03_n992 ) );
OR2_X2 _AES_ENC_us03_U336  ( .A1(_AES_ENC_us03_n617 ), .A2(_AES_ENC_us03_n735 ), .ZN(_AES_ENC_us03_n737 ) );
NAND2_X2 _AES_ENC_us03_U334  ( .A1(_AES_ENC_us03_n621 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n753 ) );
NAND2_X2 _AES_ENC_us03_U333  ( .A1(_AES_ENC_us03_n595 ), .A2(_AES_ENC_us03_n753 ), .ZN(_AES_ENC_us03_n1080 ) );
NAND2_X2 _AES_ENC_us03_U332  ( .A1(_AES_ENC_us03_n1048 ), .A2(_AES_ENC_us03_n591 ), .ZN(_AES_ENC_us03_n736 ) );
NAND2_X2 _AES_ENC_us03_U331  ( .A1(_AES_ENC_us03_n737 ), .A2(_AES_ENC_us03_n736 ), .ZN(_AES_ENC_us03_n739 ) );
NAND2_X2 _AES_ENC_us03_U330  ( .A1(_AES_ENC_us03_n739 ), .A2(_AES_ENC_us03_n738 ), .ZN(_AES_ENC_us03_n745 ) );
NAND2_X2 _AES_ENC_us03_U326  ( .A1(_AES_ENC_us03_n1096 ), .A2(_AES_ENC_us03_n602 ), .ZN(_AES_ENC_us03_n906 ) );
NAND4_X2 _AES_ENC_us03_U323  ( .A1(_AES_ENC_us03_n746 ), .A2(_AES_ENC_us03_n992 ), .A3(_AES_ENC_us03_n745 ), .A4(_AES_ENC_us03_n744 ), .ZN(_AES_ENC_us03_n747 ) );
NAND2_X2 _AES_ENC_us03_U322  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n747 ), .ZN(_AES_ENC_us03_n793 ) );
NAND2_X2 _AES_ENC_us03_U321  ( .A1(_AES_ENC_us03_n597 ), .A2(_AES_ENC_us03_n855 ), .ZN(_AES_ENC_us03_n748 ) );
NAND2_X2 _AES_ENC_us03_U320  ( .A1(_AES_ENC_us03_n956 ), .A2(_AES_ENC_us03_n748 ), .ZN(_AES_ENC_us03_n760 ) );
NAND2_X2 _AES_ENC_us03_U313  ( .A1(_AES_ENC_us03_n602 ), .A2(_AES_ENC_us03_n753 ), .ZN(_AES_ENC_us03_n1023 ) );
NAND4_X2 _AES_ENC_us03_U308  ( .A1(_AES_ENC_us03_n760 ), .A2(_AES_ENC_us03_n992 ), .A3(_AES_ENC_us03_n759 ), .A4(_AES_ENC_us03_n758 ), .ZN(_AES_ENC_us03_n761 ) );
NAND2_X2 _AES_ENC_us03_U307  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n761 ), .ZN(_AES_ENC_us03_n792 ) );
NAND2_X2 _AES_ENC_us03_U306  ( .A1(_AES_ENC_us03_n597 ), .A2(_AES_ENC_us03_n615 ), .ZN(_AES_ENC_us03_n989 ) );
NAND2_X2 _AES_ENC_us03_U305  ( .A1(_AES_ENC_us03_n1050 ), .A2(_AES_ENC_us03_n989 ), .ZN(_AES_ENC_us03_n777 ) );
NAND2_X2 _AES_ENC_us03_U304  ( .A1(_AES_ENC_us03_n1093 ), .A2(_AES_ENC_us03_n762 ), .ZN(_AES_ENC_us03_n776 ) );
XNOR2_X2 _AES_ENC_us03_U301  ( .A(_AES_ENC_sa03[7]), .B(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n959 ) );
NAND4_X2 _AES_ENC_us03_U289  ( .A1(_AES_ENC_us03_n777 ), .A2(_AES_ENC_us03_n776 ), .A3(_AES_ENC_us03_n775 ), .A4(_AES_ENC_us03_n774 ), .ZN(_AES_ENC_us03_n778 ) );
NAND2_X2 _AES_ENC_us03_U288  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n778 ), .ZN(_AES_ENC_us03_n791 ) );
NAND2_X2 _AES_ENC_us03_U287  ( .A1(_AES_ENC_us03_n1056 ), .A2(_AES_ENC_us03_n1050 ), .ZN(_AES_ENC_us03_n788 ) );
NAND2_X2 _AES_ENC_us03_U286  ( .A1(_AES_ENC_us03_n1091 ), .A2(_AES_ENC_us03_n779 ), .ZN(_AES_ENC_us03_n787 ) );
NAND2_X2 _AES_ENC_us03_U285  ( .A1(_AES_ENC_us03_n956 ), .A2(_AES_ENC_sa03[1]), .ZN(_AES_ENC_us03_n786 ) );
NAND4_X2 _AES_ENC_us03_U278  ( .A1(_AES_ENC_us03_n788 ), .A2(_AES_ENC_us03_n787 ), .A3(_AES_ENC_us03_n786 ), .A4(_AES_ENC_us03_n785 ), .ZN(_AES_ENC_us03_n789 ) );
NAND2_X2 _AES_ENC_us03_U277  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n789 ), .ZN(_AES_ENC_us03_n790 ) );
NAND4_X2 _AES_ENC_us03_U276  ( .A1(_AES_ENC_us03_n793 ), .A2(_AES_ENC_us03_n792 ), .A3(_AES_ENC_us03_n791 ), .A4(_AES_ENC_us03_n790 ), .ZN(_AES_ENC_sa03_sub[2] ) );
NAND2_X2 _AES_ENC_us03_U275  ( .A1(_AES_ENC_us03_n1059 ), .A2(_AES_ENC_us03_n794 ), .ZN(_AES_ENC_us03_n810 ) );
NAND2_X2 _AES_ENC_us03_U274  ( .A1(_AES_ENC_us03_n1049 ), .A2(_AES_ENC_us03_n956 ), .ZN(_AES_ENC_us03_n809 ) );
OR2_X2 _AES_ENC_us03_U266  ( .A1(_AES_ENC_us03_n1096 ), .A2(_AES_ENC_us03_n588 ), .ZN(_AES_ENC_us03_n802 ) );
NAND2_X2 _AES_ENC_us03_U265  ( .A1(_AES_ENC_us03_n1053 ), .A2(_AES_ENC_us03_n800 ), .ZN(_AES_ENC_us03_n801 ) );
NAND2_X2 _AES_ENC_us03_U264  ( .A1(_AES_ENC_us03_n802 ), .A2(_AES_ENC_us03_n801 ), .ZN(_AES_ENC_us03_n805 ) );
NAND4_X2 _AES_ENC_us03_U261  ( .A1(_AES_ENC_us03_n810 ), .A2(_AES_ENC_us03_n809 ), .A3(_AES_ENC_us03_n808 ), .A4(_AES_ENC_us03_n807 ), .ZN(_AES_ENC_us03_n811 ) );
NAND2_X2 _AES_ENC_us03_U260  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n811 ), .ZN(_AES_ENC_us03_n852 ) );
OR2_X2 _AES_ENC_us03_U259  ( .A1(_AES_ENC_us03_n1023 ), .A2(_AES_ENC_us03_n576 ), .ZN(_AES_ENC_us03_n819 ) );
OR2_X2 _AES_ENC_us03_U257  ( .A1(_AES_ENC_us03_n570 ), .A2(_AES_ENC_us03_n930 ), .ZN(_AES_ENC_us03_n818 ) );
NAND2_X2 _AES_ENC_us03_U256  ( .A1(_AES_ENC_us03_n1013 ), .A2(_AES_ENC_us03_n1094 ), .ZN(_AES_ENC_us03_n817 ) );
NAND4_X2 _AES_ENC_us03_U249  ( .A1(_AES_ENC_us03_n819 ), .A2(_AES_ENC_us03_n818 ), .A3(_AES_ENC_us03_n817 ), .A4(_AES_ENC_us03_n816 ), .ZN(_AES_ENC_us03_n820 ) );
NAND2_X2 _AES_ENC_us03_U248  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n820 ), .ZN(_AES_ENC_us03_n851 ) );
NAND2_X2 _AES_ENC_us03_U247  ( .A1(_AES_ENC_us03_n956 ), .A2(_AES_ENC_us03_n1080 ), .ZN(_AES_ENC_us03_n835 ) );
NAND2_X2 _AES_ENC_us03_U246  ( .A1(_AES_ENC_us03_n570 ), .A2(_AES_ENC_us03_n1030 ), .ZN(_AES_ENC_us03_n1047 ) );
OR2_X2 _AES_ENC_us03_U245  ( .A1(_AES_ENC_us03_n1047 ), .A2(_AES_ENC_us03_n583 ), .ZN(_AES_ENC_us03_n834 ) );
NAND2_X2 _AES_ENC_us03_U244  ( .A1(_AES_ENC_us03_n1072 ), .A2(_AES_ENC_us03_n601 ), .ZN(_AES_ENC_us03_n833 ) );
NAND4_X2 _AES_ENC_us03_U233  ( .A1(_AES_ENC_us03_n835 ), .A2(_AES_ENC_us03_n834 ), .A3(_AES_ENC_us03_n833 ), .A4(_AES_ENC_us03_n832 ), .ZN(_AES_ENC_us03_n836 ) );
NAND2_X2 _AES_ENC_us03_U232  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n836 ), .ZN(_AES_ENC_us03_n850 ) );
NAND2_X2 _AES_ENC_us03_U231  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n625 ), .ZN(_AES_ENC_us03_n847 ) );
NAND2_X2 _AES_ENC_us03_U230  ( .A1(_AES_ENC_us03_n1050 ), .A2(_AES_ENC_us03_n1071 ), .ZN(_AES_ENC_us03_n846 ) );
OR2_X2 _AES_ENC_us03_U224  ( .A1(_AES_ENC_us03_n1053 ), .A2(_AES_ENC_us03_n911 ), .ZN(_AES_ENC_us03_n1077 ) );
NAND4_X2 _AES_ENC_us03_U220  ( .A1(_AES_ENC_us03_n847 ), .A2(_AES_ENC_us03_n846 ), .A3(_AES_ENC_us03_n845 ), .A4(_AES_ENC_us03_n844 ), .ZN(_AES_ENC_us03_n848 ) );
NAND2_X2 _AES_ENC_us03_U219  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n848 ), .ZN(_AES_ENC_us03_n849 ) );
NAND4_X2 _AES_ENC_us03_U218  ( .A1(_AES_ENC_us03_n852 ), .A2(_AES_ENC_us03_n851 ), .A3(_AES_ENC_us03_n850 ), .A4(_AES_ENC_us03_n849 ), .ZN(_AES_ENC_sa03_sub[3] ) );
NAND2_X2 _AES_ENC_us03_U216  ( .A1(_AES_ENC_us03_n1009 ), .A2(_AES_ENC_us03_n1072 ), .ZN(_AES_ENC_us03_n862 ) );
NAND2_X2 _AES_ENC_us03_U215  ( .A1(_AES_ENC_us03_n615 ), .A2(_AES_ENC_us03_n592 ), .ZN(_AES_ENC_us03_n853 ) );
NAND2_X2 _AES_ENC_us03_U214  ( .A1(_AES_ENC_us03_n1050 ), .A2(_AES_ENC_us03_n853 ), .ZN(_AES_ENC_us03_n861 ) );
NAND4_X2 _AES_ENC_us03_U206  ( .A1(_AES_ENC_us03_n862 ), .A2(_AES_ENC_us03_n861 ), .A3(_AES_ENC_us03_n860 ), .A4(_AES_ENC_us03_n859 ), .ZN(_AES_ENC_us03_n863 ) );
NAND2_X2 _AES_ENC_us03_U205  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n863 ), .ZN(_AES_ENC_us03_n905 ) );
NAND2_X2 _AES_ENC_us03_U204  ( .A1(_AES_ENC_us03_n1010 ), .A2(_AES_ENC_us03_n989 ), .ZN(_AES_ENC_us03_n874 ) );
NAND2_X2 _AES_ENC_us03_U203  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n617 ), .ZN(_AES_ENC_us03_n864 ) );
NAND2_X2 _AES_ENC_us03_U202  ( .A1(_AES_ENC_us03_n929 ), .A2(_AES_ENC_us03_n864 ), .ZN(_AES_ENC_us03_n873 ) );
NAND4_X2 _AES_ENC_us03_U193  ( .A1(_AES_ENC_us03_n874 ), .A2(_AES_ENC_us03_n873 ), .A3(_AES_ENC_us03_n872 ), .A4(_AES_ENC_us03_n871 ), .ZN(_AES_ENC_us03_n875 ) );
NAND2_X2 _AES_ENC_us03_U192  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n875 ), .ZN(_AES_ENC_us03_n904 ) );
NAND2_X2 _AES_ENC_us03_U191  ( .A1(_AES_ENC_us03_n596 ), .A2(_AES_ENC_us03_n1050 ), .ZN(_AES_ENC_us03_n889 ) );
NAND2_X2 _AES_ENC_us03_U190  ( .A1(_AES_ENC_us03_n1093 ), .A2(_AES_ENC_us03_n599 ), .ZN(_AES_ENC_us03_n876 ) );
NAND2_X2 _AES_ENC_us03_U189  ( .A1(_AES_ENC_us03_n577 ), .A2(_AES_ENC_us03_n876 ), .ZN(_AES_ENC_us03_n877 ) );
NAND2_X2 _AES_ENC_us03_U188  ( .A1(_AES_ENC_us03_n877 ), .A2(_AES_ENC_us03_n625 ), .ZN(_AES_ENC_us03_n888 ) );
NAND4_X2 _AES_ENC_us03_U179  ( .A1(_AES_ENC_us03_n889 ), .A2(_AES_ENC_us03_n888 ), .A3(_AES_ENC_us03_n887 ), .A4(_AES_ENC_us03_n886 ), .ZN(_AES_ENC_us03_n890 ) );
NAND2_X2 _AES_ENC_us03_U178  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n890 ), .ZN(_AES_ENC_us03_n903 ) );
OR2_X2 _AES_ENC_us03_U177  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n1059 ), .ZN(_AES_ENC_us03_n900 ) );
NAND2_X2 _AES_ENC_us03_U176  ( .A1(_AES_ENC_us03_n1073 ), .A2(_AES_ENC_us03_n1047 ), .ZN(_AES_ENC_us03_n899 ) );
NAND2_X2 _AES_ENC_us03_U175  ( .A1(_AES_ENC_us03_n1094 ), .A2(_AES_ENC_us03_n607 ), .ZN(_AES_ENC_us03_n898 ) );
NAND4_X2 _AES_ENC_us03_U167  ( .A1(_AES_ENC_us03_n900 ), .A2(_AES_ENC_us03_n899 ), .A3(_AES_ENC_us03_n898 ), .A4(_AES_ENC_us03_n897 ), .ZN(_AES_ENC_us03_n901 ) );
NAND2_X2 _AES_ENC_us03_U166  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n901 ), .ZN(_AES_ENC_us03_n902 ) );
NAND4_X2 _AES_ENC_us03_U165  ( .A1(_AES_ENC_us03_n905 ), .A2(_AES_ENC_us03_n904 ), .A3(_AES_ENC_us03_n903 ), .A4(_AES_ENC_us03_n902 ), .ZN(_AES_ENC_sa03_sub[4] ) );
NAND2_X2 _AES_ENC_us03_U164  ( .A1(_AES_ENC_us03_n1094 ), .A2(_AES_ENC_us03_n611 ), .ZN(_AES_ENC_us03_n922 ) );
NAND2_X2 _AES_ENC_us03_U163  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n989 ), .ZN(_AES_ENC_us03_n921 ) );
NAND4_X2 _AES_ENC_us03_U151  ( .A1(_AES_ENC_us03_n922 ), .A2(_AES_ENC_us03_n921 ), .A3(_AES_ENC_us03_n920 ), .A4(_AES_ENC_us03_n919 ), .ZN(_AES_ENC_us03_n923 ) );
NAND2_X2 _AES_ENC_us03_U150  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n923 ), .ZN(_AES_ENC_us03_n972 ) );
NAND2_X2 _AES_ENC_us03_U149  ( .A1(_AES_ENC_us03_n595 ), .A2(_AES_ENC_us03_n621 ), .ZN(_AES_ENC_us03_n924 ) );
NAND2_X2 _AES_ENC_us03_U148  ( .A1(_AES_ENC_us03_n1073 ), .A2(_AES_ENC_us03_n924 ), .ZN(_AES_ENC_us03_n939 ) );
NAND2_X2 _AES_ENC_us03_U147  ( .A1(_AES_ENC_us03_n926 ), .A2(_AES_ENC_us03_n925 ), .ZN(_AES_ENC_us03_n927 ) );
NAND2_X2 _AES_ENC_us03_U146  ( .A1(_AES_ENC_us03_n588 ), .A2(_AES_ENC_us03_n927 ), .ZN(_AES_ENC_us03_n928 ) );
NAND2_X2 _AES_ENC_us03_U145  ( .A1(_AES_ENC_us03_n928 ), .A2(_AES_ENC_us03_n1080 ), .ZN(_AES_ENC_us03_n938 ) );
OR2_X2 _AES_ENC_us03_U144  ( .A1(_AES_ENC_us03_n1117 ), .A2(_AES_ENC_us03_n581 ), .ZN(_AES_ENC_us03_n937 ) );
NAND4_X2 _AES_ENC_us03_U139  ( .A1(_AES_ENC_us03_n939 ), .A2(_AES_ENC_us03_n938 ), .A3(_AES_ENC_us03_n937 ), .A4(_AES_ENC_us03_n936 ), .ZN(_AES_ENC_us03_n940 ) );
NAND2_X2 _AES_ENC_us03_U138  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n940 ), .ZN(_AES_ENC_us03_n971 ) );
OR2_X2 _AES_ENC_us03_U137  ( .A1(_AES_ENC_us03_n587 ), .A2(_AES_ENC_us03_n941 ), .ZN(_AES_ENC_us03_n954 ) );
NAND2_X2 _AES_ENC_us03_U136  ( .A1(_AES_ENC_us03_n1096 ), .A2(_AES_ENC_us03_n592 ), .ZN(_AES_ENC_us03_n942 ) );
NAND2_X2 _AES_ENC_us03_U135  ( .A1(_AES_ENC_us03_n1048 ), .A2(_AES_ENC_us03_n942 ), .ZN(_AES_ENC_us03_n943 ) );
NAND2_X2 _AES_ENC_us03_U134  ( .A1(_AES_ENC_us03_n583 ), .A2(_AES_ENC_us03_n943 ), .ZN(_AES_ENC_us03_n944 ) );
NAND2_X2 _AES_ENC_us03_U133  ( .A1(_AES_ENC_us03_n944 ), .A2(_AES_ENC_us03_n594 ), .ZN(_AES_ENC_us03_n953 ) );
NAND4_X2 _AES_ENC_us03_U125  ( .A1(_AES_ENC_us03_n954 ), .A2(_AES_ENC_us03_n953 ), .A3(_AES_ENC_us03_n952 ), .A4(_AES_ENC_us03_n951 ), .ZN(_AES_ENC_us03_n955 ) );
NAND2_X2 _AES_ENC_us03_U124  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n955 ), .ZN(_AES_ENC_us03_n970 ) );
NAND2_X2 _AES_ENC_us03_U123  ( .A1(_AES_ENC_us03_n1094 ), .A2(_AES_ENC_us03_n1071 ), .ZN(_AES_ENC_us03_n967 ) );
NAND2_X2 _AES_ENC_us03_U122  ( .A1(_AES_ENC_us03_n956 ), .A2(_AES_ENC_us03_n1030 ), .ZN(_AES_ENC_us03_n966 ) );
NAND4_X2 _AES_ENC_us03_U114  ( .A1(_AES_ENC_us03_n967 ), .A2(_AES_ENC_us03_n966 ), .A3(_AES_ENC_us03_n965 ), .A4(_AES_ENC_us03_n964 ), .ZN(_AES_ENC_us03_n968 ) );
NAND2_X2 _AES_ENC_us03_U113  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n968 ), .ZN(_AES_ENC_us03_n969 ) );
NAND4_X2 _AES_ENC_us03_U112  ( .A1(_AES_ENC_us03_n972 ), .A2(_AES_ENC_us03_n971 ), .A3(_AES_ENC_us03_n970 ), .A4(_AES_ENC_us03_n969 ), .ZN(_AES_ENC_sa03_sub[5] ) );
NAND2_X2 _AES_ENC_us03_U111  ( .A1(_AES_ENC_us03_n570 ), .A2(_AES_ENC_us03_n1097 ), .ZN(_AES_ENC_us03_n973 ) );
NAND2_X2 _AES_ENC_us03_U110  ( .A1(_AES_ENC_us03_n1073 ), .A2(_AES_ENC_us03_n973 ), .ZN(_AES_ENC_us03_n987 ) );
NAND2_X2 _AES_ENC_us03_U109  ( .A1(_AES_ENC_us03_n974 ), .A2(_AES_ENC_us03_n1077 ), .ZN(_AES_ENC_us03_n975 ) );
NAND2_X2 _AES_ENC_us03_U108  ( .A1(_AES_ENC_us03_n585 ), .A2(_AES_ENC_us03_n975 ), .ZN(_AES_ENC_us03_n976 ) );
NAND2_X2 _AES_ENC_us03_U107  ( .A1(_AES_ENC_us03_n977 ), .A2(_AES_ENC_us03_n976 ), .ZN(_AES_ENC_us03_n986 ) );
NAND4_X2 _AES_ENC_us03_U99  ( .A1(_AES_ENC_us03_n987 ), .A2(_AES_ENC_us03_n986 ), .A3(_AES_ENC_us03_n985 ), .A4(_AES_ENC_us03_n984 ), .ZN(_AES_ENC_us03_n988 ) );
NAND2_X2 _AES_ENC_us03_U98  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n988 ), .ZN(_AES_ENC_us03_n1044 ) );
NAND2_X2 _AES_ENC_us03_U97  ( .A1(_AES_ENC_us03_n1073 ), .A2(_AES_ENC_us03_n989 ), .ZN(_AES_ENC_us03_n1004 ) );
NAND2_X2 _AES_ENC_us03_U96  ( .A1(_AES_ENC_us03_n1092 ), .A2(_AES_ENC_us03_n621 ), .ZN(_AES_ENC_us03_n1003 ) );
NAND4_X2 _AES_ENC_us03_U85  ( .A1(_AES_ENC_us03_n1004 ), .A2(_AES_ENC_us03_n1003 ), .A3(_AES_ENC_us03_n1002 ), .A4(_AES_ENC_us03_n1001 ), .ZN(_AES_ENC_us03_n1005 ) );
NAND2_X2 _AES_ENC_us03_U84  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n1005 ), .ZN(_AES_ENC_us03_n1043 ) );
NAND2_X2 _AES_ENC_us03_U83  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n608 ), .ZN(_AES_ENC_us03_n1020 ) );
NAND2_X2 _AES_ENC_us03_U82  ( .A1(_AES_ENC_us03_n1050 ), .A2(_AES_ENC_us03_n626 ), .ZN(_AES_ENC_us03_n1019 ) );
NAND2_X2 _AES_ENC_us03_U77  ( .A1(_AES_ENC_us03_n1059 ), .A2(_AES_ENC_us03_n1114 ), .ZN(_AES_ENC_us03_n1012 ) );
NAND2_X2 _AES_ENC_us03_U76  ( .A1(_AES_ENC_us03_n1010 ), .A2(_AES_ENC_us03_n604 ), .ZN(_AES_ENC_us03_n1011 ) );
NAND2_X2 _AES_ENC_us03_U75  ( .A1(_AES_ENC_us03_n1012 ), .A2(_AES_ENC_us03_n1011 ), .ZN(_AES_ENC_us03_n1016 ) );
NAND4_X2 _AES_ENC_us03_U70  ( .A1(_AES_ENC_us03_n1020 ), .A2(_AES_ENC_us03_n1019 ), .A3(_AES_ENC_us03_n1018 ), .A4(_AES_ENC_us03_n1017 ), .ZN(_AES_ENC_us03_n1021 ) );
NAND2_X2 _AES_ENC_us03_U69  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n1021 ), .ZN(_AES_ENC_us03_n1042 ) );
NAND2_X2 _AES_ENC_us03_U68  ( .A1(_AES_ENC_us03_n1022 ), .A2(_AES_ENC_us03_n1093 ), .ZN(_AES_ENC_us03_n1039 ) );
NAND2_X2 _AES_ENC_us03_U67  ( .A1(_AES_ENC_us03_n1050 ), .A2(_AES_ENC_us03_n1023 ), .ZN(_AES_ENC_us03_n1038 ) );
NAND2_X2 _AES_ENC_us03_U66  ( .A1(_AES_ENC_us03_n1024 ), .A2(_AES_ENC_us03_n1071 ), .ZN(_AES_ENC_us03_n1037 ) );
AND2_X2 _AES_ENC_us03_U60  ( .A1(_AES_ENC_us03_n1030 ), .A2(_AES_ENC_us03_n614 ), .ZN(_AES_ENC_us03_n1078 ) );
NAND4_X2 _AES_ENC_us03_U56  ( .A1(_AES_ENC_us03_n1039 ), .A2(_AES_ENC_us03_n1038 ), .A3(_AES_ENC_us03_n1037 ), .A4(_AES_ENC_us03_n1036 ), .ZN(_AES_ENC_us03_n1040 ) );
NAND2_X2 _AES_ENC_us03_U55  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n1040 ), .ZN(_AES_ENC_us03_n1041 ) );
NAND4_X2 _AES_ENC_us03_U54  ( .A1(_AES_ENC_us03_n1044 ), .A2(_AES_ENC_us03_n1043 ), .A3(_AES_ENC_us03_n1042 ), .A4(_AES_ENC_us03_n1041 ), .ZN(_AES_ENC_sa03_sub[6] ) );
NAND2_X2 _AES_ENC_us03_U53  ( .A1(_AES_ENC_us03_n1072 ), .A2(_AES_ENC_us03_n1045 ), .ZN(_AES_ENC_us03_n1068 ) );
NAND2_X2 _AES_ENC_us03_U52  ( .A1(_AES_ENC_us03_n1046 ), .A2(_AES_ENC_us03_n595 ), .ZN(_AES_ENC_us03_n1067 ) );
NAND2_X2 _AES_ENC_us03_U51  ( .A1(_AES_ENC_us03_n1094 ), .A2(_AES_ENC_us03_n1047 ), .ZN(_AES_ENC_us03_n1066 ) );
NAND4_X2 _AES_ENC_us03_U40  ( .A1(_AES_ENC_us03_n1068 ), .A2(_AES_ENC_us03_n1067 ), .A3(_AES_ENC_us03_n1066 ), .A4(_AES_ENC_us03_n1065 ), .ZN(_AES_ENC_us03_n1069 ) );
NAND2_X2 _AES_ENC_us03_U39  ( .A1(_AES_ENC_us03_n1070 ), .A2(_AES_ENC_us03_n1069 ), .ZN(_AES_ENC_us03_n1135 ) );
NAND2_X2 _AES_ENC_us03_U38  ( .A1(_AES_ENC_us03_n1072 ), .A2(_AES_ENC_us03_n1071 ), .ZN(_AES_ENC_us03_n1088 ) );
NAND2_X2 _AES_ENC_us03_U37  ( .A1(_AES_ENC_us03_n1073 ), .A2(_AES_ENC_us03_n607 ), .ZN(_AES_ENC_us03_n1087 ) );
NAND4_X2 _AES_ENC_us03_U28  ( .A1(_AES_ENC_us03_n1088 ), .A2(_AES_ENC_us03_n1087 ), .A3(_AES_ENC_us03_n1086 ), .A4(_AES_ENC_us03_n1085 ), .ZN(_AES_ENC_us03_n1089 ) );
NAND2_X2 _AES_ENC_us03_U27  ( .A1(_AES_ENC_us03_n1090 ), .A2(_AES_ENC_us03_n1089 ), .ZN(_AES_ENC_us03_n1134 ) );
NAND2_X2 _AES_ENC_us03_U26  ( .A1(_AES_ENC_us03_n1091 ), .A2(_AES_ENC_us03_n1093 ), .ZN(_AES_ENC_us03_n1111 ) );
NAND2_X2 _AES_ENC_us03_U25  ( .A1(_AES_ENC_us03_n1092 ), .A2(_AES_ENC_us03_n1120 ), .ZN(_AES_ENC_us03_n1110 ) );
AND2_X2 _AES_ENC_us03_U22  ( .A1(_AES_ENC_us03_n1097 ), .A2(_AES_ENC_us03_n1096 ), .ZN(_AES_ENC_us03_n1098 ) );
NAND4_X2 _AES_ENC_us03_U14  ( .A1(_AES_ENC_us03_n1111 ), .A2(_AES_ENC_us03_n1110 ), .A3(_AES_ENC_us03_n1109 ), .A4(_AES_ENC_us03_n1108 ), .ZN(_AES_ENC_us03_n1112 ) );
NAND2_X2 _AES_ENC_us03_U13  ( .A1(_AES_ENC_us03_n1113 ), .A2(_AES_ENC_us03_n1112 ), .ZN(_AES_ENC_us03_n1133 ) );
NAND2_X2 _AES_ENC_us03_U12  ( .A1(_AES_ENC_us03_n1115 ), .A2(_AES_ENC_us03_n1114 ), .ZN(_AES_ENC_us03_n1129 ) );
OR2_X2 _AES_ENC_us03_U11  ( .A1(_AES_ENC_us03_n580 ), .A2(_AES_ENC_us03_n1116 ), .ZN(_AES_ENC_us03_n1128 ) );
NAND4_X2 _AES_ENC_us03_U3  ( .A1(_AES_ENC_us03_n1129 ), .A2(_AES_ENC_us03_n1128 ), .A3(_AES_ENC_us03_n1127 ), .A4(_AES_ENC_us03_n1126 ), .ZN(_AES_ENC_us03_n1130 ) );
NAND2_X2 _AES_ENC_us03_U2  ( .A1(_AES_ENC_us03_n1131 ), .A2(_AES_ENC_us03_n1130 ), .ZN(_AES_ENC_us03_n1132 ) );
NAND4_X2 _AES_ENC_us03_U1  ( .A1(_AES_ENC_us03_n1135 ), .A2(_AES_ENC_us03_n1134 ), .A3(_AES_ENC_us03_n1133 ), .A4(_AES_ENC_us03_n1132 ), .ZN(_AES_ENC_sa03_sub[7] ) );
INV_X4 _AES_ENC_us10_U575  ( .A(_AES_ENC_sa10[7]), .ZN(_AES_ENC_us10_n627 ));
INV_X4 _AES_ENC_us10_U574  ( .A(_AES_ENC_us10_n1114 ), .ZN(_AES_ENC_us10_n625 ) );
INV_X4 _AES_ENC_us10_U573  ( .A(_AES_ENC_sa10[4]), .ZN(_AES_ENC_us10_n624 ));
INV_X4 _AES_ENC_us10_U572  ( .A(_AES_ENC_us10_n1025 ), .ZN(_AES_ENC_us10_n622 ) );
INV_X4 _AES_ENC_us10_U571  ( .A(_AES_ENC_us10_n1120 ), .ZN(_AES_ENC_us10_n620 ) );
INV_X4 _AES_ENC_us10_U570  ( .A(_AES_ENC_us10_n1121 ), .ZN(_AES_ENC_us10_n619 ) );
INV_X4 _AES_ENC_us10_U569  ( .A(_AES_ENC_us10_n1048 ), .ZN(_AES_ENC_us10_n618 ) );
INV_X4 _AES_ENC_us10_U568  ( .A(_AES_ENC_us10_n974 ), .ZN(_AES_ENC_us10_n616 ) );
INV_X4 _AES_ENC_us10_U567  ( .A(_AES_ENC_us10_n794 ), .ZN(_AES_ENC_us10_n614 ) );
INV_X4 _AES_ENC_us10_U566  ( .A(_AES_ENC_sa10[2]), .ZN(_AES_ENC_us10_n611 ));
INV_X4 _AES_ENC_us10_U565  ( .A(_AES_ENC_us10_n800 ), .ZN(_AES_ENC_us10_n610 ) );
INV_X4 _AES_ENC_us10_U564  ( .A(_AES_ENC_us10_n925 ), .ZN(_AES_ENC_us10_n609 ) );
INV_X4 _AES_ENC_us10_U563  ( .A(_AES_ENC_us10_n779 ), .ZN(_AES_ENC_us10_n607 ) );
INV_X4 _AES_ENC_us10_U562  ( .A(_AES_ENC_us10_n1022 ), .ZN(_AES_ENC_us10_n603 ) );
INV_X4 _AES_ENC_us10_U561  ( .A(_AES_ENC_us10_n1102 ), .ZN(_AES_ENC_us10_n602 ) );
INV_X4 _AES_ENC_us10_U560  ( .A(_AES_ENC_us10_n929 ), .ZN(_AES_ENC_us10_n601 ) );
INV_X4 _AES_ENC_us10_U559  ( .A(_AES_ENC_us10_n1056 ), .ZN(_AES_ENC_us10_n600 ) );
INV_X4 _AES_ENC_us10_U558  ( .A(_AES_ENC_us10_n1054 ), .ZN(_AES_ENC_us10_n599 ) );
INV_X4 _AES_ENC_us10_U557  ( .A(_AES_ENC_us10_n881 ), .ZN(_AES_ENC_us10_n598 ) );
INV_X4 _AES_ENC_us10_U556  ( .A(_AES_ENC_us10_n926 ), .ZN(_AES_ENC_us10_n597 ) );
INV_X4 _AES_ENC_us10_U555  ( .A(_AES_ENC_us10_n977 ), .ZN(_AES_ENC_us10_n595 ) );
INV_X4 _AES_ENC_us10_U554  ( .A(_AES_ENC_us10_n1031 ), .ZN(_AES_ENC_us10_n594 ) );
INV_X4 _AES_ENC_us10_U553  ( .A(_AES_ENC_us10_n1103 ), .ZN(_AES_ENC_us10_n593 ) );
INV_X4 _AES_ENC_us10_U552  ( .A(_AES_ENC_us10_n1009 ), .ZN(_AES_ENC_us10_n592 ) );
INV_X4 _AES_ENC_us10_U551  ( .A(_AES_ENC_us10_n990 ), .ZN(_AES_ENC_us10_n591 ) );
INV_X4 _AES_ENC_us10_U550  ( .A(_AES_ENC_us10_n1058 ), .ZN(_AES_ENC_us10_n590 ) );
INV_X4 _AES_ENC_us10_U549  ( .A(_AES_ENC_us10_n1074 ), .ZN(_AES_ENC_us10_n589 ) );
INV_X4 _AES_ENC_us10_U548  ( .A(_AES_ENC_us10_n1053 ), .ZN(_AES_ENC_us10_n588 ) );
INV_X4 _AES_ENC_us10_U547  ( .A(_AES_ENC_us10_n826 ), .ZN(_AES_ENC_us10_n587 ) );
INV_X4 _AES_ENC_us10_U546  ( .A(_AES_ENC_us10_n992 ), .ZN(_AES_ENC_us10_n586 ) );
INV_X4 _AES_ENC_us10_U545  ( .A(_AES_ENC_us10_n821 ), .ZN(_AES_ENC_us10_n585 ) );
INV_X4 _AES_ENC_us10_U544  ( .A(_AES_ENC_us10_n910 ), .ZN(_AES_ENC_us10_n584 ) );
INV_X4 _AES_ENC_us10_U543  ( .A(_AES_ENC_us10_n906 ), .ZN(_AES_ENC_us10_n583 ) );
INV_X4 _AES_ENC_us10_U542  ( .A(_AES_ENC_us10_n880 ), .ZN(_AES_ENC_us10_n581 ) );
INV_X4 _AES_ENC_us10_U541  ( .A(_AES_ENC_us10_n1013 ), .ZN(_AES_ENC_us10_n580 ) );
INV_X4 _AES_ENC_us10_U540  ( .A(_AES_ENC_us10_n1092 ), .ZN(_AES_ENC_us10_n579 ) );
INV_X4 _AES_ENC_us10_U539  ( .A(_AES_ENC_us10_n824 ), .ZN(_AES_ENC_us10_n578 ) );
INV_X4 _AES_ENC_us10_U538  ( .A(_AES_ENC_us10_n1091 ), .ZN(_AES_ENC_us10_n577 ) );
INV_X4 _AES_ENC_us10_U537  ( .A(_AES_ENC_us10_n1080 ), .ZN(_AES_ENC_us10_n576 ) );
INV_X4 _AES_ENC_us10_U536  ( .A(_AES_ENC_us10_n959 ), .ZN(_AES_ENC_us10_n575 ) );
INV_X4 _AES_ENC_us10_U535  ( .A(_AES_ENC_sa10[0]), .ZN(_AES_ENC_us10_n574 ));
NOR2_X2 _AES_ENC_us10_U534  ( .A1(_AES_ENC_sa10[0]), .A2(_AES_ENC_sa10[6]),.ZN(_AES_ENC_us10_n1090 ) );
NOR2_X2 _AES_ENC_us10_U533  ( .A1(_AES_ENC_us10_n574 ), .A2(_AES_ENC_sa10[6]), .ZN(_AES_ENC_us10_n1070 ) );
NOR2_X2 _AES_ENC_us10_U532  ( .A1(_AES_ENC_sa10[4]), .A2(_AES_ENC_sa10[3]),.ZN(_AES_ENC_us10_n1025 ) );
INV_X4 _AES_ENC_us10_U531  ( .A(_AES_ENC_us10_n569 ), .ZN(_AES_ENC_us10_n572 ) );
NOR2_X2 _AES_ENC_us10_U530  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n765 ) );
NOR2_X2 _AES_ENC_us10_U529  ( .A1(_AES_ENC_sa10[4]), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n764 ) );
NOR2_X2 _AES_ENC_us10_U528  ( .A1(_AES_ENC_us10_n765 ), .A2(_AES_ENC_us10_n764 ), .ZN(_AES_ENC_us10_n766 ) );
NOR2_X2 _AES_ENC_us10_U527  ( .A1(_AES_ENC_us10_n766 ), .A2(_AES_ENC_us10_n575 ), .ZN(_AES_ENC_us10_n767 ) );
NOR3_X2 _AES_ENC_us10_U526  ( .A1(_AES_ENC_us10_n627 ), .A2(_AES_ENC_sa10[5]), .A3(_AES_ENC_us10_n704 ), .ZN(_AES_ENC_us10_n706 ));
NOR2_X2 _AES_ENC_us10_U525  ( .A1(_AES_ENC_us10_n1117 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n707 ) );
NOR2_X2 _AES_ENC_us10_U524  ( .A1(_AES_ENC_sa10[4]), .A2(_AES_ENC_us10_n579 ), .ZN(_AES_ENC_us10_n705 ) );
NOR3_X2 _AES_ENC_us10_U523  ( .A1(_AES_ENC_us10_n707 ), .A2(_AES_ENC_us10_n706 ), .A3(_AES_ENC_us10_n705 ), .ZN(_AES_ENC_us10_n713 ) );
INV_X4 _AES_ENC_us10_U522  ( .A(_AES_ENC_sa10[3]), .ZN(_AES_ENC_us10_n621 ));
NAND3_X2 _AES_ENC_us10_U521  ( .A1(_AES_ENC_us10_n652 ), .A2(_AES_ENC_us10_n626 ), .A3(_AES_ENC_sa10[7]), .ZN(_AES_ENC_us10_n653 ));
NOR2_X2 _AES_ENC_us10_U520  ( .A1(_AES_ENC_us10_n611 ), .A2(_AES_ENC_sa10[5]), .ZN(_AES_ENC_us10_n925 ) );
NOR2_X2 _AES_ENC_us10_U519  ( .A1(_AES_ENC_sa10[5]), .A2(_AES_ENC_sa10[2]),.ZN(_AES_ENC_us10_n974 ) );
INV_X4 _AES_ENC_us10_U518  ( .A(_AES_ENC_sa10[5]), .ZN(_AES_ENC_us10_n626 ));
NOR2_X2 _AES_ENC_us10_U517  ( .A1(_AES_ENC_us10_n611 ), .A2(_AES_ENC_sa10[7]), .ZN(_AES_ENC_us10_n779 ) );
NAND3_X2 _AES_ENC_us10_U516  ( .A1(_AES_ENC_us10_n679 ), .A2(_AES_ENC_us10_n678 ), .A3(_AES_ENC_us10_n677 ), .ZN(_AES_ENC_sa10_sub[0] ) );
NOR2_X2 _AES_ENC_us10_U515  ( .A1(_AES_ENC_us10_n626 ), .A2(_AES_ENC_sa10[2]), .ZN(_AES_ENC_us10_n1048 ) );
NOR4_X2 _AES_ENC_us10_U512  ( .A1(_AES_ENC_us10_n633 ), .A2(_AES_ENC_us10_n632 ), .A3(_AES_ENC_us10_n631 ), .A4(_AES_ENC_us10_n630 ), .ZN(_AES_ENC_us10_n634 ) );
NOR2_X2 _AES_ENC_us10_U510  ( .A1(_AES_ENC_us10_n629 ), .A2(_AES_ENC_us10_n628 ), .ZN(_AES_ENC_us10_n635 ) );
NAND3_X2 _AES_ENC_us10_U509  ( .A1(_AES_ENC_sa10[2]), .A2(_AES_ENC_sa10[7]), .A3(_AES_ENC_us10_n1059 ), .ZN(_AES_ENC_us10_n636 ) );
NOR2_X2 _AES_ENC_us10_U508  ( .A1(_AES_ENC_sa10[7]), .A2(_AES_ENC_sa10[2]),.ZN(_AES_ENC_us10_n794 ) );
NOR2_X2 _AES_ENC_us10_U507  ( .A1(_AES_ENC_sa10[4]), .A2(_AES_ENC_sa10[1]),.ZN(_AES_ENC_us10_n1102 ) );
NOR2_X2 _AES_ENC_us10_U506  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_sa10[3]), .ZN(_AES_ENC_us10_n1053 ) );
NOR2_X2 _AES_ENC_us10_U505  ( .A1(_AES_ENC_us10_n607 ), .A2(_AES_ENC_sa10[5]), .ZN(_AES_ENC_us10_n1024 ) );
NOR2_X2 _AES_ENC_us10_U504  ( .A1(_AES_ENC_us10_n625 ), .A2(_AES_ENC_sa10[2]), .ZN(_AES_ENC_us10_n1093 ) );
NOR2_X2 _AES_ENC_us10_U503  ( .A1(_AES_ENC_us10_n614 ), .A2(_AES_ENC_sa10[5]), .ZN(_AES_ENC_us10_n1094 ) );
NOR2_X2 _AES_ENC_us10_U502  ( .A1(_AES_ENC_us10_n624 ), .A2(_AES_ENC_sa10[3]), .ZN(_AES_ENC_us10_n931 ) );
INV_X4 _AES_ENC_us10_U501  ( .A(_AES_ENC_us10_n570 ), .ZN(_AES_ENC_us10_n573 ) );
NOR2_X2 _AES_ENC_us10_U500  ( .A1(_AES_ENC_us10_n1053 ), .A2(_AES_ENC_us10_n1095 ), .ZN(_AES_ENC_us10_n639 ) );
NOR3_X2 _AES_ENC_us10_U499  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n573 ), .A3(_AES_ENC_us10_n1074 ), .ZN(_AES_ENC_us10_n641 ) );
NOR2_X2 _AES_ENC_us10_U498  ( .A1(_AES_ENC_us10_n639 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n640 ) );
NOR2_X2 _AES_ENC_us10_U497  ( .A1(_AES_ENC_us10_n641 ), .A2(_AES_ENC_us10_n640 ), .ZN(_AES_ENC_us10_n646 ) );
NOR3_X2 _AES_ENC_us10_U496  ( .A1(_AES_ENC_us10_n995 ), .A2(_AES_ENC_us10_n586 ), .A3(_AES_ENC_us10_n994 ), .ZN(_AES_ENC_us10_n1002 ) );
NOR2_X2 _AES_ENC_us10_U495  ( .A1(_AES_ENC_us10_n909 ), .A2(_AES_ENC_us10_n908 ), .ZN(_AES_ENC_us10_n920 ) );
NOR2_X2 _AES_ENC_us10_U494  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n823 ) );
NOR2_X2 _AES_ENC_us10_U492  ( .A1(_AES_ENC_us10_n624 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n822 ) );
NOR2_X2 _AES_ENC_us10_U491  ( .A1(_AES_ENC_us10_n823 ), .A2(_AES_ENC_us10_n822 ), .ZN(_AES_ENC_us10_n825 ) );
NOR2_X2 _AES_ENC_us10_U490  ( .A1(_AES_ENC_sa10[1]), .A2(_AES_ENC_us10_n623 ), .ZN(_AES_ENC_us10_n913 ) );
NOR2_X2 _AES_ENC_us10_U489  ( .A1(_AES_ENC_us10_n913 ), .A2(_AES_ENC_us10_n1091 ), .ZN(_AES_ENC_us10_n914 ) );
NOR2_X2 _AES_ENC_us10_U488  ( .A1(_AES_ENC_us10_n826 ), .A2(_AES_ENC_us10_n572 ), .ZN(_AES_ENC_us10_n827 ) );
NOR3_X2 _AES_ENC_us10_U487  ( .A1(_AES_ENC_us10_n769 ), .A2(_AES_ENC_us10_n768 ), .A3(_AES_ENC_us10_n767 ), .ZN(_AES_ENC_us10_n775 ) );
NOR2_X2 _AES_ENC_us10_U486  ( .A1(_AES_ENC_us10_n1056 ), .A2(_AES_ENC_us10_n1053 ), .ZN(_AES_ENC_us10_n749 ) );
NOR2_X2 _AES_ENC_us10_U483  ( .A1(_AES_ENC_us10_n749 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n752 ) );
INV_X4 _AES_ENC_us10_U482  ( .A(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n596 ));
NOR2_X2 _AES_ENC_us10_U480  ( .A1(_AES_ENC_us10_n1054 ), .A2(_AES_ENC_us10_n1053 ), .ZN(_AES_ENC_us10_n1055 ) );
OR2_X4 _AES_ENC_us10_U479  ( .A1(_AES_ENC_us10_n1094 ), .A2(_AES_ENC_us10_n1093 ), .ZN(_AES_ENC_us10_n571 ) );
AND2_X2 _AES_ENC_us10_U478  ( .A1(_AES_ENC_us10_n571 ), .A2(_AES_ENC_us10_n1095 ), .ZN(_AES_ENC_us10_n1101 ) );
NOR2_X2 _AES_ENC_us10_U477  ( .A1(_AES_ENC_us10_n1074 ), .A2(_AES_ENC_us10_n931 ), .ZN(_AES_ENC_us10_n796 ) );
NOR2_X2 _AES_ENC_us10_U474  ( .A1(_AES_ENC_us10_n796 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n797 ) );
NOR2_X2 _AES_ENC_us10_U473  ( .A1(_AES_ENC_us10_n932 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n933 ) );
NOR2_X2 _AES_ENC_us10_U472  ( .A1(_AES_ENC_us10_n929 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n935 ) );
NOR2_X2 _AES_ENC_us10_U471  ( .A1(_AES_ENC_us10_n931 ), .A2(_AES_ENC_us10_n930 ), .ZN(_AES_ENC_us10_n934 ) );
NOR3_X2 _AES_ENC_us10_U470  ( .A1(_AES_ENC_us10_n935 ), .A2(_AES_ENC_us10_n934 ), .A3(_AES_ENC_us10_n933 ), .ZN(_AES_ENC_us10_n936 ) );
NOR2_X2 _AES_ENC_us10_U469  ( .A1(_AES_ENC_us10_n624 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n1075 ) );
NOR2_X2 _AES_ENC_us10_U468  ( .A1(_AES_ENC_us10_n572 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n949 ) );
NOR2_X2 _AES_ENC_us10_U467  ( .A1(_AES_ENC_us10_n1049 ), .A2(_AES_ENC_us10_n618 ), .ZN(_AES_ENC_us10_n1051 ) );
NOR2_X2 _AES_ENC_us10_U466  ( .A1(_AES_ENC_us10_n1051 ), .A2(_AES_ENC_us10_n1050 ), .ZN(_AES_ENC_us10_n1052 ) );
NOR2_X2 _AES_ENC_us10_U465  ( .A1(_AES_ENC_us10_n1052 ), .A2(_AES_ENC_us10_n592 ), .ZN(_AES_ENC_us10_n1064 ) );
NOR2_X2 _AES_ENC_us10_U464  ( .A1(_AES_ENC_sa10[1]), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n631 ) );
NOR2_X2 _AES_ENC_us10_U463  ( .A1(_AES_ENC_us10_n1025 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n980 ) );
NOR2_X2 _AES_ENC_us10_U462  ( .A1(_AES_ENC_us10_n1073 ), .A2(_AES_ENC_us10_n1094 ), .ZN(_AES_ENC_us10_n795 ) );
NOR2_X2 _AES_ENC_us10_U461  ( .A1(_AES_ENC_us10_n795 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n799 ) );
NOR2_X2 _AES_ENC_us10_U460  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n981 ) );
NOR2_X2 _AES_ENC_us10_U459  ( .A1(_AES_ENC_us10_n1102 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n643 ) );
NOR2_X2 _AES_ENC_us10_U458  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n621 ), .ZN(_AES_ENC_us10_n642 ) );
NOR2_X2 _AES_ENC_us10_U455  ( .A1(_AES_ENC_us10_n911 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n644 ) );
NOR4_X2 _AES_ENC_us10_U448  ( .A1(_AES_ENC_us10_n644 ), .A2(_AES_ENC_us10_n643 ), .A3(_AES_ENC_us10_n804 ), .A4(_AES_ENC_us10_n642 ), .ZN(_AES_ENC_us10_n645 ) );
NOR2_X2 _AES_ENC_us10_U447  ( .A1(_AES_ENC_us10_n1102 ), .A2(_AES_ENC_us10_n910 ), .ZN(_AES_ENC_us10_n932 ) );
NOR2_X2 _AES_ENC_us10_U442  ( .A1(_AES_ENC_us10_n1102 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n755 ) );
NOR2_X2 _AES_ENC_us10_U441  ( .A1(_AES_ENC_us10_n931 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n743 ) );
NOR2_X2 _AES_ENC_us10_U438  ( .A1(_AES_ENC_us10_n1072 ), .A2(_AES_ENC_us10_n1094 ), .ZN(_AES_ENC_us10_n930 ) );
NOR2_X2 _AES_ENC_us10_U435  ( .A1(_AES_ENC_us10_n1074 ), .A2(_AES_ENC_us10_n1025 ), .ZN(_AES_ENC_us10_n891 ) );
NOR2_X2 _AES_ENC_us10_U434  ( .A1(_AES_ENC_us10_n891 ), .A2(_AES_ENC_us10_n609 ), .ZN(_AES_ENC_us10_n894 ) );
NOR3_X2 _AES_ENC_us10_U433  ( .A1(_AES_ENC_us10_n623 ), .A2(_AES_ENC_sa10[1]), .A3(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n683 ));
INV_X4 _AES_ENC_us10_U428  ( .A(_AES_ENC_us10_n931 ), .ZN(_AES_ENC_us10_n623 ) );
NOR2_X2 _AES_ENC_us10_U427  ( .A1(_AES_ENC_us10_n996 ), .A2(_AES_ENC_us10_n931 ), .ZN(_AES_ENC_us10_n704 ) );
NOR2_X2 _AES_ENC_us10_U421  ( .A1(_AES_ENC_us10_n931 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n685 ) );
NOR2_X2 _AES_ENC_us10_U420  ( .A1(_AES_ENC_us10_n1029 ), .A2(_AES_ENC_us10_n1025 ), .ZN(_AES_ENC_us10_n1079 ) );
NOR3_X2 _AES_ENC_us10_U419  ( .A1(_AES_ENC_us10_n589 ), .A2(_AES_ENC_us10_n1025 ), .A3(_AES_ENC_us10_n616 ), .ZN(_AES_ENC_us10_n945 ) );
NOR2_X2 _AES_ENC_us10_U418  ( .A1(_AES_ENC_us10_n626 ), .A2(_AES_ENC_us10_n611 ), .ZN(_AES_ENC_us10_n800 ) );
NOR3_X2 _AES_ENC_us10_U417  ( .A1(_AES_ENC_us10_n590 ), .A2(_AES_ENC_us10_n627 ), .A3(_AES_ENC_us10_n611 ), .ZN(_AES_ENC_us10_n798 ) );
NOR3_X2 _AES_ENC_us10_U416  ( .A1(_AES_ENC_us10_n610 ), .A2(_AES_ENC_us10_n572 ), .A3(_AES_ENC_us10_n575 ), .ZN(_AES_ENC_us10_n962 ) );
NOR3_X2 _AES_ENC_us10_U415  ( .A1(_AES_ENC_us10_n959 ), .A2(_AES_ENC_us10_n572 ), .A3(_AES_ENC_us10_n609 ), .ZN(_AES_ENC_us10_n768 ) );
NOR3_X2 _AES_ENC_us10_U414  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n572 ), .A3(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n694 ) );
NOR3_X2 _AES_ENC_us10_U413  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n572 ), .A3(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n895 ) );
NOR3_X2 _AES_ENC_us10_U410  ( .A1(_AES_ENC_us10_n1008 ), .A2(_AES_ENC_us10_n1007 ), .A3(_AES_ENC_us10_n1006 ), .ZN(_AES_ENC_us10_n1018 ) );
NOR4_X2 _AES_ENC_us10_U409  ( .A1(_AES_ENC_us10_n806 ), .A2(_AES_ENC_us10_n805 ), .A3(_AES_ENC_us10_n804 ), .A4(_AES_ENC_us10_n803 ), .ZN(_AES_ENC_us10_n807 ) );
NOR3_X2 _AES_ENC_us10_U406  ( .A1(_AES_ENC_us10_n799 ), .A2(_AES_ENC_us10_n798 ), .A3(_AES_ENC_us10_n797 ), .ZN(_AES_ENC_us10_n808 ) );
NOR4_X2 _AES_ENC_us10_U405  ( .A1(_AES_ENC_us10_n843 ), .A2(_AES_ENC_us10_n842 ), .A3(_AES_ENC_us10_n841 ), .A4(_AES_ENC_us10_n840 ), .ZN(_AES_ENC_us10_n844 ) );
NOR2_X2 _AES_ENC_us10_U404  ( .A1(_AES_ENC_us10_n669 ), .A2(_AES_ENC_us10_n668 ), .ZN(_AES_ENC_us10_n673 ) );
NOR4_X2 _AES_ENC_us10_U403  ( .A1(_AES_ENC_us10_n946 ), .A2(_AES_ENC_us10_n1046 ), .A3(_AES_ENC_us10_n671 ), .A4(_AES_ENC_us10_n670 ), .ZN(_AES_ENC_us10_n672 ) );
NOR3_X2 _AES_ENC_us10_U401  ( .A1(_AES_ENC_us10_n1101 ), .A2(_AES_ENC_us10_n1100 ), .A3(_AES_ENC_us10_n1099 ), .ZN(_AES_ENC_us10_n1109 ) );
NOR4_X2 _AES_ENC_us10_U400  ( .A1(_AES_ENC_us10_n711 ), .A2(_AES_ENC_us10_n710 ), .A3(_AES_ENC_us10_n709 ), .A4(_AES_ENC_us10_n708 ), .ZN(_AES_ENC_us10_n712 ) );
NOR4_X2 _AES_ENC_us10_U399  ( .A1(_AES_ENC_us10_n963 ), .A2(_AES_ENC_us10_n962 ), .A3(_AES_ENC_us10_n961 ), .A4(_AES_ENC_us10_n960 ), .ZN(_AES_ENC_us10_n964 ) );
NOR3_X2 _AES_ENC_us10_U398  ( .A1(_AES_ENC_us10_n743 ), .A2(_AES_ENC_us10_n742 ), .A3(_AES_ENC_us10_n741 ), .ZN(_AES_ENC_us10_n744 ) );
NOR2_X2 _AES_ENC_us10_U397  ( .A1(_AES_ENC_us10_n697 ), .A2(_AES_ENC_us10_n658 ), .ZN(_AES_ENC_us10_n659 ) );
NOR2_X2 _AES_ENC_us10_U396  ( .A1(_AES_ENC_us10_n1078 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n1033 ) );
NOR2_X2 _AES_ENC_us10_U393  ( .A1(_AES_ENC_us10_n1031 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n1032 ) );
NOR3_X2 _AES_ENC_us10_U390  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n1025 ), .A3(_AES_ENC_us10_n1074 ), .ZN(_AES_ENC_us10_n1035 ) );
NOR4_X2 _AES_ENC_us10_U389  ( .A1(_AES_ENC_us10_n1035 ), .A2(_AES_ENC_us10_n1034 ), .A3(_AES_ENC_us10_n1033 ), .A4(_AES_ENC_us10_n1032 ), .ZN(_AES_ENC_us10_n1036 ) );
NOR2_X2 _AES_ENC_us10_U388  ( .A1(_AES_ENC_us10_n598 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n885 ) );
NOR2_X2 _AES_ENC_us10_U387  ( .A1(_AES_ENC_us10_n623 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n882 ) );
NOR2_X2 _AES_ENC_us10_U386  ( .A1(_AES_ENC_us10_n1053 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n884 ) );
NOR4_X2 _AES_ENC_us10_U385  ( .A1(_AES_ENC_us10_n885 ), .A2(_AES_ENC_us10_n884 ), .A3(_AES_ENC_us10_n883 ), .A4(_AES_ENC_us10_n882 ), .ZN(_AES_ENC_us10_n886 ) );
NOR2_X2 _AES_ENC_us10_U384  ( .A1(_AES_ENC_us10_n825 ), .A2(_AES_ENC_us10_n578 ), .ZN(_AES_ENC_us10_n830 ) );
NOR2_X2 _AES_ENC_us10_U383  ( .A1(_AES_ENC_us10_n827 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n829 ) );
NOR2_X2 _AES_ENC_us10_U382  ( .A1(_AES_ENC_us10_n572 ), .A2(_AES_ENC_us10_n579 ), .ZN(_AES_ENC_us10_n828 ) );
NOR4_X2 _AES_ENC_us10_U374  ( .A1(_AES_ENC_us10_n831 ), .A2(_AES_ENC_us10_n830 ), .A3(_AES_ENC_us10_n829 ), .A4(_AES_ENC_us10_n828 ), .ZN(_AES_ENC_us10_n832 ) );
NOR2_X2 _AES_ENC_us10_U373  ( .A1(_AES_ENC_us10_n606 ), .A2(_AES_ENC_us10_n582 ), .ZN(_AES_ENC_us10_n1104 ) );
NOR2_X2 _AES_ENC_us10_U372  ( .A1(_AES_ENC_us10_n1102 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n1106 ) );
NOR2_X2 _AES_ENC_us10_U370  ( .A1(_AES_ENC_us10_n1103 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n1105 ) );
NOR4_X2 _AES_ENC_us10_U369  ( .A1(_AES_ENC_us10_n1107 ), .A2(_AES_ENC_us10_n1106 ), .A3(_AES_ENC_us10_n1105 ), .A4(_AES_ENC_us10_n1104 ), .ZN(_AES_ENC_us10_n1108 ) );
NOR3_X2 _AES_ENC_us10_U368  ( .A1(_AES_ENC_us10_n959 ), .A2(_AES_ENC_us10_n621 ), .A3(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n963 ) );
NOR2_X2 _AES_ENC_us10_U367  ( .A1(_AES_ENC_us10_n626 ), .A2(_AES_ENC_us10_n627 ), .ZN(_AES_ENC_us10_n1114 ) );
INV_X4 _AES_ENC_us10_U366  ( .A(_AES_ENC_us10_n1024 ), .ZN(_AES_ENC_us10_n606 ) );
NOR3_X2 _AES_ENC_us10_U365  ( .A1(_AES_ENC_us10_n910 ), .A2(_AES_ENC_us10_n1059 ), .A3(_AES_ENC_us10_n611 ), .ZN(_AES_ENC_us10_n1115 ) );
INV_X4 _AES_ENC_us10_U364  ( .A(_AES_ENC_us10_n1094 ), .ZN(_AES_ENC_us10_n613 ) );
NOR2_X2 _AES_ENC_us10_U363  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n931 ), .ZN(_AES_ENC_us10_n1100 ) );
INV_X4 _AES_ENC_us10_U354  ( .A(_AES_ENC_us10_n1093 ), .ZN(_AES_ENC_us10_n617 ) );
NOR2_X2 _AES_ENC_us10_U353  ( .A1(_AES_ENC_us10_n569 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n929 ) );
NOR2_X2 _AES_ENC_us10_U352  ( .A1(_AES_ENC_us10_n620 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n926 ) );
NOR2_X2 _AES_ENC_us10_U351  ( .A1(_AES_ENC_us10_n572 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n1095 ) );
NOR2_X2 _AES_ENC_us10_U350  ( .A1(_AES_ENC_us10_n609 ), .A2(_AES_ENC_us10_n627 ), .ZN(_AES_ENC_us10_n1010 ) );
NOR2_X2 _AES_ENC_us10_U349  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n1103 ) );
NOR2_X2 _AES_ENC_us10_U348  ( .A1(_AES_ENC_us10_n622 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n1059 ) );
NOR2_X2 _AES_ENC_us10_U347  ( .A1(_AES_ENC_sa10[1]), .A2(_AES_ENC_us10_n1120 ), .ZN(_AES_ENC_us10_n1022 ) );
NOR2_X2 _AES_ENC_us10_U346  ( .A1(_AES_ENC_us10_n619 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n911 ) );
NOR2_X2 _AES_ENC_us10_U345  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_us10_n1025 ), .ZN(_AES_ENC_us10_n826 ) );
NOR2_X2 _AES_ENC_us10_U338  ( .A1(_AES_ENC_us10_n626 ), .A2(_AES_ENC_us10_n607 ), .ZN(_AES_ENC_us10_n1072 ) );
NOR2_X2 _AES_ENC_us10_U335  ( .A1(_AES_ENC_us10_n627 ), .A2(_AES_ENC_us10_n616 ), .ZN(_AES_ENC_us10_n956 ) );
NOR2_X2 _AES_ENC_us10_U329  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_us10_n624 ), .ZN(_AES_ENC_us10_n1121 ) );
NOR2_X2 _AES_ENC_us10_U328  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_us10_n624 ), .ZN(_AES_ENC_us10_n1058 ) );
NOR2_X2 _AES_ENC_us10_U327  ( .A1(_AES_ENC_us10_n625 ), .A2(_AES_ENC_us10_n611 ), .ZN(_AES_ENC_us10_n1073 ) );
NOR2_X2 _AES_ENC_us10_U325  ( .A1(_AES_ENC_sa10[1]), .A2(_AES_ENC_us10_n1025 ), .ZN(_AES_ENC_us10_n1054 ) );
NOR2_X2 _AES_ENC_us10_U324  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_us10_n931 ), .ZN(_AES_ENC_us10_n1029 ) );
NOR2_X2 _AES_ENC_us10_U319  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n1056 ) );
NOR2_X2 _AES_ENC_us10_U318  ( .A1(_AES_ENC_us10_n614 ), .A2(_AES_ENC_us10_n626 ), .ZN(_AES_ENC_us10_n1050 ) );
NOR2_X2 _AES_ENC_us10_U317  ( .A1(_AES_ENC_us10_n1121 ), .A2(_AES_ENC_us10_n1025 ), .ZN(_AES_ENC_us10_n1120 ) );
NOR2_X2 _AES_ENC_us10_U316  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_us10_n572 ), .ZN(_AES_ENC_us10_n1074 ) );
NOR2_X2 _AES_ENC_us10_U315  ( .A1(_AES_ENC_us10_n1058 ), .A2(_AES_ENC_us10_n1054 ), .ZN(_AES_ENC_us10_n878 ) );
NOR2_X2 _AES_ENC_us10_U314  ( .A1(_AES_ENC_us10_n878 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n879 ) );
NOR2_X2 _AES_ENC_us10_U312  ( .A1(_AES_ENC_us10_n880 ), .A2(_AES_ENC_us10_n879 ), .ZN(_AES_ENC_us10_n887 ) );
NOR2_X2 _AES_ENC_us10_U311  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n588 ), .ZN(_AES_ENC_us10_n957 ) );
NOR2_X2 _AES_ENC_us10_U310  ( .A1(_AES_ENC_us10_n958 ), .A2(_AES_ENC_us10_n957 ), .ZN(_AES_ENC_us10_n965 ) );
NOR3_X2 _AES_ENC_us10_U309  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n1091 ), .A3(_AES_ENC_us10_n1022 ), .ZN(_AES_ENC_us10_n720 ) );
NOR3_X2 _AES_ENC_us10_U303  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n1054 ), .A3(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n719 ) );
NOR2_X2 _AES_ENC_us10_U302  ( .A1(_AES_ENC_us10_n720 ), .A2(_AES_ENC_us10_n719 ), .ZN(_AES_ENC_us10_n726 ) );
NOR2_X2 _AES_ENC_us10_U300  ( .A1(_AES_ENC_us10_n614 ), .A2(_AES_ENC_us10_n591 ), .ZN(_AES_ENC_us10_n865 ) );
NOR2_X2 _AES_ENC_us10_U299  ( .A1(_AES_ENC_us10_n1059 ), .A2(_AES_ENC_us10_n1058 ), .ZN(_AES_ENC_us10_n1060 ) );
NOR2_X2 _AES_ENC_us10_U298  ( .A1(_AES_ENC_us10_n1095 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n668 ) );
NOR2_X2 _AES_ENC_us10_U297  ( .A1(_AES_ENC_us10_n911 ), .A2(_AES_ENC_us10_n910 ), .ZN(_AES_ENC_us10_n912 ) );
NOR2_X2 _AES_ENC_us10_U296  ( .A1(_AES_ENC_us10_n912 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n916 ) );
NOR2_X2 _AES_ENC_us10_U295  ( .A1(_AES_ENC_us10_n826 ), .A2(_AES_ENC_us10_n573 ), .ZN(_AES_ENC_us10_n750 ) );
NOR2_X2 _AES_ENC_us10_U294  ( .A1(_AES_ENC_us10_n750 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n751 ) );
NOR2_X2 _AES_ENC_us10_U293  ( .A1(_AES_ENC_us10_n907 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n908 ) );
NOR2_X2 _AES_ENC_us10_U292  ( .A1(_AES_ENC_us10_n990 ), .A2(_AES_ENC_us10_n926 ), .ZN(_AES_ENC_us10_n780 ) );
NOR2_X2 _AES_ENC_us10_U291  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n584 ), .ZN(_AES_ENC_us10_n838 ) );
NOR2_X2 _AES_ENC_us10_U290  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n602 ), .ZN(_AES_ENC_us10_n837 ) );
NOR2_X2 _AES_ENC_us10_U284  ( .A1(_AES_ENC_us10_n838 ), .A2(_AES_ENC_us10_n837 ), .ZN(_AES_ENC_us10_n845 ) );
NOR2_X2 _AES_ENC_us10_U283  ( .A1(_AES_ENC_us10_n1022 ), .A2(_AES_ENC_us10_n1058 ), .ZN(_AES_ENC_us10_n740 ) );
NOR2_X2 _AES_ENC_us10_U282  ( .A1(_AES_ENC_us10_n740 ), .A2(_AES_ENC_us10_n616 ), .ZN(_AES_ENC_us10_n742 ) );
NOR2_X2 _AES_ENC_us10_U281  ( .A1(_AES_ENC_us10_n1098 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n1099 ) );
NOR2_X2 _AES_ENC_us10_U280  ( .A1(_AES_ENC_us10_n1120 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n993 ) );
NOR2_X2 _AES_ENC_us10_U279  ( .A1(_AES_ENC_us10_n993 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n994 ) );
NOR2_X2 _AES_ENC_us10_U273  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n620 ), .ZN(_AES_ENC_us10_n1026 ) );
NOR2_X2 _AES_ENC_us10_U272  ( .A1(_AES_ENC_us10_n573 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n1027 ) );
NOR2_X2 _AES_ENC_us10_U271  ( .A1(_AES_ENC_us10_n1027 ), .A2(_AES_ENC_us10_n1026 ), .ZN(_AES_ENC_us10_n1028 ) );
NOR2_X2 _AES_ENC_us10_U270  ( .A1(_AES_ENC_us10_n1029 ), .A2(_AES_ENC_us10_n1028 ), .ZN(_AES_ENC_us10_n1034 ) );
NOR4_X2 _AES_ENC_us10_U269  ( .A1(_AES_ENC_us10_n757 ), .A2(_AES_ENC_us10_n756 ), .A3(_AES_ENC_us10_n755 ), .A4(_AES_ENC_us10_n754 ), .ZN(_AES_ENC_us10_n758 ) );
NOR2_X2 _AES_ENC_us10_U268  ( .A1(_AES_ENC_us10_n752 ), .A2(_AES_ENC_us10_n751 ), .ZN(_AES_ENC_us10_n759 ) );
NOR2_X2 _AES_ENC_us10_U267  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n1071 ), .ZN(_AES_ENC_us10_n669 ) );
NOR2_X2 _AES_ENC_us10_U263  ( .A1(_AES_ENC_us10_n1056 ), .A2(_AES_ENC_us10_n990 ), .ZN(_AES_ENC_us10_n991 ) );
NOR2_X2 _AES_ENC_us10_U262  ( .A1(_AES_ENC_us10_n991 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n995 ) );
NOR2_X2 _AES_ENC_us10_U258  ( .A1(_AES_ENC_us10_n607 ), .A2(_AES_ENC_us10_n590 ), .ZN(_AES_ENC_us10_n1008 ) );
NOR2_X2 _AES_ENC_us10_U255  ( .A1(_AES_ENC_us10_n839 ), .A2(_AES_ENC_us10_n582 ), .ZN(_AES_ENC_us10_n693 ) );
NOR2_X2 _AES_ENC_us10_U254  ( .A1(_AES_ENC_us10_n606 ), .A2(_AES_ENC_us10_n906 ), .ZN(_AES_ENC_us10_n741 ) );
NOR2_X2 _AES_ENC_us10_U253  ( .A1(_AES_ENC_us10_n1054 ), .A2(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n763 ) );
NOR2_X2 _AES_ENC_us10_U252  ( .A1(_AES_ENC_us10_n763 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n769 ) );
NOR2_X2 _AES_ENC_us10_U251  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n577 ), .ZN(_AES_ENC_us10_n1007 ) );
NOR2_X2 _AES_ENC_us10_U250  ( .A1(_AES_ENC_us10_n609 ), .A2(_AES_ENC_us10_n580 ), .ZN(_AES_ENC_us10_n1123 ) );
NOR2_X2 _AES_ENC_us10_U243  ( .A1(_AES_ENC_us10_n609 ), .A2(_AES_ENC_us10_n590 ), .ZN(_AES_ENC_us10_n710 ) );
INV_X4 _AES_ENC_us10_U242  ( .A(_AES_ENC_us10_n1029 ), .ZN(_AES_ENC_us10_n582 ) );
NOR2_X2 _AES_ENC_us10_U241  ( .A1(_AES_ENC_us10_n616 ), .A2(_AES_ENC_us10_n597 ), .ZN(_AES_ENC_us10_n883 ) );
NOR2_X2 _AES_ENC_us10_U240  ( .A1(_AES_ENC_us10_n593 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n1125 ) );
NOR2_X2 _AES_ENC_us10_U239  ( .A1(_AES_ENC_us10_n990 ), .A2(_AES_ENC_us10_n929 ), .ZN(_AES_ENC_us10_n892 ) );
NOR2_X2 _AES_ENC_us10_U238  ( .A1(_AES_ENC_us10_n892 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n893 ) );
NOR2_X2 _AES_ENC_us10_U237  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n602 ), .ZN(_AES_ENC_us10_n950 ) );
NOR2_X2 _AES_ENC_us10_U236  ( .A1(_AES_ENC_us10_n1079 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n1082 ) );
NOR2_X2 _AES_ENC_us10_U235  ( .A1(_AES_ENC_us10_n910 ), .A2(_AES_ENC_us10_n1056 ), .ZN(_AES_ENC_us10_n941 ) );
NOR2_X2 _AES_ENC_us10_U234  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n1077 ), .ZN(_AES_ENC_us10_n841 ) );
NOR2_X2 _AES_ENC_us10_U229  ( .A1(_AES_ENC_us10_n623 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n630 ) );
NOR2_X2 _AES_ENC_us10_U228  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n602 ), .ZN(_AES_ENC_us10_n806 ) );
NOR2_X2 _AES_ENC_us10_U227  ( .A1(_AES_ENC_us10_n623 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n948 ) );
NOR2_X2 _AES_ENC_us10_U226  ( .A1(_AES_ENC_us10_n606 ), .A2(_AES_ENC_us10_n589 ), .ZN(_AES_ENC_us10_n997 ) );
NOR2_X2 _AES_ENC_us10_U225  ( .A1(_AES_ENC_us10_n1121 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n1122 ) );
NOR2_X2 _AES_ENC_us10_U223  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n1023 ), .ZN(_AES_ENC_us10_n756 ) );
NOR2_X2 _AES_ENC_us10_U222  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n602 ), .ZN(_AES_ENC_us10_n870 ) );
NOR2_X2 _AES_ENC_us10_U221  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n569 ), .ZN(_AES_ENC_us10_n947 ) );
NOR2_X2 _AES_ENC_us10_U217  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n1077 ), .ZN(_AES_ENC_us10_n1084 ) );
NOR2_X2 _AES_ENC_us10_U213  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n855 ), .ZN(_AES_ENC_us10_n709 ) );
NOR2_X2 _AES_ENC_us10_U212  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n589 ), .ZN(_AES_ENC_us10_n868 ) );
NOR2_X2 _AES_ENC_us10_U211  ( .A1(_AES_ENC_us10_n1120 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n1124 ) );
NOR2_X2 _AES_ENC_us10_U210  ( .A1(_AES_ENC_us10_n1120 ), .A2(_AES_ENC_us10_n839 ), .ZN(_AES_ENC_us10_n842 ) );
NOR2_X2 _AES_ENC_us10_U209  ( .A1(_AES_ENC_us10_n1120 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n696 ) );
NOR2_X2 _AES_ENC_us10_U208  ( .A1(_AES_ENC_us10_n1074 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n1076 ) );
NOR2_X2 _AES_ENC_us10_U207  ( .A1(_AES_ENC_us10_n1074 ), .A2(_AES_ENC_us10_n620 ), .ZN(_AES_ENC_us10_n781 ) );
NOR3_X2 _AES_ENC_us10_U201  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n1056 ), .A3(_AES_ENC_us10_n990 ), .ZN(_AES_ENC_us10_n979 ) );
NOR3_X2 _AES_ENC_us10_U200  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n1058 ), .A3(_AES_ENC_us10_n1059 ), .ZN(_AES_ENC_us10_n854 ) );
NOR2_X2 _AES_ENC_us10_U199  ( .A1(_AES_ENC_us10_n996 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n869 ) );
NOR2_X2 _AES_ENC_us10_U198  ( .A1(_AES_ENC_us10_n1056 ), .A2(_AES_ENC_us10_n1074 ), .ZN(_AES_ENC_us10_n1057 ) );
NOR3_X2 _AES_ENC_us10_U197  ( .A1(_AES_ENC_us10_n607 ), .A2(_AES_ENC_us10_n1120 ), .A3(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n978 ) );
NOR2_X2 _AES_ENC_us10_U196  ( .A1(_AES_ENC_us10_n996 ), .A2(_AES_ENC_us10_n911 ), .ZN(_AES_ENC_us10_n1116 ) );
NOR2_X2 _AES_ENC_us10_U195  ( .A1(_AES_ENC_us10_n1074 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n754 ) );
NOR2_X2 _AES_ENC_us10_U194  ( .A1(_AES_ENC_us10_n926 ), .A2(_AES_ENC_us10_n1103 ), .ZN(_AES_ENC_us10_n977 ) );
NOR2_X2 _AES_ENC_us10_U187  ( .A1(_AES_ENC_us10_n839 ), .A2(_AES_ENC_us10_n824 ), .ZN(_AES_ENC_us10_n1092 ) );
NOR2_X2 _AES_ENC_us10_U186  ( .A1(_AES_ENC_us10_n573 ), .A2(_AES_ENC_us10_n1074 ), .ZN(_AES_ENC_us10_n684 ) );
NOR2_X2 _AES_ENC_us10_U185  ( .A1(_AES_ENC_us10_n826 ), .A2(_AES_ENC_us10_n1059 ), .ZN(_AES_ENC_us10_n907 ) );
NOR3_X2 _AES_ENC_us10_U184  ( .A1(_AES_ENC_us10_n625 ), .A2(_AES_ENC_us10_n1115 ), .A3(_AES_ENC_us10_n585 ), .ZN(_AES_ENC_us10_n831 ) );
NOR3_X2 _AES_ENC_us10_U183  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n1056 ), .A3(_AES_ENC_us10_n990 ), .ZN(_AES_ENC_us10_n896 ) );
NOR3_X2 _AES_ENC_us10_U182  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n573 ), .A3(_AES_ENC_us10_n1013 ), .ZN(_AES_ENC_us10_n670 ) );
NOR3_X2 _AES_ENC_us10_U181  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n1091 ), .A3(_AES_ENC_us10_n1022 ), .ZN(_AES_ENC_us10_n843 ) );
NOR2_X2 _AES_ENC_us10_U180  ( .A1(_AES_ENC_us10_n1029 ), .A2(_AES_ENC_us10_n1095 ), .ZN(_AES_ENC_us10_n735 ) );
NOR2_X2 _AES_ENC_us10_U174  ( .A1(_AES_ENC_us10_n1100 ), .A2(_AES_ENC_us10_n854 ), .ZN(_AES_ENC_us10_n860 ) );
NOR4_X2 _AES_ENC_us10_U173  ( .A1(_AES_ENC_us10_n1125 ), .A2(_AES_ENC_us10_n1124 ), .A3(_AES_ENC_us10_n1123 ), .A4(_AES_ENC_us10_n1122 ), .ZN(_AES_ENC_us10_n1126 ) );
NOR4_X2 _AES_ENC_us10_U172  ( .A1(_AES_ENC_us10_n1084 ), .A2(_AES_ENC_us10_n1083 ), .A3(_AES_ENC_us10_n1082 ), .A4(_AES_ENC_us10_n1081 ), .ZN(_AES_ENC_us10_n1085 ) );
NOR2_X2 _AES_ENC_us10_U171  ( .A1(_AES_ENC_us10_n1076 ), .A2(_AES_ENC_us10_n1075 ), .ZN(_AES_ENC_us10_n1086 ) );
NAND3_X2 _AES_ENC_us10_U170  ( .A1(_AES_ENC_us10_n569 ), .A2(_AES_ENC_us10_n582 ), .A3(_AES_ENC_us10_n681 ), .ZN(_AES_ENC_us10_n691 ) );
NOR2_X2 _AES_ENC_us10_U169  ( .A1(_AES_ENC_us10_n683 ), .A2(_AES_ENC_us10_n682 ), .ZN(_AES_ENC_us10_n690 ) );
NOR3_X2 _AES_ENC_us10_U168  ( .A1(_AES_ENC_us10_n695 ), .A2(_AES_ENC_us10_n694 ), .A3(_AES_ENC_us10_n693 ), .ZN(_AES_ENC_us10_n700 ) );
NOR4_X2 _AES_ENC_us10_U162  ( .A1(_AES_ENC_us10_n983 ), .A2(_AES_ENC_us10_n698 ), .A3(_AES_ENC_us10_n697 ), .A4(_AES_ENC_us10_n696 ), .ZN(_AES_ENC_us10_n699 ) );
NOR2_X2 _AES_ENC_us10_U161  ( .A1(_AES_ENC_us10_n946 ), .A2(_AES_ENC_us10_n945 ), .ZN(_AES_ENC_us10_n952 ) );
NOR4_X2 _AES_ENC_us10_U160  ( .A1(_AES_ENC_us10_n950 ), .A2(_AES_ENC_us10_n949 ), .A3(_AES_ENC_us10_n948 ), .A4(_AES_ENC_us10_n947 ), .ZN(_AES_ENC_us10_n951 ) );
NOR4_X2 _AES_ENC_us10_U159  ( .A1(_AES_ENC_us10_n983 ), .A2(_AES_ENC_us10_n982 ), .A3(_AES_ENC_us10_n981 ), .A4(_AES_ENC_us10_n980 ), .ZN(_AES_ENC_us10_n984 ) );
NOR2_X2 _AES_ENC_us10_U158  ( .A1(_AES_ENC_us10_n979 ), .A2(_AES_ENC_us10_n978 ), .ZN(_AES_ENC_us10_n985 ) );
NOR4_X2 _AES_ENC_us10_U157  ( .A1(_AES_ENC_us10_n896 ), .A2(_AES_ENC_us10_n895 ), .A3(_AES_ENC_us10_n894 ), .A4(_AES_ENC_us10_n893 ), .ZN(_AES_ENC_us10_n897 ) );
NOR2_X2 _AES_ENC_us10_U156  ( .A1(_AES_ENC_us10_n866 ), .A2(_AES_ENC_us10_n865 ), .ZN(_AES_ENC_us10_n872 ) );
NOR4_X2 _AES_ENC_us10_U155  ( .A1(_AES_ENC_us10_n870 ), .A2(_AES_ENC_us10_n869 ), .A3(_AES_ENC_us10_n868 ), .A4(_AES_ENC_us10_n867 ), .ZN(_AES_ENC_us10_n871 ) );
NOR3_X2 _AES_ENC_us10_U154  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n1054 ), .A3(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n961 ) );
NOR3_X2 _AES_ENC_us10_U153  ( .A1(_AES_ENC_us10_n620 ), .A2(_AES_ENC_us10_n1074 ), .A3(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n671 ) );
NOR2_X2 _AES_ENC_us10_U152  ( .A1(_AES_ENC_us10_n1057 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n1062 ) );
NOR2_X2 _AES_ENC_us10_U143  ( .A1(_AES_ENC_us10_n1055 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n1063 ) );
NOR2_X2 _AES_ENC_us10_U142  ( .A1(_AES_ENC_us10_n1060 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n1061 ) );
NOR4_X2 _AES_ENC_us10_U141  ( .A1(_AES_ENC_us10_n1064 ), .A2(_AES_ENC_us10_n1063 ), .A3(_AES_ENC_us10_n1062 ), .A4(_AES_ENC_us10_n1061 ), .ZN(_AES_ENC_us10_n1065 ) );
NOR3_X2 _AES_ENC_us10_U140  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n1120 ), .A3(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n918 ) );
NOR3_X2 _AES_ENC_us10_U132  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n573 ), .A3(_AES_ENC_us10_n1013 ), .ZN(_AES_ENC_us10_n917 ) );
NOR2_X2 _AES_ENC_us10_U131  ( .A1(_AES_ENC_us10_n914 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n915 ) );
NOR4_X2 _AES_ENC_us10_U130  ( .A1(_AES_ENC_us10_n918 ), .A2(_AES_ENC_us10_n917 ), .A3(_AES_ENC_us10_n916 ), .A4(_AES_ENC_us10_n915 ), .ZN(_AES_ENC_us10_n919 ) );
NOR2_X2 _AES_ENC_us10_U129  ( .A1(_AES_ENC_us10_n616 ), .A2(_AES_ENC_us10_n580 ), .ZN(_AES_ENC_us10_n771 ) );
NOR2_X2 _AES_ENC_us10_U128  ( .A1(_AES_ENC_us10_n1103 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n772 ) );
NOR2_X2 _AES_ENC_us10_U127  ( .A1(_AES_ENC_us10_n610 ), .A2(_AES_ENC_us10_n599 ), .ZN(_AES_ENC_us10_n773 ) );
NOR4_X2 _AES_ENC_us10_U126  ( .A1(_AES_ENC_us10_n773 ), .A2(_AES_ENC_us10_n772 ), .A3(_AES_ENC_us10_n771 ), .A4(_AES_ENC_us10_n770 ), .ZN(_AES_ENC_us10_n774 ) );
NOR2_X2 _AES_ENC_us10_U121  ( .A1(_AES_ENC_us10_n735 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n687 ) );
NOR2_X2 _AES_ENC_us10_U120  ( .A1(_AES_ENC_us10_n684 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n688 ) );
NOR2_X2 _AES_ENC_us10_U119  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n600 ), .ZN(_AES_ENC_us10_n686 ) );
NOR4_X2 _AES_ENC_us10_U118  ( .A1(_AES_ENC_us10_n688 ), .A2(_AES_ENC_us10_n687 ), .A3(_AES_ENC_us10_n686 ), .A4(_AES_ENC_us10_n685 ), .ZN(_AES_ENC_us10_n689 ) );
NOR2_X2 _AES_ENC_us10_U117  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n595 ), .ZN(_AES_ENC_us10_n858 ) );
NOR2_X2 _AES_ENC_us10_U116  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n855 ), .ZN(_AES_ENC_us10_n857 ) );
NOR2_X2 _AES_ENC_us10_U115  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n587 ), .ZN(_AES_ENC_us10_n856 ) );
NOR4_X2 _AES_ENC_us10_U106  ( .A1(_AES_ENC_us10_n858 ), .A2(_AES_ENC_us10_n857 ), .A3(_AES_ENC_us10_n856 ), .A4(_AES_ENC_us10_n958 ), .ZN(_AES_ENC_us10_n859 ) );
NOR2_X2 _AES_ENC_us10_U105  ( .A1(_AES_ENC_us10_n780 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n784 ) );
NOR2_X2 _AES_ENC_us10_U104  ( .A1(_AES_ENC_us10_n1117 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n782 ) );
NOR2_X2 _AES_ENC_us10_U103  ( .A1(_AES_ENC_us10_n781 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n783 ) );
NOR4_X2 _AES_ENC_us10_U102  ( .A1(_AES_ENC_us10_n880 ), .A2(_AES_ENC_us10_n784 ), .A3(_AES_ENC_us10_n783 ), .A4(_AES_ENC_us10_n782 ), .ZN(_AES_ENC_us10_n785 ) );
NOR2_X2 _AES_ENC_us10_U101  ( .A1(_AES_ENC_us10_n583 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n814 ) );
NOR2_X2 _AES_ENC_us10_U100  ( .A1(_AES_ENC_us10_n907 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n813 ) );
NOR3_X2 _AES_ENC_us10_U95  ( .A1(_AES_ENC_us10_n606 ), .A2(_AES_ENC_us10_n1058 ), .A3(_AES_ENC_us10_n1059 ), .ZN(_AES_ENC_us10_n815 ) );
NOR4_X2 _AES_ENC_us10_U94  ( .A1(_AES_ENC_us10_n815 ), .A2(_AES_ENC_us10_n814 ), .A3(_AES_ENC_us10_n813 ), .A4(_AES_ENC_us10_n812 ), .ZN(_AES_ENC_us10_n816 ) );
NOR2_X2 _AES_ENC_us10_U93  ( .A1(_AES_ENC_us10_n617 ), .A2(_AES_ENC_us10_n569 ), .ZN(_AES_ENC_us10_n721 ) );
NOR2_X2 _AES_ENC_us10_U92  ( .A1(_AES_ENC_us10_n1031 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n723 ) );
NOR2_X2 _AES_ENC_us10_U91  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n1096 ), .ZN(_AES_ENC_us10_n722 ) );
NOR4_X2 _AES_ENC_us10_U90  ( .A1(_AES_ENC_us10_n724 ), .A2(_AES_ENC_us10_n723 ), .A3(_AES_ENC_us10_n722 ), .A4(_AES_ENC_us10_n721 ), .ZN(_AES_ENC_us10_n725 ) );
NOR2_X2 _AES_ENC_us10_U89  ( .A1(_AES_ENC_us10_n911 ), .A2(_AES_ENC_us10_n990 ), .ZN(_AES_ENC_us10_n1009 ) );
NOR2_X2 _AES_ENC_us10_U88  ( .A1(_AES_ENC_us10_n1013 ), .A2(_AES_ENC_us10_n573 ), .ZN(_AES_ENC_us10_n1014 ) );
NOR2_X2 _AES_ENC_us10_U87  ( .A1(_AES_ENC_us10_n1014 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n1015 ) );
NOR4_X2 _AES_ENC_us10_U86  ( .A1(_AES_ENC_us10_n1016 ), .A2(_AES_ENC_us10_n1015 ), .A3(_AES_ENC_us10_n1119 ), .A4(_AES_ENC_us10_n1046 ), .ZN(_AES_ENC_us10_n1017 ) );
NOR2_X2 _AES_ENC_us10_U81  ( .A1(_AES_ENC_us10_n996 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n998 ) );
NOR2_X2 _AES_ENC_us10_U80  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n577 ), .ZN(_AES_ENC_us10_n1000 ) );
NOR2_X2 _AES_ENC_us10_U79  ( .A1(_AES_ENC_us10_n616 ), .A2(_AES_ENC_us10_n1096 ), .ZN(_AES_ENC_us10_n999 ) );
NOR4_X2 _AES_ENC_us10_U78  ( .A1(_AES_ENC_us10_n1000 ), .A2(_AES_ENC_us10_n999 ), .A3(_AES_ENC_us10_n998 ), .A4(_AES_ENC_us10_n997 ), .ZN(_AES_ENC_us10_n1001 ) );
NOR2_X2 _AES_ENC_us10_U74  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n1096 ), .ZN(_AES_ENC_us10_n697 ) );
NOR2_X2 _AES_ENC_us10_U73  ( .A1(_AES_ENC_us10_n620 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n958 ) );
NOR2_X2 _AES_ENC_us10_U72  ( .A1(_AES_ENC_us10_n911 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n983 ) );
NOR2_X2 _AES_ENC_us10_U71  ( .A1(_AES_ENC_us10_n1054 ), .A2(_AES_ENC_us10_n1103 ), .ZN(_AES_ENC_us10_n1031 ) );
INV_X4 _AES_ENC_us10_U65  ( .A(_AES_ENC_us10_n1050 ), .ZN(_AES_ENC_us10_n612 ) );
INV_X4 _AES_ENC_us10_U64  ( .A(_AES_ENC_us10_n1072 ), .ZN(_AES_ENC_us10_n605 ) );
INV_X4 _AES_ENC_us10_U63  ( .A(_AES_ENC_us10_n1073 ), .ZN(_AES_ENC_us10_n604 ) );
NOR2_X2 _AES_ENC_us10_U62  ( .A1(_AES_ENC_us10_n582 ), .A2(_AES_ENC_us10_n613 ), .ZN(_AES_ENC_us10_n880 ) );
NOR3_X2 _AES_ENC_us10_U61  ( .A1(_AES_ENC_us10_n826 ), .A2(_AES_ENC_us10_n1121 ), .A3(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n946 ) );
INV_X4 _AES_ENC_us10_U59  ( .A(_AES_ENC_us10_n1010 ), .ZN(_AES_ENC_us10_n608 ) );
NOR3_X2 _AES_ENC_us10_U58  ( .A1(_AES_ENC_us10_n573 ), .A2(_AES_ENC_us10_n1029 ), .A3(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n1119 ) );
INV_X4 _AES_ENC_us10_U57  ( .A(_AES_ENC_us10_n956 ), .ZN(_AES_ENC_us10_n615 ) );
NOR2_X2 _AES_ENC_us10_U50  ( .A1(_AES_ENC_us10_n623 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n1013 ) );
NOR2_X2 _AES_ENC_us10_U49  ( .A1(_AES_ENC_us10_n620 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n910 ) );
NOR2_X2 _AES_ENC_us10_U48  ( .A1(_AES_ENC_us10_n569 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n1091 ) );
NOR2_X2 _AES_ENC_us10_U47  ( .A1(_AES_ENC_us10_n622 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n990 ) );
NOR2_X2 _AES_ENC_us10_U46  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_us10_n1121 ), .ZN(_AES_ENC_us10_n996 ) );
NOR2_X2 _AES_ENC_us10_U45  ( .A1(_AES_ENC_us10_n610 ), .A2(_AES_ENC_us10_n600 ), .ZN(_AES_ENC_us10_n628 ) );
NOR2_X2 _AES_ENC_us10_U44  ( .A1(_AES_ENC_us10_n576 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n866 ) );
NOR2_X2 _AES_ENC_us10_U43  ( .A1(_AES_ENC_us10_n603 ), .A2(_AES_ENC_us10_n610 ), .ZN(_AES_ENC_us10_n1006 ) );
NOR2_X2 _AES_ENC_us10_U42  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n1117 ), .ZN(_AES_ENC_us10_n1118 ) );
NOR2_X2 _AES_ENC_us10_U41  ( .A1(_AES_ENC_us10_n1119 ), .A2(_AES_ENC_us10_n1118 ), .ZN(_AES_ENC_us10_n1127 ) );
NOR2_X2 _AES_ENC_us10_U36  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n594 ), .ZN(_AES_ENC_us10_n629 ) );
NOR2_X2 _AES_ENC_us10_U35  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n906 ), .ZN(_AES_ENC_us10_n909 ) );
NOR2_X2 _AES_ENC_us10_U34  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n597 ), .ZN(_AES_ENC_us10_n658 ) );
NOR2_X2 _AES_ENC_us10_U33  ( .A1(_AES_ENC_us10_n1116 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n695 ) );
NOR2_X2 _AES_ENC_us10_U32  ( .A1(_AES_ENC_us10_n1078 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n1083 ) );
NOR2_X2 _AES_ENC_us10_U31  ( .A1(_AES_ENC_us10_n941 ), .A2(_AES_ENC_us10_n608 ), .ZN(_AES_ENC_us10_n724 ) );
NOR2_X2 _AES_ENC_us10_U30  ( .A1(_AES_ENC_us10_n598 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n1107 ) );
NOR2_X2 _AES_ENC_us10_U29  ( .A1(_AES_ENC_us10_n576 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n840 ) );
NOR2_X2 _AES_ENC_us10_U24  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n593 ), .ZN(_AES_ENC_us10_n633 ) );
NOR2_X2 _AES_ENC_us10_U23  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n1080 ), .ZN(_AES_ENC_us10_n1081 ) );
NOR2_X2 _AES_ENC_us10_U21  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n1045 ), .ZN(_AES_ENC_us10_n812 ) );
NOR2_X2 _AES_ENC_us10_U20  ( .A1(_AES_ENC_us10_n1009 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n960 ) );
NOR2_X2 _AES_ENC_us10_U19  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n601 ), .ZN(_AES_ENC_us10_n982 ) );
NOR2_X2 _AES_ENC_us10_U18  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n594 ), .ZN(_AES_ENC_us10_n757 ) );
NOR2_X2 _AES_ENC_us10_U17  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n590 ), .ZN(_AES_ENC_us10_n698 ) );
NOR2_X2 _AES_ENC_us10_U16  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n619 ), .ZN(_AES_ENC_us10_n708 ) );
NOR2_X2 _AES_ENC_us10_U15  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n582 ), .ZN(_AES_ENC_us10_n770 ) );
NOR2_X2 _AES_ENC_us10_U10  ( .A1(_AES_ENC_us10_n619 ), .A2(_AES_ENC_us10_n604 ), .ZN(_AES_ENC_us10_n803 ) );
NOR2_X2 _AES_ENC_us10_U9  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n881 ), .ZN(_AES_ENC_us10_n711 ) );
NOR2_X2 _AES_ENC_us10_U8  ( .A1(_AES_ENC_us10_n615 ), .A2(_AES_ENC_us10_n582 ), .ZN(_AES_ENC_us10_n867 ) );
NOR2_X2 _AES_ENC_us10_U7  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n599 ), .ZN(_AES_ENC_us10_n804 ) );
NOR2_X2 _AES_ENC_us10_U6  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n620 ), .ZN(_AES_ENC_us10_n1046 ) );
OR2_X4 _AES_ENC_us10_U5  ( .A1(_AES_ENC_us10_n624 ), .A2(_AES_ENC_sa10[1]),.ZN(_AES_ENC_us10_n570 ) );
OR2_X4 _AES_ENC_us10_U4  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_sa10[4]),.ZN(_AES_ENC_us10_n569 ) );
NAND2_X2 _AES_ENC_us10_U514  ( .A1(_AES_ENC_us10_n1121 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n1030 ) );
AND2_X2 _AES_ENC_us10_U513  ( .A1(_AES_ENC_us10_n597 ), .A2(_AES_ENC_us10_n1030 ), .ZN(_AES_ENC_us10_n1049 ) );
NAND2_X2 _AES_ENC_us10_U511  ( .A1(_AES_ENC_us10_n1049 ), .A2(_AES_ENC_us10_n794 ), .ZN(_AES_ENC_us10_n637 ) );
AND2_X2 _AES_ENC_us10_U493  ( .A1(_AES_ENC_us10_n779 ), .A2(_AES_ENC_us10_n996 ), .ZN(_AES_ENC_us10_n632 ) );
NAND4_X2 _AES_ENC_us10_U485  ( .A1(_AES_ENC_us10_n637 ), .A2(_AES_ENC_us10_n636 ), .A3(_AES_ENC_us10_n635 ), .A4(_AES_ENC_us10_n634 ), .ZN(_AES_ENC_us10_n638 ) );
NAND2_X2 _AES_ENC_us10_U484  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n638 ), .ZN(_AES_ENC_us10_n679 ) );
NAND2_X2 _AES_ENC_us10_U481  ( .A1(_AES_ENC_us10_n1094 ), .A2(_AES_ENC_us10_n591 ), .ZN(_AES_ENC_us10_n648 ) );
NAND2_X2 _AES_ENC_us10_U476  ( .A1(_AES_ENC_us10_n601 ), .A2(_AES_ENC_us10_n590 ), .ZN(_AES_ENC_us10_n762 ) );
NAND2_X2 _AES_ENC_us10_U475  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n762 ), .ZN(_AES_ENC_us10_n647 ) );
NAND4_X2 _AES_ENC_us10_U457  ( .A1(_AES_ENC_us10_n648 ), .A2(_AES_ENC_us10_n647 ), .A3(_AES_ENC_us10_n646 ), .A4(_AES_ENC_us10_n645 ), .ZN(_AES_ENC_us10_n649 ) );
NAND2_X2 _AES_ENC_us10_U456  ( .A1(_AES_ENC_sa10[0]), .A2(_AES_ENC_us10_n649 ), .ZN(_AES_ENC_us10_n665 ) );
NAND2_X2 _AES_ENC_us10_U454  ( .A1(_AES_ENC_us10_n596 ), .A2(_AES_ENC_us10_n623 ), .ZN(_AES_ENC_us10_n855 ) );
NAND2_X2 _AES_ENC_us10_U453  ( .A1(_AES_ENC_us10_n587 ), .A2(_AES_ENC_us10_n855 ), .ZN(_AES_ENC_us10_n821 ) );
NAND2_X2 _AES_ENC_us10_U452  ( .A1(_AES_ENC_us10_n1093 ), .A2(_AES_ENC_us10_n821 ), .ZN(_AES_ENC_us10_n662 ) );
NAND2_X2 _AES_ENC_us10_U451  ( .A1(_AES_ENC_us10_n619 ), .A2(_AES_ENC_us10_n589 ), .ZN(_AES_ENC_us10_n650 ) );
NAND2_X2 _AES_ENC_us10_U450  ( .A1(_AES_ENC_us10_n956 ), .A2(_AES_ENC_us10_n650 ), .ZN(_AES_ENC_us10_n661 ) );
NAND2_X2 _AES_ENC_us10_U449  ( .A1(_AES_ENC_us10_n626 ), .A2(_AES_ENC_us10_n627 ), .ZN(_AES_ENC_us10_n839 ) );
OR2_X2 _AES_ENC_us10_U446  ( .A1(_AES_ENC_us10_n839 ), .A2(_AES_ENC_us10_n932 ), .ZN(_AES_ENC_us10_n656 ) );
NAND2_X2 _AES_ENC_us10_U445  ( .A1(_AES_ENC_us10_n621 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n1096 ) );
NAND2_X2 _AES_ENC_us10_U444  ( .A1(_AES_ENC_us10_n1030 ), .A2(_AES_ENC_us10_n1096 ), .ZN(_AES_ENC_us10_n651 ) );
NAND2_X2 _AES_ENC_us10_U443  ( .A1(_AES_ENC_us10_n1114 ), .A2(_AES_ENC_us10_n651 ), .ZN(_AES_ENC_us10_n655 ) );
OR3_X2 _AES_ENC_us10_U440  ( .A1(_AES_ENC_us10_n1079 ), .A2(_AES_ENC_sa10[7]), .A3(_AES_ENC_us10_n626 ), .ZN(_AES_ENC_us10_n654 ));
NAND2_X2 _AES_ENC_us10_U439  ( .A1(_AES_ENC_us10_n593 ), .A2(_AES_ENC_us10_n601 ), .ZN(_AES_ENC_us10_n652 ) );
NAND4_X2 _AES_ENC_us10_U437  ( .A1(_AES_ENC_us10_n656 ), .A2(_AES_ENC_us10_n655 ), .A3(_AES_ENC_us10_n654 ), .A4(_AES_ENC_us10_n653 ), .ZN(_AES_ENC_us10_n657 ) );
NAND2_X2 _AES_ENC_us10_U436  ( .A1(_AES_ENC_sa10[2]), .A2(_AES_ENC_us10_n657 ), .ZN(_AES_ENC_us10_n660 ) );
NAND4_X2 _AES_ENC_us10_U432  ( .A1(_AES_ENC_us10_n662 ), .A2(_AES_ENC_us10_n661 ), .A3(_AES_ENC_us10_n660 ), .A4(_AES_ENC_us10_n659 ), .ZN(_AES_ENC_us10_n663 ) );
NAND2_X2 _AES_ENC_us10_U431  ( .A1(_AES_ENC_us10_n663 ), .A2(_AES_ENC_us10_n574 ), .ZN(_AES_ENC_us10_n664 ) );
NAND2_X2 _AES_ENC_us10_U430  ( .A1(_AES_ENC_us10_n665 ), .A2(_AES_ENC_us10_n664 ), .ZN(_AES_ENC_us10_n666 ) );
NAND2_X2 _AES_ENC_us10_U429  ( .A1(_AES_ENC_sa10[6]), .A2(_AES_ENC_us10_n666 ), .ZN(_AES_ENC_us10_n678 ) );
NAND2_X2 _AES_ENC_us10_U426  ( .A1(_AES_ENC_us10_n735 ), .A2(_AES_ENC_us10_n1093 ), .ZN(_AES_ENC_us10_n675 ) );
NAND2_X2 _AES_ENC_us10_U425  ( .A1(_AES_ENC_us10_n588 ), .A2(_AES_ENC_us10_n597 ), .ZN(_AES_ENC_us10_n1045 ) );
OR2_X2 _AES_ENC_us10_U424  ( .A1(_AES_ENC_us10_n1045 ), .A2(_AES_ENC_us10_n605 ), .ZN(_AES_ENC_us10_n674 ) );
NAND2_X2 _AES_ENC_us10_U423  ( .A1(_AES_ENC_sa10[1]), .A2(_AES_ENC_us10_n620 ), .ZN(_AES_ENC_us10_n667 ) );
NAND2_X2 _AES_ENC_us10_U422  ( .A1(_AES_ENC_us10_n619 ), .A2(_AES_ENC_us10_n667 ), .ZN(_AES_ENC_us10_n1071 ) );
NAND4_X2 _AES_ENC_us10_U412  ( .A1(_AES_ENC_us10_n675 ), .A2(_AES_ENC_us10_n674 ), .A3(_AES_ENC_us10_n673 ), .A4(_AES_ENC_us10_n672 ), .ZN(_AES_ENC_us10_n676 ) );
NAND2_X2 _AES_ENC_us10_U411  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n676 ), .ZN(_AES_ENC_us10_n677 ) );
NAND2_X2 _AES_ENC_us10_U408  ( .A1(_AES_ENC_us10_n800 ), .A2(_AES_ENC_us10_n1022 ), .ZN(_AES_ENC_us10_n680 ) );
NAND2_X2 _AES_ENC_us10_U407  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n680 ), .ZN(_AES_ENC_us10_n681 ) );
AND2_X2 _AES_ENC_us10_U402  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n684 ), .ZN(_AES_ENC_us10_n682 ) );
NAND4_X2 _AES_ENC_us10_U395  ( .A1(_AES_ENC_us10_n691 ), .A2(_AES_ENC_us10_n581 ), .A3(_AES_ENC_us10_n690 ), .A4(_AES_ENC_us10_n689 ), .ZN(_AES_ENC_us10_n692 ) );
NAND2_X2 _AES_ENC_us10_U394  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n692 ), .ZN(_AES_ENC_us10_n733 ) );
NAND2_X2 _AES_ENC_us10_U392  ( .A1(_AES_ENC_us10_n977 ), .A2(_AES_ENC_us10_n1050 ), .ZN(_AES_ENC_us10_n702 ) );
NAND2_X2 _AES_ENC_us10_U391  ( .A1(_AES_ENC_us10_n1093 ), .A2(_AES_ENC_us10_n1045 ), .ZN(_AES_ENC_us10_n701 ) );
NAND4_X2 _AES_ENC_us10_U381  ( .A1(_AES_ENC_us10_n702 ), .A2(_AES_ENC_us10_n701 ), .A3(_AES_ENC_us10_n700 ), .A4(_AES_ENC_us10_n699 ), .ZN(_AES_ENC_us10_n703 ) );
NAND2_X2 _AES_ENC_us10_U380  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n703 ), .ZN(_AES_ENC_us10_n732 ) );
AND2_X2 _AES_ENC_us10_U379  ( .A1(_AES_ENC_sa10[0]), .A2(_AES_ENC_sa10[6]),.ZN(_AES_ENC_us10_n1113 ) );
NAND2_X2 _AES_ENC_us10_U378  ( .A1(_AES_ENC_us10_n601 ), .A2(_AES_ENC_us10_n1030 ), .ZN(_AES_ENC_us10_n881 ) );
NAND2_X2 _AES_ENC_us10_U377  ( .A1(_AES_ENC_us10_n1093 ), .A2(_AES_ENC_us10_n881 ), .ZN(_AES_ENC_us10_n715 ) );
NAND2_X2 _AES_ENC_us10_U376  ( .A1(_AES_ENC_us10_n1010 ), .A2(_AES_ENC_us10_n600 ), .ZN(_AES_ENC_us10_n714 ) );
NAND2_X2 _AES_ENC_us10_U375  ( .A1(_AES_ENC_us10_n855 ), .A2(_AES_ENC_us10_n588 ), .ZN(_AES_ENC_us10_n1117 ) );
XNOR2_X2 _AES_ENC_us10_U371  ( .A(_AES_ENC_us10_n611 ), .B(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n824 ) );
NAND4_X2 _AES_ENC_us10_U362  ( .A1(_AES_ENC_us10_n715 ), .A2(_AES_ENC_us10_n714 ), .A3(_AES_ENC_us10_n713 ), .A4(_AES_ENC_us10_n712 ), .ZN(_AES_ENC_us10_n716 ) );
NAND2_X2 _AES_ENC_us10_U361  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n716 ), .ZN(_AES_ENC_us10_n731 ) );
AND2_X2 _AES_ENC_us10_U360  ( .A1(_AES_ENC_sa10[6]), .A2(_AES_ENC_us10_n574 ), .ZN(_AES_ENC_us10_n1131 ) );
NAND2_X2 _AES_ENC_us10_U359  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n717 ) );
NAND2_X2 _AES_ENC_us10_U358  ( .A1(_AES_ENC_us10_n1029 ), .A2(_AES_ENC_us10_n717 ), .ZN(_AES_ENC_us10_n728 ) );
NAND2_X2 _AES_ENC_us10_U357  ( .A1(_AES_ENC_sa10[1]), .A2(_AES_ENC_us10_n624 ), .ZN(_AES_ENC_us10_n1097 ) );
NAND2_X2 _AES_ENC_us10_U356  ( .A1(_AES_ENC_us10_n603 ), .A2(_AES_ENC_us10_n1097 ), .ZN(_AES_ENC_us10_n718 ) );
NAND2_X2 _AES_ENC_us10_U355  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n718 ), .ZN(_AES_ENC_us10_n727 ) );
NAND4_X2 _AES_ENC_us10_U344  ( .A1(_AES_ENC_us10_n728 ), .A2(_AES_ENC_us10_n727 ), .A3(_AES_ENC_us10_n726 ), .A4(_AES_ENC_us10_n725 ), .ZN(_AES_ENC_us10_n729 ) );
NAND2_X2 _AES_ENC_us10_U343  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n729 ), .ZN(_AES_ENC_us10_n730 ) );
NAND4_X2 _AES_ENC_us10_U342  ( .A1(_AES_ENC_us10_n733 ), .A2(_AES_ENC_us10_n732 ), .A3(_AES_ENC_us10_n731 ), .A4(_AES_ENC_us10_n730 ), .ZN(_AES_ENC_sa10_sub[1] ) );
NAND2_X2 _AES_ENC_us10_U341  ( .A1(_AES_ENC_sa10[7]), .A2(_AES_ENC_us10_n611 ), .ZN(_AES_ENC_us10_n734 ) );
NAND2_X2 _AES_ENC_us10_U340  ( .A1(_AES_ENC_us10_n734 ), .A2(_AES_ENC_us10_n607 ), .ZN(_AES_ENC_us10_n738 ) );
OR4_X2 _AES_ENC_us10_U339  ( .A1(_AES_ENC_us10_n738 ), .A2(_AES_ENC_us10_n626 ), .A3(_AES_ENC_us10_n826 ), .A4(_AES_ENC_us10_n1121 ), .ZN(_AES_ENC_us10_n746 ) );
NAND2_X2 _AES_ENC_us10_U337  ( .A1(_AES_ENC_us10_n1100 ), .A2(_AES_ENC_us10_n587 ), .ZN(_AES_ENC_us10_n992 ) );
OR2_X2 _AES_ENC_us10_U336  ( .A1(_AES_ENC_us10_n610 ), .A2(_AES_ENC_us10_n735 ), .ZN(_AES_ENC_us10_n737 ) );
NAND2_X2 _AES_ENC_us10_U334  ( .A1(_AES_ENC_us10_n619 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n753 ) );
NAND2_X2 _AES_ENC_us10_U333  ( .A1(_AES_ENC_us10_n582 ), .A2(_AES_ENC_us10_n753 ), .ZN(_AES_ENC_us10_n1080 ) );
NAND2_X2 _AES_ENC_us10_U332  ( .A1(_AES_ENC_us10_n1048 ), .A2(_AES_ENC_us10_n576 ), .ZN(_AES_ENC_us10_n736 ) );
NAND2_X2 _AES_ENC_us10_U331  ( .A1(_AES_ENC_us10_n737 ), .A2(_AES_ENC_us10_n736 ), .ZN(_AES_ENC_us10_n739 ) );
NAND2_X2 _AES_ENC_us10_U330  ( .A1(_AES_ENC_us10_n739 ), .A2(_AES_ENC_us10_n738 ), .ZN(_AES_ENC_us10_n745 ) );
NAND2_X2 _AES_ENC_us10_U326  ( .A1(_AES_ENC_us10_n1096 ), .A2(_AES_ENC_us10_n590 ), .ZN(_AES_ENC_us10_n906 ) );
NAND4_X2 _AES_ENC_us10_U323  ( .A1(_AES_ENC_us10_n746 ), .A2(_AES_ENC_us10_n992 ), .A3(_AES_ENC_us10_n745 ), .A4(_AES_ENC_us10_n744 ), .ZN(_AES_ENC_us10_n747 ) );
NAND2_X2 _AES_ENC_us10_U322  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n747 ), .ZN(_AES_ENC_us10_n793 ) );
NAND2_X2 _AES_ENC_us10_U321  ( .A1(_AES_ENC_us10_n584 ), .A2(_AES_ENC_us10_n855 ), .ZN(_AES_ENC_us10_n748 ) );
NAND2_X2 _AES_ENC_us10_U320  ( .A1(_AES_ENC_us10_n956 ), .A2(_AES_ENC_us10_n748 ), .ZN(_AES_ENC_us10_n760 ) );
NAND2_X2 _AES_ENC_us10_U313  ( .A1(_AES_ENC_us10_n590 ), .A2(_AES_ENC_us10_n753 ), .ZN(_AES_ENC_us10_n1023 ) );
NAND4_X2 _AES_ENC_us10_U308  ( .A1(_AES_ENC_us10_n760 ), .A2(_AES_ENC_us10_n992 ), .A3(_AES_ENC_us10_n759 ), .A4(_AES_ENC_us10_n758 ), .ZN(_AES_ENC_us10_n761 ) );
NAND2_X2 _AES_ENC_us10_U307  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n761 ), .ZN(_AES_ENC_us10_n792 ) );
NAND2_X2 _AES_ENC_us10_U306  ( .A1(_AES_ENC_us10_n584 ), .A2(_AES_ENC_us10_n603 ), .ZN(_AES_ENC_us10_n989 ) );
NAND2_X2 _AES_ENC_us10_U305  ( .A1(_AES_ENC_us10_n1050 ), .A2(_AES_ENC_us10_n989 ), .ZN(_AES_ENC_us10_n777 ) );
NAND2_X2 _AES_ENC_us10_U304  ( .A1(_AES_ENC_us10_n1093 ), .A2(_AES_ENC_us10_n762 ), .ZN(_AES_ENC_us10_n776 ) );
XNOR2_X2 _AES_ENC_us10_U301  ( .A(_AES_ENC_sa10[7]), .B(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n959 ) );
NAND4_X2 _AES_ENC_us10_U289  ( .A1(_AES_ENC_us10_n777 ), .A2(_AES_ENC_us10_n776 ), .A3(_AES_ENC_us10_n775 ), .A4(_AES_ENC_us10_n774 ), .ZN(_AES_ENC_us10_n778 ) );
NAND2_X2 _AES_ENC_us10_U288  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n778 ), .ZN(_AES_ENC_us10_n791 ) );
NAND2_X2 _AES_ENC_us10_U287  ( .A1(_AES_ENC_us10_n1056 ), .A2(_AES_ENC_us10_n1050 ), .ZN(_AES_ENC_us10_n788 ) );
NAND2_X2 _AES_ENC_us10_U286  ( .A1(_AES_ENC_us10_n1091 ), .A2(_AES_ENC_us10_n779 ), .ZN(_AES_ENC_us10_n787 ) );
NAND2_X2 _AES_ENC_us10_U285  ( .A1(_AES_ENC_us10_n956 ), .A2(_AES_ENC_sa10[1]), .ZN(_AES_ENC_us10_n786 ) );
NAND4_X2 _AES_ENC_us10_U278  ( .A1(_AES_ENC_us10_n788 ), .A2(_AES_ENC_us10_n787 ), .A3(_AES_ENC_us10_n786 ), .A4(_AES_ENC_us10_n785 ), .ZN(_AES_ENC_us10_n789 ) );
NAND2_X2 _AES_ENC_us10_U277  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n789 ), .ZN(_AES_ENC_us10_n790 ) );
NAND4_X2 _AES_ENC_us10_U276  ( .A1(_AES_ENC_us10_n793 ), .A2(_AES_ENC_us10_n792 ), .A3(_AES_ENC_us10_n791 ), .A4(_AES_ENC_us10_n790 ), .ZN(_AES_ENC_sa10_sub[2] ) );
NAND2_X2 _AES_ENC_us10_U275  ( .A1(_AES_ENC_us10_n1059 ), .A2(_AES_ENC_us10_n794 ), .ZN(_AES_ENC_us10_n810 ) );
NAND2_X2 _AES_ENC_us10_U274  ( .A1(_AES_ENC_us10_n1049 ), .A2(_AES_ENC_us10_n956 ), .ZN(_AES_ENC_us10_n809 ) );
OR2_X2 _AES_ENC_us10_U266  ( .A1(_AES_ENC_us10_n1096 ), .A2(_AES_ENC_us10_n606 ), .ZN(_AES_ENC_us10_n802 ) );
NAND2_X2 _AES_ENC_us10_U265  ( .A1(_AES_ENC_us10_n1053 ), .A2(_AES_ENC_us10_n800 ), .ZN(_AES_ENC_us10_n801 ) );
NAND2_X2 _AES_ENC_us10_U264  ( .A1(_AES_ENC_us10_n802 ), .A2(_AES_ENC_us10_n801 ), .ZN(_AES_ENC_us10_n805 ) );
NAND4_X2 _AES_ENC_us10_U261  ( .A1(_AES_ENC_us10_n810 ), .A2(_AES_ENC_us10_n809 ), .A3(_AES_ENC_us10_n808 ), .A4(_AES_ENC_us10_n807 ), .ZN(_AES_ENC_us10_n811 ) );
NAND2_X2 _AES_ENC_us10_U260  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n811 ), .ZN(_AES_ENC_us10_n852 ) );
OR2_X2 _AES_ENC_us10_U259  ( .A1(_AES_ENC_us10_n1023 ), .A2(_AES_ENC_us10_n617 ), .ZN(_AES_ENC_us10_n819 ) );
OR2_X2 _AES_ENC_us10_U257  ( .A1(_AES_ENC_us10_n570 ), .A2(_AES_ENC_us10_n930 ), .ZN(_AES_ENC_us10_n818 ) );
NAND2_X2 _AES_ENC_us10_U256  ( .A1(_AES_ENC_us10_n1013 ), .A2(_AES_ENC_us10_n1094 ), .ZN(_AES_ENC_us10_n817 ) );
NAND4_X2 _AES_ENC_us10_U249  ( .A1(_AES_ENC_us10_n819 ), .A2(_AES_ENC_us10_n818 ), .A3(_AES_ENC_us10_n817 ), .A4(_AES_ENC_us10_n816 ), .ZN(_AES_ENC_us10_n820 ) );
NAND2_X2 _AES_ENC_us10_U248  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n820 ), .ZN(_AES_ENC_us10_n851 ) );
NAND2_X2 _AES_ENC_us10_U247  ( .A1(_AES_ENC_us10_n956 ), .A2(_AES_ENC_us10_n1080 ), .ZN(_AES_ENC_us10_n835 ) );
NAND2_X2 _AES_ENC_us10_U246  ( .A1(_AES_ENC_us10_n570 ), .A2(_AES_ENC_us10_n1030 ), .ZN(_AES_ENC_us10_n1047 ) );
OR2_X2 _AES_ENC_us10_U245  ( .A1(_AES_ENC_us10_n1047 ), .A2(_AES_ENC_us10_n612 ), .ZN(_AES_ENC_us10_n834 ) );
NAND2_X2 _AES_ENC_us10_U244  ( .A1(_AES_ENC_us10_n1072 ), .A2(_AES_ENC_us10_n589 ), .ZN(_AES_ENC_us10_n833 ) );
NAND4_X2 _AES_ENC_us10_U233  ( .A1(_AES_ENC_us10_n835 ), .A2(_AES_ENC_us10_n834 ), .A3(_AES_ENC_us10_n833 ), .A4(_AES_ENC_us10_n832 ), .ZN(_AES_ENC_us10_n836 ) );
NAND2_X2 _AES_ENC_us10_U232  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n836 ), .ZN(_AES_ENC_us10_n850 ) );
NAND2_X2 _AES_ENC_us10_U231  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n623 ), .ZN(_AES_ENC_us10_n847 ) );
NAND2_X2 _AES_ENC_us10_U230  ( .A1(_AES_ENC_us10_n1050 ), .A2(_AES_ENC_us10_n1071 ), .ZN(_AES_ENC_us10_n846 ) );
OR2_X2 _AES_ENC_us10_U224  ( .A1(_AES_ENC_us10_n1053 ), .A2(_AES_ENC_us10_n911 ), .ZN(_AES_ENC_us10_n1077 ) );
NAND4_X2 _AES_ENC_us10_U220  ( .A1(_AES_ENC_us10_n847 ), .A2(_AES_ENC_us10_n846 ), .A3(_AES_ENC_us10_n845 ), .A4(_AES_ENC_us10_n844 ), .ZN(_AES_ENC_us10_n848 ) );
NAND2_X2 _AES_ENC_us10_U219  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n848 ), .ZN(_AES_ENC_us10_n849 ) );
NAND4_X2 _AES_ENC_us10_U218  ( .A1(_AES_ENC_us10_n852 ), .A2(_AES_ENC_us10_n851 ), .A3(_AES_ENC_us10_n850 ), .A4(_AES_ENC_us10_n849 ), .ZN(_AES_ENC_sa10_sub[3] ) );
NAND2_X2 _AES_ENC_us10_U216  ( .A1(_AES_ENC_us10_n1009 ), .A2(_AES_ENC_us10_n1072 ), .ZN(_AES_ENC_us10_n862 ) );
NAND2_X2 _AES_ENC_us10_U215  ( .A1(_AES_ENC_us10_n603 ), .A2(_AES_ENC_us10_n577 ), .ZN(_AES_ENC_us10_n853 ) );
NAND2_X2 _AES_ENC_us10_U214  ( .A1(_AES_ENC_us10_n1050 ), .A2(_AES_ENC_us10_n853 ), .ZN(_AES_ENC_us10_n861 ) );
NAND4_X2 _AES_ENC_us10_U206  ( .A1(_AES_ENC_us10_n862 ), .A2(_AES_ENC_us10_n861 ), .A3(_AES_ENC_us10_n860 ), .A4(_AES_ENC_us10_n859 ), .ZN(_AES_ENC_us10_n863 ) );
NAND2_X2 _AES_ENC_us10_U205  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n863 ), .ZN(_AES_ENC_us10_n905 ) );
NAND2_X2 _AES_ENC_us10_U204  ( .A1(_AES_ENC_us10_n1010 ), .A2(_AES_ENC_us10_n989 ), .ZN(_AES_ENC_us10_n874 ) );
NAND2_X2 _AES_ENC_us10_U203  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n610 ), .ZN(_AES_ENC_us10_n864 ) );
NAND2_X2 _AES_ENC_us10_U202  ( .A1(_AES_ENC_us10_n929 ), .A2(_AES_ENC_us10_n864 ), .ZN(_AES_ENC_us10_n873 ) );
NAND4_X2 _AES_ENC_us10_U193  ( .A1(_AES_ENC_us10_n874 ), .A2(_AES_ENC_us10_n873 ), .A3(_AES_ENC_us10_n872 ), .A4(_AES_ENC_us10_n871 ), .ZN(_AES_ENC_us10_n875 ) );
NAND2_X2 _AES_ENC_us10_U192  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n875 ), .ZN(_AES_ENC_us10_n904 ) );
NAND2_X2 _AES_ENC_us10_U191  ( .A1(_AES_ENC_us10_n583 ), .A2(_AES_ENC_us10_n1050 ), .ZN(_AES_ENC_us10_n889 ) );
NAND2_X2 _AES_ENC_us10_U190  ( .A1(_AES_ENC_us10_n1093 ), .A2(_AES_ENC_us10_n587 ), .ZN(_AES_ENC_us10_n876 ) );
NAND2_X2 _AES_ENC_us10_U189  ( .A1(_AES_ENC_us10_n604 ), .A2(_AES_ENC_us10_n876 ), .ZN(_AES_ENC_us10_n877 ) );
NAND2_X2 _AES_ENC_us10_U188  ( .A1(_AES_ENC_us10_n877 ), .A2(_AES_ENC_us10_n623 ), .ZN(_AES_ENC_us10_n888 ) );
NAND4_X2 _AES_ENC_us10_U179  ( .A1(_AES_ENC_us10_n889 ), .A2(_AES_ENC_us10_n888 ), .A3(_AES_ENC_us10_n887 ), .A4(_AES_ENC_us10_n886 ), .ZN(_AES_ENC_us10_n890 ) );
NAND2_X2 _AES_ENC_us10_U178  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n890 ), .ZN(_AES_ENC_us10_n903 ) );
OR2_X2 _AES_ENC_us10_U177  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n1059 ), .ZN(_AES_ENC_us10_n900 ) );
NAND2_X2 _AES_ENC_us10_U176  ( .A1(_AES_ENC_us10_n1073 ), .A2(_AES_ENC_us10_n1047 ), .ZN(_AES_ENC_us10_n899 ) );
NAND2_X2 _AES_ENC_us10_U175  ( .A1(_AES_ENC_us10_n1094 ), .A2(_AES_ENC_us10_n595 ), .ZN(_AES_ENC_us10_n898 ) );
NAND4_X2 _AES_ENC_us10_U167  ( .A1(_AES_ENC_us10_n900 ), .A2(_AES_ENC_us10_n899 ), .A3(_AES_ENC_us10_n898 ), .A4(_AES_ENC_us10_n897 ), .ZN(_AES_ENC_us10_n901 ) );
NAND2_X2 _AES_ENC_us10_U166  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n901 ), .ZN(_AES_ENC_us10_n902 ) );
NAND4_X2 _AES_ENC_us10_U165  ( .A1(_AES_ENC_us10_n905 ), .A2(_AES_ENC_us10_n904 ), .A3(_AES_ENC_us10_n903 ), .A4(_AES_ENC_us10_n902 ), .ZN(_AES_ENC_sa10_sub[4] ) );
NAND2_X2 _AES_ENC_us10_U164  ( .A1(_AES_ENC_us10_n1094 ), .A2(_AES_ENC_us10_n599 ), .ZN(_AES_ENC_us10_n922 ) );
NAND2_X2 _AES_ENC_us10_U163  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n989 ), .ZN(_AES_ENC_us10_n921 ) );
NAND4_X2 _AES_ENC_us10_U151  ( .A1(_AES_ENC_us10_n922 ), .A2(_AES_ENC_us10_n921 ), .A3(_AES_ENC_us10_n920 ), .A4(_AES_ENC_us10_n919 ), .ZN(_AES_ENC_us10_n923 ) );
NAND2_X2 _AES_ENC_us10_U150  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n923 ), .ZN(_AES_ENC_us10_n972 ) );
NAND2_X2 _AES_ENC_us10_U149  ( .A1(_AES_ENC_us10_n582 ), .A2(_AES_ENC_us10_n619 ), .ZN(_AES_ENC_us10_n924 ) );
NAND2_X2 _AES_ENC_us10_U148  ( .A1(_AES_ENC_us10_n1073 ), .A2(_AES_ENC_us10_n924 ), .ZN(_AES_ENC_us10_n939 ) );
NAND2_X2 _AES_ENC_us10_U147  ( .A1(_AES_ENC_us10_n926 ), .A2(_AES_ENC_us10_n925 ), .ZN(_AES_ENC_us10_n927 ) );
NAND2_X2 _AES_ENC_us10_U146  ( .A1(_AES_ENC_us10_n606 ), .A2(_AES_ENC_us10_n927 ), .ZN(_AES_ENC_us10_n928 ) );
NAND2_X2 _AES_ENC_us10_U145  ( .A1(_AES_ENC_us10_n928 ), .A2(_AES_ENC_us10_n1080 ), .ZN(_AES_ENC_us10_n938 ) );
OR2_X2 _AES_ENC_us10_U144  ( .A1(_AES_ENC_us10_n1117 ), .A2(_AES_ENC_us10_n615 ), .ZN(_AES_ENC_us10_n937 ) );
NAND4_X2 _AES_ENC_us10_U139  ( .A1(_AES_ENC_us10_n939 ), .A2(_AES_ENC_us10_n938 ), .A3(_AES_ENC_us10_n937 ), .A4(_AES_ENC_us10_n936 ), .ZN(_AES_ENC_us10_n940 ) );
NAND2_X2 _AES_ENC_us10_U138  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n940 ), .ZN(_AES_ENC_us10_n971 ) );
OR2_X2 _AES_ENC_us10_U137  ( .A1(_AES_ENC_us10_n605 ), .A2(_AES_ENC_us10_n941 ), .ZN(_AES_ENC_us10_n954 ) );
NAND2_X2 _AES_ENC_us10_U136  ( .A1(_AES_ENC_us10_n1096 ), .A2(_AES_ENC_us10_n577 ), .ZN(_AES_ENC_us10_n942 ) );
NAND2_X2 _AES_ENC_us10_U135  ( .A1(_AES_ENC_us10_n1048 ), .A2(_AES_ENC_us10_n942 ), .ZN(_AES_ENC_us10_n943 ) );
NAND2_X2 _AES_ENC_us10_U134  ( .A1(_AES_ENC_us10_n612 ), .A2(_AES_ENC_us10_n943 ), .ZN(_AES_ENC_us10_n944 ) );
NAND2_X2 _AES_ENC_us10_U133  ( .A1(_AES_ENC_us10_n944 ), .A2(_AES_ENC_us10_n580 ), .ZN(_AES_ENC_us10_n953 ) );
NAND4_X2 _AES_ENC_us10_U125  ( .A1(_AES_ENC_us10_n954 ), .A2(_AES_ENC_us10_n953 ), .A3(_AES_ENC_us10_n952 ), .A4(_AES_ENC_us10_n951 ), .ZN(_AES_ENC_us10_n955 ) );
NAND2_X2 _AES_ENC_us10_U124  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n955 ), .ZN(_AES_ENC_us10_n970 ) );
NAND2_X2 _AES_ENC_us10_U123  ( .A1(_AES_ENC_us10_n1094 ), .A2(_AES_ENC_us10_n1071 ), .ZN(_AES_ENC_us10_n967 ) );
NAND2_X2 _AES_ENC_us10_U122  ( .A1(_AES_ENC_us10_n956 ), .A2(_AES_ENC_us10_n1030 ), .ZN(_AES_ENC_us10_n966 ) );
NAND4_X2 _AES_ENC_us10_U114  ( .A1(_AES_ENC_us10_n967 ), .A2(_AES_ENC_us10_n966 ), .A3(_AES_ENC_us10_n965 ), .A4(_AES_ENC_us10_n964 ), .ZN(_AES_ENC_us10_n968 ) );
NAND2_X2 _AES_ENC_us10_U113  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n968 ), .ZN(_AES_ENC_us10_n969 ) );
NAND4_X2 _AES_ENC_us10_U112  ( .A1(_AES_ENC_us10_n972 ), .A2(_AES_ENC_us10_n971 ), .A3(_AES_ENC_us10_n970 ), .A4(_AES_ENC_us10_n969 ), .ZN(_AES_ENC_sa10_sub[5] ) );
NAND2_X2 _AES_ENC_us10_U111  ( .A1(_AES_ENC_us10_n570 ), .A2(_AES_ENC_us10_n1097 ), .ZN(_AES_ENC_us10_n973 ) );
NAND2_X2 _AES_ENC_us10_U110  ( .A1(_AES_ENC_us10_n1073 ), .A2(_AES_ENC_us10_n973 ), .ZN(_AES_ENC_us10_n987 ) );
NAND2_X2 _AES_ENC_us10_U109  ( .A1(_AES_ENC_us10_n974 ), .A2(_AES_ENC_us10_n1077 ), .ZN(_AES_ENC_us10_n975 ) );
NAND2_X2 _AES_ENC_us10_U108  ( .A1(_AES_ENC_us10_n613 ), .A2(_AES_ENC_us10_n975 ), .ZN(_AES_ENC_us10_n976 ) );
NAND2_X2 _AES_ENC_us10_U107  ( .A1(_AES_ENC_us10_n977 ), .A2(_AES_ENC_us10_n976 ), .ZN(_AES_ENC_us10_n986 ) );
NAND4_X2 _AES_ENC_us10_U99  ( .A1(_AES_ENC_us10_n987 ), .A2(_AES_ENC_us10_n986 ), .A3(_AES_ENC_us10_n985 ), .A4(_AES_ENC_us10_n984 ), .ZN(_AES_ENC_us10_n988 ) );
NAND2_X2 _AES_ENC_us10_U98  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n988 ), .ZN(_AES_ENC_us10_n1044 ) );
NAND2_X2 _AES_ENC_us10_U97  ( .A1(_AES_ENC_us10_n1073 ), .A2(_AES_ENC_us10_n989 ), .ZN(_AES_ENC_us10_n1004 ) );
NAND2_X2 _AES_ENC_us10_U96  ( .A1(_AES_ENC_us10_n1092 ), .A2(_AES_ENC_us10_n619 ), .ZN(_AES_ENC_us10_n1003 ) );
NAND4_X2 _AES_ENC_us10_U85  ( .A1(_AES_ENC_us10_n1004 ), .A2(_AES_ENC_us10_n1003 ), .A3(_AES_ENC_us10_n1002 ), .A4(_AES_ENC_us10_n1001 ), .ZN(_AES_ENC_us10_n1005 ) );
NAND2_X2 _AES_ENC_us10_U84  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n1005 ), .ZN(_AES_ENC_us10_n1043 ) );
NAND2_X2 _AES_ENC_us10_U83  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n596 ), .ZN(_AES_ENC_us10_n1020 ) );
NAND2_X2 _AES_ENC_us10_U82  ( .A1(_AES_ENC_us10_n1050 ), .A2(_AES_ENC_us10_n624 ), .ZN(_AES_ENC_us10_n1019 ) );
NAND2_X2 _AES_ENC_us10_U77  ( .A1(_AES_ENC_us10_n1059 ), .A2(_AES_ENC_us10_n1114 ), .ZN(_AES_ENC_us10_n1012 ) );
NAND2_X2 _AES_ENC_us10_U76  ( .A1(_AES_ENC_us10_n1010 ), .A2(_AES_ENC_us10_n592 ), .ZN(_AES_ENC_us10_n1011 ) );
NAND2_X2 _AES_ENC_us10_U75  ( .A1(_AES_ENC_us10_n1012 ), .A2(_AES_ENC_us10_n1011 ), .ZN(_AES_ENC_us10_n1016 ) );
NAND4_X2 _AES_ENC_us10_U70  ( .A1(_AES_ENC_us10_n1020 ), .A2(_AES_ENC_us10_n1019 ), .A3(_AES_ENC_us10_n1018 ), .A4(_AES_ENC_us10_n1017 ), .ZN(_AES_ENC_us10_n1021 ) );
NAND2_X2 _AES_ENC_us10_U69  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n1021 ), .ZN(_AES_ENC_us10_n1042 ) );
NAND2_X2 _AES_ENC_us10_U68  ( .A1(_AES_ENC_us10_n1022 ), .A2(_AES_ENC_us10_n1093 ), .ZN(_AES_ENC_us10_n1039 ) );
NAND2_X2 _AES_ENC_us10_U67  ( .A1(_AES_ENC_us10_n1050 ), .A2(_AES_ENC_us10_n1023 ), .ZN(_AES_ENC_us10_n1038 ) );
NAND2_X2 _AES_ENC_us10_U66  ( .A1(_AES_ENC_us10_n1024 ), .A2(_AES_ENC_us10_n1071 ), .ZN(_AES_ENC_us10_n1037 ) );
AND2_X2 _AES_ENC_us10_U60  ( .A1(_AES_ENC_us10_n1030 ), .A2(_AES_ENC_us10_n602 ), .ZN(_AES_ENC_us10_n1078 ) );
NAND4_X2 _AES_ENC_us10_U56  ( .A1(_AES_ENC_us10_n1039 ), .A2(_AES_ENC_us10_n1038 ), .A3(_AES_ENC_us10_n1037 ), .A4(_AES_ENC_us10_n1036 ), .ZN(_AES_ENC_us10_n1040 ) );
NAND2_X2 _AES_ENC_us10_U55  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n1040 ), .ZN(_AES_ENC_us10_n1041 ) );
NAND4_X2 _AES_ENC_us10_U54  ( .A1(_AES_ENC_us10_n1044 ), .A2(_AES_ENC_us10_n1043 ), .A3(_AES_ENC_us10_n1042 ), .A4(_AES_ENC_us10_n1041 ), .ZN(_AES_ENC_sa10_sub[6] ) );
NAND2_X2 _AES_ENC_us10_U53  ( .A1(_AES_ENC_us10_n1072 ), .A2(_AES_ENC_us10_n1045 ), .ZN(_AES_ENC_us10_n1068 ) );
NAND2_X2 _AES_ENC_us10_U52  ( .A1(_AES_ENC_us10_n1046 ), .A2(_AES_ENC_us10_n582 ), .ZN(_AES_ENC_us10_n1067 ) );
NAND2_X2 _AES_ENC_us10_U51  ( .A1(_AES_ENC_us10_n1094 ), .A2(_AES_ENC_us10_n1047 ), .ZN(_AES_ENC_us10_n1066 ) );
NAND4_X2 _AES_ENC_us10_U40  ( .A1(_AES_ENC_us10_n1068 ), .A2(_AES_ENC_us10_n1067 ), .A3(_AES_ENC_us10_n1066 ), .A4(_AES_ENC_us10_n1065 ), .ZN(_AES_ENC_us10_n1069 ) );
NAND2_X2 _AES_ENC_us10_U39  ( .A1(_AES_ENC_us10_n1070 ), .A2(_AES_ENC_us10_n1069 ), .ZN(_AES_ENC_us10_n1135 ) );
NAND2_X2 _AES_ENC_us10_U38  ( .A1(_AES_ENC_us10_n1072 ), .A2(_AES_ENC_us10_n1071 ), .ZN(_AES_ENC_us10_n1088 ) );
NAND2_X2 _AES_ENC_us10_U37  ( .A1(_AES_ENC_us10_n1073 ), .A2(_AES_ENC_us10_n595 ), .ZN(_AES_ENC_us10_n1087 ) );
NAND4_X2 _AES_ENC_us10_U28  ( .A1(_AES_ENC_us10_n1088 ), .A2(_AES_ENC_us10_n1087 ), .A3(_AES_ENC_us10_n1086 ), .A4(_AES_ENC_us10_n1085 ), .ZN(_AES_ENC_us10_n1089 ) );
NAND2_X2 _AES_ENC_us10_U27  ( .A1(_AES_ENC_us10_n1090 ), .A2(_AES_ENC_us10_n1089 ), .ZN(_AES_ENC_us10_n1134 ) );
NAND2_X2 _AES_ENC_us10_U26  ( .A1(_AES_ENC_us10_n1091 ), .A2(_AES_ENC_us10_n1093 ), .ZN(_AES_ENC_us10_n1111 ) );
NAND2_X2 _AES_ENC_us10_U25  ( .A1(_AES_ENC_us10_n1092 ), .A2(_AES_ENC_us10_n1120 ), .ZN(_AES_ENC_us10_n1110 ) );
AND2_X2 _AES_ENC_us10_U22  ( .A1(_AES_ENC_us10_n1097 ), .A2(_AES_ENC_us10_n1096 ), .ZN(_AES_ENC_us10_n1098 ) );
NAND4_X2 _AES_ENC_us10_U14  ( .A1(_AES_ENC_us10_n1111 ), .A2(_AES_ENC_us10_n1110 ), .A3(_AES_ENC_us10_n1109 ), .A4(_AES_ENC_us10_n1108 ), .ZN(_AES_ENC_us10_n1112 ) );
NAND2_X2 _AES_ENC_us10_U13  ( .A1(_AES_ENC_us10_n1113 ), .A2(_AES_ENC_us10_n1112 ), .ZN(_AES_ENC_us10_n1133 ) );
NAND2_X2 _AES_ENC_us10_U12  ( .A1(_AES_ENC_us10_n1115 ), .A2(_AES_ENC_us10_n1114 ), .ZN(_AES_ENC_us10_n1129 ) );
OR2_X2 _AES_ENC_us10_U11  ( .A1(_AES_ENC_us10_n608 ), .A2(_AES_ENC_us10_n1116 ), .ZN(_AES_ENC_us10_n1128 ) );
NAND4_X2 _AES_ENC_us10_U3  ( .A1(_AES_ENC_us10_n1129 ), .A2(_AES_ENC_us10_n1128 ), .A3(_AES_ENC_us10_n1127 ), .A4(_AES_ENC_us10_n1126 ), .ZN(_AES_ENC_us10_n1130 ) );
NAND2_X2 _AES_ENC_us10_U2  ( .A1(_AES_ENC_us10_n1131 ), .A2(_AES_ENC_us10_n1130 ), .ZN(_AES_ENC_us10_n1132 ) );
NAND4_X2 _AES_ENC_us10_U1  ( .A1(_AES_ENC_us10_n1135 ), .A2(_AES_ENC_us10_n1134 ), .A3(_AES_ENC_us10_n1133 ), .A4(_AES_ENC_us10_n1132 ), .ZN(_AES_ENC_sa10_sub[7] ) );
INV_X4 _AES_ENC_us11_U575  ( .A(_AES_ENC_sa11[7]), .ZN(_AES_ENC_us11_n627 ));
INV_X4 _AES_ENC_us11_U574  ( .A(_AES_ENC_us11_n1114 ), .ZN(_AES_ENC_us11_n625 ) );
INV_X4 _AES_ENC_us11_U573  ( .A(_AES_ENC_sa11[4]), .ZN(_AES_ENC_us11_n624 ));
INV_X4 _AES_ENC_us11_U572  ( .A(_AES_ENC_us11_n1025 ), .ZN(_AES_ENC_us11_n622 ) );
INV_X4 _AES_ENC_us11_U571  ( .A(_AES_ENC_us11_n1120 ), .ZN(_AES_ENC_us11_n620 ) );
INV_X4 _AES_ENC_us11_U570  ( .A(_AES_ENC_us11_n1121 ), .ZN(_AES_ENC_us11_n619 ) );
INV_X4 _AES_ENC_us11_U569  ( .A(_AES_ENC_us11_n1048 ), .ZN(_AES_ENC_us11_n618 ) );
INV_X4 _AES_ENC_us11_U568  ( .A(_AES_ENC_us11_n974 ), .ZN(_AES_ENC_us11_n616 ) );
INV_X4 _AES_ENC_us11_U567  ( .A(_AES_ENC_us11_n794 ), .ZN(_AES_ENC_us11_n614 ) );
INV_X4 _AES_ENC_us11_U566  ( .A(_AES_ENC_sa11[2]), .ZN(_AES_ENC_us11_n611 ));
INV_X4 _AES_ENC_us11_U565  ( .A(_AES_ENC_us11_n800 ), .ZN(_AES_ENC_us11_n610 ) );
INV_X4 _AES_ENC_us11_U564  ( .A(_AES_ENC_us11_n925 ), .ZN(_AES_ENC_us11_n609 ) );
INV_X4 _AES_ENC_us11_U563  ( .A(_AES_ENC_us11_n779 ), .ZN(_AES_ENC_us11_n607 ) );
INV_X4 _AES_ENC_us11_U562  ( .A(_AES_ENC_us11_n1022 ), .ZN(_AES_ENC_us11_n603 ) );
INV_X4 _AES_ENC_us11_U561  ( .A(_AES_ENC_us11_n1102 ), .ZN(_AES_ENC_us11_n602 ) );
INV_X4 _AES_ENC_us11_U560  ( .A(_AES_ENC_us11_n929 ), .ZN(_AES_ENC_us11_n601 ) );
INV_X4 _AES_ENC_us11_U559  ( .A(_AES_ENC_us11_n1056 ), .ZN(_AES_ENC_us11_n600 ) );
INV_X4 _AES_ENC_us11_U558  ( .A(_AES_ENC_us11_n1054 ), .ZN(_AES_ENC_us11_n599 ) );
INV_X4 _AES_ENC_us11_U557  ( .A(_AES_ENC_us11_n881 ), .ZN(_AES_ENC_us11_n598 ) );
INV_X4 _AES_ENC_us11_U556  ( .A(_AES_ENC_us11_n926 ), .ZN(_AES_ENC_us11_n597 ) );
INV_X4 _AES_ENC_us11_U555  ( .A(_AES_ENC_us11_n977 ), .ZN(_AES_ENC_us11_n595 ) );
INV_X4 _AES_ENC_us11_U554  ( .A(_AES_ENC_us11_n1031 ), .ZN(_AES_ENC_us11_n594 ) );
INV_X4 _AES_ENC_us11_U553  ( .A(_AES_ENC_us11_n1103 ), .ZN(_AES_ENC_us11_n593 ) );
INV_X4 _AES_ENC_us11_U552  ( .A(_AES_ENC_us11_n1009 ), .ZN(_AES_ENC_us11_n592 ) );
INV_X4 _AES_ENC_us11_U551  ( .A(_AES_ENC_us11_n990 ), .ZN(_AES_ENC_us11_n591 ) );
INV_X4 _AES_ENC_us11_U550  ( .A(_AES_ENC_us11_n1058 ), .ZN(_AES_ENC_us11_n590 ) );
INV_X4 _AES_ENC_us11_U549  ( .A(_AES_ENC_us11_n1074 ), .ZN(_AES_ENC_us11_n589 ) );
INV_X4 _AES_ENC_us11_U548  ( .A(_AES_ENC_us11_n1053 ), .ZN(_AES_ENC_us11_n588 ) );
INV_X4 _AES_ENC_us11_U547  ( .A(_AES_ENC_us11_n826 ), .ZN(_AES_ENC_us11_n587 ) );
INV_X4 _AES_ENC_us11_U546  ( .A(_AES_ENC_us11_n992 ), .ZN(_AES_ENC_us11_n586 ) );
INV_X4 _AES_ENC_us11_U545  ( .A(_AES_ENC_us11_n821 ), .ZN(_AES_ENC_us11_n585 ) );
INV_X4 _AES_ENC_us11_U544  ( .A(_AES_ENC_us11_n910 ), .ZN(_AES_ENC_us11_n584 ) );
INV_X4 _AES_ENC_us11_U543  ( .A(_AES_ENC_us11_n906 ), .ZN(_AES_ENC_us11_n583 ) );
INV_X4 _AES_ENC_us11_U542  ( .A(_AES_ENC_us11_n880 ), .ZN(_AES_ENC_us11_n581 ) );
INV_X4 _AES_ENC_us11_U541  ( .A(_AES_ENC_us11_n1013 ), .ZN(_AES_ENC_us11_n580 ) );
INV_X4 _AES_ENC_us11_U540  ( .A(_AES_ENC_us11_n1092 ), .ZN(_AES_ENC_us11_n579 ) );
INV_X4 _AES_ENC_us11_U539  ( .A(_AES_ENC_us11_n824 ), .ZN(_AES_ENC_us11_n578 ) );
INV_X4 _AES_ENC_us11_U538  ( .A(_AES_ENC_us11_n1091 ), .ZN(_AES_ENC_us11_n577 ) );
INV_X4 _AES_ENC_us11_U537  ( .A(_AES_ENC_us11_n1080 ), .ZN(_AES_ENC_us11_n576 ) );
INV_X4 _AES_ENC_us11_U536  ( .A(_AES_ENC_us11_n959 ), .ZN(_AES_ENC_us11_n575 ) );
INV_X4 _AES_ENC_us11_U535  ( .A(_AES_ENC_sa11[0]), .ZN(_AES_ENC_us11_n574 ));
NOR2_X2 _AES_ENC_us11_U534  ( .A1(_AES_ENC_sa11[0]), .A2(_AES_ENC_sa11[6]),.ZN(_AES_ENC_us11_n1090 ) );
NOR2_X2 _AES_ENC_us11_U533  ( .A1(_AES_ENC_us11_n574 ), .A2(_AES_ENC_sa11[6]), .ZN(_AES_ENC_us11_n1070 ) );
NOR2_X2 _AES_ENC_us11_U532  ( .A1(_AES_ENC_sa11[4]), .A2(_AES_ENC_sa11[3]),.ZN(_AES_ENC_us11_n1025 ) );
INV_X4 _AES_ENC_us11_U531  ( .A(_AES_ENC_us11_n569 ), .ZN(_AES_ENC_us11_n572 ) );
NOR2_X2 _AES_ENC_us11_U530  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n765 ) );
NOR2_X2 _AES_ENC_us11_U529  ( .A1(_AES_ENC_sa11[4]), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n764 ) );
NOR2_X2 _AES_ENC_us11_U528  ( .A1(_AES_ENC_us11_n765 ), .A2(_AES_ENC_us11_n764 ), .ZN(_AES_ENC_us11_n766 ) );
NOR2_X2 _AES_ENC_us11_U527  ( .A1(_AES_ENC_us11_n766 ), .A2(_AES_ENC_us11_n575 ), .ZN(_AES_ENC_us11_n767 ) );
NOR3_X2 _AES_ENC_us11_U526  ( .A1(_AES_ENC_us11_n627 ), .A2(_AES_ENC_sa11[5]), .A3(_AES_ENC_us11_n704 ), .ZN(_AES_ENC_us11_n706 ));
NOR2_X2 _AES_ENC_us11_U525  ( .A1(_AES_ENC_us11_n1117 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n707 ) );
NOR2_X2 _AES_ENC_us11_U524  ( .A1(_AES_ENC_sa11[4]), .A2(_AES_ENC_us11_n579 ), .ZN(_AES_ENC_us11_n705 ) );
NOR3_X2 _AES_ENC_us11_U523  ( .A1(_AES_ENC_us11_n707 ), .A2(_AES_ENC_us11_n706 ), .A3(_AES_ENC_us11_n705 ), .ZN(_AES_ENC_us11_n713 ) );
INV_X4 _AES_ENC_us11_U522  ( .A(_AES_ENC_sa11[3]), .ZN(_AES_ENC_us11_n621 ));
NAND3_X2 _AES_ENC_us11_U521  ( .A1(_AES_ENC_us11_n652 ), .A2(_AES_ENC_us11_n626 ), .A3(_AES_ENC_sa11[7]), .ZN(_AES_ENC_us11_n653 ));
NOR2_X2 _AES_ENC_us11_U520  ( .A1(_AES_ENC_us11_n611 ), .A2(_AES_ENC_sa11[5]), .ZN(_AES_ENC_us11_n925 ) );
NOR2_X2 _AES_ENC_us11_U519  ( .A1(_AES_ENC_sa11[5]), .A2(_AES_ENC_sa11[2]),.ZN(_AES_ENC_us11_n974 ) );
INV_X4 _AES_ENC_us11_U518  ( .A(_AES_ENC_sa11[5]), .ZN(_AES_ENC_us11_n626 ));
NOR2_X2 _AES_ENC_us11_U517  ( .A1(_AES_ENC_us11_n611 ), .A2(_AES_ENC_sa11[7]), .ZN(_AES_ENC_us11_n779 ) );
NAND3_X2 _AES_ENC_us11_U516  ( .A1(_AES_ENC_us11_n679 ), .A2(_AES_ENC_us11_n678 ), .A3(_AES_ENC_us11_n677 ), .ZN(_AES_ENC_sa11_sub[0] ) );
NOR2_X2 _AES_ENC_us11_U515  ( .A1(_AES_ENC_us11_n626 ), .A2(_AES_ENC_sa11[2]), .ZN(_AES_ENC_us11_n1048 ) );
NOR4_X2 _AES_ENC_us11_U512  ( .A1(_AES_ENC_us11_n633 ), .A2(_AES_ENC_us11_n632 ), .A3(_AES_ENC_us11_n631 ), .A4(_AES_ENC_us11_n630 ), .ZN(_AES_ENC_us11_n634 ) );
NOR2_X2 _AES_ENC_us11_U510  ( .A1(_AES_ENC_us11_n629 ), .A2(_AES_ENC_us11_n628 ), .ZN(_AES_ENC_us11_n635 ) );
NAND3_X2 _AES_ENC_us11_U509  ( .A1(_AES_ENC_sa11[2]), .A2(_AES_ENC_sa11[7]), .A3(_AES_ENC_us11_n1059 ), .ZN(_AES_ENC_us11_n636 ) );
NOR2_X2 _AES_ENC_us11_U508  ( .A1(_AES_ENC_sa11[7]), .A2(_AES_ENC_sa11[2]),.ZN(_AES_ENC_us11_n794 ) );
NOR2_X2 _AES_ENC_us11_U507  ( .A1(_AES_ENC_sa11[4]), .A2(_AES_ENC_sa11[1]),.ZN(_AES_ENC_us11_n1102 ) );
NOR2_X2 _AES_ENC_us11_U506  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_sa11[3]), .ZN(_AES_ENC_us11_n1053 ) );
NOR2_X2 _AES_ENC_us11_U505  ( .A1(_AES_ENC_us11_n607 ), .A2(_AES_ENC_sa11[5]), .ZN(_AES_ENC_us11_n1024 ) );
NOR2_X2 _AES_ENC_us11_U504  ( .A1(_AES_ENC_us11_n625 ), .A2(_AES_ENC_sa11[2]), .ZN(_AES_ENC_us11_n1093 ) );
NOR2_X2 _AES_ENC_us11_U503  ( .A1(_AES_ENC_us11_n614 ), .A2(_AES_ENC_sa11[5]), .ZN(_AES_ENC_us11_n1094 ) );
NOR2_X2 _AES_ENC_us11_U502  ( .A1(_AES_ENC_us11_n624 ), .A2(_AES_ENC_sa11[3]), .ZN(_AES_ENC_us11_n931 ) );
INV_X4 _AES_ENC_us11_U501  ( .A(_AES_ENC_us11_n570 ), .ZN(_AES_ENC_us11_n573 ) );
NOR2_X2 _AES_ENC_us11_U500  ( .A1(_AES_ENC_us11_n1053 ), .A2(_AES_ENC_us11_n1095 ), .ZN(_AES_ENC_us11_n639 ) );
NOR3_X2 _AES_ENC_us11_U499  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n573 ), .A3(_AES_ENC_us11_n1074 ), .ZN(_AES_ENC_us11_n641 ) );
NOR2_X2 _AES_ENC_us11_U498  ( .A1(_AES_ENC_us11_n639 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n640 ) );
NOR2_X2 _AES_ENC_us11_U497  ( .A1(_AES_ENC_us11_n641 ), .A2(_AES_ENC_us11_n640 ), .ZN(_AES_ENC_us11_n646 ) );
NOR3_X2 _AES_ENC_us11_U496  ( .A1(_AES_ENC_us11_n995 ), .A2(_AES_ENC_us11_n586 ), .A3(_AES_ENC_us11_n994 ), .ZN(_AES_ENC_us11_n1002 ) );
NOR2_X2 _AES_ENC_us11_U495  ( .A1(_AES_ENC_us11_n909 ), .A2(_AES_ENC_us11_n908 ), .ZN(_AES_ENC_us11_n920 ) );
NOR2_X2 _AES_ENC_us11_U494  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n823 ) );
NOR2_X2 _AES_ENC_us11_U492  ( .A1(_AES_ENC_us11_n624 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n822 ) );
NOR2_X2 _AES_ENC_us11_U491  ( .A1(_AES_ENC_us11_n823 ), .A2(_AES_ENC_us11_n822 ), .ZN(_AES_ENC_us11_n825 ) );
NOR2_X2 _AES_ENC_us11_U490  ( .A1(_AES_ENC_sa11[1]), .A2(_AES_ENC_us11_n623 ), .ZN(_AES_ENC_us11_n913 ) );
NOR2_X2 _AES_ENC_us11_U489  ( .A1(_AES_ENC_us11_n913 ), .A2(_AES_ENC_us11_n1091 ), .ZN(_AES_ENC_us11_n914 ) );
NOR2_X2 _AES_ENC_us11_U488  ( .A1(_AES_ENC_us11_n826 ), .A2(_AES_ENC_us11_n572 ), .ZN(_AES_ENC_us11_n827 ) );
NOR3_X2 _AES_ENC_us11_U487  ( .A1(_AES_ENC_us11_n769 ), .A2(_AES_ENC_us11_n768 ), .A3(_AES_ENC_us11_n767 ), .ZN(_AES_ENC_us11_n775 ) );
NOR2_X2 _AES_ENC_us11_U486  ( .A1(_AES_ENC_us11_n1056 ), .A2(_AES_ENC_us11_n1053 ), .ZN(_AES_ENC_us11_n749 ) );
NOR2_X2 _AES_ENC_us11_U483  ( .A1(_AES_ENC_us11_n749 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n752 ) );
INV_X4 _AES_ENC_us11_U482  ( .A(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n596 ));
NOR2_X2 _AES_ENC_us11_U480  ( .A1(_AES_ENC_us11_n1054 ), .A2(_AES_ENC_us11_n1053 ), .ZN(_AES_ENC_us11_n1055 ) );
OR2_X4 _AES_ENC_us11_U479  ( .A1(_AES_ENC_us11_n1094 ), .A2(_AES_ENC_us11_n1093 ), .ZN(_AES_ENC_us11_n571 ) );
AND2_X2 _AES_ENC_us11_U478  ( .A1(_AES_ENC_us11_n571 ), .A2(_AES_ENC_us11_n1095 ), .ZN(_AES_ENC_us11_n1101 ) );
NOR2_X2 _AES_ENC_us11_U477  ( .A1(_AES_ENC_us11_n1074 ), .A2(_AES_ENC_us11_n931 ), .ZN(_AES_ENC_us11_n796 ) );
NOR2_X2 _AES_ENC_us11_U474  ( .A1(_AES_ENC_us11_n796 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n797 ) );
NOR2_X2 _AES_ENC_us11_U473  ( .A1(_AES_ENC_us11_n932 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n933 ) );
NOR2_X2 _AES_ENC_us11_U472  ( .A1(_AES_ENC_us11_n929 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n935 ) );
NOR2_X2 _AES_ENC_us11_U471  ( .A1(_AES_ENC_us11_n931 ), .A2(_AES_ENC_us11_n930 ), .ZN(_AES_ENC_us11_n934 ) );
NOR3_X2 _AES_ENC_us11_U470  ( .A1(_AES_ENC_us11_n935 ), .A2(_AES_ENC_us11_n934 ), .A3(_AES_ENC_us11_n933 ), .ZN(_AES_ENC_us11_n936 ) );
NOR2_X2 _AES_ENC_us11_U469  ( .A1(_AES_ENC_us11_n624 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n1075 ) );
NOR2_X2 _AES_ENC_us11_U468  ( .A1(_AES_ENC_us11_n572 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n949 ) );
NOR2_X2 _AES_ENC_us11_U467  ( .A1(_AES_ENC_us11_n1049 ), .A2(_AES_ENC_us11_n618 ), .ZN(_AES_ENC_us11_n1051 ) );
NOR2_X2 _AES_ENC_us11_U466  ( .A1(_AES_ENC_us11_n1051 ), .A2(_AES_ENC_us11_n1050 ), .ZN(_AES_ENC_us11_n1052 ) );
NOR2_X2 _AES_ENC_us11_U465  ( .A1(_AES_ENC_us11_n1052 ), .A2(_AES_ENC_us11_n592 ), .ZN(_AES_ENC_us11_n1064 ) );
NOR2_X2 _AES_ENC_us11_U464  ( .A1(_AES_ENC_sa11[1]), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n631 ) );
NOR2_X2 _AES_ENC_us11_U463  ( .A1(_AES_ENC_us11_n1025 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n980 ) );
NOR2_X2 _AES_ENC_us11_U462  ( .A1(_AES_ENC_us11_n1073 ), .A2(_AES_ENC_us11_n1094 ), .ZN(_AES_ENC_us11_n795 ) );
NOR2_X2 _AES_ENC_us11_U461  ( .A1(_AES_ENC_us11_n795 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n799 ) );
NOR2_X2 _AES_ENC_us11_U460  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n981 ) );
NOR2_X2 _AES_ENC_us11_U459  ( .A1(_AES_ENC_us11_n1102 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n643 ) );
NOR2_X2 _AES_ENC_us11_U458  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n621 ), .ZN(_AES_ENC_us11_n642 ) );
NOR2_X2 _AES_ENC_us11_U455  ( .A1(_AES_ENC_us11_n911 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n644 ) );
NOR4_X2 _AES_ENC_us11_U448  ( .A1(_AES_ENC_us11_n644 ), .A2(_AES_ENC_us11_n643 ), .A3(_AES_ENC_us11_n804 ), .A4(_AES_ENC_us11_n642 ), .ZN(_AES_ENC_us11_n645 ) );
NOR2_X2 _AES_ENC_us11_U447  ( .A1(_AES_ENC_us11_n1102 ), .A2(_AES_ENC_us11_n910 ), .ZN(_AES_ENC_us11_n932 ) );
NOR2_X2 _AES_ENC_us11_U442  ( .A1(_AES_ENC_us11_n1102 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n755 ) );
NOR2_X2 _AES_ENC_us11_U441  ( .A1(_AES_ENC_us11_n931 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n743 ) );
NOR2_X2 _AES_ENC_us11_U438  ( .A1(_AES_ENC_us11_n1072 ), .A2(_AES_ENC_us11_n1094 ), .ZN(_AES_ENC_us11_n930 ) );
NOR2_X2 _AES_ENC_us11_U435  ( .A1(_AES_ENC_us11_n1074 ), .A2(_AES_ENC_us11_n1025 ), .ZN(_AES_ENC_us11_n891 ) );
NOR2_X2 _AES_ENC_us11_U434  ( .A1(_AES_ENC_us11_n891 ), .A2(_AES_ENC_us11_n609 ), .ZN(_AES_ENC_us11_n894 ) );
NOR3_X2 _AES_ENC_us11_U433  ( .A1(_AES_ENC_us11_n623 ), .A2(_AES_ENC_sa11[1]), .A3(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n683 ));
INV_X4 _AES_ENC_us11_U428  ( .A(_AES_ENC_us11_n931 ), .ZN(_AES_ENC_us11_n623 ) );
NOR2_X2 _AES_ENC_us11_U427  ( .A1(_AES_ENC_us11_n996 ), .A2(_AES_ENC_us11_n931 ), .ZN(_AES_ENC_us11_n704 ) );
NOR2_X2 _AES_ENC_us11_U421  ( .A1(_AES_ENC_us11_n931 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n685 ) );
NOR2_X2 _AES_ENC_us11_U420  ( .A1(_AES_ENC_us11_n1029 ), .A2(_AES_ENC_us11_n1025 ), .ZN(_AES_ENC_us11_n1079 ) );
NOR3_X2 _AES_ENC_us11_U419  ( .A1(_AES_ENC_us11_n589 ), .A2(_AES_ENC_us11_n1025 ), .A3(_AES_ENC_us11_n616 ), .ZN(_AES_ENC_us11_n945 ) );
NOR2_X2 _AES_ENC_us11_U418  ( .A1(_AES_ENC_us11_n626 ), .A2(_AES_ENC_us11_n611 ), .ZN(_AES_ENC_us11_n800 ) );
NOR3_X2 _AES_ENC_us11_U417  ( .A1(_AES_ENC_us11_n590 ), .A2(_AES_ENC_us11_n627 ), .A3(_AES_ENC_us11_n611 ), .ZN(_AES_ENC_us11_n798 ) );
NOR3_X2 _AES_ENC_us11_U416  ( .A1(_AES_ENC_us11_n610 ), .A2(_AES_ENC_us11_n572 ), .A3(_AES_ENC_us11_n575 ), .ZN(_AES_ENC_us11_n962 ) );
NOR3_X2 _AES_ENC_us11_U415  ( .A1(_AES_ENC_us11_n959 ), .A2(_AES_ENC_us11_n572 ), .A3(_AES_ENC_us11_n609 ), .ZN(_AES_ENC_us11_n768 ) );
NOR3_X2 _AES_ENC_us11_U414  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n572 ), .A3(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n694 ) );
NOR3_X2 _AES_ENC_us11_U413  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n572 ), .A3(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n895 ) );
NOR3_X2 _AES_ENC_us11_U410  ( .A1(_AES_ENC_us11_n1008 ), .A2(_AES_ENC_us11_n1007 ), .A3(_AES_ENC_us11_n1006 ), .ZN(_AES_ENC_us11_n1018 ) );
NOR4_X2 _AES_ENC_us11_U409  ( .A1(_AES_ENC_us11_n806 ), .A2(_AES_ENC_us11_n805 ), .A3(_AES_ENC_us11_n804 ), .A4(_AES_ENC_us11_n803 ), .ZN(_AES_ENC_us11_n807 ) );
NOR3_X2 _AES_ENC_us11_U406  ( .A1(_AES_ENC_us11_n799 ), .A2(_AES_ENC_us11_n798 ), .A3(_AES_ENC_us11_n797 ), .ZN(_AES_ENC_us11_n808 ) );
NOR4_X2 _AES_ENC_us11_U405  ( .A1(_AES_ENC_us11_n843 ), .A2(_AES_ENC_us11_n842 ), .A3(_AES_ENC_us11_n841 ), .A4(_AES_ENC_us11_n840 ), .ZN(_AES_ENC_us11_n844 ) );
NOR2_X2 _AES_ENC_us11_U404  ( .A1(_AES_ENC_us11_n669 ), .A2(_AES_ENC_us11_n668 ), .ZN(_AES_ENC_us11_n673 ) );
NOR4_X2 _AES_ENC_us11_U403  ( .A1(_AES_ENC_us11_n946 ), .A2(_AES_ENC_us11_n1046 ), .A3(_AES_ENC_us11_n671 ), .A4(_AES_ENC_us11_n670 ), .ZN(_AES_ENC_us11_n672 ) );
NOR4_X2 _AES_ENC_us11_U401  ( .A1(_AES_ENC_us11_n711 ), .A2(_AES_ENC_us11_n710 ), .A3(_AES_ENC_us11_n709 ), .A4(_AES_ENC_us11_n708 ), .ZN(_AES_ENC_us11_n712 ) );
NOR4_X2 _AES_ENC_us11_U400  ( .A1(_AES_ENC_us11_n963 ), .A2(_AES_ENC_us11_n962 ), .A3(_AES_ENC_us11_n961 ), .A4(_AES_ENC_us11_n960 ), .ZN(_AES_ENC_us11_n964 ) );
NOR3_X2 _AES_ENC_us11_U399  ( .A1(_AES_ENC_us11_n1101 ), .A2(_AES_ENC_us11_n1100 ), .A3(_AES_ENC_us11_n1099 ), .ZN(_AES_ENC_us11_n1109 ) );
NOR3_X2 _AES_ENC_us11_U398  ( .A1(_AES_ENC_us11_n743 ), .A2(_AES_ENC_us11_n742 ), .A3(_AES_ENC_us11_n741 ), .ZN(_AES_ENC_us11_n744 ) );
NOR2_X2 _AES_ENC_us11_U397  ( .A1(_AES_ENC_us11_n697 ), .A2(_AES_ENC_us11_n658 ), .ZN(_AES_ENC_us11_n659 ) );
NOR2_X2 _AES_ENC_us11_U396  ( .A1(_AES_ENC_us11_n1078 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n1033 ) );
NOR2_X2 _AES_ENC_us11_U393  ( .A1(_AES_ENC_us11_n1031 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n1032 ) );
NOR3_X2 _AES_ENC_us11_U390  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n1025 ), .A3(_AES_ENC_us11_n1074 ), .ZN(_AES_ENC_us11_n1035 ) );
NOR4_X2 _AES_ENC_us11_U389  ( .A1(_AES_ENC_us11_n1035 ), .A2(_AES_ENC_us11_n1034 ), .A3(_AES_ENC_us11_n1033 ), .A4(_AES_ENC_us11_n1032 ), .ZN(_AES_ENC_us11_n1036 ) );
NOR2_X2 _AES_ENC_us11_U388  ( .A1(_AES_ENC_us11_n598 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n885 ) );
NOR2_X2 _AES_ENC_us11_U387  ( .A1(_AES_ENC_us11_n623 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n882 ) );
NOR2_X2 _AES_ENC_us11_U386  ( .A1(_AES_ENC_us11_n1053 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n884 ) );
NOR4_X2 _AES_ENC_us11_U385  ( .A1(_AES_ENC_us11_n885 ), .A2(_AES_ENC_us11_n884 ), .A3(_AES_ENC_us11_n883 ), .A4(_AES_ENC_us11_n882 ), .ZN(_AES_ENC_us11_n886 ) );
NOR2_X2 _AES_ENC_us11_U384  ( .A1(_AES_ENC_us11_n825 ), .A2(_AES_ENC_us11_n578 ), .ZN(_AES_ENC_us11_n830 ) );
NOR2_X2 _AES_ENC_us11_U383  ( .A1(_AES_ENC_us11_n827 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n829 ) );
NOR2_X2 _AES_ENC_us11_U382  ( .A1(_AES_ENC_us11_n572 ), .A2(_AES_ENC_us11_n579 ), .ZN(_AES_ENC_us11_n828 ) );
NOR4_X2 _AES_ENC_us11_U374  ( .A1(_AES_ENC_us11_n831 ), .A2(_AES_ENC_us11_n830 ), .A3(_AES_ENC_us11_n829 ), .A4(_AES_ENC_us11_n828 ), .ZN(_AES_ENC_us11_n832 ) );
NOR2_X2 _AES_ENC_us11_U373  ( .A1(_AES_ENC_us11_n606 ), .A2(_AES_ENC_us11_n582 ), .ZN(_AES_ENC_us11_n1104 ) );
NOR2_X2 _AES_ENC_us11_U372  ( .A1(_AES_ENC_us11_n1102 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n1106 ) );
NOR2_X2 _AES_ENC_us11_U370  ( .A1(_AES_ENC_us11_n1103 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n1105 ) );
NOR4_X2 _AES_ENC_us11_U369  ( .A1(_AES_ENC_us11_n1107 ), .A2(_AES_ENC_us11_n1106 ), .A3(_AES_ENC_us11_n1105 ), .A4(_AES_ENC_us11_n1104 ), .ZN(_AES_ENC_us11_n1108 ) );
NOR3_X2 _AES_ENC_us11_U368  ( .A1(_AES_ENC_us11_n959 ), .A2(_AES_ENC_us11_n621 ), .A3(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n963 ) );
NOR2_X2 _AES_ENC_us11_U367  ( .A1(_AES_ENC_us11_n626 ), .A2(_AES_ENC_us11_n627 ), .ZN(_AES_ENC_us11_n1114 ) );
INV_X4 _AES_ENC_us11_U366  ( .A(_AES_ENC_us11_n1024 ), .ZN(_AES_ENC_us11_n606 ) );
NOR3_X2 _AES_ENC_us11_U365  ( .A1(_AES_ENC_us11_n910 ), .A2(_AES_ENC_us11_n1059 ), .A3(_AES_ENC_us11_n611 ), .ZN(_AES_ENC_us11_n1115 ) );
INV_X4 _AES_ENC_us11_U364  ( .A(_AES_ENC_us11_n1094 ), .ZN(_AES_ENC_us11_n613 ) );
NOR2_X2 _AES_ENC_us11_U363  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n931 ), .ZN(_AES_ENC_us11_n1100 ) );
INV_X4 _AES_ENC_us11_U354  ( .A(_AES_ENC_us11_n1093 ), .ZN(_AES_ENC_us11_n617 ) );
NOR2_X2 _AES_ENC_us11_U353  ( .A1(_AES_ENC_us11_n569 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n929 ) );
NOR2_X2 _AES_ENC_us11_U352  ( .A1(_AES_ENC_us11_n620 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n926 ) );
NOR2_X2 _AES_ENC_us11_U351  ( .A1(_AES_ENC_us11_n572 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n1095 ) );
NOR2_X2 _AES_ENC_us11_U350  ( .A1(_AES_ENC_us11_n609 ), .A2(_AES_ENC_us11_n627 ), .ZN(_AES_ENC_us11_n1010 ) );
NOR2_X2 _AES_ENC_us11_U349  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n1103 ) );
NOR2_X2 _AES_ENC_us11_U348  ( .A1(_AES_ENC_us11_n622 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n1059 ) );
NOR2_X2 _AES_ENC_us11_U347  ( .A1(_AES_ENC_sa11[1]), .A2(_AES_ENC_us11_n1120 ), .ZN(_AES_ENC_us11_n1022 ) );
NOR2_X2 _AES_ENC_us11_U346  ( .A1(_AES_ENC_us11_n619 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n911 ) );
NOR2_X2 _AES_ENC_us11_U345  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_us11_n1025 ), .ZN(_AES_ENC_us11_n826 ) );
NOR2_X2 _AES_ENC_us11_U338  ( .A1(_AES_ENC_us11_n626 ), .A2(_AES_ENC_us11_n607 ), .ZN(_AES_ENC_us11_n1072 ) );
NOR2_X2 _AES_ENC_us11_U335  ( .A1(_AES_ENC_us11_n627 ), .A2(_AES_ENC_us11_n616 ), .ZN(_AES_ENC_us11_n956 ) );
NOR2_X2 _AES_ENC_us11_U329  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_us11_n624 ), .ZN(_AES_ENC_us11_n1121 ) );
NOR2_X2 _AES_ENC_us11_U328  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_us11_n624 ), .ZN(_AES_ENC_us11_n1058 ) );
NOR2_X2 _AES_ENC_us11_U327  ( .A1(_AES_ENC_us11_n625 ), .A2(_AES_ENC_us11_n611 ), .ZN(_AES_ENC_us11_n1073 ) );
NOR2_X2 _AES_ENC_us11_U325  ( .A1(_AES_ENC_sa11[1]), .A2(_AES_ENC_us11_n1025 ), .ZN(_AES_ENC_us11_n1054 ) );
NOR2_X2 _AES_ENC_us11_U324  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_us11_n931 ), .ZN(_AES_ENC_us11_n1029 ) );
NOR2_X2 _AES_ENC_us11_U319  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n1056 ) );
NOR2_X2 _AES_ENC_us11_U318  ( .A1(_AES_ENC_us11_n614 ), .A2(_AES_ENC_us11_n626 ), .ZN(_AES_ENC_us11_n1050 ) );
NOR2_X2 _AES_ENC_us11_U317  ( .A1(_AES_ENC_us11_n1121 ), .A2(_AES_ENC_us11_n1025 ), .ZN(_AES_ENC_us11_n1120 ) );
NOR2_X2 _AES_ENC_us11_U316  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_us11_n572 ), .ZN(_AES_ENC_us11_n1074 ) );
NOR2_X2 _AES_ENC_us11_U315  ( .A1(_AES_ENC_us11_n1058 ), .A2(_AES_ENC_us11_n1054 ), .ZN(_AES_ENC_us11_n878 ) );
NOR2_X2 _AES_ENC_us11_U314  ( .A1(_AES_ENC_us11_n878 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n879 ) );
NOR2_X2 _AES_ENC_us11_U312  ( .A1(_AES_ENC_us11_n880 ), .A2(_AES_ENC_us11_n879 ), .ZN(_AES_ENC_us11_n887 ) );
NOR2_X2 _AES_ENC_us11_U311  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n588 ), .ZN(_AES_ENC_us11_n957 ) );
NOR2_X2 _AES_ENC_us11_U310  ( .A1(_AES_ENC_us11_n958 ), .A2(_AES_ENC_us11_n957 ), .ZN(_AES_ENC_us11_n965 ) );
NOR3_X2 _AES_ENC_us11_U309  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n1091 ), .A3(_AES_ENC_us11_n1022 ), .ZN(_AES_ENC_us11_n720 ) );
NOR3_X2 _AES_ENC_us11_U303  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n1054 ), .A3(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n719 ) );
NOR2_X2 _AES_ENC_us11_U302  ( .A1(_AES_ENC_us11_n720 ), .A2(_AES_ENC_us11_n719 ), .ZN(_AES_ENC_us11_n726 ) );
NOR2_X2 _AES_ENC_us11_U300  ( .A1(_AES_ENC_us11_n614 ), .A2(_AES_ENC_us11_n591 ), .ZN(_AES_ENC_us11_n865 ) );
NOR2_X2 _AES_ENC_us11_U299  ( .A1(_AES_ENC_us11_n1059 ), .A2(_AES_ENC_us11_n1058 ), .ZN(_AES_ENC_us11_n1060 ) );
NOR2_X2 _AES_ENC_us11_U298  ( .A1(_AES_ENC_us11_n1095 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n668 ) );
NOR2_X2 _AES_ENC_us11_U297  ( .A1(_AES_ENC_us11_n911 ), .A2(_AES_ENC_us11_n910 ), .ZN(_AES_ENC_us11_n912 ) );
NOR2_X2 _AES_ENC_us11_U296  ( .A1(_AES_ENC_us11_n912 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n916 ) );
NOR2_X2 _AES_ENC_us11_U295  ( .A1(_AES_ENC_us11_n826 ), .A2(_AES_ENC_us11_n573 ), .ZN(_AES_ENC_us11_n750 ) );
NOR2_X2 _AES_ENC_us11_U294  ( .A1(_AES_ENC_us11_n750 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n751 ) );
NOR2_X2 _AES_ENC_us11_U293  ( .A1(_AES_ENC_us11_n907 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n908 ) );
NOR2_X2 _AES_ENC_us11_U292  ( .A1(_AES_ENC_us11_n990 ), .A2(_AES_ENC_us11_n926 ), .ZN(_AES_ENC_us11_n780 ) );
NOR2_X2 _AES_ENC_us11_U291  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n584 ), .ZN(_AES_ENC_us11_n838 ) );
NOR2_X2 _AES_ENC_us11_U290  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n602 ), .ZN(_AES_ENC_us11_n837 ) );
NOR2_X2 _AES_ENC_us11_U284  ( .A1(_AES_ENC_us11_n838 ), .A2(_AES_ENC_us11_n837 ), .ZN(_AES_ENC_us11_n845 ) );
NOR2_X2 _AES_ENC_us11_U283  ( .A1(_AES_ENC_us11_n1022 ), .A2(_AES_ENC_us11_n1058 ), .ZN(_AES_ENC_us11_n740 ) );
NOR2_X2 _AES_ENC_us11_U282  ( .A1(_AES_ENC_us11_n740 ), .A2(_AES_ENC_us11_n616 ), .ZN(_AES_ENC_us11_n742 ) );
NOR2_X2 _AES_ENC_us11_U281  ( .A1(_AES_ENC_us11_n1098 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n1099 ) );
NOR2_X2 _AES_ENC_us11_U280  ( .A1(_AES_ENC_us11_n1120 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n993 ) );
NOR2_X2 _AES_ENC_us11_U279  ( .A1(_AES_ENC_us11_n993 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n994 ) );
NOR2_X2 _AES_ENC_us11_U273  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n620 ), .ZN(_AES_ENC_us11_n1026 ) );
NOR2_X2 _AES_ENC_us11_U272  ( .A1(_AES_ENC_us11_n573 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n1027 ) );
NOR2_X2 _AES_ENC_us11_U271  ( .A1(_AES_ENC_us11_n1027 ), .A2(_AES_ENC_us11_n1026 ), .ZN(_AES_ENC_us11_n1028 ) );
NOR2_X2 _AES_ENC_us11_U270  ( .A1(_AES_ENC_us11_n1029 ), .A2(_AES_ENC_us11_n1028 ), .ZN(_AES_ENC_us11_n1034 ) );
NOR4_X2 _AES_ENC_us11_U269  ( .A1(_AES_ENC_us11_n757 ), .A2(_AES_ENC_us11_n756 ), .A3(_AES_ENC_us11_n755 ), .A4(_AES_ENC_us11_n754 ), .ZN(_AES_ENC_us11_n758 ) );
NOR2_X2 _AES_ENC_us11_U268  ( .A1(_AES_ENC_us11_n752 ), .A2(_AES_ENC_us11_n751 ), .ZN(_AES_ENC_us11_n759 ) );
NOR2_X2 _AES_ENC_us11_U267  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n1071 ), .ZN(_AES_ENC_us11_n669 ) );
NOR2_X2 _AES_ENC_us11_U263  ( .A1(_AES_ENC_us11_n1056 ), .A2(_AES_ENC_us11_n990 ), .ZN(_AES_ENC_us11_n991 ) );
NOR2_X2 _AES_ENC_us11_U262  ( .A1(_AES_ENC_us11_n991 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n995 ) );
NOR2_X2 _AES_ENC_us11_U258  ( .A1(_AES_ENC_us11_n607 ), .A2(_AES_ENC_us11_n590 ), .ZN(_AES_ENC_us11_n1008 ) );
NOR2_X2 _AES_ENC_us11_U255  ( .A1(_AES_ENC_us11_n839 ), .A2(_AES_ENC_us11_n582 ), .ZN(_AES_ENC_us11_n693 ) );
NOR2_X2 _AES_ENC_us11_U254  ( .A1(_AES_ENC_us11_n606 ), .A2(_AES_ENC_us11_n906 ), .ZN(_AES_ENC_us11_n741 ) );
NOR2_X2 _AES_ENC_us11_U253  ( .A1(_AES_ENC_us11_n1054 ), .A2(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n763 ) );
NOR2_X2 _AES_ENC_us11_U252  ( .A1(_AES_ENC_us11_n763 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n769 ) );
NOR2_X2 _AES_ENC_us11_U251  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n577 ), .ZN(_AES_ENC_us11_n1007 ) );
NOR2_X2 _AES_ENC_us11_U250  ( .A1(_AES_ENC_us11_n609 ), .A2(_AES_ENC_us11_n580 ), .ZN(_AES_ENC_us11_n1123 ) );
NOR2_X2 _AES_ENC_us11_U243  ( .A1(_AES_ENC_us11_n609 ), .A2(_AES_ENC_us11_n590 ), .ZN(_AES_ENC_us11_n710 ) );
INV_X4 _AES_ENC_us11_U242  ( .A(_AES_ENC_us11_n1029 ), .ZN(_AES_ENC_us11_n582 ) );
NOR2_X2 _AES_ENC_us11_U241  ( .A1(_AES_ENC_us11_n616 ), .A2(_AES_ENC_us11_n597 ), .ZN(_AES_ENC_us11_n883 ) );
NOR2_X2 _AES_ENC_us11_U240  ( .A1(_AES_ENC_us11_n593 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n1125 ) );
NOR2_X2 _AES_ENC_us11_U239  ( .A1(_AES_ENC_us11_n990 ), .A2(_AES_ENC_us11_n929 ), .ZN(_AES_ENC_us11_n892 ) );
NOR2_X2 _AES_ENC_us11_U238  ( .A1(_AES_ENC_us11_n892 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n893 ) );
NOR2_X2 _AES_ENC_us11_U237  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n602 ), .ZN(_AES_ENC_us11_n950 ) );
NOR2_X2 _AES_ENC_us11_U236  ( .A1(_AES_ENC_us11_n1079 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n1082 ) );
NOR2_X2 _AES_ENC_us11_U235  ( .A1(_AES_ENC_us11_n910 ), .A2(_AES_ENC_us11_n1056 ), .ZN(_AES_ENC_us11_n941 ) );
NOR2_X2 _AES_ENC_us11_U234  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n1077 ), .ZN(_AES_ENC_us11_n841 ) );
NOR2_X2 _AES_ENC_us11_U229  ( .A1(_AES_ENC_us11_n623 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n630 ) );
NOR2_X2 _AES_ENC_us11_U228  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n602 ), .ZN(_AES_ENC_us11_n806 ) );
NOR2_X2 _AES_ENC_us11_U227  ( .A1(_AES_ENC_us11_n623 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n948 ) );
NOR2_X2 _AES_ENC_us11_U226  ( .A1(_AES_ENC_us11_n606 ), .A2(_AES_ENC_us11_n589 ), .ZN(_AES_ENC_us11_n997 ) );
NOR2_X2 _AES_ENC_us11_U225  ( .A1(_AES_ENC_us11_n1121 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n1122 ) );
NOR2_X2 _AES_ENC_us11_U223  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n1023 ), .ZN(_AES_ENC_us11_n756 ) );
NOR2_X2 _AES_ENC_us11_U222  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n602 ), .ZN(_AES_ENC_us11_n870 ) );
NOR2_X2 _AES_ENC_us11_U221  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n569 ), .ZN(_AES_ENC_us11_n947 ) );
NOR2_X2 _AES_ENC_us11_U217  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n1077 ), .ZN(_AES_ENC_us11_n1084 ) );
NOR2_X2 _AES_ENC_us11_U213  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n855 ), .ZN(_AES_ENC_us11_n709 ) );
NOR2_X2 _AES_ENC_us11_U212  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n589 ), .ZN(_AES_ENC_us11_n868 ) );
NOR2_X2 _AES_ENC_us11_U211  ( .A1(_AES_ENC_us11_n1120 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n1124 ) );
NOR2_X2 _AES_ENC_us11_U210  ( .A1(_AES_ENC_us11_n1120 ), .A2(_AES_ENC_us11_n839 ), .ZN(_AES_ENC_us11_n842 ) );
NOR2_X2 _AES_ENC_us11_U209  ( .A1(_AES_ENC_us11_n1120 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n696 ) );
NOR2_X2 _AES_ENC_us11_U208  ( .A1(_AES_ENC_us11_n1074 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n1076 ) );
NOR2_X2 _AES_ENC_us11_U207  ( .A1(_AES_ENC_us11_n1074 ), .A2(_AES_ENC_us11_n620 ), .ZN(_AES_ENC_us11_n781 ) );
NOR3_X2 _AES_ENC_us11_U201  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n1056 ), .A3(_AES_ENC_us11_n990 ), .ZN(_AES_ENC_us11_n979 ) );
NOR3_X2 _AES_ENC_us11_U200  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n1058 ), .A3(_AES_ENC_us11_n1059 ), .ZN(_AES_ENC_us11_n854 ) );
NOR2_X2 _AES_ENC_us11_U199  ( .A1(_AES_ENC_us11_n996 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n869 ) );
NOR2_X2 _AES_ENC_us11_U198  ( .A1(_AES_ENC_us11_n1056 ), .A2(_AES_ENC_us11_n1074 ), .ZN(_AES_ENC_us11_n1057 ) );
NOR3_X2 _AES_ENC_us11_U197  ( .A1(_AES_ENC_us11_n607 ), .A2(_AES_ENC_us11_n1120 ), .A3(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n978 ) );
NOR2_X2 _AES_ENC_us11_U196  ( .A1(_AES_ENC_us11_n996 ), .A2(_AES_ENC_us11_n911 ), .ZN(_AES_ENC_us11_n1116 ) );
NOR2_X2 _AES_ENC_us11_U195  ( .A1(_AES_ENC_us11_n1074 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n754 ) );
NOR2_X2 _AES_ENC_us11_U194  ( .A1(_AES_ENC_us11_n926 ), .A2(_AES_ENC_us11_n1103 ), .ZN(_AES_ENC_us11_n977 ) );
NOR2_X2 _AES_ENC_us11_U187  ( .A1(_AES_ENC_us11_n839 ), .A2(_AES_ENC_us11_n824 ), .ZN(_AES_ENC_us11_n1092 ) );
NOR2_X2 _AES_ENC_us11_U186  ( .A1(_AES_ENC_us11_n573 ), .A2(_AES_ENC_us11_n1074 ), .ZN(_AES_ENC_us11_n684 ) );
NOR2_X2 _AES_ENC_us11_U185  ( .A1(_AES_ENC_us11_n826 ), .A2(_AES_ENC_us11_n1059 ), .ZN(_AES_ENC_us11_n907 ) );
NOR3_X2 _AES_ENC_us11_U184  ( .A1(_AES_ENC_us11_n625 ), .A2(_AES_ENC_us11_n1115 ), .A3(_AES_ENC_us11_n585 ), .ZN(_AES_ENC_us11_n831 ) );
NOR3_X2 _AES_ENC_us11_U183  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n1056 ), .A3(_AES_ENC_us11_n990 ), .ZN(_AES_ENC_us11_n896 ) );
NOR3_X2 _AES_ENC_us11_U182  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n573 ), .A3(_AES_ENC_us11_n1013 ), .ZN(_AES_ENC_us11_n670 ) );
NOR3_X2 _AES_ENC_us11_U181  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n1091 ), .A3(_AES_ENC_us11_n1022 ), .ZN(_AES_ENC_us11_n843 ) );
NOR2_X2 _AES_ENC_us11_U180  ( .A1(_AES_ENC_us11_n1029 ), .A2(_AES_ENC_us11_n1095 ), .ZN(_AES_ENC_us11_n735 ) );
NOR2_X2 _AES_ENC_us11_U174  ( .A1(_AES_ENC_us11_n1100 ), .A2(_AES_ENC_us11_n854 ), .ZN(_AES_ENC_us11_n860 ) );
NAND3_X2 _AES_ENC_us11_U173  ( .A1(_AES_ENC_us11_n569 ), .A2(_AES_ENC_us11_n582 ), .A3(_AES_ENC_us11_n681 ), .ZN(_AES_ENC_us11_n691 ) );
NOR2_X2 _AES_ENC_us11_U172  ( .A1(_AES_ENC_us11_n683 ), .A2(_AES_ENC_us11_n682 ), .ZN(_AES_ENC_us11_n690 ) );
NOR3_X2 _AES_ENC_us11_U171  ( .A1(_AES_ENC_us11_n695 ), .A2(_AES_ENC_us11_n694 ), .A3(_AES_ENC_us11_n693 ), .ZN(_AES_ENC_us11_n700 ) );
NOR4_X2 _AES_ENC_us11_U170  ( .A1(_AES_ENC_us11_n983 ), .A2(_AES_ENC_us11_n698 ), .A3(_AES_ENC_us11_n697 ), .A4(_AES_ENC_us11_n696 ), .ZN(_AES_ENC_us11_n699 ) );
NOR2_X2 _AES_ENC_us11_U169  ( .A1(_AES_ENC_us11_n946 ), .A2(_AES_ENC_us11_n945 ), .ZN(_AES_ENC_us11_n952 ) );
NOR4_X2 _AES_ENC_us11_U168  ( .A1(_AES_ENC_us11_n950 ), .A2(_AES_ENC_us11_n949 ), .A3(_AES_ENC_us11_n948 ), .A4(_AES_ENC_us11_n947 ), .ZN(_AES_ENC_us11_n951 ) );
NOR4_X2 _AES_ENC_us11_U162  ( .A1(_AES_ENC_us11_n896 ), .A2(_AES_ENC_us11_n895 ), .A3(_AES_ENC_us11_n894 ), .A4(_AES_ENC_us11_n893 ), .ZN(_AES_ENC_us11_n897 ) );
NOR2_X2 _AES_ENC_us11_U161  ( .A1(_AES_ENC_us11_n866 ), .A2(_AES_ENC_us11_n865 ), .ZN(_AES_ENC_us11_n872 ) );
NOR4_X2 _AES_ENC_us11_U160  ( .A1(_AES_ENC_us11_n870 ), .A2(_AES_ENC_us11_n869 ), .A3(_AES_ENC_us11_n868 ), .A4(_AES_ENC_us11_n867 ), .ZN(_AES_ENC_us11_n871 ) );
NOR4_X2 _AES_ENC_us11_U159  ( .A1(_AES_ENC_us11_n983 ), .A2(_AES_ENC_us11_n982 ), .A3(_AES_ENC_us11_n981 ), .A4(_AES_ENC_us11_n980 ), .ZN(_AES_ENC_us11_n984 ) );
NOR2_X2 _AES_ENC_us11_U158  ( .A1(_AES_ENC_us11_n979 ), .A2(_AES_ENC_us11_n978 ), .ZN(_AES_ENC_us11_n985 ) );
NOR4_X2 _AES_ENC_us11_U157  ( .A1(_AES_ENC_us11_n1125 ), .A2(_AES_ENC_us11_n1124 ), .A3(_AES_ENC_us11_n1123 ), .A4(_AES_ENC_us11_n1122 ), .ZN(_AES_ENC_us11_n1126 ) );
NOR4_X2 _AES_ENC_us11_U156  ( .A1(_AES_ENC_us11_n1084 ), .A2(_AES_ENC_us11_n1083 ), .A3(_AES_ENC_us11_n1082 ), .A4(_AES_ENC_us11_n1081 ), .ZN(_AES_ENC_us11_n1085 ) );
NOR2_X2 _AES_ENC_us11_U155  ( .A1(_AES_ENC_us11_n1076 ), .A2(_AES_ENC_us11_n1075 ), .ZN(_AES_ENC_us11_n1086 ) );
NOR3_X2 _AES_ENC_us11_U154  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n1054 ), .A3(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n961 ) );
NOR3_X2 _AES_ENC_us11_U153  ( .A1(_AES_ENC_us11_n620 ), .A2(_AES_ENC_us11_n1074 ), .A3(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n671 ) );
NOR2_X2 _AES_ENC_us11_U152  ( .A1(_AES_ENC_us11_n1057 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n1062 ) );
NOR2_X2 _AES_ENC_us11_U143  ( .A1(_AES_ENC_us11_n1055 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n1063 ) );
NOR2_X2 _AES_ENC_us11_U142  ( .A1(_AES_ENC_us11_n1060 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n1061 ) );
NOR4_X2 _AES_ENC_us11_U141  ( .A1(_AES_ENC_us11_n1064 ), .A2(_AES_ENC_us11_n1063 ), .A3(_AES_ENC_us11_n1062 ), .A4(_AES_ENC_us11_n1061 ), .ZN(_AES_ENC_us11_n1065 ) );
NOR3_X2 _AES_ENC_us11_U140  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n1120 ), .A3(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n918 ) );
NOR3_X2 _AES_ENC_us11_U132  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n573 ), .A3(_AES_ENC_us11_n1013 ), .ZN(_AES_ENC_us11_n917 ) );
NOR2_X2 _AES_ENC_us11_U131  ( .A1(_AES_ENC_us11_n914 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n915 ) );
NOR4_X2 _AES_ENC_us11_U130  ( .A1(_AES_ENC_us11_n918 ), .A2(_AES_ENC_us11_n917 ), .A3(_AES_ENC_us11_n916 ), .A4(_AES_ENC_us11_n915 ), .ZN(_AES_ENC_us11_n919 ) );
NOR2_X2 _AES_ENC_us11_U129  ( .A1(_AES_ENC_us11_n735 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n687 ) );
NOR2_X2 _AES_ENC_us11_U128  ( .A1(_AES_ENC_us11_n684 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n688 ) );
NOR2_X2 _AES_ENC_us11_U127  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n600 ), .ZN(_AES_ENC_us11_n686 ) );
NOR4_X2 _AES_ENC_us11_U126  ( .A1(_AES_ENC_us11_n688 ), .A2(_AES_ENC_us11_n687 ), .A3(_AES_ENC_us11_n686 ), .A4(_AES_ENC_us11_n685 ), .ZN(_AES_ENC_us11_n689 ) );
NOR2_X2 _AES_ENC_us11_U121  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n595 ), .ZN(_AES_ENC_us11_n858 ) );
NOR2_X2 _AES_ENC_us11_U120  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n855 ), .ZN(_AES_ENC_us11_n857 ) );
NOR2_X2 _AES_ENC_us11_U119  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n587 ), .ZN(_AES_ENC_us11_n856 ) );
NOR4_X2 _AES_ENC_us11_U118  ( .A1(_AES_ENC_us11_n858 ), .A2(_AES_ENC_us11_n857 ), .A3(_AES_ENC_us11_n856 ), .A4(_AES_ENC_us11_n958 ), .ZN(_AES_ENC_us11_n859 ) );
NOR2_X2 _AES_ENC_us11_U117  ( .A1(_AES_ENC_us11_n616 ), .A2(_AES_ENC_us11_n580 ), .ZN(_AES_ENC_us11_n771 ) );
NOR2_X2 _AES_ENC_us11_U116  ( .A1(_AES_ENC_us11_n1103 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n772 ) );
NOR2_X2 _AES_ENC_us11_U115  ( .A1(_AES_ENC_us11_n610 ), .A2(_AES_ENC_us11_n599 ), .ZN(_AES_ENC_us11_n773 ) );
NOR4_X2 _AES_ENC_us11_U106  ( .A1(_AES_ENC_us11_n773 ), .A2(_AES_ENC_us11_n772 ), .A3(_AES_ENC_us11_n771 ), .A4(_AES_ENC_us11_n770 ), .ZN(_AES_ENC_us11_n774 ) );
NOR2_X2 _AES_ENC_us11_U105  ( .A1(_AES_ENC_us11_n780 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n784 ) );
NOR2_X2 _AES_ENC_us11_U104  ( .A1(_AES_ENC_us11_n1117 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n782 ) );
NOR2_X2 _AES_ENC_us11_U103  ( .A1(_AES_ENC_us11_n781 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n783 ) );
NOR4_X2 _AES_ENC_us11_U102  ( .A1(_AES_ENC_us11_n880 ), .A2(_AES_ENC_us11_n784 ), .A3(_AES_ENC_us11_n783 ), .A4(_AES_ENC_us11_n782 ), .ZN(_AES_ENC_us11_n785 ) );
NOR2_X2 _AES_ENC_us11_U101  ( .A1(_AES_ENC_us11_n583 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n814 ) );
NOR2_X2 _AES_ENC_us11_U100  ( .A1(_AES_ENC_us11_n907 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n813 ) );
NOR3_X2 _AES_ENC_us11_U95  ( .A1(_AES_ENC_us11_n606 ), .A2(_AES_ENC_us11_n1058 ), .A3(_AES_ENC_us11_n1059 ), .ZN(_AES_ENC_us11_n815 ) );
NOR4_X2 _AES_ENC_us11_U94  ( .A1(_AES_ENC_us11_n815 ), .A2(_AES_ENC_us11_n814 ), .A3(_AES_ENC_us11_n813 ), .A4(_AES_ENC_us11_n812 ), .ZN(_AES_ENC_us11_n816 ) );
NOR2_X2 _AES_ENC_us11_U93  ( .A1(_AES_ENC_us11_n617 ), .A2(_AES_ENC_us11_n569 ), .ZN(_AES_ENC_us11_n721 ) );
NOR2_X2 _AES_ENC_us11_U92  ( .A1(_AES_ENC_us11_n1031 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n723 ) );
NOR2_X2 _AES_ENC_us11_U91  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n1096 ), .ZN(_AES_ENC_us11_n722 ) );
NOR4_X2 _AES_ENC_us11_U90  ( .A1(_AES_ENC_us11_n724 ), .A2(_AES_ENC_us11_n723 ), .A3(_AES_ENC_us11_n722 ), .A4(_AES_ENC_us11_n721 ), .ZN(_AES_ENC_us11_n725 ) );
NOR2_X2 _AES_ENC_us11_U89  ( .A1(_AES_ENC_us11_n911 ), .A2(_AES_ENC_us11_n990 ), .ZN(_AES_ENC_us11_n1009 ) );
NOR2_X2 _AES_ENC_us11_U88  ( .A1(_AES_ENC_us11_n1013 ), .A2(_AES_ENC_us11_n573 ), .ZN(_AES_ENC_us11_n1014 ) );
NOR2_X2 _AES_ENC_us11_U87  ( .A1(_AES_ENC_us11_n1014 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n1015 ) );
NOR4_X2 _AES_ENC_us11_U86  ( .A1(_AES_ENC_us11_n1016 ), .A2(_AES_ENC_us11_n1015 ), .A3(_AES_ENC_us11_n1119 ), .A4(_AES_ENC_us11_n1046 ), .ZN(_AES_ENC_us11_n1017 ) );
NOR2_X2 _AES_ENC_us11_U81  ( .A1(_AES_ENC_us11_n996 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n998 ) );
NOR2_X2 _AES_ENC_us11_U80  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n577 ), .ZN(_AES_ENC_us11_n1000 ) );
NOR2_X2 _AES_ENC_us11_U79  ( .A1(_AES_ENC_us11_n616 ), .A2(_AES_ENC_us11_n1096 ), .ZN(_AES_ENC_us11_n999 ) );
NOR4_X2 _AES_ENC_us11_U78  ( .A1(_AES_ENC_us11_n1000 ), .A2(_AES_ENC_us11_n999 ), .A3(_AES_ENC_us11_n998 ), .A4(_AES_ENC_us11_n997 ), .ZN(_AES_ENC_us11_n1001 ) );
NOR2_X2 _AES_ENC_us11_U74  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n1096 ), .ZN(_AES_ENC_us11_n697 ) );
NOR2_X2 _AES_ENC_us11_U73  ( .A1(_AES_ENC_us11_n620 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n958 ) );
NOR2_X2 _AES_ENC_us11_U72  ( .A1(_AES_ENC_us11_n911 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n983 ) );
NOR2_X2 _AES_ENC_us11_U71  ( .A1(_AES_ENC_us11_n1054 ), .A2(_AES_ENC_us11_n1103 ), .ZN(_AES_ENC_us11_n1031 ) );
INV_X4 _AES_ENC_us11_U65  ( .A(_AES_ENC_us11_n1050 ), .ZN(_AES_ENC_us11_n612 ) );
INV_X4 _AES_ENC_us11_U64  ( .A(_AES_ENC_us11_n1072 ), .ZN(_AES_ENC_us11_n605 ) );
INV_X4 _AES_ENC_us11_U63  ( .A(_AES_ENC_us11_n1073 ), .ZN(_AES_ENC_us11_n604 ) );
NOR2_X2 _AES_ENC_us11_U62  ( .A1(_AES_ENC_us11_n582 ), .A2(_AES_ENC_us11_n613 ), .ZN(_AES_ENC_us11_n880 ) );
NOR3_X2 _AES_ENC_us11_U61  ( .A1(_AES_ENC_us11_n826 ), .A2(_AES_ENC_us11_n1121 ), .A3(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n946 ) );
INV_X4 _AES_ENC_us11_U59  ( .A(_AES_ENC_us11_n1010 ), .ZN(_AES_ENC_us11_n608 ) );
NOR3_X2 _AES_ENC_us11_U58  ( .A1(_AES_ENC_us11_n573 ), .A2(_AES_ENC_us11_n1029 ), .A3(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n1119 ) );
INV_X4 _AES_ENC_us11_U57  ( .A(_AES_ENC_us11_n956 ), .ZN(_AES_ENC_us11_n615 ) );
NOR2_X2 _AES_ENC_us11_U50  ( .A1(_AES_ENC_us11_n623 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n1013 ) );
NOR2_X2 _AES_ENC_us11_U49  ( .A1(_AES_ENC_us11_n620 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n910 ) );
NOR2_X2 _AES_ENC_us11_U48  ( .A1(_AES_ENC_us11_n569 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n1091 ) );
NOR2_X2 _AES_ENC_us11_U47  ( .A1(_AES_ENC_us11_n622 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n990 ) );
NOR2_X2 _AES_ENC_us11_U46  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_us11_n1121 ), .ZN(_AES_ENC_us11_n996 ) );
NOR2_X2 _AES_ENC_us11_U45  ( .A1(_AES_ENC_us11_n610 ), .A2(_AES_ENC_us11_n600 ), .ZN(_AES_ENC_us11_n628 ) );
NOR2_X2 _AES_ENC_us11_U44  ( .A1(_AES_ENC_us11_n576 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n866 ) );
NOR2_X2 _AES_ENC_us11_U43  ( .A1(_AES_ENC_us11_n603 ), .A2(_AES_ENC_us11_n610 ), .ZN(_AES_ENC_us11_n1006 ) );
NOR2_X2 _AES_ENC_us11_U42  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n1117 ), .ZN(_AES_ENC_us11_n1118 ) );
NOR2_X2 _AES_ENC_us11_U41  ( .A1(_AES_ENC_us11_n1119 ), .A2(_AES_ENC_us11_n1118 ), .ZN(_AES_ENC_us11_n1127 ) );
NOR2_X2 _AES_ENC_us11_U36  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n594 ), .ZN(_AES_ENC_us11_n629 ) );
NOR2_X2 _AES_ENC_us11_U35  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n906 ), .ZN(_AES_ENC_us11_n909 ) );
NOR2_X2 _AES_ENC_us11_U34  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n597 ), .ZN(_AES_ENC_us11_n658 ) );
NOR2_X2 _AES_ENC_us11_U33  ( .A1(_AES_ENC_us11_n1116 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n695 ) );
NOR2_X2 _AES_ENC_us11_U32  ( .A1(_AES_ENC_us11_n1078 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n1083 ) );
NOR2_X2 _AES_ENC_us11_U31  ( .A1(_AES_ENC_us11_n941 ), .A2(_AES_ENC_us11_n608 ), .ZN(_AES_ENC_us11_n724 ) );
NOR2_X2 _AES_ENC_us11_U30  ( .A1(_AES_ENC_us11_n598 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n1107 ) );
NOR2_X2 _AES_ENC_us11_U29  ( .A1(_AES_ENC_us11_n576 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n840 ) );
NOR2_X2 _AES_ENC_us11_U24  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n593 ), .ZN(_AES_ENC_us11_n633 ) );
NOR2_X2 _AES_ENC_us11_U23  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n1080 ), .ZN(_AES_ENC_us11_n1081 ) );
NOR2_X2 _AES_ENC_us11_U21  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n1045 ), .ZN(_AES_ENC_us11_n812 ) );
NOR2_X2 _AES_ENC_us11_U20  ( .A1(_AES_ENC_us11_n1009 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n960 ) );
NOR2_X2 _AES_ENC_us11_U19  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n601 ), .ZN(_AES_ENC_us11_n982 ) );
NOR2_X2 _AES_ENC_us11_U18  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n594 ), .ZN(_AES_ENC_us11_n757 ) );
NOR2_X2 _AES_ENC_us11_U17  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n590 ), .ZN(_AES_ENC_us11_n698 ) );
NOR2_X2 _AES_ENC_us11_U16  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n619 ), .ZN(_AES_ENC_us11_n708 ) );
NOR2_X2 _AES_ENC_us11_U15  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n582 ), .ZN(_AES_ENC_us11_n770 ) );
NOR2_X2 _AES_ENC_us11_U10  ( .A1(_AES_ENC_us11_n619 ), .A2(_AES_ENC_us11_n604 ), .ZN(_AES_ENC_us11_n803 ) );
NOR2_X2 _AES_ENC_us11_U9  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n881 ), .ZN(_AES_ENC_us11_n711 ) );
NOR2_X2 _AES_ENC_us11_U8  ( .A1(_AES_ENC_us11_n615 ), .A2(_AES_ENC_us11_n582 ), .ZN(_AES_ENC_us11_n867 ) );
NOR2_X2 _AES_ENC_us11_U7  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n599 ), .ZN(_AES_ENC_us11_n804 ) );
NOR2_X2 _AES_ENC_us11_U6  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n620 ), .ZN(_AES_ENC_us11_n1046 ) );
OR2_X4 _AES_ENC_us11_U5  ( .A1(_AES_ENC_us11_n624 ), .A2(_AES_ENC_sa11[1]),.ZN(_AES_ENC_us11_n570 ) );
OR2_X4 _AES_ENC_us11_U4  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_sa11[4]),.ZN(_AES_ENC_us11_n569 ) );
NAND2_X2 _AES_ENC_us11_U514  ( .A1(_AES_ENC_us11_n1121 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n1030 ) );
AND2_X2 _AES_ENC_us11_U513  ( .A1(_AES_ENC_us11_n597 ), .A2(_AES_ENC_us11_n1030 ), .ZN(_AES_ENC_us11_n1049 ) );
NAND2_X2 _AES_ENC_us11_U511  ( .A1(_AES_ENC_us11_n1049 ), .A2(_AES_ENC_us11_n794 ), .ZN(_AES_ENC_us11_n637 ) );
AND2_X2 _AES_ENC_us11_U493  ( .A1(_AES_ENC_us11_n779 ), .A2(_AES_ENC_us11_n996 ), .ZN(_AES_ENC_us11_n632 ) );
NAND4_X2 _AES_ENC_us11_U485  ( .A1(_AES_ENC_us11_n637 ), .A2(_AES_ENC_us11_n636 ), .A3(_AES_ENC_us11_n635 ), .A4(_AES_ENC_us11_n634 ), .ZN(_AES_ENC_us11_n638 ) );
NAND2_X2 _AES_ENC_us11_U484  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n638 ), .ZN(_AES_ENC_us11_n679 ) );
NAND2_X2 _AES_ENC_us11_U481  ( .A1(_AES_ENC_us11_n1094 ), .A2(_AES_ENC_us11_n591 ), .ZN(_AES_ENC_us11_n648 ) );
NAND2_X2 _AES_ENC_us11_U476  ( .A1(_AES_ENC_us11_n601 ), .A2(_AES_ENC_us11_n590 ), .ZN(_AES_ENC_us11_n762 ) );
NAND2_X2 _AES_ENC_us11_U475  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n762 ), .ZN(_AES_ENC_us11_n647 ) );
NAND4_X2 _AES_ENC_us11_U457  ( .A1(_AES_ENC_us11_n648 ), .A2(_AES_ENC_us11_n647 ), .A3(_AES_ENC_us11_n646 ), .A4(_AES_ENC_us11_n645 ), .ZN(_AES_ENC_us11_n649 ) );
NAND2_X2 _AES_ENC_us11_U456  ( .A1(_AES_ENC_sa11[0]), .A2(_AES_ENC_us11_n649 ), .ZN(_AES_ENC_us11_n665 ) );
NAND2_X2 _AES_ENC_us11_U454  ( .A1(_AES_ENC_us11_n596 ), .A2(_AES_ENC_us11_n623 ), .ZN(_AES_ENC_us11_n855 ) );
NAND2_X2 _AES_ENC_us11_U453  ( .A1(_AES_ENC_us11_n587 ), .A2(_AES_ENC_us11_n855 ), .ZN(_AES_ENC_us11_n821 ) );
NAND2_X2 _AES_ENC_us11_U452  ( .A1(_AES_ENC_us11_n1093 ), .A2(_AES_ENC_us11_n821 ), .ZN(_AES_ENC_us11_n662 ) );
NAND2_X2 _AES_ENC_us11_U451  ( .A1(_AES_ENC_us11_n619 ), .A2(_AES_ENC_us11_n589 ), .ZN(_AES_ENC_us11_n650 ) );
NAND2_X2 _AES_ENC_us11_U450  ( .A1(_AES_ENC_us11_n956 ), .A2(_AES_ENC_us11_n650 ), .ZN(_AES_ENC_us11_n661 ) );
NAND2_X2 _AES_ENC_us11_U449  ( .A1(_AES_ENC_us11_n626 ), .A2(_AES_ENC_us11_n627 ), .ZN(_AES_ENC_us11_n839 ) );
OR2_X2 _AES_ENC_us11_U446  ( .A1(_AES_ENC_us11_n839 ), .A2(_AES_ENC_us11_n932 ), .ZN(_AES_ENC_us11_n656 ) );
NAND2_X2 _AES_ENC_us11_U445  ( .A1(_AES_ENC_us11_n621 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n1096 ) );
NAND2_X2 _AES_ENC_us11_U444  ( .A1(_AES_ENC_us11_n1030 ), .A2(_AES_ENC_us11_n1096 ), .ZN(_AES_ENC_us11_n651 ) );
NAND2_X2 _AES_ENC_us11_U443  ( .A1(_AES_ENC_us11_n1114 ), .A2(_AES_ENC_us11_n651 ), .ZN(_AES_ENC_us11_n655 ) );
OR3_X2 _AES_ENC_us11_U440  ( .A1(_AES_ENC_us11_n1079 ), .A2(_AES_ENC_sa11[7]), .A3(_AES_ENC_us11_n626 ), .ZN(_AES_ENC_us11_n654 ));
NAND2_X2 _AES_ENC_us11_U439  ( .A1(_AES_ENC_us11_n593 ), .A2(_AES_ENC_us11_n601 ), .ZN(_AES_ENC_us11_n652 ) );
NAND4_X2 _AES_ENC_us11_U437  ( .A1(_AES_ENC_us11_n656 ), .A2(_AES_ENC_us11_n655 ), .A3(_AES_ENC_us11_n654 ), .A4(_AES_ENC_us11_n653 ), .ZN(_AES_ENC_us11_n657 ) );
NAND2_X2 _AES_ENC_us11_U436  ( .A1(_AES_ENC_sa11[2]), .A2(_AES_ENC_us11_n657 ), .ZN(_AES_ENC_us11_n660 ) );
NAND4_X2 _AES_ENC_us11_U432  ( .A1(_AES_ENC_us11_n662 ), .A2(_AES_ENC_us11_n661 ), .A3(_AES_ENC_us11_n660 ), .A4(_AES_ENC_us11_n659 ), .ZN(_AES_ENC_us11_n663 ) );
NAND2_X2 _AES_ENC_us11_U431  ( .A1(_AES_ENC_us11_n663 ), .A2(_AES_ENC_us11_n574 ), .ZN(_AES_ENC_us11_n664 ) );
NAND2_X2 _AES_ENC_us11_U430  ( .A1(_AES_ENC_us11_n665 ), .A2(_AES_ENC_us11_n664 ), .ZN(_AES_ENC_us11_n666 ) );
NAND2_X2 _AES_ENC_us11_U429  ( .A1(_AES_ENC_sa11[6]), .A2(_AES_ENC_us11_n666 ), .ZN(_AES_ENC_us11_n678 ) );
NAND2_X2 _AES_ENC_us11_U426  ( .A1(_AES_ENC_us11_n735 ), .A2(_AES_ENC_us11_n1093 ), .ZN(_AES_ENC_us11_n675 ) );
NAND2_X2 _AES_ENC_us11_U425  ( .A1(_AES_ENC_us11_n588 ), .A2(_AES_ENC_us11_n597 ), .ZN(_AES_ENC_us11_n1045 ) );
OR2_X2 _AES_ENC_us11_U424  ( .A1(_AES_ENC_us11_n1045 ), .A2(_AES_ENC_us11_n605 ), .ZN(_AES_ENC_us11_n674 ) );
NAND2_X2 _AES_ENC_us11_U423  ( .A1(_AES_ENC_sa11[1]), .A2(_AES_ENC_us11_n620 ), .ZN(_AES_ENC_us11_n667 ) );
NAND2_X2 _AES_ENC_us11_U422  ( .A1(_AES_ENC_us11_n619 ), .A2(_AES_ENC_us11_n667 ), .ZN(_AES_ENC_us11_n1071 ) );
NAND4_X2 _AES_ENC_us11_U412  ( .A1(_AES_ENC_us11_n675 ), .A2(_AES_ENC_us11_n674 ), .A3(_AES_ENC_us11_n673 ), .A4(_AES_ENC_us11_n672 ), .ZN(_AES_ENC_us11_n676 ) );
NAND2_X2 _AES_ENC_us11_U411  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n676 ), .ZN(_AES_ENC_us11_n677 ) );
NAND2_X2 _AES_ENC_us11_U408  ( .A1(_AES_ENC_us11_n800 ), .A2(_AES_ENC_us11_n1022 ), .ZN(_AES_ENC_us11_n680 ) );
NAND2_X2 _AES_ENC_us11_U407  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n680 ), .ZN(_AES_ENC_us11_n681 ) );
AND2_X2 _AES_ENC_us11_U402  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n684 ), .ZN(_AES_ENC_us11_n682 ) );
NAND4_X2 _AES_ENC_us11_U395  ( .A1(_AES_ENC_us11_n691 ), .A2(_AES_ENC_us11_n581 ), .A3(_AES_ENC_us11_n690 ), .A4(_AES_ENC_us11_n689 ), .ZN(_AES_ENC_us11_n692 ) );
NAND2_X2 _AES_ENC_us11_U394  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n692 ), .ZN(_AES_ENC_us11_n733 ) );
NAND2_X2 _AES_ENC_us11_U392  ( .A1(_AES_ENC_us11_n977 ), .A2(_AES_ENC_us11_n1050 ), .ZN(_AES_ENC_us11_n702 ) );
NAND2_X2 _AES_ENC_us11_U391  ( .A1(_AES_ENC_us11_n1093 ), .A2(_AES_ENC_us11_n1045 ), .ZN(_AES_ENC_us11_n701 ) );
NAND4_X2 _AES_ENC_us11_U381  ( .A1(_AES_ENC_us11_n702 ), .A2(_AES_ENC_us11_n701 ), .A3(_AES_ENC_us11_n700 ), .A4(_AES_ENC_us11_n699 ), .ZN(_AES_ENC_us11_n703 ) );
NAND2_X2 _AES_ENC_us11_U380  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n703 ), .ZN(_AES_ENC_us11_n732 ) );
AND2_X2 _AES_ENC_us11_U379  ( .A1(_AES_ENC_sa11[0]), .A2(_AES_ENC_sa11[6]),.ZN(_AES_ENC_us11_n1113 ) );
NAND2_X2 _AES_ENC_us11_U378  ( .A1(_AES_ENC_us11_n601 ), .A2(_AES_ENC_us11_n1030 ), .ZN(_AES_ENC_us11_n881 ) );
NAND2_X2 _AES_ENC_us11_U377  ( .A1(_AES_ENC_us11_n1093 ), .A2(_AES_ENC_us11_n881 ), .ZN(_AES_ENC_us11_n715 ) );
NAND2_X2 _AES_ENC_us11_U376  ( .A1(_AES_ENC_us11_n1010 ), .A2(_AES_ENC_us11_n600 ), .ZN(_AES_ENC_us11_n714 ) );
NAND2_X2 _AES_ENC_us11_U375  ( .A1(_AES_ENC_us11_n855 ), .A2(_AES_ENC_us11_n588 ), .ZN(_AES_ENC_us11_n1117 ) );
XNOR2_X2 _AES_ENC_us11_U371  ( .A(_AES_ENC_us11_n611 ), .B(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n824 ) );
NAND4_X2 _AES_ENC_us11_U362  ( .A1(_AES_ENC_us11_n715 ), .A2(_AES_ENC_us11_n714 ), .A3(_AES_ENC_us11_n713 ), .A4(_AES_ENC_us11_n712 ), .ZN(_AES_ENC_us11_n716 ) );
NAND2_X2 _AES_ENC_us11_U361  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n716 ), .ZN(_AES_ENC_us11_n731 ) );
AND2_X2 _AES_ENC_us11_U360  ( .A1(_AES_ENC_sa11[6]), .A2(_AES_ENC_us11_n574 ), .ZN(_AES_ENC_us11_n1131 ) );
NAND2_X2 _AES_ENC_us11_U359  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n717 ) );
NAND2_X2 _AES_ENC_us11_U358  ( .A1(_AES_ENC_us11_n1029 ), .A2(_AES_ENC_us11_n717 ), .ZN(_AES_ENC_us11_n728 ) );
NAND2_X2 _AES_ENC_us11_U357  ( .A1(_AES_ENC_sa11[1]), .A2(_AES_ENC_us11_n624 ), .ZN(_AES_ENC_us11_n1097 ) );
NAND2_X2 _AES_ENC_us11_U356  ( .A1(_AES_ENC_us11_n603 ), .A2(_AES_ENC_us11_n1097 ), .ZN(_AES_ENC_us11_n718 ) );
NAND2_X2 _AES_ENC_us11_U355  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n718 ), .ZN(_AES_ENC_us11_n727 ) );
NAND4_X2 _AES_ENC_us11_U344  ( .A1(_AES_ENC_us11_n728 ), .A2(_AES_ENC_us11_n727 ), .A3(_AES_ENC_us11_n726 ), .A4(_AES_ENC_us11_n725 ), .ZN(_AES_ENC_us11_n729 ) );
NAND2_X2 _AES_ENC_us11_U343  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n729 ), .ZN(_AES_ENC_us11_n730 ) );
NAND4_X2 _AES_ENC_us11_U342  ( .A1(_AES_ENC_us11_n733 ), .A2(_AES_ENC_us11_n732 ), .A3(_AES_ENC_us11_n731 ), .A4(_AES_ENC_us11_n730 ), .ZN(_AES_ENC_sa11_sub[1] ) );
NAND2_X2 _AES_ENC_us11_U341  ( .A1(_AES_ENC_sa11[7]), .A2(_AES_ENC_us11_n611 ), .ZN(_AES_ENC_us11_n734 ) );
NAND2_X2 _AES_ENC_us11_U340  ( .A1(_AES_ENC_us11_n734 ), .A2(_AES_ENC_us11_n607 ), .ZN(_AES_ENC_us11_n738 ) );
OR4_X2 _AES_ENC_us11_U339  ( .A1(_AES_ENC_us11_n738 ), .A2(_AES_ENC_us11_n626 ), .A3(_AES_ENC_us11_n826 ), .A4(_AES_ENC_us11_n1121 ), .ZN(_AES_ENC_us11_n746 ) );
NAND2_X2 _AES_ENC_us11_U337  ( .A1(_AES_ENC_us11_n1100 ), .A2(_AES_ENC_us11_n587 ), .ZN(_AES_ENC_us11_n992 ) );
OR2_X2 _AES_ENC_us11_U336  ( .A1(_AES_ENC_us11_n610 ), .A2(_AES_ENC_us11_n735 ), .ZN(_AES_ENC_us11_n737 ) );
NAND2_X2 _AES_ENC_us11_U334  ( .A1(_AES_ENC_us11_n619 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n753 ) );
NAND2_X2 _AES_ENC_us11_U333  ( .A1(_AES_ENC_us11_n582 ), .A2(_AES_ENC_us11_n753 ), .ZN(_AES_ENC_us11_n1080 ) );
NAND2_X2 _AES_ENC_us11_U332  ( .A1(_AES_ENC_us11_n1048 ), .A2(_AES_ENC_us11_n576 ), .ZN(_AES_ENC_us11_n736 ) );
NAND2_X2 _AES_ENC_us11_U331  ( .A1(_AES_ENC_us11_n737 ), .A2(_AES_ENC_us11_n736 ), .ZN(_AES_ENC_us11_n739 ) );
NAND2_X2 _AES_ENC_us11_U330  ( .A1(_AES_ENC_us11_n739 ), .A2(_AES_ENC_us11_n738 ), .ZN(_AES_ENC_us11_n745 ) );
NAND2_X2 _AES_ENC_us11_U326  ( .A1(_AES_ENC_us11_n1096 ), .A2(_AES_ENC_us11_n590 ), .ZN(_AES_ENC_us11_n906 ) );
NAND4_X2 _AES_ENC_us11_U323  ( .A1(_AES_ENC_us11_n746 ), .A2(_AES_ENC_us11_n992 ), .A3(_AES_ENC_us11_n745 ), .A4(_AES_ENC_us11_n744 ), .ZN(_AES_ENC_us11_n747 ) );
NAND2_X2 _AES_ENC_us11_U322  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n747 ), .ZN(_AES_ENC_us11_n793 ) );
NAND2_X2 _AES_ENC_us11_U321  ( .A1(_AES_ENC_us11_n584 ), .A2(_AES_ENC_us11_n855 ), .ZN(_AES_ENC_us11_n748 ) );
NAND2_X2 _AES_ENC_us11_U320  ( .A1(_AES_ENC_us11_n956 ), .A2(_AES_ENC_us11_n748 ), .ZN(_AES_ENC_us11_n760 ) );
NAND2_X2 _AES_ENC_us11_U313  ( .A1(_AES_ENC_us11_n590 ), .A2(_AES_ENC_us11_n753 ), .ZN(_AES_ENC_us11_n1023 ) );
NAND4_X2 _AES_ENC_us11_U308  ( .A1(_AES_ENC_us11_n760 ), .A2(_AES_ENC_us11_n992 ), .A3(_AES_ENC_us11_n759 ), .A4(_AES_ENC_us11_n758 ), .ZN(_AES_ENC_us11_n761 ) );
NAND2_X2 _AES_ENC_us11_U307  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n761 ), .ZN(_AES_ENC_us11_n792 ) );
NAND2_X2 _AES_ENC_us11_U306  ( .A1(_AES_ENC_us11_n584 ), .A2(_AES_ENC_us11_n603 ), .ZN(_AES_ENC_us11_n989 ) );
NAND2_X2 _AES_ENC_us11_U305  ( .A1(_AES_ENC_us11_n1050 ), .A2(_AES_ENC_us11_n989 ), .ZN(_AES_ENC_us11_n777 ) );
NAND2_X2 _AES_ENC_us11_U304  ( .A1(_AES_ENC_us11_n1093 ), .A2(_AES_ENC_us11_n762 ), .ZN(_AES_ENC_us11_n776 ) );
XNOR2_X2 _AES_ENC_us11_U301  ( .A(_AES_ENC_sa11[7]), .B(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n959 ) );
NAND4_X2 _AES_ENC_us11_U289  ( .A1(_AES_ENC_us11_n777 ), .A2(_AES_ENC_us11_n776 ), .A3(_AES_ENC_us11_n775 ), .A4(_AES_ENC_us11_n774 ), .ZN(_AES_ENC_us11_n778 ) );
NAND2_X2 _AES_ENC_us11_U288  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n778 ), .ZN(_AES_ENC_us11_n791 ) );
NAND2_X2 _AES_ENC_us11_U287  ( .A1(_AES_ENC_us11_n1056 ), .A2(_AES_ENC_us11_n1050 ), .ZN(_AES_ENC_us11_n788 ) );
NAND2_X2 _AES_ENC_us11_U286  ( .A1(_AES_ENC_us11_n1091 ), .A2(_AES_ENC_us11_n779 ), .ZN(_AES_ENC_us11_n787 ) );
NAND2_X2 _AES_ENC_us11_U285  ( .A1(_AES_ENC_us11_n956 ), .A2(_AES_ENC_sa11[1]), .ZN(_AES_ENC_us11_n786 ) );
NAND4_X2 _AES_ENC_us11_U278  ( .A1(_AES_ENC_us11_n788 ), .A2(_AES_ENC_us11_n787 ), .A3(_AES_ENC_us11_n786 ), .A4(_AES_ENC_us11_n785 ), .ZN(_AES_ENC_us11_n789 ) );
NAND2_X2 _AES_ENC_us11_U277  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n789 ), .ZN(_AES_ENC_us11_n790 ) );
NAND4_X2 _AES_ENC_us11_U276  ( .A1(_AES_ENC_us11_n793 ), .A2(_AES_ENC_us11_n792 ), .A3(_AES_ENC_us11_n791 ), .A4(_AES_ENC_us11_n790 ), .ZN(_AES_ENC_sa11_sub[2] ) );
NAND2_X2 _AES_ENC_us11_U275  ( .A1(_AES_ENC_us11_n1059 ), .A2(_AES_ENC_us11_n794 ), .ZN(_AES_ENC_us11_n810 ) );
NAND2_X2 _AES_ENC_us11_U274  ( .A1(_AES_ENC_us11_n1049 ), .A2(_AES_ENC_us11_n956 ), .ZN(_AES_ENC_us11_n809 ) );
OR2_X2 _AES_ENC_us11_U266  ( .A1(_AES_ENC_us11_n1096 ), .A2(_AES_ENC_us11_n606 ), .ZN(_AES_ENC_us11_n802 ) );
NAND2_X2 _AES_ENC_us11_U265  ( .A1(_AES_ENC_us11_n1053 ), .A2(_AES_ENC_us11_n800 ), .ZN(_AES_ENC_us11_n801 ) );
NAND2_X2 _AES_ENC_us11_U264  ( .A1(_AES_ENC_us11_n802 ), .A2(_AES_ENC_us11_n801 ), .ZN(_AES_ENC_us11_n805 ) );
NAND4_X2 _AES_ENC_us11_U261  ( .A1(_AES_ENC_us11_n810 ), .A2(_AES_ENC_us11_n809 ), .A3(_AES_ENC_us11_n808 ), .A4(_AES_ENC_us11_n807 ), .ZN(_AES_ENC_us11_n811 ) );
NAND2_X2 _AES_ENC_us11_U260  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n811 ), .ZN(_AES_ENC_us11_n852 ) );
OR2_X2 _AES_ENC_us11_U259  ( .A1(_AES_ENC_us11_n1023 ), .A2(_AES_ENC_us11_n617 ), .ZN(_AES_ENC_us11_n819 ) );
OR2_X2 _AES_ENC_us11_U257  ( .A1(_AES_ENC_us11_n570 ), .A2(_AES_ENC_us11_n930 ), .ZN(_AES_ENC_us11_n818 ) );
NAND2_X2 _AES_ENC_us11_U256  ( .A1(_AES_ENC_us11_n1013 ), .A2(_AES_ENC_us11_n1094 ), .ZN(_AES_ENC_us11_n817 ) );
NAND4_X2 _AES_ENC_us11_U249  ( .A1(_AES_ENC_us11_n819 ), .A2(_AES_ENC_us11_n818 ), .A3(_AES_ENC_us11_n817 ), .A4(_AES_ENC_us11_n816 ), .ZN(_AES_ENC_us11_n820 ) );
NAND2_X2 _AES_ENC_us11_U248  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n820 ), .ZN(_AES_ENC_us11_n851 ) );
NAND2_X2 _AES_ENC_us11_U247  ( .A1(_AES_ENC_us11_n956 ), .A2(_AES_ENC_us11_n1080 ), .ZN(_AES_ENC_us11_n835 ) );
NAND2_X2 _AES_ENC_us11_U246  ( .A1(_AES_ENC_us11_n570 ), .A2(_AES_ENC_us11_n1030 ), .ZN(_AES_ENC_us11_n1047 ) );
OR2_X2 _AES_ENC_us11_U245  ( .A1(_AES_ENC_us11_n1047 ), .A2(_AES_ENC_us11_n612 ), .ZN(_AES_ENC_us11_n834 ) );
NAND2_X2 _AES_ENC_us11_U244  ( .A1(_AES_ENC_us11_n1072 ), .A2(_AES_ENC_us11_n589 ), .ZN(_AES_ENC_us11_n833 ) );
NAND4_X2 _AES_ENC_us11_U233  ( .A1(_AES_ENC_us11_n835 ), .A2(_AES_ENC_us11_n834 ), .A3(_AES_ENC_us11_n833 ), .A4(_AES_ENC_us11_n832 ), .ZN(_AES_ENC_us11_n836 ) );
NAND2_X2 _AES_ENC_us11_U232  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n836 ), .ZN(_AES_ENC_us11_n850 ) );
NAND2_X2 _AES_ENC_us11_U231  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n623 ), .ZN(_AES_ENC_us11_n847 ) );
NAND2_X2 _AES_ENC_us11_U230  ( .A1(_AES_ENC_us11_n1050 ), .A2(_AES_ENC_us11_n1071 ), .ZN(_AES_ENC_us11_n846 ) );
OR2_X2 _AES_ENC_us11_U224  ( .A1(_AES_ENC_us11_n1053 ), .A2(_AES_ENC_us11_n911 ), .ZN(_AES_ENC_us11_n1077 ) );
NAND4_X2 _AES_ENC_us11_U220  ( .A1(_AES_ENC_us11_n847 ), .A2(_AES_ENC_us11_n846 ), .A3(_AES_ENC_us11_n845 ), .A4(_AES_ENC_us11_n844 ), .ZN(_AES_ENC_us11_n848 ) );
NAND2_X2 _AES_ENC_us11_U219  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n848 ), .ZN(_AES_ENC_us11_n849 ) );
NAND4_X2 _AES_ENC_us11_U218  ( .A1(_AES_ENC_us11_n852 ), .A2(_AES_ENC_us11_n851 ), .A3(_AES_ENC_us11_n850 ), .A4(_AES_ENC_us11_n849 ), .ZN(_AES_ENC_sa11_sub[3] ) );
NAND2_X2 _AES_ENC_us11_U216  ( .A1(_AES_ENC_us11_n1009 ), .A2(_AES_ENC_us11_n1072 ), .ZN(_AES_ENC_us11_n862 ) );
NAND2_X2 _AES_ENC_us11_U215  ( .A1(_AES_ENC_us11_n603 ), .A2(_AES_ENC_us11_n577 ), .ZN(_AES_ENC_us11_n853 ) );
NAND2_X2 _AES_ENC_us11_U214  ( .A1(_AES_ENC_us11_n1050 ), .A2(_AES_ENC_us11_n853 ), .ZN(_AES_ENC_us11_n861 ) );
NAND4_X2 _AES_ENC_us11_U206  ( .A1(_AES_ENC_us11_n862 ), .A2(_AES_ENC_us11_n861 ), .A3(_AES_ENC_us11_n860 ), .A4(_AES_ENC_us11_n859 ), .ZN(_AES_ENC_us11_n863 ) );
NAND2_X2 _AES_ENC_us11_U205  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n863 ), .ZN(_AES_ENC_us11_n905 ) );
NAND2_X2 _AES_ENC_us11_U204  ( .A1(_AES_ENC_us11_n1010 ), .A2(_AES_ENC_us11_n989 ), .ZN(_AES_ENC_us11_n874 ) );
NAND2_X2 _AES_ENC_us11_U203  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n610 ), .ZN(_AES_ENC_us11_n864 ) );
NAND2_X2 _AES_ENC_us11_U202  ( .A1(_AES_ENC_us11_n929 ), .A2(_AES_ENC_us11_n864 ), .ZN(_AES_ENC_us11_n873 ) );
NAND4_X2 _AES_ENC_us11_U193  ( .A1(_AES_ENC_us11_n874 ), .A2(_AES_ENC_us11_n873 ), .A3(_AES_ENC_us11_n872 ), .A4(_AES_ENC_us11_n871 ), .ZN(_AES_ENC_us11_n875 ) );
NAND2_X2 _AES_ENC_us11_U192  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n875 ), .ZN(_AES_ENC_us11_n904 ) );
NAND2_X2 _AES_ENC_us11_U191  ( .A1(_AES_ENC_us11_n583 ), .A2(_AES_ENC_us11_n1050 ), .ZN(_AES_ENC_us11_n889 ) );
NAND2_X2 _AES_ENC_us11_U190  ( .A1(_AES_ENC_us11_n1093 ), .A2(_AES_ENC_us11_n587 ), .ZN(_AES_ENC_us11_n876 ) );
NAND2_X2 _AES_ENC_us11_U189  ( .A1(_AES_ENC_us11_n604 ), .A2(_AES_ENC_us11_n876 ), .ZN(_AES_ENC_us11_n877 ) );
NAND2_X2 _AES_ENC_us11_U188  ( .A1(_AES_ENC_us11_n877 ), .A2(_AES_ENC_us11_n623 ), .ZN(_AES_ENC_us11_n888 ) );
NAND4_X2 _AES_ENC_us11_U179  ( .A1(_AES_ENC_us11_n889 ), .A2(_AES_ENC_us11_n888 ), .A3(_AES_ENC_us11_n887 ), .A4(_AES_ENC_us11_n886 ), .ZN(_AES_ENC_us11_n890 ) );
NAND2_X2 _AES_ENC_us11_U178  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n890 ), .ZN(_AES_ENC_us11_n903 ) );
OR2_X2 _AES_ENC_us11_U177  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n1059 ), .ZN(_AES_ENC_us11_n900 ) );
NAND2_X2 _AES_ENC_us11_U176  ( .A1(_AES_ENC_us11_n1073 ), .A2(_AES_ENC_us11_n1047 ), .ZN(_AES_ENC_us11_n899 ) );
NAND2_X2 _AES_ENC_us11_U175  ( .A1(_AES_ENC_us11_n1094 ), .A2(_AES_ENC_us11_n595 ), .ZN(_AES_ENC_us11_n898 ) );
NAND4_X2 _AES_ENC_us11_U167  ( .A1(_AES_ENC_us11_n900 ), .A2(_AES_ENC_us11_n899 ), .A3(_AES_ENC_us11_n898 ), .A4(_AES_ENC_us11_n897 ), .ZN(_AES_ENC_us11_n901 ) );
NAND2_X2 _AES_ENC_us11_U166  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n901 ), .ZN(_AES_ENC_us11_n902 ) );
NAND4_X2 _AES_ENC_us11_U165  ( .A1(_AES_ENC_us11_n905 ), .A2(_AES_ENC_us11_n904 ), .A3(_AES_ENC_us11_n903 ), .A4(_AES_ENC_us11_n902 ), .ZN(_AES_ENC_sa11_sub[4] ) );
NAND2_X2 _AES_ENC_us11_U164  ( .A1(_AES_ENC_us11_n1094 ), .A2(_AES_ENC_us11_n599 ), .ZN(_AES_ENC_us11_n922 ) );
NAND2_X2 _AES_ENC_us11_U163  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n989 ), .ZN(_AES_ENC_us11_n921 ) );
NAND4_X2 _AES_ENC_us11_U151  ( .A1(_AES_ENC_us11_n922 ), .A2(_AES_ENC_us11_n921 ), .A3(_AES_ENC_us11_n920 ), .A4(_AES_ENC_us11_n919 ), .ZN(_AES_ENC_us11_n923 ) );
NAND2_X2 _AES_ENC_us11_U150  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n923 ), .ZN(_AES_ENC_us11_n972 ) );
NAND2_X2 _AES_ENC_us11_U149  ( .A1(_AES_ENC_us11_n582 ), .A2(_AES_ENC_us11_n619 ), .ZN(_AES_ENC_us11_n924 ) );
NAND2_X2 _AES_ENC_us11_U148  ( .A1(_AES_ENC_us11_n1073 ), .A2(_AES_ENC_us11_n924 ), .ZN(_AES_ENC_us11_n939 ) );
NAND2_X2 _AES_ENC_us11_U147  ( .A1(_AES_ENC_us11_n926 ), .A2(_AES_ENC_us11_n925 ), .ZN(_AES_ENC_us11_n927 ) );
NAND2_X2 _AES_ENC_us11_U146  ( .A1(_AES_ENC_us11_n606 ), .A2(_AES_ENC_us11_n927 ), .ZN(_AES_ENC_us11_n928 ) );
NAND2_X2 _AES_ENC_us11_U145  ( .A1(_AES_ENC_us11_n928 ), .A2(_AES_ENC_us11_n1080 ), .ZN(_AES_ENC_us11_n938 ) );
OR2_X2 _AES_ENC_us11_U144  ( .A1(_AES_ENC_us11_n1117 ), .A2(_AES_ENC_us11_n615 ), .ZN(_AES_ENC_us11_n937 ) );
NAND4_X2 _AES_ENC_us11_U139  ( .A1(_AES_ENC_us11_n939 ), .A2(_AES_ENC_us11_n938 ), .A3(_AES_ENC_us11_n937 ), .A4(_AES_ENC_us11_n936 ), .ZN(_AES_ENC_us11_n940 ) );
NAND2_X2 _AES_ENC_us11_U138  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n940 ), .ZN(_AES_ENC_us11_n971 ) );
OR2_X2 _AES_ENC_us11_U137  ( .A1(_AES_ENC_us11_n605 ), .A2(_AES_ENC_us11_n941 ), .ZN(_AES_ENC_us11_n954 ) );
NAND2_X2 _AES_ENC_us11_U136  ( .A1(_AES_ENC_us11_n1096 ), .A2(_AES_ENC_us11_n577 ), .ZN(_AES_ENC_us11_n942 ) );
NAND2_X2 _AES_ENC_us11_U135  ( .A1(_AES_ENC_us11_n1048 ), .A2(_AES_ENC_us11_n942 ), .ZN(_AES_ENC_us11_n943 ) );
NAND2_X2 _AES_ENC_us11_U134  ( .A1(_AES_ENC_us11_n612 ), .A2(_AES_ENC_us11_n943 ), .ZN(_AES_ENC_us11_n944 ) );
NAND2_X2 _AES_ENC_us11_U133  ( .A1(_AES_ENC_us11_n944 ), .A2(_AES_ENC_us11_n580 ), .ZN(_AES_ENC_us11_n953 ) );
NAND4_X2 _AES_ENC_us11_U125  ( .A1(_AES_ENC_us11_n954 ), .A2(_AES_ENC_us11_n953 ), .A3(_AES_ENC_us11_n952 ), .A4(_AES_ENC_us11_n951 ), .ZN(_AES_ENC_us11_n955 ) );
NAND2_X2 _AES_ENC_us11_U124  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n955 ), .ZN(_AES_ENC_us11_n970 ) );
NAND2_X2 _AES_ENC_us11_U123  ( .A1(_AES_ENC_us11_n1094 ), .A2(_AES_ENC_us11_n1071 ), .ZN(_AES_ENC_us11_n967 ) );
NAND2_X2 _AES_ENC_us11_U122  ( .A1(_AES_ENC_us11_n956 ), .A2(_AES_ENC_us11_n1030 ), .ZN(_AES_ENC_us11_n966 ) );
NAND4_X2 _AES_ENC_us11_U114  ( .A1(_AES_ENC_us11_n967 ), .A2(_AES_ENC_us11_n966 ), .A3(_AES_ENC_us11_n965 ), .A4(_AES_ENC_us11_n964 ), .ZN(_AES_ENC_us11_n968 ) );
NAND2_X2 _AES_ENC_us11_U113  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n968 ), .ZN(_AES_ENC_us11_n969 ) );
NAND4_X2 _AES_ENC_us11_U112  ( .A1(_AES_ENC_us11_n972 ), .A2(_AES_ENC_us11_n971 ), .A3(_AES_ENC_us11_n970 ), .A4(_AES_ENC_us11_n969 ), .ZN(_AES_ENC_sa11_sub[5] ) );
NAND2_X2 _AES_ENC_us11_U111  ( .A1(_AES_ENC_us11_n570 ), .A2(_AES_ENC_us11_n1097 ), .ZN(_AES_ENC_us11_n973 ) );
NAND2_X2 _AES_ENC_us11_U110  ( .A1(_AES_ENC_us11_n1073 ), .A2(_AES_ENC_us11_n973 ), .ZN(_AES_ENC_us11_n987 ) );
NAND2_X2 _AES_ENC_us11_U109  ( .A1(_AES_ENC_us11_n974 ), .A2(_AES_ENC_us11_n1077 ), .ZN(_AES_ENC_us11_n975 ) );
NAND2_X2 _AES_ENC_us11_U108  ( .A1(_AES_ENC_us11_n613 ), .A2(_AES_ENC_us11_n975 ), .ZN(_AES_ENC_us11_n976 ) );
NAND2_X2 _AES_ENC_us11_U107  ( .A1(_AES_ENC_us11_n977 ), .A2(_AES_ENC_us11_n976 ), .ZN(_AES_ENC_us11_n986 ) );
NAND4_X2 _AES_ENC_us11_U99  ( .A1(_AES_ENC_us11_n987 ), .A2(_AES_ENC_us11_n986 ), .A3(_AES_ENC_us11_n985 ), .A4(_AES_ENC_us11_n984 ), .ZN(_AES_ENC_us11_n988 ) );
NAND2_X2 _AES_ENC_us11_U98  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n988 ), .ZN(_AES_ENC_us11_n1044 ) );
NAND2_X2 _AES_ENC_us11_U97  ( .A1(_AES_ENC_us11_n1073 ), .A2(_AES_ENC_us11_n989 ), .ZN(_AES_ENC_us11_n1004 ) );
NAND2_X2 _AES_ENC_us11_U96  ( .A1(_AES_ENC_us11_n1092 ), .A2(_AES_ENC_us11_n619 ), .ZN(_AES_ENC_us11_n1003 ) );
NAND4_X2 _AES_ENC_us11_U85  ( .A1(_AES_ENC_us11_n1004 ), .A2(_AES_ENC_us11_n1003 ), .A3(_AES_ENC_us11_n1002 ), .A4(_AES_ENC_us11_n1001 ), .ZN(_AES_ENC_us11_n1005 ) );
NAND2_X2 _AES_ENC_us11_U84  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n1005 ), .ZN(_AES_ENC_us11_n1043 ) );
NAND2_X2 _AES_ENC_us11_U83  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n596 ), .ZN(_AES_ENC_us11_n1020 ) );
NAND2_X2 _AES_ENC_us11_U82  ( .A1(_AES_ENC_us11_n1050 ), .A2(_AES_ENC_us11_n624 ), .ZN(_AES_ENC_us11_n1019 ) );
NAND2_X2 _AES_ENC_us11_U77  ( .A1(_AES_ENC_us11_n1059 ), .A2(_AES_ENC_us11_n1114 ), .ZN(_AES_ENC_us11_n1012 ) );
NAND2_X2 _AES_ENC_us11_U76  ( .A1(_AES_ENC_us11_n1010 ), .A2(_AES_ENC_us11_n592 ), .ZN(_AES_ENC_us11_n1011 ) );
NAND2_X2 _AES_ENC_us11_U75  ( .A1(_AES_ENC_us11_n1012 ), .A2(_AES_ENC_us11_n1011 ), .ZN(_AES_ENC_us11_n1016 ) );
NAND4_X2 _AES_ENC_us11_U70  ( .A1(_AES_ENC_us11_n1020 ), .A2(_AES_ENC_us11_n1019 ), .A3(_AES_ENC_us11_n1018 ), .A4(_AES_ENC_us11_n1017 ), .ZN(_AES_ENC_us11_n1021 ) );
NAND2_X2 _AES_ENC_us11_U69  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n1021 ), .ZN(_AES_ENC_us11_n1042 ) );
NAND2_X2 _AES_ENC_us11_U68  ( .A1(_AES_ENC_us11_n1022 ), .A2(_AES_ENC_us11_n1093 ), .ZN(_AES_ENC_us11_n1039 ) );
NAND2_X2 _AES_ENC_us11_U67  ( .A1(_AES_ENC_us11_n1050 ), .A2(_AES_ENC_us11_n1023 ), .ZN(_AES_ENC_us11_n1038 ) );
NAND2_X2 _AES_ENC_us11_U66  ( .A1(_AES_ENC_us11_n1024 ), .A2(_AES_ENC_us11_n1071 ), .ZN(_AES_ENC_us11_n1037 ) );
AND2_X2 _AES_ENC_us11_U60  ( .A1(_AES_ENC_us11_n1030 ), .A2(_AES_ENC_us11_n602 ), .ZN(_AES_ENC_us11_n1078 ) );
NAND4_X2 _AES_ENC_us11_U56  ( .A1(_AES_ENC_us11_n1039 ), .A2(_AES_ENC_us11_n1038 ), .A3(_AES_ENC_us11_n1037 ), .A4(_AES_ENC_us11_n1036 ), .ZN(_AES_ENC_us11_n1040 ) );
NAND2_X2 _AES_ENC_us11_U55  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n1040 ), .ZN(_AES_ENC_us11_n1041 ) );
NAND4_X2 _AES_ENC_us11_U54  ( .A1(_AES_ENC_us11_n1044 ), .A2(_AES_ENC_us11_n1043 ), .A3(_AES_ENC_us11_n1042 ), .A4(_AES_ENC_us11_n1041 ), .ZN(_AES_ENC_sa11_sub[6] ) );
NAND2_X2 _AES_ENC_us11_U53  ( .A1(_AES_ENC_us11_n1072 ), .A2(_AES_ENC_us11_n1045 ), .ZN(_AES_ENC_us11_n1068 ) );
NAND2_X2 _AES_ENC_us11_U52  ( .A1(_AES_ENC_us11_n1046 ), .A2(_AES_ENC_us11_n582 ), .ZN(_AES_ENC_us11_n1067 ) );
NAND2_X2 _AES_ENC_us11_U51  ( .A1(_AES_ENC_us11_n1094 ), .A2(_AES_ENC_us11_n1047 ), .ZN(_AES_ENC_us11_n1066 ) );
NAND4_X2 _AES_ENC_us11_U40  ( .A1(_AES_ENC_us11_n1068 ), .A2(_AES_ENC_us11_n1067 ), .A3(_AES_ENC_us11_n1066 ), .A4(_AES_ENC_us11_n1065 ), .ZN(_AES_ENC_us11_n1069 ) );
NAND2_X2 _AES_ENC_us11_U39  ( .A1(_AES_ENC_us11_n1070 ), .A2(_AES_ENC_us11_n1069 ), .ZN(_AES_ENC_us11_n1135 ) );
NAND2_X2 _AES_ENC_us11_U38  ( .A1(_AES_ENC_us11_n1072 ), .A2(_AES_ENC_us11_n1071 ), .ZN(_AES_ENC_us11_n1088 ) );
NAND2_X2 _AES_ENC_us11_U37  ( .A1(_AES_ENC_us11_n1073 ), .A2(_AES_ENC_us11_n595 ), .ZN(_AES_ENC_us11_n1087 ) );
NAND4_X2 _AES_ENC_us11_U28  ( .A1(_AES_ENC_us11_n1088 ), .A2(_AES_ENC_us11_n1087 ), .A3(_AES_ENC_us11_n1086 ), .A4(_AES_ENC_us11_n1085 ), .ZN(_AES_ENC_us11_n1089 ) );
NAND2_X2 _AES_ENC_us11_U27  ( .A1(_AES_ENC_us11_n1090 ), .A2(_AES_ENC_us11_n1089 ), .ZN(_AES_ENC_us11_n1134 ) );
NAND2_X2 _AES_ENC_us11_U26  ( .A1(_AES_ENC_us11_n1091 ), .A2(_AES_ENC_us11_n1093 ), .ZN(_AES_ENC_us11_n1111 ) );
NAND2_X2 _AES_ENC_us11_U25  ( .A1(_AES_ENC_us11_n1092 ), .A2(_AES_ENC_us11_n1120 ), .ZN(_AES_ENC_us11_n1110 ) );
AND2_X2 _AES_ENC_us11_U22  ( .A1(_AES_ENC_us11_n1097 ), .A2(_AES_ENC_us11_n1096 ), .ZN(_AES_ENC_us11_n1098 ) );
NAND4_X2 _AES_ENC_us11_U14  ( .A1(_AES_ENC_us11_n1111 ), .A2(_AES_ENC_us11_n1110 ), .A3(_AES_ENC_us11_n1109 ), .A4(_AES_ENC_us11_n1108 ), .ZN(_AES_ENC_us11_n1112 ) );
NAND2_X2 _AES_ENC_us11_U13  ( .A1(_AES_ENC_us11_n1113 ), .A2(_AES_ENC_us11_n1112 ), .ZN(_AES_ENC_us11_n1133 ) );
NAND2_X2 _AES_ENC_us11_U12  ( .A1(_AES_ENC_us11_n1115 ), .A2(_AES_ENC_us11_n1114 ), .ZN(_AES_ENC_us11_n1129 ) );
OR2_X2 _AES_ENC_us11_U11  ( .A1(_AES_ENC_us11_n608 ), .A2(_AES_ENC_us11_n1116 ), .ZN(_AES_ENC_us11_n1128 ) );
NAND4_X2 _AES_ENC_us11_U3  ( .A1(_AES_ENC_us11_n1129 ), .A2(_AES_ENC_us11_n1128 ), .A3(_AES_ENC_us11_n1127 ), .A4(_AES_ENC_us11_n1126 ), .ZN(_AES_ENC_us11_n1130 ) );
NAND2_X2 _AES_ENC_us11_U2  ( .A1(_AES_ENC_us11_n1131 ), .A2(_AES_ENC_us11_n1130 ), .ZN(_AES_ENC_us11_n1132 ) );
NAND4_X2 _AES_ENC_us11_U1  ( .A1(_AES_ENC_us11_n1135 ), .A2(_AES_ENC_us11_n1134 ), .A3(_AES_ENC_us11_n1133 ), .A4(_AES_ENC_us11_n1132 ), .ZN(_AES_ENC_sa11_sub[7] ) );
INV_X4 _AES_ENC_us12_U575  ( .A(_AES_ENC_sa12[7]), .ZN(_AES_ENC_us12_n627 ));
INV_X4 _AES_ENC_us12_U574  ( .A(_AES_ENC_us12_n1114 ), .ZN(_AES_ENC_us12_n625 ) );
INV_X4 _AES_ENC_us12_U573  ( .A(_AES_ENC_sa12[4]), .ZN(_AES_ENC_us12_n624 ));
INV_X4 _AES_ENC_us12_U572  ( .A(_AES_ENC_us12_n1025 ), .ZN(_AES_ENC_us12_n622 ) );
INV_X4 _AES_ENC_us12_U571  ( .A(_AES_ENC_us12_n1120 ), .ZN(_AES_ENC_us12_n620 ) );
INV_X4 _AES_ENC_us12_U570  ( .A(_AES_ENC_us12_n1121 ), .ZN(_AES_ENC_us12_n619 ) );
INV_X4 _AES_ENC_us12_U569  ( .A(_AES_ENC_us12_n1048 ), .ZN(_AES_ENC_us12_n618 ) );
INV_X4 _AES_ENC_us12_U568  ( .A(_AES_ENC_us12_n974 ), .ZN(_AES_ENC_us12_n616 ) );
INV_X4 _AES_ENC_us12_U567  ( .A(_AES_ENC_us12_n794 ), .ZN(_AES_ENC_us12_n614 ) );
INV_X4 _AES_ENC_us12_U566  ( .A(_AES_ENC_sa12[2]), .ZN(_AES_ENC_us12_n611 ));
INV_X4 _AES_ENC_us12_U565  ( .A(_AES_ENC_us12_n800 ), .ZN(_AES_ENC_us12_n610 ) );
INV_X4 _AES_ENC_us12_U564  ( .A(_AES_ENC_us12_n925 ), .ZN(_AES_ENC_us12_n609 ) );
INV_X4 _AES_ENC_us12_U563  ( .A(_AES_ENC_us12_n779 ), .ZN(_AES_ENC_us12_n607 ) );
INV_X4 _AES_ENC_us12_U562  ( .A(_AES_ENC_us12_n1022 ), .ZN(_AES_ENC_us12_n603 ) );
INV_X4 _AES_ENC_us12_U561  ( .A(_AES_ENC_us12_n1102 ), .ZN(_AES_ENC_us12_n602 ) );
INV_X4 _AES_ENC_us12_U560  ( .A(_AES_ENC_us12_n929 ), .ZN(_AES_ENC_us12_n601 ) );
INV_X4 _AES_ENC_us12_U559  ( .A(_AES_ENC_us12_n1056 ), .ZN(_AES_ENC_us12_n600 ) );
INV_X4 _AES_ENC_us12_U558  ( .A(_AES_ENC_us12_n1054 ), .ZN(_AES_ENC_us12_n599 ) );
INV_X4 _AES_ENC_us12_U557  ( .A(_AES_ENC_us12_n881 ), .ZN(_AES_ENC_us12_n598 ) );
INV_X4 _AES_ENC_us12_U556  ( .A(_AES_ENC_us12_n926 ), .ZN(_AES_ENC_us12_n597 ) );
INV_X4 _AES_ENC_us12_U555  ( .A(_AES_ENC_us12_n977 ), .ZN(_AES_ENC_us12_n595 ) );
INV_X4 _AES_ENC_us12_U554  ( .A(_AES_ENC_us12_n1031 ), .ZN(_AES_ENC_us12_n594 ) );
INV_X4 _AES_ENC_us12_U553  ( .A(_AES_ENC_us12_n1103 ), .ZN(_AES_ENC_us12_n593 ) );
INV_X4 _AES_ENC_us12_U552  ( .A(_AES_ENC_us12_n1009 ), .ZN(_AES_ENC_us12_n592 ) );
INV_X4 _AES_ENC_us12_U551  ( .A(_AES_ENC_us12_n990 ), .ZN(_AES_ENC_us12_n591 ) );
INV_X4 _AES_ENC_us12_U550  ( .A(_AES_ENC_us12_n1058 ), .ZN(_AES_ENC_us12_n590 ) );
INV_X4 _AES_ENC_us12_U549  ( .A(_AES_ENC_us12_n1074 ), .ZN(_AES_ENC_us12_n589 ) );
INV_X4 _AES_ENC_us12_U548  ( .A(_AES_ENC_us12_n1053 ), .ZN(_AES_ENC_us12_n588 ) );
INV_X4 _AES_ENC_us12_U547  ( .A(_AES_ENC_us12_n826 ), .ZN(_AES_ENC_us12_n587 ) );
INV_X4 _AES_ENC_us12_U546  ( .A(_AES_ENC_us12_n992 ), .ZN(_AES_ENC_us12_n586 ) );
INV_X4 _AES_ENC_us12_U545  ( .A(_AES_ENC_us12_n821 ), .ZN(_AES_ENC_us12_n585 ) );
INV_X4 _AES_ENC_us12_U544  ( .A(_AES_ENC_us12_n910 ), .ZN(_AES_ENC_us12_n584 ) );
INV_X4 _AES_ENC_us12_U543  ( .A(_AES_ENC_us12_n906 ), .ZN(_AES_ENC_us12_n583 ) );
INV_X4 _AES_ENC_us12_U542  ( .A(_AES_ENC_us12_n880 ), .ZN(_AES_ENC_us12_n581 ) );
INV_X4 _AES_ENC_us12_U541  ( .A(_AES_ENC_us12_n1013 ), .ZN(_AES_ENC_us12_n580 ) );
INV_X4 _AES_ENC_us12_U540  ( .A(_AES_ENC_us12_n1092 ), .ZN(_AES_ENC_us12_n579 ) );
INV_X4 _AES_ENC_us12_U539  ( .A(_AES_ENC_us12_n824 ), .ZN(_AES_ENC_us12_n578 ) );
INV_X4 _AES_ENC_us12_U538  ( .A(_AES_ENC_us12_n1091 ), .ZN(_AES_ENC_us12_n577 ) );
INV_X4 _AES_ENC_us12_U537  ( .A(_AES_ENC_us12_n1080 ), .ZN(_AES_ENC_us12_n576 ) );
INV_X4 _AES_ENC_us12_U536  ( .A(_AES_ENC_us12_n959 ), .ZN(_AES_ENC_us12_n575 ) );
INV_X4 _AES_ENC_us12_U535  ( .A(_AES_ENC_sa12[0]), .ZN(_AES_ENC_us12_n574 ));
NOR2_X2 _AES_ENC_us12_U534  ( .A1(_AES_ENC_sa12[0]), .A2(_AES_ENC_sa12[6]),.ZN(_AES_ENC_us12_n1090 ) );
NOR2_X2 _AES_ENC_us12_U533  ( .A1(_AES_ENC_us12_n574 ), .A2(_AES_ENC_sa12[6]), .ZN(_AES_ENC_us12_n1070 ) );
NOR2_X2 _AES_ENC_us12_U532  ( .A1(_AES_ENC_sa12[4]), .A2(_AES_ENC_sa12[3]),.ZN(_AES_ENC_us12_n1025 ) );
INV_X4 _AES_ENC_us12_U531  ( .A(_AES_ENC_us12_n569 ), .ZN(_AES_ENC_us12_n572 ) );
NOR2_X2 _AES_ENC_us12_U530  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n765 ) );
NOR2_X2 _AES_ENC_us12_U529  ( .A1(_AES_ENC_sa12[4]), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n764 ) );
NOR2_X2 _AES_ENC_us12_U528  ( .A1(_AES_ENC_us12_n765 ), .A2(_AES_ENC_us12_n764 ), .ZN(_AES_ENC_us12_n766 ) );
NOR2_X2 _AES_ENC_us12_U527  ( .A1(_AES_ENC_us12_n766 ), .A2(_AES_ENC_us12_n575 ), .ZN(_AES_ENC_us12_n767 ) );
NOR3_X2 _AES_ENC_us12_U526  ( .A1(_AES_ENC_us12_n627 ), .A2(_AES_ENC_sa12[5]), .A3(_AES_ENC_us12_n704 ), .ZN(_AES_ENC_us12_n706 ));
NOR2_X2 _AES_ENC_us12_U525  ( .A1(_AES_ENC_us12_n1117 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n707 ) );
NOR2_X2 _AES_ENC_us12_U524  ( .A1(_AES_ENC_sa12[4]), .A2(_AES_ENC_us12_n579 ), .ZN(_AES_ENC_us12_n705 ) );
NOR3_X2 _AES_ENC_us12_U523  ( .A1(_AES_ENC_us12_n707 ), .A2(_AES_ENC_us12_n706 ), .A3(_AES_ENC_us12_n705 ), .ZN(_AES_ENC_us12_n713 ) );
INV_X4 _AES_ENC_us12_U522  ( .A(_AES_ENC_sa12[3]), .ZN(_AES_ENC_us12_n621 ));
NAND3_X2 _AES_ENC_us12_U521  ( .A1(_AES_ENC_us12_n652 ), .A2(_AES_ENC_us12_n626 ), .A3(_AES_ENC_sa12[7]), .ZN(_AES_ENC_us12_n653 ));
NOR2_X2 _AES_ENC_us12_U520  ( .A1(_AES_ENC_us12_n611 ), .A2(_AES_ENC_sa12[5]), .ZN(_AES_ENC_us12_n925 ) );
NOR2_X2 _AES_ENC_us12_U519  ( .A1(_AES_ENC_sa12[5]), .A2(_AES_ENC_sa12[2]),.ZN(_AES_ENC_us12_n974 ) );
INV_X4 _AES_ENC_us12_U518  ( .A(_AES_ENC_sa12[5]), .ZN(_AES_ENC_us12_n626 ));
NOR2_X2 _AES_ENC_us12_U517  ( .A1(_AES_ENC_us12_n611 ), .A2(_AES_ENC_sa12[7]), .ZN(_AES_ENC_us12_n779 ) );
NAND3_X2 _AES_ENC_us12_U516  ( .A1(_AES_ENC_us12_n679 ), .A2(_AES_ENC_us12_n678 ), .A3(_AES_ENC_us12_n677 ), .ZN(_AES_ENC_sa12_sub[0] ) );
NOR2_X2 _AES_ENC_us12_U515  ( .A1(_AES_ENC_us12_n626 ), .A2(_AES_ENC_sa12[2]), .ZN(_AES_ENC_us12_n1048 ) );
NOR4_X2 _AES_ENC_us12_U512  ( .A1(_AES_ENC_us12_n633 ), .A2(_AES_ENC_us12_n632 ), .A3(_AES_ENC_us12_n631 ), .A4(_AES_ENC_us12_n630 ), .ZN(_AES_ENC_us12_n634 ) );
NOR2_X2 _AES_ENC_us12_U510  ( .A1(_AES_ENC_us12_n629 ), .A2(_AES_ENC_us12_n628 ), .ZN(_AES_ENC_us12_n635 ) );
NAND3_X2 _AES_ENC_us12_U509  ( .A1(_AES_ENC_sa12[2]), .A2(_AES_ENC_sa12[7]), .A3(_AES_ENC_us12_n1059 ), .ZN(_AES_ENC_us12_n636 ) );
NOR2_X2 _AES_ENC_us12_U508  ( .A1(_AES_ENC_sa12[7]), .A2(_AES_ENC_sa12[2]),.ZN(_AES_ENC_us12_n794 ) );
NOR2_X2 _AES_ENC_us12_U507  ( .A1(_AES_ENC_sa12[4]), .A2(_AES_ENC_sa12[1]),.ZN(_AES_ENC_us12_n1102 ) );
NOR2_X2 _AES_ENC_us12_U506  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_sa12[3]), .ZN(_AES_ENC_us12_n1053 ) );
NOR2_X2 _AES_ENC_us12_U505  ( .A1(_AES_ENC_us12_n607 ), .A2(_AES_ENC_sa12[5]), .ZN(_AES_ENC_us12_n1024 ) );
NOR2_X2 _AES_ENC_us12_U504  ( .A1(_AES_ENC_us12_n625 ), .A2(_AES_ENC_sa12[2]), .ZN(_AES_ENC_us12_n1093 ) );
NOR2_X2 _AES_ENC_us12_U503  ( .A1(_AES_ENC_us12_n614 ), .A2(_AES_ENC_sa12[5]), .ZN(_AES_ENC_us12_n1094 ) );
NOR2_X2 _AES_ENC_us12_U502  ( .A1(_AES_ENC_us12_n624 ), .A2(_AES_ENC_sa12[3]), .ZN(_AES_ENC_us12_n931 ) );
INV_X4 _AES_ENC_us12_U501  ( .A(_AES_ENC_us12_n570 ), .ZN(_AES_ENC_us12_n573 ) );
NOR2_X2 _AES_ENC_us12_U500  ( .A1(_AES_ENC_us12_n1053 ), .A2(_AES_ENC_us12_n1095 ), .ZN(_AES_ENC_us12_n639 ) );
NOR3_X2 _AES_ENC_us12_U499  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n573 ), .A3(_AES_ENC_us12_n1074 ), .ZN(_AES_ENC_us12_n641 ) );
NOR2_X2 _AES_ENC_us12_U498  ( .A1(_AES_ENC_us12_n639 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n640 ) );
NOR2_X2 _AES_ENC_us12_U497  ( .A1(_AES_ENC_us12_n641 ), .A2(_AES_ENC_us12_n640 ), .ZN(_AES_ENC_us12_n646 ) );
NOR3_X2 _AES_ENC_us12_U496  ( .A1(_AES_ENC_us12_n995 ), .A2(_AES_ENC_us12_n586 ), .A3(_AES_ENC_us12_n994 ), .ZN(_AES_ENC_us12_n1002 ) );
NOR2_X2 _AES_ENC_us12_U495  ( .A1(_AES_ENC_us12_n909 ), .A2(_AES_ENC_us12_n908 ), .ZN(_AES_ENC_us12_n920 ) );
NOR2_X2 _AES_ENC_us12_U494  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n823 ) );
NOR2_X2 _AES_ENC_us12_U492  ( .A1(_AES_ENC_us12_n624 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n822 ) );
NOR2_X2 _AES_ENC_us12_U491  ( .A1(_AES_ENC_us12_n823 ), .A2(_AES_ENC_us12_n822 ), .ZN(_AES_ENC_us12_n825 ) );
NOR2_X2 _AES_ENC_us12_U490  ( .A1(_AES_ENC_sa12[1]), .A2(_AES_ENC_us12_n623 ), .ZN(_AES_ENC_us12_n913 ) );
NOR2_X2 _AES_ENC_us12_U489  ( .A1(_AES_ENC_us12_n913 ), .A2(_AES_ENC_us12_n1091 ), .ZN(_AES_ENC_us12_n914 ) );
NOR2_X2 _AES_ENC_us12_U488  ( .A1(_AES_ENC_us12_n826 ), .A2(_AES_ENC_us12_n572 ), .ZN(_AES_ENC_us12_n827 ) );
NOR3_X2 _AES_ENC_us12_U487  ( .A1(_AES_ENC_us12_n769 ), .A2(_AES_ENC_us12_n768 ), .A3(_AES_ENC_us12_n767 ), .ZN(_AES_ENC_us12_n775 ) );
NOR2_X2 _AES_ENC_us12_U486  ( .A1(_AES_ENC_us12_n1056 ), .A2(_AES_ENC_us12_n1053 ), .ZN(_AES_ENC_us12_n749 ) );
NOR2_X2 _AES_ENC_us12_U483  ( .A1(_AES_ENC_us12_n749 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n752 ) );
INV_X4 _AES_ENC_us12_U482  ( .A(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n596 ));
NOR2_X2 _AES_ENC_us12_U480  ( .A1(_AES_ENC_us12_n1054 ), .A2(_AES_ENC_us12_n1053 ), .ZN(_AES_ENC_us12_n1055 ) );
OR2_X4 _AES_ENC_us12_U479  ( .A1(_AES_ENC_us12_n1094 ), .A2(_AES_ENC_us12_n1093 ), .ZN(_AES_ENC_us12_n571 ) );
AND2_X2 _AES_ENC_us12_U478  ( .A1(_AES_ENC_us12_n571 ), .A2(_AES_ENC_us12_n1095 ), .ZN(_AES_ENC_us12_n1101 ) );
NOR2_X2 _AES_ENC_us12_U477  ( .A1(_AES_ENC_us12_n1074 ), .A2(_AES_ENC_us12_n931 ), .ZN(_AES_ENC_us12_n796 ) );
NOR2_X2 _AES_ENC_us12_U474  ( .A1(_AES_ENC_us12_n796 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n797 ) );
NOR2_X2 _AES_ENC_us12_U473  ( .A1(_AES_ENC_us12_n932 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n933 ) );
NOR2_X2 _AES_ENC_us12_U472  ( .A1(_AES_ENC_us12_n929 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n935 ) );
NOR2_X2 _AES_ENC_us12_U471  ( .A1(_AES_ENC_us12_n931 ), .A2(_AES_ENC_us12_n930 ), .ZN(_AES_ENC_us12_n934 ) );
NOR3_X2 _AES_ENC_us12_U470  ( .A1(_AES_ENC_us12_n935 ), .A2(_AES_ENC_us12_n934 ), .A3(_AES_ENC_us12_n933 ), .ZN(_AES_ENC_us12_n936 ) );
NOR2_X2 _AES_ENC_us12_U469  ( .A1(_AES_ENC_us12_n624 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n1075 ) );
NOR2_X2 _AES_ENC_us12_U468  ( .A1(_AES_ENC_us12_n572 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n949 ) );
NOR2_X2 _AES_ENC_us12_U467  ( .A1(_AES_ENC_us12_n1049 ), .A2(_AES_ENC_us12_n618 ), .ZN(_AES_ENC_us12_n1051 ) );
NOR2_X2 _AES_ENC_us12_U466  ( .A1(_AES_ENC_us12_n1051 ), .A2(_AES_ENC_us12_n1050 ), .ZN(_AES_ENC_us12_n1052 ) );
NOR2_X2 _AES_ENC_us12_U465  ( .A1(_AES_ENC_us12_n1052 ), .A2(_AES_ENC_us12_n592 ), .ZN(_AES_ENC_us12_n1064 ) );
NOR2_X2 _AES_ENC_us12_U464  ( .A1(_AES_ENC_sa12[1]), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n631 ) );
NOR2_X2 _AES_ENC_us12_U463  ( .A1(_AES_ENC_us12_n1025 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n980 ) );
NOR2_X2 _AES_ENC_us12_U462  ( .A1(_AES_ENC_us12_n1073 ), .A2(_AES_ENC_us12_n1094 ), .ZN(_AES_ENC_us12_n795 ) );
NOR2_X2 _AES_ENC_us12_U461  ( .A1(_AES_ENC_us12_n795 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n799 ) );
NOR2_X2 _AES_ENC_us12_U460  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n981 ) );
NOR2_X2 _AES_ENC_us12_U459  ( .A1(_AES_ENC_us12_n1102 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n643 ) );
NOR2_X2 _AES_ENC_us12_U458  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n621 ), .ZN(_AES_ENC_us12_n642 ) );
NOR2_X2 _AES_ENC_us12_U455  ( .A1(_AES_ENC_us12_n911 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n644 ) );
NOR4_X2 _AES_ENC_us12_U448  ( .A1(_AES_ENC_us12_n644 ), .A2(_AES_ENC_us12_n643 ), .A3(_AES_ENC_us12_n804 ), .A4(_AES_ENC_us12_n642 ), .ZN(_AES_ENC_us12_n645 ) );
NOR2_X2 _AES_ENC_us12_U447  ( .A1(_AES_ENC_us12_n1102 ), .A2(_AES_ENC_us12_n910 ), .ZN(_AES_ENC_us12_n932 ) );
NOR2_X2 _AES_ENC_us12_U442  ( .A1(_AES_ENC_us12_n1102 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n755 ) );
NOR2_X2 _AES_ENC_us12_U441  ( .A1(_AES_ENC_us12_n931 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n743 ) );
NOR2_X2 _AES_ENC_us12_U438  ( .A1(_AES_ENC_us12_n1072 ), .A2(_AES_ENC_us12_n1094 ), .ZN(_AES_ENC_us12_n930 ) );
NOR2_X2 _AES_ENC_us12_U435  ( .A1(_AES_ENC_us12_n1074 ), .A2(_AES_ENC_us12_n1025 ), .ZN(_AES_ENC_us12_n891 ) );
NOR2_X2 _AES_ENC_us12_U434  ( .A1(_AES_ENC_us12_n891 ), .A2(_AES_ENC_us12_n609 ), .ZN(_AES_ENC_us12_n894 ) );
NOR3_X2 _AES_ENC_us12_U433  ( .A1(_AES_ENC_us12_n623 ), .A2(_AES_ENC_sa12[1]), .A3(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n683 ));
INV_X4 _AES_ENC_us12_U428  ( .A(_AES_ENC_us12_n931 ), .ZN(_AES_ENC_us12_n623 ) );
NOR2_X2 _AES_ENC_us12_U427  ( .A1(_AES_ENC_us12_n996 ), .A2(_AES_ENC_us12_n931 ), .ZN(_AES_ENC_us12_n704 ) );
NOR2_X2 _AES_ENC_us12_U421  ( .A1(_AES_ENC_us12_n931 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n685 ) );
NOR2_X2 _AES_ENC_us12_U420  ( .A1(_AES_ENC_us12_n1029 ), .A2(_AES_ENC_us12_n1025 ), .ZN(_AES_ENC_us12_n1079 ) );
NOR3_X2 _AES_ENC_us12_U419  ( .A1(_AES_ENC_us12_n589 ), .A2(_AES_ENC_us12_n1025 ), .A3(_AES_ENC_us12_n616 ), .ZN(_AES_ENC_us12_n945 ) );
NOR2_X2 _AES_ENC_us12_U418  ( .A1(_AES_ENC_us12_n626 ), .A2(_AES_ENC_us12_n611 ), .ZN(_AES_ENC_us12_n800 ) );
NOR3_X2 _AES_ENC_us12_U417  ( .A1(_AES_ENC_us12_n590 ), .A2(_AES_ENC_us12_n627 ), .A3(_AES_ENC_us12_n611 ), .ZN(_AES_ENC_us12_n798 ) );
NOR3_X2 _AES_ENC_us12_U416  ( .A1(_AES_ENC_us12_n610 ), .A2(_AES_ENC_us12_n572 ), .A3(_AES_ENC_us12_n575 ), .ZN(_AES_ENC_us12_n962 ) );
NOR3_X2 _AES_ENC_us12_U415  ( .A1(_AES_ENC_us12_n959 ), .A2(_AES_ENC_us12_n572 ), .A3(_AES_ENC_us12_n609 ), .ZN(_AES_ENC_us12_n768 ) );
NOR3_X2 _AES_ENC_us12_U414  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n572 ), .A3(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n694 ) );
NOR3_X2 _AES_ENC_us12_U413  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n572 ), .A3(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n895 ) );
NOR3_X2 _AES_ENC_us12_U410  ( .A1(_AES_ENC_us12_n1008 ), .A2(_AES_ENC_us12_n1007 ), .A3(_AES_ENC_us12_n1006 ), .ZN(_AES_ENC_us12_n1018 ) );
NOR4_X2 _AES_ENC_us12_U409  ( .A1(_AES_ENC_us12_n806 ), .A2(_AES_ENC_us12_n805 ), .A3(_AES_ENC_us12_n804 ), .A4(_AES_ENC_us12_n803 ), .ZN(_AES_ENC_us12_n807 ) );
NOR3_X2 _AES_ENC_us12_U406  ( .A1(_AES_ENC_us12_n799 ), .A2(_AES_ENC_us12_n798 ), .A3(_AES_ENC_us12_n797 ), .ZN(_AES_ENC_us12_n808 ) );
NOR4_X2 _AES_ENC_us12_U405  ( .A1(_AES_ENC_us12_n843 ), .A2(_AES_ENC_us12_n842 ), .A3(_AES_ENC_us12_n841 ), .A4(_AES_ENC_us12_n840 ), .ZN(_AES_ENC_us12_n844 ) );
NOR3_X2 _AES_ENC_us12_U404  ( .A1(_AES_ENC_us12_n1101 ), .A2(_AES_ENC_us12_n1100 ), .A3(_AES_ENC_us12_n1099 ), .ZN(_AES_ENC_us12_n1109 ) );
NOR4_X2 _AES_ENC_us12_U403  ( .A1(_AES_ENC_us12_n711 ), .A2(_AES_ENC_us12_n710 ), .A3(_AES_ENC_us12_n709 ), .A4(_AES_ENC_us12_n708 ), .ZN(_AES_ENC_us12_n712 ) );
NOR4_X2 _AES_ENC_us12_U401  ( .A1(_AES_ENC_us12_n963 ), .A2(_AES_ENC_us12_n962 ), .A3(_AES_ENC_us12_n961 ), .A4(_AES_ENC_us12_n960 ), .ZN(_AES_ENC_us12_n964 ) );
NOR2_X2 _AES_ENC_us12_U400  ( .A1(_AES_ENC_us12_n669 ), .A2(_AES_ENC_us12_n668 ), .ZN(_AES_ENC_us12_n673 ) );
NOR4_X2 _AES_ENC_us12_U399  ( .A1(_AES_ENC_us12_n946 ), .A2(_AES_ENC_us12_n1046 ), .A3(_AES_ENC_us12_n671 ), .A4(_AES_ENC_us12_n670 ), .ZN(_AES_ENC_us12_n672 ) );
NOR3_X2 _AES_ENC_us12_U398  ( .A1(_AES_ENC_us12_n743 ), .A2(_AES_ENC_us12_n742 ), .A3(_AES_ENC_us12_n741 ), .ZN(_AES_ENC_us12_n744 ) );
NOR2_X2 _AES_ENC_us12_U397  ( .A1(_AES_ENC_us12_n697 ), .A2(_AES_ENC_us12_n658 ), .ZN(_AES_ENC_us12_n659 ) );
NOR2_X2 _AES_ENC_us12_U396  ( .A1(_AES_ENC_us12_n1078 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n1033 ) );
NOR2_X2 _AES_ENC_us12_U393  ( .A1(_AES_ENC_us12_n1031 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n1032 ) );
NOR3_X2 _AES_ENC_us12_U390  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n1025 ), .A3(_AES_ENC_us12_n1074 ), .ZN(_AES_ENC_us12_n1035 ) );
NOR4_X2 _AES_ENC_us12_U389  ( .A1(_AES_ENC_us12_n1035 ), .A2(_AES_ENC_us12_n1034 ), .A3(_AES_ENC_us12_n1033 ), .A4(_AES_ENC_us12_n1032 ), .ZN(_AES_ENC_us12_n1036 ) );
NOR2_X2 _AES_ENC_us12_U388  ( .A1(_AES_ENC_us12_n598 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n885 ) );
NOR2_X2 _AES_ENC_us12_U387  ( .A1(_AES_ENC_us12_n623 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n882 ) );
NOR2_X2 _AES_ENC_us12_U386  ( .A1(_AES_ENC_us12_n1053 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n884 ) );
NOR4_X2 _AES_ENC_us12_U385  ( .A1(_AES_ENC_us12_n885 ), .A2(_AES_ENC_us12_n884 ), .A3(_AES_ENC_us12_n883 ), .A4(_AES_ENC_us12_n882 ), .ZN(_AES_ENC_us12_n886 ) );
NOR2_X2 _AES_ENC_us12_U384  ( .A1(_AES_ENC_us12_n825 ), .A2(_AES_ENC_us12_n578 ), .ZN(_AES_ENC_us12_n830 ) );
NOR2_X2 _AES_ENC_us12_U383  ( .A1(_AES_ENC_us12_n827 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n829 ) );
NOR2_X2 _AES_ENC_us12_U382  ( .A1(_AES_ENC_us12_n572 ), .A2(_AES_ENC_us12_n579 ), .ZN(_AES_ENC_us12_n828 ) );
NOR4_X2 _AES_ENC_us12_U374  ( .A1(_AES_ENC_us12_n831 ), .A2(_AES_ENC_us12_n830 ), .A3(_AES_ENC_us12_n829 ), .A4(_AES_ENC_us12_n828 ), .ZN(_AES_ENC_us12_n832 ) );
NOR2_X2 _AES_ENC_us12_U373  ( .A1(_AES_ENC_us12_n606 ), .A2(_AES_ENC_us12_n582 ), .ZN(_AES_ENC_us12_n1104 ) );
NOR2_X2 _AES_ENC_us12_U372  ( .A1(_AES_ENC_us12_n1102 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n1106 ) );
NOR2_X2 _AES_ENC_us12_U370  ( .A1(_AES_ENC_us12_n1103 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n1105 ) );
NOR4_X2 _AES_ENC_us12_U369  ( .A1(_AES_ENC_us12_n1107 ), .A2(_AES_ENC_us12_n1106 ), .A3(_AES_ENC_us12_n1105 ), .A4(_AES_ENC_us12_n1104 ), .ZN(_AES_ENC_us12_n1108 ) );
NOR3_X2 _AES_ENC_us12_U368  ( .A1(_AES_ENC_us12_n959 ), .A2(_AES_ENC_us12_n621 ), .A3(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n963 ) );
NOR2_X2 _AES_ENC_us12_U367  ( .A1(_AES_ENC_us12_n626 ), .A2(_AES_ENC_us12_n627 ), .ZN(_AES_ENC_us12_n1114 ) );
INV_X4 _AES_ENC_us12_U366  ( .A(_AES_ENC_us12_n1024 ), .ZN(_AES_ENC_us12_n606 ) );
NOR3_X2 _AES_ENC_us12_U365  ( .A1(_AES_ENC_us12_n910 ), .A2(_AES_ENC_us12_n1059 ), .A3(_AES_ENC_us12_n611 ), .ZN(_AES_ENC_us12_n1115 ) );
INV_X4 _AES_ENC_us12_U364  ( .A(_AES_ENC_us12_n1094 ), .ZN(_AES_ENC_us12_n613 ) );
NOR2_X2 _AES_ENC_us12_U363  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n931 ), .ZN(_AES_ENC_us12_n1100 ) );
INV_X4 _AES_ENC_us12_U354  ( .A(_AES_ENC_us12_n1093 ), .ZN(_AES_ENC_us12_n617 ) );
NOR2_X2 _AES_ENC_us12_U353  ( .A1(_AES_ENC_us12_n569 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n929 ) );
NOR2_X2 _AES_ENC_us12_U352  ( .A1(_AES_ENC_us12_n620 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n926 ) );
NOR2_X2 _AES_ENC_us12_U351  ( .A1(_AES_ENC_us12_n572 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n1095 ) );
NOR2_X2 _AES_ENC_us12_U350  ( .A1(_AES_ENC_us12_n609 ), .A2(_AES_ENC_us12_n627 ), .ZN(_AES_ENC_us12_n1010 ) );
NOR2_X2 _AES_ENC_us12_U349  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n1103 ) );
NOR2_X2 _AES_ENC_us12_U348  ( .A1(_AES_ENC_us12_n622 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n1059 ) );
NOR2_X2 _AES_ENC_us12_U347  ( .A1(_AES_ENC_sa12[1]), .A2(_AES_ENC_us12_n1120 ), .ZN(_AES_ENC_us12_n1022 ) );
NOR2_X2 _AES_ENC_us12_U346  ( .A1(_AES_ENC_us12_n619 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n911 ) );
NOR2_X2 _AES_ENC_us12_U345  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_us12_n1025 ), .ZN(_AES_ENC_us12_n826 ) );
NOR2_X2 _AES_ENC_us12_U338  ( .A1(_AES_ENC_us12_n626 ), .A2(_AES_ENC_us12_n607 ), .ZN(_AES_ENC_us12_n1072 ) );
NOR2_X2 _AES_ENC_us12_U335  ( .A1(_AES_ENC_us12_n627 ), .A2(_AES_ENC_us12_n616 ), .ZN(_AES_ENC_us12_n956 ) );
NOR2_X2 _AES_ENC_us12_U329  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_us12_n624 ), .ZN(_AES_ENC_us12_n1121 ) );
NOR2_X2 _AES_ENC_us12_U328  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_us12_n624 ), .ZN(_AES_ENC_us12_n1058 ) );
NOR2_X2 _AES_ENC_us12_U327  ( .A1(_AES_ENC_us12_n625 ), .A2(_AES_ENC_us12_n611 ), .ZN(_AES_ENC_us12_n1073 ) );
NOR2_X2 _AES_ENC_us12_U325  ( .A1(_AES_ENC_sa12[1]), .A2(_AES_ENC_us12_n1025 ), .ZN(_AES_ENC_us12_n1054 ) );
NOR2_X2 _AES_ENC_us12_U324  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_us12_n931 ), .ZN(_AES_ENC_us12_n1029 ) );
NOR2_X2 _AES_ENC_us12_U319  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n1056 ) );
NOR2_X2 _AES_ENC_us12_U318  ( .A1(_AES_ENC_us12_n614 ), .A2(_AES_ENC_us12_n626 ), .ZN(_AES_ENC_us12_n1050 ) );
NOR2_X2 _AES_ENC_us12_U317  ( .A1(_AES_ENC_us12_n1121 ), .A2(_AES_ENC_us12_n1025 ), .ZN(_AES_ENC_us12_n1120 ) );
NOR2_X2 _AES_ENC_us12_U316  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_us12_n572 ), .ZN(_AES_ENC_us12_n1074 ) );
NOR2_X2 _AES_ENC_us12_U315  ( .A1(_AES_ENC_us12_n1058 ), .A2(_AES_ENC_us12_n1054 ), .ZN(_AES_ENC_us12_n878 ) );
NOR2_X2 _AES_ENC_us12_U314  ( .A1(_AES_ENC_us12_n878 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n879 ) );
NOR2_X2 _AES_ENC_us12_U312  ( .A1(_AES_ENC_us12_n880 ), .A2(_AES_ENC_us12_n879 ), .ZN(_AES_ENC_us12_n887 ) );
NOR2_X2 _AES_ENC_us12_U311  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n588 ), .ZN(_AES_ENC_us12_n957 ) );
NOR2_X2 _AES_ENC_us12_U310  ( .A1(_AES_ENC_us12_n958 ), .A2(_AES_ENC_us12_n957 ), .ZN(_AES_ENC_us12_n965 ) );
NOR3_X2 _AES_ENC_us12_U309  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n1091 ), .A3(_AES_ENC_us12_n1022 ), .ZN(_AES_ENC_us12_n720 ) );
NOR3_X2 _AES_ENC_us12_U303  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n1054 ), .A3(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n719 ) );
NOR2_X2 _AES_ENC_us12_U302  ( .A1(_AES_ENC_us12_n720 ), .A2(_AES_ENC_us12_n719 ), .ZN(_AES_ENC_us12_n726 ) );
NOR2_X2 _AES_ENC_us12_U300  ( .A1(_AES_ENC_us12_n614 ), .A2(_AES_ENC_us12_n591 ), .ZN(_AES_ENC_us12_n865 ) );
NOR2_X2 _AES_ENC_us12_U299  ( .A1(_AES_ENC_us12_n1059 ), .A2(_AES_ENC_us12_n1058 ), .ZN(_AES_ENC_us12_n1060 ) );
NOR2_X2 _AES_ENC_us12_U298  ( .A1(_AES_ENC_us12_n1095 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n668 ) );
NOR2_X2 _AES_ENC_us12_U297  ( .A1(_AES_ENC_us12_n911 ), .A2(_AES_ENC_us12_n910 ), .ZN(_AES_ENC_us12_n912 ) );
NOR2_X2 _AES_ENC_us12_U296  ( .A1(_AES_ENC_us12_n912 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n916 ) );
NOR2_X2 _AES_ENC_us12_U295  ( .A1(_AES_ENC_us12_n826 ), .A2(_AES_ENC_us12_n573 ), .ZN(_AES_ENC_us12_n750 ) );
NOR2_X2 _AES_ENC_us12_U294  ( .A1(_AES_ENC_us12_n750 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n751 ) );
NOR2_X2 _AES_ENC_us12_U293  ( .A1(_AES_ENC_us12_n907 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n908 ) );
NOR2_X2 _AES_ENC_us12_U292  ( .A1(_AES_ENC_us12_n990 ), .A2(_AES_ENC_us12_n926 ), .ZN(_AES_ENC_us12_n780 ) );
NOR2_X2 _AES_ENC_us12_U291  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n584 ), .ZN(_AES_ENC_us12_n838 ) );
NOR2_X2 _AES_ENC_us12_U290  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n602 ), .ZN(_AES_ENC_us12_n837 ) );
NOR2_X2 _AES_ENC_us12_U284  ( .A1(_AES_ENC_us12_n838 ), .A2(_AES_ENC_us12_n837 ), .ZN(_AES_ENC_us12_n845 ) );
NOR2_X2 _AES_ENC_us12_U283  ( .A1(_AES_ENC_us12_n1022 ), .A2(_AES_ENC_us12_n1058 ), .ZN(_AES_ENC_us12_n740 ) );
NOR2_X2 _AES_ENC_us12_U282  ( .A1(_AES_ENC_us12_n740 ), .A2(_AES_ENC_us12_n616 ), .ZN(_AES_ENC_us12_n742 ) );
NOR2_X2 _AES_ENC_us12_U281  ( .A1(_AES_ENC_us12_n1098 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n1099 ) );
NOR2_X2 _AES_ENC_us12_U280  ( .A1(_AES_ENC_us12_n1120 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n993 ) );
NOR2_X2 _AES_ENC_us12_U279  ( .A1(_AES_ENC_us12_n993 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n994 ) );
NOR2_X2 _AES_ENC_us12_U273  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n620 ), .ZN(_AES_ENC_us12_n1026 ) );
NOR2_X2 _AES_ENC_us12_U272  ( .A1(_AES_ENC_us12_n573 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n1027 ) );
NOR2_X2 _AES_ENC_us12_U271  ( .A1(_AES_ENC_us12_n1027 ), .A2(_AES_ENC_us12_n1026 ), .ZN(_AES_ENC_us12_n1028 ) );
NOR2_X2 _AES_ENC_us12_U270  ( .A1(_AES_ENC_us12_n1029 ), .A2(_AES_ENC_us12_n1028 ), .ZN(_AES_ENC_us12_n1034 ) );
NOR4_X2 _AES_ENC_us12_U269  ( .A1(_AES_ENC_us12_n757 ), .A2(_AES_ENC_us12_n756 ), .A3(_AES_ENC_us12_n755 ), .A4(_AES_ENC_us12_n754 ), .ZN(_AES_ENC_us12_n758 ) );
NOR2_X2 _AES_ENC_us12_U268  ( .A1(_AES_ENC_us12_n752 ), .A2(_AES_ENC_us12_n751 ), .ZN(_AES_ENC_us12_n759 ) );
NOR2_X2 _AES_ENC_us12_U267  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n1071 ), .ZN(_AES_ENC_us12_n669 ) );
NOR2_X2 _AES_ENC_us12_U263  ( .A1(_AES_ENC_us12_n1056 ), .A2(_AES_ENC_us12_n990 ), .ZN(_AES_ENC_us12_n991 ) );
NOR2_X2 _AES_ENC_us12_U262  ( .A1(_AES_ENC_us12_n991 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n995 ) );
NOR2_X2 _AES_ENC_us12_U258  ( .A1(_AES_ENC_us12_n607 ), .A2(_AES_ENC_us12_n590 ), .ZN(_AES_ENC_us12_n1008 ) );
NOR2_X2 _AES_ENC_us12_U255  ( .A1(_AES_ENC_us12_n839 ), .A2(_AES_ENC_us12_n582 ), .ZN(_AES_ENC_us12_n693 ) );
NOR2_X2 _AES_ENC_us12_U254  ( .A1(_AES_ENC_us12_n606 ), .A2(_AES_ENC_us12_n906 ), .ZN(_AES_ENC_us12_n741 ) );
NOR2_X2 _AES_ENC_us12_U253  ( .A1(_AES_ENC_us12_n1054 ), .A2(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n763 ) );
NOR2_X2 _AES_ENC_us12_U252  ( .A1(_AES_ENC_us12_n763 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n769 ) );
NOR2_X2 _AES_ENC_us12_U251  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n577 ), .ZN(_AES_ENC_us12_n1007 ) );
NOR2_X2 _AES_ENC_us12_U250  ( .A1(_AES_ENC_us12_n609 ), .A2(_AES_ENC_us12_n580 ), .ZN(_AES_ENC_us12_n1123 ) );
NOR2_X2 _AES_ENC_us12_U243  ( .A1(_AES_ENC_us12_n609 ), .A2(_AES_ENC_us12_n590 ), .ZN(_AES_ENC_us12_n710 ) );
INV_X4 _AES_ENC_us12_U242  ( .A(_AES_ENC_us12_n1029 ), .ZN(_AES_ENC_us12_n582 ) );
NOR2_X2 _AES_ENC_us12_U241  ( .A1(_AES_ENC_us12_n616 ), .A2(_AES_ENC_us12_n597 ), .ZN(_AES_ENC_us12_n883 ) );
NOR2_X2 _AES_ENC_us12_U240  ( .A1(_AES_ENC_us12_n593 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n1125 ) );
NOR2_X2 _AES_ENC_us12_U239  ( .A1(_AES_ENC_us12_n990 ), .A2(_AES_ENC_us12_n929 ), .ZN(_AES_ENC_us12_n892 ) );
NOR2_X2 _AES_ENC_us12_U238  ( .A1(_AES_ENC_us12_n892 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n893 ) );
NOR2_X2 _AES_ENC_us12_U237  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n602 ), .ZN(_AES_ENC_us12_n950 ) );
NOR2_X2 _AES_ENC_us12_U236  ( .A1(_AES_ENC_us12_n1079 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n1082 ) );
NOR2_X2 _AES_ENC_us12_U235  ( .A1(_AES_ENC_us12_n910 ), .A2(_AES_ENC_us12_n1056 ), .ZN(_AES_ENC_us12_n941 ) );
NOR2_X2 _AES_ENC_us12_U234  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n1077 ), .ZN(_AES_ENC_us12_n841 ) );
NOR2_X2 _AES_ENC_us12_U229  ( .A1(_AES_ENC_us12_n623 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n630 ) );
NOR2_X2 _AES_ENC_us12_U228  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n602 ), .ZN(_AES_ENC_us12_n806 ) );
NOR2_X2 _AES_ENC_us12_U227  ( .A1(_AES_ENC_us12_n623 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n948 ) );
NOR2_X2 _AES_ENC_us12_U226  ( .A1(_AES_ENC_us12_n606 ), .A2(_AES_ENC_us12_n589 ), .ZN(_AES_ENC_us12_n997 ) );
NOR2_X2 _AES_ENC_us12_U225  ( .A1(_AES_ENC_us12_n1121 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n1122 ) );
NOR2_X2 _AES_ENC_us12_U223  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n1023 ), .ZN(_AES_ENC_us12_n756 ) );
NOR2_X2 _AES_ENC_us12_U222  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n602 ), .ZN(_AES_ENC_us12_n870 ) );
NOR2_X2 _AES_ENC_us12_U221  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n569 ), .ZN(_AES_ENC_us12_n947 ) );
NOR2_X2 _AES_ENC_us12_U217  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n1077 ), .ZN(_AES_ENC_us12_n1084 ) );
NOR2_X2 _AES_ENC_us12_U213  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n855 ), .ZN(_AES_ENC_us12_n709 ) );
NOR2_X2 _AES_ENC_us12_U212  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n589 ), .ZN(_AES_ENC_us12_n868 ) );
NOR2_X2 _AES_ENC_us12_U211  ( .A1(_AES_ENC_us12_n1120 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n1124 ) );
NOR2_X2 _AES_ENC_us12_U210  ( .A1(_AES_ENC_us12_n1120 ), .A2(_AES_ENC_us12_n839 ), .ZN(_AES_ENC_us12_n842 ) );
NOR2_X2 _AES_ENC_us12_U209  ( .A1(_AES_ENC_us12_n1120 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n696 ) );
NOR2_X2 _AES_ENC_us12_U208  ( .A1(_AES_ENC_us12_n1074 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n1076 ) );
NOR2_X2 _AES_ENC_us12_U207  ( .A1(_AES_ENC_us12_n1074 ), .A2(_AES_ENC_us12_n620 ), .ZN(_AES_ENC_us12_n781 ) );
NOR3_X2 _AES_ENC_us12_U201  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n1056 ), .A3(_AES_ENC_us12_n990 ), .ZN(_AES_ENC_us12_n979 ) );
NOR3_X2 _AES_ENC_us12_U200  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n1058 ), .A3(_AES_ENC_us12_n1059 ), .ZN(_AES_ENC_us12_n854 ) );
NOR2_X2 _AES_ENC_us12_U199  ( .A1(_AES_ENC_us12_n996 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n869 ) );
NOR2_X2 _AES_ENC_us12_U198  ( .A1(_AES_ENC_us12_n1056 ), .A2(_AES_ENC_us12_n1074 ), .ZN(_AES_ENC_us12_n1057 ) );
NOR3_X2 _AES_ENC_us12_U197  ( .A1(_AES_ENC_us12_n607 ), .A2(_AES_ENC_us12_n1120 ), .A3(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n978 ) );
NOR2_X2 _AES_ENC_us12_U196  ( .A1(_AES_ENC_us12_n996 ), .A2(_AES_ENC_us12_n911 ), .ZN(_AES_ENC_us12_n1116 ) );
NOR2_X2 _AES_ENC_us12_U195  ( .A1(_AES_ENC_us12_n1074 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n754 ) );
NOR2_X2 _AES_ENC_us12_U194  ( .A1(_AES_ENC_us12_n926 ), .A2(_AES_ENC_us12_n1103 ), .ZN(_AES_ENC_us12_n977 ) );
NOR2_X2 _AES_ENC_us12_U187  ( .A1(_AES_ENC_us12_n839 ), .A2(_AES_ENC_us12_n824 ), .ZN(_AES_ENC_us12_n1092 ) );
NOR2_X2 _AES_ENC_us12_U186  ( .A1(_AES_ENC_us12_n573 ), .A2(_AES_ENC_us12_n1074 ), .ZN(_AES_ENC_us12_n684 ) );
NOR2_X2 _AES_ENC_us12_U185  ( .A1(_AES_ENC_us12_n826 ), .A2(_AES_ENC_us12_n1059 ), .ZN(_AES_ENC_us12_n907 ) );
NOR3_X2 _AES_ENC_us12_U184  ( .A1(_AES_ENC_us12_n625 ), .A2(_AES_ENC_us12_n1115 ), .A3(_AES_ENC_us12_n585 ), .ZN(_AES_ENC_us12_n831 ) );
NOR3_X2 _AES_ENC_us12_U183  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n1056 ), .A3(_AES_ENC_us12_n990 ), .ZN(_AES_ENC_us12_n896 ) );
NOR3_X2 _AES_ENC_us12_U182  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n573 ), .A3(_AES_ENC_us12_n1013 ), .ZN(_AES_ENC_us12_n670 ) );
NOR3_X2 _AES_ENC_us12_U181  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n1091 ), .A3(_AES_ENC_us12_n1022 ), .ZN(_AES_ENC_us12_n843 ) );
NOR2_X2 _AES_ENC_us12_U180  ( .A1(_AES_ENC_us12_n1029 ), .A2(_AES_ENC_us12_n1095 ), .ZN(_AES_ENC_us12_n735 ) );
NOR2_X2 _AES_ENC_us12_U174  ( .A1(_AES_ENC_us12_n1100 ), .A2(_AES_ENC_us12_n854 ), .ZN(_AES_ENC_us12_n860 ) );
NOR4_X2 _AES_ENC_us12_U173  ( .A1(_AES_ENC_us12_n1125 ), .A2(_AES_ENC_us12_n1124 ), .A3(_AES_ENC_us12_n1123 ), .A4(_AES_ENC_us12_n1122 ), .ZN(_AES_ENC_us12_n1126 ) );
NOR4_X2 _AES_ENC_us12_U172  ( .A1(_AES_ENC_us12_n1084 ), .A2(_AES_ENC_us12_n1083 ), .A3(_AES_ENC_us12_n1082 ), .A4(_AES_ENC_us12_n1081 ), .ZN(_AES_ENC_us12_n1085 ) );
NOR2_X2 _AES_ENC_us12_U171  ( .A1(_AES_ENC_us12_n1076 ), .A2(_AES_ENC_us12_n1075 ), .ZN(_AES_ENC_us12_n1086 ) );
NAND3_X2 _AES_ENC_us12_U170  ( .A1(_AES_ENC_us12_n569 ), .A2(_AES_ENC_us12_n582 ), .A3(_AES_ENC_us12_n681 ), .ZN(_AES_ENC_us12_n691 ) );
NOR2_X2 _AES_ENC_us12_U169  ( .A1(_AES_ENC_us12_n683 ), .A2(_AES_ENC_us12_n682 ), .ZN(_AES_ENC_us12_n690 ) );
NOR3_X2 _AES_ENC_us12_U168  ( .A1(_AES_ENC_us12_n695 ), .A2(_AES_ENC_us12_n694 ), .A3(_AES_ENC_us12_n693 ), .ZN(_AES_ENC_us12_n700 ) );
NOR4_X2 _AES_ENC_us12_U162  ( .A1(_AES_ENC_us12_n983 ), .A2(_AES_ENC_us12_n698 ), .A3(_AES_ENC_us12_n697 ), .A4(_AES_ENC_us12_n696 ), .ZN(_AES_ENC_us12_n699 ) );
NOR2_X2 _AES_ENC_us12_U161  ( .A1(_AES_ENC_us12_n946 ), .A2(_AES_ENC_us12_n945 ), .ZN(_AES_ENC_us12_n952 ) );
NOR4_X2 _AES_ENC_us12_U160  ( .A1(_AES_ENC_us12_n950 ), .A2(_AES_ENC_us12_n949 ), .A3(_AES_ENC_us12_n948 ), .A4(_AES_ENC_us12_n947 ), .ZN(_AES_ENC_us12_n951 ) );
NOR4_X2 _AES_ENC_us12_U159  ( .A1(_AES_ENC_us12_n983 ), .A2(_AES_ENC_us12_n982 ), .A3(_AES_ENC_us12_n981 ), .A4(_AES_ENC_us12_n980 ), .ZN(_AES_ENC_us12_n984 ) );
NOR2_X2 _AES_ENC_us12_U158  ( .A1(_AES_ENC_us12_n979 ), .A2(_AES_ENC_us12_n978 ), .ZN(_AES_ENC_us12_n985 ) );
NOR4_X2 _AES_ENC_us12_U157  ( .A1(_AES_ENC_us12_n896 ), .A2(_AES_ENC_us12_n895 ), .A3(_AES_ENC_us12_n894 ), .A4(_AES_ENC_us12_n893 ), .ZN(_AES_ENC_us12_n897 ) );
NOR2_X2 _AES_ENC_us12_U156  ( .A1(_AES_ENC_us12_n866 ), .A2(_AES_ENC_us12_n865 ), .ZN(_AES_ENC_us12_n872 ) );
NOR4_X2 _AES_ENC_us12_U155  ( .A1(_AES_ENC_us12_n870 ), .A2(_AES_ENC_us12_n869 ), .A3(_AES_ENC_us12_n868 ), .A4(_AES_ENC_us12_n867 ), .ZN(_AES_ENC_us12_n871 ) );
NOR3_X2 _AES_ENC_us12_U154  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n1054 ), .A3(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n961 ) );
NOR3_X2 _AES_ENC_us12_U153  ( .A1(_AES_ENC_us12_n620 ), .A2(_AES_ENC_us12_n1074 ), .A3(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n671 ) );
NOR2_X2 _AES_ENC_us12_U152  ( .A1(_AES_ENC_us12_n1057 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n1062 ) );
NOR2_X2 _AES_ENC_us12_U143  ( .A1(_AES_ENC_us12_n1055 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n1063 ) );
NOR2_X2 _AES_ENC_us12_U142  ( .A1(_AES_ENC_us12_n1060 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n1061 ) );
NOR4_X2 _AES_ENC_us12_U141  ( .A1(_AES_ENC_us12_n1064 ), .A2(_AES_ENC_us12_n1063 ), .A3(_AES_ENC_us12_n1062 ), .A4(_AES_ENC_us12_n1061 ), .ZN(_AES_ENC_us12_n1065 ) );
NOR3_X2 _AES_ENC_us12_U140  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n1120 ), .A3(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n918 ) );
NOR3_X2 _AES_ENC_us12_U132  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n573 ), .A3(_AES_ENC_us12_n1013 ), .ZN(_AES_ENC_us12_n917 ) );
NOR2_X2 _AES_ENC_us12_U131  ( .A1(_AES_ENC_us12_n914 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n915 ) );
NOR4_X2 _AES_ENC_us12_U130  ( .A1(_AES_ENC_us12_n918 ), .A2(_AES_ENC_us12_n917 ), .A3(_AES_ENC_us12_n916 ), .A4(_AES_ENC_us12_n915 ), .ZN(_AES_ENC_us12_n919 ) );
NOR2_X2 _AES_ENC_us12_U129  ( .A1(_AES_ENC_us12_n616 ), .A2(_AES_ENC_us12_n580 ), .ZN(_AES_ENC_us12_n771 ) );
NOR2_X2 _AES_ENC_us12_U128  ( .A1(_AES_ENC_us12_n1103 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n772 ) );
NOR2_X2 _AES_ENC_us12_U127  ( .A1(_AES_ENC_us12_n610 ), .A2(_AES_ENC_us12_n599 ), .ZN(_AES_ENC_us12_n773 ) );
NOR4_X2 _AES_ENC_us12_U126  ( .A1(_AES_ENC_us12_n773 ), .A2(_AES_ENC_us12_n772 ), .A3(_AES_ENC_us12_n771 ), .A4(_AES_ENC_us12_n770 ), .ZN(_AES_ENC_us12_n774 ) );
NOR2_X2 _AES_ENC_us12_U121  ( .A1(_AES_ENC_us12_n735 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n687 ) );
NOR2_X2 _AES_ENC_us12_U120  ( .A1(_AES_ENC_us12_n684 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n688 ) );
NOR2_X2 _AES_ENC_us12_U119  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n600 ), .ZN(_AES_ENC_us12_n686 ) );
NOR4_X2 _AES_ENC_us12_U118  ( .A1(_AES_ENC_us12_n688 ), .A2(_AES_ENC_us12_n687 ), .A3(_AES_ENC_us12_n686 ), .A4(_AES_ENC_us12_n685 ), .ZN(_AES_ENC_us12_n689 ) );
NOR2_X2 _AES_ENC_us12_U117  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n595 ), .ZN(_AES_ENC_us12_n858 ) );
NOR2_X2 _AES_ENC_us12_U116  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n855 ), .ZN(_AES_ENC_us12_n857 ) );
NOR2_X2 _AES_ENC_us12_U115  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n587 ), .ZN(_AES_ENC_us12_n856 ) );
NOR4_X2 _AES_ENC_us12_U106  ( .A1(_AES_ENC_us12_n858 ), .A2(_AES_ENC_us12_n857 ), .A3(_AES_ENC_us12_n856 ), .A4(_AES_ENC_us12_n958 ), .ZN(_AES_ENC_us12_n859 ) );
NOR2_X2 _AES_ENC_us12_U105  ( .A1(_AES_ENC_us12_n780 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n784 ) );
NOR2_X2 _AES_ENC_us12_U104  ( .A1(_AES_ENC_us12_n1117 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n782 ) );
NOR2_X2 _AES_ENC_us12_U103  ( .A1(_AES_ENC_us12_n781 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n783 ) );
NOR4_X2 _AES_ENC_us12_U102  ( .A1(_AES_ENC_us12_n880 ), .A2(_AES_ENC_us12_n784 ), .A3(_AES_ENC_us12_n783 ), .A4(_AES_ENC_us12_n782 ), .ZN(_AES_ENC_us12_n785 ) );
NOR2_X2 _AES_ENC_us12_U101  ( .A1(_AES_ENC_us12_n583 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n814 ) );
NOR2_X2 _AES_ENC_us12_U100  ( .A1(_AES_ENC_us12_n907 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n813 ) );
NOR3_X2 _AES_ENC_us12_U95  ( .A1(_AES_ENC_us12_n606 ), .A2(_AES_ENC_us12_n1058 ), .A3(_AES_ENC_us12_n1059 ), .ZN(_AES_ENC_us12_n815 ) );
NOR4_X2 _AES_ENC_us12_U94  ( .A1(_AES_ENC_us12_n815 ), .A2(_AES_ENC_us12_n814 ), .A3(_AES_ENC_us12_n813 ), .A4(_AES_ENC_us12_n812 ), .ZN(_AES_ENC_us12_n816 ) );
NOR2_X2 _AES_ENC_us12_U93  ( .A1(_AES_ENC_us12_n617 ), .A2(_AES_ENC_us12_n569 ), .ZN(_AES_ENC_us12_n721 ) );
NOR2_X2 _AES_ENC_us12_U92  ( .A1(_AES_ENC_us12_n1031 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n723 ) );
NOR2_X2 _AES_ENC_us12_U91  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n1096 ), .ZN(_AES_ENC_us12_n722 ) );
NOR4_X2 _AES_ENC_us12_U90  ( .A1(_AES_ENC_us12_n724 ), .A2(_AES_ENC_us12_n723 ), .A3(_AES_ENC_us12_n722 ), .A4(_AES_ENC_us12_n721 ), .ZN(_AES_ENC_us12_n725 ) );
NOR2_X2 _AES_ENC_us12_U89  ( .A1(_AES_ENC_us12_n911 ), .A2(_AES_ENC_us12_n990 ), .ZN(_AES_ENC_us12_n1009 ) );
NOR2_X2 _AES_ENC_us12_U88  ( .A1(_AES_ENC_us12_n1013 ), .A2(_AES_ENC_us12_n573 ), .ZN(_AES_ENC_us12_n1014 ) );
NOR2_X2 _AES_ENC_us12_U87  ( .A1(_AES_ENC_us12_n1014 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n1015 ) );
NOR4_X2 _AES_ENC_us12_U86  ( .A1(_AES_ENC_us12_n1016 ), .A2(_AES_ENC_us12_n1015 ), .A3(_AES_ENC_us12_n1119 ), .A4(_AES_ENC_us12_n1046 ), .ZN(_AES_ENC_us12_n1017 ) );
NOR2_X2 _AES_ENC_us12_U81  ( .A1(_AES_ENC_us12_n996 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n998 ) );
NOR2_X2 _AES_ENC_us12_U80  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n577 ), .ZN(_AES_ENC_us12_n1000 ) );
NOR2_X2 _AES_ENC_us12_U79  ( .A1(_AES_ENC_us12_n616 ), .A2(_AES_ENC_us12_n1096 ), .ZN(_AES_ENC_us12_n999 ) );
NOR4_X2 _AES_ENC_us12_U78  ( .A1(_AES_ENC_us12_n1000 ), .A2(_AES_ENC_us12_n999 ), .A3(_AES_ENC_us12_n998 ), .A4(_AES_ENC_us12_n997 ), .ZN(_AES_ENC_us12_n1001 ) );
NOR2_X2 _AES_ENC_us12_U74  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n1096 ), .ZN(_AES_ENC_us12_n697 ) );
NOR2_X2 _AES_ENC_us12_U73  ( .A1(_AES_ENC_us12_n620 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n958 ) );
NOR2_X2 _AES_ENC_us12_U72  ( .A1(_AES_ENC_us12_n911 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n983 ) );
NOR2_X2 _AES_ENC_us12_U71  ( .A1(_AES_ENC_us12_n1054 ), .A2(_AES_ENC_us12_n1103 ), .ZN(_AES_ENC_us12_n1031 ) );
INV_X4 _AES_ENC_us12_U65  ( .A(_AES_ENC_us12_n1050 ), .ZN(_AES_ENC_us12_n612 ) );
INV_X4 _AES_ENC_us12_U64  ( .A(_AES_ENC_us12_n1072 ), .ZN(_AES_ENC_us12_n605 ) );
INV_X4 _AES_ENC_us12_U63  ( .A(_AES_ENC_us12_n1073 ), .ZN(_AES_ENC_us12_n604 ) );
NOR2_X2 _AES_ENC_us12_U62  ( .A1(_AES_ENC_us12_n582 ), .A2(_AES_ENC_us12_n613 ), .ZN(_AES_ENC_us12_n880 ) );
NOR3_X2 _AES_ENC_us12_U61  ( .A1(_AES_ENC_us12_n826 ), .A2(_AES_ENC_us12_n1121 ), .A3(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n946 ) );
INV_X4 _AES_ENC_us12_U59  ( .A(_AES_ENC_us12_n1010 ), .ZN(_AES_ENC_us12_n608 ) );
NOR3_X2 _AES_ENC_us12_U58  ( .A1(_AES_ENC_us12_n573 ), .A2(_AES_ENC_us12_n1029 ), .A3(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n1119 ) );
INV_X4 _AES_ENC_us12_U57  ( .A(_AES_ENC_us12_n956 ), .ZN(_AES_ENC_us12_n615 ) );
NOR2_X2 _AES_ENC_us12_U50  ( .A1(_AES_ENC_us12_n623 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n1013 ) );
NOR2_X2 _AES_ENC_us12_U49  ( .A1(_AES_ENC_us12_n620 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n910 ) );
NOR2_X2 _AES_ENC_us12_U48  ( .A1(_AES_ENC_us12_n569 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n1091 ) );
NOR2_X2 _AES_ENC_us12_U47  ( .A1(_AES_ENC_us12_n622 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n990 ) );
NOR2_X2 _AES_ENC_us12_U46  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_us12_n1121 ), .ZN(_AES_ENC_us12_n996 ) );
NOR2_X2 _AES_ENC_us12_U45  ( .A1(_AES_ENC_us12_n610 ), .A2(_AES_ENC_us12_n600 ), .ZN(_AES_ENC_us12_n628 ) );
NOR2_X2 _AES_ENC_us12_U44  ( .A1(_AES_ENC_us12_n576 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n866 ) );
NOR2_X2 _AES_ENC_us12_U43  ( .A1(_AES_ENC_us12_n603 ), .A2(_AES_ENC_us12_n610 ), .ZN(_AES_ENC_us12_n1006 ) );
NOR2_X2 _AES_ENC_us12_U42  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n1117 ), .ZN(_AES_ENC_us12_n1118 ) );
NOR2_X2 _AES_ENC_us12_U41  ( .A1(_AES_ENC_us12_n1119 ), .A2(_AES_ENC_us12_n1118 ), .ZN(_AES_ENC_us12_n1127 ) );
NOR2_X2 _AES_ENC_us12_U36  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n906 ), .ZN(_AES_ENC_us12_n909 ) );
NOR2_X2 _AES_ENC_us12_U35  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n594 ), .ZN(_AES_ENC_us12_n629 ) );
NOR2_X2 _AES_ENC_us12_U34  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n597 ), .ZN(_AES_ENC_us12_n658 ) );
NOR2_X2 _AES_ENC_us12_U33  ( .A1(_AES_ENC_us12_n1116 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n695 ) );
NOR2_X2 _AES_ENC_us12_U32  ( .A1(_AES_ENC_us12_n1078 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n1083 ) );
NOR2_X2 _AES_ENC_us12_U31  ( .A1(_AES_ENC_us12_n941 ), .A2(_AES_ENC_us12_n608 ), .ZN(_AES_ENC_us12_n724 ) );
NOR2_X2 _AES_ENC_us12_U30  ( .A1(_AES_ENC_us12_n598 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n1107 ) );
NOR2_X2 _AES_ENC_us12_U29  ( .A1(_AES_ENC_us12_n576 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n840 ) );
NOR2_X2 _AES_ENC_us12_U24  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n593 ), .ZN(_AES_ENC_us12_n633 ) );
NOR2_X2 _AES_ENC_us12_U23  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n1080 ), .ZN(_AES_ENC_us12_n1081 ) );
NOR2_X2 _AES_ENC_us12_U21  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n1045 ), .ZN(_AES_ENC_us12_n812 ) );
NOR2_X2 _AES_ENC_us12_U20  ( .A1(_AES_ENC_us12_n1009 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n960 ) );
NOR2_X2 _AES_ENC_us12_U19  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n601 ), .ZN(_AES_ENC_us12_n982 ) );
NOR2_X2 _AES_ENC_us12_U18  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n594 ), .ZN(_AES_ENC_us12_n757 ) );
NOR2_X2 _AES_ENC_us12_U17  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n590 ), .ZN(_AES_ENC_us12_n698 ) );
NOR2_X2 _AES_ENC_us12_U16  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n619 ), .ZN(_AES_ENC_us12_n708 ) );
NOR2_X2 _AES_ENC_us12_U15  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n582 ), .ZN(_AES_ENC_us12_n770 ) );
NOR2_X2 _AES_ENC_us12_U10  ( .A1(_AES_ENC_us12_n619 ), .A2(_AES_ENC_us12_n604 ), .ZN(_AES_ENC_us12_n803 ) );
NOR2_X2 _AES_ENC_us12_U9  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n881 ), .ZN(_AES_ENC_us12_n711 ) );
NOR2_X2 _AES_ENC_us12_U8  ( .A1(_AES_ENC_us12_n615 ), .A2(_AES_ENC_us12_n582 ), .ZN(_AES_ENC_us12_n867 ) );
NOR2_X2 _AES_ENC_us12_U7  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n599 ), .ZN(_AES_ENC_us12_n804 ) );
NOR2_X2 _AES_ENC_us12_U6  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n620 ), .ZN(_AES_ENC_us12_n1046 ) );
OR2_X4 _AES_ENC_us12_U5  ( .A1(_AES_ENC_us12_n624 ), .A2(_AES_ENC_sa12[1]),.ZN(_AES_ENC_us12_n570 ) );
OR2_X4 _AES_ENC_us12_U4  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_sa12[4]),.ZN(_AES_ENC_us12_n569 ) );
NAND2_X2 _AES_ENC_us12_U514  ( .A1(_AES_ENC_us12_n1121 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n1030 ) );
AND2_X2 _AES_ENC_us12_U513  ( .A1(_AES_ENC_us12_n597 ), .A2(_AES_ENC_us12_n1030 ), .ZN(_AES_ENC_us12_n1049 ) );
NAND2_X2 _AES_ENC_us12_U511  ( .A1(_AES_ENC_us12_n1049 ), .A2(_AES_ENC_us12_n794 ), .ZN(_AES_ENC_us12_n637 ) );
AND2_X2 _AES_ENC_us12_U493  ( .A1(_AES_ENC_us12_n779 ), .A2(_AES_ENC_us12_n996 ), .ZN(_AES_ENC_us12_n632 ) );
NAND4_X2 _AES_ENC_us12_U485  ( .A1(_AES_ENC_us12_n637 ), .A2(_AES_ENC_us12_n636 ), .A3(_AES_ENC_us12_n635 ), .A4(_AES_ENC_us12_n634 ), .ZN(_AES_ENC_us12_n638 ) );
NAND2_X2 _AES_ENC_us12_U484  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n638 ), .ZN(_AES_ENC_us12_n679 ) );
NAND2_X2 _AES_ENC_us12_U481  ( .A1(_AES_ENC_us12_n1094 ), .A2(_AES_ENC_us12_n591 ), .ZN(_AES_ENC_us12_n648 ) );
NAND2_X2 _AES_ENC_us12_U476  ( .A1(_AES_ENC_us12_n601 ), .A2(_AES_ENC_us12_n590 ), .ZN(_AES_ENC_us12_n762 ) );
NAND2_X2 _AES_ENC_us12_U475  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n762 ), .ZN(_AES_ENC_us12_n647 ) );
NAND4_X2 _AES_ENC_us12_U457  ( .A1(_AES_ENC_us12_n648 ), .A2(_AES_ENC_us12_n647 ), .A3(_AES_ENC_us12_n646 ), .A4(_AES_ENC_us12_n645 ), .ZN(_AES_ENC_us12_n649 ) );
NAND2_X2 _AES_ENC_us12_U456  ( .A1(_AES_ENC_sa12[0]), .A2(_AES_ENC_us12_n649 ), .ZN(_AES_ENC_us12_n665 ) );
NAND2_X2 _AES_ENC_us12_U454  ( .A1(_AES_ENC_us12_n596 ), .A2(_AES_ENC_us12_n623 ), .ZN(_AES_ENC_us12_n855 ) );
NAND2_X2 _AES_ENC_us12_U453  ( .A1(_AES_ENC_us12_n587 ), .A2(_AES_ENC_us12_n855 ), .ZN(_AES_ENC_us12_n821 ) );
NAND2_X2 _AES_ENC_us12_U452  ( .A1(_AES_ENC_us12_n1093 ), .A2(_AES_ENC_us12_n821 ), .ZN(_AES_ENC_us12_n662 ) );
NAND2_X2 _AES_ENC_us12_U451  ( .A1(_AES_ENC_us12_n619 ), .A2(_AES_ENC_us12_n589 ), .ZN(_AES_ENC_us12_n650 ) );
NAND2_X2 _AES_ENC_us12_U450  ( .A1(_AES_ENC_us12_n956 ), .A2(_AES_ENC_us12_n650 ), .ZN(_AES_ENC_us12_n661 ) );
NAND2_X2 _AES_ENC_us12_U449  ( .A1(_AES_ENC_us12_n626 ), .A2(_AES_ENC_us12_n627 ), .ZN(_AES_ENC_us12_n839 ) );
OR2_X2 _AES_ENC_us12_U446  ( .A1(_AES_ENC_us12_n839 ), .A2(_AES_ENC_us12_n932 ), .ZN(_AES_ENC_us12_n656 ) );
NAND2_X2 _AES_ENC_us12_U445  ( .A1(_AES_ENC_us12_n621 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n1096 ) );
NAND2_X2 _AES_ENC_us12_U444  ( .A1(_AES_ENC_us12_n1030 ), .A2(_AES_ENC_us12_n1096 ), .ZN(_AES_ENC_us12_n651 ) );
NAND2_X2 _AES_ENC_us12_U443  ( .A1(_AES_ENC_us12_n1114 ), .A2(_AES_ENC_us12_n651 ), .ZN(_AES_ENC_us12_n655 ) );
OR3_X2 _AES_ENC_us12_U440  ( .A1(_AES_ENC_us12_n1079 ), .A2(_AES_ENC_sa12[7]), .A3(_AES_ENC_us12_n626 ), .ZN(_AES_ENC_us12_n654 ));
NAND2_X2 _AES_ENC_us12_U439  ( .A1(_AES_ENC_us12_n593 ), .A2(_AES_ENC_us12_n601 ), .ZN(_AES_ENC_us12_n652 ) );
NAND4_X2 _AES_ENC_us12_U437  ( .A1(_AES_ENC_us12_n656 ), .A2(_AES_ENC_us12_n655 ), .A3(_AES_ENC_us12_n654 ), .A4(_AES_ENC_us12_n653 ), .ZN(_AES_ENC_us12_n657 ) );
NAND2_X2 _AES_ENC_us12_U436  ( .A1(_AES_ENC_sa12[2]), .A2(_AES_ENC_us12_n657 ), .ZN(_AES_ENC_us12_n660 ) );
NAND4_X2 _AES_ENC_us12_U432  ( .A1(_AES_ENC_us12_n662 ), .A2(_AES_ENC_us12_n661 ), .A3(_AES_ENC_us12_n660 ), .A4(_AES_ENC_us12_n659 ), .ZN(_AES_ENC_us12_n663 ) );
NAND2_X2 _AES_ENC_us12_U431  ( .A1(_AES_ENC_us12_n663 ), .A2(_AES_ENC_us12_n574 ), .ZN(_AES_ENC_us12_n664 ) );
NAND2_X2 _AES_ENC_us12_U430  ( .A1(_AES_ENC_us12_n665 ), .A2(_AES_ENC_us12_n664 ), .ZN(_AES_ENC_us12_n666 ) );
NAND2_X2 _AES_ENC_us12_U429  ( .A1(_AES_ENC_sa12[6]), .A2(_AES_ENC_us12_n666 ), .ZN(_AES_ENC_us12_n678 ) );
NAND2_X2 _AES_ENC_us12_U426  ( .A1(_AES_ENC_us12_n735 ), .A2(_AES_ENC_us12_n1093 ), .ZN(_AES_ENC_us12_n675 ) );
NAND2_X2 _AES_ENC_us12_U425  ( .A1(_AES_ENC_us12_n588 ), .A2(_AES_ENC_us12_n597 ), .ZN(_AES_ENC_us12_n1045 ) );
OR2_X2 _AES_ENC_us12_U424  ( .A1(_AES_ENC_us12_n1045 ), .A2(_AES_ENC_us12_n605 ), .ZN(_AES_ENC_us12_n674 ) );
NAND2_X2 _AES_ENC_us12_U423  ( .A1(_AES_ENC_sa12[1]), .A2(_AES_ENC_us12_n620 ), .ZN(_AES_ENC_us12_n667 ) );
NAND2_X2 _AES_ENC_us12_U422  ( .A1(_AES_ENC_us12_n619 ), .A2(_AES_ENC_us12_n667 ), .ZN(_AES_ENC_us12_n1071 ) );
NAND4_X2 _AES_ENC_us12_U412  ( .A1(_AES_ENC_us12_n675 ), .A2(_AES_ENC_us12_n674 ), .A3(_AES_ENC_us12_n673 ), .A4(_AES_ENC_us12_n672 ), .ZN(_AES_ENC_us12_n676 ) );
NAND2_X2 _AES_ENC_us12_U411  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n676 ), .ZN(_AES_ENC_us12_n677 ) );
NAND2_X2 _AES_ENC_us12_U408  ( .A1(_AES_ENC_us12_n800 ), .A2(_AES_ENC_us12_n1022 ), .ZN(_AES_ENC_us12_n680 ) );
NAND2_X2 _AES_ENC_us12_U407  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n680 ), .ZN(_AES_ENC_us12_n681 ) );
AND2_X2 _AES_ENC_us12_U402  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n684 ), .ZN(_AES_ENC_us12_n682 ) );
NAND4_X2 _AES_ENC_us12_U395  ( .A1(_AES_ENC_us12_n691 ), .A2(_AES_ENC_us12_n581 ), .A3(_AES_ENC_us12_n690 ), .A4(_AES_ENC_us12_n689 ), .ZN(_AES_ENC_us12_n692 ) );
NAND2_X2 _AES_ENC_us12_U394  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n692 ), .ZN(_AES_ENC_us12_n733 ) );
NAND2_X2 _AES_ENC_us12_U392  ( .A1(_AES_ENC_us12_n977 ), .A2(_AES_ENC_us12_n1050 ), .ZN(_AES_ENC_us12_n702 ) );
NAND2_X2 _AES_ENC_us12_U391  ( .A1(_AES_ENC_us12_n1093 ), .A2(_AES_ENC_us12_n1045 ), .ZN(_AES_ENC_us12_n701 ) );
NAND4_X2 _AES_ENC_us12_U381  ( .A1(_AES_ENC_us12_n702 ), .A2(_AES_ENC_us12_n701 ), .A3(_AES_ENC_us12_n700 ), .A4(_AES_ENC_us12_n699 ), .ZN(_AES_ENC_us12_n703 ) );
NAND2_X2 _AES_ENC_us12_U380  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n703 ), .ZN(_AES_ENC_us12_n732 ) );
AND2_X2 _AES_ENC_us12_U379  ( .A1(_AES_ENC_sa12[0]), .A2(_AES_ENC_sa12[6]),.ZN(_AES_ENC_us12_n1113 ) );
NAND2_X2 _AES_ENC_us12_U378  ( .A1(_AES_ENC_us12_n601 ), .A2(_AES_ENC_us12_n1030 ), .ZN(_AES_ENC_us12_n881 ) );
NAND2_X2 _AES_ENC_us12_U377  ( .A1(_AES_ENC_us12_n1093 ), .A2(_AES_ENC_us12_n881 ), .ZN(_AES_ENC_us12_n715 ) );
NAND2_X2 _AES_ENC_us12_U376  ( .A1(_AES_ENC_us12_n1010 ), .A2(_AES_ENC_us12_n600 ), .ZN(_AES_ENC_us12_n714 ) );
NAND2_X2 _AES_ENC_us12_U375  ( .A1(_AES_ENC_us12_n855 ), .A2(_AES_ENC_us12_n588 ), .ZN(_AES_ENC_us12_n1117 ) );
XNOR2_X2 _AES_ENC_us12_U371  ( .A(_AES_ENC_us12_n611 ), .B(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n824 ) );
NAND4_X2 _AES_ENC_us12_U362  ( .A1(_AES_ENC_us12_n715 ), .A2(_AES_ENC_us12_n714 ), .A3(_AES_ENC_us12_n713 ), .A4(_AES_ENC_us12_n712 ), .ZN(_AES_ENC_us12_n716 ) );
NAND2_X2 _AES_ENC_us12_U361  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n716 ), .ZN(_AES_ENC_us12_n731 ) );
AND2_X2 _AES_ENC_us12_U360  ( .A1(_AES_ENC_sa12[6]), .A2(_AES_ENC_us12_n574 ), .ZN(_AES_ENC_us12_n1131 ) );
NAND2_X2 _AES_ENC_us12_U359  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n717 ) );
NAND2_X2 _AES_ENC_us12_U358  ( .A1(_AES_ENC_us12_n1029 ), .A2(_AES_ENC_us12_n717 ), .ZN(_AES_ENC_us12_n728 ) );
NAND2_X2 _AES_ENC_us12_U357  ( .A1(_AES_ENC_sa12[1]), .A2(_AES_ENC_us12_n624 ), .ZN(_AES_ENC_us12_n1097 ) );
NAND2_X2 _AES_ENC_us12_U356  ( .A1(_AES_ENC_us12_n603 ), .A2(_AES_ENC_us12_n1097 ), .ZN(_AES_ENC_us12_n718 ) );
NAND2_X2 _AES_ENC_us12_U355  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n718 ), .ZN(_AES_ENC_us12_n727 ) );
NAND4_X2 _AES_ENC_us12_U344  ( .A1(_AES_ENC_us12_n728 ), .A2(_AES_ENC_us12_n727 ), .A3(_AES_ENC_us12_n726 ), .A4(_AES_ENC_us12_n725 ), .ZN(_AES_ENC_us12_n729 ) );
NAND2_X2 _AES_ENC_us12_U343  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n729 ), .ZN(_AES_ENC_us12_n730 ) );
NAND4_X2 _AES_ENC_us12_U342  ( .A1(_AES_ENC_us12_n733 ), .A2(_AES_ENC_us12_n732 ), .A3(_AES_ENC_us12_n731 ), .A4(_AES_ENC_us12_n730 ), .ZN(_AES_ENC_sa12_sub[1] ) );
NAND2_X2 _AES_ENC_us12_U341  ( .A1(_AES_ENC_sa12[7]), .A2(_AES_ENC_us12_n611 ), .ZN(_AES_ENC_us12_n734 ) );
NAND2_X2 _AES_ENC_us12_U340  ( .A1(_AES_ENC_us12_n734 ), .A2(_AES_ENC_us12_n607 ), .ZN(_AES_ENC_us12_n738 ) );
OR4_X2 _AES_ENC_us12_U339  ( .A1(_AES_ENC_us12_n738 ), .A2(_AES_ENC_us12_n626 ), .A3(_AES_ENC_us12_n826 ), .A4(_AES_ENC_us12_n1121 ), .ZN(_AES_ENC_us12_n746 ) );
NAND2_X2 _AES_ENC_us12_U337  ( .A1(_AES_ENC_us12_n1100 ), .A2(_AES_ENC_us12_n587 ), .ZN(_AES_ENC_us12_n992 ) );
OR2_X2 _AES_ENC_us12_U336  ( .A1(_AES_ENC_us12_n610 ), .A2(_AES_ENC_us12_n735 ), .ZN(_AES_ENC_us12_n737 ) );
NAND2_X2 _AES_ENC_us12_U334  ( .A1(_AES_ENC_us12_n619 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n753 ) );
NAND2_X2 _AES_ENC_us12_U333  ( .A1(_AES_ENC_us12_n582 ), .A2(_AES_ENC_us12_n753 ), .ZN(_AES_ENC_us12_n1080 ) );
NAND2_X2 _AES_ENC_us12_U332  ( .A1(_AES_ENC_us12_n1048 ), .A2(_AES_ENC_us12_n576 ), .ZN(_AES_ENC_us12_n736 ) );
NAND2_X2 _AES_ENC_us12_U331  ( .A1(_AES_ENC_us12_n737 ), .A2(_AES_ENC_us12_n736 ), .ZN(_AES_ENC_us12_n739 ) );
NAND2_X2 _AES_ENC_us12_U330  ( .A1(_AES_ENC_us12_n739 ), .A2(_AES_ENC_us12_n738 ), .ZN(_AES_ENC_us12_n745 ) );
NAND2_X2 _AES_ENC_us12_U326  ( .A1(_AES_ENC_us12_n1096 ), .A2(_AES_ENC_us12_n590 ), .ZN(_AES_ENC_us12_n906 ) );
NAND4_X2 _AES_ENC_us12_U323  ( .A1(_AES_ENC_us12_n746 ), .A2(_AES_ENC_us12_n992 ), .A3(_AES_ENC_us12_n745 ), .A4(_AES_ENC_us12_n744 ), .ZN(_AES_ENC_us12_n747 ) );
NAND2_X2 _AES_ENC_us12_U322  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n747 ), .ZN(_AES_ENC_us12_n793 ) );
NAND2_X2 _AES_ENC_us12_U321  ( .A1(_AES_ENC_us12_n584 ), .A2(_AES_ENC_us12_n855 ), .ZN(_AES_ENC_us12_n748 ) );
NAND2_X2 _AES_ENC_us12_U320  ( .A1(_AES_ENC_us12_n956 ), .A2(_AES_ENC_us12_n748 ), .ZN(_AES_ENC_us12_n760 ) );
NAND2_X2 _AES_ENC_us12_U313  ( .A1(_AES_ENC_us12_n590 ), .A2(_AES_ENC_us12_n753 ), .ZN(_AES_ENC_us12_n1023 ) );
NAND4_X2 _AES_ENC_us12_U308  ( .A1(_AES_ENC_us12_n760 ), .A2(_AES_ENC_us12_n992 ), .A3(_AES_ENC_us12_n759 ), .A4(_AES_ENC_us12_n758 ), .ZN(_AES_ENC_us12_n761 ) );
NAND2_X2 _AES_ENC_us12_U307  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n761 ), .ZN(_AES_ENC_us12_n792 ) );
NAND2_X2 _AES_ENC_us12_U306  ( .A1(_AES_ENC_us12_n584 ), .A2(_AES_ENC_us12_n603 ), .ZN(_AES_ENC_us12_n989 ) );
NAND2_X2 _AES_ENC_us12_U305  ( .A1(_AES_ENC_us12_n1050 ), .A2(_AES_ENC_us12_n989 ), .ZN(_AES_ENC_us12_n777 ) );
NAND2_X2 _AES_ENC_us12_U304  ( .A1(_AES_ENC_us12_n1093 ), .A2(_AES_ENC_us12_n762 ), .ZN(_AES_ENC_us12_n776 ) );
XNOR2_X2 _AES_ENC_us12_U301  ( .A(_AES_ENC_sa12[7]), .B(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n959 ) );
NAND4_X2 _AES_ENC_us12_U289  ( .A1(_AES_ENC_us12_n777 ), .A2(_AES_ENC_us12_n776 ), .A3(_AES_ENC_us12_n775 ), .A4(_AES_ENC_us12_n774 ), .ZN(_AES_ENC_us12_n778 ) );
NAND2_X2 _AES_ENC_us12_U288  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n778 ), .ZN(_AES_ENC_us12_n791 ) );
NAND2_X2 _AES_ENC_us12_U287  ( .A1(_AES_ENC_us12_n1056 ), .A2(_AES_ENC_us12_n1050 ), .ZN(_AES_ENC_us12_n788 ) );
NAND2_X2 _AES_ENC_us12_U286  ( .A1(_AES_ENC_us12_n1091 ), .A2(_AES_ENC_us12_n779 ), .ZN(_AES_ENC_us12_n787 ) );
NAND2_X2 _AES_ENC_us12_U285  ( .A1(_AES_ENC_us12_n956 ), .A2(_AES_ENC_sa12[1]), .ZN(_AES_ENC_us12_n786 ) );
NAND4_X2 _AES_ENC_us12_U278  ( .A1(_AES_ENC_us12_n788 ), .A2(_AES_ENC_us12_n787 ), .A3(_AES_ENC_us12_n786 ), .A4(_AES_ENC_us12_n785 ), .ZN(_AES_ENC_us12_n789 ) );
NAND2_X2 _AES_ENC_us12_U277  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n789 ), .ZN(_AES_ENC_us12_n790 ) );
NAND4_X2 _AES_ENC_us12_U276  ( .A1(_AES_ENC_us12_n793 ), .A2(_AES_ENC_us12_n792 ), .A3(_AES_ENC_us12_n791 ), .A4(_AES_ENC_us12_n790 ), .ZN(_AES_ENC_sa12_sub[2] ) );
NAND2_X2 _AES_ENC_us12_U275  ( .A1(_AES_ENC_us12_n1059 ), .A2(_AES_ENC_us12_n794 ), .ZN(_AES_ENC_us12_n810 ) );
NAND2_X2 _AES_ENC_us12_U274  ( .A1(_AES_ENC_us12_n1049 ), .A2(_AES_ENC_us12_n956 ), .ZN(_AES_ENC_us12_n809 ) );
OR2_X2 _AES_ENC_us12_U266  ( .A1(_AES_ENC_us12_n1096 ), .A2(_AES_ENC_us12_n606 ), .ZN(_AES_ENC_us12_n802 ) );
NAND2_X2 _AES_ENC_us12_U265  ( .A1(_AES_ENC_us12_n1053 ), .A2(_AES_ENC_us12_n800 ), .ZN(_AES_ENC_us12_n801 ) );
NAND2_X2 _AES_ENC_us12_U264  ( .A1(_AES_ENC_us12_n802 ), .A2(_AES_ENC_us12_n801 ), .ZN(_AES_ENC_us12_n805 ) );
NAND4_X2 _AES_ENC_us12_U261  ( .A1(_AES_ENC_us12_n810 ), .A2(_AES_ENC_us12_n809 ), .A3(_AES_ENC_us12_n808 ), .A4(_AES_ENC_us12_n807 ), .ZN(_AES_ENC_us12_n811 ) );
NAND2_X2 _AES_ENC_us12_U260  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n811 ), .ZN(_AES_ENC_us12_n852 ) );
OR2_X2 _AES_ENC_us12_U259  ( .A1(_AES_ENC_us12_n1023 ), .A2(_AES_ENC_us12_n617 ), .ZN(_AES_ENC_us12_n819 ) );
OR2_X2 _AES_ENC_us12_U257  ( .A1(_AES_ENC_us12_n570 ), .A2(_AES_ENC_us12_n930 ), .ZN(_AES_ENC_us12_n818 ) );
NAND2_X2 _AES_ENC_us12_U256  ( .A1(_AES_ENC_us12_n1013 ), .A2(_AES_ENC_us12_n1094 ), .ZN(_AES_ENC_us12_n817 ) );
NAND4_X2 _AES_ENC_us12_U249  ( .A1(_AES_ENC_us12_n819 ), .A2(_AES_ENC_us12_n818 ), .A3(_AES_ENC_us12_n817 ), .A4(_AES_ENC_us12_n816 ), .ZN(_AES_ENC_us12_n820 ) );
NAND2_X2 _AES_ENC_us12_U248  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n820 ), .ZN(_AES_ENC_us12_n851 ) );
NAND2_X2 _AES_ENC_us12_U247  ( .A1(_AES_ENC_us12_n956 ), .A2(_AES_ENC_us12_n1080 ), .ZN(_AES_ENC_us12_n835 ) );
NAND2_X2 _AES_ENC_us12_U246  ( .A1(_AES_ENC_us12_n570 ), .A2(_AES_ENC_us12_n1030 ), .ZN(_AES_ENC_us12_n1047 ) );
OR2_X2 _AES_ENC_us12_U245  ( .A1(_AES_ENC_us12_n1047 ), .A2(_AES_ENC_us12_n612 ), .ZN(_AES_ENC_us12_n834 ) );
NAND2_X2 _AES_ENC_us12_U244  ( .A1(_AES_ENC_us12_n1072 ), .A2(_AES_ENC_us12_n589 ), .ZN(_AES_ENC_us12_n833 ) );
NAND4_X2 _AES_ENC_us12_U233  ( .A1(_AES_ENC_us12_n835 ), .A2(_AES_ENC_us12_n834 ), .A3(_AES_ENC_us12_n833 ), .A4(_AES_ENC_us12_n832 ), .ZN(_AES_ENC_us12_n836 ) );
NAND2_X2 _AES_ENC_us12_U232  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n836 ), .ZN(_AES_ENC_us12_n850 ) );
NAND2_X2 _AES_ENC_us12_U231  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n623 ), .ZN(_AES_ENC_us12_n847 ) );
NAND2_X2 _AES_ENC_us12_U230  ( .A1(_AES_ENC_us12_n1050 ), .A2(_AES_ENC_us12_n1071 ), .ZN(_AES_ENC_us12_n846 ) );
OR2_X2 _AES_ENC_us12_U224  ( .A1(_AES_ENC_us12_n1053 ), .A2(_AES_ENC_us12_n911 ), .ZN(_AES_ENC_us12_n1077 ) );
NAND4_X2 _AES_ENC_us12_U220  ( .A1(_AES_ENC_us12_n847 ), .A2(_AES_ENC_us12_n846 ), .A3(_AES_ENC_us12_n845 ), .A4(_AES_ENC_us12_n844 ), .ZN(_AES_ENC_us12_n848 ) );
NAND2_X2 _AES_ENC_us12_U219  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n848 ), .ZN(_AES_ENC_us12_n849 ) );
NAND4_X2 _AES_ENC_us12_U218  ( .A1(_AES_ENC_us12_n852 ), .A2(_AES_ENC_us12_n851 ), .A3(_AES_ENC_us12_n850 ), .A4(_AES_ENC_us12_n849 ), .ZN(_AES_ENC_sa12_sub[3] ) );
NAND2_X2 _AES_ENC_us12_U216  ( .A1(_AES_ENC_us12_n1009 ), .A2(_AES_ENC_us12_n1072 ), .ZN(_AES_ENC_us12_n862 ) );
NAND2_X2 _AES_ENC_us12_U215  ( .A1(_AES_ENC_us12_n603 ), .A2(_AES_ENC_us12_n577 ), .ZN(_AES_ENC_us12_n853 ) );
NAND2_X2 _AES_ENC_us12_U214  ( .A1(_AES_ENC_us12_n1050 ), .A2(_AES_ENC_us12_n853 ), .ZN(_AES_ENC_us12_n861 ) );
NAND4_X2 _AES_ENC_us12_U206  ( .A1(_AES_ENC_us12_n862 ), .A2(_AES_ENC_us12_n861 ), .A3(_AES_ENC_us12_n860 ), .A4(_AES_ENC_us12_n859 ), .ZN(_AES_ENC_us12_n863 ) );
NAND2_X2 _AES_ENC_us12_U205  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n863 ), .ZN(_AES_ENC_us12_n905 ) );
NAND2_X2 _AES_ENC_us12_U204  ( .A1(_AES_ENC_us12_n1010 ), .A2(_AES_ENC_us12_n989 ), .ZN(_AES_ENC_us12_n874 ) );
NAND2_X2 _AES_ENC_us12_U203  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n610 ), .ZN(_AES_ENC_us12_n864 ) );
NAND2_X2 _AES_ENC_us12_U202  ( .A1(_AES_ENC_us12_n929 ), .A2(_AES_ENC_us12_n864 ), .ZN(_AES_ENC_us12_n873 ) );
NAND4_X2 _AES_ENC_us12_U193  ( .A1(_AES_ENC_us12_n874 ), .A2(_AES_ENC_us12_n873 ), .A3(_AES_ENC_us12_n872 ), .A4(_AES_ENC_us12_n871 ), .ZN(_AES_ENC_us12_n875 ) );
NAND2_X2 _AES_ENC_us12_U192  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n875 ), .ZN(_AES_ENC_us12_n904 ) );
NAND2_X2 _AES_ENC_us12_U191  ( .A1(_AES_ENC_us12_n583 ), .A2(_AES_ENC_us12_n1050 ), .ZN(_AES_ENC_us12_n889 ) );
NAND2_X2 _AES_ENC_us12_U190  ( .A1(_AES_ENC_us12_n1093 ), .A2(_AES_ENC_us12_n587 ), .ZN(_AES_ENC_us12_n876 ) );
NAND2_X2 _AES_ENC_us12_U189  ( .A1(_AES_ENC_us12_n604 ), .A2(_AES_ENC_us12_n876 ), .ZN(_AES_ENC_us12_n877 ) );
NAND2_X2 _AES_ENC_us12_U188  ( .A1(_AES_ENC_us12_n877 ), .A2(_AES_ENC_us12_n623 ), .ZN(_AES_ENC_us12_n888 ) );
NAND4_X2 _AES_ENC_us12_U179  ( .A1(_AES_ENC_us12_n889 ), .A2(_AES_ENC_us12_n888 ), .A3(_AES_ENC_us12_n887 ), .A4(_AES_ENC_us12_n886 ), .ZN(_AES_ENC_us12_n890 ) );
NAND2_X2 _AES_ENC_us12_U178  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n890 ), .ZN(_AES_ENC_us12_n903 ) );
OR2_X2 _AES_ENC_us12_U177  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n1059 ), .ZN(_AES_ENC_us12_n900 ) );
NAND2_X2 _AES_ENC_us12_U176  ( .A1(_AES_ENC_us12_n1073 ), .A2(_AES_ENC_us12_n1047 ), .ZN(_AES_ENC_us12_n899 ) );
NAND2_X2 _AES_ENC_us12_U175  ( .A1(_AES_ENC_us12_n1094 ), .A2(_AES_ENC_us12_n595 ), .ZN(_AES_ENC_us12_n898 ) );
NAND4_X2 _AES_ENC_us12_U167  ( .A1(_AES_ENC_us12_n900 ), .A2(_AES_ENC_us12_n899 ), .A3(_AES_ENC_us12_n898 ), .A4(_AES_ENC_us12_n897 ), .ZN(_AES_ENC_us12_n901 ) );
NAND2_X2 _AES_ENC_us12_U166  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n901 ), .ZN(_AES_ENC_us12_n902 ) );
NAND4_X2 _AES_ENC_us12_U165  ( .A1(_AES_ENC_us12_n905 ), .A2(_AES_ENC_us12_n904 ), .A3(_AES_ENC_us12_n903 ), .A4(_AES_ENC_us12_n902 ), .ZN(_AES_ENC_sa12_sub[4] ) );
NAND2_X2 _AES_ENC_us12_U164  ( .A1(_AES_ENC_us12_n1094 ), .A2(_AES_ENC_us12_n599 ), .ZN(_AES_ENC_us12_n922 ) );
NAND2_X2 _AES_ENC_us12_U163  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n989 ), .ZN(_AES_ENC_us12_n921 ) );
NAND4_X2 _AES_ENC_us12_U151  ( .A1(_AES_ENC_us12_n922 ), .A2(_AES_ENC_us12_n921 ), .A3(_AES_ENC_us12_n920 ), .A4(_AES_ENC_us12_n919 ), .ZN(_AES_ENC_us12_n923 ) );
NAND2_X2 _AES_ENC_us12_U150  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n923 ), .ZN(_AES_ENC_us12_n972 ) );
NAND2_X2 _AES_ENC_us12_U149  ( .A1(_AES_ENC_us12_n582 ), .A2(_AES_ENC_us12_n619 ), .ZN(_AES_ENC_us12_n924 ) );
NAND2_X2 _AES_ENC_us12_U148  ( .A1(_AES_ENC_us12_n1073 ), .A2(_AES_ENC_us12_n924 ), .ZN(_AES_ENC_us12_n939 ) );
NAND2_X2 _AES_ENC_us12_U147  ( .A1(_AES_ENC_us12_n926 ), .A2(_AES_ENC_us12_n925 ), .ZN(_AES_ENC_us12_n927 ) );
NAND2_X2 _AES_ENC_us12_U146  ( .A1(_AES_ENC_us12_n606 ), .A2(_AES_ENC_us12_n927 ), .ZN(_AES_ENC_us12_n928 ) );
NAND2_X2 _AES_ENC_us12_U145  ( .A1(_AES_ENC_us12_n928 ), .A2(_AES_ENC_us12_n1080 ), .ZN(_AES_ENC_us12_n938 ) );
OR2_X2 _AES_ENC_us12_U144  ( .A1(_AES_ENC_us12_n1117 ), .A2(_AES_ENC_us12_n615 ), .ZN(_AES_ENC_us12_n937 ) );
NAND4_X2 _AES_ENC_us12_U139  ( .A1(_AES_ENC_us12_n939 ), .A2(_AES_ENC_us12_n938 ), .A3(_AES_ENC_us12_n937 ), .A4(_AES_ENC_us12_n936 ), .ZN(_AES_ENC_us12_n940 ) );
NAND2_X2 _AES_ENC_us12_U138  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n940 ), .ZN(_AES_ENC_us12_n971 ) );
OR2_X2 _AES_ENC_us12_U137  ( .A1(_AES_ENC_us12_n605 ), .A2(_AES_ENC_us12_n941 ), .ZN(_AES_ENC_us12_n954 ) );
NAND2_X2 _AES_ENC_us12_U136  ( .A1(_AES_ENC_us12_n1096 ), .A2(_AES_ENC_us12_n577 ), .ZN(_AES_ENC_us12_n942 ) );
NAND2_X2 _AES_ENC_us12_U135  ( .A1(_AES_ENC_us12_n1048 ), .A2(_AES_ENC_us12_n942 ), .ZN(_AES_ENC_us12_n943 ) );
NAND2_X2 _AES_ENC_us12_U134  ( .A1(_AES_ENC_us12_n612 ), .A2(_AES_ENC_us12_n943 ), .ZN(_AES_ENC_us12_n944 ) );
NAND2_X2 _AES_ENC_us12_U133  ( .A1(_AES_ENC_us12_n944 ), .A2(_AES_ENC_us12_n580 ), .ZN(_AES_ENC_us12_n953 ) );
NAND4_X2 _AES_ENC_us12_U125  ( .A1(_AES_ENC_us12_n954 ), .A2(_AES_ENC_us12_n953 ), .A3(_AES_ENC_us12_n952 ), .A4(_AES_ENC_us12_n951 ), .ZN(_AES_ENC_us12_n955 ) );
NAND2_X2 _AES_ENC_us12_U124  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n955 ), .ZN(_AES_ENC_us12_n970 ) );
NAND2_X2 _AES_ENC_us12_U123  ( .A1(_AES_ENC_us12_n1094 ), .A2(_AES_ENC_us12_n1071 ), .ZN(_AES_ENC_us12_n967 ) );
NAND2_X2 _AES_ENC_us12_U122  ( .A1(_AES_ENC_us12_n956 ), .A2(_AES_ENC_us12_n1030 ), .ZN(_AES_ENC_us12_n966 ) );
NAND4_X2 _AES_ENC_us12_U114  ( .A1(_AES_ENC_us12_n967 ), .A2(_AES_ENC_us12_n966 ), .A3(_AES_ENC_us12_n965 ), .A4(_AES_ENC_us12_n964 ), .ZN(_AES_ENC_us12_n968 ) );
NAND2_X2 _AES_ENC_us12_U113  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n968 ), .ZN(_AES_ENC_us12_n969 ) );
NAND4_X2 _AES_ENC_us12_U112  ( .A1(_AES_ENC_us12_n972 ), .A2(_AES_ENC_us12_n971 ), .A3(_AES_ENC_us12_n970 ), .A4(_AES_ENC_us12_n969 ), .ZN(_AES_ENC_sa12_sub[5] ) );
NAND2_X2 _AES_ENC_us12_U111  ( .A1(_AES_ENC_us12_n570 ), .A2(_AES_ENC_us12_n1097 ), .ZN(_AES_ENC_us12_n973 ) );
NAND2_X2 _AES_ENC_us12_U110  ( .A1(_AES_ENC_us12_n1073 ), .A2(_AES_ENC_us12_n973 ), .ZN(_AES_ENC_us12_n987 ) );
NAND2_X2 _AES_ENC_us12_U109  ( .A1(_AES_ENC_us12_n974 ), .A2(_AES_ENC_us12_n1077 ), .ZN(_AES_ENC_us12_n975 ) );
NAND2_X2 _AES_ENC_us12_U108  ( .A1(_AES_ENC_us12_n613 ), .A2(_AES_ENC_us12_n975 ), .ZN(_AES_ENC_us12_n976 ) );
NAND2_X2 _AES_ENC_us12_U107  ( .A1(_AES_ENC_us12_n977 ), .A2(_AES_ENC_us12_n976 ), .ZN(_AES_ENC_us12_n986 ) );
NAND4_X2 _AES_ENC_us12_U99  ( .A1(_AES_ENC_us12_n987 ), .A2(_AES_ENC_us12_n986 ), .A3(_AES_ENC_us12_n985 ), .A4(_AES_ENC_us12_n984 ), .ZN(_AES_ENC_us12_n988 ) );
NAND2_X2 _AES_ENC_us12_U98  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n988 ), .ZN(_AES_ENC_us12_n1044 ) );
NAND2_X2 _AES_ENC_us12_U97  ( .A1(_AES_ENC_us12_n1073 ), .A2(_AES_ENC_us12_n989 ), .ZN(_AES_ENC_us12_n1004 ) );
NAND2_X2 _AES_ENC_us12_U96  ( .A1(_AES_ENC_us12_n1092 ), .A2(_AES_ENC_us12_n619 ), .ZN(_AES_ENC_us12_n1003 ) );
NAND4_X2 _AES_ENC_us12_U85  ( .A1(_AES_ENC_us12_n1004 ), .A2(_AES_ENC_us12_n1003 ), .A3(_AES_ENC_us12_n1002 ), .A4(_AES_ENC_us12_n1001 ), .ZN(_AES_ENC_us12_n1005 ) );
NAND2_X2 _AES_ENC_us12_U84  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n1005 ), .ZN(_AES_ENC_us12_n1043 ) );
NAND2_X2 _AES_ENC_us12_U83  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n596 ), .ZN(_AES_ENC_us12_n1020 ) );
NAND2_X2 _AES_ENC_us12_U82  ( .A1(_AES_ENC_us12_n1050 ), .A2(_AES_ENC_us12_n624 ), .ZN(_AES_ENC_us12_n1019 ) );
NAND2_X2 _AES_ENC_us12_U77  ( .A1(_AES_ENC_us12_n1059 ), .A2(_AES_ENC_us12_n1114 ), .ZN(_AES_ENC_us12_n1012 ) );
NAND2_X2 _AES_ENC_us12_U76  ( .A1(_AES_ENC_us12_n1010 ), .A2(_AES_ENC_us12_n592 ), .ZN(_AES_ENC_us12_n1011 ) );
NAND2_X2 _AES_ENC_us12_U75  ( .A1(_AES_ENC_us12_n1012 ), .A2(_AES_ENC_us12_n1011 ), .ZN(_AES_ENC_us12_n1016 ) );
NAND4_X2 _AES_ENC_us12_U70  ( .A1(_AES_ENC_us12_n1020 ), .A2(_AES_ENC_us12_n1019 ), .A3(_AES_ENC_us12_n1018 ), .A4(_AES_ENC_us12_n1017 ), .ZN(_AES_ENC_us12_n1021 ) );
NAND2_X2 _AES_ENC_us12_U69  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n1021 ), .ZN(_AES_ENC_us12_n1042 ) );
NAND2_X2 _AES_ENC_us12_U68  ( .A1(_AES_ENC_us12_n1022 ), .A2(_AES_ENC_us12_n1093 ), .ZN(_AES_ENC_us12_n1039 ) );
NAND2_X2 _AES_ENC_us12_U67  ( .A1(_AES_ENC_us12_n1050 ), .A2(_AES_ENC_us12_n1023 ), .ZN(_AES_ENC_us12_n1038 ) );
NAND2_X2 _AES_ENC_us12_U66  ( .A1(_AES_ENC_us12_n1024 ), .A2(_AES_ENC_us12_n1071 ), .ZN(_AES_ENC_us12_n1037 ) );
AND2_X2 _AES_ENC_us12_U60  ( .A1(_AES_ENC_us12_n1030 ), .A2(_AES_ENC_us12_n602 ), .ZN(_AES_ENC_us12_n1078 ) );
NAND4_X2 _AES_ENC_us12_U56  ( .A1(_AES_ENC_us12_n1039 ), .A2(_AES_ENC_us12_n1038 ), .A3(_AES_ENC_us12_n1037 ), .A4(_AES_ENC_us12_n1036 ), .ZN(_AES_ENC_us12_n1040 ) );
NAND2_X2 _AES_ENC_us12_U55  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n1040 ), .ZN(_AES_ENC_us12_n1041 ) );
NAND4_X2 _AES_ENC_us12_U54  ( .A1(_AES_ENC_us12_n1044 ), .A2(_AES_ENC_us12_n1043 ), .A3(_AES_ENC_us12_n1042 ), .A4(_AES_ENC_us12_n1041 ), .ZN(_AES_ENC_sa12_sub[6] ) );
NAND2_X2 _AES_ENC_us12_U53  ( .A1(_AES_ENC_us12_n1072 ), .A2(_AES_ENC_us12_n1045 ), .ZN(_AES_ENC_us12_n1068 ) );
NAND2_X2 _AES_ENC_us12_U52  ( .A1(_AES_ENC_us12_n1046 ), .A2(_AES_ENC_us12_n582 ), .ZN(_AES_ENC_us12_n1067 ) );
NAND2_X2 _AES_ENC_us12_U51  ( .A1(_AES_ENC_us12_n1094 ), .A2(_AES_ENC_us12_n1047 ), .ZN(_AES_ENC_us12_n1066 ) );
NAND4_X2 _AES_ENC_us12_U40  ( .A1(_AES_ENC_us12_n1068 ), .A2(_AES_ENC_us12_n1067 ), .A3(_AES_ENC_us12_n1066 ), .A4(_AES_ENC_us12_n1065 ), .ZN(_AES_ENC_us12_n1069 ) );
NAND2_X2 _AES_ENC_us12_U39  ( .A1(_AES_ENC_us12_n1070 ), .A2(_AES_ENC_us12_n1069 ), .ZN(_AES_ENC_us12_n1135 ) );
NAND2_X2 _AES_ENC_us12_U38  ( .A1(_AES_ENC_us12_n1072 ), .A2(_AES_ENC_us12_n1071 ), .ZN(_AES_ENC_us12_n1088 ) );
NAND2_X2 _AES_ENC_us12_U37  ( .A1(_AES_ENC_us12_n1073 ), .A2(_AES_ENC_us12_n595 ), .ZN(_AES_ENC_us12_n1087 ) );
NAND4_X2 _AES_ENC_us12_U28  ( .A1(_AES_ENC_us12_n1088 ), .A2(_AES_ENC_us12_n1087 ), .A3(_AES_ENC_us12_n1086 ), .A4(_AES_ENC_us12_n1085 ), .ZN(_AES_ENC_us12_n1089 ) );
NAND2_X2 _AES_ENC_us12_U27  ( .A1(_AES_ENC_us12_n1090 ), .A2(_AES_ENC_us12_n1089 ), .ZN(_AES_ENC_us12_n1134 ) );
NAND2_X2 _AES_ENC_us12_U26  ( .A1(_AES_ENC_us12_n1091 ), .A2(_AES_ENC_us12_n1093 ), .ZN(_AES_ENC_us12_n1111 ) );
NAND2_X2 _AES_ENC_us12_U25  ( .A1(_AES_ENC_us12_n1092 ), .A2(_AES_ENC_us12_n1120 ), .ZN(_AES_ENC_us12_n1110 ) );
AND2_X2 _AES_ENC_us12_U22  ( .A1(_AES_ENC_us12_n1097 ), .A2(_AES_ENC_us12_n1096 ), .ZN(_AES_ENC_us12_n1098 ) );
NAND4_X2 _AES_ENC_us12_U14  ( .A1(_AES_ENC_us12_n1111 ), .A2(_AES_ENC_us12_n1110 ), .A3(_AES_ENC_us12_n1109 ), .A4(_AES_ENC_us12_n1108 ), .ZN(_AES_ENC_us12_n1112 ) );
NAND2_X2 _AES_ENC_us12_U13  ( .A1(_AES_ENC_us12_n1113 ), .A2(_AES_ENC_us12_n1112 ), .ZN(_AES_ENC_us12_n1133 ) );
NAND2_X2 _AES_ENC_us12_U12  ( .A1(_AES_ENC_us12_n1115 ), .A2(_AES_ENC_us12_n1114 ), .ZN(_AES_ENC_us12_n1129 ) );
OR2_X2 _AES_ENC_us12_U11  ( .A1(_AES_ENC_us12_n608 ), .A2(_AES_ENC_us12_n1116 ), .ZN(_AES_ENC_us12_n1128 ) );
NAND4_X2 _AES_ENC_us12_U3  ( .A1(_AES_ENC_us12_n1129 ), .A2(_AES_ENC_us12_n1128 ), .A3(_AES_ENC_us12_n1127 ), .A4(_AES_ENC_us12_n1126 ), .ZN(_AES_ENC_us12_n1130 ) );
NAND2_X2 _AES_ENC_us12_U2  ( .A1(_AES_ENC_us12_n1131 ), .A2(_AES_ENC_us12_n1130 ), .ZN(_AES_ENC_us12_n1132 ) );
NAND4_X2 _AES_ENC_us12_U1  ( .A1(_AES_ENC_us12_n1135 ), .A2(_AES_ENC_us12_n1134 ), .A3(_AES_ENC_us12_n1133 ), .A4(_AES_ENC_us12_n1132 ), .ZN(_AES_ENC_sa12_sub[7] ) );
INV_X4 _AES_ENC_us13_U575  ( .A(_AES_ENC_sa13[0]), .ZN(_AES_ENC_us13_n627 ));
INV_X4 _AES_ENC_us13_U574  ( .A(_AES_ENC_us13_n1053 ), .ZN(_AES_ENC_us13_n625 ) );
INV_X4 _AES_ENC_us13_U573  ( .A(_AES_ENC_us13_n1103 ), .ZN(_AES_ENC_us13_n623 ) );
INV_X4 _AES_ENC_us13_U572  ( .A(_AES_ENC_us13_n1056 ), .ZN(_AES_ENC_us13_n622 ) );
INV_X4 _AES_ENC_us13_U571  ( .A(_AES_ENC_us13_n1102 ), .ZN(_AES_ENC_us13_n621 ) );
INV_X4 _AES_ENC_us13_U570  ( .A(_AES_ENC_us13_n1074 ), .ZN(_AES_ENC_us13_n620 ) );
INV_X4 _AES_ENC_us13_U569  ( .A(_AES_ENC_us13_n929 ), .ZN(_AES_ENC_us13_n619 ) );
INV_X4 _AES_ENC_us13_U568  ( .A(_AES_ENC_us13_n1091 ), .ZN(_AES_ENC_us13_n618 ) );
INV_X4 _AES_ENC_us13_U567  ( .A(_AES_ENC_us13_n826 ), .ZN(_AES_ENC_us13_n617 ) );
INV_X4 _AES_ENC_us13_U566  ( .A(_AES_ENC_us13_n1031 ), .ZN(_AES_ENC_us13_n616 ) );
INV_X4 _AES_ENC_us13_U565  ( .A(_AES_ENC_us13_n1054 ), .ZN(_AES_ENC_us13_n615 ) );
INV_X4 _AES_ENC_us13_U564  ( .A(_AES_ENC_us13_n1025 ), .ZN(_AES_ENC_us13_n614 ) );
INV_X4 _AES_ENC_us13_U563  ( .A(_AES_ENC_us13_n990 ), .ZN(_AES_ENC_us13_n613 ) );
INV_X4 _AES_ENC_us13_U562  ( .A(_AES_ENC_sa13[4]), .ZN(_AES_ENC_us13_n612 ));
INV_X4 _AES_ENC_us13_U561  ( .A(_AES_ENC_us13_n881 ), .ZN(_AES_ENC_us13_n611 ) );
INV_X4 _AES_ENC_us13_U560  ( .A(_AES_ENC_us13_n1022 ), .ZN(_AES_ENC_us13_n610 ) );
INV_X4 _AES_ENC_us13_U559  ( .A(_AES_ENC_us13_n1120 ), .ZN(_AES_ENC_us13_n609 ) );
INV_X4 _AES_ENC_us13_U558  ( .A(_AES_ENC_us13_n977 ), .ZN(_AES_ENC_us13_n608 ) );
INV_X4 _AES_ENC_us13_U557  ( .A(_AES_ENC_us13_n926 ), .ZN(_AES_ENC_us13_n607 ) );
INV_X4 _AES_ENC_us13_U556  ( .A(_AES_ENC_us13_n910 ), .ZN(_AES_ENC_us13_n606 ) );
INV_X4 _AES_ENC_us13_U555  ( .A(_AES_ENC_us13_n1121 ), .ZN(_AES_ENC_us13_n605 ) );
INV_X4 _AES_ENC_us13_U554  ( .A(_AES_ENC_us13_n1009 ), .ZN(_AES_ENC_us13_n604 ) );
INV_X4 _AES_ENC_us13_U553  ( .A(_AES_ENC_us13_n1080 ), .ZN(_AES_ENC_us13_n602 ) );
INV_X4 _AES_ENC_us13_U552  ( .A(_AES_ENC_us13_n821 ), .ZN(_AES_ENC_us13_n600 ) );
INV_X4 _AES_ENC_us13_U551  ( .A(_AES_ENC_us13_n1013 ), .ZN(_AES_ENC_us13_n599 ) );
INV_X4 _AES_ENC_us13_U550  ( .A(_AES_ENC_us13_n1058 ), .ZN(_AES_ENC_us13_n598 ) );
INV_X4 _AES_ENC_us13_U549  ( .A(_AES_ENC_us13_n906 ), .ZN(_AES_ENC_us13_n597 ) );
INV_X4 _AES_ENC_us13_U548  ( .A(_AES_ENC_us13_n959 ), .ZN(_AES_ENC_us13_n596 ) );
INV_X4 _AES_ENC_us13_U547  ( .A(_AES_ENC_sa13[7]), .ZN(_AES_ENC_us13_n595 ));
INV_X4 _AES_ENC_us13_U546  ( .A(_AES_ENC_us13_n1114 ), .ZN(_AES_ENC_us13_n593 ) );
INV_X4 _AES_ENC_us13_U545  ( .A(_AES_ENC_us13_n1048 ), .ZN(_AES_ENC_us13_n592 ) );
INV_X4 _AES_ENC_us13_U544  ( .A(_AES_ENC_us13_n974 ), .ZN(_AES_ENC_us13_n590 ) );
INV_X4 _AES_ENC_us13_U543  ( .A(_AES_ENC_us13_n794 ), .ZN(_AES_ENC_us13_n588 ) );
INV_X4 _AES_ENC_us13_U542  ( .A(_AES_ENC_us13_n880 ), .ZN(_AES_ENC_us13_n586 ) );
INV_X4 _AES_ENC_us13_U541  ( .A(_AES_ENC_sa13[2]), .ZN(_AES_ENC_us13_n584 ));
INV_X4 _AES_ENC_us13_U540  ( .A(_AES_ENC_us13_n800 ), .ZN(_AES_ENC_us13_n583 ) );
INV_X4 _AES_ENC_us13_U539  ( .A(_AES_ENC_us13_n925 ), .ZN(_AES_ENC_us13_n582 ) );
INV_X4 _AES_ENC_us13_U538  ( .A(_AES_ENC_us13_n992 ), .ZN(_AES_ENC_us13_n580 ) );
INV_X4 _AES_ENC_us13_U537  ( .A(_AES_ENC_us13_n779 ), .ZN(_AES_ENC_us13_n579 ) );
INV_X4 _AES_ENC_us13_U536  ( .A(_AES_ENC_us13_n1092 ), .ZN(_AES_ENC_us13_n575 ) );
INV_X4 _AES_ENC_us13_U535  ( .A(_AES_ENC_us13_n824 ), .ZN(_AES_ENC_us13_n574 ) );
NOR2_X2 _AES_ENC_us13_U534  ( .A1(_AES_ENC_sa13[0]), .A2(_AES_ENC_sa13[6]),.ZN(_AES_ENC_us13_n1090 ) );
NOR2_X2 _AES_ENC_us13_U533  ( .A1(_AES_ENC_us13_n627 ), .A2(_AES_ENC_sa13[6]), .ZN(_AES_ENC_us13_n1070 ) );
NOR2_X2 _AES_ENC_us13_U532  ( .A1(_AES_ENC_sa13[4]), .A2(_AES_ENC_sa13[3]),.ZN(_AES_ENC_us13_n1025 ) );
INV_X4 _AES_ENC_us13_U531  ( .A(_AES_ENC_us13_n569 ), .ZN(_AES_ENC_us13_n572 ) );
NOR2_X2 _AES_ENC_us13_U530  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n765 ) );
NOR2_X2 _AES_ENC_us13_U529  ( .A1(_AES_ENC_sa13[4]), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n764 ) );
NOR2_X2 _AES_ENC_us13_U528  ( .A1(_AES_ENC_us13_n765 ), .A2(_AES_ENC_us13_n764 ), .ZN(_AES_ENC_us13_n766 ) );
NOR2_X2 _AES_ENC_us13_U527  ( .A1(_AES_ENC_us13_n766 ), .A2(_AES_ENC_us13_n596 ), .ZN(_AES_ENC_us13_n767 ) );
NOR3_X2 _AES_ENC_us13_U526  ( .A1(_AES_ENC_us13_n595 ), .A2(_AES_ENC_sa13[5]), .A3(_AES_ENC_us13_n704 ), .ZN(_AES_ENC_us13_n706 ));
NOR2_X2 _AES_ENC_us13_U525  ( .A1(_AES_ENC_us13_n1117 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n707 ) );
NOR2_X2 _AES_ENC_us13_U524  ( .A1(_AES_ENC_sa13[4]), .A2(_AES_ENC_us13_n575 ), .ZN(_AES_ENC_us13_n705 ) );
NOR3_X2 _AES_ENC_us13_U523  ( .A1(_AES_ENC_us13_n707 ), .A2(_AES_ENC_us13_n706 ), .A3(_AES_ENC_us13_n705 ), .ZN(_AES_ENC_us13_n713 ) );
INV_X4 _AES_ENC_us13_U522  ( .A(_AES_ENC_sa13[3]), .ZN(_AES_ENC_us13_n624 ));
NAND3_X2 _AES_ENC_us13_U521  ( .A1(_AES_ENC_us13_n652 ), .A2(_AES_ENC_us13_n594 ), .A3(_AES_ENC_sa13[7]), .ZN(_AES_ENC_us13_n653 ));
NOR2_X2 _AES_ENC_us13_U520  ( .A1(_AES_ENC_us13_n584 ), .A2(_AES_ENC_sa13[5]), .ZN(_AES_ENC_us13_n925 ) );
NOR2_X2 _AES_ENC_us13_U519  ( .A1(_AES_ENC_sa13[5]), .A2(_AES_ENC_sa13[2]),.ZN(_AES_ENC_us13_n974 ) );
INV_X4 _AES_ENC_us13_U518  ( .A(_AES_ENC_sa13[5]), .ZN(_AES_ENC_us13_n594 ));
NOR2_X2 _AES_ENC_us13_U517  ( .A1(_AES_ENC_us13_n584 ), .A2(_AES_ENC_sa13[7]), .ZN(_AES_ENC_us13_n779 ) );
NAND3_X2 _AES_ENC_us13_U516  ( .A1(_AES_ENC_us13_n679 ), .A2(_AES_ENC_us13_n678 ), .A3(_AES_ENC_us13_n677 ), .ZN(_AES_ENC_sa13_sub[0] ) );
NOR2_X2 _AES_ENC_us13_U515  ( .A1(_AES_ENC_us13_n594 ), .A2(_AES_ENC_sa13[2]), .ZN(_AES_ENC_us13_n1048 ) );
NOR4_X2 _AES_ENC_us13_U512  ( .A1(_AES_ENC_us13_n633 ), .A2(_AES_ENC_us13_n632 ), .A3(_AES_ENC_us13_n631 ), .A4(_AES_ENC_us13_n630 ), .ZN(_AES_ENC_us13_n634 ) );
NOR2_X2 _AES_ENC_us13_U510  ( .A1(_AES_ENC_us13_n629 ), .A2(_AES_ENC_us13_n628 ), .ZN(_AES_ENC_us13_n635 ) );
NAND3_X2 _AES_ENC_us13_U509  ( .A1(_AES_ENC_sa13[2]), .A2(_AES_ENC_sa13[7]), .A3(_AES_ENC_us13_n1059 ), .ZN(_AES_ENC_us13_n636 ) );
NOR2_X2 _AES_ENC_us13_U508  ( .A1(_AES_ENC_sa13[7]), .A2(_AES_ENC_sa13[2]),.ZN(_AES_ENC_us13_n794 ) );
NOR2_X2 _AES_ENC_us13_U507  ( .A1(_AES_ENC_sa13[4]), .A2(_AES_ENC_sa13[1]),.ZN(_AES_ENC_us13_n1102 ) );
NOR2_X2 _AES_ENC_us13_U506  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_sa13[3]), .ZN(_AES_ENC_us13_n1053 ) );
NOR2_X2 _AES_ENC_us13_U505  ( .A1(_AES_ENC_us13_n579 ), .A2(_AES_ENC_sa13[5]), .ZN(_AES_ENC_us13_n1024 ) );
NOR2_X2 _AES_ENC_us13_U504  ( .A1(_AES_ENC_us13_n593 ), .A2(_AES_ENC_sa13[2]), .ZN(_AES_ENC_us13_n1093 ) );
NOR2_X2 _AES_ENC_us13_U503  ( .A1(_AES_ENC_us13_n588 ), .A2(_AES_ENC_sa13[5]), .ZN(_AES_ENC_us13_n1094 ) );
NOR2_X2 _AES_ENC_us13_U502  ( .A1(_AES_ENC_us13_n612 ), .A2(_AES_ENC_sa13[3]), .ZN(_AES_ENC_us13_n931 ) );
INV_X4 _AES_ENC_us13_U501  ( .A(_AES_ENC_us13_n570 ), .ZN(_AES_ENC_us13_n573 ) );
NOR2_X2 _AES_ENC_us13_U500  ( .A1(_AES_ENC_us13_n1053 ), .A2(_AES_ENC_us13_n1095 ), .ZN(_AES_ENC_us13_n639 ) );
NOR3_X2 _AES_ENC_us13_U499  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n573 ), .A3(_AES_ENC_us13_n1074 ), .ZN(_AES_ENC_us13_n641 ) );
NOR2_X2 _AES_ENC_us13_U498  ( .A1(_AES_ENC_us13_n639 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n640 ) );
NOR2_X2 _AES_ENC_us13_U497  ( .A1(_AES_ENC_us13_n641 ), .A2(_AES_ENC_us13_n640 ), .ZN(_AES_ENC_us13_n646 ) );
NOR3_X2 _AES_ENC_us13_U496  ( .A1(_AES_ENC_us13_n995 ), .A2(_AES_ENC_us13_n580 ), .A3(_AES_ENC_us13_n994 ), .ZN(_AES_ENC_us13_n1002 ) );
NOR2_X2 _AES_ENC_us13_U495  ( .A1(_AES_ENC_us13_n909 ), .A2(_AES_ENC_us13_n908 ), .ZN(_AES_ENC_us13_n920 ) );
NOR2_X2 _AES_ENC_us13_U494  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n823 ) );
NOR2_X2 _AES_ENC_us13_U492  ( .A1(_AES_ENC_us13_n612 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n822 ) );
NOR2_X2 _AES_ENC_us13_U491  ( .A1(_AES_ENC_us13_n823 ), .A2(_AES_ENC_us13_n822 ), .ZN(_AES_ENC_us13_n825 ) );
NOR2_X2 _AES_ENC_us13_U490  ( .A1(_AES_ENC_sa13[1]), .A2(_AES_ENC_us13_n601 ), .ZN(_AES_ENC_us13_n913 ) );
NOR2_X2 _AES_ENC_us13_U489  ( .A1(_AES_ENC_us13_n913 ), .A2(_AES_ENC_us13_n1091 ), .ZN(_AES_ENC_us13_n914 ) );
NOR2_X2 _AES_ENC_us13_U488  ( .A1(_AES_ENC_us13_n826 ), .A2(_AES_ENC_us13_n572 ), .ZN(_AES_ENC_us13_n827 ) );
NOR3_X2 _AES_ENC_us13_U487  ( .A1(_AES_ENC_us13_n769 ), .A2(_AES_ENC_us13_n768 ), .A3(_AES_ENC_us13_n767 ), .ZN(_AES_ENC_us13_n775 ) );
NOR2_X2 _AES_ENC_us13_U486  ( .A1(_AES_ENC_us13_n1056 ), .A2(_AES_ENC_us13_n1053 ), .ZN(_AES_ENC_us13_n749 ) );
NOR2_X2 _AES_ENC_us13_U483  ( .A1(_AES_ENC_us13_n749 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n752 ) );
INV_X4 _AES_ENC_us13_U482  ( .A(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n626 ));
NOR2_X2 _AES_ENC_us13_U480  ( .A1(_AES_ENC_us13_n1054 ), .A2(_AES_ENC_us13_n1053 ), .ZN(_AES_ENC_us13_n1055 ) );
OR2_X4 _AES_ENC_us13_U479  ( .A1(_AES_ENC_us13_n1094 ), .A2(_AES_ENC_us13_n1093 ), .ZN(_AES_ENC_us13_n571 ) );
AND2_X2 _AES_ENC_us13_U478  ( .A1(_AES_ENC_us13_n571 ), .A2(_AES_ENC_us13_n1095 ), .ZN(_AES_ENC_us13_n1101 ) );
NOR2_X2 _AES_ENC_us13_U477  ( .A1(_AES_ENC_us13_n1074 ), .A2(_AES_ENC_us13_n931 ), .ZN(_AES_ENC_us13_n796 ) );
NOR2_X2 _AES_ENC_us13_U474  ( .A1(_AES_ENC_us13_n796 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n797 ) );
NOR2_X2 _AES_ENC_us13_U473  ( .A1(_AES_ENC_us13_n932 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n933 ) );
NOR2_X2 _AES_ENC_us13_U472  ( .A1(_AES_ENC_us13_n929 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n935 ) );
NOR2_X2 _AES_ENC_us13_U471  ( .A1(_AES_ENC_us13_n931 ), .A2(_AES_ENC_us13_n930 ), .ZN(_AES_ENC_us13_n934 ) );
NOR3_X2 _AES_ENC_us13_U470  ( .A1(_AES_ENC_us13_n935 ), .A2(_AES_ENC_us13_n934 ), .A3(_AES_ENC_us13_n933 ), .ZN(_AES_ENC_us13_n936 ) );
NOR2_X2 _AES_ENC_us13_U469  ( .A1(_AES_ENC_us13_n612 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n1075 ) );
NOR2_X2 _AES_ENC_us13_U468  ( .A1(_AES_ENC_us13_n572 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n949 ) );
NOR2_X2 _AES_ENC_us13_U467  ( .A1(_AES_ENC_us13_n1049 ), .A2(_AES_ENC_us13_n592 ), .ZN(_AES_ENC_us13_n1051 ) );
NOR2_X2 _AES_ENC_us13_U466  ( .A1(_AES_ENC_us13_n1051 ), .A2(_AES_ENC_us13_n1050 ), .ZN(_AES_ENC_us13_n1052 ) );
NOR2_X2 _AES_ENC_us13_U465  ( .A1(_AES_ENC_us13_n1052 ), .A2(_AES_ENC_us13_n604 ), .ZN(_AES_ENC_us13_n1064 ) );
NOR2_X2 _AES_ENC_us13_U464  ( .A1(_AES_ENC_sa13[1]), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n631 ) );
NOR2_X2 _AES_ENC_us13_U463  ( .A1(_AES_ENC_us13_n1025 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n980 ) );
NOR2_X2 _AES_ENC_us13_U462  ( .A1(_AES_ENC_us13_n1073 ), .A2(_AES_ENC_us13_n1094 ), .ZN(_AES_ENC_us13_n795 ) );
NOR2_X2 _AES_ENC_us13_U461  ( .A1(_AES_ENC_us13_n795 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n799 ) );
NOR2_X2 _AES_ENC_us13_U460  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n981 ) );
NOR2_X2 _AES_ENC_us13_U459  ( .A1(_AES_ENC_us13_n1102 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n643 ) );
NOR2_X2 _AES_ENC_us13_U458  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n624 ), .ZN(_AES_ENC_us13_n642 ) );
NOR2_X2 _AES_ENC_us13_U455  ( .A1(_AES_ENC_us13_n911 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n644 ) );
NOR4_X2 _AES_ENC_us13_U448  ( .A1(_AES_ENC_us13_n644 ), .A2(_AES_ENC_us13_n643 ), .A3(_AES_ENC_us13_n804 ), .A4(_AES_ENC_us13_n642 ), .ZN(_AES_ENC_us13_n645 ) );
NOR2_X2 _AES_ENC_us13_U447  ( .A1(_AES_ENC_us13_n1102 ), .A2(_AES_ENC_us13_n910 ), .ZN(_AES_ENC_us13_n932 ) );
NOR2_X2 _AES_ENC_us13_U442  ( .A1(_AES_ENC_us13_n1102 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n755 ) );
NOR2_X2 _AES_ENC_us13_U441  ( .A1(_AES_ENC_us13_n931 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n743 ) );
NOR2_X2 _AES_ENC_us13_U438  ( .A1(_AES_ENC_us13_n1072 ), .A2(_AES_ENC_us13_n1094 ), .ZN(_AES_ENC_us13_n930 ) );
NOR2_X2 _AES_ENC_us13_U435  ( .A1(_AES_ENC_us13_n1074 ), .A2(_AES_ENC_us13_n1025 ), .ZN(_AES_ENC_us13_n891 ) );
NOR2_X2 _AES_ENC_us13_U434  ( .A1(_AES_ENC_us13_n891 ), .A2(_AES_ENC_us13_n582 ), .ZN(_AES_ENC_us13_n894 ) );
NOR3_X2 _AES_ENC_us13_U433  ( .A1(_AES_ENC_us13_n601 ), .A2(_AES_ENC_sa13[1]), .A3(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n683 ));
INV_X4 _AES_ENC_us13_U428  ( .A(_AES_ENC_us13_n931 ), .ZN(_AES_ENC_us13_n601 ) );
NOR2_X2 _AES_ENC_us13_U427  ( .A1(_AES_ENC_us13_n996 ), .A2(_AES_ENC_us13_n931 ), .ZN(_AES_ENC_us13_n704 ) );
NOR2_X2 _AES_ENC_us13_U421  ( .A1(_AES_ENC_us13_n931 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n685 ) );
NOR2_X2 _AES_ENC_us13_U420  ( .A1(_AES_ENC_us13_n1029 ), .A2(_AES_ENC_us13_n1025 ), .ZN(_AES_ENC_us13_n1079 ) );
NOR3_X2 _AES_ENC_us13_U419  ( .A1(_AES_ENC_us13_n620 ), .A2(_AES_ENC_us13_n1025 ), .A3(_AES_ENC_us13_n590 ), .ZN(_AES_ENC_us13_n945 ) );
NOR2_X2 _AES_ENC_us13_U418  ( .A1(_AES_ENC_us13_n594 ), .A2(_AES_ENC_us13_n584 ), .ZN(_AES_ENC_us13_n800 ) );
NOR3_X2 _AES_ENC_us13_U417  ( .A1(_AES_ENC_us13_n598 ), .A2(_AES_ENC_us13_n595 ), .A3(_AES_ENC_us13_n584 ), .ZN(_AES_ENC_us13_n798 ) );
NOR3_X2 _AES_ENC_us13_U416  ( .A1(_AES_ENC_us13_n583 ), .A2(_AES_ENC_us13_n572 ), .A3(_AES_ENC_us13_n596 ), .ZN(_AES_ENC_us13_n962 ) );
NOR3_X2 _AES_ENC_us13_U415  ( .A1(_AES_ENC_us13_n959 ), .A2(_AES_ENC_us13_n572 ), .A3(_AES_ENC_us13_n582 ), .ZN(_AES_ENC_us13_n768 ) );
NOR3_X2 _AES_ENC_us13_U414  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n572 ), .A3(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n694 ) );
NOR3_X2 _AES_ENC_us13_U413  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n572 ), .A3(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n895 ) );
NOR3_X2 _AES_ENC_us13_U410  ( .A1(_AES_ENC_us13_n1008 ), .A2(_AES_ENC_us13_n1007 ), .A3(_AES_ENC_us13_n1006 ), .ZN(_AES_ENC_us13_n1018 ) );
NOR4_X2 _AES_ENC_us13_U409  ( .A1(_AES_ENC_us13_n806 ), .A2(_AES_ENC_us13_n805 ), .A3(_AES_ENC_us13_n804 ), .A4(_AES_ENC_us13_n803 ), .ZN(_AES_ENC_us13_n807 ) );
NOR3_X2 _AES_ENC_us13_U406  ( .A1(_AES_ENC_us13_n799 ), .A2(_AES_ENC_us13_n798 ), .A3(_AES_ENC_us13_n797 ), .ZN(_AES_ENC_us13_n808 ) );
NOR4_X2 _AES_ENC_us13_U405  ( .A1(_AES_ENC_us13_n843 ), .A2(_AES_ENC_us13_n842 ), .A3(_AES_ENC_us13_n841 ), .A4(_AES_ENC_us13_n840 ), .ZN(_AES_ENC_us13_n844 ) );
NOR2_X2 _AES_ENC_us13_U404  ( .A1(_AES_ENC_us13_n669 ), .A2(_AES_ENC_us13_n668 ), .ZN(_AES_ENC_us13_n673 ) );
NOR4_X2 _AES_ENC_us13_U403  ( .A1(_AES_ENC_us13_n946 ), .A2(_AES_ENC_us13_n1046 ), .A3(_AES_ENC_us13_n671 ), .A4(_AES_ENC_us13_n670 ), .ZN(_AES_ENC_us13_n672 ) );
NOR4_X2 _AES_ENC_us13_U401  ( .A1(_AES_ENC_us13_n711 ), .A2(_AES_ENC_us13_n710 ), .A3(_AES_ENC_us13_n709 ), .A4(_AES_ENC_us13_n708 ), .ZN(_AES_ENC_us13_n712 ) );
NOR4_X2 _AES_ENC_us13_U400  ( .A1(_AES_ENC_us13_n963 ), .A2(_AES_ENC_us13_n962 ), .A3(_AES_ENC_us13_n961 ), .A4(_AES_ENC_us13_n960 ), .ZN(_AES_ENC_us13_n964 ) );
NOR3_X2 _AES_ENC_us13_U399  ( .A1(_AES_ENC_us13_n1101 ), .A2(_AES_ENC_us13_n1100 ), .A3(_AES_ENC_us13_n1099 ), .ZN(_AES_ENC_us13_n1109 ) );
NOR3_X2 _AES_ENC_us13_U398  ( .A1(_AES_ENC_us13_n743 ), .A2(_AES_ENC_us13_n742 ), .A3(_AES_ENC_us13_n741 ), .ZN(_AES_ENC_us13_n744 ) );
NOR2_X2 _AES_ENC_us13_U397  ( .A1(_AES_ENC_us13_n697 ), .A2(_AES_ENC_us13_n658 ), .ZN(_AES_ENC_us13_n659 ) );
NOR2_X2 _AES_ENC_us13_U396  ( .A1(_AES_ENC_us13_n1078 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n1033 ) );
NOR2_X2 _AES_ENC_us13_U393  ( .A1(_AES_ENC_us13_n1031 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n1032 ) );
NOR3_X2 _AES_ENC_us13_U390  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n1025 ), .A3(_AES_ENC_us13_n1074 ), .ZN(_AES_ENC_us13_n1035 ) );
NOR4_X2 _AES_ENC_us13_U389  ( .A1(_AES_ENC_us13_n1035 ), .A2(_AES_ENC_us13_n1034 ), .A3(_AES_ENC_us13_n1033 ), .A4(_AES_ENC_us13_n1032 ), .ZN(_AES_ENC_us13_n1036 ) );
NOR2_X2 _AES_ENC_us13_U388  ( .A1(_AES_ENC_us13_n611 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n885 ) );
NOR2_X2 _AES_ENC_us13_U387  ( .A1(_AES_ENC_us13_n601 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n882 ) );
NOR2_X2 _AES_ENC_us13_U386  ( .A1(_AES_ENC_us13_n1053 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n884 ) );
NOR4_X2 _AES_ENC_us13_U385  ( .A1(_AES_ENC_us13_n885 ), .A2(_AES_ENC_us13_n884 ), .A3(_AES_ENC_us13_n883 ), .A4(_AES_ENC_us13_n882 ), .ZN(_AES_ENC_us13_n886 ) );
NOR2_X2 _AES_ENC_us13_U384  ( .A1(_AES_ENC_us13_n825 ), .A2(_AES_ENC_us13_n574 ), .ZN(_AES_ENC_us13_n830 ) );
NOR2_X2 _AES_ENC_us13_U383  ( .A1(_AES_ENC_us13_n827 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n829 ) );
NOR2_X2 _AES_ENC_us13_U382  ( .A1(_AES_ENC_us13_n572 ), .A2(_AES_ENC_us13_n575 ), .ZN(_AES_ENC_us13_n828 ) );
NOR4_X2 _AES_ENC_us13_U374  ( .A1(_AES_ENC_us13_n831 ), .A2(_AES_ENC_us13_n830 ), .A3(_AES_ENC_us13_n829 ), .A4(_AES_ENC_us13_n828 ), .ZN(_AES_ENC_us13_n832 ) );
NOR2_X2 _AES_ENC_us13_U373  ( .A1(_AES_ENC_us13_n578 ), .A2(_AES_ENC_us13_n603 ), .ZN(_AES_ENC_us13_n1104 ) );
NOR2_X2 _AES_ENC_us13_U372  ( .A1(_AES_ENC_us13_n1102 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n1106 ) );
NOR2_X2 _AES_ENC_us13_U370  ( .A1(_AES_ENC_us13_n1103 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n1105 ) );
NOR4_X2 _AES_ENC_us13_U369  ( .A1(_AES_ENC_us13_n1107 ), .A2(_AES_ENC_us13_n1106 ), .A3(_AES_ENC_us13_n1105 ), .A4(_AES_ENC_us13_n1104 ), .ZN(_AES_ENC_us13_n1108 ) );
NOR3_X2 _AES_ENC_us13_U368  ( .A1(_AES_ENC_us13_n959 ), .A2(_AES_ENC_us13_n624 ), .A3(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n963 ) );
NOR2_X2 _AES_ENC_us13_U367  ( .A1(_AES_ENC_us13_n594 ), .A2(_AES_ENC_us13_n595 ), .ZN(_AES_ENC_us13_n1114 ) );
INV_X4 _AES_ENC_us13_U366  ( .A(_AES_ENC_us13_n1024 ), .ZN(_AES_ENC_us13_n578 ) );
NOR3_X2 _AES_ENC_us13_U365  ( .A1(_AES_ENC_us13_n910 ), .A2(_AES_ENC_us13_n1059 ), .A3(_AES_ENC_us13_n584 ), .ZN(_AES_ENC_us13_n1115 ) );
INV_X4 _AES_ENC_us13_U364  ( .A(_AES_ENC_us13_n1094 ), .ZN(_AES_ENC_us13_n587 ) );
NOR2_X2 _AES_ENC_us13_U363  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n931 ), .ZN(_AES_ENC_us13_n1100 ) );
INV_X4 _AES_ENC_us13_U354  ( .A(_AES_ENC_us13_n1093 ), .ZN(_AES_ENC_us13_n591 ) );
NOR2_X2 _AES_ENC_us13_U353  ( .A1(_AES_ENC_us13_n569 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n929 ) );
NOR2_X2 _AES_ENC_us13_U352  ( .A1(_AES_ENC_us13_n609 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n926 ) );
NOR2_X2 _AES_ENC_us13_U351  ( .A1(_AES_ENC_us13_n572 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n1095 ) );
NOR2_X2 _AES_ENC_us13_U350  ( .A1(_AES_ENC_us13_n582 ), .A2(_AES_ENC_us13_n595 ), .ZN(_AES_ENC_us13_n1010 ) );
NOR2_X2 _AES_ENC_us13_U349  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n1103 ) );
NOR2_X2 _AES_ENC_us13_U348  ( .A1(_AES_ENC_us13_n614 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n1059 ) );
NOR2_X2 _AES_ENC_us13_U347  ( .A1(_AES_ENC_sa13[1]), .A2(_AES_ENC_us13_n1120 ), .ZN(_AES_ENC_us13_n1022 ) );
NOR2_X2 _AES_ENC_us13_U346  ( .A1(_AES_ENC_us13_n605 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n911 ) );
NOR2_X2 _AES_ENC_us13_U345  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_us13_n1025 ), .ZN(_AES_ENC_us13_n826 ) );
NOR2_X2 _AES_ENC_us13_U338  ( .A1(_AES_ENC_us13_n594 ), .A2(_AES_ENC_us13_n579 ), .ZN(_AES_ENC_us13_n1072 ) );
NOR2_X2 _AES_ENC_us13_U335  ( .A1(_AES_ENC_us13_n595 ), .A2(_AES_ENC_us13_n590 ), .ZN(_AES_ENC_us13_n956 ) );
NOR2_X2 _AES_ENC_us13_U329  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_us13_n612 ), .ZN(_AES_ENC_us13_n1121 ) );
NOR2_X2 _AES_ENC_us13_U328  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_us13_n612 ), .ZN(_AES_ENC_us13_n1058 ) );
NOR2_X2 _AES_ENC_us13_U327  ( .A1(_AES_ENC_us13_n593 ), .A2(_AES_ENC_us13_n584 ), .ZN(_AES_ENC_us13_n1073 ) );
NOR2_X2 _AES_ENC_us13_U325  ( .A1(_AES_ENC_sa13[1]), .A2(_AES_ENC_us13_n1025 ), .ZN(_AES_ENC_us13_n1054 ) );
NOR2_X2 _AES_ENC_us13_U324  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_us13_n931 ), .ZN(_AES_ENC_us13_n1029 ) );
NOR2_X2 _AES_ENC_us13_U319  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n1056 ) );
NOR2_X2 _AES_ENC_us13_U318  ( .A1(_AES_ENC_us13_n588 ), .A2(_AES_ENC_us13_n594 ), .ZN(_AES_ENC_us13_n1050 ) );
NOR2_X2 _AES_ENC_us13_U317  ( .A1(_AES_ENC_us13_n1121 ), .A2(_AES_ENC_us13_n1025 ), .ZN(_AES_ENC_us13_n1120 ) );
NOR2_X2 _AES_ENC_us13_U316  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_us13_n572 ), .ZN(_AES_ENC_us13_n1074 ) );
NOR2_X2 _AES_ENC_us13_U315  ( .A1(_AES_ENC_us13_n1058 ), .A2(_AES_ENC_us13_n1054 ), .ZN(_AES_ENC_us13_n878 ) );
NOR2_X2 _AES_ENC_us13_U314  ( .A1(_AES_ENC_us13_n878 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n879 ) );
NOR2_X2 _AES_ENC_us13_U312  ( .A1(_AES_ENC_us13_n880 ), .A2(_AES_ENC_us13_n879 ), .ZN(_AES_ENC_us13_n887 ) );
NOR2_X2 _AES_ENC_us13_U311  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n625 ), .ZN(_AES_ENC_us13_n957 ) );
NOR2_X2 _AES_ENC_us13_U310  ( .A1(_AES_ENC_us13_n958 ), .A2(_AES_ENC_us13_n957 ), .ZN(_AES_ENC_us13_n965 ) );
NOR3_X2 _AES_ENC_us13_U309  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n1091 ), .A3(_AES_ENC_us13_n1022 ), .ZN(_AES_ENC_us13_n720 ) );
NOR3_X2 _AES_ENC_us13_U303  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n1054 ), .A3(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n719 ) );
NOR2_X2 _AES_ENC_us13_U302  ( .A1(_AES_ENC_us13_n720 ), .A2(_AES_ENC_us13_n719 ), .ZN(_AES_ENC_us13_n726 ) );
NOR2_X2 _AES_ENC_us13_U300  ( .A1(_AES_ENC_us13_n588 ), .A2(_AES_ENC_us13_n613 ), .ZN(_AES_ENC_us13_n865 ) );
NOR2_X2 _AES_ENC_us13_U299  ( .A1(_AES_ENC_us13_n1059 ), .A2(_AES_ENC_us13_n1058 ), .ZN(_AES_ENC_us13_n1060 ) );
NOR2_X2 _AES_ENC_us13_U298  ( .A1(_AES_ENC_us13_n1095 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n668 ) );
NOR2_X2 _AES_ENC_us13_U297  ( .A1(_AES_ENC_us13_n911 ), .A2(_AES_ENC_us13_n910 ), .ZN(_AES_ENC_us13_n912 ) );
NOR2_X2 _AES_ENC_us13_U296  ( .A1(_AES_ENC_us13_n912 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n916 ) );
NOR2_X2 _AES_ENC_us13_U295  ( .A1(_AES_ENC_us13_n826 ), .A2(_AES_ENC_us13_n573 ), .ZN(_AES_ENC_us13_n750 ) );
NOR2_X2 _AES_ENC_us13_U294  ( .A1(_AES_ENC_us13_n750 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n751 ) );
NOR2_X2 _AES_ENC_us13_U293  ( .A1(_AES_ENC_us13_n907 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n908 ) );
NOR2_X2 _AES_ENC_us13_U292  ( .A1(_AES_ENC_us13_n990 ), .A2(_AES_ENC_us13_n926 ), .ZN(_AES_ENC_us13_n780 ) );
NOR2_X2 _AES_ENC_us13_U291  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n606 ), .ZN(_AES_ENC_us13_n838 ) );
NOR2_X2 _AES_ENC_us13_U290  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n621 ), .ZN(_AES_ENC_us13_n837 ) );
NOR2_X2 _AES_ENC_us13_U284  ( .A1(_AES_ENC_us13_n838 ), .A2(_AES_ENC_us13_n837 ), .ZN(_AES_ENC_us13_n845 ) );
NOR2_X2 _AES_ENC_us13_U283  ( .A1(_AES_ENC_us13_n1022 ), .A2(_AES_ENC_us13_n1058 ), .ZN(_AES_ENC_us13_n740 ) );
NOR2_X2 _AES_ENC_us13_U282  ( .A1(_AES_ENC_us13_n740 ), .A2(_AES_ENC_us13_n590 ), .ZN(_AES_ENC_us13_n742 ) );
NOR2_X2 _AES_ENC_us13_U281  ( .A1(_AES_ENC_us13_n1098 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n1099 ) );
NOR2_X2 _AES_ENC_us13_U280  ( .A1(_AES_ENC_us13_n1120 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n993 ) );
NOR2_X2 _AES_ENC_us13_U279  ( .A1(_AES_ENC_us13_n993 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n994 ) );
NOR2_X2 _AES_ENC_us13_U273  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n609 ), .ZN(_AES_ENC_us13_n1026 ) );
NOR2_X2 _AES_ENC_us13_U272  ( .A1(_AES_ENC_us13_n573 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n1027 ) );
NOR2_X2 _AES_ENC_us13_U271  ( .A1(_AES_ENC_us13_n1027 ), .A2(_AES_ENC_us13_n1026 ), .ZN(_AES_ENC_us13_n1028 ) );
NOR2_X2 _AES_ENC_us13_U270  ( .A1(_AES_ENC_us13_n1029 ), .A2(_AES_ENC_us13_n1028 ), .ZN(_AES_ENC_us13_n1034 ) );
NOR4_X2 _AES_ENC_us13_U269  ( .A1(_AES_ENC_us13_n757 ), .A2(_AES_ENC_us13_n756 ), .A3(_AES_ENC_us13_n755 ), .A4(_AES_ENC_us13_n754 ), .ZN(_AES_ENC_us13_n758 ) );
NOR2_X2 _AES_ENC_us13_U268  ( .A1(_AES_ENC_us13_n752 ), .A2(_AES_ENC_us13_n751 ), .ZN(_AES_ENC_us13_n759 ) );
NOR2_X2 _AES_ENC_us13_U267  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n1071 ), .ZN(_AES_ENC_us13_n669 ) );
NOR2_X2 _AES_ENC_us13_U263  ( .A1(_AES_ENC_us13_n1056 ), .A2(_AES_ENC_us13_n990 ), .ZN(_AES_ENC_us13_n991 ) );
NOR2_X2 _AES_ENC_us13_U262  ( .A1(_AES_ENC_us13_n991 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n995 ) );
NOR2_X2 _AES_ENC_us13_U258  ( .A1(_AES_ENC_us13_n579 ), .A2(_AES_ENC_us13_n598 ), .ZN(_AES_ENC_us13_n1008 ) );
NOR2_X2 _AES_ENC_us13_U255  ( .A1(_AES_ENC_us13_n839 ), .A2(_AES_ENC_us13_n603 ), .ZN(_AES_ENC_us13_n693 ) );
NOR2_X2 _AES_ENC_us13_U254  ( .A1(_AES_ENC_us13_n578 ), .A2(_AES_ENC_us13_n906 ), .ZN(_AES_ENC_us13_n741 ) );
NOR2_X2 _AES_ENC_us13_U253  ( .A1(_AES_ENC_us13_n1054 ), .A2(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n763 ) );
NOR2_X2 _AES_ENC_us13_U252  ( .A1(_AES_ENC_us13_n763 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n769 ) );
NOR2_X2 _AES_ENC_us13_U251  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n618 ), .ZN(_AES_ENC_us13_n1007 ) );
NOR2_X2 _AES_ENC_us13_U250  ( .A1(_AES_ENC_us13_n582 ), .A2(_AES_ENC_us13_n599 ), .ZN(_AES_ENC_us13_n1123 ) );
NOR2_X2 _AES_ENC_us13_U243  ( .A1(_AES_ENC_us13_n582 ), .A2(_AES_ENC_us13_n598 ), .ZN(_AES_ENC_us13_n710 ) );
INV_X4 _AES_ENC_us13_U242  ( .A(_AES_ENC_us13_n1029 ), .ZN(_AES_ENC_us13_n603 ) );
NOR2_X2 _AES_ENC_us13_U241  ( .A1(_AES_ENC_us13_n590 ), .A2(_AES_ENC_us13_n607 ), .ZN(_AES_ENC_us13_n883 ) );
NOR2_X2 _AES_ENC_us13_U240  ( .A1(_AES_ENC_us13_n623 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n1125 ) );
NOR2_X2 _AES_ENC_us13_U239  ( .A1(_AES_ENC_us13_n990 ), .A2(_AES_ENC_us13_n929 ), .ZN(_AES_ENC_us13_n892 ) );
NOR2_X2 _AES_ENC_us13_U238  ( .A1(_AES_ENC_us13_n892 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n893 ) );
NOR2_X2 _AES_ENC_us13_U237  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n621 ), .ZN(_AES_ENC_us13_n950 ) );
NOR2_X2 _AES_ENC_us13_U236  ( .A1(_AES_ENC_us13_n1079 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n1082 ) );
NOR2_X2 _AES_ENC_us13_U235  ( .A1(_AES_ENC_us13_n910 ), .A2(_AES_ENC_us13_n1056 ), .ZN(_AES_ENC_us13_n941 ) );
NOR2_X2 _AES_ENC_us13_U234  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n1077 ), .ZN(_AES_ENC_us13_n841 ) );
NOR2_X2 _AES_ENC_us13_U229  ( .A1(_AES_ENC_us13_n601 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n630 ) );
NOR2_X2 _AES_ENC_us13_U228  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n621 ), .ZN(_AES_ENC_us13_n806 ) );
NOR2_X2 _AES_ENC_us13_U227  ( .A1(_AES_ENC_us13_n601 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n948 ) );
NOR2_X2 _AES_ENC_us13_U226  ( .A1(_AES_ENC_us13_n578 ), .A2(_AES_ENC_us13_n620 ), .ZN(_AES_ENC_us13_n997 ) );
NOR2_X2 _AES_ENC_us13_U225  ( .A1(_AES_ENC_us13_n1121 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n1122 ) );
NOR2_X2 _AES_ENC_us13_U223  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n1023 ), .ZN(_AES_ENC_us13_n756 ) );
NOR2_X2 _AES_ENC_us13_U222  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n621 ), .ZN(_AES_ENC_us13_n870 ) );
NOR2_X2 _AES_ENC_us13_U221  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n569 ), .ZN(_AES_ENC_us13_n947 ) );
NOR2_X2 _AES_ENC_us13_U217  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n1077 ), .ZN(_AES_ENC_us13_n1084 ) );
NOR2_X2 _AES_ENC_us13_U213  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n855 ), .ZN(_AES_ENC_us13_n709 ) );
NOR2_X2 _AES_ENC_us13_U212  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n620 ), .ZN(_AES_ENC_us13_n868 ) );
NOR2_X2 _AES_ENC_us13_U211  ( .A1(_AES_ENC_us13_n1120 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n1124 ) );
NOR2_X2 _AES_ENC_us13_U210  ( .A1(_AES_ENC_us13_n1120 ), .A2(_AES_ENC_us13_n839 ), .ZN(_AES_ENC_us13_n842 ) );
NOR2_X2 _AES_ENC_us13_U209  ( .A1(_AES_ENC_us13_n1120 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n696 ) );
NOR2_X2 _AES_ENC_us13_U208  ( .A1(_AES_ENC_us13_n1074 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n1076 ) );
NOR2_X2 _AES_ENC_us13_U207  ( .A1(_AES_ENC_us13_n1074 ), .A2(_AES_ENC_us13_n609 ), .ZN(_AES_ENC_us13_n781 ) );
NOR3_X2 _AES_ENC_us13_U201  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n1056 ), .A3(_AES_ENC_us13_n990 ), .ZN(_AES_ENC_us13_n979 ) );
NOR3_X2 _AES_ENC_us13_U200  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n1058 ), .A3(_AES_ENC_us13_n1059 ), .ZN(_AES_ENC_us13_n854 ) );
NOR2_X2 _AES_ENC_us13_U199  ( .A1(_AES_ENC_us13_n996 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n869 ) );
NOR2_X2 _AES_ENC_us13_U198  ( .A1(_AES_ENC_us13_n1056 ), .A2(_AES_ENC_us13_n1074 ), .ZN(_AES_ENC_us13_n1057 ) );
NOR3_X2 _AES_ENC_us13_U197  ( .A1(_AES_ENC_us13_n579 ), .A2(_AES_ENC_us13_n1120 ), .A3(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n978 ) );
NOR2_X2 _AES_ENC_us13_U196  ( .A1(_AES_ENC_us13_n996 ), .A2(_AES_ENC_us13_n911 ), .ZN(_AES_ENC_us13_n1116 ) );
NOR2_X2 _AES_ENC_us13_U195  ( .A1(_AES_ENC_us13_n1074 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n754 ) );
NOR2_X2 _AES_ENC_us13_U194  ( .A1(_AES_ENC_us13_n926 ), .A2(_AES_ENC_us13_n1103 ), .ZN(_AES_ENC_us13_n977 ) );
NOR2_X2 _AES_ENC_us13_U187  ( .A1(_AES_ENC_us13_n839 ), .A2(_AES_ENC_us13_n824 ), .ZN(_AES_ENC_us13_n1092 ) );
NOR2_X2 _AES_ENC_us13_U186  ( .A1(_AES_ENC_us13_n573 ), .A2(_AES_ENC_us13_n1074 ), .ZN(_AES_ENC_us13_n684 ) );
NOR2_X2 _AES_ENC_us13_U185  ( .A1(_AES_ENC_us13_n826 ), .A2(_AES_ENC_us13_n1059 ), .ZN(_AES_ENC_us13_n907 ) );
NOR3_X2 _AES_ENC_us13_U184  ( .A1(_AES_ENC_us13_n593 ), .A2(_AES_ENC_us13_n1115 ), .A3(_AES_ENC_us13_n600 ), .ZN(_AES_ENC_us13_n831 ) );
NOR3_X2 _AES_ENC_us13_U183  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n1056 ), .A3(_AES_ENC_us13_n990 ), .ZN(_AES_ENC_us13_n896 ) );
NOR3_X2 _AES_ENC_us13_U182  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n573 ), .A3(_AES_ENC_us13_n1013 ), .ZN(_AES_ENC_us13_n670 ) );
NOR3_X2 _AES_ENC_us13_U181  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n1091 ), .A3(_AES_ENC_us13_n1022 ), .ZN(_AES_ENC_us13_n843 ) );
NOR2_X2 _AES_ENC_us13_U180  ( .A1(_AES_ENC_us13_n1029 ), .A2(_AES_ENC_us13_n1095 ), .ZN(_AES_ENC_us13_n735 ) );
NOR2_X2 _AES_ENC_us13_U174  ( .A1(_AES_ENC_us13_n1100 ), .A2(_AES_ENC_us13_n854 ), .ZN(_AES_ENC_us13_n860 ) );
NAND3_X2 _AES_ENC_us13_U173  ( .A1(_AES_ENC_us13_n569 ), .A2(_AES_ENC_us13_n603 ), .A3(_AES_ENC_us13_n681 ), .ZN(_AES_ENC_us13_n691 ) );
NOR2_X2 _AES_ENC_us13_U172  ( .A1(_AES_ENC_us13_n683 ), .A2(_AES_ENC_us13_n682 ), .ZN(_AES_ENC_us13_n690 ) );
NOR3_X2 _AES_ENC_us13_U171  ( .A1(_AES_ENC_us13_n695 ), .A2(_AES_ENC_us13_n694 ), .A3(_AES_ENC_us13_n693 ), .ZN(_AES_ENC_us13_n700 ) );
NOR4_X2 _AES_ENC_us13_U170  ( .A1(_AES_ENC_us13_n983 ), .A2(_AES_ENC_us13_n698 ), .A3(_AES_ENC_us13_n697 ), .A4(_AES_ENC_us13_n696 ), .ZN(_AES_ENC_us13_n699 ) );
NOR2_X2 _AES_ENC_us13_U169  ( .A1(_AES_ENC_us13_n946 ), .A2(_AES_ENC_us13_n945 ), .ZN(_AES_ENC_us13_n952 ) );
NOR4_X2 _AES_ENC_us13_U168  ( .A1(_AES_ENC_us13_n950 ), .A2(_AES_ENC_us13_n949 ), .A3(_AES_ENC_us13_n948 ), .A4(_AES_ENC_us13_n947 ), .ZN(_AES_ENC_us13_n951 ) );
NOR4_X2 _AES_ENC_us13_U162  ( .A1(_AES_ENC_us13_n983 ), .A2(_AES_ENC_us13_n982 ), .A3(_AES_ENC_us13_n981 ), .A4(_AES_ENC_us13_n980 ), .ZN(_AES_ENC_us13_n984 ) );
NOR2_X2 _AES_ENC_us13_U161  ( .A1(_AES_ENC_us13_n979 ), .A2(_AES_ENC_us13_n978 ), .ZN(_AES_ENC_us13_n985 ) );
NOR4_X2 _AES_ENC_us13_U160  ( .A1(_AES_ENC_us13_n896 ), .A2(_AES_ENC_us13_n895 ), .A3(_AES_ENC_us13_n894 ), .A4(_AES_ENC_us13_n893 ), .ZN(_AES_ENC_us13_n897 ) );
NOR2_X2 _AES_ENC_us13_U159  ( .A1(_AES_ENC_us13_n866 ), .A2(_AES_ENC_us13_n865 ), .ZN(_AES_ENC_us13_n872 ) );
NOR4_X2 _AES_ENC_us13_U158  ( .A1(_AES_ENC_us13_n870 ), .A2(_AES_ENC_us13_n869 ), .A3(_AES_ENC_us13_n868 ), .A4(_AES_ENC_us13_n867 ), .ZN(_AES_ENC_us13_n871 ) );
NOR4_X2 _AES_ENC_us13_U157  ( .A1(_AES_ENC_us13_n1125 ), .A2(_AES_ENC_us13_n1124 ), .A3(_AES_ENC_us13_n1123 ), .A4(_AES_ENC_us13_n1122 ), .ZN(_AES_ENC_us13_n1126 ) );
NOR4_X2 _AES_ENC_us13_U156  ( .A1(_AES_ENC_us13_n1084 ), .A2(_AES_ENC_us13_n1083 ), .A3(_AES_ENC_us13_n1082 ), .A4(_AES_ENC_us13_n1081 ), .ZN(_AES_ENC_us13_n1085 ) );
NOR2_X2 _AES_ENC_us13_U155  ( .A1(_AES_ENC_us13_n1076 ), .A2(_AES_ENC_us13_n1075 ), .ZN(_AES_ENC_us13_n1086 ) );
NOR3_X2 _AES_ENC_us13_U154  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n1054 ), .A3(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n961 ) );
NOR3_X2 _AES_ENC_us13_U153  ( .A1(_AES_ENC_us13_n609 ), .A2(_AES_ENC_us13_n1074 ), .A3(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n671 ) );
NOR2_X2 _AES_ENC_us13_U152  ( .A1(_AES_ENC_us13_n1057 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n1062 ) );
NOR2_X2 _AES_ENC_us13_U143  ( .A1(_AES_ENC_us13_n1055 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n1063 ) );
NOR2_X2 _AES_ENC_us13_U142  ( .A1(_AES_ENC_us13_n1060 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n1061 ) );
NOR4_X2 _AES_ENC_us13_U141  ( .A1(_AES_ENC_us13_n1064 ), .A2(_AES_ENC_us13_n1063 ), .A3(_AES_ENC_us13_n1062 ), .A4(_AES_ENC_us13_n1061 ), .ZN(_AES_ENC_us13_n1065 ) );
NOR3_X2 _AES_ENC_us13_U140  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n1120 ), .A3(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n918 ) );
NOR3_X2 _AES_ENC_us13_U132  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n573 ), .A3(_AES_ENC_us13_n1013 ), .ZN(_AES_ENC_us13_n917 ) );
NOR2_X2 _AES_ENC_us13_U131  ( .A1(_AES_ENC_us13_n914 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n915 ) );
NOR4_X2 _AES_ENC_us13_U130  ( .A1(_AES_ENC_us13_n918 ), .A2(_AES_ENC_us13_n917 ), .A3(_AES_ENC_us13_n916 ), .A4(_AES_ENC_us13_n915 ), .ZN(_AES_ENC_us13_n919 ) );
NOR2_X2 _AES_ENC_us13_U129  ( .A1(_AES_ENC_us13_n590 ), .A2(_AES_ENC_us13_n599 ), .ZN(_AES_ENC_us13_n771 ) );
NOR2_X2 _AES_ENC_us13_U128  ( .A1(_AES_ENC_us13_n1103 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n772 ) );
NOR2_X2 _AES_ENC_us13_U127  ( .A1(_AES_ENC_us13_n583 ), .A2(_AES_ENC_us13_n615 ), .ZN(_AES_ENC_us13_n773 ) );
NOR4_X2 _AES_ENC_us13_U126  ( .A1(_AES_ENC_us13_n773 ), .A2(_AES_ENC_us13_n772 ), .A3(_AES_ENC_us13_n771 ), .A4(_AES_ENC_us13_n770 ), .ZN(_AES_ENC_us13_n774 ) );
NOR2_X2 _AES_ENC_us13_U121  ( .A1(_AES_ENC_us13_n735 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n687 ) );
NOR2_X2 _AES_ENC_us13_U120  ( .A1(_AES_ENC_us13_n684 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n688 ) );
NOR2_X2 _AES_ENC_us13_U119  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n622 ), .ZN(_AES_ENC_us13_n686 ) );
NOR4_X2 _AES_ENC_us13_U118  ( .A1(_AES_ENC_us13_n688 ), .A2(_AES_ENC_us13_n687 ), .A3(_AES_ENC_us13_n686 ), .A4(_AES_ENC_us13_n685 ), .ZN(_AES_ENC_us13_n689 ) );
NOR2_X2 _AES_ENC_us13_U117  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n608 ), .ZN(_AES_ENC_us13_n858 ) );
NOR2_X2 _AES_ENC_us13_U116  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n855 ), .ZN(_AES_ENC_us13_n857 ) );
NOR2_X2 _AES_ENC_us13_U115  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n617 ), .ZN(_AES_ENC_us13_n856 ) );
NOR4_X2 _AES_ENC_us13_U106  ( .A1(_AES_ENC_us13_n858 ), .A2(_AES_ENC_us13_n857 ), .A3(_AES_ENC_us13_n856 ), .A4(_AES_ENC_us13_n958 ), .ZN(_AES_ENC_us13_n859 ) );
NOR2_X2 _AES_ENC_us13_U105  ( .A1(_AES_ENC_us13_n780 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n784 ) );
NOR2_X2 _AES_ENC_us13_U104  ( .A1(_AES_ENC_us13_n1117 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n782 ) );
NOR2_X2 _AES_ENC_us13_U103  ( .A1(_AES_ENC_us13_n781 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n783 ) );
NOR4_X2 _AES_ENC_us13_U102  ( .A1(_AES_ENC_us13_n880 ), .A2(_AES_ENC_us13_n784 ), .A3(_AES_ENC_us13_n783 ), .A4(_AES_ENC_us13_n782 ), .ZN(_AES_ENC_us13_n785 ) );
NOR2_X2 _AES_ENC_us13_U101  ( .A1(_AES_ENC_us13_n597 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n814 ) );
NOR2_X2 _AES_ENC_us13_U100  ( .A1(_AES_ENC_us13_n907 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n813 ) );
NOR3_X2 _AES_ENC_us13_U95  ( .A1(_AES_ENC_us13_n578 ), .A2(_AES_ENC_us13_n1058 ), .A3(_AES_ENC_us13_n1059 ), .ZN(_AES_ENC_us13_n815 ) );
NOR4_X2 _AES_ENC_us13_U94  ( .A1(_AES_ENC_us13_n815 ), .A2(_AES_ENC_us13_n814 ), .A3(_AES_ENC_us13_n813 ), .A4(_AES_ENC_us13_n812 ), .ZN(_AES_ENC_us13_n816 ) );
NOR2_X2 _AES_ENC_us13_U93  ( .A1(_AES_ENC_us13_n591 ), .A2(_AES_ENC_us13_n569 ), .ZN(_AES_ENC_us13_n721 ) );
NOR2_X2 _AES_ENC_us13_U92  ( .A1(_AES_ENC_us13_n1031 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n723 ) );
NOR2_X2 _AES_ENC_us13_U91  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n1096 ), .ZN(_AES_ENC_us13_n722 ) );
NOR4_X2 _AES_ENC_us13_U90  ( .A1(_AES_ENC_us13_n724 ), .A2(_AES_ENC_us13_n723 ), .A3(_AES_ENC_us13_n722 ), .A4(_AES_ENC_us13_n721 ), .ZN(_AES_ENC_us13_n725 ) );
NOR2_X2 _AES_ENC_us13_U89  ( .A1(_AES_ENC_us13_n911 ), .A2(_AES_ENC_us13_n990 ), .ZN(_AES_ENC_us13_n1009 ) );
NOR2_X2 _AES_ENC_us13_U88  ( .A1(_AES_ENC_us13_n1013 ), .A2(_AES_ENC_us13_n573 ), .ZN(_AES_ENC_us13_n1014 ) );
NOR2_X2 _AES_ENC_us13_U87  ( .A1(_AES_ENC_us13_n1014 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n1015 ) );
NOR4_X2 _AES_ENC_us13_U86  ( .A1(_AES_ENC_us13_n1016 ), .A2(_AES_ENC_us13_n1015 ), .A3(_AES_ENC_us13_n1119 ), .A4(_AES_ENC_us13_n1046 ), .ZN(_AES_ENC_us13_n1017 ) );
NOR2_X2 _AES_ENC_us13_U81  ( .A1(_AES_ENC_us13_n996 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n998 ) );
NOR2_X2 _AES_ENC_us13_U80  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n618 ), .ZN(_AES_ENC_us13_n1000 ) );
NOR2_X2 _AES_ENC_us13_U79  ( .A1(_AES_ENC_us13_n590 ), .A2(_AES_ENC_us13_n1096 ), .ZN(_AES_ENC_us13_n999 ) );
NOR4_X2 _AES_ENC_us13_U78  ( .A1(_AES_ENC_us13_n1000 ), .A2(_AES_ENC_us13_n999 ), .A3(_AES_ENC_us13_n998 ), .A4(_AES_ENC_us13_n997 ), .ZN(_AES_ENC_us13_n1001 ) );
NOR2_X2 _AES_ENC_us13_U74  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n1096 ), .ZN(_AES_ENC_us13_n697 ) );
NOR2_X2 _AES_ENC_us13_U73  ( .A1(_AES_ENC_us13_n609 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n958 ) );
NOR2_X2 _AES_ENC_us13_U72  ( .A1(_AES_ENC_us13_n911 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n983 ) );
NOR2_X2 _AES_ENC_us13_U71  ( .A1(_AES_ENC_us13_n1054 ), .A2(_AES_ENC_us13_n1103 ), .ZN(_AES_ENC_us13_n1031 ) );
INV_X4 _AES_ENC_us13_U65  ( .A(_AES_ENC_us13_n1050 ), .ZN(_AES_ENC_us13_n585 ) );
INV_X4 _AES_ENC_us13_U64  ( .A(_AES_ENC_us13_n1072 ), .ZN(_AES_ENC_us13_n577 ) );
INV_X4 _AES_ENC_us13_U63  ( .A(_AES_ENC_us13_n1073 ), .ZN(_AES_ENC_us13_n576 ) );
NOR2_X2 _AES_ENC_us13_U62  ( .A1(_AES_ENC_us13_n603 ), .A2(_AES_ENC_us13_n587 ), .ZN(_AES_ENC_us13_n880 ) );
NOR3_X2 _AES_ENC_us13_U61  ( .A1(_AES_ENC_us13_n826 ), .A2(_AES_ENC_us13_n1121 ), .A3(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n946 ) );
INV_X4 _AES_ENC_us13_U59  ( .A(_AES_ENC_us13_n1010 ), .ZN(_AES_ENC_us13_n581 ) );
NOR3_X2 _AES_ENC_us13_U58  ( .A1(_AES_ENC_us13_n573 ), .A2(_AES_ENC_us13_n1029 ), .A3(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n1119 ) );
INV_X4 _AES_ENC_us13_U57  ( .A(_AES_ENC_us13_n956 ), .ZN(_AES_ENC_us13_n589 ) );
NOR2_X2 _AES_ENC_us13_U50  ( .A1(_AES_ENC_us13_n601 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n1013 ) );
NOR2_X2 _AES_ENC_us13_U49  ( .A1(_AES_ENC_us13_n609 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n910 ) );
NOR2_X2 _AES_ENC_us13_U48  ( .A1(_AES_ENC_us13_n569 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n1091 ) );
NOR2_X2 _AES_ENC_us13_U47  ( .A1(_AES_ENC_us13_n614 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n990 ) );
NOR2_X2 _AES_ENC_us13_U46  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_us13_n1121 ), .ZN(_AES_ENC_us13_n996 ) );
NOR2_X2 _AES_ENC_us13_U45  ( .A1(_AES_ENC_us13_n583 ), .A2(_AES_ENC_us13_n622 ), .ZN(_AES_ENC_us13_n628 ) );
NOR2_X2 _AES_ENC_us13_U44  ( .A1(_AES_ENC_us13_n602 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n866 ) );
NOR2_X2 _AES_ENC_us13_U43  ( .A1(_AES_ENC_us13_n610 ), .A2(_AES_ENC_us13_n583 ), .ZN(_AES_ENC_us13_n1006 ) );
NOR2_X2 _AES_ENC_us13_U42  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n1117 ), .ZN(_AES_ENC_us13_n1118 ) );
NOR2_X2 _AES_ENC_us13_U41  ( .A1(_AES_ENC_us13_n1119 ), .A2(_AES_ENC_us13_n1118 ), .ZN(_AES_ENC_us13_n1127 ) );
NOR2_X2 _AES_ENC_us13_U36  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n616 ), .ZN(_AES_ENC_us13_n629 ) );
NOR2_X2 _AES_ENC_us13_U35  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n906 ), .ZN(_AES_ENC_us13_n909 ) );
NOR2_X2 _AES_ENC_us13_U34  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n607 ), .ZN(_AES_ENC_us13_n658 ) );
NOR2_X2 _AES_ENC_us13_U33  ( .A1(_AES_ENC_us13_n1116 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n695 ) );
NOR2_X2 _AES_ENC_us13_U32  ( .A1(_AES_ENC_us13_n1078 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n1083 ) );
NOR2_X2 _AES_ENC_us13_U31  ( .A1(_AES_ENC_us13_n941 ), .A2(_AES_ENC_us13_n581 ), .ZN(_AES_ENC_us13_n724 ) );
NOR2_X2 _AES_ENC_us13_U30  ( .A1(_AES_ENC_us13_n611 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n1107 ) );
NOR2_X2 _AES_ENC_us13_U29  ( .A1(_AES_ENC_us13_n602 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n840 ) );
NOR2_X2 _AES_ENC_us13_U24  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n623 ), .ZN(_AES_ENC_us13_n633 ) );
NOR2_X2 _AES_ENC_us13_U23  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n1080 ), .ZN(_AES_ENC_us13_n1081 ) );
NOR2_X2 _AES_ENC_us13_U21  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n1045 ), .ZN(_AES_ENC_us13_n812 ) );
NOR2_X2 _AES_ENC_us13_U20  ( .A1(_AES_ENC_us13_n1009 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n960 ) );
NOR2_X2 _AES_ENC_us13_U19  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n619 ), .ZN(_AES_ENC_us13_n982 ) );
NOR2_X2 _AES_ENC_us13_U18  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n616 ), .ZN(_AES_ENC_us13_n757 ) );
NOR2_X2 _AES_ENC_us13_U17  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n598 ), .ZN(_AES_ENC_us13_n698 ) );
NOR2_X2 _AES_ENC_us13_U16  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n605 ), .ZN(_AES_ENC_us13_n708 ) );
NOR2_X2 _AES_ENC_us13_U15  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n603 ), .ZN(_AES_ENC_us13_n770 ) );
NOR2_X2 _AES_ENC_us13_U10  ( .A1(_AES_ENC_us13_n605 ), .A2(_AES_ENC_us13_n576 ), .ZN(_AES_ENC_us13_n803 ) );
NOR2_X2 _AES_ENC_us13_U9  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n881 ), .ZN(_AES_ENC_us13_n711 ) );
NOR2_X2 _AES_ENC_us13_U8  ( .A1(_AES_ENC_us13_n589 ), .A2(_AES_ENC_us13_n603 ), .ZN(_AES_ENC_us13_n867 ) );
NOR2_X2 _AES_ENC_us13_U7  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n615 ), .ZN(_AES_ENC_us13_n804 ) );
NOR2_X2 _AES_ENC_us13_U6  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n609 ), .ZN(_AES_ENC_us13_n1046 ) );
OR2_X4 _AES_ENC_us13_U5  ( .A1(_AES_ENC_us13_n612 ), .A2(_AES_ENC_sa13[1]),.ZN(_AES_ENC_us13_n570 ) );
OR2_X4 _AES_ENC_us13_U4  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_sa13[4]),.ZN(_AES_ENC_us13_n569 ) );
NAND2_X2 _AES_ENC_us13_U514  ( .A1(_AES_ENC_us13_n1121 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n1030 ) );
AND2_X2 _AES_ENC_us13_U513  ( .A1(_AES_ENC_us13_n607 ), .A2(_AES_ENC_us13_n1030 ), .ZN(_AES_ENC_us13_n1049 ) );
NAND2_X2 _AES_ENC_us13_U511  ( .A1(_AES_ENC_us13_n1049 ), .A2(_AES_ENC_us13_n794 ), .ZN(_AES_ENC_us13_n637 ) );
AND2_X2 _AES_ENC_us13_U493  ( .A1(_AES_ENC_us13_n779 ), .A2(_AES_ENC_us13_n996 ), .ZN(_AES_ENC_us13_n632 ) );
NAND4_X2 _AES_ENC_us13_U485  ( .A1(_AES_ENC_us13_n637 ), .A2(_AES_ENC_us13_n636 ), .A3(_AES_ENC_us13_n635 ), .A4(_AES_ENC_us13_n634 ), .ZN(_AES_ENC_us13_n638 ) );
NAND2_X2 _AES_ENC_us13_U484  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n638 ), .ZN(_AES_ENC_us13_n679 ) );
NAND2_X2 _AES_ENC_us13_U481  ( .A1(_AES_ENC_us13_n1094 ), .A2(_AES_ENC_us13_n613 ), .ZN(_AES_ENC_us13_n648 ) );
NAND2_X2 _AES_ENC_us13_U476  ( .A1(_AES_ENC_us13_n619 ), .A2(_AES_ENC_us13_n598 ), .ZN(_AES_ENC_us13_n762 ) );
NAND2_X2 _AES_ENC_us13_U475  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n762 ), .ZN(_AES_ENC_us13_n647 ) );
NAND4_X2 _AES_ENC_us13_U457  ( .A1(_AES_ENC_us13_n648 ), .A2(_AES_ENC_us13_n647 ), .A3(_AES_ENC_us13_n646 ), .A4(_AES_ENC_us13_n645 ), .ZN(_AES_ENC_us13_n649 ) );
NAND2_X2 _AES_ENC_us13_U456  ( .A1(_AES_ENC_sa13[0]), .A2(_AES_ENC_us13_n649 ), .ZN(_AES_ENC_us13_n665 ) );
NAND2_X2 _AES_ENC_us13_U454  ( .A1(_AES_ENC_us13_n626 ), .A2(_AES_ENC_us13_n601 ), .ZN(_AES_ENC_us13_n855 ) );
NAND2_X2 _AES_ENC_us13_U453  ( .A1(_AES_ENC_us13_n617 ), .A2(_AES_ENC_us13_n855 ), .ZN(_AES_ENC_us13_n821 ) );
NAND2_X2 _AES_ENC_us13_U452  ( .A1(_AES_ENC_us13_n1093 ), .A2(_AES_ENC_us13_n821 ), .ZN(_AES_ENC_us13_n662 ) );
NAND2_X2 _AES_ENC_us13_U451  ( .A1(_AES_ENC_us13_n605 ), .A2(_AES_ENC_us13_n620 ), .ZN(_AES_ENC_us13_n650 ) );
NAND2_X2 _AES_ENC_us13_U450  ( .A1(_AES_ENC_us13_n956 ), .A2(_AES_ENC_us13_n650 ), .ZN(_AES_ENC_us13_n661 ) );
NAND2_X2 _AES_ENC_us13_U449  ( .A1(_AES_ENC_us13_n594 ), .A2(_AES_ENC_us13_n595 ), .ZN(_AES_ENC_us13_n839 ) );
OR2_X2 _AES_ENC_us13_U446  ( .A1(_AES_ENC_us13_n839 ), .A2(_AES_ENC_us13_n932 ), .ZN(_AES_ENC_us13_n656 ) );
NAND2_X2 _AES_ENC_us13_U445  ( .A1(_AES_ENC_us13_n624 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n1096 ) );
NAND2_X2 _AES_ENC_us13_U444  ( .A1(_AES_ENC_us13_n1030 ), .A2(_AES_ENC_us13_n1096 ), .ZN(_AES_ENC_us13_n651 ) );
NAND2_X2 _AES_ENC_us13_U443  ( .A1(_AES_ENC_us13_n1114 ), .A2(_AES_ENC_us13_n651 ), .ZN(_AES_ENC_us13_n655 ) );
OR3_X2 _AES_ENC_us13_U440  ( .A1(_AES_ENC_us13_n1079 ), .A2(_AES_ENC_sa13[7]), .A3(_AES_ENC_us13_n594 ), .ZN(_AES_ENC_us13_n654 ));
NAND2_X2 _AES_ENC_us13_U439  ( .A1(_AES_ENC_us13_n623 ), .A2(_AES_ENC_us13_n619 ), .ZN(_AES_ENC_us13_n652 ) );
NAND4_X2 _AES_ENC_us13_U437  ( .A1(_AES_ENC_us13_n656 ), .A2(_AES_ENC_us13_n655 ), .A3(_AES_ENC_us13_n654 ), .A4(_AES_ENC_us13_n653 ), .ZN(_AES_ENC_us13_n657 ) );
NAND2_X2 _AES_ENC_us13_U436  ( .A1(_AES_ENC_sa13[2]), .A2(_AES_ENC_us13_n657 ), .ZN(_AES_ENC_us13_n660 ) );
NAND4_X2 _AES_ENC_us13_U432  ( .A1(_AES_ENC_us13_n662 ), .A2(_AES_ENC_us13_n661 ), .A3(_AES_ENC_us13_n660 ), .A4(_AES_ENC_us13_n659 ), .ZN(_AES_ENC_us13_n663 ) );
NAND2_X2 _AES_ENC_us13_U431  ( .A1(_AES_ENC_us13_n663 ), .A2(_AES_ENC_us13_n627 ), .ZN(_AES_ENC_us13_n664 ) );
NAND2_X2 _AES_ENC_us13_U430  ( .A1(_AES_ENC_us13_n665 ), .A2(_AES_ENC_us13_n664 ), .ZN(_AES_ENC_us13_n666 ) );
NAND2_X2 _AES_ENC_us13_U429  ( .A1(_AES_ENC_sa13[6]), .A2(_AES_ENC_us13_n666 ), .ZN(_AES_ENC_us13_n678 ) );
NAND2_X2 _AES_ENC_us13_U426  ( .A1(_AES_ENC_us13_n735 ), .A2(_AES_ENC_us13_n1093 ), .ZN(_AES_ENC_us13_n675 ) );
NAND2_X2 _AES_ENC_us13_U425  ( .A1(_AES_ENC_us13_n625 ), .A2(_AES_ENC_us13_n607 ), .ZN(_AES_ENC_us13_n1045 ) );
OR2_X2 _AES_ENC_us13_U424  ( .A1(_AES_ENC_us13_n1045 ), .A2(_AES_ENC_us13_n577 ), .ZN(_AES_ENC_us13_n674 ) );
NAND2_X2 _AES_ENC_us13_U423  ( .A1(_AES_ENC_sa13[1]), .A2(_AES_ENC_us13_n609 ), .ZN(_AES_ENC_us13_n667 ) );
NAND2_X2 _AES_ENC_us13_U422  ( .A1(_AES_ENC_us13_n605 ), .A2(_AES_ENC_us13_n667 ), .ZN(_AES_ENC_us13_n1071 ) );
NAND4_X2 _AES_ENC_us13_U412  ( .A1(_AES_ENC_us13_n675 ), .A2(_AES_ENC_us13_n674 ), .A3(_AES_ENC_us13_n673 ), .A4(_AES_ENC_us13_n672 ), .ZN(_AES_ENC_us13_n676 ) );
NAND2_X2 _AES_ENC_us13_U411  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n676 ), .ZN(_AES_ENC_us13_n677 ) );
NAND2_X2 _AES_ENC_us13_U408  ( .A1(_AES_ENC_us13_n800 ), .A2(_AES_ENC_us13_n1022 ), .ZN(_AES_ENC_us13_n680 ) );
NAND2_X2 _AES_ENC_us13_U407  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n680 ), .ZN(_AES_ENC_us13_n681 ) );
AND2_X2 _AES_ENC_us13_U402  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n684 ), .ZN(_AES_ENC_us13_n682 ) );
NAND4_X2 _AES_ENC_us13_U395  ( .A1(_AES_ENC_us13_n691 ), .A2(_AES_ENC_us13_n586 ), .A3(_AES_ENC_us13_n690 ), .A4(_AES_ENC_us13_n689 ), .ZN(_AES_ENC_us13_n692 ) );
NAND2_X2 _AES_ENC_us13_U394  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n692 ), .ZN(_AES_ENC_us13_n733 ) );
NAND2_X2 _AES_ENC_us13_U392  ( .A1(_AES_ENC_us13_n977 ), .A2(_AES_ENC_us13_n1050 ), .ZN(_AES_ENC_us13_n702 ) );
NAND2_X2 _AES_ENC_us13_U391  ( .A1(_AES_ENC_us13_n1093 ), .A2(_AES_ENC_us13_n1045 ), .ZN(_AES_ENC_us13_n701 ) );
NAND4_X2 _AES_ENC_us13_U381  ( .A1(_AES_ENC_us13_n702 ), .A2(_AES_ENC_us13_n701 ), .A3(_AES_ENC_us13_n700 ), .A4(_AES_ENC_us13_n699 ), .ZN(_AES_ENC_us13_n703 ) );
NAND2_X2 _AES_ENC_us13_U380  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n703 ), .ZN(_AES_ENC_us13_n732 ) );
AND2_X2 _AES_ENC_us13_U379  ( .A1(_AES_ENC_sa13[0]), .A2(_AES_ENC_sa13[6]),.ZN(_AES_ENC_us13_n1113 ) );
NAND2_X2 _AES_ENC_us13_U378  ( .A1(_AES_ENC_us13_n619 ), .A2(_AES_ENC_us13_n1030 ), .ZN(_AES_ENC_us13_n881 ) );
NAND2_X2 _AES_ENC_us13_U377  ( .A1(_AES_ENC_us13_n1093 ), .A2(_AES_ENC_us13_n881 ), .ZN(_AES_ENC_us13_n715 ) );
NAND2_X2 _AES_ENC_us13_U376  ( .A1(_AES_ENC_us13_n1010 ), .A2(_AES_ENC_us13_n622 ), .ZN(_AES_ENC_us13_n714 ) );
NAND2_X2 _AES_ENC_us13_U375  ( .A1(_AES_ENC_us13_n855 ), .A2(_AES_ENC_us13_n625 ), .ZN(_AES_ENC_us13_n1117 ) );
XNOR2_X2 _AES_ENC_us13_U371  ( .A(_AES_ENC_us13_n584 ), .B(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n824 ) );
NAND4_X2 _AES_ENC_us13_U362  ( .A1(_AES_ENC_us13_n715 ), .A2(_AES_ENC_us13_n714 ), .A3(_AES_ENC_us13_n713 ), .A4(_AES_ENC_us13_n712 ), .ZN(_AES_ENC_us13_n716 ) );
NAND2_X2 _AES_ENC_us13_U361  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n716 ), .ZN(_AES_ENC_us13_n731 ) );
AND2_X2 _AES_ENC_us13_U360  ( .A1(_AES_ENC_sa13[6]), .A2(_AES_ENC_us13_n627 ), .ZN(_AES_ENC_us13_n1131 ) );
NAND2_X2 _AES_ENC_us13_U359  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n717 ) );
NAND2_X2 _AES_ENC_us13_U358  ( .A1(_AES_ENC_us13_n1029 ), .A2(_AES_ENC_us13_n717 ), .ZN(_AES_ENC_us13_n728 ) );
NAND2_X2 _AES_ENC_us13_U357  ( .A1(_AES_ENC_sa13[1]), .A2(_AES_ENC_us13_n612 ), .ZN(_AES_ENC_us13_n1097 ) );
NAND2_X2 _AES_ENC_us13_U356  ( .A1(_AES_ENC_us13_n610 ), .A2(_AES_ENC_us13_n1097 ), .ZN(_AES_ENC_us13_n718 ) );
NAND2_X2 _AES_ENC_us13_U355  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n718 ), .ZN(_AES_ENC_us13_n727 ) );
NAND4_X2 _AES_ENC_us13_U344  ( .A1(_AES_ENC_us13_n728 ), .A2(_AES_ENC_us13_n727 ), .A3(_AES_ENC_us13_n726 ), .A4(_AES_ENC_us13_n725 ), .ZN(_AES_ENC_us13_n729 ) );
NAND2_X2 _AES_ENC_us13_U343  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n729 ), .ZN(_AES_ENC_us13_n730 ) );
NAND4_X2 _AES_ENC_us13_U342  ( .A1(_AES_ENC_us13_n733 ), .A2(_AES_ENC_us13_n732 ), .A3(_AES_ENC_us13_n731 ), .A4(_AES_ENC_us13_n730 ), .ZN(_AES_ENC_sa13_sub[1] ) );
NAND2_X2 _AES_ENC_us13_U341  ( .A1(_AES_ENC_sa13[7]), .A2(_AES_ENC_us13_n584 ), .ZN(_AES_ENC_us13_n734 ) );
NAND2_X2 _AES_ENC_us13_U340  ( .A1(_AES_ENC_us13_n734 ), .A2(_AES_ENC_us13_n579 ), .ZN(_AES_ENC_us13_n738 ) );
OR4_X2 _AES_ENC_us13_U339  ( .A1(_AES_ENC_us13_n738 ), .A2(_AES_ENC_us13_n594 ), .A3(_AES_ENC_us13_n826 ), .A4(_AES_ENC_us13_n1121 ), .ZN(_AES_ENC_us13_n746 ) );
NAND2_X2 _AES_ENC_us13_U337  ( .A1(_AES_ENC_us13_n1100 ), .A2(_AES_ENC_us13_n617 ), .ZN(_AES_ENC_us13_n992 ) );
OR2_X2 _AES_ENC_us13_U336  ( .A1(_AES_ENC_us13_n583 ), .A2(_AES_ENC_us13_n735 ), .ZN(_AES_ENC_us13_n737 ) );
NAND2_X2 _AES_ENC_us13_U334  ( .A1(_AES_ENC_us13_n605 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n753 ) );
NAND2_X2 _AES_ENC_us13_U333  ( .A1(_AES_ENC_us13_n603 ), .A2(_AES_ENC_us13_n753 ), .ZN(_AES_ENC_us13_n1080 ) );
NAND2_X2 _AES_ENC_us13_U332  ( .A1(_AES_ENC_us13_n1048 ), .A2(_AES_ENC_us13_n602 ), .ZN(_AES_ENC_us13_n736 ) );
NAND2_X2 _AES_ENC_us13_U331  ( .A1(_AES_ENC_us13_n737 ), .A2(_AES_ENC_us13_n736 ), .ZN(_AES_ENC_us13_n739 ) );
NAND2_X2 _AES_ENC_us13_U330  ( .A1(_AES_ENC_us13_n739 ), .A2(_AES_ENC_us13_n738 ), .ZN(_AES_ENC_us13_n745 ) );
NAND2_X2 _AES_ENC_us13_U326  ( .A1(_AES_ENC_us13_n1096 ), .A2(_AES_ENC_us13_n598 ), .ZN(_AES_ENC_us13_n906 ) );
NAND4_X2 _AES_ENC_us13_U323  ( .A1(_AES_ENC_us13_n746 ), .A2(_AES_ENC_us13_n992 ), .A3(_AES_ENC_us13_n745 ), .A4(_AES_ENC_us13_n744 ), .ZN(_AES_ENC_us13_n747 ) );
NAND2_X2 _AES_ENC_us13_U322  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n747 ), .ZN(_AES_ENC_us13_n793 ) );
NAND2_X2 _AES_ENC_us13_U321  ( .A1(_AES_ENC_us13_n606 ), .A2(_AES_ENC_us13_n855 ), .ZN(_AES_ENC_us13_n748 ) );
NAND2_X2 _AES_ENC_us13_U320  ( .A1(_AES_ENC_us13_n956 ), .A2(_AES_ENC_us13_n748 ), .ZN(_AES_ENC_us13_n760 ) );
NAND2_X2 _AES_ENC_us13_U313  ( .A1(_AES_ENC_us13_n598 ), .A2(_AES_ENC_us13_n753 ), .ZN(_AES_ENC_us13_n1023 ) );
NAND4_X2 _AES_ENC_us13_U308  ( .A1(_AES_ENC_us13_n760 ), .A2(_AES_ENC_us13_n992 ), .A3(_AES_ENC_us13_n759 ), .A4(_AES_ENC_us13_n758 ), .ZN(_AES_ENC_us13_n761 ) );
NAND2_X2 _AES_ENC_us13_U307  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n761 ), .ZN(_AES_ENC_us13_n792 ) );
NAND2_X2 _AES_ENC_us13_U306  ( .A1(_AES_ENC_us13_n606 ), .A2(_AES_ENC_us13_n610 ), .ZN(_AES_ENC_us13_n989 ) );
NAND2_X2 _AES_ENC_us13_U305  ( .A1(_AES_ENC_us13_n1050 ), .A2(_AES_ENC_us13_n989 ), .ZN(_AES_ENC_us13_n777 ) );
NAND2_X2 _AES_ENC_us13_U304  ( .A1(_AES_ENC_us13_n1093 ), .A2(_AES_ENC_us13_n762 ), .ZN(_AES_ENC_us13_n776 ) );
XNOR2_X2 _AES_ENC_us13_U301  ( .A(_AES_ENC_sa13[7]), .B(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n959 ) );
NAND4_X2 _AES_ENC_us13_U289  ( .A1(_AES_ENC_us13_n777 ), .A2(_AES_ENC_us13_n776 ), .A3(_AES_ENC_us13_n775 ), .A4(_AES_ENC_us13_n774 ), .ZN(_AES_ENC_us13_n778 ) );
NAND2_X2 _AES_ENC_us13_U288  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n778 ), .ZN(_AES_ENC_us13_n791 ) );
NAND2_X2 _AES_ENC_us13_U287  ( .A1(_AES_ENC_us13_n1056 ), .A2(_AES_ENC_us13_n1050 ), .ZN(_AES_ENC_us13_n788 ) );
NAND2_X2 _AES_ENC_us13_U286  ( .A1(_AES_ENC_us13_n1091 ), .A2(_AES_ENC_us13_n779 ), .ZN(_AES_ENC_us13_n787 ) );
NAND2_X2 _AES_ENC_us13_U285  ( .A1(_AES_ENC_us13_n956 ), .A2(_AES_ENC_sa13[1]), .ZN(_AES_ENC_us13_n786 ) );
NAND4_X2 _AES_ENC_us13_U278  ( .A1(_AES_ENC_us13_n788 ), .A2(_AES_ENC_us13_n787 ), .A3(_AES_ENC_us13_n786 ), .A4(_AES_ENC_us13_n785 ), .ZN(_AES_ENC_us13_n789 ) );
NAND2_X2 _AES_ENC_us13_U277  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n789 ), .ZN(_AES_ENC_us13_n790 ) );
NAND4_X2 _AES_ENC_us13_U276  ( .A1(_AES_ENC_us13_n793 ), .A2(_AES_ENC_us13_n792 ), .A3(_AES_ENC_us13_n791 ), .A4(_AES_ENC_us13_n790 ), .ZN(_AES_ENC_sa13_sub[2] ) );
NAND2_X2 _AES_ENC_us13_U275  ( .A1(_AES_ENC_us13_n1059 ), .A2(_AES_ENC_us13_n794 ), .ZN(_AES_ENC_us13_n810 ) );
NAND2_X2 _AES_ENC_us13_U274  ( .A1(_AES_ENC_us13_n1049 ), .A2(_AES_ENC_us13_n956 ), .ZN(_AES_ENC_us13_n809 ) );
OR2_X2 _AES_ENC_us13_U266  ( .A1(_AES_ENC_us13_n1096 ), .A2(_AES_ENC_us13_n578 ), .ZN(_AES_ENC_us13_n802 ) );
NAND2_X2 _AES_ENC_us13_U265  ( .A1(_AES_ENC_us13_n1053 ), .A2(_AES_ENC_us13_n800 ), .ZN(_AES_ENC_us13_n801 ) );
NAND2_X2 _AES_ENC_us13_U264  ( .A1(_AES_ENC_us13_n802 ), .A2(_AES_ENC_us13_n801 ), .ZN(_AES_ENC_us13_n805 ) );
NAND4_X2 _AES_ENC_us13_U261  ( .A1(_AES_ENC_us13_n810 ), .A2(_AES_ENC_us13_n809 ), .A3(_AES_ENC_us13_n808 ), .A4(_AES_ENC_us13_n807 ), .ZN(_AES_ENC_us13_n811 ) );
NAND2_X2 _AES_ENC_us13_U260  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n811 ), .ZN(_AES_ENC_us13_n852 ) );
OR2_X2 _AES_ENC_us13_U259  ( .A1(_AES_ENC_us13_n1023 ), .A2(_AES_ENC_us13_n591 ), .ZN(_AES_ENC_us13_n819 ) );
OR2_X2 _AES_ENC_us13_U257  ( .A1(_AES_ENC_us13_n570 ), .A2(_AES_ENC_us13_n930 ), .ZN(_AES_ENC_us13_n818 ) );
NAND2_X2 _AES_ENC_us13_U256  ( .A1(_AES_ENC_us13_n1013 ), .A2(_AES_ENC_us13_n1094 ), .ZN(_AES_ENC_us13_n817 ) );
NAND4_X2 _AES_ENC_us13_U249  ( .A1(_AES_ENC_us13_n819 ), .A2(_AES_ENC_us13_n818 ), .A3(_AES_ENC_us13_n817 ), .A4(_AES_ENC_us13_n816 ), .ZN(_AES_ENC_us13_n820 ) );
NAND2_X2 _AES_ENC_us13_U248  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n820 ), .ZN(_AES_ENC_us13_n851 ) );
NAND2_X2 _AES_ENC_us13_U247  ( .A1(_AES_ENC_us13_n956 ), .A2(_AES_ENC_us13_n1080 ), .ZN(_AES_ENC_us13_n835 ) );
NAND2_X2 _AES_ENC_us13_U246  ( .A1(_AES_ENC_us13_n570 ), .A2(_AES_ENC_us13_n1030 ), .ZN(_AES_ENC_us13_n1047 ) );
OR2_X2 _AES_ENC_us13_U245  ( .A1(_AES_ENC_us13_n1047 ), .A2(_AES_ENC_us13_n585 ), .ZN(_AES_ENC_us13_n834 ) );
NAND2_X2 _AES_ENC_us13_U244  ( .A1(_AES_ENC_us13_n1072 ), .A2(_AES_ENC_us13_n620 ), .ZN(_AES_ENC_us13_n833 ) );
NAND4_X2 _AES_ENC_us13_U233  ( .A1(_AES_ENC_us13_n835 ), .A2(_AES_ENC_us13_n834 ), .A3(_AES_ENC_us13_n833 ), .A4(_AES_ENC_us13_n832 ), .ZN(_AES_ENC_us13_n836 ) );
NAND2_X2 _AES_ENC_us13_U232  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n836 ), .ZN(_AES_ENC_us13_n850 ) );
NAND2_X2 _AES_ENC_us13_U231  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n601 ), .ZN(_AES_ENC_us13_n847 ) );
NAND2_X2 _AES_ENC_us13_U230  ( .A1(_AES_ENC_us13_n1050 ), .A2(_AES_ENC_us13_n1071 ), .ZN(_AES_ENC_us13_n846 ) );
OR2_X2 _AES_ENC_us13_U224  ( .A1(_AES_ENC_us13_n1053 ), .A2(_AES_ENC_us13_n911 ), .ZN(_AES_ENC_us13_n1077 ) );
NAND4_X2 _AES_ENC_us13_U220  ( .A1(_AES_ENC_us13_n847 ), .A2(_AES_ENC_us13_n846 ), .A3(_AES_ENC_us13_n845 ), .A4(_AES_ENC_us13_n844 ), .ZN(_AES_ENC_us13_n848 ) );
NAND2_X2 _AES_ENC_us13_U219  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n848 ), .ZN(_AES_ENC_us13_n849 ) );
NAND4_X2 _AES_ENC_us13_U218  ( .A1(_AES_ENC_us13_n852 ), .A2(_AES_ENC_us13_n851 ), .A3(_AES_ENC_us13_n850 ), .A4(_AES_ENC_us13_n849 ), .ZN(_AES_ENC_sa13_sub[3] ) );
NAND2_X2 _AES_ENC_us13_U216  ( .A1(_AES_ENC_us13_n1009 ), .A2(_AES_ENC_us13_n1072 ), .ZN(_AES_ENC_us13_n862 ) );
NAND2_X2 _AES_ENC_us13_U215  ( .A1(_AES_ENC_us13_n610 ), .A2(_AES_ENC_us13_n618 ), .ZN(_AES_ENC_us13_n853 ) );
NAND2_X2 _AES_ENC_us13_U214  ( .A1(_AES_ENC_us13_n1050 ), .A2(_AES_ENC_us13_n853 ), .ZN(_AES_ENC_us13_n861 ) );
NAND4_X2 _AES_ENC_us13_U206  ( .A1(_AES_ENC_us13_n862 ), .A2(_AES_ENC_us13_n861 ), .A3(_AES_ENC_us13_n860 ), .A4(_AES_ENC_us13_n859 ), .ZN(_AES_ENC_us13_n863 ) );
NAND2_X2 _AES_ENC_us13_U205  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n863 ), .ZN(_AES_ENC_us13_n905 ) );
NAND2_X2 _AES_ENC_us13_U204  ( .A1(_AES_ENC_us13_n1010 ), .A2(_AES_ENC_us13_n989 ), .ZN(_AES_ENC_us13_n874 ) );
NAND2_X2 _AES_ENC_us13_U203  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n583 ), .ZN(_AES_ENC_us13_n864 ) );
NAND2_X2 _AES_ENC_us13_U202  ( .A1(_AES_ENC_us13_n929 ), .A2(_AES_ENC_us13_n864 ), .ZN(_AES_ENC_us13_n873 ) );
NAND4_X2 _AES_ENC_us13_U193  ( .A1(_AES_ENC_us13_n874 ), .A2(_AES_ENC_us13_n873 ), .A3(_AES_ENC_us13_n872 ), .A4(_AES_ENC_us13_n871 ), .ZN(_AES_ENC_us13_n875 ) );
NAND2_X2 _AES_ENC_us13_U192  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n875 ), .ZN(_AES_ENC_us13_n904 ) );
NAND2_X2 _AES_ENC_us13_U191  ( .A1(_AES_ENC_us13_n597 ), .A2(_AES_ENC_us13_n1050 ), .ZN(_AES_ENC_us13_n889 ) );
NAND2_X2 _AES_ENC_us13_U190  ( .A1(_AES_ENC_us13_n1093 ), .A2(_AES_ENC_us13_n617 ), .ZN(_AES_ENC_us13_n876 ) );
NAND2_X2 _AES_ENC_us13_U189  ( .A1(_AES_ENC_us13_n576 ), .A2(_AES_ENC_us13_n876 ), .ZN(_AES_ENC_us13_n877 ) );
NAND2_X2 _AES_ENC_us13_U188  ( .A1(_AES_ENC_us13_n877 ), .A2(_AES_ENC_us13_n601 ), .ZN(_AES_ENC_us13_n888 ) );
NAND4_X2 _AES_ENC_us13_U179  ( .A1(_AES_ENC_us13_n889 ), .A2(_AES_ENC_us13_n888 ), .A3(_AES_ENC_us13_n887 ), .A4(_AES_ENC_us13_n886 ), .ZN(_AES_ENC_us13_n890 ) );
NAND2_X2 _AES_ENC_us13_U178  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n890 ), .ZN(_AES_ENC_us13_n903 ) );
OR2_X2 _AES_ENC_us13_U177  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n1059 ), .ZN(_AES_ENC_us13_n900 ) );
NAND2_X2 _AES_ENC_us13_U176  ( .A1(_AES_ENC_us13_n1073 ), .A2(_AES_ENC_us13_n1047 ), .ZN(_AES_ENC_us13_n899 ) );
NAND2_X2 _AES_ENC_us13_U175  ( .A1(_AES_ENC_us13_n1094 ), .A2(_AES_ENC_us13_n608 ), .ZN(_AES_ENC_us13_n898 ) );
NAND4_X2 _AES_ENC_us13_U167  ( .A1(_AES_ENC_us13_n900 ), .A2(_AES_ENC_us13_n899 ), .A3(_AES_ENC_us13_n898 ), .A4(_AES_ENC_us13_n897 ), .ZN(_AES_ENC_us13_n901 ) );
NAND2_X2 _AES_ENC_us13_U166  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n901 ), .ZN(_AES_ENC_us13_n902 ) );
NAND4_X2 _AES_ENC_us13_U165  ( .A1(_AES_ENC_us13_n905 ), .A2(_AES_ENC_us13_n904 ), .A3(_AES_ENC_us13_n903 ), .A4(_AES_ENC_us13_n902 ), .ZN(_AES_ENC_sa13_sub[4] ) );
NAND2_X2 _AES_ENC_us13_U164  ( .A1(_AES_ENC_us13_n1094 ), .A2(_AES_ENC_us13_n615 ), .ZN(_AES_ENC_us13_n922 ) );
NAND2_X2 _AES_ENC_us13_U163  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n989 ), .ZN(_AES_ENC_us13_n921 ) );
NAND4_X2 _AES_ENC_us13_U151  ( .A1(_AES_ENC_us13_n922 ), .A2(_AES_ENC_us13_n921 ), .A3(_AES_ENC_us13_n920 ), .A4(_AES_ENC_us13_n919 ), .ZN(_AES_ENC_us13_n923 ) );
NAND2_X2 _AES_ENC_us13_U150  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n923 ), .ZN(_AES_ENC_us13_n972 ) );
NAND2_X2 _AES_ENC_us13_U149  ( .A1(_AES_ENC_us13_n603 ), .A2(_AES_ENC_us13_n605 ), .ZN(_AES_ENC_us13_n924 ) );
NAND2_X2 _AES_ENC_us13_U148  ( .A1(_AES_ENC_us13_n1073 ), .A2(_AES_ENC_us13_n924 ), .ZN(_AES_ENC_us13_n939 ) );
NAND2_X2 _AES_ENC_us13_U147  ( .A1(_AES_ENC_us13_n926 ), .A2(_AES_ENC_us13_n925 ), .ZN(_AES_ENC_us13_n927 ) );
NAND2_X2 _AES_ENC_us13_U146  ( .A1(_AES_ENC_us13_n578 ), .A2(_AES_ENC_us13_n927 ), .ZN(_AES_ENC_us13_n928 ) );
NAND2_X2 _AES_ENC_us13_U145  ( .A1(_AES_ENC_us13_n928 ), .A2(_AES_ENC_us13_n1080 ), .ZN(_AES_ENC_us13_n938 ) );
OR2_X2 _AES_ENC_us13_U144  ( .A1(_AES_ENC_us13_n1117 ), .A2(_AES_ENC_us13_n589 ), .ZN(_AES_ENC_us13_n937 ) );
NAND4_X2 _AES_ENC_us13_U139  ( .A1(_AES_ENC_us13_n939 ), .A2(_AES_ENC_us13_n938 ), .A3(_AES_ENC_us13_n937 ), .A4(_AES_ENC_us13_n936 ), .ZN(_AES_ENC_us13_n940 ) );
NAND2_X2 _AES_ENC_us13_U138  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n940 ), .ZN(_AES_ENC_us13_n971 ) );
OR2_X2 _AES_ENC_us13_U137  ( .A1(_AES_ENC_us13_n577 ), .A2(_AES_ENC_us13_n941 ), .ZN(_AES_ENC_us13_n954 ) );
NAND2_X2 _AES_ENC_us13_U136  ( .A1(_AES_ENC_us13_n1096 ), .A2(_AES_ENC_us13_n618 ), .ZN(_AES_ENC_us13_n942 ) );
NAND2_X2 _AES_ENC_us13_U135  ( .A1(_AES_ENC_us13_n1048 ), .A2(_AES_ENC_us13_n942 ), .ZN(_AES_ENC_us13_n943 ) );
NAND2_X2 _AES_ENC_us13_U134  ( .A1(_AES_ENC_us13_n585 ), .A2(_AES_ENC_us13_n943 ), .ZN(_AES_ENC_us13_n944 ) );
NAND2_X2 _AES_ENC_us13_U133  ( .A1(_AES_ENC_us13_n944 ), .A2(_AES_ENC_us13_n599 ), .ZN(_AES_ENC_us13_n953 ) );
NAND4_X2 _AES_ENC_us13_U125  ( .A1(_AES_ENC_us13_n954 ), .A2(_AES_ENC_us13_n953 ), .A3(_AES_ENC_us13_n952 ), .A4(_AES_ENC_us13_n951 ), .ZN(_AES_ENC_us13_n955 ) );
NAND2_X2 _AES_ENC_us13_U124  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n955 ), .ZN(_AES_ENC_us13_n970 ) );
NAND2_X2 _AES_ENC_us13_U123  ( .A1(_AES_ENC_us13_n1094 ), .A2(_AES_ENC_us13_n1071 ), .ZN(_AES_ENC_us13_n967 ) );
NAND2_X2 _AES_ENC_us13_U122  ( .A1(_AES_ENC_us13_n956 ), .A2(_AES_ENC_us13_n1030 ), .ZN(_AES_ENC_us13_n966 ) );
NAND4_X2 _AES_ENC_us13_U114  ( .A1(_AES_ENC_us13_n967 ), .A2(_AES_ENC_us13_n966 ), .A3(_AES_ENC_us13_n965 ), .A4(_AES_ENC_us13_n964 ), .ZN(_AES_ENC_us13_n968 ) );
NAND2_X2 _AES_ENC_us13_U113  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n968 ), .ZN(_AES_ENC_us13_n969 ) );
NAND4_X2 _AES_ENC_us13_U112  ( .A1(_AES_ENC_us13_n972 ), .A2(_AES_ENC_us13_n971 ), .A3(_AES_ENC_us13_n970 ), .A4(_AES_ENC_us13_n969 ), .ZN(_AES_ENC_sa13_sub[5] ) );
NAND2_X2 _AES_ENC_us13_U111  ( .A1(_AES_ENC_us13_n570 ), .A2(_AES_ENC_us13_n1097 ), .ZN(_AES_ENC_us13_n973 ) );
NAND2_X2 _AES_ENC_us13_U110  ( .A1(_AES_ENC_us13_n1073 ), .A2(_AES_ENC_us13_n973 ), .ZN(_AES_ENC_us13_n987 ) );
NAND2_X2 _AES_ENC_us13_U109  ( .A1(_AES_ENC_us13_n974 ), .A2(_AES_ENC_us13_n1077 ), .ZN(_AES_ENC_us13_n975 ) );
NAND2_X2 _AES_ENC_us13_U108  ( .A1(_AES_ENC_us13_n587 ), .A2(_AES_ENC_us13_n975 ), .ZN(_AES_ENC_us13_n976 ) );
NAND2_X2 _AES_ENC_us13_U107  ( .A1(_AES_ENC_us13_n977 ), .A2(_AES_ENC_us13_n976 ), .ZN(_AES_ENC_us13_n986 ) );
NAND4_X2 _AES_ENC_us13_U99  ( .A1(_AES_ENC_us13_n987 ), .A2(_AES_ENC_us13_n986 ), .A3(_AES_ENC_us13_n985 ), .A4(_AES_ENC_us13_n984 ), .ZN(_AES_ENC_us13_n988 ) );
NAND2_X2 _AES_ENC_us13_U98  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n988 ), .ZN(_AES_ENC_us13_n1044 ) );
NAND2_X2 _AES_ENC_us13_U97  ( .A1(_AES_ENC_us13_n1073 ), .A2(_AES_ENC_us13_n989 ), .ZN(_AES_ENC_us13_n1004 ) );
NAND2_X2 _AES_ENC_us13_U96  ( .A1(_AES_ENC_us13_n1092 ), .A2(_AES_ENC_us13_n605 ), .ZN(_AES_ENC_us13_n1003 ) );
NAND4_X2 _AES_ENC_us13_U85  ( .A1(_AES_ENC_us13_n1004 ), .A2(_AES_ENC_us13_n1003 ), .A3(_AES_ENC_us13_n1002 ), .A4(_AES_ENC_us13_n1001 ), .ZN(_AES_ENC_us13_n1005 ) );
NAND2_X2 _AES_ENC_us13_U84  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n1005 ), .ZN(_AES_ENC_us13_n1043 ) );
NAND2_X2 _AES_ENC_us13_U83  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n626 ), .ZN(_AES_ENC_us13_n1020 ) );
NAND2_X2 _AES_ENC_us13_U82  ( .A1(_AES_ENC_us13_n1050 ), .A2(_AES_ENC_us13_n612 ), .ZN(_AES_ENC_us13_n1019 ) );
NAND2_X2 _AES_ENC_us13_U77  ( .A1(_AES_ENC_us13_n1059 ), .A2(_AES_ENC_us13_n1114 ), .ZN(_AES_ENC_us13_n1012 ) );
NAND2_X2 _AES_ENC_us13_U76  ( .A1(_AES_ENC_us13_n1010 ), .A2(_AES_ENC_us13_n604 ), .ZN(_AES_ENC_us13_n1011 ) );
NAND2_X2 _AES_ENC_us13_U75  ( .A1(_AES_ENC_us13_n1012 ), .A2(_AES_ENC_us13_n1011 ), .ZN(_AES_ENC_us13_n1016 ) );
NAND4_X2 _AES_ENC_us13_U70  ( .A1(_AES_ENC_us13_n1020 ), .A2(_AES_ENC_us13_n1019 ), .A3(_AES_ENC_us13_n1018 ), .A4(_AES_ENC_us13_n1017 ), .ZN(_AES_ENC_us13_n1021 ) );
NAND2_X2 _AES_ENC_us13_U69  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n1021 ), .ZN(_AES_ENC_us13_n1042 ) );
NAND2_X2 _AES_ENC_us13_U68  ( .A1(_AES_ENC_us13_n1022 ), .A2(_AES_ENC_us13_n1093 ), .ZN(_AES_ENC_us13_n1039 ) );
NAND2_X2 _AES_ENC_us13_U67  ( .A1(_AES_ENC_us13_n1050 ), .A2(_AES_ENC_us13_n1023 ), .ZN(_AES_ENC_us13_n1038 ) );
NAND2_X2 _AES_ENC_us13_U66  ( .A1(_AES_ENC_us13_n1024 ), .A2(_AES_ENC_us13_n1071 ), .ZN(_AES_ENC_us13_n1037 ) );
AND2_X2 _AES_ENC_us13_U60  ( .A1(_AES_ENC_us13_n1030 ), .A2(_AES_ENC_us13_n621 ), .ZN(_AES_ENC_us13_n1078 ) );
NAND4_X2 _AES_ENC_us13_U56  ( .A1(_AES_ENC_us13_n1039 ), .A2(_AES_ENC_us13_n1038 ), .A3(_AES_ENC_us13_n1037 ), .A4(_AES_ENC_us13_n1036 ), .ZN(_AES_ENC_us13_n1040 ) );
NAND2_X2 _AES_ENC_us13_U55  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n1040 ), .ZN(_AES_ENC_us13_n1041 ) );
NAND4_X2 _AES_ENC_us13_U54  ( .A1(_AES_ENC_us13_n1044 ), .A2(_AES_ENC_us13_n1043 ), .A3(_AES_ENC_us13_n1042 ), .A4(_AES_ENC_us13_n1041 ), .ZN(_AES_ENC_sa13_sub[6] ) );
NAND2_X2 _AES_ENC_us13_U53  ( .A1(_AES_ENC_us13_n1072 ), .A2(_AES_ENC_us13_n1045 ), .ZN(_AES_ENC_us13_n1068 ) );
NAND2_X2 _AES_ENC_us13_U52  ( .A1(_AES_ENC_us13_n1046 ), .A2(_AES_ENC_us13_n603 ), .ZN(_AES_ENC_us13_n1067 ) );
NAND2_X2 _AES_ENC_us13_U51  ( .A1(_AES_ENC_us13_n1094 ), .A2(_AES_ENC_us13_n1047 ), .ZN(_AES_ENC_us13_n1066 ) );
NAND4_X2 _AES_ENC_us13_U40  ( .A1(_AES_ENC_us13_n1068 ), .A2(_AES_ENC_us13_n1067 ), .A3(_AES_ENC_us13_n1066 ), .A4(_AES_ENC_us13_n1065 ), .ZN(_AES_ENC_us13_n1069 ) );
NAND2_X2 _AES_ENC_us13_U39  ( .A1(_AES_ENC_us13_n1070 ), .A2(_AES_ENC_us13_n1069 ), .ZN(_AES_ENC_us13_n1135 ) );
NAND2_X2 _AES_ENC_us13_U38  ( .A1(_AES_ENC_us13_n1072 ), .A2(_AES_ENC_us13_n1071 ), .ZN(_AES_ENC_us13_n1088 ) );
NAND2_X2 _AES_ENC_us13_U37  ( .A1(_AES_ENC_us13_n1073 ), .A2(_AES_ENC_us13_n608 ), .ZN(_AES_ENC_us13_n1087 ) );
NAND4_X2 _AES_ENC_us13_U28  ( .A1(_AES_ENC_us13_n1088 ), .A2(_AES_ENC_us13_n1087 ), .A3(_AES_ENC_us13_n1086 ), .A4(_AES_ENC_us13_n1085 ), .ZN(_AES_ENC_us13_n1089 ) );
NAND2_X2 _AES_ENC_us13_U27  ( .A1(_AES_ENC_us13_n1090 ), .A2(_AES_ENC_us13_n1089 ), .ZN(_AES_ENC_us13_n1134 ) );
NAND2_X2 _AES_ENC_us13_U26  ( .A1(_AES_ENC_us13_n1091 ), .A2(_AES_ENC_us13_n1093 ), .ZN(_AES_ENC_us13_n1111 ) );
NAND2_X2 _AES_ENC_us13_U25  ( .A1(_AES_ENC_us13_n1092 ), .A2(_AES_ENC_us13_n1120 ), .ZN(_AES_ENC_us13_n1110 ) );
AND2_X2 _AES_ENC_us13_U22  ( .A1(_AES_ENC_us13_n1097 ), .A2(_AES_ENC_us13_n1096 ), .ZN(_AES_ENC_us13_n1098 ) );
NAND4_X2 _AES_ENC_us13_U14  ( .A1(_AES_ENC_us13_n1111 ), .A2(_AES_ENC_us13_n1110 ), .A3(_AES_ENC_us13_n1109 ), .A4(_AES_ENC_us13_n1108 ), .ZN(_AES_ENC_us13_n1112 ) );
NAND2_X2 _AES_ENC_us13_U13  ( .A1(_AES_ENC_us13_n1113 ), .A2(_AES_ENC_us13_n1112 ), .ZN(_AES_ENC_us13_n1133 ) );
NAND2_X2 _AES_ENC_us13_U12  ( .A1(_AES_ENC_us13_n1115 ), .A2(_AES_ENC_us13_n1114 ), .ZN(_AES_ENC_us13_n1129 ) );
OR2_X2 _AES_ENC_us13_U11  ( .A1(_AES_ENC_us13_n581 ), .A2(_AES_ENC_us13_n1116 ), .ZN(_AES_ENC_us13_n1128 ) );
NAND4_X2 _AES_ENC_us13_U3  ( .A1(_AES_ENC_us13_n1129 ), .A2(_AES_ENC_us13_n1128 ), .A3(_AES_ENC_us13_n1127 ), .A4(_AES_ENC_us13_n1126 ), .ZN(_AES_ENC_us13_n1130 ) );
NAND2_X2 _AES_ENC_us13_U2  ( .A1(_AES_ENC_us13_n1131 ), .A2(_AES_ENC_us13_n1130 ), .ZN(_AES_ENC_us13_n1132 ) );
NAND4_X2 _AES_ENC_us13_U1  ( .A1(_AES_ENC_us13_n1135 ), .A2(_AES_ENC_us13_n1134 ), .A3(_AES_ENC_us13_n1133 ), .A4(_AES_ENC_us13_n1132 ), .ZN(_AES_ENC_sa13_sub[7] ) );
INV_X4 _AES_ENC_us20_U575  ( .A(_AES_ENC_sa20[0]), .ZN(_AES_ENC_us20_n627 ));
INV_X4 _AES_ENC_us20_U574  ( .A(_AES_ENC_us20_n1053 ), .ZN(_AES_ENC_us20_n625 ) );
INV_X4 _AES_ENC_us20_U573  ( .A(_AES_ENC_us20_n1103 ), .ZN(_AES_ENC_us20_n623 ) );
INV_X4 _AES_ENC_us20_U572  ( .A(_AES_ENC_us20_n1056 ), .ZN(_AES_ENC_us20_n622 ) );
INV_X4 _AES_ENC_us20_U571  ( .A(_AES_ENC_us20_n1102 ), .ZN(_AES_ENC_us20_n621 ) );
INV_X4 _AES_ENC_us20_U570  ( .A(_AES_ENC_us20_n1074 ), .ZN(_AES_ENC_us20_n620 ) );
INV_X4 _AES_ENC_us20_U569  ( .A(_AES_ENC_us20_n929 ), .ZN(_AES_ENC_us20_n619 ) );
INV_X4 _AES_ENC_us20_U568  ( .A(_AES_ENC_us20_n1091 ), .ZN(_AES_ENC_us20_n618 ) );
INV_X4 _AES_ENC_us20_U567  ( .A(_AES_ENC_us20_n826 ), .ZN(_AES_ENC_us20_n617 ) );
INV_X4 _AES_ENC_us20_U566  ( .A(_AES_ENC_us20_n1031 ), .ZN(_AES_ENC_us20_n616 ) );
INV_X4 _AES_ENC_us20_U565  ( .A(_AES_ENC_us20_n1054 ), .ZN(_AES_ENC_us20_n615 ) );
INV_X4 _AES_ENC_us20_U564  ( .A(_AES_ENC_us20_n1025 ), .ZN(_AES_ENC_us20_n614 ) );
INV_X4 _AES_ENC_us20_U563  ( .A(_AES_ENC_us20_n990 ), .ZN(_AES_ENC_us20_n613 ) );
INV_X4 _AES_ENC_us20_U562  ( .A(_AES_ENC_sa20[4]), .ZN(_AES_ENC_us20_n612 ));
INV_X4 _AES_ENC_us20_U561  ( .A(_AES_ENC_us20_n881 ), .ZN(_AES_ENC_us20_n611 ) );
INV_X4 _AES_ENC_us20_U560  ( .A(_AES_ENC_us20_n1022 ), .ZN(_AES_ENC_us20_n610 ) );
INV_X4 _AES_ENC_us20_U559  ( .A(_AES_ENC_us20_n1120 ), .ZN(_AES_ENC_us20_n609 ) );
INV_X4 _AES_ENC_us20_U558  ( .A(_AES_ENC_us20_n977 ), .ZN(_AES_ENC_us20_n608 ) );
INV_X4 _AES_ENC_us20_U557  ( .A(_AES_ENC_us20_n926 ), .ZN(_AES_ENC_us20_n607 ) );
INV_X4 _AES_ENC_us20_U556  ( .A(_AES_ENC_us20_n910 ), .ZN(_AES_ENC_us20_n606 ) );
INV_X4 _AES_ENC_us20_U555  ( .A(_AES_ENC_us20_n1121 ), .ZN(_AES_ENC_us20_n605 ) );
INV_X4 _AES_ENC_us20_U554  ( .A(_AES_ENC_us20_n1009 ), .ZN(_AES_ENC_us20_n604 ) );
INV_X4 _AES_ENC_us20_U553  ( .A(_AES_ENC_us20_n1080 ), .ZN(_AES_ENC_us20_n602 ) );
INV_X4 _AES_ENC_us20_U552  ( .A(_AES_ENC_us20_n821 ), .ZN(_AES_ENC_us20_n600 ) );
INV_X4 _AES_ENC_us20_U551  ( .A(_AES_ENC_us20_n1013 ), .ZN(_AES_ENC_us20_n599 ) );
INV_X4 _AES_ENC_us20_U550  ( .A(_AES_ENC_us20_n1058 ), .ZN(_AES_ENC_us20_n598 ) );
INV_X4 _AES_ENC_us20_U549  ( .A(_AES_ENC_us20_n906 ), .ZN(_AES_ENC_us20_n597 ) );
INV_X4 _AES_ENC_us20_U548  ( .A(_AES_ENC_us20_n1048 ), .ZN(_AES_ENC_us20_n595 ) );
INV_X4 _AES_ENC_us20_U547  ( .A(_AES_ENC_us20_n974 ), .ZN(_AES_ENC_us20_n594 ) );
INV_X4 _AES_ENC_us20_U546  ( .A(_AES_ENC_sa20[2]), .ZN(_AES_ENC_us20_n593 ));
INV_X4 _AES_ENC_us20_U545  ( .A(_AES_ENC_us20_n800 ), .ZN(_AES_ENC_us20_n592 ) );
INV_X4 _AES_ENC_us20_U544  ( .A(_AES_ENC_us20_n925 ), .ZN(_AES_ENC_us20_n591 ) );
INV_X4 _AES_ENC_us20_U543  ( .A(_AES_ENC_us20_n824 ), .ZN(_AES_ENC_us20_n590 ) );
INV_X4 _AES_ENC_us20_U542  ( .A(_AES_ENC_us20_n959 ), .ZN(_AES_ENC_us20_n589 ) );
INV_X4 _AES_ENC_us20_U541  ( .A(_AES_ENC_us20_n779 ), .ZN(_AES_ENC_us20_n588 ) );
INV_X4 _AES_ENC_us20_U540  ( .A(_AES_ENC_us20_n794 ), .ZN(_AES_ENC_us20_n585 ) );
INV_X4 _AES_ENC_us20_U539  ( .A(_AES_ENC_us20_n880 ), .ZN(_AES_ENC_us20_n583 ) );
INV_X4 _AES_ENC_us20_U538  ( .A(_AES_ENC_sa20[7]), .ZN(_AES_ENC_us20_n581 ));
INV_X4 _AES_ENC_us20_U537  ( .A(_AES_ENC_us20_n992 ), .ZN(_AES_ENC_us20_n578 ) );
INV_X4 _AES_ENC_us20_U536  ( .A(_AES_ENC_us20_n1114 ), .ZN(_AES_ENC_us20_n577 ) );
INV_X4 _AES_ENC_us20_U535  ( .A(_AES_ENC_us20_n1092 ), .ZN(_AES_ENC_us20_n574 ) );
NOR2_X2 _AES_ENC_us20_U534  ( .A1(_AES_ENC_sa20[0]), .A2(_AES_ENC_sa20[6]),.ZN(_AES_ENC_us20_n1090 ) );
NOR2_X2 _AES_ENC_us20_U533  ( .A1(_AES_ENC_us20_n627 ), .A2(_AES_ENC_sa20[6]), .ZN(_AES_ENC_us20_n1070 ) );
NOR2_X2 _AES_ENC_us20_U532  ( .A1(_AES_ENC_sa20[4]), .A2(_AES_ENC_sa20[3]),.ZN(_AES_ENC_us20_n1025 ) );
INV_X4 _AES_ENC_us20_U531  ( .A(_AES_ENC_us20_n569 ), .ZN(_AES_ENC_us20_n572 ) );
NOR2_X2 _AES_ENC_us20_U530  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n765 ) );
NOR2_X2 _AES_ENC_us20_U529  ( .A1(_AES_ENC_sa20[4]), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n764 ) );
NOR2_X2 _AES_ENC_us20_U528  ( .A1(_AES_ENC_us20_n765 ), .A2(_AES_ENC_us20_n764 ), .ZN(_AES_ENC_us20_n766 ) );
NOR2_X2 _AES_ENC_us20_U527  ( .A1(_AES_ENC_us20_n766 ), .A2(_AES_ENC_us20_n589 ), .ZN(_AES_ENC_us20_n767 ) );
INV_X4 _AES_ENC_us20_U526  ( .A(_AES_ENC_sa20[3]), .ZN(_AES_ENC_us20_n624 ));
NAND3_X2 _AES_ENC_us20_U525  ( .A1(_AES_ENC_us20_n652 ), .A2(_AES_ENC_us20_n596 ), .A3(_AES_ENC_sa20[7]), .ZN(_AES_ENC_us20_n653 ));
NOR2_X2 _AES_ENC_us20_U524  ( .A1(_AES_ENC_us20_n593 ), .A2(_AES_ENC_sa20[5]), .ZN(_AES_ENC_us20_n925 ) );
NOR2_X2 _AES_ENC_us20_U523  ( .A1(_AES_ENC_sa20[5]), .A2(_AES_ENC_sa20[2]),.ZN(_AES_ENC_us20_n974 ) );
INV_X4 _AES_ENC_us20_U522  ( .A(_AES_ENC_sa20[5]), .ZN(_AES_ENC_us20_n596 ));
NOR2_X2 _AES_ENC_us20_U521  ( .A1(_AES_ENC_us20_n593 ), .A2(_AES_ENC_sa20[7]), .ZN(_AES_ENC_us20_n779 ) );
NAND3_X2 _AES_ENC_us20_U520  ( .A1(_AES_ENC_us20_n679 ), .A2(_AES_ENC_us20_n678 ), .A3(_AES_ENC_us20_n677 ), .ZN(_AES_ENC_sa20_sub[0] ) );
NOR2_X2 _AES_ENC_us20_U519  ( .A1(_AES_ENC_us20_n596 ), .A2(_AES_ENC_sa20[2]), .ZN(_AES_ENC_us20_n1048 ) );
NOR3_X2 _AES_ENC_us20_U518  ( .A1(_AES_ENC_us20_n581 ), .A2(_AES_ENC_sa20[5]), .A3(_AES_ENC_us20_n704 ), .ZN(_AES_ENC_us20_n706 ));
NOR2_X2 _AES_ENC_us20_U517  ( .A1(_AES_ENC_us20_n1117 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n707 ) );
NOR2_X2 _AES_ENC_us20_U516  ( .A1(_AES_ENC_sa20[4]), .A2(_AES_ENC_us20_n574 ), .ZN(_AES_ENC_us20_n705 ) );
NOR3_X2 _AES_ENC_us20_U515  ( .A1(_AES_ENC_us20_n707 ), .A2(_AES_ENC_us20_n706 ), .A3(_AES_ENC_us20_n705 ), .ZN(_AES_ENC_us20_n713 ) );
NOR4_X2 _AES_ENC_us20_U512  ( .A1(_AES_ENC_us20_n633 ), .A2(_AES_ENC_us20_n632 ), .A3(_AES_ENC_us20_n631 ), .A4(_AES_ENC_us20_n630 ), .ZN(_AES_ENC_us20_n634 ) );
NOR2_X2 _AES_ENC_us20_U510  ( .A1(_AES_ENC_us20_n629 ), .A2(_AES_ENC_us20_n628 ), .ZN(_AES_ENC_us20_n635 ) );
NAND3_X2 _AES_ENC_us20_U509  ( .A1(_AES_ENC_sa20[2]), .A2(_AES_ENC_sa20[7]), .A3(_AES_ENC_us20_n1059 ), .ZN(_AES_ENC_us20_n636 ) );
NOR2_X2 _AES_ENC_us20_U508  ( .A1(_AES_ENC_sa20[7]), .A2(_AES_ENC_sa20[2]),.ZN(_AES_ENC_us20_n794 ) );
NOR2_X2 _AES_ENC_us20_U507  ( .A1(_AES_ENC_sa20[4]), .A2(_AES_ENC_sa20[1]),.ZN(_AES_ENC_us20_n1102 ) );
NOR2_X2 _AES_ENC_us20_U506  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_sa20[3]), .ZN(_AES_ENC_us20_n1053 ) );
NOR2_X2 _AES_ENC_us20_U505  ( .A1(_AES_ENC_us20_n588 ), .A2(_AES_ENC_sa20[5]), .ZN(_AES_ENC_us20_n1024 ) );
NOR2_X2 _AES_ENC_us20_U504  ( .A1(_AES_ENC_us20_n577 ), .A2(_AES_ENC_sa20[2]), .ZN(_AES_ENC_us20_n1093 ) );
NOR2_X2 _AES_ENC_us20_U503  ( .A1(_AES_ENC_us20_n585 ), .A2(_AES_ENC_sa20[5]), .ZN(_AES_ENC_us20_n1094 ) );
NOR2_X2 _AES_ENC_us20_U502  ( .A1(_AES_ENC_us20_n612 ), .A2(_AES_ENC_sa20[3]), .ZN(_AES_ENC_us20_n931 ) );
INV_X4 _AES_ENC_us20_U501  ( .A(_AES_ENC_us20_n570 ), .ZN(_AES_ENC_us20_n573 ) );
NOR2_X2 _AES_ENC_us20_U500  ( .A1(_AES_ENC_us20_n1053 ), .A2(_AES_ENC_us20_n1095 ), .ZN(_AES_ENC_us20_n639 ) );
NOR3_X2 _AES_ENC_us20_U499  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n573 ), .A3(_AES_ENC_us20_n1074 ), .ZN(_AES_ENC_us20_n641 ) );
NOR2_X2 _AES_ENC_us20_U498  ( .A1(_AES_ENC_us20_n639 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n640 ) );
NOR2_X2 _AES_ENC_us20_U497  ( .A1(_AES_ENC_us20_n641 ), .A2(_AES_ENC_us20_n640 ), .ZN(_AES_ENC_us20_n646 ) );
NOR3_X2 _AES_ENC_us20_U496  ( .A1(_AES_ENC_us20_n995 ), .A2(_AES_ENC_us20_n578 ), .A3(_AES_ENC_us20_n994 ), .ZN(_AES_ENC_us20_n1002 ) );
NOR2_X2 _AES_ENC_us20_U495  ( .A1(_AES_ENC_us20_n909 ), .A2(_AES_ENC_us20_n908 ), .ZN(_AES_ENC_us20_n920 ) );
NOR2_X2 _AES_ENC_us20_U494  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n823 ) );
NOR2_X2 _AES_ENC_us20_U492  ( .A1(_AES_ENC_us20_n612 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n822 ) );
NOR2_X2 _AES_ENC_us20_U491  ( .A1(_AES_ENC_us20_n823 ), .A2(_AES_ENC_us20_n822 ), .ZN(_AES_ENC_us20_n825 ) );
NOR2_X2 _AES_ENC_us20_U490  ( .A1(_AES_ENC_sa20[1]), .A2(_AES_ENC_us20_n601 ), .ZN(_AES_ENC_us20_n913 ) );
NOR2_X2 _AES_ENC_us20_U489  ( .A1(_AES_ENC_us20_n913 ), .A2(_AES_ENC_us20_n1091 ), .ZN(_AES_ENC_us20_n914 ) );
NOR2_X2 _AES_ENC_us20_U488  ( .A1(_AES_ENC_us20_n826 ), .A2(_AES_ENC_us20_n572 ), .ZN(_AES_ENC_us20_n827 ) );
NOR3_X2 _AES_ENC_us20_U487  ( .A1(_AES_ENC_us20_n769 ), .A2(_AES_ENC_us20_n768 ), .A3(_AES_ENC_us20_n767 ), .ZN(_AES_ENC_us20_n775 ) );
NOR2_X2 _AES_ENC_us20_U486  ( .A1(_AES_ENC_us20_n1056 ), .A2(_AES_ENC_us20_n1053 ), .ZN(_AES_ENC_us20_n749 ) );
NOR2_X2 _AES_ENC_us20_U483  ( .A1(_AES_ENC_us20_n749 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n752 ) );
INV_X4 _AES_ENC_us20_U482  ( .A(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n626 ));
NOR2_X2 _AES_ENC_us20_U480  ( .A1(_AES_ENC_us20_n1054 ), .A2(_AES_ENC_us20_n1053 ), .ZN(_AES_ENC_us20_n1055 ) );
OR2_X4 _AES_ENC_us20_U479  ( .A1(_AES_ENC_us20_n1094 ), .A2(_AES_ENC_us20_n1093 ), .ZN(_AES_ENC_us20_n571 ) );
AND2_X2 _AES_ENC_us20_U478  ( .A1(_AES_ENC_us20_n571 ), .A2(_AES_ENC_us20_n1095 ), .ZN(_AES_ENC_us20_n1101 ) );
NOR2_X2 _AES_ENC_us20_U477  ( .A1(_AES_ENC_us20_n1074 ), .A2(_AES_ENC_us20_n931 ), .ZN(_AES_ENC_us20_n796 ) );
NOR2_X2 _AES_ENC_us20_U474  ( .A1(_AES_ENC_us20_n796 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n797 ) );
NOR2_X2 _AES_ENC_us20_U473  ( .A1(_AES_ENC_us20_n932 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n933 ) );
NOR2_X2 _AES_ENC_us20_U472  ( .A1(_AES_ENC_us20_n929 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n935 ) );
NOR2_X2 _AES_ENC_us20_U471  ( .A1(_AES_ENC_us20_n931 ), .A2(_AES_ENC_us20_n930 ), .ZN(_AES_ENC_us20_n934 ) );
NOR3_X2 _AES_ENC_us20_U470  ( .A1(_AES_ENC_us20_n935 ), .A2(_AES_ENC_us20_n934 ), .A3(_AES_ENC_us20_n933 ), .ZN(_AES_ENC_us20_n936 ) );
NOR2_X2 _AES_ENC_us20_U469  ( .A1(_AES_ENC_us20_n612 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n1075 ) );
NOR2_X2 _AES_ENC_us20_U468  ( .A1(_AES_ENC_us20_n572 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n949 ) );
NOR2_X2 _AES_ENC_us20_U467  ( .A1(_AES_ENC_us20_n1049 ), .A2(_AES_ENC_us20_n595 ), .ZN(_AES_ENC_us20_n1051 ) );
NOR2_X2 _AES_ENC_us20_U466  ( .A1(_AES_ENC_us20_n1051 ), .A2(_AES_ENC_us20_n1050 ), .ZN(_AES_ENC_us20_n1052 ) );
NOR2_X2 _AES_ENC_us20_U465  ( .A1(_AES_ENC_us20_n1052 ), .A2(_AES_ENC_us20_n604 ), .ZN(_AES_ENC_us20_n1064 ) );
NOR2_X2 _AES_ENC_us20_U464  ( .A1(_AES_ENC_sa20[1]), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n631 ) );
NOR2_X2 _AES_ENC_us20_U463  ( .A1(_AES_ENC_us20_n1025 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n980 ) );
NOR2_X2 _AES_ENC_us20_U462  ( .A1(_AES_ENC_us20_n1073 ), .A2(_AES_ENC_us20_n1094 ), .ZN(_AES_ENC_us20_n795 ) );
NOR2_X2 _AES_ENC_us20_U461  ( .A1(_AES_ENC_us20_n795 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n799 ) );
NOR2_X2 _AES_ENC_us20_U460  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n981 ) );
NOR2_X2 _AES_ENC_us20_U459  ( .A1(_AES_ENC_us20_n1102 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n643 ) );
NOR2_X2 _AES_ENC_us20_U458  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n624 ), .ZN(_AES_ENC_us20_n642 ) );
NOR2_X2 _AES_ENC_us20_U455  ( .A1(_AES_ENC_us20_n911 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n644 ) );
NOR4_X2 _AES_ENC_us20_U448  ( .A1(_AES_ENC_us20_n644 ), .A2(_AES_ENC_us20_n643 ), .A3(_AES_ENC_us20_n804 ), .A4(_AES_ENC_us20_n642 ), .ZN(_AES_ENC_us20_n645 ) );
NOR2_X2 _AES_ENC_us20_U447  ( .A1(_AES_ENC_us20_n1102 ), .A2(_AES_ENC_us20_n910 ), .ZN(_AES_ENC_us20_n932 ) );
NOR2_X2 _AES_ENC_us20_U442  ( .A1(_AES_ENC_us20_n1102 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n755 ) );
NOR2_X2 _AES_ENC_us20_U441  ( .A1(_AES_ENC_us20_n931 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n743 ) );
NOR2_X2 _AES_ENC_us20_U438  ( .A1(_AES_ENC_us20_n1072 ), .A2(_AES_ENC_us20_n1094 ), .ZN(_AES_ENC_us20_n930 ) );
NOR2_X2 _AES_ENC_us20_U435  ( .A1(_AES_ENC_us20_n1074 ), .A2(_AES_ENC_us20_n1025 ), .ZN(_AES_ENC_us20_n891 ) );
NOR2_X2 _AES_ENC_us20_U434  ( .A1(_AES_ENC_us20_n891 ), .A2(_AES_ENC_us20_n591 ), .ZN(_AES_ENC_us20_n894 ) );
NOR3_X2 _AES_ENC_us20_U433  ( .A1(_AES_ENC_us20_n601 ), .A2(_AES_ENC_sa20[1]), .A3(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n683 ));
INV_X4 _AES_ENC_us20_U428  ( .A(_AES_ENC_us20_n931 ), .ZN(_AES_ENC_us20_n601 ) );
NOR2_X2 _AES_ENC_us20_U427  ( .A1(_AES_ENC_us20_n996 ), .A2(_AES_ENC_us20_n931 ), .ZN(_AES_ENC_us20_n704 ) );
NOR2_X2 _AES_ENC_us20_U421  ( .A1(_AES_ENC_us20_n931 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n685 ) );
NOR2_X2 _AES_ENC_us20_U420  ( .A1(_AES_ENC_us20_n1029 ), .A2(_AES_ENC_us20_n1025 ), .ZN(_AES_ENC_us20_n1079 ) );
NOR3_X2 _AES_ENC_us20_U419  ( .A1(_AES_ENC_us20_n620 ), .A2(_AES_ENC_us20_n1025 ), .A3(_AES_ENC_us20_n594 ), .ZN(_AES_ENC_us20_n945 ) );
NOR2_X2 _AES_ENC_us20_U418  ( .A1(_AES_ENC_us20_n596 ), .A2(_AES_ENC_us20_n593 ), .ZN(_AES_ENC_us20_n800 ) );
NOR3_X2 _AES_ENC_us20_U417  ( .A1(_AES_ENC_us20_n598 ), .A2(_AES_ENC_us20_n581 ), .A3(_AES_ENC_us20_n593 ), .ZN(_AES_ENC_us20_n798 ) );
NOR3_X2 _AES_ENC_us20_U416  ( .A1(_AES_ENC_us20_n592 ), .A2(_AES_ENC_us20_n572 ), .A3(_AES_ENC_us20_n589 ), .ZN(_AES_ENC_us20_n962 ) );
NOR3_X2 _AES_ENC_us20_U415  ( .A1(_AES_ENC_us20_n959 ), .A2(_AES_ENC_us20_n572 ), .A3(_AES_ENC_us20_n591 ), .ZN(_AES_ENC_us20_n768 ) );
NOR3_X2 _AES_ENC_us20_U414  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n572 ), .A3(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n694 ) );
NOR3_X2 _AES_ENC_us20_U413  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n572 ), .A3(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n895 ) );
NOR3_X2 _AES_ENC_us20_U410  ( .A1(_AES_ENC_us20_n1008 ), .A2(_AES_ENC_us20_n1007 ), .A3(_AES_ENC_us20_n1006 ), .ZN(_AES_ENC_us20_n1018 ) );
NOR4_X2 _AES_ENC_us20_U409  ( .A1(_AES_ENC_us20_n806 ), .A2(_AES_ENC_us20_n805 ), .A3(_AES_ENC_us20_n804 ), .A4(_AES_ENC_us20_n803 ), .ZN(_AES_ENC_us20_n807 ) );
NOR3_X2 _AES_ENC_us20_U406  ( .A1(_AES_ENC_us20_n799 ), .A2(_AES_ENC_us20_n798 ), .A3(_AES_ENC_us20_n797 ), .ZN(_AES_ENC_us20_n808 ) );
NOR4_X2 _AES_ENC_us20_U405  ( .A1(_AES_ENC_us20_n843 ), .A2(_AES_ENC_us20_n842 ), .A3(_AES_ENC_us20_n841 ), .A4(_AES_ENC_us20_n840 ), .ZN(_AES_ENC_us20_n844 ) );
NOR2_X2 _AES_ENC_us20_U404  ( .A1(_AES_ENC_us20_n669 ), .A2(_AES_ENC_us20_n668 ), .ZN(_AES_ENC_us20_n673 ) );
NOR4_X2 _AES_ENC_us20_U403  ( .A1(_AES_ENC_us20_n946 ), .A2(_AES_ENC_us20_n1046 ), .A3(_AES_ENC_us20_n671 ), .A4(_AES_ENC_us20_n670 ), .ZN(_AES_ENC_us20_n672 ) );
NOR4_X2 _AES_ENC_us20_U401  ( .A1(_AES_ENC_us20_n711 ), .A2(_AES_ENC_us20_n710 ), .A3(_AES_ENC_us20_n709 ), .A4(_AES_ENC_us20_n708 ), .ZN(_AES_ENC_us20_n712 ) );
NOR4_X2 _AES_ENC_us20_U400  ( .A1(_AES_ENC_us20_n963 ), .A2(_AES_ENC_us20_n962 ), .A3(_AES_ENC_us20_n961 ), .A4(_AES_ENC_us20_n960 ), .ZN(_AES_ENC_us20_n964 ) );
NOR3_X2 _AES_ENC_us20_U399  ( .A1(_AES_ENC_us20_n1101 ), .A2(_AES_ENC_us20_n1100 ), .A3(_AES_ENC_us20_n1099 ), .ZN(_AES_ENC_us20_n1109 ) );
NOR3_X2 _AES_ENC_us20_U398  ( .A1(_AES_ENC_us20_n743 ), .A2(_AES_ENC_us20_n742 ), .A3(_AES_ENC_us20_n741 ), .ZN(_AES_ENC_us20_n744 ) );
NOR2_X2 _AES_ENC_us20_U397  ( .A1(_AES_ENC_us20_n697 ), .A2(_AES_ENC_us20_n658 ), .ZN(_AES_ENC_us20_n659 ) );
NOR2_X2 _AES_ENC_us20_U396  ( .A1(_AES_ENC_us20_n1078 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n1033 ) );
NOR2_X2 _AES_ENC_us20_U393  ( .A1(_AES_ENC_us20_n1031 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n1032 ) );
NOR3_X2 _AES_ENC_us20_U390  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n1025 ), .A3(_AES_ENC_us20_n1074 ), .ZN(_AES_ENC_us20_n1035 ) );
NOR4_X2 _AES_ENC_us20_U389  ( .A1(_AES_ENC_us20_n1035 ), .A2(_AES_ENC_us20_n1034 ), .A3(_AES_ENC_us20_n1033 ), .A4(_AES_ENC_us20_n1032 ), .ZN(_AES_ENC_us20_n1036 ) );
NOR2_X2 _AES_ENC_us20_U388  ( .A1(_AES_ENC_us20_n611 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n885 ) );
NOR2_X2 _AES_ENC_us20_U387  ( .A1(_AES_ENC_us20_n601 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n882 ) );
NOR2_X2 _AES_ENC_us20_U386  ( .A1(_AES_ENC_us20_n1053 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n884 ) );
NOR4_X2 _AES_ENC_us20_U385  ( .A1(_AES_ENC_us20_n885 ), .A2(_AES_ENC_us20_n884 ), .A3(_AES_ENC_us20_n883 ), .A4(_AES_ENC_us20_n882 ), .ZN(_AES_ENC_us20_n886 ) );
NOR2_X2 _AES_ENC_us20_U384  ( .A1(_AES_ENC_us20_n825 ), .A2(_AES_ENC_us20_n590 ), .ZN(_AES_ENC_us20_n830 ) );
NOR2_X2 _AES_ENC_us20_U383  ( .A1(_AES_ENC_us20_n827 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n829 ) );
NOR2_X2 _AES_ENC_us20_U382  ( .A1(_AES_ENC_us20_n572 ), .A2(_AES_ENC_us20_n574 ), .ZN(_AES_ENC_us20_n828 ) );
NOR4_X2 _AES_ENC_us20_U374  ( .A1(_AES_ENC_us20_n831 ), .A2(_AES_ENC_us20_n830 ), .A3(_AES_ENC_us20_n829 ), .A4(_AES_ENC_us20_n828 ), .ZN(_AES_ENC_us20_n832 ) );
NOR2_X2 _AES_ENC_us20_U373  ( .A1(_AES_ENC_us20_n587 ), .A2(_AES_ENC_us20_n603 ), .ZN(_AES_ENC_us20_n1104 ) );
NOR2_X2 _AES_ENC_us20_U372  ( .A1(_AES_ENC_us20_n1102 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n1106 ) );
NOR2_X2 _AES_ENC_us20_U370  ( .A1(_AES_ENC_us20_n1103 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n1105 ) );
NOR4_X2 _AES_ENC_us20_U369  ( .A1(_AES_ENC_us20_n1107 ), .A2(_AES_ENC_us20_n1106 ), .A3(_AES_ENC_us20_n1105 ), .A4(_AES_ENC_us20_n1104 ), .ZN(_AES_ENC_us20_n1108 ) );
NOR3_X2 _AES_ENC_us20_U368  ( .A1(_AES_ENC_us20_n959 ), .A2(_AES_ENC_us20_n624 ), .A3(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n963 ) );
NOR2_X2 _AES_ENC_us20_U367  ( .A1(_AES_ENC_us20_n596 ), .A2(_AES_ENC_us20_n581 ), .ZN(_AES_ENC_us20_n1114 ) );
INV_X4 _AES_ENC_us20_U366  ( .A(_AES_ENC_us20_n1024 ), .ZN(_AES_ENC_us20_n587 ) );
NOR3_X2 _AES_ENC_us20_U365  ( .A1(_AES_ENC_us20_n910 ), .A2(_AES_ENC_us20_n1059 ), .A3(_AES_ENC_us20_n593 ), .ZN(_AES_ENC_us20_n1115 ) );
INV_X4 _AES_ENC_us20_U364  ( .A(_AES_ENC_us20_n1094 ), .ZN(_AES_ENC_us20_n584 ) );
NOR2_X2 _AES_ENC_us20_U363  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n931 ), .ZN(_AES_ENC_us20_n1100 ) );
INV_X4 _AES_ENC_us20_U354  ( .A(_AES_ENC_us20_n1093 ), .ZN(_AES_ENC_us20_n575 ) );
NOR2_X2 _AES_ENC_us20_U353  ( .A1(_AES_ENC_us20_n569 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n929 ) );
NOR2_X2 _AES_ENC_us20_U352  ( .A1(_AES_ENC_us20_n609 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n926 ) );
NOR2_X2 _AES_ENC_us20_U351  ( .A1(_AES_ENC_us20_n572 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n1095 ) );
NOR2_X2 _AES_ENC_us20_U350  ( .A1(_AES_ENC_us20_n591 ), .A2(_AES_ENC_us20_n581 ), .ZN(_AES_ENC_us20_n1010 ) );
NOR2_X2 _AES_ENC_us20_U349  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n1103 ) );
NOR2_X2 _AES_ENC_us20_U348  ( .A1(_AES_ENC_us20_n614 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n1059 ) );
NOR2_X2 _AES_ENC_us20_U347  ( .A1(_AES_ENC_sa20[1]), .A2(_AES_ENC_us20_n1120 ), .ZN(_AES_ENC_us20_n1022 ) );
NOR2_X2 _AES_ENC_us20_U346  ( .A1(_AES_ENC_us20_n605 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n911 ) );
NOR2_X2 _AES_ENC_us20_U345  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_us20_n1025 ), .ZN(_AES_ENC_us20_n826 ) );
NOR2_X2 _AES_ENC_us20_U338  ( .A1(_AES_ENC_us20_n596 ), .A2(_AES_ENC_us20_n588 ), .ZN(_AES_ENC_us20_n1072 ) );
NOR2_X2 _AES_ENC_us20_U335  ( .A1(_AES_ENC_us20_n581 ), .A2(_AES_ENC_us20_n594 ), .ZN(_AES_ENC_us20_n956 ) );
NOR2_X2 _AES_ENC_us20_U329  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_us20_n612 ), .ZN(_AES_ENC_us20_n1121 ) );
NOR2_X2 _AES_ENC_us20_U328  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_us20_n612 ), .ZN(_AES_ENC_us20_n1058 ) );
NOR2_X2 _AES_ENC_us20_U327  ( .A1(_AES_ENC_us20_n577 ), .A2(_AES_ENC_us20_n593 ), .ZN(_AES_ENC_us20_n1073 ) );
NOR2_X2 _AES_ENC_us20_U325  ( .A1(_AES_ENC_sa20[1]), .A2(_AES_ENC_us20_n1025 ), .ZN(_AES_ENC_us20_n1054 ) );
NOR2_X2 _AES_ENC_us20_U324  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_us20_n931 ), .ZN(_AES_ENC_us20_n1029 ) );
NOR2_X2 _AES_ENC_us20_U319  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n1056 ) );
NOR2_X2 _AES_ENC_us20_U318  ( .A1(_AES_ENC_us20_n585 ), .A2(_AES_ENC_us20_n596 ), .ZN(_AES_ENC_us20_n1050 ) );
NOR2_X2 _AES_ENC_us20_U317  ( .A1(_AES_ENC_us20_n1121 ), .A2(_AES_ENC_us20_n1025 ), .ZN(_AES_ENC_us20_n1120 ) );
NOR2_X2 _AES_ENC_us20_U316  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_us20_n572 ), .ZN(_AES_ENC_us20_n1074 ) );
NOR2_X2 _AES_ENC_us20_U315  ( .A1(_AES_ENC_us20_n1058 ), .A2(_AES_ENC_us20_n1054 ), .ZN(_AES_ENC_us20_n878 ) );
NOR2_X2 _AES_ENC_us20_U314  ( .A1(_AES_ENC_us20_n878 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n879 ) );
NOR2_X2 _AES_ENC_us20_U312  ( .A1(_AES_ENC_us20_n880 ), .A2(_AES_ENC_us20_n879 ), .ZN(_AES_ENC_us20_n887 ) );
NOR2_X2 _AES_ENC_us20_U311  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n625 ), .ZN(_AES_ENC_us20_n957 ) );
NOR2_X2 _AES_ENC_us20_U310  ( .A1(_AES_ENC_us20_n958 ), .A2(_AES_ENC_us20_n957 ), .ZN(_AES_ENC_us20_n965 ) );
NOR3_X2 _AES_ENC_us20_U309  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n1091 ), .A3(_AES_ENC_us20_n1022 ), .ZN(_AES_ENC_us20_n720 ) );
NOR3_X2 _AES_ENC_us20_U303  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n1054 ), .A3(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n719 ) );
NOR2_X2 _AES_ENC_us20_U302  ( .A1(_AES_ENC_us20_n720 ), .A2(_AES_ENC_us20_n719 ), .ZN(_AES_ENC_us20_n726 ) );
NOR2_X2 _AES_ENC_us20_U300  ( .A1(_AES_ENC_us20_n585 ), .A2(_AES_ENC_us20_n613 ), .ZN(_AES_ENC_us20_n865 ) );
NOR2_X2 _AES_ENC_us20_U299  ( .A1(_AES_ENC_us20_n1059 ), .A2(_AES_ENC_us20_n1058 ), .ZN(_AES_ENC_us20_n1060 ) );
NOR2_X2 _AES_ENC_us20_U298  ( .A1(_AES_ENC_us20_n1095 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n668 ) );
NOR2_X2 _AES_ENC_us20_U297  ( .A1(_AES_ENC_us20_n826 ), .A2(_AES_ENC_us20_n573 ), .ZN(_AES_ENC_us20_n750 ) );
NOR2_X2 _AES_ENC_us20_U296  ( .A1(_AES_ENC_us20_n750 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n751 ) );
NOR2_X2 _AES_ENC_us20_U295  ( .A1(_AES_ENC_us20_n907 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n908 ) );
NOR2_X2 _AES_ENC_us20_U294  ( .A1(_AES_ENC_us20_n990 ), .A2(_AES_ENC_us20_n926 ), .ZN(_AES_ENC_us20_n780 ) );
NOR2_X2 _AES_ENC_us20_U293  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n606 ), .ZN(_AES_ENC_us20_n838 ) );
NOR2_X2 _AES_ENC_us20_U292  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n621 ), .ZN(_AES_ENC_us20_n837 ) );
NOR2_X2 _AES_ENC_us20_U291  ( .A1(_AES_ENC_us20_n838 ), .A2(_AES_ENC_us20_n837 ), .ZN(_AES_ENC_us20_n845 ) );
NOR2_X2 _AES_ENC_us20_U290  ( .A1(_AES_ENC_us20_n1022 ), .A2(_AES_ENC_us20_n1058 ), .ZN(_AES_ENC_us20_n740 ) );
NOR2_X2 _AES_ENC_us20_U284  ( .A1(_AES_ENC_us20_n740 ), .A2(_AES_ENC_us20_n594 ), .ZN(_AES_ENC_us20_n742 ) );
NOR2_X2 _AES_ENC_us20_U283  ( .A1(_AES_ENC_us20_n1098 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n1099 ) );
NOR2_X2 _AES_ENC_us20_U282  ( .A1(_AES_ENC_us20_n1120 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n993 ) );
NOR2_X2 _AES_ENC_us20_U281  ( .A1(_AES_ENC_us20_n993 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n994 ) );
NOR2_X2 _AES_ENC_us20_U280  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n609 ), .ZN(_AES_ENC_us20_n1026 ) );
NOR2_X2 _AES_ENC_us20_U279  ( .A1(_AES_ENC_us20_n573 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n1027 ) );
NOR2_X2 _AES_ENC_us20_U273  ( .A1(_AES_ENC_us20_n1027 ), .A2(_AES_ENC_us20_n1026 ), .ZN(_AES_ENC_us20_n1028 ) );
NOR2_X2 _AES_ENC_us20_U272  ( .A1(_AES_ENC_us20_n1029 ), .A2(_AES_ENC_us20_n1028 ), .ZN(_AES_ENC_us20_n1034 ) );
NOR4_X2 _AES_ENC_us20_U271  ( .A1(_AES_ENC_us20_n757 ), .A2(_AES_ENC_us20_n756 ), .A3(_AES_ENC_us20_n755 ), .A4(_AES_ENC_us20_n754 ), .ZN(_AES_ENC_us20_n758 ) );
NOR2_X2 _AES_ENC_us20_U270  ( .A1(_AES_ENC_us20_n752 ), .A2(_AES_ENC_us20_n751 ), .ZN(_AES_ENC_us20_n759 ) );
NOR2_X2 _AES_ENC_us20_U269  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n1071 ), .ZN(_AES_ENC_us20_n669 ) );
NOR2_X2 _AES_ENC_us20_U268  ( .A1(_AES_ENC_us20_n1056 ), .A2(_AES_ENC_us20_n990 ), .ZN(_AES_ENC_us20_n991 ) );
NOR2_X2 _AES_ENC_us20_U267  ( .A1(_AES_ENC_us20_n991 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n995 ) );
NOR2_X2 _AES_ENC_us20_U263  ( .A1(_AES_ENC_us20_n588 ), .A2(_AES_ENC_us20_n598 ), .ZN(_AES_ENC_us20_n1008 ) );
NOR2_X2 _AES_ENC_us20_U262  ( .A1(_AES_ENC_us20_n839 ), .A2(_AES_ENC_us20_n603 ), .ZN(_AES_ENC_us20_n693 ) );
NOR2_X2 _AES_ENC_us20_U258  ( .A1(_AES_ENC_us20_n587 ), .A2(_AES_ENC_us20_n906 ), .ZN(_AES_ENC_us20_n741 ) );
NOR2_X2 _AES_ENC_us20_U255  ( .A1(_AES_ENC_us20_n1054 ), .A2(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n763 ) );
NOR2_X2 _AES_ENC_us20_U254  ( .A1(_AES_ENC_us20_n763 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n769 ) );
NOR2_X2 _AES_ENC_us20_U253  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n618 ), .ZN(_AES_ENC_us20_n1007 ) );
NOR2_X2 _AES_ENC_us20_U252  ( .A1(_AES_ENC_us20_n591 ), .A2(_AES_ENC_us20_n599 ), .ZN(_AES_ENC_us20_n1123 ) );
NOR2_X2 _AES_ENC_us20_U251  ( .A1(_AES_ENC_us20_n591 ), .A2(_AES_ENC_us20_n598 ), .ZN(_AES_ENC_us20_n710 ) );
INV_X4 _AES_ENC_us20_U250  ( .A(_AES_ENC_us20_n1029 ), .ZN(_AES_ENC_us20_n603 ) );
NOR2_X2 _AES_ENC_us20_U243  ( .A1(_AES_ENC_us20_n594 ), .A2(_AES_ENC_us20_n607 ), .ZN(_AES_ENC_us20_n883 ) );
NOR2_X2 _AES_ENC_us20_U242  ( .A1(_AES_ENC_us20_n623 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n1125 ) );
NOR2_X2 _AES_ENC_us20_U241  ( .A1(_AES_ENC_us20_n911 ), .A2(_AES_ENC_us20_n910 ), .ZN(_AES_ENC_us20_n912 ) );
NOR2_X2 _AES_ENC_us20_U240  ( .A1(_AES_ENC_us20_n912 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n916 ) );
NOR2_X2 _AES_ENC_us20_U239  ( .A1(_AES_ENC_us20_n990 ), .A2(_AES_ENC_us20_n929 ), .ZN(_AES_ENC_us20_n892 ) );
NOR2_X2 _AES_ENC_us20_U238  ( .A1(_AES_ENC_us20_n892 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n893 ) );
NOR2_X2 _AES_ENC_us20_U237  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n621 ), .ZN(_AES_ENC_us20_n950 ) );
NOR2_X2 _AES_ENC_us20_U236  ( .A1(_AES_ENC_us20_n1079 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n1082 ) );
NOR2_X2 _AES_ENC_us20_U235  ( .A1(_AES_ENC_us20_n910 ), .A2(_AES_ENC_us20_n1056 ), .ZN(_AES_ENC_us20_n941 ) );
NOR2_X2 _AES_ENC_us20_U234  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n1077 ), .ZN(_AES_ENC_us20_n841 ) );
NOR2_X2 _AES_ENC_us20_U229  ( .A1(_AES_ENC_us20_n601 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n630 ) );
NOR2_X2 _AES_ENC_us20_U228  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n621 ), .ZN(_AES_ENC_us20_n806 ) );
NOR2_X2 _AES_ENC_us20_U227  ( .A1(_AES_ENC_us20_n601 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n948 ) );
NOR2_X2 _AES_ENC_us20_U226  ( .A1(_AES_ENC_us20_n587 ), .A2(_AES_ENC_us20_n620 ), .ZN(_AES_ENC_us20_n997 ) );
NOR2_X2 _AES_ENC_us20_U225  ( .A1(_AES_ENC_us20_n1121 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n1122 ) );
NOR2_X2 _AES_ENC_us20_U223  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n1023 ), .ZN(_AES_ENC_us20_n756 ) );
NOR2_X2 _AES_ENC_us20_U222  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n621 ), .ZN(_AES_ENC_us20_n870 ) );
NOR2_X2 _AES_ENC_us20_U221  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n569 ), .ZN(_AES_ENC_us20_n947 ) );
NOR2_X2 _AES_ENC_us20_U217  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n1077 ), .ZN(_AES_ENC_us20_n1084 ) );
NOR2_X2 _AES_ENC_us20_U213  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n855 ), .ZN(_AES_ENC_us20_n709 ) );
NOR2_X2 _AES_ENC_us20_U212  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n620 ), .ZN(_AES_ENC_us20_n868 ) );
NOR2_X2 _AES_ENC_us20_U211  ( .A1(_AES_ENC_us20_n1120 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n1124 ) );
NOR2_X2 _AES_ENC_us20_U210  ( .A1(_AES_ENC_us20_n1120 ), .A2(_AES_ENC_us20_n839 ), .ZN(_AES_ENC_us20_n842 ) );
NOR2_X2 _AES_ENC_us20_U209  ( .A1(_AES_ENC_us20_n1120 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n696 ) );
NOR2_X2 _AES_ENC_us20_U208  ( .A1(_AES_ENC_us20_n1074 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n1076 ) );
NOR2_X2 _AES_ENC_us20_U207  ( .A1(_AES_ENC_us20_n1074 ), .A2(_AES_ENC_us20_n609 ), .ZN(_AES_ENC_us20_n781 ) );
NOR3_X2 _AES_ENC_us20_U201  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n1056 ), .A3(_AES_ENC_us20_n990 ), .ZN(_AES_ENC_us20_n979 ) );
NOR3_X2 _AES_ENC_us20_U200  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n1058 ), .A3(_AES_ENC_us20_n1059 ), .ZN(_AES_ENC_us20_n854 ) );
NOR2_X2 _AES_ENC_us20_U199  ( .A1(_AES_ENC_us20_n996 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n869 ) );
NOR2_X2 _AES_ENC_us20_U198  ( .A1(_AES_ENC_us20_n1056 ), .A2(_AES_ENC_us20_n1074 ), .ZN(_AES_ENC_us20_n1057 ) );
NOR3_X2 _AES_ENC_us20_U197  ( .A1(_AES_ENC_us20_n588 ), .A2(_AES_ENC_us20_n1120 ), .A3(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n978 ) );
NOR2_X2 _AES_ENC_us20_U196  ( .A1(_AES_ENC_us20_n996 ), .A2(_AES_ENC_us20_n911 ), .ZN(_AES_ENC_us20_n1116 ) );
NOR2_X2 _AES_ENC_us20_U195  ( .A1(_AES_ENC_us20_n1074 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n754 ) );
NOR2_X2 _AES_ENC_us20_U194  ( .A1(_AES_ENC_us20_n926 ), .A2(_AES_ENC_us20_n1103 ), .ZN(_AES_ENC_us20_n977 ) );
NOR2_X2 _AES_ENC_us20_U187  ( .A1(_AES_ENC_us20_n839 ), .A2(_AES_ENC_us20_n824 ), .ZN(_AES_ENC_us20_n1092 ) );
NOR2_X2 _AES_ENC_us20_U186  ( .A1(_AES_ENC_us20_n573 ), .A2(_AES_ENC_us20_n1074 ), .ZN(_AES_ENC_us20_n684 ) );
NOR2_X2 _AES_ENC_us20_U185  ( .A1(_AES_ENC_us20_n826 ), .A2(_AES_ENC_us20_n1059 ), .ZN(_AES_ENC_us20_n907 ) );
NOR3_X2 _AES_ENC_us20_U184  ( .A1(_AES_ENC_us20_n577 ), .A2(_AES_ENC_us20_n1115 ), .A3(_AES_ENC_us20_n600 ), .ZN(_AES_ENC_us20_n831 ) );
NOR3_X2 _AES_ENC_us20_U183  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n1056 ), .A3(_AES_ENC_us20_n990 ), .ZN(_AES_ENC_us20_n896 ) );
NOR3_X2 _AES_ENC_us20_U182  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n573 ), .A3(_AES_ENC_us20_n1013 ), .ZN(_AES_ENC_us20_n670 ) );
NOR3_X2 _AES_ENC_us20_U181  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n1091 ), .A3(_AES_ENC_us20_n1022 ), .ZN(_AES_ENC_us20_n843 ) );
NOR2_X2 _AES_ENC_us20_U180  ( .A1(_AES_ENC_us20_n1029 ), .A2(_AES_ENC_us20_n1095 ), .ZN(_AES_ENC_us20_n735 ) );
NOR2_X2 _AES_ENC_us20_U174  ( .A1(_AES_ENC_us20_n1100 ), .A2(_AES_ENC_us20_n854 ), .ZN(_AES_ENC_us20_n860 ) );
NAND3_X2 _AES_ENC_us20_U173  ( .A1(_AES_ENC_us20_n569 ), .A2(_AES_ENC_us20_n603 ), .A3(_AES_ENC_us20_n681 ), .ZN(_AES_ENC_us20_n691 ) );
NOR2_X2 _AES_ENC_us20_U172  ( .A1(_AES_ENC_us20_n683 ), .A2(_AES_ENC_us20_n682 ), .ZN(_AES_ENC_us20_n690 ) );
NOR3_X2 _AES_ENC_us20_U171  ( .A1(_AES_ENC_us20_n695 ), .A2(_AES_ENC_us20_n694 ), .A3(_AES_ENC_us20_n693 ), .ZN(_AES_ENC_us20_n700 ) );
NOR4_X2 _AES_ENC_us20_U170  ( .A1(_AES_ENC_us20_n983 ), .A2(_AES_ENC_us20_n698 ), .A3(_AES_ENC_us20_n697 ), .A4(_AES_ENC_us20_n696 ), .ZN(_AES_ENC_us20_n699 ) );
NOR2_X2 _AES_ENC_us20_U169  ( .A1(_AES_ENC_us20_n946 ), .A2(_AES_ENC_us20_n945 ), .ZN(_AES_ENC_us20_n952 ) );
NOR4_X2 _AES_ENC_us20_U168  ( .A1(_AES_ENC_us20_n950 ), .A2(_AES_ENC_us20_n949 ), .A3(_AES_ENC_us20_n948 ), .A4(_AES_ENC_us20_n947 ), .ZN(_AES_ENC_us20_n951 ) );
NOR4_X2 _AES_ENC_us20_U162  ( .A1(_AES_ENC_us20_n896 ), .A2(_AES_ENC_us20_n895 ), .A3(_AES_ENC_us20_n894 ), .A4(_AES_ENC_us20_n893 ), .ZN(_AES_ENC_us20_n897 ) );
NOR2_X2 _AES_ENC_us20_U161  ( .A1(_AES_ENC_us20_n866 ), .A2(_AES_ENC_us20_n865 ), .ZN(_AES_ENC_us20_n872 ) );
NOR4_X2 _AES_ENC_us20_U160  ( .A1(_AES_ENC_us20_n870 ), .A2(_AES_ENC_us20_n869 ), .A3(_AES_ENC_us20_n868 ), .A4(_AES_ENC_us20_n867 ), .ZN(_AES_ENC_us20_n871 ) );
NOR4_X2 _AES_ENC_us20_U159  ( .A1(_AES_ENC_us20_n983 ), .A2(_AES_ENC_us20_n982 ), .A3(_AES_ENC_us20_n981 ), .A4(_AES_ENC_us20_n980 ), .ZN(_AES_ENC_us20_n984 ) );
NOR2_X2 _AES_ENC_us20_U158  ( .A1(_AES_ENC_us20_n979 ), .A2(_AES_ENC_us20_n978 ), .ZN(_AES_ENC_us20_n985 ) );
NOR4_X2 _AES_ENC_us20_U157  ( .A1(_AES_ENC_us20_n1125 ), .A2(_AES_ENC_us20_n1124 ), .A3(_AES_ENC_us20_n1123 ), .A4(_AES_ENC_us20_n1122 ), .ZN(_AES_ENC_us20_n1126 ) );
NOR4_X2 _AES_ENC_us20_U156  ( .A1(_AES_ENC_us20_n1084 ), .A2(_AES_ENC_us20_n1083 ), .A3(_AES_ENC_us20_n1082 ), .A4(_AES_ENC_us20_n1081 ), .ZN(_AES_ENC_us20_n1085 ) );
NOR2_X2 _AES_ENC_us20_U155  ( .A1(_AES_ENC_us20_n1076 ), .A2(_AES_ENC_us20_n1075 ), .ZN(_AES_ENC_us20_n1086 ) );
NOR3_X2 _AES_ENC_us20_U154  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n1054 ), .A3(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n961 ) );
NOR3_X2 _AES_ENC_us20_U153  ( .A1(_AES_ENC_us20_n609 ), .A2(_AES_ENC_us20_n1074 ), .A3(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n671 ) );
NOR2_X2 _AES_ENC_us20_U152  ( .A1(_AES_ENC_us20_n1057 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n1062 ) );
NOR2_X2 _AES_ENC_us20_U143  ( .A1(_AES_ENC_us20_n1055 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n1063 ) );
NOR2_X2 _AES_ENC_us20_U142  ( .A1(_AES_ENC_us20_n1060 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n1061 ) );
NOR4_X2 _AES_ENC_us20_U141  ( .A1(_AES_ENC_us20_n1064 ), .A2(_AES_ENC_us20_n1063 ), .A3(_AES_ENC_us20_n1062 ), .A4(_AES_ENC_us20_n1061 ), .ZN(_AES_ENC_us20_n1065 ) );
NOR3_X2 _AES_ENC_us20_U140  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n1120 ), .A3(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n918 ) );
NOR3_X2 _AES_ENC_us20_U132  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n573 ), .A3(_AES_ENC_us20_n1013 ), .ZN(_AES_ENC_us20_n917 ) );
NOR2_X2 _AES_ENC_us20_U131  ( .A1(_AES_ENC_us20_n914 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n915 ) );
NOR4_X2 _AES_ENC_us20_U130  ( .A1(_AES_ENC_us20_n918 ), .A2(_AES_ENC_us20_n917 ), .A3(_AES_ENC_us20_n916 ), .A4(_AES_ENC_us20_n915 ), .ZN(_AES_ENC_us20_n919 ) );
NOR2_X2 _AES_ENC_us20_U129  ( .A1(_AES_ENC_us20_n594 ), .A2(_AES_ENC_us20_n599 ), .ZN(_AES_ENC_us20_n771 ) );
NOR2_X2 _AES_ENC_us20_U128  ( .A1(_AES_ENC_us20_n1103 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n772 ) );
NOR2_X2 _AES_ENC_us20_U127  ( .A1(_AES_ENC_us20_n592 ), .A2(_AES_ENC_us20_n615 ), .ZN(_AES_ENC_us20_n773 ) );
NOR4_X2 _AES_ENC_us20_U126  ( .A1(_AES_ENC_us20_n773 ), .A2(_AES_ENC_us20_n772 ), .A3(_AES_ENC_us20_n771 ), .A4(_AES_ENC_us20_n770 ), .ZN(_AES_ENC_us20_n774 ) );
NOR2_X2 _AES_ENC_us20_U121  ( .A1(_AES_ENC_us20_n735 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n687 ) );
NOR2_X2 _AES_ENC_us20_U120  ( .A1(_AES_ENC_us20_n684 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n688 ) );
NOR2_X2 _AES_ENC_us20_U119  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n622 ), .ZN(_AES_ENC_us20_n686 ) );
NOR4_X2 _AES_ENC_us20_U118  ( .A1(_AES_ENC_us20_n688 ), .A2(_AES_ENC_us20_n687 ), .A3(_AES_ENC_us20_n686 ), .A4(_AES_ENC_us20_n685 ), .ZN(_AES_ENC_us20_n689 ) );
NOR2_X2 _AES_ENC_us20_U117  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n608 ), .ZN(_AES_ENC_us20_n858 ) );
NOR2_X2 _AES_ENC_us20_U116  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n855 ), .ZN(_AES_ENC_us20_n857 ) );
NOR2_X2 _AES_ENC_us20_U115  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n617 ), .ZN(_AES_ENC_us20_n856 ) );
NOR4_X2 _AES_ENC_us20_U106  ( .A1(_AES_ENC_us20_n858 ), .A2(_AES_ENC_us20_n857 ), .A3(_AES_ENC_us20_n856 ), .A4(_AES_ENC_us20_n958 ), .ZN(_AES_ENC_us20_n859 ) );
NOR2_X2 _AES_ENC_us20_U105  ( .A1(_AES_ENC_us20_n780 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n784 ) );
NOR2_X2 _AES_ENC_us20_U104  ( .A1(_AES_ENC_us20_n1117 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n782 ) );
NOR2_X2 _AES_ENC_us20_U103  ( .A1(_AES_ENC_us20_n781 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n783 ) );
NOR4_X2 _AES_ENC_us20_U102  ( .A1(_AES_ENC_us20_n880 ), .A2(_AES_ENC_us20_n784 ), .A3(_AES_ENC_us20_n783 ), .A4(_AES_ENC_us20_n782 ), .ZN(_AES_ENC_us20_n785 ) );
NOR2_X2 _AES_ENC_us20_U101  ( .A1(_AES_ENC_us20_n597 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n814 ) );
NOR2_X2 _AES_ENC_us20_U100  ( .A1(_AES_ENC_us20_n907 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n813 ) );
NOR3_X2 _AES_ENC_us20_U95  ( .A1(_AES_ENC_us20_n587 ), .A2(_AES_ENC_us20_n1058 ), .A3(_AES_ENC_us20_n1059 ), .ZN(_AES_ENC_us20_n815 ) );
NOR4_X2 _AES_ENC_us20_U94  ( .A1(_AES_ENC_us20_n815 ), .A2(_AES_ENC_us20_n814 ), .A3(_AES_ENC_us20_n813 ), .A4(_AES_ENC_us20_n812 ), .ZN(_AES_ENC_us20_n816 ) );
NOR2_X2 _AES_ENC_us20_U93  ( .A1(_AES_ENC_us20_n575 ), .A2(_AES_ENC_us20_n569 ), .ZN(_AES_ENC_us20_n721 ) );
NOR2_X2 _AES_ENC_us20_U92  ( .A1(_AES_ENC_us20_n1031 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n723 ) );
NOR2_X2 _AES_ENC_us20_U91  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n1096 ), .ZN(_AES_ENC_us20_n722 ) );
NOR4_X2 _AES_ENC_us20_U90  ( .A1(_AES_ENC_us20_n724 ), .A2(_AES_ENC_us20_n723 ), .A3(_AES_ENC_us20_n722 ), .A4(_AES_ENC_us20_n721 ), .ZN(_AES_ENC_us20_n725 ) );
NOR2_X2 _AES_ENC_us20_U89  ( .A1(_AES_ENC_us20_n911 ), .A2(_AES_ENC_us20_n990 ), .ZN(_AES_ENC_us20_n1009 ) );
NOR2_X2 _AES_ENC_us20_U88  ( .A1(_AES_ENC_us20_n1013 ), .A2(_AES_ENC_us20_n573 ), .ZN(_AES_ENC_us20_n1014 ) );
NOR2_X2 _AES_ENC_us20_U87  ( .A1(_AES_ENC_us20_n1014 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n1015 ) );
NOR4_X2 _AES_ENC_us20_U86  ( .A1(_AES_ENC_us20_n1016 ), .A2(_AES_ENC_us20_n1015 ), .A3(_AES_ENC_us20_n1119 ), .A4(_AES_ENC_us20_n1046 ), .ZN(_AES_ENC_us20_n1017 ) );
NOR2_X2 _AES_ENC_us20_U81  ( .A1(_AES_ENC_us20_n996 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n998 ) );
NOR2_X2 _AES_ENC_us20_U80  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n618 ), .ZN(_AES_ENC_us20_n1000 ) );
NOR2_X2 _AES_ENC_us20_U79  ( .A1(_AES_ENC_us20_n594 ), .A2(_AES_ENC_us20_n1096 ), .ZN(_AES_ENC_us20_n999 ) );
NOR4_X2 _AES_ENC_us20_U78  ( .A1(_AES_ENC_us20_n1000 ), .A2(_AES_ENC_us20_n999 ), .A3(_AES_ENC_us20_n998 ), .A4(_AES_ENC_us20_n997 ), .ZN(_AES_ENC_us20_n1001 ) );
NOR2_X2 _AES_ENC_us20_U74  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n1096 ), .ZN(_AES_ENC_us20_n697 ) );
NOR2_X2 _AES_ENC_us20_U73  ( .A1(_AES_ENC_us20_n609 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n958 ) );
NOR2_X2 _AES_ENC_us20_U72  ( .A1(_AES_ENC_us20_n911 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n983 ) );
NOR2_X2 _AES_ENC_us20_U71  ( .A1(_AES_ENC_us20_n1054 ), .A2(_AES_ENC_us20_n1103 ), .ZN(_AES_ENC_us20_n1031 ) );
INV_X4 _AES_ENC_us20_U65  ( .A(_AES_ENC_us20_n1050 ), .ZN(_AES_ENC_us20_n582 ) );
INV_X4 _AES_ENC_us20_U64  ( .A(_AES_ENC_us20_n1072 ), .ZN(_AES_ENC_us20_n586 ) );
INV_X4 _AES_ENC_us20_U63  ( .A(_AES_ENC_us20_n1073 ), .ZN(_AES_ENC_us20_n576 ) );
NOR2_X2 _AES_ENC_us20_U62  ( .A1(_AES_ENC_us20_n603 ), .A2(_AES_ENC_us20_n584 ), .ZN(_AES_ENC_us20_n880 ) );
NOR3_X2 _AES_ENC_us20_U61  ( .A1(_AES_ENC_us20_n826 ), .A2(_AES_ENC_us20_n1121 ), .A3(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n946 ) );
INV_X4 _AES_ENC_us20_U59  ( .A(_AES_ENC_us20_n1010 ), .ZN(_AES_ENC_us20_n579 ) );
NOR3_X2 _AES_ENC_us20_U58  ( .A1(_AES_ENC_us20_n573 ), .A2(_AES_ENC_us20_n1029 ), .A3(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n1119 ) );
INV_X4 _AES_ENC_us20_U57  ( .A(_AES_ENC_us20_n956 ), .ZN(_AES_ENC_us20_n580 ) );
NOR2_X2 _AES_ENC_us20_U50  ( .A1(_AES_ENC_us20_n601 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n1013 ) );
NOR2_X2 _AES_ENC_us20_U49  ( .A1(_AES_ENC_us20_n609 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n910 ) );
NOR2_X2 _AES_ENC_us20_U48  ( .A1(_AES_ENC_us20_n569 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n1091 ) );
NOR2_X2 _AES_ENC_us20_U47  ( .A1(_AES_ENC_us20_n614 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n990 ) );
NOR2_X2 _AES_ENC_us20_U46  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_us20_n1121 ), .ZN(_AES_ENC_us20_n996 ) );
NOR2_X2 _AES_ENC_us20_U45  ( .A1(_AES_ENC_us20_n592 ), .A2(_AES_ENC_us20_n622 ), .ZN(_AES_ENC_us20_n628 ) );
NOR2_X2 _AES_ENC_us20_U44  ( .A1(_AES_ENC_us20_n602 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n866 ) );
NOR2_X2 _AES_ENC_us20_U43  ( .A1(_AES_ENC_us20_n610 ), .A2(_AES_ENC_us20_n592 ), .ZN(_AES_ENC_us20_n1006 ) );
NOR2_X2 _AES_ENC_us20_U42  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n1117 ), .ZN(_AES_ENC_us20_n1118 ) );
NOR2_X2 _AES_ENC_us20_U41  ( .A1(_AES_ENC_us20_n1119 ), .A2(_AES_ENC_us20_n1118 ), .ZN(_AES_ENC_us20_n1127 ) );
NOR2_X2 _AES_ENC_us20_U36  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n616 ), .ZN(_AES_ENC_us20_n629 ) );
NOR2_X2 _AES_ENC_us20_U35  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n906 ), .ZN(_AES_ENC_us20_n909 ) );
NOR2_X2 _AES_ENC_us20_U34  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n607 ), .ZN(_AES_ENC_us20_n658 ) );
NOR2_X2 _AES_ENC_us20_U33  ( .A1(_AES_ENC_us20_n1116 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n695 ) );
NOR2_X2 _AES_ENC_us20_U32  ( .A1(_AES_ENC_us20_n1078 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n1083 ) );
NOR2_X2 _AES_ENC_us20_U31  ( .A1(_AES_ENC_us20_n941 ), .A2(_AES_ENC_us20_n579 ), .ZN(_AES_ENC_us20_n724 ) );
NOR2_X2 _AES_ENC_us20_U30  ( .A1(_AES_ENC_us20_n611 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n1107 ) );
NOR2_X2 _AES_ENC_us20_U29  ( .A1(_AES_ENC_us20_n602 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n840 ) );
NOR2_X2 _AES_ENC_us20_U24  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n623 ), .ZN(_AES_ENC_us20_n633 ) );
NOR2_X2 _AES_ENC_us20_U23  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n1080 ), .ZN(_AES_ENC_us20_n1081 ) );
NOR2_X2 _AES_ENC_us20_U21  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n1045 ), .ZN(_AES_ENC_us20_n812 ) );
NOR2_X2 _AES_ENC_us20_U20  ( .A1(_AES_ENC_us20_n1009 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n960 ) );
NOR2_X2 _AES_ENC_us20_U19  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n619 ), .ZN(_AES_ENC_us20_n982 ) );
NOR2_X2 _AES_ENC_us20_U18  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n616 ), .ZN(_AES_ENC_us20_n757 ) );
NOR2_X2 _AES_ENC_us20_U17  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n598 ), .ZN(_AES_ENC_us20_n698 ) );
NOR2_X2 _AES_ENC_us20_U16  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n605 ), .ZN(_AES_ENC_us20_n708 ) );
NOR2_X2 _AES_ENC_us20_U15  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n603 ), .ZN(_AES_ENC_us20_n770 ) );
NOR2_X2 _AES_ENC_us20_U10  ( .A1(_AES_ENC_us20_n605 ), .A2(_AES_ENC_us20_n576 ), .ZN(_AES_ENC_us20_n803 ) );
NOR2_X2 _AES_ENC_us20_U9  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n881 ), .ZN(_AES_ENC_us20_n711 ) );
NOR2_X2 _AES_ENC_us20_U8  ( .A1(_AES_ENC_us20_n580 ), .A2(_AES_ENC_us20_n603 ), .ZN(_AES_ENC_us20_n867 ) );
NOR2_X2 _AES_ENC_us20_U7  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n615 ), .ZN(_AES_ENC_us20_n804 ) );
NOR2_X2 _AES_ENC_us20_U6  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n609 ), .ZN(_AES_ENC_us20_n1046 ) );
OR2_X4 _AES_ENC_us20_U5  ( .A1(_AES_ENC_us20_n612 ), .A2(_AES_ENC_sa20[1]),.ZN(_AES_ENC_us20_n570 ) );
OR2_X4 _AES_ENC_us20_U4  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_sa20[4]),.ZN(_AES_ENC_us20_n569 ) );
NAND2_X2 _AES_ENC_us20_U514  ( .A1(_AES_ENC_us20_n1121 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n1030 ) );
AND2_X2 _AES_ENC_us20_U513  ( .A1(_AES_ENC_us20_n607 ), .A2(_AES_ENC_us20_n1030 ), .ZN(_AES_ENC_us20_n1049 ) );
NAND2_X2 _AES_ENC_us20_U511  ( .A1(_AES_ENC_us20_n1049 ), .A2(_AES_ENC_us20_n794 ), .ZN(_AES_ENC_us20_n637 ) );
AND2_X2 _AES_ENC_us20_U493  ( .A1(_AES_ENC_us20_n779 ), .A2(_AES_ENC_us20_n996 ), .ZN(_AES_ENC_us20_n632 ) );
NAND4_X2 _AES_ENC_us20_U485  ( .A1(_AES_ENC_us20_n637 ), .A2(_AES_ENC_us20_n636 ), .A3(_AES_ENC_us20_n635 ), .A4(_AES_ENC_us20_n634 ), .ZN(_AES_ENC_us20_n638 ) );
NAND2_X2 _AES_ENC_us20_U484  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n638 ), .ZN(_AES_ENC_us20_n679 ) );
NAND2_X2 _AES_ENC_us20_U481  ( .A1(_AES_ENC_us20_n1094 ), .A2(_AES_ENC_us20_n613 ), .ZN(_AES_ENC_us20_n648 ) );
NAND2_X2 _AES_ENC_us20_U476  ( .A1(_AES_ENC_us20_n619 ), .A2(_AES_ENC_us20_n598 ), .ZN(_AES_ENC_us20_n762 ) );
NAND2_X2 _AES_ENC_us20_U475  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n762 ), .ZN(_AES_ENC_us20_n647 ) );
NAND4_X2 _AES_ENC_us20_U457  ( .A1(_AES_ENC_us20_n648 ), .A2(_AES_ENC_us20_n647 ), .A3(_AES_ENC_us20_n646 ), .A4(_AES_ENC_us20_n645 ), .ZN(_AES_ENC_us20_n649 ) );
NAND2_X2 _AES_ENC_us20_U456  ( .A1(_AES_ENC_sa20[0]), .A2(_AES_ENC_us20_n649 ), .ZN(_AES_ENC_us20_n665 ) );
NAND2_X2 _AES_ENC_us20_U454  ( .A1(_AES_ENC_us20_n626 ), .A2(_AES_ENC_us20_n601 ), .ZN(_AES_ENC_us20_n855 ) );
NAND2_X2 _AES_ENC_us20_U453  ( .A1(_AES_ENC_us20_n617 ), .A2(_AES_ENC_us20_n855 ), .ZN(_AES_ENC_us20_n821 ) );
NAND2_X2 _AES_ENC_us20_U452  ( .A1(_AES_ENC_us20_n1093 ), .A2(_AES_ENC_us20_n821 ), .ZN(_AES_ENC_us20_n662 ) );
NAND2_X2 _AES_ENC_us20_U451  ( .A1(_AES_ENC_us20_n605 ), .A2(_AES_ENC_us20_n620 ), .ZN(_AES_ENC_us20_n650 ) );
NAND2_X2 _AES_ENC_us20_U450  ( .A1(_AES_ENC_us20_n956 ), .A2(_AES_ENC_us20_n650 ), .ZN(_AES_ENC_us20_n661 ) );
NAND2_X2 _AES_ENC_us20_U449  ( .A1(_AES_ENC_us20_n596 ), .A2(_AES_ENC_us20_n581 ), .ZN(_AES_ENC_us20_n839 ) );
OR2_X2 _AES_ENC_us20_U446  ( .A1(_AES_ENC_us20_n839 ), .A2(_AES_ENC_us20_n932 ), .ZN(_AES_ENC_us20_n656 ) );
NAND2_X2 _AES_ENC_us20_U445  ( .A1(_AES_ENC_us20_n624 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n1096 ) );
NAND2_X2 _AES_ENC_us20_U444  ( .A1(_AES_ENC_us20_n1030 ), .A2(_AES_ENC_us20_n1096 ), .ZN(_AES_ENC_us20_n651 ) );
NAND2_X2 _AES_ENC_us20_U443  ( .A1(_AES_ENC_us20_n1114 ), .A2(_AES_ENC_us20_n651 ), .ZN(_AES_ENC_us20_n655 ) );
OR3_X2 _AES_ENC_us20_U440  ( .A1(_AES_ENC_us20_n1079 ), .A2(_AES_ENC_sa20[7]), .A3(_AES_ENC_us20_n596 ), .ZN(_AES_ENC_us20_n654 ));
NAND2_X2 _AES_ENC_us20_U439  ( .A1(_AES_ENC_us20_n623 ), .A2(_AES_ENC_us20_n619 ), .ZN(_AES_ENC_us20_n652 ) );
NAND4_X2 _AES_ENC_us20_U437  ( .A1(_AES_ENC_us20_n656 ), .A2(_AES_ENC_us20_n655 ), .A3(_AES_ENC_us20_n654 ), .A4(_AES_ENC_us20_n653 ), .ZN(_AES_ENC_us20_n657 ) );
NAND2_X2 _AES_ENC_us20_U436  ( .A1(_AES_ENC_sa20[2]), .A2(_AES_ENC_us20_n657 ), .ZN(_AES_ENC_us20_n660 ) );
NAND4_X2 _AES_ENC_us20_U432  ( .A1(_AES_ENC_us20_n662 ), .A2(_AES_ENC_us20_n661 ), .A3(_AES_ENC_us20_n660 ), .A4(_AES_ENC_us20_n659 ), .ZN(_AES_ENC_us20_n663 ) );
NAND2_X2 _AES_ENC_us20_U431  ( .A1(_AES_ENC_us20_n663 ), .A2(_AES_ENC_us20_n627 ), .ZN(_AES_ENC_us20_n664 ) );
NAND2_X2 _AES_ENC_us20_U430  ( .A1(_AES_ENC_us20_n665 ), .A2(_AES_ENC_us20_n664 ), .ZN(_AES_ENC_us20_n666 ) );
NAND2_X2 _AES_ENC_us20_U429  ( .A1(_AES_ENC_sa20[6]), .A2(_AES_ENC_us20_n666 ), .ZN(_AES_ENC_us20_n678 ) );
NAND2_X2 _AES_ENC_us20_U426  ( .A1(_AES_ENC_us20_n735 ), .A2(_AES_ENC_us20_n1093 ), .ZN(_AES_ENC_us20_n675 ) );
NAND2_X2 _AES_ENC_us20_U425  ( .A1(_AES_ENC_us20_n625 ), .A2(_AES_ENC_us20_n607 ), .ZN(_AES_ENC_us20_n1045 ) );
OR2_X2 _AES_ENC_us20_U424  ( .A1(_AES_ENC_us20_n1045 ), .A2(_AES_ENC_us20_n586 ), .ZN(_AES_ENC_us20_n674 ) );
NAND2_X2 _AES_ENC_us20_U423  ( .A1(_AES_ENC_sa20[1]), .A2(_AES_ENC_us20_n609 ), .ZN(_AES_ENC_us20_n667 ) );
NAND2_X2 _AES_ENC_us20_U422  ( .A1(_AES_ENC_us20_n605 ), .A2(_AES_ENC_us20_n667 ), .ZN(_AES_ENC_us20_n1071 ) );
NAND4_X2 _AES_ENC_us20_U412  ( .A1(_AES_ENC_us20_n675 ), .A2(_AES_ENC_us20_n674 ), .A3(_AES_ENC_us20_n673 ), .A4(_AES_ENC_us20_n672 ), .ZN(_AES_ENC_us20_n676 ) );
NAND2_X2 _AES_ENC_us20_U411  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n676 ), .ZN(_AES_ENC_us20_n677 ) );
NAND2_X2 _AES_ENC_us20_U408  ( .A1(_AES_ENC_us20_n800 ), .A2(_AES_ENC_us20_n1022 ), .ZN(_AES_ENC_us20_n680 ) );
NAND2_X2 _AES_ENC_us20_U407  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n680 ), .ZN(_AES_ENC_us20_n681 ) );
AND2_X2 _AES_ENC_us20_U402  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n684 ), .ZN(_AES_ENC_us20_n682 ) );
NAND4_X2 _AES_ENC_us20_U395  ( .A1(_AES_ENC_us20_n691 ), .A2(_AES_ENC_us20_n583 ), .A3(_AES_ENC_us20_n690 ), .A4(_AES_ENC_us20_n689 ), .ZN(_AES_ENC_us20_n692 ) );
NAND2_X2 _AES_ENC_us20_U394  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n692 ), .ZN(_AES_ENC_us20_n733 ) );
NAND2_X2 _AES_ENC_us20_U392  ( .A1(_AES_ENC_us20_n977 ), .A2(_AES_ENC_us20_n1050 ), .ZN(_AES_ENC_us20_n702 ) );
NAND2_X2 _AES_ENC_us20_U391  ( .A1(_AES_ENC_us20_n1093 ), .A2(_AES_ENC_us20_n1045 ), .ZN(_AES_ENC_us20_n701 ) );
NAND4_X2 _AES_ENC_us20_U381  ( .A1(_AES_ENC_us20_n702 ), .A2(_AES_ENC_us20_n701 ), .A3(_AES_ENC_us20_n700 ), .A4(_AES_ENC_us20_n699 ), .ZN(_AES_ENC_us20_n703 ) );
NAND2_X2 _AES_ENC_us20_U380  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n703 ), .ZN(_AES_ENC_us20_n732 ) );
AND2_X2 _AES_ENC_us20_U379  ( .A1(_AES_ENC_sa20[0]), .A2(_AES_ENC_sa20[6]),.ZN(_AES_ENC_us20_n1113 ) );
NAND2_X2 _AES_ENC_us20_U378  ( .A1(_AES_ENC_us20_n619 ), .A2(_AES_ENC_us20_n1030 ), .ZN(_AES_ENC_us20_n881 ) );
NAND2_X2 _AES_ENC_us20_U377  ( .A1(_AES_ENC_us20_n1093 ), .A2(_AES_ENC_us20_n881 ), .ZN(_AES_ENC_us20_n715 ) );
NAND2_X2 _AES_ENC_us20_U376  ( .A1(_AES_ENC_us20_n1010 ), .A2(_AES_ENC_us20_n622 ), .ZN(_AES_ENC_us20_n714 ) );
NAND2_X2 _AES_ENC_us20_U375  ( .A1(_AES_ENC_us20_n855 ), .A2(_AES_ENC_us20_n625 ), .ZN(_AES_ENC_us20_n1117 ) );
XNOR2_X2 _AES_ENC_us20_U371  ( .A(_AES_ENC_us20_n593 ), .B(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n824 ) );
NAND4_X2 _AES_ENC_us20_U362  ( .A1(_AES_ENC_us20_n715 ), .A2(_AES_ENC_us20_n714 ), .A3(_AES_ENC_us20_n713 ), .A4(_AES_ENC_us20_n712 ), .ZN(_AES_ENC_us20_n716 ) );
NAND2_X2 _AES_ENC_us20_U361  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n716 ), .ZN(_AES_ENC_us20_n731 ) );
AND2_X2 _AES_ENC_us20_U360  ( .A1(_AES_ENC_sa20[6]), .A2(_AES_ENC_us20_n627 ), .ZN(_AES_ENC_us20_n1131 ) );
NAND2_X2 _AES_ENC_us20_U359  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n717 ) );
NAND2_X2 _AES_ENC_us20_U358  ( .A1(_AES_ENC_us20_n1029 ), .A2(_AES_ENC_us20_n717 ), .ZN(_AES_ENC_us20_n728 ) );
NAND2_X2 _AES_ENC_us20_U357  ( .A1(_AES_ENC_sa20[1]), .A2(_AES_ENC_us20_n612 ), .ZN(_AES_ENC_us20_n1097 ) );
NAND2_X2 _AES_ENC_us20_U356  ( .A1(_AES_ENC_us20_n610 ), .A2(_AES_ENC_us20_n1097 ), .ZN(_AES_ENC_us20_n718 ) );
NAND2_X2 _AES_ENC_us20_U355  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n718 ), .ZN(_AES_ENC_us20_n727 ) );
NAND4_X2 _AES_ENC_us20_U344  ( .A1(_AES_ENC_us20_n728 ), .A2(_AES_ENC_us20_n727 ), .A3(_AES_ENC_us20_n726 ), .A4(_AES_ENC_us20_n725 ), .ZN(_AES_ENC_us20_n729 ) );
NAND2_X2 _AES_ENC_us20_U343  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n729 ), .ZN(_AES_ENC_us20_n730 ) );
NAND4_X2 _AES_ENC_us20_U342  ( .A1(_AES_ENC_us20_n733 ), .A2(_AES_ENC_us20_n732 ), .A3(_AES_ENC_us20_n731 ), .A4(_AES_ENC_us20_n730 ), .ZN(_AES_ENC_sa20_sub[1] ) );
NAND2_X2 _AES_ENC_us20_U341  ( .A1(_AES_ENC_sa20[7]), .A2(_AES_ENC_us20_n593 ), .ZN(_AES_ENC_us20_n734 ) );
NAND2_X2 _AES_ENC_us20_U340  ( .A1(_AES_ENC_us20_n734 ), .A2(_AES_ENC_us20_n588 ), .ZN(_AES_ENC_us20_n738 ) );
OR4_X2 _AES_ENC_us20_U339  ( .A1(_AES_ENC_us20_n738 ), .A2(_AES_ENC_us20_n596 ), .A3(_AES_ENC_us20_n826 ), .A4(_AES_ENC_us20_n1121 ), .ZN(_AES_ENC_us20_n746 ) );
NAND2_X2 _AES_ENC_us20_U337  ( .A1(_AES_ENC_us20_n1100 ), .A2(_AES_ENC_us20_n617 ), .ZN(_AES_ENC_us20_n992 ) );
OR2_X2 _AES_ENC_us20_U336  ( .A1(_AES_ENC_us20_n592 ), .A2(_AES_ENC_us20_n735 ), .ZN(_AES_ENC_us20_n737 ) );
NAND2_X2 _AES_ENC_us20_U334  ( .A1(_AES_ENC_us20_n605 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n753 ) );
NAND2_X2 _AES_ENC_us20_U333  ( .A1(_AES_ENC_us20_n603 ), .A2(_AES_ENC_us20_n753 ), .ZN(_AES_ENC_us20_n1080 ) );
NAND2_X2 _AES_ENC_us20_U332  ( .A1(_AES_ENC_us20_n1048 ), .A2(_AES_ENC_us20_n602 ), .ZN(_AES_ENC_us20_n736 ) );
NAND2_X2 _AES_ENC_us20_U331  ( .A1(_AES_ENC_us20_n737 ), .A2(_AES_ENC_us20_n736 ), .ZN(_AES_ENC_us20_n739 ) );
NAND2_X2 _AES_ENC_us20_U330  ( .A1(_AES_ENC_us20_n739 ), .A2(_AES_ENC_us20_n738 ), .ZN(_AES_ENC_us20_n745 ) );
NAND2_X2 _AES_ENC_us20_U326  ( .A1(_AES_ENC_us20_n1096 ), .A2(_AES_ENC_us20_n598 ), .ZN(_AES_ENC_us20_n906 ) );
NAND4_X2 _AES_ENC_us20_U323  ( .A1(_AES_ENC_us20_n746 ), .A2(_AES_ENC_us20_n992 ), .A3(_AES_ENC_us20_n745 ), .A4(_AES_ENC_us20_n744 ), .ZN(_AES_ENC_us20_n747 ) );
NAND2_X2 _AES_ENC_us20_U322  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n747 ), .ZN(_AES_ENC_us20_n793 ) );
NAND2_X2 _AES_ENC_us20_U321  ( .A1(_AES_ENC_us20_n606 ), .A2(_AES_ENC_us20_n855 ), .ZN(_AES_ENC_us20_n748 ) );
NAND2_X2 _AES_ENC_us20_U320  ( .A1(_AES_ENC_us20_n956 ), .A2(_AES_ENC_us20_n748 ), .ZN(_AES_ENC_us20_n760 ) );
NAND2_X2 _AES_ENC_us20_U313  ( .A1(_AES_ENC_us20_n598 ), .A2(_AES_ENC_us20_n753 ), .ZN(_AES_ENC_us20_n1023 ) );
NAND4_X2 _AES_ENC_us20_U308  ( .A1(_AES_ENC_us20_n760 ), .A2(_AES_ENC_us20_n992 ), .A3(_AES_ENC_us20_n759 ), .A4(_AES_ENC_us20_n758 ), .ZN(_AES_ENC_us20_n761 ) );
NAND2_X2 _AES_ENC_us20_U307  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n761 ), .ZN(_AES_ENC_us20_n792 ) );
NAND2_X2 _AES_ENC_us20_U306  ( .A1(_AES_ENC_us20_n606 ), .A2(_AES_ENC_us20_n610 ), .ZN(_AES_ENC_us20_n989 ) );
NAND2_X2 _AES_ENC_us20_U305  ( .A1(_AES_ENC_us20_n1050 ), .A2(_AES_ENC_us20_n989 ), .ZN(_AES_ENC_us20_n777 ) );
NAND2_X2 _AES_ENC_us20_U304  ( .A1(_AES_ENC_us20_n1093 ), .A2(_AES_ENC_us20_n762 ), .ZN(_AES_ENC_us20_n776 ) );
XNOR2_X2 _AES_ENC_us20_U301  ( .A(_AES_ENC_sa20[7]), .B(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n959 ) );
NAND4_X2 _AES_ENC_us20_U289  ( .A1(_AES_ENC_us20_n777 ), .A2(_AES_ENC_us20_n776 ), .A3(_AES_ENC_us20_n775 ), .A4(_AES_ENC_us20_n774 ), .ZN(_AES_ENC_us20_n778 ) );
NAND2_X2 _AES_ENC_us20_U288  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n778 ), .ZN(_AES_ENC_us20_n791 ) );
NAND2_X2 _AES_ENC_us20_U287  ( .A1(_AES_ENC_us20_n1056 ), .A2(_AES_ENC_us20_n1050 ), .ZN(_AES_ENC_us20_n788 ) );
NAND2_X2 _AES_ENC_us20_U286  ( .A1(_AES_ENC_us20_n1091 ), .A2(_AES_ENC_us20_n779 ), .ZN(_AES_ENC_us20_n787 ) );
NAND2_X2 _AES_ENC_us20_U285  ( .A1(_AES_ENC_us20_n956 ), .A2(_AES_ENC_sa20[1]), .ZN(_AES_ENC_us20_n786 ) );
NAND4_X2 _AES_ENC_us20_U278  ( .A1(_AES_ENC_us20_n788 ), .A2(_AES_ENC_us20_n787 ), .A3(_AES_ENC_us20_n786 ), .A4(_AES_ENC_us20_n785 ), .ZN(_AES_ENC_us20_n789 ) );
NAND2_X2 _AES_ENC_us20_U277  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n789 ), .ZN(_AES_ENC_us20_n790 ) );
NAND4_X2 _AES_ENC_us20_U276  ( .A1(_AES_ENC_us20_n793 ), .A2(_AES_ENC_us20_n792 ), .A3(_AES_ENC_us20_n791 ), .A4(_AES_ENC_us20_n790 ), .ZN(_AES_ENC_sa20_sub[2] ) );
NAND2_X2 _AES_ENC_us20_U275  ( .A1(_AES_ENC_us20_n1059 ), .A2(_AES_ENC_us20_n794 ), .ZN(_AES_ENC_us20_n810 ) );
NAND2_X2 _AES_ENC_us20_U274  ( .A1(_AES_ENC_us20_n1049 ), .A2(_AES_ENC_us20_n956 ), .ZN(_AES_ENC_us20_n809 ) );
OR2_X2 _AES_ENC_us20_U266  ( .A1(_AES_ENC_us20_n1096 ), .A2(_AES_ENC_us20_n587 ), .ZN(_AES_ENC_us20_n802 ) );
NAND2_X2 _AES_ENC_us20_U265  ( .A1(_AES_ENC_us20_n1053 ), .A2(_AES_ENC_us20_n800 ), .ZN(_AES_ENC_us20_n801 ) );
NAND2_X2 _AES_ENC_us20_U264  ( .A1(_AES_ENC_us20_n802 ), .A2(_AES_ENC_us20_n801 ), .ZN(_AES_ENC_us20_n805 ) );
NAND4_X2 _AES_ENC_us20_U261  ( .A1(_AES_ENC_us20_n810 ), .A2(_AES_ENC_us20_n809 ), .A3(_AES_ENC_us20_n808 ), .A4(_AES_ENC_us20_n807 ), .ZN(_AES_ENC_us20_n811 ) );
NAND2_X2 _AES_ENC_us20_U260  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n811 ), .ZN(_AES_ENC_us20_n852 ) );
OR2_X2 _AES_ENC_us20_U259  ( .A1(_AES_ENC_us20_n1023 ), .A2(_AES_ENC_us20_n575 ), .ZN(_AES_ENC_us20_n819 ) );
OR2_X2 _AES_ENC_us20_U257  ( .A1(_AES_ENC_us20_n570 ), .A2(_AES_ENC_us20_n930 ), .ZN(_AES_ENC_us20_n818 ) );
NAND2_X2 _AES_ENC_us20_U256  ( .A1(_AES_ENC_us20_n1013 ), .A2(_AES_ENC_us20_n1094 ), .ZN(_AES_ENC_us20_n817 ) );
NAND4_X2 _AES_ENC_us20_U249  ( .A1(_AES_ENC_us20_n819 ), .A2(_AES_ENC_us20_n818 ), .A3(_AES_ENC_us20_n817 ), .A4(_AES_ENC_us20_n816 ), .ZN(_AES_ENC_us20_n820 ) );
NAND2_X2 _AES_ENC_us20_U248  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n820 ), .ZN(_AES_ENC_us20_n851 ) );
NAND2_X2 _AES_ENC_us20_U247  ( .A1(_AES_ENC_us20_n956 ), .A2(_AES_ENC_us20_n1080 ), .ZN(_AES_ENC_us20_n835 ) );
NAND2_X2 _AES_ENC_us20_U246  ( .A1(_AES_ENC_us20_n570 ), .A2(_AES_ENC_us20_n1030 ), .ZN(_AES_ENC_us20_n1047 ) );
OR2_X2 _AES_ENC_us20_U245  ( .A1(_AES_ENC_us20_n1047 ), .A2(_AES_ENC_us20_n582 ), .ZN(_AES_ENC_us20_n834 ) );
NAND2_X2 _AES_ENC_us20_U244  ( .A1(_AES_ENC_us20_n1072 ), .A2(_AES_ENC_us20_n620 ), .ZN(_AES_ENC_us20_n833 ) );
NAND4_X2 _AES_ENC_us20_U233  ( .A1(_AES_ENC_us20_n835 ), .A2(_AES_ENC_us20_n834 ), .A3(_AES_ENC_us20_n833 ), .A4(_AES_ENC_us20_n832 ), .ZN(_AES_ENC_us20_n836 ) );
NAND2_X2 _AES_ENC_us20_U232  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n836 ), .ZN(_AES_ENC_us20_n850 ) );
NAND2_X2 _AES_ENC_us20_U231  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n601 ), .ZN(_AES_ENC_us20_n847 ) );
NAND2_X2 _AES_ENC_us20_U230  ( .A1(_AES_ENC_us20_n1050 ), .A2(_AES_ENC_us20_n1071 ), .ZN(_AES_ENC_us20_n846 ) );
OR2_X2 _AES_ENC_us20_U224  ( .A1(_AES_ENC_us20_n1053 ), .A2(_AES_ENC_us20_n911 ), .ZN(_AES_ENC_us20_n1077 ) );
NAND4_X2 _AES_ENC_us20_U220  ( .A1(_AES_ENC_us20_n847 ), .A2(_AES_ENC_us20_n846 ), .A3(_AES_ENC_us20_n845 ), .A4(_AES_ENC_us20_n844 ), .ZN(_AES_ENC_us20_n848 ) );
NAND2_X2 _AES_ENC_us20_U219  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n848 ), .ZN(_AES_ENC_us20_n849 ) );
NAND4_X2 _AES_ENC_us20_U218  ( .A1(_AES_ENC_us20_n852 ), .A2(_AES_ENC_us20_n851 ), .A3(_AES_ENC_us20_n850 ), .A4(_AES_ENC_us20_n849 ), .ZN(_AES_ENC_sa20_sub[3] ) );
NAND2_X2 _AES_ENC_us20_U216  ( .A1(_AES_ENC_us20_n1009 ), .A2(_AES_ENC_us20_n1072 ), .ZN(_AES_ENC_us20_n862 ) );
NAND2_X2 _AES_ENC_us20_U215  ( .A1(_AES_ENC_us20_n610 ), .A2(_AES_ENC_us20_n618 ), .ZN(_AES_ENC_us20_n853 ) );
NAND2_X2 _AES_ENC_us20_U214  ( .A1(_AES_ENC_us20_n1050 ), .A2(_AES_ENC_us20_n853 ), .ZN(_AES_ENC_us20_n861 ) );
NAND4_X2 _AES_ENC_us20_U206  ( .A1(_AES_ENC_us20_n862 ), .A2(_AES_ENC_us20_n861 ), .A3(_AES_ENC_us20_n860 ), .A4(_AES_ENC_us20_n859 ), .ZN(_AES_ENC_us20_n863 ) );
NAND2_X2 _AES_ENC_us20_U205  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n863 ), .ZN(_AES_ENC_us20_n905 ) );
NAND2_X2 _AES_ENC_us20_U204  ( .A1(_AES_ENC_us20_n1010 ), .A2(_AES_ENC_us20_n989 ), .ZN(_AES_ENC_us20_n874 ) );
NAND2_X2 _AES_ENC_us20_U203  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n592 ), .ZN(_AES_ENC_us20_n864 ) );
NAND2_X2 _AES_ENC_us20_U202  ( .A1(_AES_ENC_us20_n929 ), .A2(_AES_ENC_us20_n864 ), .ZN(_AES_ENC_us20_n873 ) );
NAND4_X2 _AES_ENC_us20_U193  ( .A1(_AES_ENC_us20_n874 ), .A2(_AES_ENC_us20_n873 ), .A3(_AES_ENC_us20_n872 ), .A4(_AES_ENC_us20_n871 ), .ZN(_AES_ENC_us20_n875 ) );
NAND2_X2 _AES_ENC_us20_U192  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n875 ), .ZN(_AES_ENC_us20_n904 ) );
NAND2_X2 _AES_ENC_us20_U191  ( .A1(_AES_ENC_us20_n597 ), .A2(_AES_ENC_us20_n1050 ), .ZN(_AES_ENC_us20_n889 ) );
NAND2_X2 _AES_ENC_us20_U190  ( .A1(_AES_ENC_us20_n1093 ), .A2(_AES_ENC_us20_n617 ), .ZN(_AES_ENC_us20_n876 ) );
NAND2_X2 _AES_ENC_us20_U189  ( .A1(_AES_ENC_us20_n576 ), .A2(_AES_ENC_us20_n876 ), .ZN(_AES_ENC_us20_n877 ) );
NAND2_X2 _AES_ENC_us20_U188  ( .A1(_AES_ENC_us20_n877 ), .A2(_AES_ENC_us20_n601 ), .ZN(_AES_ENC_us20_n888 ) );
NAND4_X2 _AES_ENC_us20_U179  ( .A1(_AES_ENC_us20_n889 ), .A2(_AES_ENC_us20_n888 ), .A3(_AES_ENC_us20_n887 ), .A4(_AES_ENC_us20_n886 ), .ZN(_AES_ENC_us20_n890 ) );
NAND2_X2 _AES_ENC_us20_U178  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n890 ), .ZN(_AES_ENC_us20_n903 ) );
OR2_X2 _AES_ENC_us20_U177  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n1059 ), .ZN(_AES_ENC_us20_n900 ) );
NAND2_X2 _AES_ENC_us20_U176  ( .A1(_AES_ENC_us20_n1073 ), .A2(_AES_ENC_us20_n1047 ), .ZN(_AES_ENC_us20_n899 ) );
NAND2_X2 _AES_ENC_us20_U175  ( .A1(_AES_ENC_us20_n1094 ), .A2(_AES_ENC_us20_n608 ), .ZN(_AES_ENC_us20_n898 ) );
NAND4_X2 _AES_ENC_us20_U167  ( .A1(_AES_ENC_us20_n900 ), .A2(_AES_ENC_us20_n899 ), .A3(_AES_ENC_us20_n898 ), .A4(_AES_ENC_us20_n897 ), .ZN(_AES_ENC_us20_n901 ) );
NAND2_X2 _AES_ENC_us20_U166  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n901 ), .ZN(_AES_ENC_us20_n902 ) );
NAND4_X2 _AES_ENC_us20_U165  ( .A1(_AES_ENC_us20_n905 ), .A2(_AES_ENC_us20_n904 ), .A3(_AES_ENC_us20_n903 ), .A4(_AES_ENC_us20_n902 ), .ZN(_AES_ENC_sa20_sub[4] ) );
NAND2_X2 _AES_ENC_us20_U164  ( .A1(_AES_ENC_us20_n1094 ), .A2(_AES_ENC_us20_n615 ), .ZN(_AES_ENC_us20_n922 ) );
NAND2_X2 _AES_ENC_us20_U163  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n989 ), .ZN(_AES_ENC_us20_n921 ) );
NAND4_X2 _AES_ENC_us20_U151  ( .A1(_AES_ENC_us20_n922 ), .A2(_AES_ENC_us20_n921 ), .A3(_AES_ENC_us20_n920 ), .A4(_AES_ENC_us20_n919 ), .ZN(_AES_ENC_us20_n923 ) );
NAND2_X2 _AES_ENC_us20_U150  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n923 ), .ZN(_AES_ENC_us20_n972 ) );
NAND2_X2 _AES_ENC_us20_U149  ( .A1(_AES_ENC_us20_n603 ), .A2(_AES_ENC_us20_n605 ), .ZN(_AES_ENC_us20_n924 ) );
NAND2_X2 _AES_ENC_us20_U148  ( .A1(_AES_ENC_us20_n1073 ), .A2(_AES_ENC_us20_n924 ), .ZN(_AES_ENC_us20_n939 ) );
NAND2_X2 _AES_ENC_us20_U147  ( .A1(_AES_ENC_us20_n926 ), .A2(_AES_ENC_us20_n925 ), .ZN(_AES_ENC_us20_n927 ) );
NAND2_X2 _AES_ENC_us20_U146  ( .A1(_AES_ENC_us20_n587 ), .A2(_AES_ENC_us20_n927 ), .ZN(_AES_ENC_us20_n928 ) );
NAND2_X2 _AES_ENC_us20_U145  ( .A1(_AES_ENC_us20_n928 ), .A2(_AES_ENC_us20_n1080 ), .ZN(_AES_ENC_us20_n938 ) );
OR2_X2 _AES_ENC_us20_U144  ( .A1(_AES_ENC_us20_n1117 ), .A2(_AES_ENC_us20_n580 ), .ZN(_AES_ENC_us20_n937 ) );
NAND4_X2 _AES_ENC_us20_U139  ( .A1(_AES_ENC_us20_n939 ), .A2(_AES_ENC_us20_n938 ), .A3(_AES_ENC_us20_n937 ), .A4(_AES_ENC_us20_n936 ), .ZN(_AES_ENC_us20_n940 ) );
NAND2_X2 _AES_ENC_us20_U138  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n940 ), .ZN(_AES_ENC_us20_n971 ) );
OR2_X2 _AES_ENC_us20_U137  ( .A1(_AES_ENC_us20_n586 ), .A2(_AES_ENC_us20_n941 ), .ZN(_AES_ENC_us20_n954 ) );
NAND2_X2 _AES_ENC_us20_U136  ( .A1(_AES_ENC_us20_n1096 ), .A2(_AES_ENC_us20_n618 ), .ZN(_AES_ENC_us20_n942 ) );
NAND2_X2 _AES_ENC_us20_U135  ( .A1(_AES_ENC_us20_n1048 ), .A2(_AES_ENC_us20_n942 ), .ZN(_AES_ENC_us20_n943 ) );
NAND2_X2 _AES_ENC_us20_U134  ( .A1(_AES_ENC_us20_n582 ), .A2(_AES_ENC_us20_n943 ), .ZN(_AES_ENC_us20_n944 ) );
NAND2_X2 _AES_ENC_us20_U133  ( .A1(_AES_ENC_us20_n944 ), .A2(_AES_ENC_us20_n599 ), .ZN(_AES_ENC_us20_n953 ) );
NAND4_X2 _AES_ENC_us20_U125  ( .A1(_AES_ENC_us20_n954 ), .A2(_AES_ENC_us20_n953 ), .A3(_AES_ENC_us20_n952 ), .A4(_AES_ENC_us20_n951 ), .ZN(_AES_ENC_us20_n955 ) );
NAND2_X2 _AES_ENC_us20_U124  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n955 ), .ZN(_AES_ENC_us20_n970 ) );
NAND2_X2 _AES_ENC_us20_U123  ( .A1(_AES_ENC_us20_n1094 ), .A2(_AES_ENC_us20_n1071 ), .ZN(_AES_ENC_us20_n967 ) );
NAND2_X2 _AES_ENC_us20_U122  ( .A1(_AES_ENC_us20_n956 ), .A2(_AES_ENC_us20_n1030 ), .ZN(_AES_ENC_us20_n966 ) );
NAND4_X2 _AES_ENC_us20_U114  ( .A1(_AES_ENC_us20_n967 ), .A2(_AES_ENC_us20_n966 ), .A3(_AES_ENC_us20_n965 ), .A4(_AES_ENC_us20_n964 ), .ZN(_AES_ENC_us20_n968 ) );
NAND2_X2 _AES_ENC_us20_U113  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n968 ), .ZN(_AES_ENC_us20_n969 ) );
NAND4_X2 _AES_ENC_us20_U112  ( .A1(_AES_ENC_us20_n972 ), .A2(_AES_ENC_us20_n971 ), .A3(_AES_ENC_us20_n970 ), .A4(_AES_ENC_us20_n969 ), .ZN(_AES_ENC_sa20_sub[5] ) );
NAND2_X2 _AES_ENC_us20_U111  ( .A1(_AES_ENC_us20_n570 ), .A2(_AES_ENC_us20_n1097 ), .ZN(_AES_ENC_us20_n973 ) );
NAND2_X2 _AES_ENC_us20_U110  ( .A1(_AES_ENC_us20_n1073 ), .A2(_AES_ENC_us20_n973 ), .ZN(_AES_ENC_us20_n987 ) );
NAND2_X2 _AES_ENC_us20_U109  ( .A1(_AES_ENC_us20_n974 ), .A2(_AES_ENC_us20_n1077 ), .ZN(_AES_ENC_us20_n975 ) );
NAND2_X2 _AES_ENC_us20_U108  ( .A1(_AES_ENC_us20_n584 ), .A2(_AES_ENC_us20_n975 ), .ZN(_AES_ENC_us20_n976 ) );
NAND2_X2 _AES_ENC_us20_U107  ( .A1(_AES_ENC_us20_n977 ), .A2(_AES_ENC_us20_n976 ), .ZN(_AES_ENC_us20_n986 ) );
NAND4_X2 _AES_ENC_us20_U99  ( .A1(_AES_ENC_us20_n987 ), .A2(_AES_ENC_us20_n986 ), .A3(_AES_ENC_us20_n985 ), .A4(_AES_ENC_us20_n984 ), .ZN(_AES_ENC_us20_n988 ) );
NAND2_X2 _AES_ENC_us20_U98  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n988 ), .ZN(_AES_ENC_us20_n1044 ) );
NAND2_X2 _AES_ENC_us20_U97  ( .A1(_AES_ENC_us20_n1073 ), .A2(_AES_ENC_us20_n989 ), .ZN(_AES_ENC_us20_n1004 ) );
NAND2_X2 _AES_ENC_us20_U96  ( .A1(_AES_ENC_us20_n1092 ), .A2(_AES_ENC_us20_n605 ), .ZN(_AES_ENC_us20_n1003 ) );
NAND4_X2 _AES_ENC_us20_U85  ( .A1(_AES_ENC_us20_n1004 ), .A2(_AES_ENC_us20_n1003 ), .A3(_AES_ENC_us20_n1002 ), .A4(_AES_ENC_us20_n1001 ), .ZN(_AES_ENC_us20_n1005 ) );
NAND2_X2 _AES_ENC_us20_U84  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n1005 ), .ZN(_AES_ENC_us20_n1043 ) );
NAND2_X2 _AES_ENC_us20_U83  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n626 ), .ZN(_AES_ENC_us20_n1020 ) );
NAND2_X2 _AES_ENC_us20_U82  ( .A1(_AES_ENC_us20_n1050 ), .A2(_AES_ENC_us20_n612 ), .ZN(_AES_ENC_us20_n1019 ) );
NAND2_X2 _AES_ENC_us20_U77  ( .A1(_AES_ENC_us20_n1059 ), .A2(_AES_ENC_us20_n1114 ), .ZN(_AES_ENC_us20_n1012 ) );
NAND2_X2 _AES_ENC_us20_U76  ( .A1(_AES_ENC_us20_n1010 ), .A2(_AES_ENC_us20_n604 ), .ZN(_AES_ENC_us20_n1011 ) );
NAND2_X2 _AES_ENC_us20_U75  ( .A1(_AES_ENC_us20_n1012 ), .A2(_AES_ENC_us20_n1011 ), .ZN(_AES_ENC_us20_n1016 ) );
NAND4_X2 _AES_ENC_us20_U70  ( .A1(_AES_ENC_us20_n1020 ), .A2(_AES_ENC_us20_n1019 ), .A3(_AES_ENC_us20_n1018 ), .A4(_AES_ENC_us20_n1017 ), .ZN(_AES_ENC_us20_n1021 ) );
NAND2_X2 _AES_ENC_us20_U69  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n1021 ), .ZN(_AES_ENC_us20_n1042 ) );
NAND2_X2 _AES_ENC_us20_U68  ( .A1(_AES_ENC_us20_n1022 ), .A2(_AES_ENC_us20_n1093 ), .ZN(_AES_ENC_us20_n1039 ) );
NAND2_X2 _AES_ENC_us20_U67  ( .A1(_AES_ENC_us20_n1050 ), .A2(_AES_ENC_us20_n1023 ), .ZN(_AES_ENC_us20_n1038 ) );
NAND2_X2 _AES_ENC_us20_U66  ( .A1(_AES_ENC_us20_n1024 ), .A2(_AES_ENC_us20_n1071 ), .ZN(_AES_ENC_us20_n1037 ) );
AND2_X2 _AES_ENC_us20_U60  ( .A1(_AES_ENC_us20_n1030 ), .A2(_AES_ENC_us20_n621 ), .ZN(_AES_ENC_us20_n1078 ) );
NAND4_X2 _AES_ENC_us20_U56  ( .A1(_AES_ENC_us20_n1039 ), .A2(_AES_ENC_us20_n1038 ), .A3(_AES_ENC_us20_n1037 ), .A4(_AES_ENC_us20_n1036 ), .ZN(_AES_ENC_us20_n1040 ) );
NAND2_X2 _AES_ENC_us20_U55  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n1040 ), .ZN(_AES_ENC_us20_n1041 ) );
NAND4_X2 _AES_ENC_us20_U54  ( .A1(_AES_ENC_us20_n1044 ), .A2(_AES_ENC_us20_n1043 ), .A3(_AES_ENC_us20_n1042 ), .A4(_AES_ENC_us20_n1041 ), .ZN(_AES_ENC_sa20_sub[6] ) );
NAND2_X2 _AES_ENC_us20_U53  ( .A1(_AES_ENC_us20_n1072 ), .A2(_AES_ENC_us20_n1045 ), .ZN(_AES_ENC_us20_n1068 ) );
NAND2_X2 _AES_ENC_us20_U52  ( .A1(_AES_ENC_us20_n1046 ), .A2(_AES_ENC_us20_n603 ), .ZN(_AES_ENC_us20_n1067 ) );
NAND2_X2 _AES_ENC_us20_U51  ( .A1(_AES_ENC_us20_n1094 ), .A2(_AES_ENC_us20_n1047 ), .ZN(_AES_ENC_us20_n1066 ) );
NAND4_X2 _AES_ENC_us20_U40  ( .A1(_AES_ENC_us20_n1068 ), .A2(_AES_ENC_us20_n1067 ), .A3(_AES_ENC_us20_n1066 ), .A4(_AES_ENC_us20_n1065 ), .ZN(_AES_ENC_us20_n1069 ) );
NAND2_X2 _AES_ENC_us20_U39  ( .A1(_AES_ENC_us20_n1070 ), .A2(_AES_ENC_us20_n1069 ), .ZN(_AES_ENC_us20_n1135 ) );
NAND2_X2 _AES_ENC_us20_U38  ( .A1(_AES_ENC_us20_n1072 ), .A2(_AES_ENC_us20_n1071 ), .ZN(_AES_ENC_us20_n1088 ) );
NAND2_X2 _AES_ENC_us20_U37  ( .A1(_AES_ENC_us20_n1073 ), .A2(_AES_ENC_us20_n608 ), .ZN(_AES_ENC_us20_n1087 ) );
NAND4_X2 _AES_ENC_us20_U28  ( .A1(_AES_ENC_us20_n1088 ), .A2(_AES_ENC_us20_n1087 ), .A3(_AES_ENC_us20_n1086 ), .A4(_AES_ENC_us20_n1085 ), .ZN(_AES_ENC_us20_n1089 ) );
NAND2_X2 _AES_ENC_us20_U27  ( .A1(_AES_ENC_us20_n1090 ), .A2(_AES_ENC_us20_n1089 ), .ZN(_AES_ENC_us20_n1134 ) );
NAND2_X2 _AES_ENC_us20_U26  ( .A1(_AES_ENC_us20_n1091 ), .A2(_AES_ENC_us20_n1093 ), .ZN(_AES_ENC_us20_n1111 ) );
NAND2_X2 _AES_ENC_us20_U25  ( .A1(_AES_ENC_us20_n1092 ), .A2(_AES_ENC_us20_n1120 ), .ZN(_AES_ENC_us20_n1110 ) );
AND2_X2 _AES_ENC_us20_U22  ( .A1(_AES_ENC_us20_n1097 ), .A2(_AES_ENC_us20_n1096 ), .ZN(_AES_ENC_us20_n1098 ) );
NAND4_X2 _AES_ENC_us20_U14  ( .A1(_AES_ENC_us20_n1111 ), .A2(_AES_ENC_us20_n1110 ), .A3(_AES_ENC_us20_n1109 ), .A4(_AES_ENC_us20_n1108 ), .ZN(_AES_ENC_us20_n1112 ) );
NAND2_X2 _AES_ENC_us20_U13  ( .A1(_AES_ENC_us20_n1113 ), .A2(_AES_ENC_us20_n1112 ), .ZN(_AES_ENC_us20_n1133 ) );
NAND2_X2 _AES_ENC_us20_U12  ( .A1(_AES_ENC_us20_n1115 ), .A2(_AES_ENC_us20_n1114 ), .ZN(_AES_ENC_us20_n1129 ) );
OR2_X2 _AES_ENC_us20_U11  ( .A1(_AES_ENC_us20_n579 ), .A2(_AES_ENC_us20_n1116 ), .ZN(_AES_ENC_us20_n1128 ) );
NAND4_X2 _AES_ENC_us20_U3  ( .A1(_AES_ENC_us20_n1129 ), .A2(_AES_ENC_us20_n1128 ), .A3(_AES_ENC_us20_n1127 ), .A4(_AES_ENC_us20_n1126 ), .ZN(_AES_ENC_us20_n1130 ) );
NAND2_X2 _AES_ENC_us20_U2  ( .A1(_AES_ENC_us20_n1131 ), .A2(_AES_ENC_us20_n1130 ), .ZN(_AES_ENC_us20_n1132 ) );
NAND4_X2 _AES_ENC_us20_U1  ( .A1(_AES_ENC_us20_n1135 ), .A2(_AES_ENC_us20_n1134 ), .A3(_AES_ENC_us20_n1133 ), .A4(_AES_ENC_us20_n1132 ), .ZN(_AES_ENC_sa20_sub[7] ) );
INV_X4 _AES_ENC_us21_U575  ( .A(_AES_ENC_sa21[0]), .ZN(_AES_ENC_us21_n627 ));
INV_X4 _AES_ENC_us21_U574  ( .A(_AES_ENC_us21_n1053 ), .ZN(_AES_ENC_us21_n625 ) );
INV_X4 _AES_ENC_us21_U573  ( .A(_AES_ENC_us21_n1103 ), .ZN(_AES_ENC_us21_n623 ) );
INV_X4 _AES_ENC_us21_U572  ( .A(_AES_ENC_us21_n1056 ), .ZN(_AES_ENC_us21_n622 ) );
INV_X4 _AES_ENC_us21_U571  ( .A(_AES_ENC_us21_n1102 ), .ZN(_AES_ENC_us21_n621 ) );
INV_X4 _AES_ENC_us21_U570  ( .A(_AES_ENC_us21_n1074 ), .ZN(_AES_ENC_us21_n620 ) );
INV_X4 _AES_ENC_us21_U569  ( .A(_AES_ENC_us21_n929 ), .ZN(_AES_ENC_us21_n619 ) );
INV_X4 _AES_ENC_us21_U568  ( .A(_AES_ENC_us21_n1091 ), .ZN(_AES_ENC_us21_n618 ) );
INV_X4 _AES_ENC_us21_U567  ( .A(_AES_ENC_us21_n826 ), .ZN(_AES_ENC_us21_n617 ) );
INV_X4 _AES_ENC_us21_U566  ( .A(_AES_ENC_us21_n1031 ), .ZN(_AES_ENC_us21_n616 ) );
INV_X4 _AES_ENC_us21_U565  ( .A(_AES_ENC_us21_n1054 ), .ZN(_AES_ENC_us21_n615 ) );
INV_X4 _AES_ENC_us21_U564  ( .A(_AES_ENC_us21_n1025 ), .ZN(_AES_ENC_us21_n614 ) );
INV_X4 _AES_ENC_us21_U563  ( .A(_AES_ENC_us21_n990 ), .ZN(_AES_ENC_us21_n613 ) );
INV_X4 _AES_ENC_us21_U562  ( .A(_AES_ENC_sa21[4]), .ZN(_AES_ENC_us21_n612 ));
INV_X4 _AES_ENC_us21_U561  ( .A(_AES_ENC_us21_n881 ), .ZN(_AES_ENC_us21_n611 ) );
INV_X4 _AES_ENC_us21_U560  ( .A(_AES_ENC_us21_n1022 ), .ZN(_AES_ENC_us21_n610 ) );
INV_X4 _AES_ENC_us21_U559  ( .A(_AES_ENC_us21_n1120 ), .ZN(_AES_ENC_us21_n609 ) );
INV_X4 _AES_ENC_us21_U558  ( .A(_AES_ENC_us21_n977 ), .ZN(_AES_ENC_us21_n608 ) );
INV_X4 _AES_ENC_us21_U557  ( .A(_AES_ENC_us21_n926 ), .ZN(_AES_ENC_us21_n607 ) );
INV_X4 _AES_ENC_us21_U556  ( .A(_AES_ENC_us21_n910 ), .ZN(_AES_ENC_us21_n606 ) );
INV_X4 _AES_ENC_us21_U555  ( .A(_AES_ENC_us21_n1121 ), .ZN(_AES_ENC_us21_n605 ) );
INV_X4 _AES_ENC_us21_U554  ( .A(_AES_ENC_us21_n1009 ), .ZN(_AES_ENC_us21_n604 ) );
INV_X4 _AES_ENC_us21_U553  ( .A(_AES_ENC_us21_n1080 ), .ZN(_AES_ENC_us21_n602 ) );
INV_X4 _AES_ENC_us21_U552  ( .A(_AES_ENC_us21_n821 ), .ZN(_AES_ENC_us21_n600 ) );
INV_X4 _AES_ENC_us21_U551  ( .A(_AES_ENC_us21_n1013 ), .ZN(_AES_ENC_us21_n599 ) );
INV_X4 _AES_ENC_us21_U550  ( .A(_AES_ENC_us21_n1058 ), .ZN(_AES_ENC_us21_n598 ) );
INV_X4 _AES_ENC_us21_U549  ( .A(_AES_ENC_us21_n906 ), .ZN(_AES_ENC_us21_n597 ) );
INV_X4 _AES_ENC_us21_U548  ( .A(_AES_ENC_us21_n959 ), .ZN(_AES_ENC_us21_n596 ) );
INV_X4 _AES_ENC_us21_U547  ( .A(_AES_ENC_sa21[7]), .ZN(_AES_ENC_us21_n595 ));
INV_X4 _AES_ENC_us21_U546  ( .A(_AES_ENC_us21_n1114 ), .ZN(_AES_ENC_us21_n593 ) );
INV_X4 _AES_ENC_us21_U545  ( .A(_AES_ENC_us21_n1048 ), .ZN(_AES_ENC_us21_n592 ) );
INV_X4 _AES_ENC_us21_U544  ( .A(_AES_ENC_us21_n974 ), .ZN(_AES_ENC_us21_n590 ) );
INV_X4 _AES_ENC_us21_U543  ( .A(_AES_ENC_us21_n794 ), .ZN(_AES_ENC_us21_n588 ) );
INV_X4 _AES_ENC_us21_U542  ( .A(_AES_ENC_us21_n880 ), .ZN(_AES_ENC_us21_n586 ) );
INV_X4 _AES_ENC_us21_U541  ( .A(_AES_ENC_sa21[2]), .ZN(_AES_ENC_us21_n584 ));
INV_X4 _AES_ENC_us21_U540  ( .A(_AES_ENC_us21_n800 ), .ZN(_AES_ENC_us21_n583 ) );
INV_X4 _AES_ENC_us21_U539  ( .A(_AES_ENC_us21_n925 ), .ZN(_AES_ENC_us21_n582 ) );
INV_X4 _AES_ENC_us21_U538  ( .A(_AES_ENC_us21_n992 ), .ZN(_AES_ENC_us21_n580 ) );
INV_X4 _AES_ENC_us21_U537  ( .A(_AES_ENC_us21_n779 ), .ZN(_AES_ENC_us21_n579 ) );
INV_X4 _AES_ENC_us21_U536  ( .A(_AES_ENC_us21_n1092 ), .ZN(_AES_ENC_us21_n575 ) );
INV_X4 _AES_ENC_us21_U535  ( .A(_AES_ENC_us21_n824 ), .ZN(_AES_ENC_us21_n574 ) );
NOR2_X2 _AES_ENC_us21_U534  ( .A1(_AES_ENC_sa21[0]), .A2(_AES_ENC_sa21[6]),.ZN(_AES_ENC_us21_n1090 ) );
NOR2_X2 _AES_ENC_us21_U533  ( .A1(_AES_ENC_us21_n627 ), .A2(_AES_ENC_sa21[6]), .ZN(_AES_ENC_us21_n1070 ) );
NOR2_X2 _AES_ENC_us21_U532  ( .A1(_AES_ENC_sa21[4]), .A2(_AES_ENC_sa21[3]),.ZN(_AES_ENC_us21_n1025 ) );
INV_X4 _AES_ENC_us21_U531  ( .A(_AES_ENC_us21_n569 ), .ZN(_AES_ENC_us21_n572 ) );
NOR2_X2 _AES_ENC_us21_U530  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n765 ) );
NOR2_X2 _AES_ENC_us21_U529  ( .A1(_AES_ENC_sa21[4]), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n764 ) );
NOR2_X2 _AES_ENC_us21_U528  ( .A1(_AES_ENC_us21_n765 ), .A2(_AES_ENC_us21_n764 ), .ZN(_AES_ENC_us21_n766 ) );
NOR2_X2 _AES_ENC_us21_U527  ( .A1(_AES_ENC_us21_n766 ), .A2(_AES_ENC_us21_n596 ), .ZN(_AES_ENC_us21_n767 ) );
NOR3_X2 _AES_ENC_us21_U526  ( .A1(_AES_ENC_us21_n595 ), .A2(_AES_ENC_sa21[5]), .A3(_AES_ENC_us21_n704 ), .ZN(_AES_ENC_us21_n706 ));
NOR2_X2 _AES_ENC_us21_U525  ( .A1(_AES_ENC_us21_n1117 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n707 ) );
NOR2_X2 _AES_ENC_us21_U524  ( .A1(_AES_ENC_sa21[4]), .A2(_AES_ENC_us21_n575 ), .ZN(_AES_ENC_us21_n705 ) );
NOR3_X2 _AES_ENC_us21_U523  ( .A1(_AES_ENC_us21_n707 ), .A2(_AES_ENC_us21_n706 ), .A3(_AES_ENC_us21_n705 ), .ZN(_AES_ENC_us21_n713 ) );
INV_X4 _AES_ENC_us21_U522  ( .A(_AES_ENC_sa21[3]), .ZN(_AES_ENC_us21_n624 ));
NAND3_X2 _AES_ENC_us21_U521  ( .A1(_AES_ENC_us21_n652 ), .A2(_AES_ENC_us21_n594 ), .A3(_AES_ENC_sa21[7]), .ZN(_AES_ENC_us21_n653 ));
NOR2_X2 _AES_ENC_us21_U520  ( .A1(_AES_ENC_us21_n584 ), .A2(_AES_ENC_sa21[5]), .ZN(_AES_ENC_us21_n925 ) );
NOR2_X2 _AES_ENC_us21_U519  ( .A1(_AES_ENC_sa21[5]), .A2(_AES_ENC_sa21[2]),.ZN(_AES_ENC_us21_n974 ) );
INV_X4 _AES_ENC_us21_U518  ( .A(_AES_ENC_sa21[5]), .ZN(_AES_ENC_us21_n594 ));
NOR2_X2 _AES_ENC_us21_U517  ( .A1(_AES_ENC_us21_n584 ), .A2(_AES_ENC_sa21[7]), .ZN(_AES_ENC_us21_n779 ) );
NAND3_X2 _AES_ENC_us21_U516  ( .A1(_AES_ENC_us21_n679 ), .A2(_AES_ENC_us21_n678 ), .A3(_AES_ENC_us21_n677 ), .ZN(_AES_ENC_sa21_sub[0] ) );
NOR2_X2 _AES_ENC_us21_U515  ( .A1(_AES_ENC_us21_n594 ), .A2(_AES_ENC_sa21[2]), .ZN(_AES_ENC_us21_n1048 ) );
NOR4_X2 _AES_ENC_us21_U512  ( .A1(_AES_ENC_us21_n633 ), .A2(_AES_ENC_us21_n632 ), .A3(_AES_ENC_us21_n631 ), .A4(_AES_ENC_us21_n630 ), .ZN(_AES_ENC_us21_n634 ) );
NOR2_X2 _AES_ENC_us21_U510  ( .A1(_AES_ENC_us21_n629 ), .A2(_AES_ENC_us21_n628 ), .ZN(_AES_ENC_us21_n635 ) );
NAND3_X2 _AES_ENC_us21_U509  ( .A1(_AES_ENC_sa21[2]), .A2(_AES_ENC_sa21[7]), .A3(_AES_ENC_us21_n1059 ), .ZN(_AES_ENC_us21_n636 ) );
NOR2_X2 _AES_ENC_us21_U508  ( .A1(_AES_ENC_sa21[7]), .A2(_AES_ENC_sa21[2]),.ZN(_AES_ENC_us21_n794 ) );
NOR2_X2 _AES_ENC_us21_U507  ( .A1(_AES_ENC_sa21[4]), .A2(_AES_ENC_sa21[1]),.ZN(_AES_ENC_us21_n1102 ) );
NOR2_X2 _AES_ENC_us21_U506  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_sa21[3]), .ZN(_AES_ENC_us21_n1053 ) );
NOR2_X2 _AES_ENC_us21_U505  ( .A1(_AES_ENC_us21_n579 ), .A2(_AES_ENC_sa21[5]), .ZN(_AES_ENC_us21_n1024 ) );
NOR2_X2 _AES_ENC_us21_U504  ( .A1(_AES_ENC_us21_n593 ), .A2(_AES_ENC_sa21[2]), .ZN(_AES_ENC_us21_n1093 ) );
NOR2_X2 _AES_ENC_us21_U503  ( .A1(_AES_ENC_us21_n588 ), .A2(_AES_ENC_sa21[5]), .ZN(_AES_ENC_us21_n1094 ) );
NOR2_X2 _AES_ENC_us21_U502  ( .A1(_AES_ENC_us21_n612 ), .A2(_AES_ENC_sa21[3]), .ZN(_AES_ENC_us21_n931 ) );
INV_X4 _AES_ENC_us21_U501  ( .A(_AES_ENC_us21_n570 ), .ZN(_AES_ENC_us21_n573 ) );
NOR2_X2 _AES_ENC_us21_U500  ( .A1(_AES_ENC_us21_n1053 ), .A2(_AES_ENC_us21_n1095 ), .ZN(_AES_ENC_us21_n639 ) );
NOR3_X2 _AES_ENC_us21_U499  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n573 ), .A3(_AES_ENC_us21_n1074 ), .ZN(_AES_ENC_us21_n641 ) );
NOR2_X2 _AES_ENC_us21_U498  ( .A1(_AES_ENC_us21_n639 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n640 ) );
NOR2_X2 _AES_ENC_us21_U497  ( .A1(_AES_ENC_us21_n641 ), .A2(_AES_ENC_us21_n640 ), .ZN(_AES_ENC_us21_n646 ) );
NOR3_X2 _AES_ENC_us21_U496  ( .A1(_AES_ENC_us21_n995 ), .A2(_AES_ENC_us21_n580 ), .A3(_AES_ENC_us21_n994 ), .ZN(_AES_ENC_us21_n1002 ) );
NOR2_X2 _AES_ENC_us21_U495  ( .A1(_AES_ENC_us21_n909 ), .A2(_AES_ENC_us21_n908 ), .ZN(_AES_ENC_us21_n920 ) );
NOR2_X2 _AES_ENC_us21_U494  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n823 ) );
NOR2_X2 _AES_ENC_us21_U492  ( .A1(_AES_ENC_us21_n612 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n822 ) );
NOR2_X2 _AES_ENC_us21_U491  ( .A1(_AES_ENC_us21_n823 ), .A2(_AES_ENC_us21_n822 ), .ZN(_AES_ENC_us21_n825 ) );
NOR2_X2 _AES_ENC_us21_U490  ( .A1(_AES_ENC_sa21[1]), .A2(_AES_ENC_us21_n601 ), .ZN(_AES_ENC_us21_n913 ) );
NOR2_X2 _AES_ENC_us21_U489  ( .A1(_AES_ENC_us21_n913 ), .A2(_AES_ENC_us21_n1091 ), .ZN(_AES_ENC_us21_n914 ) );
NOR2_X2 _AES_ENC_us21_U488  ( .A1(_AES_ENC_us21_n826 ), .A2(_AES_ENC_us21_n572 ), .ZN(_AES_ENC_us21_n827 ) );
NOR3_X2 _AES_ENC_us21_U487  ( .A1(_AES_ENC_us21_n769 ), .A2(_AES_ENC_us21_n768 ), .A3(_AES_ENC_us21_n767 ), .ZN(_AES_ENC_us21_n775 ) );
NOR2_X2 _AES_ENC_us21_U486  ( .A1(_AES_ENC_us21_n1056 ), .A2(_AES_ENC_us21_n1053 ), .ZN(_AES_ENC_us21_n749 ) );
NOR2_X2 _AES_ENC_us21_U483  ( .A1(_AES_ENC_us21_n749 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n752 ) );
INV_X4 _AES_ENC_us21_U482  ( .A(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n626 ));
NOR2_X2 _AES_ENC_us21_U480  ( .A1(_AES_ENC_us21_n1054 ), .A2(_AES_ENC_us21_n1053 ), .ZN(_AES_ENC_us21_n1055 ) );
OR2_X4 _AES_ENC_us21_U479  ( .A1(_AES_ENC_us21_n1094 ), .A2(_AES_ENC_us21_n1093 ), .ZN(_AES_ENC_us21_n571 ) );
AND2_X2 _AES_ENC_us21_U478  ( .A1(_AES_ENC_us21_n571 ), .A2(_AES_ENC_us21_n1095 ), .ZN(_AES_ENC_us21_n1101 ) );
NOR2_X2 _AES_ENC_us21_U477  ( .A1(_AES_ENC_us21_n1074 ), .A2(_AES_ENC_us21_n931 ), .ZN(_AES_ENC_us21_n796 ) );
NOR2_X2 _AES_ENC_us21_U474  ( .A1(_AES_ENC_us21_n796 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n797 ) );
NOR2_X2 _AES_ENC_us21_U473  ( .A1(_AES_ENC_us21_n932 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n933 ) );
NOR2_X2 _AES_ENC_us21_U472  ( .A1(_AES_ENC_us21_n929 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n935 ) );
NOR2_X2 _AES_ENC_us21_U471  ( .A1(_AES_ENC_us21_n931 ), .A2(_AES_ENC_us21_n930 ), .ZN(_AES_ENC_us21_n934 ) );
NOR3_X2 _AES_ENC_us21_U470  ( .A1(_AES_ENC_us21_n935 ), .A2(_AES_ENC_us21_n934 ), .A3(_AES_ENC_us21_n933 ), .ZN(_AES_ENC_us21_n936 ) );
NOR2_X2 _AES_ENC_us21_U469  ( .A1(_AES_ENC_us21_n612 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n1075 ) );
NOR2_X2 _AES_ENC_us21_U468  ( .A1(_AES_ENC_us21_n572 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n949 ) );
NOR2_X2 _AES_ENC_us21_U467  ( .A1(_AES_ENC_us21_n1049 ), .A2(_AES_ENC_us21_n592 ), .ZN(_AES_ENC_us21_n1051 ) );
NOR2_X2 _AES_ENC_us21_U466  ( .A1(_AES_ENC_us21_n1051 ), .A2(_AES_ENC_us21_n1050 ), .ZN(_AES_ENC_us21_n1052 ) );
NOR2_X2 _AES_ENC_us21_U465  ( .A1(_AES_ENC_us21_n1052 ), .A2(_AES_ENC_us21_n604 ), .ZN(_AES_ENC_us21_n1064 ) );
NOR2_X2 _AES_ENC_us21_U464  ( .A1(_AES_ENC_sa21[1]), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n631 ) );
NOR2_X2 _AES_ENC_us21_U463  ( .A1(_AES_ENC_us21_n1025 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n980 ) );
NOR2_X2 _AES_ENC_us21_U462  ( .A1(_AES_ENC_us21_n1073 ), .A2(_AES_ENC_us21_n1094 ), .ZN(_AES_ENC_us21_n795 ) );
NOR2_X2 _AES_ENC_us21_U461  ( .A1(_AES_ENC_us21_n795 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n799 ) );
NOR2_X2 _AES_ENC_us21_U460  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n981 ) );
NOR2_X2 _AES_ENC_us21_U459  ( .A1(_AES_ENC_us21_n1102 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n643 ) );
NOR2_X2 _AES_ENC_us21_U458  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n624 ), .ZN(_AES_ENC_us21_n642 ) );
NOR2_X2 _AES_ENC_us21_U455  ( .A1(_AES_ENC_us21_n911 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n644 ) );
NOR4_X2 _AES_ENC_us21_U448  ( .A1(_AES_ENC_us21_n644 ), .A2(_AES_ENC_us21_n643 ), .A3(_AES_ENC_us21_n804 ), .A4(_AES_ENC_us21_n642 ), .ZN(_AES_ENC_us21_n645 ) );
NOR2_X2 _AES_ENC_us21_U447  ( .A1(_AES_ENC_us21_n1102 ), .A2(_AES_ENC_us21_n910 ), .ZN(_AES_ENC_us21_n932 ) );
NOR2_X2 _AES_ENC_us21_U442  ( .A1(_AES_ENC_us21_n1102 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n755 ) );
NOR2_X2 _AES_ENC_us21_U441  ( .A1(_AES_ENC_us21_n931 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n743 ) );
NOR2_X2 _AES_ENC_us21_U438  ( .A1(_AES_ENC_us21_n1072 ), .A2(_AES_ENC_us21_n1094 ), .ZN(_AES_ENC_us21_n930 ) );
NOR2_X2 _AES_ENC_us21_U435  ( .A1(_AES_ENC_us21_n1074 ), .A2(_AES_ENC_us21_n1025 ), .ZN(_AES_ENC_us21_n891 ) );
NOR2_X2 _AES_ENC_us21_U434  ( .A1(_AES_ENC_us21_n891 ), .A2(_AES_ENC_us21_n582 ), .ZN(_AES_ENC_us21_n894 ) );
NOR3_X2 _AES_ENC_us21_U433  ( .A1(_AES_ENC_us21_n601 ), .A2(_AES_ENC_sa21[1]), .A3(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n683 ));
INV_X4 _AES_ENC_us21_U428  ( .A(_AES_ENC_us21_n931 ), .ZN(_AES_ENC_us21_n601 ) );
NOR2_X2 _AES_ENC_us21_U427  ( .A1(_AES_ENC_us21_n996 ), .A2(_AES_ENC_us21_n931 ), .ZN(_AES_ENC_us21_n704 ) );
NOR2_X2 _AES_ENC_us21_U421  ( .A1(_AES_ENC_us21_n931 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n685 ) );
NOR2_X2 _AES_ENC_us21_U420  ( .A1(_AES_ENC_us21_n1029 ), .A2(_AES_ENC_us21_n1025 ), .ZN(_AES_ENC_us21_n1079 ) );
NOR3_X2 _AES_ENC_us21_U419  ( .A1(_AES_ENC_us21_n620 ), .A2(_AES_ENC_us21_n1025 ), .A3(_AES_ENC_us21_n590 ), .ZN(_AES_ENC_us21_n945 ) );
NOR2_X2 _AES_ENC_us21_U418  ( .A1(_AES_ENC_us21_n594 ), .A2(_AES_ENC_us21_n584 ), .ZN(_AES_ENC_us21_n800 ) );
NOR3_X2 _AES_ENC_us21_U417  ( .A1(_AES_ENC_us21_n598 ), .A2(_AES_ENC_us21_n595 ), .A3(_AES_ENC_us21_n584 ), .ZN(_AES_ENC_us21_n798 ) );
NOR3_X2 _AES_ENC_us21_U416  ( .A1(_AES_ENC_us21_n583 ), .A2(_AES_ENC_us21_n572 ), .A3(_AES_ENC_us21_n596 ), .ZN(_AES_ENC_us21_n962 ) );
NOR3_X2 _AES_ENC_us21_U415  ( .A1(_AES_ENC_us21_n959 ), .A2(_AES_ENC_us21_n572 ), .A3(_AES_ENC_us21_n582 ), .ZN(_AES_ENC_us21_n768 ) );
NOR3_X2 _AES_ENC_us21_U414  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n572 ), .A3(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n694 ) );
NOR3_X2 _AES_ENC_us21_U413  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n572 ), .A3(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n895 ) );
NOR3_X2 _AES_ENC_us21_U410  ( .A1(_AES_ENC_us21_n1008 ), .A2(_AES_ENC_us21_n1007 ), .A3(_AES_ENC_us21_n1006 ), .ZN(_AES_ENC_us21_n1018 ) );
NOR4_X2 _AES_ENC_us21_U409  ( .A1(_AES_ENC_us21_n806 ), .A2(_AES_ENC_us21_n805 ), .A3(_AES_ENC_us21_n804 ), .A4(_AES_ENC_us21_n803 ), .ZN(_AES_ENC_us21_n807 ) );
NOR3_X2 _AES_ENC_us21_U406  ( .A1(_AES_ENC_us21_n799 ), .A2(_AES_ENC_us21_n798 ), .A3(_AES_ENC_us21_n797 ), .ZN(_AES_ENC_us21_n808 ) );
NOR4_X2 _AES_ENC_us21_U405  ( .A1(_AES_ENC_us21_n843 ), .A2(_AES_ENC_us21_n842 ), .A3(_AES_ENC_us21_n841 ), .A4(_AES_ENC_us21_n840 ), .ZN(_AES_ENC_us21_n844 ) );
NOR2_X2 _AES_ENC_us21_U404  ( .A1(_AES_ENC_us21_n669 ), .A2(_AES_ENC_us21_n668 ), .ZN(_AES_ENC_us21_n673 ) );
NOR4_X2 _AES_ENC_us21_U403  ( .A1(_AES_ENC_us21_n946 ), .A2(_AES_ENC_us21_n1046 ), .A3(_AES_ENC_us21_n671 ), .A4(_AES_ENC_us21_n670 ), .ZN(_AES_ENC_us21_n672 ) );
NOR4_X2 _AES_ENC_us21_U401  ( .A1(_AES_ENC_us21_n711 ), .A2(_AES_ENC_us21_n710 ), .A3(_AES_ENC_us21_n709 ), .A4(_AES_ENC_us21_n708 ), .ZN(_AES_ENC_us21_n712 ) );
NOR4_X2 _AES_ENC_us21_U400  ( .A1(_AES_ENC_us21_n963 ), .A2(_AES_ENC_us21_n962 ), .A3(_AES_ENC_us21_n961 ), .A4(_AES_ENC_us21_n960 ), .ZN(_AES_ENC_us21_n964 ) );
NOR3_X2 _AES_ENC_us21_U399  ( .A1(_AES_ENC_us21_n1101 ), .A2(_AES_ENC_us21_n1100 ), .A3(_AES_ENC_us21_n1099 ), .ZN(_AES_ENC_us21_n1109 ) );
NOR3_X2 _AES_ENC_us21_U398  ( .A1(_AES_ENC_us21_n743 ), .A2(_AES_ENC_us21_n742 ), .A3(_AES_ENC_us21_n741 ), .ZN(_AES_ENC_us21_n744 ) );
NOR2_X2 _AES_ENC_us21_U397  ( .A1(_AES_ENC_us21_n697 ), .A2(_AES_ENC_us21_n658 ), .ZN(_AES_ENC_us21_n659 ) );
NOR2_X2 _AES_ENC_us21_U396  ( .A1(_AES_ENC_us21_n1078 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n1033 ) );
NOR2_X2 _AES_ENC_us21_U393  ( .A1(_AES_ENC_us21_n1031 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n1032 ) );
NOR3_X2 _AES_ENC_us21_U390  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n1025 ), .A3(_AES_ENC_us21_n1074 ), .ZN(_AES_ENC_us21_n1035 ) );
NOR4_X2 _AES_ENC_us21_U389  ( .A1(_AES_ENC_us21_n1035 ), .A2(_AES_ENC_us21_n1034 ), .A3(_AES_ENC_us21_n1033 ), .A4(_AES_ENC_us21_n1032 ), .ZN(_AES_ENC_us21_n1036 ) );
NOR2_X2 _AES_ENC_us21_U388  ( .A1(_AES_ENC_us21_n611 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n885 ) );
NOR2_X2 _AES_ENC_us21_U387  ( .A1(_AES_ENC_us21_n601 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n882 ) );
NOR2_X2 _AES_ENC_us21_U386  ( .A1(_AES_ENC_us21_n1053 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n884 ) );
NOR4_X2 _AES_ENC_us21_U385  ( .A1(_AES_ENC_us21_n885 ), .A2(_AES_ENC_us21_n884 ), .A3(_AES_ENC_us21_n883 ), .A4(_AES_ENC_us21_n882 ), .ZN(_AES_ENC_us21_n886 ) );
NOR2_X2 _AES_ENC_us21_U384  ( .A1(_AES_ENC_us21_n825 ), .A2(_AES_ENC_us21_n574 ), .ZN(_AES_ENC_us21_n830 ) );
NOR2_X2 _AES_ENC_us21_U383  ( .A1(_AES_ENC_us21_n827 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n829 ) );
NOR2_X2 _AES_ENC_us21_U382  ( .A1(_AES_ENC_us21_n572 ), .A2(_AES_ENC_us21_n575 ), .ZN(_AES_ENC_us21_n828 ) );
NOR4_X2 _AES_ENC_us21_U374  ( .A1(_AES_ENC_us21_n831 ), .A2(_AES_ENC_us21_n830 ), .A3(_AES_ENC_us21_n829 ), .A4(_AES_ENC_us21_n828 ), .ZN(_AES_ENC_us21_n832 ) );
NOR2_X2 _AES_ENC_us21_U373  ( .A1(_AES_ENC_us21_n578 ), .A2(_AES_ENC_us21_n603 ), .ZN(_AES_ENC_us21_n1104 ) );
NOR2_X2 _AES_ENC_us21_U372  ( .A1(_AES_ENC_us21_n1102 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n1106 ) );
NOR2_X2 _AES_ENC_us21_U370  ( .A1(_AES_ENC_us21_n1103 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n1105 ) );
NOR4_X2 _AES_ENC_us21_U369  ( .A1(_AES_ENC_us21_n1107 ), .A2(_AES_ENC_us21_n1106 ), .A3(_AES_ENC_us21_n1105 ), .A4(_AES_ENC_us21_n1104 ), .ZN(_AES_ENC_us21_n1108 ) );
NOR3_X2 _AES_ENC_us21_U368  ( .A1(_AES_ENC_us21_n959 ), .A2(_AES_ENC_us21_n624 ), .A3(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n963 ) );
NOR2_X2 _AES_ENC_us21_U367  ( .A1(_AES_ENC_us21_n594 ), .A2(_AES_ENC_us21_n595 ), .ZN(_AES_ENC_us21_n1114 ) );
INV_X4 _AES_ENC_us21_U366  ( .A(_AES_ENC_us21_n1024 ), .ZN(_AES_ENC_us21_n578 ) );
NOR3_X2 _AES_ENC_us21_U365  ( .A1(_AES_ENC_us21_n910 ), .A2(_AES_ENC_us21_n1059 ), .A3(_AES_ENC_us21_n584 ), .ZN(_AES_ENC_us21_n1115 ) );
INV_X4 _AES_ENC_us21_U364  ( .A(_AES_ENC_us21_n1094 ), .ZN(_AES_ENC_us21_n587 ) );
NOR2_X2 _AES_ENC_us21_U363  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n931 ), .ZN(_AES_ENC_us21_n1100 ) );
INV_X4 _AES_ENC_us21_U354  ( .A(_AES_ENC_us21_n1093 ), .ZN(_AES_ENC_us21_n591 ) );
NOR2_X2 _AES_ENC_us21_U353  ( .A1(_AES_ENC_us21_n569 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n929 ) );
NOR2_X2 _AES_ENC_us21_U352  ( .A1(_AES_ENC_us21_n609 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n926 ) );
NOR2_X2 _AES_ENC_us21_U351  ( .A1(_AES_ENC_us21_n572 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n1095 ) );
NOR2_X2 _AES_ENC_us21_U350  ( .A1(_AES_ENC_us21_n582 ), .A2(_AES_ENC_us21_n595 ), .ZN(_AES_ENC_us21_n1010 ) );
NOR2_X2 _AES_ENC_us21_U349  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n1103 ) );
NOR2_X2 _AES_ENC_us21_U348  ( .A1(_AES_ENC_us21_n614 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n1059 ) );
NOR2_X2 _AES_ENC_us21_U347  ( .A1(_AES_ENC_sa21[1]), .A2(_AES_ENC_us21_n1120 ), .ZN(_AES_ENC_us21_n1022 ) );
NOR2_X2 _AES_ENC_us21_U346  ( .A1(_AES_ENC_us21_n605 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n911 ) );
NOR2_X2 _AES_ENC_us21_U345  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_us21_n1025 ), .ZN(_AES_ENC_us21_n826 ) );
NOR2_X2 _AES_ENC_us21_U338  ( .A1(_AES_ENC_us21_n594 ), .A2(_AES_ENC_us21_n579 ), .ZN(_AES_ENC_us21_n1072 ) );
NOR2_X2 _AES_ENC_us21_U335  ( .A1(_AES_ENC_us21_n595 ), .A2(_AES_ENC_us21_n590 ), .ZN(_AES_ENC_us21_n956 ) );
NOR2_X2 _AES_ENC_us21_U329  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_us21_n612 ), .ZN(_AES_ENC_us21_n1121 ) );
NOR2_X2 _AES_ENC_us21_U328  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_us21_n612 ), .ZN(_AES_ENC_us21_n1058 ) );
NOR2_X2 _AES_ENC_us21_U327  ( .A1(_AES_ENC_us21_n593 ), .A2(_AES_ENC_us21_n584 ), .ZN(_AES_ENC_us21_n1073 ) );
NOR2_X2 _AES_ENC_us21_U325  ( .A1(_AES_ENC_sa21[1]), .A2(_AES_ENC_us21_n1025 ), .ZN(_AES_ENC_us21_n1054 ) );
NOR2_X2 _AES_ENC_us21_U324  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_us21_n931 ), .ZN(_AES_ENC_us21_n1029 ) );
NOR2_X2 _AES_ENC_us21_U319  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n1056 ) );
NOR2_X2 _AES_ENC_us21_U318  ( .A1(_AES_ENC_us21_n588 ), .A2(_AES_ENC_us21_n594 ), .ZN(_AES_ENC_us21_n1050 ) );
NOR2_X2 _AES_ENC_us21_U317  ( .A1(_AES_ENC_us21_n1121 ), .A2(_AES_ENC_us21_n1025 ), .ZN(_AES_ENC_us21_n1120 ) );
NOR2_X2 _AES_ENC_us21_U316  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_us21_n572 ), .ZN(_AES_ENC_us21_n1074 ) );
NOR2_X2 _AES_ENC_us21_U315  ( .A1(_AES_ENC_us21_n1058 ), .A2(_AES_ENC_us21_n1054 ), .ZN(_AES_ENC_us21_n878 ) );
NOR2_X2 _AES_ENC_us21_U314  ( .A1(_AES_ENC_us21_n878 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n879 ) );
NOR2_X2 _AES_ENC_us21_U312  ( .A1(_AES_ENC_us21_n880 ), .A2(_AES_ENC_us21_n879 ), .ZN(_AES_ENC_us21_n887 ) );
NOR2_X2 _AES_ENC_us21_U311  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n625 ), .ZN(_AES_ENC_us21_n957 ) );
NOR2_X2 _AES_ENC_us21_U310  ( .A1(_AES_ENC_us21_n958 ), .A2(_AES_ENC_us21_n957 ), .ZN(_AES_ENC_us21_n965 ) );
NOR3_X2 _AES_ENC_us21_U309  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n1091 ), .A3(_AES_ENC_us21_n1022 ), .ZN(_AES_ENC_us21_n720 ) );
NOR3_X2 _AES_ENC_us21_U303  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n1054 ), .A3(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n719 ) );
NOR2_X2 _AES_ENC_us21_U302  ( .A1(_AES_ENC_us21_n720 ), .A2(_AES_ENC_us21_n719 ), .ZN(_AES_ENC_us21_n726 ) );
NOR2_X2 _AES_ENC_us21_U300  ( .A1(_AES_ENC_us21_n588 ), .A2(_AES_ENC_us21_n613 ), .ZN(_AES_ENC_us21_n865 ) );
NOR2_X2 _AES_ENC_us21_U299  ( .A1(_AES_ENC_us21_n1059 ), .A2(_AES_ENC_us21_n1058 ), .ZN(_AES_ENC_us21_n1060 ) );
NOR2_X2 _AES_ENC_us21_U298  ( .A1(_AES_ENC_us21_n1095 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n668 ) );
NOR2_X2 _AES_ENC_us21_U297  ( .A1(_AES_ENC_us21_n826 ), .A2(_AES_ENC_us21_n573 ), .ZN(_AES_ENC_us21_n750 ) );
NOR2_X2 _AES_ENC_us21_U296  ( .A1(_AES_ENC_us21_n750 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n751 ) );
NOR2_X2 _AES_ENC_us21_U295  ( .A1(_AES_ENC_us21_n907 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n908 ) );
NOR2_X2 _AES_ENC_us21_U294  ( .A1(_AES_ENC_us21_n990 ), .A2(_AES_ENC_us21_n926 ), .ZN(_AES_ENC_us21_n780 ) );
NOR2_X2 _AES_ENC_us21_U293  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n606 ), .ZN(_AES_ENC_us21_n838 ) );
NOR2_X2 _AES_ENC_us21_U292  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n621 ), .ZN(_AES_ENC_us21_n837 ) );
NOR2_X2 _AES_ENC_us21_U291  ( .A1(_AES_ENC_us21_n838 ), .A2(_AES_ENC_us21_n837 ), .ZN(_AES_ENC_us21_n845 ) );
NOR2_X2 _AES_ENC_us21_U290  ( .A1(_AES_ENC_us21_n1022 ), .A2(_AES_ENC_us21_n1058 ), .ZN(_AES_ENC_us21_n740 ) );
NOR2_X2 _AES_ENC_us21_U284  ( .A1(_AES_ENC_us21_n740 ), .A2(_AES_ENC_us21_n590 ), .ZN(_AES_ENC_us21_n742 ) );
NOR2_X2 _AES_ENC_us21_U283  ( .A1(_AES_ENC_us21_n1098 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n1099 ) );
NOR2_X2 _AES_ENC_us21_U282  ( .A1(_AES_ENC_us21_n1120 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n993 ) );
NOR2_X2 _AES_ENC_us21_U281  ( .A1(_AES_ENC_us21_n993 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n994 ) );
NOR2_X2 _AES_ENC_us21_U280  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n609 ), .ZN(_AES_ENC_us21_n1026 ) );
NOR2_X2 _AES_ENC_us21_U279  ( .A1(_AES_ENC_us21_n573 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n1027 ) );
NOR2_X2 _AES_ENC_us21_U273  ( .A1(_AES_ENC_us21_n1027 ), .A2(_AES_ENC_us21_n1026 ), .ZN(_AES_ENC_us21_n1028 ) );
NOR2_X2 _AES_ENC_us21_U272  ( .A1(_AES_ENC_us21_n1029 ), .A2(_AES_ENC_us21_n1028 ), .ZN(_AES_ENC_us21_n1034 ) );
NOR4_X2 _AES_ENC_us21_U271  ( .A1(_AES_ENC_us21_n757 ), .A2(_AES_ENC_us21_n756 ), .A3(_AES_ENC_us21_n755 ), .A4(_AES_ENC_us21_n754 ), .ZN(_AES_ENC_us21_n758 ) );
NOR2_X2 _AES_ENC_us21_U270  ( .A1(_AES_ENC_us21_n752 ), .A2(_AES_ENC_us21_n751 ), .ZN(_AES_ENC_us21_n759 ) );
NOR2_X2 _AES_ENC_us21_U269  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n1071 ), .ZN(_AES_ENC_us21_n669 ) );
NOR2_X2 _AES_ENC_us21_U268  ( .A1(_AES_ENC_us21_n1056 ), .A2(_AES_ENC_us21_n990 ), .ZN(_AES_ENC_us21_n991 ) );
NOR2_X2 _AES_ENC_us21_U267  ( .A1(_AES_ENC_us21_n991 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n995 ) );
NOR2_X2 _AES_ENC_us21_U263  ( .A1(_AES_ENC_us21_n579 ), .A2(_AES_ENC_us21_n598 ), .ZN(_AES_ENC_us21_n1008 ) );
NOR2_X2 _AES_ENC_us21_U262  ( .A1(_AES_ENC_us21_n839 ), .A2(_AES_ENC_us21_n603 ), .ZN(_AES_ENC_us21_n693 ) );
NOR2_X2 _AES_ENC_us21_U258  ( .A1(_AES_ENC_us21_n578 ), .A2(_AES_ENC_us21_n906 ), .ZN(_AES_ENC_us21_n741 ) );
NOR2_X2 _AES_ENC_us21_U255  ( .A1(_AES_ENC_us21_n1054 ), .A2(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n763 ) );
NOR2_X2 _AES_ENC_us21_U254  ( .A1(_AES_ENC_us21_n763 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n769 ) );
NOR2_X2 _AES_ENC_us21_U253  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n618 ), .ZN(_AES_ENC_us21_n1007 ) );
NOR2_X2 _AES_ENC_us21_U252  ( .A1(_AES_ENC_us21_n582 ), .A2(_AES_ENC_us21_n599 ), .ZN(_AES_ENC_us21_n1123 ) );
NOR2_X2 _AES_ENC_us21_U251  ( .A1(_AES_ENC_us21_n582 ), .A2(_AES_ENC_us21_n598 ), .ZN(_AES_ENC_us21_n710 ) );
INV_X4 _AES_ENC_us21_U250  ( .A(_AES_ENC_us21_n1029 ), .ZN(_AES_ENC_us21_n603 ) );
NOR2_X2 _AES_ENC_us21_U243  ( .A1(_AES_ENC_us21_n590 ), .A2(_AES_ENC_us21_n607 ), .ZN(_AES_ENC_us21_n883 ) );
NOR2_X2 _AES_ENC_us21_U242  ( .A1(_AES_ENC_us21_n623 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n1125 ) );
NOR2_X2 _AES_ENC_us21_U241  ( .A1(_AES_ENC_us21_n911 ), .A2(_AES_ENC_us21_n910 ), .ZN(_AES_ENC_us21_n912 ) );
NOR2_X2 _AES_ENC_us21_U240  ( .A1(_AES_ENC_us21_n912 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n916 ) );
NOR2_X2 _AES_ENC_us21_U239  ( .A1(_AES_ENC_us21_n990 ), .A2(_AES_ENC_us21_n929 ), .ZN(_AES_ENC_us21_n892 ) );
NOR2_X2 _AES_ENC_us21_U238  ( .A1(_AES_ENC_us21_n892 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n893 ) );
NOR2_X2 _AES_ENC_us21_U237  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n621 ), .ZN(_AES_ENC_us21_n950 ) );
NOR2_X2 _AES_ENC_us21_U236  ( .A1(_AES_ENC_us21_n1079 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n1082 ) );
NOR2_X2 _AES_ENC_us21_U235  ( .A1(_AES_ENC_us21_n910 ), .A2(_AES_ENC_us21_n1056 ), .ZN(_AES_ENC_us21_n941 ) );
NOR2_X2 _AES_ENC_us21_U234  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n1077 ), .ZN(_AES_ENC_us21_n841 ) );
NOR2_X2 _AES_ENC_us21_U229  ( .A1(_AES_ENC_us21_n601 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n630 ) );
NOR2_X2 _AES_ENC_us21_U228  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n621 ), .ZN(_AES_ENC_us21_n806 ) );
NOR2_X2 _AES_ENC_us21_U227  ( .A1(_AES_ENC_us21_n601 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n948 ) );
NOR2_X2 _AES_ENC_us21_U226  ( .A1(_AES_ENC_us21_n578 ), .A2(_AES_ENC_us21_n620 ), .ZN(_AES_ENC_us21_n997 ) );
NOR2_X2 _AES_ENC_us21_U225  ( .A1(_AES_ENC_us21_n1121 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n1122 ) );
NOR2_X2 _AES_ENC_us21_U223  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n1023 ), .ZN(_AES_ENC_us21_n756 ) );
NOR2_X2 _AES_ENC_us21_U222  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n621 ), .ZN(_AES_ENC_us21_n870 ) );
NOR2_X2 _AES_ENC_us21_U221  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n569 ), .ZN(_AES_ENC_us21_n947 ) );
NOR2_X2 _AES_ENC_us21_U217  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n1077 ), .ZN(_AES_ENC_us21_n1084 ) );
NOR2_X2 _AES_ENC_us21_U213  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n855 ), .ZN(_AES_ENC_us21_n709 ) );
NOR2_X2 _AES_ENC_us21_U212  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n620 ), .ZN(_AES_ENC_us21_n868 ) );
NOR2_X2 _AES_ENC_us21_U211  ( .A1(_AES_ENC_us21_n1120 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n1124 ) );
NOR2_X2 _AES_ENC_us21_U210  ( .A1(_AES_ENC_us21_n1120 ), .A2(_AES_ENC_us21_n839 ), .ZN(_AES_ENC_us21_n842 ) );
NOR2_X2 _AES_ENC_us21_U209  ( .A1(_AES_ENC_us21_n1120 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n696 ) );
NOR2_X2 _AES_ENC_us21_U208  ( .A1(_AES_ENC_us21_n1074 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n1076 ) );
NOR2_X2 _AES_ENC_us21_U207  ( .A1(_AES_ENC_us21_n1074 ), .A2(_AES_ENC_us21_n609 ), .ZN(_AES_ENC_us21_n781 ) );
NOR3_X2 _AES_ENC_us21_U201  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n1056 ), .A3(_AES_ENC_us21_n990 ), .ZN(_AES_ENC_us21_n979 ) );
NOR3_X2 _AES_ENC_us21_U200  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n1058 ), .A3(_AES_ENC_us21_n1059 ), .ZN(_AES_ENC_us21_n854 ) );
NOR2_X2 _AES_ENC_us21_U199  ( .A1(_AES_ENC_us21_n996 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n869 ) );
NOR2_X2 _AES_ENC_us21_U198  ( .A1(_AES_ENC_us21_n1056 ), .A2(_AES_ENC_us21_n1074 ), .ZN(_AES_ENC_us21_n1057 ) );
NOR3_X2 _AES_ENC_us21_U197  ( .A1(_AES_ENC_us21_n579 ), .A2(_AES_ENC_us21_n1120 ), .A3(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n978 ) );
NOR2_X2 _AES_ENC_us21_U196  ( .A1(_AES_ENC_us21_n996 ), .A2(_AES_ENC_us21_n911 ), .ZN(_AES_ENC_us21_n1116 ) );
NOR2_X2 _AES_ENC_us21_U195  ( .A1(_AES_ENC_us21_n1074 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n754 ) );
NOR2_X2 _AES_ENC_us21_U194  ( .A1(_AES_ENC_us21_n926 ), .A2(_AES_ENC_us21_n1103 ), .ZN(_AES_ENC_us21_n977 ) );
NOR2_X2 _AES_ENC_us21_U187  ( .A1(_AES_ENC_us21_n839 ), .A2(_AES_ENC_us21_n824 ), .ZN(_AES_ENC_us21_n1092 ) );
NOR2_X2 _AES_ENC_us21_U186  ( .A1(_AES_ENC_us21_n573 ), .A2(_AES_ENC_us21_n1074 ), .ZN(_AES_ENC_us21_n684 ) );
NOR2_X2 _AES_ENC_us21_U185  ( .A1(_AES_ENC_us21_n826 ), .A2(_AES_ENC_us21_n1059 ), .ZN(_AES_ENC_us21_n907 ) );
NOR3_X2 _AES_ENC_us21_U184  ( .A1(_AES_ENC_us21_n593 ), .A2(_AES_ENC_us21_n1115 ), .A3(_AES_ENC_us21_n600 ), .ZN(_AES_ENC_us21_n831 ) );
NOR3_X2 _AES_ENC_us21_U183  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n1056 ), .A3(_AES_ENC_us21_n990 ), .ZN(_AES_ENC_us21_n896 ) );
NOR3_X2 _AES_ENC_us21_U182  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n573 ), .A3(_AES_ENC_us21_n1013 ), .ZN(_AES_ENC_us21_n670 ) );
NOR3_X2 _AES_ENC_us21_U181  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n1091 ), .A3(_AES_ENC_us21_n1022 ), .ZN(_AES_ENC_us21_n843 ) );
NOR2_X2 _AES_ENC_us21_U180  ( .A1(_AES_ENC_us21_n1029 ), .A2(_AES_ENC_us21_n1095 ), .ZN(_AES_ENC_us21_n735 ) );
NOR2_X2 _AES_ENC_us21_U174  ( .A1(_AES_ENC_us21_n1100 ), .A2(_AES_ENC_us21_n854 ), .ZN(_AES_ENC_us21_n860 ) );
NAND3_X2 _AES_ENC_us21_U173  ( .A1(_AES_ENC_us21_n569 ), .A2(_AES_ENC_us21_n603 ), .A3(_AES_ENC_us21_n681 ), .ZN(_AES_ENC_us21_n691 ) );
NOR2_X2 _AES_ENC_us21_U172  ( .A1(_AES_ENC_us21_n683 ), .A2(_AES_ENC_us21_n682 ), .ZN(_AES_ENC_us21_n690 ) );
NOR3_X2 _AES_ENC_us21_U171  ( .A1(_AES_ENC_us21_n695 ), .A2(_AES_ENC_us21_n694 ), .A3(_AES_ENC_us21_n693 ), .ZN(_AES_ENC_us21_n700 ) );
NOR4_X2 _AES_ENC_us21_U170  ( .A1(_AES_ENC_us21_n983 ), .A2(_AES_ENC_us21_n698 ), .A3(_AES_ENC_us21_n697 ), .A4(_AES_ENC_us21_n696 ), .ZN(_AES_ENC_us21_n699 ) );
NOR2_X2 _AES_ENC_us21_U169  ( .A1(_AES_ENC_us21_n946 ), .A2(_AES_ENC_us21_n945 ), .ZN(_AES_ENC_us21_n952 ) );
NOR4_X2 _AES_ENC_us21_U168  ( .A1(_AES_ENC_us21_n950 ), .A2(_AES_ENC_us21_n949 ), .A3(_AES_ENC_us21_n948 ), .A4(_AES_ENC_us21_n947 ), .ZN(_AES_ENC_us21_n951 ) );
NOR4_X2 _AES_ENC_us21_U162  ( .A1(_AES_ENC_us21_n896 ), .A2(_AES_ENC_us21_n895 ), .A3(_AES_ENC_us21_n894 ), .A4(_AES_ENC_us21_n893 ), .ZN(_AES_ENC_us21_n897 ) );
NOR2_X2 _AES_ENC_us21_U161  ( .A1(_AES_ENC_us21_n866 ), .A2(_AES_ENC_us21_n865 ), .ZN(_AES_ENC_us21_n872 ) );
NOR4_X2 _AES_ENC_us21_U160  ( .A1(_AES_ENC_us21_n870 ), .A2(_AES_ENC_us21_n869 ), .A3(_AES_ENC_us21_n868 ), .A4(_AES_ENC_us21_n867 ), .ZN(_AES_ENC_us21_n871 ) );
NOR4_X2 _AES_ENC_us21_U159  ( .A1(_AES_ENC_us21_n983 ), .A2(_AES_ENC_us21_n982 ), .A3(_AES_ENC_us21_n981 ), .A4(_AES_ENC_us21_n980 ), .ZN(_AES_ENC_us21_n984 ) );
NOR2_X2 _AES_ENC_us21_U158  ( .A1(_AES_ENC_us21_n979 ), .A2(_AES_ENC_us21_n978 ), .ZN(_AES_ENC_us21_n985 ) );
NOR4_X2 _AES_ENC_us21_U157  ( .A1(_AES_ENC_us21_n1125 ), .A2(_AES_ENC_us21_n1124 ), .A3(_AES_ENC_us21_n1123 ), .A4(_AES_ENC_us21_n1122 ), .ZN(_AES_ENC_us21_n1126 ) );
NOR4_X2 _AES_ENC_us21_U156  ( .A1(_AES_ENC_us21_n1084 ), .A2(_AES_ENC_us21_n1083 ), .A3(_AES_ENC_us21_n1082 ), .A4(_AES_ENC_us21_n1081 ), .ZN(_AES_ENC_us21_n1085 ) );
NOR2_X2 _AES_ENC_us21_U155  ( .A1(_AES_ENC_us21_n1076 ), .A2(_AES_ENC_us21_n1075 ), .ZN(_AES_ENC_us21_n1086 ) );
NOR3_X2 _AES_ENC_us21_U154  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n1054 ), .A3(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n961 ) );
NOR3_X2 _AES_ENC_us21_U153  ( .A1(_AES_ENC_us21_n609 ), .A2(_AES_ENC_us21_n1074 ), .A3(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n671 ) );
NOR2_X2 _AES_ENC_us21_U152  ( .A1(_AES_ENC_us21_n1057 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n1062 ) );
NOR2_X2 _AES_ENC_us21_U143  ( .A1(_AES_ENC_us21_n1055 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n1063 ) );
NOR2_X2 _AES_ENC_us21_U142  ( .A1(_AES_ENC_us21_n1060 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n1061 ) );
NOR4_X2 _AES_ENC_us21_U141  ( .A1(_AES_ENC_us21_n1064 ), .A2(_AES_ENC_us21_n1063 ), .A3(_AES_ENC_us21_n1062 ), .A4(_AES_ENC_us21_n1061 ), .ZN(_AES_ENC_us21_n1065 ) );
NOR3_X2 _AES_ENC_us21_U140  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n1120 ), .A3(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n918 ) );
NOR3_X2 _AES_ENC_us21_U132  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n573 ), .A3(_AES_ENC_us21_n1013 ), .ZN(_AES_ENC_us21_n917 ) );
NOR2_X2 _AES_ENC_us21_U131  ( .A1(_AES_ENC_us21_n914 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n915 ) );
NOR4_X2 _AES_ENC_us21_U130  ( .A1(_AES_ENC_us21_n918 ), .A2(_AES_ENC_us21_n917 ), .A3(_AES_ENC_us21_n916 ), .A4(_AES_ENC_us21_n915 ), .ZN(_AES_ENC_us21_n919 ) );
NOR2_X2 _AES_ENC_us21_U129  ( .A1(_AES_ENC_us21_n590 ), .A2(_AES_ENC_us21_n599 ), .ZN(_AES_ENC_us21_n771 ) );
NOR2_X2 _AES_ENC_us21_U128  ( .A1(_AES_ENC_us21_n1103 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n772 ) );
NOR2_X2 _AES_ENC_us21_U127  ( .A1(_AES_ENC_us21_n583 ), .A2(_AES_ENC_us21_n615 ), .ZN(_AES_ENC_us21_n773 ) );
NOR4_X2 _AES_ENC_us21_U126  ( .A1(_AES_ENC_us21_n773 ), .A2(_AES_ENC_us21_n772 ), .A3(_AES_ENC_us21_n771 ), .A4(_AES_ENC_us21_n770 ), .ZN(_AES_ENC_us21_n774 ) );
NOR2_X2 _AES_ENC_us21_U121  ( .A1(_AES_ENC_us21_n735 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n687 ) );
NOR2_X2 _AES_ENC_us21_U120  ( .A1(_AES_ENC_us21_n684 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n688 ) );
NOR2_X2 _AES_ENC_us21_U119  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n622 ), .ZN(_AES_ENC_us21_n686 ) );
NOR4_X2 _AES_ENC_us21_U118  ( .A1(_AES_ENC_us21_n688 ), .A2(_AES_ENC_us21_n687 ), .A3(_AES_ENC_us21_n686 ), .A4(_AES_ENC_us21_n685 ), .ZN(_AES_ENC_us21_n689 ) );
NOR2_X2 _AES_ENC_us21_U117  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n608 ), .ZN(_AES_ENC_us21_n858 ) );
NOR2_X2 _AES_ENC_us21_U116  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n855 ), .ZN(_AES_ENC_us21_n857 ) );
NOR2_X2 _AES_ENC_us21_U115  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n617 ), .ZN(_AES_ENC_us21_n856 ) );
NOR4_X2 _AES_ENC_us21_U106  ( .A1(_AES_ENC_us21_n858 ), .A2(_AES_ENC_us21_n857 ), .A3(_AES_ENC_us21_n856 ), .A4(_AES_ENC_us21_n958 ), .ZN(_AES_ENC_us21_n859 ) );
NOR2_X2 _AES_ENC_us21_U105  ( .A1(_AES_ENC_us21_n780 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n784 ) );
NOR2_X2 _AES_ENC_us21_U104  ( .A1(_AES_ENC_us21_n1117 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n782 ) );
NOR2_X2 _AES_ENC_us21_U103  ( .A1(_AES_ENC_us21_n781 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n783 ) );
NOR4_X2 _AES_ENC_us21_U102  ( .A1(_AES_ENC_us21_n880 ), .A2(_AES_ENC_us21_n784 ), .A3(_AES_ENC_us21_n783 ), .A4(_AES_ENC_us21_n782 ), .ZN(_AES_ENC_us21_n785 ) );
NOR2_X2 _AES_ENC_us21_U101  ( .A1(_AES_ENC_us21_n597 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n814 ) );
NOR2_X2 _AES_ENC_us21_U100  ( .A1(_AES_ENC_us21_n907 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n813 ) );
NOR3_X2 _AES_ENC_us21_U95  ( .A1(_AES_ENC_us21_n578 ), .A2(_AES_ENC_us21_n1058 ), .A3(_AES_ENC_us21_n1059 ), .ZN(_AES_ENC_us21_n815 ) );
NOR4_X2 _AES_ENC_us21_U94  ( .A1(_AES_ENC_us21_n815 ), .A2(_AES_ENC_us21_n814 ), .A3(_AES_ENC_us21_n813 ), .A4(_AES_ENC_us21_n812 ), .ZN(_AES_ENC_us21_n816 ) );
NOR2_X2 _AES_ENC_us21_U93  ( .A1(_AES_ENC_us21_n591 ), .A2(_AES_ENC_us21_n569 ), .ZN(_AES_ENC_us21_n721 ) );
NOR2_X2 _AES_ENC_us21_U92  ( .A1(_AES_ENC_us21_n1031 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n723 ) );
NOR2_X2 _AES_ENC_us21_U91  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n1096 ), .ZN(_AES_ENC_us21_n722 ) );
NOR4_X2 _AES_ENC_us21_U90  ( .A1(_AES_ENC_us21_n724 ), .A2(_AES_ENC_us21_n723 ), .A3(_AES_ENC_us21_n722 ), .A4(_AES_ENC_us21_n721 ), .ZN(_AES_ENC_us21_n725 ) );
NOR2_X2 _AES_ENC_us21_U89  ( .A1(_AES_ENC_us21_n911 ), .A2(_AES_ENC_us21_n990 ), .ZN(_AES_ENC_us21_n1009 ) );
NOR2_X2 _AES_ENC_us21_U88  ( .A1(_AES_ENC_us21_n1013 ), .A2(_AES_ENC_us21_n573 ), .ZN(_AES_ENC_us21_n1014 ) );
NOR2_X2 _AES_ENC_us21_U87  ( .A1(_AES_ENC_us21_n1014 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n1015 ) );
NOR4_X2 _AES_ENC_us21_U86  ( .A1(_AES_ENC_us21_n1016 ), .A2(_AES_ENC_us21_n1015 ), .A3(_AES_ENC_us21_n1119 ), .A4(_AES_ENC_us21_n1046 ), .ZN(_AES_ENC_us21_n1017 ) );
NOR2_X2 _AES_ENC_us21_U81  ( .A1(_AES_ENC_us21_n996 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n998 ) );
NOR2_X2 _AES_ENC_us21_U80  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n618 ), .ZN(_AES_ENC_us21_n1000 ) );
NOR2_X2 _AES_ENC_us21_U79  ( .A1(_AES_ENC_us21_n590 ), .A2(_AES_ENC_us21_n1096 ), .ZN(_AES_ENC_us21_n999 ) );
NOR4_X2 _AES_ENC_us21_U78  ( .A1(_AES_ENC_us21_n1000 ), .A2(_AES_ENC_us21_n999 ), .A3(_AES_ENC_us21_n998 ), .A4(_AES_ENC_us21_n997 ), .ZN(_AES_ENC_us21_n1001 ) );
NOR2_X2 _AES_ENC_us21_U74  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n1096 ), .ZN(_AES_ENC_us21_n697 ) );
NOR2_X2 _AES_ENC_us21_U73  ( .A1(_AES_ENC_us21_n609 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n958 ) );
NOR2_X2 _AES_ENC_us21_U72  ( .A1(_AES_ENC_us21_n911 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n983 ) );
NOR2_X2 _AES_ENC_us21_U71  ( .A1(_AES_ENC_us21_n1054 ), .A2(_AES_ENC_us21_n1103 ), .ZN(_AES_ENC_us21_n1031 ) );
INV_X4 _AES_ENC_us21_U65  ( .A(_AES_ENC_us21_n1050 ), .ZN(_AES_ENC_us21_n585 ) );
INV_X4 _AES_ENC_us21_U64  ( .A(_AES_ENC_us21_n1072 ), .ZN(_AES_ENC_us21_n577 ) );
INV_X4 _AES_ENC_us21_U63  ( .A(_AES_ENC_us21_n1073 ), .ZN(_AES_ENC_us21_n576 ) );
NOR2_X2 _AES_ENC_us21_U62  ( .A1(_AES_ENC_us21_n603 ), .A2(_AES_ENC_us21_n587 ), .ZN(_AES_ENC_us21_n880 ) );
NOR3_X2 _AES_ENC_us21_U61  ( .A1(_AES_ENC_us21_n826 ), .A2(_AES_ENC_us21_n1121 ), .A3(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n946 ) );
INV_X4 _AES_ENC_us21_U59  ( .A(_AES_ENC_us21_n1010 ), .ZN(_AES_ENC_us21_n581 ) );
NOR3_X2 _AES_ENC_us21_U58  ( .A1(_AES_ENC_us21_n573 ), .A2(_AES_ENC_us21_n1029 ), .A3(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n1119 ) );
INV_X4 _AES_ENC_us21_U57  ( .A(_AES_ENC_us21_n956 ), .ZN(_AES_ENC_us21_n589 ) );
NOR2_X2 _AES_ENC_us21_U50  ( .A1(_AES_ENC_us21_n601 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n1013 ) );
NOR2_X2 _AES_ENC_us21_U49  ( .A1(_AES_ENC_us21_n609 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n910 ) );
NOR2_X2 _AES_ENC_us21_U48  ( .A1(_AES_ENC_us21_n569 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n1091 ) );
NOR2_X2 _AES_ENC_us21_U47  ( .A1(_AES_ENC_us21_n614 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n990 ) );
NOR2_X2 _AES_ENC_us21_U46  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_us21_n1121 ), .ZN(_AES_ENC_us21_n996 ) );
NOR2_X2 _AES_ENC_us21_U45  ( .A1(_AES_ENC_us21_n583 ), .A2(_AES_ENC_us21_n622 ), .ZN(_AES_ENC_us21_n628 ) );
NOR2_X2 _AES_ENC_us21_U44  ( .A1(_AES_ENC_us21_n602 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n866 ) );
NOR2_X2 _AES_ENC_us21_U43  ( .A1(_AES_ENC_us21_n610 ), .A2(_AES_ENC_us21_n583 ), .ZN(_AES_ENC_us21_n1006 ) );
NOR2_X2 _AES_ENC_us21_U42  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n1117 ), .ZN(_AES_ENC_us21_n1118 ) );
NOR2_X2 _AES_ENC_us21_U41  ( .A1(_AES_ENC_us21_n1119 ), .A2(_AES_ENC_us21_n1118 ), .ZN(_AES_ENC_us21_n1127 ) );
NOR2_X2 _AES_ENC_us21_U36  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n616 ), .ZN(_AES_ENC_us21_n629 ) );
NOR2_X2 _AES_ENC_us21_U35  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n906 ), .ZN(_AES_ENC_us21_n909 ) );
NOR2_X2 _AES_ENC_us21_U34  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n607 ), .ZN(_AES_ENC_us21_n658 ) );
NOR2_X2 _AES_ENC_us21_U33  ( .A1(_AES_ENC_us21_n1116 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n695 ) );
NOR2_X2 _AES_ENC_us21_U32  ( .A1(_AES_ENC_us21_n1078 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n1083 ) );
NOR2_X2 _AES_ENC_us21_U31  ( .A1(_AES_ENC_us21_n941 ), .A2(_AES_ENC_us21_n581 ), .ZN(_AES_ENC_us21_n724 ) );
NOR2_X2 _AES_ENC_us21_U30  ( .A1(_AES_ENC_us21_n611 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n1107 ) );
NOR2_X2 _AES_ENC_us21_U29  ( .A1(_AES_ENC_us21_n602 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n840 ) );
NOR2_X2 _AES_ENC_us21_U24  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n623 ), .ZN(_AES_ENC_us21_n633 ) );
NOR2_X2 _AES_ENC_us21_U23  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n1080 ), .ZN(_AES_ENC_us21_n1081 ) );
NOR2_X2 _AES_ENC_us21_U21  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n1045 ), .ZN(_AES_ENC_us21_n812 ) );
NOR2_X2 _AES_ENC_us21_U20  ( .A1(_AES_ENC_us21_n1009 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n960 ) );
NOR2_X2 _AES_ENC_us21_U19  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n619 ), .ZN(_AES_ENC_us21_n982 ) );
NOR2_X2 _AES_ENC_us21_U18  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n616 ), .ZN(_AES_ENC_us21_n757 ) );
NOR2_X2 _AES_ENC_us21_U17  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n598 ), .ZN(_AES_ENC_us21_n698 ) );
NOR2_X2 _AES_ENC_us21_U16  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n605 ), .ZN(_AES_ENC_us21_n708 ) );
NOR2_X2 _AES_ENC_us21_U15  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n603 ), .ZN(_AES_ENC_us21_n770 ) );
NOR2_X2 _AES_ENC_us21_U10  ( .A1(_AES_ENC_us21_n605 ), .A2(_AES_ENC_us21_n576 ), .ZN(_AES_ENC_us21_n803 ) );
NOR2_X2 _AES_ENC_us21_U9  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n881 ), .ZN(_AES_ENC_us21_n711 ) );
NOR2_X2 _AES_ENC_us21_U8  ( .A1(_AES_ENC_us21_n589 ), .A2(_AES_ENC_us21_n603 ), .ZN(_AES_ENC_us21_n867 ) );
NOR2_X2 _AES_ENC_us21_U7  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n615 ), .ZN(_AES_ENC_us21_n804 ) );
NOR2_X2 _AES_ENC_us21_U6  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n609 ), .ZN(_AES_ENC_us21_n1046 ) );
OR2_X4 _AES_ENC_us21_U5  ( .A1(_AES_ENC_us21_n612 ), .A2(_AES_ENC_sa21[1]),.ZN(_AES_ENC_us21_n570 ) );
OR2_X4 _AES_ENC_us21_U4  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_sa21[4]),.ZN(_AES_ENC_us21_n569 ) );
NAND2_X2 _AES_ENC_us21_U514  ( .A1(_AES_ENC_us21_n1121 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n1030 ) );
AND2_X2 _AES_ENC_us21_U513  ( .A1(_AES_ENC_us21_n607 ), .A2(_AES_ENC_us21_n1030 ), .ZN(_AES_ENC_us21_n1049 ) );
NAND2_X2 _AES_ENC_us21_U511  ( .A1(_AES_ENC_us21_n1049 ), .A2(_AES_ENC_us21_n794 ), .ZN(_AES_ENC_us21_n637 ) );
AND2_X2 _AES_ENC_us21_U493  ( .A1(_AES_ENC_us21_n779 ), .A2(_AES_ENC_us21_n996 ), .ZN(_AES_ENC_us21_n632 ) );
NAND4_X2 _AES_ENC_us21_U485  ( .A1(_AES_ENC_us21_n637 ), .A2(_AES_ENC_us21_n636 ), .A3(_AES_ENC_us21_n635 ), .A4(_AES_ENC_us21_n634 ), .ZN(_AES_ENC_us21_n638 ) );
NAND2_X2 _AES_ENC_us21_U484  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n638 ), .ZN(_AES_ENC_us21_n679 ) );
NAND2_X2 _AES_ENC_us21_U481  ( .A1(_AES_ENC_us21_n1094 ), .A2(_AES_ENC_us21_n613 ), .ZN(_AES_ENC_us21_n648 ) );
NAND2_X2 _AES_ENC_us21_U476  ( .A1(_AES_ENC_us21_n619 ), .A2(_AES_ENC_us21_n598 ), .ZN(_AES_ENC_us21_n762 ) );
NAND2_X2 _AES_ENC_us21_U475  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n762 ), .ZN(_AES_ENC_us21_n647 ) );
NAND4_X2 _AES_ENC_us21_U457  ( .A1(_AES_ENC_us21_n648 ), .A2(_AES_ENC_us21_n647 ), .A3(_AES_ENC_us21_n646 ), .A4(_AES_ENC_us21_n645 ), .ZN(_AES_ENC_us21_n649 ) );
NAND2_X2 _AES_ENC_us21_U456  ( .A1(_AES_ENC_sa21[0]), .A2(_AES_ENC_us21_n649 ), .ZN(_AES_ENC_us21_n665 ) );
NAND2_X2 _AES_ENC_us21_U454  ( .A1(_AES_ENC_us21_n626 ), .A2(_AES_ENC_us21_n601 ), .ZN(_AES_ENC_us21_n855 ) );
NAND2_X2 _AES_ENC_us21_U453  ( .A1(_AES_ENC_us21_n617 ), .A2(_AES_ENC_us21_n855 ), .ZN(_AES_ENC_us21_n821 ) );
NAND2_X2 _AES_ENC_us21_U452  ( .A1(_AES_ENC_us21_n1093 ), .A2(_AES_ENC_us21_n821 ), .ZN(_AES_ENC_us21_n662 ) );
NAND2_X2 _AES_ENC_us21_U451  ( .A1(_AES_ENC_us21_n605 ), .A2(_AES_ENC_us21_n620 ), .ZN(_AES_ENC_us21_n650 ) );
NAND2_X2 _AES_ENC_us21_U450  ( .A1(_AES_ENC_us21_n956 ), .A2(_AES_ENC_us21_n650 ), .ZN(_AES_ENC_us21_n661 ) );
NAND2_X2 _AES_ENC_us21_U449  ( .A1(_AES_ENC_us21_n594 ), .A2(_AES_ENC_us21_n595 ), .ZN(_AES_ENC_us21_n839 ) );
OR2_X2 _AES_ENC_us21_U446  ( .A1(_AES_ENC_us21_n839 ), .A2(_AES_ENC_us21_n932 ), .ZN(_AES_ENC_us21_n656 ) );
NAND2_X2 _AES_ENC_us21_U445  ( .A1(_AES_ENC_us21_n624 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n1096 ) );
NAND2_X2 _AES_ENC_us21_U444  ( .A1(_AES_ENC_us21_n1030 ), .A2(_AES_ENC_us21_n1096 ), .ZN(_AES_ENC_us21_n651 ) );
NAND2_X2 _AES_ENC_us21_U443  ( .A1(_AES_ENC_us21_n1114 ), .A2(_AES_ENC_us21_n651 ), .ZN(_AES_ENC_us21_n655 ) );
OR3_X2 _AES_ENC_us21_U440  ( .A1(_AES_ENC_us21_n1079 ), .A2(_AES_ENC_sa21[7]), .A3(_AES_ENC_us21_n594 ), .ZN(_AES_ENC_us21_n654 ));
NAND2_X2 _AES_ENC_us21_U439  ( .A1(_AES_ENC_us21_n623 ), .A2(_AES_ENC_us21_n619 ), .ZN(_AES_ENC_us21_n652 ) );
NAND4_X2 _AES_ENC_us21_U437  ( .A1(_AES_ENC_us21_n656 ), .A2(_AES_ENC_us21_n655 ), .A3(_AES_ENC_us21_n654 ), .A4(_AES_ENC_us21_n653 ), .ZN(_AES_ENC_us21_n657 ) );
NAND2_X2 _AES_ENC_us21_U436  ( .A1(_AES_ENC_sa21[2]), .A2(_AES_ENC_us21_n657 ), .ZN(_AES_ENC_us21_n660 ) );
NAND4_X2 _AES_ENC_us21_U432  ( .A1(_AES_ENC_us21_n662 ), .A2(_AES_ENC_us21_n661 ), .A3(_AES_ENC_us21_n660 ), .A4(_AES_ENC_us21_n659 ), .ZN(_AES_ENC_us21_n663 ) );
NAND2_X2 _AES_ENC_us21_U431  ( .A1(_AES_ENC_us21_n663 ), .A2(_AES_ENC_us21_n627 ), .ZN(_AES_ENC_us21_n664 ) );
NAND2_X2 _AES_ENC_us21_U430  ( .A1(_AES_ENC_us21_n665 ), .A2(_AES_ENC_us21_n664 ), .ZN(_AES_ENC_us21_n666 ) );
NAND2_X2 _AES_ENC_us21_U429  ( .A1(_AES_ENC_sa21[6]), .A2(_AES_ENC_us21_n666 ), .ZN(_AES_ENC_us21_n678 ) );
NAND2_X2 _AES_ENC_us21_U426  ( .A1(_AES_ENC_us21_n735 ), .A2(_AES_ENC_us21_n1093 ), .ZN(_AES_ENC_us21_n675 ) );
NAND2_X2 _AES_ENC_us21_U425  ( .A1(_AES_ENC_us21_n625 ), .A2(_AES_ENC_us21_n607 ), .ZN(_AES_ENC_us21_n1045 ) );
OR2_X2 _AES_ENC_us21_U424  ( .A1(_AES_ENC_us21_n1045 ), .A2(_AES_ENC_us21_n577 ), .ZN(_AES_ENC_us21_n674 ) );
NAND2_X2 _AES_ENC_us21_U423  ( .A1(_AES_ENC_sa21[1]), .A2(_AES_ENC_us21_n609 ), .ZN(_AES_ENC_us21_n667 ) );
NAND2_X2 _AES_ENC_us21_U422  ( .A1(_AES_ENC_us21_n605 ), .A2(_AES_ENC_us21_n667 ), .ZN(_AES_ENC_us21_n1071 ) );
NAND4_X2 _AES_ENC_us21_U412  ( .A1(_AES_ENC_us21_n675 ), .A2(_AES_ENC_us21_n674 ), .A3(_AES_ENC_us21_n673 ), .A4(_AES_ENC_us21_n672 ), .ZN(_AES_ENC_us21_n676 ) );
NAND2_X2 _AES_ENC_us21_U411  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n676 ), .ZN(_AES_ENC_us21_n677 ) );
NAND2_X2 _AES_ENC_us21_U408  ( .A1(_AES_ENC_us21_n800 ), .A2(_AES_ENC_us21_n1022 ), .ZN(_AES_ENC_us21_n680 ) );
NAND2_X2 _AES_ENC_us21_U407  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n680 ), .ZN(_AES_ENC_us21_n681 ) );
AND2_X2 _AES_ENC_us21_U402  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n684 ), .ZN(_AES_ENC_us21_n682 ) );
NAND4_X2 _AES_ENC_us21_U395  ( .A1(_AES_ENC_us21_n691 ), .A2(_AES_ENC_us21_n586 ), .A3(_AES_ENC_us21_n690 ), .A4(_AES_ENC_us21_n689 ), .ZN(_AES_ENC_us21_n692 ) );
NAND2_X2 _AES_ENC_us21_U394  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n692 ), .ZN(_AES_ENC_us21_n733 ) );
NAND2_X2 _AES_ENC_us21_U392  ( .A1(_AES_ENC_us21_n977 ), .A2(_AES_ENC_us21_n1050 ), .ZN(_AES_ENC_us21_n702 ) );
NAND2_X2 _AES_ENC_us21_U391  ( .A1(_AES_ENC_us21_n1093 ), .A2(_AES_ENC_us21_n1045 ), .ZN(_AES_ENC_us21_n701 ) );
NAND4_X2 _AES_ENC_us21_U381  ( .A1(_AES_ENC_us21_n702 ), .A2(_AES_ENC_us21_n701 ), .A3(_AES_ENC_us21_n700 ), .A4(_AES_ENC_us21_n699 ), .ZN(_AES_ENC_us21_n703 ) );
NAND2_X2 _AES_ENC_us21_U380  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n703 ), .ZN(_AES_ENC_us21_n732 ) );
AND2_X2 _AES_ENC_us21_U379  ( .A1(_AES_ENC_sa21[0]), .A2(_AES_ENC_sa21[6]),.ZN(_AES_ENC_us21_n1113 ) );
NAND2_X2 _AES_ENC_us21_U378  ( .A1(_AES_ENC_us21_n619 ), .A2(_AES_ENC_us21_n1030 ), .ZN(_AES_ENC_us21_n881 ) );
NAND2_X2 _AES_ENC_us21_U377  ( .A1(_AES_ENC_us21_n1093 ), .A2(_AES_ENC_us21_n881 ), .ZN(_AES_ENC_us21_n715 ) );
NAND2_X2 _AES_ENC_us21_U376  ( .A1(_AES_ENC_us21_n1010 ), .A2(_AES_ENC_us21_n622 ), .ZN(_AES_ENC_us21_n714 ) );
NAND2_X2 _AES_ENC_us21_U375  ( .A1(_AES_ENC_us21_n855 ), .A2(_AES_ENC_us21_n625 ), .ZN(_AES_ENC_us21_n1117 ) );
XNOR2_X2 _AES_ENC_us21_U371  ( .A(_AES_ENC_us21_n584 ), .B(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n824 ) );
NAND4_X2 _AES_ENC_us21_U362  ( .A1(_AES_ENC_us21_n715 ), .A2(_AES_ENC_us21_n714 ), .A3(_AES_ENC_us21_n713 ), .A4(_AES_ENC_us21_n712 ), .ZN(_AES_ENC_us21_n716 ) );
NAND2_X2 _AES_ENC_us21_U361  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n716 ), .ZN(_AES_ENC_us21_n731 ) );
AND2_X2 _AES_ENC_us21_U360  ( .A1(_AES_ENC_sa21[6]), .A2(_AES_ENC_us21_n627 ), .ZN(_AES_ENC_us21_n1131 ) );
NAND2_X2 _AES_ENC_us21_U359  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n717 ) );
NAND2_X2 _AES_ENC_us21_U358  ( .A1(_AES_ENC_us21_n1029 ), .A2(_AES_ENC_us21_n717 ), .ZN(_AES_ENC_us21_n728 ) );
NAND2_X2 _AES_ENC_us21_U357  ( .A1(_AES_ENC_sa21[1]), .A2(_AES_ENC_us21_n612 ), .ZN(_AES_ENC_us21_n1097 ) );
NAND2_X2 _AES_ENC_us21_U356  ( .A1(_AES_ENC_us21_n610 ), .A2(_AES_ENC_us21_n1097 ), .ZN(_AES_ENC_us21_n718 ) );
NAND2_X2 _AES_ENC_us21_U355  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n718 ), .ZN(_AES_ENC_us21_n727 ) );
NAND4_X2 _AES_ENC_us21_U344  ( .A1(_AES_ENC_us21_n728 ), .A2(_AES_ENC_us21_n727 ), .A3(_AES_ENC_us21_n726 ), .A4(_AES_ENC_us21_n725 ), .ZN(_AES_ENC_us21_n729 ) );
NAND2_X2 _AES_ENC_us21_U343  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n729 ), .ZN(_AES_ENC_us21_n730 ) );
NAND4_X2 _AES_ENC_us21_U342  ( .A1(_AES_ENC_us21_n733 ), .A2(_AES_ENC_us21_n732 ), .A3(_AES_ENC_us21_n731 ), .A4(_AES_ENC_us21_n730 ), .ZN(_AES_ENC_sa21_sub[1] ) );
NAND2_X2 _AES_ENC_us21_U341  ( .A1(_AES_ENC_sa21[7]), .A2(_AES_ENC_us21_n584 ), .ZN(_AES_ENC_us21_n734 ) );
NAND2_X2 _AES_ENC_us21_U340  ( .A1(_AES_ENC_us21_n734 ), .A2(_AES_ENC_us21_n579 ), .ZN(_AES_ENC_us21_n738 ) );
OR4_X2 _AES_ENC_us21_U339  ( .A1(_AES_ENC_us21_n738 ), .A2(_AES_ENC_us21_n594 ), .A3(_AES_ENC_us21_n826 ), .A4(_AES_ENC_us21_n1121 ), .ZN(_AES_ENC_us21_n746 ) );
NAND2_X2 _AES_ENC_us21_U337  ( .A1(_AES_ENC_us21_n1100 ), .A2(_AES_ENC_us21_n617 ), .ZN(_AES_ENC_us21_n992 ) );
OR2_X2 _AES_ENC_us21_U336  ( .A1(_AES_ENC_us21_n583 ), .A2(_AES_ENC_us21_n735 ), .ZN(_AES_ENC_us21_n737 ) );
NAND2_X2 _AES_ENC_us21_U334  ( .A1(_AES_ENC_us21_n605 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n753 ) );
NAND2_X2 _AES_ENC_us21_U333  ( .A1(_AES_ENC_us21_n603 ), .A2(_AES_ENC_us21_n753 ), .ZN(_AES_ENC_us21_n1080 ) );
NAND2_X2 _AES_ENC_us21_U332  ( .A1(_AES_ENC_us21_n1048 ), .A2(_AES_ENC_us21_n602 ), .ZN(_AES_ENC_us21_n736 ) );
NAND2_X2 _AES_ENC_us21_U331  ( .A1(_AES_ENC_us21_n737 ), .A2(_AES_ENC_us21_n736 ), .ZN(_AES_ENC_us21_n739 ) );
NAND2_X2 _AES_ENC_us21_U330  ( .A1(_AES_ENC_us21_n739 ), .A2(_AES_ENC_us21_n738 ), .ZN(_AES_ENC_us21_n745 ) );
NAND2_X2 _AES_ENC_us21_U326  ( .A1(_AES_ENC_us21_n1096 ), .A2(_AES_ENC_us21_n598 ), .ZN(_AES_ENC_us21_n906 ) );
NAND4_X2 _AES_ENC_us21_U323  ( .A1(_AES_ENC_us21_n746 ), .A2(_AES_ENC_us21_n992 ), .A3(_AES_ENC_us21_n745 ), .A4(_AES_ENC_us21_n744 ), .ZN(_AES_ENC_us21_n747 ) );
NAND2_X2 _AES_ENC_us21_U322  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n747 ), .ZN(_AES_ENC_us21_n793 ) );
NAND2_X2 _AES_ENC_us21_U321  ( .A1(_AES_ENC_us21_n606 ), .A2(_AES_ENC_us21_n855 ), .ZN(_AES_ENC_us21_n748 ) );
NAND2_X2 _AES_ENC_us21_U320  ( .A1(_AES_ENC_us21_n956 ), .A2(_AES_ENC_us21_n748 ), .ZN(_AES_ENC_us21_n760 ) );
NAND2_X2 _AES_ENC_us21_U313  ( .A1(_AES_ENC_us21_n598 ), .A2(_AES_ENC_us21_n753 ), .ZN(_AES_ENC_us21_n1023 ) );
NAND4_X2 _AES_ENC_us21_U308  ( .A1(_AES_ENC_us21_n760 ), .A2(_AES_ENC_us21_n992 ), .A3(_AES_ENC_us21_n759 ), .A4(_AES_ENC_us21_n758 ), .ZN(_AES_ENC_us21_n761 ) );
NAND2_X2 _AES_ENC_us21_U307  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n761 ), .ZN(_AES_ENC_us21_n792 ) );
NAND2_X2 _AES_ENC_us21_U306  ( .A1(_AES_ENC_us21_n606 ), .A2(_AES_ENC_us21_n610 ), .ZN(_AES_ENC_us21_n989 ) );
NAND2_X2 _AES_ENC_us21_U305  ( .A1(_AES_ENC_us21_n1050 ), .A2(_AES_ENC_us21_n989 ), .ZN(_AES_ENC_us21_n777 ) );
NAND2_X2 _AES_ENC_us21_U304  ( .A1(_AES_ENC_us21_n1093 ), .A2(_AES_ENC_us21_n762 ), .ZN(_AES_ENC_us21_n776 ) );
XNOR2_X2 _AES_ENC_us21_U301  ( .A(_AES_ENC_sa21[7]), .B(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n959 ) );
NAND4_X2 _AES_ENC_us21_U289  ( .A1(_AES_ENC_us21_n777 ), .A2(_AES_ENC_us21_n776 ), .A3(_AES_ENC_us21_n775 ), .A4(_AES_ENC_us21_n774 ), .ZN(_AES_ENC_us21_n778 ) );
NAND2_X2 _AES_ENC_us21_U288  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n778 ), .ZN(_AES_ENC_us21_n791 ) );
NAND2_X2 _AES_ENC_us21_U287  ( .A1(_AES_ENC_us21_n1056 ), .A2(_AES_ENC_us21_n1050 ), .ZN(_AES_ENC_us21_n788 ) );
NAND2_X2 _AES_ENC_us21_U286  ( .A1(_AES_ENC_us21_n1091 ), .A2(_AES_ENC_us21_n779 ), .ZN(_AES_ENC_us21_n787 ) );
NAND2_X2 _AES_ENC_us21_U285  ( .A1(_AES_ENC_us21_n956 ), .A2(_AES_ENC_sa21[1]), .ZN(_AES_ENC_us21_n786 ) );
NAND4_X2 _AES_ENC_us21_U278  ( .A1(_AES_ENC_us21_n788 ), .A2(_AES_ENC_us21_n787 ), .A3(_AES_ENC_us21_n786 ), .A4(_AES_ENC_us21_n785 ), .ZN(_AES_ENC_us21_n789 ) );
NAND2_X2 _AES_ENC_us21_U277  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n789 ), .ZN(_AES_ENC_us21_n790 ) );
NAND4_X2 _AES_ENC_us21_U276  ( .A1(_AES_ENC_us21_n793 ), .A2(_AES_ENC_us21_n792 ), .A3(_AES_ENC_us21_n791 ), .A4(_AES_ENC_us21_n790 ), .ZN(_AES_ENC_sa21_sub[2] ) );
NAND2_X2 _AES_ENC_us21_U275  ( .A1(_AES_ENC_us21_n1059 ), .A2(_AES_ENC_us21_n794 ), .ZN(_AES_ENC_us21_n810 ) );
NAND2_X2 _AES_ENC_us21_U274  ( .A1(_AES_ENC_us21_n1049 ), .A2(_AES_ENC_us21_n956 ), .ZN(_AES_ENC_us21_n809 ) );
OR2_X2 _AES_ENC_us21_U266  ( .A1(_AES_ENC_us21_n1096 ), .A2(_AES_ENC_us21_n578 ), .ZN(_AES_ENC_us21_n802 ) );
NAND2_X2 _AES_ENC_us21_U265  ( .A1(_AES_ENC_us21_n1053 ), .A2(_AES_ENC_us21_n800 ), .ZN(_AES_ENC_us21_n801 ) );
NAND2_X2 _AES_ENC_us21_U264  ( .A1(_AES_ENC_us21_n802 ), .A2(_AES_ENC_us21_n801 ), .ZN(_AES_ENC_us21_n805 ) );
NAND4_X2 _AES_ENC_us21_U261  ( .A1(_AES_ENC_us21_n810 ), .A2(_AES_ENC_us21_n809 ), .A3(_AES_ENC_us21_n808 ), .A4(_AES_ENC_us21_n807 ), .ZN(_AES_ENC_us21_n811 ) );
NAND2_X2 _AES_ENC_us21_U260  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n811 ), .ZN(_AES_ENC_us21_n852 ) );
OR2_X2 _AES_ENC_us21_U259  ( .A1(_AES_ENC_us21_n1023 ), .A2(_AES_ENC_us21_n591 ), .ZN(_AES_ENC_us21_n819 ) );
OR2_X2 _AES_ENC_us21_U257  ( .A1(_AES_ENC_us21_n570 ), .A2(_AES_ENC_us21_n930 ), .ZN(_AES_ENC_us21_n818 ) );
NAND2_X2 _AES_ENC_us21_U256  ( .A1(_AES_ENC_us21_n1013 ), .A2(_AES_ENC_us21_n1094 ), .ZN(_AES_ENC_us21_n817 ) );
NAND4_X2 _AES_ENC_us21_U249  ( .A1(_AES_ENC_us21_n819 ), .A2(_AES_ENC_us21_n818 ), .A3(_AES_ENC_us21_n817 ), .A4(_AES_ENC_us21_n816 ), .ZN(_AES_ENC_us21_n820 ) );
NAND2_X2 _AES_ENC_us21_U248  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n820 ), .ZN(_AES_ENC_us21_n851 ) );
NAND2_X2 _AES_ENC_us21_U247  ( .A1(_AES_ENC_us21_n956 ), .A2(_AES_ENC_us21_n1080 ), .ZN(_AES_ENC_us21_n835 ) );
NAND2_X2 _AES_ENC_us21_U246  ( .A1(_AES_ENC_us21_n570 ), .A2(_AES_ENC_us21_n1030 ), .ZN(_AES_ENC_us21_n1047 ) );
OR2_X2 _AES_ENC_us21_U245  ( .A1(_AES_ENC_us21_n1047 ), .A2(_AES_ENC_us21_n585 ), .ZN(_AES_ENC_us21_n834 ) );
NAND2_X2 _AES_ENC_us21_U244  ( .A1(_AES_ENC_us21_n1072 ), .A2(_AES_ENC_us21_n620 ), .ZN(_AES_ENC_us21_n833 ) );
NAND4_X2 _AES_ENC_us21_U233  ( .A1(_AES_ENC_us21_n835 ), .A2(_AES_ENC_us21_n834 ), .A3(_AES_ENC_us21_n833 ), .A4(_AES_ENC_us21_n832 ), .ZN(_AES_ENC_us21_n836 ) );
NAND2_X2 _AES_ENC_us21_U232  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n836 ), .ZN(_AES_ENC_us21_n850 ) );
NAND2_X2 _AES_ENC_us21_U231  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n601 ), .ZN(_AES_ENC_us21_n847 ) );
NAND2_X2 _AES_ENC_us21_U230  ( .A1(_AES_ENC_us21_n1050 ), .A2(_AES_ENC_us21_n1071 ), .ZN(_AES_ENC_us21_n846 ) );
OR2_X2 _AES_ENC_us21_U224  ( .A1(_AES_ENC_us21_n1053 ), .A2(_AES_ENC_us21_n911 ), .ZN(_AES_ENC_us21_n1077 ) );
NAND4_X2 _AES_ENC_us21_U220  ( .A1(_AES_ENC_us21_n847 ), .A2(_AES_ENC_us21_n846 ), .A3(_AES_ENC_us21_n845 ), .A4(_AES_ENC_us21_n844 ), .ZN(_AES_ENC_us21_n848 ) );
NAND2_X2 _AES_ENC_us21_U219  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n848 ), .ZN(_AES_ENC_us21_n849 ) );
NAND4_X2 _AES_ENC_us21_U218  ( .A1(_AES_ENC_us21_n852 ), .A2(_AES_ENC_us21_n851 ), .A3(_AES_ENC_us21_n850 ), .A4(_AES_ENC_us21_n849 ), .ZN(_AES_ENC_sa21_sub[3] ) );
NAND2_X2 _AES_ENC_us21_U216  ( .A1(_AES_ENC_us21_n1009 ), .A2(_AES_ENC_us21_n1072 ), .ZN(_AES_ENC_us21_n862 ) );
NAND2_X2 _AES_ENC_us21_U215  ( .A1(_AES_ENC_us21_n610 ), .A2(_AES_ENC_us21_n618 ), .ZN(_AES_ENC_us21_n853 ) );
NAND2_X2 _AES_ENC_us21_U214  ( .A1(_AES_ENC_us21_n1050 ), .A2(_AES_ENC_us21_n853 ), .ZN(_AES_ENC_us21_n861 ) );
NAND4_X2 _AES_ENC_us21_U206  ( .A1(_AES_ENC_us21_n862 ), .A2(_AES_ENC_us21_n861 ), .A3(_AES_ENC_us21_n860 ), .A4(_AES_ENC_us21_n859 ), .ZN(_AES_ENC_us21_n863 ) );
NAND2_X2 _AES_ENC_us21_U205  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n863 ), .ZN(_AES_ENC_us21_n905 ) );
NAND2_X2 _AES_ENC_us21_U204  ( .A1(_AES_ENC_us21_n1010 ), .A2(_AES_ENC_us21_n989 ), .ZN(_AES_ENC_us21_n874 ) );
NAND2_X2 _AES_ENC_us21_U203  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n583 ), .ZN(_AES_ENC_us21_n864 ) );
NAND2_X2 _AES_ENC_us21_U202  ( .A1(_AES_ENC_us21_n929 ), .A2(_AES_ENC_us21_n864 ), .ZN(_AES_ENC_us21_n873 ) );
NAND4_X2 _AES_ENC_us21_U193  ( .A1(_AES_ENC_us21_n874 ), .A2(_AES_ENC_us21_n873 ), .A3(_AES_ENC_us21_n872 ), .A4(_AES_ENC_us21_n871 ), .ZN(_AES_ENC_us21_n875 ) );
NAND2_X2 _AES_ENC_us21_U192  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n875 ), .ZN(_AES_ENC_us21_n904 ) );
NAND2_X2 _AES_ENC_us21_U191  ( .A1(_AES_ENC_us21_n597 ), .A2(_AES_ENC_us21_n1050 ), .ZN(_AES_ENC_us21_n889 ) );
NAND2_X2 _AES_ENC_us21_U190  ( .A1(_AES_ENC_us21_n1093 ), .A2(_AES_ENC_us21_n617 ), .ZN(_AES_ENC_us21_n876 ) );
NAND2_X2 _AES_ENC_us21_U189  ( .A1(_AES_ENC_us21_n576 ), .A2(_AES_ENC_us21_n876 ), .ZN(_AES_ENC_us21_n877 ) );
NAND2_X2 _AES_ENC_us21_U188  ( .A1(_AES_ENC_us21_n877 ), .A2(_AES_ENC_us21_n601 ), .ZN(_AES_ENC_us21_n888 ) );
NAND4_X2 _AES_ENC_us21_U179  ( .A1(_AES_ENC_us21_n889 ), .A2(_AES_ENC_us21_n888 ), .A3(_AES_ENC_us21_n887 ), .A4(_AES_ENC_us21_n886 ), .ZN(_AES_ENC_us21_n890 ) );
NAND2_X2 _AES_ENC_us21_U178  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n890 ), .ZN(_AES_ENC_us21_n903 ) );
OR2_X2 _AES_ENC_us21_U177  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n1059 ), .ZN(_AES_ENC_us21_n900 ) );
NAND2_X2 _AES_ENC_us21_U176  ( .A1(_AES_ENC_us21_n1073 ), .A2(_AES_ENC_us21_n1047 ), .ZN(_AES_ENC_us21_n899 ) );
NAND2_X2 _AES_ENC_us21_U175  ( .A1(_AES_ENC_us21_n1094 ), .A2(_AES_ENC_us21_n608 ), .ZN(_AES_ENC_us21_n898 ) );
NAND4_X2 _AES_ENC_us21_U167  ( .A1(_AES_ENC_us21_n900 ), .A2(_AES_ENC_us21_n899 ), .A3(_AES_ENC_us21_n898 ), .A4(_AES_ENC_us21_n897 ), .ZN(_AES_ENC_us21_n901 ) );
NAND2_X2 _AES_ENC_us21_U166  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n901 ), .ZN(_AES_ENC_us21_n902 ) );
NAND4_X2 _AES_ENC_us21_U165  ( .A1(_AES_ENC_us21_n905 ), .A2(_AES_ENC_us21_n904 ), .A3(_AES_ENC_us21_n903 ), .A4(_AES_ENC_us21_n902 ), .ZN(_AES_ENC_sa21_sub[4] ) );
NAND2_X2 _AES_ENC_us21_U164  ( .A1(_AES_ENC_us21_n1094 ), .A2(_AES_ENC_us21_n615 ), .ZN(_AES_ENC_us21_n922 ) );
NAND2_X2 _AES_ENC_us21_U163  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n989 ), .ZN(_AES_ENC_us21_n921 ) );
NAND4_X2 _AES_ENC_us21_U151  ( .A1(_AES_ENC_us21_n922 ), .A2(_AES_ENC_us21_n921 ), .A3(_AES_ENC_us21_n920 ), .A4(_AES_ENC_us21_n919 ), .ZN(_AES_ENC_us21_n923 ) );
NAND2_X2 _AES_ENC_us21_U150  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n923 ), .ZN(_AES_ENC_us21_n972 ) );
NAND2_X2 _AES_ENC_us21_U149  ( .A1(_AES_ENC_us21_n603 ), .A2(_AES_ENC_us21_n605 ), .ZN(_AES_ENC_us21_n924 ) );
NAND2_X2 _AES_ENC_us21_U148  ( .A1(_AES_ENC_us21_n1073 ), .A2(_AES_ENC_us21_n924 ), .ZN(_AES_ENC_us21_n939 ) );
NAND2_X2 _AES_ENC_us21_U147  ( .A1(_AES_ENC_us21_n926 ), .A2(_AES_ENC_us21_n925 ), .ZN(_AES_ENC_us21_n927 ) );
NAND2_X2 _AES_ENC_us21_U146  ( .A1(_AES_ENC_us21_n578 ), .A2(_AES_ENC_us21_n927 ), .ZN(_AES_ENC_us21_n928 ) );
NAND2_X2 _AES_ENC_us21_U145  ( .A1(_AES_ENC_us21_n928 ), .A2(_AES_ENC_us21_n1080 ), .ZN(_AES_ENC_us21_n938 ) );
OR2_X2 _AES_ENC_us21_U144  ( .A1(_AES_ENC_us21_n1117 ), .A2(_AES_ENC_us21_n589 ), .ZN(_AES_ENC_us21_n937 ) );
NAND4_X2 _AES_ENC_us21_U139  ( .A1(_AES_ENC_us21_n939 ), .A2(_AES_ENC_us21_n938 ), .A3(_AES_ENC_us21_n937 ), .A4(_AES_ENC_us21_n936 ), .ZN(_AES_ENC_us21_n940 ) );
NAND2_X2 _AES_ENC_us21_U138  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n940 ), .ZN(_AES_ENC_us21_n971 ) );
OR2_X2 _AES_ENC_us21_U137  ( .A1(_AES_ENC_us21_n577 ), .A2(_AES_ENC_us21_n941 ), .ZN(_AES_ENC_us21_n954 ) );
NAND2_X2 _AES_ENC_us21_U136  ( .A1(_AES_ENC_us21_n1096 ), .A2(_AES_ENC_us21_n618 ), .ZN(_AES_ENC_us21_n942 ) );
NAND2_X2 _AES_ENC_us21_U135  ( .A1(_AES_ENC_us21_n1048 ), .A2(_AES_ENC_us21_n942 ), .ZN(_AES_ENC_us21_n943 ) );
NAND2_X2 _AES_ENC_us21_U134  ( .A1(_AES_ENC_us21_n585 ), .A2(_AES_ENC_us21_n943 ), .ZN(_AES_ENC_us21_n944 ) );
NAND2_X2 _AES_ENC_us21_U133  ( .A1(_AES_ENC_us21_n944 ), .A2(_AES_ENC_us21_n599 ), .ZN(_AES_ENC_us21_n953 ) );
NAND4_X2 _AES_ENC_us21_U125  ( .A1(_AES_ENC_us21_n954 ), .A2(_AES_ENC_us21_n953 ), .A3(_AES_ENC_us21_n952 ), .A4(_AES_ENC_us21_n951 ), .ZN(_AES_ENC_us21_n955 ) );
NAND2_X2 _AES_ENC_us21_U124  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n955 ), .ZN(_AES_ENC_us21_n970 ) );
NAND2_X2 _AES_ENC_us21_U123  ( .A1(_AES_ENC_us21_n1094 ), .A2(_AES_ENC_us21_n1071 ), .ZN(_AES_ENC_us21_n967 ) );
NAND2_X2 _AES_ENC_us21_U122  ( .A1(_AES_ENC_us21_n956 ), .A2(_AES_ENC_us21_n1030 ), .ZN(_AES_ENC_us21_n966 ) );
NAND4_X2 _AES_ENC_us21_U114  ( .A1(_AES_ENC_us21_n967 ), .A2(_AES_ENC_us21_n966 ), .A3(_AES_ENC_us21_n965 ), .A4(_AES_ENC_us21_n964 ), .ZN(_AES_ENC_us21_n968 ) );
NAND2_X2 _AES_ENC_us21_U113  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n968 ), .ZN(_AES_ENC_us21_n969 ) );
NAND4_X2 _AES_ENC_us21_U112  ( .A1(_AES_ENC_us21_n972 ), .A2(_AES_ENC_us21_n971 ), .A3(_AES_ENC_us21_n970 ), .A4(_AES_ENC_us21_n969 ), .ZN(_AES_ENC_sa21_sub[5] ) );
NAND2_X2 _AES_ENC_us21_U111  ( .A1(_AES_ENC_us21_n570 ), .A2(_AES_ENC_us21_n1097 ), .ZN(_AES_ENC_us21_n973 ) );
NAND2_X2 _AES_ENC_us21_U110  ( .A1(_AES_ENC_us21_n1073 ), .A2(_AES_ENC_us21_n973 ), .ZN(_AES_ENC_us21_n987 ) );
NAND2_X2 _AES_ENC_us21_U109  ( .A1(_AES_ENC_us21_n974 ), .A2(_AES_ENC_us21_n1077 ), .ZN(_AES_ENC_us21_n975 ) );
NAND2_X2 _AES_ENC_us21_U108  ( .A1(_AES_ENC_us21_n587 ), .A2(_AES_ENC_us21_n975 ), .ZN(_AES_ENC_us21_n976 ) );
NAND2_X2 _AES_ENC_us21_U107  ( .A1(_AES_ENC_us21_n977 ), .A2(_AES_ENC_us21_n976 ), .ZN(_AES_ENC_us21_n986 ) );
NAND4_X2 _AES_ENC_us21_U99  ( .A1(_AES_ENC_us21_n987 ), .A2(_AES_ENC_us21_n986 ), .A3(_AES_ENC_us21_n985 ), .A4(_AES_ENC_us21_n984 ), .ZN(_AES_ENC_us21_n988 ) );
NAND2_X2 _AES_ENC_us21_U98  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n988 ), .ZN(_AES_ENC_us21_n1044 ) );
NAND2_X2 _AES_ENC_us21_U97  ( .A1(_AES_ENC_us21_n1073 ), .A2(_AES_ENC_us21_n989 ), .ZN(_AES_ENC_us21_n1004 ) );
NAND2_X2 _AES_ENC_us21_U96  ( .A1(_AES_ENC_us21_n1092 ), .A2(_AES_ENC_us21_n605 ), .ZN(_AES_ENC_us21_n1003 ) );
NAND4_X2 _AES_ENC_us21_U85  ( .A1(_AES_ENC_us21_n1004 ), .A2(_AES_ENC_us21_n1003 ), .A3(_AES_ENC_us21_n1002 ), .A4(_AES_ENC_us21_n1001 ), .ZN(_AES_ENC_us21_n1005 ) );
NAND2_X2 _AES_ENC_us21_U84  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n1005 ), .ZN(_AES_ENC_us21_n1043 ) );
NAND2_X2 _AES_ENC_us21_U83  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n626 ), .ZN(_AES_ENC_us21_n1020 ) );
NAND2_X2 _AES_ENC_us21_U82  ( .A1(_AES_ENC_us21_n1050 ), .A2(_AES_ENC_us21_n612 ), .ZN(_AES_ENC_us21_n1019 ) );
NAND2_X2 _AES_ENC_us21_U77  ( .A1(_AES_ENC_us21_n1059 ), .A2(_AES_ENC_us21_n1114 ), .ZN(_AES_ENC_us21_n1012 ) );
NAND2_X2 _AES_ENC_us21_U76  ( .A1(_AES_ENC_us21_n1010 ), .A2(_AES_ENC_us21_n604 ), .ZN(_AES_ENC_us21_n1011 ) );
NAND2_X2 _AES_ENC_us21_U75  ( .A1(_AES_ENC_us21_n1012 ), .A2(_AES_ENC_us21_n1011 ), .ZN(_AES_ENC_us21_n1016 ) );
NAND4_X2 _AES_ENC_us21_U70  ( .A1(_AES_ENC_us21_n1020 ), .A2(_AES_ENC_us21_n1019 ), .A3(_AES_ENC_us21_n1018 ), .A4(_AES_ENC_us21_n1017 ), .ZN(_AES_ENC_us21_n1021 ) );
NAND2_X2 _AES_ENC_us21_U69  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n1021 ), .ZN(_AES_ENC_us21_n1042 ) );
NAND2_X2 _AES_ENC_us21_U68  ( .A1(_AES_ENC_us21_n1022 ), .A2(_AES_ENC_us21_n1093 ), .ZN(_AES_ENC_us21_n1039 ) );
NAND2_X2 _AES_ENC_us21_U67  ( .A1(_AES_ENC_us21_n1050 ), .A2(_AES_ENC_us21_n1023 ), .ZN(_AES_ENC_us21_n1038 ) );
NAND2_X2 _AES_ENC_us21_U66  ( .A1(_AES_ENC_us21_n1024 ), .A2(_AES_ENC_us21_n1071 ), .ZN(_AES_ENC_us21_n1037 ) );
AND2_X2 _AES_ENC_us21_U60  ( .A1(_AES_ENC_us21_n1030 ), .A2(_AES_ENC_us21_n621 ), .ZN(_AES_ENC_us21_n1078 ) );
NAND4_X2 _AES_ENC_us21_U56  ( .A1(_AES_ENC_us21_n1039 ), .A2(_AES_ENC_us21_n1038 ), .A3(_AES_ENC_us21_n1037 ), .A4(_AES_ENC_us21_n1036 ), .ZN(_AES_ENC_us21_n1040 ) );
NAND2_X2 _AES_ENC_us21_U55  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n1040 ), .ZN(_AES_ENC_us21_n1041 ) );
NAND4_X2 _AES_ENC_us21_U54  ( .A1(_AES_ENC_us21_n1044 ), .A2(_AES_ENC_us21_n1043 ), .A3(_AES_ENC_us21_n1042 ), .A4(_AES_ENC_us21_n1041 ), .ZN(_AES_ENC_sa21_sub[6] ) );
NAND2_X2 _AES_ENC_us21_U53  ( .A1(_AES_ENC_us21_n1072 ), .A2(_AES_ENC_us21_n1045 ), .ZN(_AES_ENC_us21_n1068 ) );
NAND2_X2 _AES_ENC_us21_U52  ( .A1(_AES_ENC_us21_n1046 ), .A2(_AES_ENC_us21_n603 ), .ZN(_AES_ENC_us21_n1067 ) );
NAND2_X2 _AES_ENC_us21_U51  ( .A1(_AES_ENC_us21_n1094 ), .A2(_AES_ENC_us21_n1047 ), .ZN(_AES_ENC_us21_n1066 ) );
NAND4_X2 _AES_ENC_us21_U40  ( .A1(_AES_ENC_us21_n1068 ), .A2(_AES_ENC_us21_n1067 ), .A3(_AES_ENC_us21_n1066 ), .A4(_AES_ENC_us21_n1065 ), .ZN(_AES_ENC_us21_n1069 ) );
NAND2_X2 _AES_ENC_us21_U39  ( .A1(_AES_ENC_us21_n1070 ), .A2(_AES_ENC_us21_n1069 ), .ZN(_AES_ENC_us21_n1135 ) );
NAND2_X2 _AES_ENC_us21_U38  ( .A1(_AES_ENC_us21_n1072 ), .A2(_AES_ENC_us21_n1071 ), .ZN(_AES_ENC_us21_n1088 ) );
NAND2_X2 _AES_ENC_us21_U37  ( .A1(_AES_ENC_us21_n1073 ), .A2(_AES_ENC_us21_n608 ), .ZN(_AES_ENC_us21_n1087 ) );
NAND4_X2 _AES_ENC_us21_U28  ( .A1(_AES_ENC_us21_n1088 ), .A2(_AES_ENC_us21_n1087 ), .A3(_AES_ENC_us21_n1086 ), .A4(_AES_ENC_us21_n1085 ), .ZN(_AES_ENC_us21_n1089 ) );
NAND2_X2 _AES_ENC_us21_U27  ( .A1(_AES_ENC_us21_n1090 ), .A2(_AES_ENC_us21_n1089 ), .ZN(_AES_ENC_us21_n1134 ) );
NAND2_X2 _AES_ENC_us21_U26  ( .A1(_AES_ENC_us21_n1091 ), .A2(_AES_ENC_us21_n1093 ), .ZN(_AES_ENC_us21_n1111 ) );
NAND2_X2 _AES_ENC_us21_U25  ( .A1(_AES_ENC_us21_n1092 ), .A2(_AES_ENC_us21_n1120 ), .ZN(_AES_ENC_us21_n1110 ) );
AND2_X2 _AES_ENC_us21_U22  ( .A1(_AES_ENC_us21_n1097 ), .A2(_AES_ENC_us21_n1096 ), .ZN(_AES_ENC_us21_n1098 ) );
NAND4_X2 _AES_ENC_us21_U14  ( .A1(_AES_ENC_us21_n1111 ), .A2(_AES_ENC_us21_n1110 ), .A3(_AES_ENC_us21_n1109 ), .A4(_AES_ENC_us21_n1108 ), .ZN(_AES_ENC_us21_n1112 ) );
NAND2_X2 _AES_ENC_us21_U13  ( .A1(_AES_ENC_us21_n1113 ), .A2(_AES_ENC_us21_n1112 ), .ZN(_AES_ENC_us21_n1133 ) );
NAND2_X2 _AES_ENC_us21_U12  ( .A1(_AES_ENC_us21_n1115 ), .A2(_AES_ENC_us21_n1114 ), .ZN(_AES_ENC_us21_n1129 ) );
OR2_X2 _AES_ENC_us21_U11  ( .A1(_AES_ENC_us21_n581 ), .A2(_AES_ENC_us21_n1116 ), .ZN(_AES_ENC_us21_n1128 ) );
NAND4_X2 _AES_ENC_us21_U3  ( .A1(_AES_ENC_us21_n1129 ), .A2(_AES_ENC_us21_n1128 ), .A3(_AES_ENC_us21_n1127 ), .A4(_AES_ENC_us21_n1126 ), .ZN(_AES_ENC_us21_n1130 ) );
NAND2_X2 _AES_ENC_us21_U2  ( .A1(_AES_ENC_us21_n1131 ), .A2(_AES_ENC_us21_n1130 ), .ZN(_AES_ENC_us21_n1132 ) );
NAND4_X2 _AES_ENC_us21_U1  ( .A1(_AES_ENC_us21_n1135 ), .A2(_AES_ENC_us21_n1134 ), .A3(_AES_ENC_us21_n1133 ), .A4(_AES_ENC_us21_n1132 ), .ZN(_AES_ENC_sa21_sub[7] ) );
INV_X4 _AES_ENC_us22_U575  ( .A(_AES_ENC_sa22[7]), .ZN(_AES_ENC_us22_n627 ));
INV_X4 _AES_ENC_us22_U574  ( .A(_AES_ENC_us22_n1114 ), .ZN(_AES_ENC_us22_n625 ) );
INV_X4 _AES_ENC_us22_U573  ( .A(_AES_ENC_sa22[4]), .ZN(_AES_ENC_us22_n624 ));
INV_X4 _AES_ENC_us22_U572  ( .A(_AES_ENC_us22_n1025 ), .ZN(_AES_ENC_us22_n622 ) );
INV_X4 _AES_ENC_us22_U571  ( .A(_AES_ENC_us22_n1120 ), .ZN(_AES_ENC_us22_n620 ) );
INV_X4 _AES_ENC_us22_U570  ( .A(_AES_ENC_us22_n1121 ), .ZN(_AES_ENC_us22_n619 ) );
INV_X4 _AES_ENC_us22_U569  ( .A(_AES_ENC_us22_n1048 ), .ZN(_AES_ENC_us22_n618 ) );
INV_X4 _AES_ENC_us22_U568  ( .A(_AES_ENC_us22_n974 ), .ZN(_AES_ENC_us22_n616 ) );
INV_X4 _AES_ENC_us22_U567  ( .A(_AES_ENC_us22_n794 ), .ZN(_AES_ENC_us22_n614 ) );
INV_X4 _AES_ENC_us22_U566  ( .A(_AES_ENC_sa22[2]), .ZN(_AES_ENC_us22_n611 ));
INV_X4 _AES_ENC_us22_U565  ( .A(_AES_ENC_us22_n800 ), .ZN(_AES_ENC_us22_n610 ) );
INV_X4 _AES_ENC_us22_U564  ( .A(_AES_ENC_us22_n925 ), .ZN(_AES_ENC_us22_n609 ) );
INV_X4 _AES_ENC_us22_U563  ( .A(_AES_ENC_us22_n779 ), .ZN(_AES_ENC_us22_n607 ) );
INV_X4 _AES_ENC_us22_U562  ( .A(_AES_ENC_us22_n1022 ), .ZN(_AES_ENC_us22_n603 ) );
INV_X4 _AES_ENC_us22_U561  ( .A(_AES_ENC_us22_n1102 ), .ZN(_AES_ENC_us22_n602 ) );
INV_X4 _AES_ENC_us22_U560  ( .A(_AES_ENC_us22_n929 ), .ZN(_AES_ENC_us22_n601 ) );
INV_X4 _AES_ENC_us22_U559  ( .A(_AES_ENC_us22_n1056 ), .ZN(_AES_ENC_us22_n600 ) );
INV_X4 _AES_ENC_us22_U558  ( .A(_AES_ENC_us22_n1054 ), .ZN(_AES_ENC_us22_n599 ) );
INV_X4 _AES_ENC_us22_U557  ( .A(_AES_ENC_us22_n881 ), .ZN(_AES_ENC_us22_n598 ) );
INV_X4 _AES_ENC_us22_U556  ( .A(_AES_ENC_us22_n926 ), .ZN(_AES_ENC_us22_n597 ) );
INV_X4 _AES_ENC_us22_U555  ( .A(_AES_ENC_us22_n977 ), .ZN(_AES_ENC_us22_n595 ) );
INV_X4 _AES_ENC_us22_U554  ( .A(_AES_ENC_us22_n1031 ), .ZN(_AES_ENC_us22_n594 ) );
INV_X4 _AES_ENC_us22_U553  ( .A(_AES_ENC_us22_n1103 ), .ZN(_AES_ENC_us22_n593 ) );
INV_X4 _AES_ENC_us22_U552  ( .A(_AES_ENC_us22_n1009 ), .ZN(_AES_ENC_us22_n592 ) );
INV_X4 _AES_ENC_us22_U551  ( .A(_AES_ENC_us22_n990 ), .ZN(_AES_ENC_us22_n591 ) );
INV_X4 _AES_ENC_us22_U550  ( .A(_AES_ENC_us22_n1058 ), .ZN(_AES_ENC_us22_n590 ) );
INV_X4 _AES_ENC_us22_U549  ( .A(_AES_ENC_us22_n1074 ), .ZN(_AES_ENC_us22_n589 ) );
INV_X4 _AES_ENC_us22_U548  ( .A(_AES_ENC_us22_n1053 ), .ZN(_AES_ENC_us22_n588 ) );
INV_X4 _AES_ENC_us22_U547  ( .A(_AES_ENC_us22_n826 ), .ZN(_AES_ENC_us22_n587 ) );
INV_X4 _AES_ENC_us22_U546  ( .A(_AES_ENC_us22_n992 ), .ZN(_AES_ENC_us22_n586 ) );
INV_X4 _AES_ENC_us22_U545  ( .A(_AES_ENC_us22_n821 ), .ZN(_AES_ENC_us22_n585 ) );
INV_X4 _AES_ENC_us22_U544  ( .A(_AES_ENC_us22_n910 ), .ZN(_AES_ENC_us22_n584 ) );
INV_X4 _AES_ENC_us22_U543  ( .A(_AES_ENC_us22_n906 ), .ZN(_AES_ENC_us22_n583 ) );
INV_X4 _AES_ENC_us22_U542  ( .A(_AES_ENC_us22_n880 ), .ZN(_AES_ENC_us22_n581 ) );
INV_X4 _AES_ENC_us22_U541  ( .A(_AES_ENC_us22_n1013 ), .ZN(_AES_ENC_us22_n580 ) );
INV_X4 _AES_ENC_us22_U540  ( .A(_AES_ENC_us22_n1092 ), .ZN(_AES_ENC_us22_n579 ) );
INV_X4 _AES_ENC_us22_U539  ( .A(_AES_ENC_us22_n824 ), .ZN(_AES_ENC_us22_n578 ) );
INV_X4 _AES_ENC_us22_U538  ( .A(_AES_ENC_us22_n1091 ), .ZN(_AES_ENC_us22_n577 ) );
INV_X4 _AES_ENC_us22_U537  ( .A(_AES_ENC_us22_n1080 ), .ZN(_AES_ENC_us22_n576 ) );
INV_X4 _AES_ENC_us22_U536  ( .A(_AES_ENC_us22_n959 ), .ZN(_AES_ENC_us22_n575 ) );
INV_X4 _AES_ENC_us22_U535  ( .A(_AES_ENC_sa22[0]), .ZN(_AES_ENC_us22_n574 ));
NOR2_X2 _AES_ENC_us22_U534  ( .A1(_AES_ENC_sa22[0]), .A2(_AES_ENC_sa22[6]),.ZN(_AES_ENC_us22_n1090 ) );
NOR2_X2 _AES_ENC_us22_U533  ( .A1(_AES_ENC_us22_n574 ), .A2(_AES_ENC_sa22[6]), .ZN(_AES_ENC_us22_n1070 ) );
NOR2_X2 _AES_ENC_us22_U532  ( .A1(_AES_ENC_sa22[4]), .A2(_AES_ENC_sa22[3]),.ZN(_AES_ENC_us22_n1025 ) );
INV_X4 _AES_ENC_us22_U531  ( .A(_AES_ENC_us22_n569 ), .ZN(_AES_ENC_us22_n572 ) );
NOR2_X2 _AES_ENC_us22_U530  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n765 ) );
NOR2_X2 _AES_ENC_us22_U529  ( .A1(_AES_ENC_sa22[4]), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n764 ) );
NOR2_X2 _AES_ENC_us22_U528  ( .A1(_AES_ENC_us22_n765 ), .A2(_AES_ENC_us22_n764 ), .ZN(_AES_ENC_us22_n766 ) );
NOR2_X2 _AES_ENC_us22_U527  ( .A1(_AES_ENC_us22_n766 ), .A2(_AES_ENC_us22_n575 ), .ZN(_AES_ENC_us22_n767 ) );
INV_X4 _AES_ENC_us22_U526  ( .A(_AES_ENC_sa22[3]), .ZN(_AES_ENC_us22_n621 ));
NAND3_X2 _AES_ENC_us22_U525  ( .A1(_AES_ENC_us22_n652 ), .A2(_AES_ENC_us22_n626 ), .A3(_AES_ENC_sa22[7]), .ZN(_AES_ENC_us22_n653 ));
NOR2_X2 _AES_ENC_us22_U524  ( .A1(_AES_ENC_us22_n611 ), .A2(_AES_ENC_sa22[5]), .ZN(_AES_ENC_us22_n925 ) );
NOR2_X2 _AES_ENC_us22_U523  ( .A1(_AES_ENC_sa22[5]), .A2(_AES_ENC_sa22[2]),.ZN(_AES_ENC_us22_n974 ) );
INV_X4 _AES_ENC_us22_U522  ( .A(_AES_ENC_sa22[5]), .ZN(_AES_ENC_us22_n626 ));
NOR2_X2 _AES_ENC_us22_U521  ( .A1(_AES_ENC_us22_n611 ), .A2(_AES_ENC_sa22[7]), .ZN(_AES_ENC_us22_n779 ) );
NAND3_X2 _AES_ENC_us22_U520  ( .A1(_AES_ENC_us22_n679 ), .A2(_AES_ENC_us22_n678 ), .A3(_AES_ENC_us22_n677 ), .ZN(_AES_ENC_sa22_sub[0] ) );
NOR2_X2 _AES_ENC_us22_U519  ( .A1(_AES_ENC_us22_n626 ), .A2(_AES_ENC_sa22[2]), .ZN(_AES_ENC_us22_n1048 ) );
NOR3_X2 _AES_ENC_us22_U518  ( .A1(_AES_ENC_us22_n627 ), .A2(_AES_ENC_sa22[5]), .A3(_AES_ENC_us22_n704 ), .ZN(_AES_ENC_us22_n706 ));
NOR2_X2 _AES_ENC_us22_U517  ( .A1(_AES_ENC_us22_n1117 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n707 ) );
NOR2_X2 _AES_ENC_us22_U516  ( .A1(_AES_ENC_sa22[4]), .A2(_AES_ENC_us22_n579 ), .ZN(_AES_ENC_us22_n705 ) );
NOR3_X2 _AES_ENC_us22_U515  ( .A1(_AES_ENC_us22_n707 ), .A2(_AES_ENC_us22_n706 ), .A3(_AES_ENC_us22_n705 ), .ZN(_AES_ENC_us22_n713 ) );
NOR4_X2 _AES_ENC_us22_U512  ( .A1(_AES_ENC_us22_n633 ), .A2(_AES_ENC_us22_n632 ), .A3(_AES_ENC_us22_n631 ), .A4(_AES_ENC_us22_n630 ), .ZN(_AES_ENC_us22_n634 ) );
NOR2_X2 _AES_ENC_us22_U510  ( .A1(_AES_ENC_us22_n629 ), .A2(_AES_ENC_us22_n628 ), .ZN(_AES_ENC_us22_n635 ) );
NAND3_X2 _AES_ENC_us22_U509  ( .A1(_AES_ENC_sa22[2]), .A2(_AES_ENC_sa22[7]), .A3(_AES_ENC_us22_n1059 ), .ZN(_AES_ENC_us22_n636 ) );
NOR2_X2 _AES_ENC_us22_U508  ( .A1(_AES_ENC_sa22[7]), .A2(_AES_ENC_sa22[2]),.ZN(_AES_ENC_us22_n794 ) );
NOR2_X2 _AES_ENC_us22_U507  ( .A1(_AES_ENC_sa22[4]), .A2(_AES_ENC_sa22[1]),.ZN(_AES_ENC_us22_n1102 ) );
NOR2_X2 _AES_ENC_us22_U506  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_sa22[3]), .ZN(_AES_ENC_us22_n1053 ) );
NOR2_X2 _AES_ENC_us22_U505  ( .A1(_AES_ENC_us22_n607 ), .A2(_AES_ENC_sa22[5]), .ZN(_AES_ENC_us22_n1024 ) );
NOR2_X2 _AES_ENC_us22_U504  ( .A1(_AES_ENC_us22_n625 ), .A2(_AES_ENC_sa22[2]), .ZN(_AES_ENC_us22_n1093 ) );
NOR2_X2 _AES_ENC_us22_U503  ( .A1(_AES_ENC_us22_n614 ), .A2(_AES_ENC_sa22[5]), .ZN(_AES_ENC_us22_n1094 ) );
NOR2_X2 _AES_ENC_us22_U502  ( .A1(_AES_ENC_us22_n624 ), .A2(_AES_ENC_sa22[3]), .ZN(_AES_ENC_us22_n931 ) );
INV_X4 _AES_ENC_us22_U501  ( .A(_AES_ENC_us22_n570 ), .ZN(_AES_ENC_us22_n573 ) );
NOR2_X2 _AES_ENC_us22_U500  ( .A1(_AES_ENC_us22_n1053 ), .A2(_AES_ENC_us22_n1095 ), .ZN(_AES_ENC_us22_n639 ) );
NOR3_X2 _AES_ENC_us22_U499  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n573 ), .A3(_AES_ENC_us22_n1074 ), .ZN(_AES_ENC_us22_n641 ) );
NOR2_X2 _AES_ENC_us22_U498  ( .A1(_AES_ENC_us22_n639 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n640 ) );
NOR2_X2 _AES_ENC_us22_U497  ( .A1(_AES_ENC_us22_n641 ), .A2(_AES_ENC_us22_n640 ), .ZN(_AES_ENC_us22_n646 ) );
NOR3_X2 _AES_ENC_us22_U496  ( .A1(_AES_ENC_us22_n995 ), .A2(_AES_ENC_us22_n586 ), .A3(_AES_ENC_us22_n994 ), .ZN(_AES_ENC_us22_n1002 ) );
NOR2_X2 _AES_ENC_us22_U495  ( .A1(_AES_ENC_us22_n909 ), .A2(_AES_ENC_us22_n908 ), .ZN(_AES_ENC_us22_n920 ) );
NOR2_X2 _AES_ENC_us22_U494  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n823 ) );
NOR2_X2 _AES_ENC_us22_U492  ( .A1(_AES_ENC_us22_n624 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n822 ) );
NOR2_X2 _AES_ENC_us22_U491  ( .A1(_AES_ENC_us22_n823 ), .A2(_AES_ENC_us22_n822 ), .ZN(_AES_ENC_us22_n825 ) );
NOR2_X2 _AES_ENC_us22_U490  ( .A1(_AES_ENC_sa22[1]), .A2(_AES_ENC_us22_n623 ), .ZN(_AES_ENC_us22_n913 ) );
NOR2_X2 _AES_ENC_us22_U489  ( .A1(_AES_ENC_us22_n913 ), .A2(_AES_ENC_us22_n1091 ), .ZN(_AES_ENC_us22_n914 ) );
NOR2_X2 _AES_ENC_us22_U488  ( .A1(_AES_ENC_us22_n826 ), .A2(_AES_ENC_us22_n572 ), .ZN(_AES_ENC_us22_n827 ) );
NOR3_X2 _AES_ENC_us22_U487  ( .A1(_AES_ENC_us22_n769 ), .A2(_AES_ENC_us22_n768 ), .A3(_AES_ENC_us22_n767 ), .ZN(_AES_ENC_us22_n775 ) );
NOR2_X2 _AES_ENC_us22_U486  ( .A1(_AES_ENC_us22_n1056 ), .A2(_AES_ENC_us22_n1053 ), .ZN(_AES_ENC_us22_n749 ) );
NOR2_X2 _AES_ENC_us22_U483  ( .A1(_AES_ENC_us22_n749 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n752 ) );
INV_X4 _AES_ENC_us22_U482  ( .A(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n596 ));
NOR2_X2 _AES_ENC_us22_U480  ( .A1(_AES_ENC_us22_n1054 ), .A2(_AES_ENC_us22_n1053 ), .ZN(_AES_ENC_us22_n1055 ) );
OR2_X4 _AES_ENC_us22_U479  ( .A1(_AES_ENC_us22_n1094 ), .A2(_AES_ENC_us22_n1093 ), .ZN(_AES_ENC_us22_n571 ) );
AND2_X2 _AES_ENC_us22_U478  ( .A1(_AES_ENC_us22_n571 ), .A2(_AES_ENC_us22_n1095 ), .ZN(_AES_ENC_us22_n1101 ) );
NOR2_X2 _AES_ENC_us22_U477  ( .A1(_AES_ENC_us22_n1074 ), .A2(_AES_ENC_us22_n931 ), .ZN(_AES_ENC_us22_n796 ) );
NOR2_X2 _AES_ENC_us22_U474  ( .A1(_AES_ENC_us22_n796 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n797 ) );
NOR2_X2 _AES_ENC_us22_U473  ( .A1(_AES_ENC_us22_n932 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n933 ) );
NOR2_X2 _AES_ENC_us22_U472  ( .A1(_AES_ENC_us22_n929 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n935 ) );
NOR2_X2 _AES_ENC_us22_U471  ( .A1(_AES_ENC_us22_n931 ), .A2(_AES_ENC_us22_n930 ), .ZN(_AES_ENC_us22_n934 ) );
NOR3_X2 _AES_ENC_us22_U470  ( .A1(_AES_ENC_us22_n935 ), .A2(_AES_ENC_us22_n934 ), .A3(_AES_ENC_us22_n933 ), .ZN(_AES_ENC_us22_n936 ) );
NOR2_X2 _AES_ENC_us22_U469  ( .A1(_AES_ENC_us22_n624 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n1075 ) );
NOR2_X2 _AES_ENC_us22_U468  ( .A1(_AES_ENC_us22_n572 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n949 ) );
NOR2_X2 _AES_ENC_us22_U467  ( .A1(_AES_ENC_us22_n1049 ), .A2(_AES_ENC_us22_n618 ), .ZN(_AES_ENC_us22_n1051 ) );
NOR2_X2 _AES_ENC_us22_U466  ( .A1(_AES_ENC_us22_n1051 ), .A2(_AES_ENC_us22_n1050 ), .ZN(_AES_ENC_us22_n1052 ) );
NOR2_X2 _AES_ENC_us22_U465  ( .A1(_AES_ENC_us22_n1052 ), .A2(_AES_ENC_us22_n592 ), .ZN(_AES_ENC_us22_n1064 ) );
NOR2_X2 _AES_ENC_us22_U464  ( .A1(_AES_ENC_sa22[1]), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n631 ) );
NOR2_X2 _AES_ENC_us22_U463  ( .A1(_AES_ENC_us22_n1025 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n980 ) );
NOR2_X2 _AES_ENC_us22_U462  ( .A1(_AES_ENC_us22_n1073 ), .A2(_AES_ENC_us22_n1094 ), .ZN(_AES_ENC_us22_n795 ) );
NOR2_X2 _AES_ENC_us22_U461  ( .A1(_AES_ENC_us22_n795 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n799 ) );
NOR2_X2 _AES_ENC_us22_U460  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n981 ) );
NOR2_X2 _AES_ENC_us22_U459  ( .A1(_AES_ENC_us22_n1102 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n643 ) );
NOR2_X2 _AES_ENC_us22_U458  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n621 ), .ZN(_AES_ENC_us22_n642 ) );
NOR2_X2 _AES_ENC_us22_U455  ( .A1(_AES_ENC_us22_n911 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n644 ) );
NOR4_X2 _AES_ENC_us22_U448  ( .A1(_AES_ENC_us22_n644 ), .A2(_AES_ENC_us22_n643 ), .A3(_AES_ENC_us22_n804 ), .A4(_AES_ENC_us22_n642 ), .ZN(_AES_ENC_us22_n645 ) );
NOR2_X2 _AES_ENC_us22_U447  ( .A1(_AES_ENC_us22_n1102 ), .A2(_AES_ENC_us22_n910 ), .ZN(_AES_ENC_us22_n932 ) );
NOR2_X2 _AES_ENC_us22_U442  ( .A1(_AES_ENC_us22_n1102 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n755 ) );
NOR2_X2 _AES_ENC_us22_U441  ( .A1(_AES_ENC_us22_n931 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n743 ) );
NOR2_X2 _AES_ENC_us22_U438  ( .A1(_AES_ENC_us22_n1072 ), .A2(_AES_ENC_us22_n1094 ), .ZN(_AES_ENC_us22_n930 ) );
NOR2_X2 _AES_ENC_us22_U435  ( .A1(_AES_ENC_us22_n1074 ), .A2(_AES_ENC_us22_n1025 ), .ZN(_AES_ENC_us22_n891 ) );
NOR2_X2 _AES_ENC_us22_U434  ( .A1(_AES_ENC_us22_n891 ), .A2(_AES_ENC_us22_n609 ), .ZN(_AES_ENC_us22_n894 ) );
NOR3_X2 _AES_ENC_us22_U433  ( .A1(_AES_ENC_us22_n623 ), .A2(_AES_ENC_sa22[1]), .A3(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n683 ));
INV_X4 _AES_ENC_us22_U428  ( .A(_AES_ENC_us22_n931 ), .ZN(_AES_ENC_us22_n623 ) );
NOR2_X2 _AES_ENC_us22_U427  ( .A1(_AES_ENC_us22_n996 ), .A2(_AES_ENC_us22_n931 ), .ZN(_AES_ENC_us22_n704 ) );
NOR2_X2 _AES_ENC_us22_U421  ( .A1(_AES_ENC_us22_n931 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n685 ) );
NOR2_X2 _AES_ENC_us22_U420  ( .A1(_AES_ENC_us22_n1029 ), .A2(_AES_ENC_us22_n1025 ), .ZN(_AES_ENC_us22_n1079 ) );
NOR3_X2 _AES_ENC_us22_U419  ( .A1(_AES_ENC_us22_n589 ), .A2(_AES_ENC_us22_n1025 ), .A3(_AES_ENC_us22_n616 ), .ZN(_AES_ENC_us22_n945 ) );
NOR2_X2 _AES_ENC_us22_U418  ( .A1(_AES_ENC_us22_n626 ), .A2(_AES_ENC_us22_n611 ), .ZN(_AES_ENC_us22_n800 ) );
NOR3_X2 _AES_ENC_us22_U417  ( .A1(_AES_ENC_us22_n590 ), .A2(_AES_ENC_us22_n627 ), .A3(_AES_ENC_us22_n611 ), .ZN(_AES_ENC_us22_n798 ) );
NOR3_X2 _AES_ENC_us22_U416  ( .A1(_AES_ENC_us22_n610 ), .A2(_AES_ENC_us22_n572 ), .A3(_AES_ENC_us22_n575 ), .ZN(_AES_ENC_us22_n962 ) );
NOR3_X2 _AES_ENC_us22_U415  ( .A1(_AES_ENC_us22_n959 ), .A2(_AES_ENC_us22_n572 ), .A3(_AES_ENC_us22_n609 ), .ZN(_AES_ENC_us22_n768 ) );
NOR3_X2 _AES_ENC_us22_U414  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n572 ), .A3(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n694 ) );
NOR3_X2 _AES_ENC_us22_U413  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n572 ), .A3(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n895 ) );
NOR3_X2 _AES_ENC_us22_U410  ( .A1(_AES_ENC_us22_n1008 ), .A2(_AES_ENC_us22_n1007 ), .A3(_AES_ENC_us22_n1006 ), .ZN(_AES_ENC_us22_n1018 ) );
NOR4_X2 _AES_ENC_us22_U409  ( .A1(_AES_ENC_us22_n806 ), .A2(_AES_ENC_us22_n805 ), .A3(_AES_ENC_us22_n804 ), .A4(_AES_ENC_us22_n803 ), .ZN(_AES_ENC_us22_n807 ) );
NOR3_X2 _AES_ENC_us22_U406  ( .A1(_AES_ENC_us22_n799 ), .A2(_AES_ENC_us22_n798 ), .A3(_AES_ENC_us22_n797 ), .ZN(_AES_ENC_us22_n808 ) );
NOR4_X2 _AES_ENC_us22_U405  ( .A1(_AES_ENC_us22_n843 ), .A2(_AES_ENC_us22_n842 ), .A3(_AES_ENC_us22_n841 ), .A4(_AES_ENC_us22_n840 ), .ZN(_AES_ENC_us22_n844 ) );
NOR2_X2 _AES_ENC_us22_U404  ( .A1(_AES_ENC_us22_n669 ), .A2(_AES_ENC_us22_n668 ), .ZN(_AES_ENC_us22_n673 ) );
NOR4_X2 _AES_ENC_us22_U403  ( .A1(_AES_ENC_us22_n946 ), .A2(_AES_ENC_us22_n1046 ), .A3(_AES_ENC_us22_n671 ), .A4(_AES_ENC_us22_n670 ), .ZN(_AES_ENC_us22_n672 ) );
NOR4_X2 _AES_ENC_us22_U401  ( .A1(_AES_ENC_us22_n711 ), .A2(_AES_ENC_us22_n710 ), .A3(_AES_ENC_us22_n709 ), .A4(_AES_ENC_us22_n708 ), .ZN(_AES_ENC_us22_n712 ) );
NOR4_X2 _AES_ENC_us22_U400  ( .A1(_AES_ENC_us22_n963 ), .A2(_AES_ENC_us22_n962 ), .A3(_AES_ENC_us22_n961 ), .A4(_AES_ENC_us22_n960 ), .ZN(_AES_ENC_us22_n964 ) );
NOR3_X2 _AES_ENC_us22_U399  ( .A1(_AES_ENC_us22_n1101 ), .A2(_AES_ENC_us22_n1100 ), .A3(_AES_ENC_us22_n1099 ), .ZN(_AES_ENC_us22_n1109 ) );
NOR3_X2 _AES_ENC_us22_U398  ( .A1(_AES_ENC_us22_n743 ), .A2(_AES_ENC_us22_n742 ), .A3(_AES_ENC_us22_n741 ), .ZN(_AES_ENC_us22_n744 ) );
NOR2_X2 _AES_ENC_us22_U397  ( .A1(_AES_ENC_us22_n697 ), .A2(_AES_ENC_us22_n658 ), .ZN(_AES_ENC_us22_n659 ) );
NOR2_X2 _AES_ENC_us22_U396  ( .A1(_AES_ENC_us22_n1078 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n1033 ) );
NOR2_X2 _AES_ENC_us22_U393  ( .A1(_AES_ENC_us22_n1031 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n1032 ) );
NOR3_X2 _AES_ENC_us22_U390  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n1025 ), .A3(_AES_ENC_us22_n1074 ), .ZN(_AES_ENC_us22_n1035 ) );
NOR4_X2 _AES_ENC_us22_U389  ( .A1(_AES_ENC_us22_n1035 ), .A2(_AES_ENC_us22_n1034 ), .A3(_AES_ENC_us22_n1033 ), .A4(_AES_ENC_us22_n1032 ), .ZN(_AES_ENC_us22_n1036 ) );
NOR2_X2 _AES_ENC_us22_U388  ( .A1(_AES_ENC_us22_n598 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n885 ) );
NOR2_X2 _AES_ENC_us22_U387  ( .A1(_AES_ENC_us22_n623 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n882 ) );
NOR2_X2 _AES_ENC_us22_U386  ( .A1(_AES_ENC_us22_n1053 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n884 ) );
NOR4_X2 _AES_ENC_us22_U385  ( .A1(_AES_ENC_us22_n885 ), .A2(_AES_ENC_us22_n884 ), .A3(_AES_ENC_us22_n883 ), .A4(_AES_ENC_us22_n882 ), .ZN(_AES_ENC_us22_n886 ) );
NOR2_X2 _AES_ENC_us22_U384  ( .A1(_AES_ENC_us22_n825 ), .A2(_AES_ENC_us22_n578 ), .ZN(_AES_ENC_us22_n830 ) );
NOR2_X2 _AES_ENC_us22_U383  ( .A1(_AES_ENC_us22_n827 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n829 ) );
NOR2_X2 _AES_ENC_us22_U382  ( .A1(_AES_ENC_us22_n572 ), .A2(_AES_ENC_us22_n579 ), .ZN(_AES_ENC_us22_n828 ) );
NOR4_X2 _AES_ENC_us22_U374  ( .A1(_AES_ENC_us22_n831 ), .A2(_AES_ENC_us22_n830 ), .A3(_AES_ENC_us22_n829 ), .A4(_AES_ENC_us22_n828 ), .ZN(_AES_ENC_us22_n832 ) );
NOR2_X2 _AES_ENC_us22_U373  ( .A1(_AES_ENC_us22_n606 ), .A2(_AES_ENC_us22_n582 ), .ZN(_AES_ENC_us22_n1104 ) );
NOR2_X2 _AES_ENC_us22_U372  ( .A1(_AES_ENC_us22_n1102 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n1106 ) );
NOR2_X2 _AES_ENC_us22_U370  ( .A1(_AES_ENC_us22_n1103 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n1105 ) );
NOR4_X2 _AES_ENC_us22_U369  ( .A1(_AES_ENC_us22_n1107 ), .A2(_AES_ENC_us22_n1106 ), .A3(_AES_ENC_us22_n1105 ), .A4(_AES_ENC_us22_n1104 ), .ZN(_AES_ENC_us22_n1108 ) );
NOR3_X2 _AES_ENC_us22_U368  ( .A1(_AES_ENC_us22_n959 ), .A2(_AES_ENC_us22_n621 ), .A3(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n963 ) );
NOR2_X2 _AES_ENC_us22_U367  ( .A1(_AES_ENC_us22_n626 ), .A2(_AES_ENC_us22_n627 ), .ZN(_AES_ENC_us22_n1114 ) );
INV_X4 _AES_ENC_us22_U366  ( .A(_AES_ENC_us22_n1024 ), .ZN(_AES_ENC_us22_n606 ) );
NOR3_X2 _AES_ENC_us22_U365  ( .A1(_AES_ENC_us22_n910 ), .A2(_AES_ENC_us22_n1059 ), .A3(_AES_ENC_us22_n611 ), .ZN(_AES_ENC_us22_n1115 ) );
INV_X4 _AES_ENC_us22_U364  ( .A(_AES_ENC_us22_n1094 ), .ZN(_AES_ENC_us22_n613 ) );
NOR2_X2 _AES_ENC_us22_U363  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n931 ), .ZN(_AES_ENC_us22_n1100 ) );
INV_X4 _AES_ENC_us22_U354  ( .A(_AES_ENC_us22_n1093 ), .ZN(_AES_ENC_us22_n617 ) );
NOR2_X2 _AES_ENC_us22_U353  ( .A1(_AES_ENC_us22_n569 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n929 ) );
NOR2_X2 _AES_ENC_us22_U352  ( .A1(_AES_ENC_us22_n620 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n926 ) );
NOR2_X2 _AES_ENC_us22_U351  ( .A1(_AES_ENC_us22_n572 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n1095 ) );
NOR2_X2 _AES_ENC_us22_U350  ( .A1(_AES_ENC_us22_n609 ), .A2(_AES_ENC_us22_n627 ), .ZN(_AES_ENC_us22_n1010 ) );
NOR2_X2 _AES_ENC_us22_U349  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n1103 ) );
NOR2_X2 _AES_ENC_us22_U348  ( .A1(_AES_ENC_us22_n622 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n1059 ) );
NOR2_X2 _AES_ENC_us22_U347  ( .A1(_AES_ENC_sa22[1]), .A2(_AES_ENC_us22_n1120 ), .ZN(_AES_ENC_us22_n1022 ) );
NOR2_X2 _AES_ENC_us22_U346  ( .A1(_AES_ENC_us22_n619 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n911 ) );
NOR2_X2 _AES_ENC_us22_U345  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_us22_n1025 ), .ZN(_AES_ENC_us22_n826 ) );
NOR2_X2 _AES_ENC_us22_U338  ( .A1(_AES_ENC_us22_n626 ), .A2(_AES_ENC_us22_n607 ), .ZN(_AES_ENC_us22_n1072 ) );
NOR2_X2 _AES_ENC_us22_U335  ( .A1(_AES_ENC_us22_n627 ), .A2(_AES_ENC_us22_n616 ), .ZN(_AES_ENC_us22_n956 ) );
NOR2_X2 _AES_ENC_us22_U329  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_us22_n624 ), .ZN(_AES_ENC_us22_n1121 ) );
NOR2_X2 _AES_ENC_us22_U328  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_us22_n624 ), .ZN(_AES_ENC_us22_n1058 ) );
NOR2_X2 _AES_ENC_us22_U327  ( .A1(_AES_ENC_us22_n625 ), .A2(_AES_ENC_us22_n611 ), .ZN(_AES_ENC_us22_n1073 ) );
NOR2_X2 _AES_ENC_us22_U325  ( .A1(_AES_ENC_sa22[1]), .A2(_AES_ENC_us22_n1025 ), .ZN(_AES_ENC_us22_n1054 ) );
NOR2_X2 _AES_ENC_us22_U324  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_us22_n931 ), .ZN(_AES_ENC_us22_n1029 ) );
NOR2_X2 _AES_ENC_us22_U319  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n1056 ) );
NOR2_X2 _AES_ENC_us22_U318  ( .A1(_AES_ENC_us22_n614 ), .A2(_AES_ENC_us22_n626 ), .ZN(_AES_ENC_us22_n1050 ) );
NOR2_X2 _AES_ENC_us22_U317  ( .A1(_AES_ENC_us22_n1121 ), .A2(_AES_ENC_us22_n1025 ), .ZN(_AES_ENC_us22_n1120 ) );
NOR2_X2 _AES_ENC_us22_U316  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_us22_n572 ), .ZN(_AES_ENC_us22_n1074 ) );
NOR2_X2 _AES_ENC_us22_U315  ( .A1(_AES_ENC_us22_n1058 ), .A2(_AES_ENC_us22_n1054 ), .ZN(_AES_ENC_us22_n878 ) );
NOR2_X2 _AES_ENC_us22_U314  ( .A1(_AES_ENC_us22_n878 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n879 ) );
NOR2_X2 _AES_ENC_us22_U312  ( .A1(_AES_ENC_us22_n880 ), .A2(_AES_ENC_us22_n879 ), .ZN(_AES_ENC_us22_n887 ) );
NOR2_X2 _AES_ENC_us22_U311  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n588 ), .ZN(_AES_ENC_us22_n957 ) );
NOR2_X2 _AES_ENC_us22_U310  ( .A1(_AES_ENC_us22_n958 ), .A2(_AES_ENC_us22_n957 ), .ZN(_AES_ENC_us22_n965 ) );
NOR3_X2 _AES_ENC_us22_U309  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n1091 ), .A3(_AES_ENC_us22_n1022 ), .ZN(_AES_ENC_us22_n720 ) );
NOR3_X2 _AES_ENC_us22_U303  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n1054 ), .A3(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n719 ) );
NOR2_X2 _AES_ENC_us22_U302  ( .A1(_AES_ENC_us22_n720 ), .A2(_AES_ENC_us22_n719 ), .ZN(_AES_ENC_us22_n726 ) );
NOR2_X2 _AES_ENC_us22_U300  ( .A1(_AES_ENC_us22_n614 ), .A2(_AES_ENC_us22_n591 ), .ZN(_AES_ENC_us22_n865 ) );
NOR2_X2 _AES_ENC_us22_U299  ( .A1(_AES_ENC_us22_n1059 ), .A2(_AES_ENC_us22_n1058 ), .ZN(_AES_ENC_us22_n1060 ) );
NOR2_X2 _AES_ENC_us22_U298  ( .A1(_AES_ENC_us22_n1095 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n668 ) );
NOR2_X2 _AES_ENC_us22_U297  ( .A1(_AES_ENC_us22_n826 ), .A2(_AES_ENC_us22_n573 ), .ZN(_AES_ENC_us22_n750 ) );
NOR2_X2 _AES_ENC_us22_U296  ( .A1(_AES_ENC_us22_n750 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n751 ) );
NOR2_X2 _AES_ENC_us22_U295  ( .A1(_AES_ENC_us22_n907 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n908 ) );
NOR2_X2 _AES_ENC_us22_U294  ( .A1(_AES_ENC_us22_n990 ), .A2(_AES_ENC_us22_n926 ), .ZN(_AES_ENC_us22_n780 ) );
NOR2_X2 _AES_ENC_us22_U293  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n584 ), .ZN(_AES_ENC_us22_n838 ) );
NOR2_X2 _AES_ENC_us22_U292  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n602 ), .ZN(_AES_ENC_us22_n837 ) );
NOR2_X2 _AES_ENC_us22_U291  ( .A1(_AES_ENC_us22_n838 ), .A2(_AES_ENC_us22_n837 ), .ZN(_AES_ENC_us22_n845 ) );
NOR2_X2 _AES_ENC_us22_U290  ( .A1(_AES_ENC_us22_n1022 ), .A2(_AES_ENC_us22_n1058 ), .ZN(_AES_ENC_us22_n740 ) );
NOR2_X2 _AES_ENC_us22_U284  ( .A1(_AES_ENC_us22_n740 ), .A2(_AES_ENC_us22_n616 ), .ZN(_AES_ENC_us22_n742 ) );
NOR2_X2 _AES_ENC_us22_U283  ( .A1(_AES_ENC_us22_n1098 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n1099 ) );
NOR2_X2 _AES_ENC_us22_U282  ( .A1(_AES_ENC_us22_n1120 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n993 ) );
NOR2_X2 _AES_ENC_us22_U281  ( .A1(_AES_ENC_us22_n993 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n994 ) );
NOR2_X2 _AES_ENC_us22_U280  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n620 ), .ZN(_AES_ENC_us22_n1026 ) );
NOR2_X2 _AES_ENC_us22_U279  ( .A1(_AES_ENC_us22_n573 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n1027 ) );
NOR2_X2 _AES_ENC_us22_U273  ( .A1(_AES_ENC_us22_n1027 ), .A2(_AES_ENC_us22_n1026 ), .ZN(_AES_ENC_us22_n1028 ) );
NOR2_X2 _AES_ENC_us22_U272  ( .A1(_AES_ENC_us22_n1029 ), .A2(_AES_ENC_us22_n1028 ), .ZN(_AES_ENC_us22_n1034 ) );
NOR4_X2 _AES_ENC_us22_U271  ( .A1(_AES_ENC_us22_n757 ), .A2(_AES_ENC_us22_n756 ), .A3(_AES_ENC_us22_n755 ), .A4(_AES_ENC_us22_n754 ), .ZN(_AES_ENC_us22_n758 ) );
NOR2_X2 _AES_ENC_us22_U270  ( .A1(_AES_ENC_us22_n752 ), .A2(_AES_ENC_us22_n751 ), .ZN(_AES_ENC_us22_n759 ) );
NOR2_X2 _AES_ENC_us22_U269  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n1071 ), .ZN(_AES_ENC_us22_n669 ) );
NOR2_X2 _AES_ENC_us22_U268  ( .A1(_AES_ENC_us22_n1056 ), .A2(_AES_ENC_us22_n990 ), .ZN(_AES_ENC_us22_n991 ) );
NOR2_X2 _AES_ENC_us22_U267  ( .A1(_AES_ENC_us22_n991 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n995 ) );
NOR2_X2 _AES_ENC_us22_U263  ( .A1(_AES_ENC_us22_n607 ), .A2(_AES_ENC_us22_n590 ), .ZN(_AES_ENC_us22_n1008 ) );
NOR2_X2 _AES_ENC_us22_U262  ( .A1(_AES_ENC_us22_n839 ), .A2(_AES_ENC_us22_n582 ), .ZN(_AES_ENC_us22_n693 ) );
NOR2_X2 _AES_ENC_us22_U258  ( .A1(_AES_ENC_us22_n606 ), .A2(_AES_ENC_us22_n906 ), .ZN(_AES_ENC_us22_n741 ) );
NOR2_X2 _AES_ENC_us22_U255  ( .A1(_AES_ENC_us22_n1054 ), .A2(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n763 ) );
NOR2_X2 _AES_ENC_us22_U254  ( .A1(_AES_ENC_us22_n763 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n769 ) );
NOR2_X2 _AES_ENC_us22_U253  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n577 ), .ZN(_AES_ENC_us22_n1007 ) );
NOR2_X2 _AES_ENC_us22_U252  ( .A1(_AES_ENC_us22_n609 ), .A2(_AES_ENC_us22_n580 ), .ZN(_AES_ENC_us22_n1123 ) );
NOR2_X2 _AES_ENC_us22_U251  ( .A1(_AES_ENC_us22_n609 ), .A2(_AES_ENC_us22_n590 ), .ZN(_AES_ENC_us22_n710 ) );
INV_X4 _AES_ENC_us22_U250  ( .A(_AES_ENC_us22_n1029 ), .ZN(_AES_ENC_us22_n582 ) );
NOR2_X2 _AES_ENC_us22_U243  ( .A1(_AES_ENC_us22_n616 ), .A2(_AES_ENC_us22_n597 ), .ZN(_AES_ENC_us22_n883 ) );
NOR2_X2 _AES_ENC_us22_U242  ( .A1(_AES_ENC_us22_n593 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n1125 ) );
NOR2_X2 _AES_ENC_us22_U241  ( .A1(_AES_ENC_us22_n911 ), .A2(_AES_ENC_us22_n910 ), .ZN(_AES_ENC_us22_n912 ) );
NOR2_X2 _AES_ENC_us22_U240  ( .A1(_AES_ENC_us22_n912 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n916 ) );
NOR2_X2 _AES_ENC_us22_U239  ( .A1(_AES_ENC_us22_n990 ), .A2(_AES_ENC_us22_n929 ), .ZN(_AES_ENC_us22_n892 ) );
NOR2_X2 _AES_ENC_us22_U238  ( .A1(_AES_ENC_us22_n892 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n893 ) );
NOR2_X2 _AES_ENC_us22_U237  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n602 ), .ZN(_AES_ENC_us22_n950 ) );
NOR2_X2 _AES_ENC_us22_U236  ( .A1(_AES_ENC_us22_n1079 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n1082 ) );
NOR2_X2 _AES_ENC_us22_U235  ( .A1(_AES_ENC_us22_n910 ), .A2(_AES_ENC_us22_n1056 ), .ZN(_AES_ENC_us22_n941 ) );
NOR2_X2 _AES_ENC_us22_U234  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n1077 ), .ZN(_AES_ENC_us22_n841 ) );
NOR2_X2 _AES_ENC_us22_U229  ( .A1(_AES_ENC_us22_n623 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n630 ) );
NOR2_X2 _AES_ENC_us22_U228  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n602 ), .ZN(_AES_ENC_us22_n806 ) );
NOR2_X2 _AES_ENC_us22_U227  ( .A1(_AES_ENC_us22_n623 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n948 ) );
NOR2_X2 _AES_ENC_us22_U226  ( .A1(_AES_ENC_us22_n606 ), .A2(_AES_ENC_us22_n589 ), .ZN(_AES_ENC_us22_n997 ) );
NOR2_X2 _AES_ENC_us22_U225  ( .A1(_AES_ENC_us22_n1121 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n1122 ) );
NOR2_X2 _AES_ENC_us22_U223  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n1023 ), .ZN(_AES_ENC_us22_n756 ) );
NOR2_X2 _AES_ENC_us22_U222  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n602 ), .ZN(_AES_ENC_us22_n870 ) );
NOR2_X2 _AES_ENC_us22_U221  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n569 ), .ZN(_AES_ENC_us22_n947 ) );
NOR2_X2 _AES_ENC_us22_U217  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n1077 ), .ZN(_AES_ENC_us22_n1084 ) );
NOR2_X2 _AES_ENC_us22_U213  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n855 ), .ZN(_AES_ENC_us22_n709 ) );
NOR2_X2 _AES_ENC_us22_U212  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n589 ), .ZN(_AES_ENC_us22_n868 ) );
NOR2_X2 _AES_ENC_us22_U211  ( .A1(_AES_ENC_us22_n1120 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n1124 ) );
NOR2_X2 _AES_ENC_us22_U210  ( .A1(_AES_ENC_us22_n1120 ), .A2(_AES_ENC_us22_n839 ), .ZN(_AES_ENC_us22_n842 ) );
NOR2_X2 _AES_ENC_us22_U209  ( .A1(_AES_ENC_us22_n1120 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n696 ) );
NOR2_X2 _AES_ENC_us22_U208  ( .A1(_AES_ENC_us22_n1074 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n1076 ) );
NOR2_X2 _AES_ENC_us22_U207  ( .A1(_AES_ENC_us22_n1074 ), .A2(_AES_ENC_us22_n620 ), .ZN(_AES_ENC_us22_n781 ) );
NOR3_X2 _AES_ENC_us22_U201  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n1056 ), .A3(_AES_ENC_us22_n990 ), .ZN(_AES_ENC_us22_n979 ) );
NOR3_X2 _AES_ENC_us22_U200  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n1058 ), .A3(_AES_ENC_us22_n1059 ), .ZN(_AES_ENC_us22_n854 ) );
NOR2_X2 _AES_ENC_us22_U199  ( .A1(_AES_ENC_us22_n996 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n869 ) );
NOR2_X2 _AES_ENC_us22_U198  ( .A1(_AES_ENC_us22_n1056 ), .A2(_AES_ENC_us22_n1074 ), .ZN(_AES_ENC_us22_n1057 ) );
NOR3_X2 _AES_ENC_us22_U197  ( .A1(_AES_ENC_us22_n607 ), .A2(_AES_ENC_us22_n1120 ), .A3(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n978 ) );
NOR2_X2 _AES_ENC_us22_U196  ( .A1(_AES_ENC_us22_n996 ), .A2(_AES_ENC_us22_n911 ), .ZN(_AES_ENC_us22_n1116 ) );
NOR2_X2 _AES_ENC_us22_U195  ( .A1(_AES_ENC_us22_n1074 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n754 ) );
NOR2_X2 _AES_ENC_us22_U194  ( .A1(_AES_ENC_us22_n926 ), .A2(_AES_ENC_us22_n1103 ), .ZN(_AES_ENC_us22_n977 ) );
NOR2_X2 _AES_ENC_us22_U187  ( .A1(_AES_ENC_us22_n839 ), .A2(_AES_ENC_us22_n824 ), .ZN(_AES_ENC_us22_n1092 ) );
NOR2_X2 _AES_ENC_us22_U186  ( .A1(_AES_ENC_us22_n573 ), .A2(_AES_ENC_us22_n1074 ), .ZN(_AES_ENC_us22_n684 ) );
NOR2_X2 _AES_ENC_us22_U185  ( .A1(_AES_ENC_us22_n826 ), .A2(_AES_ENC_us22_n1059 ), .ZN(_AES_ENC_us22_n907 ) );
NOR3_X2 _AES_ENC_us22_U184  ( .A1(_AES_ENC_us22_n625 ), .A2(_AES_ENC_us22_n1115 ), .A3(_AES_ENC_us22_n585 ), .ZN(_AES_ENC_us22_n831 ) );
NOR3_X2 _AES_ENC_us22_U183  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n1056 ), .A3(_AES_ENC_us22_n990 ), .ZN(_AES_ENC_us22_n896 ) );
NOR3_X2 _AES_ENC_us22_U182  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n573 ), .A3(_AES_ENC_us22_n1013 ), .ZN(_AES_ENC_us22_n670 ) );
NOR3_X2 _AES_ENC_us22_U181  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n1091 ), .A3(_AES_ENC_us22_n1022 ), .ZN(_AES_ENC_us22_n843 ) );
NOR2_X2 _AES_ENC_us22_U180  ( .A1(_AES_ENC_us22_n1029 ), .A2(_AES_ENC_us22_n1095 ), .ZN(_AES_ENC_us22_n735 ) );
NOR2_X2 _AES_ENC_us22_U174  ( .A1(_AES_ENC_us22_n1100 ), .A2(_AES_ENC_us22_n854 ), .ZN(_AES_ENC_us22_n860 ) );
NAND3_X2 _AES_ENC_us22_U173  ( .A1(_AES_ENC_us22_n569 ), .A2(_AES_ENC_us22_n582 ), .A3(_AES_ENC_us22_n681 ), .ZN(_AES_ENC_us22_n691 ) );
NOR2_X2 _AES_ENC_us22_U172  ( .A1(_AES_ENC_us22_n683 ), .A2(_AES_ENC_us22_n682 ), .ZN(_AES_ENC_us22_n690 ) );
NOR3_X2 _AES_ENC_us22_U171  ( .A1(_AES_ENC_us22_n695 ), .A2(_AES_ENC_us22_n694 ), .A3(_AES_ENC_us22_n693 ), .ZN(_AES_ENC_us22_n700 ) );
NOR4_X2 _AES_ENC_us22_U170  ( .A1(_AES_ENC_us22_n983 ), .A2(_AES_ENC_us22_n698 ), .A3(_AES_ENC_us22_n697 ), .A4(_AES_ENC_us22_n696 ), .ZN(_AES_ENC_us22_n699 ) );
NOR4_X2 _AES_ENC_us22_U169  ( .A1(_AES_ENC_us22_n896 ), .A2(_AES_ENC_us22_n895 ), .A3(_AES_ENC_us22_n894 ), .A4(_AES_ENC_us22_n893 ), .ZN(_AES_ENC_us22_n897 ) );
NOR2_X2 _AES_ENC_us22_U168  ( .A1(_AES_ENC_us22_n866 ), .A2(_AES_ENC_us22_n865 ), .ZN(_AES_ENC_us22_n872 ) );
NOR4_X2 _AES_ENC_us22_U162  ( .A1(_AES_ENC_us22_n870 ), .A2(_AES_ENC_us22_n869 ), .A3(_AES_ENC_us22_n868 ), .A4(_AES_ENC_us22_n867 ), .ZN(_AES_ENC_us22_n871 ) );
NOR2_X2 _AES_ENC_us22_U161  ( .A1(_AES_ENC_us22_n946 ), .A2(_AES_ENC_us22_n945 ), .ZN(_AES_ENC_us22_n952 ) );
NOR4_X2 _AES_ENC_us22_U160  ( .A1(_AES_ENC_us22_n950 ), .A2(_AES_ENC_us22_n949 ), .A3(_AES_ENC_us22_n948 ), .A4(_AES_ENC_us22_n947 ), .ZN(_AES_ENC_us22_n951 ) );
NOR4_X2 _AES_ENC_us22_U159  ( .A1(_AES_ENC_us22_n983 ), .A2(_AES_ENC_us22_n982 ), .A3(_AES_ENC_us22_n981 ), .A4(_AES_ENC_us22_n980 ), .ZN(_AES_ENC_us22_n984 ) );
NOR2_X2 _AES_ENC_us22_U158  ( .A1(_AES_ENC_us22_n979 ), .A2(_AES_ENC_us22_n978 ), .ZN(_AES_ENC_us22_n985 ) );
NOR4_X2 _AES_ENC_us22_U157  ( .A1(_AES_ENC_us22_n1125 ), .A2(_AES_ENC_us22_n1124 ), .A3(_AES_ENC_us22_n1123 ), .A4(_AES_ENC_us22_n1122 ), .ZN(_AES_ENC_us22_n1126 ) );
NOR4_X2 _AES_ENC_us22_U156  ( .A1(_AES_ENC_us22_n1084 ), .A2(_AES_ENC_us22_n1083 ), .A3(_AES_ENC_us22_n1082 ), .A4(_AES_ENC_us22_n1081 ), .ZN(_AES_ENC_us22_n1085 ) );
NOR2_X2 _AES_ENC_us22_U155  ( .A1(_AES_ENC_us22_n1076 ), .A2(_AES_ENC_us22_n1075 ), .ZN(_AES_ENC_us22_n1086 ) );
NOR3_X2 _AES_ENC_us22_U154  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n1054 ), .A3(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n961 ) );
NOR3_X2 _AES_ENC_us22_U153  ( .A1(_AES_ENC_us22_n620 ), .A2(_AES_ENC_us22_n1074 ), .A3(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n671 ) );
NOR2_X2 _AES_ENC_us22_U152  ( .A1(_AES_ENC_us22_n1057 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n1062 ) );
NOR2_X2 _AES_ENC_us22_U143  ( .A1(_AES_ENC_us22_n1055 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n1063 ) );
NOR2_X2 _AES_ENC_us22_U142  ( .A1(_AES_ENC_us22_n1060 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n1061 ) );
NOR4_X2 _AES_ENC_us22_U141  ( .A1(_AES_ENC_us22_n1064 ), .A2(_AES_ENC_us22_n1063 ), .A3(_AES_ENC_us22_n1062 ), .A4(_AES_ENC_us22_n1061 ), .ZN(_AES_ENC_us22_n1065 ) );
NOR3_X2 _AES_ENC_us22_U140  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n1120 ), .A3(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n918 ) );
NOR3_X2 _AES_ENC_us22_U132  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n573 ), .A3(_AES_ENC_us22_n1013 ), .ZN(_AES_ENC_us22_n917 ) );
NOR2_X2 _AES_ENC_us22_U131  ( .A1(_AES_ENC_us22_n914 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n915 ) );
NOR4_X2 _AES_ENC_us22_U130  ( .A1(_AES_ENC_us22_n918 ), .A2(_AES_ENC_us22_n917 ), .A3(_AES_ENC_us22_n916 ), .A4(_AES_ENC_us22_n915 ), .ZN(_AES_ENC_us22_n919 ) );
NOR2_X2 _AES_ENC_us22_U129  ( .A1(_AES_ENC_us22_n616 ), .A2(_AES_ENC_us22_n580 ), .ZN(_AES_ENC_us22_n771 ) );
NOR2_X2 _AES_ENC_us22_U128  ( .A1(_AES_ENC_us22_n1103 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n772 ) );
NOR2_X2 _AES_ENC_us22_U127  ( .A1(_AES_ENC_us22_n610 ), .A2(_AES_ENC_us22_n599 ), .ZN(_AES_ENC_us22_n773 ) );
NOR4_X2 _AES_ENC_us22_U126  ( .A1(_AES_ENC_us22_n773 ), .A2(_AES_ENC_us22_n772 ), .A3(_AES_ENC_us22_n771 ), .A4(_AES_ENC_us22_n770 ), .ZN(_AES_ENC_us22_n774 ) );
NOR2_X2 _AES_ENC_us22_U121  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n595 ), .ZN(_AES_ENC_us22_n858 ) );
NOR2_X2 _AES_ENC_us22_U120  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n855 ), .ZN(_AES_ENC_us22_n857 ) );
NOR2_X2 _AES_ENC_us22_U119  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n587 ), .ZN(_AES_ENC_us22_n856 ) );
NOR4_X2 _AES_ENC_us22_U118  ( .A1(_AES_ENC_us22_n858 ), .A2(_AES_ENC_us22_n857 ), .A3(_AES_ENC_us22_n856 ), .A4(_AES_ENC_us22_n958 ), .ZN(_AES_ENC_us22_n859 ) );
NOR2_X2 _AES_ENC_us22_U117  ( .A1(_AES_ENC_us22_n735 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n687 ) );
NOR2_X2 _AES_ENC_us22_U116  ( .A1(_AES_ENC_us22_n684 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n688 ) );
NOR2_X2 _AES_ENC_us22_U115  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n600 ), .ZN(_AES_ENC_us22_n686 ) );
NOR4_X2 _AES_ENC_us22_U106  ( .A1(_AES_ENC_us22_n688 ), .A2(_AES_ENC_us22_n687 ), .A3(_AES_ENC_us22_n686 ), .A4(_AES_ENC_us22_n685 ), .ZN(_AES_ENC_us22_n689 ) );
NOR2_X2 _AES_ENC_us22_U105  ( .A1(_AES_ENC_us22_n780 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n784 ) );
NOR2_X2 _AES_ENC_us22_U104  ( .A1(_AES_ENC_us22_n1117 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n782 ) );
NOR2_X2 _AES_ENC_us22_U103  ( .A1(_AES_ENC_us22_n781 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n783 ) );
NOR4_X2 _AES_ENC_us22_U102  ( .A1(_AES_ENC_us22_n880 ), .A2(_AES_ENC_us22_n784 ), .A3(_AES_ENC_us22_n783 ), .A4(_AES_ENC_us22_n782 ), .ZN(_AES_ENC_us22_n785 ) );
NOR2_X2 _AES_ENC_us22_U101  ( .A1(_AES_ENC_us22_n583 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n814 ) );
NOR2_X2 _AES_ENC_us22_U100  ( .A1(_AES_ENC_us22_n907 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n813 ) );
NOR3_X2 _AES_ENC_us22_U95  ( .A1(_AES_ENC_us22_n606 ), .A2(_AES_ENC_us22_n1058 ), .A3(_AES_ENC_us22_n1059 ), .ZN(_AES_ENC_us22_n815 ) );
NOR4_X2 _AES_ENC_us22_U94  ( .A1(_AES_ENC_us22_n815 ), .A2(_AES_ENC_us22_n814 ), .A3(_AES_ENC_us22_n813 ), .A4(_AES_ENC_us22_n812 ), .ZN(_AES_ENC_us22_n816 ) );
NOR2_X2 _AES_ENC_us22_U93  ( .A1(_AES_ENC_us22_n617 ), .A2(_AES_ENC_us22_n569 ), .ZN(_AES_ENC_us22_n721 ) );
NOR2_X2 _AES_ENC_us22_U92  ( .A1(_AES_ENC_us22_n1031 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n723 ) );
NOR2_X2 _AES_ENC_us22_U91  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n1096 ), .ZN(_AES_ENC_us22_n722 ) );
NOR4_X2 _AES_ENC_us22_U90  ( .A1(_AES_ENC_us22_n724 ), .A2(_AES_ENC_us22_n723 ), .A3(_AES_ENC_us22_n722 ), .A4(_AES_ENC_us22_n721 ), .ZN(_AES_ENC_us22_n725 ) );
NOR2_X2 _AES_ENC_us22_U89  ( .A1(_AES_ENC_us22_n911 ), .A2(_AES_ENC_us22_n990 ), .ZN(_AES_ENC_us22_n1009 ) );
NOR2_X2 _AES_ENC_us22_U88  ( .A1(_AES_ENC_us22_n1013 ), .A2(_AES_ENC_us22_n573 ), .ZN(_AES_ENC_us22_n1014 ) );
NOR2_X2 _AES_ENC_us22_U87  ( .A1(_AES_ENC_us22_n1014 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n1015 ) );
NOR4_X2 _AES_ENC_us22_U86  ( .A1(_AES_ENC_us22_n1016 ), .A2(_AES_ENC_us22_n1015 ), .A3(_AES_ENC_us22_n1119 ), .A4(_AES_ENC_us22_n1046 ), .ZN(_AES_ENC_us22_n1017 ) );
NOR2_X2 _AES_ENC_us22_U81  ( .A1(_AES_ENC_us22_n996 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n998 ) );
NOR2_X2 _AES_ENC_us22_U80  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n577 ), .ZN(_AES_ENC_us22_n1000 ) );
NOR2_X2 _AES_ENC_us22_U79  ( .A1(_AES_ENC_us22_n616 ), .A2(_AES_ENC_us22_n1096 ), .ZN(_AES_ENC_us22_n999 ) );
NOR4_X2 _AES_ENC_us22_U78  ( .A1(_AES_ENC_us22_n1000 ), .A2(_AES_ENC_us22_n999 ), .A3(_AES_ENC_us22_n998 ), .A4(_AES_ENC_us22_n997 ), .ZN(_AES_ENC_us22_n1001 ) );
NOR2_X2 _AES_ENC_us22_U74  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n1096 ), .ZN(_AES_ENC_us22_n697 ) );
NOR2_X2 _AES_ENC_us22_U73  ( .A1(_AES_ENC_us22_n620 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n958 ) );
NOR2_X2 _AES_ENC_us22_U72  ( .A1(_AES_ENC_us22_n911 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n983 ) );
NOR2_X2 _AES_ENC_us22_U71  ( .A1(_AES_ENC_us22_n1054 ), .A2(_AES_ENC_us22_n1103 ), .ZN(_AES_ENC_us22_n1031 ) );
INV_X4 _AES_ENC_us22_U65  ( .A(_AES_ENC_us22_n1050 ), .ZN(_AES_ENC_us22_n612 ) );
INV_X4 _AES_ENC_us22_U64  ( .A(_AES_ENC_us22_n1072 ), .ZN(_AES_ENC_us22_n605 ) );
INV_X4 _AES_ENC_us22_U63  ( .A(_AES_ENC_us22_n1073 ), .ZN(_AES_ENC_us22_n604 ) );
NOR2_X2 _AES_ENC_us22_U62  ( .A1(_AES_ENC_us22_n582 ), .A2(_AES_ENC_us22_n613 ), .ZN(_AES_ENC_us22_n880 ) );
NOR3_X2 _AES_ENC_us22_U61  ( .A1(_AES_ENC_us22_n826 ), .A2(_AES_ENC_us22_n1121 ), .A3(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n946 ) );
INV_X4 _AES_ENC_us22_U59  ( .A(_AES_ENC_us22_n1010 ), .ZN(_AES_ENC_us22_n608 ) );
NOR3_X2 _AES_ENC_us22_U58  ( .A1(_AES_ENC_us22_n573 ), .A2(_AES_ENC_us22_n1029 ), .A3(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n1119 ) );
INV_X4 _AES_ENC_us22_U57  ( .A(_AES_ENC_us22_n956 ), .ZN(_AES_ENC_us22_n615 ) );
NOR2_X2 _AES_ENC_us22_U50  ( .A1(_AES_ENC_us22_n623 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n1013 ) );
NOR2_X2 _AES_ENC_us22_U49  ( .A1(_AES_ENC_us22_n620 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n910 ) );
NOR2_X2 _AES_ENC_us22_U48  ( .A1(_AES_ENC_us22_n569 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n1091 ) );
NOR2_X2 _AES_ENC_us22_U47  ( .A1(_AES_ENC_us22_n622 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n990 ) );
NOR2_X2 _AES_ENC_us22_U46  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_us22_n1121 ), .ZN(_AES_ENC_us22_n996 ) );
NOR2_X2 _AES_ENC_us22_U45  ( .A1(_AES_ENC_us22_n610 ), .A2(_AES_ENC_us22_n600 ), .ZN(_AES_ENC_us22_n628 ) );
NOR2_X2 _AES_ENC_us22_U44  ( .A1(_AES_ENC_us22_n576 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n866 ) );
NOR2_X2 _AES_ENC_us22_U43  ( .A1(_AES_ENC_us22_n603 ), .A2(_AES_ENC_us22_n610 ), .ZN(_AES_ENC_us22_n1006 ) );
NOR2_X2 _AES_ENC_us22_U42  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n1117 ), .ZN(_AES_ENC_us22_n1118 ) );
NOR2_X2 _AES_ENC_us22_U41  ( .A1(_AES_ENC_us22_n1119 ), .A2(_AES_ENC_us22_n1118 ), .ZN(_AES_ENC_us22_n1127 ) );
NOR2_X2 _AES_ENC_us22_U36  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n594 ), .ZN(_AES_ENC_us22_n629 ) );
NOR2_X2 _AES_ENC_us22_U35  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n906 ), .ZN(_AES_ENC_us22_n909 ) );
NOR2_X2 _AES_ENC_us22_U34  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n597 ), .ZN(_AES_ENC_us22_n658 ) );
NOR2_X2 _AES_ENC_us22_U33  ( .A1(_AES_ENC_us22_n1116 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n695 ) );
NOR2_X2 _AES_ENC_us22_U32  ( .A1(_AES_ENC_us22_n1078 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n1083 ) );
NOR2_X2 _AES_ENC_us22_U31  ( .A1(_AES_ENC_us22_n941 ), .A2(_AES_ENC_us22_n608 ), .ZN(_AES_ENC_us22_n724 ) );
NOR2_X2 _AES_ENC_us22_U30  ( .A1(_AES_ENC_us22_n598 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n1107 ) );
NOR2_X2 _AES_ENC_us22_U29  ( .A1(_AES_ENC_us22_n576 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n840 ) );
NOR2_X2 _AES_ENC_us22_U24  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n593 ), .ZN(_AES_ENC_us22_n633 ) );
NOR2_X2 _AES_ENC_us22_U23  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n1080 ), .ZN(_AES_ENC_us22_n1081 ) );
NOR2_X2 _AES_ENC_us22_U21  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n1045 ), .ZN(_AES_ENC_us22_n812 ) );
NOR2_X2 _AES_ENC_us22_U20  ( .A1(_AES_ENC_us22_n1009 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n960 ) );
NOR2_X2 _AES_ENC_us22_U19  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n601 ), .ZN(_AES_ENC_us22_n982 ) );
NOR2_X2 _AES_ENC_us22_U18  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n594 ), .ZN(_AES_ENC_us22_n757 ) );
NOR2_X2 _AES_ENC_us22_U17  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n590 ), .ZN(_AES_ENC_us22_n698 ) );
NOR2_X2 _AES_ENC_us22_U16  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n619 ), .ZN(_AES_ENC_us22_n708 ) );
NOR2_X2 _AES_ENC_us22_U15  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n582 ), .ZN(_AES_ENC_us22_n770 ) );
NOR2_X2 _AES_ENC_us22_U10  ( .A1(_AES_ENC_us22_n619 ), .A2(_AES_ENC_us22_n604 ), .ZN(_AES_ENC_us22_n803 ) );
NOR2_X2 _AES_ENC_us22_U9  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n881 ), .ZN(_AES_ENC_us22_n711 ) );
NOR2_X2 _AES_ENC_us22_U8  ( .A1(_AES_ENC_us22_n615 ), .A2(_AES_ENC_us22_n582 ), .ZN(_AES_ENC_us22_n867 ) );
NOR2_X2 _AES_ENC_us22_U7  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n599 ), .ZN(_AES_ENC_us22_n804 ) );
NOR2_X2 _AES_ENC_us22_U6  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n620 ), .ZN(_AES_ENC_us22_n1046 ) );
OR2_X4 _AES_ENC_us22_U5  ( .A1(_AES_ENC_us22_n624 ), .A2(_AES_ENC_sa22[1]),.ZN(_AES_ENC_us22_n570 ) );
OR2_X4 _AES_ENC_us22_U4  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_sa22[4]),.ZN(_AES_ENC_us22_n569 ) );
NAND2_X2 _AES_ENC_us22_U514  ( .A1(_AES_ENC_us22_n1121 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n1030 ) );
AND2_X2 _AES_ENC_us22_U513  ( .A1(_AES_ENC_us22_n597 ), .A2(_AES_ENC_us22_n1030 ), .ZN(_AES_ENC_us22_n1049 ) );
NAND2_X2 _AES_ENC_us22_U511  ( .A1(_AES_ENC_us22_n1049 ), .A2(_AES_ENC_us22_n794 ), .ZN(_AES_ENC_us22_n637 ) );
AND2_X2 _AES_ENC_us22_U493  ( .A1(_AES_ENC_us22_n779 ), .A2(_AES_ENC_us22_n996 ), .ZN(_AES_ENC_us22_n632 ) );
NAND4_X2 _AES_ENC_us22_U485  ( .A1(_AES_ENC_us22_n637 ), .A2(_AES_ENC_us22_n636 ), .A3(_AES_ENC_us22_n635 ), .A4(_AES_ENC_us22_n634 ), .ZN(_AES_ENC_us22_n638 ) );
NAND2_X2 _AES_ENC_us22_U484  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n638 ), .ZN(_AES_ENC_us22_n679 ) );
NAND2_X2 _AES_ENC_us22_U481  ( .A1(_AES_ENC_us22_n1094 ), .A2(_AES_ENC_us22_n591 ), .ZN(_AES_ENC_us22_n648 ) );
NAND2_X2 _AES_ENC_us22_U476  ( .A1(_AES_ENC_us22_n601 ), .A2(_AES_ENC_us22_n590 ), .ZN(_AES_ENC_us22_n762 ) );
NAND2_X2 _AES_ENC_us22_U475  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n762 ), .ZN(_AES_ENC_us22_n647 ) );
NAND4_X2 _AES_ENC_us22_U457  ( .A1(_AES_ENC_us22_n648 ), .A2(_AES_ENC_us22_n647 ), .A3(_AES_ENC_us22_n646 ), .A4(_AES_ENC_us22_n645 ), .ZN(_AES_ENC_us22_n649 ) );
NAND2_X2 _AES_ENC_us22_U456  ( .A1(_AES_ENC_sa22[0]), .A2(_AES_ENC_us22_n649 ), .ZN(_AES_ENC_us22_n665 ) );
NAND2_X2 _AES_ENC_us22_U454  ( .A1(_AES_ENC_us22_n596 ), .A2(_AES_ENC_us22_n623 ), .ZN(_AES_ENC_us22_n855 ) );
NAND2_X2 _AES_ENC_us22_U453  ( .A1(_AES_ENC_us22_n587 ), .A2(_AES_ENC_us22_n855 ), .ZN(_AES_ENC_us22_n821 ) );
NAND2_X2 _AES_ENC_us22_U452  ( .A1(_AES_ENC_us22_n1093 ), .A2(_AES_ENC_us22_n821 ), .ZN(_AES_ENC_us22_n662 ) );
NAND2_X2 _AES_ENC_us22_U451  ( .A1(_AES_ENC_us22_n619 ), .A2(_AES_ENC_us22_n589 ), .ZN(_AES_ENC_us22_n650 ) );
NAND2_X2 _AES_ENC_us22_U450  ( .A1(_AES_ENC_us22_n956 ), .A2(_AES_ENC_us22_n650 ), .ZN(_AES_ENC_us22_n661 ) );
NAND2_X2 _AES_ENC_us22_U449  ( .A1(_AES_ENC_us22_n626 ), .A2(_AES_ENC_us22_n627 ), .ZN(_AES_ENC_us22_n839 ) );
OR2_X2 _AES_ENC_us22_U446  ( .A1(_AES_ENC_us22_n839 ), .A2(_AES_ENC_us22_n932 ), .ZN(_AES_ENC_us22_n656 ) );
NAND2_X2 _AES_ENC_us22_U445  ( .A1(_AES_ENC_us22_n621 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n1096 ) );
NAND2_X2 _AES_ENC_us22_U444  ( .A1(_AES_ENC_us22_n1030 ), .A2(_AES_ENC_us22_n1096 ), .ZN(_AES_ENC_us22_n651 ) );
NAND2_X2 _AES_ENC_us22_U443  ( .A1(_AES_ENC_us22_n1114 ), .A2(_AES_ENC_us22_n651 ), .ZN(_AES_ENC_us22_n655 ) );
OR3_X2 _AES_ENC_us22_U440  ( .A1(_AES_ENC_us22_n1079 ), .A2(_AES_ENC_sa22[7]), .A3(_AES_ENC_us22_n626 ), .ZN(_AES_ENC_us22_n654 ));
NAND2_X2 _AES_ENC_us22_U439  ( .A1(_AES_ENC_us22_n593 ), .A2(_AES_ENC_us22_n601 ), .ZN(_AES_ENC_us22_n652 ) );
NAND4_X2 _AES_ENC_us22_U437  ( .A1(_AES_ENC_us22_n656 ), .A2(_AES_ENC_us22_n655 ), .A3(_AES_ENC_us22_n654 ), .A4(_AES_ENC_us22_n653 ), .ZN(_AES_ENC_us22_n657 ) );
NAND2_X2 _AES_ENC_us22_U436  ( .A1(_AES_ENC_sa22[2]), .A2(_AES_ENC_us22_n657 ), .ZN(_AES_ENC_us22_n660 ) );
NAND4_X2 _AES_ENC_us22_U432  ( .A1(_AES_ENC_us22_n662 ), .A2(_AES_ENC_us22_n661 ), .A3(_AES_ENC_us22_n660 ), .A4(_AES_ENC_us22_n659 ), .ZN(_AES_ENC_us22_n663 ) );
NAND2_X2 _AES_ENC_us22_U431  ( .A1(_AES_ENC_us22_n663 ), .A2(_AES_ENC_us22_n574 ), .ZN(_AES_ENC_us22_n664 ) );
NAND2_X2 _AES_ENC_us22_U430  ( .A1(_AES_ENC_us22_n665 ), .A2(_AES_ENC_us22_n664 ), .ZN(_AES_ENC_us22_n666 ) );
NAND2_X2 _AES_ENC_us22_U429  ( .A1(_AES_ENC_sa22[6]), .A2(_AES_ENC_us22_n666 ), .ZN(_AES_ENC_us22_n678 ) );
NAND2_X2 _AES_ENC_us22_U426  ( .A1(_AES_ENC_us22_n735 ), .A2(_AES_ENC_us22_n1093 ), .ZN(_AES_ENC_us22_n675 ) );
NAND2_X2 _AES_ENC_us22_U425  ( .A1(_AES_ENC_us22_n588 ), .A2(_AES_ENC_us22_n597 ), .ZN(_AES_ENC_us22_n1045 ) );
OR2_X2 _AES_ENC_us22_U424  ( .A1(_AES_ENC_us22_n1045 ), .A2(_AES_ENC_us22_n605 ), .ZN(_AES_ENC_us22_n674 ) );
NAND2_X2 _AES_ENC_us22_U423  ( .A1(_AES_ENC_sa22[1]), .A2(_AES_ENC_us22_n620 ), .ZN(_AES_ENC_us22_n667 ) );
NAND2_X2 _AES_ENC_us22_U422  ( .A1(_AES_ENC_us22_n619 ), .A2(_AES_ENC_us22_n667 ), .ZN(_AES_ENC_us22_n1071 ) );
NAND4_X2 _AES_ENC_us22_U412  ( .A1(_AES_ENC_us22_n675 ), .A2(_AES_ENC_us22_n674 ), .A3(_AES_ENC_us22_n673 ), .A4(_AES_ENC_us22_n672 ), .ZN(_AES_ENC_us22_n676 ) );
NAND2_X2 _AES_ENC_us22_U411  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n676 ), .ZN(_AES_ENC_us22_n677 ) );
NAND2_X2 _AES_ENC_us22_U408  ( .A1(_AES_ENC_us22_n800 ), .A2(_AES_ENC_us22_n1022 ), .ZN(_AES_ENC_us22_n680 ) );
NAND2_X2 _AES_ENC_us22_U407  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n680 ), .ZN(_AES_ENC_us22_n681 ) );
AND2_X2 _AES_ENC_us22_U402  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n684 ), .ZN(_AES_ENC_us22_n682 ) );
NAND4_X2 _AES_ENC_us22_U395  ( .A1(_AES_ENC_us22_n691 ), .A2(_AES_ENC_us22_n581 ), .A3(_AES_ENC_us22_n690 ), .A4(_AES_ENC_us22_n689 ), .ZN(_AES_ENC_us22_n692 ) );
NAND2_X2 _AES_ENC_us22_U394  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n692 ), .ZN(_AES_ENC_us22_n733 ) );
NAND2_X2 _AES_ENC_us22_U392  ( .A1(_AES_ENC_us22_n977 ), .A2(_AES_ENC_us22_n1050 ), .ZN(_AES_ENC_us22_n702 ) );
NAND2_X2 _AES_ENC_us22_U391  ( .A1(_AES_ENC_us22_n1093 ), .A2(_AES_ENC_us22_n1045 ), .ZN(_AES_ENC_us22_n701 ) );
NAND4_X2 _AES_ENC_us22_U381  ( .A1(_AES_ENC_us22_n702 ), .A2(_AES_ENC_us22_n701 ), .A3(_AES_ENC_us22_n700 ), .A4(_AES_ENC_us22_n699 ), .ZN(_AES_ENC_us22_n703 ) );
NAND2_X2 _AES_ENC_us22_U380  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n703 ), .ZN(_AES_ENC_us22_n732 ) );
AND2_X2 _AES_ENC_us22_U379  ( .A1(_AES_ENC_sa22[0]), .A2(_AES_ENC_sa22[6]),.ZN(_AES_ENC_us22_n1113 ) );
NAND2_X2 _AES_ENC_us22_U378  ( .A1(_AES_ENC_us22_n601 ), .A2(_AES_ENC_us22_n1030 ), .ZN(_AES_ENC_us22_n881 ) );
NAND2_X2 _AES_ENC_us22_U377  ( .A1(_AES_ENC_us22_n1093 ), .A2(_AES_ENC_us22_n881 ), .ZN(_AES_ENC_us22_n715 ) );
NAND2_X2 _AES_ENC_us22_U376  ( .A1(_AES_ENC_us22_n1010 ), .A2(_AES_ENC_us22_n600 ), .ZN(_AES_ENC_us22_n714 ) );
NAND2_X2 _AES_ENC_us22_U375  ( .A1(_AES_ENC_us22_n855 ), .A2(_AES_ENC_us22_n588 ), .ZN(_AES_ENC_us22_n1117 ) );
XNOR2_X2 _AES_ENC_us22_U371  ( .A(_AES_ENC_us22_n611 ), .B(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n824 ) );
NAND4_X2 _AES_ENC_us22_U362  ( .A1(_AES_ENC_us22_n715 ), .A2(_AES_ENC_us22_n714 ), .A3(_AES_ENC_us22_n713 ), .A4(_AES_ENC_us22_n712 ), .ZN(_AES_ENC_us22_n716 ) );
NAND2_X2 _AES_ENC_us22_U361  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n716 ), .ZN(_AES_ENC_us22_n731 ) );
AND2_X2 _AES_ENC_us22_U360  ( .A1(_AES_ENC_sa22[6]), .A2(_AES_ENC_us22_n574 ), .ZN(_AES_ENC_us22_n1131 ) );
NAND2_X2 _AES_ENC_us22_U359  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n717 ) );
NAND2_X2 _AES_ENC_us22_U358  ( .A1(_AES_ENC_us22_n1029 ), .A2(_AES_ENC_us22_n717 ), .ZN(_AES_ENC_us22_n728 ) );
NAND2_X2 _AES_ENC_us22_U357  ( .A1(_AES_ENC_sa22[1]), .A2(_AES_ENC_us22_n624 ), .ZN(_AES_ENC_us22_n1097 ) );
NAND2_X2 _AES_ENC_us22_U356  ( .A1(_AES_ENC_us22_n603 ), .A2(_AES_ENC_us22_n1097 ), .ZN(_AES_ENC_us22_n718 ) );
NAND2_X2 _AES_ENC_us22_U355  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n718 ), .ZN(_AES_ENC_us22_n727 ) );
NAND4_X2 _AES_ENC_us22_U344  ( .A1(_AES_ENC_us22_n728 ), .A2(_AES_ENC_us22_n727 ), .A3(_AES_ENC_us22_n726 ), .A4(_AES_ENC_us22_n725 ), .ZN(_AES_ENC_us22_n729 ) );
NAND2_X2 _AES_ENC_us22_U343  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n729 ), .ZN(_AES_ENC_us22_n730 ) );
NAND4_X2 _AES_ENC_us22_U342  ( .A1(_AES_ENC_us22_n733 ), .A2(_AES_ENC_us22_n732 ), .A3(_AES_ENC_us22_n731 ), .A4(_AES_ENC_us22_n730 ), .ZN(_AES_ENC_sa22_sub[1] ) );
NAND2_X2 _AES_ENC_us22_U341  ( .A1(_AES_ENC_sa22[7]), .A2(_AES_ENC_us22_n611 ), .ZN(_AES_ENC_us22_n734 ) );
NAND2_X2 _AES_ENC_us22_U340  ( .A1(_AES_ENC_us22_n734 ), .A2(_AES_ENC_us22_n607 ), .ZN(_AES_ENC_us22_n738 ) );
OR4_X2 _AES_ENC_us22_U339  ( .A1(_AES_ENC_us22_n738 ), .A2(_AES_ENC_us22_n626 ), .A3(_AES_ENC_us22_n826 ), .A4(_AES_ENC_us22_n1121 ), .ZN(_AES_ENC_us22_n746 ) );
NAND2_X2 _AES_ENC_us22_U337  ( .A1(_AES_ENC_us22_n1100 ), .A2(_AES_ENC_us22_n587 ), .ZN(_AES_ENC_us22_n992 ) );
OR2_X2 _AES_ENC_us22_U336  ( .A1(_AES_ENC_us22_n610 ), .A2(_AES_ENC_us22_n735 ), .ZN(_AES_ENC_us22_n737 ) );
NAND2_X2 _AES_ENC_us22_U334  ( .A1(_AES_ENC_us22_n619 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n753 ) );
NAND2_X2 _AES_ENC_us22_U333  ( .A1(_AES_ENC_us22_n582 ), .A2(_AES_ENC_us22_n753 ), .ZN(_AES_ENC_us22_n1080 ) );
NAND2_X2 _AES_ENC_us22_U332  ( .A1(_AES_ENC_us22_n1048 ), .A2(_AES_ENC_us22_n576 ), .ZN(_AES_ENC_us22_n736 ) );
NAND2_X2 _AES_ENC_us22_U331  ( .A1(_AES_ENC_us22_n737 ), .A2(_AES_ENC_us22_n736 ), .ZN(_AES_ENC_us22_n739 ) );
NAND2_X2 _AES_ENC_us22_U330  ( .A1(_AES_ENC_us22_n739 ), .A2(_AES_ENC_us22_n738 ), .ZN(_AES_ENC_us22_n745 ) );
NAND2_X2 _AES_ENC_us22_U326  ( .A1(_AES_ENC_us22_n1096 ), .A2(_AES_ENC_us22_n590 ), .ZN(_AES_ENC_us22_n906 ) );
NAND4_X2 _AES_ENC_us22_U323  ( .A1(_AES_ENC_us22_n746 ), .A2(_AES_ENC_us22_n992 ), .A3(_AES_ENC_us22_n745 ), .A4(_AES_ENC_us22_n744 ), .ZN(_AES_ENC_us22_n747 ) );
NAND2_X2 _AES_ENC_us22_U322  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n747 ), .ZN(_AES_ENC_us22_n793 ) );
NAND2_X2 _AES_ENC_us22_U321  ( .A1(_AES_ENC_us22_n584 ), .A2(_AES_ENC_us22_n855 ), .ZN(_AES_ENC_us22_n748 ) );
NAND2_X2 _AES_ENC_us22_U320  ( .A1(_AES_ENC_us22_n956 ), .A2(_AES_ENC_us22_n748 ), .ZN(_AES_ENC_us22_n760 ) );
NAND2_X2 _AES_ENC_us22_U313  ( .A1(_AES_ENC_us22_n590 ), .A2(_AES_ENC_us22_n753 ), .ZN(_AES_ENC_us22_n1023 ) );
NAND4_X2 _AES_ENC_us22_U308  ( .A1(_AES_ENC_us22_n760 ), .A2(_AES_ENC_us22_n992 ), .A3(_AES_ENC_us22_n759 ), .A4(_AES_ENC_us22_n758 ), .ZN(_AES_ENC_us22_n761 ) );
NAND2_X2 _AES_ENC_us22_U307  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n761 ), .ZN(_AES_ENC_us22_n792 ) );
NAND2_X2 _AES_ENC_us22_U306  ( .A1(_AES_ENC_us22_n584 ), .A2(_AES_ENC_us22_n603 ), .ZN(_AES_ENC_us22_n989 ) );
NAND2_X2 _AES_ENC_us22_U305  ( .A1(_AES_ENC_us22_n1050 ), .A2(_AES_ENC_us22_n989 ), .ZN(_AES_ENC_us22_n777 ) );
NAND2_X2 _AES_ENC_us22_U304  ( .A1(_AES_ENC_us22_n1093 ), .A2(_AES_ENC_us22_n762 ), .ZN(_AES_ENC_us22_n776 ) );
XNOR2_X2 _AES_ENC_us22_U301  ( .A(_AES_ENC_sa22[7]), .B(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n959 ) );
NAND4_X2 _AES_ENC_us22_U289  ( .A1(_AES_ENC_us22_n777 ), .A2(_AES_ENC_us22_n776 ), .A3(_AES_ENC_us22_n775 ), .A4(_AES_ENC_us22_n774 ), .ZN(_AES_ENC_us22_n778 ) );
NAND2_X2 _AES_ENC_us22_U288  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n778 ), .ZN(_AES_ENC_us22_n791 ) );
NAND2_X2 _AES_ENC_us22_U287  ( .A1(_AES_ENC_us22_n1056 ), .A2(_AES_ENC_us22_n1050 ), .ZN(_AES_ENC_us22_n788 ) );
NAND2_X2 _AES_ENC_us22_U286  ( .A1(_AES_ENC_us22_n1091 ), .A2(_AES_ENC_us22_n779 ), .ZN(_AES_ENC_us22_n787 ) );
NAND2_X2 _AES_ENC_us22_U285  ( .A1(_AES_ENC_us22_n956 ), .A2(_AES_ENC_sa22[1]), .ZN(_AES_ENC_us22_n786 ) );
NAND4_X2 _AES_ENC_us22_U278  ( .A1(_AES_ENC_us22_n788 ), .A2(_AES_ENC_us22_n787 ), .A3(_AES_ENC_us22_n786 ), .A4(_AES_ENC_us22_n785 ), .ZN(_AES_ENC_us22_n789 ) );
NAND2_X2 _AES_ENC_us22_U277  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n789 ), .ZN(_AES_ENC_us22_n790 ) );
NAND4_X2 _AES_ENC_us22_U276  ( .A1(_AES_ENC_us22_n793 ), .A2(_AES_ENC_us22_n792 ), .A3(_AES_ENC_us22_n791 ), .A4(_AES_ENC_us22_n790 ), .ZN(_AES_ENC_sa22_sub[2] ) );
NAND2_X2 _AES_ENC_us22_U275  ( .A1(_AES_ENC_us22_n1059 ), .A2(_AES_ENC_us22_n794 ), .ZN(_AES_ENC_us22_n810 ) );
NAND2_X2 _AES_ENC_us22_U274  ( .A1(_AES_ENC_us22_n1049 ), .A2(_AES_ENC_us22_n956 ), .ZN(_AES_ENC_us22_n809 ) );
OR2_X2 _AES_ENC_us22_U266  ( .A1(_AES_ENC_us22_n1096 ), .A2(_AES_ENC_us22_n606 ), .ZN(_AES_ENC_us22_n802 ) );
NAND2_X2 _AES_ENC_us22_U265  ( .A1(_AES_ENC_us22_n1053 ), .A2(_AES_ENC_us22_n800 ), .ZN(_AES_ENC_us22_n801 ) );
NAND2_X2 _AES_ENC_us22_U264  ( .A1(_AES_ENC_us22_n802 ), .A2(_AES_ENC_us22_n801 ), .ZN(_AES_ENC_us22_n805 ) );
NAND4_X2 _AES_ENC_us22_U261  ( .A1(_AES_ENC_us22_n810 ), .A2(_AES_ENC_us22_n809 ), .A3(_AES_ENC_us22_n808 ), .A4(_AES_ENC_us22_n807 ), .ZN(_AES_ENC_us22_n811 ) );
NAND2_X2 _AES_ENC_us22_U260  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n811 ), .ZN(_AES_ENC_us22_n852 ) );
OR2_X2 _AES_ENC_us22_U259  ( .A1(_AES_ENC_us22_n1023 ), .A2(_AES_ENC_us22_n617 ), .ZN(_AES_ENC_us22_n819 ) );
OR2_X2 _AES_ENC_us22_U257  ( .A1(_AES_ENC_us22_n570 ), .A2(_AES_ENC_us22_n930 ), .ZN(_AES_ENC_us22_n818 ) );
NAND2_X2 _AES_ENC_us22_U256  ( .A1(_AES_ENC_us22_n1013 ), .A2(_AES_ENC_us22_n1094 ), .ZN(_AES_ENC_us22_n817 ) );
NAND4_X2 _AES_ENC_us22_U249  ( .A1(_AES_ENC_us22_n819 ), .A2(_AES_ENC_us22_n818 ), .A3(_AES_ENC_us22_n817 ), .A4(_AES_ENC_us22_n816 ), .ZN(_AES_ENC_us22_n820 ) );
NAND2_X2 _AES_ENC_us22_U248  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n820 ), .ZN(_AES_ENC_us22_n851 ) );
NAND2_X2 _AES_ENC_us22_U247  ( .A1(_AES_ENC_us22_n956 ), .A2(_AES_ENC_us22_n1080 ), .ZN(_AES_ENC_us22_n835 ) );
NAND2_X2 _AES_ENC_us22_U246  ( .A1(_AES_ENC_us22_n570 ), .A2(_AES_ENC_us22_n1030 ), .ZN(_AES_ENC_us22_n1047 ) );
OR2_X2 _AES_ENC_us22_U245  ( .A1(_AES_ENC_us22_n1047 ), .A2(_AES_ENC_us22_n612 ), .ZN(_AES_ENC_us22_n834 ) );
NAND2_X2 _AES_ENC_us22_U244  ( .A1(_AES_ENC_us22_n1072 ), .A2(_AES_ENC_us22_n589 ), .ZN(_AES_ENC_us22_n833 ) );
NAND4_X2 _AES_ENC_us22_U233  ( .A1(_AES_ENC_us22_n835 ), .A2(_AES_ENC_us22_n834 ), .A3(_AES_ENC_us22_n833 ), .A4(_AES_ENC_us22_n832 ), .ZN(_AES_ENC_us22_n836 ) );
NAND2_X2 _AES_ENC_us22_U232  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n836 ), .ZN(_AES_ENC_us22_n850 ) );
NAND2_X2 _AES_ENC_us22_U231  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n623 ), .ZN(_AES_ENC_us22_n847 ) );
NAND2_X2 _AES_ENC_us22_U230  ( .A1(_AES_ENC_us22_n1050 ), .A2(_AES_ENC_us22_n1071 ), .ZN(_AES_ENC_us22_n846 ) );
OR2_X2 _AES_ENC_us22_U224  ( .A1(_AES_ENC_us22_n1053 ), .A2(_AES_ENC_us22_n911 ), .ZN(_AES_ENC_us22_n1077 ) );
NAND4_X2 _AES_ENC_us22_U220  ( .A1(_AES_ENC_us22_n847 ), .A2(_AES_ENC_us22_n846 ), .A3(_AES_ENC_us22_n845 ), .A4(_AES_ENC_us22_n844 ), .ZN(_AES_ENC_us22_n848 ) );
NAND2_X2 _AES_ENC_us22_U219  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n848 ), .ZN(_AES_ENC_us22_n849 ) );
NAND4_X2 _AES_ENC_us22_U218  ( .A1(_AES_ENC_us22_n852 ), .A2(_AES_ENC_us22_n851 ), .A3(_AES_ENC_us22_n850 ), .A4(_AES_ENC_us22_n849 ), .ZN(_AES_ENC_sa22_sub[3] ) );
NAND2_X2 _AES_ENC_us22_U216  ( .A1(_AES_ENC_us22_n1009 ), .A2(_AES_ENC_us22_n1072 ), .ZN(_AES_ENC_us22_n862 ) );
NAND2_X2 _AES_ENC_us22_U215  ( .A1(_AES_ENC_us22_n603 ), .A2(_AES_ENC_us22_n577 ), .ZN(_AES_ENC_us22_n853 ) );
NAND2_X2 _AES_ENC_us22_U214  ( .A1(_AES_ENC_us22_n1050 ), .A2(_AES_ENC_us22_n853 ), .ZN(_AES_ENC_us22_n861 ) );
NAND4_X2 _AES_ENC_us22_U206  ( .A1(_AES_ENC_us22_n862 ), .A2(_AES_ENC_us22_n861 ), .A3(_AES_ENC_us22_n860 ), .A4(_AES_ENC_us22_n859 ), .ZN(_AES_ENC_us22_n863 ) );
NAND2_X2 _AES_ENC_us22_U205  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n863 ), .ZN(_AES_ENC_us22_n905 ) );
NAND2_X2 _AES_ENC_us22_U204  ( .A1(_AES_ENC_us22_n1010 ), .A2(_AES_ENC_us22_n989 ), .ZN(_AES_ENC_us22_n874 ) );
NAND2_X2 _AES_ENC_us22_U203  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n610 ), .ZN(_AES_ENC_us22_n864 ) );
NAND2_X2 _AES_ENC_us22_U202  ( .A1(_AES_ENC_us22_n929 ), .A2(_AES_ENC_us22_n864 ), .ZN(_AES_ENC_us22_n873 ) );
NAND4_X2 _AES_ENC_us22_U193  ( .A1(_AES_ENC_us22_n874 ), .A2(_AES_ENC_us22_n873 ), .A3(_AES_ENC_us22_n872 ), .A4(_AES_ENC_us22_n871 ), .ZN(_AES_ENC_us22_n875 ) );
NAND2_X2 _AES_ENC_us22_U192  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n875 ), .ZN(_AES_ENC_us22_n904 ) );
NAND2_X2 _AES_ENC_us22_U191  ( .A1(_AES_ENC_us22_n583 ), .A2(_AES_ENC_us22_n1050 ), .ZN(_AES_ENC_us22_n889 ) );
NAND2_X2 _AES_ENC_us22_U190  ( .A1(_AES_ENC_us22_n1093 ), .A2(_AES_ENC_us22_n587 ), .ZN(_AES_ENC_us22_n876 ) );
NAND2_X2 _AES_ENC_us22_U189  ( .A1(_AES_ENC_us22_n604 ), .A2(_AES_ENC_us22_n876 ), .ZN(_AES_ENC_us22_n877 ) );
NAND2_X2 _AES_ENC_us22_U188  ( .A1(_AES_ENC_us22_n877 ), .A2(_AES_ENC_us22_n623 ), .ZN(_AES_ENC_us22_n888 ) );
NAND4_X2 _AES_ENC_us22_U179  ( .A1(_AES_ENC_us22_n889 ), .A2(_AES_ENC_us22_n888 ), .A3(_AES_ENC_us22_n887 ), .A4(_AES_ENC_us22_n886 ), .ZN(_AES_ENC_us22_n890 ) );
NAND2_X2 _AES_ENC_us22_U178  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n890 ), .ZN(_AES_ENC_us22_n903 ) );
OR2_X2 _AES_ENC_us22_U177  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n1059 ), .ZN(_AES_ENC_us22_n900 ) );
NAND2_X2 _AES_ENC_us22_U176  ( .A1(_AES_ENC_us22_n1073 ), .A2(_AES_ENC_us22_n1047 ), .ZN(_AES_ENC_us22_n899 ) );
NAND2_X2 _AES_ENC_us22_U175  ( .A1(_AES_ENC_us22_n1094 ), .A2(_AES_ENC_us22_n595 ), .ZN(_AES_ENC_us22_n898 ) );
NAND4_X2 _AES_ENC_us22_U167  ( .A1(_AES_ENC_us22_n900 ), .A2(_AES_ENC_us22_n899 ), .A3(_AES_ENC_us22_n898 ), .A4(_AES_ENC_us22_n897 ), .ZN(_AES_ENC_us22_n901 ) );
NAND2_X2 _AES_ENC_us22_U166  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n901 ), .ZN(_AES_ENC_us22_n902 ) );
NAND4_X2 _AES_ENC_us22_U165  ( .A1(_AES_ENC_us22_n905 ), .A2(_AES_ENC_us22_n904 ), .A3(_AES_ENC_us22_n903 ), .A4(_AES_ENC_us22_n902 ), .ZN(_AES_ENC_sa22_sub[4] ) );
NAND2_X2 _AES_ENC_us22_U164  ( .A1(_AES_ENC_us22_n1094 ), .A2(_AES_ENC_us22_n599 ), .ZN(_AES_ENC_us22_n922 ) );
NAND2_X2 _AES_ENC_us22_U163  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n989 ), .ZN(_AES_ENC_us22_n921 ) );
NAND4_X2 _AES_ENC_us22_U151  ( .A1(_AES_ENC_us22_n922 ), .A2(_AES_ENC_us22_n921 ), .A3(_AES_ENC_us22_n920 ), .A4(_AES_ENC_us22_n919 ), .ZN(_AES_ENC_us22_n923 ) );
NAND2_X2 _AES_ENC_us22_U150  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n923 ), .ZN(_AES_ENC_us22_n972 ) );
NAND2_X2 _AES_ENC_us22_U149  ( .A1(_AES_ENC_us22_n582 ), .A2(_AES_ENC_us22_n619 ), .ZN(_AES_ENC_us22_n924 ) );
NAND2_X2 _AES_ENC_us22_U148  ( .A1(_AES_ENC_us22_n1073 ), .A2(_AES_ENC_us22_n924 ), .ZN(_AES_ENC_us22_n939 ) );
NAND2_X2 _AES_ENC_us22_U147  ( .A1(_AES_ENC_us22_n926 ), .A2(_AES_ENC_us22_n925 ), .ZN(_AES_ENC_us22_n927 ) );
NAND2_X2 _AES_ENC_us22_U146  ( .A1(_AES_ENC_us22_n606 ), .A2(_AES_ENC_us22_n927 ), .ZN(_AES_ENC_us22_n928 ) );
NAND2_X2 _AES_ENC_us22_U145  ( .A1(_AES_ENC_us22_n928 ), .A2(_AES_ENC_us22_n1080 ), .ZN(_AES_ENC_us22_n938 ) );
OR2_X2 _AES_ENC_us22_U144  ( .A1(_AES_ENC_us22_n1117 ), .A2(_AES_ENC_us22_n615 ), .ZN(_AES_ENC_us22_n937 ) );
NAND4_X2 _AES_ENC_us22_U139  ( .A1(_AES_ENC_us22_n939 ), .A2(_AES_ENC_us22_n938 ), .A3(_AES_ENC_us22_n937 ), .A4(_AES_ENC_us22_n936 ), .ZN(_AES_ENC_us22_n940 ) );
NAND2_X2 _AES_ENC_us22_U138  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n940 ), .ZN(_AES_ENC_us22_n971 ) );
OR2_X2 _AES_ENC_us22_U137  ( .A1(_AES_ENC_us22_n605 ), .A2(_AES_ENC_us22_n941 ), .ZN(_AES_ENC_us22_n954 ) );
NAND2_X2 _AES_ENC_us22_U136  ( .A1(_AES_ENC_us22_n1096 ), .A2(_AES_ENC_us22_n577 ), .ZN(_AES_ENC_us22_n942 ) );
NAND2_X2 _AES_ENC_us22_U135  ( .A1(_AES_ENC_us22_n1048 ), .A2(_AES_ENC_us22_n942 ), .ZN(_AES_ENC_us22_n943 ) );
NAND2_X2 _AES_ENC_us22_U134  ( .A1(_AES_ENC_us22_n612 ), .A2(_AES_ENC_us22_n943 ), .ZN(_AES_ENC_us22_n944 ) );
NAND2_X2 _AES_ENC_us22_U133  ( .A1(_AES_ENC_us22_n944 ), .A2(_AES_ENC_us22_n580 ), .ZN(_AES_ENC_us22_n953 ) );
NAND4_X2 _AES_ENC_us22_U125  ( .A1(_AES_ENC_us22_n954 ), .A2(_AES_ENC_us22_n953 ), .A3(_AES_ENC_us22_n952 ), .A4(_AES_ENC_us22_n951 ), .ZN(_AES_ENC_us22_n955 ) );
NAND2_X2 _AES_ENC_us22_U124  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n955 ), .ZN(_AES_ENC_us22_n970 ) );
NAND2_X2 _AES_ENC_us22_U123  ( .A1(_AES_ENC_us22_n1094 ), .A2(_AES_ENC_us22_n1071 ), .ZN(_AES_ENC_us22_n967 ) );
NAND2_X2 _AES_ENC_us22_U122  ( .A1(_AES_ENC_us22_n956 ), .A2(_AES_ENC_us22_n1030 ), .ZN(_AES_ENC_us22_n966 ) );
NAND4_X2 _AES_ENC_us22_U114  ( .A1(_AES_ENC_us22_n967 ), .A2(_AES_ENC_us22_n966 ), .A3(_AES_ENC_us22_n965 ), .A4(_AES_ENC_us22_n964 ), .ZN(_AES_ENC_us22_n968 ) );
NAND2_X2 _AES_ENC_us22_U113  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n968 ), .ZN(_AES_ENC_us22_n969 ) );
NAND4_X2 _AES_ENC_us22_U112  ( .A1(_AES_ENC_us22_n972 ), .A2(_AES_ENC_us22_n971 ), .A3(_AES_ENC_us22_n970 ), .A4(_AES_ENC_us22_n969 ), .ZN(_AES_ENC_sa22_sub[5] ) );
NAND2_X2 _AES_ENC_us22_U111  ( .A1(_AES_ENC_us22_n570 ), .A2(_AES_ENC_us22_n1097 ), .ZN(_AES_ENC_us22_n973 ) );
NAND2_X2 _AES_ENC_us22_U110  ( .A1(_AES_ENC_us22_n1073 ), .A2(_AES_ENC_us22_n973 ), .ZN(_AES_ENC_us22_n987 ) );
NAND2_X2 _AES_ENC_us22_U109  ( .A1(_AES_ENC_us22_n974 ), .A2(_AES_ENC_us22_n1077 ), .ZN(_AES_ENC_us22_n975 ) );
NAND2_X2 _AES_ENC_us22_U108  ( .A1(_AES_ENC_us22_n613 ), .A2(_AES_ENC_us22_n975 ), .ZN(_AES_ENC_us22_n976 ) );
NAND2_X2 _AES_ENC_us22_U107  ( .A1(_AES_ENC_us22_n977 ), .A2(_AES_ENC_us22_n976 ), .ZN(_AES_ENC_us22_n986 ) );
NAND4_X2 _AES_ENC_us22_U99  ( .A1(_AES_ENC_us22_n987 ), .A2(_AES_ENC_us22_n986 ), .A3(_AES_ENC_us22_n985 ), .A4(_AES_ENC_us22_n984 ), .ZN(_AES_ENC_us22_n988 ) );
NAND2_X2 _AES_ENC_us22_U98  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n988 ), .ZN(_AES_ENC_us22_n1044 ) );
NAND2_X2 _AES_ENC_us22_U97  ( .A1(_AES_ENC_us22_n1073 ), .A2(_AES_ENC_us22_n989 ), .ZN(_AES_ENC_us22_n1004 ) );
NAND2_X2 _AES_ENC_us22_U96  ( .A1(_AES_ENC_us22_n1092 ), .A2(_AES_ENC_us22_n619 ), .ZN(_AES_ENC_us22_n1003 ) );
NAND4_X2 _AES_ENC_us22_U85  ( .A1(_AES_ENC_us22_n1004 ), .A2(_AES_ENC_us22_n1003 ), .A3(_AES_ENC_us22_n1002 ), .A4(_AES_ENC_us22_n1001 ), .ZN(_AES_ENC_us22_n1005 ) );
NAND2_X2 _AES_ENC_us22_U84  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n1005 ), .ZN(_AES_ENC_us22_n1043 ) );
NAND2_X2 _AES_ENC_us22_U83  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n596 ), .ZN(_AES_ENC_us22_n1020 ) );
NAND2_X2 _AES_ENC_us22_U82  ( .A1(_AES_ENC_us22_n1050 ), .A2(_AES_ENC_us22_n624 ), .ZN(_AES_ENC_us22_n1019 ) );
NAND2_X2 _AES_ENC_us22_U77  ( .A1(_AES_ENC_us22_n1059 ), .A2(_AES_ENC_us22_n1114 ), .ZN(_AES_ENC_us22_n1012 ) );
NAND2_X2 _AES_ENC_us22_U76  ( .A1(_AES_ENC_us22_n1010 ), .A2(_AES_ENC_us22_n592 ), .ZN(_AES_ENC_us22_n1011 ) );
NAND2_X2 _AES_ENC_us22_U75  ( .A1(_AES_ENC_us22_n1012 ), .A2(_AES_ENC_us22_n1011 ), .ZN(_AES_ENC_us22_n1016 ) );
NAND4_X2 _AES_ENC_us22_U70  ( .A1(_AES_ENC_us22_n1020 ), .A2(_AES_ENC_us22_n1019 ), .A3(_AES_ENC_us22_n1018 ), .A4(_AES_ENC_us22_n1017 ), .ZN(_AES_ENC_us22_n1021 ) );
NAND2_X2 _AES_ENC_us22_U69  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n1021 ), .ZN(_AES_ENC_us22_n1042 ) );
NAND2_X2 _AES_ENC_us22_U68  ( .A1(_AES_ENC_us22_n1022 ), .A2(_AES_ENC_us22_n1093 ), .ZN(_AES_ENC_us22_n1039 ) );
NAND2_X2 _AES_ENC_us22_U67  ( .A1(_AES_ENC_us22_n1050 ), .A2(_AES_ENC_us22_n1023 ), .ZN(_AES_ENC_us22_n1038 ) );
NAND2_X2 _AES_ENC_us22_U66  ( .A1(_AES_ENC_us22_n1024 ), .A2(_AES_ENC_us22_n1071 ), .ZN(_AES_ENC_us22_n1037 ) );
AND2_X2 _AES_ENC_us22_U60  ( .A1(_AES_ENC_us22_n1030 ), .A2(_AES_ENC_us22_n602 ), .ZN(_AES_ENC_us22_n1078 ) );
NAND4_X2 _AES_ENC_us22_U56  ( .A1(_AES_ENC_us22_n1039 ), .A2(_AES_ENC_us22_n1038 ), .A3(_AES_ENC_us22_n1037 ), .A4(_AES_ENC_us22_n1036 ), .ZN(_AES_ENC_us22_n1040 ) );
NAND2_X2 _AES_ENC_us22_U55  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n1040 ), .ZN(_AES_ENC_us22_n1041 ) );
NAND4_X2 _AES_ENC_us22_U54  ( .A1(_AES_ENC_us22_n1044 ), .A2(_AES_ENC_us22_n1043 ), .A3(_AES_ENC_us22_n1042 ), .A4(_AES_ENC_us22_n1041 ), .ZN(_AES_ENC_sa22_sub[6] ) );
NAND2_X2 _AES_ENC_us22_U53  ( .A1(_AES_ENC_us22_n1072 ), .A2(_AES_ENC_us22_n1045 ), .ZN(_AES_ENC_us22_n1068 ) );
NAND2_X2 _AES_ENC_us22_U52  ( .A1(_AES_ENC_us22_n1046 ), .A2(_AES_ENC_us22_n582 ), .ZN(_AES_ENC_us22_n1067 ) );
NAND2_X2 _AES_ENC_us22_U51  ( .A1(_AES_ENC_us22_n1094 ), .A2(_AES_ENC_us22_n1047 ), .ZN(_AES_ENC_us22_n1066 ) );
NAND4_X2 _AES_ENC_us22_U40  ( .A1(_AES_ENC_us22_n1068 ), .A2(_AES_ENC_us22_n1067 ), .A3(_AES_ENC_us22_n1066 ), .A4(_AES_ENC_us22_n1065 ), .ZN(_AES_ENC_us22_n1069 ) );
NAND2_X2 _AES_ENC_us22_U39  ( .A1(_AES_ENC_us22_n1070 ), .A2(_AES_ENC_us22_n1069 ), .ZN(_AES_ENC_us22_n1135 ) );
NAND2_X2 _AES_ENC_us22_U38  ( .A1(_AES_ENC_us22_n1072 ), .A2(_AES_ENC_us22_n1071 ), .ZN(_AES_ENC_us22_n1088 ) );
NAND2_X2 _AES_ENC_us22_U37  ( .A1(_AES_ENC_us22_n1073 ), .A2(_AES_ENC_us22_n595 ), .ZN(_AES_ENC_us22_n1087 ) );
NAND4_X2 _AES_ENC_us22_U28  ( .A1(_AES_ENC_us22_n1088 ), .A2(_AES_ENC_us22_n1087 ), .A3(_AES_ENC_us22_n1086 ), .A4(_AES_ENC_us22_n1085 ), .ZN(_AES_ENC_us22_n1089 ) );
NAND2_X2 _AES_ENC_us22_U27  ( .A1(_AES_ENC_us22_n1090 ), .A2(_AES_ENC_us22_n1089 ), .ZN(_AES_ENC_us22_n1134 ) );
NAND2_X2 _AES_ENC_us22_U26  ( .A1(_AES_ENC_us22_n1091 ), .A2(_AES_ENC_us22_n1093 ), .ZN(_AES_ENC_us22_n1111 ) );
NAND2_X2 _AES_ENC_us22_U25  ( .A1(_AES_ENC_us22_n1092 ), .A2(_AES_ENC_us22_n1120 ), .ZN(_AES_ENC_us22_n1110 ) );
AND2_X2 _AES_ENC_us22_U22  ( .A1(_AES_ENC_us22_n1097 ), .A2(_AES_ENC_us22_n1096 ), .ZN(_AES_ENC_us22_n1098 ) );
NAND4_X2 _AES_ENC_us22_U14  ( .A1(_AES_ENC_us22_n1111 ), .A2(_AES_ENC_us22_n1110 ), .A3(_AES_ENC_us22_n1109 ), .A4(_AES_ENC_us22_n1108 ), .ZN(_AES_ENC_us22_n1112 ) );
NAND2_X2 _AES_ENC_us22_U13  ( .A1(_AES_ENC_us22_n1113 ), .A2(_AES_ENC_us22_n1112 ), .ZN(_AES_ENC_us22_n1133 ) );
NAND2_X2 _AES_ENC_us22_U12  ( .A1(_AES_ENC_us22_n1115 ), .A2(_AES_ENC_us22_n1114 ), .ZN(_AES_ENC_us22_n1129 ) );
OR2_X2 _AES_ENC_us22_U11  ( .A1(_AES_ENC_us22_n608 ), .A2(_AES_ENC_us22_n1116 ), .ZN(_AES_ENC_us22_n1128 ) );
NAND4_X2 _AES_ENC_us22_U3  ( .A1(_AES_ENC_us22_n1129 ), .A2(_AES_ENC_us22_n1128 ), .A3(_AES_ENC_us22_n1127 ), .A4(_AES_ENC_us22_n1126 ), .ZN(_AES_ENC_us22_n1130 ) );
NAND2_X2 _AES_ENC_us22_U2  ( .A1(_AES_ENC_us22_n1131 ), .A2(_AES_ENC_us22_n1130 ), .ZN(_AES_ENC_us22_n1132 ) );
NAND4_X2 _AES_ENC_us22_U1  ( .A1(_AES_ENC_us22_n1135 ), .A2(_AES_ENC_us22_n1134 ), .A3(_AES_ENC_us22_n1133 ), .A4(_AES_ENC_us22_n1132 ), .ZN(_AES_ENC_sa22_sub[7] ) );
INV_X4 _AES_ENC_us23_U575  ( .A(_AES_ENC_sa23[0]), .ZN(_AES_ENC_us23_n627 ));
INV_X4 _AES_ENC_us23_U574  ( .A(_AES_ENC_us23_n1053 ), .ZN(_AES_ENC_us23_n625 ) );
INV_X4 _AES_ENC_us23_U573  ( .A(_AES_ENC_us23_n1103 ), .ZN(_AES_ENC_us23_n623 ) );
INV_X4 _AES_ENC_us23_U572  ( .A(_AES_ENC_us23_n1056 ), .ZN(_AES_ENC_us23_n622 ) );
INV_X4 _AES_ENC_us23_U571  ( .A(_AES_ENC_us23_n1102 ), .ZN(_AES_ENC_us23_n621 ) );
INV_X4 _AES_ENC_us23_U570  ( .A(_AES_ENC_us23_n1074 ), .ZN(_AES_ENC_us23_n620 ) );
INV_X4 _AES_ENC_us23_U569  ( .A(_AES_ENC_us23_n929 ), .ZN(_AES_ENC_us23_n619 ) );
INV_X4 _AES_ENC_us23_U568  ( .A(_AES_ENC_us23_n1091 ), .ZN(_AES_ENC_us23_n618 ) );
INV_X4 _AES_ENC_us23_U567  ( .A(_AES_ENC_us23_n826 ), .ZN(_AES_ENC_us23_n617 ) );
INV_X4 _AES_ENC_us23_U566  ( .A(_AES_ENC_us23_n1031 ), .ZN(_AES_ENC_us23_n616 ) );
INV_X4 _AES_ENC_us23_U565  ( .A(_AES_ENC_us23_n1054 ), .ZN(_AES_ENC_us23_n615 ) );
INV_X4 _AES_ENC_us23_U564  ( .A(_AES_ENC_us23_n1025 ), .ZN(_AES_ENC_us23_n614 ) );
INV_X4 _AES_ENC_us23_U563  ( .A(_AES_ENC_us23_n990 ), .ZN(_AES_ENC_us23_n613 ) );
INV_X4 _AES_ENC_us23_U562  ( .A(_AES_ENC_sa23[4]), .ZN(_AES_ENC_us23_n612 ));
INV_X4 _AES_ENC_us23_U561  ( .A(_AES_ENC_us23_n881 ), .ZN(_AES_ENC_us23_n611 ) );
INV_X4 _AES_ENC_us23_U560  ( .A(_AES_ENC_us23_n1022 ), .ZN(_AES_ENC_us23_n610 ) );
INV_X4 _AES_ENC_us23_U559  ( .A(_AES_ENC_us23_n1120 ), .ZN(_AES_ENC_us23_n609 ) );
INV_X4 _AES_ENC_us23_U558  ( .A(_AES_ENC_us23_n977 ), .ZN(_AES_ENC_us23_n608 ) );
INV_X4 _AES_ENC_us23_U557  ( .A(_AES_ENC_us23_n926 ), .ZN(_AES_ENC_us23_n607 ) );
INV_X4 _AES_ENC_us23_U556  ( .A(_AES_ENC_us23_n910 ), .ZN(_AES_ENC_us23_n606 ) );
INV_X4 _AES_ENC_us23_U555  ( .A(_AES_ENC_us23_n1121 ), .ZN(_AES_ENC_us23_n605 ) );
INV_X4 _AES_ENC_us23_U554  ( .A(_AES_ENC_us23_n1009 ), .ZN(_AES_ENC_us23_n604 ) );
INV_X4 _AES_ENC_us23_U553  ( .A(_AES_ENC_us23_n1080 ), .ZN(_AES_ENC_us23_n602 ) );
INV_X4 _AES_ENC_us23_U552  ( .A(_AES_ENC_us23_n821 ), .ZN(_AES_ENC_us23_n600 ) );
INV_X4 _AES_ENC_us23_U551  ( .A(_AES_ENC_us23_n1013 ), .ZN(_AES_ENC_us23_n599 ) );
INV_X4 _AES_ENC_us23_U550  ( .A(_AES_ENC_us23_n1058 ), .ZN(_AES_ENC_us23_n598 ) );
INV_X4 _AES_ENC_us23_U549  ( .A(_AES_ENC_us23_n906 ), .ZN(_AES_ENC_us23_n597 ) );
INV_X4 _AES_ENC_us23_U548  ( .A(_AES_ENC_us23_n1048 ), .ZN(_AES_ENC_us23_n595 ) );
INV_X4 _AES_ENC_us23_U547  ( .A(_AES_ENC_us23_n974 ), .ZN(_AES_ENC_us23_n594 ) );
INV_X4 _AES_ENC_us23_U546  ( .A(_AES_ENC_sa23[2]), .ZN(_AES_ENC_us23_n593 ));
INV_X4 _AES_ENC_us23_U545  ( .A(_AES_ENC_us23_n800 ), .ZN(_AES_ENC_us23_n592 ) );
INV_X4 _AES_ENC_us23_U544  ( .A(_AES_ENC_us23_n925 ), .ZN(_AES_ENC_us23_n591 ) );
INV_X4 _AES_ENC_us23_U543  ( .A(_AES_ENC_us23_n824 ), .ZN(_AES_ENC_us23_n590 ) );
INV_X4 _AES_ENC_us23_U542  ( .A(_AES_ENC_us23_n959 ), .ZN(_AES_ENC_us23_n589 ) );
INV_X4 _AES_ENC_us23_U541  ( .A(_AES_ENC_us23_n779 ), .ZN(_AES_ENC_us23_n588 ) );
INV_X4 _AES_ENC_us23_U540  ( .A(_AES_ENC_us23_n794 ), .ZN(_AES_ENC_us23_n585 ) );
INV_X4 _AES_ENC_us23_U539  ( .A(_AES_ENC_us23_n880 ), .ZN(_AES_ENC_us23_n583 ) );
INV_X4 _AES_ENC_us23_U538  ( .A(_AES_ENC_sa23[7]), .ZN(_AES_ENC_us23_n581 ));
INV_X4 _AES_ENC_us23_U537  ( .A(_AES_ENC_us23_n992 ), .ZN(_AES_ENC_us23_n578 ) );
INV_X4 _AES_ENC_us23_U536  ( .A(_AES_ENC_us23_n1114 ), .ZN(_AES_ENC_us23_n577 ) );
INV_X4 _AES_ENC_us23_U535  ( .A(_AES_ENC_us23_n1092 ), .ZN(_AES_ENC_us23_n574 ) );
NOR2_X2 _AES_ENC_us23_U534  ( .A1(_AES_ENC_sa23[0]), .A2(_AES_ENC_sa23[6]),.ZN(_AES_ENC_us23_n1090 ) );
NOR2_X2 _AES_ENC_us23_U533  ( .A1(_AES_ENC_us23_n627 ), .A2(_AES_ENC_sa23[6]), .ZN(_AES_ENC_us23_n1070 ) );
NOR2_X2 _AES_ENC_us23_U532  ( .A1(_AES_ENC_sa23[4]), .A2(_AES_ENC_sa23[3]),.ZN(_AES_ENC_us23_n1025 ) );
INV_X4 _AES_ENC_us23_U531  ( .A(_AES_ENC_us23_n569 ), .ZN(_AES_ENC_us23_n572 ) );
NOR2_X2 _AES_ENC_us23_U530  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n765 ) );
NOR2_X2 _AES_ENC_us23_U529  ( .A1(_AES_ENC_sa23[4]), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n764 ) );
NOR2_X2 _AES_ENC_us23_U528  ( .A1(_AES_ENC_us23_n765 ), .A2(_AES_ENC_us23_n764 ), .ZN(_AES_ENC_us23_n766 ) );
NOR2_X2 _AES_ENC_us23_U527  ( .A1(_AES_ENC_us23_n766 ), .A2(_AES_ENC_us23_n589 ), .ZN(_AES_ENC_us23_n767 ) );
INV_X4 _AES_ENC_us23_U526  ( .A(_AES_ENC_sa23[3]), .ZN(_AES_ENC_us23_n624 ));
NAND3_X2 _AES_ENC_us23_U525  ( .A1(_AES_ENC_us23_n652 ), .A2(_AES_ENC_us23_n596 ), .A3(_AES_ENC_sa23[7]), .ZN(_AES_ENC_us23_n653 ));
NOR2_X2 _AES_ENC_us23_U524  ( .A1(_AES_ENC_us23_n593 ), .A2(_AES_ENC_sa23[5]), .ZN(_AES_ENC_us23_n925 ) );
NOR2_X2 _AES_ENC_us23_U523  ( .A1(_AES_ENC_sa23[5]), .A2(_AES_ENC_sa23[2]),.ZN(_AES_ENC_us23_n974 ) );
INV_X4 _AES_ENC_us23_U522  ( .A(_AES_ENC_sa23[5]), .ZN(_AES_ENC_us23_n596 ));
NOR2_X2 _AES_ENC_us23_U521  ( .A1(_AES_ENC_us23_n593 ), .A2(_AES_ENC_sa23[7]), .ZN(_AES_ENC_us23_n779 ) );
NAND3_X2 _AES_ENC_us23_U520  ( .A1(_AES_ENC_us23_n679 ), .A2(_AES_ENC_us23_n678 ), .A3(_AES_ENC_us23_n677 ), .ZN(_AES_ENC_sa23_sub[0] ) );
NOR2_X2 _AES_ENC_us23_U519  ( .A1(_AES_ENC_us23_n596 ), .A2(_AES_ENC_sa23[2]), .ZN(_AES_ENC_us23_n1048 ) );
NOR3_X2 _AES_ENC_us23_U518  ( .A1(_AES_ENC_us23_n581 ), .A2(_AES_ENC_sa23[5]), .A3(_AES_ENC_us23_n704 ), .ZN(_AES_ENC_us23_n706 ));
NOR2_X2 _AES_ENC_us23_U517  ( .A1(_AES_ENC_us23_n1117 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n707 ) );
NOR2_X2 _AES_ENC_us23_U516  ( .A1(_AES_ENC_sa23[4]), .A2(_AES_ENC_us23_n574 ), .ZN(_AES_ENC_us23_n705 ) );
NOR3_X2 _AES_ENC_us23_U515  ( .A1(_AES_ENC_us23_n707 ), .A2(_AES_ENC_us23_n706 ), .A3(_AES_ENC_us23_n705 ), .ZN(_AES_ENC_us23_n713 ) );
NOR4_X2 _AES_ENC_us23_U512  ( .A1(_AES_ENC_us23_n633 ), .A2(_AES_ENC_us23_n632 ), .A3(_AES_ENC_us23_n631 ), .A4(_AES_ENC_us23_n630 ), .ZN(_AES_ENC_us23_n634 ) );
NOR2_X2 _AES_ENC_us23_U510  ( .A1(_AES_ENC_us23_n629 ), .A2(_AES_ENC_us23_n628 ), .ZN(_AES_ENC_us23_n635 ) );
NAND3_X2 _AES_ENC_us23_U509  ( .A1(_AES_ENC_sa23[2]), .A2(_AES_ENC_sa23[7]), .A3(_AES_ENC_us23_n1059 ), .ZN(_AES_ENC_us23_n636 ) );
NOR2_X2 _AES_ENC_us23_U508  ( .A1(_AES_ENC_sa23[7]), .A2(_AES_ENC_sa23[2]),.ZN(_AES_ENC_us23_n794 ) );
NOR2_X2 _AES_ENC_us23_U507  ( .A1(_AES_ENC_sa23[4]), .A2(_AES_ENC_sa23[1]),.ZN(_AES_ENC_us23_n1102 ) );
NOR2_X2 _AES_ENC_us23_U506  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_sa23[3]), .ZN(_AES_ENC_us23_n1053 ) );
NOR2_X2 _AES_ENC_us23_U505  ( .A1(_AES_ENC_us23_n588 ), .A2(_AES_ENC_sa23[5]), .ZN(_AES_ENC_us23_n1024 ) );
NOR2_X2 _AES_ENC_us23_U504  ( .A1(_AES_ENC_us23_n577 ), .A2(_AES_ENC_sa23[2]), .ZN(_AES_ENC_us23_n1093 ) );
NOR2_X2 _AES_ENC_us23_U503  ( .A1(_AES_ENC_us23_n585 ), .A2(_AES_ENC_sa23[5]), .ZN(_AES_ENC_us23_n1094 ) );
NOR2_X2 _AES_ENC_us23_U502  ( .A1(_AES_ENC_us23_n612 ), .A2(_AES_ENC_sa23[3]), .ZN(_AES_ENC_us23_n931 ) );
INV_X4 _AES_ENC_us23_U501  ( .A(_AES_ENC_us23_n570 ), .ZN(_AES_ENC_us23_n573 ) );
NOR2_X2 _AES_ENC_us23_U500  ( .A1(_AES_ENC_us23_n1053 ), .A2(_AES_ENC_us23_n1095 ), .ZN(_AES_ENC_us23_n639 ) );
NOR3_X2 _AES_ENC_us23_U499  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n573 ), .A3(_AES_ENC_us23_n1074 ), .ZN(_AES_ENC_us23_n641 ) );
NOR2_X2 _AES_ENC_us23_U498  ( .A1(_AES_ENC_us23_n639 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n640 ) );
NOR2_X2 _AES_ENC_us23_U497  ( .A1(_AES_ENC_us23_n641 ), .A2(_AES_ENC_us23_n640 ), .ZN(_AES_ENC_us23_n646 ) );
NOR3_X2 _AES_ENC_us23_U496  ( .A1(_AES_ENC_us23_n995 ), .A2(_AES_ENC_us23_n578 ), .A3(_AES_ENC_us23_n994 ), .ZN(_AES_ENC_us23_n1002 ) );
NOR2_X2 _AES_ENC_us23_U495  ( .A1(_AES_ENC_us23_n909 ), .A2(_AES_ENC_us23_n908 ), .ZN(_AES_ENC_us23_n920 ) );
NOR2_X2 _AES_ENC_us23_U494  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n823 ) );
NOR2_X2 _AES_ENC_us23_U492  ( .A1(_AES_ENC_us23_n612 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n822 ) );
NOR2_X2 _AES_ENC_us23_U491  ( .A1(_AES_ENC_us23_n823 ), .A2(_AES_ENC_us23_n822 ), .ZN(_AES_ENC_us23_n825 ) );
NOR2_X2 _AES_ENC_us23_U490  ( .A1(_AES_ENC_sa23[1]), .A2(_AES_ENC_us23_n601 ), .ZN(_AES_ENC_us23_n913 ) );
NOR2_X2 _AES_ENC_us23_U489  ( .A1(_AES_ENC_us23_n913 ), .A2(_AES_ENC_us23_n1091 ), .ZN(_AES_ENC_us23_n914 ) );
NOR2_X2 _AES_ENC_us23_U488  ( .A1(_AES_ENC_us23_n826 ), .A2(_AES_ENC_us23_n572 ), .ZN(_AES_ENC_us23_n827 ) );
NOR3_X2 _AES_ENC_us23_U487  ( .A1(_AES_ENC_us23_n769 ), .A2(_AES_ENC_us23_n768 ), .A3(_AES_ENC_us23_n767 ), .ZN(_AES_ENC_us23_n775 ) );
NOR2_X2 _AES_ENC_us23_U486  ( .A1(_AES_ENC_us23_n1056 ), .A2(_AES_ENC_us23_n1053 ), .ZN(_AES_ENC_us23_n749 ) );
NOR2_X2 _AES_ENC_us23_U483  ( .A1(_AES_ENC_us23_n749 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n752 ) );
INV_X4 _AES_ENC_us23_U482  ( .A(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n626 ));
NOR2_X2 _AES_ENC_us23_U480  ( .A1(_AES_ENC_us23_n1054 ), .A2(_AES_ENC_us23_n1053 ), .ZN(_AES_ENC_us23_n1055 ) );
OR2_X4 _AES_ENC_us23_U479  ( .A1(_AES_ENC_us23_n1094 ), .A2(_AES_ENC_us23_n1093 ), .ZN(_AES_ENC_us23_n571 ) );
AND2_X2 _AES_ENC_us23_U478  ( .A1(_AES_ENC_us23_n571 ), .A2(_AES_ENC_us23_n1095 ), .ZN(_AES_ENC_us23_n1101 ) );
NOR2_X2 _AES_ENC_us23_U477  ( .A1(_AES_ENC_us23_n1074 ), .A2(_AES_ENC_us23_n931 ), .ZN(_AES_ENC_us23_n796 ) );
NOR2_X2 _AES_ENC_us23_U474  ( .A1(_AES_ENC_us23_n796 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n797 ) );
NOR2_X2 _AES_ENC_us23_U473  ( .A1(_AES_ENC_us23_n932 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n933 ) );
NOR2_X2 _AES_ENC_us23_U472  ( .A1(_AES_ENC_us23_n929 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n935 ) );
NOR2_X2 _AES_ENC_us23_U471  ( .A1(_AES_ENC_us23_n931 ), .A2(_AES_ENC_us23_n930 ), .ZN(_AES_ENC_us23_n934 ) );
NOR3_X2 _AES_ENC_us23_U470  ( .A1(_AES_ENC_us23_n935 ), .A2(_AES_ENC_us23_n934 ), .A3(_AES_ENC_us23_n933 ), .ZN(_AES_ENC_us23_n936 ) );
NOR2_X2 _AES_ENC_us23_U469  ( .A1(_AES_ENC_us23_n612 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n1075 ) );
NOR2_X2 _AES_ENC_us23_U468  ( .A1(_AES_ENC_us23_n572 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n949 ) );
NOR2_X2 _AES_ENC_us23_U467  ( .A1(_AES_ENC_us23_n1049 ), .A2(_AES_ENC_us23_n595 ), .ZN(_AES_ENC_us23_n1051 ) );
NOR2_X2 _AES_ENC_us23_U466  ( .A1(_AES_ENC_us23_n1051 ), .A2(_AES_ENC_us23_n1050 ), .ZN(_AES_ENC_us23_n1052 ) );
NOR2_X2 _AES_ENC_us23_U465  ( .A1(_AES_ENC_us23_n1052 ), .A2(_AES_ENC_us23_n604 ), .ZN(_AES_ENC_us23_n1064 ) );
NOR2_X2 _AES_ENC_us23_U464  ( .A1(_AES_ENC_sa23[1]), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n631 ) );
NOR2_X2 _AES_ENC_us23_U463  ( .A1(_AES_ENC_us23_n1025 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n980 ) );
NOR2_X2 _AES_ENC_us23_U462  ( .A1(_AES_ENC_us23_n1073 ), .A2(_AES_ENC_us23_n1094 ), .ZN(_AES_ENC_us23_n795 ) );
NOR2_X2 _AES_ENC_us23_U461  ( .A1(_AES_ENC_us23_n795 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n799 ) );
NOR2_X2 _AES_ENC_us23_U460  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n981 ) );
NOR2_X2 _AES_ENC_us23_U459  ( .A1(_AES_ENC_us23_n1102 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n643 ) );
NOR2_X2 _AES_ENC_us23_U458  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n624 ), .ZN(_AES_ENC_us23_n642 ) );
NOR2_X2 _AES_ENC_us23_U455  ( .A1(_AES_ENC_us23_n911 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n644 ) );
NOR4_X2 _AES_ENC_us23_U448  ( .A1(_AES_ENC_us23_n644 ), .A2(_AES_ENC_us23_n643 ), .A3(_AES_ENC_us23_n804 ), .A4(_AES_ENC_us23_n642 ), .ZN(_AES_ENC_us23_n645 ) );
NOR2_X2 _AES_ENC_us23_U447  ( .A1(_AES_ENC_us23_n1102 ), .A2(_AES_ENC_us23_n910 ), .ZN(_AES_ENC_us23_n932 ) );
NOR2_X2 _AES_ENC_us23_U442  ( .A1(_AES_ENC_us23_n1102 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n755 ) );
NOR2_X2 _AES_ENC_us23_U441  ( .A1(_AES_ENC_us23_n931 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n743 ) );
NOR2_X2 _AES_ENC_us23_U438  ( .A1(_AES_ENC_us23_n1072 ), .A2(_AES_ENC_us23_n1094 ), .ZN(_AES_ENC_us23_n930 ) );
NOR2_X2 _AES_ENC_us23_U435  ( .A1(_AES_ENC_us23_n1074 ), .A2(_AES_ENC_us23_n1025 ), .ZN(_AES_ENC_us23_n891 ) );
NOR2_X2 _AES_ENC_us23_U434  ( .A1(_AES_ENC_us23_n891 ), .A2(_AES_ENC_us23_n591 ), .ZN(_AES_ENC_us23_n894 ) );
NOR3_X2 _AES_ENC_us23_U433  ( .A1(_AES_ENC_us23_n601 ), .A2(_AES_ENC_sa23[1]), .A3(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n683 ));
INV_X4 _AES_ENC_us23_U428  ( .A(_AES_ENC_us23_n931 ), .ZN(_AES_ENC_us23_n601 ) );
NOR2_X2 _AES_ENC_us23_U427  ( .A1(_AES_ENC_us23_n996 ), .A2(_AES_ENC_us23_n931 ), .ZN(_AES_ENC_us23_n704 ) );
NOR2_X2 _AES_ENC_us23_U421  ( .A1(_AES_ENC_us23_n931 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n685 ) );
NOR2_X2 _AES_ENC_us23_U420  ( .A1(_AES_ENC_us23_n1029 ), .A2(_AES_ENC_us23_n1025 ), .ZN(_AES_ENC_us23_n1079 ) );
NOR3_X2 _AES_ENC_us23_U419  ( .A1(_AES_ENC_us23_n620 ), .A2(_AES_ENC_us23_n1025 ), .A3(_AES_ENC_us23_n594 ), .ZN(_AES_ENC_us23_n945 ) );
NOR2_X2 _AES_ENC_us23_U418  ( .A1(_AES_ENC_us23_n596 ), .A2(_AES_ENC_us23_n593 ), .ZN(_AES_ENC_us23_n800 ) );
NOR3_X2 _AES_ENC_us23_U417  ( .A1(_AES_ENC_us23_n598 ), .A2(_AES_ENC_us23_n581 ), .A3(_AES_ENC_us23_n593 ), .ZN(_AES_ENC_us23_n798 ) );
NOR3_X2 _AES_ENC_us23_U416  ( .A1(_AES_ENC_us23_n592 ), .A2(_AES_ENC_us23_n572 ), .A3(_AES_ENC_us23_n589 ), .ZN(_AES_ENC_us23_n962 ) );
NOR3_X2 _AES_ENC_us23_U415  ( .A1(_AES_ENC_us23_n959 ), .A2(_AES_ENC_us23_n572 ), .A3(_AES_ENC_us23_n591 ), .ZN(_AES_ENC_us23_n768 ) );
NOR3_X2 _AES_ENC_us23_U414  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n572 ), .A3(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n694 ) );
NOR3_X2 _AES_ENC_us23_U413  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n572 ), .A3(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n895 ) );
NOR3_X2 _AES_ENC_us23_U410  ( .A1(_AES_ENC_us23_n1008 ), .A2(_AES_ENC_us23_n1007 ), .A3(_AES_ENC_us23_n1006 ), .ZN(_AES_ENC_us23_n1018 ) );
NOR4_X2 _AES_ENC_us23_U409  ( .A1(_AES_ENC_us23_n806 ), .A2(_AES_ENC_us23_n805 ), .A3(_AES_ENC_us23_n804 ), .A4(_AES_ENC_us23_n803 ), .ZN(_AES_ENC_us23_n807 ) );
NOR3_X2 _AES_ENC_us23_U406  ( .A1(_AES_ENC_us23_n799 ), .A2(_AES_ENC_us23_n798 ), .A3(_AES_ENC_us23_n797 ), .ZN(_AES_ENC_us23_n808 ) );
NOR4_X2 _AES_ENC_us23_U405  ( .A1(_AES_ENC_us23_n843 ), .A2(_AES_ENC_us23_n842 ), .A3(_AES_ENC_us23_n841 ), .A4(_AES_ENC_us23_n840 ), .ZN(_AES_ENC_us23_n844 ) );
NOR2_X2 _AES_ENC_us23_U404  ( .A1(_AES_ENC_us23_n669 ), .A2(_AES_ENC_us23_n668 ), .ZN(_AES_ENC_us23_n673 ) );
NOR4_X2 _AES_ENC_us23_U403  ( .A1(_AES_ENC_us23_n946 ), .A2(_AES_ENC_us23_n1046 ), .A3(_AES_ENC_us23_n671 ), .A4(_AES_ENC_us23_n670 ), .ZN(_AES_ENC_us23_n672 ) );
NOR4_X2 _AES_ENC_us23_U401  ( .A1(_AES_ENC_us23_n711 ), .A2(_AES_ENC_us23_n710 ), .A3(_AES_ENC_us23_n709 ), .A4(_AES_ENC_us23_n708 ), .ZN(_AES_ENC_us23_n712 ) );
NOR4_X2 _AES_ENC_us23_U400  ( .A1(_AES_ENC_us23_n963 ), .A2(_AES_ENC_us23_n962 ), .A3(_AES_ENC_us23_n961 ), .A4(_AES_ENC_us23_n960 ), .ZN(_AES_ENC_us23_n964 ) );
NOR3_X2 _AES_ENC_us23_U399  ( .A1(_AES_ENC_us23_n1101 ), .A2(_AES_ENC_us23_n1100 ), .A3(_AES_ENC_us23_n1099 ), .ZN(_AES_ENC_us23_n1109 ) );
NOR3_X2 _AES_ENC_us23_U398  ( .A1(_AES_ENC_us23_n743 ), .A2(_AES_ENC_us23_n742 ), .A3(_AES_ENC_us23_n741 ), .ZN(_AES_ENC_us23_n744 ) );
NOR2_X2 _AES_ENC_us23_U397  ( .A1(_AES_ENC_us23_n697 ), .A2(_AES_ENC_us23_n658 ), .ZN(_AES_ENC_us23_n659 ) );
NOR2_X2 _AES_ENC_us23_U396  ( .A1(_AES_ENC_us23_n1078 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n1033 ) );
NOR2_X2 _AES_ENC_us23_U393  ( .A1(_AES_ENC_us23_n1031 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n1032 ) );
NOR3_X2 _AES_ENC_us23_U390  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n1025 ), .A3(_AES_ENC_us23_n1074 ), .ZN(_AES_ENC_us23_n1035 ) );
NOR4_X2 _AES_ENC_us23_U389  ( .A1(_AES_ENC_us23_n1035 ), .A2(_AES_ENC_us23_n1034 ), .A3(_AES_ENC_us23_n1033 ), .A4(_AES_ENC_us23_n1032 ), .ZN(_AES_ENC_us23_n1036 ) );
NOR2_X2 _AES_ENC_us23_U388  ( .A1(_AES_ENC_us23_n611 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n885 ) );
NOR2_X2 _AES_ENC_us23_U387  ( .A1(_AES_ENC_us23_n601 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n882 ) );
NOR2_X2 _AES_ENC_us23_U386  ( .A1(_AES_ENC_us23_n1053 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n884 ) );
NOR4_X2 _AES_ENC_us23_U385  ( .A1(_AES_ENC_us23_n885 ), .A2(_AES_ENC_us23_n884 ), .A3(_AES_ENC_us23_n883 ), .A4(_AES_ENC_us23_n882 ), .ZN(_AES_ENC_us23_n886 ) );
NOR2_X2 _AES_ENC_us23_U384  ( .A1(_AES_ENC_us23_n825 ), .A2(_AES_ENC_us23_n590 ), .ZN(_AES_ENC_us23_n830 ) );
NOR2_X2 _AES_ENC_us23_U383  ( .A1(_AES_ENC_us23_n827 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n829 ) );
NOR2_X2 _AES_ENC_us23_U382  ( .A1(_AES_ENC_us23_n572 ), .A2(_AES_ENC_us23_n574 ), .ZN(_AES_ENC_us23_n828 ) );
NOR4_X2 _AES_ENC_us23_U374  ( .A1(_AES_ENC_us23_n831 ), .A2(_AES_ENC_us23_n830 ), .A3(_AES_ENC_us23_n829 ), .A4(_AES_ENC_us23_n828 ), .ZN(_AES_ENC_us23_n832 ) );
NOR2_X2 _AES_ENC_us23_U373  ( .A1(_AES_ENC_us23_n587 ), .A2(_AES_ENC_us23_n603 ), .ZN(_AES_ENC_us23_n1104 ) );
NOR2_X2 _AES_ENC_us23_U372  ( .A1(_AES_ENC_us23_n1102 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n1106 ) );
NOR2_X2 _AES_ENC_us23_U370  ( .A1(_AES_ENC_us23_n1103 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n1105 ) );
NOR4_X2 _AES_ENC_us23_U369  ( .A1(_AES_ENC_us23_n1107 ), .A2(_AES_ENC_us23_n1106 ), .A3(_AES_ENC_us23_n1105 ), .A4(_AES_ENC_us23_n1104 ), .ZN(_AES_ENC_us23_n1108 ) );
NOR3_X2 _AES_ENC_us23_U368  ( .A1(_AES_ENC_us23_n959 ), .A2(_AES_ENC_us23_n624 ), .A3(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n963 ) );
NOR2_X2 _AES_ENC_us23_U367  ( .A1(_AES_ENC_us23_n596 ), .A2(_AES_ENC_us23_n581 ), .ZN(_AES_ENC_us23_n1114 ) );
INV_X4 _AES_ENC_us23_U366  ( .A(_AES_ENC_us23_n1024 ), .ZN(_AES_ENC_us23_n587 ) );
NOR3_X2 _AES_ENC_us23_U365  ( .A1(_AES_ENC_us23_n910 ), .A2(_AES_ENC_us23_n1059 ), .A3(_AES_ENC_us23_n593 ), .ZN(_AES_ENC_us23_n1115 ) );
INV_X4 _AES_ENC_us23_U364  ( .A(_AES_ENC_us23_n1094 ), .ZN(_AES_ENC_us23_n584 ) );
NOR2_X2 _AES_ENC_us23_U363  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n931 ), .ZN(_AES_ENC_us23_n1100 ) );
INV_X4 _AES_ENC_us23_U354  ( .A(_AES_ENC_us23_n1093 ), .ZN(_AES_ENC_us23_n575 ) );
NOR2_X2 _AES_ENC_us23_U353  ( .A1(_AES_ENC_us23_n569 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n929 ) );
NOR2_X2 _AES_ENC_us23_U352  ( .A1(_AES_ENC_us23_n609 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n926 ) );
NOR2_X2 _AES_ENC_us23_U351  ( .A1(_AES_ENC_us23_n572 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n1095 ) );
NOR2_X2 _AES_ENC_us23_U350  ( .A1(_AES_ENC_us23_n591 ), .A2(_AES_ENC_us23_n581 ), .ZN(_AES_ENC_us23_n1010 ) );
NOR2_X2 _AES_ENC_us23_U349  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n1103 ) );
NOR2_X2 _AES_ENC_us23_U348  ( .A1(_AES_ENC_us23_n614 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n1059 ) );
NOR2_X2 _AES_ENC_us23_U347  ( .A1(_AES_ENC_sa23[1]), .A2(_AES_ENC_us23_n1120 ), .ZN(_AES_ENC_us23_n1022 ) );
NOR2_X2 _AES_ENC_us23_U346  ( .A1(_AES_ENC_us23_n605 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n911 ) );
NOR2_X2 _AES_ENC_us23_U345  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_us23_n1025 ), .ZN(_AES_ENC_us23_n826 ) );
NOR2_X2 _AES_ENC_us23_U338  ( .A1(_AES_ENC_us23_n596 ), .A2(_AES_ENC_us23_n588 ), .ZN(_AES_ENC_us23_n1072 ) );
NOR2_X2 _AES_ENC_us23_U335  ( .A1(_AES_ENC_us23_n581 ), .A2(_AES_ENC_us23_n594 ), .ZN(_AES_ENC_us23_n956 ) );
NOR2_X2 _AES_ENC_us23_U329  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_us23_n612 ), .ZN(_AES_ENC_us23_n1121 ) );
NOR2_X2 _AES_ENC_us23_U328  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_us23_n612 ), .ZN(_AES_ENC_us23_n1058 ) );
NOR2_X2 _AES_ENC_us23_U327  ( .A1(_AES_ENC_us23_n577 ), .A2(_AES_ENC_us23_n593 ), .ZN(_AES_ENC_us23_n1073 ) );
NOR2_X2 _AES_ENC_us23_U325  ( .A1(_AES_ENC_sa23[1]), .A2(_AES_ENC_us23_n1025 ), .ZN(_AES_ENC_us23_n1054 ) );
NOR2_X2 _AES_ENC_us23_U324  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_us23_n931 ), .ZN(_AES_ENC_us23_n1029 ) );
NOR2_X2 _AES_ENC_us23_U319  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n1056 ) );
NOR2_X2 _AES_ENC_us23_U318  ( .A1(_AES_ENC_us23_n585 ), .A2(_AES_ENC_us23_n596 ), .ZN(_AES_ENC_us23_n1050 ) );
NOR2_X2 _AES_ENC_us23_U317  ( .A1(_AES_ENC_us23_n1121 ), .A2(_AES_ENC_us23_n1025 ), .ZN(_AES_ENC_us23_n1120 ) );
NOR2_X2 _AES_ENC_us23_U316  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_us23_n572 ), .ZN(_AES_ENC_us23_n1074 ) );
NOR2_X2 _AES_ENC_us23_U315  ( .A1(_AES_ENC_us23_n1058 ), .A2(_AES_ENC_us23_n1054 ), .ZN(_AES_ENC_us23_n878 ) );
NOR2_X2 _AES_ENC_us23_U314  ( .A1(_AES_ENC_us23_n878 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n879 ) );
NOR2_X2 _AES_ENC_us23_U312  ( .A1(_AES_ENC_us23_n880 ), .A2(_AES_ENC_us23_n879 ), .ZN(_AES_ENC_us23_n887 ) );
NOR2_X2 _AES_ENC_us23_U311  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n625 ), .ZN(_AES_ENC_us23_n957 ) );
NOR2_X2 _AES_ENC_us23_U310  ( .A1(_AES_ENC_us23_n958 ), .A2(_AES_ENC_us23_n957 ), .ZN(_AES_ENC_us23_n965 ) );
NOR3_X2 _AES_ENC_us23_U309  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n1091 ), .A3(_AES_ENC_us23_n1022 ), .ZN(_AES_ENC_us23_n720 ) );
NOR3_X2 _AES_ENC_us23_U303  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n1054 ), .A3(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n719 ) );
NOR2_X2 _AES_ENC_us23_U302  ( .A1(_AES_ENC_us23_n720 ), .A2(_AES_ENC_us23_n719 ), .ZN(_AES_ENC_us23_n726 ) );
NOR2_X2 _AES_ENC_us23_U300  ( .A1(_AES_ENC_us23_n585 ), .A2(_AES_ENC_us23_n613 ), .ZN(_AES_ENC_us23_n865 ) );
NOR2_X2 _AES_ENC_us23_U299  ( .A1(_AES_ENC_us23_n1059 ), .A2(_AES_ENC_us23_n1058 ), .ZN(_AES_ENC_us23_n1060 ) );
NOR2_X2 _AES_ENC_us23_U298  ( .A1(_AES_ENC_us23_n1095 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n668 ) );
NOR2_X2 _AES_ENC_us23_U297  ( .A1(_AES_ENC_us23_n826 ), .A2(_AES_ENC_us23_n573 ), .ZN(_AES_ENC_us23_n750 ) );
NOR2_X2 _AES_ENC_us23_U296  ( .A1(_AES_ENC_us23_n750 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n751 ) );
NOR2_X2 _AES_ENC_us23_U295  ( .A1(_AES_ENC_us23_n907 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n908 ) );
NOR2_X2 _AES_ENC_us23_U294  ( .A1(_AES_ENC_us23_n990 ), .A2(_AES_ENC_us23_n926 ), .ZN(_AES_ENC_us23_n780 ) );
NOR2_X2 _AES_ENC_us23_U293  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n606 ), .ZN(_AES_ENC_us23_n838 ) );
NOR2_X2 _AES_ENC_us23_U292  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n621 ), .ZN(_AES_ENC_us23_n837 ) );
NOR2_X2 _AES_ENC_us23_U291  ( .A1(_AES_ENC_us23_n838 ), .A2(_AES_ENC_us23_n837 ), .ZN(_AES_ENC_us23_n845 ) );
NOR2_X2 _AES_ENC_us23_U290  ( .A1(_AES_ENC_us23_n1022 ), .A2(_AES_ENC_us23_n1058 ), .ZN(_AES_ENC_us23_n740 ) );
NOR2_X2 _AES_ENC_us23_U284  ( .A1(_AES_ENC_us23_n740 ), .A2(_AES_ENC_us23_n594 ), .ZN(_AES_ENC_us23_n742 ) );
NOR2_X2 _AES_ENC_us23_U283  ( .A1(_AES_ENC_us23_n1098 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n1099 ) );
NOR2_X2 _AES_ENC_us23_U282  ( .A1(_AES_ENC_us23_n1120 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n993 ) );
NOR2_X2 _AES_ENC_us23_U281  ( .A1(_AES_ENC_us23_n993 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n994 ) );
NOR2_X2 _AES_ENC_us23_U280  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n609 ), .ZN(_AES_ENC_us23_n1026 ) );
NOR2_X2 _AES_ENC_us23_U279  ( .A1(_AES_ENC_us23_n573 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n1027 ) );
NOR2_X2 _AES_ENC_us23_U273  ( .A1(_AES_ENC_us23_n1027 ), .A2(_AES_ENC_us23_n1026 ), .ZN(_AES_ENC_us23_n1028 ) );
NOR2_X2 _AES_ENC_us23_U272  ( .A1(_AES_ENC_us23_n1029 ), .A2(_AES_ENC_us23_n1028 ), .ZN(_AES_ENC_us23_n1034 ) );
NOR4_X2 _AES_ENC_us23_U271  ( .A1(_AES_ENC_us23_n757 ), .A2(_AES_ENC_us23_n756 ), .A3(_AES_ENC_us23_n755 ), .A4(_AES_ENC_us23_n754 ), .ZN(_AES_ENC_us23_n758 ) );
NOR2_X2 _AES_ENC_us23_U270  ( .A1(_AES_ENC_us23_n752 ), .A2(_AES_ENC_us23_n751 ), .ZN(_AES_ENC_us23_n759 ) );
NOR2_X2 _AES_ENC_us23_U269  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n1071 ), .ZN(_AES_ENC_us23_n669 ) );
NOR2_X2 _AES_ENC_us23_U268  ( .A1(_AES_ENC_us23_n1056 ), .A2(_AES_ENC_us23_n990 ), .ZN(_AES_ENC_us23_n991 ) );
NOR2_X2 _AES_ENC_us23_U267  ( .A1(_AES_ENC_us23_n991 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n995 ) );
NOR2_X2 _AES_ENC_us23_U263  ( .A1(_AES_ENC_us23_n588 ), .A2(_AES_ENC_us23_n598 ), .ZN(_AES_ENC_us23_n1008 ) );
NOR2_X2 _AES_ENC_us23_U262  ( .A1(_AES_ENC_us23_n839 ), .A2(_AES_ENC_us23_n603 ), .ZN(_AES_ENC_us23_n693 ) );
NOR2_X2 _AES_ENC_us23_U258  ( .A1(_AES_ENC_us23_n587 ), .A2(_AES_ENC_us23_n906 ), .ZN(_AES_ENC_us23_n741 ) );
NOR2_X2 _AES_ENC_us23_U255  ( .A1(_AES_ENC_us23_n1054 ), .A2(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n763 ) );
NOR2_X2 _AES_ENC_us23_U254  ( .A1(_AES_ENC_us23_n763 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n769 ) );
NOR2_X2 _AES_ENC_us23_U253  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n618 ), .ZN(_AES_ENC_us23_n1007 ) );
NOR2_X2 _AES_ENC_us23_U252  ( .A1(_AES_ENC_us23_n591 ), .A2(_AES_ENC_us23_n599 ), .ZN(_AES_ENC_us23_n1123 ) );
NOR2_X2 _AES_ENC_us23_U251  ( .A1(_AES_ENC_us23_n591 ), .A2(_AES_ENC_us23_n598 ), .ZN(_AES_ENC_us23_n710 ) );
INV_X4 _AES_ENC_us23_U250  ( .A(_AES_ENC_us23_n1029 ), .ZN(_AES_ENC_us23_n603 ) );
NOR2_X2 _AES_ENC_us23_U243  ( .A1(_AES_ENC_us23_n594 ), .A2(_AES_ENC_us23_n607 ), .ZN(_AES_ENC_us23_n883 ) );
NOR2_X2 _AES_ENC_us23_U242  ( .A1(_AES_ENC_us23_n623 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n1125 ) );
NOR2_X2 _AES_ENC_us23_U241  ( .A1(_AES_ENC_us23_n911 ), .A2(_AES_ENC_us23_n910 ), .ZN(_AES_ENC_us23_n912 ) );
NOR2_X2 _AES_ENC_us23_U240  ( .A1(_AES_ENC_us23_n912 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n916 ) );
NOR2_X2 _AES_ENC_us23_U239  ( .A1(_AES_ENC_us23_n990 ), .A2(_AES_ENC_us23_n929 ), .ZN(_AES_ENC_us23_n892 ) );
NOR2_X2 _AES_ENC_us23_U238  ( .A1(_AES_ENC_us23_n892 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n893 ) );
NOR2_X2 _AES_ENC_us23_U237  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n621 ), .ZN(_AES_ENC_us23_n950 ) );
NOR2_X2 _AES_ENC_us23_U236  ( .A1(_AES_ENC_us23_n1079 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n1082 ) );
NOR2_X2 _AES_ENC_us23_U235  ( .A1(_AES_ENC_us23_n910 ), .A2(_AES_ENC_us23_n1056 ), .ZN(_AES_ENC_us23_n941 ) );
NOR2_X2 _AES_ENC_us23_U234  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n1077 ), .ZN(_AES_ENC_us23_n841 ) );
NOR2_X2 _AES_ENC_us23_U229  ( .A1(_AES_ENC_us23_n601 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n630 ) );
NOR2_X2 _AES_ENC_us23_U228  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n621 ), .ZN(_AES_ENC_us23_n806 ) );
NOR2_X2 _AES_ENC_us23_U227  ( .A1(_AES_ENC_us23_n601 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n948 ) );
NOR2_X2 _AES_ENC_us23_U226  ( .A1(_AES_ENC_us23_n587 ), .A2(_AES_ENC_us23_n620 ), .ZN(_AES_ENC_us23_n997 ) );
NOR2_X2 _AES_ENC_us23_U225  ( .A1(_AES_ENC_us23_n1121 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n1122 ) );
NOR2_X2 _AES_ENC_us23_U223  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n1023 ), .ZN(_AES_ENC_us23_n756 ) );
NOR2_X2 _AES_ENC_us23_U222  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n621 ), .ZN(_AES_ENC_us23_n870 ) );
NOR2_X2 _AES_ENC_us23_U221  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n569 ), .ZN(_AES_ENC_us23_n947 ) );
NOR2_X2 _AES_ENC_us23_U217  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n1077 ), .ZN(_AES_ENC_us23_n1084 ) );
NOR2_X2 _AES_ENC_us23_U213  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n855 ), .ZN(_AES_ENC_us23_n709 ) );
NOR2_X2 _AES_ENC_us23_U212  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n620 ), .ZN(_AES_ENC_us23_n868 ) );
NOR2_X2 _AES_ENC_us23_U211  ( .A1(_AES_ENC_us23_n1120 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n1124 ) );
NOR2_X2 _AES_ENC_us23_U210  ( .A1(_AES_ENC_us23_n1120 ), .A2(_AES_ENC_us23_n839 ), .ZN(_AES_ENC_us23_n842 ) );
NOR2_X2 _AES_ENC_us23_U209  ( .A1(_AES_ENC_us23_n1120 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n696 ) );
NOR2_X2 _AES_ENC_us23_U208  ( .A1(_AES_ENC_us23_n1074 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n1076 ) );
NOR2_X2 _AES_ENC_us23_U207  ( .A1(_AES_ENC_us23_n1074 ), .A2(_AES_ENC_us23_n609 ), .ZN(_AES_ENC_us23_n781 ) );
NOR3_X2 _AES_ENC_us23_U201  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n1056 ), .A3(_AES_ENC_us23_n990 ), .ZN(_AES_ENC_us23_n979 ) );
NOR3_X2 _AES_ENC_us23_U200  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n1058 ), .A3(_AES_ENC_us23_n1059 ), .ZN(_AES_ENC_us23_n854 ) );
NOR2_X2 _AES_ENC_us23_U199  ( .A1(_AES_ENC_us23_n996 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n869 ) );
NOR2_X2 _AES_ENC_us23_U198  ( .A1(_AES_ENC_us23_n1056 ), .A2(_AES_ENC_us23_n1074 ), .ZN(_AES_ENC_us23_n1057 ) );
NOR3_X2 _AES_ENC_us23_U197  ( .A1(_AES_ENC_us23_n588 ), .A2(_AES_ENC_us23_n1120 ), .A3(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n978 ) );
NOR2_X2 _AES_ENC_us23_U196  ( .A1(_AES_ENC_us23_n996 ), .A2(_AES_ENC_us23_n911 ), .ZN(_AES_ENC_us23_n1116 ) );
NOR2_X2 _AES_ENC_us23_U195  ( .A1(_AES_ENC_us23_n1074 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n754 ) );
NOR2_X2 _AES_ENC_us23_U194  ( .A1(_AES_ENC_us23_n926 ), .A2(_AES_ENC_us23_n1103 ), .ZN(_AES_ENC_us23_n977 ) );
NOR2_X2 _AES_ENC_us23_U187  ( .A1(_AES_ENC_us23_n839 ), .A2(_AES_ENC_us23_n824 ), .ZN(_AES_ENC_us23_n1092 ) );
NOR2_X2 _AES_ENC_us23_U186  ( .A1(_AES_ENC_us23_n573 ), .A2(_AES_ENC_us23_n1074 ), .ZN(_AES_ENC_us23_n684 ) );
NOR2_X2 _AES_ENC_us23_U185  ( .A1(_AES_ENC_us23_n826 ), .A2(_AES_ENC_us23_n1059 ), .ZN(_AES_ENC_us23_n907 ) );
NOR3_X2 _AES_ENC_us23_U184  ( .A1(_AES_ENC_us23_n577 ), .A2(_AES_ENC_us23_n1115 ), .A3(_AES_ENC_us23_n600 ), .ZN(_AES_ENC_us23_n831 ) );
NOR3_X2 _AES_ENC_us23_U183  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n1056 ), .A3(_AES_ENC_us23_n990 ), .ZN(_AES_ENC_us23_n896 ) );
NOR3_X2 _AES_ENC_us23_U182  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n573 ), .A3(_AES_ENC_us23_n1013 ), .ZN(_AES_ENC_us23_n670 ) );
NOR3_X2 _AES_ENC_us23_U181  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n1091 ), .A3(_AES_ENC_us23_n1022 ), .ZN(_AES_ENC_us23_n843 ) );
NOR2_X2 _AES_ENC_us23_U180  ( .A1(_AES_ENC_us23_n1029 ), .A2(_AES_ENC_us23_n1095 ), .ZN(_AES_ENC_us23_n735 ) );
NOR2_X2 _AES_ENC_us23_U174  ( .A1(_AES_ENC_us23_n1100 ), .A2(_AES_ENC_us23_n854 ), .ZN(_AES_ENC_us23_n860 ) );
NAND3_X2 _AES_ENC_us23_U173  ( .A1(_AES_ENC_us23_n569 ), .A2(_AES_ENC_us23_n603 ), .A3(_AES_ENC_us23_n681 ), .ZN(_AES_ENC_us23_n691 ) );
NOR2_X2 _AES_ENC_us23_U172  ( .A1(_AES_ENC_us23_n683 ), .A2(_AES_ENC_us23_n682 ), .ZN(_AES_ENC_us23_n690 ) );
NOR3_X2 _AES_ENC_us23_U171  ( .A1(_AES_ENC_us23_n695 ), .A2(_AES_ENC_us23_n694 ), .A3(_AES_ENC_us23_n693 ), .ZN(_AES_ENC_us23_n700 ) );
NOR4_X2 _AES_ENC_us23_U170  ( .A1(_AES_ENC_us23_n983 ), .A2(_AES_ENC_us23_n698 ), .A3(_AES_ENC_us23_n697 ), .A4(_AES_ENC_us23_n696 ), .ZN(_AES_ENC_us23_n699 ) );
NOR2_X2 _AES_ENC_us23_U169  ( .A1(_AES_ENC_us23_n946 ), .A2(_AES_ENC_us23_n945 ), .ZN(_AES_ENC_us23_n952 ) );
NOR4_X2 _AES_ENC_us23_U168  ( .A1(_AES_ENC_us23_n950 ), .A2(_AES_ENC_us23_n949 ), .A3(_AES_ENC_us23_n948 ), .A4(_AES_ENC_us23_n947 ), .ZN(_AES_ENC_us23_n951 ) );
NOR4_X2 _AES_ENC_us23_U162  ( .A1(_AES_ENC_us23_n896 ), .A2(_AES_ENC_us23_n895 ), .A3(_AES_ENC_us23_n894 ), .A4(_AES_ENC_us23_n893 ), .ZN(_AES_ENC_us23_n897 ) );
NOR2_X2 _AES_ENC_us23_U161  ( .A1(_AES_ENC_us23_n866 ), .A2(_AES_ENC_us23_n865 ), .ZN(_AES_ENC_us23_n872 ) );
NOR4_X2 _AES_ENC_us23_U160  ( .A1(_AES_ENC_us23_n870 ), .A2(_AES_ENC_us23_n869 ), .A3(_AES_ENC_us23_n868 ), .A4(_AES_ENC_us23_n867 ), .ZN(_AES_ENC_us23_n871 ) );
NOR4_X2 _AES_ENC_us23_U159  ( .A1(_AES_ENC_us23_n983 ), .A2(_AES_ENC_us23_n982 ), .A3(_AES_ENC_us23_n981 ), .A4(_AES_ENC_us23_n980 ), .ZN(_AES_ENC_us23_n984 ) );
NOR2_X2 _AES_ENC_us23_U158  ( .A1(_AES_ENC_us23_n979 ), .A2(_AES_ENC_us23_n978 ), .ZN(_AES_ENC_us23_n985 ) );
NOR4_X2 _AES_ENC_us23_U157  ( .A1(_AES_ENC_us23_n1125 ), .A2(_AES_ENC_us23_n1124 ), .A3(_AES_ENC_us23_n1123 ), .A4(_AES_ENC_us23_n1122 ), .ZN(_AES_ENC_us23_n1126 ) );
NOR4_X2 _AES_ENC_us23_U156  ( .A1(_AES_ENC_us23_n1084 ), .A2(_AES_ENC_us23_n1083 ), .A3(_AES_ENC_us23_n1082 ), .A4(_AES_ENC_us23_n1081 ), .ZN(_AES_ENC_us23_n1085 ) );
NOR2_X2 _AES_ENC_us23_U155  ( .A1(_AES_ENC_us23_n1076 ), .A2(_AES_ENC_us23_n1075 ), .ZN(_AES_ENC_us23_n1086 ) );
NOR3_X2 _AES_ENC_us23_U154  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n1054 ), .A3(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n961 ) );
NOR3_X2 _AES_ENC_us23_U153  ( .A1(_AES_ENC_us23_n609 ), .A2(_AES_ENC_us23_n1074 ), .A3(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n671 ) );
NOR2_X2 _AES_ENC_us23_U152  ( .A1(_AES_ENC_us23_n1057 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n1062 ) );
NOR2_X2 _AES_ENC_us23_U143  ( .A1(_AES_ENC_us23_n1055 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n1063 ) );
NOR2_X2 _AES_ENC_us23_U142  ( .A1(_AES_ENC_us23_n1060 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n1061 ) );
NOR4_X2 _AES_ENC_us23_U141  ( .A1(_AES_ENC_us23_n1064 ), .A2(_AES_ENC_us23_n1063 ), .A3(_AES_ENC_us23_n1062 ), .A4(_AES_ENC_us23_n1061 ), .ZN(_AES_ENC_us23_n1065 ) );
NOR3_X2 _AES_ENC_us23_U140  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n1120 ), .A3(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n918 ) );
NOR3_X2 _AES_ENC_us23_U132  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n573 ), .A3(_AES_ENC_us23_n1013 ), .ZN(_AES_ENC_us23_n917 ) );
NOR2_X2 _AES_ENC_us23_U131  ( .A1(_AES_ENC_us23_n914 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n915 ) );
NOR4_X2 _AES_ENC_us23_U130  ( .A1(_AES_ENC_us23_n918 ), .A2(_AES_ENC_us23_n917 ), .A3(_AES_ENC_us23_n916 ), .A4(_AES_ENC_us23_n915 ), .ZN(_AES_ENC_us23_n919 ) );
NOR2_X2 _AES_ENC_us23_U129  ( .A1(_AES_ENC_us23_n594 ), .A2(_AES_ENC_us23_n599 ), .ZN(_AES_ENC_us23_n771 ) );
NOR2_X2 _AES_ENC_us23_U128  ( .A1(_AES_ENC_us23_n1103 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n772 ) );
NOR2_X2 _AES_ENC_us23_U127  ( .A1(_AES_ENC_us23_n592 ), .A2(_AES_ENC_us23_n615 ), .ZN(_AES_ENC_us23_n773 ) );
NOR4_X2 _AES_ENC_us23_U126  ( .A1(_AES_ENC_us23_n773 ), .A2(_AES_ENC_us23_n772 ), .A3(_AES_ENC_us23_n771 ), .A4(_AES_ENC_us23_n770 ), .ZN(_AES_ENC_us23_n774 ) );
NOR2_X2 _AES_ENC_us23_U121  ( .A1(_AES_ENC_us23_n735 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n687 ) );
NOR2_X2 _AES_ENC_us23_U120  ( .A1(_AES_ENC_us23_n684 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n688 ) );
NOR2_X2 _AES_ENC_us23_U119  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n622 ), .ZN(_AES_ENC_us23_n686 ) );
NOR4_X2 _AES_ENC_us23_U118  ( .A1(_AES_ENC_us23_n688 ), .A2(_AES_ENC_us23_n687 ), .A3(_AES_ENC_us23_n686 ), .A4(_AES_ENC_us23_n685 ), .ZN(_AES_ENC_us23_n689 ) );
NOR2_X2 _AES_ENC_us23_U117  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n608 ), .ZN(_AES_ENC_us23_n858 ) );
NOR2_X2 _AES_ENC_us23_U116  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n855 ), .ZN(_AES_ENC_us23_n857 ) );
NOR2_X2 _AES_ENC_us23_U115  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n617 ), .ZN(_AES_ENC_us23_n856 ) );
NOR4_X2 _AES_ENC_us23_U106  ( .A1(_AES_ENC_us23_n858 ), .A2(_AES_ENC_us23_n857 ), .A3(_AES_ENC_us23_n856 ), .A4(_AES_ENC_us23_n958 ), .ZN(_AES_ENC_us23_n859 ) );
NOR2_X2 _AES_ENC_us23_U105  ( .A1(_AES_ENC_us23_n780 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n784 ) );
NOR2_X2 _AES_ENC_us23_U104  ( .A1(_AES_ENC_us23_n1117 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n782 ) );
NOR2_X2 _AES_ENC_us23_U103  ( .A1(_AES_ENC_us23_n781 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n783 ) );
NOR4_X2 _AES_ENC_us23_U102  ( .A1(_AES_ENC_us23_n880 ), .A2(_AES_ENC_us23_n784 ), .A3(_AES_ENC_us23_n783 ), .A4(_AES_ENC_us23_n782 ), .ZN(_AES_ENC_us23_n785 ) );
NOR2_X2 _AES_ENC_us23_U101  ( .A1(_AES_ENC_us23_n597 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n814 ) );
NOR2_X2 _AES_ENC_us23_U100  ( .A1(_AES_ENC_us23_n907 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n813 ) );
NOR3_X2 _AES_ENC_us23_U95  ( .A1(_AES_ENC_us23_n587 ), .A2(_AES_ENC_us23_n1058 ), .A3(_AES_ENC_us23_n1059 ), .ZN(_AES_ENC_us23_n815 ) );
NOR4_X2 _AES_ENC_us23_U94  ( .A1(_AES_ENC_us23_n815 ), .A2(_AES_ENC_us23_n814 ), .A3(_AES_ENC_us23_n813 ), .A4(_AES_ENC_us23_n812 ), .ZN(_AES_ENC_us23_n816 ) );
NOR2_X2 _AES_ENC_us23_U93  ( .A1(_AES_ENC_us23_n575 ), .A2(_AES_ENC_us23_n569 ), .ZN(_AES_ENC_us23_n721 ) );
NOR2_X2 _AES_ENC_us23_U92  ( .A1(_AES_ENC_us23_n1031 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n723 ) );
NOR2_X2 _AES_ENC_us23_U91  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n1096 ), .ZN(_AES_ENC_us23_n722 ) );
NOR4_X2 _AES_ENC_us23_U90  ( .A1(_AES_ENC_us23_n724 ), .A2(_AES_ENC_us23_n723 ), .A3(_AES_ENC_us23_n722 ), .A4(_AES_ENC_us23_n721 ), .ZN(_AES_ENC_us23_n725 ) );
NOR2_X2 _AES_ENC_us23_U89  ( .A1(_AES_ENC_us23_n911 ), .A2(_AES_ENC_us23_n990 ), .ZN(_AES_ENC_us23_n1009 ) );
NOR2_X2 _AES_ENC_us23_U88  ( .A1(_AES_ENC_us23_n1013 ), .A2(_AES_ENC_us23_n573 ), .ZN(_AES_ENC_us23_n1014 ) );
NOR2_X2 _AES_ENC_us23_U87  ( .A1(_AES_ENC_us23_n1014 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n1015 ) );
NOR4_X2 _AES_ENC_us23_U86  ( .A1(_AES_ENC_us23_n1016 ), .A2(_AES_ENC_us23_n1015 ), .A3(_AES_ENC_us23_n1119 ), .A4(_AES_ENC_us23_n1046 ), .ZN(_AES_ENC_us23_n1017 ) );
NOR2_X2 _AES_ENC_us23_U81  ( .A1(_AES_ENC_us23_n996 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n998 ) );
NOR2_X2 _AES_ENC_us23_U80  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n618 ), .ZN(_AES_ENC_us23_n1000 ) );
NOR2_X2 _AES_ENC_us23_U79  ( .A1(_AES_ENC_us23_n594 ), .A2(_AES_ENC_us23_n1096 ), .ZN(_AES_ENC_us23_n999 ) );
NOR4_X2 _AES_ENC_us23_U78  ( .A1(_AES_ENC_us23_n1000 ), .A2(_AES_ENC_us23_n999 ), .A3(_AES_ENC_us23_n998 ), .A4(_AES_ENC_us23_n997 ), .ZN(_AES_ENC_us23_n1001 ) );
NOR2_X2 _AES_ENC_us23_U74  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n1096 ), .ZN(_AES_ENC_us23_n697 ) );
NOR2_X2 _AES_ENC_us23_U73  ( .A1(_AES_ENC_us23_n609 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n958 ) );
NOR2_X2 _AES_ENC_us23_U72  ( .A1(_AES_ENC_us23_n911 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n983 ) );
NOR2_X2 _AES_ENC_us23_U71  ( .A1(_AES_ENC_us23_n1054 ), .A2(_AES_ENC_us23_n1103 ), .ZN(_AES_ENC_us23_n1031 ) );
INV_X4 _AES_ENC_us23_U65  ( .A(_AES_ENC_us23_n1050 ), .ZN(_AES_ENC_us23_n582 ) );
INV_X4 _AES_ENC_us23_U64  ( .A(_AES_ENC_us23_n1072 ), .ZN(_AES_ENC_us23_n586 ) );
INV_X4 _AES_ENC_us23_U63  ( .A(_AES_ENC_us23_n1073 ), .ZN(_AES_ENC_us23_n576 ) );
NOR2_X2 _AES_ENC_us23_U62  ( .A1(_AES_ENC_us23_n603 ), .A2(_AES_ENC_us23_n584 ), .ZN(_AES_ENC_us23_n880 ) );
NOR3_X2 _AES_ENC_us23_U61  ( .A1(_AES_ENC_us23_n826 ), .A2(_AES_ENC_us23_n1121 ), .A3(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n946 ) );
INV_X4 _AES_ENC_us23_U59  ( .A(_AES_ENC_us23_n1010 ), .ZN(_AES_ENC_us23_n579 ) );
NOR3_X2 _AES_ENC_us23_U58  ( .A1(_AES_ENC_us23_n573 ), .A2(_AES_ENC_us23_n1029 ), .A3(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n1119 ) );
INV_X4 _AES_ENC_us23_U57  ( .A(_AES_ENC_us23_n956 ), .ZN(_AES_ENC_us23_n580 ) );
NOR2_X2 _AES_ENC_us23_U50  ( .A1(_AES_ENC_us23_n601 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n1013 ) );
NOR2_X2 _AES_ENC_us23_U49  ( .A1(_AES_ENC_us23_n609 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n910 ) );
NOR2_X2 _AES_ENC_us23_U48  ( .A1(_AES_ENC_us23_n569 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n1091 ) );
NOR2_X2 _AES_ENC_us23_U47  ( .A1(_AES_ENC_us23_n614 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n990 ) );
NOR2_X2 _AES_ENC_us23_U46  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_us23_n1121 ), .ZN(_AES_ENC_us23_n996 ) );
NOR2_X2 _AES_ENC_us23_U45  ( .A1(_AES_ENC_us23_n592 ), .A2(_AES_ENC_us23_n622 ), .ZN(_AES_ENC_us23_n628 ) );
NOR2_X2 _AES_ENC_us23_U44  ( .A1(_AES_ENC_us23_n602 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n866 ) );
NOR2_X2 _AES_ENC_us23_U43  ( .A1(_AES_ENC_us23_n610 ), .A2(_AES_ENC_us23_n592 ), .ZN(_AES_ENC_us23_n1006 ) );
NOR2_X2 _AES_ENC_us23_U42  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n1117 ), .ZN(_AES_ENC_us23_n1118 ) );
NOR2_X2 _AES_ENC_us23_U41  ( .A1(_AES_ENC_us23_n1119 ), .A2(_AES_ENC_us23_n1118 ), .ZN(_AES_ENC_us23_n1127 ) );
NOR2_X2 _AES_ENC_us23_U36  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n616 ), .ZN(_AES_ENC_us23_n629 ) );
NOR2_X2 _AES_ENC_us23_U35  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n906 ), .ZN(_AES_ENC_us23_n909 ) );
NOR2_X2 _AES_ENC_us23_U34  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n607 ), .ZN(_AES_ENC_us23_n658 ) );
NOR2_X2 _AES_ENC_us23_U33  ( .A1(_AES_ENC_us23_n1116 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n695 ) );
NOR2_X2 _AES_ENC_us23_U32  ( .A1(_AES_ENC_us23_n1078 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n1083 ) );
NOR2_X2 _AES_ENC_us23_U31  ( .A1(_AES_ENC_us23_n941 ), .A2(_AES_ENC_us23_n579 ), .ZN(_AES_ENC_us23_n724 ) );
NOR2_X2 _AES_ENC_us23_U30  ( .A1(_AES_ENC_us23_n611 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n1107 ) );
NOR2_X2 _AES_ENC_us23_U29  ( .A1(_AES_ENC_us23_n602 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n840 ) );
NOR2_X2 _AES_ENC_us23_U24  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n623 ), .ZN(_AES_ENC_us23_n633 ) );
NOR2_X2 _AES_ENC_us23_U23  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n1080 ), .ZN(_AES_ENC_us23_n1081 ) );
NOR2_X2 _AES_ENC_us23_U21  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n1045 ), .ZN(_AES_ENC_us23_n812 ) );
NOR2_X2 _AES_ENC_us23_U20  ( .A1(_AES_ENC_us23_n1009 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n960 ) );
NOR2_X2 _AES_ENC_us23_U19  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n619 ), .ZN(_AES_ENC_us23_n982 ) );
NOR2_X2 _AES_ENC_us23_U18  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n616 ), .ZN(_AES_ENC_us23_n757 ) );
NOR2_X2 _AES_ENC_us23_U17  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n598 ), .ZN(_AES_ENC_us23_n698 ) );
NOR2_X2 _AES_ENC_us23_U16  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n605 ), .ZN(_AES_ENC_us23_n708 ) );
NOR2_X2 _AES_ENC_us23_U15  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n603 ), .ZN(_AES_ENC_us23_n770 ) );
NOR2_X2 _AES_ENC_us23_U10  ( .A1(_AES_ENC_us23_n605 ), .A2(_AES_ENC_us23_n576 ), .ZN(_AES_ENC_us23_n803 ) );
NOR2_X2 _AES_ENC_us23_U9  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n881 ), .ZN(_AES_ENC_us23_n711 ) );
NOR2_X2 _AES_ENC_us23_U8  ( .A1(_AES_ENC_us23_n580 ), .A2(_AES_ENC_us23_n603 ), .ZN(_AES_ENC_us23_n867 ) );
NOR2_X2 _AES_ENC_us23_U7  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n615 ), .ZN(_AES_ENC_us23_n804 ) );
NOR2_X2 _AES_ENC_us23_U6  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n609 ), .ZN(_AES_ENC_us23_n1046 ) );
OR2_X4 _AES_ENC_us23_U5  ( .A1(_AES_ENC_us23_n612 ), .A2(_AES_ENC_sa23[1]),.ZN(_AES_ENC_us23_n570 ) );
OR2_X4 _AES_ENC_us23_U4  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_sa23[4]),.ZN(_AES_ENC_us23_n569 ) );
NAND2_X2 _AES_ENC_us23_U514  ( .A1(_AES_ENC_us23_n1121 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n1030 ) );
AND2_X2 _AES_ENC_us23_U513  ( .A1(_AES_ENC_us23_n607 ), .A2(_AES_ENC_us23_n1030 ), .ZN(_AES_ENC_us23_n1049 ) );
NAND2_X2 _AES_ENC_us23_U511  ( .A1(_AES_ENC_us23_n1049 ), .A2(_AES_ENC_us23_n794 ), .ZN(_AES_ENC_us23_n637 ) );
AND2_X2 _AES_ENC_us23_U493  ( .A1(_AES_ENC_us23_n779 ), .A2(_AES_ENC_us23_n996 ), .ZN(_AES_ENC_us23_n632 ) );
NAND4_X2 _AES_ENC_us23_U485  ( .A1(_AES_ENC_us23_n637 ), .A2(_AES_ENC_us23_n636 ), .A3(_AES_ENC_us23_n635 ), .A4(_AES_ENC_us23_n634 ), .ZN(_AES_ENC_us23_n638 ) );
NAND2_X2 _AES_ENC_us23_U484  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n638 ), .ZN(_AES_ENC_us23_n679 ) );
NAND2_X2 _AES_ENC_us23_U481  ( .A1(_AES_ENC_us23_n1094 ), .A2(_AES_ENC_us23_n613 ), .ZN(_AES_ENC_us23_n648 ) );
NAND2_X2 _AES_ENC_us23_U476  ( .A1(_AES_ENC_us23_n619 ), .A2(_AES_ENC_us23_n598 ), .ZN(_AES_ENC_us23_n762 ) );
NAND2_X2 _AES_ENC_us23_U475  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n762 ), .ZN(_AES_ENC_us23_n647 ) );
NAND4_X2 _AES_ENC_us23_U457  ( .A1(_AES_ENC_us23_n648 ), .A2(_AES_ENC_us23_n647 ), .A3(_AES_ENC_us23_n646 ), .A4(_AES_ENC_us23_n645 ), .ZN(_AES_ENC_us23_n649 ) );
NAND2_X2 _AES_ENC_us23_U456  ( .A1(_AES_ENC_sa23[0]), .A2(_AES_ENC_us23_n649 ), .ZN(_AES_ENC_us23_n665 ) );
NAND2_X2 _AES_ENC_us23_U454  ( .A1(_AES_ENC_us23_n626 ), .A2(_AES_ENC_us23_n601 ), .ZN(_AES_ENC_us23_n855 ) );
NAND2_X2 _AES_ENC_us23_U453  ( .A1(_AES_ENC_us23_n617 ), .A2(_AES_ENC_us23_n855 ), .ZN(_AES_ENC_us23_n821 ) );
NAND2_X2 _AES_ENC_us23_U452  ( .A1(_AES_ENC_us23_n1093 ), .A2(_AES_ENC_us23_n821 ), .ZN(_AES_ENC_us23_n662 ) );
NAND2_X2 _AES_ENC_us23_U451  ( .A1(_AES_ENC_us23_n605 ), .A2(_AES_ENC_us23_n620 ), .ZN(_AES_ENC_us23_n650 ) );
NAND2_X2 _AES_ENC_us23_U450  ( .A1(_AES_ENC_us23_n956 ), .A2(_AES_ENC_us23_n650 ), .ZN(_AES_ENC_us23_n661 ) );
NAND2_X2 _AES_ENC_us23_U449  ( .A1(_AES_ENC_us23_n596 ), .A2(_AES_ENC_us23_n581 ), .ZN(_AES_ENC_us23_n839 ) );
OR2_X2 _AES_ENC_us23_U446  ( .A1(_AES_ENC_us23_n839 ), .A2(_AES_ENC_us23_n932 ), .ZN(_AES_ENC_us23_n656 ) );
NAND2_X2 _AES_ENC_us23_U445  ( .A1(_AES_ENC_us23_n624 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n1096 ) );
NAND2_X2 _AES_ENC_us23_U444  ( .A1(_AES_ENC_us23_n1030 ), .A2(_AES_ENC_us23_n1096 ), .ZN(_AES_ENC_us23_n651 ) );
NAND2_X2 _AES_ENC_us23_U443  ( .A1(_AES_ENC_us23_n1114 ), .A2(_AES_ENC_us23_n651 ), .ZN(_AES_ENC_us23_n655 ) );
OR3_X2 _AES_ENC_us23_U440  ( .A1(_AES_ENC_us23_n1079 ), .A2(_AES_ENC_sa23[7]), .A3(_AES_ENC_us23_n596 ), .ZN(_AES_ENC_us23_n654 ));
NAND2_X2 _AES_ENC_us23_U439  ( .A1(_AES_ENC_us23_n623 ), .A2(_AES_ENC_us23_n619 ), .ZN(_AES_ENC_us23_n652 ) );
NAND4_X2 _AES_ENC_us23_U437  ( .A1(_AES_ENC_us23_n656 ), .A2(_AES_ENC_us23_n655 ), .A3(_AES_ENC_us23_n654 ), .A4(_AES_ENC_us23_n653 ), .ZN(_AES_ENC_us23_n657 ) );
NAND2_X2 _AES_ENC_us23_U436  ( .A1(_AES_ENC_sa23[2]), .A2(_AES_ENC_us23_n657 ), .ZN(_AES_ENC_us23_n660 ) );
NAND4_X2 _AES_ENC_us23_U432  ( .A1(_AES_ENC_us23_n662 ), .A2(_AES_ENC_us23_n661 ), .A3(_AES_ENC_us23_n660 ), .A4(_AES_ENC_us23_n659 ), .ZN(_AES_ENC_us23_n663 ) );
NAND2_X2 _AES_ENC_us23_U431  ( .A1(_AES_ENC_us23_n663 ), .A2(_AES_ENC_us23_n627 ), .ZN(_AES_ENC_us23_n664 ) );
NAND2_X2 _AES_ENC_us23_U430  ( .A1(_AES_ENC_us23_n665 ), .A2(_AES_ENC_us23_n664 ), .ZN(_AES_ENC_us23_n666 ) );
NAND2_X2 _AES_ENC_us23_U429  ( .A1(_AES_ENC_sa23[6]), .A2(_AES_ENC_us23_n666 ), .ZN(_AES_ENC_us23_n678 ) );
NAND2_X2 _AES_ENC_us23_U426  ( .A1(_AES_ENC_us23_n735 ), .A2(_AES_ENC_us23_n1093 ), .ZN(_AES_ENC_us23_n675 ) );
NAND2_X2 _AES_ENC_us23_U425  ( .A1(_AES_ENC_us23_n625 ), .A2(_AES_ENC_us23_n607 ), .ZN(_AES_ENC_us23_n1045 ) );
OR2_X2 _AES_ENC_us23_U424  ( .A1(_AES_ENC_us23_n1045 ), .A2(_AES_ENC_us23_n586 ), .ZN(_AES_ENC_us23_n674 ) );
NAND2_X2 _AES_ENC_us23_U423  ( .A1(_AES_ENC_sa23[1]), .A2(_AES_ENC_us23_n609 ), .ZN(_AES_ENC_us23_n667 ) );
NAND2_X2 _AES_ENC_us23_U422  ( .A1(_AES_ENC_us23_n605 ), .A2(_AES_ENC_us23_n667 ), .ZN(_AES_ENC_us23_n1071 ) );
NAND4_X2 _AES_ENC_us23_U412  ( .A1(_AES_ENC_us23_n675 ), .A2(_AES_ENC_us23_n674 ), .A3(_AES_ENC_us23_n673 ), .A4(_AES_ENC_us23_n672 ), .ZN(_AES_ENC_us23_n676 ) );
NAND2_X2 _AES_ENC_us23_U411  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n676 ), .ZN(_AES_ENC_us23_n677 ) );
NAND2_X2 _AES_ENC_us23_U408  ( .A1(_AES_ENC_us23_n800 ), .A2(_AES_ENC_us23_n1022 ), .ZN(_AES_ENC_us23_n680 ) );
NAND2_X2 _AES_ENC_us23_U407  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n680 ), .ZN(_AES_ENC_us23_n681 ) );
AND2_X2 _AES_ENC_us23_U402  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n684 ), .ZN(_AES_ENC_us23_n682 ) );
NAND4_X2 _AES_ENC_us23_U395  ( .A1(_AES_ENC_us23_n691 ), .A2(_AES_ENC_us23_n583 ), .A3(_AES_ENC_us23_n690 ), .A4(_AES_ENC_us23_n689 ), .ZN(_AES_ENC_us23_n692 ) );
NAND2_X2 _AES_ENC_us23_U394  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n692 ), .ZN(_AES_ENC_us23_n733 ) );
NAND2_X2 _AES_ENC_us23_U392  ( .A1(_AES_ENC_us23_n977 ), .A2(_AES_ENC_us23_n1050 ), .ZN(_AES_ENC_us23_n702 ) );
NAND2_X2 _AES_ENC_us23_U391  ( .A1(_AES_ENC_us23_n1093 ), .A2(_AES_ENC_us23_n1045 ), .ZN(_AES_ENC_us23_n701 ) );
NAND4_X2 _AES_ENC_us23_U381  ( .A1(_AES_ENC_us23_n702 ), .A2(_AES_ENC_us23_n701 ), .A3(_AES_ENC_us23_n700 ), .A4(_AES_ENC_us23_n699 ), .ZN(_AES_ENC_us23_n703 ) );
NAND2_X2 _AES_ENC_us23_U380  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n703 ), .ZN(_AES_ENC_us23_n732 ) );
AND2_X2 _AES_ENC_us23_U379  ( .A1(_AES_ENC_sa23[0]), .A2(_AES_ENC_sa23[6]),.ZN(_AES_ENC_us23_n1113 ) );
NAND2_X2 _AES_ENC_us23_U378  ( .A1(_AES_ENC_us23_n619 ), .A2(_AES_ENC_us23_n1030 ), .ZN(_AES_ENC_us23_n881 ) );
NAND2_X2 _AES_ENC_us23_U377  ( .A1(_AES_ENC_us23_n1093 ), .A2(_AES_ENC_us23_n881 ), .ZN(_AES_ENC_us23_n715 ) );
NAND2_X2 _AES_ENC_us23_U376  ( .A1(_AES_ENC_us23_n1010 ), .A2(_AES_ENC_us23_n622 ), .ZN(_AES_ENC_us23_n714 ) );
NAND2_X2 _AES_ENC_us23_U375  ( .A1(_AES_ENC_us23_n855 ), .A2(_AES_ENC_us23_n625 ), .ZN(_AES_ENC_us23_n1117 ) );
XNOR2_X2 _AES_ENC_us23_U371  ( .A(_AES_ENC_us23_n593 ), .B(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n824 ) );
NAND4_X2 _AES_ENC_us23_U362  ( .A1(_AES_ENC_us23_n715 ), .A2(_AES_ENC_us23_n714 ), .A3(_AES_ENC_us23_n713 ), .A4(_AES_ENC_us23_n712 ), .ZN(_AES_ENC_us23_n716 ) );
NAND2_X2 _AES_ENC_us23_U361  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n716 ), .ZN(_AES_ENC_us23_n731 ) );
AND2_X2 _AES_ENC_us23_U360  ( .A1(_AES_ENC_sa23[6]), .A2(_AES_ENC_us23_n627 ), .ZN(_AES_ENC_us23_n1131 ) );
NAND2_X2 _AES_ENC_us23_U359  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n717 ) );
NAND2_X2 _AES_ENC_us23_U358  ( .A1(_AES_ENC_us23_n1029 ), .A2(_AES_ENC_us23_n717 ), .ZN(_AES_ENC_us23_n728 ) );
NAND2_X2 _AES_ENC_us23_U357  ( .A1(_AES_ENC_sa23[1]), .A2(_AES_ENC_us23_n612 ), .ZN(_AES_ENC_us23_n1097 ) );
NAND2_X2 _AES_ENC_us23_U356  ( .A1(_AES_ENC_us23_n610 ), .A2(_AES_ENC_us23_n1097 ), .ZN(_AES_ENC_us23_n718 ) );
NAND2_X2 _AES_ENC_us23_U355  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n718 ), .ZN(_AES_ENC_us23_n727 ) );
NAND4_X2 _AES_ENC_us23_U344  ( .A1(_AES_ENC_us23_n728 ), .A2(_AES_ENC_us23_n727 ), .A3(_AES_ENC_us23_n726 ), .A4(_AES_ENC_us23_n725 ), .ZN(_AES_ENC_us23_n729 ) );
NAND2_X2 _AES_ENC_us23_U343  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n729 ), .ZN(_AES_ENC_us23_n730 ) );
NAND4_X2 _AES_ENC_us23_U342  ( .A1(_AES_ENC_us23_n733 ), .A2(_AES_ENC_us23_n732 ), .A3(_AES_ENC_us23_n731 ), .A4(_AES_ENC_us23_n730 ), .ZN(_AES_ENC_sa23_sub[1] ) );
NAND2_X2 _AES_ENC_us23_U341  ( .A1(_AES_ENC_sa23[7]), .A2(_AES_ENC_us23_n593 ), .ZN(_AES_ENC_us23_n734 ) );
NAND2_X2 _AES_ENC_us23_U340  ( .A1(_AES_ENC_us23_n734 ), .A2(_AES_ENC_us23_n588 ), .ZN(_AES_ENC_us23_n738 ) );
OR4_X2 _AES_ENC_us23_U339  ( .A1(_AES_ENC_us23_n738 ), .A2(_AES_ENC_us23_n596 ), .A3(_AES_ENC_us23_n826 ), .A4(_AES_ENC_us23_n1121 ), .ZN(_AES_ENC_us23_n746 ) );
NAND2_X2 _AES_ENC_us23_U337  ( .A1(_AES_ENC_us23_n1100 ), .A2(_AES_ENC_us23_n617 ), .ZN(_AES_ENC_us23_n992 ) );
OR2_X2 _AES_ENC_us23_U336  ( .A1(_AES_ENC_us23_n592 ), .A2(_AES_ENC_us23_n735 ), .ZN(_AES_ENC_us23_n737 ) );
NAND2_X2 _AES_ENC_us23_U334  ( .A1(_AES_ENC_us23_n605 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n753 ) );
NAND2_X2 _AES_ENC_us23_U333  ( .A1(_AES_ENC_us23_n603 ), .A2(_AES_ENC_us23_n753 ), .ZN(_AES_ENC_us23_n1080 ) );
NAND2_X2 _AES_ENC_us23_U332  ( .A1(_AES_ENC_us23_n1048 ), .A2(_AES_ENC_us23_n602 ), .ZN(_AES_ENC_us23_n736 ) );
NAND2_X2 _AES_ENC_us23_U331  ( .A1(_AES_ENC_us23_n737 ), .A2(_AES_ENC_us23_n736 ), .ZN(_AES_ENC_us23_n739 ) );
NAND2_X2 _AES_ENC_us23_U330  ( .A1(_AES_ENC_us23_n739 ), .A2(_AES_ENC_us23_n738 ), .ZN(_AES_ENC_us23_n745 ) );
NAND2_X2 _AES_ENC_us23_U326  ( .A1(_AES_ENC_us23_n1096 ), .A2(_AES_ENC_us23_n598 ), .ZN(_AES_ENC_us23_n906 ) );
NAND4_X2 _AES_ENC_us23_U323  ( .A1(_AES_ENC_us23_n746 ), .A2(_AES_ENC_us23_n992 ), .A3(_AES_ENC_us23_n745 ), .A4(_AES_ENC_us23_n744 ), .ZN(_AES_ENC_us23_n747 ) );
NAND2_X2 _AES_ENC_us23_U322  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n747 ), .ZN(_AES_ENC_us23_n793 ) );
NAND2_X2 _AES_ENC_us23_U321  ( .A1(_AES_ENC_us23_n606 ), .A2(_AES_ENC_us23_n855 ), .ZN(_AES_ENC_us23_n748 ) );
NAND2_X2 _AES_ENC_us23_U320  ( .A1(_AES_ENC_us23_n956 ), .A2(_AES_ENC_us23_n748 ), .ZN(_AES_ENC_us23_n760 ) );
NAND2_X2 _AES_ENC_us23_U313  ( .A1(_AES_ENC_us23_n598 ), .A2(_AES_ENC_us23_n753 ), .ZN(_AES_ENC_us23_n1023 ) );
NAND4_X2 _AES_ENC_us23_U308  ( .A1(_AES_ENC_us23_n760 ), .A2(_AES_ENC_us23_n992 ), .A3(_AES_ENC_us23_n759 ), .A4(_AES_ENC_us23_n758 ), .ZN(_AES_ENC_us23_n761 ) );
NAND2_X2 _AES_ENC_us23_U307  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n761 ), .ZN(_AES_ENC_us23_n792 ) );
NAND2_X2 _AES_ENC_us23_U306  ( .A1(_AES_ENC_us23_n606 ), .A2(_AES_ENC_us23_n610 ), .ZN(_AES_ENC_us23_n989 ) );
NAND2_X2 _AES_ENC_us23_U305  ( .A1(_AES_ENC_us23_n1050 ), .A2(_AES_ENC_us23_n989 ), .ZN(_AES_ENC_us23_n777 ) );
NAND2_X2 _AES_ENC_us23_U304  ( .A1(_AES_ENC_us23_n1093 ), .A2(_AES_ENC_us23_n762 ), .ZN(_AES_ENC_us23_n776 ) );
XNOR2_X2 _AES_ENC_us23_U301  ( .A(_AES_ENC_sa23[7]), .B(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n959 ) );
NAND4_X2 _AES_ENC_us23_U289  ( .A1(_AES_ENC_us23_n777 ), .A2(_AES_ENC_us23_n776 ), .A3(_AES_ENC_us23_n775 ), .A4(_AES_ENC_us23_n774 ), .ZN(_AES_ENC_us23_n778 ) );
NAND2_X2 _AES_ENC_us23_U288  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n778 ), .ZN(_AES_ENC_us23_n791 ) );
NAND2_X2 _AES_ENC_us23_U287  ( .A1(_AES_ENC_us23_n1056 ), .A2(_AES_ENC_us23_n1050 ), .ZN(_AES_ENC_us23_n788 ) );
NAND2_X2 _AES_ENC_us23_U286  ( .A1(_AES_ENC_us23_n1091 ), .A2(_AES_ENC_us23_n779 ), .ZN(_AES_ENC_us23_n787 ) );
NAND2_X2 _AES_ENC_us23_U285  ( .A1(_AES_ENC_us23_n956 ), .A2(_AES_ENC_sa23[1]), .ZN(_AES_ENC_us23_n786 ) );
NAND4_X2 _AES_ENC_us23_U278  ( .A1(_AES_ENC_us23_n788 ), .A2(_AES_ENC_us23_n787 ), .A3(_AES_ENC_us23_n786 ), .A4(_AES_ENC_us23_n785 ), .ZN(_AES_ENC_us23_n789 ) );
NAND2_X2 _AES_ENC_us23_U277  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n789 ), .ZN(_AES_ENC_us23_n790 ) );
NAND4_X2 _AES_ENC_us23_U276  ( .A1(_AES_ENC_us23_n793 ), .A2(_AES_ENC_us23_n792 ), .A3(_AES_ENC_us23_n791 ), .A4(_AES_ENC_us23_n790 ), .ZN(_AES_ENC_sa23_sub[2] ) );
NAND2_X2 _AES_ENC_us23_U275  ( .A1(_AES_ENC_us23_n1059 ), .A2(_AES_ENC_us23_n794 ), .ZN(_AES_ENC_us23_n810 ) );
NAND2_X2 _AES_ENC_us23_U274  ( .A1(_AES_ENC_us23_n1049 ), .A2(_AES_ENC_us23_n956 ), .ZN(_AES_ENC_us23_n809 ) );
OR2_X2 _AES_ENC_us23_U266  ( .A1(_AES_ENC_us23_n1096 ), .A2(_AES_ENC_us23_n587 ), .ZN(_AES_ENC_us23_n802 ) );
NAND2_X2 _AES_ENC_us23_U265  ( .A1(_AES_ENC_us23_n1053 ), .A2(_AES_ENC_us23_n800 ), .ZN(_AES_ENC_us23_n801 ) );
NAND2_X2 _AES_ENC_us23_U264  ( .A1(_AES_ENC_us23_n802 ), .A2(_AES_ENC_us23_n801 ), .ZN(_AES_ENC_us23_n805 ) );
NAND4_X2 _AES_ENC_us23_U261  ( .A1(_AES_ENC_us23_n810 ), .A2(_AES_ENC_us23_n809 ), .A3(_AES_ENC_us23_n808 ), .A4(_AES_ENC_us23_n807 ), .ZN(_AES_ENC_us23_n811 ) );
NAND2_X2 _AES_ENC_us23_U260  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n811 ), .ZN(_AES_ENC_us23_n852 ) );
OR2_X2 _AES_ENC_us23_U259  ( .A1(_AES_ENC_us23_n1023 ), .A2(_AES_ENC_us23_n575 ), .ZN(_AES_ENC_us23_n819 ) );
OR2_X2 _AES_ENC_us23_U257  ( .A1(_AES_ENC_us23_n570 ), .A2(_AES_ENC_us23_n930 ), .ZN(_AES_ENC_us23_n818 ) );
NAND2_X2 _AES_ENC_us23_U256  ( .A1(_AES_ENC_us23_n1013 ), .A2(_AES_ENC_us23_n1094 ), .ZN(_AES_ENC_us23_n817 ) );
NAND4_X2 _AES_ENC_us23_U249  ( .A1(_AES_ENC_us23_n819 ), .A2(_AES_ENC_us23_n818 ), .A3(_AES_ENC_us23_n817 ), .A4(_AES_ENC_us23_n816 ), .ZN(_AES_ENC_us23_n820 ) );
NAND2_X2 _AES_ENC_us23_U248  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n820 ), .ZN(_AES_ENC_us23_n851 ) );
NAND2_X2 _AES_ENC_us23_U247  ( .A1(_AES_ENC_us23_n956 ), .A2(_AES_ENC_us23_n1080 ), .ZN(_AES_ENC_us23_n835 ) );
NAND2_X2 _AES_ENC_us23_U246  ( .A1(_AES_ENC_us23_n570 ), .A2(_AES_ENC_us23_n1030 ), .ZN(_AES_ENC_us23_n1047 ) );
OR2_X2 _AES_ENC_us23_U245  ( .A1(_AES_ENC_us23_n1047 ), .A2(_AES_ENC_us23_n582 ), .ZN(_AES_ENC_us23_n834 ) );
NAND2_X2 _AES_ENC_us23_U244  ( .A1(_AES_ENC_us23_n1072 ), .A2(_AES_ENC_us23_n620 ), .ZN(_AES_ENC_us23_n833 ) );
NAND4_X2 _AES_ENC_us23_U233  ( .A1(_AES_ENC_us23_n835 ), .A2(_AES_ENC_us23_n834 ), .A3(_AES_ENC_us23_n833 ), .A4(_AES_ENC_us23_n832 ), .ZN(_AES_ENC_us23_n836 ) );
NAND2_X2 _AES_ENC_us23_U232  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n836 ), .ZN(_AES_ENC_us23_n850 ) );
NAND2_X2 _AES_ENC_us23_U231  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n601 ), .ZN(_AES_ENC_us23_n847 ) );
NAND2_X2 _AES_ENC_us23_U230  ( .A1(_AES_ENC_us23_n1050 ), .A2(_AES_ENC_us23_n1071 ), .ZN(_AES_ENC_us23_n846 ) );
OR2_X2 _AES_ENC_us23_U224  ( .A1(_AES_ENC_us23_n1053 ), .A2(_AES_ENC_us23_n911 ), .ZN(_AES_ENC_us23_n1077 ) );
NAND4_X2 _AES_ENC_us23_U220  ( .A1(_AES_ENC_us23_n847 ), .A2(_AES_ENC_us23_n846 ), .A3(_AES_ENC_us23_n845 ), .A4(_AES_ENC_us23_n844 ), .ZN(_AES_ENC_us23_n848 ) );
NAND2_X2 _AES_ENC_us23_U219  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n848 ), .ZN(_AES_ENC_us23_n849 ) );
NAND4_X2 _AES_ENC_us23_U218  ( .A1(_AES_ENC_us23_n852 ), .A2(_AES_ENC_us23_n851 ), .A3(_AES_ENC_us23_n850 ), .A4(_AES_ENC_us23_n849 ), .ZN(_AES_ENC_sa23_sub[3] ) );
NAND2_X2 _AES_ENC_us23_U216  ( .A1(_AES_ENC_us23_n1009 ), .A2(_AES_ENC_us23_n1072 ), .ZN(_AES_ENC_us23_n862 ) );
NAND2_X2 _AES_ENC_us23_U215  ( .A1(_AES_ENC_us23_n610 ), .A2(_AES_ENC_us23_n618 ), .ZN(_AES_ENC_us23_n853 ) );
NAND2_X2 _AES_ENC_us23_U214  ( .A1(_AES_ENC_us23_n1050 ), .A2(_AES_ENC_us23_n853 ), .ZN(_AES_ENC_us23_n861 ) );
NAND4_X2 _AES_ENC_us23_U206  ( .A1(_AES_ENC_us23_n862 ), .A2(_AES_ENC_us23_n861 ), .A3(_AES_ENC_us23_n860 ), .A4(_AES_ENC_us23_n859 ), .ZN(_AES_ENC_us23_n863 ) );
NAND2_X2 _AES_ENC_us23_U205  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n863 ), .ZN(_AES_ENC_us23_n905 ) );
NAND2_X2 _AES_ENC_us23_U204  ( .A1(_AES_ENC_us23_n1010 ), .A2(_AES_ENC_us23_n989 ), .ZN(_AES_ENC_us23_n874 ) );
NAND2_X2 _AES_ENC_us23_U203  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n592 ), .ZN(_AES_ENC_us23_n864 ) );
NAND2_X2 _AES_ENC_us23_U202  ( .A1(_AES_ENC_us23_n929 ), .A2(_AES_ENC_us23_n864 ), .ZN(_AES_ENC_us23_n873 ) );
NAND4_X2 _AES_ENC_us23_U193  ( .A1(_AES_ENC_us23_n874 ), .A2(_AES_ENC_us23_n873 ), .A3(_AES_ENC_us23_n872 ), .A4(_AES_ENC_us23_n871 ), .ZN(_AES_ENC_us23_n875 ) );
NAND2_X2 _AES_ENC_us23_U192  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n875 ), .ZN(_AES_ENC_us23_n904 ) );
NAND2_X2 _AES_ENC_us23_U191  ( .A1(_AES_ENC_us23_n597 ), .A2(_AES_ENC_us23_n1050 ), .ZN(_AES_ENC_us23_n889 ) );
NAND2_X2 _AES_ENC_us23_U190  ( .A1(_AES_ENC_us23_n1093 ), .A2(_AES_ENC_us23_n617 ), .ZN(_AES_ENC_us23_n876 ) );
NAND2_X2 _AES_ENC_us23_U189  ( .A1(_AES_ENC_us23_n576 ), .A2(_AES_ENC_us23_n876 ), .ZN(_AES_ENC_us23_n877 ) );
NAND2_X2 _AES_ENC_us23_U188  ( .A1(_AES_ENC_us23_n877 ), .A2(_AES_ENC_us23_n601 ), .ZN(_AES_ENC_us23_n888 ) );
NAND4_X2 _AES_ENC_us23_U179  ( .A1(_AES_ENC_us23_n889 ), .A2(_AES_ENC_us23_n888 ), .A3(_AES_ENC_us23_n887 ), .A4(_AES_ENC_us23_n886 ), .ZN(_AES_ENC_us23_n890 ) );
NAND2_X2 _AES_ENC_us23_U178  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n890 ), .ZN(_AES_ENC_us23_n903 ) );
OR2_X2 _AES_ENC_us23_U177  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n1059 ), .ZN(_AES_ENC_us23_n900 ) );
NAND2_X2 _AES_ENC_us23_U176  ( .A1(_AES_ENC_us23_n1073 ), .A2(_AES_ENC_us23_n1047 ), .ZN(_AES_ENC_us23_n899 ) );
NAND2_X2 _AES_ENC_us23_U175  ( .A1(_AES_ENC_us23_n1094 ), .A2(_AES_ENC_us23_n608 ), .ZN(_AES_ENC_us23_n898 ) );
NAND4_X2 _AES_ENC_us23_U167  ( .A1(_AES_ENC_us23_n900 ), .A2(_AES_ENC_us23_n899 ), .A3(_AES_ENC_us23_n898 ), .A4(_AES_ENC_us23_n897 ), .ZN(_AES_ENC_us23_n901 ) );
NAND2_X2 _AES_ENC_us23_U166  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n901 ), .ZN(_AES_ENC_us23_n902 ) );
NAND4_X2 _AES_ENC_us23_U165  ( .A1(_AES_ENC_us23_n905 ), .A2(_AES_ENC_us23_n904 ), .A3(_AES_ENC_us23_n903 ), .A4(_AES_ENC_us23_n902 ), .ZN(_AES_ENC_sa23_sub[4] ) );
NAND2_X2 _AES_ENC_us23_U164  ( .A1(_AES_ENC_us23_n1094 ), .A2(_AES_ENC_us23_n615 ), .ZN(_AES_ENC_us23_n922 ) );
NAND2_X2 _AES_ENC_us23_U163  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n989 ), .ZN(_AES_ENC_us23_n921 ) );
NAND4_X2 _AES_ENC_us23_U151  ( .A1(_AES_ENC_us23_n922 ), .A2(_AES_ENC_us23_n921 ), .A3(_AES_ENC_us23_n920 ), .A4(_AES_ENC_us23_n919 ), .ZN(_AES_ENC_us23_n923 ) );
NAND2_X2 _AES_ENC_us23_U150  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n923 ), .ZN(_AES_ENC_us23_n972 ) );
NAND2_X2 _AES_ENC_us23_U149  ( .A1(_AES_ENC_us23_n603 ), .A2(_AES_ENC_us23_n605 ), .ZN(_AES_ENC_us23_n924 ) );
NAND2_X2 _AES_ENC_us23_U148  ( .A1(_AES_ENC_us23_n1073 ), .A2(_AES_ENC_us23_n924 ), .ZN(_AES_ENC_us23_n939 ) );
NAND2_X2 _AES_ENC_us23_U147  ( .A1(_AES_ENC_us23_n926 ), .A2(_AES_ENC_us23_n925 ), .ZN(_AES_ENC_us23_n927 ) );
NAND2_X2 _AES_ENC_us23_U146  ( .A1(_AES_ENC_us23_n587 ), .A2(_AES_ENC_us23_n927 ), .ZN(_AES_ENC_us23_n928 ) );
NAND2_X2 _AES_ENC_us23_U145  ( .A1(_AES_ENC_us23_n928 ), .A2(_AES_ENC_us23_n1080 ), .ZN(_AES_ENC_us23_n938 ) );
OR2_X2 _AES_ENC_us23_U144  ( .A1(_AES_ENC_us23_n1117 ), .A2(_AES_ENC_us23_n580 ), .ZN(_AES_ENC_us23_n937 ) );
NAND4_X2 _AES_ENC_us23_U139  ( .A1(_AES_ENC_us23_n939 ), .A2(_AES_ENC_us23_n938 ), .A3(_AES_ENC_us23_n937 ), .A4(_AES_ENC_us23_n936 ), .ZN(_AES_ENC_us23_n940 ) );
NAND2_X2 _AES_ENC_us23_U138  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n940 ), .ZN(_AES_ENC_us23_n971 ) );
OR2_X2 _AES_ENC_us23_U137  ( .A1(_AES_ENC_us23_n586 ), .A2(_AES_ENC_us23_n941 ), .ZN(_AES_ENC_us23_n954 ) );
NAND2_X2 _AES_ENC_us23_U136  ( .A1(_AES_ENC_us23_n1096 ), .A2(_AES_ENC_us23_n618 ), .ZN(_AES_ENC_us23_n942 ) );
NAND2_X2 _AES_ENC_us23_U135  ( .A1(_AES_ENC_us23_n1048 ), .A2(_AES_ENC_us23_n942 ), .ZN(_AES_ENC_us23_n943 ) );
NAND2_X2 _AES_ENC_us23_U134  ( .A1(_AES_ENC_us23_n582 ), .A2(_AES_ENC_us23_n943 ), .ZN(_AES_ENC_us23_n944 ) );
NAND2_X2 _AES_ENC_us23_U133  ( .A1(_AES_ENC_us23_n944 ), .A2(_AES_ENC_us23_n599 ), .ZN(_AES_ENC_us23_n953 ) );
NAND4_X2 _AES_ENC_us23_U125  ( .A1(_AES_ENC_us23_n954 ), .A2(_AES_ENC_us23_n953 ), .A3(_AES_ENC_us23_n952 ), .A4(_AES_ENC_us23_n951 ), .ZN(_AES_ENC_us23_n955 ) );
NAND2_X2 _AES_ENC_us23_U124  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n955 ), .ZN(_AES_ENC_us23_n970 ) );
NAND2_X2 _AES_ENC_us23_U123  ( .A1(_AES_ENC_us23_n1094 ), .A2(_AES_ENC_us23_n1071 ), .ZN(_AES_ENC_us23_n967 ) );
NAND2_X2 _AES_ENC_us23_U122  ( .A1(_AES_ENC_us23_n956 ), .A2(_AES_ENC_us23_n1030 ), .ZN(_AES_ENC_us23_n966 ) );
NAND4_X2 _AES_ENC_us23_U114  ( .A1(_AES_ENC_us23_n967 ), .A2(_AES_ENC_us23_n966 ), .A3(_AES_ENC_us23_n965 ), .A4(_AES_ENC_us23_n964 ), .ZN(_AES_ENC_us23_n968 ) );
NAND2_X2 _AES_ENC_us23_U113  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n968 ), .ZN(_AES_ENC_us23_n969 ) );
NAND4_X2 _AES_ENC_us23_U112  ( .A1(_AES_ENC_us23_n972 ), .A2(_AES_ENC_us23_n971 ), .A3(_AES_ENC_us23_n970 ), .A4(_AES_ENC_us23_n969 ), .ZN(_AES_ENC_sa23_sub[5] ) );
NAND2_X2 _AES_ENC_us23_U111  ( .A1(_AES_ENC_us23_n570 ), .A2(_AES_ENC_us23_n1097 ), .ZN(_AES_ENC_us23_n973 ) );
NAND2_X2 _AES_ENC_us23_U110  ( .A1(_AES_ENC_us23_n1073 ), .A2(_AES_ENC_us23_n973 ), .ZN(_AES_ENC_us23_n987 ) );
NAND2_X2 _AES_ENC_us23_U109  ( .A1(_AES_ENC_us23_n974 ), .A2(_AES_ENC_us23_n1077 ), .ZN(_AES_ENC_us23_n975 ) );
NAND2_X2 _AES_ENC_us23_U108  ( .A1(_AES_ENC_us23_n584 ), .A2(_AES_ENC_us23_n975 ), .ZN(_AES_ENC_us23_n976 ) );
NAND2_X2 _AES_ENC_us23_U107  ( .A1(_AES_ENC_us23_n977 ), .A2(_AES_ENC_us23_n976 ), .ZN(_AES_ENC_us23_n986 ) );
NAND4_X2 _AES_ENC_us23_U99  ( .A1(_AES_ENC_us23_n987 ), .A2(_AES_ENC_us23_n986 ), .A3(_AES_ENC_us23_n985 ), .A4(_AES_ENC_us23_n984 ), .ZN(_AES_ENC_us23_n988 ) );
NAND2_X2 _AES_ENC_us23_U98  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n988 ), .ZN(_AES_ENC_us23_n1044 ) );
NAND2_X2 _AES_ENC_us23_U97  ( .A1(_AES_ENC_us23_n1073 ), .A2(_AES_ENC_us23_n989 ), .ZN(_AES_ENC_us23_n1004 ) );
NAND2_X2 _AES_ENC_us23_U96  ( .A1(_AES_ENC_us23_n1092 ), .A2(_AES_ENC_us23_n605 ), .ZN(_AES_ENC_us23_n1003 ) );
NAND4_X2 _AES_ENC_us23_U85  ( .A1(_AES_ENC_us23_n1004 ), .A2(_AES_ENC_us23_n1003 ), .A3(_AES_ENC_us23_n1002 ), .A4(_AES_ENC_us23_n1001 ), .ZN(_AES_ENC_us23_n1005 ) );
NAND2_X2 _AES_ENC_us23_U84  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n1005 ), .ZN(_AES_ENC_us23_n1043 ) );
NAND2_X2 _AES_ENC_us23_U83  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n626 ), .ZN(_AES_ENC_us23_n1020 ) );
NAND2_X2 _AES_ENC_us23_U82  ( .A1(_AES_ENC_us23_n1050 ), .A2(_AES_ENC_us23_n612 ), .ZN(_AES_ENC_us23_n1019 ) );
NAND2_X2 _AES_ENC_us23_U77  ( .A1(_AES_ENC_us23_n1059 ), .A2(_AES_ENC_us23_n1114 ), .ZN(_AES_ENC_us23_n1012 ) );
NAND2_X2 _AES_ENC_us23_U76  ( .A1(_AES_ENC_us23_n1010 ), .A2(_AES_ENC_us23_n604 ), .ZN(_AES_ENC_us23_n1011 ) );
NAND2_X2 _AES_ENC_us23_U75  ( .A1(_AES_ENC_us23_n1012 ), .A2(_AES_ENC_us23_n1011 ), .ZN(_AES_ENC_us23_n1016 ) );
NAND4_X2 _AES_ENC_us23_U70  ( .A1(_AES_ENC_us23_n1020 ), .A2(_AES_ENC_us23_n1019 ), .A3(_AES_ENC_us23_n1018 ), .A4(_AES_ENC_us23_n1017 ), .ZN(_AES_ENC_us23_n1021 ) );
NAND2_X2 _AES_ENC_us23_U69  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n1021 ), .ZN(_AES_ENC_us23_n1042 ) );
NAND2_X2 _AES_ENC_us23_U68  ( .A1(_AES_ENC_us23_n1022 ), .A2(_AES_ENC_us23_n1093 ), .ZN(_AES_ENC_us23_n1039 ) );
NAND2_X2 _AES_ENC_us23_U67  ( .A1(_AES_ENC_us23_n1050 ), .A2(_AES_ENC_us23_n1023 ), .ZN(_AES_ENC_us23_n1038 ) );
NAND2_X2 _AES_ENC_us23_U66  ( .A1(_AES_ENC_us23_n1024 ), .A2(_AES_ENC_us23_n1071 ), .ZN(_AES_ENC_us23_n1037 ) );
AND2_X2 _AES_ENC_us23_U60  ( .A1(_AES_ENC_us23_n1030 ), .A2(_AES_ENC_us23_n621 ), .ZN(_AES_ENC_us23_n1078 ) );
NAND4_X2 _AES_ENC_us23_U56  ( .A1(_AES_ENC_us23_n1039 ), .A2(_AES_ENC_us23_n1038 ), .A3(_AES_ENC_us23_n1037 ), .A4(_AES_ENC_us23_n1036 ), .ZN(_AES_ENC_us23_n1040 ) );
NAND2_X2 _AES_ENC_us23_U55  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n1040 ), .ZN(_AES_ENC_us23_n1041 ) );
NAND4_X2 _AES_ENC_us23_U54  ( .A1(_AES_ENC_us23_n1044 ), .A2(_AES_ENC_us23_n1043 ), .A3(_AES_ENC_us23_n1042 ), .A4(_AES_ENC_us23_n1041 ), .ZN(_AES_ENC_sa23_sub[6] ) );
NAND2_X2 _AES_ENC_us23_U53  ( .A1(_AES_ENC_us23_n1072 ), .A2(_AES_ENC_us23_n1045 ), .ZN(_AES_ENC_us23_n1068 ) );
NAND2_X2 _AES_ENC_us23_U52  ( .A1(_AES_ENC_us23_n1046 ), .A2(_AES_ENC_us23_n603 ), .ZN(_AES_ENC_us23_n1067 ) );
NAND2_X2 _AES_ENC_us23_U51  ( .A1(_AES_ENC_us23_n1094 ), .A2(_AES_ENC_us23_n1047 ), .ZN(_AES_ENC_us23_n1066 ) );
NAND4_X2 _AES_ENC_us23_U40  ( .A1(_AES_ENC_us23_n1068 ), .A2(_AES_ENC_us23_n1067 ), .A3(_AES_ENC_us23_n1066 ), .A4(_AES_ENC_us23_n1065 ), .ZN(_AES_ENC_us23_n1069 ) );
NAND2_X2 _AES_ENC_us23_U39  ( .A1(_AES_ENC_us23_n1070 ), .A2(_AES_ENC_us23_n1069 ), .ZN(_AES_ENC_us23_n1135 ) );
NAND2_X2 _AES_ENC_us23_U38  ( .A1(_AES_ENC_us23_n1072 ), .A2(_AES_ENC_us23_n1071 ), .ZN(_AES_ENC_us23_n1088 ) );
NAND2_X2 _AES_ENC_us23_U37  ( .A1(_AES_ENC_us23_n1073 ), .A2(_AES_ENC_us23_n608 ), .ZN(_AES_ENC_us23_n1087 ) );
NAND4_X2 _AES_ENC_us23_U28  ( .A1(_AES_ENC_us23_n1088 ), .A2(_AES_ENC_us23_n1087 ), .A3(_AES_ENC_us23_n1086 ), .A4(_AES_ENC_us23_n1085 ), .ZN(_AES_ENC_us23_n1089 ) );
NAND2_X2 _AES_ENC_us23_U27  ( .A1(_AES_ENC_us23_n1090 ), .A2(_AES_ENC_us23_n1089 ), .ZN(_AES_ENC_us23_n1134 ) );
NAND2_X2 _AES_ENC_us23_U26  ( .A1(_AES_ENC_us23_n1091 ), .A2(_AES_ENC_us23_n1093 ), .ZN(_AES_ENC_us23_n1111 ) );
NAND2_X2 _AES_ENC_us23_U25  ( .A1(_AES_ENC_us23_n1092 ), .A2(_AES_ENC_us23_n1120 ), .ZN(_AES_ENC_us23_n1110 ) );
AND2_X2 _AES_ENC_us23_U22  ( .A1(_AES_ENC_us23_n1097 ), .A2(_AES_ENC_us23_n1096 ), .ZN(_AES_ENC_us23_n1098 ) );
NAND4_X2 _AES_ENC_us23_U14  ( .A1(_AES_ENC_us23_n1111 ), .A2(_AES_ENC_us23_n1110 ), .A3(_AES_ENC_us23_n1109 ), .A4(_AES_ENC_us23_n1108 ), .ZN(_AES_ENC_us23_n1112 ) );
NAND2_X2 _AES_ENC_us23_U13  ( .A1(_AES_ENC_us23_n1113 ), .A2(_AES_ENC_us23_n1112 ), .ZN(_AES_ENC_us23_n1133 ) );
NAND2_X2 _AES_ENC_us23_U12  ( .A1(_AES_ENC_us23_n1115 ), .A2(_AES_ENC_us23_n1114 ), .ZN(_AES_ENC_us23_n1129 ) );
OR2_X2 _AES_ENC_us23_U11  ( .A1(_AES_ENC_us23_n579 ), .A2(_AES_ENC_us23_n1116 ), .ZN(_AES_ENC_us23_n1128 ) );
NAND4_X2 _AES_ENC_us23_U3  ( .A1(_AES_ENC_us23_n1129 ), .A2(_AES_ENC_us23_n1128 ), .A3(_AES_ENC_us23_n1127 ), .A4(_AES_ENC_us23_n1126 ), .ZN(_AES_ENC_us23_n1130 ) );
NAND2_X2 _AES_ENC_us23_U2  ( .A1(_AES_ENC_us23_n1131 ), .A2(_AES_ENC_us23_n1130 ), .ZN(_AES_ENC_us23_n1132 ) );
NAND4_X2 _AES_ENC_us23_U1  ( .A1(_AES_ENC_us23_n1135 ), .A2(_AES_ENC_us23_n1134 ), .A3(_AES_ENC_us23_n1133 ), .A4(_AES_ENC_us23_n1132 ), .ZN(_AES_ENC_sa23_sub[7] ) );
INV_X4 _AES_ENC_us30_U575  ( .A(_AES_ENC_sa30[7]), .ZN(_AES_ENC_us30_n627 ));
INV_X4 _AES_ENC_us30_U574  ( .A(_AES_ENC_us30_n1114 ), .ZN(_AES_ENC_us30_n625 ) );
INV_X4 _AES_ENC_us30_U573  ( .A(_AES_ENC_sa30[4]), .ZN(_AES_ENC_us30_n624 ));
INV_X4 _AES_ENC_us30_U572  ( .A(_AES_ENC_us30_n1025 ), .ZN(_AES_ENC_us30_n622 ) );
INV_X4 _AES_ENC_us30_U571  ( .A(_AES_ENC_us30_n1120 ), .ZN(_AES_ENC_us30_n620 ) );
INV_X4 _AES_ENC_us30_U570  ( .A(_AES_ENC_us30_n1121 ), .ZN(_AES_ENC_us30_n619 ) );
INV_X4 _AES_ENC_us30_U569  ( .A(_AES_ENC_us30_n1048 ), .ZN(_AES_ENC_us30_n618 ) );
INV_X4 _AES_ENC_us30_U568  ( .A(_AES_ENC_us30_n974 ), .ZN(_AES_ENC_us30_n616 ) );
INV_X4 _AES_ENC_us30_U567  ( .A(_AES_ENC_us30_n794 ), .ZN(_AES_ENC_us30_n614 ) );
INV_X4 _AES_ENC_us30_U566  ( .A(_AES_ENC_sa30[2]), .ZN(_AES_ENC_us30_n611 ));
INV_X4 _AES_ENC_us30_U565  ( .A(_AES_ENC_us30_n800 ), .ZN(_AES_ENC_us30_n610 ) );
INV_X4 _AES_ENC_us30_U564  ( .A(_AES_ENC_us30_n925 ), .ZN(_AES_ENC_us30_n609 ) );
INV_X4 _AES_ENC_us30_U563  ( .A(_AES_ENC_us30_n779 ), .ZN(_AES_ENC_us30_n607 ) );
INV_X4 _AES_ENC_us30_U562  ( .A(_AES_ENC_us30_n1022 ), .ZN(_AES_ENC_us30_n603 ) );
INV_X4 _AES_ENC_us30_U561  ( .A(_AES_ENC_us30_n1102 ), .ZN(_AES_ENC_us30_n602 ) );
INV_X4 _AES_ENC_us30_U560  ( .A(_AES_ENC_us30_n929 ), .ZN(_AES_ENC_us30_n601 ) );
INV_X4 _AES_ENC_us30_U559  ( .A(_AES_ENC_us30_n1056 ), .ZN(_AES_ENC_us30_n600 ) );
INV_X4 _AES_ENC_us30_U558  ( .A(_AES_ENC_us30_n1054 ), .ZN(_AES_ENC_us30_n599 ) );
INV_X4 _AES_ENC_us30_U557  ( .A(_AES_ENC_us30_n881 ), .ZN(_AES_ENC_us30_n598 ) );
INV_X4 _AES_ENC_us30_U556  ( .A(_AES_ENC_us30_n926 ), .ZN(_AES_ENC_us30_n597 ) );
INV_X4 _AES_ENC_us30_U555  ( .A(_AES_ENC_us30_n977 ), .ZN(_AES_ENC_us30_n595 ) );
INV_X4 _AES_ENC_us30_U554  ( .A(_AES_ENC_us30_n1031 ), .ZN(_AES_ENC_us30_n594 ) );
INV_X4 _AES_ENC_us30_U553  ( .A(_AES_ENC_us30_n1103 ), .ZN(_AES_ENC_us30_n593 ) );
INV_X4 _AES_ENC_us30_U552  ( .A(_AES_ENC_us30_n1009 ), .ZN(_AES_ENC_us30_n592 ) );
INV_X4 _AES_ENC_us30_U551  ( .A(_AES_ENC_us30_n990 ), .ZN(_AES_ENC_us30_n591 ) );
INV_X4 _AES_ENC_us30_U550  ( .A(_AES_ENC_us30_n1058 ), .ZN(_AES_ENC_us30_n590 ) );
INV_X4 _AES_ENC_us30_U549  ( .A(_AES_ENC_us30_n1074 ), .ZN(_AES_ENC_us30_n589 ) );
INV_X4 _AES_ENC_us30_U548  ( .A(_AES_ENC_us30_n1053 ), .ZN(_AES_ENC_us30_n588 ) );
INV_X4 _AES_ENC_us30_U547  ( .A(_AES_ENC_us30_n826 ), .ZN(_AES_ENC_us30_n587 ) );
INV_X4 _AES_ENC_us30_U546  ( .A(_AES_ENC_us30_n992 ), .ZN(_AES_ENC_us30_n586 ) );
INV_X4 _AES_ENC_us30_U545  ( .A(_AES_ENC_us30_n821 ), .ZN(_AES_ENC_us30_n585 ) );
INV_X4 _AES_ENC_us30_U544  ( .A(_AES_ENC_us30_n910 ), .ZN(_AES_ENC_us30_n584 ) );
INV_X4 _AES_ENC_us30_U543  ( .A(_AES_ENC_us30_n906 ), .ZN(_AES_ENC_us30_n583 ) );
INV_X4 _AES_ENC_us30_U542  ( .A(_AES_ENC_us30_n880 ), .ZN(_AES_ENC_us30_n581 ) );
INV_X4 _AES_ENC_us30_U541  ( .A(_AES_ENC_us30_n1013 ), .ZN(_AES_ENC_us30_n580 ) );
INV_X4 _AES_ENC_us30_U540  ( .A(_AES_ENC_us30_n1092 ), .ZN(_AES_ENC_us30_n579 ) );
INV_X4 _AES_ENC_us30_U539  ( .A(_AES_ENC_us30_n824 ), .ZN(_AES_ENC_us30_n578 ) );
INV_X4 _AES_ENC_us30_U538  ( .A(_AES_ENC_us30_n1091 ), .ZN(_AES_ENC_us30_n577 ) );
INV_X4 _AES_ENC_us30_U537  ( .A(_AES_ENC_us30_n1080 ), .ZN(_AES_ENC_us30_n576 ) );
INV_X4 _AES_ENC_us30_U536  ( .A(_AES_ENC_us30_n959 ), .ZN(_AES_ENC_us30_n575 ) );
INV_X4 _AES_ENC_us30_U535  ( .A(_AES_ENC_sa30[0]), .ZN(_AES_ENC_us30_n574 ));
NOR2_X2 _AES_ENC_us30_U534  ( .A1(_AES_ENC_us30_n574 ), .A2(_AES_ENC_sa30[6]), .ZN(_AES_ENC_us30_n1070 ) );
NOR2_X2 _AES_ENC_us30_U533  ( .A1(_AES_ENC_sa30[0]), .A2(_AES_ENC_sa30[6]),.ZN(_AES_ENC_us30_n1090 ) );
NOR2_X2 _AES_ENC_us30_U532  ( .A1(_AES_ENC_sa30[4]), .A2(_AES_ENC_sa30[3]),.ZN(_AES_ENC_us30_n1025 ) );
INV_X4 _AES_ENC_us30_U531  ( .A(_AES_ENC_us30_n569 ), .ZN(_AES_ENC_us30_n572 ) );
NOR2_X2 _AES_ENC_us30_U530  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n765 ) );
NOR2_X2 _AES_ENC_us30_U529  ( .A1(_AES_ENC_sa30[4]), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n764 ) );
NOR2_X2 _AES_ENC_us30_U528  ( .A1(_AES_ENC_us30_n765 ), .A2(_AES_ENC_us30_n764 ), .ZN(_AES_ENC_us30_n766 ) );
NOR2_X2 _AES_ENC_us30_U527  ( .A1(_AES_ENC_us30_n766 ), .A2(_AES_ENC_us30_n575 ), .ZN(_AES_ENC_us30_n767 ) );
NOR3_X2 _AES_ENC_us30_U526  ( .A1(_AES_ENC_us30_n627 ), .A2(_AES_ENC_sa30[5]), .A3(_AES_ENC_us30_n704 ), .ZN(_AES_ENC_us30_n706 ));
NOR2_X2 _AES_ENC_us30_U525  ( .A1(_AES_ENC_us30_n1117 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n707 ) );
NOR2_X2 _AES_ENC_us30_U524  ( .A1(_AES_ENC_sa30[4]), .A2(_AES_ENC_us30_n579 ), .ZN(_AES_ENC_us30_n705 ) );
NOR3_X2 _AES_ENC_us30_U523  ( .A1(_AES_ENC_us30_n707 ), .A2(_AES_ENC_us30_n706 ), .A3(_AES_ENC_us30_n705 ), .ZN(_AES_ENC_us30_n713 ) );
INV_X4 _AES_ENC_us30_U522  ( .A(_AES_ENC_sa30[3]), .ZN(_AES_ENC_us30_n621 ));
NAND3_X2 _AES_ENC_us30_U521  ( .A1(_AES_ENC_us30_n652 ), .A2(_AES_ENC_us30_n626 ), .A3(_AES_ENC_sa30[7]), .ZN(_AES_ENC_us30_n653 ));
NOR2_X2 _AES_ENC_us30_U520  ( .A1(_AES_ENC_us30_n611 ), .A2(_AES_ENC_sa30[5]), .ZN(_AES_ENC_us30_n925 ) );
NOR2_X2 _AES_ENC_us30_U519  ( .A1(_AES_ENC_sa30[5]), .A2(_AES_ENC_sa30[2]),.ZN(_AES_ENC_us30_n974 ) );
INV_X4 _AES_ENC_us30_U518  ( .A(_AES_ENC_sa30[5]), .ZN(_AES_ENC_us30_n626 ));
NOR2_X2 _AES_ENC_us30_U517  ( .A1(_AES_ENC_us30_n611 ), .A2(_AES_ENC_sa30[7]), .ZN(_AES_ENC_us30_n779 ) );
NAND3_X2 _AES_ENC_us30_U516  ( .A1(_AES_ENC_us30_n679 ), .A2(_AES_ENC_us30_n678 ), .A3(_AES_ENC_us30_n677 ), .ZN(_AES_ENC_sa30_sub[0] ) );
NOR2_X2 _AES_ENC_us30_U515  ( .A1(_AES_ENC_us30_n626 ), .A2(_AES_ENC_sa30[2]), .ZN(_AES_ENC_us30_n1048 ) );
NOR4_X2 _AES_ENC_us30_U512  ( .A1(_AES_ENC_us30_n633 ), .A2(_AES_ENC_us30_n632 ), .A3(_AES_ENC_us30_n631 ), .A4(_AES_ENC_us30_n630 ), .ZN(_AES_ENC_us30_n634 ) );
NOR2_X2 _AES_ENC_us30_U510  ( .A1(_AES_ENC_us30_n629 ), .A2(_AES_ENC_us30_n628 ), .ZN(_AES_ENC_us30_n635 ) );
NAND3_X2 _AES_ENC_us30_U509  ( .A1(_AES_ENC_sa30[2]), .A2(_AES_ENC_sa30[7]), .A3(_AES_ENC_us30_n1059 ), .ZN(_AES_ENC_us30_n636 ) );
NOR2_X2 _AES_ENC_us30_U508  ( .A1(_AES_ENC_sa30[7]), .A2(_AES_ENC_sa30[2]),.ZN(_AES_ENC_us30_n794 ) );
NOR2_X2 _AES_ENC_us30_U507  ( .A1(_AES_ENC_sa30[4]), .A2(_AES_ENC_sa30[1]),.ZN(_AES_ENC_us30_n1102 ) );
NOR2_X2 _AES_ENC_us30_U506  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_sa30[3]), .ZN(_AES_ENC_us30_n1053 ) );
NOR2_X2 _AES_ENC_us30_U505  ( .A1(_AES_ENC_us30_n607 ), .A2(_AES_ENC_sa30[5]), .ZN(_AES_ENC_us30_n1024 ) );
NOR2_X2 _AES_ENC_us30_U504  ( .A1(_AES_ENC_us30_n625 ), .A2(_AES_ENC_sa30[2]), .ZN(_AES_ENC_us30_n1093 ) );
NOR2_X2 _AES_ENC_us30_U503  ( .A1(_AES_ENC_us30_n614 ), .A2(_AES_ENC_sa30[5]), .ZN(_AES_ENC_us30_n1094 ) );
NOR2_X2 _AES_ENC_us30_U502  ( .A1(_AES_ENC_us30_n624 ), .A2(_AES_ENC_sa30[3]), .ZN(_AES_ENC_us30_n931 ) );
INV_X4 _AES_ENC_us30_U501  ( .A(_AES_ENC_us30_n570 ), .ZN(_AES_ENC_us30_n573 ) );
NOR2_X2 _AES_ENC_us30_U500  ( .A1(_AES_ENC_us30_n1053 ), .A2(_AES_ENC_us30_n1095 ), .ZN(_AES_ENC_us30_n639 ) );
NOR3_X2 _AES_ENC_us30_U499  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n573 ), .A3(_AES_ENC_us30_n1074 ), .ZN(_AES_ENC_us30_n641 ) );
NOR2_X2 _AES_ENC_us30_U498  ( .A1(_AES_ENC_us30_n639 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n640 ) );
NOR2_X2 _AES_ENC_us30_U497  ( .A1(_AES_ENC_us30_n641 ), .A2(_AES_ENC_us30_n640 ), .ZN(_AES_ENC_us30_n646 ) );
NOR3_X2 _AES_ENC_us30_U496  ( .A1(_AES_ENC_us30_n995 ), .A2(_AES_ENC_us30_n586 ), .A3(_AES_ENC_us30_n994 ), .ZN(_AES_ENC_us30_n1002 ) );
NOR2_X2 _AES_ENC_us30_U495  ( .A1(_AES_ENC_us30_n909 ), .A2(_AES_ENC_us30_n908 ), .ZN(_AES_ENC_us30_n920 ) );
NOR2_X2 _AES_ENC_us30_U494  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n823 ) );
NOR2_X2 _AES_ENC_us30_U492  ( .A1(_AES_ENC_us30_n624 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n822 ) );
NOR2_X2 _AES_ENC_us30_U491  ( .A1(_AES_ENC_us30_n823 ), .A2(_AES_ENC_us30_n822 ), .ZN(_AES_ENC_us30_n825 ) );
NOR2_X2 _AES_ENC_us30_U490  ( .A1(_AES_ENC_sa30[1]), .A2(_AES_ENC_us30_n623 ), .ZN(_AES_ENC_us30_n913 ) );
NOR2_X2 _AES_ENC_us30_U489  ( .A1(_AES_ENC_us30_n913 ), .A2(_AES_ENC_us30_n1091 ), .ZN(_AES_ENC_us30_n914 ) );
NOR2_X2 _AES_ENC_us30_U488  ( .A1(_AES_ENC_us30_n826 ), .A2(_AES_ENC_us30_n572 ), .ZN(_AES_ENC_us30_n827 ) );
NOR3_X2 _AES_ENC_us30_U487  ( .A1(_AES_ENC_us30_n769 ), .A2(_AES_ENC_us30_n768 ), .A3(_AES_ENC_us30_n767 ), .ZN(_AES_ENC_us30_n775 ) );
NOR2_X2 _AES_ENC_us30_U486  ( .A1(_AES_ENC_us30_n1056 ), .A2(_AES_ENC_us30_n1053 ), .ZN(_AES_ENC_us30_n749 ) );
NOR2_X2 _AES_ENC_us30_U483  ( .A1(_AES_ENC_us30_n749 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n752 ) );
INV_X4 _AES_ENC_us30_U482  ( .A(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n596 ));
NOR2_X2 _AES_ENC_us30_U480  ( .A1(_AES_ENC_us30_n1054 ), .A2(_AES_ENC_us30_n1053 ), .ZN(_AES_ENC_us30_n1055 ) );
OR2_X4 _AES_ENC_us30_U479  ( .A1(_AES_ENC_us30_n1094 ), .A2(_AES_ENC_us30_n1093 ), .ZN(_AES_ENC_us30_n571 ) );
AND2_X2 _AES_ENC_us30_U478  ( .A1(_AES_ENC_us30_n571 ), .A2(_AES_ENC_us30_n1095 ), .ZN(_AES_ENC_us30_n1101 ) );
NOR2_X2 _AES_ENC_us30_U477  ( .A1(_AES_ENC_us30_n1074 ), .A2(_AES_ENC_us30_n931 ), .ZN(_AES_ENC_us30_n796 ) );
NOR2_X2 _AES_ENC_us30_U474  ( .A1(_AES_ENC_us30_n796 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n797 ) );
NOR2_X2 _AES_ENC_us30_U473  ( .A1(_AES_ENC_us30_n932 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n933 ) );
NOR2_X2 _AES_ENC_us30_U472  ( .A1(_AES_ENC_us30_n929 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n935 ) );
NOR2_X2 _AES_ENC_us30_U471  ( .A1(_AES_ENC_us30_n931 ), .A2(_AES_ENC_us30_n930 ), .ZN(_AES_ENC_us30_n934 ) );
NOR3_X2 _AES_ENC_us30_U470  ( .A1(_AES_ENC_us30_n935 ), .A2(_AES_ENC_us30_n934 ), .A3(_AES_ENC_us30_n933 ), .ZN(_AES_ENC_us30_n936 ) );
NOR2_X2 _AES_ENC_us30_U469  ( .A1(_AES_ENC_us30_n624 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n1075 ) );
NOR2_X2 _AES_ENC_us30_U468  ( .A1(_AES_ENC_us30_n572 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n949 ) );
NOR2_X2 _AES_ENC_us30_U467  ( .A1(_AES_ENC_us30_n1049 ), .A2(_AES_ENC_us30_n618 ), .ZN(_AES_ENC_us30_n1051 ) );
NOR2_X2 _AES_ENC_us30_U466  ( .A1(_AES_ENC_us30_n1051 ), .A2(_AES_ENC_us30_n1050 ), .ZN(_AES_ENC_us30_n1052 ) );
NOR2_X2 _AES_ENC_us30_U465  ( .A1(_AES_ENC_us30_n1052 ), .A2(_AES_ENC_us30_n592 ), .ZN(_AES_ENC_us30_n1064 ) );
NOR2_X2 _AES_ENC_us30_U464  ( .A1(_AES_ENC_sa30[1]), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n631 ) );
NOR2_X2 _AES_ENC_us30_U463  ( .A1(_AES_ENC_us30_n1025 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n980 ) );
NOR2_X2 _AES_ENC_us30_U462  ( .A1(_AES_ENC_us30_n1073 ), .A2(_AES_ENC_us30_n1094 ), .ZN(_AES_ENC_us30_n795 ) );
NOR2_X2 _AES_ENC_us30_U461  ( .A1(_AES_ENC_us30_n795 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n799 ) );
NOR2_X2 _AES_ENC_us30_U460  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n981 ) );
NOR2_X2 _AES_ENC_us30_U459  ( .A1(_AES_ENC_us30_n1102 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n643 ) );
NOR2_X2 _AES_ENC_us30_U458  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n621 ), .ZN(_AES_ENC_us30_n642 ) );
NOR2_X2 _AES_ENC_us30_U455  ( .A1(_AES_ENC_us30_n911 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n644 ) );
NOR4_X2 _AES_ENC_us30_U448  ( .A1(_AES_ENC_us30_n644 ), .A2(_AES_ENC_us30_n643 ), .A3(_AES_ENC_us30_n804 ), .A4(_AES_ENC_us30_n642 ), .ZN(_AES_ENC_us30_n645 ) );
NOR2_X2 _AES_ENC_us30_U447  ( .A1(_AES_ENC_us30_n1102 ), .A2(_AES_ENC_us30_n910 ), .ZN(_AES_ENC_us30_n932 ) );
NOR2_X2 _AES_ENC_us30_U442  ( .A1(_AES_ENC_us30_n1102 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n755 ) );
NOR2_X2 _AES_ENC_us30_U441  ( .A1(_AES_ENC_us30_n931 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n743 ) );
NOR2_X2 _AES_ENC_us30_U438  ( .A1(_AES_ENC_us30_n1072 ), .A2(_AES_ENC_us30_n1094 ), .ZN(_AES_ENC_us30_n930 ) );
NOR2_X2 _AES_ENC_us30_U435  ( .A1(_AES_ENC_us30_n1074 ), .A2(_AES_ENC_us30_n1025 ), .ZN(_AES_ENC_us30_n891 ) );
NOR2_X2 _AES_ENC_us30_U434  ( .A1(_AES_ENC_us30_n891 ), .A2(_AES_ENC_us30_n609 ), .ZN(_AES_ENC_us30_n894 ) );
NOR3_X2 _AES_ENC_us30_U433  ( .A1(_AES_ENC_us30_n623 ), .A2(_AES_ENC_sa30[1]), .A3(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n683 ));
INV_X4 _AES_ENC_us30_U428  ( .A(_AES_ENC_us30_n931 ), .ZN(_AES_ENC_us30_n623 ) );
NOR2_X2 _AES_ENC_us30_U427  ( .A1(_AES_ENC_us30_n996 ), .A2(_AES_ENC_us30_n931 ), .ZN(_AES_ENC_us30_n704 ) );
NOR2_X2 _AES_ENC_us30_U421  ( .A1(_AES_ENC_us30_n931 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n685 ) );
NOR2_X2 _AES_ENC_us30_U420  ( .A1(_AES_ENC_us30_n1029 ), .A2(_AES_ENC_us30_n1025 ), .ZN(_AES_ENC_us30_n1079 ) );
NOR3_X2 _AES_ENC_us30_U419  ( .A1(_AES_ENC_us30_n589 ), .A2(_AES_ENC_us30_n1025 ), .A3(_AES_ENC_us30_n616 ), .ZN(_AES_ENC_us30_n945 ) );
NOR2_X2 _AES_ENC_us30_U418  ( .A1(_AES_ENC_us30_n626 ), .A2(_AES_ENC_us30_n611 ), .ZN(_AES_ENC_us30_n800 ) );
NOR3_X2 _AES_ENC_us30_U417  ( .A1(_AES_ENC_us30_n590 ), .A2(_AES_ENC_us30_n627 ), .A3(_AES_ENC_us30_n611 ), .ZN(_AES_ENC_us30_n798 ) );
NOR3_X2 _AES_ENC_us30_U416  ( .A1(_AES_ENC_us30_n610 ), .A2(_AES_ENC_us30_n572 ), .A3(_AES_ENC_us30_n575 ), .ZN(_AES_ENC_us30_n962 ) );
NOR3_X2 _AES_ENC_us30_U415  ( .A1(_AES_ENC_us30_n959 ), .A2(_AES_ENC_us30_n572 ), .A3(_AES_ENC_us30_n609 ), .ZN(_AES_ENC_us30_n768 ) );
NOR3_X2 _AES_ENC_us30_U414  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n572 ), .A3(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n694 ) );
NOR3_X2 _AES_ENC_us30_U413  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n572 ), .A3(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n895 ) );
NOR3_X2 _AES_ENC_us30_U410  ( .A1(_AES_ENC_us30_n1008 ), .A2(_AES_ENC_us30_n1007 ), .A3(_AES_ENC_us30_n1006 ), .ZN(_AES_ENC_us30_n1018 ) );
NOR4_X2 _AES_ENC_us30_U409  ( .A1(_AES_ENC_us30_n806 ), .A2(_AES_ENC_us30_n805 ), .A3(_AES_ENC_us30_n804 ), .A4(_AES_ENC_us30_n803 ), .ZN(_AES_ENC_us30_n807 ) );
NOR3_X2 _AES_ENC_us30_U406  ( .A1(_AES_ENC_us30_n799 ), .A2(_AES_ENC_us30_n798 ), .A3(_AES_ENC_us30_n797 ), .ZN(_AES_ENC_us30_n808 ) );
NOR4_X2 _AES_ENC_us30_U405  ( .A1(_AES_ENC_us30_n711 ), .A2(_AES_ENC_us30_n710 ), .A3(_AES_ENC_us30_n709 ), .A4(_AES_ENC_us30_n708 ), .ZN(_AES_ENC_us30_n712 ) );
NOR4_X2 _AES_ENC_us30_U404  ( .A1(_AES_ENC_us30_n963 ), .A2(_AES_ENC_us30_n962 ), .A3(_AES_ENC_us30_n961 ), .A4(_AES_ENC_us30_n960 ), .ZN(_AES_ENC_us30_n964 ) );
NOR3_X2 _AES_ENC_us30_U403  ( .A1(_AES_ENC_us30_n1101 ), .A2(_AES_ENC_us30_n1100 ), .A3(_AES_ENC_us30_n1099 ), .ZN(_AES_ENC_us30_n1109 ) );
NOR2_X2 _AES_ENC_us30_U401  ( .A1(_AES_ENC_us30_n669 ), .A2(_AES_ENC_us30_n668 ), .ZN(_AES_ENC_us30_n673 ) );
NOR4_X2 _AES_ENC_us30_U400  ( .A1(_AES_ENC_us30_n946 ), .A2(_AES_ENC_us30_n1046 ), .A3(_AES_ENC_us30_n671 ), .A4(_AES_ENC_us30_n670 ), .ZN(_AES_ENC_us30_n672 ) );
NOR4_X2 _AES_ENC_us30_U399  ( .A1(_AES_ENC_us30_n843 ), .A2(_AES_ENC_us30_n842 ), .A3(_AES_ENC_us30_n841 ), .A4(_AES_ENC_us30_n840 ), .ZN(_AES_ENC_us30_n844 ) );
NOR3_X2 _AES_ENC_us30_U398  ( .A1(_AES_ENC_us30_n743 ), .A2(_AES_ENC_us30_n742 ), .A3(_AES_ENC_us30_n741 ), .ZN(_AES_ENC_us30_n744 ) );
NOR2_X2 _AES_ENC_us30_U397  ( .A1(_AES_ENC_us30_n697 ), .A2(_AES_ENC_us30_n658 ), .ZN(_AES_ENC_us30_n659 ) );
NOR2_X2 _AES_ENC_us30_U396  ( .A1(_AES_ENC_us30_n1078 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n1033 ) );
NOR2_X2 _AES_ENC_us30_U393  ( .A1(_AES_ENC_us30_n1031 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n1032 ) );
NOR3_X2 _AES_ENC_us30_U390  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n1025 ), .A3(_AES_ENC_us30_n1074 ), .ZN(_AES_ENC_us30_n1035 ) );
NOR4_X2 _AES_ENC_us30_U389  ( .A1(_AES_ENC_us30_n1035 ), .A2(_AES_ENC_us30_n1034 ), .A3(_AES_ENC_us30_n1033 ), .A4(_AES_ENC_us30_n1032 ), .ZN(_AES_ENC_us30_n1036 ) );
NOR2_X2 _AES_ENC_us30_U388  ( .A1(_AES_ENC_us30_n598 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n885 ) );
NOR2_X2 _AES_ENC_us30_U387  ( .A1(_AES_ENC_us30_n623 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n882 ) );
NOR2_X2 _AES_ENC_us30_U386  ( .A1(_AES_ENC_us30_n1053 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n884 ) );
NOR4_X2 _AES_ENC_us30_U385  ( .A1(_AES_ENC_us30_n885 ), .A2(_AES_ENC_us30_n884 ), .A3(_AES_ENC_us30_n883 ), .A4(_AES_ENC_us30_n882 ), .ZN(_AES_ENC_us30_n886 ) );
NOR2_X2 _AES_ENC_us30_U384  ( .A1(_AES_ENC_us30_n825 ), .A2(_AES_ENC_us30_n578 ), .ZN(_AES_ENC_us30_n830 ) );
NOR2_X2 _AES_ENC_us30_U383  ( .A1(_AES_ENC_us30_n827 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n829 ) );
NOR2_X2 _AES_ENC_us30_U382  ( .A1(_AES_ENC_us30_n572 ), .A2(_AES_ENC_us30_n579 ), .ZN(_AES_ENC_us30_n828 ) );
NOR4_X2 _AES_ENC_us30_U374  ( .A1(_AES_ENC_us30_n831 ), .A2(_AES_ENC_us30_n830 ), .A3(_AES_ENC_us30_n829 ), .A4(_AES_ENC_us30_n828 ), .ZN(_AES_ENC_us30_n832 ) );
NOR2_X2 _AES_ENC_us30_U373  ( .A1(_AES_ENC_us30_n606 ), .A2(_AES_ENC_us30_n582 ), .ZN(_AES_ENC_us30_n1104 ) );
NOR2_X2 _AES_ENC_us30_U372  ( .A1(_AES_ENC_us30_n1102 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n1106 ) );
NOR2_X2 _AES_ENC_us30_U370  ( .A1(_AES_ENC_us30_n1103 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n1105 ) );
NOR4_X2 _AES_ENC_us30_U369  ( .A1(_AES_ENC_us30_n1107 ), .A2(_AES_ENC_us30_n1106 ), .A3(_AES_ENC_us30_n1105 ), .A4(_AES_ENC_us30_n1104 ), .ZN(_AES_ENC_us30_n1108 ) );
NOR3_X2 _AES_ENC_us30_U368  ( .A1(_AES_ENC_us30_n959 ), .A2(_AES_ENC_us30_n621 ), .A3(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n963 ) );
NOR2_X2 _AES_ENC_us30_U367  ( .A1(_AES_ENC_us30_n626 ), .A2(_AES_ENC_us30_n627 ), .ZN(_AES_ENC_us30_n1114 ) );
INV_X4 _AES_ENC_us30_U366  ( .A(_AES_ENC_us30_n1024 ), .ZN(_AES_ENC_us30_n606 ) );
NOR3_X2 _AES_ENC_us30_U365  ( .A1(_AES_ENC_us30_n910 ), .A2(_AES_ENC_us30_n1059 ), .A3(_AES_ENC_us30_n611 ), .ZN(_AES_ENC_us30_n1115 ) );
INV_X4 _AES_ENC_us30_U364  ( .A(_AES_ENC_us30_n1094 ), .ZN(_AES_ENC_us30_n613 ) );
NOR2_X2 _AES_ENC_us30_U363  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n931 ), .ZN(_AES_ENC_us30_n1100 ) );
INV_X4 _AES_ENC_us30_U354  ( .A(_AES_ENC_us30_n1093 ), .ZN(_AES_ENC_us30_n617 ) );
NOR2_X2 _AES_ENC_us30_U353  ( .A1(_AES_ENC_us30_n569 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n929 ) );
NOR2_X2 _AES_ENC_us30_U352  ( .A1(_AES_ENC_us30_n620 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n926 ) );
NOR2_X2 _AES_ENC_us30_U351  ( .A1(_AES_ENC_us30_n572 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n1095 ) );
NOR2_X2 _AES_ENC_us30_U350  ( .A1(_AES_ENC_us30_n609 ), .A2(_AES_ENC_us30_n627 ), .ZN(_AES_ENC_us30_n1010 ) );
NOR2_X2 _AES_ENC_us30_U349  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n1103 ) );
NOR2_X2 _AES_ENC_us30_U348  ( .A1(_AES_ENC_us30_n622 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n1059 ) );
NOR2_X2 _AES_ENC_us30_U347  ( .A1(_AES_ENC_sa30[1]), .A2(_AES_ENC_us30_n1120 ), .ZN(_AES_ENC_us30_n1022 ) );
NOR2_X2 _AES_ENC_us30_U346  ( .A1(_AES_ENC_us30_n619 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n911 ) );
NOR2_X2 _AES_ENC_us30_U345  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_us30_n1025 ), .ZN(_AES_ENC_us30_n826 ) );
NOR2_X2 _AES_ENC_us30_U338  ( .A1(_AES_ENC_us30_n626 ), .A2(_AES_ENC_us30_n607 ), .ZN(_AES_ENC_us30_n1072 ) );
NOR2_X2 _AES_ENC_us30_U335  ( .A1(_AES_ENC_us30_n627 ), .A2(_AES_ENC_us30_n616 ), .ZN(_AES_ENC_us30_n956 ) );
NOR2_X2 _AES_ENC_us30_U329  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_us30_n624 ), .ZN(_AES_ENC_us30_n1121 ) );
NOR2_X2 _AES_ENC_us30_U328  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_us30_n624 ), .ZN(_AES_ENC_us30_n1058 ) );
NOR2_X2 _AES_ENC_us30_U327  ( .A1(_AES_ENC_us30_n625 ), .A2(_AES_ENC_us30_n611 ), .ZN(_AES_ENC_us30_n1073 ) );
NOR2_X2 _AES_ENC_us30_U325  ( .A1(_AES_ENC_sa30[1]), .A2(_AES_ENC_us30_n1025 ), .ZN(_AES_ENC_us30_n1054 ) );
NOR2_X2 _AES_ENC_us30_U324  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_us30_n931 ), .ZN(_AES_ENC_us30_n1029 ) );
NOR2_X2 _AES_ENC_us30_U319  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n1056 ) );
NOR2_X2 _AES_ENC_us30_U318  ( .A1(_AES_ENC_us30_n614 ), .A2(_AES_ENC_us30_n626 ), .ZN(_AES_ENC_us30_n1050 ) );
NOR2_X2 _AES_ENC_us30_U317  ( .A1(_AES_ENC_us30_n1121 ), .A2(_AES_ENC_us30_n1025 ), .ZN(_AES_ENC_us30_n1120 ) );
NOR2_X2 _AES_ENC_us30_U316  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_us30_n572 ), .ZN(_AES_ENC_us30_n1074 ) );
NOR2_X2 _AES_ENC_us30_U315  ( .A1(_AES_ENC_us30_n1058 ), .A2(_AES_ENC_us30_n1054 ), .ZN(_AES_ENC_us30_n878 ) );
NOR2_X2 _AES_ENC_us30_U314  ( .A1(_AES_ENC_us30_n878 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n879 ) );
NOR2_X2 _AES_ENC_us30_U312  ( .A1(_AES_ENC_us30_n880 ), .A2(_AES_ENC_us30_n879 ), .ZN(_AES_ENC_us30_n887 ) );
NOR2_X2 _AES_ENC_us30_U311  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n588 ), .ZN(_AES_ENC_us30_n957 ) );
NOR2_X2 _AES_ENC_us30_U310  ( .A1(_AES_ENC_us30_n958 ), .A2(_AES_ENC_us30_n957 ), .ZN(_AES_ENC_us30_n965 ) );
NOR3_X2 _AES_ENC_us30_U309  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n1091 ), .A3(_AES_ENC_us30_n1022 ), .ZN(_AES_ENC_us30_n720 ) );
NOR3_X2 _AES_ENC_us30_U303  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n1054 ), .A3(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n719 ) );
NOR2_X2 _AES_ENC_us30_U302  ( .A1(_AES_ENC_us30_n720 ), .A2(_AES_ENC_us30_n719 ), .ZN(_AES_ENC_us30_n726 ) );
NOR2_X2 _AES_ENC_us30_U300  ( .A1(_AES_ENC_us30_n614 ), .A2(_AES_ENC_us30_n591 ), .ZN(_AES_ENC_us30_n865 ) );
NOR2_X2 _AES_ENC_us30_U299  ( .A1(_AES_ENC_us30_n1059 ), .A2(_AES_ENC_us30_n1058 ), .ZN(_AES_ENC_us30_n1060 ) );
NOR2_X2 _AES_ENC_us30_U298  ( .A1(_AES_ENC_us30_n1095 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n668 ) );
NOR2_X2 _AES_ENC_us30_U297  ( .A1(_AES_ENC_us30_n911 ), .A2(_AES_ENC_us30_n910 ), .ZN(_AES_ENC_us30_n912 ) );
NOR2_X2 _AES_ENC_us30_U296  ( .A1(_AES_ENC_us30_n912 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n916 ) );
NOR2_X2 _AES_ENC_us30_U295  ( .A1(_AES_ENC_us30_n826 ), .A2(_AES_ENC_us30_n573 ), .ZN(_AES_ENC_us30_n750 ) );
NOR2_X2 _AES_ENC_us30_U294  ( .A1(_AES_ENC_us30_n750 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n751 ) );
NOR2_X2 _AES_ENC_us30_U293  ( .A1(_AES_ENC_us30_n907 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n908 ) );
NOR2_X2 _AES_ENC_us30_U292  ( .A1(_AES_ENC_us30_n990 ), .A2(_AES_ENC_us30_n926 ), .ZN(_AES_ENC_us30_n780 ) );
NOR2_X2 _AES_ENC_us30_U291  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n584 ), .ZN(_AES_ENC_us30_n838 ) );
NOR2_X2 _AES_ENC_us30_U290  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n602 ), .ZN(_AES_ENC_us30_n837 ) );
NOR2_X2 _AES_ENC_us30_U284  ( .A1(_AES_ENC_us30_n838 ), .A2(_AES_ENC_us30_n837 ), .ZN(_AES_ENC_us30_n845 ) );
NOR2_X2 _AES_ENC_us30_U283  ( .A1(_AES_ENC_us30_n1022 ), .A2(_AES_ENC_us30_n1058 ), .ZN(_AES_ENC_us30_n740 ) );
NOR2_X2 _AES_ENC_us30_U282  ( .A1(_AES_ENC_us30_n740 ), .A2(_AES_ENC_us30_n616 ), .ZN(_AES_ENC_us30_n742 ) );
NOR2_X2 _AES_ENC_us30_U281  ( .A1(_AES_ENC_us30_n1098 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n1099 ) );
NOR2_X2 _AES_ENC_us30_U280  ( .A1(_AES_ENC_us30_n1120 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n993 ) );
NOR2_X2 _AES_ENC_us30_U279  ( .A1(_AES_ENC_us30_n993 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n994 ) );
NOR2_X2 _AES_ENC_us30_U273  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n620 ), .ZN(_AES_ENC_us30_n1026 ) );
NOR2_X2 _AES_ENC_us30_U272  ( .A1(_AES_ENC_us30_n573 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n1027 ) );
NOR2_X2 _AES_ENC_us30_U271  ( .A1(_AES_ENC_us30_n1027 ), .A2(_AES_ENC_us30_n1026 ), .ZN(_AES_ENC_us30_n1028 ) );
NOR2_X2 _AES_ENC_us30_U270  ( .A1(_AES_ENC_us30_n1029 ), .A2(_AES_ENC_us30_n1028 ), .ZN(_AES_ENC_us30_n1034 ) );
NOR4_X2 _AES_ENC_us30_U269  ( .A1(_AES_ENC_us30_n757 ), .A2(_AES_ENC_us30_n756 ), .A3(_AES_ENC_us30_n755 ), .A4(_AES_ENC_us30_n754 ), .ZN(_AES_ENC_us30_n758 ) );
NOR2_X2 _AES_ENC_us30_U268  ( .A1(_AES_ENC_us30_n752 ), .A2(_AES_ENC_us30_n751 ), .ZN(_AES_ENC_us30_n759 ) );
NOR2_X2 _AES_ENC_us30_U267  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n1071 ), .ZN(_AES_ENC_us30_n669 ) );
NOR2_X2 _AES_ENC_us30_U263  ( .A1(_AES_ENC_us30_n1056 ), .A2(_AES_ENC_us30_n990 ), .ZN(_AES_ENC_us30_n991 ) );
NOR2_X2 _AES_ENC_us30_U262  ( .A1(_AES_ENC_us30_n991 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n995 ) );
NOR2_X2 _AES_ENC_us30_U258  ( .A1(_AES_ENC_us30_n607 ), .A2(_AES_ENC_us30_n590 ), .ZN(_AES_ENC_us30_n1008 ) );
NOR2_X2 _AES_ENC_us30_U255  ( .A1(_AES_ENC_us30_n839 ), .A2(_AES_ENC_us30_n582 ), .ZN(_AES_ENC_us30_n693 ) );
NOR2_X2 _AES_ENC_us30_U254  ( .A1(_AES_ENC_us30_n606 ), .A2(_AES_ENC_us30_n906 ), .ZN(_AES_ENC_us30_n741 ) );
NOR2_X2 _AES_ENC_us30_U253  ( .A1(_AES_ENC_us30_n1054 ), .A2(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n763 ) );
NOR2_X2 _AES_ENC_us30_U252  ( .A1(_AES_ENC_us30_n763 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n769 ) );
NOR2_X2 _AES_ENC_us30_U251  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n577 ), .ZN(_AES_ENC_us30_n1007 ) );
NOR2_X2 _AES_ENC_us30_U250  ( .A1(_AES_ENC_us30_n609 ), .A2(_AES_ENC_us30_n580 ), .ZN(_AES_ENC_us30_n1123 ) );
NOR2_X2 _AES_ENC_us30_U243  ( .A1(_AES_ENC_us30_n609 ), .A2(_AES_ENC_us30_n590 ), .ZN(_AES_ENC_us30_n710 ) );
INV_X4 _AES_ENC_us30_U242  ( .A(_AES_ENC_us30_n1029 ), .ZN(_AES_ENC_us30_n582 ) );
NOR2_X2 _AES_ENC_us30_U241  ( .A1(_AES_ENC_us30_n616 ), .A2(_AES_ENC_us30_n597 ), .ZN(_AES_ENC_us30_n883 ) );
NOR2_X2 _AES_ENC_us30_U240  ( .A1(_AES_ENC_us30_n593 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n1125 ) );
NOR2_X2 _AES_ENC_us30_U239  ( .A1(_AES_ENC_us30_n990 ), .A2(_AES_ENC_us30_n929 ), .ZN(_AES_ENC_us30_n892 ) );
NOR2_X2 _AES_ENC_us30_U238  ( .A1(_AES_ENC_us30_n892 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n893 ) );
NOR2_X2 _AES_ENC_us30_U237  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n602 ), .ZN(_AES_ENC_us30_n950 ) );
NOR2_X2 _AES_ENC_us30_U236  ( .A1(_AES_ENC_us30_n1079 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n1082 ) );
NOR2_X2 _AES_ENC_us30_U235  ( .A1(_AES_ENC_us30_n910 ), .A2(_AES_ENC_us30_n1056 ), .ZN(_AES_ENC_us30_n941 ) );
NOR2_X2 _AES_ENC_us30_U234  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n1077 ), .ZN(_AES_ENC_us30_n841 ) );
NOR2_X2 _AES_ENC_us30_U229  ( .A1(_AES_ENC_us30_n623 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n630 ) );
NOR2_X2 _AES_ENC_us30_U228  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n602 ), .ZN(_AES_ENC_us30_n806 ) );
NOR2_X2 _AES_ENC_us30_U227  ( .A1(_AES_ENC_us30_n623 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n948 ) );
NOR2_X2 _AES_ENC_us30_U226  ( .A1(_AES_ENC_us30_n606 ), .A2(_AES_ENC_us30_n589 ), .ZN(_AES_ENC_us30_n997 ) );
NOR2_X2 _AES_ENC_us30_U225  ( .A1(_AES_ENC_us30_n1121 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n1122 ) );
NOR2_X2 _AES_ENC_us30_U223  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n1023 ), .ZN(_AES_ENC_us30_n756 ) );
NOR2_X2 _AES_ENC_us30_U222  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n602 ), .ZN(_AES_ENC_us30_n870 ) );
NOR2_X2 _AES_ENC_us30_U221  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n569 ), .ZN(_AES_ENC_us30_n947 ) );
NOR2_X2 _AES_ENC_us30_U217  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n1077 ), .ZN(_AES_ENC_us30_n1084 ) );
NOR2_X2 _AES_ENC_us30_U213  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n855 ), .ZN(_AES_ENC_us30_n709 ) );
NOR2_X2 _AES_ENC_us30_U212  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n589 ), .ZN(_AES_ENC_us30_n868 ) );
NOR2_X2 _AES_ENC_us30_U211  ( .A1(_AES_ENC_us30_n1120 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n1124 ) );
NOR2_X2 _AES_ENC_us30_U210  ( .A1(_AES_ENC_us30_n1120 ), .A2(_AES_ENC_us30_n839 ), .ZN(_AES_ENC_us30_n842 ) );
NOR2_X2 _AES_ENC_us30_U209  ( .A1(_AES_ENC_us30_n1120 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n696 ) );
NOR2_X2 _AES_ENC_us30_U208  ( .A1(_AES_ENC_us30_n1074 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n1076 ) );
NOR2_X2 _AES_ENC_us30_U207  ( .A1(_AES_ENC_us30_n1074 ), .A2(_AES_ENC_us30_n620 ), .ZN(_AES_ENC_us30_n781 ) );
NOR3_X2 _AES_ENC_us30_U201  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n1056 ), .A3(_AES_ENC_us30_n990 ), .ZN(_AES_ENC_us30_n979 ) );
NOR3_X2 _AES_ENC_us30_U200  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n1058 ), .A3(_AES_ENC_us30_n1059 ), .ZN(_AES_ENC_us30_n854 ) );
NOR2_X2 _AES_ENC_us30_U199  ( .A1(_AES_ENC_us30_n996 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n869 ) );
NOR2_X2 _AES_ENC_us30_U198  ( .A1(_AES_ENC_us30_n1056 ), .A2(_AES_ENC_us30_n1074 ), .ZN(_AES_ENC_us30_n1057 ) );
NOR3_X2 _AES_ENC_us30_U197  ( .A1(_AES_ENC_us30_n607 ), .A2(_AES_ENC_us30_n1120 ), .A3(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n978 ) );
NOR2_X2 _AES_ENC_us30_U196  ( .A1(_AES_ENC_us30_n996 ), .A2(_AES_ENC_us30_n911 ), .ZN(_AES_ENC_us30_n1116 ) );
NOR2_X2 _AES_ENC_us30_U195  ( .A1(_AES_ENC_us30_n1074 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n754 ) );
NOR2_X2 _AES_ENC_us30_U194  ( .A1(_AES_ENC_us30_n926 ), .A2(_AES_ENC_us30_n1103 ), .ZN(_AES_ENC_us30_n977 ) );
NOR2_X2 _AES_ENC_us30_U187  ( .A1(_AES_ENC_us30_n839 ), .A2(_AES_ENC_us30_n824 ), .ZN(_AES_ENC_us30_n1092 ) );
NOR2_X2 _AES_ENC_us30_U186  ( .A1(_AES_ENC_us30_n573 ), .A2(_AES_ENC_us30_n1074 ), .ZN(_AES_ENC_us30_n684 ) );
NOR2_X2 _AES_ENC_us30_U185  ( .A1(_AES_ENC_us30_n826 ), .A2(_AES_ENC_us30_n1059 ), .ZN(_AES_ENC_us30_n907 ) );
NOR3_X2 _AES_ENC_us30_U184  ( .A1(_AES_ENC_us30_n625 ), .A2(_AES_ENC_us30_n1115 ), .A3(_AES_ENC_us30_n585 ), .ZN(_AES_ENC_us30_n831 ) );
NOR3_X2 _AES_ENC_us30_U183  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n1056 ), .A3(_AES_ENC_us30_n990 ), .ZN(_AES_ENC_us30_n896 ) );
NOR3_X2 _AES_ENC_us30_U182  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n573 ), .A3(_AES_ENC_us30_n1013 ), .ZN(_AES_ENC_us30_n670 ) );
NOR3_X2 _AES_ENC_us30_U181  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n1091 ), .A3(_AES_ENC_us30_n1022 ), .ZN(_AES_ENC_us30_n843 ) );
NOR2_X2 _AES_ENC_us30_U180  ( .A1(_AES_ENC_us30_n1029 ), .A2(_AES_ENC_us30_n1095 ), .ZN(_AES_ENC_us30_n735 ) );
NOR2_X2 _AES_ENC_us30_U174  ( .A1(_AES_ENC_us30_n1100 ), .A2(_AES_ENC_us30_n854 ), .ZN(_AES_ENC_us30_n860 ) );
NAND3_X2 _AES_ENC_us30_U173  ( .A1(_AES_ENC_us30_n569 ), .A2(_AES_ENC_us30_n582 ), .A3(_AES_ENC_us30_n681 ), .ZN(_AES_ENC_us30_n691 ) );
NOR2_X2 _AES_ENC_us30_U172  ( .A1(_AES_ENC_us30_n683 ), .A2(_AES_ENC_us30_n682 ), .ZN(_AES_ENC_us30_n690 ) );
NOR3_X2 _AES_ENC_us30_U171  ( .A1(_AES_ENC_us30_n695 ), .A2(_AES_ENC_us30_n694 ), .A3(_AES_ENC_us30_n693 ), .ZN(_AES_ENC_us30_n700 ) );
NOR4_X2 _AES_ENC_us30_U170  ( .A1(_AES_ENC_us30_n983 ), .A2(_AES_ENC_us30_n698 ), .A3(_AES_ENC_us30_n697 ), .A4(_AES_ENC_us30_n696 ), .ZN(_AES_ENC_us30_n699 ) );
NOR2_X2 _AES_ENC_us30_U169  ( .A1(_AES_ENC_us30_n946 ), .A2(_AES_ENC_us30_n945 ), .ZN(_AES_ENC_us30_n952 ) );
NOR4_X2 _AES_ENC_us30_U168  ( .A1(_AES_ENC_us30_n950 ), .A2(_AES_ENC_us30_n949 ), .A3(_AES_ENC_us30_n948 ), .A4(_AES_ENC_us30_n947 ), .ZN(_AES_ENC_us30_n951 ) );
NOR4_X2 _AES_ENC_us30_U162  ( .A1(_AES_ENC_us30_n896 ), .A2(_AES_ENC_us30_n895 ), .A3(_AES_ENC_us30_n894 ), .A4(_AES_ENC_us30_n893 ), .ZN(_AES_ENC_us30_n897 ) );
NOR2_X2 _AES_ENC_us30_U161  ( .A1(_AES_ENC_us30_n866 ), .A2(_AES_ENC_us30_n865 ), .ZN(_AES_ENC_us30_n872 ) );
NOR4_X2 _AES_ENC_us30_U160  ( .A1(_AES_ENC_us30_n870 ), .A2(_AES_ENC_us30_n869 ), .A3(_AES_ENC_us30_n868 ), .A4(_AES_ENC_us30_n867 ), .ZN(_AES_ENC_us30_n871 ) );
NOR4_X2 _AES_ENC_us30_U159  ( .A1(_AES_ENC_us30_n983 ), .A2(_AES_ENC_us30_n982 ), .A3(_AES_ENC_us30_n981 ), .A4(_AES_ENC_us30_n980 ), .ZN(_AES_ENC_us30_n984 ) );
NOR2_X2 _AES_ENC_us30_U158  ( .A1(_AES_ENC_us30_n979 ), .A2(_AES_ENC_us30_n978 ), .ZN(_AES_ENC_us30_n985 ) );
NOR4_X2 _AES_ENC_us30_U157  ( .A1(_AES_ENC_us30_n1125 ), .A2(_AES_ENC_us30_n1124 ), .A3(_AES_ENC_us30_n1123 ), .A4(_AES_ENC_us30_n1122 ), .ZN(_AES_ENC_us30_n1126 ) );
NOR4_X2 _AES_ENC_us30_U156  ( .A1(_AES_ENC_us30_n1084 ), .A2(_AES_ENC_us30_n1083 ), .A3(_AES_ENC_us30_n1082 ), .A4(_AES_ENC_us30_n1081 ), .ZN(_AES_ENC_us30_n1085 ) );
NOR2_X2 _AES_ENC_us30_U155  ( .A1(_AES_ENC_us30_n1076 ), .A2(_AES_ENC_us30_n1075 ), .ZN(_AES_ENC_us30_n1086 ) );
NOR3_X2 _AES_ENC_us30_U154  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n1054 ), .A3(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n961 ) );
NOR3_X2 _AES_ENC_us30_U153  ( .A1(_AES_ENC_us30_n620 ), .A2(_AES_ENC_us30_n1074 ), .A3(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n671 ) );
NOR2_X2 _AES_ENC_us30_U152  ( .A1(_AES_ENC_us30_n1057 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n1062 ) );
NOR2_X2 _AES_ENC_us30_U143  ( .A1(_AES_ENC_us30_n1055 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n1063 ) );
NOR2_X2 _AES_ENC_us30_U142  ( .A1(_AES_ENC_us30_n1060 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n1061 ) );
NOR4_X2 _AES_ENC_us30_U141  ( .A1(_AES_ENC_us30_n1064 ), .A2(_AES_ENC_us30_n1063 ), .A3(_AES_ENC_us30_n1062 ), .A4(_AES_ENC_us30_n1061 ), .ZN(_AES_ENC_us30_n1065 ) );
NOR3_X2 _AES_ENC_us30_U140  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n1120 ), .A3(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n918 ) );
NOR3_X2 _AES_ENC_us30_U132  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n573 ), .A3(_AES_ENC_us30_n1013 ), .ZN(_AES_ENC_us30_n917 ) );
NOR2_X2 _AES_ENC_us30_U131  ( .A1(_AES_ENC_us30_n914 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n915 ) );
NOR4_X2 _AES_ENC_us30_U130  ( .A1(_AES_ENC_us30_n918 ), .A2(_AES_ENC_us30_n917 ), .A3(_AES_ENC_us30_n916 ), .A4(_AES_ENC_us30_n915 ), .ZN(_AES_ENC_us30_n919 ) );
NOR2_X2 _AES_ENC_us30_U129  ( .A1(_AES_ENC_us30_n616 ), .A2(_AES_ENC_us30_n580 ), .ZN(_AES_ENC_us30_n771 ) );
NOR2_X2 _AES_ENC_us30_U128  ( .A1(_AES_ENC_us30_n1103 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n772 ) );
NOR2_X2 _AES_ENC_us30_U127  ( .A1(_AES_ENC_us30_n610 ), .A2(_AES_ENC_us30_n599 ), .ZN(_AES_ENC_us30_n773 ) );
NOR4_X2 _AES_ENC_us30_U126  ( .A1(_AES_ENC_us30_n773 ), .A2(_AES_ENC_us30_n772 ), .A3(_AES_ENC_us30_n771 ), .A4(_AES_ENC_us30_n770 ), .ZN(_AES_ENC_us30_n774 ) );
NOR2_X2 _AES_ENC_us30_U121  ( .A1(_AES_ENC_us30_n735 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n687 ) );
NOR2_X2 _AES_ENC_us30_U120  ( .A1(_AES_ENC_us30_n684 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n688 ) );
NOR2_X2 _AES_ENC_us30_U119  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n600 ), .ZN(_AES_ENC_us30_n686 ) );
NOR4_X2 _AES_ENC_us30_U118  ( .A1(_AES_ENC_us30_n688 ), .A2(_AES_ENC_us30_n687 ), .A3(_AES_ENC_us30_n686 ), .A4(_AES_ENC_us30_n685 ), .ZN(_AES_ENC_us30_n689 ) );
NOR2_X2 _AES_ENC_us30_U117  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n595 ), .ZN(_AES_ENC_us30_n858 ) );
NOR2_X2 _AES_ENC_us30_U116  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n855 ), .ZN(_AES_ENC_us30_n857 ) );
NOR2_X2 _AES_ENC_us30_U115  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n587 ), .ZN(_AES_ENC_us30_n856 ) );
NOR4_X2 _AES_ENC_us30_U106  ( .A1(_AES_ENC_us30_n858 ), .A2(_AES_ENC_us30_n857 ), .A3(_AES_ENC_us30_n856 ), .A4(_AES_ENC_us30_n958 ), .ZN(_AES_ENC_us30_n859 ) );
NOR2_X2 _AES_ENC_us30_U105  ( .A1(_AES_ENC_us30_n780 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n784 ) );
NOR2_X2 _AES_ENC_us30_U104  ( .A1(_AES_ENC_us30_n1117 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n782 ) );
NOR2_X2 _AES_ENC_us30_U103  ( .A1(_AES_ENC_us30_n781 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n783 ) );
NOR4_X2 _AES_ENC_us30_U102  ( .A1(_AES_ENC_us30_n880 ), .A2(_AES_ENC_us30_n784 ), .A3(_AES_ENC_us30_n783 ), .A4(_AES_ENC_us30_n782 ), .ZN(_AES_ENC_us30_n785 ) );
NOR2_X2 _AES_ENC_us30_U101  ( .A1(_AES_ENC_us30_n583 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n814 ) );
NOR2_X2 _AES_ENC_us30_U100  ( .A1(_AES_ENC_us30_n907 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n813 ) );
NOR3_X2 _AES_ENC_us30_U95  ( .A1(_AES_ENC_us30_n606 ), .A2(_AES_ENC_us30_n1058 ), .A3(_AES_ENC_us30_n1059 ), .ZN(_AES_ENC_us30_n815 ) );
NOR4_X2 _AES_ENC_us30_U94  ( .A1(_AES_ENC_us30_n815 ), .A2(_AES_ENC_us30_n814 ), .A3(_AES_ENC_us30_n813 ), .A4(_AES_ENC_us30_n812 ), .ZN(_AES_ENC_us30_n816 ) );
NOR2_X2 _AES_ENC_us30_U93  ( .A1(_AES_ENC_us30_n617 ), .A2(_AES_ENC_us30_n569 ), .ZN(_AES_ENC_us30_n721 ) );
NOR2_X2 _AES_ENC_us30_U92  ( .A1(_AES_ENC_us30_n1031 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n723 ) );
NOR2_X2 _AES_ENC_us30_U91  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n1096 ), .ZN(_AES_ENC_us30_n722 ) );
NOR4_X2 _AES_ENC_us30_U90  ( .A1(_AES_ENC_us30_n724 ), .A2(_AES_ENC_us30_n723 ), .A3(_AES_ENC_us30_n722 ), .A4(_AES_ENC_us30_n721 ), .ZN(_AES_ENC_us30_n725 ) );
NOR2_X2 _AES_ENC_us30_U89  ( .A1(_AES_ENC_us30_n911 ), .A2(_AES_ENC_us30_n990 ), .ZN(_AES_ENC_us30_n1009 ) );
NOR2_X2 _AES_ENC_us30_U88  ( .A1(_AES_ENC_us30_n1013 ), .A2(_AES_ENC_us30_n573 ), .ZN(_AES_ENC_us30_n1014 ) );
NOR2_X2 _AES_ENC_us30_U87  ( .A1(_AES_ENC_us30_n1014 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n1015 ) );
NOR4_X2 _AES_ENC_us30_U86  ( .A1(_AES_ENC_us30_n1016 ), .A2(_AES_ENC_us30_n1015 ), .A3(_AES_ENC_us30_n1119 ), .A4(_AES_ENC_us30_n1046 ), .ZN(_AES_ENC_us30_n1017 ) );
NOR2_X2 _AES_ENC_us30_U81  ( .A1(_AES_ENC_us30_n996 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n998 ) );
NOR2_X2 _AES_ENC_us30_U80  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n577 ), .ZN(_AES_ENC_us30_n1000 ) );
NOR2_X2 _AES_ENC_us30_U79  ( .A1(_AES_ENC_us30_n616 ), .A2(_AES_ENC_us30_n1096 ), .ZN(_AES_ENC_us30_n999 ) );
NOR4_X2 _AES_ENC_us30_U78  ( .A1(_AES_ENC_us30_n1000 ), .A2(_AES_ENC_us30_n999 ), .A3(_AES_ENC_us30_n998 ), .A4(_AES_ENC_us30_n997 ), .ZN(_AES_ENC_us30_n1001 ) );
NOR2_X2 _AES_ENC_us30_U74  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n1096 ), .ZN(_AES_ENC_us30_n697 ) );
NOR2_X2 _AES_ENC_us30_U73  ( .A1(_AES_ENC_us30_n620 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n958 ) );
NOR2_X2 _AES_ENC_us30_U72  ( .A1(_AES_ENC_us30_n911 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n983 ) );
NOR2_X2 _AES_ENC_us30_U71  ( .A1(_AES_ENC_us30_n1054 ), .A2(_AES_ENC_us30_n1103 ), .ZN(_AES_ENC_us30_n1031 ) );
INV_X4 _AES_ENC_us30_U65  ( .A(_AES_ENC_us30_n1050 ), .ZN(_AES_ENC_us30_n612 ) );
INV_X4 _AES_ENC_us30_U64  ( .A(_AES_ENC_us30_n1072 ), .ZN(_AES_ENC_us30_n605 ) );
INV_X4 _AES_ENC_us30_U63  ( .A(_AES_ENC_us30_n1073 ), .ZN(_AES_ENC_us30_n604 ) );
NOR2_X2 _AES_ENC_us30_U62  ( .A1(_AES_ENC_us30_n582 ), .A2(_AES_ENC_us30_n613 ), .ZN(_AES_ENC_us30_n880 ) );
NOR3_X2 _AES_ENC_us30_U61  ( .A1(_AES_ENC_us30_n826 ), .A2(_AES_ENC_us30_n1121 ), .A3(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n946 ) );
INV_X4 _AES_ENC_us30_U59  ( .A(_AES_ENC_us30_n1010 ), .ZN(_AES_ENC_us30_n608 ) );
NOR3_X2 _AES_ENC_us30_U58  ( .A1(_AES_ENC_us30_n573 ), .A2(_AES_ENC_us30_n1029 ), .A3(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n1119 ) );
INV_X4 _AES_ENC_us30_U57  ( .A(_AES_ENC_us30_n956 ), .ZN(_AES_ENC_us30_n615 ) );
NOR2_X2 _AES_ENC_us30_U50  ( .A1(_AES_ENC_us30_n623 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n1013 ) );
NOR2_X2 _AES_ENC_us30_U49  ( .A1(_AES_ENC_us30_n620 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n910 ) );
NOR2_X2 _AES_ENC_us30_U48  ( .A1(_AES_ENC_us30_n569 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n1091 ) );
NOR2_X2 _AES_ENC_us30_U47  ( .A1(_AES_ENC_us30_n622 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n990 ) );
NOR2_X2 _AES_ENC_us30_U46  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_us30_n1121 ), .ZN(_AES_ENC_us30_n996 ) );
NOR2_X2 _AES_ENC_us30_U45  ( .A1(_AES_ENC_us30_n610 ), .A2(_AES_ENC_us30_n600 ), .ZN(_AES_ENC_us30_n628 ) );
NOR2_X2 _AES_ENC_us30_U44  ( .A1(_AES_ENC_us30_n576 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n866 ) );
NOR2_X2 _AES_ENC_us30_U43  ( .A1(_AES_ENC_us30_n603 ), .A2(_AES_ENC_us30_n610 ), .ZN(_AES_ENC_us30_n1006 ) );
NOR2_X2 _AES_ENC_us30_U42  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n1117 ), .ZN(_AES_ENC_us30_n1118 ) );
NOR2_X2 _AES_ENC_us30_U41  ( .A1(_AES_ENC_us30_n1119 ), .A2(_AES_ENC_us30_n1118 ), .ZN(_AES_ENC_us30_n1127 ) );
NOR2_X2 _AES_ENC_us30_U36  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n906 ), .ZN(_AES_ENC_us30_n909 ) );
NOR2_X2 _AES_ENC_us30_U35  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n594 ), .ZN(_AES_ENC_us30_n629 ) );
NOR2_X2 _AES_ENC_us30_U34  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n597 ), .ZN(_AES_ENC_us30_n658 ) );
NOR2_X2 _AES_ENC_us30_U33  ( .A1(_AES_ENC_us30_n1116 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n695 ) );
NOR2_X2 _AES_ENC_us30_U32  ( .A1(_AES_ENC_us30_n1078 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n1083 ) );
NOR2_X2 _AES_ENC_us30_U31  ( .A1(_AES_ENC_us30_n941 ), .A2(_AES_ENC_us30_n608 ), .ZN(_AES_ENC_us30_n724 ) );
NOR2_X2 _AES_ENC_us30_U30  ( .A1(_AES_ENC_us30_n598 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n1107 ) );
NOR2_X2 _AES_ENC_us30_U29  ( .A1(_AES_ENC_us30_n576 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n840 ) );
NOR2_X2 _AES_ENC_us30_U24  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n593 ), .ZN(_AES_ENC_us30_n633 ) );
NOR2_X2 _AES_ENC_us30_U23  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n1080 ), .ZN(_AES_ENC_us30_n1081 ) );
NOR2_X2 _AES_ENC_us30_U21  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n1045 ), .ZN(_AES_ENC_us30_n812 ) );
NOR2_X2 _AES_ENC_us30_U20  ( .A1(_AES_ENC_us30_n1009 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n960 ) );
NOR2_X2 _AES_ENC_us30_U19  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n601 ), .ZN(_AES_ENC_us30_n982 ) );
NOR2_X2 _AES_ENC_us30_U18  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n594 ), .ZN(_AES_ENC_us30_n757 ) );
NOR2_X2 _AES_ENC_us30_U17  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n590 ), .ZN(_AES_ENC_us30_n698 ) );
NOR2_X2 _AES_ENC_us30_U16  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n619 ), .ZN(_AES_ENC_us30_n708 ) );
NOR2_X2 _AES_ENC_us30_U15  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n582 ), .ZN(_AES_ENC_us30_n770 ) );
NOR2_X2 _AES_ENC_us30_U10  ( .A1(_AES_ENC_us30_n619 ), .A2(_AES_ENC_us30_n604 ), .ZN(_AES_ENC_us30_n803 ) );
NOR2_X2 _AES_ENC_us30_U9  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n881 ), .ZN(_AES_ENC_us30_n711 ) );
NOR2_X2 _AES_ENC_us30_U8  ( .A1(_AES_ENC_us30_n615 ), .A2(_AES_ENC_us30_n582 ), .ZN(_AES_ENC_us30_n867 ) );
NOR2_X2 _AES_ENC_us30_U7  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n599 ), .ZN(_AES_ENC_us30_n804 ) );
NOR2_X2 _AES_ENC_us30_U6  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n620 ), .ZN(_AES_ENC_us30_n1046 ) );
OR2_X4 _AES_ENC_us30_U5  ( .A1(_AES_ENC_us30_n624 ), .A2(_AES_ENC_sa30[1]),.ZN(_AES_ENC_us30_n570 ) );
OR2_X4 _AES_ENC_us30_U4  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_sa30[4]),.ZN(_AES_ENC_us30_n569 ) );
NAND2_X2 _AES_ENC_us30_U514  ( .A1(_AES_ENC_us30_n1121 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n1030 ) );
AND2_X2 _AES_ENC_us30_U513  ( .A1(_AES_ENC_us30_n597 ), .A2(_AES_ENC_us30_n1030 ), .ZN(_AES_ENC_us30_n1049 ) );
NAND2_X2 _AES_ENC_us30_U511  ( .A1(_AES_ENC_us30_n1049 ), .A2(_AES_ENC_us30_n794 ), .ZN(_AES_ENC_us30_n637 ) );
AND2_X2 _AES_ENC_us30_U493  ( .A1(_AES_ENC_us30_n779 ), .A2(_AES_ENC_us30_n996 ), .ZN(_AES_ENC_us30_n632 ) );
NAND4_X2 _AES_ENC_us30_U485  ( .A1(_AES_ENC_us30_n637 ), .A2(_AES_ENC_us30_n636 ), .A3(_AES_ENC_us30_n635 ), .A4(_AES_ENC_us30_n634 ), .ZN(_AES_ENC_us30_n638 ) );
NAND2_X2 _AES_ENC_us30_U484  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n638 ), .ZN(_AES_ENC_us30_n679 ) );
NAND2_X2 _AES_ENC_us30_U481  ( .A1(_AES_ENC_us30_n1094 ), .A2(_AES_ENC_us30_n591 ), .ZN(_AES_ENC_us30_n648 ) );
NAND2_X2 _AES_ENC_us30_U476  ( .A1(_AES_ENC_us30_n601 ), .A2(_AES_ENC_us30_n590 ), .ZN(_AES_ENC_us30_n762 ) );
NAND2_X2 _AES_ENC_us30_U475  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n762 ), .ZN(_AES_ENC_us30_n647 ) );
NAND4_X2 _AES_ENC_us30_U457  ( .A1(_AES_ENC_us30_n648 ), .A2(_AES_ENC_us30_n647 ), .A3(_AES_ENC_us30_n646 ), .A4(_AES_ENC_us30_n645 ), .ZN(_AES_ENC_us30_n649 ) );
NAND2_X2 _AES_ENC_us30_U456  ( .A1(_AES_ENC_sa30[0]), .A2(_AES_ENC_us30_n649 ), .ZN(_AES_ENC_us30_n665 ) );
NAND2_X2 _AES_ENC_us30_U454  ( .A1(_AES_ENC_us30_n596 ), .A2(_AES_ENC_us30_n623 ), .ZN(_AES_ENC_us30_n855 ) );
NAND2_X2 _AES_ENC_us30_U453  ( .A1(_AES_ENC_us30_n587 ), .A2(_AES_ENC_us30_n855 ), .ZN(_AES_ENC_us30_n821 ) );
NAND2_X2 _AES_ENC_us30_U452  ( .A1(_AES_ENC_us30_n1093 ), .A2(_AES_ENC_us30_n821 ), .ZN(_AES_ENC_us30_n662 ) );
NAND2_X2 _AES_ENC_us30_U451  ( .A1(_AES_ENC_us30_n619 ), .A2(_AES_ENC_us30_n589 ), .ZN(_AES_ENC_us30_n650 ) );
NAND2_X2 _AES_ENC_us30_U450  ( .A1(_AES_ENC_us30_n956 ), .A2(_AES_ENC_us30_n650 ), .ZN(_AES_ENC_us30_n661 ) );
NAND2_X2 _AES_ENC_us30_U449  ( .A1(_AES_ENC_us30_n626 ), .A2(_AES_ENC_us30_n627 ), .ZN(_AES_ENC_us30_n839 ) );
OR2_X2 _AES_ENC_us30_U446  ( .A1(_AES_ENC_us30_n839 ), .A2(_AES_ENC_us30_n932 ), .ZN(_AES_ENC_us30_n656 ) );
NAND2_X2 _AES_ENC_us30_U445  ( .A1(_AES_ENC_us30_n621 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n1096 ) );
NAND2_X2 _AES_ENC_us30_U444  ( .A1(_AES_ENC_us30_n1030 ), .A2(_AES_ENC_us30_n1096 ), .ZN(_AES_ENC_us30_n651 ) );
NAND2_X2 _AES_ENC_us30_U443  ( .A1(_AES_ENC_us30_n1114 ), .A2(_AES_ENC_us30_n651 ), .ZN(_AES_ENC_us30_n655 ) );
OR3_X2 _AES_ENC_us30_U440  ( .A1(_AES_ENC_us30_n1079 ), .A2(_AES_ENC_sa30[7]), .A3(_AES_ENC_us30_n626 ), .ZN(_AES_ENC_us30_n654 ));
NAND2_X2 _AES_ENC_us30_U439  ( .A1(_AES_ENC_us30_n593 ), .A2(_AES_ENC_us30_n601 ), .ZN(_AES_ENC_us30_n652 ) );
NAND4_X2 _AES_ENC_us30_U437  ( .A1(_AES_ENC_us30_n656 ), .A2(_AES_ENC_us30_n655 ), .A3(_AES_ENC_us30_n654 ), .A4(_AES_ENC_us30_n653 ), .ZN(_AES_ENC_us30_n657 ) );
NAND2_X2 _AES_ENC_us30_U436  ( .A1(_AES_ENC_sa30[2]), .A2(_AES_ENC_us30_n657 ), .ZN(_AES_ENC_us30_n660 ) );
NAND4_X2 _AES_ENC_us30_U432  ( .A1(_AES_ENC_us30_n662 ), .A2(_AES_ENC_us30_n661 ), .A3(_AES_ENC_us30_n660 ), .A4(_AES_ENC_us30_n659 ), .ZN(_AES_ENC_us30_n663 ) );
NAND2_X2 _AES_ENC_us30_U431  ( .A1(_AES_ENC_us30_n663 ), .A2(_AES_ENC_us30_n574 ), .ZN(_AES_ENC_us30_n664 ) );
NAND2_X2 _AES_ENC_us30_U430  ( .A1(_AES_ENC_us30_n665 ), .A2(_AES_ENC_us30_n664 ), .ZN(_AES_ENC_us30_n666 ) );
NAND2_X2 _AES_ENC_us30_U429  ( .A1(_AES_ENC_sa30[6]), .A2(_AES_ENC_us30_n666 ), .ZN(_AES_ENC_us30_n678 ) );
NAND2_X2 _AES_ENC_us30_U426  ( .A1(_AES_ENC_us30_n735 ), .A2(_AES_ENC_us30_n1093 ), .ZN(_AES_ENC_us30_n675 ) );
NAND2_X2 _AES_ENC_us30_U425  ( .A1(_AES_ENC_us30_n588 ), .A2(_AES_ENC_us30_n597 ), .ZN(_AES_ENC_us30_n1045 ) );
OR2_X2 _AES_ENC_us30_U424  ( .A1(_AES_ENC_us30_n1045 ), .A2(_AES_ENC_us30_n605 ), .ZN(_AES_ENC_us30_n674 ) );
NAND2_X2 _AES_ENC_us30_U423  ( .A1(_AES_ENC_sa30[1]), .A2(_AES_ENC_us30_n620 ), .ZN(_AES_ENC_us30_n667 ) );
NAND2_X2 _AES_ENC_us30_U422  ( .A1(_AES_ENC_us30_n619 ), .A2(_AES_ENC_us30_n667 ), .ZN(_AES_ENC_us30_n1071 ) );
NAND4_X2 _AES_ENC_us30_U412  ( .A1(_AES_ENC_us30_n675 ), .A2(_AES_ENC_us30_n674 ), .A3(_AES_ENC_us30_n673 ), .A4(_AES_ENC_us30_n672 ), .ZN(_AES_ENC_us30_n676 ) );
NAND2_X2 _AES_ENC_us30_U411  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n676 ), .ZN(_AES_ENC_us30_n677 ) );
NAND2_X2 _AES_ENC_us30_U408  ( .A1(_AES_ENC_us30_n800 ), .A2(_AES_ENC_us30_n1022 ), .ZN(_AES_ENC_us30_n680 ) );
NAND2_X2 _AES_ENC_us30_U407  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n680 ), .ZN(_AES_ENC_us30_n681 ) );
AND2_X2 _AES_ENC_us30_U402  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n684 ), .ZN(_AES_ENC_us30_n682 ) );
NAND4_X2 _AES_ENC_us30_U395  ( .A1(_AES_ENC_us30_n691 ), .A2(_AES_ENC_us30_n581 ), .A3(_AES_ENC_us30_n690 ), .A4(_AES_ENC_us30_n689 ), .ZN(_AES_ENC_us30_n692 ) );
NAND2_X2 _AES_ENC_us30_U394  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n692 ), .ZN(_AES_ENC_us30_n733 ) );
NAND2_X2 _AES_ENC_us30_U392  ( .A1(_AES_ENC_us30_n977 ), .A2(_AES_ENC_us30_n1050 ), .ZN(_AES_ENC_us30_n702 ) );
NAND2_X2 _AES_ENC_us30_U391  ( .A1(_AES_ENC_us30_n1093 ), .A2(_AES_ENC_us30_n1045 ), .ZN(_AES_ENC_us30_n701 ) );
NAND4_X2 _AES_ENC_us30_U381  ( .A1(_AES_ENC_us30_n702 ), .A2(_AES_ENC_us30_n701 ), .A3(_AES_ENC_us30_n700 ), .A4(_AES_ENC_us30_n699 ), .ZN(_AES_ENC_us30_n703 ) );
NAND2_X2 _AES_ENC_us30_U380  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n703 ), .ZN(_AES_ENC_us30_n732 ) );
AND2_X2 _AES_ENC_us30_U379  ( .A1(_AES_ENC_sa30[0]), .A2(_AES_ENC_sa30[6]),.ZN(_AES_ENC_us30_n1113 ) );
NAND2_X2 _AES_ENC_us30_U378  ( .A1(_AES_ENC_us30_n601 ), .A2(_AES_ENC_us30_n1030 ), .ZN(_AES_ENC_us30_n881 ) );
NAND2_X2 _AES_ENC_us30_U377  ( .A1(_AES_ENC_us30_n1093 ), .A2(_AES_ENC_us30_n881 ), .ZN(_AES_ENC_us30_n715 ) );
NAND2_X2 _AES_ENC_us30_U376  ( .A1(_AES_ENC_us30_n1010 ), .A2(_AES_ENC_us30_n600 ), .ZN(_AES_ENC_us30_n714 ) );
NAND2_X2 _AES_ENC_us30_U375  ( .A1(_AES_ENC_us30_n855 ), .A2(_AES_ENC_us30_n588 ), .ZN(_AES_ENC_us30_n1117 ) );
XNOR2_X2 _AES_ENC_us30_U371  ( .A(_AES_ENC_us30_n611 ), .B(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n824 ) );
NAND4_X2 _AES_ENC_us30_U362  ( .A1(_AES_ENC_us30_n715 ), .A2(_AES_ENC_us30_n714 ), .A3(_AES_ENC_us30_n713 ), .A4(_AES_ENC_us30_n712 ), .ZN(_AES_ENC_us30_n716 ) );
NAND2_X2 _AES_ENC_us30_U361  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n716 ), .ZN(_AES_ENC_us30_n731 ) );
AND2_X2 _AES_ENC_us30_U360  ( .A1(_AES_ENC_sa30[6]), .A2(_AES_ENC_us30_n574 ), .ZN(_AES_ENC_us30_n1131 ) );
NAND2_X2 _AES_ENC_us30_U359  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n717 ) );
NAND2_X2 _AES_ENC_us30_U358  ( .A1(_AES_ENC_us30_n1029 ), .A2(_AES_ENC_us30_n717 ), .ZN(_AES_ENC_us30_n728 ) );
NAND2_X2 _AES_ENC_us30_U357  ( .A1(_AES_ENC_sa30[1]), .A2(_AES_ENC_us30_n624 ), .ZN(_AES_ENC_us30_n1097 ) );
NAND2_X2 _AES_ENC_us30_U356  ( .A1(_AES_ENC_us30_n603 ), .A2(_AES_ENC_us30_n1097 ), .ZN(_AES_ENC_us30_n718 ) );
NAND2_X2 _AES_ENC_us30_U355  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n718 ), .ZN(_AES_ENC_us30_n727 ) );
NAND4_X2 _AES_ENC_us30_U344  ( .A1(_AES_ENC_us30_n728 ), .A2(_AES_ENC_us30_n727 ), .A3(_AES_ENC_us30_n726 ), .A4(_AES_ENC_us30_n725 ), .ZN(_AES_ENC_us30_n729 ) );
NAND2_X2 _AES_ENC_us30_U343  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n729 ), .ZN(_AES_ENC_us30_n730 ) );
NAND4_X2 _AES_ENC_us30_U342  ( .A1(_AES_ENC_us30_n733 ), .A2(_AES_ENC_us30_n732 ), .A3(_AES_ENC_us30_n731 ), .A4(_AES_ENC_us30_n730 ), .ZN(_AES_ENC_sa30_sub[1] ) );
NAND2_X2 _AES_ENC_us30_U341  ( .A1(_AES_ENC_sa30[7]), .A2(_AES_ENC_us30_n611 ), .ZN(_AES_ENC_us30_n734 ) );
NAND2_X2 _AES_ENC_us30_U340  ( .A1(_AES_ENC_us30_n734 ), .A2(_AES_ENC_us30_n607 ), .ZN(_AES_ENC_us30_n738 ) );
OR4_X2 _AES_ENC_us30_U339  ( .A1(_AES_ENC_us30_n738 ), .A2(_AES_ENC_us30_n626 ), .A3(_AES_ENC_us30_n826 ), .A4(_AES_ENC_us30_n1121 ), .ZN(_AES_ENC_us30_n746 ) );
NAND2_X2 _AES_ENC_us30_U337  ( .A1(_AES_ENC_us30_n1100 ), .A2(_AES_ENC_us30_n587 ), .ZN(_AES_ENC_us30_n992 ) );
OR2_X2 _AES_ENC_us30_U336  ( .A1(_AES_ENC_us30_n610 ), .A2(_AES_ENC_us30_n735 ), .ZN(_AES_ENC_us30_n737 ) );
NAND2_X2 _AES_ENC_us30_U334  ( .A1(_AES_ENC_us30_n619 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n753 ) );
NAND2_X2 _AES_ENC_us30_U333  ( .A1(_AES_ENC_us30_n582 ), .A2(_AES_ENC_us30_n753 ), .ZN(_AES_ENC_us30_n1080 ) );
NAND2_X2 _AES_ENC_us30_U332  ( .A1(_AES_ENC_us30_n1048 ), .A2(_AES_ENC_us30_n576 ), .ZN(_AES_ENC_us30_n736 ) );
NAND2_X2 _AES_ENC_us30_U331  ( .A1(_AES_ENC_us30_n737 ), .A2(_AES_ENC_us30_n736 ), .ZN(_AES_ENC_us30_n739 ) );
NAND2_X2 _AES_ENC_us30_U330  ( .A1(_AES_ENC_us30_n739 ), .A2(_AES_ENC_us30_n738 ), .ZN(_AES_ENC_us30_n745 ) );
NAND2_X2 _AES_ENC_us30_U326  ( .A1(_AES_ENC_us30_n1096 ), .A2(_AES_ENC_us30_n590 ), .ZN(_AES_ENC_us30_n906 ) );
NAND4_X2 _AES_ENC_us30_U323  ( .A1(_AES_ENC_us30_n746 ), .A2(_AES_ENC_us30_n992 ), .A3(_AES_ENC_us30_n745 ), .A4(_AES_ENC_us30_n744 ), .ZN(_AES_ENC_us30_n747 ) );
NAND2_X2 _AES_ENC_us30_U322  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n747 ), .ZN(_AES_ENC_us30_n793 ) );
NAND2_X2 _AES_ENC_us30_U321  ( .A1(_AES_ENC_us30_n584 ), .A2(_AES_ENC_us30_n855 ), .ZN(_AES_ENC_us30_n748 ) );
NAND2_X2 _AES_ENC_us30_U320  ( .A1(_AES_ENC_us30_n956 ), .A2(_AES_ENC_us30_n748 ), .ZN(_AES_ENC_us30_n760 ) );
NAND2_X2 _AES_ENC_us30_U313  ( .A1(_AES_ENC_us30_n590 ), .A2(_AES_ENC_us30_n753 ), .ZN(_AES_ENC_us30_n1023 ) );
NAND4_X2 _AES_ENC_us30_U308  ( .A1(_AES_ENC_us30_n760 ), .A2(_AES_ENC_us30_n992 ), .A3(_AES_ENC_us30_n759 ), .A4(_AES_ENC_us30_n758 ), .ZN(_AES_ENC_us30_n761 ) );
NAND2_X2 _AES_ENC_us30_U307  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n761 ), .ZN(_AES_ENC_us30_n792 ) );
NAND2_X2 _AES_ENC_us30_U306  ( .A1(_AES_ENC_us30_n584 ), .A2(_AES_ENC_us30_n603 ), .ZN(_AES_ENC_us30_n989 ) );
NAND2_X2 _AES_ENC_us30_U305  ( .A1(_AES_ENC_us30_n1050 ), .A2(_AES_ENC_us30_n989 ), .ZN(_AES_ENC_us30_n777 ) );
NAND2_X2 _AES_ENC_us30_U304  ( .A1(_AES_ENC_us30_n1093 ), .A2(_AES_ENC_us30_n762 ), .ZN(_AES_ENC_us30_n776 ) );
XNOR2_X2 _AES_ENC_us30_U301  ( .A(_AES_ENC_sa30[7]), .B(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n959 ) );
NAND4_X2 _AES_ENC_us30_U289  ( .A1(_AES_ENC_us30_n777 ), .A2(_AES_ENC_us30_n776 ), .A3(_AES_ENC_us30_n775 ), .A4(_AES_ENC_us30_n774 ), .ZN(_AES_ENC_us30_n778 ) );
NAND2_X2 _AES_ENC_us30_U288  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n778 ), .ZN(_AES_ENC_us30_n791 ) );
NAND2_X2 _AES_ENC_us30_U287  ( .A1(_AES_ENC_us30_n1056 ), .A2(_AES_ENC_us30_n1050 ), .ZN(_AES_ENC_us30_n788 ) );
NAND2_X2 _AES_ENC_us30_U286  ( .A1(_AES_ENC_us30_n1091 ), .A2(_AES_ENC_us30_n779 ), .ZN(_AES_ENC_us30_n787 ) );
NAND2_X2 _AES_ENC_us30_U285  ( .A1(_AES_ENC_us30_n956 ), .A2(_AES_ENC_sa30[1]), .ZN(_AES_ENC_us30_n786 ) );
NAND4_X2 _AES_ENC_us30_U278  ( .A1(_AES_ENC_us30_n788 ), .A2(_AES_ENC_us30_n787 ), .A3(_AES_ENC_us30_n786 ), .A4(_AES_ENC_us30_n785 ), .ZN(_AES_ENC_us30_n789 ) );
NAND2_X2 _AES_ENC_us30_U277  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n789 ), .ZN(_AES_ENC_us30_n790 ) );
NAND4_X2 _AES_ENC_us30_U276  ( .A1(_AES_ENC_us30_n793 ), .A2(_AES_ENC_us30_n792 ), .A3(_AES_ENC_us30_n791 ), .A4(_AES_ENC_us30_n790 ), .ZN(_AES_ENC_sa30_sub[2] ) );
NAND2_X2 _AES_ENC_us30_U275  ( .A1(_AES_ENC_us30_n1059 ), .A2(_AES_ENC_us30_n794 ), .ZN(_AES_ENC_us30_n810 ) );
NAND2_X2 _AES_ENC_us30_U274  ( .A1(_AES_ENC_us30_n1049 ), .A2(_AES_ENC_us30_n956 ), .ZN(_AES_ENC_us30_n809 ) );
OR2_X2 _AES_ENC_us30_U266  ( .A1(_AES_ENC_us30_n1096 ), .A2(_AES_ENC_us30_n606 ), .ZN(_AES_ENC_us30_n802 ) );
NAND2_X2 _AES_ENC_us30_U265  ( .A1(_AES_ENC_us30_n1053 ), .A2(_AES_ENC_us30_n800 ), .ZN(_AES_ENC_us30_n801 ) );
NAND2_X2 _AES_ENC_us30_U264  ( .A1(_AES_ENC_us30_n802 ), .A2(_AES_ENC_us30_n801 ), .ZN(_AES_ENC_us30_n805 ) );
NAND4_X2 _AES_ENC_us30_U261  ( .A1(_AES_ENC_us30_n810 ), .A2(_AES_ENC_us30_n809 ), .A3(_AES_ENC_us30_n808 ), .A4(_AES_ENC_us30_n807 ), .ZN(_AES_ENC_us30_n811 ) );
NAND2_X2 _AES_ENC_us30_U260  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n811 ), .ZN(_AES_ENC_us30_n852 ) );
OR2_X2 _AES_ENC_us30_U259  ( .A1(_AES_ENC_us30_n1023 ), .A2(_AES_ENC_us30_n617 ), .ZN(_AES_ENC_us30_n819 ) );
OR2_X2 _AES_ENC_us30_U257  ( .A1(_AES_ENC_us30_n570 ), .A2(_AES_ENC_us30_n930 ), .ZN(_AES_ENC_us30_n818 ) );
NAND2_X2 _AES_ENC_us30_U256  ( .A1(_AES_ENC_us30_n1013 ), .A2(_AES_ENC_us30_n1094 ), .ZN(_AES_ENC_us30_n817 ) );
NAND4_X2 _AES_ENC_us30_U249  ( .A1(_AES_ENC_us30_n819 ), .A2(_AES_ENC_us30_n818 ), .A3(_AES_ENC_us30_n817 ), .A4(_AES_ENC_us30_n816 ), .ZN(_AES_ENC_us30_n820 ) );
NAND2_X2 _AES_ENC_us30_U248  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n820 ), .ZN(_AES_ENC_us30_n851 ) );
NAND2_X2 _AES_ENC_us30_U247  ( .A1(_AES_ENC_us30_n956 ), .A2(_AES_ENC_us30_n1080 ), .ZN(_AES_ENC_us30_n835 ) );
NAND2_X2 _AES_ENC_us30_U246  ( .A1(_AES_ENC_us30_n570 ), .A2(_AES_ENC_us30_n1030 ), .ZN(_AES_ENC_us30_n1047 ) );
OR2_X2 _AES_ENC_us30_U245  ( .A1(_AES_ENC_us30_n1047 ), .A2(_AES_ENC_us30_n612 ), .ZN(_AES_ENC_us30_n834 ) );
NAND2_X2 _AES_ENC_us30_U244  ( .A1(_AES_ENC_us30_n1072 ), .A2(_AES_ENC_us30_n589 ), .ZN(_AES_ENC_us30_n833 ) );
NAND4_X2 _AES_ENC_us30_U233  ( .A1(_AES_ENC_us30_n835 ), .A2(_AES_ENC_us30_n834 ), .A3(_AES_ENC_us30_n833 ), .A4(_AES_ENC_us30_n832 ), .ZN(_AES_ENC_us30_n836 ) );
NAND2_X2 _AES_ENC_us30_U232  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n836 ), .ZN(_AES_ENC_us30_n850 ) );
NAND2_X2 _AES_ENC_us30_U231  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n623 ), .ZN(_AES_ENC_us30_n847 ) );
NAND2_X2 _AES_ENC_us30_U230  ( .A1(_AES_ENC_us30_n1050 ), .A2(_AES_ENC_us30_n1071 ), .ZN(_AES_ENC_us30_n846 ) );
OR2_X2 _AES_ENC_us30_U224  ( .A1(_AES_ENC_us30_n1053 ), .A2(_AES_ENC_us30_n911 ), .ZN(_AES_ENC_us30_n1077 ) );
NAND4_X2 _AES_ENC_us30_U220  ( .A1(_AES_ENC_us30_n847 ), .A2(_AES_ENC_us30_n846 ), .A3(_AES_ENC_us30_n845 ), .A4(_AES_ENC_us30_n844 ), .ZN(_AES_ENC_us30_n848 ) );
NAND2_X2 _AES_ENC_us30_U219  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n848 ), .ZN(_AES_ENC_us30_n849 ) );
NAND4_X2 _AES_ENC_us30_U218  ( .A1(_AES_ENC_us30_n852 ), .A2(_AES_ENC_us30_n851 ), .A3(_AES_ENC_us30_n850 ), .A4(_AES_ENC_us30_n849 ), .ZN(_AES_ENC_sa30_sub[3] ) );
NAND2_X2 _AES_ENC_us30_U216  ( .A1(_AES_ENC_us30_n1009 ), .A2(_AES_ENC_us30_n1072 ), .ZN(_AES_ENC_us30_n862 ) );
NAND2_X2 _AES_ENC_us30_U215  ( .A1(_AES_ENC_us30_n603 ), .A2(_AES_ENC_us30_n577 ), .ZN(_AES_ENC_us30_n853 ) );
NAND2_X2 _AES_ENC_us30_U214  ( .A1(_AES_ENC_us30_n1050 ), .A2(_AES_ENC_us30_n853 ), .ZN(_AES_ENC_us30_n861 ) );
NAND4_X2 _AES_ENC_us30_U206  ( .A1(_AES_ENC_us30_n862 ), .A2(_AES_ENC_us30_n861 ), .A3(_AES_ENC_us30_n860 ), .A4(_AES_ENC_us30_n859 ), .ZN(_AES_ENC_us30_n863 ) );
NAND2_X2 _AES_ENC_us30_U205  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n863 ), .ZN(_AES_ENC_us30_n905 ) );
NAND2_X2 _AES_ENC_us30_U204  ( .A1(_AES_ENC_us30_n1010 ), .A2(_AES_ENC_us30_n989 ), .ZN(_AES_ENC_us30_n874 ) );
NAND2_X2 _AES_ENC_us30_U203  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n610 ), .ZN(_AES_ENC_us30_n864 ) );
NAND2_X2 _AES_ENC_us30_U202  ( .A1(_AES_ENC_us30_n929 ), .A2(_AES_ENC_us30_n864 ), .ZN(_AES_ENC_us30_n873 ) );
NAND4_X2 _AES_ENC_us30_U193  ( .A1(_AES_ENC_us30_n874 ), .A2(_AES_ENC_us30_n873 ), .A3(_AES_ENC_us30_n872 ), .A4(_AES_ENC_us30_n871 ), .ZN(_AES_ENC_us30_n875 ) );
NAND2_X2 _AES_ENC_us30_U192  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n875 ), .ZN(_AES_ENC_us30_n904 ) );
NAND2_X2 _AES_ENC_us30_U191  ( .A1(_AES_ENC_us30_n583 ), .A2(_AES_ENC_us30_n1050 ), .ZN(_AES_ENC_us30_n889 ) );
NAND2_X2 _AES_ENC_us30_U190  ( .A1(_AES_ENC_us30_n1093 ), .A2(_AES_ENC_us30_n587 ), .ZN(_AES_ENC_us30_n876 ) );
NAND2_X2 _AES_ENC_us30_U189  ( .A1(_AES_ENC_us30_n604 ), .A2(_AES_ENC_us30_n876 ), .ZN(_AES_ENC_us30_n877 ) );
NAND2_X2 _AES_ENC_us30_U188  ( .A1(_AES_ENC_us30_n877 ), .A2(_AES_ENC_us30_n623 ), .ZN(_AES_ENC_us30_n888 ) );
NAND4_X2 _AES_ENC_us30_U179  ( .A1(_AES_ENC_us30_n889 ), .A2(_AES_ENC_us30_n888 ), .A3(_AES_ENC_us30_n887 ), .A4(_AES_ENC_us30_n886 ), .ZN(_AES_ENC_us30_n890 ) );
NAND2_X2 _AES_ENC_us30_U178  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n890 ), .ZN(_AES_ENC_us30_n903 ) );
OR2_X2 _AES_ENC_us30_U177  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n1059 ), .ZN(_AES_ENC_us30_n900 ) );
NAND2_X2 _AES_ENC_us30_U176  ( .A1(_AES_ENC_us30_n1073 ), .A2(_AES_ENC_us30_n1047 ), .ZN(_AES_ENC_us30_n899 ) );
NAND2_X2 _AES_ENC_us30_U175  ( .A1(_AES_ENC_us30_n1094 ), .A2(_AES_ENC_us30_n595 ), .ZN(_AES_ENC_us30_n898 ) );
NAND4_X2 _AES_ENC_us30_U167  ( .A1(_AES_ENC_us30_n900 ), .A2(_AES_ENC_us30_n899 ), .A3(_AES_ENC_us30_n898 ), .A4(_AES_ENC_us30_n897 ), .ZN(_AES_ENC_us30_n901 ) );
NAND2_X2 _AES_ENC_us30_U166  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n901 ), .ZN(_AES_ENC_us30_n902 ) );
NAND4_X2 _AES_ENC_us30_U165  ( .A1(_AES_ENC_us30_n905 ), .A2(_AES_ENC_us30_n904 ), .A3(_AES_ENC_us30_n903 ), .A4(_AES_ENC_us30_n902 ), .ZN(_AES_ENC_sa30_sub[4] ) );
NAND2_X2 _AES_ENC_us30_U164  ( .A1(_AES_ENC_us30_n1094 ), .A2(_AES_ENC_us30_n599 ), .ZN(_AES_ENC_us30_n922 ) );
NAND2_X2 _AES_ENC_us30_U163  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n989 ), .ZN(_AES_ENC_us30_n921 ) );
NAND4_X2 _AES_ENC_us30_U151  ( .A1(_AES_ENC_us30_n922 ), .A2(_AES_ENC_us30_n921 ), .A3(_AES_ENC_us30_n920 ), .A4(_AES_ENC_us30_n919 ), .ZN(_AES_ENC_us30_n923 ) );
NAND2_X2 _AES_ENC_us30_U150  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n923 ), .ZN(_AES_ENC_us30_n972 ) );
NAND2_X2 _AES_ENC_us30_U149  ( .A1(_AES_ENC_us30_n582 ), .A2(_AES_ENC_us30_n619 ), .ZN(_AES_ENC_us30_n924 ) );
NAND2_X2 _AES_ENC_us30_U148  ( .A1(_AES_ENC_us30_n1073 ), .A2(_AES_ENC_us30_n924 ), .ZN(_AES_ENC_us30_n939 ) );
NAND2_X2 _AES_ENC_us30_U147  ( .A1(_AES_ENC_us30_n926 ), .A2(_AES_ENC_us30_n925 ), .ZN(_AES_ENC_us30_n927 ) );
NAND2_X2 _AES_ENC_us30_U146  ( .A1(_AES_ENC_us30_n606 ), .A2(_AES_ENC_us30_n927 ), .ZN(_AES_ENC_us30_n928 ) );
NAND2_X2 _AES_ENC_us30_U145  ( .A1(_AES_ENC_us30_n928 ), .A2(_AES_ENC_us30_n1080 ), .ZN(_AES_ENC_us30_n938 ) );
OR2_X2 _AES_ENC_us30_U144  ( .A1(_AES_ENC_us30_n1117 ), .A2(_AES_ENC_us30_n615 ), .ZN(_AES_ENC_us30_n937 ) );
NAND4_X2 _AES_ENC_us30_U139  ( .A1(_AES_ENC_us30_n939 ), .A2(_AES_ENC_us30_n938 ), .A3(_AES_ENC_us30_n937 ), .A4(_AES_ENC_us30_n936 ), .ZN(_AES_ENC_us30_n940 ) );
NAND2_X2 _AES_ENC_us30_U138  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n940 ), .ZN(_AES_ENC_us30_n971 ) );
OR2_X2 _AES_ENC_us30_U137  ( .A1(_AES_ENC_us30_n605 ), .A2(_AES_ENC_us30_n941 ), .ZN(_AES_ENC_us30_n954 ) );
NAND2_X2 _AES_ENC_us30_U136  ( .A1(_AES_ENC_us30_n1096 ), .A2(_AES_ENC_us30_n577 ), .ZN(_AES_ENC_us30_n942 ) );
NAND2_X2 _AES_ENC_us30_U135  ( .A1(_AES_ENC_us30_n1048 ), .A2(_AES_ENC_us30_n942 ), .ZN(_AES_ENC_us30_n943 ) );
NAND2_X2 _AES_ENC_us30_U134  ( .A1(_AES_ENC_us30_n612 ), .A2(_AES_ENC_us30_n943 ), .ZN(_AES_ENC_us30_n944 ) );
NAND2_X2 _AES_ENC_us30_U133  ( .A1(_AES_ENC_us30_n944 ), .A2(_AES_ENC_us30_n580 ), .ZN(_AES_ENC_us30_n953 ) );
NAND4_X2 _AES_ENC_us30_U125  ( .A1(_AES_ENC_us30_n954 ), .A2(_AES_ENC_us30_n953 ), .A3(_AES_ENC_us30_n952 ), .A4(_AES_ENC_us30_n951 ), .ZN(_AES_ENC_us30_n955 ) );
NAND2_X2 _AES_ENC_us30_U124  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n955 ), .ZN(_AES_ENC_us30_n970 ) );
NAND2_X2 _AES_ENC_us30_U123  ( .A1(_AES_ENC_us30_n1094 ), .A2(_AES_ENC_us30_n1071 ), .ZN(_AES_ENC_us30_n967 ) );
NAND2_X2 _AES_ENC_us30_U122  ( .A1(_AES_ENC_us30_n956 ), .A2(_AES_ENC_us30_n1030 ), .ZN(_AES_ENC_us30_n966 ) );
NAND4_X2 _AES_ENC_us30_U114  ( .A1(_AES_ENC_us30_n967 ), .A2(_AES_ENC_us30_n966 ), .A3(_AES_ENC_us30_n965 ), .A4(_AES_ENC_us30_n964 ), .ZN(_AES_ENC_us30_n968 ) );
NAND2_X2 _AES_ENC_us30_U113  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n968 ), .ZN(_AES_ENC_us30_n969 ) );
NAND4_X2 _AES_ENC_us30_U112  ( .A1(_AES_ENC_us30_n972 ), .A2(_AES_ENC_us30_n971 ), .A3(_AES_ENC_us30_n970 ), .A4(_AES_ENC_us30_n969 ), .ZN(_AES_ENC_sa30_sub[5] ) );
NAND2_X2 _AES_ENC_us30_U111  ( .A1(_AES_ENC_us30_n570 ), .A2(_AES_ENC_us30_n1097 ), .ZN(_AES_ENC_us30_n973 ) );
NAND2_X2 _AES_ENC_us30_U110  ( .A1(_AES_ENC_us30_n1073 ), .A2(_AES_ENC_us30_n973 ), .ZN(_AES_ENC_us30_n987 ) );
NAND2_X2 _AES_ENC_us30_U109  ( .A1(_AES_ENC_us30_n974 ), .A2(_AES_ENC_us30_n1077 ), .ZN(_AES_ENC_us30_n975 ) );
NAND2_X2 _AES_ENC_us30_U108  ( .A1(_AES_ENC_us30_n613 ), .A2(_AES_ENC_us30_n975 ), .ZN(_AES_ENC_us30_n976 ) );
NAND2_X2 _AES_ENC_us30_U107  ( .A1(_AES_ENC_us30_n977 ), .A2(_AES_ENC_us30_n976 ), .ZN(_AES_ENC_us30_n986 ) );
NAND4_X2 _AES_ENC_us30_U99  ( .A1(_AES_ENC_us30_n987 ), .A2(_AES_ENC_us30_n986 ), .A3(_AES_ENC_us30_n985 ), .A4(_AES_ENC_us30_n984 ), .ZN(_AES_ENC_us30_n988 ) );
NAND2_X2 _AES_ENC_us30_U98  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n988 ), .ZN(_AES_ENC_us30_n1044 ) );
NAND2_X2 _AES_ENC_us30_U97  ( .A1(_AES_ENC_us30_n1073 ), .A2(_AES_ENC_us30_n989 ), .ZN(_AES_ENC_us30_n1004 ) );
NAND2_X2 _AES_ENC_us30_U96  ( .A1(_AES_ENC_us30_n1092 ), .A2(_AES_ENC_us30_n619 ), .ZN(_AES_ENC_us30_n1003 ) );
NAND4_X2 _AES_ENC_us30_U85  ( .A1(_AES_ENC_us30_n1004 ), .A2(_AES_ENC_us30_n1003 ), .A3(_AES_ENC_us30_n1002 ), .A4(_AES_ENC_us30_n1001 ), .ZN(_AES_ENC_us30_n1005 ) );
NAND2_X2 _AES_ENC_us30_U84  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n1005 ), .ZN(_AES_ENC_us30_n1043 ) );
NAND2_X2 _AES_ENC_us30_U83  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n596 ), .ZN(_AES_ENC_us30_n1020 ) );
NAND2_X2 _AES_ENC_us30_U82  ( .A1(_AES_ENC_us30_n1050 ), .A2(_AES_ENC_us30_n624 ), .ZN(_AES_ENC_us30_n1019 ) );
NAND2_X2 _AES_ENC_us30_U77  ( .A1(_AES_ENC_us30_n1059 ), .A2(_AES_ENC_us30_n1114 ), .ZN(_AES_ENC_us30_n1012 ) );
NAND2_X2 _AES_ENC_us30_U76  ( .A1(_AES_ENC_us30_n1010 ), .A2(_AES_ENC_us30_n592 ), .ZN(_AES_ENC_us30_n1011 ) );
NAND2_X2 _AES_ENC_us30_U75  ( .A1(_AES_ENC_us30_n1012 ), .A2(_AES_ENC_us30_n1011 ), .ZN(_AES_ENC_us30_n1016 ) );
NAND4_X2 _AES_ENC_us30_U70  ( .A1(_AES_ENC_us30_n1020 ), .A2(_AES_ENC_us30_n1019 ), .A3(_AES_ENC_us30_n1018 ), .A4(_AES_ENC_us30_n1017 ), .ZN(_AES_ENC_us30_n1021 ) );
NAND2_X2 _AES_ENC_us30_U69  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n1021 ), .ZN(_AES_ENC_us30_n1042 ) );
NAND2_X2 _AES_ENC_us30_U68  ( .A1(_AES_ENC_us30_n1022 ), .A2(_AES_ENC_us30_n1093 ), .ZN(_AES_ENC_us30_n1039 ) );
NAND2_X2 _AES_ENC_us30_U67  ( .A1(_AES_ENC_us30_n1050 ), .A2(_AES_ENC_us30_n1023 ), .ZN(_AES_ENC_us30_n1038 ) );
NAND2_X2 _AES_ENC_us30_U66  ( .A1(_AES_ENC_us30_n1024 ), .A2(_AES_ENC_us30_n1071 ), .ZN(_AES_ENC_us30_n1037 ) );
AND2_X2 _AES_ENC_us30_U60  ( .A1(_AES_ENC_us30_n1030 ), .A2(_AES_ENC_us30_n602 ), .ZN(_AES_ENC_us30_n1078 ) );
NAND4_X2 _AES_ENC_us30_U56  ( .A1(_AES_ENC_us30_n1039 ), .A2(_AES_ENC_us30_n1038 ), .A3(_AES_ENC_us30_n1037 ), .A4(_AES_ENC_us30_n1036 ), .ZN(_AES_ENC_us30_n1040 ) );
NAND2_X2 _AES_ENC_us30_U55  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n1040 ), .ZN(_AES_ENC_us30_n1041 ) );
NAND4_X2 _AES_ENC_us30_U54  ( .A1(_AES_ENC_us30_n1044 ), .A2(_AES_ENC_us30_n1043 ), .A3(_AES_ENC_us30_n1042 ), .A4(_AES_ENC_us30_n1041 ), .ZN(_AES_ENC_sa30_sub[6] ) );
NAND2_X2 _AES_ENC_us30_U53  ( .A1(_AES_ENC_us30_n1072 ), .A2(_AES_ENC_us30_n1045 ), .ZN(_AES_ENC_us30_n1068 ) );
NAND2_X2 _AES_ENC_us30_U52  ( .A1(_AES_ENC_us30_n1046 ), .A2(_AES_ENC_us30_n582 ), .ZN(_AES_ENC_us30_n1067 ) );
NAND2_X2 _AES_ENC_us30_U51  ( .A1(_AES_ENC_us30_n1094 ), .A2(_AES_ENC_us30_n1047 ), .ZN(_AES_ENC_us30_n1066 ) );
NAND4_X2 _AES_ENC_us30_U40  ( .A1(_AES_ENC_us30_n1068 ), .A2(_AES_ENC_us30_n1067 ), .A3(_AES_ENC_us30_n1066 ), .A4(_AES_ENC_us30_n1065 ), .ZN(_AES_ENC_us30_n1069 ) );
NAND2_X2 _AES_ENC_us30_U39  ( .A1(_AES_ENC_us30_n1070 ), .A2(_AES_ENC_us30_n1069 ), .ZN(_AES_ENC_us30_n1135 ) );
NAND2_X2 _AES_ENC_us30_U38  ( .A1(_AES_ENC_us30_n1072 ), .A2(_AES_ENC_us30_n1071 ), .ZN(_AES_ENC_us30_n1088 ) );
NAND2_X2 _AES_ENC_us30_U37  ( .A1(_AES_ENC_us30_n1073 ), .A2(_AES_ENC_us30_n595 ), .ZN(_AES_ENC_us30_n1087 ) );
NAND4_X2 _AES_ENC_us30_U28  ( .A1(_AES_ENC_us30_n1088 ), .A2(_AES_ENC_us30_n1087 ), .A3(_AES_ENC_us30_n1086 ), .A4(_AES_ENC_us30_n1085 ), .ZN(_AES_ENC_us30_n1089 ) );
NAND2_X2 _AES_ENC_us30_U27  ( .A1(_AES_ENC_us30_n1090 ), .A2(_AES_ENC_us30_n1089 ), .ZN(_AES_ENC_us30_n1134 ) );
NAND2_X2 _AES_ENC_us30_U26  ( .A1(_AES_ENC_us30_n1091 ), .A2(_AES_ENC_us30_n1093 ), .ZN(_AES_ENC_us30_n1111 ) );
NAND2_X2 _AES_ENC_us30_U25  ( .A1(_AES_ENC_us30_n1092 ), .A2(_AES_ENC_us30_n1120 ), .ZN(_AES_ENC_us30_n1110 ) );
AND2_X2 _AES_ENC_us30_U22  ( .A1(_AES_ENC_us30_n1097 ), .A2(_AES_ENC_us30_n1096 ), .ZN(_AES_ENC_us30_n1098 ) );
NAND4_X2 _AES_ENC_us30_U14  ( .A1(_AES_ENC_us30_n1111 ), .A2(_AES_ENC_us30_n1110 ), .A3(_AES_ENC_us30_n1109 ), .A4(_AES_ENC_us30_n1108 ), .ZN(_AES_ENC_us30_n1112 ) );
NAND2_X2 _AES_ENC_us30_U13  ( .A1(_AES_ENC_us30_n1113 ), .A2(_AES_ENC_us30_n1112 ), .ZN(_AES_ENC_us30_n1133 ) );
NAND2_X2 _AES_ENC_us30_U12  ( .A1(_AES_ENC_us30_n1115 ), .A2(_AES_ENC_us30_n1114 ), .ZN(_AES_ENC_us30_n1129 ) );
OR2_X2 _AES_ENC_us30_U11  ( .A1(_AES_ENC_us30_n608 ), .A2(_AES_ENC_us30_n1116 ), .ZN(_AES_ENC_us30_n1128 ) );
NAND4_X2 _AES_ENC_us30_U3  ( .A1(_AES_ENC_us30_n1129 ), .A2(_AES_ENC_us30_n1128 ), .A3(_AES_ENC_us30_n1127 ), .A4(_AES_ENC_us30_n1126 ), .ZN(_AES_ENC_us30_n1130 ) );
NAND2_X2 _AES_ENC_us30_U2  ( .A1(_AES_ENC_us30_n1131 ), .A2(_AES_ENC_us30_n1130 ), .ZN(_AES_ENC_us30_n1132 ) );
NAND4_X2 _AES_ENC_us30_U1  ( .A1(_AES_ENC_us30_n1135 ), .A2(_AES_ENC_us30_n1134 ), .A3(_AES_ENC_us30_n1133 ), .A4(_AES_ENC_us30_n1132 ), .ZN(_AES_ENC_sa30_sub[7] ) );
INV_X4 _AES_ENC_us31_U575  ( .A(_AES_ENC_sa31[7]), .ZN(_AES_ENC_us31_n627 ));
INV_X4 _AES_ENC_us31_U574  ( .A(_AES_ENC_us31_n1114 ), .ZN(_AES_ENC_us31_n625 ) );
INV_X4 _AES_ENC_us31_U573  ( .A(_AES_ENC_sa31[4]), .ZN(_AES_ENC_us31_n624 ));
INV_X4 _AES_ENC_us31_U572  ( .A(_AES_ENC_us31_n1025 ), .ZN(_AES_ENC_us31_n622 ) );
INV_X4 _AES_ENC_us31_U571  ( .A(_AES_ENC_us31_n1120 ), .ZN(_AES_ENC_us31_n620 ) );
INV_X4 _AES_ENC_us31_U570  ( .A(_AES_ENC_us31_n1121 ), .ZN(_AES_ENC_us31_n619 ) );
INV_X4 _AES_ENC_us31_U569  ( .A(_AES_ENC_us31_n1048 ), .ZN(_AES_ENC_us31_n618 ) );
INV_X4 _AES_ENC_us31_U568  ( .A(_AES_ENC_us31_n974 ), .ZN(_AES_ENC_us31_n616 ) );
INV_X4 _AES_ENC_us31_U567  ( .A(_AES_ENC_us31_n794 ), .ZN(_AES_ENC_us31_n614 ) );
INV_X4 _AES_ENC_us31_U566  ( .A(_AES_ENC_sa31[2]), .ZN(_AES_ENC_us31_n611 ));
INV_X4 _AES_ENC_us31_U565  ( .A(_AES_ENC_us31_n800 ), .ZN(_AES_ENC_us31_n610 ) );
INV_X4 _AES_ENC_us31_U564  ( .A(_AES_ENC_us31_n925 ), .ZN(_AES_ENC_us31_n609 ) );
INV_X4 _AES_ENC_us31_U563  ( .A(_AES_ENC_us31_n779 ), .ZN(_AES_ENC_us31_n607 ) );
INV_X4 _AES_ENC_us31_U562  ( .A(_AES_ENC_us31_n1022 ), .ZN(_AES_ENC_us31_n603 ) );
INV_X4 _AES_ENC_us31_U561  ( .A(_AES_ENC_us31_n1102 ), .ZN(_AES_ENC_us31_n602 ) );
INV_X4 _AES_ENC_us31_U560  ( .A(_AES_ENC_us31_n929 ), .ZN(_AES_ENC_us31_n601 ) );
INV_X4 _AES_ENC_us31_U559  ( .A(_AES_ENC_us31_n1056 ), .ZN(_AES_ENC_us31_n600 ) );
INV_X4 _AES_ENC_us31_U558  ( .A(_AES_ENC_us31_n1054 ), .ZN(_AES_ENC_us31_n599 ) );
INV_X4 _AES_ENC_us31_U557  ( .A(_AES_ENC_us31_n881 ), .ZN(_AES_ENC_us31_n598 ) );
INV_X4 _AES_ENC_us31_U556  ( .A(_AES_ENC_us31_n926 ), .ZN(_AES_ENC_us31_n597 ) );
INV_X4 _AES_ENC_us31_U555  ( .A(_AES_ENC_us31_n977 ), .ZN(_AES_ENC_us31_n595 ) );
INV_X4 _AES_ENC_us31_U554  ( .A(_AES_ENC_us31_n1031 ), .ZN(_AES_ENC_us31_n594 ) );
INV_X4 _AES_ENC_us31_U553  ( .A(_AES_ENC_us31_n1103 ), .ZN(_AES_ENC_us31_n593 ) );
INV_X4 _AES_ENC_us31_U552  ( .A(_AES_ENC_us31_n1009 ), .ZN(_AES_ENC_us31_n592 ) );
INV_X4 _AES_ENC_us31_U551  ( .A(_AES_ENC_us31_n990 ), .ZN(_AES_ENC_us31_n591 ) );
INV_X4 _AES_ENC_us31_U550  ( .A(_AES_ENC_us31_n1058 ), .ZN(_AES_ENC_us31_n590 ) );
INV_X4 _AES_ENC_us31_U549  ( .A(_AES_ENC_us31_n1074 ), .ZN(_AES_ENC_us31_n589 ) );
INV_X4 _AES_ENC_us31_U548  ( .A(_AES_ENC_us31_n1053 ), .ZN(_AES_ENC_us31_n588 ) );
INV_X4 _AES_ENC_us31_U547  ( .A(_AES_ENC_us31_n826 ), .ZN(_AES_ENC_us31_n587 ) );
INV_X4 _AES_ENC_us31_U546  ( .A(_AES_ENC_us31_n992 ), .ZN(_AES_ENC_us31_n586 ) );
INV_X4 _AES_ENC_us31_U545  ( .A(_AES_ENC_us31_n821 ), .ZN(_AES_ENC_us31_n585 ) );
INV_X4 _AES_ENC_us31_U544  ( .A(_AES_ENC_us31_n910 ), .ZN(_AES_ENC_us31_n584 ) );
INV_X4 _AES_ENC_us31_U543  ( .A(_AES_ENC_us31_n906 ), .ZN(_AES_ENC_us31_n583 ) );
INV_X4 _AES_ENC_us31_U542  ( .A(_AES_ENC_us31_n880 ), .ZN(_AES_ENC_us31_n581 ) );
INV_X4 _AES_ENC_us31_U541  ( .A(_AES_ENC_us31_n1013 ), .ZN(_AES_ENC_us31_n580 ) );
INV_X4 _AES_ENC_us31_U540  ( .A(_AES_ENC_us31_n1092 ), .ZN(_AES_ENC_us31_n579 ) );
INV_X4 _AES_ENC_us31_U539  ( .A(_AES_ENC_us31_n824 ), .ZN(_AES_ENC_us31_n578 ) );
INV_X4 _AES_ENC_us31_U538  ( .A(_AES_ENC_us31_n1091 ), .ZN(_AES_ENC_us31_n577 ) );
INV_X4 _AES_ENC_us31_U537  ( .A(_AES_ENC_us31_n1080 ), .ZN(_AES_ENC_us31_n576 ) );
INV_X4 _AES_ENC_us31_U536  ( .A(_AES_ENC_us31_n959 ), .ZN(_AES_ENC_us31_n575 ) );
INV_X4 _AES_ENC_us31_U535  ( .A(_AES_ENC_sa31[0]), .ZN(_AES_ENC_us31_n574 ));
NOR2_X2 _AES_ENC_us31_U534  ( .A1(_AES_ENC_sa31[0]), .A2(_AES_ENC_sa31[6]),.ZN(_AES_ENC_us31_n1090 ) );
NOR2_X2 _AES_ENC_us31_U533  ( .A1(_AES_ENC_us31_n574 ), .A2(_AES_ENC_sa31[6]), .ZN(_AES_ENC_us31_n1070 ) );
NOR2_X2 _AES_ENC_us31_U532  ( .A1(_AES_ENC_sa31[4]), .A2(_AES_ENC_sa31[3]),.ZN(_AES_ENC_us31_n1025 ) );
INV_X4 _AES_ENC_us31_U531  ( .A(_AES_ENC_us31_n569 ), .ZN(_AES_ENC_us31_n572 ) );
NOR2_X2 _AES_ENC_us31_U530  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n765 ) );
NOR2_X2 _AES_ENC_us31_U529  ( .A1(_AES_ENC_sa31[4]), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n764 ) );
NOR2_X2 _AES_ENC_us31_U528  ( .A1(_AES_ENC_us31_n765 ), .A2(_AES_ENC_us31_n764 ), .ZN(_AES_ENC_us31_n766 ) );
NOR2_X2 _AES_ENC_us31_U527  ( .A1(_AES_ENC_us31_n766 ), .A2(_AES_ENC_us31_n575 ), .ZN(_AES_ENC_us31_n767 ) );
NOR3_X2 _AES_ENC_us31_U526  ( .A1(_AES_ENC_us31_n627 ), .A2(_AES_ENC_sa31[5]), .A3(_AES_ENC_us31_n704 ), .ZN(_AES_ENC_us31_n706 ));
NOR2_X2 _AES_ENC_us31_U525  ( .A1(_AES_ENC_us31_n1117 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n707 ) );
NOR2_X2 _AES_ENC_us31_U524  ( .A1(_AES_ENC_sa31[4]), .A2(_AES_ENC_us31_n579 ), .ZN(_AES_ENC_us31_n705 ) );
NOR3_X2 _AES_ENC_us31_U523  ( .A1(_AES_ENC_us31_n707 ), .A2(_AES_ENC_us31_n706 ), .A3(_AES_ENC_us31_n705 ), .ZN(_AES_ENC_us31_n713 ) );
INV_X4 _AES_ENC_us31_U522  ( .A(_AES_ENC_sa31[3]), .ZN(_AES_ENC_us31_n621 ));
NAND3_X2 _AES_ENC_us31_U521  ( .A1(_AES_ENC_us31_n652 ), .A2(_AES_ENC_us31_n626 ), .A3(_AES_ENC_sa31[7]), .ZN(_AES_ENC_us31_n653 ));
NOR2_X2 _AES_ENC_us31_U520  ( .A1(_AES_ENC_us31_n611 ), .A2(_AES_ENC_sa31[5]), .ZN(_AES_ENC_us31_n925 ) );
NOR2_X2 _AES_ENC_us31_U519  ( .A1(_AES_ENC_sa31[5]), .A2(_AES_ENC_sa31[2]),.ZN(_AES_ENC_us31_n974 ) );
INV_X4 _AES_ENC_us31_U518  ( .A(_AES_ENC_sa31[5]), .ZN(_AES_ENC_us31_n626 ));
NOR2_X2 _AES_ENC_us31_U517  ( .A1(_AES_ENC_us31_n611 ), .A2(_AES_ENC_sa31[7]), .ZN(_AES_ENC_us31_n779 ) );
NAND3_X2 _AES_ENC_us31_U516  ( .A1(_AES_ENC_us31_n679 ), .A2(_AES_ENC_us31_n678 ), .A3(_AES_ENC_us31_n677 ), .ZN(_AES_ENC_sa31_sub[0] ) );
NOR2_X2 _AES_ENC_us31_U515  ( .A1(_AES_ENC_us31_n626 ), .A2(_AES_ENC_sa31[2]), .ZN(_AES_ENC_us31_n1048 ) );
NOR4_X2 _AES_ENC_us31_U512  ( .A1(_AES_ENC_us31_n633 ), .A2(_AES_ENC_us31_n632 ), .A3(_AES_ENC_us31_n631 ), .A4(_AES_ENC_us31_n630 ), .ZN(_AES_ENC_us31_n634 ) );
NOR2_X2 _AES_ENC_us31_U510  ( .A1(_AES_ENC_us31_n629 ), .A2(_AES_ENC_us31_n628 ), .ZN(_AES_ENC_us31_n635 ) );
NAND3_X2 _AES_ENC_us31_U509  ( .A1(_AES_ENC_sa31[2]), .A2(_AES_ENC_sa31[7]), .A3(_AES_ENC_us31_n1059 ), .ZN(_AES_ENC_us31_n636 ) );
NOR2_X2 _AES_ENC_us31_U508  ( .A1(_AES_ENC_sa31[7]), .A2(_AES_ENC_sa31[2]),.ZN(_AES_ENC_us31_n794 ) );
NOR2_X2 _AES_ENC_us31_U507  ( .A1(_AES_ENC_sa31[4]), .A2(_AES_ENC_sa31[1]),.ZN(_AES_ENC_us31_n1102 ) );
NOR2_X2 _AES_ENC_us31_U506  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_sa31[3]), .ZN(_AES_ENC_us31_n1053 ) );
NOR2_X2 _AES_ENC_us31_U505  ( .A1(_AES_ENC_us31_n607 ), .A2(_AES_ENC_sa31[5]), .ZN(_AES_ENC_us31_n1024 ) );
NOR2_X2 _AES_ENC_us31_U504  ( .A1(_AES_ENC_us31_n625 ), .A2(_AES_ENC_sa31[2]), .ZN(_AES_ENC_us31_n1093 ) );
NOR2_X2 _AES_ENC_us31_U503  ( .A1(_AES_ENC_us31_n614 ), .A2(_AES_ENC_sa31[5]), .ZN(_AES_ENC_us31_n1094 ) );
NOR2_X2 _AES_ENC_us31_U502  ( .A1(_AES_ENC_us31_n624 ), .A2(_AES_ENC_sa31[3]), .ZN(_AES_ENC_us31_n931 ) );
INV_X4 _AES_ENC_us31_U501  ( .A(_AES_ENC_us31_n570 ), .ZN(_AES_ENC_us31_n573 ) );
NOR2_X2 _AES_ENC_us31_U500  ( .A1(_AES_ENC_us31_n1053 ), .A2(_AES_ENC_us31_n1095 ), .ZN(_AES_ENC_us31_n639 ) );
NOR3_X2 _AES_ENC_us31_U499  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n573 ), .A3(_AES_ENC_us31_n1074 ), .ZN(_AES_ENC_us31_n641 ) );
NOR2_X2 _AES_ENC_us31_U498  ( .A1(_AES_ENC_us31_n639 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n640 ) );
NOR2_X2 _AES_ENC_us31_U497  ( .A1(_AES_ENC_us31_n641 ), .A2(_AES_ENC_us31_n640 ), .ZN(_AES_ENC_us31_n646 ) );
NOR3_X2 _AES_ENC_us31_U496  ( .A1(_AES_ENC_us31_n995 ), .A2(_AES_ENC_us31_n586 ), .A3(_AES_ENC_us31_n994 ), .ZN(_AES_ENC_us31_n1002 ) );
NOR2_X2 _AES_ENC_us31_U495  ( .A1(_AES_ENC_us31_n909 ), .A2(_AES_ENC_us31_n908 ), .ZN(_AES_ENC_us31_n920 ) );
NOR2_X2 _AES_ENC_us31_U494  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n823 ) );
NOR2_X2 _AES_ENC_us31_U492  ( .A1(_AES_ENC_us31_n624 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n822 ) );
NOR2_X2 _AES_ENC_us31_U491  ( .A1(_AES_ENC_us31_n823 ), .A2(_AES_ENC_us31_n822 ), .ZN(_AES_ENC_us31_n825 ) );
NOR2_X2 _AES_ENC_us31_U490  ( .A1(_AES_ENC_sa31[1]), .A2(_AES_ENC_us31_n623 ), .ZN(_AES_ENC_us31_n913 ) );
NOR2_X2 _AES_ENC_us31_U489  ( .A1(_AES_ENC_us31_n913 ), .A2(_AES_ENC_us31_n1091 ), .ZN(_AES_ENC_us31_n914 ) );
NOR2_X2 _AES_ENC_us31_U488  ( .A1(_AES_ENC_us31_n826 ), .A2(_AES_ENC_us31_n572 ), .ZN(_AES_ENC_us31_n827 ) );
NOR3_X2 _AES_ENC_us31_U487  ( .A1(_AES_ENC_us31_n769 ), .A2(_AES_ENC_us31_n768 ), .A3(_AES_ENC_us31_n767 ), .ZN(_AES_ENC_us31_n775 ) );
NOR2_X2 _AES_ENC_us31_U486  ( .A1(_AES_ENC_us31_n1056 ), .A2(_AES_ENC_us31_n1053 ), .ZN(_AES_ENC_us31_n749 ) );
NOR2_X2 _AES_ENC_us31_U483  ( .A1(_AES_ENC_us31_n749 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n752 ) );
INV_X4 _AES_ENC_us31_U482  ( .A(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n596 ));
NOR2_X2 _AES_ENC_us31_U480  ( .A1(_AES_ENC_us31_n1054 ), .A2(_AES_ENC_us31_n1053 ), .ZN(_AES_ENC_us31_n1055 ) );
OR2_X4 _AES_ENC_us31_U479  ( .A1(_AES_ENC_us31_n1094 ), .A2(_AES_ENC_us31_n1093 ), .ZN(_AES_ENC_us31_n571 ) );
AND2_X2 _AES_ENC_us31_U478  ( .A1(_AES_ENC_us31_n571 ), .A2(_AES_ENC_us31_n1095 ), .ZN(_AES_ENC_us31_n1101 ) );
NOR2_X2 _AES_ENC_us31_U477  ( .A1(_AES_ENC_us31_n1074 ), .A2(_AES_ENC_us31_n931 ), .ZN(_AES_ENC_us31_n796 ) );
NOR2_X2 _AES_ENC_us31_U474  ( .A1(_AES_ENC_us31_n796 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n797 ) );
NOR2_X2 _AES_ENC_us31_U473  ( .A1(_AES_ENC_us31_n932 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n933 ) );
NOR2_X2 _AES_ENC_us31_U472  ( .A1(_AES_ENC_us31_n929 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n935 ) );
NOR2_X2 _AES_ENC_us31_U471  ( .A1(_AES_ENC_us31_n931 ), .A2(_AES_ENC_us31_n930 ), .ZN(_AES_ENC_us31_n934 ) );
NOR3_X2 _AES_ENC_us31_U470  ( .A1(_AES_ENC_us31_n935 ), .A2(_AES_ENC_us31_n934 ), .A3(_AES_ENC_us31_n933 ), .ZN(_AES_ENC_us31_n936 ) );
NOR2_X2 _AES_ENC_us31_U469  ( .A1(_AES_ENC_us31_n624 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n1075 ) );
NOR2_X2 _AES_ENC_us31_U468  ( .A1(_AES_ENC_us31_n572 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n949 ) );
NOR2_X2 _AES_ENC_us31_U467  ( .A1(_AES_ENC_us31_n1049 ), .A2(_AES_ENC_us31_n618 ), .ZN(_AES_ENC_us31_n1051 ) );
NOR2_X2 _AES_ENC_us31_U466  ( .A1(_AES_ENC_us31_n1051 ), .A2(_AES_ENC_us31_n1050 ), .ZN(_AES_ENC_us31_n1052 ) );
NOR2_X2 _AES_ENC_us31_U465  ( .A1(_AES_ENC_us31_n1052 ), .A2(_AES_ENC_us31_n592 ), .ZN(_AES_ENC_us31_n1064 ) );
NOR2_X2 _AES_ENC_us31_U464  ( .A1(_AES_ENC_sa31[1]), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n631 ) );
NOR2_X2 _AES_ENC_us31_U463  ( .A1(_AES_ENC_us31_n1025 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n980 ) );
NOR2_X2 _AES_ENC_us31_U462  ( .A1(_AES_ENC_us31_n1073 ), .A2(_AES_ENC_us31_n1094 ), .ZN(_AES_ENC_us31_n795 ) );
NOR2_X2 _AES_ENC_us31_U461  ( .A1(_AES_ENC_us31_n795 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n799 ) );
NOR2_X2 _AES_ENC_us31_U460  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n981 ) );
NOR2_X2 _AES_ENC_us31_U459  ( .A1(_AES_ENC_us31_n1102 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n643 ) );
NOR2_X2 _AES_ENC_us31_U458  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n621 ), .ZN(_AES_ENC_us31_n642 ) );
NOR2_X2 _AES_ENC_us31_U455  ( .A1(_AES_ENC_us31_n911 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n644 ) );
NOR4_X2 _AES_ENC_us31_U448  ( .A1(_AES_ENC_us31_n644 ), .A2(_AES_ENC_us31_n643 ), .A3(_AES_ENC_us31_n804 ), .A4(_AES_ENC_us31_n642 ), .ZN(_AES_ENC_us31_n645 ) );
NOR2_X2 _AES_ENC_us31_U447  ( .A1(_AES_ENC_us31_n1102 ), .A2(_AES_ENC_us31_n910 ), .ZN(_AES_ENC_us31_n932 ) );
NOR2_X2 _AES_ENC_us31_U442  ( .A1(_AES_ENC_us31_n1102 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n755 ) );
NOR2_X2 _AES_ENC_us31_U441  ( .A1(_AES_ENC_us31_n931 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n743 ) );
NOR2_X2 _AES_ENC_us31_U438  ( .A1(_AES_ENC_us31_n1072 ), .A2(_AES_ENC_us31_n1094 ), .ZN(_AES_ENC_us31_n930 ) );
NOR2_X2 _AES_ENC_us31_U435  ( .A1(_AES_ENC_us31_n1074 ), .A2(_AES_ENC_us31_n1025 ), .ZN(_AES_ENC_us31_n891 ) );
NOR2_X2 _AES_ENC_us31_U434  ( .A1(_AES_ENC_us31_n891 ), .A2(_AES_ENC_us31_n609 ), .ZN(_AES_ENC_us31_n894 ) );
NOR3_X2 _AES_ENC_us31_U433  ( .A1(_AES_ENC_us31_n623 ), .A2(_AES_ENC_sa31[1]), .A3(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n683 ));
INV_X4 _AES_ENC_us31_U428  ( .A(_AES_ENC_us31_n931 ), .ZN(_AES_ENC_us31_n623 ) );
NOR2_X2 _AES_ENC_us31_U427  ( .A1(_AES_ENC_us31_n996 ), .A2(_AES_ENC_us31_n931 ), .ZN(_AES_ENC_us31_n704 ) );
NOR2_X2 _AES_ENC_us31_U421  ( .A1(_AES_ENC_us31_n931 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n685 ) );
NOR2_X2 _AES_ENC_us31_U420  ( .A1(_AES_ENC_us31_n1029 ), .A2(_AES_ENC_us31_n1025 ), .ZN(_AES_ENC_us31_n1079 ) );
NOR3_X2 _AES_ENC_us31_U419  ( .A1(_AES_ENC_us31_n589 ), .A2(_AES_ENC_us31_n1025 ), .A3(_AES_ENC_us31_n616 ), .ZN(_AES_ENC_us31_n945 ) );
NOR2_X2 _AES_ENC_us31_U418  ( .A1(_AES_ENC_us31_n626 ), .A2(_AES_ENC_us31_n611 ), .ZN(_AES_ENC_us31_n800 ) );
NOR3_X2 _AES_ENC_us31_U417  ( .A1(_AES_ENC_us31_n590 ), .A2(_AES_ENC_us31_n627 ), .A3(_AES_ENC_us31_n611 ), .ZN(_AES_ENC_us31_n798 ) );
NOR3_X2 _AES_ENC_us31_U416  ( .A1(_AES_ENC_us31_n610 ), .A2(_AES_ENC_us31_n572 ), .A3(_AES_ENC_us31_n575 ), .ZN(_AES_ENC_us31_n962 ) );
NOR3_X2 _AES_ENC_us31_U415  ( .A1(_AES_ENC_us31_n959 ), .A2(_AES_ENC_us31_n572 ), .A3(_AES_ENC_us31_n609 ), .ZN(_AES_ENC_us31_n768 ) );
NOR3_X2 _AES_ENC_us31_U414  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n572 ), .A3(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n694 ) );
NOR3_X2 _AES_ENC_us31_U413  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n572 ), .A3(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n895 ) );
NOR3_X2 _AES_ENC_us31_U410  ( .A1(_AES_ENC_us31_n1008 ), .A2(_AES_ENC_us31_n1007 ), .A3(_AES_ENC_us31_n1006 ), .ZN(_AES_ENC_us31_n1018 ) );
NOR4_X2 _AES_ENC_us31_U409  ( .A1(_AES_ENC_us31_n806 ), .A2(_AES_ENC_us31_n805 ), .A3(_AES_ENC_us31_n804 ), .A4(_AES_ENC_us31_n803 ), .ZN(_AES_ENC_us31_n807 ) );
NOR3_X2 _AES_ENC_us31_U406  ( .A1(_AES_ENC_us31_n799 ), .A2(_AES_ENC_us31_n798 ), .A3(_AES_ENC_us31_n797 ), .ZN(_AES_ENC_us31_n808 ) );
NOR2_X2 _AES_ENC_us31_U405  ( .A1(_AES_ENC_us31_n669 ), .A2(_AES_ENC_us31_n668 ), .ZN(_AES_ENC_us31_n673 ) );
NOR4_X2 _AES_ENC_us31_U404  ( .A1(_AES_ENC_us31_n946 ), .A2(_AES_ENC_us31_n1046 ), .A3(_AES_ENC_us31_n671 ), .A4(_AES_ENC_us31_n670 ), .ZN(_AES_ENC_us31_n672 ) );
NOR4_X2 _AES_ENC_us31_U403  ( .A1(_AES_ENC_us31_n711 ), .A2(_AES_ENC_us31_n710 ), .A3(_AES_ENC_us31_n709 ), .A4(_AES_ENC_us31_n708 ), .ZN(_AES_ENC_us31_n712 ) );
NOR4_X2 _AES_ENC_us31_U401  ( .A1(_AES_ENC_us31_n963 ), .A2(_AES_ENC_us31_n962 ), .A3(_AES_ENC_us31_n961 ), .A4(_AES_ENC_us31_n960 ), .ZN(_AES_ENC_us31_n964 ) );
NOR3_X2 _AES_ENC_us31_U400  ( .A1(_AES_ENC_us31_n1101 ), .A2(_AES_ENC_us31_n1100 ), .A3(_AES_ENC_us31_n1099 ), .ZN(_AES_ENC_us31_n1109 ) );
NOR4_X2 _AES_ENC_us31_U399  ( .A1(_AES_ENC_us31_n843 ), .A2(_AES_ENC_us31_n842 ), .A3(_AES_ENC_us31_n841 ), .A4(_AES_ENC_us31_n840 ), .ZN(_AES_ENC_us31_n844 ) );
NOR3_X2 _AES_ENC_us31_U398  ( .A1(_AES_ENC_us31_n743 ), .A2(_AES_ENC_us31_n742 ), .A3(_AES_ENC_us31_n741 ), .ZN(_AES_ENC_us31_n744 ) );
NOR2_X2 _AES_ENC_us31_U397  ( .A1(_AES_ENC_us31_n697 ), .A2(_AES_ENC_us31_n658 ), .ZN(_AES_ENC_us31_n659 ) );
NOR2_X2 _AES_ENC_us31_U396  ( .A1(_AES_ENC_us31_n1078 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n1033 ) );
NOR2_X2 _AES_ENC_us31_U393  ( .A1(_AES_ENC_us31_n1031 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n1032 ) );
NOR3_X2 _AES_ENC_us31_U390  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n1025 ), .A3(_AES_ENC_us31_n1074 ), .ZN(_AES_ENC_us31_n1035 ) );
NOR4_X2 _AES_ENC_us31_U389  ( .A1(_AES_ENC_us31_n1035 ), .A2(_AES_ENC_us31_n1034 ), .A3(_AES_ENC_us31_n1033 ), .A4(_AES_ENC_us31_n1032 ), .ZN(_AES_ENC_us31_n1036 ) );
NOR2_X2 _AES_ENC_us31_U388  ( .A1(_AES_ENC_us31_n598 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n885 ) );
NOR2_X2 _AES_ENC_us31_U387  ( .A1(_AES_ENC_us31_n623 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n882 ) );
NOR2_X2 _AES_ENC_us31_U386  ( .A1(_AES_ENC_us31_n1053 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n884 ) );
NOR4_X2 _AES_ENC_us31_U385  ( .A1(_AES_ENC_us31_n885 ), .A2(_AES_ENC_us31_n884 ), .A3(_AES_ENC_us31_n883 ), .A4(_AES_ENC_us31_n882 ), .ZN(_AES_ENC_us31_n886 ) );
NOR2_X2 _AES_ENC_us31_U384  ( .A1(_AES_ENC_us31_n825 ), .A2(_AES_ENC_us31_n578 ), .ZN(_AES_ENC_us31_n830 ) );
NOR2_X2 _AES_ENC_us31_U383  ( .A1(_AES_ENC_us31_n827 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n829 ) );
NOR2_X2 _AES_ENC_us31_U382  ( .A1(_AES_ENC_us31_n572 ), .A2(_AES_ENC_us31_n579 ), .ZN(_AES_ENC_us31_n828 ) );
NOR4_X2 _AES_ENC_us31_U374  ( .A1(_AES_ENC_us31_n831 ), .A2(_AES_ENC_us31_n830 ), .A3(_AES_ENC_us31_n829 ), .A4(_AES_ENC_us31_n828 ), .ZN(_AES_ENC_us31_n832 ) );
NOR2_X2 _AES_ENC_us31_U373  ( .A1(_AES_ENC_us31_n606 ), .A2(_AES_ENC_us31_n582 ), .ZN(_AES_ENC_us31_n1104 ) );
NOR2_X2 _AES_ENC_us31_U372  ( .A1(_AES_ENC_us31_n1102 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n1106 ) );
NOR2_X2 _AES_ENC_us31_U370  ( .A1(_AES_ENC_us31_n1103 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n1105 ) );
NOR4_X2 _AES_ENC_us31_U369  ( .A1(_AES_ENC_us31_n1107 ), .A2(_AES_ENC_us31_n1106 ), .A3(_AES_ENC_us31_n1105 ), .A4(_AES_ENC_us31_n1104 ), .ZN(_AES_ENC_us31_n1108 ) );
NOR3_X2 _AES_ENC_us31_U368  ( .A1(_AES_ENC_us31_n959 ), .A2(_AES_ENC_us31_n621 ), .A3(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n963 ) );
NOR2_X2 _AES_ENC_us31_U367  ( .A1(_AES_ENC_us31_n626 ), .A2(_AES_ENC_us31_n627 ), .ZN(_AES_ENC_us31_n1114 ) );
INV_X4 _AES_ENC_us31_U366  ( .A(_AES_ENC_us31_n1024 ), .ZN(_AES_ENC_us31_n606 ) );
NOR3_X2 _AES_ENC_us31_U365  ( .A1(_AES_ENC_us31_n910 ), .A2(_AES_ENC_us31_n1059 ), .A3(_AES_ENC_us31_n611 ), .ZN(_AES_ENC_us31_n1115 ) );
INV_X4 _AES_ENC_us31_U364  ( .A(_AES_ENC_us31_n1094 ), .ZN(_AES_ENC_us31_n613 ) );
NOR2_X2 _AES_ENC_us31_U363  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n931 ), .ZN(_AES_ENC_us31_n1100 ) );
INV_X4 _AES_ENC_us31_U354  ( .A(_AES_ENC_us31_n1093 ), .ZN(_AES_ENC_us31_n617 ) );
NOR2_X2 _AES_ENC_us31_U353  ( .A1(_AES_ENC_us31_n569 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n929 ) );
NOR2_X2 _AES_ENC_us31_U352  ( .A1(_AES_ENC_us31_n620 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n926 ) );
NOR2_X2 _AES_ENC_us31_U351  ( .A1(_AES_ENC_us31_n572 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n1095 ) );
NOR2_X2 _AES_ENC_us31_U350  ( .A1(_AES_ENC_us31_n609 ), .A2(_AES_ENC_us31_n627 ), .ZN(_AES_ENC_us31_n1010 ) );
NOR2_X2 _AES_ENC_us31_U349  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n1103 ) );
NOR2_X2 _AES_ENC_us31_U348  ( .A1(_AES_ENC_us31_n622 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n1059 ) );
NOR2_X2 _AES_ENC_us31_U347  ( .A1(_AES_ENC_sa31[1]), .A2(_AES_ENC_us31_n1120 ), .ZN(_AES_ENC_us31_n1022 ) );
NOR2_X2 _AES_ENC_us31_U346  ( .A1(_AES_ENC_us31_n619 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n911 ) );
NOR2_X2 _AES_ENC_us31_U345  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_us31_n1025 ), .ZN(_AES_ENC_us31_n826 ) );
NOR2_X2 _AES_ENC_us31_U338  ( .A1(_AES_ENC_us31_n626 ), .A2(_AES_ENC_us31_n607 ), .ZN(_AES_ENC_us31_n1072 ) );
NOR2_X2 _AES_ENC_us31_U335  ( .A1(_AES_ENC_us31_n627 ), .A2(_AES_ENC_us31_n616 ), .ZN(_AES_ENC_us31_n956 ) );
NOR2_X2 _AES_ENC_us31_U329  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_us31_n624 ), .ZN(_AES_ENC_us31_n1121 ) );
NOR2_X2 _AES_ENC_us31_U328  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_us31_n624 ), .ZN(_AES_ENC_us31_n1058 ) );
NOR2_X2 _AES_ENC_us31_U327  ( .A1(_AES_ENC_us31_n625 ), .A2(_AES_ENC_us31_n611 ), .ZN(_AES_ENC_us31_n1073 ) );
NOR2_X2 _AES_ENC_us31_U325  ( .A1(_AES_ENC_sa31[1]), .A2(_AES_ENC_us31_n1025 ), .ZN(_AES_ENC_us31_n1054 ) );
NOR2_X2 _AES_ENC_us31_U324  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_us31_n931 ), .ZN(_AES_ENC_us31_n1029 ) );
NOR2_X2 _AES_ENC_us31_U319  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n1056 ) );
NOR2_X2 _AES_ENC_us31_U318  ( .A1(_AES_ENC_us31_n614 ), .A2(_AES_ENC_us31_n626 ), .ZN(_AES_ENC_us31_n1050 ) );
NOR2_X2 _AES_ENC_us31_U317  ( .A1(_AES_ENC_us31_n1121 ), .A2(_AES_ENC_us31_n1025 ), .ZN(_AES_ENC_us31_n1120 ) );
NOR2_X2 _AES_ENC_us31_U316  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_us31_n572 ), .ZN(_AES_ENC_us31_n1074 ) );
NOR2_X2 _AES_ENC_us31_U315  ( .A1(_AES_ENC_us31_n1058 ), .A2(_AES_ENC_us31_n1054 ), .ZN(_AES_ENC_us31_n878 ) );
NOR2_X2 _AES_ENC_us31_U314  ( .A1(_AES_ENC_us31_n878 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n879 ) );
NOR2_X2 _AES_ENC_us31_U312  ( .A1(_AES_ENC_us31_n880 ), .A2(_AES_ENC_us31_n879 ), .ZN(_AES_ENC_us31_n887 ) );
NOR2_X2 _AES_ENC_us31_U311  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n588 ), .ZN(_AES_ENC_us31_n957 ) );
NOR2_X2 _AES_ENC_us31_U310  ( .A1(_AES_ENC_us31_n958 ), .A2(_AES_ENC_us31_n957 ), .ZN(_AES_ENC_us31_n965 ) );
NOR3_X2 _AES_ENC_us31_U309  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n1091 ), .A3(_AES_ENC_us31_n1022 ), .ZN(_AES_ENC_us31_n720 ) );
NOR3_X2 _AES_ENC_us31_U303  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n1054 ), .A3(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n719 ) );
NOR2_X2 _AES_ENC_us31_U302  ( .A1(_AES_ENC_us31_n720 ), .A2(_AES_ENC_us31_n719 ), .ZN(_AES_ENC_us31_n726 ) );
NOR2_X2 _AES_ENC_us31_U300  ( .A1(_AES_ENC_us31_n614 ), .A2(_AES_ENC_us31_n591 ), .ZN(_AES_ENC_us31_n865 ) );
NOR2_X2 _AES_ENC_us31_U299  ( .A1(_AES_ENC_us31_n1059 ), .A2(_AES_ENC_us31_n1058 ), .ZN(_AES_ENC_us31_n1060 ) );
NOR2_X2 _AES_ENC_us31_U298  ( .A1(_AES_ENC_us31_n1095 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n668 ) );
NOR2_X2 _AES_ENC_us31_U297  ( .A1(_AES_ENC_us31_n911 ), .A2(_AES_ENC_us31_n910 ), .ZN(_AES_ENC_us31_n912 ) );
NOR2_X2 _AES_ENC_us31_U296  ( .A1(_AES_ENC_us31_n912 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n916 ) );
NOR2_X2 _AES_ENC_us31_U295  ( .A1(_AES_ENC_us31_n826 ), .A2(_AES_ENC_us31_n573 ), .ZN(_AES_ENC_us31_n750 ) );
NOR2_X2 _AES_ENC_us31_U294  ( .A1(_AES_ENC_us31_n750 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n751 ) );
NOR2_X2 _AES_ENC_us31_U293  ( .A1(_AES_ENC_us31_n907 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n908 ) );
NOR2_X2 _AES_ENC_us31_U292  ( .A1(_AES_ENC_us31_n990 ), .A2(_AES_ENC_us31_n926 ), .ZN(_AES_ENC_us31_n780 ) );
NOR2_X2 _AES_ENC_us31_U291  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n584 ), .ZN(_AES_ENC_us31_n838 ) );
NOR2_X2 _AES_ENC_us31_U290  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n602 ), .ZN(_AES_ENC_us31_n837 ) );
NOR2_X2 _AES_ENC_us31_U284  ( .A1(_AES_ENC_us31_n838 ), .A2(_AES_ENC_us31_n837 ), .ZN(_AES_ENC_us31_n845 ) );
NOR2_X2 _AES_ENC_us31_U283  ( .A1(_AES_ENC_us31_n1022 ), .A2(_AES_ENC_us31_n1058 ), .ZN(_AES_ENC_us31_n740 ) );
NOR2_X2 _AES_ENC_us31_U282  ( .A1(_AES_ENC_us31_n740 ), .A2(_AES_ENC_us31_n616 ), .ZN(_AES_ENC_us31_n742 ) );
NOR2_X2 _AES_ENC_us31_U281  ( .A1(_AES_ENC_us31_n1098 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n1099 ) );
NOR2_X2 _AES_ENC_us31_U280  ( .A1(_AES_ENC_us31_n1120 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n993 ) );
NOR2_X2 _AES_ENC_us31_U279  ( .A1(_AES_ENC_us31_n993 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n994 ) );
NOR2_X2 _AES_ENC_us31_U273  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n620 ), .ZN(_AES_ENC_us31_n1026 ) );
NOR2_X2 _AES_ENC_us31_U272  ( .A1(_AES_ENC_us31_n573 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n1027 ) );
NOR2_X2 _AES_ENC_us31_U271  ( .A1(_AES_ENC_us31_n1027 ), .A2(_AES_ENC_us31_n1026 ), .ZN(_AES_ENC_us31_n1028 ) );
NOR2_X2 _AES_ENC_us31_U270  ( .A1(_AES_ENC_us31_n1029 ), .A2(_AES_ENC_us31_n1028 ), .ZN(_AES_ENC_us31_n1034 ) );
NOR4_X2 _AES_ENC_us31_U269  ( .A1(_AES_ENC_us31_n757 ), .A2(_AES_ENC_us31_n756 ), .A3(_AES_ENC_us31_n755 ), .A4(_AES_ENC_us31_n754 ), .ZN(_AES_ENC_us31_n758 ) );
NOR2_X2 _AES_ENC_us31_U268  ( .A1(_AES_ENC_us31_n752 ), .A2(_AES_ENC_us31_n751 ), .ZN(_AES_ENC_us31_n759 ) );
NOR2_X2 _AES_ENC_us31_U267  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n1071 ), .ZN(_AES_ENC_us31_n669 ) );
NOR2_X2 _AES_ENC_us31_U263  ( .A1(_AES_ENC_us31_n1056 ), .A2(_AES_ENC_us31_n990 ), .ZN(_AES_ENC_us31_n991 ) );
NOR2_X2 _AES_ENC_us31_U262  ( .A1(_AES_ENC_us31_n991 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n995 ) );
NOR2_X2 _AES_ENC_us31_U258  ( .A1(_AES_ENC_us31_n607 ), .A2(_AES_ENC_us31_n590 ), .ZN(_AES_ENC_us31_n1008 ) );
NOR2_X2 _AES_ENC_us31_U255  ( .A1(_AES_ENC_us31_n839 ), .A2(_AES_ENC_us31_n582 ), .ZN(_AES_ENC_us31_n693 ) );
NOR2_X2 _AES_ENC_us31_U254  ( .A1(_AES_ENC_us31_n606 ), .A2(_AES_ENC_us31_n906 ), .ZN(_AES_ENC_us31_n741 ) );
NOR2_X2 _AES_ENC_us31_U253  ( .A1(_AES_ENC_us31_n1054 ), .A2(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n763 ) );
NOR2_X2 _AES_ENC_us31_U252  ( .A1(_AES_ENC_us31_n763 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n769 ) );
NOR2_X2 _AES_ENC_us31_U251  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n577 ), .ZN(_AES_ENC_us31_n1007 ) );
NOR2_X2 _AES_ENC_us31_U250  ( .A1(_AES_ENC_us31_n609 ), .A2(_AES_ENC_us31_n580 ), .ZN(_AES_ENC_us31_n1123 ) );
NOR2_X2 _AES_ENC_us31_U243  ( .A1(_AES_ENC_us31_n609 ), .A2(_AES_ENC_us31_n590 ), .ZN(_AES_ENC_us31_n710 ) );
INV_X4 _AES_ENC_us31_U242  ( .A(_AES_ENC_us31_n1029 ), .ZN(_AES_ENC_us31_n582 ) );
NOR2_X2 _AES_ENC_us31_U241  ( .A1(_AES_ENC_us31_n616 ), .A2(_AES_ENC_us31_n597 ), .ZN(_AES_ENC_us31_n883 ) );
NOR2_X2 _AES_ENC_us31_U240  ( .A1(_AES_ENC_us31_n593 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n1125 ) );
NOR2_X2 _AES_ENC_us31_U239  ( .A1(_AES_ENC_us31_n990 ), .A2(_AES_ENC_us31_n929 ), .ZN(_AES_ENC_us31_n892 ) );
NOR2_X2 _AES_ENC_us31_U238  ( .A1(_AES_ENC_us31_n892 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n893 ) );
NOR2_X2 _AES_ENC_us31_U237  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n602 ), .ZN(_AES_ENC_us31_n950 ) );
NOR2_X2 _AES_ENC_us31_U236  ( .A1(_AES_ENC_us31_n1079 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n1082 ) );
NOR2_X2 _AES_ENC_us31_U235  ( .A1(_AES_ENC_us31_n910 ), .A2(_AES_ENC_us31_n1056 ), .ZN(_AES_ENC_us31_n941 ) );
NOR2_X2 _AES_ENC_us31_U234  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n1077 ), .ZN(_AES_ENC_us31_n841 ) );
NOR2_X2 _AES_ENC_us31_U229  ( .A1(_AES_ENC_us31_n623 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n630 ) );
NOR2_X2 _AES_ENC_us31_U228  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n602 ), .ZN(_AES_ENC_us31_n806 ) );
NOR2_X2 _AES_ENC_us31_U227  ( .A1(_AES_ENC_us31_n623 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n948 ) );
NOR2_X2 _AES_ENC_us31_U226  ( .A1(_AES_ENC_us31_n606 ), .A2(_AES_ENC_us31_n589 ), .ZN(_AES_ENC_us31_n997 ) );
NOR2_X2 _AES_ENC_us31_U225  ( .A1(_AES_ENC_us31_n1121 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n1122 ) );
NOR2_X2 _AES_ENC_us31_U223  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n1023 ), .ZN(_AES_ENC_us31_n756 ) );
NOR2_X2 _AES_ENC_us31_U222  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n602 ), .ZN(_AES_ENC_us31_n870 ) );
NOR2_X2 _AES_ENC_us31_U221  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n569 ), .ZN(_AES_ENC_us31_n947 ) );
NOR2_X2 _AES_ENC_us31_U217  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n1077 ), .ZN(_AES_ENC_us31_n1084 ) );
NOR2_X2 _AES_ENC_us31_U213  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n855 ), .ZN(_AES_ENC_us31_n709 ) );
NOR2_X2 _AES_ENC_us31_U212  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n589 ), .ZN(_AES_ENC_us31_n868 ) );
NOR2_X2 _AES_ENC_us31_U211  ( .A1(_AES_ENC_us31_n1120 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n1124 ) );
NOR2_X2 _AES_ENC_us31_U210  ( .A1(_AES_ENC_us31_n1120 ), .A2(_AES_ENC_us31_n839 ), .ZN(_AES_ENC_us31_n842 ) );
NOR2_X2 _AES_ENC_us31_U209  ( .A1(_AES_ENC_us31_n1120 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n696 ) );
NOR2_X2 _AES_ENC_us31_U208  ( .A1(_AES_ENC_us31_n1074 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n1076 ) );
NOR2_X2 _AES_ENC_us31_U207  ( .A1(_AES_ENC_us31_n1074 ), .A2(_AES_ENC_us31_n620 ), .ZN(_AES_ENC_us31_n781 ) );
NOR3_X2 _AES_ENC_us31_U201  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n1056 ), .A3(_AES_ENC_us31_n990 ), .ZN(_AES_ENC_us31_n979 ) );
NOR3_X2 _AES_ENC_us31_U200  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n1058 ), .A3(_AES_ENC_us31_n1059 ), .ZN(_AES_ENC_us31_n854 ) );
NOR2_X2 _AES_ENC_us31_U199  ( .A1(_AES_ENC_us31_n996 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n869 ) );
NOR2_X2 _AES_ENC_us31_U198  ( .A1(_AES_ENC_us31_n1056 ), .A2(_AES_ENC_us31_n1074 ), .ZN(_AES_ENC_us31_n1057 ) );
NOR3_X2 _AES_ENC_us31_U197  ( .A1(_AES_ENC_us31_n607 ), .A2(_AES_ENC_us31_n1120 ), .A3(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n978 ) );
NOR2_X2 _AES_ENC_us31_U196  ( .A1(_AES_ENC_us31_n996 ), .A2(_AES_ENC_us31_n911 ), .ZN(_AES_ENC_us31_n1116 ) );
NOR2_X2 _AES_ENC_us31_U195  ( .A1(_AES_ENC_us31_n1074 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n754 ) );
NOR2_X2 _AES_ENC_us31_U194  ( .A1(_AES_ENC_us31_n926 ), .A2(_AES_ENC_us31_n1103 ), .ZN(_AES_ENC_us31_n977 ) );
NOR2_X2 _AES_ENC_us31_U187  ( .A1(_AES_ENC_us31_n839 ), .A2(_AES_ENC_us31_n824 ), .ZN(_AES_ENC_us31_n1092 ) );
NOR2_X2 _AES_ENC_us31_U186  ( .A1(_AES_ENC_us31_n573 ), .A2(_AES_ENC_us31_n1074 ), .ZN(_AES_ENC_us31_n684 ) );
NOR2_X2 _AES_ENC_us31_U185  ( .A1(_AES_ENC_us31_n826 ), .A2(_AES_ENC_us31_n1059 ), .ZN(_AES_ENC_us31_n907 ) );
NOR3_X2 _AES_ENC_us31_U184  ( .A1(_AES_ENC_us31_n625 ), .A2(_AES_ENC_us31_n1115 ), .A3(_AES_ENC_us31_n585 ), .ZN(_AES_ENC_us31_n831 ) );
NOR3_X2 _AES_ENC_us31_U183  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n1056 ), .A3(_AES_ENC_us31_n990 ), .ZN(_AES_ENC_us31_n896 ) );
NOR3_X2 _AES_ENC_us31_U182  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n573 ), .A3(_AES_ENC_us31_n1013 ), .ZN(_AES_ENC_us31_n670 ) );
NOR3_X2 _AES_ENC_us31_U181  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n1091 ), .A3(_AES_ENC_us31_n1022 ), .ZN(_AES_ENC_us31_n843 ) );
NOR2_X2 _AES_ENC_us31_U180  ( .A1(_AES_ENC_us31_n1029 ), .A2(_AES_ENC_us31_n1095 ), .ZN(_AES_ENC_us31_n735 ) );
NOR2_X2 _AES_ENC_us31_U174  ( .A1(_AES_ENC_us31_n1100 ), .A2(_AES_ENC_us31_n854 ), .ZN(_AES_ENC_us31_n860 ) );
NAND3_X2 _AES_ENC_us31_U173  ( .A1(_AES_ENC_us31_n569 ), .A2(_AES_ENC_us31_n582 ), .A3(_AES_ENC_us31_n681 ), .ZN(_AES_ENC_us31_n691 ) );
NOR2_X2 _AES_ENC_us31_U172  ( .A1(_AES_ENC_us31_n683 ), .A2(_AES_ENC_us31_n682 ), .ZN(_AES_ENC_us31_n690 ) );
NOR3_X2 _AES_ENC_us31_U171  ( .A1(_AES_ENC_us31_n695 ), .A2(_AES_ENC_us31_n694 ), .A3(_AES_ENC_us31_n693 ), .ZN(_AES_ENC_us31_n700 ) );
NOR4_X2 _AES_ENC_us31_U170  ( .A1(_AES_ENC_us31_n983 ), .A2(_AES_ENC_us31_n698 ), .A3(_AES_ENC_us31_n697 ), .A4(_AES_ENC_us31_n696 ), .ZN(_AES_ENC_us31_n699 ) );
NOR2_X2 _AES_ENC_us31_U169  ( .A1(_AES_ENC_us31_n946 ), .A2(_AES_ENC_us31_n945 ), .ZN(_AES_ENC_us31_n952 ) );
NOR4_X2 _AES_ENC_us31_U168  ( .A1(_AES_ENC_us31_n950 ), .A2(_AES_ENC_us31_n949 ), .A3(_AES_ENC_us31_n948 ), .A4(_AES_ENC_us31_n947 ), .ZN(_AES_ENC_us31_n951 ) );
NOR4_X2 _AES_ENC_us31_U162  ( .A1(_AES_ENC_us31_n896 ), .A2(_AES_ENC_us31_n895 ), .A3(_AES_ENC_us31_n894 ), .A4(_AES_ENC_us31_n893 ), .ZN(_AES_ENC_us31_n897 ) );
NOR2_X2 _AES_ENC_us31_U161  ( .A1(_AES_ENC_us31_n866 ), .A2(_AES_ENC_us31_n865 ), .ZN(_AES_ENC_us31_n872 ) );
NOR4_X2 _AES_ENC_us31_U160  ( .A1(_AES_ENC_us31_n870 ), .A2(_AES_ENC_us31_n869 ), .A3(_AES_ENC_us31_n868 ), .A4(_AES_ENC_us31_n867 ), .ZN(_AES_ENC_us31_n871 ) );
NOR4_X2 _AES_ENC_us31_U159  ( .A1(_AES_ENC_us31_n983 ), .A2(_AES_ENC_us31_n982 ), .A3(_AES_ENC_us31_n981 ), .A4(_AES_ENC_us31_n980 ), .ZN(_AES_ENC_us31_n984 ) );
NOR2_X2 _AES_ENC_us31_U158  ( .A1(_AES_ENC_us31_n979 ), .A2(_AES_ENC_us31_n978 ), .ZN(_AES_ENC_us31_n985 ) );
NOR4_X2 _AES_ENC_us31_U157  ( .A1(_AES_ENC_us31_n1125 ), .A2(_AES_ENC_us31_n1124 ), .A3(_AES_ENC_us31_n1123 ), .A4(_AES_ENC_us31_n1122 ), .ZN(_AES_ENC_us31_n1126 ) );
NOR4_X2 _AES_ENC_us31_U156  ( .A1(_AES_ENC_us31_n1084 ), .A2(_AES_ENC_us31_n1083 ), .A3(_AES_ENC_us31_n1082 ), .A4(_AES_ENC_us31_n1081 ), .ZN(_AES_ENC_us31_n1085 ) );
NOR2_X2 _AES_ENC_us31_U155  ( .A1(_AES_ENC_us31_n1076 ), .A2(_AES_ENC_us31_n1075 ), .ZN(_AES_ENC_us31_n1086 ) );
NOR3_X2 _AES_ENC_us31_U154  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n1054 ), .A3(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n961 ) );
NOR3_X2 _AES_ENC_us31_U153  ( .A1(_AES_ENC_us31_n620 ), .A2(_AES_ENC_us31_n1074 ), .A3(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n671 ) );
NOR2_X2 _AES_ENC_us31_U152  ( .A1(_AES_ENC_us31_n1057 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n1062 ) );
NOR2_X2 _AES_ENC_us31_U143  ( .A1(_AES_ENC_us31_n1055 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n1063 ) );
NOR2_X2 _AES_ENC_us31_U142  ( .A1(_AES_ENC_us31_n1060 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n1061 ) );
NOR4_X2 _AES_ENC_us31_U141  ( .A1(_AES_ENC_us31_n1064 ), .A2(_AES_ENC_us31_n1063 ), .A3(_AES_ENC_us31_n1062 ), .A4(_AES_ENC_us31_n1061 ), .ZN(_AES_ENC_us31_n1065 ) );
NOR3_X2 _AES_ENC_us31_U140  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n1120 ), .A3(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n918 ) );
NOR3_X2 _AES_ENC_us31_U132  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n573 ), .A3(_AES_ENC_us31_n1013 ), .ZN(_AES_ENC_us31_n917 ) );
NOR2_X2 _AES_ENC_us31_U131  ( .A1(_AES_ENC_us31_n914 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n915 ) );
NOR4_X2 _AES_ENC_us31_U130  ( .A1(_AES_ENC_us31_n918 ), .A2(_AES_ENC_us31_n917 ), .A3(_AES_ENC_us31_n916 ), .A4(_AES_ENC_us31_n915 ), .ZN(_AES_ENC_us31_n919 ) );
NOR2_X2 _AES_ENC_us31_U129  ( .A1(_AES_ENC_us31_n616 ), .A2(_AES_ENC_us31_n580 ), .ZN(_AES_ENC_us31_n771 ) );
NOR2_X2 _AES_ENC_us31_U128  ( .A1(_AES_ENC_us31_n1103 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n772 ) );
NOR2_X2 _AES_ENC_us31_U127  ( .A1(_AES_ENC_us31_n610 ), .A2(_AES_ENC_us31_n599 ), .ZN(_AES_ENC_us31_n773 ) );
NOR4_X2 _AES_ENC_us31_U126  ( .A1(_AES_ENC_us31_n773 ), .A2(_AES_ENC_us31_n772 ), .A3(_AES_ENC_us31_n771 ), .A4(_AES_ENC_us31_n770 ), .ZN(_AES_ENC_us31_n774 ) );
NOR2_X2 _AES_ENC_us31_U121  ( .A1(_AES_ENC_us31_n735 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n687 ) );
NOR2_X2 _AES_ENC_us31_U120  ( .A1(_AES_ENC_us31_n684 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n688 ) );
NOR2_X2 _AES_ENC_us31_U119  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n600 ), .ZN(_AES_ENC_us31_n686 ) );
NOR4_X2 _AES_ENC_us31_U118  ( .A1(_AES_ENC_us31_n688 ), .A2(_AES_ENC_us31_n687 ), .A3(_AES_ENC_us31_n686 ), .A4(_AES_ENC_us31_n685 ), .ZN(_AES_ENC_us31_n689 ) );
NOR2_X2 _AES_ENC_us31_U117  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n595 ), .ZN(_AES_ENC_us31_n858 ) );
NOR2_X2 _AES_ENC_us31_U116  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n855 ), .ZN(_AES_ENC_us31_n857 ) );
NOR2_X2 _AES_ENC_us31_U115  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n587 ), .ZN(_AES_ENC_us31_n856 ) );
NOR4_X2 _AES_ENC_us31_U106  ( .A1(_AES_ENC_us31_n858 ), .A2(_AES_ENC_us31_n857 ), .A3(_AES_ENC_us31_n856 ), .A4(_AES_ENC_us31_n958 ), .ZN(_AES_ENC_us31_n859 ) );
NOR2_X2 _AES_ENC_us31_U105  ( .A1(_AES_ENC_us31_n780 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n784 ) );
NOR2_X2 _AES_ENC_us31_U104  ( .A1(_AES_ENC_us31_n1117 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n782 ) );
NOR2_X2 _AES_ENC_us31_U103  ( .A1(_AES_ENC_us31_n781 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n783 ) );
NOR4_X2 _AES_ENC_us31_U102  ( .A1(_AES_ENC_us31_n880 ), .A2(_AES_ENC_us31_n784 ), .A3(_AES_ENC_us31_n783 ), .A4(_AES_ENC_us31_n782 ), .ZN(_AES_ENC_us31_n785 ) );
NOR2_X2 _AES_ENC_us31_U101  ( .A1(_AES_ENC_us31_n583 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n814 ) );
NOR2_X2 _AES_ENC_us31_U100  ( .A1(_AES_ENC_us31_n907 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n813 ) );
NOR3_X2 _AES_ENC_us31_U95  ( .A1(_AES_ENC_us31_n606 ), .A2(_AES_ENC_us31_n1058 ), .A3(_AES_ENC_us31_n1059 ), .ZN(_AES_ENC_us31_n815 ) );
NOR4_X2 _AES_ENC_us31_U94  ( .A1(_AES_ENC_us31_n815 ), .A2(_AES_ENC_us31_n814 ), .A3(_AES_ENC_us31_n813 ), .A4(_AES_ENC_us31_n812 ), .ZN(_AES_ENC_us31_n816 ) );
NOR2_X2 _AES_ENC_us31_U93  ( .A1(_AES_ENC_us31_n617 ), .A2(_AES_ENC_us31_n569 ), .ZN(_AES_ENC_us31_n721 ) );
NOR2_X2 _AES_ENC_us31_U92  ( .A1(_AES_ENC_us31_n1031 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n723 ) );
NOR2_X2 _AES_ENC_us31_U91  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n1096 ), .ZN(_AES_ENC_us31_n722 ) );
NOR4_X2 _AES_ENC_us31_U90  ( .A1(_AES_ENC_us31_n724 ), .A2(_AES_ENC_us31_n723 ), .A3(_AES_ENC_us31_n722 ), .A4(_AES_ENC_us31_n721 ), .ZN(_AES_ENC_us31_n725 ) );
NOR2_X2 _AES_ENC_us31_U89  ( .A1(_AES_ENC_us31_n911 ), .A2(_AES_ENC_us31_n990 ), .ZN(_AES_ENC_us31_n1009 ) );
NOR2_X2 _AES_ENC_us31_U88  ( .A1(_AES_ENC_us31_n1013 ), .A2(_AES_ENC_us31_n573 ), .ZN(_AES_ENC_us31_n1014 ) );
NOR2_X2 _AES_ENC_us31_U87  ( .A1(_AES_ENC_us31_n1014 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n1015 ) );
NOR4_X2 _AES_ENC_us31_U86  ( .A1(_AES_ENC_us31_n1016 ), .A2(_AES_ENC_us31_n1015 ), .A3(_AES_ENC_us31_n1119 ), .A4(_AES_ENC_us31_n1046 ), .ZN(_AES_ENC_us31_n1017 ) );
NOR2_X2 _AES_ENC_us31_U81  ( .A1(_AES_ENC_us31_n996 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n998 ) );
NOR2_X2 _AES_ENC_us31_U80  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n577 ), .ZN(_AES_ENC_us31_n1000 ) );
NOR2_X2 _AES_ENC_us31_U79  ( .A1(_AES_ENC_us31_n616 ), .A2(_AES_ENC_us31_n1096 ), .ZN(_AES_ENC_us31_n999 ) );
NOR4_X2 _AES_ENC_us31_U78  ( .A1(_AES_ENC_us31_n1000 ), .A2(_AES_ENC_us31_n999 ), .A3(_AES_ENC_us31_n998 ), .A4(_AES_ENC_us31_n997 ), .ZN(_AES_ENC_us31_n1001 ) );
NOR2_X2 _AES_ENC_us31_U74  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n1096 ), .ZN(_AES_ENC_us31_n697 ) );
NOR2_X2 _AES_ENC_us31_U73  ( .A1(_AES_ENC_us31_n620 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n958 ) );
NOR2_X2 _AES_ENC_us31_U72  ( .A1(_AES_ENC_us31_n911 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n983 ) );
NOR2_X2 _AES_ENC_us31_U71  ( .A1(_AES_ENC_us31_n1054 ), .A2(_AES_ENC_us31_n1103 ), .ZN(_AES_ENC_us31_n1031 ) );
INV_X4 _AES_ENC_us31_U65  ( .A(_AES_ENC_us31_n1050 ), .ZN(_AES_ENC_us31_n612 ) );
INV_X4 _AES_ENC_us31_U64  ( .A(_AES_ENC_us31_n1072 ), .ZN(_AES_ENC_us31_n605 ) );
INV_X4 _AES_ENC_us31_U63  ( .A(_AES_ENC_us31_n1073 ), .ZN(_AES_ENC_us31_n604 ) );
NOR2_X2 _AES_ENC_us31_U62  ( .A1(_AES_ENC_us31_n582 ), .A2(_AES_ENC_us31_n613 ), .ZN(_AES_ENC_us31_n880 ) );
NOR3_X2 _AES_ENC_us31_U61  ( .A1(_AES_ENC_us31_n826 ), .A2(_AES_ENC_us31_n1121 ), .A3(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n946 ) );
INV_X4 _AES_ENC_us31_U59  ( .A(_AES_ENC_us31_n1010 ), .ZN(_AES_ENC_us31_n608 ) );
NOR3_X2 _AES_ENC_us31_U58  ( .A1(_AES_ENC_us31_n573 ), .A2(_AES_ENC_us31_n1029 ), .A3(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n1119 ) );
INV_X4 _AES_ENC_us31_U57  ( .A(_AES_ENC_us31_n956 ), .ZN(_AES_ENC_us31_n615 ) );
NOR2_X2 _AES_ENC_us31_U50  ( .A1(_AES_ENC_us31_n623 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n1013 ) );
NOR2_X2 _AES_ENC_us31_U49  ( .A1(_AES_ENC_us31_n620 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n910 ) );
NOR2_X2 _AES_ENC_us31_U48  ( .A1(_AES_ENC_us31_n569 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n1091 ) );
NOR2_X2 _AES_ENC_us31_U47  ( .A1(_AES_ENC_us31_n622 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n990 ) );
NOR2_X2 _AES_ENC_us31_U46  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_us31_n1121 ), .ZN(_AES_ENC_us31_n996 ) );
NOR2_X2 _AES_ENC_us31_U45  ( .A1(_AES_ENC_us31_n610 ), .A2(_AES_ENC_us31_n600 ), .ZN(_AES_ENC_us31_n628 ) );
NOR2_X2 _AES_ENC_us31_U44  ( .A1(_AES_ENC_us31_n576 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n866 ) );
NOR2_X2 _AES_ENC_us31_U43  ( .A1(_AES_ENC_us31_n603 ), .A2(_AES_ENC_us31_n610 ), .ZN(_AES_ENC_us31_n1006 ) );
NOR2_X2 _AES_ENC_us31_U42  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n1117 ), .ZN(_AES_ENC_us31_n1118 ) );
NOR2_X2 _AES_ENC_us31_U41  ( .A1(_AES_ENC_us31_n1119 ), .A2(_AES_ENC_us31_n1118 ), .ZN(_AES_ENC_us31_n1127 ) );
NOR2_X2 _AES_ENC_us31_U36  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n594 ), .ZN(_AES_ENC_us31_n629 ) );
NOR2_X2 _AES_ENC_us31_U35  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n906 ), .ZN(_AES_ENC_us31_n909 ) );
NOR2_X2 _AES_ENC_us31_U34  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n597 ), .ZN(_AES_ENC_us31_n658 ) );
NOR2_X2 _AES_ENC_us31_U33  ( .A1(_AES_ENC_us31_n1116 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n695 ) );
NOR2_X2 _AES_ENC_us31_U32  ( .A1(_AES_ENC_us31_n1078 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n1083 ) );
NOR2_X2 _AES_ENC_us31_U31  ( .A1(_AES_ENC_us31_n941 ), .A2(_AES_ENC_us31_n608 ), .ZN(_AES_ENC_us31_n724 ) );
NOR2_X2 _AES_ENC_us31_U30  ( .A1(_AES_ENC_us31_n598 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n1107 ) );
NOR2_X2 _AES_ENC_us31_U29  ( .A1(_AES_ENC_us31_n576 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n840 ) );
NOR2_X2 _AES_ENC_us31_U24  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n593 ), .ZN(_AES_ENC_us31_n633 ) );
NOR2_X2 _AES_ENC_us31_U23  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n1080 ), .ZN(_AES_ENC_us31_n1081 ) );
NOR2_X2 _AES_ENC_us31_U21  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n1045 ), .ZN(_AES_ENC_us31_n812 ) );
NOR2_X2 _AES_ENC_us31_U20  ( .A1(_AES_ENC_us31_n1009 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n960 ) );
NOR2_X2 _AES_ENC_us31_U19  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n601 ), .ZN(_AES_ENC_us31_n982 ) );
NOR2_X2 _AES_ENC_us31_U18  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n594 ), .ZN(_AES_ENC_us31_n757 ) );
NOR2_X2 _AES_ENC_us31_U17  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n590 ), .ZN(_AES_ENC_us31_n698 ) );
NOR2_X2 _AES_ENC_us31_U16  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n619 ), .ZN(_AES_ENC_us31_n708 ) );
NOR2_X2 _AES_ENC_us31_U15  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n582 ), .ZN(_AES_ENC_us31_n770 ) );
NOR2_X2 _AES_ENC_us31_U10  ( .A1(_AES_ENC_us31_n619 ), .A2(_AES_ENC_us31_n604 ), .ZN(_AES_ENC_us31_n803 ) );
NOR2_X2 _AES_ENC_us31_U9  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n881 ), .ZN(_AES_ENC_us31_n711 ) );
NOR2_X2 _AES_ENC_us31_U8  ( .A1(_AES_ENC_us31_n615 ), .A2(_AES_ENC_us31_n582 ), .ZN(_AES_ENC_us31_n867 ) );
NOR2_X2 _AES_ENC_us31_U7  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n599 ), .ZN(_AES_ENC_us31_n804 ) );
NOR2_X2 _AES_ENC_us31_U6  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n620 ), .ZN(_AES_ENC_us31_n1046 ) );
OR2_X4 _AES_ENC_us31_U5  ( .A1(_AES_ENC_us31_n624 ), .A2(_AES_ENC_sa31[1]),.ZN(_AES_ENC_us31_n570 ) );
OR2_X4 _AES_ENC_us31_U4  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_sa31[4]),.ZN(_AES_ENC_us31_n569 ) );
NAND2_X2 _AES_ENC_us31_U514  ( .A1(_AES_ENC_us31_n1121 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n1030 ) );
AND2_X2 _AES_ENC_us31_U513  ( .A1(_AES_ENC_us31_n597 ), .A2(_AES_ENC_us31_n1030 ), .ZN(_AES_ENC_us31_n1049 ) );
NAND2_X2 _AES_ENC_us31_U511  ( .A1(_AES_ENC_us31_n1049 ), .A2(_AES_ENC_us31_n794 ), .ZN(_AES_ENC_us31_n637 ) );
AND2_X2 _AES_ENC_us31_U493  ( .A1(_AES_ENC_us31_n779 ), .A2(_AES_ENC_us31_n996 ), .ZN(_AES_ENC_us31_n632 ) );
NAND4_X2 _AES_ENC_us31_U485  ( .A1(_AES_ENC_us31_n637 ), .A2(_AES_ENC_us31_n636 ), .A3(_AES_ENC_us31_n635 ), .A4(_AES_ENC_us31_n634 ), .ZN(_AES_ENC_us31_n638 ) );
NAND2_X2 _AES_ENC_us31_U484  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n638 ), .ZN(_AES_ENC_us31_n679 ) );
NAND2_X2 _AES_ENC_us31_U481  ( .A1(_AES_ENC_us31_n1094 ), .A2(_AES_ENC_us31_n591 ), .ZN(_AES_ENC_us31_n648 ) );
NAND2_X2 _AES_ENC_us31_U476  ( .A1(_AES_ENC_us31_n601 ), .A2(_AES_ENC_us31_n590 ), .ZN(_AES_ENC_us31_n762 ) );
NAND2_X2 _AES_ENC_us31_U475  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n762 ), .ZN(_AES_ENC_us31_n647 ) );
NAND4_X2 _AES_ENC_us31_U457  ( .A1(_AES_ENC_us31_n648 ), .A2(_AES_ENC_us31_n647 ), .A3(_AES_ENC_us31_n646 ), .A4(_AES_ENC_us31_n645 ), .ZN(_AES_ENC_us31_n649 ) );
NAND2_X2 _AES_ENC_us31_U456  ( .A1(_AES_ENC_sa31[0]), .A2(_AES_ENC_us31_n649 ), .ZN(_AES_ENC_us31_n665 ) );
NAND2_X2 _AES_ENC_us31_U454  ( .A1(_AES_ENC_us31_n596 ), .A2(_AES_ENC_us31_n623 ), .ZN(_AES_ENC_us31_n855 ) );
NAND2_X2 _AES_ENC_us31_U453  ( .A1(_AES_ENC_us31_n587 ), .A2(_AES_ENC_us31_n855 ), .ZN(_AES_ENC_us31_n821 ) );
NAND2_X2 _AES_ENC_us31_U452  ( .A1(_AES_ENC_us31_n1093 ), .A2(_AES_ENC_us31_n821 ), .ZN(_AES_ENC_us31_n662 ) );
NAND2_X2 _AES_ENC_us31_U451  ( .A1(_AES_ENC_us31_n619 ), .A2(_AES_ENC_us31_n589 ), .ZN(_AES_ENC_us31_n650 ) );
NAND2_X2 _AES_ENC_us31_U450  ( .A1(_AES_ENC_us31_n956 ), .A2(_AES_ENC_us31_n650 ), .ZN(_AES_ENC_us31_n661 ) );
NAND2_X2 _AES_ENC_us31_U449  ( .A1(_AES_ENC_us31_n626 ), .A2(_AES_ENC_us31_n627 ), .ZN(_AES_ENC_us31_n839 ) );
OR2_X2 _AES_ENC_us31_U446  ( .A1(_AES_ENC_us31_n839 ), .A2(_AES_ENC_us31_n932 ), .ZN(_AES_ENC_us31_n656 ) );
NAND2_X2 _AES_ENC_us31_U445  ( .A1(_AES_ENC_us31_n621 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n1096 ) );
NAND2_X2 _AES_ENC_us31_U444  ( .A1(_AES_ENC_us31_n1030 ), .A2(_AES_ENC_us31_n1096 ), .ZN(_AES_ENC_us31_n651 ) );
NAND2_X2 _AES_ENC_us31_U443  ( .A1(_AES_ENC_us31_n1114 ), .A2(_AES_ENC_us31_n651 ), .ZN(_AES_ENC_us31_n655 ) );
OR3_X2 _AES_ENC_us31_U440  ( .A1(_AES_ENC_us31_n1079 ), .A2(_AES_ENC_sa31[7]), .A3(_AES_ENC_us31_n626 ), .ZN(_AES_ENC_us31_n654 ));
NAND2_X2 _AES_ENC_us31_U439  ( .A1(_AES_ENC_us31_n593 ), .A2(_AES_ENC_us31_n601 ), .ZN(_AES_ENC_us31_n652 ) );
NAND4_X2 _AES_ENC_us31_U437  ( .A1(_AES_ENC_us31_n656 ), .A2(_AES_ENC_us31_n655 ), .A3(_AES_ENC_us31_n654 ), .A4(_AES_ENC_us31_n653 ), .ZN(_AES_ENC_us31_n657 ) );
NAND2_X2 _AES_ENC_us31_U436  ( .A1(_AES_ENC_sa31[2]), .A2(_AES_ENC_us31_n657 ), .ZN(_AES_ENC_us31_n660 ) );
NAND4_X2 _AES_ENC_us31_U432  ( .A1(_AES_ENC_us31_n662 ), .A2(_AES_ENC_us31_n661 ), .A3(_AES_ENC_us31_n660 ), .A4(_AES_ENC_us31_n659 ), .ZN(_AES_ENC_us31_n663 ) );
NAND2_X2 _AES_ENC_us31_U431  ( .A1(_AES_ENC_us31_n663 ), .A2(_AES_ENC_us31_n574 ), .ZN(_AES_ENC_us31_n664 ) );
NAND2_X2 _AES_ENC_us31_U430  ( .A1(_AES_ENC_us31_n665 ), .A2(_AES_ENC_us31_n664 ), .ZN(_AES_ENC_us31_n666 ) );
NAND2_X2 _AES_ENC_us31_U429  ( .A1(_AES_ENC_sa31[6]), .A2(_AES_ENC_us31_n666 ), .ZN(_AES_ENC_us31_n678 ) );
NAND2_X2 _AES_ENC_us31_U426  ( .A1(_AES_ENC_us31_n735 ), .A2(_AES_ENC_us31_n1093 ), .ZN(_AES_ENC_us31_n675 ) );
NAND2_X2 _AES_ENC_us31_U425  ( .A1(_AES_ENC_us31_n588 ), .A2(_AES_ENC_us31_n597 ), .ZN(_AES_ENC_us31_n1045 ) );
OR2_X2 _AES_ENC_us31_U424  ( .A1(_AES_ENC_us31_n1045 ), .A2(_AES_ENC_us31_n605 ), .ZN(_AES_ENC_us31_n674 ) );
NAND2_X2 _AES_ENC_us31_U423  ( .A1(_AES_ENC_sa31[1]), .A2(_AES_ENC_us31_n620 ), .ZN(_AES_ENC_us31_n667 ) );
NAND2_X2 _AES_ENC_us31_U422  ( .A1(_AES_ENC_us31_n619 ), .A2(_AES_ENC_us31_n667 ), .ZN(_AES_ENC_us31_n1071 ) );
NAND4_X2 _AES_ENC_us31_U412  ( .A1(_AES_ENC_us31_n675 ), .A2(_AES_ENC_us31_n674 ), .A3(_AES_ENC_us31_n673 ), .A4(_AES_ENC_us31_n672 ), .ZN(_AES_ENC_us31_n676 ) );
NAND2_X2 _AES_ENC_us31_U411  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n676 ), .ZN(_AES_ENC_us31_n677 ) );
NAND2_X2 _AES_ENC_us31_U408  ( .A1(_AES_ENC_us31_n800 ), .A2(_AES_ENC_us31_n1022 ), .ZN(_AES_ENC_us31_n680 ) );
NAND2_X2 _AES_ENC_us31_U407  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n680 ), .ZN(_AES_ENC_us31_n681 ) );
AND2_X2 _AES_ENC_us31_U402  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n684 ), .ZN(_AES_ENC_us31_n682 ) );
NAND4_X2 _AES_ENC_us31_U395  ( .A1(_AES_ENC_us31_n691 ), .A2(_AES_ENC_us31_n581 ), .A3(_AES_ENC_us31_n690 ), .A4(_AES_ENC_us31_n689 ), .ZN(_AES_ENC_us31_n692 ) );
NAND2_X2 _AES_ENC_us31_U394  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n692 ), .ZN(_AES_ENC_us31_n733 ) );
NAND2_X2 _AES_ENC_us31_U392  ( .A1(_AES_ENC_us31_n977 ), .A2(_AES_ENC_us31_n1050 ), .ZN(_AES_ENC_us31_n702 ) );
NAND2_X2 _AES_ENC_us31_U391  ( .A1(_AES_ENC_us31_n1093 ), .A2(_AES_ENC_us31_n1045 ), .ZN(_AES_ENC_us31_n701 ) );
NAND4_X2 _AES_ENC_us31_U381  ( .A1(_AES_ENC_us31_n702 ), .A2(_AES_ENC_us31_n701 ), .A3(_AES_ENC_us31_n700 ), .A4(_AES_ENC_us31_n699 ), .ZN(_AES_ENC_us31_n703 ) );
NAND2_X2 _AES_ENC_us31_U380  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n703 ), .ZN(_AES_ENC_us31_n732 ) );
AND2_X2 _AES_ENC_us31_U379  ( .A1(_AES_ENC_sa31[0]), .A2(_AES_ENC_sa31[6]),.ZN(_AES_ENC_us31_n1113 ) );
NAND2_X2 _AES_ENC_us31_U378  ( .A1(_AES_ENC_us31_n601 ), .A2(_AES_ENC_us31_n1030 ), .ZN(_AES_ENC_us31_n881 ) );
NAND2_X2 _AES_ENC_us31_U377  ( .A1(_AES_ENC_us31_n1093 ), .A2(_AES_ENC_us31_n881 ), .ZN(_AES_ENC_us31_n715 ) );
NAND2_X2 _AES_ENC_us31_U376  ( .A1(_AES_ENC_us31_n1010 ), .A2(_AES_ENC_us31_n600 ), .ZN(_AES_ENC_us31_n714 ) );
NAND2_X2 _AES_ENC_us31_U375  ( .A1(_AES_ENC_us31_n855 ), .A2(_AES_ENC_us31_n588 ), .ZN(_AES_ENC_us31_n1117 ) );
XNOR2_X2 _AES_ENC_us31_U371  ( .A(_AES_ENC_us31_n611 ), .B(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n824 ) );
NAND4_X2 _AES_ENC_us31_U362  ( .A1(_AES_ENC_us31_n715 ), .A2(_AES_ENC_us31_n714 ), .A3(_AES_ENC_us31_n713 ), .A4(_AES_ENC_us31_n712 ), .ZN(_AES_ENC_us31_n716 ) );
NAND2_X2 _AES_ENC_us31_U361  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n716 ), .ZN(_AES_ENC_us31_n731 ) );
AND2_X2 _AES_ENC_us31_U360  ( .A1(_AES_ENC_sa31[6]), .A2(_AES_ENC_us31_n574 ), .ZN(_AES_ENC_us31_n1131 ) );
NAND2_X2 _AES_ENC_us31_U359  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n717 ) );
NAND2_X2 _AES_ENC_us31_U358  ( .A1(_AES_ENC_us31_n1029 ), .A2(_AES_ENC_us31_n717 ), .ZN(_AES_ENC_us31_n728 ) );
NAND2_X2 _AES_ENC_us31_U357  ( .A1(_AES_ENC_sa31[1]), .A2(_AES_ENC_us31_n624 ), .ZN(_AES_ENC_us31_n1097 ) );
NAND2_X2 _AES_ENC_us31_U356  ( .A1(_AES_ENC_us31_n603 ), .A2(_AES_ENC_us31_n1097 ), .ZN(_AES_ENC_us31_n718 ) );
NAND2_X2 _AES_ENC_us31_U355  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n718 ), .ZN(_AES_ENC_us31_n727 ) );
NAND4_X2 _AES_ENC_us31_U344  ( .A1(_AES_ENC_us31_n728 ), .A2(_AES_ENC_us31_n727 ), .A3(_AES_ENC_us31_n726 ), .A4(_AES_ENC_us31_n725 ), .ZN(_AES_ENC_us31_n729 ) );
NAND2_X2 _AES_ENC_us31_U343  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n729 ), .ZN(_AES_ENC_us31_n730 ) );
NAND4_X2 _AES_ENC_us31_U342  ( .A1(_AES_ENC_us31_n733 ), .A2(_AES_ENC_us31_n732 ), .A3(_AES_ENC_us31_n731 ), .A4(_AES_ENC_us31_n730 ), .ZN(_AES_ENC_sa31_sub[1] ) );
NAND2_X2 _AES_ENC_us31_U341  ( .A1(_AES_ENC_sa31[7]), .A2(_AES_ENC_us31_n611 ), .ZN(_AES_ENC_us31_n734 ) );
NAND2_X2 _AES_ENC_us31_U340  ( .A1(_AES_ENC_us31_n734 ), .A2(_AES_ENC_us31_n607 ), .ZN(_AES_ENC_us31_n738 ) );
OR4_X2 _AES_ENC_us31_U339  ( .A1(_AES_ENC_us31_n738 ), .A2(_AES_ENC_us31_n626 ), .A3(_AES_ENC_us31_n826 ), .A4(_AES_ENC_us31_n1121 ), .ZN(_AES_ENC_us31_n746 ) );
NAND2_X2 _AES_ENC_us31_U337  ( .A1(_AES_ENC_us31_n1100 ), .A2(_AES_ENC_us31_n587 ), .ZN(_AES_ENC_us31_n992 ) );
OR2_X2 _AES_ENC_us31_U336  ( .A1(_AES_ENC_us31_n610 ), .A2(_AES_ENC_us31_n735 ), .ZN(_AES_ENC_us31_n737 ) );
NAND2_X2 _AES_ENC_us31_U334  ( .A1(_AES_ENC_us31_n619 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n753 ) );
NAND2_X2 _AES_ENC_us31_U333  ( .A1(_AES_ENC_us31_n582 ), .A2(_AES_ENC_us31_n753 ), .ZN(_AES_ENC_us31_n1080 ) );
NAND2_X2 _AES_ENC_us31_U332  ( .A1(_AES_ENC_us31_n1048 ), .A2(_AES_ENC_us31_n576 ), .ZN(_AES_ENC_us31_n736 ) );
NAND2_X2 _AES_ENC_us31_U331  ( .A1(_AES_ENC_us31_n737 ), .A2(_AES_ENC_us31_n736 ), .ZN(_AES_ENC_us31_n739 ) );
NAND2_X2 _AES_ENC_us31_U330  ( .A1(_AES_ENC_us31_n739 ), .A2(_AES_ENC_us31_n738 ), .ZN(_AES_ENC_us31_n745 ) );
NAND2_X2 _AES_ENC_us31_U326  ( .A1(_AES_ENC_us31_n1096 ), .A2(_AES_ENC_us31_n590 ), .ZN(_AES_ENC_us31_n906 ) );
NAND4_X2 _AES_ENC_us31_U323  ( .A1(_AES_ENC_us31_n746 ), .A2(_AES_ENC_us31_n992 ), .A3(_AES_ENC_us31_n745 ), .A4(_AES_ENC_us31_n744 ), .ZN(_AES_ENC_us31_n747 ) );
NAND2_X2 _AES_ENC_us31_U322  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n747 ), .ZN(_AES_ENC_us31_n793 ) );
NAND2_X2 _AES_ENC_us31_U321  ( .A1(_AES_ENC_us31_n584 ), .A2(_AES_ENC_us31_n855 ), .ZN(_AES_ENC_us31_n748 ) );
NAND2_X2 _AES_ENC_us31_U320  ( .A1(_AES_ENC_us31_n956 ), .A2(_AES_ENC_us31_n748 ), .ZN(_AES_ENC_us31_n760 ) );
NAND2_X2 _AES_ENC_us31_U313  ( .A1(_AES_ENC_us31_n590 ), .A2(_AES_ENC_us31_n753 ), .ZN(_AES_ENC_us31_n1023 ) );
NAND4_X2 _AES_ENC_us31_U308  ( .A1(_AES_ENC_us31_n760 ), .A2(_AES_ENC_us31_n992 ), .A3(_AES_ENC_us31_n759 ), .A4(_AES_ENC_us31_n758 ), .ZN(_AES_ENC_us31_n761 ) );
NAND2_X2 _AES_ENC_us31_U307  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n761 ), .ZN(_AES_ENC_us31_n792 ) );
NAND2_X2 _AES_ENC_us31_U306  ( .A1(_AES_ENC_us31_n584 ), .A2(_AES_ENC_us31_n603 ), .ZN(_AES_ENC_us31_n989 ) );
NAND2_X2 _AES_ENC_us31_U305  ( .A1(_AES_ENC_us31_n1050 ), .A2(_AES_ENC_us31_n989 ), .ZN(_AES_ENC_us31_n777 ) );
NAND2_X2 _AES_ENC_us31_U304  ( .A1(_AES_ENC_us31_n1093 ), .A2(_AES_ENC_us31_n762 ), .ZN(_AES_ENC_us31_n776 ) );
XNOR2_X2 _AES_ENC_us31_U301  ( .A(_AES_ENC_sa31[7]), .B(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n959 ) );
NAND4_X2 _AES_ENC_us31_U289  ( .A1(_AES_ENC_us31_n777 ), .A2(_AES_ENC_us31_n776 ), .A3(_AES_ENC_us31_n775 ), .A4(_AES_ENC_us31_n774 ), .ZN(_AES_ENC_us31_n778 ) );
NAND2_X2 _AES_ENC_us31_U288  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n778 ), .ZN(_AES_ENC_us31_n791 ) );
NAND2_X2 _AES_ENC_us31_U287  ( .A1(_AES_ENC_us31_n1056 ), .A2(_AES_ENC_us31_n1050 ), .ZN(_AES_ENC_us31_n788 ) );
NAND2_X2 _AES_ENC_us31_U286  ( .A1(_AES_ENC_us31_n1091 ), .A2(_AES_ENC_us31_n779 ), .ZN(_AES_ENC_us31_n787 ) );
NAND2_X2 _AES_ENC_us31_U285  ( .A1(_AES_ENC_us31_n956 ), .A2(_AES_ENC_sa31[1]), .ZN(_AES_ENC_us31_n786 ) );
NAND4_X2 _AES_ENC_us31_U278  ( .A1(_AES_ENC_us31_n788 ), .A2(_AES_ENC_us31_n787 ), .A3(_AES_ENC_us31_n786 ), .A4(_AES_ENC_us31_n785 ), .ZN(_AES_ENC_us31_n789 ) );
NAND2_X2 _AES_ENC_us31_U277  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n789 ), .ZN(_AES_ENC_us31_n790 ) );
NAND4_X2 _AES_ENC_us31_U276  ( .A1(_AES_ENC_us31_n793 ), .A2(_AES_ENC_us31_n792 ), .A3(_AES_ENC_us31_n791 ), .A4(_AES_ENC_us31_n790 ), .ZN(_AES_ENC_sa31_sub[2] ) );
NAND2_X2 _AES_ENC_us31_U275  ( .A1(_AES_ENC_us31_n1059 ), .A2(_AES_ENC_us31_n794 ), .ZN(_AES_ENC_us31_n810 ) );
NAND2_X2 _AES_ENC_us31_U274  ( .A1(_AES_ENC_us31_n1049 ), .A2(_AES_ENC_us31_n956 ), .ZN(_AES_ENC_us31_n809 ) );
OR2_X2 _AES_ENC_us31_U266  ( .A1(_AES_ENC_us31_n1096 ), .A2(_AES_ENC_us31_n606 ), .ZN(_AES_ENC_us31_n802 ) );
NAND2_X2 _AES_ENC_us31_U265  ( .A1(_AES_ENC_us31_n1053 ), .A2(_AES_ENC_us31_n800 ), .ZN(_AES_ENC_us31_n801 ) );
NAND2_X2 _AES_ENC_us31_U264  ( .A1(_AES_ENC_us31_n802 ), .A2(_AES_ENC_us31_n801 ), .ZN(_AES_ENC_us31_n805 ) );
NAND4_X2 _AES_ENC_us31_U261  ( .A1(_AES_ENC_us31_n810 ), .A2(_AES_ENC_us31_n809 ), .A3(_AES_ENC_us31_n808 ), .A4(_AES_ENC_us31_n807 ), .ZN(_AES_ENC_us31_n811 ) );
NAND2_X2 _AES_ENC_us31_U260  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n811 ), .ZN(_AES_ENC_us31_n852 ) );
OR2_X2 _AES_ENC_us31_U259  ( .A1(_AES_ENC_us31_n1023 ), .A2(_AES_ENC_us31_n617 ), .ZN(_AES_ENC_us31_n819 ) );
OR2_X2 _AES_ENC_us31_U257  ( .A1(_AES_ENC_us31_n570 ), .A2(_AES_ENC_us31_n930 ), .ZN(_AES_ENC_us31_n818 ) );
NAND2_X2 _AES_ENC_us31_U256  ( .A1(_AES_ENC_us31_n1013 ), .A2(_AES_ENC_us31_n1094 ), .ZN(_AES_ENC_us31_n817 ) );
NAND4_X2 _AES_ENC_us31_U249  ( .A1(_AES_ENC_us31_n819 ), .A2(_AES_ENC_us31_n818 ), .A3(_AES_ENC_us31_n817 ), .A4(_AES_ENC_us31_n816 ), .ZN(_AES_ENC_us31_n820 ) );
NAND2_X2 _AES_ENC_us31_U248  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n820 ), .ZN(_AES_ENC_us31_n851 ) );
NAND2_X2 _AES_ENC_us31_U247  ( .A1(_AES_ENC_us31_n956 ), .A2(_AES_ENC_us31_n1080 ), .ZN(_AES_ENC_us31_n835 ) );
NAND2_X2 _AES_ENC_us31_U246  ( .A1(_AES_ENC_us31_n570 ), .A2(_AES_ENC_us31_n1030 ), .ZN(_AES_ENC_us31_n1047 ) );
OR2_X2 _AES_ENC_us31_U245  ( .A1(_AES_ENC_us31_n1047 ), .A2(_AES_ENC_us31_n612 ), .ZN(_AES_ENC_us31_n834 ) );
NAND2_X2 _AES_ENC_us31_U244  ( .A1(_AES_ENC_us31_n1072 ), .A2(_AES_ENC_us31_n589 ), .ZN(_AES_ENC_us31_n833 ) );
NAND4_X2 _AES_ENC_us31_U233  ( .A1(_AES_ENC_us31_n835 ), .A2(_AES_ENC_us31_n834 ), .A3(_AES_ENC_us31_n833 ), .A4(_AES_ENC_us31_n832 ), .ZN(_AES_ENC_us31_n836 ) );
NAND2_X2 _AES_ENC_us31_U232  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n836 ), .ZN(_AES_ENC_us31_n850 ) );
NAND2_X2 _AES_ENC_us31_U231  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n623 ), .ZN(_AES_ENC_us31_n847 ) );
NAND2_X2 _AES_ENC_us31_U230  ( .A1(_AES_ENC_us31_n1050 ), .A2(_AES_ENC_us31_n1071 ), .ZN(_AES_ENC_us31_n846 ) );
OR2_X2 _AES_ENC_us31_U224  ( .A1(_AES_ENC_us31_n1053 ), .A2(_AES_ENC_us31_n911 ), .ZN(_AES_ENC_us31_n1077 ) );
NAND4_X2 _AES_ENC_us31_U220  ( .A1(_AES_ENC_us31_n847 ), .A2(_AES_ENC_us31_n846 ), .A3(_AES_ENC_us31_n845 ), .A4(_AES_ENC_us31_n844 ), .ZN(_AES_ENC_us31_n848 ) );
NAND2_X2 _AES_ENC_us31_U219  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n848 ), .ZN(_AES_ENC_us31_n849 ) );
NAND4_X2 _AES_ENC_us31_U218  ( .A1(_AES_ENC_us31_n852 ), .A2(_AES_ENC_us31_n851 ), .A3(_AES_ENC_us31_n850 ), .A4(_AES_ENC_us31_n849 ), .ZN(_AES_ENC_sa31_sub[3] ) );
NAND2_X2 _AES_ENC_us31_U216  ( .A1(_AES_ENC_us31_n1009 ), .A2(_AES_ENC_us31_n1072 ), .ZN(_AES_ENC_us31_n862 ) );
NAND2_X2 _AES_ENC_us31_U215  ( .A1(_AES_ENC_us31_n603 ), .A2(_AES_ENC_us31_n577 ), .ZN(_AES_ENC_us31_n853 ) );
NAND2_X2 _AES_ENC_us31_U214  ( .A1(_AES_ENC_us31_n1050 ), .A2(_AES_ENC_us31_n853 ), .ZN(_AES_ENC_us31_n861 ) );
NAND4_X2 _AES_ENC_us31_U206  ( .A1(_AES_ENC_us31_n862 ), .A2(_AES_ENC_us31_n861 ), .A3(_AES_ENC_us31_n860 ), .A4(_AES_ENC_us31_n859 ), .ZN(_AES_ENC_us31_n863 ) );
NAND2_X2 _AES_ENC_us31_U205  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n863 ), .ZN(_AES_ENC_us31_n905 ) );
NAND2_X2 _AES_ENC_us31_U204  ( .A1(_AES_ENC_us31_n1010 ), .A2(_AES_ENC_us31_n989 ), .ZN(_AES_ENC_us31_n874 ) );
NAND2_X2 _AES_ENC_us31_U203  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n610 ), .ZN(_AES_ENC_us31_n864 ) );
NAND2_X2 _AES_ENC_us31_U202  ( .A1(_AES_ENC_us31_n929 ), .A2(_AES_ENC_us31_n864 ), .ZN(_AES_ENC_us31_n873 ) );
NAND4_X2 _AES_ENC_us31_U193  ( .A1(_AES_ENC_us31_n874 ), .A2(_AES_ENC_us31_n873 ), .A3(_AES_ENC_us31_n872 ), .A4(_AES_ENC_us31_n871 ), .ZN(_AES_ENC_us31_n875 ) );
NAND2_X2 _AES_ENC_us31_U192  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n875 ), .ZN(_AES_ENC_us31_n904 ) );
NAND2_X2 _AES_ENC_us31_U191  ( .A1(_AES_ENC_us31_n583 ), .A2(_AES_ENC_us31_n1050 ), .ZN(_AES_ENC_us31_n889 ) );
NAND2_X2 _AES_ENC_us31_U190  ( .A1(_AES_ENC_us31_n1093 ), .A2(_AES_ENC_us31_n587 ), .ZN(_AES_ENC_us31_n876 ) );
NAND2_X2 _AES_ENC_us31_U189  ( .A1(_AES_ENC_us31_n604 ), .A2(_AES_ENC_us31_n876 ), .ZN(_AES_ENC_us31_n877 ) );
NAND2_X2 _AES_ENC_us31_U188  ( .A1(_AES_ENC_us31_n877 ), .A2(_AES_ENC_us31_n623 ), .ZN(_AES_ENC_us31_n888 ) );
NAND4_X2 _AES_ENC_us31_U179  ( .A1(_AES_ENC_us31_n889 ), .A2(_AES_ENC_us31_n888 ), .A3(_AES_ENC_us31_n887 ), .A4(_AES_ENC_us31_n886 ), .ZN(_AES_ENC_us31_n890 ) );
NAND2_X2 _AES_ENC_us31_U178  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n890 ), .ZN(_AES_ENC_us31_n903 ) );
OR2_X2 _AES_ENC_us31_U177  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n1059 ), .ZN(_AES_ENC_us31_n900 ) );
NAND2_X2 _AES_ENC_us31_U176  ( .A1(_AES_ENC_us31_n1073 ), .A2(_AES_ENC_us31_n1047 ), .ZN(_AES_ENC_us31_n899 ) );
NAND2_X2 _AES_ENC_us31_U175  ( .A1(_AES_ENC_us31_n1094 ), .A2(_AES_ENC_us31_n595 ), .ZN(_AES_ENC_us31_n898 ) );
NAND4_X2 _AES_ENC_us31_U167  ( .A1(_AES_ENC_us31_n900 ), .A2(_AES_ENC_us31_n899 ), .A3(_AES_ENC_us31_n898 ), .A4(_AES_ENC_us31_n897 ), .ZN(_AES_ENC_us31_n901 ) );
NAND2_X2 _AES_ENC_us31_U166  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n901 ), .ZN(_AES_ENC_us31_n902 ) );
NAND4_X2 _AES_ENC_us31_U165  ( .A1(_AES_ENC_us31_n905 ), .A2(_AES_ENC_us31_n904 ), .A3(_AES_ENC_us31_n903 ), .A4(_AES_ENC_us31_n902 ), .ZN(_AES_ENC_sa31_sub[4] ) );
NAND2_X2 _AES_ENC_us31_U164  ( .A1(_AES_ENC_us31_n1094 ), .A2(_AES_ENC_us31_n599 ), .ZN(_AES_ENC_us31_n922 ) );
NAND2_X2 _AES_ENC_us31_U163  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n989 ), .ZN(_AES_ENC_us31_n921 ) );
NAND4_X2 _AES_ENC_us31_U151  ( .A1(_AES_ENC_us31_n922 ), .A2(_AES_ENC_us31_n921 ), .A3(_AES_ENC_us31_n920 ), .A4(_AES_ENC_us31_n919 ), .ZN(_AES_ENC_us31_n923 ) );
NAND2_X2 _AES_ENC_us31_U150  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n923 ), .ZN(_AES_ENC_us31_n972 ) );
NAND2_X2 _AES_ENC_us31_U149  ( .A1(_AES_ENC_us31_n582 ), .A2(_AES_ENC_us31_n619 ), .ZN(_AES_ENC_us31_n924 ) );
NAND2_X2 _AES_ENC_us31_U148  ( .A1(_AES_ENC_us31_n1073 ), .A2(_AES_ENC_us31_n924 ), .ZN(_AES_ENC_us31_n939 ) );
NAND2_X2 _AES_ENC_us31_U147  ( .A1(_AES_ENC_us31_n926 ), .A2(_AES_ENC_us31_n925 ), .ZN(_AES_ENC_us31_n927 ) );
NAND2_X2 _AES_ENC_us31_U146  ( .A1(_AES_ENC_us31_n606 ), .A2(_AES_ENC_us31_n927 ), .ZN(_AES_ENC_us31_n928 ) );
NAND2_X2 _AES_ENC_us31_U145  ( .A1(_AES_ENC_us31_n928 ), .A2(_AES_ENC_us31_n1080 ), .ZN(_AES_ENC_us31_n938 ) );
OR2_X2 _AES_ENC_us31_U144  ( .A1(_AES_ENC_us31_n1117 ), .A2(_AES_ENC_us31_n615 ), .ZN(_AES_ENC_us31_n937 ) );
NAND4_X2 _AES_ENC_us31_U139  ( .A1(_AES_ENC_us31_n939 ), .A2(_AES_ENC_us31_n938 ), .A3(_AES_ENC_us31_n937 ), .A4(_AES_ENC_us31_n936 ), .ZN(_AES_ENC_us31_n940 ) );
NAND2_X2 _AES_ENC_us31_U138  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n940 ), .ZN(_AES_ENC_us31_n971 ) );
OR2_X2 _AES_ENC_us31_U137  ( .A1(_AES_ENC_us31_n605 ), .A2(_AES_ENC_us31_n941 ), .ZN(_AES_ENC_us31_n954 ) );
NAND2_X2 _AES_ENC_us31_U136  ( .A1(_AES_ENC_us31_n1096 ), .A2(_AES_ENC_us31_n577 ), .ZN(_AES_ENC_us31_n942 ) );
NAND2_X2 _AES_ENC_us31_U135  ( .A1(_AES_ENC_us31_n1048 ), .A2(_AES_ENC_us31_n942 ), .ZN(_AES_ENC_us31_n943 ) );
NAND2_X2 _AES_ENC_us31_U134  ( .A1(_AES_ENC_us31_n612 ), .A2(_AES_ENC_us31_n943 ), .ZN(_AES_ENC_us31_n944 ) );
NAND2_X2 _AES_ENC_us31_U133  ( .A1(_AES_ENC_us31_n944 ), .A2(_AES_ENC_us31_n580 ), .ZN(_AES_ENC_us31_n953 ) );
NAND4_X2 _AES_ENC_us31_U125  ( .A1(_AES_ENC_us31_n954 ), .A2(_AES_ENC_us31_n953 ), .A3(_AES_ENC_us31_n952 ), .A4(_AES_ENC_us31_n951 ), .ZN(_AES_ENC_us31_n955 ) );
NAND2_X2 _AES_ENC_us31_U124  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n955 ), .ZN(_AES_ENC_us31_n970 ) );
NAND2_X2 _AES_ENC_us31_U123  ( .A1(_AES_ENC_us31_n1094 ), .A2(_AES_ENC_us31_n1071 ), .ZN(_AES_ENC_us31_n967 ) );
NAND2_X2 _AES_ENC_us31_U122  ( .A1(_AES_ENC_us31_n956 ), .A2(_AES_ENC_us31_n1030 ), .ZN(_AES_ENC_us31_n966 ) );
NAND4_X2 _AES_ENC_us31_U114  ( .A1(_AES_ENC_us31_n967 ), .A2(_AES_ENC_us31_n966 ), .A3(_AES_ENC_us31_n965 ), .A4(_AES_ENC_us31_n964 ), .ZN(_AES_ENC_us31_n968 ) );
NAND2_X2 _AES_ENC_us31_U113  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n968 ), .ZN(_AES_ENC_us31_n969 ) );
NAND4_X2 _AES_ENC_us31_U112  ( .A1(_AES_ENC_us31_n972 ), .A2(_AES_ENC_us31_n971 ), .A3(_AES_ENC_us31_n970 ), .A4(_AES_ENC_us31_n969 ), .ZN(_AES_ENC_sa31_sub[5] ) );
NAND2_X2 _AES_ENC_us31_U111  ( .A1(_AES_ENC_us31_n570 ), .A2(_AES_ENC_us31_n1097 ), .ZN(_AES_ENC_us31_n973 ) );
NAND2_X2 _AES_ENC_us31_U110  ( .A1(_AES_ENC_us31_n1073 ), .A2(_AES_ENC_us31_n973 ), .ZN(_AES_ENC_us31_n987 ) );
NAND2_X2 _AES_ENC_us31_U109  ( .A1(_AES_ENC_us31_n974 ), .A2(_AES_ENC_us31_n1077 ), .ZN(_AES_ENC_us31_n975 ) );
NAND2_X2 _AES_ENC_us31_U108  ( .A1(_AES_ENC_us31_n613 ), .A2(_AES_ENC_us31_n975 ), .ZN(_AES_ENC_us31_n976 ) );
NAND2_X2 _AES_ENC_us31_U107  ( .A1(_AES_ENC_us31_n977 ), .A2(_AES_ENC_us31_n976 ), .ZN(_AES_ENC_us31_n986 ) );
NAND4_X2 _AES_ENC_us31_U99  ( .A1(_AES_ENC_us31_n987 ), .A2(_AES_ENC_us31_n986 ), .A3(_AES_ENC_us31_n985 ), .A4(_AES_ENC_us31_n984 ), .ZN(_AES_ENC_us31_n988 ) );
NAND2_X2 _AES_ENC_us31_U98  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n988 ), .ZN(_AES_ENC_us31_n1044 ) );
NAND2_X2 _AES_ENC_us31_U97  ( .A1(_AES_ENC_us31_n1073 ), .A2(_AES_ENC_us31_n989 ), .ZN(_AES_ENC_us31_n1004 ) );
NAND2_X2 _AES_ENC_us31_U96  ( .A1(_AES_ENC_us31_n1092 ), .A2(_AES_ENC_us31_n619 ), .ZN(_AES_ENC_us31_n1003 ) );
NAND4_X2 _AES_ENC_us31_U85  ( .A1(_AES_ENC_us31_n1004 ), .A2(_AES_ENC_us31_n1003 ), .A3(_AES_ENC_us31_n1002 ), .A4(_AES_ENC_us31_n1001 ), .ZN(_AES_ENC_us31_n1005 ) );
NAND2_X2 _AES_ENC_us31_U84  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n1005 ), .ZN(_AES_ENC_us31_n1043 ) );
NAND2_X2 _AES_ENC_us31_U83  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n596 ), .ZN(_AES_ENC_us31_n1020 ) );
NAND2_X2 _AES_ENC_us31_U82  ( .A1(_AES_ENC_us31_n1050 ), .A2(_AES_ENC_us31_n624 ), .ZN(_AES_ENC_us31_n1019 ) );
NAND2_X2 _AES_ENC_us31_U77  ( .A1(_AES_ENC_us31_n1059 ), .A2(_AES_ENC_us31_n1114 ), .ZN(_AES_ENC_us31_n1012 ) );
NAND2_X2 _AES_ENC_us31_U76  ( .A1(_AES_ENC_us31_n1010 ), .A2(_AES_ENC_us31_n592 ), .ZN(_AES_ENC_us31_n1011 ) );
NAND2_X2 _AES_ENC_us31_U75  ( .A1(_AES_ENC_us31_n1012 ), .A2(_AES_ENC_us31_n1011 ), .ZN(_AES_ENC_us31_n1016 ) );
NAND4_X2 _AES_ENC_us31_U70  ( .A1(_AES_ENC_us31_n1020 ), .A2(_AES_ENC_us31_n1019 ), .A3(_AES_ENC_us31_n1018 ), .A4(_AES_ENC_us31_n1017 ), .ZN(_AES_ENC_us31_n1021 ) );
NAND2_X2 _AES_ENC_us31_U69  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n1021 ), .ZN(_AES_ENC_us31_n1042 ) );
NAND2_X2 _AES_ENC_us31_U68  ( .A1(_AES_ENC_us31_n1022 ), .A2(_AES_ENC_us31_n1093 ), .ZN(_AES_ENC_us31_n1039 ) );
NAND2_X2 _AES_ENC_us31_U67  ( .A1(_AES_ENC_us31_n1050 ), .A2(_AES_ENC_us31_n1023 ), .ZN(_AES_ENC_us31_n1038 ) );
NAND2_X2 _AES_ENC_us31_U66  ( .A1(_AES_ENC_us31_n1024 ), .A2(_AES_ENC_us31_n1071 ), .ZN(_AES_ENC_us31_n1037 ) );
AND2_X2 _AES_ENC_us31_U60  ( .A1(_AES_ENC_us31_n1030 ), .A2(_AES_ENC_us31_n602 ), .ZN(_AES_ENC_us31_n1078 ) );
NAND4_X2 _AES_ENC_us31_U56  ( .A1(_AES_ENC_us31_n1039 ), .A2(_AES_ENC_us31_n1038 ), .A3(_AES_ENC_us31_n1037 ), .A4(_AES_ENC_us31_n1036 ), .ZN(_AES_ENC_us31_n1040 ) );
NAND2_X2 _AES_ENC_us31_U55  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n1040 ), .ZN(_AES_ENC_us31_n1041 ) );
NAND4_X2 _AES_ENC_us31_U54  ( .A1(_AES_ENC_us31_n1044 ), .A2(_AES_ENC_us31_n1043 ), .A3(_AES_ENC_us31_n1042 ), .A4(_AES_ENC_us31_n1041 ), .ZN(_AES_ENC_sa31_sub[6] ) );
NAND2_X2 _AES_ENC_us31_U53  ( .A1(_AES_ENC_us31_n1072 ), .A2(_AES_ENC_us31_n1045 ), .ZN(_AES_ENC_us31_n1068 ) );
NAND2_X2 _AES_ENC_us31_U52  ( .A1(_AES_ENC_us31_n1046 ), .A2(_AES_ENC_us31_n582 ), .ZN(_AES_ENC_us31_n1067 ) );
NAND2_X2 _AES_ENC_us31_U51  ( .A1(_AES_ENC_us31_n1094 ), .A2(_AES_ENC_us31_n1047 ), .ZN(_AES_ENC_us31_n1066 ) );
NAND4_X2 _AES_ENC_us31_U40  ( .A1(_AES_ENC_us31_n1068 ), .A2(_AES_ENC_us31_n1067 ), .A3(_AES_ENC_us31_n1066 ), .A4(_AES_ENC_us31_n1065 ), .ZN(_AES_ENC_us31_n1069 ) );
NAND2_X2 _AES_ENC_us31_U39  ( .A1(_AES_ENC_us31_n1070 ), .A2(_AES_ENC_us31_n1069 ), .ZN(_AES_ENC_us31_n1135 ) );
NAND2_X2 _AES_ENC_us31_U38  ( .A1(_AES_ENC_us31_n1072 ), .A2(_AES_ENC_us31_n1071 ), .ZN(_AES_ENC_us31_n1088 ) );
NAND2_X2 _AES_ENC_us31_U37  ( .A1(_AES_ENC_us31_n1073 ), .A2(_AES_ENC_us31_n595 ), .ZN(_AES_ENC_us31_n1087 ) );
NAND4_X2 _AES_ENC_us31_U28  ( .A1(_AES_ENC_us31_n1088 ), .A2(_AES_ENC_us31_n1087 ), .A3(_AES_ENC_us31_n1086 ), .A4(_AES_ENC_us31_n1085 ), .ZN(_AES_ENC_us31_n1089 ) );
NAND2_X2 _AES_ENC_us31_U27  ( .A1(_AES_ENC_us31_n1090 ), .A2(_AES_ENC_us31_n1089 ), .ZN(_AES_ENC_us31_n1134 ) );
NAND2_X2 _AES_ENC_us31_U26  ( .A1(_AES_ENC_us31_n1091 ), .A2(_AES_ENC_us31_n1093 ), .ZN(_AES_ENC_us31_n1111 ) );
NAND2_X2 _AES_ENC_us31_U25  ( .A1(_AES_ENC_us31_n1092 ), .A2(_AES_ENC_us31_n1120 ), .ZN(_AES_ENC_us31_n1110 ) );
AND2_X2 _AES_ENC_us31_U22  ( .A1(_AES_ENC_us31_n1097 ), .A2(_AES_ENC_us31_n1096 ), .ZN(_AES_ENC_us31_n1098 ) );
NAND4_X2 _AES_ENC_us31_U14  ( .A1(_AES_ENC_us31_n1111 ), .A2(_AES_ENC_us31_n1110 ), .A3(_AES_ENC_us31_n1109 ), .A4(_AES_ENC_us31_n1108 ), .ZN(_AES_ENC_us31_n1112 ) );
NAND2_X2 _AES_ENC_us31_U13  ( .A1(_AES_ENC_us31_n1113 ), .A2(_AES_ENC_us31_n1112 ), .ZN(_AES_ENC_us31_n1133 ) );
NAND2_X2 _AES_ENC_us31_U12  ( .A1(_AES_ENC_us31_n1115 ), .A2(_AES_ENC_us31_n1114 ), .ZN(_AES_ENC_us31_n1129 ) );
OR2_X2 _AES_ENC_us31_U11  ( .A1(_AES_ENC_us31_n608 ), .A2(_AES_ENC_us31_n1116 ), .ZN(_AES_ENC_us31_n1128 ) );
NAND4_X2 _AES_ENC_us31_U3  ( .A1(_AES_ENC_us31_n1129 ), .A2(_AES_ENC_us31_n1128 ), .A3(_AES_ENC_us31_n1127 ), .A4(_AES_ENC_us31_n1126 ), .ZN(_AES_ENC_us31_n1130 ) );
NAND2_X2 _AES_ENC_us31_U2  ( .A1(_AES_ENC_us31_n1131 ), .A2(_AES_ENC_us31_n1130 ), .ZN(_AES_ENC_us31_n1132 ) );
NAND4_X2 _AES_ENC_us31_U1  ( .A1(_AES_ENC_us31_n1135 ), .A2(_AES_ENC_us31_n1134 ), .A3(_AES_ENC_us31_n1133 ), .A4(_AES_ENC_us31_n1132 ), .ZN(_AES_ENC_sa31_sub[7] ) );
INV_X4 _AES_ENC_us32_U575  ( .A(_AES_ENC_sa32[7]), .ZN(_AES_ENC_us32_n627 ));
INV_X4 _AES_ENC_us32_U574  ( .A(_AES_ENC_us32_n1114 ), .ZN(_AES_ENC_us32_n625 ) );
INV_X4 _AES_ENC_us32_U573  ( .A(_AES_ENC_sa32[4]), .ZN(_AES_ENC_us32_n624 ));
INV_X4 _AES_ENC_us32_U572  ( .A(_AES_ENC_us32_n1025 ), .ZN(_AES_ENC_us32_n622 ) );
INV_X4 _AES_ENC_us32_U571  ( .A(_AES_ENC_us32_n1120 ), .ZN(_AES_ENC_us32_n620 ) );
INV_X4 _AES_ENC_us32_U570  ( .A(_AES_ENC_us32_n1121 ), .ZN(_AES_ENC_us32_n619 ) );
INV_X4 _AES_ENC_us32_U569  ( .A(_AES_ENC_us32_n1048 ), .ZN(_AES_ENC_us32_n618 ) );
INV_X4 _AES_ENC_us32_U568  ( .A(_AES_ENC_us32_n974 ), .ZN(_AES_ENC_us32_n616 ) );
INV_X4 _AES_ENC_us32_U567  ( .A(_AES_ENC_us32_n794 ), .ZN(_AES_ENC_us32_n614 ) );
INV_X4 _AES_ENC_us32_U566  ( .A(_AES_ENC_sa32[2]), .ZN(_AES_ENC_us32_n611 ));
INV_X4 _AES_ENC_us32_U565  ( .A(_AES_ENC_us32_n800 ), .ZN(_AES_ENC_us32_n610 ) );
INV_X4 _AES_ENC_us32_U564  ( .A(_AES_ENC_us32_n925 ), .ZN(_AES_ENC_us32_n609 ) );
INV_X4 _AES_ENC_us32_U563  ( .A(_AES_ENC_us32_n779 ), .ZN(_AES_ENC_us32_n607 ) );
INV_X4 _AES_ENC_us32_U562  ( .A(_AES_ENC_us32_n1022 ), .ZN(_AES_ENC_us32_n603 ) );
INV_X4 _AES_ENC_us32_U561  ( .A(_AES_ENC_us32_n1102 ), .ZN(_AES_ENC_us32_n602 ) );
INV_X4 _AES_ENC_us32_U560  ( .A(_AES_ENC_us32_n929 ), .ZN(_AES_ENC_us32_n601 ) );
INV_X4 _AES_ENC_us32_U559  ( .A(_AES_ENC_us32_n1056 ), .ZN(_AES_ENC_us32_n600 ) );
INV_X4 _AES_ENC_us32_U558  ( .A(_AES_ENC_us32_n1054 ), .ZN(_AES_ENC_us32_n599 ) );
INV_X4 _AES_ENC_us32_U557  ( .A(_AES_ENC_us32_n881 ), .ZN(_AES_ENC_us32_n598 ) );
INV_X4 _AES_ENC_us32_U556  ( .A(_AES_ENC_us32_n926 ), .ZN(_AES_ENC_us32_n597 ) );
INV_X4 _AES_ENC_us32_U555  ( .A(_AES_ENC_us32_n977 ), .ZN(_AES_ENC_us32_n595 ) );
INV_X4 _AES_ENC_us32_U554  ( .A(_AES_ENC_us32_n1031 ), .ZN(_AES_ENC_us32_n594 ) );
INV_X4 _AES_ENC_us32_U553  ( .A(_AES_ENC_us32_n1103 ), .ZN(_AES_ENC_us32_n593 ) );
INV_X4 _AES_ENC_us32_U552  ( .A(_AES_ENC_us32_n1009 ), .ZN(_AES_ENC_us32_n592 ) );
INV_X4 _AES_ENC_us32_U551  ( .A(_AES_ENC_us32_n990 ), .ZN(_AES_ENC_us32_n591 ) );
INV_X4 _AES_ENC_us32_U550  ( .A(_AES_ENC_us32_n1058 ), .ZN(_AES_ENC_us32_n590 ) );
INV_X4 _AES_ENC_us32_U549  ( .A(_AES_ENC_us32_n1074 ), .ZN(_AES_ENC_us32_n589 ) );
INV_X4 _AES_ENC_us32_U548  ( .A(_AES_ENC_us32_n1053 ), .ZN(_AES_ENC_us32_n588 ) );
INV_X4 _AES_ENC_us32_U547  ( .A(_AES_ENC_us32_n826 ), .ZN(_AES_ENC_us32_n587 ) );
INV_X4 _AES_ENC_us32_U546  ( .A(_AES_ENC_us32_n992 ), .ZN(_AES_ENC_us32_n586 ) );
INV_X4 _AES_ENC_us32_U545  ( .A(_AES_ENC_us32_n821 ), .ZN(_AES_ENC_us32_n585 ) );
INV_X4 _AES_ENC_us32_U544  ( .A(_AES_ENC_us32_n910 ), .ZN(_AES_ENC_us32_n584 ) );
INV_X4 _AES_ENC_us32_U543  ( .A(_AES_ENC_us32_n906 ), .ZN(_AES_ENC_us32_n583 ) );
INV_X4 _AES_ENC_us32_U542  ( .A(_AES_ENC_us32_n880 ), .ZN(_AES_ENC_us32_n581 ) );
INV_X4 _AES_ENC_us32_U541  ( .A(_AES_ENC_us32_n1013 ), .ZN(_AES_ENC_us32_n580 ) );
INV_X4 _AES_ENC_us32_U540  ( .A(_AES_ENC_us32_n1092 ), .ZN(_AES_ENC_us32_n579 ) );
INV_X4 _AES_ENC_us32_U539  ( .A(_AES_ENC_us32_n824 ), .ZN(_AES_ENC_us32_n578 ) );
INV_X4 _AES_ENC_us32_U538  ( .A(_AES_ENC_us32_n1091 ), .ZN(_AES_ENC_us32_n577 ) );
INV_X4 _AES_ENC_us32_U537  ( .A(_AES_ENC_us32_n1080 ), .ZN(_AES_ENC_us32_n576 ) );
INV_X4 _AES_ENC_us32_U536  ( .A(_AES_ENC_us32_n959 ), .ZN(_AES_ENC_us32_n575 ) );
INV_X4 _AES_ENC_us32_U535  ( .A(_AES_ENC_sa32[0]), .ZN(_AES_ENC_us32_n574 ));
NOR2_X2 _AES_ENC_us32_U534  ( .A1(_AES_ENC_sa32[0]), .A2(_AES_ENC_sa32[6]),.ZN(_AES_ENC_us32_n1090 ) );
NOR2_X2 _AES_ENC_us32_U533  ( .A1(_AES_ENC_us32_n574 ), .A2(_AES_ENC_sa32[6]), .ZN(_AES_ENC_us32_n1070 ) );
NOR2_X2 _AES_ENC_us32_U532  ( .A1(_AES_ENC_sa32[4]), .A2(_AES_ENC_sa32[3]),.ZN(_AES_ENC_us32_n1025 ) );
INV_X4 _AES_ENC_us32_U531  ( .A(_AES_ENC_us32_n569 ), .ZN(_AES_ENC_us32_n572 ) );
NOR2_X2 _AES_ENC_us32_U530  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n765 ) );
NOR2_X2 _AES_ENC_us32_U529  ( .A1(_AES_ENC_sa32[4]), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n764 ) );
NOR2_X2 _AES_ENC_us32_U528  ( .A1(_AES_ENC_us32_n765 ), .A2(_AES_ENC_us32_n764 ), .ZN(_AES_ENC_us32_n766 ) );
NOR2_X2 _AES_ENC_us32_U527  ( .A1(_AES_ENC_us32_n766 ), .A2(_AES_ENC_us32_n575 ), .ZN(_AES_ENC_us32_n767 ) );
INV_X4 _AES_ENC_us32_U526  ( .A(_AES_ENC_sa32[3]), .ZN(_AES_ENC_us32_n621 ));
NAND3_X2 _AES_ENC_us32_U525  ( .A1(_AES_ENC_us32_n652 ), .A2(_AES_ENC_us32_n626 ), .A3(_AES_ENC_sa32[7]), .ZN(_AES_ENC_us32_n653 ));
NOR2_X2 _AES_ENC_us32_U524  ( .A1(_AES_ENC_us32_n611 ), .A2(_AES_ENC_sa32[5]), .ZN(_AES_ENC_us32_n925 ) );
NOR2_X2 _AES_ENC_us32_U523  ( .A1(_AES_ENC_sa32[5]), .A2(_AES_ENC_sa32[2]),.ZN(_AES_ENC_us32_n974 ) );
INV_X4 _AES_ENC_us32_U522  ( .A(_AES_ENC_sa32[5]), .ZN(_AES_ENC_us32_n626 ));
NOR2_X2 _AES_ENC_us32_U521  ( .A1(_AES_ENC_us32_n611 ), .A2(_AES_ENC_sa32[7]), .ZN(_AES_ENC_us32_n779 ) );
NAND3_X2 _AES_ENC_us32_U520  ( .A1(_AES_ENC_us32_n679 ), .A2(_AES_ENC_us32_n678 ), .A3(_AES_ENC_us32_n677 ), .ZN(_AES_ENC_sa32_sub[0] ) );
NOR2_X2 _AES_ENC_us32_U519  ( .A1(_AES_ENC_us32_n626 ), .A2(_AES_ENC_sa32[2]), .ZN(_AES_ENC_us32_n1048 ) );
NOR3_X2 _AES_ENC_us32_U518  ( .A1(_AES_ENC_us32_n627 ), .A2(_AES_ENC_sa32[5]), .A3(_AES_ENC_us32_n704 ), .ZN(_AES_ENC_us32_n706 ));
NOR2_X2 _AES_ENC_us32_U517  ( .A1(_AES_ENC_us32_n1117 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n707 ) );
NOR2_X2 _AES_ENC_us32_U516  ( .A1(_AES_ENC_sa32[4]), .A2(_AES_ENC_us32_n579 ), .ZN(_AES_ENC_us32_n705 ) );
NOR3_X2 _AES_ENC_us32_U515  ( .A1(_AES_ENC_us32_n707 ), .A2(_AES_ENC_us32_n706 ), .A3(_AES_ENC_us32_n705 ), .ZN(_AES_ENC_us32_n713 ) );
NOR4_X2 _AES_ENC_us32_U512  ( .A1(_AES_ENC_us32_n633 ), .A2(_AES_ENC_us32_n632 ), .A3(_AES_ENC_us32_n631 ), .A4(_AES_ENC_us32_n630 ), .ZN(_AES_ENC_us32_n634 ) );
NOR2_X2 _AES_ENC_us32_U510  ( .A1(_AES_ENC_us32_n629 ), .A2(_AES_ENC_us32_n628 ), .ZN(_AES_ENC_us32_n635 ) );
NAND3_X2 _AES_ENC_us32_U509  ( .A1(_AES_ENC_sa32[2]), .A2(_AES_ENC_sa32[7]), .A3(_AES_ENC_us32_n1059 ), .ZN(_AES_ENC_us32_n636 ) );
NOR2_X2 _AES_ENC_us32_U508  ( .A1(_AES_ENC_sa32[7]), .A2(_AES_ENC_sa32[2]),.ZN(_AES_ENC_us32_n794 ) );
NOR2_X2 _AES_ENC_us32_U507  ( .A1(_AES_ENC_sa32[4]), .A2(_AES_ENC_sa32[1]),.ZN(_AES_ENC_us32_n1102 ) );
NOR2_X2 _AES_ENC_us32_U506  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_sa32[3]), .ZN(_AES_ENC_us32_n1053 ) );
NOR2_X2 _AES_ENC_us32_U505  ( .A1(_AES_ENC_us32_n607 ), .A2(_AES_ENC_sa32[5]), .ZN(_AES_ENC_us32_n1024 ) );
NOR2_X2 _AES_ENC_us32_U504  ( .A1(_AES_ENC_us32_n625 ), .A2(_AES_ENC_sa32[2]), .ZN(_AES_ENC_us32_n1093 ) );
NOR2_X2 _AES_ENC_us32_U503  ( .A1(_AES_ENC_us32_n614 ), .A2(_AES_ENC_sa32[5]), .ZN(_AES_ENC_us32_n1094 ) );
NOR2_X2 _AES_ENC_us32_U502  ( .A1(_AES_ENC_us32_n624 ), .A2(_AES_ENC_sa32[3]), .ZN(_AES_ENC_us32_n931 ) );
INV_X4 _AES_ENC_us32_U501  ( .A(_AES_ENC_us32_n570 ), .ZN(_AES_ENC_us32_n573 ) );
NOR2_X2 _AES_ENC_us32_U500  ( .A1(_AES_ENC_us32_n1053 ), .A2(_AES_ENC_us32_n1095 ), .ZN(_AES_ENC_us32_n639 ) );
NOR3_X2 _AES_ENC_us32_U499  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n573 ), .A3(_AES_ENC_us32_n1074 ), .ZN(_AES_ENC_us32_n641 ) );
NOR2_X2 _AES_ENC_us32_U498  ( .A1(_AES_ENC_us32_n639 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n640 ) );
NOR2_X2 _AES_ENC_us32_U497  ( .A1(_AES_ENC_us32_n641 ), .A2(_AES_ENC_us32_n640 ), .ZN(_AES_ENC_us32_n646 ) );
NOR3_X2 _AES_ENC_us32_U496  ( .A1(_AES_ENC_us32_n995 ), .A2(_AES_ENC_us32_n586 ), .A3(_AES_ENC_us32_n994 ), .ZN(_AES_ENC_us32_n1002 ) );
NOR2_X2 _AES_ENC_us32_U495  ( .A1(_AES_ENC_us32_n909 ), .A2(_AES_ENC_us32_n908 ), .ZN(_AES_ENC_us32_n920 ) );
NOR2_X2 _AES_ENC_us32_U494  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n823 ) );
NOR2_X2 _AES_ENC_us32_U492  ( .A1(_AES_ENC_us32_n624 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n822 ) );
NOR2_X2 _AES_ENC_us32_U491  ( .A1(_AES_ENC_us32_n823 ), .A2(_AES_ENC_us32_n822 ), .ZN(_AES_ENC_us32_n825 ) );
NOR2_X2 _AES_ENC_us32_U490  ( .A1(_AES_ENC_sa32[1]), .A2(_AES_ENC_us32_n623 ), .ZN(_AES_ENC_us32_n913 ) );
NOR2_X2 _AES_ENC_us32_U489  ( .A1(_AES_ENC_us32_n913 ), .A2(_AES_ENC_us32_n1091 ), .ZN(_AES_ENC_us32_n914 ) );
NOR2_X2 _AES_ENC_us32_U488  ( .A1(_AES_ENC_us32_n826 ), .A2(_AES_ENC_us32_n572 ), .ZN(_AES_ENC_us32_n827 ) );
NOR3_X2 _AES_ENC_us32_U487  ( .A1(_AES_ENC_us32_n769 ), .A2(_AES_ENC_us32_n768 ), .A3(_AES_ENC_us32_n767 ), .ZN(_AES_ENC_us32_n775 ) );
NOR2_X2 _AES_ENC_us32_U486  ( .A1(_AES_ENC_us32_n1056 ), .A2(_AES_ENC_us32_n1053 ), .ZN(_AES_ENC_us32_n749 ) );
NOR2_X2 _AES_ENC_us32_U483  ( .A1(_AES_ENC_us32_n749 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n752 ) );
INV_X4 _AES_ENC_us32_U482  ( .A(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n596 ));
NOR2_X2 _AES_ENC_us32_U480  ( .A1(_AES_ENC_us32_n1054 ), .A2(_AES_ENC_us32_n1053 ), .ZN(_AES_ENC_us32_n1055 ) );
OR2_X4 _AES_ENC_us32_U479  ( .A1(_AES_ENC_us32_n1094 ), .A2(_AES_ENC_us32_n1093 ), .ZN(_AES_ENC_us32_n571 ) );
AND2_X2 _AES_ENC_us32_U478  ( .A1(_AES_ENC_us32_n571 ), .A2(_AES_ENC_us32_n1095 ), .ZN(_AES_ENC_us32_n1101 ) );
NOR2_X2 _AES_ENC_us32_U477  ( .A1(_AES_ENC_us32_n1074 ), .A2(_AES_ENC_us32_n931 ), .ZN(_AES_ENC_us32_n796 ) );
NOR2_X2 _AES_ENC_us32_U474  ( .A1(_AES_ENC_us32_n796 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n797 ) );
NOR2_X2 _AES_ENC_us32_U473  ( .A1(_AES_ENC_us32_n932 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n933 ) );
NOR2_X2 _AES_ENC_us32_U472  ( .A1(_AES_ENC_us32_n929 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n935 ) );
NOR2_X2 _AES_ENC_us32_U471  ( .A1(_AES_ENC_us32_n931 ), .A2(_AES_ENC_us32_n930 ), .ZN(_AES_ENC_us32_n934 ) );
NOR3_X2 _AES_ENC_us32_U470  ( .A1(_AES_ENC_us32_n935 ), .A2(_AES_ENC_us32_n934 ), .A3(_AES_ENC_us32_n933 ), .ZN(_AES_ENC_us32_n936 ) );
NOR2_X2 _AES_ENC_us32_U469  ( .A1(_AES_ENC_us32_n624 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n1075 ) );
NOR2_X2 _AES_ENC_us32_U468  ( .A1(_AES_ENC_us32_n572 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n949 ) );
NOR2_X2 _AES_ENC_us32_U467  ( .A1(_AES_ENC_us32_n1049 ), .A2(_AES_ENC_us32_n618 ), .ZN(_AES_ENC_us32_n1051 ) );
NOR2_X2 _AES_ENC_us32_U466  ( .A1(_AES_ENC_us32_n1051 ), .A2(_AES_ENC_us32_n1050 ), .ZN(_AES_ENC_us32_n1052 ) );
NOR2_X2 _AES_ENC_us32_U465  ( .A1(_AES_ENC_us32_n1052 ), .A2(_AES_ENC_us32_n592 ), .ZN(_AES_ENC_us32_n1064 ) );
NOR2_X2 _AES_ENC_us32_U464  ( .A1(_AES_ENC_sa32[1]), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n631 ) );
NOR2_X2 _AES_ENC_us32_U463  ( .A1(_AES_ENC_us32_n1025 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n980 ) );
NOR2_X2 _AES_ENC_us32_U462  ( .A1(_AES_ENC_us32_n1073 ), .A2(_AES_ENC_us32_n1094 ), .ZN(_AES_ENC_us32_n795 ) );
NOR2_X2 _AES_ENC_us32_U461  ( .A1(_AES_ENC_us32_n795 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n799 ) );
NOR2_X2 _AES_ENC_us32_U460  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n981 ) );
NOR2_X2 _AES_ENC_us32_U459  ( .A1(_AES_ENC_us32_n1102 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n643 ) );
NOR2_X2 _AES_ENC_us32_U458  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n621 ), .ZN(_AES_ENC_us32_n642 ) );
NOR2_X2 _AES_ENC_us32_U455  ( .A1(_AES_ENC_us32_n911 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n644 ) );
NOR4_X2 _AES_ENC_us32_U448  ( .A1(_AES_ENC_us32_n644 ), .A2(_AES_ENC_us32_n643 ), .A3(_AES_ENC_us32_n804 ), .A4(_AES_ENC_us32_n642 ), .ZN(_AES_ENC_us32_n645 ) );
NOR2_X2 _AES_ENC_us32_U447  ( .A1(_AES_ENC_us32_n1102 ), .A2(_AES_ENC_us32_n910 ), .ZN(_AES_ENC_us32_n932 ) );
NOR2_X2 _AES_ENC_us32_U442  ( .A1(_AES_ENC_us32_n1102 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n755 ) );
NOR2_X2 _AES_ENC_us32_U441  ( .A1(_AES_ENC_us32_n931 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n743 ) );
NOR2_X2 _AES_ENC_us32_U438  ( .A1(_AES_ENC_us32_n1072 ), .A2(_AES_ENC_us32_n1094 ), .ZN(_AES_ENC_us32_n930 ) );
NOR2_X2 _AES_ENC_us32_U435  ( .A1(_AES_ENC_us32_n1074 ), .A2(_AES_ENC_us32_n1025 ), .ZN(_AES_ENC_us32_n891 ) );
NOR2_X2 _AES_ENC_us32_U434  ( .A1(_AES_ENC_us32_n891 ), .A2(_AES_ENC_us32_n609 ), .ZN(_AES_ENC_us32_n894 ) );
NOR3_X2 _AES_ENC_us32_U433  ( .A1(_AES_ENC_us32_n623 ), .A2(_AES_ENC_sa32[1]), .A3(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n683 ));
INV_X4 _AES_ENC_us32_U428  ( .A(_AES_ENC_us32_n931 ), .ZN(_AES_ENC_us32_n623 ) );
NOR2_X2 _AES_ENC_us32_U427  ( .A1(_AES_ENC_us32_n996 ), .A2(_AES_ENC_us32_n931 ), .ZN(_AES_ENC_us32_n704 ) );
NOR2_X2 _AES_ENC_us32_U421  ( .A1(_AES_ENC_us32_n931 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n685 ) );
NOR2_X2 _AES_ENC_us32_U420  ( .A1(_AES_ENC_us32_n1029 ), .A2(_AES_ENC_us32_n1025 ), .ZN(_AES_ENC_us32_n1079 ) );
NOR3_X2 _AES_ENC_us32_U419  ( .A1(_AES_ENC_us32_n589 ), .A2(_AES_ENC_us32_n1025 ), .A3(_AES_ENC_us32_n616 ), .ZN(_AES_ENC_us32_n945 ) );
NOR2_X2 _AES_ENC_us32_U418  ( .A1(_AES_ENC_us32_n626 ), .A2(_AES_ENC_us32_n611 ), .ZN(_AES_ENC_us32_n800 ) );
NOR3_X2 _AES_ENC_us32_U417  ( .A1(_AES_ENC_us32_n590 ), .A2(_AES_ENC_us32_n627 ), .A3(_AES_ENC_us32_n611 ), .ZN(_AES_ENC_us32_n798 ) );
NOR3_X2 _AES_ENC_us32_U416  ( .A1(_AES_ENC_us32_n610 ), .A2(_AES_ENC_us32_n572 ), .A3(_AES_ENC_us32_n575 ), .ZN(_AES_ENC_us32_n962 ) );
NOR3_X2 _AES_ENC_us32_U415  ( .A1(_AES_ENC_us32_n959 ), .A2(_AES_ENC_us32_n572 ), .A3(_AES_ENC_us32_n609 ), .ZN(_AES_ENC_us32_n768 ) );
NOR3_X2 _AES_ENC_us32_U414  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n572 ), .A3(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n694 ) );
NOR3_X2 _AES_ENC_us32_U413  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n572 ), .A3(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n895 ) );
NOR3_X2 _AES_ENC_us32_U410  ( .A1(_AES_ENC_us32_n1008 ), .A2(_AES_ENC_us32_n1007 ), .A3(_AES_ENC_us32_n1006 ), .ZN(_AES_ENC_us32_n1018 ) );
NOR4_X2 _AES_ENC_us32_U409  ( .A1(_AES_ENC_us32_n806 ), .A2(_AES_ENC_us32_n805 ), .A3(_AES_ENC_us32_n804 ), .A4(_AES_ENC_us32_n803 ), .ZN(_AES_ENC_us32_n807 ) );
NOR3_X2 _AES_ENC_us32_U406  ( .A1(_AES_ENC_us32_n799 ), .A2(_AES_ENC_us32_n798 ), .A3(_AES_ENC_us32_n797 ), .ZN(_AES_ENC_us32_n808 ) );
NOR4_X2 _AES_ENC_us32_U405  ( .A1(_AES_ENC_us32_n843 ), .A2(_AES_ENC_us32_n842 ), .A3(_AES_ENC_us32_n841 ), .A4(_AES_ENC_us32_n840 ), .ZN(_AES_ENC_us32_n844 ) );
NOR3_X2 _AES_ENC_us32_U404  ( .A1(_AES_ENC_us32_n1101 ), .A2(_AES_ENC_us32_n1100 ), .A3(_AES_ENC_us32_n1099 ), .ZN(_AES_ENC_us32_n1109 ) );
NOR4_X2 _AES_ENC_us32_U403  ( .A1(_AES_ENC_us32_n711 ), .A2(_AES_ENC_us32_n710 ), .A3(_AES_ENC_us32_n709 ), .A4(_AES_ENC_us32_n708 ), .ZN(_AES_ENC_us32_n712 ) );
NOR4_X2 _AES_ENC_us32_U401  ( .A1(_AES_ENC_us32_n963 ), .A2(_AES_ENC_us32_n962 ), .A3(_AES_ENC_us32_n961 ), .A4(_AES_ENC_us32_n960 ), .ZN(_AES_ENC_us32_n964 ) );
NOR2_X2 _AES_ENC_us32_U400  ( .A1(_AES_ENC_us32_n669 ), .A2(_AES_ENC_us32_n668 ), .ZN(_AES_ENC_us32_n673 ) );
NOR4_X2 _AES_ENC_us32_U399  ( .A1(_AES_ENC_us32_n946 ), .A2(_AES_ENC_us32_n1046 ), .A3(_AES_ENC_us32_n671 ), .A4(_AES_ENC_us32_n670 ), .ZN(_AES_ENC_us32_n672 ) );
NOR3_X2 _AES_ENC_us32_U398  ( .A1(_AES_ENC_us32_n743 ), .A2(_AES_ENC_us32_n742 ), .A3(_AES_ENC_us32_n741 ), .ZN(_AES_ENC_us32_n744 ) );
NOR2_X2 _AES_ENC_us32_U397  ( .A1(_AES_ENC_us32_n697 ), .A2(_AES_ENC_us32_n658 ), .ZN(_AES_ENC_us32_n659 ) );
NOR2_X2 _AES_ENC_us32_U396  ( .A1(_AES_ENC_us32_n1078 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n1033 ) );
NOR2_X2 _AES_ENC_us32_U393  ( .A1(_AES_ENC_us32_n1031 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n1032 ) );
NOR3_X2 _AES_ENC_us32_U390  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n1025 ), .A3(_AES_ENC_us32_n1074 ), .ZN(_AES_ENC_us32_n1035 ) );
NOR4_X2 _AES_ENC_us32_U389  ( .A1(_AES_ENC_us32_n1035 ), .A2(_AES_ENC_us32_n1034 ), .A3(_AES_ENC_us32_n1033 ), .A4(_AES_ENC_us32_n1032 ), .ZN(_AES_ENC_us32_n1036 ) );
NOR2_X2 _AES_ENC_us32_U388  ( .A1(_AES_ENC_us32_n598 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n885 ) );
NOR2_X2 _AES_ENC_us32_U387  ( .A1(_AES_ENC_us32_n623 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n882 ) );
NOR2_X2 _AES_ENC_us32_U386  ( .A1(_AES_ENC_us32_n1053 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n884 ) );
NOR4_X2 _AES_ENC_us32_U385  ( .A1(_AES_ENC_us32_n885 ), .A2(_AES_ENC_us32_n884 ), .A3(_AES_ENC_us32_n883 ), .A4(_AES_ENC_us32_n882 ), .ZN(_AES_ENC_us32_n886 ) );
NOR2_X2 _AES_ENC_us32_U384  ( .A1(_AES_ENC_us32_n825 ), .A2(_AES_ENC_us32_n578 ), .ZN(_AES_ENC_us32_n830 ) );
NOR2_X2 _AES_ENC_us32_U383  ( .A1(_AES_ENC_us32_n827 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n829 ) );
NOR2_X2 _AES_ENC_us32_U382  ( .A1(_AES_ENC_us32_n572 ), .A2(_AES_ENC_us32_n579 ), .ZN(_AES_ENC_us32_n828 ) );
NOR4_X2 _AES_ENC_us32_U374  ( .A1(_AES_ENC_us32_n831 ), .A2(_AES_ENC_us32_n830 ), .A3(_AES_ENC_us32_n829 ), .A4(_AES_ENC_us32_n828 ), .ZN(_AES_ENC_us32_n832 ) );
NOR2_X2 _AES_ENC_us32_U373  ( .A1(_AES_ENC_us32_n606 ), .A2(_AES_ENC_us32_n582 ), .ZN(_AES_ENC_us32_n1104 ) );
NOR2_X2 _AES_ENC_us32_U372  ( .A1(_AES_ENC_us32_n1102 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n1106 ) );
NOR2_X2 _AES_ENC_us32_U370  ( .A1(_AES_ENC_us32_n1103 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n1105 ) );
NOR4_X2 _AES_ENC_us32_U369  ( .A1(_AES_ENC_us32_n1107 ), .A2(_AES_ENC_us32_n1106 ), .A3(_AES_ENC_us32_n1105 ), .A4(_AES_ENC_us32_n1104 ), .ZN(_AES_ENC_us32_n1108 ) );
NOR3_X2 _AES_ENC_us32_U368  ( .A1(_AES_ENC_us32_n959 ), .A2(_AES_ENC_us32_n621 ), .A3(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n963 ) );
NOR2_X2 _AES_ENC_us32_U367  ( .A1(_AES_ENC_us32_n626 ), .A2(_AES_ENC_us32_n627 ), .ZN(_AES_ENC_us32_n1114 ) );
INV_X4 _AES_ENC_us32_U366  ( .A(_AES_ENC_us32_n1024 ), .ZN(_AES_ENC_us32_n606 ) );
NOR3_X2 _AES_ENC_us32_U365  ( .A1(_AES_ENC_us32_n910 ), .A2(_AES_ENC_us32_n1059 ), .A3(_AES_ENC_us32_n611 ), .ZN(_AES_ENC_us32_n1115 ) );
INV_X4 _AES_ENC_us32_U364  ( .A(_AES_ENC_us32_n1094 ), .ZN(_AES_ENC_us32_n613 ) );
NOR2_X2 _AES_ENC_us32_U363  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n931 ), .ZN(_AES_ENC_us32_n1100 ) );
INV_X4 _AES_ENC_us32_U354  ( .A(_AES_ENC_us32_n1093 ), .ZN(_AES_ENC_us32_n617 ) );
NOR2_X2 _AES_ENC_us32_U353  ( .A1(_AES_ENC_us32_n569 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n929 ) );
NOR2_X2 _AES_ENC_us32_U352  ( .A1(_AES_ENC_us32_n620 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n926 ) );
NOR2_X2 _AES_ENC_us32_U351  ( .A1(_AES_ENC_us32_n572 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n1095 ) );
NOR2_X2 _AES_ENC_us32_U350  ( .A1(_AES_ENC_us32_n609 ), .A2(_AES_ENC_us32_n627 ), .ZN(_AES_ENC_us32_n1010 ) );
NOR2_X2 _AES_ENC_us32_U349  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n1103 ) );
NOR2_X2 _AES_ENC_us32_U348  ( .A1(_AES_ENC_us32_n622 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n1059 ) );
NOR2_X2 _AES_ENC_us32_U347  ( .A1(_AES_ENC_sa32[1]), .A2(_AES_ENC_us32_n1120 ), .ZN(_AES_ENC_us32_n1022 ) );
NOR2_X2 _AES_ENC_us32_U346  ( .A1(_AES_ENC_us32_n619 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n911 ) );
NOR2_X2 _AES_ENC_us32_U345  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_us32_n1025 ), .ZN(_AES_ENC_us32_n826 ) );
NOR2_X2 _AES_ENC_us32_U338  ( .A1(_AES_ENC_us32_n626 ), .A2(_AES_ENC_us32_n607 ), .ZN(_AES_ENC_us32_n1072 ) );
NOR2_X2 _AES_ENC_us32_U335  ( .A1(_AES_ENC_us32_n627 ), .A2(_AES_ENC_us32_n616 ), .ZN(_AES_ENC_us32_n956 ) );
NOR2_X2 _AES_ENC_us32_U329  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_us32_n624 ), .ZN(_AES_ENC_us32_n1121 ) );
NOR2_X2 _AES_ENC_us32_U328  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_us32_n624 ), .ZN(_AES_ENC_us32_n1058 ) );
NOR2_X2 _AES_ENC_us32_U327  ( .A1(_AES_ENC_us32_n625 ), .A2(_AES_ENC_us32_n611 ), .ZN(_AES_ENC_us32_n1073 ) );
NOR2_X2 _AES_ENC_us32_U325  ( .A1(_AES_ENC_sa32[1]), .A2(_AES_ENC_us32_n1025 ), .ZN(_AES_ENC_us32_n1054 ) );
NOR2_X2 _AES_ENC_us32_U324  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_us32_n931 ), .ZN(_AES_ENC_us32_n1029 ) );
NOR2_X2 _AES_ENC_us32_U319  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n1056 ) );
NOR2_X2 _AES_ENC_us32_U318  ( .A1(_AES_ENC_us32_n614 ), .A2(_AES_ENC_us32_n626 ), .ZN(_AES_ENC_us32_n1050 ) );
NOR2_X2 _AES_ENC_us32_U317  ( .A1(_AES_ENC_us32_n1121 ), .A2(_AES_ENC_us32_n1025 ), .ZN(_AES_ENC_us32_n1120 ) );
NOR2_X2 _AES_ENC_us32_U316  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_us32_n572 ), .ZN(_AES_ENC_us32_n1074 ) );
NOR2_X2 _AES_ENC_us32_U315  ( .A1(_AES_ENC_us32_n1058 ), .A2(_AES_ENC_us32_n1054 ), .ZN(_AES_ENC_us32_n878 ) );
NOR2_X2 _AES_ENC_us32_U314  ( .A1(_AES_ENC_us32_n878 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n879 ) );
NOR2_X2 _AES_ENC_us32_U312  ( .A1(_AES_ENC_us32_n880 ), .A2(_AES_ENC_us32_n879 ), .ZN(_AES_ENC_us32_n887 ) );
NOR2_X2 _AES_ENC_us32_U311  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n588 ), .ZN(_AES_ENC_us32_n957 ) );
NOR2_X2 _AES_ENC_us32_U310  ( .A1(_AES_ENC_us32_n958 ), .A2(_AES_ENC_us32_n957 ), .ZN(_AES_ENC_us32_n965 ) );
NOR3_X2 _AES_ENC_us32_U309  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n1091 ), .A3(_AES_ENC_us32_n1022 ), .ZN(_AES_ENC_us32_n720 ) );
NOR3_X2 _AES_ENC_us32_U303  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n1054 ), .A3(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n719 ) );
NOR2_X2 _AES_ENC_us32_U302  ( .A1(_AES_ENC_us32_n720 ), .A2(_AES_ENC_us32_n719 ), .ZN(_AES_ENC_us32_n726 ) );
NOR2_X2 _AES_ENC_us32_U300  ( .A1(_AES_ENC_us32_n614 ), .A2(_AES_ENC_us32_n591 ), .ZN(_AES_ENC_us32_n865 ) );
NOR2_X2 _AES_ENC_us32_U299  ( .A1(_AES_ENC_us32_n1059 ), .A2(_AES_ENC_us32_n1058 ), .ZN(_AES_ENC_us32_n1060 ) );
NOR2_X2 _AES_ENC_us32_U298  ( .A1(_AES_ENC_us32_n1095 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n668 ) );
NOR2_X2 _AES_ENC_us32_U297  ( .A1(_AES_ENC_us32_n911 ), .A2(_AES_ENC_us32_n910 ), .ZN(_AES_ENC_us32_n912 ) );
NOR2_X2 _AES_ENC_us32_U296  ( .A1(_AES_ENC_us32_n912 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n916 ) );
NOR2_X2 _AES_ENC_us32_U295  ( .A1(_AES_ENC_us32_n826 ), .A2(_AES_ENC_us32_n573 ), .ZN(_AES_ENC_us32_n750 ) );
NOR2_X2 _AES_ENC_us32_U294  ( .A1(_AES_ENC_us32_n750 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n751 ) );
NOR2_X2 _AES_ENC_us32_U293  ( .A1(_AES_ENC_us32_n907 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n908 ) );
NOR2_X2 _AES_ENC_us32_U292  ( .A1(_AES_ENC_us32_n990 ), .A2(_AES_ENC_us32_n926 ), .ZN(_AES_ENC_us32_n780 ) );
NOR2_X2 _AES_ENC_us32_U291  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n584 ), .ZN(_AES_ENC_us32_n838 ) );
NOR2_X2 _AES_ENC_us32_U290  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n602 ), .ZN(_AES_ENC_us32_n837 ) );
NOR2_X2 _AES_ENC_us32_U284  ( .A1(_AES_ENC_us32_n838 ), .A2(_AES_ENC_us32_n837 ), .ZN(_AES_ENC_us32_n845 ) );
NOR2_X2 _AES_ENC_us32_U283  ( .A1(_AES_ENC_us32_n1022 ), .A2(_AES_ENC_us32_n1058 ), .ZN(_AES_ENC_us32_n740 ) );
NOR2_X2 _AES_ENC_us32_U282  ( .A1(_AES_ENC_us32_n740 ), .A2(_AES_ENC_us32_n616 ), .ZN(_AES_ENC_us32_n742 ) );
NOR2_X2 _AES_ENC_us32_U281  ( .A1(_AES_ENC_us32_n1098 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n1099 ) );
NOR2_X2 _AES_ENC_us32_U280  ( .A1(_AES_ENC_us32_n1120 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n993 ) );
NOR2_X2 _AES_ENC_us32_U279  ( .A1(_AES_ENC_us32_n993 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n994 ) );
NOR2_X2 _AES_ENC_us32_U273  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n620 ), .ZN(_AES_ENC_us32_n1026 ) );
NOR2_X2 _AES_ENC_us32_U272  ( .A1(_AES_ENC_us32_n573 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n1027 ) );
NOR2_X2 _AES_ENC_us32_U271  ( .A1(_AES_ENC_us32_n1027 ), .A2(_AES_ENC_us32_n1026 ), .ZN(_AES_ENC_us32_n1028 ) );
NOR2_X2 _AES_ENC_us32_U270  ( .A1(_AES_ENC_us32_n1029 ), .A2(_AES_ENC_us32_n1028 ), .ZN(_AES_ENC_us32_n1034 ) );
NOR4_X2 _AES_ENC_us32_U269  ( .A1(_AES_ENC_us32_n757 ), .A2(_AES_ENC_us32_n756 ), .A3(_AES_ENC_us32_n755 ), .A4(_AES_ENC_us32_n754 ), .ZN(_AES_ENC_us32_n758 ) );
NOR2_X2 _AES_ENC_us32_U268  ( .A1(_AES_ENC_us32_n752 ), .A2(_AES_ENC_us32_n751 ), .ZN(_AES_ENC_us32_n759 ) );
NOR2_X2 _AES_ENC_us32_U267  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n1071 ), .ZN(_AES_ENC_us32_n669 ) );
NOR2_X2 _AES_ENC_us32_U263  ( .A1(_AES_ENC_us32_n1056 ), .A2(_AES_ENC_us32_n990 ), .ZN(_AES_ENC_us32_n991 ) );
NOR2_X2 _AES_ENC_us32_U262  ( .A1(_AES_ENC_us32_n991 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n995 ) );
NOR2_X2 _AES_ENC_us32_U258  ( .A1(_AES_ENC_us32_n607 ), .A2(_AES_ENC_us32_n590 ), .ZN(_AES_ENC_us32_n1008 ) );
NOR2_X2 _AES_ENC_us32_U255  ( .A1(_AES_ENC_us32_n839 ), .A2(_AES_ENC_us32_n582 ), .ZN(_AES_ENC_us32_n693 ) );
NOR2_X2 _AES_ENC_us32_U254  ( .A1(_AES_ENC_us32_n606 ), .A2(_AES_ENC_us32_n906 ), .ZN(_AES_ENC_us32_n741 ) );
NOR2_X2 _AES_ENC_us32_U253  ( .A1(_AES_ENC_us32_n1054 ), .A2(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n763 ) );
NOR2_X2 _AES_ENC_us32_U252  ( .A1(_AES_ENC_us32_n763 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n769 ) );
NOR2_X2 _AES_ENC_us32_U251  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n577 ), .ZN(_AES_ENC_us32_n1007 ) );
NOR2_X2 _AES_ENC_us32_U250  ( .A1(_AES_ENC_us32_n609 ), .A2(_AES_ENC_us32_n580 ), .ZN(_AES_ENC_us32_n1123 ) );
NOR2_X2 _AES_ENC_us32_U243  ( .A1(_AES_ENC_us32_n609 ), .A2(_AES_ENC_us32_n590 ), .ZN(_AES_ENC_us32_n710 ) );
INV_X4 _AES_ENC_us32_U242  ( .A(_AES_ENC_us32_n1029 ), .ZN(_AES_ENC_us32_n582 ) );
NOR2_X2 _AES_ENC_us32_U241  ( .A1(_AES_ENC_us32_n616 ), .A2(_AES_ENC_us32_n597 ), .ZN(_AES_ENC_us32_n883 ) );
NOR2_X2 _AES_ENC_us32_U240  ( .A1(_AES_ENC_us32_n593 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n1125 ) );
NOR2_X2 _AES_ENC_us32_U239  ( .A1(_AES_ENC_us32_n990 ), .A2(_AES_ENC_us32_n929 ), .ZN(_AES_ENC_us32_n892 ) );
NOR2_X2 _AES_ENC_us32_U238  ( .A1(_AES_ENC_us32_n892 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n893 ) );
NOR2_X2 _AES_ENC_us32_U237  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n602 ), .ZN(_AES_ENC_us32_n950 ) );
NOR2_X2 _AES_ENC_us32_U236  ( .A1(_AES_ENC_us32_n1079 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n1082 ) );
NOR2_X2 _AES_ENC_us32_U235  ( .A1(_AES_ENC_us32_n910 ), .A2(_AES_ENC_us32_n1056 ), .ZN(_AES_ENC_us32_n941 ) );
NOR2_X2 _AES_ENC_us32_U234  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n1077 ), .ZN(_AES_ENC_us32_n841 ) );
NOR2_X2 _AES_ENC_us32_U229  ( .A1(_AES_ENC_us32_n623 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n630 ) );
NOR2_X2 _AES_ENC_us32_U228  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n602 ), .ZN(_AES_ENC_us32_n806 ) );
NOR2_X2 _AES_ENC_us32_U227  ( .A1(_AES_ENC_us32_n623 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n948 ) );
NOR2_X2 _AES_ENC_us32_U226  ( .A1(_AES_ENC_us32_n606 ), .A2(_AES_ENC_us32_n589 ), .ZN(_AES_ENC_us32_n997 ) );
NOR2_X2 _AES_ENC_us32_U225  ( .A1(_AES_ENC_us32_n1121 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n1122 ) );
NOR2_X2 _AES_ENC_us32_U223  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n1023 ), .ZN(_AES_ENC_us32_n756 ) );
NOR2_X2 _AES_ENC_us32_U222  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n602 ), .ZN(_AES_ENC_us32_n870 ) );
NOR2_X2 _AES_ENC_us32_U221  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n569 ), .ZN(_AES_ENC_us32_n947 ) );
NOR2_X2 _AES_ENC_us32_U217  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n1077 ), .ZN(_AES_ENC_us32_n1084 ) );
NOR2_X2 _AES_ENC_us32_U213  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n855 ), .ZN(_AES_ENC_us32_n709 ) );
NOR2_X2 _AES_ENC_us32_U212  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n589 ), .ZN(_AES_ENC_us32_n868 ) );
NOR2_X2 _AES_ENC_us32_U211  ( .A1(_AES_ENC_us32_n1120 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n1124 ) );
NOR2_X2 _AES_ENC_us32_U210  ( .A1(_AES_ENC_us32_n1120 ), .A2(_AES_ENC_us32_n839 ), .ZN(_AES_ENC_us32_n842 ) );
NOR2_X2 _AES_ENC_us32_U209  ( .A1(_AES_ENC_us32_n1120 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n696 ) );
NOR2_X2 _AES_ENC_us32_U208  ( .A1(_AES_ENC_us32_n1074 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n1076 ) );
NOR2_X2 _AES_ENC_us32_U207  ( .A1(_AES_ENC_us32_n1074 ), .A2(_AES_ENC_us32_n620 ), .ZN(_AES_ENC_us32_n781 ) );
NOR3_X2 _AES_ENC_us32_U201  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n1056 ), .A3(_AES_ENC_us32_n990 ), .ZN(_AES_ENC_us32_n979 ) );
NOR3_X2 _AES_ENC_us32_U200  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n1058 ), .A3(_AES_ENC_us32_n1059 ), .ZN(_AES_ENC_us32_n854 ) );
NOR2_X2 _AES_ENC_us32_U199  ( .A1(_AES_ENC_us32_n996 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n869 ) );
NOR2_X2 _AES_ENC_us32_U198  ( .A1(_AES_ENC_us32_n1056 ), .A2(_AES_ENC_us32_n1074 ), .ZN(_AES_ENC_us32_n1057 ) );
NOR3_X2 _AES_ENC_us32_U197  ( .A1(_AES_ENC_us32_n607 ), .A2(_AES_ENC_us32_n1120 ), .A3(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n978 ) );
NOR2_X2 _AES_ENC_us32_U196  ( .A1(_AES_ENC_us32_n996 ), .A2(_AES_ENC_us32_n911 ), .ZN(_AES_ENC_us32_n1116 ) );
NOR2_X2 _AES_ENC_us32_U195  ( .A1(_AES_ENC_us32_n1074 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n754 ) );
NOR2_X2 _AES_ENC_us32_U194  ( .A1(_AES_ENC_us32_n926 ), .A2(_AES_ENC_us32_n1103 ), .ZN(_AES_ENC_us32_n977 ) );
NOR2_X2 _AES_ENC_us32_U187  ( .A1(_AES_ENC_us32_n839 ), .A2(_AES_ENC_us32_n824 ), .ZN(_AES_ENC_us32_n1092 ) );
NOR2_X2 _AES_ENC_us32_U186  ( .A1(_AES_ENC_us32_n573 ), .A2(_AES_ENC_us32_n1074 ), .ZN(_AES_ENC_us32_n684 ) );
NOR2_X2 _AES_ENC_us32_U185  ( .A1(_AES_ENC_us32_n826 ), .A2(_AES_ENC_us32_n1059 ), .ZN(_AES_ENC_us32_n907 ) );
NOR3_X2 _AES_ENC_us32_U184  ( .A1(_AES_ENC_us32_n625 ), .A2(_AES_ENC_us32_n1115 ), .A3(_AES_ENC_us32_n585 ), .ZN(_AES_ENC_us32_n831 ) );
NOR3_X2 _AES_ENC_us32_U183  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n1056 ), .A3(_AES_ENC_us32_n990 ), .ZN(_AES_ENC_us32_n896 ) );
NOR3_X2 _AES_ENC_us32_U182  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n573 ), .A3(_AES_ENC_us32_n1013 ), .ZN(_AES_ENC_us32_n670 ) );
NOR3_X2 _AES_ENC_us32_U181  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n1091 ), .A3(_AES_ENC_us32_n1022 ), .ZN(_AES_ENC_us32_n843 ) );
NOR2_X2 _AES_ENC_us32_U180  ( .A1(_AES_ENC_us32_n1029 ), .A2(_AES_ENC_us32_n1095 ), .ZN(_AES_ENC_us32_n735 ) );
NOR2_X2 _AES_ENC_us32_U174  ( .A1(_AES_ENC_us32_n1100 ), .A2(_AES_ENC_us32_n854 ), .ZN(_AES_ENC_us32_n860 ) );
NOR4_X2 _AES_ENC_us32_U173  ( .A1(_AES_ENC_us32_n1125 ), .A2(_AES_ENC_us32_n1124 ), .A3(_AES_ENC_us32_n1123 ), .A4(_AES_ENC_us32_n1122 ), .ZN(_AES_ENC_us32_n1126 ) );
NOR4_X2 _AES_ENC_us32_U172  ( .A1(_AES_ENC_us32_n1084 ), .A2(_AES_ENC_us32_n1083 ), .A3(_AES_ENC_us32_n1082 ), .A4(_AES_ENC_us32_n1081 ), .ZN(_AES_ENC_us32_n1085 ) );
NOR2_X2 _AES_ENC_us32_U171  ( .A1(_AES_ENC_us32_n1076 ), .A2(_AES_ENC_us32_n1075 ), .ZN(_AES_ENC_us32_n1086 ) );
NAND3_X2 _AES_ENC_us32_U170  ( .A1(_AES_ENC_us32_n569 ), .A2(_AES_ENC_us32_n582 ), .A3(_AES_ENC_us32_n681 ), .ZN(_AES_ENC_us32_n691 ) );
NOR2_X2 _AES_ENC_us32_U169  ( .A1(_AES_ENC_us32_n683 ), .A2(_AES_ENC_us32_n682 ), .ZN(_AES_ENC_us32_n690 ) );
NOR3_X2 _AES_ENC_us32_U168  ( .A1(_AES_ENC_us32_n695 ), .A2(_AES_ENC_us32_n694 ), .A3(_AES_ENC_us32_n693 ), .ZN(_AES_ENC_us32_n700 ) );
NOR4_X2 _AES_ENC_us32_U162  ( .A1(_AES_ENC_us32_n983 ), .A2(_AES_ENC_us32_n698 ), .A3(_AES_ENC_us32_n697 ), .A4(_AES_ENC_us32_n696 ), .ZN(_AES_ENC_us32_n699 ) );
NOR2_X2 _AES_ENC_us32_U161  ( .A1(_AES_ENC_us32_n946 ), .A2(_AES_ENC_us32_n945 ), .ZN(_AES_ENC_us32_n952 ) );
NOR4_X2 _AES_ENC_us32_U160  ( .A1(_AES_ENC_us32_n950 ), .A2(_AES_ENC_us32_n949 ), .A3(_AES_ENC_us32_n948 ), .A4(_AES_ENC_us32_n947 ), .ZN(_AES_ENC_us32_n951 ) );
NOR4_X2 _AES_ENC_us32_U159  ( .A1(_AES_ENC_us32_n896 ), .A2(_AES_ENC_us32_n895 ), .A3(_AES_ENC_us32_n894 ), .A4(_AES_ENC_us32_n893 ), .ZN(_AES_ENC_us32_n897 ) );
NOR2_X2 _AES_ENC_us32_U158  ( .A1(_AES_ENC_us32_n866 ), .A2(_AES_ENC_us32_n865 ), .ZN(_AES_ENC_us32_n872 ) );
NOR4_X2 _AES_ENC_us32_U157  ( .A1(_AES_ENC_us32_n870 ), .A2(_AES_ENC_us32_n869 ), .A3(_AES_ENC_us32_n868 ), .A4(_AES_ENC_us32_n867 ), .ZN(_AES_ENC_us32_n871 ) );
NOR4_X2 _AES_ENC_us32_U156  ( .A1(_AES_ENC_us32_n983 ), .A2(_AES_ENC_us32_n982 ), .A3(_AES_ENC_us32_n981 ), .A4(_AES_ENC_us32_n980 ), .ZN(_AES_ENC_us32_n984 ) );
NOR2_X2 _AES_ENC_us32_U155  ( .A1(_AES_ENC_us32_n979 ), .A2(_AES_ENC_us32_n978 ), .ZN(_AES_ENC_us32_n985 ) );
NOR3_X2 _AES_ENC_us32_U154  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n1054 ), .A3(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n961 ) );
NOR3_X2 _AES_ENC_us32_U153  ( .A1(_AES_ENC_us32_n620 ), .A2(_AES_ENC_us32_n1074 ), .A3(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n671 ) );
NOR2_X2 _AES_ENC_us32_U152  ( .A1(_AES_ENC_us32_n1057 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n1062 ) );
NOR2_X2 _AES_ENC_us32_U143  ( .A1(_AES_ENC_us32_n1055 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n1063 ) );
NOR2_X2 _AES_ENC_us32_U142  ( .A1(_AES_ENC_us32_n1060 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n1061 ) );
NOR4_X2 _AES_ENC_us32_U141  ( .A1(_AES_ENC_us32_n1064 ), .A2(_AES_ENC_us32_n1063 ), .A3(_AES_ENC_us32_n1062 ), .A4(_AES_ENC_us32_n1061 ), .ZN(_AES_ENC_us32_n1065 ) );
NOR3_X2 _AES_ENC_us32_U140  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n1120 ), .A3(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n918 ) );
NOR3_X2 _AES_ENC_us32_U132  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n573 ), .A3(_AES_ENC_us32_n1013 ), .ZN(_AES_ENC_us32_n917 ) );
NOR2_X2 _AES_ENC_us32_U131  ( .A1(_AES_ENC_us32_n914 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n915 ) );
NOR4_X2 _AES_ENC_us32_U130  ( .A1(_AES_ENC_us32_n918 ), .A2(_AES_ENC_us32_n917 ), .A3(_AES_ENC_us32_n916 ), .A4(_AES_ENC_us32_n915 ), .ZN(_AES_ENC_us32_n919 ) );
NOR2_X2 _AES_ENC_us32_U129  ( .A1(_AES_ENC_us32_n616 ), .A2(_AES_ENC_us32_n580 ), .ZN(_AES_ENC_us32_n771 ) );
NOR2_X2 _AES_ENC_us32_U128  ( .A1(_AES_ENC_us32_n1103 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n772 ) );
NOR2_X2 _AES_ENC_us32_U127  ( .A1(_AES_ENC_us32_n610 ), .A2(_AES_ENC_us32_n599 ), .ZN(_AES_ENC_us32_n773 ) );
NOR4_X2 _AES_ENC_us32_U126  ( .A1(_AES_ENC_us32_n773 ), .A2(_AES_ENC_us32_n772 ), .A3(_AES_ENC_us32_n771 ), .A4(_AES_ENC_us32_n770 ), .ZN(_AES_ENC_us32_n774 ) );
NOR2_X2 _AES_ENC_us32_U121  ( .A1(_AES_ENC_us32_n735 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n687 ) );
NOR2_X2 _AES_ENC_us32_U120  ( .A1(_AES_ENC_us32_n684 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n688 ) );
NOR2_X2 _AES_ENC_us32_U119  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n600 ), .ZN(_AES_ENC_us32_n686 ) );
NOR4_X2 _AES_ENC_us32_U118  ( .A1(_AES_ENC_us32_n688 ), .A2(_AES_ENC_us32_n687 ), .A3(_AES_ENC_us32_n686 ), .A4(_AES_ENC_us32_n685 ), .ZN(_AES_ENC_us32_n689 ) );
NOR2_X2 _AES_ENC_us32_U117  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n595 ), .ZN(_AES_ENC_us32_n858 ) );
NOR2_X2 _AES_ENC_us32_U116  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n855 ), .ZN(_AES_ENC_us32_n857 ) );
NOR2_X2 _AES_ENC_us32_U115  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n587 ), .ZN(_AES_ENC_us32_n856 ) );
NOR4_X2 _AES_ENC_us32_U106  ( .A1(_AES_ENC_us32_n858 ), .A2(_AES_ENC_us32_n857 ), .A3(_AES_ENC_us32_n856 ), .A4(_AES_ENC_us32_n958 ), .ZN(_AES_ENC_us32_n859 ) );
NOR2_X2 _AES_ENC_us32_U105  ( .A1(_AES_ENC_us32_n780 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n784 ) );
NOR2_X2 _AES_ENC_us32_U104  ( .A1(_AES_ENC_us32_n1117 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n782 ) );
NOR2_X2 _AES_ENC_us32_U103  ( .A1(_AES_ENC_us32_n781 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n783 ) );
NOR4_X2 _AES_ENC_us32_U102  ( .A1(_AES_ENC_us32_n880 ), .A2(_AES_ENC_us32_n784 ), .A3(_AES_ENC_us32_n783 ), .A4(_AES_ENC_us32_n782 ), .ZN(_AES_ENC_us32_n785 ) );
NOR2_X2 _AES_ENC_us32_U101  ( .A1(_AES_ENC_us32_n583 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n814 ) );
NOR2_X2 _AES_ENC_us32_U100  ( .A1(_AES_ENC_us32_n907 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n813 ) );
NOR3_X2 _AES_ENC_us32_U95  ( .A1(_AES_ENC_us32_n606 ), .A2(_AES_ENC_us32_n1058 ), .A3(_AES_ENC_us32_n1059 ), .ZN(_AES_ENC_us32_n815 ) );
NOR4_X2 _AES_ENC_us32_U94  ( .A1(_AES_ENC_us32_n815 ), .A2(_AES_ENC_us32_n814 ), .A3(_AES_ENC_us32_n813 ), .A4(_AES_ENC_us32_n812 ), .ZN(_AES_ENC_us32_n816 ) );
NOR2_X2 _AES_ENC_us32_U93  ( .A1(_AES_ENC_us32_n617 ), .A2(_AES_ENC_us32_n569 ), .ZN(_AES_ENC_us32_n721 ) );
NOR2_X2 _AES_ENC_us32_U92  ( .A1(_AES_ENC_us32_n1031 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n723 ) );
NOR2_X2 _AES_ENC_us32_U91  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n1096 ), .ZN(_AES_ENC_us32_n722 ) );
NOR4_X2 _AES_ENC_us32_U90  ( .A1(_AES_ENC_us32_n724 ), .A2(_AES_ENC_us32_n723 ), .A3(_AES_ENC_us32_n722 ), .A4(_AES_ENC_us32_n721 ), .ZN(_AES_ENC_us32_n725 ) );
NOR2_X2 _AES_ENC_us32_U89  ( .A1(_AES_ENC_us32_n911 ), .A2(_AES_ENC_us32_n990 ), .ZN(_AES_ENC_us32_n1009 ) );
NOR2_X2 _AES_ENC_us32_U88  ( .A1(_AES_ENC_us32_n1013 ), .A2(_AES_ENC_us32_n573 ), .ZN(_AES_ENC_us32_n1014 ) );
NOR2_X2 _AES_ENC_us32_U87  ( .A1(_AES_ENC_us32_n1014 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n1015 ) );
NOR4_X2 _AES_ENC_us32_U86  ( .A1(_AES_ENC_us32_n1016 ), .A2(_AES_ENC_us32_n1015 ), .A3(_AES_ENC_us32_n1119 ), .A4(_AES_ENC_us32_n1046 ), .ZN(_AES_ENC_us32_n1017 ) );
NOR2_X2 _AES_ENC_us32_U81  ( .A1(_AES_ENC_us32_n996 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n998 ) );
NOR2_X2 _AES_ENC_us32_U80  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n577 ), .ZN(_AES_ENC_us32_n1000 ) );
NOR2_X2 _AES_ENC_us32_U79  ( .A1(_AES_ENC_us32_n616 ), .A2(_AES_ENC_us32_n1096 ), .ZN(_AES_ENC_us32_n999 ) );
NOR4_X2 _AES_ENC_us32_U78  ( .A1(_AES_ENC_us32_n1000 ), .A2(_AES_ENC_us32_n999 ), .A3(_AES_ENC_us32_n998 ), .A4(_AES_ENC_us32_n997 ), .ZN(_AES_ENC_us32_n1001 ) );
NOR2_X2 _AES_ENC_us32_U74  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n1096 ), .ZN(_AES_ENC_us32_n697 ) );
NOR2_X2 _AES_ENC_us32_U73  ( .A1(_AES_ENC_us32_n620 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n958 ) );
NOR2_X2 _AES_ENC_us32_U72  ( .A1(_AES_ENC_us32_n911 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n983 ) );
NOR2_X2 _AES_ENC_us32_U71  ( .A1(_AES_ENC_us32_n1054 ), .A2(_AES_ENC_us32_n1103 ), .ZN(_AES_ENC_us32_n1031 ) );
INV_X4 _AES_ENC_us32_U65  ( .A(_AES_ENC_us32_n1050 ), .ZN(_AES_ENC_us32_n612 ) );
INV_X4 _AES_ENC_us32_U64  ( .A(_AES_ENC_us32_n1072 ), .ZN(_AES_ENC_us32_n605 ) );
INV_X4 _AES_ENC_us32_U63  ( .A(_AES_ENC_us32_n1073 ), .ZN(_AES_ENC_us32_n604 ) );
NOR2_X2 _AES_ENC_us32_U62  ( .A1(_AES_ENC_us32_n582 ), .A2(_AES_ENC_us32_n613 ), .ZN(_AES_ENC_us32_n880 ) );
NOR3_X2 _AES_ENC_us32_U61  ( .A1(_AES_ENC_us32_n826 ), .A2(_AES_ENC_us32_n1121 ), .A3(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n946 ) );
INV_X4 _AES_ENC_us32_U59  ( .A(_AES_ENC_us32_n1010 ), .ZN(_AES_ENC_us32_n608 ) );
NOR3_X2 _AES_ENC_us32_U58  ( .A1(_AES_ENC_us32_n573 ), .A2(_AES_ENC_us32_n1029 ), .A3(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n1119 ) );
INV_X4 _AES_ENC_us32_U57  ( .A(_AES_ENC_us32_n956 ), .ZN(_AES_ENC_us32_n615 ) );
NOR2_X2 _AES_ENC_us32_U50  ( .A1(_AES_ENC_us32_n623 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n1013 ) );
NOR2_X2 _AES_ENC_us32_U49  ( .A1(_AES_ENC_us32_n620 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n910 ) );
NOR2_X2 _AES_ENC_us32_U48  ( .A1(_AES_ENC_us32_n569 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n1091 ) );
NOR2_X2 _AES_ENC_us32_U47  ( .A1(_AES_ENC_us32_n622 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n990 ) );
NOR2_X2 _AES_ENC_us32_U46  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_us32_n1121 ), .ZN(_AES_ENC_us32_n996 ) );
NOR2_X2 _AES_ENC_us32_U45  ( .A1(_AES_ENC_us32_n610 ), .A2(_AES_ENC_us32_n600 ), .ZN(_AES_ENC_us32_n628 ) );
NOR2_X2 _AES_ENC_us32_U44  ( .A1(_AES_ENC_us32_n576 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n866 ) );
NOR2_X2 _AES_ENC_us32_U43  ( .A1(_AES_ENC_us32_n603 ), .A2(_AES_ENC_us32_n610 ), .ZN(_AES_ENC_us32_n1006 ) );
NOR2_X2 _AES_ENC_us32_U42  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n1117 ), .ZN(_AES_ENC_us32_n1118 ) );
NOR2_X2 _AES_ENC_us32_U41  ( .A1(_AES_ENC_us32_n1119 ), .A2(_AES_ENC_us32_n1118 ), .ZN(_AES_ENC_us32_n1127 ) );
NOR2_X2 _AES_ENC_us32_U36  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n906 ), .ZN(_AES_ENC_us32_n909 ) );
NOR2_X2 _AES_ENC_us32_U35  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n594 ), .ZN(_AES_ENC_us32_n629 ) );
NOR2_X2 _AES_ENC_us32_U34  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n597 ), .ZN(_AES_ENC_us32_n658 ) );
NOR2_X2 _AES_ENC_us32_U33  ( .A1(_AES_ENC_us32_n1116 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n695 ) );
NOR2_X2 _AES_ENC_us32_U32  ( .A1(_AES_ENC_us32_n1078 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n1083 ) );
NOR2_X2 _AES_ENC_us32_U31  ( .A1(_AES_ENC_us32_n941 ), .A2(_AES_ENC_us32_n608 ), .ZN(_AES_ENC_us32_n724 ) );
NOR2_X2 _AES_ENC_us32_U30  ( .A1(_AES_ENC_us32_n598 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n1107 ) );
NOR2_X2 _AES_ENC_us32_U29  ( .A1(_AES_ENC_us32_n576 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n840 ) );
NOR2_X2 _AES_ENC_us32_U24  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n593 ), .ZN(_AES_ENC_us32_n633 ) );
NOR2_X2 _AES_ENC_us32_U23  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n1080 ), .ZN(_AES_ENC_us32_n1081 ) );
NOR2_X2 _AES_ENC_us32_U21  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n1045 ), .ZN(_AES_ENC_us32_n812 ) );
NOR2_X2 _AES_ENC_us32_U20  ( .A1(_AES_ENC_us32_n1009 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n960 ) );
NOR2_X2 _AES_ENC_us32_U19  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n601 ), .ZN(_AES_ENC_us32_n982 ) );
NOR2_X2 _AES_ENC_us32_U18  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n594 ), .ZN(_AES_ENC_us32_n757 ) );
NOR2_X2 _AES_ENC_us32_U17  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n590 ), .ZN(_AES_ENC_us32_n698 ) );
NOR2_X2 _AES_ENC_us32_U16  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n619 ), .ZN(_AES_ENC_us32_n708 ) );
NOR2_X2 _AES_ENC_us32_U15  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n582 ), .ZN(_AES_ENC_us32_n770 ) );
NOR2_X2 _AES_ENC_us32_U10  ( .A1(_AES_ENC_us32_n619 ), .A2(_AES_ENC_us32_n604 ), .ZN(_AES_ENC_us32_n803 ) );
NOR2_X2 _AES_ENC_us32_U9  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n881 ), .ZN(_AES_ENC_us32_n711 ) );
NOR2_X2 _AES_ENC_us32_U8  ( .A1(_AES_ENC_us32_n615 ), .A2(_AES_ENC_us32_n582 ), .ZN(_AES_ENC_us32_n867 ) );
NOR2_X2 _AES_ENC_us32_U7  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n599 ), .ZN(_AES_ENC_us32_n804 ) );
NOR2_X2 _AES_ENC_us32_U6  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n620 ), .ZN(_AES_ENC_us32_n1046 ) );
OR2_X4 _AES_ENC_us32_U5  ( .A1(_AES_ENC_us32_n624 ), .A2(_AES_ENC_sa32[1]),.ZN(_AES_ENC_us32_n570 ) );
OR2_X4 _AES_ENC_us32_U4  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_sa32[4]),.ZN(_AES_ENC_us32_n569 ) );
NAND2_X2 _AES_ENC_us32_U514  ( .A1(_AES_ENC_us32_n1121 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n1030 ) );
AND2_X2 _AES_ENC_us32_U513  ( .A1(_AES_ENC_us32_n597 ), .A2(_AES_ENC_us32_n1030 ), .ZN(_AES_ENC_us32_n1049 ) );
NAND2_X2 _AES_ENC_us32_U511  ( .A1(_AES_ENC_us32_n1049 ), .A2(_AES_ENC_us32_n794 ), .ZN(_AES_ENC_us32_n637 ) );
AND2_X2 _AES_ENC_us32_U493  ( .A1(_AES_ENC_us32_n779 ), .A2(_AES_ENC_us32_n996 ), .ZN(_AES_ENC_us32_n632 ) );
NAND4_X2 _AES_ENC_us32_U485  ( .A1(_AES_ENC_us32_n637 ), .A2(_AES_ENC_us32_n636 ), .A3(_AES_ENC_us32_n635 ), .A4(_AES_ENC_us32_n634 ), .ZN(_AES_ENC_us32_n638 ) );
NAND2_X2 _AES_ENC_us32_U484  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n638 ), .ZN(_AES_ENC_us32_n679 ) );
NAND2_X2 _AES_ENC_us32_U481  ( .A1(_AES_ENC_us32_n1094 ), .A2(_AES_ENC_us32_n591 ), .ZN(_AES_ENC_us32_n648 ) );
NAND2_X2 _AES_ENC_us32_U476  ( .A1(_AES_ENC_us32_n601 ), .A2(_AES_ENC_us32_n590 ), .ZN(_AES_ENC_us32_n762 ) );
NAND2_X2 _AES_ENC_us32_U475  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n762 ), .ZN(_AES_ENC_us32_n647 ) );
NAND4_X2 _AES_ENC_us32_U457  ( .A1(_AES_ENC_us32_n648 ), .A2(_AES_ENC_us32_n647 ), .A3(_AES_ENC_us32_n646 ), .A4(_AES_ENC_us32_n645 ), .ZN(_AES_ENC_us32_n649 ) );
NAND2_X2 _AES_ENC_us32_U456  ( .A1(_AES_ENC_sa32[0]), .A2(_AES_ENC_us32_n649 ), .ZN(_AES_ENC_us32_n665 ) );
NAND2_X2 _AES_ENC_us32_U454  ( .A1(_AES_ENC_us32_n596 ), .A2(_AES_ENC_us32_n623 ), .ZN(_AES_ENC_us32_n855 ) );
NAND2_X2 _AES_ENC_us32_U453  ( .A1(_AES_ENC_us32_n587 ), .A2(_AES_ENC_us32_n855 ), .ZN(_AES_ENC_us32_n821 ) );
NAND2_X2 _AES_ENC_us32_U452  ( .A1(_AES_ENC_us32_n1093 ), .A2(_AES_ENC_us32_n821 ), .ZN(_AES_ENC_us32_n662 ) );
NAND2_X2 _AES_ENC_us32_U451  ( .A1(_AES_ENC_us32_n619 ), .A2(_AES_ENC_us32_n589 ), .ZN(_AES_ENC_us32_n650 ) );
NAND2_X2 _AES_ENC_us32_U450  ( .A1(_AES_ENC_us32_n956 ), .A2(_AES_ENC_us32_n650 ), .ZN(_AES_ENC_us32_n661 ) );
NAND2_X2 _AES_ENC_us32_U449  ( .A1(_AES_ENC_us32_n626 ), .A2(_AES_ENC_us32_n627 ), .ZN(_AES_ENC_us32_n839 ) );
OR2_X2 _AES_ENC_us32_U446  ( .A1(_AES_ENC_us32_n839 ), .A2(_AES_ENC_us32_n932 ), .ZN(_AES_ENC_us32_n656 ) );
NAND2_X2 _AES_ENC_us32_U445  ( .A1(_AES_ENC_us32_n621 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n1096 ) );
NAND2_X2 _AES_ENC_us32_U444  ( .A1(_AES_ENC_us32_n1030 ), .A2(_AES_ENC_us32_n1096 ), .ZN(_AES_ENC_us32_n651 ) );
NAND2_X2 _AES_ENC_us32_U443  ( .A1(_AES_ENC_us32_n1114 ), .A2(_AES_ENC_us32_n651 ), .ZN(_AES_ENC_us32_n655 ) );
OR3_X2 _AES_ENC_us32_U440  ( .A1(_AES_ENC_us32_n1079 ), .A2(_AES_ENC_sa32[7]), .A3(_AES_ENC_us32_n626 ), .ZN(_AES_ENC_us32_n654 ));
NAND2_X2 _AES_ENC_us32_U439  ( .A1(_AES_ENC_us32_n593 ), .A2(_AES_ENC_us32_n601 ), .ZN(_AES_ENC_us32_n652 ) );
NAND4_X2 _AES_ENC_us32_U437  ( .A1(_AES_ENC_us32_n656 ), .A2(_AES_ENC_us32_n655 ), .A3(_AES_ENC_us32_n654 ), .A4(_AES_ENC_us32_n653 ), .ZN(_AES_ENC_us32_n657 ) );
NAND2_X2 _AES_ENC_us32_U436  ( .A1(_AES_ENC_sa32[2]), .A2(_AES_ENC_us32_n657 ), .ZN(_AES_ENC_us32_n660 ) );
NAND4_X2 _AES_ENC_us32_U432  ( .A1(_AES_ENC_us32_n662 ), .A2(_AES_ENC_us32_n661 ), .A3(_AES_ENC_us32_n660 ), .A4(_AES_ENC_us32_n659 ), .ZN(_AES_ENC_us32_n663 ) );
NAND2_X2 _AES_ENC_us32_U431  ( .A1(_AES_ENC_us32_n663 ), .A2(_AES_ENC_us32_n574 ), .ZN(_AES_ENC_us32_n664 ) );
NAND2_X2 _AES_ENC_us32_U430  ( .A1(_AES_ENC_us32_n665 ), .A2(_AES_ENC_us32_n664 ), .ZN(_AES_ENC_us32_n666 ) );
NAND2_X2 _AES_ENC_us32_U429  ( .A1(_AES_ENC_sa32[6]), .A2(_AES_ENC_us32_n666 ), .ZN(_AES_ENC_us32_n678 ) );
NAND2_X2 _AES_ENC_us32_U426  ( .A1(_AES_ENC_us32_n735 ), .A2(_AES_ENC_us32_n1093 ), .ZN(_AES_ENC_us32_n675 ) );
NAND2_X2 _AES_ENC_us32_U425  ( .A1(_AES_ENC_us32_n588 ), .A2(_AES_ENC_us32_n597 ), .ZN(_AES_ENC_us32_n1045 ) );
OR2_X2 _AES_ENC_us32_U424  ( .A1(_AES_ENC_us32_n1045 ), .A2(_AES_ENC_us32_n605 ), .ZN(_AES_ENC_us32_n674 ) );
NAND2_X2 _AES_ENC_us32_U423  ( .A1(_AES_ENC_sa32[1]), .A2(_AES_ENC_us32_n620 ), .ZN(_AES_ENC_us32_n667 ) );
NAND2_X2 _AES_ENC_us32_U422  ( .A1(_AES_ENC_us32_n619 ), .A2(_AES_ENC_us32_n667 ), .ZN(_AES_ENC_us32_n1071 ) );
NAND4_X2 _AES_ENC_us32_U412  ( .A1(_AES_ENC_us32_n675 ), .A2(_AES_ENC_us32_n674 ), .A3(_AES_ENC_us32_n673 ), .A4(_AES_ENC_us32_n672 ), .ZN(_AES_ENC_us32_n676 ) );
NAND2_X2 _AES_ENC_us32_U411  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n676 ), .ZN(_AES_ENC_us32_n677 ) );
NAND2_X2 _AES_ENC_us32_U408  ( .A1(_AES_ENC_us32_n800 ), .A2(_AES_ENC_us32_n1022 ), .ZN(_AES_ENC_us32_n680 ) );
NAND2_X2 _AES_ENC_us32_U407  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n680 ), .ZN(_AES_ENC_us32_n681 ) );
AND2_X2 _AES_ENC_us32_U402  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n684 ), .ZN(_AES_ENC_us32_n682 ) );
NAND4_X2 _AES_ENC_us32_U395  ( .A1(_AES_ENC_us32_n691 ), .A2(_AES_ENC_us32_n581 ), .A3(_AES_ENC_us32_n690 ), .A4(_AES_ENC_us32_n689 ), .ZN(_AES_ENC_us32_n692 ) );
NAND2_X2 _AES_ENC_us32_U394  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n692 ), .ZN(_AES_ENC_us32_n733 ) );
NAND2_X2 _AES_ENC_us32_U392  ( .A1(_AES_ENC_us32_n977 ), .A2(_AES_ENC_us32_n1050 ), .ZN(_AES_ENC_us32_n702 ) );
NAND2_X2 _AES_ENC_us32_U391  ( .A1(_AES_ENC_us32_n1093 ), .A2(_AES_ENC_us32_n1045 ), .ZN(_AES_ENC_us32_n701 ) );
NAND4_X2 _AES_ENC_us32_U381  ( .A1(_AES_ENC_us32_n702 ), .A2(_AES_ENC_us32_n701 ), .A3(_AES_ENC_us32_n700 ), .A4(_AES_ENC_us32_n699 ), .ZN(_AES_ENC_us32_n703 ) );
NAND2_X2 _AES_ENC_us32_U380  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n703 ), .ZN(_AES_ENC_us32_n732 ) );
AND2_X2 _AES_ENC_us32_U379  ( .A1(_AES_ENC_sa32[0]), .A2(_AES_ENC_sa32[6]),.ZN(_AES_ENC_us32_n1113 ) );
NAND2_X2 _AES_ENC_us32_U378  ( .A1(_AES_ENC_us32_n601 ), .A2(_AES_ENC_us32_n1030 ), .ZN(_AES_ENC_us32_n881 ) );
NAND2_X2 _AES_ENC_us32_U377  ( .A1(_AES_ENC_us32_n1093 ), .A2(_AES_ENC_us32_n881 ), .ZN(_AES_ENC_us32_n715 ) );
NAND2_X2 _AES_ENC_us32_U376  ( .A1(_AES_ENC_us32_n1010 ), .A2(_AES_ENC_us32_n600 ), .ZN(_AES_ENC_us32_n714 ) );
NAND2_X2 _AES_ENC_us32_U375  ( .A1(_AES_ENC_us32_n855 ), .A2(_AES_ENC_us32_n588 ), .ZN(_AES_ENC_us32_n1117 ) );
XNOR2_X2 _AES_ENC_us32_U371  ( .A(_AES_ENC_us32_n611 ), .B(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n824 ) );
NAND4_X2 _AES_ENC_us32_U362  ( .A1(_AES_ENC_us32_n715 ), .A2(_AES_ENC_us32_n714 ), .A3(_AES_ENC_us32_n713 ), .A4(_AES_ENC_us32_n712 ), .ZN(_AES_ENC_us32_n716 ) );
NAND2_X2 _AES_ENC_us32_U361  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n716 ), .ZN(_AES_ENC_us32_n731 ) );
AND2_X2 _AES_ENC_us32_U360  ( .A1(_AES_ENC_sa32[6]), .A2(_AES_ENC_us32_n574 ), .ZN(_AES_ENC_us32_n1131 ) );
NAND2_X2 _AES_ENC_us32_U359  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n717 ) );
NAND2_X2 _AES_ENC_us32_U358  ( .A1(_AES_ENC_us32_n1029 ), .A2(_AES_ENC_us32_n717 ), .ZN(_AES_ENC_us32_n728 ) );
NAND2_X2 _AES_ENC_us32_U357  ( .A1(_AES_ENC_sa32[1]), .A2(_AES_ENC_us32_n624 ), .ZN(_AES_ENC_us32_n1097 ) );
NAND2_X2 _AES_ENC_us32_U356  ( .A1(_AES_ENC_us32_n603 ), .A2(_AES_ENC_us32_n1097 ), .ZN(_AES_ENC_us32_n718 ) );
NAND2_X2 _AES_ENC_us32_U355  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n718 ), .ZN(_AES_ENC_us32_n727 ) );
NAND4_X2 _AES_ENC_us32_U344  ( .A1(_AES_ENC_us32_n728 ), .A2(_AES_ENC_us32_n727 ), .A3(_AES_ENC_us32_n726 ), .A4(_AES_ENC_us32_n725 ), .ZN(_AES_ENC_us32_n729 ) );
NAND2_X2 _AES_ENC_us32_U343  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n729 ), .ZN(_AES_ENC_us32_n730 ) );
NAND4_X2 _AES_ENC_us32_U342  ( .A1(_AES_ENC_us32_n733 ), .A2(_AES_ENC_us32_n732 ), .A3(_AES_ENC_us32_n731 ), .A4(_AES_ENC_us32_n730 ), .ZN(_AES_ENC_sa32_sub[1] ) );
NAND2_X2 _AES_ENC_us32_U341  ( .A1(_AES_ENC_sa32[7]), .A2(_AES_ENC_us32_n611 ), .ZN(_AES_ENC_us32_n734 ) );
NAND2_X2 _AES_ENC_us32_U340  ( .A1(_AES_ENC_us32_n734 ), .A2(_AES_ENC_us32_n607 ), .ZN(_AES_ENC_us32_n738 ) );
OR4_X2 _AES_ENC_us32_U339  ( .A1(_AES_ENC_us32_n738 ), .A2(_AES_ENC_us32_n626 ), .A3(_AES_ENC_us32_n826 ), .A4(_AES_ENC_us32_n1121 ), .ZN(_AES_ENC_us32_n746 ) );
NAND2_X2 _AES_ENC_us32_U337  ( .A1(_AES_ENC_us32_n1100 ), .A2(_AES_ENC_us32_n587 ), .ZN(_AES_ENC_us32_n992 ) );
OR2_X2 _AES_ENC_us32_U336  ( .A1(_AES_ENC_us32_n610 ), .A2(_AES_ENC_us32_n735 ), .ZN(_AES_ENC_us32_n737 ) );
NAND2_X2 _AES_ENC_us32_U334  ( .A1(_AES_ENC_us32_n619 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n753 ) );
NAND2_X2 _AES_ENC_us32_U333  ( .A1(_AES_ENC_us32_n582 ), .A2(_AES_ENC_us32_n753 ), .ZN(_AES_ENC_us32_n1080 ) );
NAND2_X2 _AES_ENC_us32_U332  ( .A1(_AES_ENC_us32_n1048 ), .A2(_AES_ENC_us32_n576 ), .ZN(_AES_ENC_us32_n736 ) );
NAND2_X2 _AES_ENC_us32_U331  ( .A1(_AES_ENC_us32_n737 ), .A2(_AES_ENC_us32_n736 ), .ZN(_AES_ENC_us32_n739 ) );
NAND2_X2 _AES_ENC_us32_U330  ( .A1(_AES_ENC_us32_n739 ), .A2(_AES_ENC_us32_n738 ), .ZN(_AES_ENC_us32_n745 ) );
NAND2_X2 _AES_ENC_us32_U326  ( .A1(_AES_ENC_us32_n1096 ), .A2(_AES_ENC_us32_n590 ), .ZN(_AES_ENC_us32_n906 ) );
NAND4_X2 _AES_ENC_us32_U323  ( .A1(_AES_ENC_us32_n746 ), .A2(_AES_ENC_us32_n992 ), .A3(_AES_ENC_us32_n745 ), .A4(_AES_ENC_us32_n744 ), .ZN(_AES_ENC_us32_n747 ) );
NAND2_X2 _AES_ENC_us32_U322  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n747 ), .ZN(_AES_ENC_us32_n793 ) );
NAND2_X2 _AES_ENC_us32_U321  ( .A1(_AES_ENC_us32_n584 ), .A2(_AES_ENC_us32_n855 ), .ZN(_AES_ENC_us32_n748 ) );
NAND2_X2 _AES_ENC_us32_U320  ( .A1(_AES_ENC_us32_n956 ), .A2(_AES_ENC_us32_n748 ), .ZN(_AES_ENC_us32_n760 ) );
NAND2_X2 _AES_ENC_us32_U313  ( .A1(_AES_ENC_us32_n590 ), .A2(_AES_ENC_us32_n753 ), .ZN(_AES_ENC_us32_n1023 ) );
NAND4_X2 _AES_ENC_us32_U308  ( .A1(_AES_ENC_us32_n760 ), .A2(_AES_ENC_us32_n992 ), .A3(_AES_ENC_us32_n759 ), .A4(_AES_ENC_us32_n758 ), .ZN(_AES_ENC_us32_n761 ) );
NAND2_X2 _AES_ENC_us32_U307  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n761 ), .ZN(_AES_ENC_us32_n792 ) );
NAND2_X2 _AES_ENC_us32_U306  ( .A1(_AES_ENC_us32_n584 ), .A2(_AES_ENC_us32_n603 ), .ZN(_AES_ENC_us32_n989 ) );
NAND2_X2 _AES_ENC_us32_U305  ( .A1(_AES_ENC_us32_n1050 ), .A2(_AES_ENC_us32_n989 ), .ZN(_AES_ENC_us32_n777 ) );
NAND2_X2 _AES_ENC_us32_U304  ( .A1(_AES_ENC_us32_n1093 ), .A2(_AES_ENC_us32_n762 ), .ZN(_AES_ENC_us32_n776 ) );
XNOR2_X2 _AES_ENC_us32_U301  ( .A(_AES_ENC_sa32[7]), .B(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n959 ) );
NAND4_X2 _AES_ENC_us32_U289  ( .A1(_AES_ENC_us32_n777 ), .A2(_AES_ENC_us32_n776 ), .A3(_AES_ENC_us32_n775 ), .A4(_AES_ENC_us32_n774 ), .ZN(_AES_ENC_us32_n778 ) );
NAND2_X2 _AES_ENC_us32_U288  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n778 ), .ZN(_AES_ENC_us32_n791 ) );
NAND2_X2 _AES_ENC_us32_U287  ( .A1(_AES_ENC_us32_n1056 ), .A2(_AES_ENC_us32_n1050 ), .ZN(_AES_ENC_us32_n788 ) );
NAND2_X2 _AES_ENC_us32_U286  ( .A1(_AES_ENC_us32_n1091 ), .A2(_AES_ENC_us32_n779 ), .ZN(_AES_ENC_us32_n787 ) );
NAND2_X2 _AES_ENC_us32_U285  ( .A1(_AES_ENC_us32_n956 ), .A2(_AES_ENC_sa32[1]), .ZN(_AES_ENC_us32_n786 ) );
NAND4_X2 _AES_ENC_us32_U278  ( .A1(_AES_ENC_us32_n788 ), .A2(_AES_ENC_us32_n787 ), .A3(_AES_ENC_us32_n786 ), .A4(_AES_ENC_us32_n785 ), .ZN(_AES_ENC_us32_n789 ) );
NAND2_X2 _AES_ENC_us32_U277  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n789 ), .ZN(_AES_ENC_us32_n790 ) );
NAND4_X2 _AES_ENC_us32_U276  ( .A1(_AES_ENC_us32_n793 ), .A2(_AES_ENC_us32_n792 ), .A3(_AES_ENC_us32_n791 ), .A4(_AES_ENC_us32_n790 ), .ZN(_AES_ENC_sa32_sub[2] ) );
NAND2_X2 _AES_ENC_us32_U275  ( .A1(_AES_ENC_us32_n1059 ), .A2(_AES_ENC_us32_n794 ), .ZN(_AES_ENC_us32_n810 ) );
NAND2_X2 _AES_ENC_us32_U274  ( .A1(_AES_ENC_us32_n1049 ), .A2(_AES_ENC_us32_n956 ), .ZN(_AES_ENC_us32_n809 ) );
OR2_X2 _AES_ENC_us32_U266  ( .A1(_AES_ENC_us32_n1096 ), .A2(_AES_ENC_us32_n606 ), .ZN(_AES_ENC_us32_n802 ) );
NAND2_X2 _AES_ENC_us32_U265  ( .A1(_AES_ENC_us32_n1053 ), .A2(_AES_ENC_us32_n800 ), .ZN(_AES_ENC_us32_n801 ) );
NAND2_X2 _AES_ENC_us32_U264  ( .A1(_AES_ENC_us32_n802 ), .A2(_AES_ENC_us32_n801 ), .ZN(_AES_ENC_us32_n805 ) );
NAND4_X2 _AES_ENC_us32_U261  ( .A1(_AES_ENC_us32_n810 ), .A2(_AES_ENC_us32_n809 ), .A3(_AES_ENC_us32_n808 ), .A4(_AES_ENC_us32_n807 ), .ZN(_AES_ENC_us32_n811 ) );
NAND2_X2 _AES_ENC_us32_U260  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n811 ), .ZN(_AES_ENC_us32_n852 ) );
OR2_X2 _AES_ENC_us32_U259  ( .A1(_AES_ENC_us32_n1023 ), .A2(_AES_ENC_us32_n617 ), .ZN(_AES_ENC_us32_n819 ) );
OR2_X2 _AES_ENC_us32_U257  ( .A1(_AES_ENC_us32_n570 ), .A2(_AES_ENC_us32_n930 ), .ZN(_AES_ENC_us32_n818 ) );
NAND2_X2 _AES_ENC_us32_U256  ( .A1(_AES_ENC_us32_n1013 ), .A2(_AES_ENC_us32_n1094 ), .ZN(_AES_ENC_us32_n817 ) );
NAND4_X2 _AES_ENC_us32_U249  ( .A1(_AES_ENC_us32_n819 ), .A2(_AES_ENC_us32_n818 ), .A3(_AES_ENC_us32_n817 ), .A4(_AES_ENC_us32_n816 ), .ZN(_AES_ENC_us32_n820 ) );
NAND2_X2 _AES_ENC_us32_U248  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n820 ), .ZN(_AES_ENC_us32_n851 ) );
NAND2_X2 _AES_ENC_us32_U247  ( .A1(_AES_ENC_us32_n956 ), .A2(_AES_ENC_us32_n1080 ), .ZN(_AES_ENC_us32_n835 ) );
NAND2_X2 _AES_ENC_us32_U246  ( .A1(_AES_ENC_us32_n570 ), .A2(_AES_ENC_us32_n1030 ), .ZN(_AES_ENC_us32_n1047 ) );
OR2_X2 _AES_ENC_us32_U245  ( .A1(_AES_ENC_us32_n1047 ), .A2(_AES_ENC_us32_n612 ), .ZN(_AES_ENC_us32_n834 ) );
NAND2_X2 _AES_ENC_us32_U244  ( .A1(_AES_ENC_us32_n1072 ), .A2(_AES_ENC_us32_n589 ), .ZN(_AES_ENC_us32_n833 ) );
NAND4_X2 _AES_ENC_us32_U233  ( .A1(_AES_ENC_us32_n835 ), .A2(_AES_ENC_us32_n834 ), .A3(_AES_ENC_us32_n833 ), .A4(_AES_ENC_us32_n832 ), .ZN(_AES_ENC_us32_n836 ) );
NAND2_X2 _AES_ENC_us32_U232  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n836 ), .ZN(_AES_ENC_us32_n850 ) );
NAND2_X2 _AES_ENC_us32_U231  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n623 ), .ZN(_AES_ENC_us32_n847 ) );
NAND2_X2 _AES_ENC_us32_U230  ( .A1(_AES_ENC_us32_n1050 ), .A2(_AES_ENC_us32_n1071 ), .ZN(_AES_ENC_us32_n846 ) );
OR2_X2 _AES_ENC_us32_U224  ( .A1(_AES_ENC_us32_n1053 ), .A2(_AES_ENC_us32_n911 ), .ZN(_AES_ENC_us32_n1077 ) );
NAND4_X2 _AES_ENC_us32_U220  ( .A1(_AES_ENC_us32_n847 ), .A2(_AES_ENC_us32_n846 ), .A3(_AES_ENC_us32_n845 ), .A4(_AES_ENC_us32_n844 ), .ZN(_AES_ENC_us32_n848 ) );
NAND2_X2 _AES_ENC_us32_U219  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n848 ), .ZN(_AES_ENC_us32_n849 ) );
NAND4_X2 _AES_ENC_us32_U218  ( .A1(_AES_ENC_us32_n852 ), .A2(_AES_ENC_us32_n851 ), .A3(_AES_ENC_us32_n850 ), .A4(_AES_ENC_us32_n849 ), .ZN(_AES_ENC_sa32_sub[3] ) );
NAND2_X2 _AES_ENC_us32_U216  ( .A1(_AES_ENC_us32_n1009 ), .A2(_AES_ENC_us32_n1072 ), .ZN(_AES_ENC_us32_n862 ) );
NAND2_X2 _AES_ENC_us32_U215  ( .A1(_AES_ENC_us32_n603 ), .A2(_AES_ENC_us32_n577 ), .ZN(_AES_ENC_us32_n853 ) );
NAND2_X2 _AES_ENC_us32_U214  ( .A1(_AES_ENC_us32_n1050 ), .A2(_AES_ENC_us32_n853 ), .ZN(_AES_ENC_us32_n861 ) );
NAND4_X2 _AES_ENC_us32_U206  ( .A1(_AES_ENC_us32_n862 ), .A2(_AES_ENC_us32_n861 ), .A3(_AES_ENC_us32_n860 ), .A4(_AES_ENC_us32_n859 ), .ZN(_AES_ENC_us32_n863 ) );
NAND2_X2 _AES_ENC_us32_U205  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n863 ), .ZN(_AES_ENC_us32_n905 ) );
NAND2_X2 _AES_ENC_us32_U204  ( .A1(_AES_ENC_us32_n1010 ), .A2(_AES_ENC_us32_n989 ), .ZN(_AES_ENC_us32_n874 ) );
NAND2_X2 _AES_ENC_us32_U203  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n610 ), .ZN(_AES_ENC_us32_n864 ) );
NAND2_X2 _AES_ENC_us32_U202  ( .A1(_AES_ENC_us32_n929 ), .A2(_AES_ENC_us32_n864 ), .ZN(_AES_ENC_us32_n873 ) );
NAND4_X2 _AES_ENC_us32_U193  ( .A1(_AES_ENC_us32_n874 ), .A2(_AES_ENC_us32_n873 ), .A3(_AES_ENC_us32_n872 ), .A4(_AES_ENC_us32_n871 ), .ZN(_AES_ENC_us32_n875 ) );
NAND2_X2 _AES_ENC_us32_U192  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n875 ), .ZN(_AES_ENC_us32_n904 ) );
NAND2_X2 _AES_ENC_us32_U191  ( .A1(_AES_ENC_us32_n583 ), .A2(_AES_ENC_us32_n1050 ), .ZN(_AES_ENC_us32_n889 ) );
NAND2_X2 _AES_ENC_us32_U190  ( .A1(_AES_ENC_us32_n1093 ), .A2(_AES_ENC_us32_n587 ), .ZN(_AES_ENC_us32_n876 ) );
NAND2_X2 _AES_ENC_us32_U189  ( .A1(_AES_ENC_us32_n604 ), .A2(_AES_ENC_us32_n876 ), .ZN(_AES_ENC_us32_n877 ) );
NAND2_X2 _AES_ENC_us32_U188  ( .A1(_AES_ENC_us32_n877 ), .A2(_AES_ENC_us32_n623 ), .ZN(_AES_ENC_us32_n888 ) );
NAND4_X2 _AES_ENC_us32_U179  ( .A1(_AES_ENC_us32_n889 ), .A2(_AES_ENC_us32_n888 ), .A3(_AES_ENC_us32_n887 ), .A4(_AES_ENC_us32_n886 ), .ZN(_AES_ENC_us32_n890 ) );
NAND2_X2 _AES_ENC_us32_U178  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n890 ), .ZN(_AES_ENC_us32_n903 ) );
OR2_X2 _AES_ENC_us32_U177  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n1059 ), .ZN(_AES_ENC_us32_n900 ) );
NAND2_X2 _AES_ENC_us32_U176  ( .A1(_AES_ENC_us32_n1073 ), .A2(_AES_ENC_us32_n1047 ), .ZN(_AES_ENC_us32_n899 ) );
NAND2_X2 _AES_ENC_us32_U175  ( .A1(_AES_ENC_us32_n1094 ), .A2(_AES_ENC_us32_n595 ), .ZN(_AES_ENC_us32_n898 ) );
NAND4_X2 _AES_ENC_us32_U167  ( .A1(_AES_ENC_us32_n900 ), .A2(_AES_ENC_us32_n899 ), .A3(_AES_ENC_us32_n898 ), .A4(_AES_ENC_us32_n897 ), .ZN(_AES_ENC_us32_n901 ) );
NAND2_X2 _AES_ENC_us32_U166  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n901 ), .ZN(_AES_ENC_us32_n902 ) );
NAND4_X2 _AES_ENC_us32_U165  ( .A1(_AES_ENC_us32_n905 ), .A2(_AES_ENC_us32_n904 ), .A3(_AES_ENC_us32_n903 ), .A4(_AES_ENC_us32_n902 ), .ZN(_AES_ENC_sa32_sub[4] ) );
NAND2_X2 _AES_ENC_us32_U164  ( .A1(_AES_ENC_us32_n1094 ), .A2(_AES_ENC_us32_n599 ), .ZN(_AES_ENC_us32_n922 ) );
NAND2_X2 _AES_ENC_us32_U163  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n989 ), .ZN(_AES_ENC_us32_n921 ) );
NAND4_X2 _AES_ENC_us32_U151  ( .A1(_AES_ENC_us32_n922 ), .A2(_AES_ENC_us32_n921 ), .A3(_AES_ENC_us32_n920 ), .A4(_AES_ENC_us32_n919 ), .ZN(_AES_ENC_us32_n923 ) );
NAND2_X2 _AES_ENC_us32_U150  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n923 ), .ZN(_AES_ENC_us32_n972 ) );
NAND2_X2 _AES_ENC_us32_U149  ( .A1(_AES_ENC_us32_n582 ), .A2(_AES_ENC_us32_n619 ), .ZN(_AES_ENC_us32_n924 ) );
NAND2_X2 _AES_ENC_us32_U148  ( .A1(_AES_ENC_us32_n1073 ), .A2(_AES_ENC_us32_n924 ), .ZN(_AES_ENC_us32_n939 ) );
NAND2_X2 _AES_ENC_us32_U147  ( .A1(_AES_ENC_us32_n926 ), .A2(_AES_ENC_us32_n925 ), .ZN(_AES_ENC_us32_n927 ) );
NAND2_X2 _AES_ENC_us32_U146  ( .A1(_AES_ENC_us32_n606 ), .A2(_AES_ENC_us32_n927 ), .ZN(_AES_ENC_us32_n928 ) );
NAND2_X2 _AES_ENC_us32_U145  ( .A1(_AES_ENC_us32_n928 ), .A2(_AES_ENC_us32_n1080 ), .ZN(_AES_ENC_us32_n938 ) );
OR2_X2 _AES_ENC_us32_U144  ( .A1(_AES_ENC_us32_n1117 ), .A2(_AES_ENC_us32_n615 ), .ZN(_AES_ENC_us32_n937 ) );
NAND4_X2 _AES_ENC_us32_U139  ( .A1(_AES_ENC_us32_n939 ), .A2(_AES_ENC_us32_n938 ), .A3(_AES_ENC_us32_n937 ), .A4(_AES_ENC_us32_n936 ), .ZN(_AES_ENC_us32_n940 ) );
NAND2_X2 _AES_ENC_us32_U138  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n940 ), .ZN(_AES_ENC_us32_n971 ) );
OR2_X2 _AES_ENC_us32_U137  ( .A1(_AES_ENC_us32_n605 ), .A2(_AES_ENC_us32_n941 ), .ZN(_AES_ENC_us32_n954 ) );
NAND2_X2 _AES_ENC_us32_U136  ( .A1(_AES_ENC_us32_n1096 ), .A2(_AES_ENC_us32_n577 ), .ZN(_AES_ENC_us32_n942 ) );
NAND2_X2 _AES_ENC_us32_U135  ( .A1(_AES_ENC_us32_n1048 ), .A2(_AES_ENC_us32_n942 ), .ZN(_AES_ENC_us32_n943 ) );
NAND2_X2 _AES_ENC_us32_U134  ( .A1(_AES_ENC_us32_n612 ), .A2(_AES_ENC_us32_n943 ), .ZN(_AES_ENC_us32_n944 ) );
NAND2_X2 _AES_ENC_us32_U133  ( .A1(_AES_ENC_us32_n944 ), .A2(_AES_ENC_us32_n580 ), .ZN(_AES_ENC_us32_n953 ) );
NAND4_X2 _AES_ENC_us32_U125  ( .A1(_AES_ENC_us32_n954 ), .A2(_AES_ENC_us32_n953 ), .A3(_AES_ENC_us32_n952 ), .A4(_AES_ENC_us32_n951 ), .ZN(_AES_ENC_us32_n955 ) );
NAND2_X2 _AES_ENC_us32_U124  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n955 ), .ZN(_AES_ENC_us32_n970 ) );
NAND2_X2 _AES_ENC_us32_U123  ( .A1(_AES_ENC_us32_n1094 ), .A2(_AES_ENC_us32_n1071 ), .ZN(_AES_ENC_us32_n967 ) );
NAND2_X2 _AES_ENC_us32_U122  ( .A1(_AES_ENC_us32_n956 ), .A2(_AES_ENC_us32_n1030 ), .ZN(_AES_ENC_us32_n966 ) );
NAND4_X2 _AES_ENC_us32_U114  ( .A1(_AES_ENC_us32_n967 ), .A2(_AES_ENC_us32_n966 ), .A3(_AES_ENC_us32_n965 ), .A4(_AES_ENC_us32_n964 ), .ZN(_AES_ENC_us32_n968 ) );
NAND2_X2 _AES_ENC_us32_U113  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n968 ), .ZN(_AES_ENC_us32_n969 ) );
NAND4_X2 _AES_ENC_us32_U112  ( .A1(_AES_ENC_us32_n972 ), .A2(_AES_ENC_us32_n971 ), .A3(_AES_ENC_us32_n970 ), .A4(_AES_ENC_us32_n969 ), .ZN(_AES_ENC_sa32_sub[5] ) );
NAND2_X2 _AES_ENC_us32_U111  ( .A1(_AES_ENC_us32_n570 ), .A2(_AES_ENC_us32_n1097 ), .ZN(_AES_ENC_us32_n973 ) );
NAND2_X2 _AES_ENC_us32_U110  ( .A1(_AES_ENC_us32_n1073 ), .A2(_AES_ENC_us32_n973 ), .ZN(_AES_ENC_us32_n987 ) );
NAND2_X2 _AES_ENC_us32_U109  ( .A1(_AES_ENC_us32_n974 ), .A2(_AES_ENC_us32_n1077 ), .ZN(_AES_ENC_us32_n975 ) );
NAND2_X2 _AES_ENC_us32_U108  ( .A1(_AES_ENC_us32_n613 ), .A2(_AES_ENC_us32_n975 ), .ZN(_AES_ENC_us32_n976 ) );
NAND2_X2 _AES_ENC_us32_U107  ( .A1(_AES_ENC_us32_n977 ), .A2(_AES_ENC_us32_n976 ), .ZN(_AES_ENC_us32_n986 ) );
NAND4_X2 _AES_ENC_us32_U99  ( .A1(_AES_ENC_us32_n987 ), .A2(_AES_ENC_us32_n986 ), .A3(_AES_ENC_us32_n985 ), .A4(_AES_ENC_us32_n984 ), .ZN(_AES_ENC_us32_n988 ) );
NAND2_X2 _AES_ENC_us32_U98  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n988 ), .ZN(_AES_ENC_us32_n1044 ) );
NAND2_X2 _AES_ENC_us32_U97  ( .A1(_AES_ENC_us32_n1073 ), .A2(_AES_ENC_us32_n989 ), .ZN(_AES_ENC_us32_n1004 ) );
NAND2_X2 _AES_ENC_us32_U96  ( .A1(_AES_ENC_us32_n1092 ), .A2(_AES_ENC_us32_n619 ), .ZN(_AES_ENC_us32_n1003 ) );
NAND4_X2 _AES_ENC_us32_U85  ( .A1(_AES_ENC_us32_n1004 ), .A2(_AES_ENC_us32_n1003 ), .A3(_AES_ENC_us32_n1002 ), .A4(_AES_ENC_us32_n1001 ), .ZN(_AES_ENC_us32_n1005 ) );
NAND2_X2 _AES_ENC_us32_U84  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n1005 ), .ZN(_AES_ENC_us32_n1043 ) );
NAND2_X2 _AES_ENC_us32_U83  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n596 ), .ZN(_AES_ENC_us32_n1020 ) );
NAND2_X2 _AES_ENC_us32_U82  ( .A1(_AES_ENC_us32_n1050 ), .A2(_AES_ENC_us32_n624 ), .ZN(_AES_ENC_us32_n1019 ) );
NAND2_X2 _AES_ENC_us32_U77  ( .A1(_AES_ENC_us32_n1059 ), .A2(_AES_ENC_us32_n1114 ), .ZN(_AES_ENC_us32_n1012 ) );
NAND2_X2 _AES_ENC_us32_U76  ( .A1(_AES_ENC_us32_n1010 ), .A2(_AES_ENC_us32_n592 ), .ZN(_AES_ENC_us32_n1011 ) );
NAND2_X2 _AES_ENC_us32_U75  ( .A1(_AES_ENC_us32_n1012 ), .A2(_AES_ENC_us32_n1011 ), .ZN(_AES_ENC_us32_n1016 ) );
NAND4_X2 _AES_ENC_us32_U70  ( .A1(_AES_ENC_us32_n1020 ), .A2(_AES_ENC_us32_n1019 ), .A3(_AES_ENC_us32_n1018 ), .A4(_AES_ENC_us32_n1017 ), .ZN(_AES_ENC_us32_n1021 ) );
NAND2_X2 _AES_ENC_us32_U69  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n1021 ), .ZN(_AES_ENC_us32_n1042 ) );
NAND2_X2 _AES_ENC_us32_U68  ( .A1(_AES_ENC_us32_n1022 ), .A2(_AES_ENC_us32_n1093 ), .ZN(_AES_ENC_us32_n1039 ) );
NAND2_X2 _AES_ENC_us32_U67  ( .A1(_AES_ENC_us32_n1050 ), .A2(_AES_ENC_us32_n1023 ), .ZN(_AES_ENC_us32_n1038 ) );
NAND2_X2 _AES_ENC_us32_U66  ( .A1(_AES_ENC_us32_n1024 ), .A2(_AES_ENC_us32_n1071 ), .ZN(_AES_ENC_us32_n1037 ) );
AND2_X2 _AES_ENC_us32_U60  ( .A1(_AES_ENC_us32_n1030 ), .A2(_AES_ENC_us32_n602 ), .ZN(_AES_ENC_us32_n1078 ) );
NAND4_X2 _AES_ENC_us32_U56  ( .A1(_AES_ENC_us32_n1039 ), .A2(_AES_ENC_us32_n1038 ), .A3(_AES_ENC_us32_n1037 ), .A4(_AES_ENC_us32_n1036 ), .ZN(_AES_ENC_us32_n1040 ) );
NAND2_X2 _AES_ENC_us32_U55  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n1040 ), .ZN(_AES_ENC_us32_n1041 ) );
NAND4_X2 _AES_ENC_us32_U54  ( .A1(_AES_ENC_us32_n1044 ), .A2(_AES_ENC_us32_n1043 ), .A3(_AES_ENC_us32_n1042 ), .A4(_AES_ENC_us32_n1041 ), .ZN(_AES_ENC_sa32_sub[6] ) );
NAND2_X2 _AES_ENC_us32_U53  ( .A1(_AES_ENC_us32_n1072 ), .A2(_AES_ENC_us32_n1045 ), .ZN(_AES_ENC_us32_n1068 ) );
NAND2_X2 _AES_ENC_us32_U52  ( .A1(_AES_ENC_us32_n1046 ), .A2(_AES_ENC_us32_n582 ), .ZN(_AES_ENC_us32_n1067 ) );
NAND2_X2 _AES_ENC_us32_U51  ( .A1(_AES_ENC_us32_n1094 ), .A2(_AES_ENC_us32_n1047 ), .ZN(_AES_ENC_us32_n1066 ) );
NAND4_X2 _AES_ENC_us32_U40  ( .A1(_AES_ENC_us32_n1068 ), .A2(_AES_ENC_us32_n1067 ), .A3(_AES_ENC_us32_n1066 ), .A4(_AES_ENC_us32_n1065 ), .ZN(_AES_ENC_us32_n1069 ) );
NAND2_X2 _AES_ENC_us32_U39  ( .A1(_AES_ENC_us32_n1070 ), .A2(_AES_ENC_us32_n1069 ), .ZN(_AES_ENC_us32_n1135 ) );
NAND2_X2 _AES_ENC_us32_U38  ( .A1(_AES_ENC_us32_n1072 ), .A2(_AES_ENC_us32_n1071 ), .ZN(_AES_ENC_us32_n1088 ) );
NAND2_X2 _AES_ENC_us32_U37  ( .A1(_AES_ENC_us32_n1073 ), .A2(_AES_ENC_us32_n595 ), .ZN(_AES_ENC_us32_n1087 ) );
NAND4_X2 _AES_ENC_us32_U28  ( .A1(_AES_ENC_us32_n1088 ), .A2(_AES_ENC_us32_n1087 ), .A3(_AES_ENC_us32_n1086 ), .A4(_AES_ENC_us32_n1085 ), .ZN(_AES_ENC_us32_n1089 ) );
NAND2_X2 _AES_ENC_us32_U27  ( .A1(_AES_ENC_us32_n1090 ), .A2(_AES_ENC_us32_n1089 ), .ZN(_AES_ENC_us32_n1134 ) );
NAND2_X2 _AES_ENC_us32_U26  ( .A1(_AES_ENC_us32_n1091 ), .A2(_AES_ENC_us32_n1093 ), .ZN(_AES_ENC_us32_n1111 ) );
NAND2_X2 _AES_ENC_us32_U25  ( .A1(_AES_ENC_us32_n1092 ), .A2(_AES_ENC_us32_n1120 ), .ZN(_AES_ENC_us32_n1110 ) );
AND2_X2 _AES_ENC_us32_U22  ( .A1(_AES_ENC_us32_n1097 ), .A2(_AES_ENC_us32_n1096 ), .ZN(_AES_ENC_us32_n1098 ) );
NAND4_X2 _AES_ENC_us32_U14  ( .A1(_AES_ENC_us32_n1111 ), .A2(_AES_ENC_us32_n1110 ), .A3(_AES_ENC_us32_n1109 ), .A4(_AES_ENC_us32_n1108 ), .ZN(_AES_ENC_us32_n1112 ) );
NAND2_X2 _AES_ENC_us32_U13  ( .A1(_AES_ENC_us32_n1113 ), .A2(_AES_ENC_us32_n1112 ), .ZN(_AES_ENC_us32_n1133 ) );
NAND2_X2 _AES_ENC_us32_U12  ( .A1(_AES_ENC_us32_n1115 ), .A2(_AES_ENC_us32_n1114 ), .ZN(_AES_ENC_us32_n1129 ) );
OR2_X2 _AES_ENC_us32_U11  ( .A1(_AES_ENC_us32_n608 ), .A2(_AES_ENC_us32_n1116 ), .ZN(_AES_ENC_us32_n1128 ) );
NAND4_X2 _AES_ENC_us32_U3  ( .A1(_AES_ENC_us32_n1129 ), .A2(_AES_ENC_us32_n1128 ), .A3(_AES_ENC_us32_n1127 ), .A4(_AES_ENC_us32_n1126 ), .ZN(_AES_ENC_us32_n1130 ) );
NAND2_X2 _AES_ENC_us32_U2  ( .A1(_AES_ENC_us32_n1131 ), .A2(_AES_ENC_us32_n1130 ), .ZN(_AES_ENC_us32_n1132 ) );
NAND4_X2 _AES_ENC_us32_U1  ( .A1(_AES_ENC_us32_n1135 ), .A2(_AES_ENC_us32_n1134 ), .A3(_AES_ENC_us32_n1133 ), .A4(_AES_ENC_us32_n1132 ), .ZN(_AES_ENC_sa32_sub[7] ) );
INV_X4 _AES_ENC_us33_U575  ( .A(_AES_ENC_sa33[7]), .ZN(_AES_ENC_us33_n627 ));
INV_X4 _AES_ENC_us33_U574  ( .A(_AES_ENC_us33_n1114 ), .ZN(_AES_ENC_us33_n625 ) );
INV_X4 _AES_ENC_us33_U573  ( .A(_AES_ENC_sa33[4]), .ZN(_AES_ENC_us33_n624 ));
INV_X4 _AES_ENC_us33_U572  ( .A(_AES_ENC_us33_n1025 ), .ZN(_AES_ENC_us33_n622 ) );
INV_X4 _AES_ENC_us33_U571  ( .A(_AES_ENC_us33_n1120 ), .ZN(_AES_ENC_us33_n620 ) );
INV_X4 _AES_ENC_us33_U570  ( .A(_AES_ENC_us33_n1121 ), .ZN(_AES_ENC_us33_n619 ) );
INV_X4 _AES_ENC_us33_U569  ( .A(_AES_ENC_us33_n1048 ), .ZN(_AES_ENC_us33_n618 ) );
INV_X4 _AES_ENC_us33_U568  ( .A(_AES_ENC_us33_n974 ), .ZN(_AES_ENC_us33_n616 ) );
INV_X4 _AES_ENC_us33_U567  ( .A(_AES_ENC_us33_n794 ), .ZN(_AES_ENC_us33_n614 ) );
INV_X4 _AES_ENC_us33_U566  ( .A(_AES_ENC_sa33[2]), .ZN(_AES_ENC_us33_n611 ));
INV_X4 _AES_ENC_us33_U565  ( .A(_AES_ENC_us33_n800 ), .ZN(_AES_ENC_us33_n610 ) );
INV_X4 _AES_ENC_us33_U564  ( .A(_AES_ENC_us33_n925 ), .ZN(_AES_ENC_us33_n609 ) );
INV_X4 _AES_ENC_us33_U563  ( .A(_AES_ENC_us33_n779 ), .ZN(_AES_ENC_us33_n607 ) );
INV_X4 _AES_ENC_us33_U562  ( .A(_AES_ENC_us33_n1022 ), .ZN(_AES_ENC_us33_n603 ) );
INV_X4 _AES_ENC_us33_U561  ( .A(_AES_ENC_us33_n1102 ), .ZN(_AES_ENC_us33_n602 ) );
INV_X4 _AES_ENC_us33_U560  ( .A(_AES_ENC_us33_n929 ), .ZN(_AES_ENC_us33_n601 ) );
INV_X4 _AES_ENC_us33_U559  ( .A(_AES_ENC_us33_n1056 ), .ZN(_AES_ENC_us33_n600 ) );
INV_X4 _AES_ENC_us33_U558  ( .A(_AES_ENC_us33_n1054 ), .ZN(_AES_ENC_us33_n599 ) );
INV_X4 _AES_ENC_us33_U557  ( .A(_AES_ENC_us33_n881 ), .ZN(_AES_ENC_us33_n598 ) );
INV_X4 _AES_ENC_us33_U556  ( .A(_AES_ENC_us33_n926 ), .ZN(_AES_ENC_us33_n597 ) );
INV_X4 _AES_ENC_us33_U555  ( .A(_AES_ENC_us33_n977 ), .ZN(_AES_ENC_us33_n595 ) );
INV_X4 _AES_ENC_us33_U554  ( .A(_AES_ENC_us33_n1031 ), .ZN(_AES_ENC_us33_n594 ) );
INV_X4 _AES_ENC_us33_U553  ( .A(_AES_ENC_us33_n1103 ), .ZN(_AES_ENC_us33_n593 ) );
INV_X4 _AES_ENC_us33_U552  ( .A(_AES_ENC_us33_n1009 ), .ZN(_AES_ENC_us33_n592 ) );
INV_X4 _AES_ENC_us33_U551  ( .A(_AES_ENC_us33_n990 ), .ZN(_AES_ENC_us33_n591 ) );
INV_X4 _AES_ENC_us33_U550  ( .A(_AES_ENC_us33_n1058 ), .ZN(_AES_ENC_us33_n590 ) );
INV_X4 _AES_ENC_us33_U549  ( .A(_AES_ENC_us33_n1074 ), .ZN(_AES_ENC_us33_n589 ) );
INV_X4 _AES_ENC_us33_U548  ( .A(_AES_ENC_us33_n1053 ), .ZN(_AES_ENC_us33_n588 ) );
INV_X4 _AES_ENC_us33_U547  ( .A(_AES_ENC_us33_n826 ), .ZN(_AES_ENC_us33_n587 ) );
INV_X4 _AES_ENC_us33_U546  ( .A(_AES_ENC_us33_n992 ), .ZN(_AES_ENC_us33_n586 ) );
INV_X4 _AES_ENC_us33_U545  ( .A(_AES_ENC_us33_n821 ), .ZN(_AES_ENC_us33_n585 ) );
INV_X4 _AES_ENC_us33_U544  ( .A(_AES_ENC_us33_n910 ), .ZN(_AES_ENC_us33_n584 ) );
INV_X4 _AES_ENC_us33_U543  ( .A(_AES_ENC_us33_n906 ), .ZN(_AES_ENC_us33_n583 ) );
INV_X4 _AES_ENC_us33_U542  ( .A(_AES_ENC_us33_n880 ), .ZN(_AES_ENC_us33_n581 ) );
INV_X4 _AES_ENC_us33_U541  ( .A(_AES_ENC_us33_n1013 ), .ZN(_AES_ENC_us33_n580 ) );
INV_X4 _AES_ENC_us33_U540  ( .A(_AES_ENC_us33_n1092 ), .ZN(_AES_ENC_us33_n579 ) );
INV_X4 _AES_ENC_us33_U539  ( .A(_AES_ENC_us33_n824 ), .ZN(_AES_ENC_us33_n578 ) );
INV_X4 _AES_ENC_us33_U538  ( .A(_AES_ENC_us33_n1091 ), .ZN(_AES_ENC_us33_n577 ) );
INV_X4 _AES_ENC_us33_U537  ( .A(_AES_ENC_us33_n1080 ), .ZN(_AES_ENC_us33_n576 ) );
INV_X4 _AES_ENC_us33_U536  ( .A(_AES_ENC_us33_n959 ), .ZN(_AES_ENC_us33_n575 ) );
INV_X4 _AES_ENC_us33_U535  ( .A(_AES_ENC_sa33[0]), .ZN(_AES_ENC_us33_n574 ));
NOR2_X2 _AES_ENC_us33_U534  ( .A1(_AES_ENC_sa33[0]), .A2(_AES_ENC_sa33[6]),.ZN(_AES_ENC_us33_n1090 ) );
NOR2_X2 _AES_ENC_us33_U533  ( .A1(_AES_ENC_us33_n574 ), .A2(_AES_ENC_sa33[6]), .ZN(_AES_ENC_us33_n1070 ) );
NOR2_X2 _AES_ENC_us33_U532  ( .A1(_AES_ENC_sa33[4]), .A2(_AES_ENC_sa33[3]),.ZN(_AES_ENC_us33_n1025 ) );
INV_X4 _AES_ENC_us33_U531  ( .A(_AES_ENC_us33_n569 ), .ZN(_AES_ENC_us33_n572 ) );
NOR2_X2 _AES_ENC_us33_U530  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n765 ) );
NOR2_X2 _AES_ENC_us33_U529  ( .A1(_AES_ENC_sa33[4]), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n764 ) );
NOR2_X2 _AES_ENC_us33_U528  ( .A1(_AES_ENC_us33_n765 ), .A2(_AES_ENC_us33_n764 ), .ZN(_AES_ENC_us33_n766 ) );
NOR2_X2 _AES_ENC_us33_U527  ( .A1(_AES_ENC_us33_n766 ), .A2(_AES_ENC_us33_n575 ), .ZN(_AES_ENC_us33_n767 ) );
NOR3_X2 _AES_ENC_us33_U526  ( .A1(_AES_ENC_us33_n627 ), .A2(_AES_ENC_sa33[5]), .A3(_AES_ENC_us33_n704 ), .ZN(_AES_ENC_us33_n706 ));
NOR2_X2 _AES_ENC_us33_U525  ( .A1(_AES_ENC_us33_n1117 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n707 ) );
NOR2_X2 _AES_ENC_us33_U524  ( .A1(_AES_ENC_sa33[4]), .A2(_AES_ENC_us33_n579 ), .ZN(_AES_ENC_us33_n705 ) );
NOR3_X2 _AES_ENC_us33_U523  ( .A1(_AES_ENC_us33_n707 ), .A2(_AES_ENC_us33_n706 ), .A3(_AES_ENC_us33_n705 ), .ZN(_AES_ENC_us33_n713 ) );
INV_X4 _AES_ENC_us33_U522  ( .A(_AES_ENC_sa33[3]), .ZN(_AES_ENC_us33_n621 ));
NAND3_X2 _AES_ENC_us33_U521  ( .A1(_AES_ENC_us33_n652 ), .A2(_AES_ENC_us33_n626 ), .A3(_AES_ENC_sa33[7]), .ZN(_AES_ENC_us33_n653 ));
NOR2_X2 _AES_ENC_us33_U520  ( .A1(_AES_ENC_us33_n611 ), .A2(_AES_ENC_sa33[5]), .ZN(_AES_ENC_us33_n925 ) );
NOR2_X2 _AES_ENC_us33_U519  ( .A1(_AES_ENC_sa33[5]), .A2(_AES_ENC_sa33[2]),.ZN(_AES_ENC_us33_n974 ) );
INV_X4 _AES_ENC_us33_U518  ( .A(_AES_ENC_sa33[5]), .ZN(_AES_ENC_us33_n626 ));
NOR2_X2 _AES_ENC_us33_U517  ( .A1(_AES_ENC_us33_n611 ), .A2(_AES_ENC_sa33[7]), .ZN(_AES_ENC_us33_n779 ) );
NAND3_X2 _AES_ENC_us33_U516  ( .A1(_AES_ENC_us33_n679 ), .A2(_AES_ENC_us33_n678 ), .A3(_AES_ENC_us33_n677 ), .ZN(_AES_ENC_sa33_sub[0] ) );
NOR2_X2 _AES_ENC_us33_U515  ( .A1(_AES_ENC_us33_n626 ), .A2(_AES_ENC_sa33[2]), .ZN(_AES_ENC_us33_n1048 ) );
NOR4_X2 _AES_ENC_us33_U512  ( .A1(_AES_ENC_us33_n633 ), .A2(_AES_ENC_us33_n632 ), .A3(_AES_ENC_us33_n631 ), .A4(_AES_ENC_us33_n630 ), .ZN(_AES_ENC_us33_n634 ) );
NOR2_X2 _AES_ENC_us33_U510  ( .A1(_AES_ENC_us33_n629 ), .A2(_AES_ENC_us33_n628 ), .ZN(_AES_ENC_us33_n635 ) );
NAND3_X2 _AES_ENC_us33_U509  ( .A1(_AES_ENC_sa33[2]), .A2(_AES_ENC_sa33[7]), .A3(_AES_ENC_us33_n1059 ), .ZN(_AES_ENC_us33_n636 ) );
NOR2_X2 _AES_ENC_us33_U508  ( .A1(_AES_ENC_sa33[7]), .A2(_AES_ENC_sa33[2]),.ZN(_AES_ENC_us33_n794 ) );
NOR2_X2 _AES_ENC_us33_U507  ( .A1(_AES_ENC_sa33[4]), .A2(_AES_ENC_sa33[1]),.ZN(_AES_ENC_us33_n1102 ) );
NOR2_X2 _AES_ENC_us33_U506  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_sa33[3]), .ZN(_AES_ENC_us33_n1053 ) );
NOR2_X2 _AES_ENC_us33_U505  ( .A1(_AES_ENC_us33_n607 ), .A2(_AES_ENC_sa33[5]), .ZN(_AES_ENC_us33_n1024 ) );
NOR2_X2 _AES_ENC_us33_U504  ( .A1(_AES_ENC_us33_n625 ), .A2(_AES_ENC_sa33[2]), .ZN(_AES_ENC_us33_n1093 ) );
NOR2_X2 _AES_ENC_us33_U503  ( .A1(_AES_ENC_us33_n614 ), .A2(_AES_ENC_sa33[5]), .ZN(_AES_ENC_us33_n1094 ) );
NOR2_X2 _AES_ENC_us33_U502  ( .A1(_AES_ENC_us33_n624 ), .A2(_AES_ENC_sa33[3]), .ZN(_AES_ENC_us33_n931 ) );
INV_X4 _AES_ENC_us33_U501  ( .A(_AES_ENC_us33_n570 ), .ZN(_AES_ENC_us33_n573 ) );
NOR2_X2 _AES_ENC_us33_U500  ( .A1(_AES_ENC_us33_n1053 ), .A2(_AES_ENC_us33_n1095 ), .ZN(_AES_ENC_us33_n639 ) );
NOR3_X2 _AES_ENC_us33_U499  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n573 ), .A3(_AES_ENC_us33_n1074 ), .ZN(_AES_ENC_us33_n641 ) );
NOR2_X2 _AES_ENC_us33_U498  ( .A1(_AES_ENC_us33_n639 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n640 ) );
NOR2_X2 _AES_ENC_us33_U497  ( .A1(_AES_ENC_us33_n641 ), .A2(_AES_ENC_us33_n640 ), .ZN(_AES_ENC_us33_n646 ) );
NOR3_X2 _AES_ENC_us33_U496  ( .A1(_AES_ENC_us33_n995 ), .A2(_AES_ENC_us33_n586 ), .A3(_AES_ENC_us33_n994 ), .ZN(_AES_ENC_us33_n1002 ) );
NOR2_X2 _AES_ENC_us33_U495  ( .A1(_AES_ENC_us33_n909 ), .A2(_AES_ENC_us33_n908 ), .ZN(_AES_ENC_us33_n920 ) );
NOR2_X2 _AES_ENC_us33_U494  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n823 ) );
NOR2_X2 _AES_ENC_us33_U492  ( .A1(_AES_ENC_us33_n624 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n822 ) );
NOR2_X2 _AES_ENC_us33_U491  ( .A1(_AES_ENC_us33_n823 ), .A2(_AES_ENC_us33_n822 ), .ZN(_AES_ENC_us33_n825 ) );
NOR2_X2 _AES_ENC_us33_U490  ( .A1(_AES_ENC_sa33[1]), .A2(_AES_ENC_us33_n623 ), .ZN(_AES_ENC_us33_n913 ) );
NOR2_X2 _AES_ENC_us33_U489  ( .A1(_AES_ENC_us33_n913 ), .A2(_AES_ENC_us33_n1091 ), .ZN(_AES_ENC_us33_n914 ) );
NOR2_X2 _AES_ENC_us33_U488  ( .A1(_AES_ENC_us33_n826 ), .A2(_AES_ENC_us33_n572 ), .ZN(_AES_ENC_us33_n827 ) );
NOR3_X2 _AES_ENC_us33_U487  ( .A1(_AES_ENC_us33_n769 ), .A2(_AES_ENC_us33_n768 ), .A3(_AES_ENC_us33_n767 ), .ZN(_AES_ENC_us33_n775 ) );
NOR2_X2 _AES_ENC_us33_U486  ( .A1(_AES_ENC_us33_n1056 ), .A2(_AES_ENC_us33_n1053 ), .ZN(_AES_ENC_us33_n749 ) );
NOR2_X2 _AES_ENC_us33_U483  ( .A1(_AES_ENC_us33_n749 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n752 ) );
INV_X4 _AES_ENC_us33_U482  ( .A(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n596 ));
NOR2_X2 _AES_ENC_us33_U480  ( .A1(_AES_ENC_us33_n1054 ), .A2(_AES_ENC_us33_n1053 ), .ZN(_AES_ENC_us33_n1055 ) );
OR2_X4 _AES_ENC_us33_U479  ( .A1(_AES_ENC_us33_n1094 ), .A2(_AES_ENC_us33_n1093 ), .ZN(_AES_ENC_us33_n571 ) );
AND2_X2 _AES_ENC_us33_U478  ( .A1(_AES_ENC_us33_n571 ), .A2(_AES_ENC_us33_n1095 ), .ZN(_AES_ENC_us33_n1101 ) );
NOR2_X2 _AES_ENC_us33_U477  ( .A1(_AES_ENC_us33_n1074 ), .A2(_AES_ENC_us33_n931 ), .ZN(_AES_ENC_us33_n796 ) );
NOR2_X2 _AES_ENC_us33_U474  ( .A1(_AES_ENC_us33_n796 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n797 ) );
NOR2_X2 _AES_ENC_us33_U473  ( .A1(_AES_ENC_us33_n932 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n933 ) );
NOR2_X2 _AES_ENC_us33_U472  ( .A1(_AES_ENC_us33_n929 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n935 ) );
NOR2_X2 _AES_ENC_us33_U471  ( .A1(_AES_ENC_us33_n931 ), .A2(_AES_ENC_us33_n930 ), .ZN(_AES_ENC_us33_n934 ) );
NOR3_X2 _AES_ENC_us33_U470  ( .A1(_AES_ENC_us33_n935 ), .A2(_AES_ENC_us33_n934 ), .A3(_AES_ENC_us33_n933 ), .ZN(_AES_ENC_us33_n936 ) );
NOR2_X2 _AES_ENC_us33_U469  ( .A1(_AES_ENC_us33_n624 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n1075 ) );
NOR2_X2 _AES_ENC_us33_U468  ( .A1(_AES_ENC_us33_n572 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n949 ) );
NOR2_X2 _AES_ENC_us33_U467  ( .A1(_AES_ENC_us33_n1049 ), .A2(_AES_ENC_us33_n618 ), .ZN(_AES_ENC_us33_n1051 ) );
NOR2_X2 _AES_ENC_us33_U466  ( .A1(_AES_ENC_us33_n1051 ), .A2(_AES_ENC_us33_n1050 ), .ZN(_AES_ENC_us33_n1052 ) );
NOR2_X2 _AES_ENC_us33_U465  ( .A1(_AES_ENC_us33_n1052 ), .A2(_AES_ENC_us33_n592 ), .ZN(_AES_ENC_us33_n1064 ) );
NOR2_X2 _AES_ENC_us33_U464  ( .A1(_AES_ENC_sa33[1]), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n631 ) );
NOR2_X2 _AES_ENC_us33_U463  ( .A1(_AES_ENC_us33_n1025 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n980 ) );
NOR2_X2 _AES_ENC_us33_U462  ( .A1(_AES_ENC_us33_n1073 ), .A2(_AES_ENC_us33_n1094 ), .ZN(_AES_ENC_us33_n795 ) );
NOR2_X2 _AES_ENC_us33_U461  ( .A1(_AES_ENC_us33_n795 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n799 ) );
NOR2_X2 _AES_ENC_us33_U460  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n981 ) );
NOR2_X2 _AES_ENC_us33_U459  ( .A1(_AES_ENC_us33_n1102 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n643 ) );
NOR2_X2 _AES_ENC_us33_U458  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n621 ), .ZN(_AES_ENC_us33_n642 ) );
NOR2_X2 _AES_ENC_us33_U455  ( .A1(_AES_ENC_us33_n911 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n644 ) );
NOR4_X2 _AES_ENC_us33_U448  ( .A1(_AES_ENC_us33_n644 ), .A2(_AES_ENC_us33_n643 ), .A3(_AES_ENC_us33_n804 ), .A4(_AES_ENC_us33_n642 ), .ZN(_AES_ENC_us33_n645 ) );
NOR2_X2 _AES_ENC_us33_U447  ( .A1(_AES_ENC_us33_n1102 ), .A2(_AES_ENC_us33_n910 ), .ZN(_AES_ENC_us33_n932 ) );
NOR2_X2 _AES_ENC_us33_U442  ( .A1(_AES_ENC_us33_n1102 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n755 ) );
NOR2_X2 _AES_ENC_us33_U441  ( .A1(_AES_ENC_us33_n931 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n743 ) );
NOR2_X2 _AES_ENC_us33_U438  ( .A1(_AES_ENC_us33_n1072 ), .A2(_AES_ENC_us33_n1094 ), .ZN(_AES_ENC_us33_n930 ) );
NOR2_X2 _AES_ENC_us33_U435  ( .A1(_AES_ENC_us33_n1074 ), .A2(_AES_ENC_us33_n1025 ), .ZN(_AES_ENC_us33_n891 ) );
NOR2_X2 _AES_ENC_us33_U434  ( .A1(_AES_ENC_us33_n891 ), .A2(_AES_ENC_us33_n609 ), .ZN(_AES_ENC_us33_n894 ) );
NOR3_X2 _AES_ENC_us33_U433  ( .A1(_AES_ENC_us33_n623 ), .A2(_AES_ENC_sa33[1]), .A3(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n683 ));
INV_X4 _AES_ENC_us33_U428  ( .A(_AES_ENC_us33_n931 ), .ZN(_AES_ENC_us33_n623 ) );
NOR2_X2 _AES_ENC_us33_U427  ( .A1(_AES_ENC_us33_n996 ), .A2(_AES_ENC_us33_n931 ), .ZN(_AES_ENC_us33_n704 ) );
NOR2_X2 _AES_ENC_us33_U421  ( .A1(_AES_ENC_us33_n931 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n685 ) );
NOR2_X2 _AES_ENC_us33_U420  ( .A1(_AES_ENC_us33_n1029 ), .A2(_AES_ENC_us33_n1025 ), .ZN(_AES_ENC_us33_n1079 ) );
NOR3_X2 _AES_ENC_us33_U419  ( .A1(_AES_ENC_us33_n589 ), .A2(_AES_ENC_us33_n1025 ), .A3(_AES_ENC_us33_n616 ), .ZN(_AES_ENC_us33_n945 ) );
NOR2_X2 _AES_ENC_us33_U418  ( .A1(_AES_ENC_us33_n626 ), .A2(_AES_ENC_us33_n611 ), .ZN(_AES_ENC_us33_n800 ) );
NOR3_X2 _AES_ENC_us33_U417  ( .A1(_AES_ENC_us33_n590 ), .A2(_AES_ENC_us33_n627 ), .A3(_AES_ENC_us33_n611 ), .ZN(_AES_ENC_us33_n798 ) );
NOR3_X2 _AES_ENC_us33_U416  ( .A1(_AES_ENC_us33_n610 ), .A2(_AES_ENC_us33_n572 ), .A3(_AES_ENC_us33_n575 ), .ZN(_AES_ENC_us33_n962 ) );
NOR3_X2 _AES_ENC_us33_U415  ( .A1(_AES_ENC_us33_n959 ), .A2(_AES_ENC_us33_n572 ), .A3(_AES_ENC_us33_n609 ), .ZN(_AES_ENC_us33_n768 ) );
NOR3_X2 _AES_ENC_us33_U414  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n572 ), .A3(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n694 ) );
NOR3_X2 _AES_ENC_us33_U413  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n572 ), .A3(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n895 ) );
NOR3_X2 _AES_ENC_us33_U410  ( .A1(_AES_ENC_us33_n1008 ), .A2(_AES_ENC_us33_n1007 ), .A3(_AES_ENC_us33_n1006 ), .ZN(_AES_ENC_us33_n1018 ) );
NOR4_X2 _AES_ENC_us33_U409  ( .A1(_AES_ENC_us33_n806 ), .A2(_AES_ENC_us33_n805 ), .A3(_AES_ENC_us33_n804 ), .A4(_AES_ENC_us33_n803 ), .ZN(_AES_ENC_us33_n807 ) );
NOR3_X2 _AES_ENC_us33_U406  ( .A1(_AES_ENC_us33_n799 ), .A2(_AES_ENC_us33_n798 ), .A3(_AES_ENC_us33_n797 ), .ZN(_AES_ENC_us33_n808 ) );
NOR4_X2 _AES_ENC_us33_U405  ( .A1(_AES_ENC_us33_n843 ), .A2(_AES_ENC_us33_n842 ), .A3(_AES_ENC_us33_n841 ), .A4(_AES_ENC_us33_n840 ), .ZN(_AES_ENC_us33_n844 ) );
NOR3_X2 _AES_ENC_us33_U404  ( .A1(_AES_ENC_us33_n1101 ), .A2(_AES_ENC_us33_n1100 ), .A3(_AES_ENC_us33_n1099 ), .ZN(_AES_ENC_us33_n1109 ) );
NOR4_X2 _AES_ENC_us33_U403  ( .A1(_AES_ENC_us33_n711 ), .A2(_AES_ENC_us33_n710 ), .A3(_AES_ENC_us33_n709 ), .A4(_AES_ENC_us33_n708 ), .ZN(_AES_ENC_us33_n712 ) );
NOR4_X2 _AES_ENC_us33_U401  ( .A1(_AES_ENC_us33_n963 ), .A2(_AES_ENC_us33_n962 ), .A3(_AES_ENC_us33_n961 ), .A4(_AES_ENC_us33_n960 ), .ZN(_AES_ENC_us33_n964 ) );
NOR2_X2 _AES_ENC_us33_U400  ( .A1(_AES_ENC_us33_n669 ), .A2(_AES_ENC_us33_n668 ), .ZN(_AES_ENC_us33_n673 ) );
NOR4_X2 _AES_ENC_us33_U399  ( .A1(_AES_ENC_us33_n946 ), .A2(_AES_ENC_us33_n1046 ), .A3(_AES_ENC_us33_n671 ), .A4(_AES_ENC_us33_n670 ), .ZN(_AES_ENC_us33_n672 ) );
NOR3_X2 _AES_ENC_us33_U398  ( .A1(_AES_ENC_us33_n743 ), .A2(_AES_ENC_us33_n742 ), .A3(_AES_ENC_us33_n741 ), .ZN(_AES_ENC_us33_n744 ) );
NOR2_X2 _AES_ENC_us33_U397  ( .A1(_AES_ENC_us33_n697 ), .A2(_AES_ENC_us33_n658 ), .ZN(_AES_ENC_us33_n659 ) );
NOR2_X2 _AES_ENC_us33_U396  ( .A1(_AES_ENC_us33_n1078 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n1033 ) );
NOR2_X2 _AES_ENC_us33_U393  ( .A1(_AES_ENC_us33_n1031 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n1032 ) );
NOR3_X2 _AES_ENC_us33_U390  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n1025 ), .A3(_AES_ENC_us33_n1074 ), .ZN(_AES_ENC_us33_n1035 ) );
NOR4_X2 _AES_ENC_us33_U389  ( .A1(_AES_ENC_us33_n1035 ), .A2(_AES_ENC_us33_n1034 ), .A3(_AES_ENC_us33_n1033 ), .A4(_AES_ENC_us33_n1032 ), .ZN(_AES_ENC_us33_n1036 ) );
NOR2_X2 _AES_ENC_us33_U388  ( .A1(_AES_ENC_us33_n598 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n885 ) );
NOR2_X2 _AES_ENC_us33_U387  ( .A1(_AES_ENC_us33_n623 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n882 ) );
NOR2_X2 _AES_ENC_us33_U386  ( .A1(_AES_ENC_us33_n1053 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n884 ) );
NOR4_X2 _AES_ENC_us33_U385  ( .A1(_AES_ENC_us33_n885 ), .A2(_AES_ENC_us33_n884 ), .A3(_AES_ENC_us33_n883 ), .A4(_AES_ENC_us33_n882 ), .ZN(_AES_ENC_us33_n886 ) );
NOR2_X2 _AES_ENC_us33_U384  ( .A1(_AES_ENC_us33_n825 ), .A2(_AES_ENC_us33_n578 ), .ZN(_AES_ENC_us33_n830 ) );
NOR2_X2 _AES_ENC_us33_U383  ( .A1(_AES_ENC_us33_n827 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n829 ) );
NOR2_X2 _AES_ENC_us33_U382  ( .A1(_AES_ENC_us33_n572 ), .A2(_AES_ENC_us33_n579 ), .ZN(_AES_ENC_us33_n828 ) );
NOR4_X2 _AES_ENC_us33_U374  ( .A1(_AES_ENC_us33_n831 ), .A2(_AES_ENC_us33_n830 ), .A3(_AES_ENC_us33_n829 ), .A4(_AES_ENC_us33_n828 ), .ZN(_AES_ENC_us33_n832 ) );
NOR2_X2 _AES_ENC_us33_U373  ( .A1(_AES_ENC_us33_n606 ), .A2(_AES_ENC_us33_n582 ), .ZN(_AES_ENC_us33_n1104 ) );
NOR2_X2 _AES_ENC_us33_U372  ( .A1(_AES_ENC_us33_n1102 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n1106 ) );
NOR2_X2 _AES_ENC_us33_U370  ( .A1(_AES_ENC_us33_n1103 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n1105 ) );
NOR4_X2 _AES_ENC_us33_U369  ( .A1(_AES_ENC_us33_n1107 ), .A2(_AES_ENC_us33_n1106 ), .A3(_AES_ENC_us33_n1105 ), .A4(_AES_ENC_us33_n1104 ), .ZN(_AES_ENC_us33_n1108 ) );
NOR3_X2 _AES_ENC_us33_U368  ( .A1(_AES_ENC_us33_n959 ), .A2(_AES_ENC_us33_n621 ), .A3(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n963 ) );
NOR2_X2 _AES_ENC_us33_U367  ( .A1(_AES_ENC_us33_n626 ), .A2(_AES_ENC_us33_n627 ), .ZN(_AES_ENC_us33_n1114 ) );
INV_X4 _AES_ENC_us33_U366  ( .A(_AES_ENC_us33_n1024 ), .ZN(_AES_ENC_us33_n606 ) );
NOR3_X2 _AES_ENC_us33_U365  ( .A1(_AES_ENC_us33_n910 ), .A2(_AES_ENC_us33_n1059 ), .A3(_AES_ENC_us33_n611 ), .ZN(_AES_ENC_us33_n1115 ) );
INV_X4 _AES_ENC_us33_U364  ( .A(_AES_ENC_us33_n1094 ), .ZN(_AES_ENC_us33_n613 ) );
NOR2_X2 _AES_ENC_us33_U363  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n931 ), .ZN(_AES_ENC_us33_n1100 ) );
INV_X4 _AES_ENC_us33_U354  ( .A(_AES_ENC_us33_n1093 ), .ZN(_AES_ENC_us33_n617 ) );
NOR2_X2 _AES_ENC_us33_U353  ( .A1(_AES_ENC_us33_n569 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n929 ) );
NOR2_X2 _AES_ENC_us33_U352  ( .A1(_AES_ENC_us33_n620 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n926 ) );
NOR2_X2 _AES_ENC_us33_U351  ( .A1(_AES_ENC_us33_n572 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n1095 ) );
NOR2_X2 _AES_ENC_us33_U350  ( .A1(_AES_ENC_us33_n609 ), .A2(_AES_ENC_us33_n627 ), .ZN(_AES_ENC_us33_n1010 ) );
NOR2_X2 _AES_ENC_us33_U349  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n1103 ) );
NOR2_X2 _AES_ENC_us33_U348  ( .A1(_AES_ENC_us33_n622 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n1059 ) );
NOR2_X2 _AES_ENC_us33_U347  ( .A1(_AES_ENC_sa33[1]), .A2(_AES_ENC_us33_n1120 ), .ZN(_AES_ENC_us33_n1022 ) );
NOR2_X2 _AES_ENC_us33_U346  ( .A1(_AES_ENC_us33_n619 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n911 ) );
NOR2_X2 _AES_ENC_us33_U345  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_us33_n1025 ), .ZN(_AES_ENC_us33_n826 ) );
NOR2_X2 _AES_ENC_us33_U338  ( .A1(_AES_ENC_us33_n626 ), .A2(_AES_ENC_us33_n607 ), .ZN(_AES_ENC_us33_n1072 ) );
NOR2_X2 _AES_ENC_us33_U335  ( .A1(_AES_ENC_us33_n627 ), .A2(_AES_ENC_us33_n616 ), .ZN(_AES_ENC_us33_n956 ) );
NOR2_X2 _AES_ENC_us33_U329  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_us33_n624 ), .ZN(_AES_ENC_us33_n1121 ) );
NOR2_X2 _AES_ENC_us33_U328  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_us33_n624 ), .ZN(_AES_ENC_us33_n1058 ) );
NOR2_X2 _AES_ENC_us33_U327  ( .A1(_AES_ENC_us33_n625 ), .A2(_AES_ENC_us33_n611 ), .ZN(_AES_ENC_us33_n1073 ) );
NOR2_X2 _AES_ENC_us33_U325  ( .A1(_AES_ENC_sa33[1]), .A2(_AES_ENC_us33_n1025 ), .ZN(_AES_ENC_us33_n1054 ) );
NOR2_X2 _AES_ENC_us33_U324  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_us33_n931 ), .ZN(_AES_ENC_us33_n1029 ) );
NOR2_X2 _AES_ENC_us33_U319  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n1056 ) );
NOR2_X2 _AES_ENC_us33_U318  ( .A1(_AES_ENC_us33_n614 ), .A2(_AES_ENC_us33_n626 ), .ZN(_AES_ENC_us33_n1050 ) );
NOR2_X2 _AES_ENC_us33_U317  ( .A1(_AES_ENC_us33_n1121 ), .A2(_AES_ENC_us33_n1025 ), .ZN(_AES_ENC_us33_n1120 ) );
NOR2_X2 _AES_ENC_us33_U316  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_us33_n572 ), .ZN(_AES_ENC_us33_n1074 ) );
NOR2_X2 _AES_ENC_us33_U315  ( .A1(_AES_ENC_us33_n1058 ), .A2(_AES_ENC_us33_n1054 ), .ZN(_AES_ENC_us33_n878 ) );
NOR2_X2 _AES_ENC_us33_U314  ( .A1(_AES_ENC_us33_n878 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n879 ) );
NOR2_X2 _AES_ENC_us33_U312  ( .A1(_AES_ENC_us33_n880 ), .A2(_AES_ENC_us33_n879 ), .ZN(_AES_ENC_us33_n887 ) );
NOR2_X2 _AES_ENC_us33_U311  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n588 ), .ZN(_AES_ENC_us33_n957 ) );
NOR2_X2 _AES_ENC_us33_U310  ( .A1(_AES_ENC_us33_n958 ), .A2(_AES_ENC_us33_n957 ), .ZN(_AES_ENC_us33_n965 ) );
NOR3_X2 _AES_ENC_us33_U309  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n1091 ), .A3(_AES_ENC_us33_n1022 ), .ZN(_AES_ENC_us33_n720 ) );
NOR3_X2 _AES_ENC_us33_U303  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n1054 ), .A3(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n719 ) );
NOR2_X2 _AES_ENC_us33_U302  ( .A1(_AES_ENC_us33_n720 ), .A2(_AES_ENC_us33_n719 ), .ZN(_AES_ENC_us33_n726 ) );
NOR2_X2 _AES_ENC_us33_U300  ( .A1(_AES_ENC_us33_n614 ), .A2(_AES_ENC_us33_n591 ), .ZN(_AES_ENC_us33_n865 ) );
NOR2_X2 _AES_ENC_us33_U299  ( .A1(_AES_ENC_us33_n1059 ), .A2(_AES_ENC_us33_n1058 ), .ZN(_AES_ENC_us33_n1060 ) );
NOR2_X2 _AES_ENC_us33_U298  ( .A1(_AES_ENC_us33_n1095 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n668 ) );
NOR2_X2 _AES_ENC_us33_U297  ( .A1(_AES_ENC_us33_n911 ), .A2(_AES_ENC_us33_n910 ), .ZN(_AES_ENC_us33_n912 ) );
NOR2_X2 _AES_ENC_us33_U296  ( .A1(_AES_ENC_us33_n912 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n916 ) );
NOR2_X2 _AES_ENC_us33_U295  ( .A1(_AES_ENC_us33_n826 ), .A2(_AES_ENC_us33_n573 ), .ZN(_AES_ENC_us33_n750 ) );
NOR2_X2 _AES_ENC_us33_U294  ( .A1(_AES_ENC_us33_n750 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n751 ) );
NOR2_X2 _AES_ENC_us33_U293  ( .A1(_AES_ENC_us33_n907 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n908 ) );
NOR2_X2 _AES_ENC_us33_U292  ( .A1(_AES_ENC_us33_n990 ), .A2(_AES_ENC_us33_n926 ), .ZN(_AES_ENC_us33_n780 ) );
NOR2_X2 _AES_ENC_us33_U291  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n584 ), .ZN(_AES_ENC_us33_n838 ) );
NOR2_X2 _AES_ENC_us33_U290  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n602 ), .ZN(_AES_ENC_us33_n837 ) );
NOR2_X2 _AES_ENC_us33_U284  ( .A1(_AES_ENC_us33_n838 ), .A2(_AES_ENC_us33_n837 ), .ZN(_AES_ENC_us33_n845 ) );
NOR2_X2 _AES_ENC_us33_U283  ( .A1(_AES_ENC_us33_n1022 ), .A2(_AES_ENC_us33_n1058 ), .ZN(_AES_ENC_us33_n740 ) );
NOR2_X2 _AES_ENC_us33_U282  ( .A1(_AES_ENC_us33_n740 ), .A2(_AES_ENC_us33_n616 ), .ZN(_AES_ENC_us33_n742 ) );
NOR2_X2 _AES_ENC_us33_U281  ( .A1(_AES_ENC_us33_n1098 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n1099 ) );
NOR2_X2 _AES_ENC_us33_U280  ( .A1(_AES_ENC_us33_n1120 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n993 ) );
NOR2_X2 _AES_ENC_us33_U279  ( .A1(_AES_ENC_us33_n993 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n994 ) );
NOR2_X2 _AES_ENC_us33_U273  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n620 ), .ZN(_AES_ENC_us33_n1026 ) );
NOR2_X2 _AES_ENC_us33_U272  ( .A1(_AES_ENC_us33_n573 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n1027 ) );
NOR2_X2 _AES_ENC_us33_U271  ( .A1(_AES_ENC_us33_n1027 ), .A2(_AES_ENC_us33_n1026 ), .ZN(_AES_ENC_us33_n1028 ) );
NOR2_X2 _AES_ENC_us33_U270  ( .A1(_AES_ENC_us33_n1029 ), .A2(_AES_ENC_us33_n1028 ), .ZN(_AES_ENC_us33_n1034 ) );
NOR4_X2 _AES_ENC_us33_U269  ( .A1(_AES_ENC_us33_n757 ), .A2(_AES_ENC_us33_n756 ), .A3(_AES_ENC_us33_n755 ), .A4(_AES_ENC_us33_n754 ), .ZN(_AES_ENC_us33_n758 ) );
NOR2_X2 _AES_ENC_us33_U268  ( .A1(_AES_ENC_us33_n752 ), .A2(_AES_ENC_us33_n751 ), .ZN(_AES_ENC_us33_n759 ) );
NOR2_X2 _AES_ENC_us33_U267  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n1071 ), .ZN(_AES_ENC_us33_n669 ) );
NOR2_X2 _AES_ENC_us33_U263  ( .A1(_AES_ENC_us33_n1056 ), .A2(_AES_ENC_us33_n990 ), .ZN(_AES_ENC_us33_n991 ) );
NOR2_X2 _AES_ENC_us33_U262  ( .A1(_AES_ENC_us33_n991 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n995 ) );
NOR2_X2 _AES_ENC_us33_U258  ( .A1(_AES_ENC_us33_n607 ), .A2(_AES_ENC_us33_n590 ), .ZN(_AES_ENC_us33_n1008 ) );
NOR2_X2 _AES_ENC_us33_U255  ( .A1(_AES_ENC_us33_n839 ), .A2(_AES_ENC_us33_n582 ), .ZN(_AES_ENC_us33_n693 ) );
NOR2_X2 _AES_ENC_us33_U254  ( .A1(_AES_ENC_us33_n606 ), .A2(_AES_ENC_us33_n906 ), .ZN(_AES_ENC_us33_n741 ) );
NOR2_X2 _AES_ENC_us33_U253  ( .A1(_AES_ENC_us33_n1054 ), .A2(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n763 ) );
NOR2_X2 _AES_ENC_us33_U252  ( .A1(_AES_ENC_us33_n763 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n769 ) );
NOR2_X2 _AES_ENC_us33_U251  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n577 ), .ZN(_AES_ENC_us33_n1007 ) );
NOR2_X2 _AES_ENC_us33_U250  ( .A1(_AES_ENC_us33_n609 ), .A2(_AES_ENC_us33_n580 ), .ZN(_AES_ENC_us33_n1123 ) );
NOR2_X2 _AES_ENC_us33_U243  ( .A1(_AES_ENC_us33_n609 ), .A2(_AES_ENC_us33_n590 ), .ZN(_AES_ENC_us33_n710 ) );
INV_X4 _AES_ENC_us33_U242  ( .A(_AES_ENC_us33_n1029 ), .ZN(_AES_ENC_us33_n582 ) );
NOR2_X2 _AES_ENC_us33_U241  ( .A1(_AES_ENC_us33_n616 ), .A2(_AES_ENC_us33_n597 ), .ZN(_AES_ENC_us33_n883 ) );
NOR2_X2 _AES_ENC_us33_U240  ( .A1(_AES_ENC_us33_n593 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n1125 ) );
NOR2_X2 _AES_ENC_us33_U239  ( .A1(_AES_ENC_us33_n990 ), .A2(_AES_ENC_us33_n929 ), .ZN(_AES_ENC_us33_n892 ) );
NOR2_X2 _AES_ENC_us33_U238  ( .A1(_AES_ENC_us33_n892 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n893 ) );
NOR2_X2 _AES_ENC_us33_U237  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n602 ), .ZN(_AES_ENC_us33_n950 ) );
NOR2_X2 _AES_ENC_us33_U236  ( .A1(_AES_ENC_us33_n1079 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n1082 ) );
NOR2_X2 _AES_ENC_us33_U235  ( .A1(_AES_ENC_us33_n910 ), .A2(_AES_ENC_us33_n1056 ), .ZN(_AES_ENC_us33_n941 ) );
NOR2_X2 _AES_ENC_us33_U234  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n1077 ), .ZN(_AES_ENC_us33_n841 ) );
NOR2_X2 _AES_ENC_us33_U229  ( .A1(_AES_ENC_us33_n623 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n630 ) );
NOR2_X2 _AES_ENC_us33_U228  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n602 ), .ZN(_AES_ENC_us33_n806 ) );
NOR2_X2 _AES_ENC_us33_U227  ( .A1(_AES_ENC_us33_n623 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n948 ) );
NOR2_X2 _AES_ENC_us33_U226  ( .A1(_AES_ENC_us33_n606 ), .A2(_AES_ENC_us33_n589 ), .ZN(_AES_ENC_us33_n997 ) );
NOR2_X2 _AES_ENC_us33_U225  ( .A1(_AES_ENC_us33_n1121 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n1122 ) );
NOR2_X2 _AES_ENC_us33_U223  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n1023 ), .ZN(_AES_ENC_us33_n756 ) );
NOR2_X2 _AES_ENC_us33_U222  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n602 ), .ZN(_AES_ENC_us33_n870 ) );
NOR2_X2 _AES_ENC_us33_U221  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n569 ), .ZN(_AES_ENC_us33_n947 ) );
NOR2_X2 _AES_ENC_us33_U217  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n1077 ), .ZN(_AES_ENC_us33_n1084 ) );
NOR2_X2 _AES_ENC_us33_U213  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n855 ), .ZN(_AES_ENC_us33_n709 ) );
NOR2_X2 _AES_ENC_us33_U212  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n589 ), .ZN(_AES_ENC_us33_n868 ) );
NOR2_X2 _AES_ENC_us33_U211  ( .A1(_AES_ENC_us33_n1120 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n1124 ) );
NOR2_X2 _AES_ENC_us33_U210  ( .A1(_AES_ENC_us33_n1120 ), .A2(_AES_ENC_us33_n839 ), .ZN(_AES_ENC_us33_n842 ) );
NOR2_X2 _AES_ENC_us33_U209  ( .A1(_AES_ENC_us33_n1120 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n696 ) );
NOR2_X2 _AES_ENC_us33_U208  ( .A1(_AES_ENC_us33_n1074 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n1076 ) );
NOR2_X2 _AES_ENC_us33_U207  ( .A1(_AES_ENC_us33_n1074 ), .A2(_AES_ENC_us33_n620 ), .ZN(_AES_ENC_us33_n781 ) );
NOR3_X2 _AES_ENC_us33_U201  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n1056 ), .A3(_AES_ENC_us33_n990 ), .ZN(_AES_ENC_us33_n979 ) );
NOR3_X2 _AES_ENC_us33_U200  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n1058 ), .A3(_AES_ENC_us33_n1059 ), .ZN(_AES_ENC_us33_n854 ) );
NOR2_X2 _AES_ENC_us33_U199  ( .A1(_AES_ENC_us33_n996 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n869 ) );
NOR2_X2 _AES_ENC_us33_U198  ( .A1(_AES_ENC_us33_n1056 ), .A2(_AES_ENC_us33_n1074 ), .ZN(_AES_ENC_us33_n1057 ) );
NOR3_X2 _AES_ENC_us33_U197  ( .A1(_AES_ENC_us33_n607 ), .A2(_AES_ENC_us33_n1120 ), .A3(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n978 ) );
NOR2_X2 _AES_ENC_us33_U196  ( .A1(_AES_ENC_us33_n996 ), .A2(_AES_ENC_us33_n911 ), .ZN(_AES_ENC_us33_n1116 ) );
NOR2_X2 _AES_ENC_us33_U195  ( .A1(_AES_ENC_us33_n1074 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n754 ) );
NOR2_X2 _AES_ENC_us33_U194  ( .A1(_AES_ENC_us33_n926 ), .A2(_AES_ENC_us33_n1103 ), .ZN(_AES_ENC_us33_n977 ) );
NOR2_X2 _AES_ENC_us33_U187  ( .A1(_AES_ENC_us33_n839 ), .A2(_AES_ENC_us33_n824 ), .ZN(_AES_ENC_us33_n1092 ) );
NOR2_X2 _AES_ENC_us33_U186  ( .A1(_AES_ENC_us33_n573 ), .A2(_AES_ENC_us33_n1074 ), .ZN(_AES_ENC_us33_n684 ) );
NOR2_X2 _AES_ENC_us33_U185  ( .A1(_AES_ENC_us33_n826 ), .A2(_AES_ENC_us33_n1059 ), .ZN(_AES_ENC_us33_n907 ) );
NOR3_X2 _AES_ENC_us33_U184  ( .A1(_AES_ENC_us33_n625 ), .A2(_AES_ENC_us33_n1115 ), .A3(_AES_ENC_us33_n585 ), .ZN(_AES_ENC_us33_n831 ) );
NOR3_X2 _AES_ENC_us33_U183  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n1056 ), .A3(_AES_ENC_us33_n990 ), .ZN(_AES_ENC_us33_n896 ) );
NOR3_X2 _AES_ENC_us33_U182  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n573 ), .A3(_AES_ENC_us33_n1013 ), .ZN(_AES_ENC_us33_n670 ) );
NOR3_X2 _AES_ENC_us33_U181  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n1091 ), .A3(_AES_ENC_us33_n1022 ), .ZN(_AES_ENC_us33_n843 ) );
NOR2_X2 _AES_ENC_us33_U180  ( .A1(_AES_ENC_us33_n1029 ), .A2(_AES_ENC_us33_n1095 ), .ZN(_AES_ENC_us33_n735 ) );
NOR2_X2 _AES_ENC_us33_U174  ( .A1(_AES_ENC_us33_n1100 ), .A2(_AES_ENC_us33_n854 ), .ZN(_AES_ENC_us33_n860 ) );
NOR4_X2 _AES_ENC_us33_U173  ( .A1(_AES_ENC_us33_n1125 ), .A2(_AES_ENC_us33_n1124 ), .A3(_AES_ENC_us33_n1123 ), .A4(_AES_ENC_us33_n1122 ), .ZN(_AES_ENC_us33_n1126 ) );
NOR4_X2 _AES_ENC_us33_U172  ( .A1(_AES_ENC_us33_n1084 ), .A2(_AES_ENC_us33_n1083 ), .A3(_AES_ENC_us33_n1082 ), .A4(_AES_ENC_us33_n1081 ), .ZN(_AES_ENC_us33_n1085 ) );
NOR2_X2 _AES_ENC_us33_U171  ( .A1(_AES_ENC_us33_n1076 ), .A2(_AES_ENC_us33_n1075 ), .ZN(_AES_ENC_us33_n1086 ) );
NAND3_X2 _AES_ENC_us33_U170  ( .A1(_AES_ENC_us33_n569 ), .A2(_AES_ENC_us33_n582 ), .A3(_AES_ENC_us33_n681 ), .ZN(_AES_ENC_us33_n691 ) );
NOR2_X2 _AES_ENC_us33_U169  ( .A1(_AES_ENC_us33_n683 ), .A2(_AES_ENC_us33_n682 ), .ZN(_AES_ENC_us33_n690 ) );
NOR3_X2 _AES_ENC_us33_U168  ( .A1(_AES_ENC_us33_n695 ), .A2(_AES_ENC_us33_n694 ), .A3(_AES_ENC_us33_n693 ), .ZN(_AES_ENC_us33_n700 ) );
NOR4_X2 _AES_ENC_us33_U162  ( .A1(_AES_ENC_us33_n983 ), .A2(_AES_ENC_us33_n698 ), .A3(_AES_ENC_us33_n697 ), .A4(_AES_ENC_us33_n696 ), .ZN(_AES_ENC_us33_n699 ) );
NOR2_X2 _AES_ENC_us33_U161  ( .A1(_AES_ENC_us33_n946 ), .A2(_AES_ENC_us33_n945 ), .ZN(_AES_ENC_us33_n952 ) );
NOR4_X2 _AES_ENC_us33_U160  ( .A1(_AES_ENC_us33_n950 ), .A2(_AES_ENC_us33_n949 ), .A3(_AES_ENC_us33_n948 ), .A4(_AES_ENC_us33_n947 ), .ZN(_AES_ENC_us33_n951 ) );
NOR4_X2 _AES_ENC_us33_U159  ( .A1(_AES_ENC_us33_n983 ), .A2(_AES_ENC_us33_n982 ), .A3(_AES_ENC_us33_n981 ), .A4(_AES_ENC_us33_n980 ), .ZN(_AES_ENC_us33_n984 ) );
NOR2_X2 _AES_ENC_us33_U158  ( .A1(_AES_ENC_us33_n979 ), .A2(_AES_ENC_us33_n978 ), .ZN(_AES_ENC_us33_n985 ) );
NOR4_X2 _AES_ENC_us33_U157  ( .A1(_AES_ENC_us33_n896 ), .A2(_AES_ENC_us33_n895 ), .A3(_AES_ENC_us33_n894 ), .A4(_AES_ENC_us33_n893 ), .ZN(_AES_ENC_us33_n897 ) );
NOR2_X2 _AES_ENC_us33_U156  ( .A1(_AES_ENC_us33_n866 ), .A2(_AES_ENC_us33_n865 ), .ZN(_AES_ENC_us33_n872 ) );
NOR4_X2 _AES_ENC_us33_U155  ( .A1(_AES_ENC_us33_n870 ), .A2(_AES_ENC_us33_n869 ), .A3(_AES_ENC_us33_n868 ), .A4(_AES_ENC_us33_n867 ), .ZN(_AES_ENC_us33_n871 ) );
NOR3_X2 _AES_ENC_us33_U154  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n1054 ), .A3(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n961 ) );
NOR3_X2 _AES_ENC_us33_U153  ( .A1(_AES_ENC_us33_n620 ), .A2(_AES_ENC_us33_n1074 ), .A3(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n671 ) );
NOR2_X2 _AES_ENC_us33_U152  ( .A1(_AES_ENC_us33_n1057 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n1062 ) );
NOR2_X2 _AES_ENC_us33_U143  ( .A1(_AES_ENC_us33_n1055 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n1063 ) );
NOR2_X2 _AES_ENC_us33_U142  ( .A1(_AES_ENC_us33_n1060 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n1061 ) );
NOR4_X2 _AES_ENC_us33_U141  ( .A1(_AES_ENC_us33_n1064 ), .A2(_AES_ENC_us33_n1063 ), .A3(_AES_ENC_us33_n1062 ), .A4(_AES_ENC_us33_n1061 ), .ZN(_AES_ENC_us33_n1065 ) );
NOR3_X2 _AES_ENC_us33_U140  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n1120 ), .A3(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n918 ) );
NOR3_X2 _AES_ENC_us33_U132  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n573 ), .A3(_AES_ENC_us33_n1013 ), .ZN(_AES_ENC_us33_n917 ) );
NOR2_X2 _AES_ENC_us33_U131  ( .A1(_AES_ENC_us33_n914 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n915 ) );
NOR4_X2 _AES_ENC_us33_U130  ( .A1(_AES_ENC_us33_n918 ), .A2(_AES_ENC_us33_n917 ), .A3(_AES_ENC_us33_n916 ), .A4(_AES_ENC_us33_n915 ), .ZN(_AES_ENC_us33_n919 ) );
NOR2_X2 _AES_ENC_us33_U129  ( .A1(_AES_ENC_us33_n735 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n687 ) );
NOR2_X2 _AES_ENC_us33_U128  ( .A1(_AES_ENC_us33_n684 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n688 ) );
NOR2_X2 _AES_ENC_us33_U127  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n600 ), .ZN(_AES_ENC_us33_n686 ) );
NOR4_X2 _AES_ENC_us33_U126  ( .A1(_AES_ENC_us33_n688 ), .A2(_AES_ENC_us33_n687 ), .A3(_AES_ENC_us33_n686 ), .A4(_AES_ENC_us33_n685 ), .ZN(_AES_ENC_us33_n689 ) );
NOR2_X2 _AES_ENC_us33_U121  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n595 ), .ZN(_AES_ENC_us33_n858 ) );
NOR2_X2 _AES_ENC_us33_U120  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n855 ), .ZN(_AES_ENC_us33_n857 ) );
NOR2_X2 _AES_ENC_us33_U119  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n587 ), .ZN(_AES_ENC_us33_n856 ) );
NOR4_X2 _AES_ENC_us33_U118  ( .A1(_AES_ENC_us33_n858 ), .A2(_AES_ENC_us33_n857 ), .A3(_AES_ENC_us33_n856 ), .A4(_AES_ENC_us33_n958 ), .ZN(_AES_ENC_us33_n859 ) );
NOR2_X2 _AES_ENC_us33_U117  ( .A1(_AES_ENC_us33_n616 ), .A2(_AES_ENC_us33_n580 ), .ZN(_AES_ENC_us33_n771 ) );
NOR2_X2 _AES_ENC_us33_U116  ( .A1(_AES_ENC_us33_n1103 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n772 ) );
NOR2_X2 _AES_ENC_us33_U115  ( .A1(_AES_ENC_us33_n610 ), .A2(_AES_ENC_us33_n599 ), .ZN(_AES_ENC_us33_n773 ) );
NOR4_X2 _AES_ENC_us33_U106  ( .A1(_AES_ENC_us33_n773 ), .A2(_AES_ENC_us33_n772 ), .A3(_AES_ENC_us33_n771 ), .A4(_AES_ENC_us33_n770 ), .ZN(_AES_ENC_us33_n774 ) );
NOR2_X2 _AES_ENC_us33_U105  ( .A1(_AES_ENC_us33_n780 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n784 ) );
NOR2_X2 _AES_ENC_us33_U104  ( .A1(_AES_ENC_us33_n1117 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n782 ) );
NOR2_X2 _AES_ENC_us33_U103  ( .A1(_AES_ENC_us33_n781 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n783 ) );
NOR4_X2 _AES_ENC_us33_U102  ( .A1(_AES_ENC_us33_n880 ), .A2(_AES_ENC_us33_n784 ), .A3(_AES_ENC_us33_n783 ), .A4(_AES_ENC_us33_n782 ), .ZN(_AES_ENC_us33_n785 ) );
NOR2_X2 _AES_ENC_us33_U101  ( .A1(_AES_ENC_us33_n583 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n814 ) );
NOR2_X2 _AES_ENC_us33_U100  ( .A1(_AES_ENC_us33_n907 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n813 ) );
NOR3_X2 _AES_ENC_us33_U95  ( .A1(_AES_ENC_us33_n606 ), .A2(_AES_ENC_us33_n1058 ), .A3(_AES_ENC_us33_n1059 ), .ZN(_AES_ENC_us33_n815 ) );
NOR4_X2 _AES_ENC_us33_U94  ( .A1(_AES_ENC_us33_n815 ), .A2(_AES_ENC_us33_n814 ), .A3(_AES_ENC_us33_n813 ), .A4(_AES_ENC_us33_n812 ), .ZN(_AES_ENC_us33_n816 ) );
NOR2_X2 _AES_ENC_us33_U93  ( .A1(_AES_ENC_us33_n617 ), .A2(_AES_ENC_us33_n569 ), .ZN(_AES_ENC_us33_n721 ) );
NOR2_X2 _AES_ENC_us33_U92  ( .A1(_AES_ENC_us33_n1031 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n723 ) );
NOR2_X2 _AES_ENC_us33_U91  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n1096 ), .ZN(_AES_ENC_us33_n722 ) );
NOR4_X2 _AES_ENC_us33_U90  ( .A1(_AES_ENC_us33_n724 ), .A2(_AES_ENC_us33_n723 ), .A3(_AES_ENC_us33_n722 ), .A4(_AES_ENC_us33_n721 ), .ZN(_AES_ENC_us33_n725 ) );
NOR2_X2 _AES_ENC_us33_U89  ( .A1(_AES_ENC_us33_n911 ), .A2(_AES_ENC_us33_n990 ), .ZN(_AES_ENC_us33_n1009 ) );
NOR2_X2 _AES_ENC_us33_U88  ( .A1(_AES_ENC_us33_n1013 ), .A2(_AES_ENC_us33_n573 ), .ZN(_AES_ENC_us33_n1014 ) );
NOR2_X2 _AES_ENC_us33_U87  ( .A1(_AES_ENC_us33_n1014 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n1015 ) );
NOR4_X2 _AES_ENC_us33_U86  ( .A1(_AES_ENC_us33_n1016 ), .A2(_AES_ENC_us33_n1015 ), .A3(_AES_ENC_us33_n1119 ), .A4(_AES_ENC_us33_n1046 ), .ZN(_AES_ENC_us33_n1017 ) );
NOR2_X2 _AES_ENC_us33_U81  ( .A1(_AES_ENC_us33_n996 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n998 ) );
NOR2_X2 _AES_ENC_us33_U80  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n577 ), .ZN(_AES_ENC_us33_n1000 ) );
NOR2_X2 _AES_ENC_us33_U79  ( .A1(_AES_ENC_us33_n616 ), .A2(_AES_ENC_us33_n1096 ), .ZN(_AES_ENC_us33_n999 ) );
NOR4_X2 _AES_ENC_us33_U78  ( .A1(_AES_ENC_us33_n1000 ), .A2(_AES_ENC_us33_n999 ), .A3(_AES_ENC_us33_n998 ), .A4(_AES_ENC_us33_n997 ), .ZN(_AES_ENC_us33_n1001 ) );
NOR2_X2 _AES_ENC_us33_U74  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n1096 ), .ZN(_AES_ENC_us33_n697 ) );
NOR2_X2 _AES_ENC_us33_U73  ( .A1(_AES_ENC_us33_n620 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n958 ) );
NOR2_X2 _AES_ENC_us33_U72  ( .A1(_AES_ENC_us33_n911 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n983 ) );
NOR2_X2 _AES_ENC_us33_U71  ( .A1(_AES_ENC_us33_n1054 ), .A2(_AES_ENC_us33_n1103 ), .ZN(_AES_ENC_us33_n1031 ) );
INV_X4 _AES_ENC_us33_U65  ( .A(_AES_ENC_us33_n1050 ), .ZN(_AES_ENC_us33_n612 ) );
INV_X4 _AES_ENC_us33_U64  ( .A(_AES_ENC_us33_n1072 ), .ZN(_AES_ENC_us33_n605 ) );
INV_X4 _AES_ENC_us33_U63  ( .A(_AES_ENC_us33_n1073 ), .ZN(_AES_ENC_us33_n604 ) );
NOR2_X2 _AES_ENC_us33_U62  ( .A1(_AES_ENC_us33_n582 ), .A2(_AES_ENC_us33_n613 ), .ZN(_AES_ENC_us33_n880 ) );
NOR3_X2 _AES_ENC_us33_U61  ( .A1(_AES_ENC_us33_n826 ), .A2(_AES_ENC_us33_n1121 ), .A3(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n946 ) );
INV_X4 _AES_ENC_us33_U59  ( .A(_AES_ENC_us33_n1010 ), .ZN(_AES_ENC_us33_n608 ) );
NOR3_X2 _AES_ENC_us33_U58  ( .A1(_AES_ENC_us33_n573 ), .A2(_AES_ENC_us33_n1029 ), .A3(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n1119 ) );
INV_X4 _AES_ENC_us33_U57  ( .A(_AES_ENC_us33_n956 ), .ZN(_AES_ENC_us33_n615 ) );
NOR2_X2 _AES_ENC_us33_U50  ( .A1(_AES_ENC_us33_n623 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n1013 ) );
NOR2_X2 _AES_ENC_us33_U49  ( .A1(_AES_ENC_us33_n620 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n910 ) );
NOR2_X2 _AES_ENC_us33_U48  ( .A1(_AES_ENC_us33_n569 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n1091 ) );
NOR2_X2 _AES_ENC_us33_U47  ( .A1(_AES_ENC_us33_n622 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n990 ) );
NOR2_X2 _AES_ENC_us33_U46  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_us33_n1121 ), .ZN(_AES_ENC_us33_n996 ) );
NOR2_X2 _AES_ENC_us33_U45  ( .A1(_AES_ENC_us33_n610 ), .A2(_AES_ENC_us33_n600 ), .ZN(_AES_ENC_us33_n628 ) );
NOR2_X2 _AES_ENC_us33_U44  ( .A1(_AES_ENC_us33_n576 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n866 ) );
NOR2_X2 _AES_ENC_us33_U43  ( .A1(_AES_ENC_us33_n603 ), .A2(_AES_ENC_us33_n610 ), .ZN(_AES_ENC_us33_n1006 ) );
NOR2_X2 _AES_ENC_us33_U42  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n1117 ), .ZN(_AES_ENC_us33_n1118 ) );
NOR2_X2 _AES_ENC_us33_U41  ( .A1(_AES_ENC_us33_n1119 ), .A2(_AES_ENC_us33_n1118 ), .ZN(_AES_ENC_us33_n1127 ) );
NOR2_X2 _AES_ENC_us33_U36  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n906 ), .ZN(_AES_ENC_us33_n909 ) );
NOR2_X2 _AES_ENC_us33_U35  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n594 ), .ZN(_AES_ENC_us33_n629 ) );
NOR2_X2 _AES_ENC_us33_U34  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n597 ), .ZN(_AES_ENC_us33_n658 ) );
NOR2_X2 _AES_ENC_us33_U33  ( .A1(_AES_ENC_us33_n1116 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n695 ) );
NOR2_X2 _AES_ENC_us33_U32  ( .A1(_AES_ENC_us33_n1078 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n1083 ) );
NOR2_X2 _AES_ENC_us33_U31  ( .A1(_AES_ENC_us33_n941 ), .A2(_AES_ENC_us33_n608 ), .ZN(_AES_ENC_us33_n724 ) );
NOR2_X2 _AES_ENC_us33_U30  ( .A1(_AES_ENC_us33_n598 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n1107 ) );
NOR2_X2 _AES_ENC_us33_U29  ( .A1(_AES_ENC_us33_n576 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n840 ) );
NOR2_X2 _AES_ENC_us33_U24  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n593 ), .ZN(_AES_ENC_us33_n633 ) );
NOR2_X2 _AES_ENC_us33_U23  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n1080 ), .ZN(_AES_ENC_us33_n1081 ) );
NOR2_X2 _AES_ENC_us33_U21  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n1045 ), .ZN(_AES_ENC_us33_n812 ) );
NOR2_X2 _AES_ENC_us33_U20  ( .A1(_AES_ENC_us33_n1009 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n960 ) );
NOR2_X2 _AES_ENC_us33_U19  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n601 ), .ZN(_AES_ENC_us33_n982 ) );
NOR2_X2 _AES_ENC_us33_U18  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n594 ), .ZN(_AES_ENC_us33_n757 ) );
NOR2_X2 _AES_ENC_us33_U17  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n590 ), .ZN(_AES_ENC_us33_n698 ) );
NOR2_X2 _AES_ENC_us33_U16  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n619 ), .ZN(_AES_ENC_us33_n708 ) );
NOR2_X2 _AES_ENC_us33_U15  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n582 ), .ZN(_AES_ENC_us33_n770 ) );
NOR2_X2 _AES_ENC_us33_U10  ( .A1(_AES_ENC_us33_n619 ), .A2(_AES_ENC_us33_n604 ), .ZN(_AES_ENC_us33_n803 ) );
NOR2_X2 _AES_ENC_us33_U9  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n881 ), .ZN(_AES_ENC_us33_n711 ) );
NOR2_X2 _AES_ENC_us33_U8  ( .A1(_AES_ENC_us33_n615 ), .A2(_AES_ENC_us33_n582 ), .ZN(_AES_ENC_us33_n867 ) );
NOR2_X2 _AES_ENC_us33_U7  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n599 ), .ZN(_AES_ENC_us33_n804 ) );
NOR2_X2 _AES_ENC_us33_U6  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n620 ), .ZN(_AES_ENC_us33_n1046 ) );
OR2_X4 _AES_ENC_us33_U5  ( .A1(_AES_ENC_us33_n624 ), .A2(_AES_ENC_sa33[1]),.ZN(_AES_ENC_us33_n570 ) );
OR2_X4 _AES_ENC_us33_U4  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_sa33[4]),.ZN(_AES_ENC_us33_n569 ) );
NAND2_X2 _AES_ENC_us33_U514  ( .A1(_AES_ENC_us33_n1121 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n1030 ) );
AND2_X2 _AES_ENC_us33_U513  ( .A1(_AES_ENC_us33_n597 ), .A2(_AES_ENC_us33_n1030 ), .ZN(_AES_ENC_us33_n1049 ) );
NAND2_X2 _AES_ENC_us33_U511  ( .A1(_AES_ENC_us33_n1049 ), .A2(_AES_ENC_us33_n794 ), .ZN(_AES_ENC_us33_n637 ) );
AND2_X2 _AES_ENC_us33_U493  ( .A1(_AES_ENC_us33_n779 ), .A2(_AES_ENC_us33_n996 ), .ZN(_AES_ENC_us33_n632 ) );
NAND4_X2 _AES_ENC_us33_U485  ( .A1(_AES_ENC_us33_n637 ), .A2(_AES_ENC_us33_n636 ), .A3(_AES_ENC_us33_n635 ), .A4(_AES_ENC_us33_n634 ), .ZN(_AES_ENC_us33_n638 ) );
NAND2_X2 _AES_ENC_us33_U484  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n638 ), .ZN(_AES_ENC_us33_n679 ) );
NAND2_X2 _AES_ENC_us33_U481  ( .A1(_AES_ENC_us33_n1094 ), .A2(_AES_ENC_us33_n591 ), .ZN(_AES_ENC_us33_n648 ) );
NAND2_X2 _AES_ENC_us33_U476  ( .A1(_AES_ENC_us33_n601 ), .A2(_AES_ENC_us33_n590 ), .ZN(_AES_ENC_us33_n762 ) );
NAND2_X2 _AES_ENC_us33_U475  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n762 ), .ZN(_AES_ENC_us33_n647 ) );
NAND4_X2 _AES_ENC_us33_U457  ( .A1(_AES_ENC_us33_n648 ), .A2(_AES_ENC_us33_n647 ), .A3(_AES_ENC_us33_n646 ), .A4(_AES_ENC_us33_n645 ), .ZN(_AES_ENC_us33_n649 ) );
NAND2_X2 _AES_ENC_us33_U456  ( .A1(_AES_ENC_sa33[0]), .A2(_AES_ENC_us33_n649 ), .ZN(_AES_ENC_us33_n665 ) );
NAND2_X2 _AES_ENC_us33_U454  ( .A1(_AES_ENC_us33_n596 ), .A2(_AES_ENC_us33_n623 ), .ZN(_AES_ENC_us33_n855 ) );
NAND2_X2 _AES_ENC_us33_U453  ( .A1(_AES_ENC_us33_n587 ), .A2(_AES_ENC_us33_n855 ), .ZN(_AES_ENC_us33_n821 ) );
NAND2_X2 _AES_ENC_us33_U452  ( .A1(_AES_ENC_us33_n1093 ), .A2(_AES_ENC_us33_n821 ), .ZN(_AES_ENC_us33_n662 ) );
NAND2_X2 _AES_ENC_us33_U451  ( .A1(_AES_ENC_us33_n619 ), .A2(_AES_ENC_us33_n589 ), .ZN(_AES_ENC_us33_n650 ) );
NAND2_X2 _AES_ENC_us33_U450  ( .A1(_AES_ENC_us33_n956 ), .A2(_AES_ENC_us33_n650 ), .ZN(_AES_ENC_us33_n661 ) );
NAND2_X2 _AES_ENC_us33_U449  ( .A1(_AES_ENC_us33_n626 ), .A2(_AES_ENC_us33_n627 ), .ZN(_AES_ENC_us33_n839 ) );
OR2_X2 _AES_ENC_us33_U446  ( .A1(_AES_ENC_us33_n839 ), .A2(_AES_ENC_us33_n932 ), .ZN(_AES_ENC_us33_n656 ) );
NAND2_X2 _AES_ENC_us33_U445  ( .A1(_AES_ENC_us33_n621 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n1096 ) );
NAND2_X2 _AES_ENC_us33_U444  ( .A1(_AES_ENC_us33_n1030 ), .A2(_AES_ENC_us33_n1096 ), .ZN(_AES_ENC_us33_n651 ) );
NAND2_X2 _AES_ENC_us33_U443  ( .A1(_AES_ENC_us33_n1114 ), .A2(_AES_ENC_us33_n651 ), .ZN(_AES_ENC_us33_n655 ) );
OR3_X2 _AES_ENC_us33_U440  ( .A1(_AES_ENC_us33_n1079 ), .A2(_AES_ENC_sa33[7]), .A3(_AES_ENC_us33_n626 ), .ZN(_AES_ENC_us33_n654 ));
NAND2_X2 _AES_ENC_us33_U439  ( .A1(_AES_ENC_us33_n593 ), .A2(_AES_ENC_us33_n601 ), .ZN(_AES_ENC_us33_n652 ) );
NAND4_X2 _AES_ENC_us33_U437  ( .A1(_AES_ENC_us33_n656 ), .A2(_AES_ENC_us33_n655 ), .A3(_AES_ENC_us33_n654 ), .A4(_AES_ENC_us33_n653 ), .ZN(_AES_ENC_us33_n657 ) );
NAND2_X2 _AES_ENC_us33_U436  ( .A1(_AES_ENC_sa33[2]), .A2(_AES_ENC_us33_n657 ), .ZN(_AES_ENC_us33_n660 ) );
NAND4_X2 _AES_ENC_us33_U432  ( .A1(_AES_ENC_us33_n662 ), .A2(_AES_ENC_us33_n661 ), .A3(_AES_ENC_us33_n660 ), .A4(_AES_ENC_us33_n659 ), .ZN(_AES_ENC_us33_n663 ) );
NAND2_X2 _AES_ENC_us33_U431  ( .A1(_AES_ENC_us33_n663 ), .A2(_AES_ENC_us33_n574 ), .ZN(_AES_ENC_us33_n664 ) );
NAND2_X2 _AES_ENC_us33_U430  ( .A1(_AES_ENC_us33_n665 ), .A2(_AES_ENC_us33_n664 ), .ZN(_AES_ENC_us33_n666 ) );
NAND2_X2 _AES_ENC_us33_U429  ( .A1(_AES_ENC_sa33[6]), .A2(_AES_ENC_us33_n666 ), .ZN(_AES_ENC_us33_n678 ) );
NAND2_X2 _AES_ENC_us33_U426  ( .A1(_AES_ENC_us33_n735 ), .A2(_AES_ENC_us33_n1093 ), .ZN(_AES_ENC_us33_n675 ) );
NAND2_X2 _AES_ENC_us33_U425  ( .A1(_AES_ENC_us33_n588 ), .A2(_AES_ENC_us33_n597 ), .ZN(_AES_ENC_us33_n1045 ) );
OR2_X2 _AES_ENC_us33_U424  ( .A1(_AES_ENC_us33_n1045 ), .A2(_AES_ENC_us33_n605 ), .ZN(_AES_ENC_us33_n674 ) );
NAND2_X2 _AES_ENC_us33_U423  ( .A1(_AES_ENC_sa33[1]), .A2(_AES_ENC_us33_n620 ), .ZN(_AES_ENC_us33_n667 ) );
NAND2_X2 _AES_ENC_us33_U422  ( .A1(_AES_ENC_us33_n619 ), .A2(_AES_ENC_us33_n667 ), .ZN(_AES_ENC_us33_n1071 ) );
NAND4_X2 _AES_ENC_us33_U412  ( .A1(_AES_ENC_us33_n675 ), .A2(_AES_ENC_us33_n674 ), .A3(_AES_ENC_us33_n673 ), .A4(_AES_ENC_us33_n672 ), .ZN(_AES_ENC_us33_n676 ) );
NAND2_X2 _AES_ENC_us33_U411  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n676 ), .ZN(_AES_ENC_us33_n677 ) );
NAND2_X2 _AES_ENC_us33_U408  ( .A1(_AES_ENC_us33_n800 ), .A2(_AES_ENC_us33_n1022 ), .ZN(_AES_ENC_us33_n680 ) );
NAND2_X2 _AES_ENC_us33_U407  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n680 ), .ZN(_AES_ENC_us33_n681 ) );
AND2_X2 _AES_ENC_us33_U402  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n684 ), .ZN(_AES_ENC_us33_n682 ) );
NAND4_X2 _AES_ENC_us33_U395  ( .A1(_AES_ENC_us33_n691 ), .A2(_AES_ENC_us33_n581 ), .A3(_AES_ENC_us33_n690 ), .A4(_AES_ENC_us33_n689 ), .ZN(_AES_ENC_us33_n692 ) );
NAND2_X2 _AES_ENC_us33_U394  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n692 ), .ZN(_AES_ENC_us33_n733 ) );
NAND2_X2 _AES_ENC_us33_U392  ( .A1(_AES_ENC_us33_n977 ), .A2(_AES_ENC_us33_n1050 ), .ZN(_AES_ENC_us33_n702 ) );
NAND2_X2 _AES_ENC_us33_U391  ( .A1(_AES_ENC_us33_n1093 ), .A2(_AES_ENC_us33_n1045 ), .ZN(_AES_ENC_us33_n701 ) );
NAND4_X2 _AES_ENC_us33_U381  ( .A1(_AES_ENC_us33_n702 ), .A2(_AES_ENC_us33_n701 ), .A3(_AES_ENC_us33_n700 ), .A4(_AES_ENC_us33_n699 ), .ZN(_AES_ENC_us33_n703 ) );
NAND2_X2 _AES_ENC_us33_U380  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n703 ), .ZN(_AES_ENC_us33_n732 ) );
AND2_X2 _AES_ENC_us33_U379  ( .A1(_AES_ENC_sa33[0]), .A2(_AES_ENC_sa33[6]),.ZN(_AES_ENC_us33_n1113 ) );
NAND2_X2 _AES_ENC_us33_U378  ( .A1(_AES_ENC_us33_n601 ), .A2(_AES_ENC_us33_n1030 ), .ZN(_AES_ENC_us33_n881 ) );
NAND2_X2 _AES_ENC_us33_U377  ( .A1(_AES_ENC_us33_n1093 ), .A2(_AES_ENC_us33_n881 ), .ZN(_AES_ENC_us33_n715 ) );
NAND2_X2 _AES_ENC_us33_U376  ( .A1(_AES_ENC_us33_n1010 ), .A2(_AES_ENC_us33_n600 ), .ZN(_AES_ENC_us33_n714 ) );
NAND2_X2 _AES_ENC_us33_U375  ( .A1(_AES_ENC_us33_n855 ), .A2(_AES_ENC_us33_n588 ), .ZN(_AES_ENC_us33_n1117 ) );
XNOR2_X2 _AES_ENC_us33_U371  ( .A(_AES_ENC_us33_n611 ), .B(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n824 ) );
NAND4_X2 _AES_ENC_us33_U362  ( .A1(_AES_ENC_us33_n715 ), .A2(_AES_ENC_us33_n714 ), .A3(_AES_ENC_us33_n713 ), .A4(_AES_ENC_us33_n712 ), .ZN(_AES_ENC_us33_n716 ) );
NAND2_X2 _AES_ENC_us33_U361  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n716 ), .ZN(_AES_ENC_us33_n731 ) );
AND2_X2 _AES_ENC_us33_U360  ( .A1(_AES_ENC_sa33[6]), .A2(_AES_ENC_us33_n574 ), .ZN(_AES_ENC_us33_n1131 ) );
NAND2_X2 _AES_ENC_us33_U359  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n717 ) );
NAND2_X2 _AES_ENC_us33_U358  ( .A1(_AES_ENC_us33_n1029 ), .A2(_AES_ENC_us33_n717 ), .ZN(_AES_ENC_us33_n728 ) );
NAND2_X2 _AES_ENC_us33_U357  ( .A1(_AES_ENC_sa33[1]), .A2(_AES_ENC_us33_n624 ), .ZN(_AES_ENC_us33_n1097 ) );
NAND2_X2 _AES_ENC_us33_U356  ( .A1(_AES_ENC_us33_n603 ), .A2(_AES_ENC_us33_n1097 ), .ZN(_AES_ENC_us33_n718 ) );
NAND2_X2 _AES_ENC_us33_U355  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n718 ), .ZN(_AES_ENC_us33_n727 ) );
NAND4_X2 _AES_ENC_us33_U344  ( .A1(_AES_ENC_us33_n728 ), .A2(_AES_ENC_us33_n727 ), .A3(_AES_ENC_us33_n726 ), .A4(_AES_ENC_us33_n725 ), .ZN(_AES_ENC_us33_n729 ) );
NAND2_X2 _AES_ENC_us33_U343  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n729 ), .ZN(_AES_ENC_us33_n730 ) );
NAND4_X2 _AES_ENC_us33_U342  ( .A1(_AES_ENC_us33_n733 ), .A2(_AES_ENC_us33_n732 ), .A3(_AES_ENC_us33_n731 ), .A4(_AES_ENC_us33_n730 ), .ZN(_AES_ENC_sa33_sub[1] ) );
NAND2_X2 _AES_ENC_us33_U341  ( .A1(_AES_ENC_sa33[7]), .A2(_AES_ENC_us33_n611 ), .ZN(_AES_ENC_us33_n734 ) );
NAND2_X2 _AES_ENC_us33_U340  ( .A1(_AES_ENC_us33_n734 ), .A2(_AES_ENC_us33_n607 ), .ZN(_AES_ENC_us33_n738 ) );
OR4_X2 _AES_ENC_us33_U339  ( .A1(_AES_ENC_us33_n738 ), .A2(_AES_ENC_us33_n626 ), .A3(_AES_ENC_us33_n826 ), .A4(_AES_ENC_us33_n1121 ), .ZN(_AES_ENC_us33_n746 ) );
NAND2_X2 _AES_ENC_us33_U337  ( .A1(_AES_ENC_us33_n1100 ), .A2(_AES_ENC_us33_n587 ), .ZN(_AES_ENC_us33_n992 ) );
OR2_X2 _AES_ENC_us33_U336  ( .A1(_AES_ENC_us33_n610 ), .A2(_AES_ENC_us33_n735 ), .ZN(_AES_ENC_us33_n737 ) );
NAND2_X2 _AES_ENC_us33_U334  ( .A1(_AES_ENC_us33_n619 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n753 ) );
NAND2_X2 _AES_ENC_us33_U333  ( .A1(_AES_ENC_us33_n582 ), .A2(_AES_ENC_us33_n753 ), .ZN(_AES_ENC_us33_n1080 ) );
NAND2_X2 _AES_ENC_us33_U332  ( .A1(_AES_ENC_us33_n1048 ), .A2(_AES_ENC_us33_n576 ), .ZN(_AES_ENC_us33_n736 ) );
NAND2_X2 _AES_ENC_us33_U331  ( .A1(_AES_ENC_us33_n737 ), .A2(_AES_ENC_us33_n736 ), .ZN(_AES_ENC_us33_n739 ) );
NAND2_X2 _AES_ENC_us33_U330  ( .A1(_AES_ENC_us33_n739 ), .A2(_AES_ENC_us33_n738 ), .ZN(_AES_ENC_us33_n745 ) );
NAND2_X2 _AES_ENC_us33_U326  ( .A1(_AES_ENC_us33_n1096 ), .A2(_AES_ENC_us33_n590 ), .ZN(_AES_ENC_us33_n906 ) );
NAND4_X2 _AES_ENC_us33_U323  ( .A1(_AES_ENC_us33_n746 ), .A2(_AES_ENC_us33_n992 ), .A3(_AES_ENC_us33_n745 ), .A4(_AES_ENC_us33_n744 ), .ZN(_AES_ENC_us33_n747 ) );
NAND2_X2 _AES_ENC_us33_U322  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n747 ), .ZN(_AES_ENC_us33_n793 ) );
NAND2_X2 _AES_ENC_us33_U321  ( .A1(_AES_ENC_us33_n584 ), .A2(_AES_ENC_us33_n855 ), .ZN(_AES_ENC_us33_n748 ) );
NAND2_X2 _AES_ENC_us33_U320  ( .A1(_AES_ENC_us33_n956 ), .A2(_AES_ENC_us33_n748 ), .ZN(_AES_ENC_us33_n760 ) );
NAND2_X2 _AES_ENC_us33_U313  ( .A1(_AES_ENC_us33_n590 ), .A2(_AES_ENC_us33_n753 ), .ZN(_AES_ENC_us33_n1023 ) );
NAND4_X2 _AES_ENC_us33_U308  ( .A1(_AES_ENC_us33_n760 ), .A2(_AES_ENC_us33_n992 ), .A3(_AES_ENC_us33_n759 ), .A4(_AES_ENC_us33_n758 ), .ZN(_AES_ENC_us33_n761 ) );
NAND2_X2 _AES_ENC_us33_U307  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n761 ), .ZN(_AES_ENC_us33_n792 ) );
NAND2_X2 _AES_ENC_us33_U306  ( .A1(_AES_ENC_us33_n584 ), .A2(_AES_ENC_us33_n603 ), .ZN(_AES_ENC_us33_n989 ) );
NAND2_X2 _AES_ENC_us33_U305  ( .A1(_AES_ENC_us33_n1050 ), .A2(_AES_ENC_us33_n989 ), .ZN(_AES_ENC_us33_n777 ) );
NAND2_X2 _AES_ENC_us33_U304  ( .A1(_AES_ENC_us33_n1093 ), .A2(_AES_ENC_us33_n762 ), .ZN(_AES_ENC_us33_n776 ) );
XNOR2_X2 _AES_ENC_us33_U301  ( .A(_AES_ENC_sa33[7]), .B(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n959 ) );
NAND4_X2 _AES_ENC_us33_U289  ( .A1(_AES_ENC_us33_n777 ), .A2(_AES_ENC_us33_n776 ), .A3(_AES_ENC_us33_n775 ), .A4(_AES_ENC_us33_n774 ), .ZN(_AES_ENC_us33_n778 ) );
NAND2_X2 _AES_ENC_us33_U288  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n778 ), .ZN(_AES_ENC_us33_n791 ) );
NAND2_X2 _AES_ENC_us33_U287  ( .A1(_AES_ENC_us33_n1056 ), .A2(_AES_ENC_us33_n1050 ), .ZN(_AES_ENC_us33_n788 ) );
NAND2_X2 _AES_ENC_us33_U286  ( .A1(_AES_ENC_us33_n1091 ), .A2(_AES_ENC_us33_n779 ), .ZN(_AES_ENC_us33_n787 ) );
NAND2_X2 _AES_ENC_us33_U285  ( .A1(_AES_ENC_us33_n956 ), .A2(_AES_ENC_sa33[1]), .ZN(_AES_ENC_us33_n786 ) );
NAND4_X2 _AES_ENC_us33_U278  ( .A1(_AES_ENC_us33_n788 ), .A2(_AES_ENC_us33_n787 ), .A3(_AES_ENC_us33_n786 ), .A4(_AES_ENC_us33_n785 ), .ZN(_AES_ENC_us33_n789 ) );
NAND2_X2 _AES_ENC_us33_U277  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n789 ), .ZN(_AES_ENC_us33_n790 ) );
NAND4_X2 _AES_ENC_us33_U276  ( .A1(_AES_ENC_us33_n793 ), .A2(_AES_ENC_us33_n792 ), .A3(_AES_ENC_us33_n791 ), .A4(_AES_ENC_us33_n790 ), .ZN(_AES_ENC_sa33_sub[2] ) );
NAND2_X2 _AES_ENC_us33_U275  ( .A1(_AES_ENC_us33_n1059 ), .A2(_AES_ENC_us33_n794 ), .ZN(_AES_ENC_us33_n810 ) );
NAND2_X2 _AES_ENC_us33_U274  ( .A1(_AES_ENC_us33_n1049 ), .A2(_AES_ENC_us33_n956 ), .ZN(_AES_ENC_us33_n809 ) );
OR2_X2 _AES_ENC_us33_U266  ( .A1(_AES_ENC_us33_n1096 ), .A2(_AES_ENC_us33_n606 ), .ZN(_AES_ENC_us33_n802 ) );
NAND2_X2 _AES_ENC_us33_U265  ( .A1(_AES_ENC_us33_n1053 ), .A2(_AES_ENC_us33_n800 ), .ZN(_AES_ENC_us33_n801 ) );
NAND2_X2 _AES_ENC_us33_U264  ( .A1(_AES_ENC_us33_n802 ), .A2(_AES_ENC_us33_n801 ), .ZN(_AES_ENC_us33_n805 ) );
NAND4_X2 _AES_ENC_us33_U261  ( .A1(_AES_ENC_us33_n810 ), .A2(_AES_ENC_us33_n809 ), .A3(_AES_ENC_us33_n808 ), .A4(_AES_ENC_us33_n807 ), .ZN(_AES_ENC_us33_n811 ) );
NAND2_X2 _AES_ENC_us33_U260  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n811 ), .ZN(_AES_ENC_us33_n852 ) );
OR2_X2 _AES_ENC_us33_U259  ( .A1(_AES_ENC_us33_n1023 ), .A2(_AES_ENC_us33_n617 ), .ZN(_AES_ENC_us33_n819 ) );
OR2_X2 _AES_ENC_us33_U257  ( .A1(_AES_ENC_us33_n570 ), .A2(_AES_ENC_us33_n930 ), .ZN(_AES_ENC_us33_n818 ) );
NAND2_X2 _AES_ENC_us33_U256  ( .A1(_AES_ENC_us33_n1013 ), .A2(_AES_ENC_us33_n1094 ), .ZN(_AES_ENC_us33_n817 ) );
NAND4_X2 _AES_ENC_us33_U249  ( .A1(_AES_ENC_us33_n819 ), .A2(_AES_ENC_us33_n818 ), .A3(_AES_ENC_us33_n817 ), .A4(_AES_ENC_us33_n816 ), .ZN(_AES_ENC_us33_n820 ) );
NAND2_X2 _AES_ENC_us33_U248  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n820 ), .ZN(_AES_ENC_us33_n851 ) );
NAND2_X2 _AES_ENC_us33_U247  ( .A1(_AES_ENC_us33_n956 ), .A2(_AES_ENC_us33_n1080 ), .ZN(_AES_ENC_us33_n835 ) );
NAND2_X2 _AES_ENC_us33_U246  ( .A1(_AES_ENC_us33_n570 ), .A2(_AES_ENC_us33_n1030 ), .ZN(_AES_ENC_us33_n1047 ) );
OR2_X2 _AES_ENC_us33_U245  ( .A1(_AES_ENC_us33_n1047 ), .A2(_AES_ENC_us33_n612 ), .ZN(_AES_ENC_us33_n834 ) );
NAND2_X2 _AES_ENC_us33_U244  ( .A1(_AES_ENC_us33_n1072 ), .A2(_AES_ENC_us33_n589 ), .ZN(_AES_ENC_us33_n833 ) );
NAND4_X2 _AES_ENC_us33_U233  ( .A1(_AES_ENC_us33_n835 ), .A2(_AES_ENC_us33_n834 ), .A3(_AES_ENC_us33_n833 ), .A4(_AES_ENC_us33_n832 ), .ZN(_AES_ENC_us33_n836 ) );
NAND2_X2 _AES_ENC_us33_U232  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n836 ), .ZN(_AES_ENC_us33_n850 ) );
NAND2_X2 _AES_ENC_us33_U231  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n623 ), .ZN(_AES_ENC_us33_n847 ) );
NAND2_X2 _AES_ENC_us33_U230  ( .A1(_AES_ENC_us33_n1050 ), .A2(_AES_ENC_us33_n1071 ), .ZN(_AES_ENC_us33_n846 ) );
OR2_X2 _AES_ENC_us33_U224  ( .A1(_AES_ENC_us33_n1053 ), .A2(_AES_ENC_us33_n911 ), .ZN(_AES_ENC_us33_n1077 ) );
NAND4_X2 _AES_ENC_us33_U220  ( .A1(_AES_ENC_us33_n847 ), .A2(_AES_ENC_us33_n846 ), .A3(_AES_ENC_us33_n845 ), .A4(_AES_ENC_us33_n844 ), .ZN(_AES_ENC_us33_n848 ) );
NAND2_X2 _AES_ENC_us33_U219  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n848 ), .ZN(_AES_ENC_us33_n849 ) );
NAND4_X2 _AES_ENC_us33_U218  ( .A1(_AES_ENC_us33_n852 ), .A2(_AES_ENC_us33_n851 ), .A3(_AES_ENC_us33_n850 ), .A4(_AES_ENC_us33_n849 ), .ZN(_AES_ENC_sa33_sub[3] ) );
NAND2_X2 _AES_ENC_us33_U216  ( .A1(_AES_ENC_us33_n1009 ), .A2(_AES_ENC_us33_n1072 ), .ZN(_AES_ENC_us33_n862 ) );
NAND2_X2 _AES_ENC_us33_U215  ( .A1(_AES_ENC_us33_n603 ), .A2(_AES_ENC_us33_n577 ), .ZN(_AES_ENC_us33_n853 ) );
NAND2_X2 _AES_ENC_us33_U214  ( .A1(_AES_ENC_us33_n1050 ), .A2(_AES_ENC_us33_n853 ), .ZN(_AES_ENC_us33_n861 ) );
NAND4_X2 _AES_ENC_us33_U206  ( .A1(_AES_ENC_us33_n862 ), .A2(_AES_ENC_us33_n861 ), .A3(_AES_ENC_us33_n860 ), .A4(_AES_ENC_us33_n859 ), .ZN(_AES_ENC_us33_n863 ) );
NAND2_X2 _AES_ENC_us33_U205  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n863 ), .ZN(_AES_ENC_us33_n905 ) );
NAND2_X2 _AES_ENC_us33_U204  ( .A1(_AES_ENC_us33_n1010 ), .A2(_AES_ENC_us33_n989 ), .ZN(_AES_ENC_us33_n874 ) );
NAND2_X2 _AES_ENC_us33_U203  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n610 ), .ZN(_AES_ENC_us33_n864 ) );
NAND2_X2 _AES_ENC_us33_U202  ( .A1(_AES_ENC_us33_n929 ), .A2(_AES_ENC_us33_n864 ), .ZN(_AES_ENC_us33_n873 ) );
NAND4_X2 _AES_ENC_us33_U193  ( .A1(_AES_ENC_us33_n874 ), .A2(_AES_ENC_us33_n873 ), .A3(_AES_ENC_us33_n872 ), .A4(_AES_ENC_us33_n871 ), .ZN(_AES_ENC_us33_n875 ) );
NAND2_X2 _AES_ENC_us33_U192  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n875 ), .ZN(_AES_ENC_us33_n904 ) );
NAND2_X2 _AES_ENC_us33_U191  ( .A1(_AES_ENC_us33_n583 ), .A2(_AES_ENC_us33_n1050 ), .ZN(_AES_ENC_us33_n889 ) );
NAND2_X2 _AES_ENC_us33_U190  ( .A1(_AES_ENC_us33_n1093 ), .A2(_AES_ENC_us33_n587 ), .ZN(_AES_ENC_us33_n876 ) );
NAND2_X2 _AES_ENC_us33_U189  ( .A1(_AES_ENC_us33_n604 ), .A2(_AES_ENC_us33_n876 ), .ZN(_AES_ENC_us33_n877 ) );
NAND2_X2 _AES_ENC_us33_U188  ( .A1(_AES_ENC_us33_n877 ), .A2(_AES_ENC_us33_n623 ), .ZN(_AES_ENC_us33_n888 ) );
NAND4_X2 _AES_ENC_us33_U179  ( .A1(_AES_ENC_us33_n889 ), .A2(_AES_ENC_us33_n888 ), .A3(_AES_ENC_us33_n887 ), .A4(_AES_ENC_us33_n886 ), .ZN(_AES_ENC_us33_n890 ) );
NAND2_X2 _AES_ENC_us33_U178  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n890 ), .ZN(_AES_ENC_us33_n903 ) );
OR2_X2 _AES_ENC_us33_U177  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n1059 ), .ZN(_AES_ENC_us33_n900 ) );
NAND2_X2 _AES_ENC_us33_U176  ( .A1(_AES_ENC_us33_n1073 ), .A2(_AES_ENC_us33_n1047 ), .ZN(_AES_ENC_us33_n899 ) );
NAND2_X2 _AES_ENC_us33_U175  ( .A1(_AES_ENC_us33_n1094 ), .A2(_AES_ENC_us33_n595 ), .ZN(_AES_ENC_us33_n898 ) );
NAND4_X2 _AES_ENC_us33_U167  ( .A1(_AES_ENC_us33_n900 ), .A2(_AES_ENC_us33_n899 ), .A3(_AES_ENC_us33_n898 ), .A4(_AES_ENC_us33_n897 ), .ZN(_AES_ENC_us33_n901 ) );
NAND2_X2 _AES_ENC_us33_U166  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n901 ), .ZN(_AES_ENC_us33_n902 ) );
NAND4_X2 _AES_ENC_us33_U165  ( .A1(_AES_ENC_us33_n905 ), .A2(_AES_ENC_us33_n904 ), .A3(_AES_ENC_us33_n903 ), .A4(_AES_ENC_us33_n902 ), .ZN(_AES_ENC_sa33_sub[4] ) );
NAND2_X2 _AES_ENC_us33_U164  ( .A1(_AES_ENC_us33_n1094 ), .A2(_AES_ENC_us33_n599 ), .ZN(_AES_ENC_us33_n922 ) );
NAND2_X2 _AES_ENC_us33_U163  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n989 ), .ZN(_AES_ENC_us33_n921 ) );
NAND4_X2 _AES_ENC_us33_U151  ( .A1(_AES_ENC_us33_n922 ), .A2(_AES_ENC_us33_n921 ), .A3(_AES_ENC_us33_n920 ), .A4(_AES_ENC_us33_n919 ), .ZN(_AES_ENC_us33_n923 ) );
NAND2_X2 _AES_ENC_us33_U150  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n923 ), .ZN(_AES_ENC_us33_n972 ) );
NAND2_X2 _AES_ENC_us33_U149  ( .A1(_AES_ENC_us33_n582 ), .A2(_AES_ENC_us33_n619 ), .ZN(_AES_ENC_us33_n924 ) );
NAND2_X2 _AES_ENC_us33_U148  ( .A1(_AES_ENC_us33_n1073 ), .A2(_AES_ENC_us33_n924 ), .ZN(_AES_ENC_us33_n939 ) );
NAND2_X2 _AES_ENC_us33_U147  ( .A1(_AES_ENC_us33_n926 ), .A2(_AES_ENC_us33_n925 ), .ZN(_AES_ENC_us33_n927 ) );
NAND2_X2 _AES_ENC_us33_U146  ( .A1(_AES_ENC_us33_n606 ), .A2(_AES_ENC_us33_n927 ), .ZN(_AES_ENC_us33_n928 ) );
NAND2_X2 _AES_ENC_us33_U145  ( .A1(_AES_ENC_us33_n928 ), .A2(_AES_ENC_us33_n1080 ), .ZN(_AES_ENC_us33_n938 ) );
OR2_X2 _AES_ENC_us33_U144  ( .A1(_AES_ENC_us33_n1117 ), .A2(_AES_ENC_us33_n615 ), .ZN(_AES_ENC_us33_n937 ) );
NAND4_X2 _AES_ENC_us33_U139  ( .A1(_AES_ENC_us33_n939 ), .A2(_AES_ENC_us33_n938 ), .A3(_AES_ENC_us33_n937 ), .A4(_AES_ENC_us33_n936 ), .ZN(_AES_ENC_us33_n940 ) );
NAND2_X2 _AES_ENC_us33_U138  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n940 ), .ZN(_AES_ENC_us33_n971 ) );
OR2_X2 _AES_ENC_us33_U137  ( .A1(_AES_ENC_us33_n605 ), .A2(_AES_ENC_us33_n941 ), .ZN(_AES_ENC_us33_n954 ) );
NAND2_X2 _AES_ENC_us33_U136  ( .A1(_AES_ENC_us33_n1096 ), .A2(_AES_ENC_us33_n577 ), .ZN(_AES_ENC_us33_n942 ) );
NAND2_X2 _AES_ENC_us33_U135  ( .A1(_AES_ENC_us33_n1048 ), .A2(_AES_ENC_us33_n942 ), .ZN(_AES_ENC_us33_n943 ) );
NAND2_X2 _AES_ENC_us33_U134  ( .A1(_AES_ENC_us33_n612 ), .A2(_AES_ENC_us33_n943 ), .ZN(_AES_ENC_us33_n944 ) );
NAND2_X2 _AES_ENC_us33_U133  ( .A1(_AES_ENC_us33_n944 ), .A2(_AES_ENC_us33_n580 ), .ZN(_AES_ENC_us33_n953 ) );
NAND4_X2 _AES_ENC_us33_U125  ( .A1(_AES_ENC_us33_n954 ), .A2(_AES_ENC_us33_n953 ), .A3(_AES_ENC_us33_n952 ), .A4(_AES_ENC_us33_n951 ), .ZN(_AES_ENC_us33_n955 ) );
NAND2_X2 _AES_ENC_us33_U124  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n955 ), .ZN(_AES_ENC_us33_n970 ) );
NAND2_X2 _AES_ENC_us33_U123  ( .A1(_AES_ENC_us33_n1094 ), .A2(_AES_ENC_us33_n1071 ), .ZN(_AES_ENC_us33_n967 ) );
NAND2_X2 _AES_ENC_us33_U122  ( .A1(_AES_ENC_us33_n956 ), .A2(_AES_ENC_us33_n1030 ), .ZN(_AES_ENC_us33_n966 ) );
NAND4_X2 _AES_ENC_us33_U114  ( .A1(_AES_ENC_us33_n967 ), .A2(_AES_ENC_us33_n966 ), .A3(_AES_ENC_us33_n965 ), .A4(_AES_ENC_us33_n964 ), .ZN(_AES_ENC_us33_n968 ) );
NAND2_X2 _AES_ENC_us33_U113  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n968 ), .ZN(_AES_ENC_us33_n969 ) );
NAND4_X2 _AES_ENC_us33_U112  ( .A1(_AES_ENC_us33_n972 ), .A2(_AES_ENC_us33_n971 ), .A3(_AES_ENC_us33_n970 ), .A4(_AES_ENC_us33_n969 ), .ZN(_AES_ENC_sa33_sub[5] ) );
NAND2_X2 _AES_ENC_us33_U111  ( .A1(_AES_ENC_us33_n570 ), .A2(_AES_ENC_us33_n1097 ), .ZN(_AES_ENC_us33_n973 ) );
NAND2_X2 _AES_ENC_us33_U110  ( .A1(_AES_ENC_us33_n1073 ), .A2(_AES_ENC_us33_n973 ), .ZN(_AES_ENC_us33_n987 ) );
NAND2_X2 _AES_ENC_us33_U109  ( .A1(_AES_ENC_us33_n974 ), .A2(_AES_ENC_us33_n1077 ), .ZN(_AES_ENC_us33_n975 ) );
NAND2_X2 _AES_ENC_us33_U108  ( .A1(_AES_ENC_us33_n613 ), .A2(_AES_ENC_us33_n975 ), .ZN(_AES_ENC_us33_n976 ) );
NAND2_X2 _AES_ENC_us33_U107  ( .A1(_AES_ENC_us33_n977 ), .A2(_AES_ENC_us33_n976 ), .ZN(_AES_ENC_us33_n986 ) );
NAND4_X2 _AES_ENC_us33_U99  ( .A1(_AES_ENC_us33_n987 ), .A2(_AES_ENC_us33_n986 ), .A3(_AES_ENC_us33_n985 ), .A4(_AES_ENC_us33_n984 ), .ZN(_AES_ENC_us33_n988 ) );
NAND2_X2 _AES_ENC_us33_U98  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n988 ), .ZN(_AES_ENC_us33_n1044 ) );
NAND2_X2 _AES_ENC_us33_U97  ( .A1(_AES_ENC_us33_n1073 ), .A2(_AES_ENC_us33_n989 ), .ZN(_AES_ENC_us33_n1004 ) );
NAND2_X2 _AES_ENC_us33_U96  ( .A1(_AES_ENC_us33_n1092 ), .A2(_AES_ENC_us33_n619 ), .ZN(_AES_ENC_us33_n1003 ) );
NAND4_X2 _AES_ENC_us33_U85  ( .A1(_AES_ENC_us33_n1004 ), .A2(_AES_ENC_us33_n1003 ), .A3(_AES_ENC_us33_n1002 ), .A4(_AES_ENC_us33_n1001 ), .ZN(_AES_ENC_us33_n1005 ) );
NAND2_X2 _AES_ENC_us33_U84  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n1005 ), .ZN(_AES_ENC_us33_n1043 ) );
NAND2_X2 _AES_ENC_us33_U83  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n596 ), .ZN(_AES_ENC_us33_n1020 ) );
NAND2_X2 _AES_ENC_us33_U82  ( .A1(_AES_ENC_us33_n1050 ), .A2(_AES_ENC_us33_n624 ), .ZN(_AES_ENC_us33_n1019 ) );
NAND2_X2 _AES_ENC_us33_U77  ( .A1(_AES_ENC_us33_n1059 ), .A2(_AES_ENC_us33_n1114 ), .ZN(_AES_ENC_us33_n1012 ) );
NAND2_X2 _AES_ENC_us33_U76  ( .A1(_AES_ENC_us33_n1010 ), .A2(_AES_ENC_us33_n592 ), .ZN(_AES_ENC_us33_n1011 ) );
NAND2_X2 _AES_ENC_us33_U75  ( .A1(_AES_ENC_us33_n1012 ), .A2(_AES_ENC_us33_n1011 ), .ZN(_AES_ENC_us33_n1016 ) );
NAND4_X2 _AES_ENC_us33_U70  ( .A1(_AES_ENC_us33_n1020 ), .A2(_AES_ENC_us33_n1019 ), .A3(_AES_ENC_us33_n1018 ), .A4(_AES_ENC_us33_n1017 ), .ZN(_AES_ENC_us33_n1021 ) );
NAND2_X2 _AES_ENC_us33_U69  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n1021 ), .ZN(_AES_ENC_us33_n1042 ) );
NAND2_X2 _AES_ENC_us33_U68  ( .A1(_AES_ENC_us33_n1022 ), .A2(_AES_ENC_us33_n1093 ), .ZN(_AES_ENC_us33_n1039 ) );
NAND2_X2 _AES_ENC_us33_U67  ( .A1(_AES_ENC_us33_n1050 ), .A2(_AES_ENC_us33_n1023 ), .ZN(_AES_ENC_us33_n1038 ) );
NAND2_X2 _AES_ENC_us33_U66  ( .A1(_AES_ENC_us33_n1024 ), .A2(_AES_ENC_us33_n1071 ), .ZN(_AES_ENC_us33_n1037 ) );
AND2_X2 _AES_ENC_us33_U60  ( .A1(_AES_ENC_us33_n1030 ), .A2(_AES_ENC_us33_n602 ), .ZN(_AES_ENC_us33_n1078 ) );
NAND4_X2 _AES_ENC_us33_U56  ( .A1(_AES_ENC_us33_n1039 ), .A2(_AES_ENC_us33_n1038 ), .A3(_AES_ENC_us33_n1037 ), .A4(_AES_ENC_us33_n1036 ), .ZN(_AES_ENC_us33_n1040 ) );
NAND2_X2 _AES_ENC_us33_U55  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n1040 ), .ZN(_AES_ENC_us33_n1041 ) );
NAND4_X2 _AES_ENC_us33_U54  ( .A1(_AES_ENC_us33_n1044 ), .A2(_AES_ENC_us33_n1043 ), .A3(_AES_ENC_us33_n1042 ), .A4(_AES_ENC_us33_n1041 ), .ZN(_AES_ENC_sa33_sub[6] ) );
NAND2_X2 _AES_ENC_us33_U53  ( .A1(_AES_ENC_us33_n1072 ), .A2(_AES_ENC_us33_n1045 ), .ZN(_AES_ENC_us33_n1068 ) );
NAND2_X2 _AES_ENC_us33_U52  ( .A1(_AES_ENC_us33_n1046 ), .A2(_AES_ENC_us33_n582 ), .ZN(_AES_ENC_us33_n1067 ) );
NAND2_X2 _AES_ENC_us33_U51  ( .A1(_AES_ENC_us33_n1094 ), .A2(_AES_ENC_us33_n1047 ), .ZN(_AES_ENC_us33_n1066 ) );
NAND4_X2 _AES_ENC_us33_U40  ( .A1(_AES_ENC_us33_n1068 ), .A2(_AES_ENC_us33_n1067 ), .A3(_AES_ENC_us33_n1066 ), .A4(_AES_ENC_us33_n1065 ), .ZN(_AES_ENC_us33_n1069 ) );
NAND2_X2 _AES_ENC_us33_U39  ( .A1(_AES_ENC_us33_n1070 ), .A2(_AES_ENC_us33_n1069 ), .ZN(_AES_ENC_us33_n1135 ) );
NAND2_X2 _AES_ENC_us33_U38  ( .A1(_AES_ENC_us33_n1072 ), .A2(_AES_ENC_us33_n1071 ), .ZN(_AES_ENC_us33_n1088 ) );
NAND2_X2 _AES_ENC_us33_U37  ( .A1(_AES_ENC_us33_n1073 ), .A2(_AES_ENC_us33_n595 ), .ZN(_AES_ENC_us33_n1087 ) );
NAND4_X2 _AES_ENC_us33_U28  ( .A1(_AES_ENC_us33_n1088 ), .A2(_AES_ENC_us33_n1087 ), .A3(_AES_ENC_us33_n1086 ), .A4(_AES_ENC_us33_n1085 ), .ZN(_AES_ENC_us33_n1089 ) );
NAND2_X2 _AES_ENC_us33_U27  ( .A1(_AES_ENC_us33_n1090 ), .A2(_AES_ENC_us33_n1089 ), .ZN(_AES_ENC_us33_n1134 ) );
NAND2_X2 _AES_ENC_us33_U26  ( .A1(_AES_ENC_us33_n1091 ), .A2(_AES_ENC_us33_n1093 ), .ZN(_AES_ENC_us33_n1111 ) );
NAND2_X2 _AES_ENC_us33_U25  ( .A1(_AES_ENC_us33_n1092 ), .A2(_AES_ENC_us33_n1120 ), .ZN(_AES_ENC_us33_n1110 ) );
AND2_X2 _AES_ENC_us33_U22  ( .A1(_AES_ENC_us33_n1097 ), .A2(_AES_ENC_us33_n1096 ), .ZN(_AES_ENC_us33_n1098 ) );
NAND4_X2 _AES_ENC_us33_U14  ( .A1(_AES_ENC_us33_n1111 ), .A2(_AES_ENC_us33_n1110 ), .A3(_AES_ENC_us33_n1109 ), .A4(_AES_ENC_us33_n1108 ), .ZN(_AES_ENC_us33_n1112 ) );
NAND2_X2 _AES_ENC_us33_U13  ( .A1(_AES_ENC_us33_n1113 ), .A2(_AES_ENC_us33_n1112 ), .ZN(_AES_ENC_us33_n1133 ) );
NAND2_X2 _AES_ENC_us33_U12  ( .A1(_AES_ENC_us33_n1115 ), .A2(_AES_ENC_us33_n1114 ), .ZN(_AES_ENC_us33_n1129 ) );
OR2_X2 _AES_ENC_us33_U11  ( .A1(_AES_ENC_us33_n608 ), .A2(_AES_ENC_us33_n1116 ), .ZN(_AES_ENC_us33_n1128 ) );
NAND4_X2 _AES_ENC_us33_U3  ( .A1(_AES_ENC_us33_n1129 ), .A2(_AES_ENC_us33_n1128 ), .A3(_AES_ENC_us33_n1127 ), .A4(_AES_ENC_us33_n1126 ), .ZN(_AES_ENC_us33_n1130 ) );
NAND2_X2 _AES_ENC_us33_U2  ( .A1(_AES_ENC_us33_n1131 ), .A2(_AES_ENC_us33_n1130 ), .ZN(_AES_ENC_us33_n1132 ) );
NAND4_X2 _AES_ENC_us33_U1  ( .A1(_AES_ENC_us33_n1135 ), .A2(_AES_ENC_us33_n1134 ), .A3(_AES_ENC_us33_n1133 ), .A4(_AES_ENC_us33_n1132 ), .ZN(_AES_ENC_sa33_sub[7] ) );
INV_X4 _add_506_U775  ( .A(n18589), .ZN(N2027) );
NAND2_X2 _add_506_U774  ( .A1(n18233), .A2(n18237), .ZN(_add_506_n646 ) );
NAND2_X2 _add_506_U773  ( .A1(n18225), .A2(n18229), .ZN(_add_506_n647 ) );
NAND2_X2 _add_506_U772  ( .A1(n18249), .A2(n18253), .ZN(_add_506_n644 ) );
NAND2_X2 _add_506_U771  ( .A1(n18241), .A2(n18245), .ZN(_add_506_n645 ) );
NAND4_X2 _add_506_U770  ( .A1(n18273), .A2(n18277), .A3(n18281), .A4(n18285),.ZN(_add_506_n642 ) );
NAND4_X2 _add_506_U769  ( .A1(n18257), .A2(n18261), .A3(n18265), .A4(n18269),.ZN(_add_506_n643 ) );
INV_X4 _add_506_U768  ( .A(_add_506_n37 ), .ZN(_add_506_n63 ) );
NAND4_X2 _add_506_U767  ( .A1(n18301), .A2(n18305), .A3(n18309), .A4(n18313),.ZN(_add_506_n637 ) );
NAND4_X2 _add_506_U766  ( .A1(n18329), .A2(n18333), .A3(n18337), .A4(n18341),.ZN(_add_506_n635 ) );
NAND4_X2 _add_506_U765  ( .A1(n18357), .A2(n18361), .A3(n18365), .A4(n18369),.ZN(_add_506_n633 ) );
NAND4_X2 _add_506_U764  ( .A1(n18385), .A2(n18389), .A3(n18393), .A4(n18397),.ZN(_add_506_n631 ) );
NAND2_X2 _add_506_U763  ( .A1(n18409), .A2(n18413), .ZN(_add_506_n625 ) );
NAND2_X2 _add_506_U762  ( .A1(n18401), .A2(n18405), .ZN(_add_506_n626 ) );
NAND2_X2 _add_506_U761  ( .A1(n18425), .A2(n18429), .ZN(_add_506_n623 ) );
NAND2_X2 _add_506_U760  ( .A1(n18417), .A2(n18421), .ZN(_add_506_n624 ) );
NAND4_X2 _add_506_U759  ( .A1(n18449), .A2(n18453), .A3(n18457), .A4(n18461),.ZN(_add_506_n621 ) );
NAND4_X2 _add_506_U758  ( .A1(n18433), .A2(n18437), .A3(n18441), .A4(n18445),.ZN(_add_506_n622 ) );
INV_X4 _add_506_U757  ( .A(n18197), .ZN(_add_506_n617 ) );
INV_X4 _add_506_U756  ( .A(n18193), .ZN(_add_506_n31 ) );
INV_X4 _add_506_U755  ( .A(n18205), .ZN(_add_506_n39 ) );
INV_X4 _add_506_U754  ( .A(n18201), .ZN(_add_506_n616 ) );
NAND2_X2 _add_506_U753  ( .A1(n18217), .A2(n18221), .ZN(_add_506_n614 ) );
NAND2_X2 _add_506_U752  ( .A1(n18209), .A2(n18213), .ZN(_add_506_n615 ) );
NAND4_X2 _add_506_U751  ( .A1(n18481), .A2(n18485), .A3(n18489), .A4(n18493),.ZN(_add_506_n609 ) );
NAND4_X2 _add_506_U750  ( .A1(n18465), .A2(n18469), .A3(n18473), .A4(n18477),.ZN(_add_506_n610 ) );
NAND4_X2 _add_506_U749  ( .A1(n18513), .A2(n18517), .A3(n18521), .A4(n18525),.ZN(_add_506_n607 ) );
NAND4_X2 _add_506_U748  ( .A1(n18497), .A2(n18501), .A3(n18505), .A4(n18509),.ZN(_add_506_n608 ) );
NAND2_X2 _add_506_U747  ( .A1(n18569), .A2(n18573), .ZN(_add_506_n605 ) );
NAND2_X2 _add_506_U746  ( .A1(n18561), .A2(n18565), .ZN(_add_506_n606 ) );
NAND2_X2 _add_506_U745  ( .A1(n18585), .A2(n18589), .ZN(_add_506_n603 ) );
NAND2_X2 _add_506_U744  ( .A1(n18577), .A2(n18581), .ZN(_add_506_n604 ) );
NAND2_X2 _add_506_U743  ( .A1(_add_506_n601 ), .A2(_add_506_n602 ), .ZN(_add_506_n598 ) );
NAND4_X2 _add_506_U742  ( .A1(n18545), .A2(n18549), .A3(n18553), .A4(n18557),.ZN(_add_506_n599 ) );
NAND4_X2 _add_506_U741  ( .A1(n18529), .A2(n18533), .A3(n18537), .A4(n18541),.ZN(_add_506_n600 ) );
NAND4_X2 _add_506_U740  ( .A1(_add_506_n63 ), .A2(_add_506_n20 ), .A3(_add_506_n594 ), .A4(_add_506_n15 ), .ZN(_add_506_n593 ) );
XNOR2_X2 _add_506_U739  ( .A(_add_506_n593 ), .B(n18189), .ZN(N2127) );
INV_X4 _add_506_U738  ( .A(_add_506_n584 ), .ZN(_add_506_n592 ) );
NAND2_X2 _add_506_U737  ( .A1(n18189), .A2(_add_506_n592 ), .ZN(_add_506_n591 ) );
NAND4_X2 _add_506_U736  ( .A1(_add_506_n63 ), .A2(_add_506_n20 ), .A3(_add_506_n590 ), .A4(_add_506_n15 ), .ZN(_add_506_n589 ) );
XNOR2_X2 _add_506_U735  ( .A(_add_506_n589 ), .B(n18185), .ZN(N2128) );
NAND2_X2 _add_506_U734  ( .A1(n18185), .A2(n18189), .ZN(_add_506_n588 ) );
NAND4_X2 _add_506_U733  ( .A1(_add_506_n63 ), .A2(_add_506_n16 ), .A3(_add_506_n587 ), .A4(_add_506_n19 ), .ZN(_add_506_n586 ) );
XNOR2_X2 _add_506_U732  ( .A(_add_506_n586 ), .B(n18181), .ZN(N2129) );
NAND4_X2 _add_506_U731  ( .A1(_add_506_n63 ), .A2(_add_506_n17 ), .A3(_add_506_n583 ), .A4(_add_506_n19 ), .ZN(_add_506_n582 ) );
XNOR2_X2 _add_506_U730  ( .A(_add_506_n582 ), .B(n18177), .ZN(N2130) );
NAND2_X2 _add_506_U729  ( .A1(n18217), .A2(n18221), .ZN(_add_506_n580 ) );
NAND2_X2 _add_506_U728  ( .A1(n18209), .A2(n18213), .ZN(_add_506_n581 ) );
NAND4_X2 _add_506_U727  ( .A1(n18193), .A2(n18197), .A3(n18201), .A4(n18205),.ZN(_add_506_n578 ) );
NAND4_X2 _add_506_U726  ( .A1(n18177), .A2(n18181), .A3(n18185), .A4(n18189),.ZN(_add_506_n579 ) );
NAND4_X2 _add_506_U725  ( .A1(_add_506_n576 ), .A2(_add_506_n20 ), .A3(_add_506_n16 ), .A4(_add_506_n577 ), .ZN(_add_506_n575 ) );
XNOR2_X2 _add_506_U724  ( .A(_add_506_n575 ), .B(n18173), .ZN(N2131) );
NAND4_X2 _add_506_U723  ( .A1(n18209), .A2(n18221), .A3(n18217), .A4(n18213),.ZN(_add_506_n572 ) );
NAND4_X2 _add_506_U722  ( .A1(n18189), .A2(n18193), .A3(n18197), .A4(n18201),.ZN(_add_506_n573 ) );
NAND4_X2 _add_506_U721  ( .A1(n18173), .A2(n18177), .A3(n18181), .A4(n18185),.ZN(_add_506_n574 ) );
NAND4_X2 _add_506_U720  ( .A1(_add_506_n19 ), .A2(_add_506_n570 ), .A3(_add_506_n16 ), .A4(_add_506_n571 ), .ZN(_add_506_n569 ) );
XNOR2_X2 _add_506_U719  ( .A(_add_506_n569 ), .B(n18169), .ZN(N2132) );
INV_X4 _add_506_U718  ( .A(n18173), .ZN(_add_506_n555 ) );
INV_X4 _add_506_U717  ( .A(n18169), .ZN(_add_506_n556 ) );
INV_X4 _add_506_U716  ( .A(n18181), .ZN(_add_506_n553 ) );
INV_X4 _add_506_U715  ( .A(n18177), .ZN(_add_506_n554 ) );
INV_X4 _add_506_U714  ( .A(n18189), .ZN(_add_506_n568 ) );
INV_X4 _add_506_U713  ( .A(n18185), .ZN(_add_506_n552 ) );
NAND3_X2 _add_506_U712  ( .A1(_add_506_n565 ), .A2(_add_506_n566 ), .A3(_add_506_n567 ), .ZN(_add_506_n562 ) );
NAND4_X2 _add_506_U711  ( .A1(n18209), .A2(n18221), .A3(n18217), .A4(n18213),.ZN(_add_506_n563 ) );
NAND4_X2 _add_506_U710  ( .A1(_add_506_n19 ), .A2(_add_506_n560 ), .A3(_add_506_n16 ), .A4(_add_506_n561 ), .ZN(_add_506_n559 ) );
XNOR2_X2 _add_506_U709  ( .A(_add_506_n559 ), .B(n18165), .ZN(N2133) );
NAND2_X2 _add_506_U708  ( .A1(n18201), .A2(n18205), .ZN(_add_506_n558 ) );
INV_X4 _add_506_U707  ( .A(n18165), .ZN(_add_506_n557 ) );
NAND3_X2 _add_506_U706  ( .A1(_add_506_n549 ), .A2(_add_506_n550 ), .A3(_add_506_n551 ), .ZN(_add_506_n546 ) );
NAND4_X2 _add_506_U705  ( .A1(n18209), .A2(n18221), .A3(n18217), .A4(n18213),.ZN(_add_506_n547 ) );
NAND4_X2 _add_506_U704  ( .A1(_add_506_n20 ), .A2(_add_506_n544 ), .A3(_add_506_n16 ), .A4(_add_506_n545 ), .ZN(_add_506_n543 ) );
XNOR2_X2 _add_506_U703  ( .A(_add_506_n543 ), .B(n18161), .ZN(N2134) );
NAND4_X2 _add_506_U702  ( .A1(n18177), .A2(n18181), .A3(n18185), .A4(n18189),.ZN(_add_506_n541 ) );
NAND4_X2 _add_506_U701  ( .A1(n18161), .A2(n18165), .A3(n18169), .A4(n18173),.ZN(_add_506_n542 ) );
NAND4_X2 _add_506_U700  ( .A1(n18209), .A2(n18213), .A3(n18217), .A4(n18221),.ZN(_add_506_n539 ) );
NAND4_X2 _add_506_U699  ( .A1(n18193), .A2(n18197), .A3(n18201), .A4(n18205),.ZN(_add_506_n540 ) );
NAND2_X2 _add_506_U698  ( .A1(n18265), .A2(n18269), .ZN(_add_506_n537 ) );
NAND2_X2 _add_506_U697  ( .A1(n18257), .A2(n18261), .ZN(_add_506_n538 ) );
NAND2_X2 _add_506_U696  ( .A1(n18281), .A2(n18285), .ZN(_add_506_n535 ) );
NAND2_X2 _add_506_U695  ( .A1(n18273), .A2(n18277), .ZN(_add_506_n536 ) );
NAND2_X2 _add_506_U694  ( .A1(_add_506_n533 ), .A2(_add_506_n534 ), .ZN(_add_506_n530 ) );
NAND4_X2 _add_506_U693  ( .A1(n18241), .A2(n18245), .A3(n18249), .A4(n18253),.ZN(_add_506_n531 ) );
NAND4_X2 _add_506_U692  ( .A1(n18225), .A2(n18229), .A3(n18233), .A4(n18237),.ZN(_add_506_n532 ) );
NAND4_X2 _add_506_U691  ( .A1(_add_506_n398 ), .A2(_add_506_n27 ), .A3(_add_506_n19 ), .A4(_add_506_n15 ), .ZN(_add_506_n526 ) );
XNOR2_X2 _add_506_U690  ( .A(_add_506_n526 ), .B(n18157), .ZN(N2135) );
INV_X4 _add_506_U689  ( .A(n18153), .ZN(_add_506_n427 ) );
NAND3_X2 _add_506_U688  ( .A1(n18157), .A2(_add_506_n398 ), .A3(_add_506_n17 ), .ZN(_add_506_n524 ) );
NAND2_X2 _add_506_U687  ( .A1(_add_506_n22 ), .A2(_add_506_n28 ), .ZN(_add_506_n525 ) );
XNOR2_X2 _add_506_U686  ( .A(_add_506_n427 ), .B(_add_506_n523 ), .ZN(N2136));
NAND2_X2 _add_506_U685  ( .A1(n18565), .A2(n18561), .ZN(_add_506_n520 ) );
NAND4_X2 _add_506_U684  ( .A1(n18577), .A2(n18581), .A3(n18585), .A4(n18589),.ZN(_add_506_n521 ) );
NAND2_X2 _add_506_U683  ( .A1(n18569), .A2(n18573), .ZN(_add_506_n522 ) );
NAND2_X2 _add_506_U682  ( .A1(_add_506_n3 ), .A2(_add_506_n30 ), .ZN(_add_506_n519 ) );
XNOR2_X2 _add_506_U681  ( .A(_add_506_n519 ), .B(n18549), .ZN(N2037) );
NAND3_X2 _add_506_U680  ( .A1(_add_506_n518 ), .A2(_add_506_n398 ), .A3(_add_506_n17 ), .ZN(_add_506_n516 ) );
NAND2_X2 _add_506_U679  ( .A1(_add_506_n22 ), .A2(_add_506_n28 ), .ZN(_add_506_n517 ) );
NAND4_X2 _add_506_U678  ( .A1(_add_506_n20 ), .A2(_add_506_n16 ), .A3(_add_506_n514 ), .A4(_add_506_n398 ), .ZN(_add_506_n513 ) );
XNOR2_X2 _add_506_U677  ( .A(_add_506_n513 ), .B(n18145), .ZN(N2138) );
INV_X4 _add_506_U676  ( .A(n18141), .ZN(_add_506_n493 ) );
NAND4_X2 _add_506_U675  ( .A1(n18145), .A2(n18149), .A3(n18153), .A4(n18157),.ZN(_add_506_n505 ) );
INV_X4 _add_506_U674  ( .A(_add_506_n505 ), .ZN(_add_506_n500 ) );
NAND3_X2 _add_506_U673  ( .A1(_add_506_n500 ), .A2(_add_506_n398 ), .A3(_add_506_n17 ), .ZN(_add_506_n511 ) );
NAND2_X2 _add_506_U672  ( .A1(_add_506_n22 ), .A2(_add_506_n28 ), .ZN(_add_506_n512 ) );
XNOR2_X2 _add_506_U671  ( .A(_add_506_n493 ), .B(_add_506_n510 ), .ZN(N2139));
INV_X4 _add_506_U670  ( .A(n18137), .ZN(_add_506_n494 ) );
NAND3_X2 _add_506_U669  ( .A1(_add_506_n509 ), .A2(_add_506_n398 ), .A3(_add_506_n17 ), .ZN(_add_506_n507 ) );
NAND2_X2 _add_506_U668  ( .A1(_add_506_n22 ), .A2(_add_506_n28 ), .ZN(_add_506_n508 ) );
XNOR2_X2 _add_506_U667  ( .A(_add_506_n494 ), .B(_add_506_n506 ), .ZN(N2140));
NAND4_X2 _add_506_U666  ( .A1(_add_506_n503 ), .A2(_add_506_n27 ), .A3(_add_506_n398 ), .A4(_add_506_n504 ), .ZN(_add_506_n502 ) );
XNOR2_X2 _add_506_U665  ( .A(_add_506_n502 ), .B(n18133), .ZN(N2141) );
NAND2_X2 _add_506_U664  ( .A1(n18137), .A2(n18133), .ZN(_add_506_n501 ) );
NAND2_X2 _add_506_U663  ( .A1(_add_506_n499 ), .A2(_add_506_n500 ), .ZN(_add_506_n498 ) );
NAND4_X2 _add_506_U662  ( .A1(_add_506_n20 ), .A2(_add_506_n16 ), .A3(_add_506_n497 ), .A4(_add_506_n398 ), .ZN(_add_506_n496 ) );
XNOR2_X2 _add_506_U661  ( .A(_add_506_n496 ), .B(n18129), .ZN(N2142) );
INV_X4 _add_506_U660  ( .A(n18125), .ZN(_add_506_n465 ) );
INV_X4 _add_506_U659  ( .A(n18133), .ZN(_add_506_n495 ) );
NAND2_X2 _add_506_U658  ( .A1(n18153), .A2(n18157), .ZN(_add_506_n491 ) );
NAND2_X2 _add_506_U657  ( .A1(n18145), .A2(n18149), .ZN(_add_506_n492 ) );
INV_X4 _add_506_U656  ( .A(_add_506_n474 ), .ZN(_add_506_n481 ) );
NAND3_X2 _add_506_U655  ( .A1(_add_506_n481 ), .A2(_add_506_n398 ), .A3(_add_506_n17 ), .ZN(_add_506_n486 ) );
NAND2_X2 _add_506_U654  ( .A1(_add_506_n22 ), .A2(_add_506_n27 ), .ZN(_add_506_n487 ) );
XNOR2_X2 _add_506_U653  ( .A(_add_506_n465 ), .B(_add_506_n485 ), .ZN(N2143));
INV_X4 _add_506_U652  ( .A(n18121), .ZN(_add_506_n475 ) );
NAND4_X2 _add_506_U651  ( .A1(_add_506_n398 ), .A2(_add_506_n16 ), .A3(_add_506_n481 ), .A4(n18125), .ZN(_add_506_n483 ) );
NAND2_X2 _add_506_U650  ( .A1(_add_506_n22 ), .A2(_add_506_n27 ), .ZN(_add_506_n484 ) );
XNOR2_X2 _add_506_U649  ( .A(_add_506_n475 ), .B(_add_506_n482 ), .ZN(N2144));
INV_X4 _add_506_U648  ( .A(n18117), .ZN(_add_506_n473 ) );
AND2_X2 _add_506_U647  ( .A1(_add_506_n481 ), .A2(n18121), .ZN(_add_506_n480 ) );
NAND3_X2 _add_506_U646  ( .A1(_add_506_n480 ), .A2(_add_506_n398 ), .A3(_add_506_n17 ), .ZN(_add_506_n477 ) );
NAND2_X2 _add_506_U645  ( .A1(_add_506_n21 ), .A2(_add_506_n479 ), .ZN(_add_506_n478 ) );
XNOR2_X2 _add_506_U644  ( .A(_add_506_n473 ), .B(_add_506_n476 ), .ZN(N2145));
NAND4_X2 _add_506_U643  ( .A1(_add_506_n398 ), .A2(_add_506_n16 ), .A3(_add_506_n471 ), .A4(_add_506_n472 ), .ZN(_add_506_n470 ) );
XNOR2_X2 _add_506_U642  ( .A(_add_506_n470 ), .B(n18113), .ZN(N2146) );
XNOR2_X2 _add_506_U641  ( .A(_add_506_n469 ), .B(n18545), .ZN(N2038) );
NAND4_X2 _add_506_U640  ( .A1(n18145), .A2(n18149), .A3(n18153), .A4(n18157),.ZN(_add_506_n466 ) );
NAND4_X2 _add_506_U639  ( .A1(n18129), .A2(n18133), .A3(n18137), .A4(n18141),.ZN(_add_506_n467 ) );
NAND2_X2 _add_506_U638  ( .A1(_add_506_n27 ), .A2(_add_506_n464 ), .ZN(_add_506_n463 ) );
NAND3_X2 _add_506_U637  ( .A1(_add_506_n17 ), .A2(_add_506_n461 ), .A3(_add_506_n462 ), .ZN(_add_506_n460 ) );
XNOR2_X2 _add_506_U636  ( .A(_add_506_n460 ), .B(n18109), .ZN(N2147) );
NAND2_X2 _add_506_U635  ( .A1(n18137), .A2(n18145), .ZN(_add_506_n459 ) );
NAND4_X2 _add_506_U634  ( .A1(_add_506_n20 ), .A2(_add_506_n454 ), .A3(_add_506_n455 ), .A4(_add_506_n456 ), .ZN(_add_506_n453 ) );
XNOR2_X2 _add_506_U633  ( .A(n18105), .B(_add_506_n453 ), .ZN(N2148) );
NAND2_X2 _add_506_U632  ( .A1(n18157), .A2(n18153), .ZN(_add_506_n452 ) );
NAND4_X2 _add_506_U631  ( .A1(n18129), .A2(n18133), .A3(n18145), .A4(n18149),.ZN(_add_506_n449 ) );
NAND2_X2 _add_506_U630  ( .A1(n18137), .A2(n18141), .ZN(_add_506_n450 ) );
NOR2_X2 _add_506_U629  ( .A1(_add_506_n449 ), .A2(_add_506_n450 ), .ZN(_add_506_n448 ) );
INV_X4 _add_506_U628  ( .A(_add_506_n8 ), .ZN(_add_506_n436 ) );
NAND2_X2 _add_506_U627  ( .A1(_add_506_n448 ), .A2(_add_506_n436 ), .ZN(_add_506_n447 ) );
INV_X4 _add_506_U626  ( .A(n18105), .ZN(_add_506_n434 ) );
NAND2_X2 _add_506_U625  ( .A1(_add_506_n27 ), .A2(_add_506_n446 ), .ZN(_add_506_n445 ) );
NAND3_X2 _add_506_U624  ( .A1(_add_506_n17 ), .A2(_add_506_n443 ), .A3(_add_506_n444 ), .ZN(_add_506_n442 ) );
XNOR2_X2 _add_506_U623  ( .A(_add_506_n442 ), .B(n18101), .ZN(N2149) );
NAND2_X2 _add_506_U622  ( .A1(n18153), .A2(n18101), .ZN(_add_506_n441 ) );
NAND2_X2 _add_506_U621  ( .A1(_add_506_n398 ), .A2(_add_506_n440 ), .ZN(_add_506_n439 ) );
NAND4_X2 _add_506_U620  ( .A1(n18129), .A2(n18133), .A3(n18145), .A4(n18149),.ZN(_add_506_n437 ) );
NAND2_X2 _add_506_U619  ( .A1(n18137), .A2(n18141), .ZN(_add_506_n438 ) );
NOR2_X2 _add_506_U618  ( .A1(_add_506_n437 ), .A2(_add_506_n438 ), .ZN(_add_506_n435 ) );
NAND2_X2 _add_506_U617  ( .A1(_add_506_n435 ), .A2(_add_506_n436 ), .ZN(_add_506_n433 ) );
NAND2_X2 _add_506_U616  ( .A1(_add_506_n27 ), .A2(_add_506_n432 ), .ZN(_add_506_n431 ) );
NAND2_X2 _add_506_U615  ( .A1(_add_506_n429 ), .A2(_add_506_n430 ), .ZN(_add_506_n428 ) );
XNOR2_X2 _add_506_U614  ( .A(_add_506_n428 ), .B(n18097), .ZN(N2150) );
NAND2_X2 _add_506_U613  ( .A1(_add_506_n426 ), .A2(_add_506_n398 ), .ZN(_add_506_n425 ) );
NAND2_X2 _add_506_U612  ( .A1(n18101), .A2(n18097), .ZN(_add_506_n422 ) );
NAND4_X2 _add_506_U611  ( .A1(n18113), .A2(n18117), .A3(n18121), .A4(n18125),.ZN(_add_506_n423 ) );
NAND2_X2 _add_506_U610  ( .A1(n18105), .A2(n18109), .ZN(_add_506_n424 ) );
NAND2_X2 _add_506_U609  ( .A1(_add_506_n401 ), .A2(_add_506_n419 ), .ZN(_add_506_n418 ) );
NAND2_X2 _add_506_U608  ( .A1(_add_506_n416 ), .A2(_add_506_n417 ), .ZN(_add_506_n415 ) );
XNOR2_X2 _add_506_U607  ( .A(_add_506_n415 ), .B(n18093), .ZN(N2151) );
INV_X4 _add_506_U606  ( .A(_add_506_n401 ), .ZN(_add_506_n412 ) );
NAND4_X2 _add_506_U605  ( .A1(n18137), .A2(n18141), .A3(n18145), .A4(n18149),.ZN(_add_506_n413 ) );
NAND4_X2 _add_506_U604  ( .A1(_add_506_n409 ), .A2(_add_506_n22 ), .A3(_add_506_n26 ), .A4(_add_506_n410 ), .ZN(_add_506_n408 ) );
XNOR2_X2 _add_506_U603  ( .A(_add_506_n408 ), .B(n18089), .ZN(N2152) );
NAND4_X2 _add_506_U602  ( .A1(n18133), .A2(n18137), .A3(n18141), .A4(n18145),.ZN(_add_506_n406 ) );
NAND4_X2 _add_506_U601  ( .A1(n18149), .A2(n18153), .A3(n18157), .A4(_add_506_n398 ), .ZN(_add_506_n405 ) );
NAND4_X2 _add_506_U600  ( .A1(_add_506_n403 ), .A2(_add_506_n19 ), .A3(_add_506_n26 ), .A4(_add_506_n404 ), .ZN(_add_506_n402 ) );
XNOR2_X2 _add_506_U599  ( .A(_add_506_n402 ), .B(n18082), .ZN(N2153) );
NAND4_X2 _add_506_U598  ( .A1(n18133), .A2(n18137), .A3(n18141), .A4(n18145),.ZN(_add_506_n399 ) );
NAND4_X2 _add_506_U597  ( .A1(n18082), .A2(n18089), .A3(n18093), .A4(n18129),.ZN(_add_506_n400 ) );
NAND4_X2 _add_506_U596  ( .A1(n18149), .A2(n18153), .A3(n18157), .A4(_add_506_n398 ), .ZN(_add_506_n397 ) );
NAND4_X2 _add_506_U595  ( .A1(_add_506_n395 ), .A2(_add_506_n21 ), .A3(_add_506_n26 ), .A4(_add_506_n396 ), .ZN(_add_506_n394 ) );
XNOR2_X2 _add_506_U594  ( .A(_add_506_n394 ), .B(n18593), .ZN(N2154) );
NAND2_X2 _add_506_U593  ( .A1(_add_506_n2 ), .A2(_add_506_n30 ), .ZN(_add_506_n393 ) );
XNOR2_X2 _add_506_U592  ( .A(_add_506_n393 ), .B(n18541), .ZN(N2039) );
XNOR2_X2 _add_506_U591  ( .A(_add_506_n392 ), .B(n18537), .ZN(N2040) );
NAND2_X2 _add_506_U590  ( .A1(_add_506_n30 ), .A2(_add_506_n389 ), .ZN(_add_506_n388 ) );
XNOR2_X2 _add_506_U589  ( .A(_add_506_n388 ), .B(n18533), .ZN(N2041) );
NAND4_X2 _add_506_U588  ( .A1(n18533), .A2(n18537), .A3(n18541), .A4(n18545),.ZN(_add_506_n387 ) );
NAND2_X2 _add_506_U587  ( .A1(_add_506_n30 ), .A2(_add_506_n385 ), .ZN(_add_506_n384 ) );
XNOR2_X2 _add_506_U586  ( .A(_add_506_n384 ), .B(n18529), .ZN(N2042) );
NAND2_X2 _add_506_U585  ( .A1(n18537), .A2(n18541), .ZN(_add_506_n382 ) );
NAND2_X2 _add_506_U584  ( .A1(n18529), .A2(n18533), .ZN(_add_506_n383 ) );
NAND2_X2 _add_506_U583  ( .A1(n18553), .A2(n18557), .ZN(_add_506_n380 ) );
NAND2_X2 _add_506_U582  ( .A1(n18545), .A2(n18549), .ZN(_add_506_n381 ) );
NAND4_X2 _add_506_U581  ( .A1(n18577), .A2(n18581), .A3(n18585), .A4(n18589),.ZN(_add_506_n378 ) );
NAND4_X2 _add_506_U580  ( .A1(n18561), .A2(n18565), .A3(n18569), .A4(n18573),.ZN(_add_506_n379 ) );
XNOR2_X2 _add_506_U579  ( .A(_add_506_n374 ), .B(n18525), .ZN(N2043) );
NAND2_X2 _add_506_U578  ( .A1(_add_506_n337 ), .A2(n18525), .ZN(_add_506_n373 ) );
XNOR2_X2 _add_506_U577  ( .A(_add_506_n373 ), .B(n18521), .ZN(N2044) );
XNOR2_X2 _add_506_U576  ( .A(_add_506_n372 ), .B(n18517), .ZN(N2045) );
NAND4_X2 _add_506_U575  ( .A1(n18521), .A2(n18517), .A3(n18525), .A4(_add_506_n337 ), .ZN(_add_506_n371 ) );
XNOR2_X2 _add_506_U574  ( .A(_add_506_n371 ), .B(n18513), .ZN(N2046) );
NAND2_X2 _add_506_U573  ( .A1(_add_506_n337 ), .A2(_add_506_n362 ), .ZN(_add_506_n370 ) );
XNOR2_X2 _add_506_U572  ( .A(_add_506_n370 ), .B(n18509), .ZN(N2047) );
XNOR2_X2 _add_506_U571  ( .A(_add_506_n369 ), .B(n18505), .ZN(N2048) );
NAND4_X2 _add_506_U570  ( .A1(n18505), .A2(n18509), .A3(_add_506_n362 ),.A4(_add_506_n337 ), .ZN(_add_506_n368 ) );
XNOR2_X2 _add_506_U569  ( .A(_add_506_n368 ), .B(n18501), .ZN(N2049) );
NAND2_X2 _add_506_U568  ( .A1(_add_506_n366 ), .A2(_add_506_n337 ), .ZN(_add_506_n365 ) );
XNOR2_X2 _add_506_U567  ( .A(_add_506_n365 ), .B(n18497), .ZN(N2050) );
NAND4_X2 _add_506_U566  ( .A1(n18497), .A2(n18501), .A3(n18505), .A4(n18509),.ZN(_add_506_n339 ) );
NAND2_X2 _add_506_U565  ( .A1(_add_506_n364 ), .A2(_add_506_n337 ), .ZN(_add_506_n363 ) );
XNOR2_X2 _add_506_U564  ( .A(_add_506_n363 ), .B(n18493), .ZN(N2051) );
INV_X4 _add_506_U563  ( .A(_add_506_n339 ), .ZN(_add_506_n361 ) );
INV_X4 _add_506_U562  ( .A(_add_506_n607 ), .ZN(_add_506_n362 ) );
NAND4_X2 _add_506_U561  ( .A1(_add_506_n361 ), .A2(_add_506_n362 ), .A3(n18493), .A4(_add_506_n337 ), .ZN(_add_506_n360 ) );
XNOR2_X2 _add_506_U560  ( .A(_add_506_n360 ), .B(n18489), .ZN(N2052) );
NAND4_X2 _add_506_U559  ( .A1(n18489), .A2(n18493), .A3(_add_506_n359 ),.A4(_add_506_n337 ), .ZN(_add_506_n358 ) );
XNOR2_X2 _add_506_U558  ( .A(_add_506_n358 ), .B(n18485), .ZN(N2053) );
NAND2_X2 _add_506_U557  ( .A1(_add_506_n356 ), .A2(_add_506_n337 ), .ZN(_add_506_n355 ) );
XNOR2_X2 _add_506_U556  ( .A(_add_506_n355 ), .B(n18481), .ZN(N2054) );
NAND4_X2 _add_506_U555  ( .A1(n18481), .A2(n18485), .A3(n18489), .A4(n18493),.ZN(_add_506_n352 ) );
NAND2_X2 _add_506_U554  ( .A1(_add_506_n354 ), .A2(_add_506_n337 ), .ZN(_add_506_n353 ) );
XNOR2_X2 _add_506_U553  ( .A(_add_506_n353 ), .B(n18477), .ZN(N2055) );
INV_X4 _add_506_U552  ( .A(_add_506_n352 ), .ZN(_add_506_n341 ) );
NAND2_X2 _add_506_U551  ( .A1(_add_506_n341 ), .A2(n18477), .ZN(_add_506_n351 ) );
NAND2_X2 _add_506_U550  ( .A1(_add_506_n350 ), .A2(_add_506_n337 ), .ZN(_add_506_n349 ) );
XNOR2_X2 _add_506_U549  ( .A(_add_506_n349 ), .B(n18473), .ZN(N2056) );
NAND2_X2 _add_506_U548  ( .A1(n18585), .A2(n18589), .ZN(_add_506_n304 ) );
XNOR2_X2 _add_506_U547  ( .A(_add_506_n304 ), .B(n18581), .ZN(N2029) );
INV_X4 _add_506_U546  ( .A(n18477), .ZN(_add_506_n342 ) );
INV_X4 _add_506_U545  ( .A(n18473), .ZN(_add_506_n348 ) );
NAND2_X2 _add_506_U544  ( .A1(_add_506_n347 ), .A2(_add_506_n341 ), .ZN(_add_506_n346 ) );
NAND2_X2 _add_506_U543  ( .A1(_add_506_n345 ), .A2(_add_506_n337 ), .ZN(_add_506_n344 ) );
XNOR2_X2 _add_506_U542  ( .A(_add_506_n344 ), .B(n18469), .ZN(N2057) );
NAND2_X2 _add_506_U541  ( .A1(n18473), .A2(n18469), .ZN(_add_506_n343 ) );
NAND2_X2 _add_506_U540  ( .A1(_add_506_n340 ), .A2(_add_506_n341 ), .ZN(_add_506_n338 ) );
NAND2_X2 _add_506_U539  ( .A1(_add_506_n336 ), .A2(_add_506_n337 ), .ZN(_add_506_n335 ) );
XNOR2_X2 _add_506_U538  ( .A(_add_506_n335 ), .B(n18465), .ZN(N2058) );
NAND2_X2 _add_506_U537  ( .A1(n18505), .A2(n18509), .ZN(_add_506_n333 ) );
NAND2_X2 _add_506_U536  ( .A1(n18497), .A2(n18501), .ZN(_add_506_n334 ) );
NAND2_X2 _add_506_U535  ( .A1(n18521), .A2(n18525), .ZN(_add_506_n331 ) );
NAND2_X2 _add_506_U534  ( .A1(n18513), .A2(n18517), .ZN(_add_506_n332 ) );
NAND2_X2 _add_506_U533  ( .A1(_add_506_n329 ), .A2(_add_506_n330 ), .ZN(_add_506_n326 ) );
NAND4_X2 _add_506_U532  ( .A1(n18481), .A2(n18485), .A3(n18489), .A4(n18493),.ZN(_add_506_n327 ) );
NAND4_X2 _add_506_U531  ( .A1(n18465), .A2(n18469), .A3(n18473), .A4(n18477),.ZN(_add_506_n328 ) );
NAND2_X2 _add_506_U530  ( .A1(n18569), .A2(n18573), .ZN(_add_506_n324 ) );
NAND2_X2 _add_506_U529  ( .A1(n18561), .A2(n18565), .ZN(_add_506_n325 ) );
NAND2_X2 _add_506_U528  ( .A1(n18585), .A2(n18589), .ZN(_add_506_n322 ) );
NAND2_X2 _add_506_U527  ( .A1(n18577), .A2(n18581), .ZN(_add_506_n323 ) );
NAND2_X2 _add_506_U526  ( .A1(_add_506_n320 ), .A2(_add_506_n321 ), .ZN(_add_506_n317 ) );
NAND4_X2 _add_506_U525  ( .A1(n18545), .A2(n18549), .A3(n18553), .A4(n18557),.ZN(_add_506_n318 ) );
NAND4_X2 _add_506_U524  ( .A1(n18529), .A2(n18533), .A3(n18537), .A4(n18541),.ZN(_add_506_n319 ) );
NAND2_X2 _add_506_U523  ( .A1(_add_506_n315 ), .A2(_add_506_n316 ), .ZN(_add_506_n314 ) );
XNOR2_X2 _add_506_U522  ( .A(_add_506_n314 ), .B(n18461), .ZN(N2059) );
NAND2_X2 _add_506_U521  ( .A1(_add_506_n17 ), .A2(n18461), .ZN(_add_506_n313 ) );
XNOR2_X2 _add_506_U520  ( .A(_add_506_n313 ), .B(n18457), .ZN(N2060) );
XNOR2_X2 _add_506_U519  ( .A(_add_506_n312 ), .B(n18453), .ZN(N2061) );
NAND4_X2 _add_506_U518  ( .A1(n18457), .A2(n18453), .A3(n18461), .A4(_add_506_n15 ), .ZN(_add_506_n311 ) );
XNOR2_X2 _add_506_U517  ( .A(_add_506_n311 ), .B(n18449), .ZN(N2062) );
NAND2_X2 _add_506_U516  ( .A1(_add_506_n267 ), .A2(_add_506_n18 ), .ZN(_add_506_n310 ) );
XNOR2_X2 _add_506_U515  ( .A(_add_506_n310 ), .B(n18445), .ZN(N2063) );
INV_X4 _add_506_U514  ( .A(n18445), .ZN(_add_506_n280 ) );
NAND2_X2 _add_506_U513  ( .A1(_add_506_n309 ), .A2(_add_506_n18 ), .ZN(_add_506_n308 ) );
XNOR2_X2 _add_506_U512  ( .A(_add_506_n308 ), .B(n18441), .ZN(N2064) );
NAND4_X2 _add_506_U511  ( .A1(n18445), .A2(_add_506_n267 ), .A3(n18441),.A4(_add_506_n15 ), .ZN(_add_506_n307 ) );
XNOR2_X2 _add_506_U510  ( .A(_add_506_n307 ), .B(n18437), .ZN(N2065) );
NAND4_X2 _add_506_U509  ( .A1(n18441), .A2(n18437), .A3(_add_506_n306 ),.A4(_add_506_n15 ), .ZN(_add_506_n305 ) );
XNOR2_X2 _add_506_U508  ( .A(_add_506_n305 ), .B(n18433), .ZN(N2066) );
INV_X4 _add_506_U507  ( .A(_add_506_n304 ), .ZN(_add_506_n303 ) );
NAND2_X2 _add_506_U506  ( .A1(n18581), .A2(_add_506_n303 ), .ZN(_add_506_n302 ) );
XNOR2_X2 _add_506_U505  ( .A(_add_506_n302 ), .B(n18577), .ZN(N2030) );
NAND4_X2 _add_506_U504  ( .A1(n18433), .A2(n18437), .A3(n18441), .A4(n18445),.ZN(_add_506_n288 ) );
NAND2_X2 _add_506_U503  ( .A1(_add_506_n301 ), .A2(_add_506_n18 ), .ZN(_add_506_n300 ) );
XNOR2_X2 _add_506_U502  ( .A(_add_506_n300 ), .B(n18429), .ZN(N2067) );
INV_X4 _add_506_U501  ( .A(_add_506_n288 ), .ZN(_add_506_n299 ) );
NAND4_X2 _add_506_U500  ( .A1(n18429), .A2(_add_506_n267 ), .A3(_add_506_n299 ), .A4(_add_506_n15 ), .ZN(_add_506_n298 ) );
XNOR2_X2 _add_506_U499  ( .A(_add_506_n298 ), .B(n18425), .ZN(N2068) );
NAND2_X2 _add_506_U498  ( .A1(n18425), .A2(n18429), .ZN(_add_506_n297 ) );
NAND2_X2 _add_506_U497  ( .A1(_add_506_n17 ), .A2(_add_506_n296 ), .ZN(_add_506_n295 ) );
XNOR2_X2 _add_506_U496  ( .A(_add_506_n295 ), .B(n18421), .ZN(N2069) );
NAND2_X2 _add_506_U495  ( .A1(_add_506_n293 ), .A2(_add_506_n18 ), .ZN(_add_506_n292 ) );
XNOR2_X2 _add_506_U494  ( .A(_add_506_n292 ), .B(n18417), .ZN(N2070) );
NAND4_X2 _add_506_U493  ( .A1(n18417), .A2(n18421), .A3(n18425), .A4(n18429),.ZN(_add_506_n291 ) );
NAND2_X2 _add_506_U492  ( .A1(_add_506_n290 ), .A2(_add_506_n18 ), .ZN(_add_506_n289 ) );
XNOR2_X2 _add_506_U491  ( .A(_add_506_n289 ), .B(n18413), .ZN(N2071) );
NAND2_X2 _add_506_U490  ( .A1(_add_506_n299 ), .A2(n18413), .ZN(_add_506_n286 ) );
NAND4_X2 _add_506_U489  ( .A1(n18417), .A2(n18421), .A3(n18425), .A4(n18429),.ZN(_add_506_n287 ) );
NAND2_X2 _add_506_U488  ( .A1(_add_506_n285 ), .A2(_add_506_n18 ), .ZN(_add_506_n284 ) );
XNOR2_X2 _add_506_U487  ( .A(_add_506_n284 ), .B(n18409), .ZN(N2072) );
INV_X4 _add_506_U486  ( .A(n18429), .ZN(_add_506_n282 ) );
NAND2_X2 _add_506_U485  ( .A1(n18425), .A2(n18433), .ZN(_add_506_n283 ) );
NAND2_X2 _add_506_U484  ( .A1(n18441), .A2(n18437), .ZN(_add_506_n281 ) );
NAND2_X2 _add_506_U483  ( .A1(_add_506_n278 ), .A2(_add_506_n279 ), .ZN(_add_506_n276 ) );
NAND4_X2 _add_506_U482  ( .A1(n18409), .A2(n18421), .A3(n18417), .A4(n18413),.ZN(_add_506_n277 ) );
NAND2_X2 _add_506_U481  ( .A1(_add_506_n275 ), .A2(_add_506_n17 ), .ZN(_add_506_n274 ) );
XNOR2_X2 _add_506_U480  ( .A(_add_506_n274 ), .B(n18405), .ZN(N2073) );
INV_X4 _add_506_U479  ( .A(_add_506_n621 ), .ZN(_add_506_n267 ) );
NAND4_X2 _add_506_U478  ( .A1(n18433), .A2(n18437), .A3(n18441), .A4(n18445),.ZN(_add_506_n272 ) );
NAND2_X2 _add_506_U477  ( .A1(n18413), .A2(n18409), .ZN(_add_506_n270 ) );
NAND2_X2 _add_506_U476  ( .A1(n18405), .A2(n18417), .ZN(_add_506_n271 ) );
NAND4_X2 _add_506_U475  ( .A1(_add_506_n267 ), .A2(_add_506_n268 ), .A3(_add_506_n269 ), .A4(_add_506_n16 ), .ZN(_add_506_n266 ) );
XNOR2_X2 _add_506_U474  ( .A(_add_506_n266 ), .B(n18401), .ZN(N2074) );
NAND2_X2 _add_506_U473  ( .A1(_add_506_n27 ), .A2(_add_506_n17 ), .ZN(_add_506_n265 ) );
XNOR2_X2 _add_506_U472  ( .A(_add_506_n265 ), .B(n18397), .ZN(N2075) );
INV_X4 _add_506_U471  ( .A(n18397), .ZN(_add_506_n234 ) );
NAND2_X2 _add_506_U470  ( .A1(_add_506_n264 ), .A2(_add_506_n18 ), .ZN(_add_506_n263 ) );
XNOR2_X2 _add_506_U469  ( .A(_add_506_n263 ), .B(n18393), .ZN(N2076) );
INV_X4 _add_506_U468  ( .A(n18573), .ZN(_add_506_n262 ) );
XNOR2_X2 _add_506_U467  ( .A(_add_506_n262 ), .B(_add_506_n4 ), .ZN(N2031));
NAND4_X2 _add_506_U466  ( .A1(n18397), .A2(_add_506_n27 ), .A3(n18393), .A4(_add_506_n16 ), .ZN(_add_506_n261 ) );
XNOR2_X2 _add_506_U465  ( .A(_add_506_n261 ), .B(n18389), .ZN(N2077) );
NAND4_X2 _add_506_U464  ( .A1(n18393), .A2(n18389), .A3(_add_506_n260 ),.A4(_add_506_n16 ), .ZN(_add_506_n259 ) );
XNOR2_X2 _add_506_U463  ( .A(_add_506_n259 ), .B(n18385), .ZN(N2078) );
NAND4_X2 _add_506_U462  ( .A1(n18385), .A2(n18389), .A3(n18393), .A4(n18397),.ZN(_add_506_n244 ) );
NAND2_X2 _add_506_U461  ( .A1(_add_506_n258 ), .A2(_add_506_n17 ), .ZN(_add_506_n257 ) );
XNOR2_X2 _add_506_U460  ( .A(_add_506_n257 ), .B(n18381), .ZN(N2079) );
INV_X4 _add_506_U459  ( .A(_add_506_n244 ), .ZN(_add_506_n247 ) );
NAND4_X2 _add_506_U458  ( .A1(_add_506_n247 ), .A2(n18381), .A3(_add_506_n26 ), .A4(_add_506_n16 ), .ZN(_add_506_n256 ) );
XNOR2_X2 _add_506_U457  ( .A(_add_506_n256 ), .B(n18377), .ZN(N2080) );
NAND2_X2 _add_506_U456  ( .A1(n18377), .A2(n18381), .ZN(_add_506_n255 ) );
NAND2_X2 _add_506_U455  ( .A1(_add_506_n17 ), .A2(_add_506_n254 ), .ZN(_add_506_n253 ) );
XNOR2_X2 _add_506_U454  ( .A(_add_506_n253 ), .B(n18373), .ZN(N2081) );
INV_X4 _add_506_U453  ( .A(n18381), .ZN(_add_506_n236 ) );
NAND2_X2 _add_506_U452  ( .A1(n18377), .A2(n18373), .ZN(_add_506_n252 ) );
NAND4_X2 _add_506_U451  ( .A1(_add_506_n251 ), .A2(_add_506_n247 ), .A3(_add_506_n26 ), .A4(_add_506_n16 ), .ZN(_add_506_n250 ) );
XNOR2_X2 _add_506_U450  ( .A(_add_506_n250 ), .B(n18369), .ZN(N2082) );
NAND2_X2 _add_506_U449  ( .A1(n18377), .A2(n18381), .ZN(_add_506_n248 ) );
NAND2_X2 _add_506_U448  ( .A1(n18369), .A2(n18373), .ZN(_add_506_n249 ) );
NAND4_X2 _add_506_U447  ( .A1(_add_506_n246 ), .A2(_add_506_n247 ), .A3(_add_506_n26 ), .A4(_add_506_n16 ), .ZN(_add_506_n245 ) );
XNOR2_X2 _add_506_U446  ( .A(_add_506_n245 ), .B(n18365), .ZN(N2083) );
INV_X4 _add_506_U445  ( .A(n18365), .ZN(_add_506_n243 ) );
NAND2_X2 _add_506_U444  ( .A1(n18377), .A2(n18381), .ZN(_add_506_n241 ) );
NAND2_X2 _add_506_U443  ( .A1(n18373), .A2(n18369), .ZN(_add_506_n242 ) );
NAND4_X2 _add_506_U442  ( .A1(_add_506_n239 ), .A2(_add_506_n240 ), .A3(_add_506_n26 ), .A4(_add_506_n16 ), .ZN(_add_506_n238 ) );
XNOR2_X2 _add_506_U441  ( .A(_add_506_n238 ), .B(n18361), .ZN(N2084) );
NAND2_X2 _add_506_U440  ( .A1(n18377), .A2(n18385), .ZN(_add_506_n237 ) );
NAND2_X2 _add_506_U439  ( .A1(n18393), .A2(n18389), .ZN(_add_506_n235 ) );
NAND2_X2 _add_506_U438  ( .A1(_add_506_n232 ), .A2(_add_506_n233 ), .ZN(_add_506_n230 ) );
NAND4_X2 _add_506_U437  ( .A1(n18361), .A2(n18373), .A3(n18369), .A4(n18365),.ZN(_add_506_n231 ) );
NAND2_X2 _add_506_U436  ( .A1(_add_506_n229 ), .A2(_add_506_n18 ), .ZN(_add_506_n228 ) );
XNOR2_X2 _add_506_U435  ( .A(_add_506_n228 ), .B(n18357), .ZN(N2085) );
NAND4_X2 _add_506_U434  ( .A1(n18385), .A2(n18389), .A3(n18393), .A4(n18397),.ZN(_add_506_n226 ) );
NAND2_X2 _add_506_U433  ( .A1(n18365), .A2(n18361), .ZN(_add_506_n224 ) );
NAND2_X2 _add_506_U432  ( .A1(n18357), .A2(n18369), .ZN(_add_506_n225 ) );
NAND4_X2 _add_506_U431  ( .A1(_add_506_n222 ), .A2(_add_506_n27 ), .A3(_add_506_n223 ), .A4(_add_506_n16 ), .ZN(_add_506_n221 ) );
XNOR2_X2 _add_506_U430  ( .A(_add_506_n221 ), .B(n18353), .ZN(N2086) );
NAND2_X2 _add_506_U429  ( .A1(_add_506_n4 ), .A2(n18573), .ZN(_add_506_n220 ) );
XNOR2_X2 _add_506_U428  ( .A(_add_506_n220 ), .B(n18569), .ZN(N2032) );
NAND2_X2 _add_506_U427  ( .A1(_add_506_n213 ), .A2(_add_506_n18 ), .ZN(_add_506_n212 ) );
XNOR2_X2 _add_506_U426  ( .A(_add_506_n212 ), .B(n18349), .ZN(N2087) );
INV_X4 _add_506_U425  ( .A(_add_506_n135 ), .ZN(_add_506_n211 ) );
NAND4_X2 _add_506_U424  ( .A1(_add_506_n211 ), .A2(_add_506_n27 ), .A3(n18349), .A4(_add_506_n15 ), .ZN(_add_506_n210 ) );
XNOR2_X2 _add_506_U423  ( .A(_add_506_n210 ), .B(n18345), .ZN(N2088) );
NAND2_X2 _add_506_U422  ( .A1(n18345), .A2(n18349), .ZN(_add_506_n209 ) );
NAND2_X2 _add_506_U421  ( .A1(_add_506_n17 ), .A2(_add_506_n208 ), .ZN(_add_506_n207 ) );
XNOR2_X2 _add_506_U420  ( .A(_add_506_n207 ), .B(n18341), .ZN(N2089) );
NAND2_X2 _add_506_U419  ( .A1(_add_506_n205 ), .A2(_add_506_n18 ), .ZN(_add_506_n204 ) );
XNOR2_X2 _add_506_U418  ( .A(_add_506_n204 ), .B(n18337), .ZN(N2090) );
NAND4_X2 _add_506_U417  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(_add_506_n199 ) );
NAND2_X2 _add_506_U416  ( .A1(_add_506_n17 ), .A2(_add_506_n203 ), .ZN(_add_506_n202 ) );
XNOR2_X2 _add_506_U415  ( .A(_add_506_n202 ), .B(n18333), .ZN(N2091) );
NAND4_X2 _add_506_U414  ( .A1(_add_506_n201 ), .A2(_add_506_n17 ), .A3(_add_506_n26 ), .A4(n18333), .ZN(_add_506_n200 ) );
XNOR2_X2 _add_506_U413  ( .A(_add_506_n200 ), .B(n18329), .ZN(N2092) );
NAND3_X2 _add_506_U412  ( .A1(_add_506_n197 ), .A2(_add_506_n17 ), .A3(_add_506_n198 ), .ZN(_add_506_n196 ) );
XNOR2_X2 _add_506_U411  ( .A(_add_506_n196 ), .B(n18325), .ZN(N2093) );
NAND2_X2 _add_506_U410  ( .A1(n18345), .A2(n18341), .ZN(_add_506_n195 ) );
INV_X4 _add_506_U409  ( .A(n18325), .ZN(_add_506_n187 ) );
NAND4_X2 _add_506_U408  ( .A1(_add_506_n16 ), .A2(_add_506_n192 ), .A3(_add_506_n26 ), .A4(_add_506_n193 ), .ZN(_add_506_n191 ) );
XNOR2_X2 _add_506_U407  ( .A(_add_506_n191 ), .B(n18321), .ZN(N2094) );
INV_X4 _add_506_U406  ( .A(n18321), .ZN(_add_506_n188 ) );
NAND4_X2 _add_506_U405  ( .A1(_add_506_n16 ), .A2(_add_506_n185 ), .A3(_add_506_n26 ), .A4(_add_506_n186 ), .ZN(_add_506_n184 ) );
XNOR2_X2 _add_506_U404  ( .A(_add_506_n184 ), .B(n18317), .ZN(N2095) );
NAND3_X2 _add_506_U403  ( .A1(_add_506_n179 ), .A2(_add_506_n17 ), .A3(_add_506_n180 ), .ZN(_add_506_n178 ) );
XNOR2_X2 _add_506_U402  ( .A(_add_506_n178 ), .B(n18313), .ZN(N2096) );
XNOR2_X2 _add_506_U401  ( .A(_add_506_n177 ), .B(n18565), .ZN(N2033) );
NAND4_X2 _add_506_U400  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(_add_506_n175 ) );
NAND3_X2 _add_506_U399  ( .A1(_add_506_n172 ), .A2(_add_506_n17 ), .A3(_add_506_n173 ), .ZN(_add_506_n171 ) );
XNOR2_X2 _add_506_U398  ( .A(_add_506_n171 ), .B(n18309), .ZN(N2097) );
NAND4_X2 _add_506_U397  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(_add_506_n169 ) );
NAND4_X2 _add_506_U396  ( .A1(n18309), .A2(n18313), .A3(n18317), .A4(n18321),.ZN(_add_506_n168 ) );
NAND3_X2 _add_506_U395  ( .A1(_add_506_n166 ), .A2(_add_506_n17 ), .A3(_add_506_n167 ), .ZN(_add_506_n165 ) );
XNOR2_X2 _add_506_U394  ( .A(_add_506_n165 ), .B(n18305), .ZN(N2098) );
NAND4_X2 _add_506_U393  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(_add_506_n163 ) );
NAND4_X2 _add_506_U392  ( .A1(n18321), .A2(n18325), .A3(n18329), .A4(n18333),.ZN(_add_506_n164 ) );
NAND4_X2 _add_506_U391  ( .A1(n18305), .A2(n18309), .A3(n18313), .A4(n18317),.ZN(_add_506_n162 ) );
NAND3_X2 _add_506_U390  ( .A1(_add_506_n160 ), .A2(_add_506_n17 ), .A3(_add_506_n161 ), .ZN(_add_506_n159 ) );
XNOR2_X2 _add_506_U389  ( .A(_add_506_n159 ), .B(n18301), .ZN(N2099) );
NAND2_X2 _add_506_U388  ( .A1(n18329), .A2(n18333), .ZN(_add_506_n157 ) );
NAND2_X2 _add_506_U387  ( .A1(n18321), .A2(n18325), .ZN(_add_506_n158 ) );
NAND2_X2 _add_506_U386  ( .A1(n18345), .A2(n18349), .ZN(_add_506_n155 ) );
NAND2_X2 _add_506_U385  ( .A1(n18337), .A2(n18341), .ZN(_add_506_n156 ) );
INV_X4 _add_506_U384  ( .A(n18301), .ZN(_add_506_n154 ) );
NAND4_X2 _add_506_U383  ( .A1(_add_506_n151 ), .A2(_add_506_n152 ), .A3(_add_506_n26 ), .A4(_add_506_n153 ), .ZN(_add_506_n149 ) );
NAND4_X2 _add_506_U382  ( .A1(n18305), .A2(n18309), .A3(n18313), .A4(n18317),.ZN(_add_506_n150 ) );
NAND2_X2 _add_506_U381  ( .A1(n18341), .A2(n18345), .ZN(_add_506_n146 ) );
NAND4_X2 _add_506_U380  ( .A1(n18317), .A2(n18321), .A3(n18325), .A4(n18329),.ZN(_add_506_n148 ) );
INV_X4 _add_506_U379  ( .A(n18297), .ZN(_add_506_n145 ) );
NAND4_X2 _add_506_U378  ( .A1(n18301), .A2(n18305), .A3(n18309), .A4(n18313),.ZN(_add_506_n144 ) );
NAND4_X2 _add_506_U377  ( .A1(_add_506_n141 ), .A2(_add_506_n27 ), .A3(_add_506_n142 ), .A4(_add_506_n143 ), .ZN(_add_506_n140 ) );
XNOR2_X2 _add_506_U376  ( .A(_add_506_n140 ), .B(n18293), .ZN(N2101) );
NAND2_X2 _add_506_U375  ( .A1(n18345), .A2(n18341), .ZN(_add_506_n137 ) );
NAND4_X2 _add_506_U374  ( .A1(n18317), .A2(n18321), .A3(n18325), .A4(n18329),.ZN(_add_506_n139 ) );
INV_X4 _add_506_U373  ( .A(n18293), .ZN(_add_506_n136 ) );
NAND2_X2 _add_506_U372  ( .A1(n18309), .A2(n18305), .ZN(_add_506_n134 ) );
NAND4_X2 _add_506_U371  ( .A1(_add_506_n130 ), .A2(_add_506_n27 ), .A3(_add_506_n131 ), .A4(_add_506_n132 ), .ZN(_add_506_n129 ) );
XNOR2_X2 _add_506_U370  ( .A(_add_506_n129 ), .B(n18289), .ZN(N2102) );
NAND3_X2 _add_506_U369  ( .A1(_add_506_n21 ), .A2(_add_506_n27 ), .A3(_add_506_n17 ), .ZN(_add_506_n128 ) );
XNOR2_X2 _add_506_U368  ( .A(_add_506_n128 ), .B(n18285), .ZN(N2103) );
NAND4_X2 _add_506_U367  ( .A1(_add_506_n26 ), .A2(_add_506_n20 ), .A3(_add_506_n16 ), .A4(n18285), .ZN(_add_506_n127 ) );
XNOR2_X2 _add_506_U366  ( .A(_add_506_n127 ), .B(n18281), .ZN(N2104) );
INV_X4 _add_506_U365  ( .A(n18285), .ZN(_add_506_n122 ) );
INV_X4 _add_506_U364  ( .A(n18281), .ZN(_add_506_n126 ) );
NAND4_X2 _add_506_U363  ( .A1(_add_506_n27 ), .A2(_add_506_n20 ), .A3(_add_506_n125 ), .A4(_add_506_n15 ), .ZN(_add_506_n124 ) );
XNOR2_X2 _add_506_U362  ( .A(_add_506_n124 ), .B(n18277), .ZN(N2105) );
NAND2_X2 _add_506_U361  ( .A1(n18281), .A2(n18277), .ZN(_add_506_n123 ) );
NAND4_X2 _add_506_U360  ( .A1(_add_506_n121 ), .A2(_add_506_n16 ), .A3(_add_506_n19 ), .A4(_add_506_n26 ), .ZN(_add_506_n120 ) );
XNOR2_X2 _add_506_U359  ( .A(_add_506_n120 ), .B(n18273), .ZN(N2106) );
NAND4_X2 _add_506_U358  ( .A1(n18569), .A2(n18565), .A3(n18573), .A4(_add_506_n4 ), .ZN(_add_506_n119 ) );
XNOR2_X2 _add_506_U357  ( .A(_add_506_n119 ), .B(n18561), .ZN(N2034) );
NAND4_X2 _add_506_U356  ( .A1(n18273), .A2(n18277), .A3(n18281), .A4(n18285),.ZN(_add_506_n114 ) );
NAND3_X2 _add_506_U355  ( .A1(_add_506_n21 ), .A2(_add_506_n118 ), .A3(_add_506_n17 ), .ZN(_add_506_n117 ) );
XNOR2_X2 _add_506_U354  ( .A(_add_506_n117 ), .B(n18269), .ZN(N2107) );
NAND4_X2 _add_506_U353  ( .A1(_add_506_n20 ), .A2(n18269), .A3(_add_506_n116 ), .A4(_add_506_n16 ), .ZN(_add_506_n115 ) );
XNOR2_X2 _add_506_U352  ( .A(_add_506_n115 ), .B(n18265), .ZN(N2108) );
INV_X4 _add_506_U351  ( .A(n18269), .ZN(_add_506_n102 ) );
INV_X4 _add_506_U350  ( .A(n18265), .ZN(_add_506_n103 ) );
NAND4_X2 _add_506_U349  ( .A1(_add_506_n112 ), .A2(_add_506_n20 ), .A3(_add_506_n113 ), .A4(_add_506_n15 ), .ZN(_add_506_n111 ) );
XNOR2_X2 _add_506_U348  ( .A(_add_506_n111 ), .B(n18261), .ZN(N2109) );
NAND2_X2 _add_506_U347  ( .A1(n18281), .A2(n18277), .ZN(_add_506_n110 ) );
INV_X4 _add_506_U346  ( .A(n18261), .ZN(_add_506_n104 ) );
NAND4_X2 _add_506_U345  ( .A1(_add_506_n107 ), .A2(_add_506_n21 ), .A3(_add_506_n108 ), .A4(_add_506_n16 ), .ZN(_add_506_n106 ) );
XNOR2_X2 _add_506_U344  ( .A(_add_506_n106 ), .B(n18257), .ZN(N2110) );
INV_X4 _add_506_U343  ( .A(n18257), .ZN(_add_506_n105 ) );
NAND2_X2 _add_506_U342  ( .A1(n18281), .A2(n18285), .ZN(_add_506_n100 ) );
NAND2_X2 _add_506_U341  ( .A1(n18273), .A2(n18277), .ZN(_add_506_n101 ) );
NAND3_X2 _add_506_U340  ( .A1(_add_506_n21 ), .A2(_add_506_n96 ), .A3(_add_506_n17 ), .ZN(_add_506_n95 ) );
XNOR2_X2 _add_506_U339  ( .A(_add_506_n95 ), .B(n18253), .ZN(N2111) );
NAND4_X2 _add_506_U338  ( .A1(_add_506_n19 ), .A2(n18253), .A3(_add_506_n94 ), .A4(_add_506_n15 ), .ZN(_add_506_n93 ) );
XNOR2_X2 _add_506_U337  ( .A(_add_506_n93 ), .B(n18249), .ZN(N2112) );
INV_X4 _add_506_U336  ( .A(n18253), .ZN(_add_506_n87 ) );
INV_X4 _add_506_U335  ( .A(n18249), .ZN(_add_506_n92 ) );
NAND4_X2 _add_506_U334  ( .A1(_add_506_n90 ), .A2(_add_506_n21 ), .A3(_add_506_n91 ), .A4(_add_506_n15 ), .ZN(_add_506_n89 ) );
XNOR2_X2 _add_506_U333  ( .A(_add_506_n89 ), .B(n18245), .ZN(N2113) );
NAND2_X2 _add_506_U332  ( .A1(n18249), .A2(n18245), .ZN(_add_506_n88 ) );
NAND4_X2 _add_506_U331  ( .A1(_add_506_n85 ), .A2(_add_506_n21 ), .A3(_add_506_n86 ), .A4(_add_506_n15 ), .ZN(_add_506_n84 ) );
XNOR2_X2 _add_506_U330  ( .A(_add_506_n84 ), .B(n18241), .ZN(N2114) );
INV_X4 _add_506_U329  ( .A(_add_506_n75 ), .ZN(_add_506_n70 ) );
NAND4_X2 _add_506_U328  ( .A1(n18241), .A2(n18245), .A3(n18249), .A4(n18253),.ZN(_add_506_n76 ) );
INV_X4 _add_506_U327  ( .A(_add_506_n76 ), .ZN(_add_506_n71 ) );
AND2_X2 _add_506_U326  ( .A1(_add_506_n70 ), .A2(_add_506_n71 ), .ZN(_add_506_n83 ) );
NAND4_X2 _add_506_U325  ( .A1(_add_506_n19 ), .A2(_add_506_n27 ), .A3(_add_506_n83 ), .A4(_add_506_n15 ), .ZN(_add_506_n82 ) );
XNOR2_X2 _add_506_U324  ( .A(_add_506_n82 ), .B(n18237), .ZN(N2115) );
NAND2_X2 _add_506_U323  ( .A1(_add_506_n71 ), .A2(_add_506_n70 ), .ZN(_add_506_n81 ) );
NAND4_X2 _add_506_U322  ( .A1(_add_506_n19 ), .A2(n18237), .A3(_add_506_n80 ), .A4(_add_506_n15 ), .ZN(_add_506_n79 ) );
XNOR2_X2 _add_506_U321  ( .A(_add_506_n79 ), .B(n18233), .ZN(N2116) );
INV_X4 _add_506_U320  ( .A(n18557), .ZN(_add_506_n78 ) );
XNOR2_X2 _add_506_U319  ( .A(_add_506_n78 ), .B(_add_506_n30 ), .ZN(N2035));
INV_X4 _add_506_U318  ( .A(n18237), .ZN(_add_506_n67 ) );
INV_X4 _add_506_U317  ( .A(n18233), .ZN(_add_506_n77 ) );
NAND4_X2 _add_506_U316  ( .A1(_add_506_n19 ), .A2(_add_506_n73 ), .A3(_add_506_n74 ), .A4(_add_506_n15 ), .ZN(_add_506_n72 ) );
XNOR2_X2 _add_506_U315  ( .A(_add_506_n72 ), .B(n18229), .ZN(N2117) );
NAND2_X2 _add_506_U314  ( .A1(_add_506_n70 ), .A2(_add_506_n71 ), .ZN(_add_506_n69 ) );
NAND2_X2 _add_506_U313  ( .A1(n18233), .A2(n18229), .ZN(_add_506_n68 ) );
NAND4_X2 _add_506_U312  ( .A1(_add_506_n19 ), .A2(_add_506_n65 ), .A3(_add_506_n66 ), .A4(_add_506_n15 ), .ZN(_add_506_n64 ) );
XNOR2_X2 _add_506_U311  ( .A(_add_506_n64 ), .B(n18225), .ZN(N2118) );
NAND4_X2 _add_506_U310  ( .A1(_add_506_n27 ), .A2(_add_506_n21 ), .A3(_add_506_n63 ), .A4(_add_506_n15 ), .ZN(_add_506_n62 ) );
XNOR2_X2 _add_506_U309  ( .A(_add_506_n62 ), .B(n18221), .ZN(N2119) );
INV_X4 _add_506_U308  ( .A(n18221), .ZN(_add_506_n52 ) );
NAND4_X2 _add_506_U307  ( .A1(_add_506_n27 ), .A2(_add_506_n20 ), .A3(_add_506_n61 ), .A4(_add_506_n15 ), .ZN(_add_506_n60 ) );
XNOR2_X2 _add_506_U306  ( .A(_add_506_n60 ), .B(n18217), .ZN(N2120) );
NAND2_X2 _add_506_U305  ( .A1(n18217), .A2(n18221), .ZN(_add_506_n58 ) );
NAND2_X2 _add_506_U304  ( .A1(_add_506_n55 ), .A2(_add_506_n56 ), .ZN(_add_506_n54 ) );
XNOR2_X2 _add_506_U303  ( .A(_add_506_n54 ), .B(n18213), .ZN(N2121) );
NAND2_X2 _add_506_U302  ( .A1(n18217), .A2(n18213), .ZN(_add_506_n53 ) );
NAND4_X2 _add_506_U301  ( .A1(_add_506_n50 ), .A2(_add_506_n21 ), .A3(_add_506_n51 ), .A4(_add_506_n15 ), .ZN(_add_506_n49 ) );
XNOR2_X2 _add_506_U300  ( .A(_add_506_n49 ), .B(n18209), .ZN(N2122) );
NAND4_X2 _add_506_U299  ( .A1(n18209), .A2(n18213), .A3(n18217), .A4(n18221),.ZN(_add_506_n43 ) );
NAND4_X2 _add_506_U298  ( .A1(_add_506_n27 ), .A2(_add_506_n21 ), .A3(_add_506_n48 ), .A4(_add_506_n15 ), .ZN(_add_506_n47 ) );
XNOR2_X2 _add_506_U297  ( .A(_add_506_n47 ), .B(n18205), .ZN(N2123) );
NAND4_X2 _add_506_U296  ( .A1(_add_506_n45 ), .A2(_add_506_n21 ), .A3(_add_506_n46 ), .A4(_add_506_n15 ), .ZN(_add_506_n44 ) );
XNOR2_X2 _add_506_U295  ( .A(_add_506_n44 ), .B(n18201), .ZN(N2124) );
INV_X4 _add_506_U294  ( .A(_add_506_n43 ), .ZN(_add_506_n35 ) );
NAND2_X2 _add_506_U293  ( .A1(n18205), .A2(n18201), .ZN(_add_506_n42 ) );
NAND4_X2 _add_506_U292  ( .A1(_add_506_n35 ), .A2(_add_506_n16 ), .A3(_add_506_n41 ), .A4(_add_506_n19 ), .ZN(_add_506_n40 ) );
XNOR2_X2 _add_506_U291  ( .A(_add_506_n40 ), .B(n18197), .ZN(N2125) );
NAND2_X2 _add_506_U290  ( .A1(n18197), .A2(n18201), .ZN(_add_506_n38 ) );
NAND3_X2 _add_506_U289  ( .A1(_add_506_n36 ), .A2(_add_506_n27 ), .A3(_add_506_n21 ), .ZN(_add_506_n33 ) );
NAND2_X2 _add_506_U288  ( .A1(_add_506_n35 ), .A2(_add_506_n18 ), .ZN(_add_506_n34 ) );
XNOR2_X2 _add_506_U287  ( .A(_add_506_n31 ), .B(_add_506_n32 ), .ZN(N2126));
NAND2_X2 _add_506_U286  ( .A1(n18557), .A2(_add_506_n30 ), .ZN(_add_506_n29 ) );
XNOR2_X2 _add_506_U285  ( .A(_add_506_n29 ), .B(n18553), .ZN(N2036) );
INV_X4 _add_506_U284  ( .A(n18129), .ZN(_add_506_n14 ) );
INV_X4 _add_506_U283  ( .A(n18329), .ZN(_add_506_n12 ) );
NOR2_X2 _add_506_U282  ( .A1(_add_506_n342 ), .A2(_add_506_n348 ), .ZN(_add_506_n347 ) );
NOR2_X2 _add_506_U281  ( .A1(_add_506_n342 ), .A2(_add_506_n343 ), .ZN(_add_506_n340 ) );
NAND3_X2 _add_506_U280  ( .A1(n18149), .A2(n18157), .A3(n18153), .ZN(_add_506_n457 ) );
NOR2_X2 _add_506_U279  ( .A1(_add_506_n25 ), .A2(_add_506_n457 ), .ZN(_add_506_n456 ) );
INV_X4 _add_506_U278  ( .A(n18157), .ZN(_add_506_n13 ) );
INV_X4 _add_506_U277  ( .A(n18333), .ZN(_add_506_n11 ) );
NAND3_X2 _add_506_U276  ( .A1(n18345), .A2(n18353), .A3(n18349), .ZN(_add_506_n634 ) );
NAND3_X2 _add_506_U275  ( .A1(n18089), .A2(n18129), .A3(n18093), .ZN(_add_506_n407 ) );
NOR2_X2 _add_506_U274  ( .A1(_add_506_n144 ), .A2(_add_506_n57 ), .ZN(_add_506_n143 ) );
NOR2_X2 _add_506_U273  ( .A1(_add_506_n405 ), .A2(_add_506_n57 ), .ZN(_add_506_n404 ) );
NOR2_X2 _add_506_U272  ( .A1(_add_506_n397 ), .A2(_add_506_n57 ), .ZN(_add_506_n396 ) );
NAND3_X2 _add_506_U271  ( .A1(n18377), .A2(n18385), .A3(n18381), .ZN(_add_506_n217 ) );
NAND3_X2 _add_506_U270  ( .A1(n18393), .A2(n18389), .A3(n18397), .ZN(_add_506_n216 ) );
NOR2_X2 _add_506_U269  ( .A1(_add_506_n216 ), .A2(_add_506_n217 ), .ZN(_add_506_n215 ) );
NAND3_X2 _add_506_U268  ( .A1(n18357), .A2(n18353), .A3(n18361), .ZN(_add_506_n219 ) );
NOR2_X2 _add_506_U267  ( .A1(_add_506_n288 ), .A2(_add_506_n621 ), .ZN(_add_506_n301 ) );
NAND3_X2 _add_506_U266  ( .A1(n18425), .A2(n18421), .A3(n18429), .ZN(_add_506_n294 ) );
NOR3_X2 _add_506_U265  ( .A1(_add_506_n621 ), .A2(_add_506_n288 ), .A3(_add_506_n294 ), .ZN(_add_506_n293 ) );
NOR3_X2 _add_506_U264  ( .A1(_add_506_n621 ), .A2(_add_506_n288 ), .A3(_add_506_n291 ), .ZN(_add_506_n290 ) );
NOR2_X2 _add_506_U263  ( .A1(_add_506_n234 ), .A2(_add_506_n24 ), .ZN(_add_506_n264 ) );
NOR3_X2 _add_506_U262  ( .A1(_add_506_n24 ), .A2(_add_506_n230 ), .A3(_add_506_n231 ), .ZN(_add_506_n229 ) );
NOR3_X2 _add_506_U261  ( .A1(_add_506_n276 ), .A2(_add_506_n621 ), .A3(_add_506_n277 ), .ZN(_add_506_n275 ) );
NOR2_X2 _add_506_U260  ( .A1(_add_506_n244 ), .A2(_add_506_n24 ), .ZN(_add_506_n258 ) );
NOR2_X2 _add_506_U259  ( .A1(_add_506_n439 ), .A2(_add_506_n57 ), .ZN(_add_506_n429 ) );
NOR2_X2 _add_506_U258  ( .A1(_add_506_n59 ), .A2(_add_506_n431 ), .ZN(_add_506_n430 ) );
NOR2_X2 _add_506_U257  ( .A1(_add_506_n425 ), .A2(_add_506_n57 ), .ZN(_add_506_n416 ) );
NOR3_X2 _add_506_U256  ( .A1(_add_506_n59 ), .A2(_add_506_n418 ), .A3(_add_506_n23 ), .ZN(_add_506_n417 ) );
NAND3_X2 _add_506_U255  ( .A1(n18505), .A2(n18501), .A3(n18509), .ZN(_add_506_n367 ) );
NOR2_X2 _add_506_U254  ( .A1(_add_506_n607 ), .A2(_add_506_n367 ), .ZN(_add_506_n366 ) );
NAND3_X2 _add_506_U253  ( .A1(n18489), .A2(n18485), .A3(n18493), .ZN(_add_506_n357 ) );
NOR3_X2 _add_506_U252  ( .A1(_add_506_n607 ), .A2(_add_506_n339 ), .A3(_add_506_n357 ), .ZN(_add_506_n356 ) );
NOR3_X2 _add_506_U251  ( .A1(_add_506_n338 ), .A2(_add_506_n339 ), .A3(_add_506_n607 ), .ZN(_add_506_n336 ) );
NOR3_X2 _add_506_U250  ( .A1(_add_506_n59 ), .A2(_add_506_n37 ), .A3(_add_506_n23 ), .ZN(_add_506_n55 ) );
NOR2_X2 _add_506_U249  ( .A1(_add_506_n57 ), .A2(_add_506_n58 ), .ZN(_add_506_n56 ) );
NOR3_X2 _add_506_U248  ( .A1(_add_506_n607 ), .A2(_add_506_n352 ), .A3(_add_506_n339 ), .ZN(_add_506_n354 ) );
NOR3_X2 _add_506_U247  ( .A1(_add_506_n37 ), .A2(_add_506_n38 ), .A3(_add_506_n39 ), .ZN(_add_506_n36 ) );
NAND3_X2 _add_506_U246  ( .A1(n18457), .A2(n18461), .A3(_add_506_n15 ), .ZN(_add_506_n312 ) );
NAND3_X2 _add_506_U245  ( .A1(n18117), .A2(n18113), .A3(n18121), .ZN(_add_506_n468 ) );
NOR2_X2 _add_506_U244  ( .A1(_add_506_n13 ), .A2(_add_506_n441 ), .ZN(_add_506_n440 ) );
NOR3_X2 _add_506_U243  ( .A1(_add_506_n465 ), .A2(_add_506_n466 ), .A3(_add_506_n467 ), .ZN(_add_506_n464 ) );
NAND3_X2 _add_506_U242  ( .A1(n18569), .A2(n18573), .A3(_add_506_n4 ), .ZN(_add_506_n177 ) );
AND3_X4 _add_506_U241  ( .A1(n18121), .A2(n18117), .A3(n18125), .ZN(_add_506_n10 ) );
AND2_X4 _add_506_U240  ( .A1(n18109), .A2(n18113), .ZN(_add_506_n9 ) );
NAND2_X2 _add_506_U239  ( .A1(_add_506_n9 ), .A2(_add_506_n10 ), .ZN(_add_506_n8 ) );
NAND3_X2 _add_506_U238  ( .A1(n18269), .A2(n18273), .A3(n18285), .ZN(_add_506_n109 ) );
NOR2_X2 _add_506_U237  ( .A1(_add_506_n644 ), .A2(_add_506_n645 ), .ZN(_add_506_n640 ) );
NOR2_X2 _add_506_U236  ( .A1(_add_506_n642 ), .A2(_add_506_n643 ), .ZN(_add_506_n641 ) );
NAND3_X2 _add_506_U235  ( .A1(n18369), .A2(n18365), .A3(n18373), .ZN(_add_506_n218 ) );
NAND3_X2 _add_506_U234  ( .A1(n18133), .A2(n18129), .A3(n18137), .ZN(_add_506_n421 ) );
NAND3_X2 _add_506_U233  ( .A1(n18145), .A2(n18149), .A3(n18141), .ZN(_add_506_n420 ) );
NOR2_X2 _add_506_U232  ( .A1(_add_506_n420 ), .A2(_add_506_n421 ), .ZN(_add_506_n419 ) );
NOR2_X2 _add_506_U231  ( .A1(_add_506_n236 ), .A2(_add_506_n237 ), .ZN(_add_506_n232 ) );
NOR2_X2 _add_506_U230  ( .A1(_add_506_n234 ), .A2(_add_506_n235 ), .ZN(_add_506_n233 ) );
NAND3_X2 _add_506_U229  ( .A1(n18541), .A2(_add_506_n2 ), .A3(_add_506_n30 ),.ZN(_add_506_n392 ) );
NOR2_X2 _add_506_U228  ( .A1(_add_506_n331 ), .A2(_add_506_n332 ), .ZN(_add_506_n330 ) );
NOR2_X2 _add_506_U227  ( .A1(_add_506_n333 ), .A2(_add_506_n334 ), .ZN(_add_506_n329 ) );
NOR2_X2 _add_506_U226  ( .A1(_add_506_n324 ), .A2(_add_506_n325 ), .ZN(_add_506_n320 ) );
NOR2_X2 _add_506_U225  ( .A1(_add_506_n322 ), .A2(_add_506_n323 ), .ZN(_add_506_n321 ) );
NOR2_X2 _add_506_U224  ( .A1(_add_506_n282 ), .A2(_add_506_n283 ), .ZN(_add_506_n278 ) );
NOR2_X2 _add_506_U223  ( .A1(_add_506_n280 ), .A2(_add_506_n281 ), .ZN(_add_506_n279 ) );
NOR2_X2 _add_506_U222  ( .A1(_add_506_n605 ), .A2(_add_506_n606 ), .ZN(_add_506_n601 ) );
NOR2_X2 _add_506_U221  ( .A1(_add_506_n603 ), .A2(_add_506_n604 ), .ZN(_add_506_n602 ) );
NOR2_X2 _add_506_U220  ( .A1(_add_506_n535 ), .A2(_add_506_n536 ), .ZN(_add_506_n534 ) );
NOR2_X2 _add_506_U219  ( .A1(_add_506_n537 ), .A2(_add_506_n538 ), .ZN(_add_506_n533 ) );
NAND3_X2 _add_506_U218  ( .A1(n18193), .A2(n18197), .A3(n18189), .ZN(_add_506_n548 ) );
NAND3_X2 _add_506_U217  ( .A1(n18301), .A2(n18313), .A3(n18297), .ZN(_add_506_n133 ) );
NOR3_X2 _add_506_U216  ( .A1(_add_506_n57 ), .A2(_add_506_n133 ), .A3(_add_506_n134 ), .ZN(_add_506_n132 ) );
NOR3_X2 _add_506_U215  ( .A1(_add_506_n23 ), .A2(_add_506_n135 ), .A3(_add_506_n181 ), .ZN(_add_506_n180 ) );
NOR2_X2 _add_506_U214  ( .A1(_add_506_n182 ), .A2(_add_506_n183 ), .ZN(_add_506_n179 ) );
NOR3_X2 _add_506_U213  ( .A1(_add_506_n23 ), .A2(_add_506_n135 ), .A3(_add_506_n174 ), .ZN(_add_506_n173 ) );
NOR2_X2 _add_506_U212  ( .A1(_add_506_n175 ), .A2(_add_506_n176 ), .ZN(_add_506_n172 ) );
NOR3_X2 _add_506_U211  ( .A1(_add_506_n23 ), .A2(_add_506_n135 ), .A3(_add_506_n162 ), .ZN(_add_506_n161 ) );
NOR2_X2 _add_506_U210  ( .A1(_add_506_n163 ), .A2(_add_506_n164 ), .ZN(_add_506_n160 ) );
NOR2_X2 _add_506_U209  ( .A1(_add_506_n25 ), .A2(_add_506_n114 ), .ZN(_add_506_n118 ) );
NOR2_X2 _add_506_U208  ( .A1(_add_506_n25 ), .A2(_add_506_n75 ), .ZN(_add_506_n96 ) );
NOR3_X2 _add_506_U207  ( .A1(_add_506_n412 ), .A2(_add_506_n399 ), .A3(_add_506_n400 ), .ZN(_add_506_n395 ) );
OR3_X4 _add_506_U206  ( .A1(_add_506_n149 ), .A2(_add_506_n150 ), .A3(_add_506_n57 ), .ZN(_add_506_n7 ) );
XNOR2_X2 _add_506_U205  ( .A(n18297), .B(_add_506_n7 ), .ZN(N2100) );
NOR3_X2 _add_506_U204  ( .A1(_add_506_n412 ), .A2(_add_506_n406 ), .A3(_add_506_n407 ), .ZN(_add_506_n403 ) );
NOR2_X2 _add_506_U203  ( .A1(_add_506_n59 ), .A2(_add_506_n463 ), .ZN(_add_506_n462 ) );
NOR2_X2 _add_506_U202  ( .A1(_add_506_n451 ), .A2(_add_506_n468 ), .ZN(_add_506_n461 ) );
NOR2_X2 _add_506_U201  ( .A1(_add_506_n59 ), .A2(_add_506_n445 ), .ZN(_add_506_n444 ) );
NOR2_X2 _add_506_U200  ( .A1(_add_506_n451 ), .A2(_add_506_n452 ), .ZN(_add_506_n443 ) );
NOR3_X2 _add_506_U199  ( .A1(_add_506_n24 ), .A2(_add_506_n37 ), .A3(_add_506_n39 ), .ZN(_add_506_n570 ) );
NOR3_X2 _add_506_U198  ( .A1(_add_506_n572 ), .A2(_add_506_n573 ), .A3(_add_506_n574 ), .ZN(_add_506_n571 ) );
NOR3_X2 _add_506_U197  ( .A1(_add_506_n24 ), .A2(_add_506_n37 ), .A3(_add_506_n39 ), .ZN(_add_506_n560 ) );
NOR3_X2 _add_506_U196  ( .A1(_add_506_n562 ), .A2(_add_506_n563 ), .A3(_add_506_n564 ), .ZN(_add_506_n561 ) );
NOR3_X2 _add_506_U195  ( .A1(_add_506_n286 ), .A2(_add_506_n621 ), .A3(_add_506_n287 ), .ZN(_add_506_n285 ) );
NOR3_X2 _add_506_U194  ( .A1(_add_506_n346 ), .A2(_add_506_n339 ), .A3(_add_506_n607 ), .ZN(_add_506_n345 ) );
NOR3_X2 _add_506_U193  ( .A1(_add_506_n412 ), .A2(_add_506_n413 ), .A3(_add_506_n414 ), .ZN(_add_506_n409 ) );
NOR2_X2 _add_506_U192  ( .A1(_add_506_n483 ), .A2(_add_506_n484 ), .ZN(_add_506_n482 ) );
NOR2_X2 _add_506_U191  ( .A1(_add_506_n135 ), .A2(_add_506_n145 ), .ZN(_add_506_n142 ) );
NOR3_X2 _add_506_U190  ( .A1(_add_506_n146 ), .A2(_add_506_n147 ), .A3(_add_506_n148 ), .ZN(_add_506_n141 ) );
NOR3_X2 _add_506_U189  ( .A1(_add_506_n351 ), .A2(_add_506_n339 ), .A3(_add_506_n607 ), .ZN(_add_506_n350 ) );
NOR3_X2 _add_506_U188  ( .A1(_add_506_n59 ), .A2(_add_506_n23 ), .A3(_add_506_n465 ), .ZN(_add_506_n472 ) );
NOR3_X2 _add_506_U187  ( .A1(_add_506_n473 ), .A2(_add_506_n474 ), .A3(_add_506_n475 ), .ZN(_add_506_n471 ) );
NAND3_X2 _add_506_U186  ( .A1(n18185), .A2(n18181), .A3(n18189), .ZN(_add_506_n585 ) );
NOR3_X2 _add_506_U185  ( .A1(_add_506_n24 ), .A2(_add_506_n584 ), .A3(_add_506_n585 ), .ZN(_add_506_n583 ) );
NOR3_X2 _add_506_U184  ( .A1(_add_506_n23 ), .A2(_add_506_n135 ), .A3(_add_506_n168 ), .ZN(_add_506_n167 ) );
NOR2_X2 _add_506_U183  ( .A1(_add_506_n169 ), .A2(_add_506_n170 ), .ZN(_add_506_n166 ) );
NOR2_X2 _add_506_U182  ( .A1(_add_506_n57 ), .A2(_add_506_n451 ), .ZN(_add_506_n455 ) );
NOR3_X2 _add_506_U181  ( .A1(_add_506_n8 ), .A2(_add_506_n458 ), .A3(_add_506_n459 ), .ZN(_add_506_n454 ) );
NAND3_X2 _add_506_U180  ( .A1(n18525), .A2(n18521), .A3(_add_506_n337 ),.ZN(_add_506_n372 ) );
NAND3_X2 _add_506_U179  ( .A1(n18541), .A2(n18545), .A3(n18537), .ZN(_add_506_n391 ) );
NOR2_X2 _add_506_U178  ( .A1(_add_506_n390 ), .A2(_add_506_n391 ), .ZN(_add_506_n389 ) );
NAND3_X2 _add_506_U177  ( .A1(n18549), .A2(n18553), .A3(n18557), .ZN(_add_506_n386 ) );
NOR2_X2 _add_506_U176  ( .A1(_add_506_n386 ), .A2(_add_506_n387 ), .ZN(_add_506_n385 ) );
NOR2_X2 _add_506_U175  ( .A1(_add_506_n280 ), .A2(_add_506_n621 ), .ZN(_add_506_n309 ) );
NAND3_X2 _add_506_U174  ( .A1(n18509), .A2(_add_506_n362 ), .A3(_add_506_n337 ), .ZN(_add_506_n369 ) );
NOR2_X2 _add_506_U173  ( .A1(_add_506_n122 ), .A2(_add_506_n123 ), .ZN(_add_506_n121 ) );
NOR3_X2 _add_506_U172  ( .A1(_add_506_n24 ), .A2(_add_506_n584 ), .A3(_add_506_n588 ), .ZN(_add_506_n587 ) );
NAND3_X2 _add_506_U171  ( .A1(n18425), .A2(n18421), .A3(n18429), .ZN(_add_506_n273 ) );
NOR3_X2 _add_506_U170  ( .A1(_add_506_n317 ), .A2(_add_506_n318 ), .A3(_add_506_n319 ), .ZN(_add_506_n316 ) );
NOR3_X2 _add_506_U169  ( .A1(_add_506_n326 ), .A2(_add_506_n327 ), .A3(_add_506_n328 ), .ZN(_add_506_n315 ) );
NOR2_X2 _add_506_U168  ( .A1(_add_506_n339 ), .A2(_add_506_n607 ), .ZN(_add_506_n364 ) );
NAND3_X2 _add_506_U167  ( .A1(n18157), .A2(n18153), .A3(_add_506_n398 ),.ZN(_add_506_n411 ) );
NOR2_X2 _add_506_U166  ( .A1(_add_506_n411 ), .A2(_add_506_n57 ), .ZN(_add_506_n410 ) );
NAND3_X2 _add_506_U165  ( .A1(n18549), .A2(_add_506_n3 ), .A3(_add_506_n30 ),.ZN(_add_506_n469 ) );
NOR3_X2 _add_506_U164  ( .A1(_add_506_n621 ), .A2(_add_506_n297 ), .A3(_add_506_n288 ), .ZN(_add_506_n296 ) );
NAND3_X2 _add_506_U163  ( .A1(n18197), .A2(n18193), .A3(n18201), .ZN(_add_506_n564 ) );
NAND3_X2 _add_506_U162  ( .A1(n18093), .A2(n18133), .A3(n18129), .ZN(_add_506_n414 ) );
NAND3_X2 _add_506_U161  ( .A1(n18549), .A2(n18553), .A3(n18557), .ZN(_add_506_n390 ) );
NOR3_X2 _add_506_U160  ( .A1(_add_506_n23 ), .A2(_add_506_n37 ), .A3(_add_506_n42 ), .ZN(_add_506_n41 ) );
NOR2_X2 _add_506_U159  ( .A1(_add_506_n493 ), .A2(_add_506_n501 ), .ZN(_add_506_n499 ) );
NAND3_X2 _add_506_U158  ( .A1(n18377), .A2(n18373), .A3(n18381), .ZN(_add_506_n227 ) );
NOR3_X2 _add_506_U157  ( .A1(_add_506_n24 ), .A2(_add_506_n255 ), .A3(_add_506_n244 ), .ZN(_add_506_n254 ) );
NAND3_X2 _add_506_U156  ( .A1(n18153), .A2(n18149), .A3(n18157), .ZN(_add_506_n515 ) );
NOR2_X2 _add_506_U155  ( .A1(_add_506_n25 ), .A2(_add_506_n515 ), .ZN(_add_506_n514 ) );
NAND3_X2 _add_506_U154  ( .A1(n18317), .A2(n18313), .A3(n18321), .ZN(_add_506_n174 ) );
NOR2_X2 _add_506_U153  ( .A1(_add_506_n135 ), .A2(_add_506_n136 ), .ZN(_add_506_n131 ) );
NOR3_X2 _add_506_U152  ( .A1(_add_506_n137 ), .A2(_add_506_n138 ), .A3(_add_506_n139 ), .ZN(_add_506_n130 ) );
NOR3_X2 _add_506_U151  ( .A1(_add_506_n24 ), .A2(_add_506_n580 ), .A3(_add_506_n581 ), .ZN(_add_506_n576 ) );
NOR3_X2 _add_506_U150  ( .A1(_add_506_n37 ), .A2(_add_506_n578 ), .A3(_add_506_n579 ), .ZN(_add_506_n577 ) );
NOR2_X2 _add_506_U149  ( .A1(_add_506_n607 ), .A2(_add_506_n339 ), .ZN(_add_506_n359 ) );
NOR3_X2 _add_506_U148  ( .A1(_add_506_n24 ), .A2(_add_506_n37 ), .A3(_add_506_n558 ), .ZN(_add_506_n544 ) );
NOR3_X2 _add_506_U147  ( .A1(_add_506_n546 ), .A2(_add_506_n547 ), .A3(_add_506_n548 ), .ZN(_add_506_n545 ) );
NOR2_X2 _add_506_U146  ( .A1(_add_506_n226 ), .A2(_add_506_n227 ), .ZN(_add_506_n222 ) );
NOR2_X2 _add_506_U145  ( .A1(_add_506_n224 ), .A2(_add_506_n225 ), .ZN(_add_506_n223 ) );
NOR3_X2 _add_506_U144  ( .A1(_add_506_n135 ), .A2(_add_506_n12 ), .A3(_add_506_n187 ), .ZN(_add_506_n193 ) );
NOR2_X2 _add_506_U143  ( .A1(_add_506_n194 ), .A2(_add_506_n195 ), .ZN(_add_506_n192 ) );
NOR2_X2 _add_506_U142  ( .A1(_add_506_n621 ), .A2(_add_506_n280 ), .ZN(_add_506_n306 ) );
NOR2_X2 _add_506_U141  ( .A1(_add_506_n272 ), .A2(_add_506_n273 ), .ZN(_add_506_n268 ) );
NOR2_X2 _add_506_U140  ( .A1(_add_506_n270 ), .A2(_add_506_n271 ), .ZN(_add_506_n269 ) );
NOR2_X2 _add_506_U139  ( .A1(_add_506_n25 ), .A2(_add_506_n234 ), .ZN(_add_506_n260 ) );
NOR2_X2 _add_506_U138  ( .A1(_add_506_n236 ), .A2(_add_506_n252 ), .ZN(_add_506_n251 ) );
NOR2_X2 _add_506_U137  ( .A1(_add_506_n248 ), .A2(_add_506_n249 ), .ZN(_add_506_n246 ) );
NOR2_X2 _add_506_U136  ( .A1(_add_506_n243 ), .A2(_add_506_n244 ), .ZN(_add_506_n239 ) );
NOR2_X2 _add_506_U135  ( .A1(_add_506_n241 ), .A2(_add_506_n242 ), .ZN(_add_506_n240 ) );
NOR3_X2 _add_506_U134  ( .A1(_add_506_n135 ), .A2(_add_506_n187 ), .A3(_add_506_n188 ), .ZN(_add_506_n186 ) );
NOR2_X2 _add_506_U133  ( .A1(_add_506_n189 ), .A2(_add_506_n190 ), .ZN(_add_506_n185 ) );
NOR2_X2 _add_506_U132  ( .A1(_add_506_n122 ), .A2(_add_506_n126 ), .ZN(_add_506_n125 ) );
NOR2_X2 _add_506_U131  ( .A1(_add_506_n25 ), .A2(_add_506_n114 ), .ZN(_add_506_n116 ) );
NOR2_X2 _add_506_U130  ( .A1(_add_506_n114 ), .A2(_add_506_n24 ), .ZN(_add_506_n112 ) );
NOR2_X2 _add_506_U129  ( .A1(_add_506_n102 ), .A2(_add_506_n103 ), .ZN(_add_506_n113 ) );
NOR3_X2 _add_506_U128  ( .A1(_add_506_n23 ), .A2(_add_506_n109 ), .A3(_add_506_n110 ), .ZN(_add_506_n107 ) );
NOR2_X2 _add_506_U127  ( .A1(_add_506_n103 ), .A2(_add_506_n104 ), .ZN(_add_506_n108 ) );
NOR2_X2 _add_506_U126  ( .A1(_add_506_n25 ), .A2(_add_506_n75 ), .ZN(_add_506_n94 ) );
NOR2_X2 _add_506_U125  ( .A1(_add_506_n75 ), .A2(_add_506_n25 ), .ZN(_add_506_n90 ) );
NOR2_X2 _add_506_U124  ( .A1(_add_506_n87 ), .A2(_add_506_n92 ), .ZN(_add_506_n91 ) );
NOR2_X2 _add_506_U123  ( .A1(_add_506_n75 ), .A2(_add_506_n25 ), .ZN(_add_506_n85 ) );
NOR2_X2 _add_506_U122  ( .A1(_add_506_n87 ), .A2(_add_506_n88 ), .ZN(_add_506_n86 ) );
NOR2_X2 _add_506_U121  ( .A1(_add_506_n1 ), .A2(_add_506_n81 ), .ZN(_add_506_n80 ) );
NOR3_X2 _add_506_U120  ( .A1(_add_506_n23 ), .A2(_add_506_n75 ), .A3(_add_506_n76 ), .ZN(_add_506_n74 ) );
NOR2_X2 _add_506_U119  ( .A1(_add_506_n67 ), .A2(_add_506_n77 ), .ZN(_add_506_n73 ) );
NOR2_X2 _add_506_U118  ( .A1(_add_506_n69 ), .A2(_add_506_n25 ), .ZN(_add_506_n65 ) );
NOR2_X2 _add_506_U117  ( .A1(_add_506_n67 ), .A2(_add_506_n68 ), .ZN(_add_506_n66 ) );
NOR2_X2 _add_506_U116  ( .A1(_add_506_n52 ), .A2(_add_506_n37 ), .ZN(_add_506_n61 ) );
NOR2_X2 _add_506_U115  ( .A1(_add_506_n37 ), .A2(_add_506_n25 ), .ZN(_add_506_n50 ) );
NOR2_X2 _add_506_U114  ( .A1(_add_506_n52 ), .A2(_add_506_n53 ), .ZN(_add_506_n51 ) );
NOR2_X2 _add_506_U113  ( .A1(_add_506_n37 ), .A2(_add_506_n43 ), .ZN(_add_506_n48 ) );
NOR2_X2 _add_506_U112  ( .A1(_add_506_n39 ), .A2(_add_506_n25 ), .ZN(_add_506_n45 ) );
NOR2_X2 _add_506_U111  ( .A1(_add_506_n37 ), .A2(_add_506_n43 ), .ZN(_add_506_n46 ) );
NOR2_X2 _add_506_U110  ( .A1(_add_506_n1 ), .A2(_add_506_n584 ), .ZN(_add_506_n594 ) );
NOR2_X2 _add_506_U109  ( .A1(_add_506_n1 ), .A2(_add_506_n591 ), .ZN(_add_506_n590 ) );
NAND3_X2 _add_506_U108  ( .A1(n18321), .A2(n18317), .A3(n18325), .ZN(_add_506_n181 ) );
NAND3_X2 _add_506_U107  ( .A1(n18133), .A2(n18141), .A3(n18129), .ZN(_add_506_n458 ) );
NOR2_X2 _add_506_U106  ( .A1(_add_506_n57 ), .A2(_add_506_n59 ), .ZN(_add_506_n504 ) );
NOR3_X2 _add_506_U105  ( .A1(_add_506_n505 ), .A2(_add_506_n493 ), .A3(_add_506_n494 ), .ZN(_add_506_n503 ) );
NAND3_X2 _add_506_U104  ( .A1(n18321), .A2(n18317), .A3(n18325), .ZN(_add_506_n636 ) );
NOR2_X2 _add_506_U103  ( .A1(_add_506_n635 ), .A2(_add_506_n636 ), .ZN(_add_506_n628 ) );
NOR2_X2 _add_506_U102  ( .A1(_add_506_n621 ), .A2(_add_506_n622 ), .ZN(_add_506_n620 ) );
NAND3_X2 _add_506_U101  ( .A1(n18377), .A2(n18373), .A3(n18381), .ZN(_add_506_n632 ) );
NOR2_X2 _add_506_U100  ( .A1(_add_506_n631 ), .A2(_add_506_n632 ), .ZN(_add_506_n630 ) );
NAND3_X2 _add_506_U99  ( .A1(n18293), .A2(n18289), .A3(n18297), .ZN(_add_506_n638 ) );
NOR2_X2 _add_506_U98  ( .A1(_add_506_n637 ), .A2(_add_506_n638 ), .ZN(_add_506_n627 ) );
NOR3_X2 _add_506_U97  ( .A1(_add_506_n422 ), .A2(_add_506_n423 ), .A3(_add_506_n424 ), .ZN(_add_506_n401 ) );
NOR3_X2 _add_506_U96  ( .A1(_add_506_n520 ), .A2(_add_506_n521 ), .A3(_add_506_n522 ), .ZN(_add_506_n30 ) );
NOR2_X2 _add_506_U95  ( .A1(_add_506_n633 ), .A2(_add_506_n634 ), .ZN(_add_506_n629 ) );
NAND4_X2 _add_506_U94  ( .A1(_add_506_n627 ), .A2(_add_506_n628 ), .A3(_add_506_n629 ), .A4(_add_506_n630 ), .ZN(_add_506_n59 ) );
NAND3_X2 _add_506_U93  ( .A1(n18333), .A2(n18337), .A3(n18349), .ZN(_add_506_n194 ) );
NAND3_X2 _add_506_U92  ( .A1(n18345), .A2(n18341), .A3(n18349), .ZN(_add_506_n189 ) );
NAND3_X2 _add_506_U91  ( .A1(n18345), .A2(n18341), .A3(n18349), .ZN(_add_506_n182 ) );
NAND3_X2 _add_506_U90  ( .A1(n18329), .A2(n18337), .A3(n18333), .ZN(_add_506_n190 ) );
NAND3_X2 _add_506_U89  ( .A1(n18329), .A2(n18337), .A3(n18333), .ZN(_add_506_n183 ) );
NAND3_X2 _add_506_U88  ( .A1(n18329), .A2(n18325), .A3(n18333), .ZN(_add_506_n176 ) );
NAND3_X2 _add_506_U87  ( .A1(n18329), .A2(n18325), .A3(n18333), .ZN(_add_506_n170 ) );
NAND3_X2 _add_506_U86  ( .A1(n18333), .A2(n18337), .A3(n18349), .ZN(_add_506_n147 ) );
NAND3_X2 _add_506_U85  ( .A1(n18333), .A2(n18337), .A3(n18349), .ZN(_add_506_n138 ) );
NOR2_X2 _add_506_U84  ( .A1(_add_506_n646 ), .A2(_add_506_n647 ), .ZN(_add_506_n639 ) );
NAND3_X2 _add_506_U83  ( .A1(_add_506_n639 ), .A2(_add_506_n640 ), .A3(_add_506_n641 ), .ZN(_add_506_n37 ) );
NOR2_X2 _add_506_U82  ( .A1(_add_506_n25 ), .A2(_add_506_n465 ), .ZN(_add_506_n479 ) );
NOR2_X2 _add_506_U81  ( .A1(_add_506_n135 ), .A2(_add_506_n154 ), .ZN(_add_506_n153 ) );
NOR2_X2 _add_506_U80  ( .A1(_add_506_n157 ), .A2(_add_506_n158 ), .ZN(_add_506_n151 ) );
NOR2_X2 _add_506_U79  ( .A1(_add_506_n155 ), .A2(_add_506_n156 ), .ZN(_add_506_n152 ) );
NOR2_X2 _add_506_U78  ( .A1(_add_506_n33 ), .A2(_add_506_n34 ), .ZN(_add_506_n32 ) );
NOR2_X2 _add_506_U77  ( .A1(_add_506_n491 ), .A2(_add_506_n492 ), .ZN(_add_506_n490 ) );
NOR2_X2 _add_506_U76  ( .A1(_add_506_n493 ), .A2(_add_506_n494 ), .ZN(_add_506_n489 ) );
NOR2_X2 _add_506_U75  ( .A1(_add_506_n495 ), .A2(_add_506_n14 ), .ZN(_add_506_n488 ) );
NAND3_X2 _add_506_U74  ( .A1(_add_506_n488 ), .A2(_add_506_n489 ), .A3(_add_506_n490 ), .ZN(_add_506_n474 ) );
NOR2_X2 _add_506_U73  ( .A1(_add_506_n218 ), .A2(_add_506_n219 ), .ZN(_add_506_n214 ) );
NAND2_X2 _add_506_U72  ( .A1(_add_506_n214 ), .A2(_add_506_n215 ), .ZN(_add_506_n135 ) );
NOR2_X2 _add_506_U71  ( .A1(_add_506_n135 ), .A2(_add_506_n24 ), .ZN(_add_506_n213 ) );
NAND3_X2 _add_506_U70  ( .A1(n18345), .A2(n18341), .A3(n18349), .ZN(_add_506_n206 ) );
NOR3_X2 _add_506_U69  ( .A1(_add_506_n24 ), .A2(_add_506_n135 ), .A3(_add_506_n206 ), .ZN(_add_506_n205 ) );
NOR3_X2 _add_506_U68  ( .A1(_add_506_n23 ), .A2(_add_506_n209 ), .A3(_add_506_n135 ), .ZN(_add_506_n208 ) );
NOR3_X2 _add_506_U67  ( .A1(_add_506_n23 ), .A2(_add_506_n135 ), .A3(_add_506_n199 ), .ZN(_add_506_n203 ) );
NOR2_X2 _add_506_U66  ( .A1(_add_506_n505 ), .A2(_add_506_n493 ), .ZN(_add_506_n509 ) );
NOR2_X2 _add_506_U65  ( .A1(_add_506_n378 ), .A2(_add_506_n379 ), .ZN(_add_506_n377 ) );
NOR2_X2 _add_506_U64  ( .A1(_add_506_n380 ), .A2(_add_506_n381 ), .ZN(_add_506_n376 ) );
NOR2_X2 _add_506_U63  ( .A1(_add_506_n382 ), .A2(_add_506_n383 ), .ZN(_add_506_n375 ) );
NAND3_X2 _add_506_U62  ( .A1(_add_506_n375 ), .A2(_add_506_n376 ), .A3(_add_506_n377 ), .ZN(_add_506_n374 ) );
NOR2_X2 _add_506_U61  ( .A1(_add_506_n427 ), .A2(_add_506_n13 ), .ZN(_add_506_n426 ) );
NOR2_X2 _add_506_U60  ( .A1(_add_506_n447 ), .A2(_add_506_n434 ), .ZN(_add_506_n446 ) );
NOR2_X2 _add_506_U59  ( .A1(_add_506_n433 ), .A2(_add_506_n434 ), .ZN(_add_506_n432 ) );
NOR2_X2 _add_506_U58  ( .A1(_add_506_n614 ), .A2(_add_506_n615 ), .ZN(_add_506_n613 ) );
NOR2_X2 _add_506_U57  ( .A1(_add_506_n39 ), .A2(_add_506_n616 ), .ZN(_add_506_n612 ) );
NOR2_X2 _add_506_U56  ( .A1(_add_506_n617 ), .A2(_add_506_n31 ), .ZN(_add_506_n611 ) );
NAND3_X2 _add_506_U55  ( .A1(_add_506_n611 ), .A2(_add_506_n612 ), .A3(_add_506_n613 ), .ZN(_add_506_n584 ) );
NOR3_X2 _add_506_U54  ( .A1(_add_506_n23 ), .A2(_add_506_n199 ), .A3(_add_506_n135 ), .ZN(_add_506_n198 ) );
NOR2_X2 _add_506_U53  ( .A1(_add_506_n11 ), .A2(_add_506_n12 ), .ZN(_add_506_n197 ) );
NOR2_X2 _add_506_U52  ( .A1(_add_506_n623 ), .A2(_add_506_n624 ), .ZN(_add_506_n619 ) );
NOR2_X2 _add_506_U51  ( .A1(_add_506_n625 ), .A2(_add_506_n626 ), .ZN(_add_506_n618 ) );
NOR2_X2 _add_506_U50  ( .A1(_add_506_n135 ), .A2(_add_506_n199 ), .ZN(_add_506_n201 ) );
NOR2_X2 _add_506_U49  ( .A1(_add_506_n25 ), .A2(_add_506_n498 ), .ZN(_add_506_n497 ) );
OR2_X4 _add_506_U48  ( .A1(_add_506_n516 ), .A2(_add_506_n517 ), .ZN(_add_506_n6 ) );
XNOR2_X2 _add_506_U47  ( .A(n18149), .B(_add_506_n6 ), .ZN(N2137) );
NOR2_X2 _add_506_U46  ( .A1(_add_506_n477 ), .A2(_add_506_n478 ), .ZN(_add_506_n476 ) );
NOR2_X2 _add_506_U45  ( .A1(_add_506_n486 ), .A2(_add_506_n487 ), .ZN(_add_506_n485 ) );
NOR2_X2 _add_506_U44  ( .A1(_add_506_n507 ), .A2(_add_506_n508 ), .ZN(_add_506_n506 ) );
NOR2_X2 _add_506_U43  ( .A1(_add_506_n524 ), .A2(_add_506_n525 ), .ZN(_add_506_n523 ) );
NOR2_X2 _add_506_U42  ( .A1(_add_506_n511 ), .A2(_add_506_n512 ), .ZN(_add_506_n510 ) );
NOR3_X2 _add_506_U41  ( .A1(_add_506_n530 ), .A2(_add_506_n531 ), .A3(_add_506_n532 ), .ZN(_add_506_n529 ) );
NOR2_X2 _add_506_U40  ( .A1(_add_506_n541 ), .A2(_add_506_n542 ), .ZN(_add_506_n527 ) );
NOR2_X2 _add_506_U39  ( .A1(_add_506_n539 ), .A2(_add_506_n540 ), .ZN(_add_506_n528 ) );
NAND3_X2 _add_506_U38  ( .A1(_add_506_n527 ), .A2(_add_506_n528 ), .A3(_add_506_n529 ), .ZN(_add_506_n451 ) );
NOR2_X2 _add_506_U37  ( .A1(_add_506_n427 ), .A2(_add_506_n13 ), .ZN(_add_506_n518 ) );
NOR2_X2 _add_506_U36  ( .A1(_add_506_n100 ), .A2(_add_506_n101 ), .ZN(_add_506_n99 ) );
NOR2_X2 _add_506_U35  ( .A1(_add_506_n102 ), .A2(_add_506_n103 ), .ZN(_add_506_n98 ) );
NOR2_X2 _add_506_U34  ( .A1(_add_506_n104 ), .A2(_add_506_n105 ), .ZN(_add_506_n97 ) );
NAND3_X2 _add_506_U33  ( .A1(_add_506_n97 ), .A2(_add_506_n98 ), .A3(_add_506_n99 ), .ZN(_add_506_n75 ) );
NOR2_X2 _add_506_U32  ( .A1(_add_506_n568 ), .A2(_add_506_n552 ), .ZN(_add_506_n567 ) );
NOR2_X2 _add_506_U31  ( .A1(_add_506_n553 ), .A2(_add_506_n554 ), .ZN(_add_506_n566 ) );
NOR2_X2 _add_506_U30  ( .A1(_add_506_n555 ), .A2(_add_506_n556 ), .ZN(_add_506_n565 ) );
NOR2_X2 _add_506_U29  ( .A1(_add_506_n552 ), .A2(_add_506_n553 ), .ZN(_add_506_n551 ) );
NOR2_X2 _add_506_U28  ( .A1(_add_506_n554 ), .A2(_add_506_n555 ), .ZN(_add_506_n550 ) );
NOR2_X2 _add_506_U27  ( .A1(_add_506_n556 ), .A2(_add_506_n557 ), .ZN(_add_506_n549 ) );
NOR3_X2 _add_506_U26  ( .A1(_add_506_n598 ), .A2(_add_506_n599 ), .A3(_add_506_n600 ), .ZN(_add_506_n597 ) );
NOR2_X2 _add_506_U25  ( .A1(_add_506_n607 ), .A2(_add_506_n608 ), .ZN(_add_506_n596 ) );
NOR2_X2 _add_506_U24  ( .A1(_add_506_n609 ), .A2(_add_506_n610 ), .ZN(_add_506_n595 ) );
NAND3_X2 _add_506_U23  ( .A1(_add_506_n595 ), .A2(_add_506_n596 ), .A3(_add_506_n597 ), .ZN(_add_506_n57 ) );
INV_X4 _add_506_U22  ( .A(_add_506_n1 ), .ZN(_add_506_n28 ) );
INV_X4 _add_506_U21  ( .A(_add_506_n374 ), .ZN(_add_506_n337 ) );
INV_X4 _add_506_U20  ( .A(_add_506_n451 ), .ZN(_add_506_n398 ) );
INV_X4 _add_506_U19  ( .A(_add_506_n57 ), .ZN(_add_506_n15 ) );
INV_X4 _add_506_U18  ( .A(_add_506_n59 ), .ZN(_add_506_n19 ) );
INV_X4 _add_506_U17  ( .A(_add_506_n1 ), .ZN(_add_506_n27 ) );
INV_X4 _add_506_U16  ( .A(_add_506_n1 ), .ZN(_add_506_n26 ) );
INV_X4 _add_506_U15  ( .A(_add_506_n59 ), .ZN(_add_506_n22 ) );
INV_X4 _add_506_U14  ( .A(_add_506_n57 ), .ZN(_add_506_n18 ) );
INV_X4 _add_506_U13  ( .A(_add_506_n59 ), .ZN(_add_506_n21 ) );
INV_X4 _add_506_U12  ( .A(_add_506_n59 ), .ZN(_add_506_n20 ) );
INV_X4 _add_506_U11  ( .A(_add_506_n28 ), .ZN(_add_506_n25 ) );
INV_X4 _add_506_U10  ( .A(_add_506_n28 ), .ZN(_add_506_n24 ) );
INV_X4 _add_506_U9  ( .A(_add_506_n26 ), .ZN(_add_506_n23 ) );
INV_X4 _add_506_U8  ( .A(_add_506_n57 ), .ZN(_add_506_n16 ) );
INV_X4 _add_506_U7  ( .A(_add_506_n57 ), .ZN(_add_506_n17 ) );
XOR2_X2 _add_506_U6  ( .A(n18585), .B(n18589), .Z(N2028) );
AND4_X4 _add_506_U5  ( .A1(n18577), .A2(n18581), .A3(n18585), .A4(n18589),.ZN(_add_506_n4 ) );
AND2_X4 _add_506_U4  ( .A1(n18553), .A2(n18557), .ZN(_add_506_n3 ) );
AND4_X4 _add_506_U3  ( .A1(n18545), .A2(n18549), .A3(n18553), .A4(n18557),.ZN(_add_506_n2 ) );
NAND3_X2 _add_506_U2  ( .A1(_add_506_n618 ), .A2(_add_506_n619 ), .A3(_add_506_n620 ), .ZN(_add_506_n1 ) );
NAND2_X2 _add_1_root_add_519_2_U289  ( .A1(n17750), .A2(aad_byte_cnt[0]),.ZN(_add_1_root_add_519_2_n185 ) );
NAND2_X2 _add_1_root_add_519_2_U288  ( .A1(_add_1_root_add_519_2_n185 ),.A2(_add_1_root_add_519_2_n210 ), .ZN(N2479) );
INV_X4 _add_1_root_add_519_2_U287  ( .A(aad_byte_cnt[7]), .ZN(_add_1_root_add_519_2_n224 ) );
INV_X4 _add_1_root_add_519_2_U286  ( .A(_add_1_root_add_519_2_n198 ), .ZN(_add_1_root_add_519_2_n194 ) );
NAND2_X2 _add_1_root_add_519_2_U285  ( .A1(_add_1_root_add_519_2_n219 ),.A2(_add_1_root_add_519_2_n220 ), .ZN(_add_1_root_add_519_2_n214 ) );
NAND2_X2 _add_1_root_add_519_2_U284  ( .A1(dii_data_size[2]), .A2(aad_byte_cnt[2]), .ZN(_add_1_root_add_519_2_n142 ) );
INV_X4 _add_1_root_add_519_2_U283  ( .A(_add_1_root_add_519_2_n142 ), .ZN(_add_1_root_add_519_2_n217 ) );
NAND2_X2 _add_1_root_add_519_2_U282  ( .A1(n18074), .A2(aad_byte_cnt[3]),.ZN(_add_1_root_add_519_2_n139 ) );
INV_X4 _add_1_root_add_519_2_U281  ( .A(_add_1_root_add_519_2_n139 ), .ZN(_add_1_root_add_519_2_n218 ) );
INV_X4 _add_1_root_add_519_2_U280  ( .A(aad_byte_cnt[3]), .ZN(_add_1_root_add_519_2_n213 ) );
NAND2_X2 _add_1_root_add_519_2_U279  ( .A1(_add_1_root_add_519_2_n61 ), .A2(_add_1_root_add_519_2_n213 ), .ZN(_add_1_root_add_519_2_n140 ) );
NAND2_X2 _add_1_root_add_519_2_U278  ( .A1(_add_1_root_add_519_2_n193 ),.A2(_add_1_root_add_519_2_n140 ), .ZN(_add_1_root_add_519_2_n209 ) );
INV_X4 _add_1_root_add_519_2_U277  ( .A(_add_1_root_add_519_2_n140 ), .ZN(_add_1_root_add_519_2_n212 ) );
NAND2_X2 _add_1_root_add_519_2_U276  ( .A1(_add_1_root_add_519_2_n209 ),.A2(_add_1_root_add_519_2_n200 ), .ZN(_add_1_root_add_519_2_n80 ) );
NAND2_X2 _add_1_root_add_519_2_U275  ( .A1(_add_1_root_add_519_2_n194 ),.A2(_add_1_root_add_519_2_n80 ), .ZN(_add_1_root_add_519_2_n208 ) );
XNOR2_X2 _add_1_root_add_519_2_U274  ( .A(_add_1_root_add_519_2_n59 ), .B(aad_byte_cnt[10]), .ZN(N2489) );
INV_X4 _add_1_root_add_519_2_U273  ( .A(aad_byte_cnt[11]), .ZN(_add_1_root_add_519_2_n207 ) );
XNOR2_X2 _add_1_root_add_519_2_U272  ( .A(_add_1_root_add_519_2_n32 ), .B(aad_byte_cnt[11]), .ZN(N2490) );
INV_X4 _add_1_root_add_519_2_U271  ( .A(aad_byte_cnt[12]), .ZN(_add_1_root_add_519_2_n204 ) );
XNOR2_X2 _add_1_root_add_519_2_U270  ( .A(_add_1_root_add_519_2_n5 ), .B(_add_1_root_add_519_2_n204 ), .ZN(N2491) );
INV_X4 _add_1_root_add_519_2_U269  ( .A(aad_byte_cnt[13]), .ZN(_add_1_root_add_519_2_n203 ) );
XNOR2_X2 _add_1_root_add_519_2_U268  ( .A(_add_1_root_add_519_2_n6 ), .B(_add_1_root_add_519_2_n203 ), .ZN(N2492) );
INV_X4 _add_1_root_add_519_2_U267  ( .A(aad_byte_cnt[14]), .ZN(_add_1_root_add_519_2_n202 ) );
XNOR2_X2 _add_1_root_add_519_2_U266  ( .A(_add_1_root_add_519_2_n9 ), .B(_add_1_root_add_519_2_n202 ), .ZN(N2493) );
INV_X4 _add_1_root_add_519_2_U265  ( .A(aad_byte_cnt[15]), .ZN(_add_1_root_add_519_2_n201 ) );
XNOR2_X2 _add_1_root_add_519_2_U264  ( .A(_add_1_root_add_519_2_n30 ), .B(_add_1_root_add_519_2_n201 ), .ZN(N2494) );
NAND2_X2 _add_1_root_add_519_2_U263  ( .A1(_add_1_root_add_519_2_n196 ),.A2(_add_1_root_add_519_2_n197 ), .ZN(_add_1_root_add_519_2_n195 ) );
XNOR2_X2 _add_1_root_add_519_2_U262  ( .A(_add_1_root_add_519_2_n152 ), .B(aad_byte_cnt[16]), .ZN(N2495) );
XNOR2_X2 _add_1_root_add_519_2_U261  ( .A(_add_1_root_add_519_2_n189 ), .B(_add_1_root_add_519_2_n4 ), .ZN(N2496) );
NAND2_X2 _add_1_root_add_519_2_U260  ( .A1(_add_1_root_add_519_2_n4 ), .A2(aad_byte_cnt[17]), .ZN(_add_1_root_add_519_2_n188 ) );
XNOR2_X2 _add_1_root_add_519_2_U259  ( .A(_add_1_root_add_519_2_n188 ), .B(aad_byte_cnt[18]), .ZN(N2497) );
INV_X4 _add_1_root_add_519_2_U258  ( .A(aad_byte_cnt[19]), .ZN(_add_1_root_add_519_2_n187 ) );
XNOR2_X2 _add_1_root_add_519_2_U257  ( .A(_add_1_root_add_519_2_n40 ), .B(aad_byte_cnt[19]), .ZN(N2498) );
NAND2_X2 _add_1_root_add_519_2_U256  ( .A1(dii_data_size[1]), .A2(aad_byte_cnt[1]), .ZN(_add_1_root_add_519_2_n164 ) );
INV_X4 _add_1_root_add_519_2_U255  ( .A(_add_1_root_add_519_2_n164 ), .ZN(_add_1_root_add_519_2_n184 ) );
XNOR2_X2 _add_1_root_add_519_2_U254  ( .A(_add_1_root_add_519_2_n166 ), .B(_add_1_root_add_519_2_n183 ), .ZN(N2480) );
INV_X4 _add_1_root_add_519_2_U253  ( .A(_add_1_root_add_519_2_n45 ), .ZN(_add_1_root_add_519_2_n178 ) );
XNOR2_X2 _add_1_root_add_519_2_U252  ( .A(_add_1_root_add_519_2_n179 ), .B(_add_1_root_add_519_2_n178 ), .ZN(N2499) );
NAND2_X2 _add_1_root_add_519_2_U251  ( .A1(_add_1_root_add_519_2_n178 ),.A2(aad_byte_cnt[20]), .ZN(_add_1_root_add_519_2_n177 ) );
XNOR2_X2 _add_1_root_add_519_2_U250  ( .A(_add_1_root_add_519_2_n177 ), .B(aad_byte_cnt[21]), .ZN(N2500) );
XNOR2_X2 _add_1_root_add_519_2_U249  ( .A(_add_1_root_add_519_2_n52 ), .B(aad_byte_cnt[22]), .ZN(N2501) );
XNOR2_X2 _add_1_root_add_519_2_U248  ( .A(_add_1_root_add_519_2_n27 ), .B(aad_byte_cnt[23]), .ZN(N2502) );
XNOR2_X2 _add_1_root_add_519_2_U247  ( .A(_add_1_root_add_519_2_n43 ), .B(aad_byte_cnt[24]), .ZN(N2503) );
XNOR2_X2 _add_1_root_add_519_2_U246  ( .A(_add_1_root_add_519_2_n50 ), .B(aad_byte_cnt[25]), .ZN(N2504) );
XNOR2_X2 _add_1_root_add_519_2_U245  ( .A(_add_1_root_add_519_2_n51 ), .B(aad_byte_cnt[26]), .ZN(N2505) );
INV_X4 _add_1_root_add_519_2_U244  ( .A(aad_byte_cnt[27]), .ZN(_add_1_root_add_519_2_n172 ) );
XNOR2_X2 _add_1_root_add_519_2_U243  ( .A(_add_1_root_add_519_2_n28 ), .B(aad_byte_cnt[27]), .ZN(N2506) );
INV_X4 _add_1_root_add_519_2_U242  ( .A(aad_byte_cnt[28]), .ZN(_add_1_root_add_519_2_n159 ) );
XNOR2_X2 _add_1_root_add_519_2_U241  ( .A(_add_1_root_add_519_2_n47 ), .B(aad_byte_cnt[28]), .ZN(N2507) );
INV_X4 _add_1_root_add_519_2_U240  ( .A(aad_byte_cnt[29]), .ZN(_add_1_root_add_519_2_n167 ) );
XNOR2_X2 _add_1_root_add_519_2_U239  ( .A(_add_1_root_add_519_2_n21 ), .B(aad_byte_cnt[29]), .ZN(N2508) );
NAND2_X2 _add_1_root_add_519_2_U238  ( .A1(_add_1_root_add_519_2_n60 ), .A2(_add_1_root_add_519_2_n142 ), .ZN(_add_1_root_add_519_2_n163 ) );
NAND2_X2 _add_1_root_add_519_2_U237  ( .A1(_add_1_root_add_519_2_n57 ), .A2(_add_1_root_add_519_2_n164 ), .ZN(_add_1_root_add_519_2_n143 ) );
INV_X4 _add_1_root_add_519_2_U236  ( .A(_add_1_root_add_519_2_n53 ), .ZN(_add_1_root_add_519_2_n161 ) );
INV_X4 _add_1_root_add_519_2_U235  ( .A(aad_byte_cnt[30]), .ZN(_add_1_root_add_519_2_n162 ) );
XNOR2_X2 _add_1_root_add_519_2_U234  ( .A(_add_1_root_add_519_2_n161 ), .B(_add_1_root_add_519_2_n162 ), .ZN(N2509) );
INV_X4 _add_1_root_add_519_2_U233  ( .A(aad_byte_cnt[31]), .ZN(_add_1_root_add_519_2_n160 ) );
XNOR2_X2 _add_1_root_add_519_2_U232  ( .A(_add_1_root_add_519_2_n17 ), .B(_add_1_root_add_519_2_n160 ), .ZN(N2510) );
INV_X4 _add_1_root_add_519_2_U231  ( .A(_add_1_root_add_519_2_n93 ), .ZN(_add_1_root_add_519_2_n148 ) );
INV_X4 _add_1_root_add_519_2_U230  ( .A(_add_1_root_add_519_2_n94 ), .ZN(_add_1_root_add_519_2_n147 ) );
NAND2_X2 _add_1_root_add_519_2_U229  ( .A1(_add_1_root_add_519_2_n148 ),.A2(_add_1_root_add_519_2_n147 ), .ZN(_add_1_root_add_519_2_n107 ) );
XNOR2_X2 _add_1_root_add_519_2_U228  ( .A(_add_1_root_add_519_2_n157 ), .B(aad_byte_cnt[32]), .ZN(N2511) );
XNOR2_X2 _add_1_root_add_519_2_U227  ( .A(_add_1_root_add_519_2_n34 ), .B(_add_1_root_add_519_2_n151 ), .ZN(N2512) );
XNOR2_X2 _add_1_root_add_519_2_U226  ( .A(_add_1_root_add_519_2_n3 ), .B(_add_1_root_add_519_2_n150 ), .ZN(N2513) );
INV_X4 _add_1_root_add_519_2_U225  ( .A(aad_byte_cnt[35]), .ZN(_add_1_root_add_519_2_n154 ) );
XNOR2_X2 _add_1_root_add_519_2_U224  ( .A(_add_1_root_add_519_2_n7 ), .B(_add_1_root_add_519_2_n154 ), .ZN(N2514) );
NAND2_X2 _add_1_root_add_519_2_U223  ( .A1(_add_1_root_add_519_2_n148 ),.A2(_add_1_root_add_519_2_n8 ), .ZN(_add_1_root_add_519_2_n145 ) );
INV_X4 _add_1_root_add_519_2_U222  ( .A(_add_1_root_add_519_2_n108 ), .ZN(_add_1_root_add_519_2_n78 ) );
NAND2_X2 _add_1_root_add_519_2_U221  ( .A1(_add_1_root_add_519_2_n78 ), .A2(_add_1_root_add_519_2_n147 ), .ZN(_add_1_root_add_519_2_n146 ) );
XNOR2_X2 _add_1_root_add_519_2_U220  ( .A(_add_1_root_add_519_2_n2 ), .B(aad_byte_cnt[36]), .ZN(N2515) );
XNOR2_X2 _add_1_root_add_519_2_U219  ( .A(_add_1_root_add_519_2_n39 ), .B(aad_byte_cnt[37]), .ZN(N2516) );
XNOR2_X2 _add_1_root_add_519_2_U218  ( .A(_add_1_root_add_519_2_n54 ), .B(aad_byte_cnt[38]), .ZN(N2517) );
INV_X4 _add_1_root_add_519_2_U217  ( .A(aad_byte_cnt[39]), .ZN(_add_1_root_add_519_2_n144 ) );
XNOR2_X2 _add_1_root_add_519_2_U216  ( .A(_add_1_root_add_519_2_n38 ), .B(aad_byte_cnt[39]), .ZN(N2518) );
NAND2_X2 _add_1_root_add_519_2_U215  ( .A1(_add_1_root_add_519_2_n143 ),.A2(_add_1_root_add_519_2_n60 ), .ZN(_add_1_root_add_519_2_n141 ) );
NAND2_X2 _add_1_root_add_519_2_U214  ( .A1(_add_1_root_add_519_2_n141 ),.A2(_add_1_root_add_519_2_n142 ), .ZN(_add_1_root_add_519_2_n137 ) );
NAND2_X2 _add_1_root_add_519_2_U213  ( .A1(_add_1_root_add_519_2_n139 ),.A2(_add_1_root_add_519_2_n140 ), .ZN(_add_1_root_add_519_2_n138 ) );
XNOR2_X2 _add_1_root_add_519_2_U212  ( .A(_add_1_root_add_519_2_n137 ), .B(_add_1_root_add_519_2_n138 ), .ZN(N2482) );
INV_X4 _add_1_root_add_519_2_U211  ( .A(_add_1_root_add_519_2_n111 ), .ZN(_add_1_root_add_519_2_n132 ) );
NAND2_X2 _add_1_root_add_519_2_U210  ( .A1(_add_1_root_add_519_2_n132 ),.A2(_add_1_root_add_519_2_n8 ), .ZN(_add_1_root_add_519_2_n131 ) );
XNOR2_X2 _add_1_root_add_519_2_U209  ( .A(_add_1_root_add_519_2_n24 ), .B(aad_byte_cnt[40]), .ZN(N2519) );
INV_X4 _add_1_root_add_519_2_U208  ( .A(_add_1_root_add_519_2_n131 ), .ZN(_add_1_root_add_519_2_n124 ) );
NAND2_X2 _add_1_root_add_519_2_U207  ( .A1(_add_1_root_add_519_2_n124 ),.A2(aad_byte_cnt[40]), .ZN(_add_1_root_add_519_2_n130 ) );
XNOR2_X2 _add_1_root_add_519_2_U206  ( .A(_add_1_root_add_519_2_n23 ), .B(aad_byte_cnt[41]), .ZN(N2520) );
INV_X4 _add_1_root_add_519_2_U205  ( .A(_add_1_root_add_519_2_n130 ), .ZN(_add_1_root_add_519_2_n129 ) );
XNOR2_X2 _add_1_root_add_519_2_U204  ( .A(_add_1_root_add_519_2_n128 ), .B(aad_byte_cnt[42]), .ZN(N2521) );
INV_X4 _add_1_root_add_519_2_U203  ( .A(aad_byte_cnt[43]), .ZN(_add_1_root_add_519_2_n126 ) );
XNOR2_X2 _add_1_root_add_519_2_U202  ( .A(_add_1_root_add_519_2_n26 ), .B(_add_1_root_add_519_2_n126 ), .ZN(N2522) );
NAND4_X2 _add_1_root_add_519_2_U201  ( .A1(aad_byte_cnt[43]), .A2(aad_byte_cnt[42]), .A3(aad_byte_cnt[40]), .A4(aad_byte_cnt[41]), .ZN(_add_1_root_add_519_2_n112 ) );
INV_X4 _add_1_root_add_519_2_U200  ( .A(_add_1_root_add_519_2_n112 ), .ZN(_add_1_root_add_519_2_n125 ) );
NAND2_X2 _add_1_root_add_519_2_U199  ( .A1(_add_1_root_add_519_2_n124 ),.A2(_add_1_root_add_519_2_n125 ), .ZN(_add_1_root_add_519_2_n122 ) );
INV_X4 _add_1_root_add_519_2_U198  ( .A(aad_byte_cnt[44]), .ZN(_add_1_root_add_519_2_n123 ) );
XNOR2_X2 _add_1_root_add_519_2_U197  ( .A(_add_1_root_add_519_2_n36 ), .B(aad_byte_cnt[44]), .ZN(N2523) );
INV_X4 _add_1_root_add_519_2_U196  ( .A(_add_1_root_add_519_2_n122 ), .ZN(_add_1_root_add_519_2_n121 ) );
NAND2_X2 _add_1_root_add_519_2_U195  ( .A1(_add_1_root_add_519_2_n121 ),.A2(aad_byte_cnt[44]), .ZN(_add_1_root_add_519_2_n119 ) );
INV_X4 _add_1_root_add_519_2_U194  ( .A(aad_byte_cnt[45]), .ZN(_add_1_root_add_519_2_n120 ) );
XNOR2_X2 _add_1_root_add_519_2_U193  ( .A(_add_1_root_add_519_2_n22 ), .B(aad_byte_cnt[45]), .ZN(N2524) );
INV_X4 _add_1_root_add_519_2_U192  ( .A(_add_1_root_add_519_2_n119 ), .ZN(_add_1_root_add_519_2_n118 ) );
INV_X4 _add_1_root_add_519_2_U191  ( .A(aad_byte_cnt[46]), .ZN(_add_1_root_add_519_2_n117 ) );
XNOR2_X2 _add_1_root_add_519_2_U190  ( .A(_add_1_root_add_519_2_n116 ), .B(_add_1_root_add_519_2_n117 ), .ZN(N2525) );
INV_X4 _add_1_root_add_519_2_U189  ( .A(aad_byte_cnt[47]), .ZN(_add_1_root_add_519_2_n115 ) );
XNOR2_X2 _add_1_root_add_519_2_U188  ( .A(_add_1_root_add_519_2_n25 ), .B(_add_1_root_add_519_2_n115 ), .ZN(N2526) );
NAND2_X2 _add_1_root_add_519_2_U187  ( .A1(aad_byte_cnt[47]), .A2(aad_byte_cnt[46]), .ZN(_add_1_root_add_519_2_n113 ) );
XNOR2_X2 _add_1_root_add_519_2_U186  ( .A(_add_1_root_add_519_2_n20 ), .B(aad_byte_cnt[48]), .ZN(N2527) );
INV_X4 _add_1_root_add_519_2_U185  ( .A(_add_1_root_add_519_2_n105 ), .ZN(_add_1_root_add_519_2_n92 ) );
INV_X4 _add_1_root_add_519_2_U184  ( .A(_add_1_root_add_519_2_n55 ), .ZN(_add_1_root_add_519_2_n104 ) );
XNOR2_X2 _add_1_root_add_519_2_U183  ( .A(_add_1_root_add_519_2_n104 ), .B(_add_1_root_add_519_2_n101 ), .ZN(N2528) );
XNOR2_X2 _add_1_root_add_519_2_U182  ( .A(_add_1_root_add_519_2_n103 ), .B(_add_1_root_add_519_2_n80 ), .ZN(N2483) );
INV_X4 _add_1_root_add_519_2_U181  ( .A(aad_byte_cnt[49]), .ZN(_add_1_root_add_519_2_n101 ) );
INV_X4 _add_1_root_add_519_2_U180  ( .A(aad_byte_cnt[50]), .ZN(_add_1_root_add_519_2_n102 ) );
XNOR2_X2 _add_1_root_add_519_2_U179  ( .A(_add_1_root_add_519_2_n37 ), .B(_add_1_root_add_519_2_n102 ), .ZN(N2529) );
INV_X4 _add_1_root_add_519_2_U178  ( .A(_add_1_root_add_519_2_n99 ), .ZN(_add_1_root_add_519_2_n100 ) );
XNOR2_X2 _add_1_root_add_519_2_U177  ( .A(_add_1_root_add_519_2_n12 ), .B(aad_byte_cnt[51]), .ZN(N2530) );
NAND2_X2 _add_1_root_add_519_2_U176  ( .A1(_add_1_root_add_519_2_n99 ), .A2(aad_byte_cnt[51]), .ZN(_add_1_root_add_519_2_n98 ) );
XNOR2_X2 _add_1_root_add_519_2_U175  ( .A(_add_1_root_add_519_2_n11 ), .B(aad_byte_cnt[52]), .ZN(N2531) );
INV_X4 _add_1_root_add_519_2_U174  ( .A(_add_1_root_add_519_2_n98 ), .ZN(_add_1_root_add_519_2_n97 ) );
NAND2_X2 _add_1_root_add_519_2_U173  ( .A1(_add_1_root_add_519_2_n97 ), .A2(aad_byte_cnt[52]), .ZN(_add_1_root_add_519_2_n96 ) );
XNOR2_X2 _add_1_root_add_519_2_U172  ( .A(_add_1_root_add_519_2_n10 ), .B(aad_byte_cnt[53]), .ZN(N2532) );
INV_X4 _add_1_root_add_519_2_U171  ( .A(_add_1_root_add_519_2_n96 ), .ZN(_add_1_root_add_519_2_n77 ) );
NAND2_X2 _add_1_root_add_519_2_U170  ( .A1(_add_1_root_add_519_2_n77 ), .A2(_add_1_root_add_519_2_n78 ), .ZN(_add_1_root_add_519_2_n90 ) );
NAND2_X2 _add_1_root_add_519_2_U169  ( .A1(aad_byte_cnt[48]), .A2(aad_byte_cnt[53]), .ZN(_add_1_root_add_519_2_n95 ) );
NAND2_X2 _add_1_root_add_519_2_U168  ( .A1(_add_1_root_add_519_2_n91 ), .A2(_add_1_root_add_519_2_n92 ), .ZN(_add_1_root_add_519_2_n76 ) );
INV_X4 _add_1_root_add_519_2_U167  ( .A(aad_byte_cnt[54]), .ZN(_add_1_root_add_519_2_n89 ) );
XNOR2_X2 _add_1_root_add_519_2_U166  ( .A(_add_1_root_add_519_2_n1 ), .B(aad_byte_cnt[54]), .ZN(N2533) );
INV_X4 _add_1_root_add_519_2_U165  ( .A(aad_byte_cnt[55]), .ZN(_add_1_root_add_519_2_n88 ) );
XNOR2_X2 _add_1_root_add_519_2_U164  ( .A(_add_1_root_add_519_2_n35 ), .B(aad_byte_cnt[55]), .ZN(N2534) );
INV_X4 _add_1_root_add_519_2_U163  ( .A(_add_1_root_add_519_2_n86 ), .ZN(_add_1_root_add_519_2_n87 ) );
XNOR2_X2 _add_1_root_add_519_2_U162  ( .A(_add_1_root_add_519_2_n16 ), .B(aad_byte_cnt[56]), .ZN(N2535) );
NAND2_X2 _add_1_root_add_519_2_U161  ( .A1(_add_1_root_add_519_2_n86 ), .A2(aad_byte_cnt[56]), .ZN(_add_1_root_add_519_2_n85 ) );
XNOR2_X2 _add_1_root_add_519_2_U160  ( .A(_add_1_root_add_519_2_n15 ), .B(aad_byte_cnt[57]), .ZN(N2536) );
INV_X4 _add_1_root_add_519_2_U159  ( .A(_add_1_root_add_519_2_n85 ), .ZN(_add_1_root_add_519_2_n84 ) );
NAND2_X2 _add_1_root_add_519_2_U158  ( .A1(_add_1_root_add_519_2_n84 ), .A2(aad_byte_cnt[57]), .ZN(_add_1_root_add_519_2_n83 ) );
XNOR2_X2 _add_1_root_add_519_2_U157  ( .A(_add_1_root_add_519_2_n14 ), .B(aad_byte_cnt[58]), .ZN(N2537) );
INV_X4 _add_1_root_add_519_2_U156  ( .A(_add_1_root_add_519_2_n83 ), .ZN(_add_1_root_add_519_2_n82 ) );
NAND2_X2 _add_1_root_add_519_2_U155  ( .A1(_add_1_root_add_519_2_n82 ), .A2(aad_byte_cnt[58]), .ZN(_add_1_root_add_519_2_n74 ) );
XNOR2_X2 _add_1_root_add_519_2_U154  ( .A(_add_1_root_add_519_2_n13 ), .B(aad_byte_cnt[59]), .ZN(N2538) );
XNOR2_X2 _add_1_root_add_519_2_U153  ( .A(_add_1_root_add_519_2_n81 ), .B(_add_1_root_add_519_2_n18 ), .ZN(N2484) );
INV_X4 _add_1_root_add_519_2_U152  ( .A(aad_byte_cnt[60]), .ZN(_add_1_root_add_519_2_n79 ) );
NAND2_X2 _add_1_root_add_519_2_U151  ( .A1(_add_1_root_add_519_2_n77 ), .A2(_add_1_root_add_519_2_n78 ), .ZN(_add_1_root_add_519_2_n75 ) );
INV_X4 _add_1_root_add_519_2_U150  ( .A(_add_1_root_add_519_2_n74 ), .ZN(_add_1_root_add_519_2_n73 ) );
NAND2_X2 _add_1_root_add_519_2_U149  ( .A1(_add_1_root_add_519_2_n73 ), .A2(aad_byte_cnt[59]), .ZN(_add_1_root_add_519_2_n70 ) );
XNOR2_X2 _add_1_root_add_519_2_U148  ( .A(_add_1_root_add_519_2_n79 ), .B(_add_1_root_add_519_2_n19 ), .ZN(N2539) );
INV_X4 _add_1_root_add_519_2_U147  ( .A(aad_byte_cnt[61]), .ZN(_add_1_root_add_519_2_n72 ) );
XNOR2_X2 _add_1_root_add_519_2_U146  ( .A(_add_1_root_add_519_2_n31 ), .B(_add_1_root_add_519_2_n72 ), .ZN(N2540) );
INV_X4 _add_1_root_add_519_2_U145  ( .A(aad_byte_cnt[62]), .ZN(_add_1_root_add_519_2_n71 ) );
XNOR2_X2 _add_1_root_add_519_2_U144  ( .A(_add_1_root_add_519_2_n29 ), .B(_add_1_root_add_519_2_n71 ), .ZN(N2541) );
NAND2_X2 _add_1_root_add_519_2_U143  ( .A1(_add_1_root_add_519_2_n69 ), .A2(aad_byte_cnt[62]), .ZN(_add_1_root_add_519_2_n68 ) );
NAND2_X2 _add_1_root_add_519_2_U142  ( .A1(_add_1_root_add_519_2_n18 ), .A2(aad_byte_cnt[5]), .ZN(_add_1_root_add_519_2_n66 ) );
XNOR2_X2 _add_1_root_add_519_2_U141  ( .A(_add_1_root_add_519_2_n66 ), .B(aad_byte_cnt[6]), .ZN(N2485) );
XNOR2_X2 _add_1_root_add_519_2_U140  ( .A(_add_1_root_add_519_2_n33 ), .B(aad_byte_cnt[7]), .ZN(N2486) );
XNOR2_X2 _add_1_root_add_519_2_U139  ( .A(_add_1_root_add_519_2_n63 ), .B(_add_1_root_add_519_2_n64 ), .ZN(N2487) );
XNOR2_X2 _add_1_root_add_519_2_U138  ( .A(_add_1_root_add_519_2_n58 ), .B(aad_byte_cnt[9]), .ZN(N2488) );
INV_X4 _add_1_root_add_519_2_U137  ( .A(aad_byte_cnt[38]), .ZN(_add_1_root_add_519_2_n134 ) );
INV_X4 _add_1_root_add_519_2_U136  ( .A(aad_byte_cnt[37]), .ZN(_add_1_root_add_519_2_n136 ) );
INV_X4 _add_1_root_add_519_2_U135  ( .A(aad_byte_cnt[36]), .ZN(_add_1_root_add_519_2_n135 ) );
INV_X4 _add_1_root_add_519_2_U134  ( .A(aad_byte_cnt[34]), .ZN(_add_1_root_add_519_2_n150 ) );
INV_X4 _add_1_root_add_519_2_U133  ( .A(aad_byte_cnt[33]), .ZN(_add_1_root_add_519_2_n151 ) );
INV_X4 _add_1_root_add_519_2_U132  ( .A(aad_byte_cnt[32]), .ZN(_add_1_root_add_519_2_n156 ) );
INV_X4 _add_1_root_add_519_2_U131  ( .A(aad_byte_cnt[26]), .ZN(_add_1_root_add_519_2_n169 ) );
INV_X4 _add_1_root_add_519_2_U130  ( .A(aad_byte_cnt[25]), .ZN(_add_1_root_add_519_2_n171 ) );
INV_X4 _add_1_root_add_519_2_U129  ( .A(aad_byte_cnt[24]), .ZN(_add_1_root_add_519_2_n170 ) );
INV_X4 _add_1_root_add_519_2_U128  ( .A(aad_byte_cnt[23]), .ZN(_add_1_root_add_519_2_n175 ) );
INV_X4 _add_1_root_add_519_2_U127  ( .A(aad_byte_cnt[22]), .ZN(_add_1_root_add_519_2_n174 ) );
INV_X4 _add_1_root_add_519_2_U126  ( .A(aad_byte_cnt[21]), .ZN(_add_1_root_add_519_2_n176 ) );
INV_X4 _add_1_root_add_519_2_U125  ( .A(aad_byte_cnt[20]), .ZN(_add_1_root_add_519_2_n179 ) );
INV_X4 _add_1_root_add_519_2_U124  ( .A(aad_byte_cnt[18]), .ZN(_add_1_root_add_519_2_n181 ) );
INV_X4 _add_1_root_add_519_2_U123  ( .A(aad_byte_cnt[17]), .ZN(_add_1_root_add_519_2_n189 ) );
INV_X4 _add_1_root_add_519_2_U122  ( .A(aad_byte_cnt[16]), .ZN(_add_1_root_add_519_2_n182 ) );
INV_X4 _add_1_root_add_519_2_U121  ( .A(aad_byte_cnt[10]), .ZN(_add_1_root_add_519_2_n206 ) );
INV_X4 _add_1_root_add_519_2_U120  ( .A(aad_byte_cnt[9]), .ZN(_add_1_root_add_519_2_n62 ) );
INV_X4 _add_1_root_add_519_2_U119  ( .A(aad_byte_cnt[8]), .ZN(_add_1_root_add_519_2_n64 ) );
INV_X4 _add_1_root_add_519_2_U118  ( .A(aad_byte_cnt[6]), .ZN(_add_1_root_add_519_2_n65 ) );
INV_X4 _add_1_root_add_519_2_U117  ( .A(aad_byte_cnt[4]), .ZN(_add_1_root_add_519_2_n103 ) );
INV_X4 _add_1_root_add_519_2_U116  ( .A(aad_byte_cnt[5]), .ZN(_add_1_root_add_519_2_n81 ) );
INV_X4 _add_1_root_add_519_2_U115  ( .A(_add_1_root_add_519_2_n186 ), .ZN(_add_1_root_add_519_2_n210 ) );
INV_X4 _add_1_root_add_519_2_U114  ( .A(_add_1_root_add_519_2_n114 ), .ZN(_add_1_root_add_519_2_n157 ) );
INV_X4 _add_1_root_add_519_2_U113  ( .A(_add_1_root_add_519_2_n127 ), .ZN(_add_1_root_add_519_2_n128 ) );
INV_X4 _add_1_root_add_519_2_U112  ( .A(_add_1_root_add_519_2_n208 ), .ZN(_add_1_root_add_519_2_n63 ) );
OR2_X2 _add_1_root_add_519_2_U111  ( .A1(aad_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(_add_1_root_add_519_2_n60 ) );
NOR2_X2 _add_1_root_add_519_2_U110  ( .A1(_add_1_root_add_519_2_n48 ), .A2(_add_1_root_add_519_2_n68 ), .ZN(_add_1_root_add_519_2_n67 ) );
XOR2_X2 _add_1_root_add_519_2_U109  ( .A(_add_1_root_add_519_2_n67 ), .B(aad_byte_cnt[63]), .Z(N2542) );
AND2_X2 _add_1_root_add_519_2_U108  ( .A1(aad_byte_cnt[0]), .A2(n17750),.ZN(_add_1_root_add_519_2_n219 ) );
NOR2_X2 _add_1_root_add_519_2_U107  ( .A1(_add_1_root_add_519_2_n217 ), .A2(_add_1_root_add_519_2_n218 ), .ZN(_add_1_root_add_519_2_n216 ) );
NAND3_X2 _add_1_root_add_519_2_U106  ( .A1(dii_data_size[1]), .A2(_add_1_root_add_519_2_n60 ), .A3(aad_byte_cnt[1]), .ZN(_add_1_root_add_519_2_n215 ) );
NAND3_X2 _add_1_root_add_519_2_U105  ( .A1(_add_1_root_add_519_2_n214 ),.A2(_add_1_root_add_519_2_n215 ), .A3(_add_1_root_add_519_2_n216 ),.ZN(_add_1_root_add_519_2_n193 ) );
NOR2_X2 _add_1_root_add_519_2_U104  ( .A1(aad_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(_add_1_root_add_519_2_n222 ) );
NOR2_X2 _add_1_root_add_519_2_U103  ( .A1(aad_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(_add_1_root_add_519_2_n221 ) );
NOR2_X2 _add_1_root_add_519_2_U102  ( .A1(_add_1_root_add_519_2_n221 ), .A2(_add_1_root_add_519_2_n222 ), .ZN(_add_1_root_add_519_2_n220 ) );
NOR2_X2 _add_1_root_add_519_2_U101  ( .A1(aad_byte_cnt[0]), .A2(n17750),.ZN(_add_1_root_add_519_2_n186 ) );
NOR2_X2 _add_1_root_add_519_2_U100  ( .A1(aad_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(_add_1_root_add_519_2_n165 ) );
INV_X4 _add_1_root_add_519_2_U99  ( .A(n18074), .ZN(_add_1_root_add_519_2_n61 ) );
AND2_X2 _add_1_root_add_519_2_U98  ( .A1(_add_1_root_add_519_2_n186 ), .A2(_add_1_root_add_519_2_n185 ), .ZN(_add_1_root_add_519_2_n166 ) );
NOR2_X2 _add_1_root_add_519_2_U97  ( .A1(_add_1_root_add_519_2_n154 ), .A2(_add_1_root_add_519_2_n150 ), .ZN(_add_1_root_add_519_2_n149 ) );
OR2_X2 _add_1_root_add_519_2_U96  ( .A1(_add_1_root_add_519_2_n58 ), .A2(_add_1_root_add_519_2_n62 ), .ZN(_add_1_root_add_519_2_n59 ) );
NOR2_X2 _add_1_root_add_519_2_U95  ( .A1(_add_1_root_add_519_2_n134 ), .A2(_add_1_root_add_519_2_n144 ), .ZN(_add_1_root_add_519_2_n133 ) );
NAND3_X2 _add_1_root_add_519_2_U94  ( .A1(aad_byte_cnt[37]), .A2(aad_byte_cnt[36]), .A3(_add_1_root_add_519_2_n133 ), .ZN(_add_1_root_add_519_2_n111 ) );
OR2_X2 _add_1_root_add_519_2_U93  ( .A1(_add_1_root_add_519_2_n208 ), .A2(_add_1_root_add_519_2_n64 ), .ZN(_add_1_root_add_519_2_n58 ) );
NOR2_X2 _add_1_root_add_519_2_U92  ( .A1(_add_1_root_add_519_2_n167 ), .A2(_add_1_root_add_519_2_n159 ), .ZN(_add_1_root_add_519_2_n158 ) );
NAND3_X2 _add_1_root_add_519_2_U91  ( .A1(aad_byte_cnt[30]), .A2(aad_byte_cnt[31]), .A3(_add_1_root_add_519_2_n158 ), .ZN(_add_1_root_add_519_2_n93 ) );
NOR2_X2 _add_1_root_add_519_2_U90  ( .A1(_add_1_root_add_519_2_n184 ), .A2(_add_1_root_add_519_2_n165 ), .ZN(_add_1_root_add_519_2_n183 ) );
NOR2_X2 _add_1_root_add_519_2_U89  ( .A1(_add_1_root_add_519_2_n151 ), .A2(_add_1_root_add_519_2_n156 ), .ZN(_add_1_root_add_519_2_n155 ) );
AND2_X2 _add_1_root_add_519_2_U88  ( .A1(aad_byte_cnt[61]), .A2(aad_byte_cnt[60]), .ZN(_add_1_root_add_519_2_n69 ) );
NOR2_X2 _add_1_root_add_519_2_U87  ( .A1(_add_1_root_add_519_2_n169 ), .A2(_add_1_root_add_519_2_n172 ), .ZN(_add_1_root_add_519_2_n168 ) );
NAND3_X2 _add_1_root_add_519_2_U86  ( .A1(aad_byte_cnt[25]), .A2(aad_byte_cnt[24]), .A3(_add_1_root_add_519_2_n168 ), .ZN(_add_1_root_add_519_2_n94 ) );
NOR2_X2 _add_1_root_add_519_2_U85  ( .A1(_add_1_root_add_519_2_n102 ), .A2(_add_1_root_add_519_2_n101 ), .ZN(_add_1_root_add_519_2_n99 ) );
NOR2_X2 _add_1_root_add_519_2_U84  ( .A1(_add_1_root_add_519_2_n88 ), .A2(_add_1_root_add_519_2_n89 ), .ZN(_add_1_root_add_519_2_n86 ) );
NOR2_X2 _add_1_root_add_519_2_U83  ( .A1(_add_1_root_add_519_2_n187 ), .A2(_add_1_root_add_519_2_n181 ), .ZN(_add_1_root_add_519_2_n180 ) );
NAND3_X2 _add_1_root_add_519_2_U82  ( .A1(aad_byte_cnt[16]), .A2(aad_byte_cnt[17]), .A3(_add_1_root_add_519_2_n180 ), .ZN(_add_1_root_add_519_2_n153 ) );
NOR2_X2 _add_1_root_add_519_2_U81  ( .A1(_add_1_root_add_519_2_n174 ), .A2(_add_1_root_add_519_2_n175 ), .ZN(_add_1_root_add_519_2_n173 ) );
NAND3_X2 _add_1_root_add_519_2_U80  ( .A1(aad_byte_cnt[21]), .A2(aad_byte_cnt[20]), .A3(_add_1_root_add_519_2_n173 ), .ZN(_add_1_root_add_519_2_n108 ) );
OR2_X2 _add_1_root_add_519_2_U79  ( .A1(_add_1_root_add_519_2_n165 ), .A2(_add_1_root_add_519_2_n166 ), .ZN(_add_1_root_add_519_2_n57 ) );
NOR3_X2 _add_1_root_add_519_2_U78  ( .A1(_add_1_root_add_519_2_n93 ), .A2(_add_1_root_add_519_2_n94 ), .A3(_add_1_root_add_519_2_n95 ), .ZN(_add_1_root_add_519_2_n91 ) );
AND2_X4 _add_1_root_add_519_2_U77  ( .A1(_add_1_root_add_519_2_n92 ), .A2(aad_byte_cnt[48]), .ZN(_add_1_root_add_519_2_n56 ) );
NAND2_X2 _add_1_root_add_519_2_U76  ( .A1(_add_1_root_add_519_2_n106 ), .A2(_add_1_root_add_519_2_n56 ), .ZN(_add_1_root_add_519_2_n55 ) );
NOR2_X2 _add_1_root_add_519_2_U75  ( .A1(_add_1_root_add_519_2_n212 ), .A2(_add_1_root_add_519_2_n165 ), .ZN(_add_1_root_add_519_2_n211 ) );
NAND3_X2 _add_1_root_add_519_2_U74  ( .A1(_add_1_root_add_519_2_n210 ), .A2(_add_1_root_add_519_2_n60 ), .A3(_add_1_root_add_519_2_n211 ), .ZN(_add_1_root_add_519_2_n200 ) );
OR3_X2 _add_1_root_add_519_2_U73  ( .A1(_add_1_root_add_519_2_n2 ), .A2(_add_1_root_add_519_2_n135 ), .A3(_add_1_root_add_519_2_n136 ), .ZN(_add_1_root_add_519_2_n54 ) );
OR3_X2 _add_1_root_add_519_2_U72  ( .A1(_add_1_root_add_519_2_n47 ), .A2(_add_1_root_add_519_2_n167 ), .A3(_add_1_root_add_519_2_n159 ), .ZN(_add_1_root_add_519_2_n53 ) );
NOR2_X2 _add_1_root_add_519_2_U71  ( .A1(_add_1_root_add_519_2_n65 ), .A2(_add_1_root_add_519_2_n224 ), .ZN(_add_1_root_add_519_2_n223 ) );
NAND3_X2 _add_1_root_add_519_2_U70  ( .A1(aad_byte_cnt[5]), .A2(aad_byte_cnt[4]), .A3(_add_1_root_add_519_2_n223 ), .ZN(_add_1_root_add_519_2_n198 ) );
OR2_X2 _add_1_root_add_519_2_U69  ( .A1(_add_1_root_add_519_2_n176 ), .A2(_add_1_root_add_519_2_n177 ), .ZN(_add_1_root_add_519_2_n52 ) );
OR2_X2 _add_1_root_add_519_2_U68  ( .A1(_add_1_root_add_519_2_n171 ), .A2(_add_1_root_add_519_2_n50 ), .ZN(_add_1_root_add_519_2_n51 ) );
OR2_X2 _add_1_root_add_519_2_U67  ( .A1(_add_1_root_add_519_2_n170 ), .A2(_add_1_root_add_519_2_n43 ), .ZN(_add_1_root_add_519_2_n50 ) );
AND2_X2 _add_1_root_add_519_2_U66  ( .A1(aad_byte_cnt[13]), .A2(aad_byte_cnt[12]), .ZN(_add_1_root_add_519_2_n199 ) );
AND2_X4 _add_1_root_add_519_2_U65  ( .A1(_add_1_root_add_519_2_n118 ), .A2(aad_byte_cnt[45]), .ZN(_add_1_root_add_519_2_n49 ) );
AND2_X2 _add_1_root_add_519_2_U64  ( .A1(_add_1_root_add_519_2_n114 ), .A2(_add_1_root_add_519_2_n49 ), .ZN(_add_1_root_add_519_2_n116 ) );
NOR2_X2 _add_1_root_add_519_2_U63  ( .A1(_add_1_root_add_519_2_n206 ), .A2(_add_1_root_add_519_2_n207 ), .ZN(_add_1_root_add_519_2_n205 ) );
NAND3_X2 _add_1_root_add_519_2_U62  ( .A1(aad_byte_cnt[9]), .A2(aad_byte_cnt[8]), .A3(_add_1_root_add_519_2_n205 ), .ZN(_add_1_root_add_519_2_n192 ) );
NAND3_X2 _add_1_root_add_519_2_U61  ( .A1(_add_1_root_add_519_2_n140 ), .A2(_add_1_root_add_519_2_n193 ), .A3(_add_1_root_add_519_2_n194 ), .ZN(_add_1_root_add_519_2_n190 ) );
NOR2_X2 _add_1_root_add_519_2_U60  ( .A1(_add_1_root_add_519_2_n111 ), .A2(_add_1_root_add_519_2_n112 ), .ZN(_add_1_root_add_519_2_n110 ) );
NOR3_X2 _add_1_root_add_519_2_U59  ( .A1(_add_1_root_add_519_2_n113 ), .A2(_add_1_root_add_519_2_n120 ), .A3(_add_1_root_add_519_2_n123 ), .ZN(_add_1_root_add_519_2_n109 ) );
NAND3_X2 _add_1_root_add_519_2_U58  ( .A1(_add_1_root_add_519_2_n109 ), .A2(_add_1_root_add_519_2_n8 ), .A3(_add_1_root_add_519_2_n110 ), .ZN(_add_1_root_add_519_2_n105 ) );
AND2_X2 _add_1_root_add_519_2_U57  ( .A1(_add_1_root_add_519_2_n195 ), .A2(_add_1_root_add_519_2_n42 ), .ZN(_add_1_root_add_519_2_n152 ) );
OR2_X2 _add_1_root_add_519_2_U56  ( .A1(_add_1_root_add_519_2_n1 ), .A2(_add_1_root_add_519_2_n70 ), .ZN(_add_1_root_add_519_2_n48 ) );
NOR2_X2 _add_1_root_add_519_2_U55  ( .A1(_add_1_root_add_519_2_n198 ), .A2(_add_1_root_add_519_2_n191 ), .ZN(_add_1_root_add_519_2_n197 ) );
NOR2_X2 _add_1_root_add_519_2_U54  ( .A1(_add_1_root_add_519_2_n192 ), .A2(_add_1_root_add_519_2_n200 ), .ZN(_add_1_root_add_519_2_n196 ) );
OR2_X2 _add_1_root_add_519_2_U53  ( .A1(_add_1_root_add_519_2_n43 ), .A2(_add_1_root_add_519_2_n94 ), .ZN(_add_1_root_add_519_2_n47 ) );
OR2_X2 _add_1_root_add_519_2_U52  ( .A1(_add_1_root_add_519_2_n152 ), .A2(_add_1_root_add_519_2_n153 ), .ZN(_add_1_root_add_519_2_n46 ) );
OR2_X2 _add_1_root_add_519_2_U51  ( .A1(_add_1_root_add_519_2_n152 ), .A2(_add_1_root_add_519_2_n153 ), .ZN(_add_1_root_add_519_2_n45 ) );
AND2_X4 _add_1_root_add_519_2_U50  ( .A1(_add_1_root_add_519_2_n129 ), .A2(aad_byte_cnt[41]), .ZN(_add_1_root_add_519_2_n44 ) );
AND2_X2 _add_1_root_add_519_2_U49  ( .A1(_add_1_root_add_519_2_n114 ), .A2(_add_1_root_add_519_2_n44 ), .ZN(_add_1_root_add_519_2_n127 ) );
OR3_X2 _add_1_root_add_519_2_U48  ( .A1(_add_1_root_add_519_2_n152 ), .A2(_add_1_root_add_519_2_n153 ), .A3(_add_1_root_add_519_2_n108 ), .ZN(_add_1_root_add_519_2_n43 ) );
NOR3_X2 _add_1_root_add_519_2_U47  ( .A1(_add_1_root_add_519_2_n46 ), .A2(_add_1_root_add_519_2_n107 ), .A3(_add_1_root_add_519_2_n108 ), .ZN(_add_1_root_add_519_2_n106 ) );
NOR3_X2 _add_1_root_add_519_2_U46  ( .A1(_add_1_root_add_519_2_n107 ), .A2(_add_1_root_add_519_2_n45 ), .A3(_add_1_root_add_519_2_n108 ), .ZN(_add_1_root_add_519_2_n114 ) );
XNOR2_X1 _add_1_root_add_519_2_U45  ( .A(_add_1_root_add_519_2_n163 ), .B(_add_1_root_add_519_2_n143 ), .ZN(N2481) );
OR3_X4 _add_1_root_add_519_2_U44  ( .A1(_add_1_root_add_519_2_n190 ), .A2(_add_1_root_add_519_2_n191 ), .A3(_add_1_root_add_519_2_n192 ), .ZN(_add_1_root_add_519_2_n42 ) );
OR3_X4 _add_1_root_add_519_2_U43  ( .A1(_add_1_root_add_519_2_n46 ), .A2(_add_1_root_add_519_2_n75 ), .A3(_add_1_root_add_519_2_n76 ), .ZN(_add_1_root_add_519_2_n41 ) );
OR2_X4 _add_1_root_add_519_2_U42  ( .A1(_add_1_root_add_519_2_n181 ), .A2(_add_1_root_add_519_2_n188 ), .ZN(_add_1_root_add_519_2_n40 ) );
OR2_X4 _add_1_root_add_519_2_U41  ( .A1(_add_1_root_add_519_2_n135 ), .A2(_add_1_root_add_519_2_n2 ), .ZN(_add_1_root_add_519_2_n39 ) );
OR2_X4 _add_1_root_add_519_2_U40  ( .A1(_add_1_root_add_519_2_n134 ), .A2(_add_1_root_add_519_2_n54 ), .ZN(_add_1_root_add_519_2_n38 ) );
NOR2_X2 _add_1_root_add_519_2_U39  ( .A1(_add_1_root_add_519_2_n101 ), .A2(_add_1_root_add_519_2_n55 ), .ZN(_add_1_root_add_519_2_n37 ) );
OR2_X4 _add_1_root_add_519_2_U38  ( .A1(_add_1_root_add_519_2_n157 ), .A2(_add_1_root_add_519_2_n122 ), .ZN(_add_1_root_add_519_2_n36 ) );
OR2_X4 _add_1_root_add_519_2_U37  ( .A1(_add_1_root_add_519_2_n89 ), .A2(_add_1_root_add_519_2_n1 ), .ZN(_add_1_root_add_519_2_n35 ) );
AND2_X4 _add_1_root_add_519_2_U36  ( .A1(_add_1_root_add_519_2_n114 ), .A2(aad_byte_cnt[32]), .ZN(_add_1_root_add_519_2_n34 ) );
OR2_X4 _add_1_root_add_519_2_U35  ( .A1(_add_1_root_add_519_2_n65 ), .A2(_add_1_root_add_519_2_n66 ), .ZN(_add_1_root_add_519_2_n33 ) );
OR2_X4 _add_1_root_add_519_2_U34  ( .A1(_add_1_root_add_519_2_n206 ), .A2(_add_1_root_add_519_2_n59 ), .ZN(_add_1_root_add_519_2_n32 ) );
AND2_X4 _add_1_root_add_519_2_U33  ( .A1(aad_byte_cnt[60]), .A2(_add_1_root_add_519_2_n19 ), .ZN(_add_1_root_add_519_2_n31 ) );
AND2_X4 _add_1_root_add_519_2_U32  ( .A1(aad_byte_cnt[14]), .A2(_add_1_root_add_519_2_n9 ), .ZN(_add_1_root_add_519_2_n30 ) );
AND2_X4 _add_1_root_add_519_2_U31  ( .A1(_add_1_root_add_519_2_n69 ), .A2(_add_1_root_add_519_2_n19 ), .ZN(_add_1_root_add_519_2_n29 ) );
OR2_X4 _add_1_root_add_519_2_U30  ( .A1(_add_1_root_add_519_2_n169 ), .A2(_add_1_root_add_519_2_n51 ), .ZN(_add_1_root_add_519_2_n28 ) );
OR2_X4 _add_1_root_add_519_2_U29  ( .A1(_add_1_root_add_519_2_n174 ), .A2(_add_1_root_add_519_2_n52 ), .ZN(_add_1_root_add_519_2_n27 ) );
AND2_X4 _add_1_root_add_519_2_U28  ( .A1(_add_1_root_add_519_2_n127 ), .A2(aad_byte_cnt[42]), .ZN(_add_1_root_add_519_2_n26 ) );
AND2_X4 _add_1_root_add_519_2_U27  ( .A1(_add_1_root_add_519_2_n116 ), .A2(aad_byte_cnt[46]), .ZN(_add_1_root_add_519_2_n25 ) );
OR2_X4 _add_1_root_add_519_2_U26  ( .A1(_add_1_root_add_519_2_n157 ), .A2(_add_1_root_add_519_2_n131 ), .ZN(_add_1_root_add_519_2_n24 ) );
OR2_X4 _add_1_root_add_519_2_U25  ( .A1(_add_1_root_add_519_2_n157 ), .A2(_add_1_root_add_519_2_n130 ), .ZN(_add_1_root_add_519_2_n23 ) );
OR2_X4 _add_1_root_add_519_2_U24  ( .A1(_add_1_root_add_519_2_n157 ), .A2(_add_1_root_add_519_2_n119 ), .ZN(_add_1_root_add_519_2_n22 ) );
OR2_X4 _add_1_root_add_519_2_U23  ( .A1(_add_1_root_add_519_2_n159 ), .A2(_add_1_root_add_519_2_n47 ), .ZN(_add_1_root_add_519_2_n21 ) );
OR2_X4 _add_1_root_add_519_2_U22  ( .A1(_add_1_root_add_519_2_n157 ), .A2(_add_1_root_add_519_2_n105 ), .ZN(_add_1_root_add_519_2_n20 ) );
NOR2_X2 _add_1_root_add_519_2_U21  ( .A1(_add_1_root_add_519_2_n41 ), .A2(_add_1_root_add_519_2_n70 ), .ZN(_add_1_root_add_519_2_n19 ) );
AND2_X4 _add_1_root_add_519_2_U20  ( .A1(aad_byte_cnt[4]), .A2(_add_1_root_add_519_2_n80 ), .ZN(_add_1_root_add_519_2_n18 ) );
NOR2_X2 _add_1_root_add_519_2_U19  ( .A1(_add_1_root_add_519_2_n162 ), .A2(_add_1_root_add_519_2_n53 ), .ZN(_add_1_root_add_519_2_n17 ) );
OR2_X4 _add_1_root_add_519_2_U18  ( .A1(_add_1_root_add_519_2_n1 ), .A2(_add_1_root_add_519_2_n87 ), .ZN(_add_1_root_add_519_2_n16 ) );
OR2_X4 _add_1_root_add_519_2_U17  ( .A1(_add_1_root_add_519_2_n1 ), .A2(_add_1_root_add_519_2_n85 ), .ZN(_add_1_root_add_519_2_n15 ) );
OR2_X4 _add_1_root_add_519_2_U16  ( .A1(_add_1_root_add_519_2_n1 ), .A2(_add_1_root_add_519_2_n83 ), .ZN(_add_1_root_add_519_2_n14 ) );
OR2_X4 _add_1_root_add_519_2_U15  ( .A1(_add_1_root_add_519_2_n1 ), .A2(_add_1_root_add_519_2_n74 ), .ZN(_add_1_root_add_519_2_n13 ) );
OR2_X4 _add_1_root_add_519_2_U14  ( .A1(_add_1_root_add_519_2_n55 ), .A2(_add_1_root_add_519_2_n100 ), .ZN(_add_1_root_add_519_2_n12 ) );
OR2_X4 _add_1_root_add_519_2_U13  ( .A1(_add_1_root_add_519_2_n55 ), .A2(_add_1_root_add_519_2_n98 ), .ZN(_add_1_root_add_519_2_n11 ) );
OR2_X4 _add_1_root_add_519_2_U12  ( .A1(_add_1_root_add_519_2_n55 ), .A2(_add_1_root_add_519_2_n96 ), .ZN(_add_1_root_add_519_2_n10 ) );
AND2_X4 _add_1_root_add_519_2_U11  ( .A1(_add_1_root_add_519_2_n6 ), .A2(aad_byte_cnt[13]), .ZN(_add_1_root_add_519_2_n9 ) );
AND3_X4 _add_1_root_add_519_2_U10  ( .A1(aad_byte_cnt[32]), .A2(aad_byte_cnt[33]), .A3(_add_1_root_add_519_2_n149 ), .ZN(_add_1_root_add_519_2_n8 ) );
AND2_X4 _add_1_root_add_519_2_U9  ( .A1(_add_1_root_add_519_2_n3 ), .A2(aad_byte_cnt[34]), .ZN(_add_1_root_add_519_2_n7 ) );
AND2_X4 _add_1_root_add_519_2_U8  ( .A1(_add_1_root_add_519_2_n5 ), .A2(aad_byte_cnt[12]), .ZN(_add_1_root_add_519_2_n6 ) );
NOR2_X2 _add_1_root_add_519_2_U7  ( .A1(_add_1_root_add_519_2_n208 ), .A2(_add_1_root_add_519_2_n192 ), .ZN(_add_1_root_add_519_2_n5 ) );
NOR2_X2 _add_1_root_add_519_2_U6  ( .A1(_add_1_root_add_519_2_n152 ), .A2(_add_1_root_add_519_2_n182 ), .ZN(_add_1_root_add_519_2_n4 ) );
AND2_X4 _add_1_root_add_519_2_U5  ( .A1(_add_1_root_add_519_2_n114 ), .A2(_add_1_root_add_519_2_n155 ), .ZN(_add_1_root_add_519_2_n3 ) );
OR3_X4 _add_1_root_add_519_2_U4  ( .A1(_add_1_root_add_519_2_n46 ), .A2(_add_1_root_add_519_2_n145 ), .A3(_add_1_root_add_519_2_n146 ), .ZN(_add_1_root_add_519_2_n2 ) );
OR3_X4 _add_1_root_add_519_2_U3  ( .A1(_add_1_root_add_519_2_n46 ), .A2(_add_1_root_add_519_2_n90 ), .A3(_add_1_root_add_519_2_n76 ), .ZN(_add_1_root_add_519_2_n1 ) );
NAND3_X2 _add_1_root_add_519_2_U2  ( .A1(aad_byte_cnt[14]), .A2(aad_byte_cnt[15]), .A3(_add_1_root_add_519_2_n199 ), .ZN(_add_1_root_add_519_2_n191 ) );
INV_X4 _add_1_root_add_513_2_U289  ( .A(enc_byte_cnt[7]), .ZN(_add_1_root_add_513_2_n224 ) );
INV_X4 _add_1_root_add_513_2_U288  ( .A(_add_1_root_add_513_2_n198 ), .ZN(_add_1_root_add_513_2_n194 ) );
NAND2_X2 _add_1_root_add_513_2_U287  ( .A1(_add_1_root_add_513_2_n219 ),.A2(_add_1_root_add_513_2_n220 ), .ZN(_add_1_root_add_513_2_n214 ) );
NAND2_X2 _add_1_root_add_513_2_U286  ( .A1(dii_data_size[2]), .A2(enc_byte_cnt[2]), .ZN(_add_1_root_add_513_2_n142 ) );
INV_X4 _add_1_root_add_513_2_U285  ( .A(_add_1_root_add_513_2_n142 ), .ZN(_add_1_root_add_513_2_n217 ) );
NAND2_X2 _add_1_root_add_513_2_U284  ( .A1(n18074), .A2(enc_byte_cnt[3]),.ZN(_add_1_root_add_513_2_n139 ) );
INV_X4 _add_1_root_add_513_2_U283  ( .A(_add_1_root_add_513_2_n139 ), .ZN(_add_1_root_add_513_2_n218 ) );
INV_X4 _add_1_root_add_513_2_U282  ( .A(enc_byte_cnt[3]), .ZN(_add_1_root_add_513_2_n213 ) );
NAND2_X2 _add_1_root_add_513_2_U281  ( .A1(_add_1_root_add_513_2_n61 ), .A2(_add_1_root_add_513_2_n213 ), .ZN(_add_1_root_add_513_2_n140 ) );
NAND2_X2 _add_1_root_add_513_2_U280  ( .A1(_add_1_root_add_513_2_n193 ),.A2(_add_1_root_add_513_2_n140 ), .ZN(_add_1_root_add_513_2_n209 ) );
INV_X4 _add_1_root_add_513_2_U279  ( .A(_add_1_root_add_513_2_n140 ), .ZN(_add_1_root_add_513_2_n212 ) );
NAND2_X2 _add_1_root_add_513_2_U278  ( .A1(_add_1_root_add_513_2_n209 ),.A2(_add_1_root_add_513_2_n200 ), .ZN(_add_1_root_add_513_2_n80 ) );
NAND2_X2 _add_1_root_add_513_2_U277  ( .A1(_add_1_root_add_513_2_n194 ),.A2(_add_1_root_add_513_2_n80 ), .ZN(_add_1_root_add_513_2_n208 ) );
XNOR2_X2 _add_1_root_add_513_2_U276  ( .A(_add_1_root_add_513_2_n59 ), .B(enc_byte_cnt[10]), .ZN(N2359) );
INV_X4 _add_1_root_add_513_2_U275  ( .A(enc_byte_cnt[11]), .ZN(_add_1_root_add_513_2_n207 ) );
XNOR2_X2 _add_1_root_add_513_2_U274  ( .A(_add_1_root_add_513_2_n28 ), .B(enc_byte_cnt[11]), .ZN(N2360) );
INV_X4 _add_1_root_add_513_2_U273  ( .A(enc_byte_cnt[12]), .ZN(_add_1_root_add_513_2_n204 ) );
XNOR2_X2 _add_1_root_add_513_2_U272  ( .A(_add_1_root_add_513_2_n3 ), .B(_add_1_root_add_513_2_n204 ), .ZN(N2361) );
INV_X4 _add_1_root_add_513_2_U271  ( .A(enc_byte_cnt[13]), .ZN(_add_1_root_add_513_2_n203 ) );
XNOR2_X2 _add_1_root_add_513_2_U270  ( .A(_add_1_root_add_513_2_n4 ), .B(_add_1_root_add_513_2_n203 ), .ZN(N2362) );
INV_X4 _add_1_root_add_513_2_U269  ( .A(enc_byte_cnt[14]), .ZN(_add_1_root_add_513_2_n202 ) );
XNOR2_X2 _add_1_root_add_513_2_U268  ( .A(_add_1_root_add_513_2_n7 ), .B(_add_1_root_add_513_2_n202 ), .ZN(N2363) );
INV_X4 _add_1_root_add_513_2_U267  ( .A(enc_byte_cnt[15]), .ZN(_add_1_root_add_513_2_n201 ) );
XNOR2_X2 _add_1_root_add_513_2_U266  ( .A(_add_1_root_add_513_2_n26 ), .B(_add_1_root_add_513_2_n201 ), .ZN(N2364) );
NAND2_X2 _add_1_root_add_513_2_U265  ( .A1(_add_1_root_add_513_2_n196 ),.A2(_add_1_root_add_513_2_n197 ), .ZN(_add_1_root_add_513_2_n195 ) );
XNOR2_X2 _add_1_root_add_513_2_U264  ( .A(_add_1_root_add_513_2_n152 ), .B(enc_byte_cnt[16]), .ZN(N2365) );
XNOR2_X2 _add_1_root_add_513_2_U263  ( .A(_add_1_root_add_513_2_n189 ), .B(_add_1_root_add_513_2_n2 ), .ZN(N2366) );
NAND2_X2 _add_1_root_add_513_2_U262  ( .A1(_add_1_root_add_513_2_n2 ), .A2(enc_byte_cnt[17]), .ZN(_add_1_root_add_513_2_n188 ) );
XNOR2_X2 _add_1_root_add_513_2_U261  ( .A(_add_1_root_add_513_2_n188 ), .B(enc_byte_cnt[18]), .ZN(N2367) );
INV_X4 _add_1_root_add_513_2_U260  ( .A(enc_byte_cnt[19]), .ZN(_add_1_root_add_513_2_n187 ) );
XNOR2_X2 _add_1_root_add_513_2_U259  ( .A(_add_1_root_add_513_2_n48 ), .B(enc_byte_cnt[19]), .ZN(N2368) );
NAND2_X2 _add_1_root_add_513_2_U258  ( .A1(dii_data_size[1]), .A2(enc_byte_cnt[1]), .ZN(_add_1_root_add_513_2_n164 ) );
INV_X4 _add_1_root_add_513_2_U257  ( .A(_add_1_root_add_513_2_n164 ), .ZN(_add_1_root_add_513_2_n184 ) );
XNOR2_X2 _add_1_root_add_513_2_U256  ( .A(_add_1_root_add_513_2_n166 ), .B(_add_1_root_add_513_2_n183 ), .ZN(N2350) );
INV_X4 _add_1_root_add_513_2_U255  ( .A(_add_1_root_add_513_2_n41 ), .ZN(_add_1_root_add_513_2_n178 ) );
XNOR2_X2 _add_1_root_add_513_2_U254  ( .A(_add_1_root_add_513_2_n179 ), .B(_add_1_root_add_513_2_n178 ), .ZN(N2369) );
NAND2_X2 _add_1_root_add_513_2_U253  ( .A1(_add_1_root_add_513_2_n178 ),.A2(enc_byte_cnt[20]), .ZN(_add_1_root_add_513_2_n177 ) );
XNOR2_X2 _add_1_root_add_513_2_U252  ( .A(_add_1_root_add_513_2_n177 ), .B(enc_byte_cnt[21]), .ZN(N2370) );
XNOR2_X2 _add_1_root_add_513_2_U251  ( .A(_add_1_root_add_513_2_n51 ), .B(enc_byte_cnt[22]), .ZN(N2371) );
XNOR2_X2 _add_1_root_add_513_2_U250  ( .A(_add_1_root_add_513_2_n23 ), .B(enc_byte_cnt[23]), .ZN(N2372) );
XNOR2_X2 _add_1_root_add_513_2_U249  ( .A(_add_1_root_add_513_2_n38 ), .B(enc_byte_cnt[24]), .ZN(N2373) );
XNOR2_X2 _add_1_root_add_513_2_U248  ( .A(_add_1_root_add_513_2_n49 ), .B(enc_byte_cnt[25]), .ZN(N2374) );
XNOR2_X2 _add_1_root_add_513_2_U247  ( .A(_add_1_root_add_513_2_n50 ), .B(enc_byte_cnt[26]), .ZN(N2375) );
INV_X4 _add_1_root_add_513_2_U246  ( .A(enc_byte_cnt[27]), .ZN(_add_1_root_add_513_2_n172 ) );
XNOR2_X2 _add_1_root_add_513_2_U245  ( .A(_add_1_root_add_513_2_n24 ), .B(enc_byte_cnt[27]), .ZN(N2376) );
INV_X4 _add_1_root_add_513_2_U244  ( .A(enc_byte_cnt[28]), .ZN(_add_1_root_add_513_2_n159 ) );
XNOR2_X2 _add_1_root_add_513_2_U243  ( .A(_add_1_root_add_513_2_n42 ), .B(enc_byte_cnt[28]), .ZN(N2377) );
INV_X4 _add_1_root_add_513_2_U242  ( .A(enc_byte_cnt[29]), .ZN(_add_1_root_add_513_2_n167 ) );
XNOR2_X2 _add_1_root_add_513_2_U241  ( .A(_add_1_root_add_513_2_n52 ), .B(enc_byte_cnt[29]), .ZN(N2378) );
NAND2_X2 _add_1_root_add_513_2_U240  ( .A1(_add_1_root_add_513_2_n60 ), .A2(_add_1_root_add_513_2_n142 ), .ZN(_add_1_root_add_513_2_n163 ) );
NAND2_X2 _add_1_root_add_513_2_U239  ( .A1(_add_1_root_add_513_2_n57 ), .A2(_add_1_root_add_513_2_n164 ), .ZN(_add_1_root_add_513_2_n143 ) );
INV_X4 _add_1_root_add_513_2_U238  ( .A(_add_1_root_add_513_2_n53 ), .ZN(_add_1_root_add_513_2_n161 ) );
INV_X4 _add_1_root_add_513_2_U237  ( .A(enc_byte_cnt[30]), .ZN(_add_1_root_add_513_2_n162 ) );
XNOR2_X2 _add_1_root_add_513_2_U236  ( .A(_add_1_root_add_513_2_n161 ), .B(_add_1_root_add_513_2_n162 ), .ZN(N2379) );
INV_X4 _add_1_root_add_513_2_U235  ( .A(enc_byte_cnt[31]), .ZN(_add_1_root_add_513_2_n160 ) );
XNOR2_X2 _add_1_root_add_513_2_U234  ( .A(_add_1_root_add_513_2_n13 ), .B(_add_1_root_add_513_2_n160 ), .ZN(N2380) );
INV_X4 _add_1_root_add_513_2_U233  ( .A(_add_1_root_add_513_2_n93 ), .ZN(_add_1_root_add_513_2_n148 ) );
INV_X4 _add_1_root_add_513_2_U232  ( .A(_add_1_root_add_513_2_n94 ), .ZN(_add_1_root_add_513_2_n147 ) );
NAND2_X2 _add_1_root_add_513_2_U231  ( .A1(_add_1_root_add_513_2_n148 ),.A2(_add_1_root_add_513_2_n147 ), .ZN(_add_1_root_add_513_2_n107 ) );
XNOR2_X2 _add_1_root_add_513_2_U230  ( .A(_add_1_root_add_513_2_n157 ), .B(enc_byte_cnt[32]), .ZN(N2381) );
XNOR2_X2 _add_1_root_add_513_2_U229  ( .A(_add_1_root_add_513_2_n18 ), .B(_add_1_root_add_513_2_n151 ), .ZN(N2382) );
XNOR2_X2 _add_1_root_add_513_2_U228  ( .A(_add_1_root_add_513_2_n6 ), .B(_add_1_root_add_513_2_n150 ), .ZN(N2383) );
INV_X4 _add_1_root_add_513_2_U227  ( .A(enc_byte_cnt[35]), .ZN(_add_1_root_add_513_2_n154 ) );
XNOR2_X2 _add_1_root_add_513_2_U226  ( .A(_add_1_root_add_513_2_n34 ), .B(_add_1_root_add_513_2_n154 ), .ZN(N2384) );
NAND2_X2 _add_1_root_add_513_2_U225  ( .A1(_add_1_root_add_513_2_n148 ),.A2(_add_1_root_add_513_2_n15 ), .ZN(_add_1_root_add_513_2_n145 ) );
INV_X4 _add_1_root_add_513_2_U224  ( .A(_add_1_root_add_513_2_n108 ), .ZN(_add_1_root_add_513_2_n78 ) );
NAND2_X2 _add_1_root_add_513_2_U223  ( .A1(_add_1_root_add_513_2_n78 ), .A2(_add_1_root_add_513_2_n147 ), .ZN(_add_1_root_add_513_2_n146 ) );
XNOR2_X2 _add_1_root_add_513_2_U222  ( .A(_add_1_root_add_513_2_n5 ), .B(enc_byte_cnt[36]), .ZN(N2385) );
XNOR2_X2 _add_1_root_add_513_2_U221  ( .A(_add_1_root_add_513_2_n14 ), .B(enc_byte_cnt[37]), .ZN(N2386) );
XNOR2_X2 _add_1_root_add_513_2_U220  ( .A(_add_1_root_add_513_2_n54 ), .B(enc_byte_cnt[38]), .ZN(N2387) );
INV_X4 _add_1_root_add_513_2_U219  ( .A(enc_byte_cnt[39]), .ZN(_add_1_root_add_513_2_n144 ) );
XNOR2_X2 _add_1_root_add_513_2_U218  ( .A(_add_1_root_add_513_2_n33 ), .B(enc_byte_cnt[39]), .ZN(N2388) );
NAND2_X2 _add_1_root_add_513_2_U217  ( .A1(_add_1_root_add_513_2_n143 ),.A2(_add_1_root_add_513_2_n60 ), .ZN(_add_1_root_add_513_2_n141 ) );
NAND2_X2 _add_1_root_add_513_2_U216  ( .A1(_add_1_root_add_513_2_n141 ),.A2(_add_1_root_add_513_2_n142 ), .ZN(_add_1_root_add_513_2_n137 ) );
NAND2_X2 _add_1_root_add_513_2_U215  ( .A1(_add_1_root_add_513_2_n139 ),.A2(_add_1_root_add_513_2_n140 ), .ZN(_add_1_root_add_513_2_n138 ) );
XNOR2_X2 _add_1_root_add_513_2_U214  ( .A(_add_1_root_add_513_2_n137 ), .B(_add_1_root_add_513_2_n138 ), .ZN(N2352) );
INV_X4 _add_1_root_add_513_2_U213  ( .A(_add_1_root_add_513_2_n111 ), .ZN(_add_1_root_add_513_2_n132 ) );
NAND2_X2 _add_1_root_add_513_2_U212  ( .A1(_add_1_root_add_513_2_n132 ),.A2(_add_1_root_add_513_2_n15 ), .ZN(_add_1_root_add_513_2_n131 ) );
XNOR2_X2 _add_1_root_add_513_2_U211  ( .A(_add_1_root_add_513_2_n20 ), .B(enc_byte_cnt[40]), .ZN(N2389) );
INV_X4 _add_1_root_add_513_2_U210  ( .A(_add_1_root_add_513_2_n131 ), .ZN(_add_1_root_add_513_2_n124 ) );
NAND2_X2 _add_1_root_add_513_2_U209  ( .A1(_add_1_root_add_513_2_n124 ),.A2(enc_byte_cnt[40]), .ZN(_add_1_root_add_513_2_n130 ) );
XNOR2_X2 _add_1_root_add_513_2_U208  ( .A(_add_1_root_add_513_2_n19 ), .B(enc_byte_cnt[41]), .ZN(N2390) );
INV_X4 _add_1_root_add_513_2_U207  ( .A(_add_1_root_add_513_2_n130 ), .ZN(_add_1_root_add_513_2_n129 ) );
XNOR2_X2 _add_1_root_add_513_2_U206  ( .A(_add_1_root_add_513_2_n128 ), .B(enc_byte_cnt[42]), .ZN(N2391) );
INV_X4 _add_1_root_add_513_2_U205  ( .A(enc_byte_cnt[43]), .ZN(_add_1_root_add_513_2_n126 ) );
XNOR2_X2 _add_1_root_add_513_2_U204  ( .A(_add_1_root_add_513_2_n22 ), .B(_add_1_root_add_513_2_n126 ), .ZN(N2392) );
NAND4_X2 _add_1_root_add_513_2_U203  ( .A1(enc_byte_cnt[43]), .A2(enc_byte_cnt[42]), .A3(enc_byte_cnt[40]), .A4(enc_byte_cnt[41]), .ZN(_add_1_root_add_513_2_n112 ) );
INV_X4 _add_1_root_add_513_2_U202  ( .A(_add_1_root_add_513_2_n112 ), .ZN(_add_1_root_add_513_2_n125 ) );
NAND2_X2 _add_1_root_add_513_2_U201  ( .A1(_add_1_root_add_513_2_n124 ),.A2(_add_1_root_add_513_2_n125 ), .ZN(_add_1_root_add_513_2_n122 ) );
INV_X4 _add_1_root_add_513_2_U200  ( .A(enc_byte_cnt[44]), .ZN(_add_1_root_add_513_2_n123 ) );
XNOR2_X2 _add_1_root_add_513_2_U199  ( .A(_add_1_root_add_513_2_n31 ), .B(enc_byte_cnt[44]), .ZN(N2393) );
INV_X4 _add_1_root_add_513_2_U198  ( .A(_add_1_root_add_513_2_n122 ), .ZN(_add_1_root_add_513_2_n121 ) );
NAND2_X2 _add_1_root_add_513_2_U197  ( .A1(_add_1_root_add_513_2_n121 ),.A2(enc_byte_cnt[44]), .ZN(_add_1_root_add_513_2_n119 ) );
INV_X4 _add_1_root_add_513_2_U196  ( .A(enc_byte_cnt[45]), .ZN(_add_1_root_add_513_2_n120 ) );
XNOR2_X2 _add_1_root_add_513_2_U195  ( .A(_add_1_root_add_513_2_n45 ), .B(enc_byte_cnt[45]), .ZN(N2394) );
INV_X4 _add_1_root_add_513_2_U194  ( .A(_add_1_root_add_513_2_n119 ), .ZN(_add_1_root_add_513_2_n118 ) );
INV_X4 _add_1_root_add_513_2_U193  ( .A(enc_byte_cnt[46]), .ZN(_add_1_root_add_513_2_n117 ) );
XNOR2_X2 _add_1_root_add_513_2_U192  ( .A(_add_1_root_add_513_2_n116 ), .B(_add_1_root_add_513_2_n117 ), .ZN(N2395) );
INV_X4 _add_1_root_add_513_2_U191  ( .A(enc_byte_cnt[47]), .ZN(_add_1_root_add_513_2_n115 ) );
XNOR2_X2 _add_1_root_add_513_2_U190  ( .A(_add_1_root_add_513_2_n21 ), .B(_add_1_root_add_513_2_n115 ), .ZN(N2396) );
NAND2_X2 _add_1_root_add_513_2_U189  ( .A1(enc_byte_cnt[47]), .A2(enc_byte_cnt[46]), .ZN(_add_1_root_add_513_2_n113 ) );
XNOR2_X2 _add_1_root_add_513_2_U188  ( .A(_add_1_root_add_513_2_n37 ), .B(enc_byte_cnt[48]), .ZN(N2397) );
INV_X4 _add_1_root_add_513_2_U187  ( .A(_add_1_root_add_513_2_n105 ), .ZN(_add_1_root_add_513_2_n92 ) );
INV_X4 _add_1_root_add_513_2_U186  ( .A(_add_1_root_add_513_2_n55 ), .ZN(_add_1_root_add_513_2_n104 ) );
XNOR2_X2 _add_1_root_add_513_2_U185  ( .A(_add_1_root_add_513_2_n104 ), .B(_add_1_root_add_513_2_n101 ), .ZN(N2398) );
XNOR2_X2 _add_1_root_add_513_2_U184  ( .A(_add_1_root_add_513_2_n103 ), .B(_add_1_root_add_513_2_n80 ), .ZN(N2353) );
INV_X4 _add_1_root_add_513_2_U183  ( .A(enc_byte_cnt[49]), .ZN(_add_1_root_add_513_2_n101 ) );
INV_X4 _add_1_root_add_513_2_U182  ( .A(enc_byte_cnt[50]), .ZN(_add_1_root_add_513_2_n102 ) );
XNOR2_X2 _add_1_root_add_513_2_U181  ( .A(_add_1_root_add_513_2_n32 ), .B(_add_1_root_add_513_2_n102 ), .ZN(N2399) );
INV_X4 _add_1_root_add_513_2_U180  ( .A(_add_1_root_add_513_2_n99 ), .ZN(_add_1_root_add_513_2_n100 ) );
XNOR2_X2 _add_1_root_add_513_2_U179  ( .A(_add_1_root_add_513_2_n46 ), .B(enc_byte_cnt[51]), .ZN(N2400) );
NAND2_X2 _add_1_root_add_513_2_U178  ( .A1(_add_1_root_add_513_2_n99 ), .A2(enc_byte_cnt[51]), .ZN(_add_1_root_add_513_2_n98 ) );
XNOR2_X2 _add_1_root_add_513_2_U177  ( .A(_add_1_root_add_513_2_n43 ), .B(enc_byte_cnt[52]), .ZN(N2401) );
INV_X4 _add_1_root_add_513_2_U176  ( .A(_add_1_root_add_513_2_n98 ), .ZN(_add_1_root_add_513_2_n97 ) );
NAND2_X2 _add_1_root_add_513_2_U175  ( .A1(_add_1_root_add_513_2_n97 ), .A2(enc_byte_cnt[52]), .ZN(_add_1_root_add_513_2_n96 ) );
XNOR2_X2 _add_1_root_add_513_2_U174  ( .A(_add_1_root_add_513_2_n8 ), .B(enc_byte_cnt[53]), .ZN(N2402) );
INV_X4 _add_1_root_add_513_2_U173  ( .A(_add_1_root_add_513_2_n96 ), .ZN(_add_1_root_add_513_2_n77 ) );
NAND2_X2 _add_1_root_add_513_2_U172  ( .A1(_add_1_root_add_513_2_n77 ), .A2(_add_1_root_add_513_2_n78 ), .ZN(_add_1_root_add_513_2_n90 ) );
NAND2_X2 _add_1_root_add_513_2_U171  ( .A1(enc_byte_cnt[48]), .A2(enc_byte_cnt[53]), .ZN(_add_1_root_add_513_2_n95 ) );
NAND2_X2 _add_1_root_add_513_2_U170  ( .A1(_add_1_root_add_513_2_n91 ), .A2(_add_1_root_add_513_2_n92 ), .ZN(_add_1_root_add_513_2_n76 ) );
INV_X4 _add_1_root_add_513_2_U169  ( .A(enc_byte_cnt[54]), .ZN(_add_1_root_add_513_2_n89 ) );
XNOR2_X2 _add_1_root_add_513_2_U168  ( .A(_add_1_root_add_513_2_n1 ), .B(enc_byte_cnt[54]), .ZN(N2403) );
INV_X4 _add_1_root_add_513_2_U167  ( .A(enc_byte_cnt[55]), .ZN(_add_1_root_add_513_2_n88 ) );
XNOR2_X2 _add_1_root_add_513_2_U166  ( .A(_add_1_root_add_513_2_n30 ), .B(enc_byte_cnt[55]), .ZN(N2404) );
INV_X4 _add_1_root_add_513_2_U165  ( .A(_add_1_root_add_513_2_n86 ), .ZN(_add_1_root_add_513_2_n87 ) );
XNOR2_X2 _add_1_root_add_513_2_U164  ( .A(_add_1_root_add_513_2_n12 ), .B(enc_byte_cnt[56]), .ZN(N2405) );
NAND2_X2 _add_1_root_add_513_2_U163  ( .A1(_add_1_root_add_513_2_n86 ), .A2(enc_byte_cnt[56]), .ZN(_add_1_root_add_513_2_n85 ) );
XNOR2_X2 _add_1_root_add_513_2_U162  ( .A(_add_1_root_add_513_2_n11 ), .B(enc_byte_cnt[57]), .ZN(N2406) );
INV_X4 _add_1_root_add_513_2_U161  ( .A(_add_1_root_add_513_2_n85 ), .ZN(_add_1_root_add_513_2_n84 ) );
NAND2_X2 _add_1_root_add_513_2_U160  ( .A1(_add_1_root_add_513_2_n84 ), .A2(enc_byte_cnt[57]), .ZN(_add_1_root_add_513_2_n83 ) );
XNOR2_X2 _add_1_root_add_513_2_U159  ( .A(_add_1_root_add_513_2_n10 ), .B(enc_byte_cnt[58]), .ZN(N2407) );
INV_X4 _add_1_root_add_513_2_U158  ( .A(_add_1_root_add_513_2_n83 ), .ZN(_add_1_root_add_513_2_n82 ) );
NAND2_X2 _add_1_root_add_513_2_U157  ( .A1(_add_1_root_add_513_2_n82 ), .A2(enc_byte_cnt[58]), .ZN(_add_1_root_add_513_2_n74 ) );
XNOR2_X2 _add_1_root_add_513_2_U156  ( .A(_add_1_root_add_513_2_n9 ), .B(enc_byte_cnt[59]), .ZN(N2408) );
XNOR2_X2 _add_1_root_add_513_2_U155  ( .A(_add_1_root_add_513_2_n81 ), .B(_add_1_root_add_513_2_n16 ), .ZN(N2354) );
INV_X4 _add_1_root_add_513_2_U154  ( .A(enc_byte_cnt[60]), .ZN(_add_1_root_add_513_2_n79 ) );
NAND2_X2 _add_1_root_add_513_2_U153  ( .A1(_add_1_root_add_513_2_n77 ), .A2(_add_1_root_add_513_2_n78 ), .ZN(_add_1_root_add_513_2_n75 ) );
INV_X4 _add_1_root_add_513_2_U152  ( .A(_add_1_root_add_513_2_n74 ), .ZN(_add_1_root_add_513_2_n73 ) );
NAND2_X2 _add_1_root_add_513_2_U151  ( .A1(_add_1_root_add_513_2_n73 ), .A2(enc_byte_cnt[59]), .ZN(_add_1_root_add_513_2_n70 ) );
XNOR2_X2 _add_1_root_add_513_2_U150  ( .A(_add_1_root_add_513_2_n79 ), .B(_add_1_root_add_513_2_n17 ), .ZN(N2409) );
INV_X4 _add_1_root_add_513_2_U149  ( .A(enc_byte_cnt[61]), .ZN(_add_1_root_add_513_2_n72 ) );
XNOR2_X2 _add_1_root_add_513_2_U148  ( .A(_add_1_root_add_513_2_n27 ), .B(_add_1_root_add_513_2_n72 ), .ZN(N2410) );
INV_X4 _add_1_root_add_513_2_U147  ( .A(enc_byte_cnt[62]), .ZN(_add_1_root_add_513_2_n71 ) );
XNOR2_X2 _add_1_root_add_513_2_U146  ( .A(_add_1_root_add_513_2_n25 ), .B(_add_1_root_add_513_2_n71 ), .ZN(N2411) );
NAND2_X2 _add_1_root_add_513_2_U145  ( .A1(_add_1_root_add_513_2_n69 ), .A2(enc_byte_cnt[62]), .ZN(_add_1_root_add_513_2_n68 ) );
NAND2_X2 _add_1_root_add_513_2_U144  ( .A1(_add_1_root_add_513_2_n16 ), .A2(enc_byte_cnt[5]), .ZN(_add_1_root_add_513_2_n66 ) );
XNOR2_X2 _add_1_root_add_513_2_U143  ( .A(_add_1_root_add_513_2_n66 ), .B(enc_byte_cnt[6]), .ZN(N2355) );
XNOR2_X2 _add_1_root_add_513_2_U142  ( .A(_add_1_root_add_513_2_n29 ), .B(enc_byte_cnt[7]), .ZN(N2356) );
XNOR2_X2 _add_1_root_add_513_2_U141  ( .A(_add_1_root_add_513_2_n63 ), .B(_add_1_root_add_513_2_n64 ), .ZN(N2357) );
XNOR2_X2 _add_1_root_add_513_2_U140  ( .A(_add_1_root_add_513_2_n58 ), .B(enc_byte_cnt[9]), .ZN(N2358) );
INV_X4 _add_1_root_add_513_2_U139  ( .A(enc_byte_cnt[38]), .ZN(_add_1_root_add_513_2_n134 ) );
INV_X4 _add_1_root_add_513_2_U138  ( .A(enc_byte_cnt[37]), .ZN(_add_1_root_add_513_2_n136 ) );
INV_X4 _add_1_root_add_513_2_U137  ( .A(enc_byte_cnt[36]), .ZN(_add_1_root_add_513_2_n135 ) );
INV_X4 _add_1_root_add_513_2_U136  ( .A(enc_byte_cnt[34]), .ZN(_add_1_root_add_513_2_n150 ) );
INV_X4 _add_1_root_add_513_2_U135  ( .A(enc_byte_cnt[33]), .ZN(_add_1_root_add_513_2_n151 ) );
INV_X4 _add_1_root_add_513_2_U134  ( .A(enc_byte_cnt[32]), .ZN(_add_1_root_add_513_2_n156 ) );
INV_X4 _add_1_root_add_513_2_U133  ( .A(enc_byte_cnt[26]), .ZN(_add_1_root_add_513_2_n169 ) );
INV_X4 _add_1_root_add_513_2_U132  ( .A(enc_byte_cnt[25]), .ZN(_add_1_root_add_513_2_n171 ) );
INV_X4 _add_1_root_add_513_2_U131  ( .A(enc_byte_cnt[24]), .ZN(_add_1_root_add_513_2_n170 ) );
INV_X4 _add_1_root_add_513_2_U130  ( .A(enc_byte_cnt[23]), .ZN(_add_1_root_add_513_2_n175 ) );
INV_X4 _add_1_root_add_513_2_U129  ( .A(enc_byte_cnt[22]), .ZN(_add_1_root_add_513_2_n174 ) );
INV_X4 _add_1_root_add_513_2_U128  ( .A(enc_byte_cnt[21]), .ZN(_add_1_root_add_513_2_n176 ) );
INV_X4 _add_1_root_add_513_2_U127  ( .A(enc_byte_cnt[20]), .ZN(_add_1_root_add_513_2_n179 ) );
INV_X4 _add_1_root_add_513_2_U126  ( .A(enc_byte_cnt[18]), .ZN(_add_1_root_add_513_2_n181 ) );
INV_X4 _add_1_root_add_513_2_U125  ( .A(enc_byte_cnt[17]), .ZN(_add_1_root_add_513_2_n189 ) );
INV_X4 _add_1_root_add_513_2_U124  ( .A(enc_byte_cnt[16]), .ZN(_add_1_root_add_513_2_n182 ) );
INV_X4 _add_1_root_add_513_2_U123  ( .A(enc_byte_cnt[10]), .ZN(_add_1_root_add_513_2_n206 ) );
INV_X4 _add_1_root_add_513_2_U122  ( .A(enc_byte_cnt[9]), .ZN(_add_1_root_add_513_2_n62 ) );
INV_X4 _add_1_root_add_513_2_U121  ( .A(enc_byte_cnt[8]), .ZN(_add_1_root_add_513_2_n64 ) );
INV_X4 _add_1_root_add_513_2_U120  ( .A(enc_byte_cnt[6]), .ZN(_add_1_root_add_513_2_n65 ) );
INV_X4 _add_1_root_add_513_2_U119  ( .A(enc_byte_cnt[4]), .ZN(_add_1_root_add_513_2_n103 ) );
INV_X4 _add_1_root_add_513_2_U118  ( .A(enc_byte_cnt[5]), .ZN(_add_1_root_add_513_2_n81 ) );
INV_X4 _add_1_root_add_513_2_U117  ( .A(_add_1_root_add_513_2_n186 ), .ZN(_add_1_root_add_513_2_n210 ) );
INV_X4 _add_1_root_add_513_2_U116  ( .A(_add_1_root_add_513_2_n114 ), .ZN(_add_1_root_add_513_2_n157 ) );
INV_X4 _add_1_root_add_513_2_U115  ( .A(_add_1_root_add_513_2_n127 ), .ZN(_add_1_root_add_513_2_n128 ) );
INV_X4 _add_1_root_add_513_2_U114  ( .A(_add_1_root_add_513_2_n208 ), .ZN(_add_1_root_add_513_2_n63 ) );
NOR2_X2 _add_1_root_add_513_2_U113  ( .A1(_add_1_root_add_513_2_n184 ), .A2(_add_1_root_add_513_2_n165 ), .ZN(_add_1_root_add_513_2_n183 ) );
OR2_X2 _add_1_root_add_513_2_U112  ( .A1(enc_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(_add_1_root_add_513_2_n60 ) );
NOR2_X2 _add_1_root_add_513_2_U111  ( .A1(_add_1_root_add_513_2_n44 ), .A2(_add_1_root_add_513_2_n68 ), .ZN(_add_1_root_add_513_2_n67 ) );
XOR2_X2 _add_1_root_add_513_2_U110  ( .A(_add_1_root_add_513_2_n67 ), .B(enc_byte_cnt[63]), .Z(N2412) );
AND2_X2 _add_1_root_add_513_2_U109  ( .A1(enc_byte_cnt[0]), .A2(n17750),.ZN(_add_1_root_add_513_2_n219 ) );
NOR2_X2 _add_1_root_add_513_2_U108  ( .A1(_add_1_root_add_513_2_n217 ), .A2(_add_1_root_add_513_2_n218 ), .ZN(_add_1_root_add_513_2_n216 ) );
NAND3_X2 _add_1_root_add_513_2_U107  ( .A1(dii_data_size[1]), .A2(_add_1_root_add_513_2_n60 ), .A3(enc_byte_cnt[1]), .ZN(_add_1_root_add_513_2_n215 ) );
NAND3_X2 _add_1_root_add_513_2_U106  ( .A1(_add_1_root_add_513_2_n214 ),.A2(_add_1_root_add_513_2_n215 ), .A3(_add_1_root_add_513_2_n216 ),.ZN(_add_1_root_add_513_2_n193 ) );
NOR2_X2 _add_1_root_add_513_2_U105  ( .A1(enc_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(_add_1_root_add_513_2_n222 ) );
NOR2_X2 _add_1_root_add_513_2_U104  ( .A1(enc_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(_add_1_root_add_513_2_n221 ) );
NOR2_X2 _add_1_root_add_513_2_U103  ( .A1(_add_1_root_add_513_2_n221 ), .A2(_add_1_root_add_513_2_n222 ), .ZN(_add_1_root_add_513_2_n220 ) );
NOR2_X2 _add_1_root_add_513_2_U102  ( .A1(enc_byte_cnt[0]), .A2(n17750),.ZN(_add_1_root_add_513_2_n186 ) );
NOR2_X2 _add_1_root_add_513_2_U101  ( .A1(enc_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(_add_1_root_add_513_2_n165 ) );
INV_X4 _add_1_root_add_513_2_U100  ( .A(n18074), .ZN(_add_1_root_add_513_2_n61 ) );
AND2_X2 _add_1_root_add_513_2_U99  ( .A1(_add_1_root_add_513_2_n186 ), .A2(_add_1_root_add_513_2_n185 ), .ZN(_add_1_root_add_513_2_n166 ) );
NOR2_X2 _add_1_root_add_513_2_U98  ( .A1(_add_1_root_add_513_2_n154 ), .A2(_add_1_root_add_513_2_n150 ), .ZN(_add_1_root_add_513_2_n149 ) );
OR2_X2 _add_1_root_add_513_2_U97  ( .A1(_add_1_root_add_513_2_n58 ), .A2(_add_1_root_add_513_2_n62 ), .ZN(_add_1_root_add_513_2_n59 ) );
NOR2_X2 _add_1_root_add_513_2_U96  ( .A1(_add_1_root_add_513_2_n134 ), .A2(_add_1_root_add_513_2_n144 ), .ZN(_add_1_root_add_513_2_n133 ) );
NAND3_X2 _add_1_root_add_513_2_U95  ( .A1(enc_byte_cnt[37]), .A2(enc_byte_cnt[36]), .A3(_add_1_root_add_513_2_n133 ), .ZN(_add_1_root_add_513_2_n111 ) );
OR2_X2 _add_1_root_add_513_2_U94  ( .A1(_add_1_root_add_513_2_n208 ), .A2(_add_1_root_add_513_2_n64 ), .ZN(_add_1_root_add_513_2_n58 ) );
NOR2_X2 _add_1_root_add_513_2_U93  ( .A1(_add_1_root_add_513_2_n167 ), .A2(_add_1_root_add_513_2_n159 ), .ZN(_add_1_root_add_513_2_n158 ) );
NAND3_X2 _add_1_root_add_513_2_U92  ( .A1(enc_byte_cnt[30]), .A2(enc_byte_cnt[31]), .A3(_add_1_root_add_513_2_n158 ), .ZN(_add_1_root_add_513_2_n93 ) );
NOR2_X2 _add_1_root_add_513_2_U91  ( .A1(_add_1_root_add_513_2_n151 ), .A2(_add_1_root_add_513_2_n156 ), .ZN(_add_1_root_add_513_2_n155 ) );
AND2_X2 _add_1_root_add_513_2_U90  ( .A1(enc_byte_cnt[61]), .A2(enc_byte_cnt[60]), .ZN(_add_1_root_add_513_2_n69 ) );
NOR2_X2 _add_1_root_add_513_2_U89  ( .A1(_add_1_root_add_513_2_n169 ), .A2(_add_1_root_add_513_2_n172 ), .ZN(_add_1_root_add_513_2_n168 ) );
NAND3_X2 _add_1_root_add_513_2_U88  ( .A1(enc_byte_cnt[25]), .A2(enc_byte_cnt[24]), .A3(_add_1_root_add_513_2_n168 ), .ZN(_add_1_root_add_513_2_n94 ) );
NOR2_X2 _add_1_root_add_513_2_U87  ( .A1(_add_1_root_add_513_2_n102 ), .A2(_add_1_root_add_513_2_n101 ), .ZN(_add_1_root_add_513_2_n99 ) );
NOR2_X2 _add_1_root_add_513_2_U86  ( .A1(_add_1_root_add_513_2_n88 ), .A2(_add_1_root_add_513_2_n89 ), .ZN(_add_1_root_add_513_2_n86 ) );
NOR2_X2 _add_1_root_add_513_2_U85  ( .A1(_add_1_root_add_513_2_n187 ), .A2(_add_1_root_add_513_2_n181 ), .ZN(_add_1_root_add_513_2_n180 ) );
NAND3_X2 _add_1_root_add_513_2_U84  ( .A1(enc_byte_cnt[16]), .A2(enc_byte_cnt[17]), .A3(_add_1_root_add_513_2_n180 ), .ZN(_add_1_root_add_513_2_n153 ) );
NOR2_X2 _add_1_root_add_513_2_U83  ( .A1(_add_1_root_add_513_2_n174 ), .A2(_add_1_root_add_513_2_n175 ), .ZN(_add_1_root_add_513_2_n173 ) );
NAND3_X2 _add_1_root_add_513_2_U82  ( .A1(enc_byte_cnt[21]), .A2(enc_byte_cnt[20]), .A3(_add_1_root_add_513_2_n173 ), .ZN(_add_1_root_add_513_2_n108 ) );
OR2_X2 _add_1_root_add_513_2_U81  ( .A1(_add_1_root_add_513_2_n165 ), .A2(_add_1_root_add_513_2_n166 ), .ZN(_add_1_root_add_513_2_n57 ) );
NOR3_X2 _add_1_root_add_513_2_U80  ( .A1(_add_1_root_add_513_2_n93 ), .A2(_add_1_root_add_513_2_n94 ), .A3(_add_1_root_add_513_2_n95 ), .ZN(_add_1_root_add_513_2_n91 ) );
AND2_X4 _add_1_root_add_513_2_U79  ( .A1(_add_1_root_add_513_2_n92 ), .A2(enc_byte_cnt[48]), .ZN(_add_1_root_add_513_2_n56 ) );
NAND2_X2 _add_1_root_add_513_2_U78  ( .A1(_add_1_root_add_513_2_n106 ), .A2(_add_1_root_add_513_2_n56 ), .ZN(_add_1_root_add_513_2_n55 ) );
NOR2_X2 _add_1_root_add_513_2_U77  ( .A1(_add_1_root_add_513_2_n212 ), .A2(_add_1_root_add_513_2_n165 ), .ZN(_add_1_root_add_513_2_n211 ) );
NAND3_X2 _add_1_root_add_513_2_U76  ( .A1(_add_1_root_add_513_2_n210 ), .A2(_add_1_root_add_513_2_n60 ), .A3(_add_1_root_add_513_2_n211 ), .ZN(_add_1_root_add_513_2_n200 ) );
OR3_X2 _add_1_root_add_513_2_U75  ( .A1(_add_1_root_add_513_2_n5 ), .A2(_add_1_root_add_513_2_n135 ), .A3(_add_1_root_add_513_2_n136 ), .ZN(_add_1_root_add_513_2_n54 ) );
OR3_X2 _add_1_root_add_513_2_U74  ( .A1(_add_1_root_add_513_2_n42 ), .A2(_add_1_root_add_513_2_n167 ), .A3(_add_1_root_add_513_2_n159 ), .ZN(_add_1_root_add_513_2_n53 ) );
NOR2_X2 _add_1_root_add_513_2_U73  ( .A1(_add_1_root_add_513_2_n65 ), .A2(_add_1_root_add_513_2_n224 ), .ZN(_add_1_root_add_513_2_n223 ) );
NAND3_X2 _add_1_root_add_513_2_U72  ( .A1(enc_byte_cnt[5]), .A2(enc_byte_cnt[4]), .A3(_add_1_root_add_513_2_n223 ), .ZN(_add_1_root_add_513_2_n198 ) );
OR2_X2 _add_1_root_add_513_2_U71  ( .A1(_add_1_root_add_513_2_n159 ), .A2(_add_1_root_add_513_2_n42 ), .ZN(_add_1_root_add_513_2_n52 ) );
OR2_X2 _add_1_root_add_513_2_U70  ( .A1(_add_1_root_add_513_2_n176 ), .A2(_add_1_root_add_513_2_n177 ), .ZN(_add_1_root_add_513_2_n51 ) );
OR2_X2 _add_1_root_add_513_2_U69  ( .A1(_add_1_root_add_513_2_n171 ), .A2(_add_1_root_add_513_2_n49 ), .ZN(_add_1_root_add_513_2_n50 ) );
OR2_X2 _add_1_root_add_513_2_U68  ( .A1(_add_1_root_add_513_2_n170 ), .A2(_add_1_root_add_513_2_n38 ), .ZN(_add_1_root_add_513_2_n49 ) );
OR2_X2 _add_1_root_add_513_2_U67  ( .A1(_add_1_root_add_513_2_n181 ), .A2(_add_1_root_add_513_2_n188 ), .ZN(_add_1_root_add_513_2_n48 ) );
AND2_X2 _add_1_root_add_513_2_U66  ( .A1(enc_byte_cnt[13]), .A2(enc_byte_cnt[12]), .ZN(_add_1_root_add_513_2_n199 ) );
AND2_X4 _add_1_root_add_513_2_U65  ( .A1(_add_1_root_add_513_2_n118 ), .A2(enc_byte_cnt[45]), .ZN(_add_1_root_add_513_2_n47 ) );
AND2_X2 _add_1_root_add_513_2_U64  ( .A1(_add_1_root_add_513_2_n114 ), .A2(_add_1_root_add_513_2_n47 ), .ZN(_add_1_root_add_513_2_n116 ) );
NOR2_X2 _add_1_root_add_513_2_U63  ( .A1(_add_1_root_add_513_2_n206 ), .A2(_add_1_root_add_513_2_n207 ), .ZN(_add_1_root_add_513_2_n205 ) );
NAND3_X2 _add_1_root_add_513_2_U62  ( .A1(enc_byte_cnt[9]), .A2(enc_byte_cnt[8]), .A3(_add_1_root_add_513_2_n205 ), .ZN(_add_1_root_add_513_2_n192 ) );
NAND3_X2 _add_1_root_add_513_2_U61  ( .A1(_add_1_root_add_513_2_n140 ), .A2(_add_1_root_add_513_2_n193 ), .A3(_add_1_root_add_513_2_n194 ), .ZN(_add_1_root_add_513_2_n190 ) );
NOR2_X2 _add_1_root_add_513_2_U60  ( .A1(_add_1_root_add_513_2_n111 ), .A2(_add_1_root_add_513_2_n112 ), .ZN(_add_1_root_add_513_2_n110 ) );
NOR3_X2 _add_1_root_add_513_2_U59  ( .A1(_add_1_root_add_513_2_n113 ), .A2(_add_1_root_add_513_2_n120 ), .A3(_add_1_root_add_513_2_n123 ), .ZN(_add_1_root_add_513_2_n109 ) );
NAND3_X2 _add_1_root_add_513_2_U58  ( .A1(_add_1_root_add_513_2_n109 ), .A2(_add_1_root_add_513_2_n15 ), .A3(_add_1_root_add_513_2_n110 ), .ZN(_add_1_root_add_513_2_n105 ) );
OR2_X2 _add_1_root_add_513_2_U57  ( .A1(_add_1_root_add_513_2_n55 ), .A2(_add_1_root_add_513_2_n100 ), .ZN(_add_1_root_add_513_2_n46 ) );
OR2_X2 _add_1_root_add_513_2_U56  ( .A1(_add_1_root_add_513_2_n157 ), .A2(_add_1_root_add_513_2_n119 ), .ZN(_add_1_root_add_513_2_n45 ) );
AND2_X2 _add_1_root_add_513_2_U55  ( .A1(_add_1_root_add_513_2_n195 ), .A2(_add_1_root_add_513_2_n36 ), .ZN(_add_1_root_add_513_2_n152 ) );
OR2_X2 _add_1_root_add_513_2_U54  ( .A1(_add_1_root_add_513_2_n1 ), .A2(_add_1_root_add_513_2_n70 ), .ZN(_add_1_root_add_513_2_n44 ) );
NOR2_X2 _add_1_root_add_513_2_U53  ( .A1(_add_1_root_add_513_2_n198 ), .A2(_add_1_root_add_513_2_n191 ), .ZN(_add_1_root_add_513_2_n197 ) );
NOR2_X2 _add_1_root_add_513_2_U52  ( .A1(_add_1_root_add_513_2_n192 ), .A2(_add_1_root_add_513_2_n200 ), .ZN(_add_1_root_add_513_2_n196 ) );
OR2_X2 _add_1_root_add_513_2_U51  ( .A1(_add_1_root_add_513_2_n55 ), .A2(_add_1_root_add_513_2_n98 ), .ZN(_add_1_root_add_513_2_n43 ) );
OR2_X2 _add_1_root_add_513_2_U50  ( .A1(_add_1_root_add_513_2_n38 ), .A2(_add_1_root_add_513_2_n94 ), .ZN(_add_1_root_add_513_2_n42 ) );
OR2_X2 _add_1_root_add_513_2_U49  ( .A1(_add_1_root_add_513_2_n152 ), .A2(_add_1_root_add_513_2_n153 ), .ZN(_add_1_root_add_513_2_n41 ) );
OR2_X2 _add_1_root_add_513_2_U48  ( .A1(_add_1_root_add_513_2_n152 ), .A2(_add_1_root_add_513_2_n153 ), .ZN(_add_1_root_add_513_2_n40 ) );
AND2_X4 _add_1_root_add_513_2_U47  ( .A1(_add_1_root_add_513_2_n129 ), .A2(enc_byte_cnt[41]), .ZN(_add_1_root_add_513_2_n39 ) );
AND2_X2 _add_1_root_add_513_2_U46  ( .A1(_add_1_root_add_513_2_n114 ), .A2(_add_1_root_add_513_2_n39 ), .ZN(_add_1_root_add_513_2_n127 ) );
OR3_X2 _add_1_root_add_513_2_U45  ( .A1(_add_1_root_add_513_2_n152 ), .A2(_add_1_root_add_513_2_n153 ), .A3(_add_1_root_add_513_2_n108 ), .ZN(_add_1_root_add_513_2_n38 ) );
NOR3_X2 _add_1_root_add_513_2_U44  ( .A1(_add_1_root_add_513_2_n40 ), .A2(_add_1_root_add_513_2_n107 ), .A3(_add_1_root_add_513_2_n108 ), .ZN(_add_1_root_add_513_2_n106 ) );
NOR3_X2 _add_1_root_add_513_2_U43  ( .A1(_add_1_root_add_513_2_n107 ), .A2(_add_1_root_add_513_2_n41 ), .A3(_add_1_root_add_513_2_n108 ), .ZN(_add_1_root_add_513_2_n114 ) );
OR2_X2 _add_1_root_add_513_2_U42  ( .A1(_add_1_root_add_513_2_n157 ), .A2(_add_1_root_add_513_2_n105 ), .ZN(_add_1_root_add_513_2_n37 ) );
XNOR2_X1 _add_1_root_add_513_2_U41  ( .A(_add_1_root_add_513_2_n163 ), .B(_add_1_root_add_513_2_n143 ), .ZN(N2351) );
NAND2_X1 _add_1_root_add_513_2_U40  ( .A1(n17750), .A2(enc_byte_cnt[0]),.ZN(_add_1_root_add_513_2_n185 ) );
NAND2_X1 _add_1_root_add_513_2_U39  ( .A1(_add_1_root_add_513_2_n185 ), .A2(_add_1_root_add_513_2_n210 ), .ZN(N2349) );
OR3_X4 _add_1_root_add_513_2_U38  ( .A1(_add_1_root_add_513_2_n190 ), .A2(_add_1_root_add_513_2_n191 ), .A3(_add_1_root_add_513_2_n192 ), .ZN(_add_1_root_add_513_2_n36 ) );
OR3_X4 _add_1_root_add_513_2_U37  ( .A1(_add_1_root_add_513_2_n40 ), .A2(_add_1_root_add_513_2_n75 ), .A3(_add_1_root_add_513_2_n76 ), .ZN(_add_1_root_add_513_2_n35 ) );
AND2_X4 _add_1_root_add_513_2_U36  ( .A1(_add_1_root_add_513_2_n6 ), .A2(enc_byte_cnt[34]), .ZN(_add_1_root_add_513_2_n34 ) );
OR2_X4 _add_1_root_add_513_2_U35  ( .A1(_add_1_root_add_513_2_n134 ), .A2(_add_1_root_add_513_2_n54 ), .ZN(_add_1_root_add_513_2_n33 ) );
NOR2_X2 _add_1_root_add_513_2_U34  ( .A1(_add_1_root_add_513_2_n101 ), .A2(_add_1_root_add_513_2_n55 ), .ZN(_add_1_root_add_513_2_n32 ) );
OR2_X4 _add_1_root_add_513_2_U33  ( .A1(_add_1_root_add_513_2_n157 ), .A2(_add_1_root_add_513_2_n122 ), .ZN(_add_1_root_add_513_2_n31 ) );
OR2_X4 _add_1_root_add_513_2_U32  ( .A1(_add_1_root_add_513_2_n89 ), .A2(_add_1_root_add_513_2_n1 ), .ZN(_add_1_root_add_513_2_n30 ) );
OR2_X4 _add_1_root_add_513_2_U31  ( .A1(_add_1_root_add_513_2_n65 ), .A2(_add_1_root_add_513_2_n66 ), .ZN(_add_1_root_add_513_2_n29 ) );
OR2_X4 _add_1_root_add_513_2_U30  ( .A1(_add_1_root_add_513_2_n206 ), .A2(_add_1_root_add_513_2_n59 ), .ZN(_add_1_root_add_513_2_n28 ) );
AND2_X4 _add_1_root_add_513_2_U29  ( .A1(enc_byte_cnt[60]), .A2(_add_1_root_add_513_2_n17 ), .ZN(_add_1_root_add_513_2_n27 ) );
AND2_X4 _add_1_root_add_513_2_U28  ( .A1(enc_byte_cnt[14]), .A2(_add_1_root_add_513_2_n7 ), .ZN(_add_1_root_add_513_2_n26 ) );
AND2_X4 _add_1_root_add_513_2_U27  ( .A1(_add_1_root_add_513_2_n69 ), .A2(_add_1_root_add_513_2_n17 ), .ZN(_add_1_root_add_513_2_n25 ) );
OR2_X4 _add_1_root_add_513_2_U26  ( .A1(_add_1_root_add_513_2_n169 ), .A2(_add_1_root_add_513_2_n50 ), .ZN(_add_1_root_add_513_2_n24 ) );
OR2_X4 _add_1_root_add_513_2_U25  ( .A1(_add_1_root_add_513_2_n174 ), .A2(_add_1_root_add_513_2_n51 ), .ZN(_add_1_root_add_513_2_n23 ) );
AND2_X4 _add_1_root_add_513_2_U24  ( .A1(_add_1_root_add_513_2_n127 ), .A2(enc_byte_cnt[42]), .ZN(_add_1_root_add_513_2_n22 ) );
AND2_X4 _add_1_root_add_513_2_U23  ( .A1(_add_1_root_add_513_2_n116 ), .A2(enc_byte_cnt[46]), .ZN(_add_1_root_add_513_2_n21 ) );
OR2_X4 _add_1_root_add_513_2_U22  ( .A1(_add_1_root_add_513_2_n157 ), .A2(_add_1_root_add_513_2_n131 ), .ZN(_add_1_root_add_513_2_n20 ) );
OR2_X4 _add_1_root_add_513_2_U21  ( .A1(_add_1_root_add_513_2_n157 ), .A2(_add_1_root_add_513_2_n130 ), .ZN(_add_1_root_add_513_2_n19 ) );
AND2_X4 _add_1_root_add_513_2_U20  ( .A1(_add_1_root_add_513_2_n114 ), .A2(enc_byte_cnt[32]), .ZN(_add_1_root_add_513_2_n18 ) );
NOR2_X2 _add_1_root_add_513_2_U19  ( .A1(_add_1_root_add_513_2_n35 ), .A2(_add_1_root_add_513_2_n70 ), .ZN(_add_1_root_add_513_2_n17 ) );
AND2_X4 _add_1_root_add_513_2_U18  ( .A1(enc_byte_cnt[4]), .A2(_add_1_root_add_513_2_n80 ), .ZN(_add_1_root_add_513_2_n16 ) );
AND3_X4 _add_1_root_add_513_2_U17  ( .A1(enc_byte_cnt[32]), .A2(enc_byte_cnt[33]), .A3(_add_1_root_add_513_2_n149 ), .ZN(_add_1_root_add_513_2_n15 ) );
OR2_X4 _add_1_root_add_513_2_U16  ( .A1(_add_1_root_add_513_2_n135 ), .A2(_add_1_root_add_513_2_n5 ), .ZN(_add_1_root_add_513_2_n14 ) );
NOR2_X2 _add_1_root_add_513_2_U15  ( .A1(_add_1_root_add_513_2_n162 ), .A2(_add_1_root_add_513_2_n53 ), .ZN(_add_1_root_add_513_2_n13 ) );
OR2_X4 _add_1_root_add_513_2_U14  ( .A1(_add_1_root_add_513_2_n1 ), .A2(_add_1_root_add_513_2_n87 ), .ZN(_add_1_root_add_513_2_n12 ) );
OR2_X4 _add_1_root_add_513_2_U13  ( .A1(_add_1_root_add_513_2_n1 ), .A2(_add_1_root_add_513_2_n85 ), .ZN(_add_1_root_add_513_2_n11 ) );
OR2_X4 _add_1_root_add_513_2_U12  ( .A1(_add_1_root_add_513_2_n1 ), .A2(_add_1_root_add_513_2_n83 ), .ZN(_add_1_root_add_513_2_n10 ) );
OR2_X4 _add_1_root_add_513_2_U11  ( .A1(_add_1_root_add_513_2_n1 ), .A2(_add_1_root_add_513_2_n74 ), .ZN(_add_1_root_add_513_2_n9 ) );
OR2_X4 _add_1_root_add_513_2_U10  ( .A1(_add_1_root_add_513_2_n55 ), .A2(_add_1_root_add_513_2_n96 ), .ZN(_add_1_root_add_513_2_n8 ) );
AND2_X4 _add_1_root_add_513_2_U9  ( .A1(_add_1_root_add_513_2_n4 ), .A2(enc_byte_cnt[13]), .ZN(_add_1_root_add_513_2_n7 ) );
AND2_X4 _add_1_root_add_513_2_U8  ( .A1(_add_1_root_add_513_2_n114 ), .A2(_add_1_root_add_513_2_n155 ), .ZN(_add_1_root_add_513_2_n6 ) );
OR3_X4 _add_1_root_add_513_2_U7  ( .A1(_add_1_root_add_513_2_n40 ), .A2(_add_1_root_add_513_2_n145 ), .A3(_add_1_root_add_513_2_n146 ), .ZN(_add_1_root_add_513_2_n5 ) );
AND2_X4 _add_1_root_add_513_2_U6  ( .A1(_add_1_root_add_513_2_n3 ), .A2(enc_byte_cnt[12]), .ZN(_add_1_root_add_513_2_n4 ) );
NOR2_X2 _add_1_root_add_513_2_U5  ( .A1(_add_1_root_add_513_2_n208 ), .A2(_add_1_root_add_513_2_n192 ), .ZN(_add_1_root_add_513_2_n3 ) );
NOR2_X2 _add_1_root_add_513_2_U4  ( .A1(_add_1_root_add_513_2_n152 ), .A2(_add_1_root_add_513_2_n182 ), .ZN(_add_1_root_add_513_2_n2 ) );
OR3_X4 _add_1_root_add_513_2_U3  ( .A1(_add_1_root_add_513_2_n40 ), .A2(_add_1_root_add_513_2_n90 ), .A3(_add_1_root_add_513_2_n76 ), .ZN(_add_1_root_add_513_2_n1 ) );
NAND3_X2 _add_1_root_add_513_2_U2  ( .A1(enc_byte_cnt[14]), .A2(enc_byte_cnt[15]), .A3(_add_1_root_add_513_2_n199 ), .ZN(_add_1_root_add_513_2_n191 ) );
endmodule
