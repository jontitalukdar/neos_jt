module b22(clock, reset, si, so, rd, wr, d_out_1, qn_in_1, d_out_2, qn_in_2, d_out_3, q_in_3, d_out_4, q_in_4, d_out_5, q_in_5, d_out_6, q_in_6, d_out_7, qn_in_7, d_out_8, qn_in_8, d_out_9, q_in_9, d_out_10, q_in_10, d_out_11, q_in_11, d_out_12, q_in_12, d_out_13, q_in_13, d_out_14, q_in_14, d_out_15, q_in_15, d_out_16, q_in_16, d_out_17, qn_in_17, d_out_18, q_in_18, d_out_19, q_in_19, d_out_20, q_in_20, d_out_21, qn_in_21, d_out_22, q_in_22, d_out_23, qn_in_23, d_out_24, qn_in_24, d_out_25, qn_in_25, d_out_26, qn_in_26, d_out_27, q_in_27, d_out_28, q_in_28, d_out_29, q_in_29, d_out_30, q_in_30, d_out_31, q_in_31, d_out_32, qn_in_32, d_out_33, q_in_33, d_out_34, q_in_34, d_out_35, qn_in_35, d_out_36, qn_in_36, d_out_37, qn_in_37, d_out_38, qn_in_38, d_out_39, q_in_39, d_out_40, q_in_40, d_out_41, q_in_41, d_out_42, q_in_42, d_out_43, qn_in_43, d_out_44, q_in_44, d_out_45, q_in_45, d_out_46, qn_in_46, d_out_47, qn_in_47, d_out_48, qn_in_48, d_out_49, qn_in_49, d_out_50, qn_in_50, d_out_51, qn_in_51, d_out_52, q_in_52, d_out_53, q_in_53, d_out_54, q_in_54, d_out_55, q_in_55, d_out_56, q_in_56, d_out_57, q_in_57, d_out_58, q_in_58, d_out_59, q_in_59, d_out_60, q_in_60, d_out_61, qn_in_61, d_out_62, q_in_62, d_out_63, q_in_63, d_out_64, q_in_64, d_out_65, q_in_65, d_out_66, q_in_66, d_out_67, q_in_67, d_out_68, q_in_68, d_out_69, q_in_69, d_out_70, q_in_70, d_out_71, q_in_71, d_out_72, q_in_72, d_out_73, q_in_73, d_out_74, q_in_74, d_out_75, q_in_75, d_out_76, q_in_76, d_out_77, q_in_77, d_out_78, q_in_78, d_out_79, q_in_79, d_out_80, q_in_80, d_out_81, q_in_81, d_out_82, q_in_82, d_out_83, q_in_83, d_out_84, qn_in_84, d_out_85, qn_in_85, d_out_86, qn_in_86, d_out_87, q_in_87, d_out_88, qn_in_88, d_out_89, q_in_89, d_out_90, q_in_90, d_out_91, q_in_91, d_out_92, q_in_92, d_out_93, q_in_93, d_out_94, q_in_94, d_out_95, q_in_95, d_out_96, q_in_96, d_out_97, q_in_97, d_out_98, q_in_98, d_out_99, q_in_99, d_out_100, q_in_100, d_out_101, q_in_101, d_out_102, q_in_102, d_out_103, q_in_103, d_out_104, q_in_104, d_out_105, q_in_105, d_out_106, q_in_106, d_out_107, q_in_107, d_out_108, q_in_108, d_out_109, q_in_109, d_out_110, q_in_110, d_out_111, q_in_111, d_out_112, qn_in_112, d_out_113, q_in_113, d_out_114, q_in_114, d_out_115, q_in_115, d_out_116, q_in_116, d_out_117, q_in_117, d_out_118, q_in_118, d_out_119, q_in_119, d_out_120, q_in_120, d_out_121, q_in_121, d_out_122, q_in_122, d_out_123, q_in_123, d_out_124, q_in_124, d_out_125, q_in_125, d_out_126, q_in_126, d_out_127, q_in_127, d_out_128, q_in_128, d_out_129, q_in_129, d_out_130, q_in_130, d_out_131, q_in_131, d_out_132, q_in_132, d_out_133, q_in_133, d_out_134, q_in_134, d_out_135, q_in_135, d_out_136, q_in_136, d_out_137, q_in_137, d_out_138, q_in_138, d_out_139, qn_in_139, d_out_140, q_in_140, d_out_141, q_in_141, d_out_142, q_in_142, d_out_143, qn_in_143, d_out_144, qn_in_144, d_out_145, q_in_145, d_out_146, q_in_146, d_out_147, q_in_147, d_out_148, q_in_148, d_out_149, q_in_149, d_out_150, q_in_150, d_out_151, q_in_151, d_out_152, q_in_152, d_out_153, q_in_153, d_out_154, q_in_154, d_out_155, q_in_155, d_out_156, q_in_156, d_out_157, q_in_157, d_out_158, q_in_158, d_out_159, q_in_159, d_out_160, q_in_160, d_out_161, q_in_161, d_out_162, q_in_162, d_out_163, q_in_163, d_out_164, q_in_164, d_out_165, q_in_165, d_out_166, q_in_166, d_out_167, q_in_167, d_out_168, q_in_168, d_out_169, q_in_169, d_out_170, q_in_170, d_out_171, q_in_171, d_out_172, q_in_172, d_out_173, q_in_173, d_out_174, q_in_174, d_out_175, q_in_175, d_out_176, q_in_176, d_out_177, q_in_177, d_out_178, q_in_178, d_out_179, q_in_179, d_out_180, q_in_180, d_out_181, q_in_181, d_out_182, qn_in_182, d_out_183, q_in_183, d_out_184, q_in_184, d_out_185, q_in_185, d_out_186, q_in_186, d_out_187, q_in_187, d_out_188, q_in_188, d_out_189, q_in_189, d_out_190, q_in_190, d_out_191, q_in_191, d_out_192, q_in_192, d_out_193, q_in_193, d_out_194, q_in_194, d_out_195, q_in_195, d_out_196, q_in_196, d_out_197, q_in_197, d_out_198, q_in_198, d_out_199, q_in_199, d_out_200, q_in_200, d_out_201, q_in_201, d_out_202, q_in_202, d_out_203, q_in_203, d_out_204, q_in_204, d_out_205, q_in_205, d_out_206, q_in_206, d_out_207, q_in_207, d_out_208, q_in_208, d_out_209, q_in_209, d_out_210, q_in_210, d_out_211, q_in_211, d_out_212, q_in_212, d_out_213, q_in_213, d_out_214, q_in_214, d_out_215, q_in_215, d_out_216, q_in_216, d_out_217, q_in_217, d_out_218, q_in_218, d_out_219, q_in_219, d_out_220, q_in_220, d_out_221, q_in_221, d_out_222, q_in_222, d_out_223, q_in_223, d_out_224, q_in_224, d_out_225, q_in_225, d_out_226, q_in_226, d_out_227, q_in_227, d_out_228, q_in_228, d_out_229, q_in_229, d_out_230, q_in_230, d_out_231, qn_in_231, d_out_232, q_in_232, d_out_233, qn_in_233, d_out_234, q_in_234, d_out_235, q_in_235, d_out_236, q_in_236, d_out_237, q_in_237, d_out_238, q_in_238, d_out_239, q_in_239, d_out_240, q_in_240, d_out_241, q_in_241, d_out_242, q_in_242, d_out_243, q_in_243, d_out_244, q_in_244, d_out_245, q_in_245, d_out_246, q_in_246, d_out_247, q_in_247, d_out_248, q_in_248, d_out_249, q_in_249, d_out_250, q_in_250, d_out_251, q_in_251, d_out_252, q_in_252, d_out_253, q_in_253, d_out_254, qn_in_254, d_out_255, q_in_255, d_out_256, q_in_256, d_out_257, q_in_257, d_out_258, q_in_258, d_out_259, q_in_259, d_out_260, q_in_260, d_out_261, q_in_261, d_out_262, q_in_262, d_out_263, q_in_263, d_out_264, q_in_264, d_out_265, q_in_265, d_out_266, q_in_266, d_out_267, q_in_267, d_out_268, q_in_268, d_out_269, q_in_269, d_out_270, q_in_270, d_out_271, q_in_271, d_out_272, q_in_272, d_out_273, qn_in_273, d_out_274, qn_in_274, d_out_275, qn_in_275, d_out_276, q_in_276, d_out_277, q_in_277, d_out_278, q_in_278, d_out_279, q_in_279, d_out_280, q_in_280, d_out_281, q_in_281, d_out_282, q_in_282, d_out_283, q_in_283, d_out_284, q_in_284, d_out_285, q_in_285, d_out_286, q_in_286, d_out_287, q_in_287, d_out_288, q_in_288, d_out_289, qn_in_289, d_out_290, q_in_290, d_out_291, q_in_291, d_out_292, q_in_292, d_out_293, q_in_293, d_out_294, q_in_294, d_out_295, q_in_295, d_out_296, q_in_296, d_out_297, q_in_297, d_out_298, q_in_298, d_out_299, q_in_299, d_out_300, q_in_300, d_out_301, q_in_301, d_out_302, q_in_302, d_out_303, q_in_303, d_out_304, q_in_304, d_out_305, q_in_305, d_out_306, q_in_306, d_out_307, q_in_307, d_out_308, q_in_308, d_out_309, q_in_309, d_out_310, q_in_310, d_out_311, q_in_311, d_out_312, q_in_312, d_out_313, q_in_313, d_out_314, q_in_314, d_out_315, q_in_315, d_out_316, q_in_316, d_out_317, q_in_317, d_out_318, q_in_318, d_out_319, q_in_319, d_out_320, q_in_320, d_out_321, q_in_321, d_out_322, q_in_322, d_out_323, q_in_323, d_out_324, q_in_324, d_out_325, q_in_325, d_out_326, q_in_326, d_out_327, q_in_327, d_out_328, q_in_328, d_out_329, q_in_329, d_out_330, q_in_330, d_out_331, q_in_331, d_out_332, q_in_332, d_out_333, q_in_333, d_out_334, q_in_334, d_out_335, q_in_335, d_out_336, q_in_336, d_out_337, q_in_337, d_out_338, q_in_338, d_out_339, q_in_339, d_out_340, q_in_340, d_out_341, q_in_341, d_out_342, q_in_342, d_out_343, q_in_343, d_out_344, q_in_344, d_out_345, q_in_345, d_out_346, q_in_346, d_out_347, q_in_347, d_out_348, q_in_348, d_out_349, q_in_349, d_out_350, q_in_350, d_out_351, q_in_351, d_out_352, q_in_352, d_out_353, q_in_353, d_out_354, q_in_354, d_out_355, q_in_355, d_out_356, q_in_356, d_out_357, q_in_357, d_out_358, q_in_358, d_out_359, q_in_359, d_out_360, q_in_360, d_out_361, q_in_361, d_out_362, q_in_362, d_out_363, q_in_363, d_out_364, q_in_364, d_out_365, q_in_365, d_out_366, q_in_366, d_out_367, q_in_367, d_out_368, q_in_368, d_out_369, q_in_369, d_out_370, q_in_370, d_out_371, q_in_371, d_out_372, q_in_372, d_out_373, q_in_373, d_out_374, q_in_374, d_out_375, q_in_375, d_out_376, q_in_376, d_out_377, q_in_377, d_out_378, q_in_378, d_out_379, q_in_379, d_out_380, q_in_380, d_out_381, q_in_381, d_out_382, q_in_382, d_out_383, q_in_383, d_out_384, q_in_384, d_out_385, q_in_385, d_out_386, q_in_386, d_out_387, q_in_387, d_out_388, q_in_388, d_out_389, q_in_389, d_out_390, q_in_390, d_out_391, q_in_391, d_out_392, q_in_392, d_out_393, q_in_393, d_out_394, q_in_394, d_out_395, q_in_395, d_out_396, q_in_396, d_out_397, q_in_397, d_out_398, q_in_398, d_out_399, q_in_399, d_out_400, q_in_400, d_out_401, q_in_401, d_out_402, q_in_402, d_out_403, q_in_403, d_out_404, q_in_404, d_out_405, q_in_405, d_out_406, q_in_406, d_out_407, q_in_407, d_out_408, q_in_408, d_out_409, q_in_409, d_out_410, q_in_410, d_out_411, q_in_411, d_out_412, q_in_412, d_out_413, q_in_413, d_out_414, q_in_414, d_out_415, q_in_415, d_out_416, q_in_416, d_out_417, q_in_417, d_out_418, q_in_418, d_out_419, q_in_419, d_out_420, q_in_420, d_out_421, q_in_421, d_out_422, q_in_422, d_out_423, q_in_423, d_out_424, q_in_424, d_out_425, q_in_425, d_out_426, q_in_426, d_out_427, q_in_427, d_out_428, q_in_428, d_out_429, q_in_429, d_out_430, q_in_430, d_out_431, q_in_431, d_out_432, q_in_432, d_out_433, q_in_433, d_out_434, q_in_434, d_out_435, q_in_435, d_out_436, q_in_436, d_out_437, q_in_437, d_out_438, q_in_438, d_out_439, q_in_439, d_out_440, q_in_440, d_out_441, q_in_441, d_out_442, q_in_442, d_out_443, q_in_443, d_out_444, q_in_444, d_out_445, q_in_445, d_out_446, q_in_446, d_out_447, q_in_447, d_out_448, q_in_448, d_out_449, q_in_449, d_out_450, q_in_450, d_out_451, q_in_451, d_out_452, q_in_452, d_out_453, q_in_453, d_out_454, q_in_454, d_out_455, q_in_455, d_out_456, q_in_456, d_out_457, q_in_457, d_out_458, q_in_458, d_out_459, q_in_459, d_out_460, q_in_460, d_out_461, q_in_461, d_out_462, q_in_462, d_out_463, q_in_463, d_out_464, q_in_464, d_out_465, q_in_465, d_out_466, q_in_466, d_out_467, q_in_467, d_out_468, q_in_468, d_out_469, q_in_469, d_out_470, q_in_470, d_out_471, q_in_471, d_out_472, q_in_472, d_out_473, q_in_473, d_out_474, q_in_474, d_out_475, qn_in_475, d_out_476, qn_in_476, d_out_477, q_in_477, d_out_478, qn_in_478, d_out_479, qn_in_479, d_out_480, q_in_480, d_out_481, q_in_481, d_out_482, q_in_482, d_out_483, q_in_483, d_out_484, q_in_484, d_out_485, q_in_485, d_out_486, q_in_486, d_out_487, q_in_487, d_out_488, q_in_488, d_out_489, q_in_489, d_out_490, q_in_490, d_out_491, q_in_491, d_out_492, q_in_492, d_out_493, q_in_493, d_out_494, q_in_494, d_out_495, q_in_495, d_out_496, q_in_496, d_out_497, qn_in_497, d_out_498, q_in_498, d_out_499, qn_in_499, d_out_500, q_in_500, d_out_501, q_in_501, d_out_502, qn_in_502, d_out_503, q_in_503, d_out_504, q_in_504, d_out_505, q_in_505, d_out_506, q_in_506, d_out_507, q_in_507, d_out_508, q_in_508, d_out_509, q_in_509, d_out_510, q_in_510, d_out_511, q_in_511, d_out_512, q_in_512, d_out_513, q_in_513, d_out_514, q_in_514, d_out_515, q_in_515, d_out_516, q_in_516, d_out_517, q_in_517, d_out_518, q_in_518, d_out_519, q_in_519, d_out_520, q_in_520, d_out_521, q_in_521, d_out_522, q_in_522, d_out_523, q_in_523, d_out_524, q_in_524, d_out_525, q_in_525, d_out_526, q_in_526, d_out_527, q_in_527, d_out_528, q_in_528, d_out_529, q_in_529, d_out_530, q_in_530, d_out_531, q_in_531, d_out_532, q_in_532, d_out_533, q_in_533, d_out_534, q_in_534, d_out_535, q_in_535, d_out_536, q_in_536, d_out_537, q_in_537, d_out_538, q_in_538, d_out_539, q_in_539, d_out_540, q_in_540, d_out_541, q_in_541, d_out_542, q_in_542, d_out_543, qn_in_543, d_out_544, q_in_544, d_out_545, q_in_545, d_out_546, q_in_546, d_out_547, q_in_547, d_out_548, q_in_548, d_out_549, q_in_549, d_out_550, q_in_550, d_out_551, q_in_551, d_out_552, q_in_552, d_out_553, q_in_553, d_out_554, q_in_554, d_out_555, q_in_555, d_out_556, q_in_556, d_out_557, q_in_557, d_out_558, q_in_558, d_out_559, q_in_559, d_out_560, q_in_560, d_out_561, q_in_561, d_out_562, q_in_562, d_out_563, q_in_563, d_out_564, q_in_564, d_out_565, q_in_565, d_out_566, q_in_566, d_out_567, q_in_567, d_out_568, q_in_568, d_out_569, q_in_569, d_out_570, q_in_570, d_out_571, q_in_571, d_out_572, q_in_572, d_out_573, q_in_573, d_out_574, q_in_574, d_out_575, q_in_575, d_out_576, q_in_576, d_out_577, q_in_577, d_out_578, q_in_578, d_out_579, q_in_579, d_out_580, q_in_580, d_out_581, q_in_581, d_out_582, q_in_582, d_out_583, q_in_583, d_out_584, q_in_584, d_out_585, q_in_585, d_out_586, q_in_586, d_out_587, q_in_587, d_out_588, q_in_588, d_out_589, q_in_589, d_out_590, q_in_590, d_out_591, q_in_591, d_out_592, q_in_592, d_out_593, q_in_593, d_out_594, q_in_594, d_out_595, q_in_595, d_out_596, q_in_596, d_out_597, q_in_597, d_out_598, q_in_598, d_out_599, q_in_599, d_out_600, q_in_600, d_out_601, q_in_601, d_out_602, q_in_602, d_out_603, q_in_603, d_out_604, q_in_604, d_out_605, q_in_605, d_out_606, q_in_606, d_out_607, q_in_607, d_out_608, q_in_608, d_out_609, q_in_609, d_out_610, q_in_610, d_out_611, q_in_611, d_out_612, q_in_612, d_out_613, q_in_613, d_out_614, q_in_614, d_out_615, q_in_615, d_out_616, q_in_616, d_out_617, q_in_617, d_out_618, q_in_618, d_out_619, q_in_619, d_out_620, q_in_620, d_out_621, q_in_621, d_out_622, q_in_622, d_out_623, q_in_623, d_out_624, q_in_624, d_out_625, q_in_625, d_out_626, q_in_626, d_out_627, q_in_627, d_out_628, q_in_628, d_out_629, q_in_629, d_out_630, q_in_630, d_out_631, q_in_631, d_out_632, q_in_632, d_out_633, q_in_633, d_out_634, q_in_634, d_out_635, q_in_635, d_out_636, q_in_636, d_out_637, q_in_637, d_out_638, q_in_638, d_out_639, q_in_639, d_out_640, q_in_640, d_out_641, q_in_641, d_out_642, q_in_642, d_out_643, q_in_643, d_out_644, q_in_644, d_out_645, q_in_645, d_out_646, q_in_646, d_out_647, q_in_647, d_out_648, q_in_648, d_out_649, q_in_649, d_out_650, q_in_650, d_out_651, q_in_651, d_out_652, q_in_652, d_out_653, q_in_653, d_out_654, q_in_654, d_out_655, q_in_655, d_out_656, q_in_656, d_out_657, q_in_657, d_out_658, q_in_658, d_out_659, q_in_659, d_out_660, q_in_660, d_out_661, q_in_661, d_out_662, q_in_662, d_out_663, q_in_663, d_out_664, q_in_664, d_out_665, q_in_665, d_out_666, q_in_666, d_out_667, q_in_667, d_out_668, q_in_668, d_out_669, q_in_669, d_out_670, q_in_670, d_out_671, q_in_671, d_out_672, q_in_672, d_out_673, q_in_673, d_out_674, q_in_674, d_out_675, q_in_675, d_out_676, q_in_676, d_out_677, q_in_677, d_out_678, q_in_678, d_out_679, q_in_679, d_out_680, q_in_680, d_out_681, q_in_681, d_out_682, q_in_682, d_out_683, q_in_683, d_out_684, q_in_684, d_out_685, q_in_685, d_out_686, q_in_686, d_out_687, q_in_687, d_out_688, q_in_688, d_out_689, q_in_689, d_out_690, q_in_690, d_out_691, q_in_691, d_out_692, q_in_692, d_out_693, q_in_693, d_out_694, q_in_694, d_out_695, q_in_695, d_out_696, q_in_696, d_out_697, q_in_697, d_out_698, qn_in_698, d_out_699, qn_in_699, d_out_700, qn_in_700, d_out_701, qn_in_701, d_out_702, qn_in_702, d_out_703, qn_in_703);
input q_in_405;
input q_in_217;
input q_in_664;
input q_in_404;
input q_in_403;
input q_in_402;
input q_in_401;
input q_in_400;
input q_in_399;
input q_in_398;
input q_in_397;
input q_in_663;
input q_in_216;
input q_in_215;
input q_in_214;
input q_in_213;
input q_in_212;
input q_in_211;
input q_in_210;
input q_in_209;
input q_in_208;
input q_in_207;
input q_in_206;
input q_in_205;
input q_in_204;
input q_in_203;
input q_in_202;
input q_in_201;
input q_in_200;
input q_in_199;
input q_in_198;
input q_in_197;
input q_in_196;
input q_in_195;
input q_in_194;
input q_in_690;
input q_in_696;
input q_in_396;
input q_in_193;
input q_in_192;
input q_in_191;
input q_in_190;
input q_in_189;
input q_in_188;
input q_in_187;
input q_in_186;
input q_in_185;
input q_in_184;
input q_in_183;
input qn_in_182;
input q_in_181;
input q_in_180;
input q_in_179;
input q_in_178;
input q_in_177;
input q_in_176;
input q_in_175;
input q_in_174;
input q_in_173;
input q_in_172;
input q_in_171;
input q_in_170;
input q_in_169;
input q_in_168;
input q_in_688;
input q_in_695;
input q_in_694;
input q_in_693;
input q_in_351;
input q_in_350;
input q_in_349;
input q_in_348;
input q_in_347;
input q_in_167;
input q_in_166;
input q_in_165;
input q_in_164;
input q_in_163;
input q_in_162;
input q_in_161;
input q_in_160;
input q_in_159;
input q_in_158;
input q_in_157;
input q_in_156;
input q_in_155;
input q_in_154;
input q_in_153;
input q_in_152;
input q_in_151;
input q_in_150;
input q_in_149;
input q_in_148;
input q_in_147;
input q_in_146;
input q_in_145;
input qn_in_144;
input qn_in_143;
input qn_in_702;
input q_in_394;
input q_in_393;
input q_in_392;
input q_in_391;
input q_in_390;
input q_in_142;
input q_in_141;
input q_in_140;
input qn_in_139;
input q_in_138;
input q_in_137;
input q_in_136;
input q_in_135;
input q_in_134;
input q_in_133;
input q_in_132;
input q_in_131;
input q_in_130;
input q_in_129;
input q_in_128;
input q_in_127;
input q_in_126;
input q_in_125;
input q_in_124;
input q_in_123;
input q_in_122;
input q_in_121;
input q_in_120;
input q_in_119;
input q_in_118;
input q_in_117;
input q_in_116;
input q_in_115;
input q_in_114;
input q_in_113;
input qn_in_112;
input q_in_687;
input q_in_686;
input q_in_364;
input q_in_561;
input q_in_560;
input q_in_111;
input q_in_110;
input q_in_109;
input q_in_108;
input q_in_107;
input q_in_106;
input q_in_105;
input q_in_104;
input q_in_103;
input q_in_102;
input q_in_101;
input q_in_100;
input q_in_99;
input q_in_98;
input q_in_97;
input q_in_96;
input q_in_95;
input q_in_94;
input q_in_93;
input q_in_92;
input q_in_91;
input q_in_90;
input q_in_89;
input qn_in_88;
input q_in_87;
input qn_in_86;
input qn_in_85;
input qn_in_84;
input q_in_83;
input qn_in_703;
input q_in_554;
input q_in_685;
input q_in_684;
input q_in_683;
input q_in_682;
input q_in_681;
input q_in_680;
input q_in_679;
input q_in_678;
input q_in_677;
input q_in_676;
input q_in_675;
input q_in_674;
input q_in_673;
input q_in_672;
input q_in_671;
input q_in_670;
input q_in_669;
input q_in_82;
input q_in_81;
input q_in_80;
input q_in_79;
input q_in_78;
input q_in_77;
input q_in_76;
input q_in_75;
input q_in_74;
input q_in_73;
input q_in_72;
input q_in_71;
input q_in_70;
input q_in_69;
input q_in_68;
input q_in_67;
input q_in_66;
input q_in_65;
input q_in_64;
input q_in_63;
input q_in_661;
input q_in_660;
input q_in_659;
input q_in_62;
input qn_in_61;
input q_in_60;
input q_in_59;
input q_in_58;
input q_in_57;
input q_in_56;
input q_in_55;
input q_in_54;
input q_in_53;
input q_in_52;
input qn_in_51;
input qn_in_50;
input qn_in_49;
input qn_in_48;
input qn_in_47;
input qn_in_46;
input q_in_45;
input q_in_44;
input q_in_668;
input q_in_658;
input q_in_667;
input qn_in_43;
input q_in_42;
input q_in_41;
input q_in_40;
input q_in_39;
input qn_in_38;
input qn_in_37;
input qn_in_36;
input qn_in_35;
input q_in_34;
input q_in_33;
input qn_in_32;
input q_in_31;
input q_in_341;
input q_in_340;
input q_in_30;
input q_in_29;
input q_in_28;
input q_in_27;
input qn_in_26;
input qn_in_25;
input qn_in_24;
input qn_in_23;
input q_in_22;
input qn_in_21;
input q_in_20;
input q_in_19;
input q_in_18;
input q_in_653;
input q_in_652;
input q_in_651;
input q_in_650;
input qn_in_17;
input q_in_16;
input q_in_15;
input q_in_14;
input q_in_13;
input q_in_12;
input q_in_643;
input q_in_642;
input q_in_11;
input q_in_10;
input q_in_9;
input qn_in_8;
input qn_in_7;
input q_in_6;
input q_in_5;
input q_in_4;
input q_in_3;
input qn_in_2;
input qn_in_1;
input q_in_630;
input q_in_629;
input q_in_628;
input q_in_627;
input q_in_626;
input q_in_625;
input q_in_389;
input q_in_624;
input q_in_623;
input q_in_662;
input q_in_388;
input q_in_387;
input q_in_386;
input q_in_385;
input q_in_384;
input q_in_383;
input q_in_636;
input q_in_622;
input q_in_621;
input q_in_620;
input q_in_619;
input q_in_618;
input q_in_617;
input q_in_616;
input q_in_615;
input q_in_614;
input q_in_613;
input q_in_612;
input q_in_611;
input q_in_610;
input q_in_609;
input q_in_608;
input q_in_607;
input q_in_606;
input q_in_605;
input q_in_604;
input q_in_603;
input q_in_602;
input q_in_601;
input q_in_600;
input q_in_599;
input q_in_598;
input q_in_597;
input q_in_596;
input q_in_595;
input q_in_594;
input q_in_593;
input q_in_592;
input q_in_591;
input q_in_590;
input q_in_589;
input q_in_588;
input q_in_431;
input q_in_587;
input q_in_586;
input q_in_585;
input q_in_584;
input q_in_583;
input q_in_582;
input q_in_581;
input q_in_580;
input q_in_579;
input q_in_578;
input q_in_577;
input q_in_576;
input q_in_575;
input q_in_574;
input q_in_573;
input q_in_572;
input q_in_571;
input q_in_570;
input q_in_569;
input q_in_568;
input q_in_567;
input q_in_566;
input q_in_565;
input q_in_564;
input q_in_563;
input q_in_562;
input q_in_339;
input q_in_338;
input q_in_337;
input q_in_336;
input q_in_335;
input q_in_334;
input q_in_333;
input q_in_332;
input qn_in_701;
input q_in_553;
input q_in_552;
input q_in_461;
input q_in_551;
input q_in_331;
input q_in_550;
input q_in_549;
input q_in_548;
input q_in_547;
input q_in_546;
input q_in_545;
input q_in_544;
input q_in_697;
input qn_in_543;
input q_in_542;
input q_in_541;
input q_in_540;
input q_in_539;
input q_in_382;
input q_in_538;
input q_in_537;
input q_in_536;
input q_in_535;
input q_in_534;
input q_in_533;
input q_in_532;
input q_in_531;
input q_in_441;
input q_in_529;
input q_in_528;
input q_in_343;
input q_in_527;
input q_in_342;
input q_in_330;
input q_in_380;
input q_in_526;
input q_in_525;
input q_in_524;
input q_in_523;
input q_in_522;
input q_in_521;
input q_in_520;
input q_in_519;
input q_in_329;
input q_in_328;
input q_in_327;
input q_in_326;
input q_in_325;
input q_in_324;
input q_in_323;
input q_in_322;
input q_in_321;
input q_in_510;
input q_in_509;
input q_in_508;
input q_in_507;
input q_in_506;
input q_in_505;
input q_in_504;
input q_in_503;
input qn_in_502;
input q_in_501;
input q_in_500;
input q_in_657;
input q_in_656;
input q_in_655;
input q_in_654;
input q_in_378;
input q_in_518;
input q_in_498;
input qn_in_497;
input q_in_320;
input q_in_517;
input q_in_649;
input q_in_474;
input q_in_648;
input q_in_647;
input q_in_646;
input q_in_645;
input q_in_516;
input q_in_644;
input q_in_641;
input q_in_640;
input q_in_515;
input q_in_639;
input q_in_363;
input q_in_638;
input q_in_637;
input q_in_473;
input q_in_472;
input q_in_471;
input q_in_470;
input q_in_469;
input q_in_468;
input q_in_467;
input q_in_466;
input q_in_635;
input q_in_514;
input q_in_634;
input q_in_496;
input q_in_495;
input q_in_494;
input q_in_493;
input q_in_492;
input q_in_491;
input q_in_319;
input q_in_318;
input q_in_317;
input q_in_316;
input q_in_315;
input q_in_314;
input q_in_313;
input q_in_483;
input q_in_482;
input q_in_631;
input q_in_481;
input q_in_558;
input q_in_464;
input q_in_463;
input q_in_462;
input q_in_465;
input q_in_377;
input q_in_376;
input q_in_489;
input q_in_557;
input q_in_460;
input q_in_488;
input q_in_459;
input q_in_458;
input q_in_487;
input q_in_457;
input q_in_486;
input q_in_485;
input q_in_484;
input q_in_556;
input q_in_312;
input q_in_555;
input qn_in_700;
input q_in_346;
input q_in_456;
input q_in_530;
input q_in_345;
input q_in_311;
input q_in_310;
input q_in_309;
input q_in_308;
input q_in_307;
input q_in_455;
input q_in_454;
input q_in_453;
input q_in_452;
input q_in_451;
input q_in_450;
input q_in_449;
input q_in_448;
input q_in_447;
input q_in_446;
input q_in_445;
input q_in_444;
input q_in_443;
input q_in_442;
input q_in_306;
input q_in_440;
input q_in_439;
input q_in_438;
input q_in_437;
input q_in_436;
input q_in_435;
input q_in_434;
input q_in_433;
input q_in_432;
input q_in_480;
input q_in_305;
input q_in_395;
input q_in_633;
input q_in_344;
input q_in_632;
input q_in_304;
input q_in_430;
input q_in_429;
input q_in_428;
input q_in_427;
input q_in_426;
input q_in_303;
input q_in_302;
input q_in_301;
input q_in_300;
input q_in_299;
input q_in_298;
input q_in_297;
input q_in_296;
input q_in_295;
input q_in_294;
input q_in_293;
input q_in_292;
input q_in_291;
input q_in_425;
input q_in_424;
input q_in_423;
input q_in_422;
input q_in_421;
input qn_in_479;
input q_in_290;
input qn_in_478;
input q_in_477;
input qn_in_476;
input qn_in_475;
input q_in_375;
input q_in_374;
input q_in_420;
input qn_in_289;
input q_in_288;
input q_in_287;
input q_in_286;
input q_in_285;
input q_in_284;
input q_in_283;
input q_in_282;
input q_in_281;
input q_in_280;
input q_in_362;
input q_in_361;
input q_in_360;
input q_in_359;
input q_in_358;
input q_in_419;
input q_in_279;
input q_in_417;
input q_in_490;
input q_in_416;
input q_in_415;
input q_in_414;
input q_in_413;
input q_in_357;
input qn_in_699;
input q_in_379;
input q_in_373;
input q_in_418;
input q_in_356;
input q_in_355;
input q_in_354;
input qn_in_499;
input q_in_278;
input q_in_692;
input q_in_691;
input q_in_277;
input q_in_276;
input qn_in_275;
input qn_in_274;
input qn_in_273;
input q_in_272;
input q_in_271;
input q_in_270;
input q_in_269;
input q_in_268;
input q_in_267;
input q_in_266;
input q_in_689;
input q_in_412;
input q_in_411;
input q_in_265;
input q_in_410;
input q_in_409;
input q_in_408;
input q_in_407;
input q_in_264;
input q_in_666;
input qn_in_698;
input q_in_665;
input q_in_263;
input q_in_262;
input q_in_261;
input q_in_260;
input q_in_259;
input q_in_258;
input q_in_257;
input q_in_256;
input q_in_255;
input qn_in_254;
input q_in_253;
input q_in_252;
input q_in_251;
input q_in_250;
input q_in_249;
input q_in_248;
input q_in_366;
input q_in_365;
input q_in_247;
input q_in_372;
input q_in_371;
input q_in_370;
input q_in_369;
input q_in_368;
input q_in_381;
input q_in_559;
input q_in_246;
input q_in_245;
input q_in_244;
input q_in_243;
input q_in_242;
input q_in_241;
input q_in_240;
input q_in_239;
input q_in_238;
input q_in_237;
input q_in_236;
input q_in_235;
input q_in_234;
input qn_in_233;
input q_in_232;
input qn_in_231;
input q_in_230;
input q_in_229;
input q_in_228;
input q_in_227;
input q_in_226;
input q_in_225;
input q_in_224;
input q_in_223;
input q_in_222;
input q_in_221;
input q_in_220;
input q_in_513;
input q_in_219;
input q_in_512;
input q_in_353;
input q_in_511;
input q_in_406;
input q_in_218;
input q_in_352;
input q_in_367;
input [31:0] si;
input clock, reset;
output d_out_405;
output d_out_217;
output d_out_664;
output d_out_404;
output d_out_403;
output d_out_402;
output d_out_401;
output d_out_400;
output d_out_399;
output d_out_398;
output d_out_397;
output d_out_663;
output d_out_216;
output d_out_215;
output d_out_214;
output d_out_213;
output d_out_212;
output d_out_211;
output d_out_210;
output d_out_209;
output d_out_208;
output d_out_207;
output d_out_206;
output d_out_205;
output d_out_204;
output d_out_203;
output d_out_202;
output d_out_201;
output d_out_200;
output d_out_199;
output d_out_198;
output d_out_197;
output d_out_196;
output d_out_195;
output d_out_194;
output d_out_690;
output d_out_696;
output d_out_396;
output d_out_193;
output d_out_192;
output d_out_191;
output d_out_190;
output d_out_189;
output d_out_188;
output d_out_187;
output d_out_186;
output d_out_185;
output d_out_184;
output d_out_183;
output d_out_182;
output d_out_181;
output d_out_180;
output d_out_179;
output d_out_178;
output d_out_177;
output d_out_176;
output d_out_175;
output d_out_174;
output d_out_173;
output d_out_172;
output d_out_171;
output d_out_170;
output d_out_169;
output d_out_168;
output d_out_688;
output d_out_695;
output d_out_694;
output d_out_693;
output d_out_351;
output d_out_350;
output d_out_349;
output d_out_348;
output d_out_347;
output d_out_167;
output d_out_166;
output d_out_165;
output d_out_164;
output d_out_163;
output d_out_162;
output d_out_161;
output d_out_160;
output d_out_159;
output d_out_158;
output d_out_157;
output d_out_156;
output d_out_155;
output d_out_154;
output d_out_153;
output d_out_152;
output d_out_151;
output d_out_150;
output d_out_149;
output d_out_148;
output d_out_147;
output d_out_146;
output d_out_145;
output d_out_144;
output d_out_143;
output d_out_702;
output d_out_394;
output d_out_393;
output d_out_392;
output d_out_391;
output d_out_390;
output d_out_142;
output d_out_141;
output d_out_140;
output d_out_139;
output d_out_138;
output d_out_137;
output d_out_136;
output d_out_135;
output d_out_134;
output d_out_133;
output d_out_132;
output d_out_131;
output d_out_130;
output d_out_129;
output d_out_128;
output d_out_127;
output d_out_126;
output d_out_125;
output d_out_124;
output d_out_123;
output d_out_122;
output d_out_121;
output d_out_120;
output d_out_119;
output d_out_118;
output d_out_117;
output d_out_116;
output d_out_115;
output d_out_114;
output d_out_113;
output d_out_112;
output d_out_687;
output d_out_686;
output d_out_364;
output d_out_561;
output d_out_560;
output d_out_111;
output d_out_110;
output d_out_109;
output d_out_108;
output d_out_107;
output d_out_106;
output d_out_105;
output d_out_104;
output d_out_103;
output d_out_102;
output d_out_101;
output d_out_100;
output d_out_99;
output d_out_98;
output d_out_97;
output d_out_96;
output d_out_95;
output d_out_94;
output d_out_93;
output d_out_92;
output d_out_91;
output d_out_90;
output d_out_89;
output d_out_88;
output d_out_87;
output d_out_86;
output d_out_85;
output d_out_84;
output d_out_83;
output d_out_703;
output d_out_554;
output d_out_685;
output d_out_684;
output d_out_683;
output d_out_682;
output d_out_681;
output d_out_680;
output d_out_679;
output d_out_678;
output d_out_677;
output d_out_676;
output d_out_675;
output d_out_674;
output d_out_673;
output d_out_672;
output d_out_671;
output d_out_670;
output d_out_669;
output d_out_82;
output d_out_81;
output d_out_80;
output d_out_79;
output d_out_78;
output d_out_77;
output d_out_76;
output d_out_75;
output d_out_74;
output d_out_73;
output d_out_72;
output d_out_71;
output d_out_70;
output d_out_69;
output d_out_68;
output d_out_67;
output d_out_66;
output d_out_65;
output d_out_64;
output d_out_63;
output d_out_661;
output d_out_660;
output d_out_659;
output d_out_62;
output d_out_61;
output d_out_60;
output d_out_59;
output d_out_58;
output d_out_57;
output d_out_56;
output d_out_55;
output d_out_54;
output d_out_53;
output d_out_52;
output d_out_51;
output d_out_50;
output d_out_49;
output d_out_48;
output d_out_47;
output d_out_46;
output d_out_45;
output d_out_44;
output d_out_668;
output d_out_658;
output d_out_667;
output d_out_43;
output d_out_42;
output d_out_41;
output d_out_40;
output d_out_39;
output d_out_38;
output d_out_37;
output d_out_36;
output d_out_35;
output d_out_34;
output d_out_33;
output d_out_32;
output d_out_31;
output d_out_341;
output d_out_340;
output d_out_30;
output d_out_29;
output d_out_28;
output d_out_27;
output d_out_26;
output d_out_25;
output d_out_24;
output d_out_23;
output d_out_22;
output d_out_21;
output d_out_20;
output d_out_19;
output d_out_18;
output d_out_653;
output d_out_652;
output d_out_651;
output d_out_650;
output d_out_17;
output d_out_16;
output d_out_15;
output d_out_14;
output d_out_13;
output d_out_12;
output d_out_643;
output d_out_642;
output d_out_11;
output d_out_10;
output d_out_9;
output d_out_8;
output d_out_7;
output d_out_6;
output d_out_5;
output d_out_4;
output d_out_3;
output d_out_2;
output d_out_1;
output d_out_630;
output d_out_629;
output d_out_628;
output d_out_627;
output d_out_626;
output d_out_511;
output d_out_625;
output d_out_389;
output d_out_624;
output d_out_623;
output d_out_662;
output d_out_388;
output d_out_387;
output d_out_386;
output d_out_385;
output d_out_384;
output d_out_383;
output d_out_636;
output d_out_622;
output d_out_621;
output d_out_620;
output d_out_619;
output d_out_618;
output d_out_617;
output d_out_616;
output d_out_615;
output d_out_614;
output d_out_613;
output d_out_612;
output d_out_611;
output d_out_610;
output d_out_609;
output d_out_608;
output d_out_607;
output d_out_606;
output d_out_605;
output d_out_604;
output d_out_603;
output d_out_602;
output d_out_601;
output d_out_600;
output d_out_599;
output d_out_598;
output d_out_597;
output d_out_596;
output d_out_595;
output d_out_594;
output d_out_593;
output d_out_592;
output d_out_591;
output d_out_590;
output d_out_589;
output d_out_588;
output d_out_431;
output d_out_587;
output d_out_586;
output d_out_585;
output d_out_584;
output d_out_583;
output d_out_582;
output d_out_581;
output d_out_580;
output d_out_579;
output d_out_578;
output d_out_577;
output d_out_576;
output d_out_575;
output d_out_574;
output d_out_573;
output d_out_572;
output d_out_571;
output d_out_570;
output d_out_569;
output d_out_568;
output d_out_567;
output d_out_566;
output d_out_565;
output d_out_564;
output d_out_563;
output d_out_562;
output d_out_339;
output d_out_338;
output d_out_337;
output d_out_336;
output d_out_335;
output d_out_334;
output d_out_333;
output d_out_332;
output d_out_701;
output d_out_553;
output d_out_552;
output d_out_461;
output d_out_551;
output d_out_331;
output d_out_550;
output d_out_549;
output d_out_548;
output d_out_547;
output d_out_546;
output d_out_545;
output d_out_544;
output d_out_697;
output d_out_543;
output d_out_542;
output d_out_541;
output d_out_540;
output d_out_539;
output d_out_382;
output d_out_538;
output d_out_537;
output d_out_536;
output d_out_535;
output d_out_534;
output d_out_533;
output d_out_532;
output d_out_531;
output d_out_441;
output d_out_529;
output d_out_528;
output d_out_343;
output d_out_527;
output d_out_342;
output d_out_330;
output d_out_380;
output d_out_526;
output d_out_525;
output d_out_524;
output d_out_523;
output d_out_522;
output d_out_521;
output d_out_520;
output d_out_519;
output d_out_329;
output d_out_328;
output d_out_327;
output d_out_326;
output d_out_325;
output d_out_324;
output d_out_323;
output d_out_322;
output d_out_321;
output d_out_510;
output d_out_509;
output d_out_508;
output d_out_507;
output d_out_506;
output d_out_505;
output d_out_504;
output d_out_503;
output d_out_502;
output d_out_501;
output d_out_500;
output d_out_657;
output d_out_656;
output d_out_655;
output d_out_654;
output d_out_378;
output d_out_518;
output d_out_498;
output d_out_497;
output d_out_320;
output d_out_517;
output d_out_649;
output d_out_474;
output d_out_648;
output d_out_647;
output d_out_646;
output d_out_645;
output d_out_516;
output d_out_644;
output d_out_641;
output d_out_640;
output d_out_515;
output d_out_639;
output d_out_363;
output d_out_638;
output d_out_637;
output d_out_473;
output d_out_472;
output d_out_471;
output d_out_470;
output d_out_469;
output d_out_468;
output d_out_467;
output d_out_466;
output d_out_635;
output d_out_514;
output d_out_634;
output d_out_496;
output d_out_495;
output d_out_494;
output d_out_493;
output d_out_492;
output d_out_491;
output d_out_319;
output d_out_318;
output d_out_317;
output d_out_316;
output d_out_315;
output d_out_314;
output d_out_313;
output d_out_483;
output d_out_482;
output d_out_631;
output d_out_481;
output d_out_558;
output d_out_464;
output d_out_463;
output d_out_462;
output d_out_465;
output d_out_377;
output d_out_376;
output d_out_489;
output d_out_557;
output d_out_460;
output d_out_488;
output d_out_459;
output d_out_458;
output d_out_487;
output d_out_457;
output d_out_486;
output d_out_485;
output d_out_484;
output d_out_556;
output d_out_312;
output d_out_555;
output d_out_700;
output d_out_346;
output d_out_456;
output d_out_530;
output d_out_345;
output d_out_311;
output d_out_310;
output d_out_309;
output d_out_308;
output d_out_307;
output d_out_455;
output d_out_454;
output d_out_453;
output d_out_452;
output d_out_451;
output d_out_450;
output d_out_449;
output d_out_448;
output d_out_447;
output d_out_446;
output d_out_445;
output d_out_444;
output d_out_443;
output d_out_442;
output d_out_306;
output d_out_440;
output d_out_439;
output d_out_438;
output d_out_437;
output d_out_436;
output d_out_435;
output d_out_434;
output d_out_433;
output d_out_432;
output d_out_480;
output d_out_305;
output d_out_395;
output d_out_633;
output d_out_344;
output d_out_632;
output d_out_304;
output d_out_430;
output d_out_429;
output d_out_428;
output d_out_427;
output d_out_426;
output d_out_303;
output d_out_302;
output d_out_301;
output d_out_300;
output d_out_299;
output d_out_298;
output d_out_297;
output d_out_296;
output d_out_295;
output d_out_294;
output d_out_293;
output d_out_292;
output d_out_291;
output d_out_425;
output d_out_424;
output d_out_423;
output d_out_422;
output d_out_421;
output d_out_479;
output d_out_290;
output d_out_478;
output d_out_477;
output d_out_476;
output d_out_475;
output d_out_375;
output d_out_374;
output d_out_420;
output d_out_289;
output d_out_288;
output d_out_287;
output d_out_286;
output d_out_285;
output d_out_284;
output d_out_283;
output d_out_282;
output d_out_281;
output d_out_280;
output d_out_362;
output d_out_361;
output d_out_360;
output d_out_359;
output d_out_358;
output d_out_419;
output d_out_279;
output d_out_417;
output d_out_490;
output d_out_416;
output d_out_415;
output d_out_414;
output d_out_413;
output d_out_357;
output d_out_699;
output d_out_379;
output d_out_373;
output d_out_418;
output d_out_356;
output d_out_355;
output d_out_354;
output d_out_499;
output d_out_278;
output d_out_692;
output d_out_691;
output d_out_277;
output d_out_276;
output d_out_275;
output d_out_274;
output d_out_273;
output d_out_272;
output d_out_271;
output d_out_270;
output d_out_269;
output d_out_268;
output d_out_267;
output d_out_266;
output d_out_689;
output d_out_412;
output d_out_411;
output d_out_265;
output d_out_410;
output d_out_409;
output d_out_408;
output d_out_407;
output d_out_264;
output d_out_666;
output d_out_698;
output d_out_665;
output d_out_263;
output d_out_262;
output d_out_261;
output d_out_260;
output d_out_259;
output d_out_258;
output d_out_257;
output d_out_256;
output d_out_255;
output d_out_254;
output d_out_253;
output d_out_252;
output d_out_251;
output d_out_250;
output d_out_249;
output d_out_248;
output d_out_366;
output d_out_365;
output d_out_247;
output d_out_372;
output d_out_371;
output d_out_370;
output d_out_369;
output d_out_368;
output d_out_381;
output d_out_559;
output d_out_246;
output d_out_245;
output d_out_244;
output d_out_243;
output d_out_242;
output d_out_241;
output d_out_240;
output d_out_239;
output d_out_238;
output d_out_237;
output d_out_236;
output d_out_235;
output d_out_234;
output d_out_233;
output d_out_232;
output d_out_231;
output d_out_230;
output d_out_229;
output d_out_228;
output d_out_227;
output d_out_226;
output d_out_225;
output d_out_224;
output d_out_223;
output d_out_222;
output d_out_221;
output d_out_220;
output d_out_513;
output d_out_219;
output d_out_512;
output d_out_353;
output d_out_367;
output d_out_218;
output d_out_352;
output rd, wr;
output [19:0] so;
output d_out_406;
wire wr_3;
wire n_35950, n_35951, n_35952, rd_1, rd_2, rd_3, wr_1, wr_2;
wire n_35941, n_35942, n_35943, n_35944, n_35945, n_35946, n_35947, n_35949;
wire n_35933, n_35934, n_35935, n_35936, n_35937, n_35938, n_35939, n_35940;
wire n_35925, n_35926, n_35927, n_35928, n_35929, n_35930, n_35931, n_35932;
wire n_35917, n_35918, n_35919, n_35920, n_35921, n_35922, n_35923, n_35924;
wire n_35906, n_35907, n_35908, n_35909, n_35912, n_35913, n_35914, n_35915;
wire n_35898, n_35899, n_35900, n_35901, n_35902, n_35903, n_35904, n_35905;
wire n_35884, n_35885, n_35886, n_35889, n_35890, n_35895, n_35896, n_35897;
wire n_35876, n_35877, n_35878, n_35879, n_35880, n_35881, n_35882, n_35883;
wire n_35868, n_35869, n_35870, n_35871, n_35872, n_35873, n_35874, n_35875;
wire n_35849, n_35850, n_35860, n_35861, n_35863, n_35864, n_35865, n_35867;
wire n_35822, n_35824, n_35829, n_35830, n_35834, n_35840, n_35842, n_35844;
wire n_35771, n_35775, n_35776, n_35790, n_35794, n_35813, n_35816, n_35818;
wire n_35718, n_35719, n_35736, n_35744, n_35761, n_35766, n_35767, n_35768;
wire n_35710, n_35711, n_35712, n_35713, n_35714, n_35715, n_35716, n_35717;
wire n_35702, n_35703, n_35704, n_35705, n_35706, n_35707, n_35708, n_35709;
wire n_35693, n_35694, n_35695, n_35696, n_35697, n_35698, n_35699, n_35700;
wire n_35675, n_35679, n_35686, n_35688, n_35689, n_35690, n_35691, n_35692;
wire n_35666, n_35667, n_35668, n_35669, n_35670, n_35671, n_35672, n_35674;
wire n_35657, n_35658, n_35659, n_35660, n_35661, n_35662, n_35663, n_35665;
wire n_35648, n_35649, n_35650, n_35651, n_35652, n_35653, n_35655, n_35656;
wire n_35638, n_35639, n_35640, n_35641, n_35644, n_35645, n_35646, n_35647;
wire n_35630, n_35631, n_35632, n_35633, n_35634, n_35635, n_35636, n_35637;
wire n_35621, n_35622, n_35623, n_35624, n_35625, n_35626, n_35627, n_35629;
wire n_35613, n_35614, n_35615, n_35616, n_35617, n_35618, n_35619, n_35620;
wire n_35602, n_35606, n_35607, n_35608, n_35609, n_35610, n_35611, n_35612;
wire n_35572, n_35576, n_35578, n_35580, n_35583, n_35590, n_35596, n_35600;
wire n_35529, n_35532, n_35537, n_35538, n_35540, n_35546, n_35555, n_35570;
wire n_35508, n_35514, n_35515, n_35519, n_35520, n_35523, n_35524, n_35528;
wire n_35468, n_35473, n_35478, n_35479, n_35485, n_35494, n_35500, n_35505;
wire n_35456, n_35457, n_35459, n_35462, n_35463, n_35464, n_35466, n_35467;
wire n_35447, n_35448, n_35449, n_35450, n_35452, n_35453, n_35454, n_35455;
wire n_35439, n_35440, n_35441, n_35442, n_35443, n_35444, n_35445, n_35446;
wire n_35430, n_35431, n_35432, n_35433, n_35434, n_35435, n_35436, n_35438;
wire n_35416, n_35417, n_35420, n_35423, n_35425, n_35426, n_35427, n_35429;
wire n_35408, n_35409, n_35410, n_35411, n_35412, n_35413, n_35414, n_35415;
wire n_35398, n_35399, n_35400, n_35401, n_35402, n_35403, n_35404, n_35407;
wire n_35390, n_35391, n_35392, n_35393, n_35394, n_35395, n_35396, n_35397;
wire n_35382, n_35383, n_35384, n_35385, n_35386, n_35387, n_35388, n_35389;
wire n_35359, n_35360, n_35361, n_35364, n_35366, n_35368, n_35380, n_35381;
wire n_35350, n_35351, n_35352, n_35353, n_35354, n_35355, n_35356, n_35357;
wire n_35342, n_35343, n_35344, n_35345, n_35346, n_35347, n_35348, n_35349;
wire n_35334, n_35335, n_35336, n_35337, n_35338, n_35339, n_35340, n_35341;
wire n_35324, n_35325, n_35326, n_35329, n_35330, n_35331, n_35332, n_35333;
wire n_35309, n_35310, n_35311, n_35313, n_35314, n_35315, n_35318, n_35321;
wire n_35301, n_35302, n_35303, n_35304, n_35305, n_35306, n_35307, n_35308;
wire n_35291, n_35292, n_35293, n_35295, n_35296, n_35298, n_35299, n_35300;
wire n_35283, n_35284, n_35285, n_35286, n_35287, n_35288, n_35289, n_35290;
wire n_35275, n_35276, n_35277, n_35278, n_35279, n_35280, n_35281, n_35282;
wire n_35267, n_35268, n_35269, n_35270, n_35271, n_35272, n_35273, n_35274;
wire n_35259, n_35260, n_35261, n_35262, n_35263, n_35264, n_35265, n_35266;
wire n_35250, n_35251, n_35252, n_35253, n_35254, n_35255, n_35256, n_35258;
wire n_35230, n_35231, n_35233, n_35244, n_35245, n_35247, n_35248, n_35249;
wire n_35215, n_35216, n_35217, n_35218, n_35221, n_35223, n_35224, n_35225;
wire n_35201, n_35202, n_35203, n_35205, n_35206, n_35208, n_35212, n_35214;
wire n_35179, n_35180, n_35188, n_35195, n_35196, n_35197, n_35198, n_35199;
wire n_35167, n_35168, n_35170, n_35171, n_35173, n_35174, n_35175, n_35176;
wire n_35159, n_35160, n_35161, n_35162, n_35163, n_35164, n_35165, n_35166;
wire n_35151, n_35152, n_35153, n_35154, n_35155, n_35156, n_35157, n_35158;
wire n_35142, n_35143, n_35144, n_35145, n_35146, n_35147, n_35148, n_35150;
wire n_35134, n_35135, n_35136, n_35137, n_35138, n_35139, n_35140, n_35141;
wire n_35124, n_35125, n_35126, n_35127, n_35128, n_35131, n_35132, n_35133;
wire n_35116, n_35117, n_35118, n_35119, n_35120, n_35121, n_35122, n_35123;
wire n_35108, n_35109, n_35110, n_35111, n_35112, n_35113, n_35114, n_35115;
wire n_35097, n_35098, n_35101, n_35102, n_35103, n_35104, n_35105, n_35107;
wire n_35089, n_35090, n_35091, n_35092, n_35093, n_35094, n_35095, n_35096;
wire n_35080, n_35081, n_35082, n_35084, n_35085, n_35086, n_35087, n_35088;
wire n_35063, n_35073, n_35074, n_35075, n_35076, n_35077, n_35078, n_35079;
wire n_35055, n_35056, n_35057, n_35058, n_35059, n_35060, n_35061, n_35062;
wire n_35047, n_35048, n_35049, n_35050, n_35051, n_35052, n_35053, n_35054;
wire n_35039, n_35040, n_35041, n_35042, n_35043, n_35044, n_35045, n_35046;
wire n_35021, n_35022, n_35023, n_35024, n_35035, n_35036, n_35037, n_35038;
wire n_35013, n_35014, n_35015, n_35016, n_35017, n_35018, n_35019, n_35020;
wire n_35005, n_35006, n_35007, n_35008, n_35009, n_35010, n_35011, n_35012;
wire n_34996, n_34997, n_34998, n_34999, n_35000, n_35001, n_35002, n_35003;
wire n_34985, n_34986, n_34987, n_34989, n_34991, n_34992, n_34993, n_34995;
wire n_34976, n_34977, n_34978, n_34979, n_34981, n_34982, n_34983, n_34984;
wire n_34961, n_34962, n_34963, n_34971, n_34972, n_34973, n_34974, n_34975;
wire n_34953, n_34954, n_34955, n_34956, n_34957, n_34958, n_34959, n_34960;
wire n_34944, n_34945, n_34946, n_34947, n_34948, n_34950, n_34951, n_34952;
wire n_34936, n_34937, n_34938, n_34939, n_34940, n_34941, n_34942, n_34943;
wire n_34928, n_34929, n_34930, n_34931, n_34932, n_34933, n_34934, n_34935;
wire n_34919, n_34920, n_34921, n_34923, n_34924, n_34925, n_34926, n_34927;
wire n_34874, n_34875, n_34912, n_34913, n_34915, n_34916, n_34917, n_34918;
wire n_34866, n_34867, n_34868, n_34869, n_34870, n_34871, n_34872, n_34873;
wire n_34858, n_34859, n_34860, n_34861, n_34862, n_34863, n_34864, n_34865;
wire n_34850, n_34851, n_34852, n_34853, n_34854, n_34855, n_34856, n_34857;
wire n_34837, n_34838, n_34841, n_34842, n_34843, n_34844, n_34845, n_34849;
wire n_34829, n_34830, n_34831, n_34832, n_34833, n_34834, n_34835, n_34836;
wire n_34821, n_34822, n_34823, n_34824, n_34825, n_34826, n_34827, n_34828;
wire n_34812, n_34813, n_34814, n_34815, n_34816, n_34817, n_34819, n_34820;
wire n_34803, n_34804, n_34805, n_34806, n_34807, n_34808, n_34809, n_34810;
wire n_34779, n_34780, n_34781, n_34784, n_34799, n_34800, n_34801, n_34802;
wire n_34769, n_34770, n_34771, n_34772, n_34773, n_34774, n_34775, n_34776;
wire n_34761, n_34762, n_34763, n_34764, n_34765, n_34766, n_34767, n_34768;
wire n_34749, n_34751, n_34752, n_34753, n_34756, n_34757, n_34758, n_34760;
wire n_34739, n_34740, n_34741, n_34742, n_34743, n_34744, n_34745, n_34746;
wire n_34725, n_34726, n_34731, n_34732, n_34733, n_34736, n_34737, n_34738;
wire n_34717, n_34718, n_34719, n_34720, n_34721, n_34722, n_34723, n_34724;
wire n_34708, n_34709, n_34711, n_34712, n_34713, n_34714, n_34715, n_34716;
wire n_34698, n_34699, n_34700, n_34701, n_34702, n_34703, n_34704, n_34706;
wire n_34690, n_34691, n_34692, n_34693, n_34694, n_34695, n_34696, n_34697;
wire n_34682, n_34683, n_34684, n_34685, n_34686, n_34687, n_34688, n_34689;
wire n_34674, n_34675, n_34676, n_34677, n_34678, n_34679, n_34680, n_34681;
wire n_34650, n_34651, n_34668, n_34669, n_34670, n_34671, n_34672, n_34673;
wire n_34617, n_34641, n_34642, n_34645, n_34646, n_34647, n_34648, n_34649;
wire n_34609, n_34610, n_34611, n_34612, n_34613, n_34614, n_34615, n_34616;
wire n_34601, n_34602, n_34603, n_34604, n_34605, n_34606, n_34607, n_34608;
wire n_34591, n_34592, n_34595, n_34596, n_34597, n_34598, n_34599, n_34600;
wire n_34583, n_34584, n_34585, n_34586, n_34587, n_34588, n_34589, n_34590;
wire n_34574, n_34575, n_34577, n_34578, n_34579, n_34580, n_34581, n_34582;
wire n_34555, n_34557, n_34568, n_34569, n_34570, n_34571, n_34572, n_34573;
wire n_34545, n_34546, n_34547, n_34548, n_34549, n_34551, n_34552, n_34554;
wire n_34537, n_34538, n_34539, n_34540, n_34541, n_34542, n_34543, n_34544;
wire n_34529, n_34530, n_34531, n_34532, n_34533, n_34534, n_34535, n_34536;
wire n_34520, n_34521, n_34522, n_34524, n_34525, n_34526, n_34527, n_34528;
wire n_34512, n_34513, n_34514, n_34515, n_34516, n_34517, n_34518, n_34519;
wire n_34503, n_34504, n_34505, n_34506, n_34507, n_34508, n_34509, n_34511;
wire n_34495, n_34496, n_34497, n_34498, n_34499, n_34500, n_34501, n_34502;
wire n_34487, n_34488, n_34489, n_34490, n_34491, n_34492, n_34493, n_34494;
wire n_34469, n_34470, n_34471, n_34472, n_34482, n_34483, n_34484, n_34485;
wire n_34451, n_34452, n_34453, n_34455, n_34465, n_34466, n_34467, n_34468;
wire n_34437, n_34438, n_34439, n_34440, n_34441, n_34445, n_34446, n_34450;
wire n_34428, n_34429, n_34430, n_34431, n_34432, n_34433, n_34434, n_34435;
wire n_34420, n_34421, n_34422, n_34423, n_34424, n_34425, n_34426, n_34427;
wire n_34410, n_34411, n_34412, n_34413, n_34415, n_34416, n_34417, n_34418;
wire n_34399, n_34400, n_34401, n_34403, n_34405, n_34407, n_34408, n_34409;
wire n_34389, n_34390, n_34391, n_34392, n_34393, n_34395, n_34396, n_34398;
wire n_34381, n_34382, n_34383, n_34384, n_34385, n_34386, n_34387, n_34388;
wire n_34363, n_34364, n_34372, n_34375, n_34377, n_34378, n_34379, n_34380;
wire n_34353, n_34354, n_34355, n_34356, n_34357, n_34358, n_34359, n_34362;
wire n_34324, n_34326, n_34330, n_34336, n_34349, n_34350, n_34351, n_34352;
wire n_34314, n_34317, n_34318, n_34319, n_34320, n_34321, n_34322, n_34323;
wire n_34304, n_34305, n_34306, n_34307, n_34308, n_34309, n_34310, n_34312;
wire n_34296, n_34297, n_34298, n_34299, n_34300, n_34301, n_34302, n_34303;
wire n_34286, n_34287, n_34288, n_34289, n_34290, n_34291, n_34292, n_34293;
wire n_34259, n_34264, n_34280, n_34281, n_34282, n_34283, n_34284, n_34285;
wire n_34230, n_34231, n_34232, n_34234, n_34235, n_34236, n_34237, n_34258;
wire n_34222, n_34223, n_34224, n_34225, n_34226, n_34227, n_34228, n_34229;
wire n_34211, n_34212, n_34213, n_34214, n_34215, n_34216, n_34220, n_34221;
wire n_34201, n_34203, n_34205, n_34206, n_34207, n_34208, n_34209, n_34210;
wire n_34190, n_34191, n_34192, n_34193, n_34194, n_34195, n_34196, n_34199;
wire n_34177, n_34178, n_34179, n_34180, n_34181, n_34187, n_34188, n_34189;
wire n_34163, n_34167, n_34171, n_34172, n_34173, n_34174, n_34175, n_34176;
wire n_34115, n_34116, n_34117, n_34118, n_34119, n_34120, n_34159, n_34160;
wire n_34106, n_34107, n_34108, n_34109, n_34110, n_34111, n_34112, n_34114;
wire n_34095, n_34096, n_34097, n_34098, n_34099, n_34100, n_34101, n_34104;
wire n_34087, n_34088, n_34089, n_34090, n_34091, n_34092, n_34093, n_34094;
wire n_34076, n_34077, n_34078, n_34079, n_34080, n_34081, n_34082, n_34086;
wire n_34067, n_34068, n_34069, n_34070, n_34071, n_34072, n_34073, n_34075;
wire n_34014, n_34015, n_34016, n_34062, n_34063, n_34064, n_34065, n_34066;
wire n_34005, n_34006, n_34007, n_34008, n_34009, n_34010, n_34011, n_34012;
wire n_33997, n_33998, n_33999, n_34000, n_34001, n_34002, n_34003, n_34004;
wire n_33985, n_33986, n_33989, n_33991, n_33993, n_33994, n_33995, n_33996;
wire n_33973, n_33976, n_33977, n_33979, n_33980, n_33981, n_33982, n_33983;
wire n_33963, n_33964, n_33967, n_33968, n_33969, n_33970, n_33971, n_33972;
wire n_33918, n_33920, n_33921, n_33922, n_33923, n_33924, n_33961, n_33962;
wire n_33909, n_33910, n_33911, n_33912, n_33914, n_33915, n_33916, n_33917;
wire n_33901, n_33902, n_33903, n_33904, n_33905, n_33906, n_33907, n_33908;
wire n_33859, n_33860, n_33894, n_33895, n_33896, n_33897, n_33898, n_33899;
wire n_33815, n_33816, n_33851, n_33852, n_33853, n_33854, n_33857, n_33858;
wire n_33807, n_33808, n_33809, n_33810, n_33811, n_33812, n_33813, n_33814;
wire n_33793, n_33799, n_33800, n_33801, n_33802, n_33803, n_33805, n_33806;
wire n_33784, n_33785, n_33786, n_33787, n_33788, n_33789, n_33790, n_33792;
wire n_33775, n_33776, n_33777, n_33778, n_33780, n_33781, n_33782, n_33783;
wire n_33755, n_33767, n_33768, n_33769, n_33770, n_33771, n_33772, n_33774;
wire n_33746, n_33748, n_33749, n_33750, n_33751, n_33752, n_33753, n_33754;
wire n_33734, n_33736, n_33737, n_33738, n_33739, n_33741, n_33744, n_33745;
wire n_33725, n_33726, n_33727, n_33728, n_33730, n_33731, n_33732, n_33733;
wire n_33717, n_33718, n_33719, n_33720, n_33721, n_33722, n_33723, n_33724;
wire n_33707, n_33708, n_33709, n_33710, n_33711, n_33712, n_33713, n_33716;
wire n_33677, n_33678, n_33679, n_33680, n_33681, n_33703, n_33705, n_33706;
wire n_33668, n_33670, n_33671, n_33672, n_33673, n_33674, n_33675, n_33676;
wire n_33658, n_33659, n_33661, n_33662, n_33663, n_33664, n_33665, n_33666;
wire n_33650, n_33651, n_33652, n_33653, n_33654, n_33655, n_33656, n_33657;
wire n_33642, n_33643, n_33644, n_33645, n_33646, n_33647, n_33648, n_33649;
wire n_33633, n_33634, n_33635, n_33636, n_33637, n_33638, n_33640, n_33641;
wire n_33624, n_33625, n_33626, n_33627, n_33629, n_33630, n_33631, n_33632;
wire n_33616, n_33617, n_33618, n_33619, n_33620, n_33621, n_33622, n_33623;
wire n_33608, n_33609, n_33610, n_33611, n_33612, n_33613, n_33614, n_33615;
wire n_33584, n_33585, n_33586, n_33587, n_33588, n_33589, n_33590, n_33592;
wire n_33576, n_33577, n_33578, n_33579, n_33580, n_33581, n_33582, n_33583;
wire n_33566, n_33567, n_33568, n_33570, n_33571, n_33572, n_33573, n_33574;
wire n_33557, n_33558, n_33559, n_33560, n_33561, n_33562, n_33563, n_33564;
wire n_33548, n_33550, n_33551, n_33552, n_33553, n_33554, n_33555, n_33556;
wire n_33540, n_33541, n_33542, n_33543, n_33544, n_33545, n_33546, n_33547;
wire n_33507, n_33509, n_33510, n_33511, n_33512, n_33513, n_33535, n_33536;
wire n_33498, n_33499, n_33500, n_33501, n_33503, n_33504, n_33505, n_33506;
wire n_33479, n_33480, n_33481, n_33485, n_33492, n_33494, n_33495, n_33496;
wire n_33457, n_33458, n_33473, n_33474, n_33475, n_33476, n_33477, n_33478;
wire n_33445, n_33446, n_33447, n_33448, n_33450, n_33454, n_33455, n_33456;
wire n_33429, n_33430, n_33431, n_33432, n_33433, n_33434, n_33436, n_33444;
wire n_33411, n_33412, n_33415, n_33416, n_33419, n_33420, n_33426, n_33427;
wire n_33403, n_33404, n_33405, n_33406, n_33407, n_33408, n_33409, n_33410;
wire n_33377, n_33378, n_33379, n_33380, n_33381, n_33382, n_33401, n_33402;
wire n_33368, n_33369, n_33370, n_33371, n_33373, n_33374, n_33375, n_33376;
wire n_33358, n_33361, n_33362, n_33363, n_33364, n_33365, n_33366, n_33367;
wire n_33350, n_33351, n_33352, n_33353, n_33354, n_33355, n_33356, n_33357;
wire n_33339, n_33340, n_33341, n_33345, n_33346, n_33347, n_33348, n_33349;
wire n_33330, n_33331, n_33332, n_33333, n_33335, n_33336, n_33337, n_33338;
wire n_33313, n_33314, n_33315, n_33316, n_33317, n_33318, n_33319, n_33329;
wire n_33302, n_33303, n_33304, n_33305, n_33309, n_33310, n_33311, n_33312;
wire n_33293, n_33295, n_33296, n_33297, n_33298, n_33299, n_33300, n_33301;
wire n_33280, n_33281, n_33286, n_33287, n_33288, n_33290, n_33291, n_33292;
wire n_33270, n_33271, n_33272, n_33273, n_33274, n_33275, n_33276, n_33277;
wire n_33250, n_33257, n_33261, n_33264, n_33265, n_33267, n_33268, n_33269;
wire n_33238, n_33239, n_33242, n_33243, n_33244, n_33245, n_33246, n_33247;
wire n_33227, n_33228, n_33230, n_33231, n_33232, n_33233, n_33234, n_33237;
wire n_33216, n_33217, n_33218, n_33220, n_33221, n_33222, n_33225, n_33226;
wire n_33198, n_33199, n_33200, n_33201, n_33209, n_33213, n_33214, n_33215;
wire n_33183, n_33184, n_33185, n_33188, n_33194, n_33195, n_33196, n_33197;
wire n_33170, n_33172, n_33173, n_33174, n_33175, n_33176, n_33180, n_33181;
wire n_33159, n_33161, n_33163, n_33164, n_33165, n_33166, n_33167, n_33168;
wire n_33135, n_33136, n_33138, n_33139, n_33140, n_33141, n_33156, n_33157;
wire n_33123, n_33124, n_33125, n_33127, n_33129, n_33131, n_33132, n_33133;
wire n_33114, n_33115, n_33116, n_33117, n_33118, n_33119, n_33120, n_33121;
wire n_33095, n_33097, n_33098, n_33099, n_33110, n_33111, n_33112, n_33113;
wire n_33085, n_33086, n_33088, n_33089, n_33091, n_33092, n_33093, n_33094;
wire n_33072, n_33077, n_33078, n_33079, n_33080, n_33081, n_33082, n_33084;
wire n_33051, n_33052, n_33053, n_33055, n_33058, n_33059, n_33068, n_33071;
wire n_33025, n_33026, n_33027, n_33031, n_33032, n_33034, n_33042, n_33046;
wire n_33009, n_33010, n_33011, n_33012, n_33015, n_33016, n_33017, n_33024;
wire n_32984, n_32992, n_32995, n_33000, n_33004, n_33006, n_33007, n_33008;
wire n_32969, n_32970, n_32971, n_32976, n_32977, n_32978, n_32979, n_32982;
wire n_32950, n_32951, n_32954, n_32956, n_32957, n_32959, n_32967, n_32968;
wire n_32935, n_32936, n_32938, n_32941, n_32944, n_32945, n_32947, n_32949;
wire n_32926, n_32927, n_32928, n_32929, n_32930, n_32932, n_32933, n_32934;
wire n_32918, n_32919, n_32920, n_32921, n_32922, n_32923, n_32924, n_32925;
wire n_32905, n_32908, n_32909, n_32913, n_32914, n_32915, n_32916, n_32917;
wire n_32893, n_32894, n_32899, n_32900, n_32901, n_32902, n_32903, n_32904;
wire n_32885, n_32886, n_32887, n_32888, n_32889, n_32890, n_32891, n_32892;
wire n_32877, n_32878, n_32879, n_32880, n_32881, n_32882, n_32883, n_32884;
wire n_32869, n_32870, n_32871, n_32872, n_32873, n_32874, n_32875, n_32876;
wire n_32856, n_32857, n_32858, n_32859, n_32862, n_32864, n_32867, n_32868;
wire n_32839, n_32841, n_32843, n_32844, n_32845, n_32847, n_32850, n_32851;
wire n_32817, n_32818, n_32827, n_32834, n_32835, n_32836, n_32837, n_32838;
wire n_32786, n_32791, n_32794, n_32798, n_32802, n_32803, n_32812, n_32815;
wire n_32764, n_32765, n_32767, n_32768, n_32770, n_32774, n_32777, n_32784;
wire n_32719, n_32720, n_32723, n_32728, n_32739, n_32745, n_32746, n_32748;
wire n_32697, n_32698, n_32707, n_32709, n_32710, n_32711, n_32715, n_32718;
wire n_32664, n_32669, n_32673, n_32675, n_32677, n_32683, n_32685, n_32690;
wire n_32642, n_32644, n_32646, n_32648, n_32649, n_32652, n_32654, n_32662;
wire n_32614, n_32615, n_32616, n_32620, n_32621, n_32637, n_32639, n_32641;
wire n_32599, n_32601, n_32602, n_32606, n_32607, n_32611, n_32612, n_32613;
wire n_32589, n_32590, n_32591, n_32592, n_32593, n_32596, n_32597, n_32598;
wire n_32571, n_32575, n_32576, n_32577, n_32578, n_32579, n_32580, n_32582;
wire n_32562, n_32563, n_32564, n_32565, n_32566, n_32568, n_32569, n_32570;
wire n_32544, n_32548, n_32550, n_32552, n_32556, n_32557, n_32560, n_32561;
wire n_32505, n_32509, n_32517, n_32532, n_32533, n_32535, n_32537, n_32543;
wire n_32487, n_32488, n_32489, n_32490, n_32496, n_32500, n_32501, n_32503;
wire n_32479, n_32480, n_32481, n_32482, n_32483, n_32484, n_32485, n_32486;
wire n_32448, n_32449, n_32450, n_32452, n_32453, n_32473, n_32475, n_32476;
wire n_32429, n_32430, n_32431, n_32432, n_32433, n_32435, n_32442, n_32445;
wire n_32401, n_32406, n_32409, n_32411, n_32412, n_32417, n_32426, n_32428;
wire n_32386, n_32388, n_32394, n_32395, n_32397, n_32398, n_32399, n_32400;
wire n_32371, n_32373, n_32374, n_32375, n_32378, n_32379, n_32381, n_32382;
wire n_32362, n_32363, n_32364, n_32365, n_32366, n_32367, n_32368, n_32369;
wire n_32343, n_32344, n_32349, n_32350, n_32356, n_32358, n_32359, n_32361;
wire n_32320, n_32321, n_32325, n_32334, n_32339, n_32340, n_32341, n_32342;
wire n_32308, n_32311, n_32313, n_32314, n_32315, n_32316, n_32317, n_32318;
wire n_32297, n_32299, n_32300, n_32301, n_32302, n_32303, n_32304, n_32307;
wire n_32287, n_32289, n_32290, n_32291, n_32293, n_32294, n_32295, n_32296;
wire n_32278, n_32279, n_32280, n_32281, n_32282, n_32283, n_32284, n_32286;
wire n_32270, n_32271, n_32272, n_32273, n_32274, n_32275, n_32276, n_32277;
wire n_32255, n_32260, n_32261, n_32263, n_32264, n_32265, n_32266, n_32269;
wire n_32245, n_32248, n_32249, n_32250, n_32251, n_32252, n_32253, n_32254;
wire n_32237, n_32238, n_32239, n_32240, n_32241, n_32242, n_32243, n_32244;
wire n_32222, n_32223, n_32224, n_32226, n_32230, n_32231, n_32235, n_32236;
wire n_32214, n_32215, n_32216, n_32217, n_32218, n_32219, n_32220, n_32221;
wire n_32204, n_32205, n_32206, n_32209, n_32210, n_32211, n_32212, n_32213;
wire n_32196, n_32197, n_32198, n_32199, n_32200, n_32201, n_32202, n_32203;
wire n_32172, n_32173, n_32174, n_32175, n_32180, n_32187, n_32188, n_32189;
wire n_32160, n_32161, n_32162, n_32163, n_32164, n_32166, n_32167, n_32171;
wire n_32150, n_32151, n_32152, n_32153, n_32156, n_32157, n_32158, n_32159;
wire n_32141, n_32142, n_32144, n_32145, n_32146, n_32147, n_32148, n_32149;
wire n_32132, n_32133, n_32134, n_32135, n_32136, n_32137, n_32138, n_32139;
wire n_32118, n_32119, n_32120, n_32121, n_32123, n_32125, n_32128, n_32129;
wire n_32109, n_32110, n_32112, n_32113, n_32114, n_32115, n_32116, n_32117;
wire n_32099, n_32100, n_32103, n_32104, n_32105, n_32106, n_32107, n_32108;
wire n_32089, n_32091, n_32092, n_32093, n_32094, n_32095, n_32096, n_32097;
wire n_32081, n_32082, n_32083, n_32084, n_32085, n_32086, n_32087, n_32088;
wire n_32070, n_32071, n_32072, n_32073, n_32076, n_32078, n_32079, n_32080;
wire n_32061, n_32062, n_32063, n_32064, n_32066, n_32067, n_32068, n_32069;
wire n_32052, n_32054, n_32055, n_32056, n_32057, n_32058, n_32059, n_32060;
wire n_32041, n_32042, n_32043, n_32045, n_32046, n_32049, n_32050, n_32051;
wire n_32020, n_32021, n_32022, n_32023, n_32028, n_32029, n_32039, n_32040;
wire n_32007, n_32008, n_32009, n_32010, n_32011, n_32015, n_32016, n_32019;
wire n_31998, n_31999, n_32000, n_32001, n_32002, n_32004, n_32005, n_32006;
wire n_31985, n_31986, n_31987, n_31988, n_31989, n_31990, n_31992, n_31993;
wire n_31974, n_31975, n_31976, n_31979, n_31980, n_31981, n_31983, n_31984;
wire n_31962, n_31965, n_31968, n_31969, n_31970, n_31971, n_31972, n_31973;
wire n_31948, n_31949, n_31950, n_31951, n_31954, n_31955, n_31958, n_31959;
wire n_31932, n_31933, n_31936, n_31937, n_31939, n_31942, n_31945, n_31946;
wire n_31923, n_31924, n_31925, n_31926, n_31927, n_31928, n_31929, n_31930;
wire n_31914, n_31915, n_31916, n_31917, n_31919, n_31920, n_31921, n_31922;
wire n_31904, n_31905, n_31907, n_31909, n_31910, n_31911, n_31912, n_31913;
wire n_31894, n_31895, n_31896, n_31897, n_31900, n_31901, n_31902, n_31903;
wire n_31882, n_31885, n_31886, n_31887, n_31888, n_31890, n_31891, n_31893;
wire n_31873, n_31874, n_31875, n_31876, n_31877, n_31878, n_31879, n_31881;
wire n_31862, n_31863, n_31865, n_31867, n_31868, n_31869, n_31871, n_31872;
wire n_31854, n_31855, n_31856, n_31857, n_31858, n_31859, n_31860, n_31861;
wire n_31845, n_31846, n_31847, n_31848, n_31849, n_31850, n_31851, n_31853;
wire n_31834, n_31835, n_31836, n_31837, n_31838, n_31840, n_31841, n_31844;
wire n_31820, n_31821, n_31822, n_31824, n_31825, n_31826, n_31827, n_31829;
wire n_31806, n_31810, n_31812, n_31813, n_31815, n_31816, n_31817, n_31819;
wire n_31798, n_31799, n_31800, n_31801, n_31802, n_31803, n_31804, n_31805;
wire n_31790, n_31791, n_31792, n_31793, n_31794, n_31795, n_31796, n_31797;
wire n_31781, n_31783, n_31784, n_31785, n_31786, n_31787, n_31788, n_31789;
wire n_31772, n_31773, n_31774, n_31776, n_31777, n_31778, n_31779, n_31780;
wire n_31763, n_31764, n_31765, n_31766, n_31767, n_31768, n_31769, n_31771;
wire n_31753, n_31754, n_31756, n_31758, n_31759, n_31760, n_31761, n_31762;
wire n_31741, n_31742, n_31744, n_31745, n_31746, n_31747, n_31748, n_31752;
wire n_31731, n_31732, n_31733, n_31734, n_31735, n_31736, n_31738, n_31740;
wire n_31723, n_31724, n_31725, n_31726, n_31727, n_31728, n_31729, n_31730;
wire n_31714, n_31715, n_31716, n_31717, n_31718, n_31719, n_31720, n_31722;
wire n_31705, n_31706, n_31707, n_31708, n_31710, n_31711, n_31712, n_31713;
wire n_31697, n_31698, n_31699, n_31700, n_31701, n_31702, n_31703, n_31704;
wire n_31689, n_31690, n_31691, n_31692, n_31693, n_31694, n_31695, n_31696;
wire n_31678, n_31679, n_31680, n_31681, n_31683, n_31685, n_31687, n_31688;
wire n_31668, n_31669, n_31670, n_31671, n_31672, n_31673, n_31676, n_31677;
wire n_31657, n_31658, n_31659, n_31660, n_31661, n_31664, n_31666, n_31667;
wire n_31649, n_31650, n_31651, n_31652, n_31653, n_31654, n_31655, n_31656;
wire n_31640, n_31641, n_31642, n_31644, n_31645, n_31646, n_31647, n_31648;
wire n_31630, n_31631, n_31632, n_31634, n_31636, n_31637, n_31638, n_31639;
wire n_31618, n_31619, n_31620, n_31621, n_31622, n_31623, n_31628, n_31629;
wire n_31608, n_31609, n_31610, n_31611, n_31613, n_31614, n_31616, n_31617;
wire n_31600, n_31601, n_31602, n_31603, n_31604, n_31605, n_31606, n_31607;
wire n_31590, n_31591, n_31592, n_31593, n_31594, n_31595, n_31596, n_31599;
wire n_31582, n_31583, n_31584, n_31585, n_31586, n_31587, n_31588, n_31589;
wire n_31574, n_31575, n_31576, n_31577, n_31578, n_31579, n_31580, n_31581;
wire n_31564, n_31566, n_31567, n_31568, n_31569, n_31570, n_31572, n_31573;
wire n_31556, n_31557, n_31558, n_31559, n_31560, n_31561, n_31562, n_31563;
wire n_31544, n_31545, n_31548, n_31549, n_31552, n_31553, n_31554, n_31555;
wire n_31534, n_31536, n_31538, n_31539, n_31540, n_31541, n_31542, n_31543;
wire n_31526, n_31527, n_31528, n_31529, n_31530, n_31531, n_31532, n_31533;
wire n_31517, n_31518, n_31520, n_31521, n_31522, n_31523, n_31524, n_31525;
wire n_31506, n_31507, n_31508, n_31509, n_31510, n_31511, n_31513, n_31514;
wire n_31498, n_31499, n_31500, n_31501, n_31502, n_31503, n_31504, n_31505;
wire n_31488, n_31489, n_31490, n_31491, n_31492, n_31493, n_31495, n_31497;
wire n_31479, n_31480, n_31481, n_31482, n_31483, n_31485, n_31486, n_31487;
wire n_31470, n_31471, n_31472, n_31473, n_31474, n_31475, n_31477, n_31478;
wire n_31458, n_31459, n_31460, n_31462, n_31463, n_31466, n_31467, n_31469;
wire n_31449, n_31450, n_31451, n_31452, n_31453, n_31454, n_31455, n_31457;
wire n_31437, n_31439, n_31441, n_31443, n_31444, n_31445, n_31446, n_31447;
wire n_31426, n_31428, n_31430, n_31431, n_31432, n_31434, n_31435, n_31436;
wire n_31416, n_31417, n_31418, n_31419, n_31420, n_31422, n_31423, n_31424;
wire n_31407, n_31408, n_31410, n_31411, n_31412, n_31413, n_31414, n_31415;
wire n_31399, n_31400, n_31401, n_31402, n_31403, n_31404, n_31405, n_31406;
wire n_31391, n_31392, n_31393, n_31394, n_31395, n_31396, n_31397, n_31398;
wire n_31383, n_31384, n_31385, n_31386, n_31387, n_31388, n_31389, n_31390;
wire n_31374, n_31375, n_31376, n_31377, n_31378, n_31379, n_31381, n_31382;
wire n_31365, n_31366, n_31367, n_31368, n_31369, n_31370, n_31371, n_31372;
wire n_31354, n_31356, n_31357, n_31358, n_31359, n_31360, n_31361, n_31362;
wire n_31346, n_31347, n_31348, n_31349, n_31350, n_31351, n_31352, n_31353;
wire n_31337, n_31338, n_31339, n_31340, n_31341, n_31343, n_31344, n_31345;
wire n_31329, n_31330, n_31331, n_31332, n_31333, n_31334, n_31335, n_31336;
wire n_31321, n_31322, n_31323, n_31324, n_31325, n_31326, n_31327, n_31328;
wire n_31311, n_31313, n_31314, n_31315, n_31316, n_31318, n_31319, n_31320;
wire n_31302, n_31303, n_31304, n_31305, n_31306, n_31307, n_31309, n_31310;
wire n_31294, n_31295, n_31296, n_31297, n_31298, n_31299, n_31300, n_31301;
wire n_31286, n_31287, n_31288, n_31289, n_31290, n_31291, n_31292, n_31293;
wire n_31278, n_31279, n_31280, n_31281, n_31282, n_31283, n_31284, n_31285;
wire n_31270, n_31271, n_31272, n_31273, n_31274, n_31275, n_31276, n_31277;
wire n_31262, n_31263, n_31264, n_31265, n_31266, n_31267, n_31268, n_31269;
wire n_31253, n_31255, n_31256, n_31257, n_31258, n_31259, n_31260, n_31261;
wire n_31245, n_31246, n_31247, n_31248, n_31249, n_31250, n_31251, n_31252;
wire n_31237, n_31238, n_31239, n_31240, n_31241, n_31242, n_31243, n_31244;
wire n_31227, n_31228, n_31229, n_31230, n_31232, n_31233, n_31234, n_31236;
wire n_31218, n_31220, n_31221, n_31222, n_31223, n_31224, n_31225, n_31226;
wire n_31208, n_31209, n_31210, n_31211, n_31212, n_31213, n_31214, n_31215;
wire n_31200, n_31201, n_31202, n_31203, n_31204, n_31205, n_31206, n_31207;
wire n_31190, n_31192, n_31193, n_31195, n_31196, n_31197, n_31198, n_31199;
wire n_31181, n_31182, n_31183, n_31184, n_31186, n_31187, n_31188, n_31189;
wire n_31173, n_31174, n_31175, n_31176, n_31177, n_31178, n_31179, n_31180;
wire n_31162, n_31164, n_31165, n_31167, n_31168, n_31169, n_31170, n_31171;
wire n_31154, n_31155, n_31156, n_31157, n_31158, n_31159, n_31160, n_31161;
wire n_31146, n_31147, n_31148, n_31149, n_31150, n_31151, n_31152, n_31153;
wire n_31135, n_31137, n_31138, n_31139, n_31141, n_31143, n_31144, n_31145;
wire n_31127, n_31128, n_31129, n_31130, n_31131, n_31132, n_31133, n_31134;
wire n_31119, n_31120, n_31121, n_31122, n_31123, n_31124, n_31125, n_31126;
wire n_31111, n_31112, n_31113, n_31114, n_31115, n_31116, n_31117, n_31118;
wire n_31103, n_31104, n_31105, n_31106, n_31107, n_31108, n_31109, n_31110;
wire n_31094, n_31095, n_31096, n_31097, n_31099, n_31100, n_31101, n_31102;
wire n_31083, n_31084, n_31085, n_31089, n_31090, n_31091, n_31092, n_31093;
wire n_31072, n_31073, n_31074, n_31075, n_31076, n_31079, n_31081, n_31082;
wire n_31064, n_31065, n_31066, n_31067, n_31068, n_31069, n_31070, n_31071;
wire n_31055, n_31056, n_31058, n_31059, n_31060, n_31061, n_31062, n_31063;
wire n_31045, n_31046, n_31047, n_31048, n_31049, n_31051, n_31052, n_31054;
wire n_31034, n_31035, n_31036, n_31037, n_31038, n_31040, n_31041, n_31043;
wire n_31023, n_31024, n_31025, n_31027, n_31028, n_31031, n_31032, n_31033;
wire n_31014, n_31015, n_31016, n_31017, n_31018, n_31019, n_31020, n_31021;
wire n_31004, n_31006, n_31007, n_31008, n_31009, n_31010, n_31012, n_31013;
wire n_30995, n_30996, n_30998, n_30999, n_31000, n_31001, n_31002, n_31003;
wire n_30987, n_30988, n_30989, n_30990, n_30991, n_30992, n_30993, n_30994;
wire n_30978, n_30979, n_30980, n_30981, n_30982, n_30983, n_30984, n_30986;
wire n_30968, n_30969, n_30970, n_30972, n_30974, n_30975, n_30976, n_30977;
wire n_30959, n_30960, n_30961, n_30962, n_30964, n_30965, n_30966, n_30967;
wire n_30951, n_30952, n_30953, n_30954, n_30955, n_30956, n_30957, n_30958;
wire n_30941, n_30942, n_30944, n_30945, n_30946, n_30947, n_30948, n_30949;
wire n_30933, n_30934, n_30935, n_30936, n_30937, n_30938, n_30939, n_30940;
wire n_30921, n_30924, n_30926, n_30927, n_30929, n_30930, n_30931, n_30932;
wire n_30910, n_30912, n_30913, n_30914, n_30915, n_30916, n_30917, n_30919;
wire n_30902, n_30903, n_30904, n_30905, n_30906, n_30907, n_30908, n_30909;
wire n_30894, n_30895, n_30896, n_30897, n_30898, n_30899, n_30900, n_30901;
wire n_30885, n_30886, n_30887, n_30888, n_30889, n_30890, n_30891, n_30893;
wire n_30876, n_30878, n_30879, n_30880, n_30881, n_30882, n_30883, n_30884;
wire n_30866, n_30867, n_30868, n_30869, n_30870, n_30873, n_30874, n_30875;
wire n_30856, n_30857, n_30858, n_30859, n_30860, n_30862, n_30864, n_30865;
wire n_30844, n_30846, n_30847, n_30848, n_30850, n_30851, n_30853, n_30854;
wire n_30835, n_30836, n_30837, n_30838, n_30839, n_30840, n_30841, n_30842;
wire n_30827, n_30828, n_30829, n_30830, n_30831, n_30832, n_30833, n_30834;
wire n_30817, n_30818, n_30819, n_30820, n_30823, n_30824, n_30825, n_30826;
wire n_30809, n_30810, n_30811, n_30812, n_30813, n_30814, n_30815, n_30816;
wire n_30799, n_30800, n_30801, n_30803, n_30804, n_30805, n_30807, n_30808;
wire n_30788, n_30789, n_30790, n_30791, n_30792, n_30793, n_30794, n_30795;
wire n_30780, n_30781, n_30782, n_30783, n_30784, n_30785, n_30786, n_30787;
wire n_30772, n_30773, n_30774, n_30775, n_30776, n_30777, n_30778, n_30779;
wire n_30764, n_30765, n_30766, n_30767, n_30768, n_30769, n_30770, n_30771;
wire n_30752, n_30753, n_30754, n_30755, n_30757, n_30759, n_30761, n_30762;
wire n_30743, n_30744, n_30745, n_30746, n_30747, n_30748, n_30750, n_30751;
wire n_30735, n_30736, n_30737, n_30738, n_30739, n_30740, n_30741, n_30742;
wire n_30727, n_30728, n_30729, n_30730, n_30731, n_30732, n_30733, n_30734;
wire n_30717, n_30718, n_30719, n_30720, n_30721, n_30722, n_30723, n_30726;
wire n_30708, n_30709, n_30711, n_30712, n_30713, n_30714, n_30715, n_30716;
wire n_30700, n_30701, n_30702, n_30703, n_30704, n_30705, n_30706, n_30707;
wire n_30691, n_30692, n_30694, n_30695, n_30696, n_30697, n_30698, n_30699;
wire n_30681, n_30682, n_30683, n_30684, n_30685, n_30686, n_30687, n_30689;
wire n_30668, n_30669, n_30673, n_30674, n_30675, n_30676, n_30678, n_30679;
wire n_30659, n_30660, n_30661, n_30662, n_30664, n_30665, n_30666, n_30667;
wire n_30650, n_30651, n_30652, n_30653, n_30655, n_30656, n_30657, n_30658;
wire n_30642, n_30643, n_30644, n_30645, n_30646, n_30647, n_30648, n_30649;
wire n_30634, n_30635, n_30636, n_30637, n_30638, n_30639, n_30640, n_30641;
wire n_30624, n_30626, n_30627, n_30628, n_30629, n_30630, n_30631, n_30632;
wire n_30615, n_30616, n_30617, n_30619, n_30620, n_30621, n_30622, n_30623;
wire n_30605, n_30606, n_30608, n_30610, n_30611, n_30612, n_30613, n_30614;
wire n_30595, n_30596, n_30597, n_30598, n_30599, n_30600, n_30601, n_30604;
wire n_30583, n_30584, n_30585, n_30586, n_30589, n_30590, n_30591, n_30594;
wire n_30575, n_30576, n_30577, n_30578, n_30579, n_30580, n_30581, n_30582;
wire n_30566, n_30567, n_30568, n_30569, n_30570, n_30571, n_30572, n_30573;
wire n_30554, n_30555, n_30557, n_30559, n_30561, n_30562, n_30563, n_30565;
wire n_30540, n_30541, n_30542, n_30543, n_30548, n_30549, n_30552, n_30553;
wire n_30530, n_30531, n_30533, n_30534, n_30535, n_30537, n_30538, n_30539;
wire n_30522, n_30523, n_30524, n_30525, n_30526, n_30527, n_30528, n_30529;
wire n_30512, n_30514, n_30515, n_30516, n_30517, n_30518, n_30520, n_30521;
wire n_30497, n_30498, n_30500, n_30501, n_30502, n_30504, n_30505, n_30507;
wire n_30488, n_30489, n_30491, n_30492, n_30493, n_30494, n_30495, n_30496;
wire n_30475, n_30476, n_30478, n_30480, n_30481, n_30482, n_30485, n_30487;
wire n_30467, n_30468, n_30469, n_30470, n_30471, n_30472, n_30473, n_30474;
wire n_30457, n_30459, n_30460, n_30461, n_30462, n_30463, n_30465, n_30466;
wire n_30449, n_30450, n_30451, n_30452, n_30453, n_30454, n_30455, n_30456;
wire n_30441, n_30442, n_30443, n_30444, n_30445, n_30446, n_30447, n_30448;
wire n_30432, n_30433, n_30435, n_30436, n_30437, n_30438, n_30439, n_30440;
wire n_30423, n_30424, n_30425, n_30427, n_30428, n_30429, n_30430, n_30431;
wire n_30415, n_30416, n_30417, n_30418, n_30419, n_30420, n_30421, n_30422;
wire n_30407, n_30408, n_30409, n_30410, n_30411, n_30412, n_30413, n_30414;
wire n_30394, n_30395, n_30397, n_30399, n_30403, n_30404, n_30405, n_30406;
wire n_30386, n_30387, n_30388, n_30389, n_30390, n_30391, n_30392, n_30393;
wire n_30378, n_30379, n_30380, n_30381, n_30382, n_30383, n_30384, n_30385;
wire n_30366, n_30368, n_30369, n_30373, n_30374, n_30375, n_30376, n_30377;
wire n_30355, n_30356, n_30360, n_30361, n_30362, n_30363, n_30364, n_30365;
wire n_30347, n_30348, n_30349, n_30350, n_30351, n_30352, n_30353, n_30354;
wire n_30336, n_30337, n_30338, n_30339, n_30341, n_30342, n_30345, n_30346;
wire n_30328, n_30329, n_30330, n_30331, n_30332, n_30333, n_30334, n_30335;
wire n_30320, n_30321, n_30322, n_30323, n_30324, n_30325, n_30326, n_30327;
wire n_30309, n_30311, n_30314, n_30315, n_30316, n_30317, n_30318, n_30319;
wire n_30298, n_30299, n_30300, n_30301, n_30302, n_30303, n_30304, n_30307;
wire n_30287, n_30288, n_30291, n_30292, n_30294, n_30295, n_30296, n_30297;
wire n_30278, n_30279, n_30280, n_30281, n_30282, n_30283, n_30285, n_30286;
wire n_30268, n_30269, n_30270, n_30271, n_30272, n_30273, n_30274, n_30277;
wire n_30260, n_30261, n_30262, n_30263, n_30264, n_30265, n_30266, n_30267;
wire n_30251, n_30253, n_30254, n_30255, n_30256, n_30257, n_30258, n_30259;
wire n_30240, n_30241, n_30242, n_30243, n_30244, n_30246, n_30247, n_30248;
wire n_30230, n_30232, n_30233, n_30234, n_30235, n_30237, n_30238, n_30239;
wire n_30222, n_30223, n_30224, n_30225, n_30226, n_30227, n_30228, n_30229;
wire n_30214, n_30215, n_30216, n_30217, n_30218, n_30219, n_30220, n_30221;
wire n_30200, n_30201, n_30203, n_30208, n_30210, n_30211, n_30212, n_30213;
wire n_30189, n_30190, n_30191, n_30192, n_30194, n_30195, n_30196, n_30197;
wire n_30180, n_30181, n_30182, n_30183, n_30184, n_30185, n_30187, n_30188;
wire n_30171, n_30172, n_30173, n_30174, n_30175, n_30176, n_30177, n_30179;
wire n_30163, n_30164, n_30165, n_30166, n_30167, n_30168, n_30169, n_30170;
wire n_30152, n_30153, n_30157, n_30158, n_30159, n_30160, n_30161, n_30162;
wire n_30143, n_30145, n_30146, n_30147, n_30148, n_30149, n_30150, n_30151;
wire n_30135, n_30136, n_30137, n_30138, n_30139, n_30140, n_30141, n_30142;
wire n_30126, n_30127, n_30128, n_30129, n_30130, n_30132, n_30133, n_30134;
wire n_30116, n_30117, n_30118, n_30119, n_30120, n_30121, n_30122, n_30125;
wire n_30106, n_30107, n_30108, n_30109, n_30110, n_30111, n_30113, n_30115;
wire n_30096, n_30097, n_30098, n_30099, n_30100, n_30103, n_30104, n_30105;
wire n_30085, n_30086, n_30087, n_30088, n_30090, n_30093, n_30094, n_30095;
wire n_30072, n_30075, n_30076, n_30079, n_30081, n_30082, n_30083, n_30084;
wire n_30062, n_30063, n_30064, n_30065, n_30066, n_30068, n_30070, n_30071;
wire n_30053, n_30054, n_30055, n_30056, n_30057, n_30058, n_30059, n_30061;
wire n_30045, n_30046, n_30047, n_30048, n_30049, n_30050, n_30051, n_30052;
wire n_30037, n_30038, n_30039, n_30040, n_30041, n_30042, n_30043, n_30044;
wire n_30027, n_30028, n_30029, n_30030, n_30033, n_30034, n_30035, n_30036;
wire n_30017, n_30018, n_30020, n_30022, n_30023, n_30024, n_30025, n_30026;
wire n_30005, n_30007, n_30008, n_30009, n_30010, n_30012, n_30013, n_30015;
wire n_29996, n_29997, n_29998, n_29999, n_30000, n_30002, n_30003, n_30004;
wire n_29985, n_29986, n_29988, n_29990, n_29991, n_29993, n_29994, n_29995;
wire n_29975, n_29976, n_29978, n_29980, n_29981, n_29982, n_29983, n_29984;
wire n_29966, n_29967, n_29968, n_29969, n_29970, n_29971, n_29972, n_29973;
wire n_29954, n_29955, n_29957, n_29958, n_29959, n_29960, n_29961, n_29962;
wire n_29944, n_29945, n_29947, n_29948, n_29950, n_29951, n_29952, n_29953;
wire n_29935, n_29936, n_29937, n_29938, n_29940, n_29941, n_29942, n_29943;
wire n_29925, n_29926, n_29927, n_29930, n_29931, n_29932, n_29933, n_29934;
wire n_29913, n_29915, n_29916, n_29917, n_29919, n_29920, n_29923, n_29924;
wire n_29904, n_29905, n_29906, n_29907, n_29908, n_29909, n_29910, n_29911;
wire n_29892, n_29893, n_29894, n_29898, n_29899, n_29900, n_29901, n_29902;
wire n_29883, n_29884, n_29885, n_29886, n_29887, n_29888, n_29889, n_29891;
wire n_29870, n_29871, n_29872, n_29873, n_29875, n_29878, n_29880, n_29881;
wire n_29862, n_29863, n_29864, n_29865, n_29866, n_29867, n_29868, n_29869;
wire n_29852, n_29853, n_29854, n_29855, n_29856, n_29859, n_29860, n_29861;
wire n_29841, n_29842, n_29843, n_29845, n_29848, n_29849, n_29850, n_29851;
wire n_29831, n_29832, n_29833, n_29834, n_29835, n_29836, n_29839, n_29840;
wire n_29819, n_29820, n_29822, n_29823, n_29825, n_29826, n_29827, n_29829;
wire n_29810, n_29811, n_29813, n_29814, n_29815, n_29816, n_29817, n_29818;
wire n_29802, n_29803, n_29804, n_29805, n_29806, n_29807, n_29808, n_29809;
wire n_29793, n_29794, n_29795, n_29796, n_29797, n_29798, n_29799, n_29801;
wire n_29785, n_29786, n_29787, n_29788, n_29789, n_29790, n_29791, n_29792;
wire n_29777, n_29778, n_29779, n_29780, n_29781, n_29782, n_29783, n_29784;
wire n_29766, n_29767, n_29768, n_29769, n_29770, n_29771, n_29775, n_29776;
wire n_29755, n_29758, n_29759, n_29760, n_29761, n_29762, n_29763, n_29765;
wire n_29744, n_29745, n_29746, n_29747, n_29749, n_29750, n_29751, n_29753;
wire n_29734, n_29736, n_29737, n_29738, n_29740, n_29741, n_29742, n_29743;
wire n_29724, n_29725, n_29726, n_29727, n_29729, n_29730, n_29732, n_29733;
wire n_29716, n_29717, n_29718, n_29719, n_29720, n_29721, n_29722, n_29723;
wire n_29707, n_29708, n_29709, n_29710, n_29711, n_29712, n_29714, n_29715;
wire n_29699, n_29700, n_29701, n_29702, n_29703, n_29704, n_29705, n_29706;
wire n_29688, n_29689, n_29690, n_29692, n_29693, n_29694, n_29695, n_29697;
wire n_29680, n_29681, n_29682, n_29683, n_29684, n_29685, n_29686, n_29687;
wire n_29671, n_29672, n_29673, n_29674, n_29676, n_29677, n_29678, n_29679;
wire n_29662, n_29663, n_29664, n_29665, n_29666, n_29667, n_29669, n_29670;
wire n_29654, n_29655, n_29656, n_29657, n_29658, n_29659, n_29660, n_29661;
wire n_29646, n_29647, n_29648, n_29649, n_29650, n_29651, n_29652, n_29653;
wire n_29637, n_29639, n_29640, n_29641, n_29642, n_29643, n_29644, n_29645;
wire n_29626, n_29627, n_29630, n_29632, n_29633, n_29634, n_29635, n_29636;
wire n_29618, n_29619, n_29620, n_29621, n_29622, n_29623, n_29624, n_29625;
wire n_29606, n_29607, n_29610, n_29611, n_29612, n_29613, n_29615, n_29616;
wire n_29594, n_29595, n_29596, n_29597, n_29598, n_29601, n_29604, n_29605;
wire n_29586, n_29587, n_29588, n_29589, n_29590, n_29591, n_29592, n_29593;
wire n_29576, n_29577, n_29578, n_29580, n_29582, n_29583, n_29584, n_29585;
wire n_29568, n_29569, n_29570, n_29571, n_29572, n_29573, n_29574, n_29575;
wire n_29559, n_29560, n_29561, n_29562, n_29563, n_29565, n_29566, n_29567;
wire n_29551, n_29552, n_29553, n_29554, n_29555, n_29556, n_29557, n_29558;
wire n_29538, n_29539, n_29540, n_29543, n_29544, n_29545, n_29547, n_29548;
wire n_29528, n_29530, n_29532, n_29533, n_29534, n_29535, n_29536, n_29537;
wire n_29519, n_29520, n_29521, n_29522, n_29523, n_29524, n_29526, n_29527;
wire n_29510, n_29511, n_29513, n_29514, n_29515, n_29516, n_29517, n_29518;
wire n_29501, n_29502, n_29503, n_29504, n_29505, n_29506, n_29507, n_29509;
wire n_29490, n_29491, n_29493, n_29494, n_29495, n_29496, n_29498, n_29500;
wire n_29480, n_29481, n_29482, n_29484, n_29485, n_29486, n_29487, n_29489;
wire n_29472, n_29473, n_29474, n_29475, n_29476, n_29477, n_29478, n_29479;
wire n_29462, n_29464, n_29465, n_29466, n_29467, n_29468, n_29470, n_29471;
wire n_29451, n_29453, n_29454, n_29455, n_29457, n_29458, n_29460, n_29461;
wire n_29441, n_29442, n_29443, n_29444, n_29445, n_29446, n_29447, n_29450;
wire n_29432, n_29433, n_29435, n_29436, n_29437, n_29438, n_29439, n_29440;
wire n_29423, n_29425, n_29426, n_29427, n_29428, n_29429, n_29430, n_29431;
wire n_29411, n_29412, n_29413, n_29415, n_29417, n_29419, n_29421, n_29422;
wire n_29400, n_29401, n_29404, n_29405, n_29406, n_29408, n_29409, n_29410;
wire n_29390, n_29391, n_29392, n_29394, n_29395, n_29396, n_29398, n_29399;
wire n_29381, n_29382, n_29383, n_29384, n_29385, n_29387, n_29388, n_29389;
wire n_29371, n_29372, n_29373, n_29374, n_29376, n_29378, n_29379, n_29380;
wire n_29363, n_29364, n_29365, n_29366, n_29367, n_29368, n_29369, n_29370;
wire n_29352, n_29353, n_29355, n_29356, n_29357, n_29359, n_29360, n_29361;
wire n_29342, n_29343, n_29344, n_29345, n_29346, n_29347, n_29348, n_29350;
wire n_29331, n_29332, n_29335, n_29337, n_29338, n_29339, n_29340, n_29341;
wire n_29323, n_29324, n_29325, n_29326, n_29327, n_29328, n_29329, n_29330;
wire n_29314, n_29315, n_29316, n_29317, n_29318, n_29319, n_29320, n_29321;
wire n_29306, n_29307, n_29308, n_29309, n_29310, n_29311, n_29312, n_29313;
wire n_29294, n_29295, n_29297, n_29298, n_29300, n_29302, n_29303, n_29305;
wire n_29285, n_29286, n_29287, n_29288, n_29290, n_29291, n_29292, n_29293;
wire n_29275, n_29276, n_29277, n_29278, n_29279, n_29282, n_29283, n_29284;
wire n_29263, n_29265, n_29267, n_29268, n_29269, n_29270, n_29272, n_29273;
wire n_29255, n_29256, n_29257, n_29258, n_29259, n_29260, n_29261, n_29262;
wire n_29244, n_29247, n_29248, n_29250, n_29251, n_29252, n_29253, n_29254;
wire n_29235, n_29236, n_29238, n_29239, n_29240, n_29241, n_29242, n_29243;
wire n_29226, n_29227, n_29228, n_29229, n_29230, n_29232, n_29233, n_29234;
wire n_29218, n_29219, n_29220, n_29221, n_29222, n_29223, n_29224, n_29225;
wire n_29209, n_29211, n_29212, n_29213, n_29214, n_29215, n_29216, n_29217;
wire n_29198, n_29199, n_29200, n_29201, n_29202, n_29204, n_29206, n_29208;
wire n_29190, n_29191, n_29192, n_29193, n_29194, n_29195, n_29196, n_29197;
wire n_29182, n_29183, n_29184, n_29185, n_29186, n_29187, n_29188, n_29189;
wire n_29172, n_29173, n_29174, n_29175, n_29177, n_29178, n_29179, n_29181;
wire n_29164, n_29165, n_29166, n_29167, n_29168, n_29169, n_29170, n_29171;
wire n_29156, n_29157, n_29158, n_29159, n_29160, n_29161, n_29162, n_29163;
wire n_29147, n_29148, n_29149, n_29150, n_29151, n_29153, n_29154, n_29155;
wire n_29139, n_29140, n_29141, n_29142, n_29143, n_29144, n_29145, n_29146;
wire n_29129, n_29131, n_29132, n_29133, n_29134, n_29135, n_29136, n_29138;
wire n_29119, n_29120, n_29121, n_29122, n_29123, n_29125, n_29127, n_29128;
wire n_29111, n_29112, n_29113, n_29114, n_29115, n_29116, n_29117, n_29118;
wire n_29100, n_29101, n_29103, n_29104, n_29105, n_29106, n_29108, n_29109;
wire n_29090, n_29091, n_29092, n_29093, n_29096, n_29097, n_29098, n_29099;
wire n_29081, n_29082, n_29083, n_29084, n_29085, n_29086, n_29088, n_29089;
wire n_29073, n_29074, n_29075, n_29076, n_29077, n_29078, n_29079, n_29080;
wire n_29064, n_29065, n_29066, n_29067, n_29068, n_29070, n_29071, n_29072;
wire n_29056, n_29057, n_29058, n_29059, n_29060, n_29061, n_29062, n_29063;
wire n_29047, n_29048, n_29049, n_29051, n_29052, n_29053, n_29054, n_29055;
wire n_29038, n_29039, n_29040, n_29042, n_29043, n_29044, n_29045, n_29046;
wire n_29028, n_29029, n_29032, n_29033, n_29034, n_29035, n_29036, n_29037;
wire n_29018, n_29019, n_29020, n_29023, n_29024, n_29025, n_29026, n_29027;
wire n_29007, n_29008, n_29009, n_29010, n_29011, n_29012, n_29014, n_29015;
wire n_28999, n_29000, n_29001, n_29002, n_29003, n_29004, n_29005, n_29006;
wire n_28990, n_28991, n_28992, n_28993, n_28994, n_28995, n_28996, n_28997;
wire n_28980, n_28982, n_28983, n_28984, n_28985, n_28986, n_28987, n_28988;
wire n_28971, n_28972, n_28974, n_28975, n_28976, n_28977, n_28978, n_28979;
wire n_28962, n_28963, n_28964, n_28965, n_28966, n_28967, n_28969, n_28970;
wire n_28953, n_28954, n_28955, n_28956, n_28957, n_28958, n_28959, n_28961;
wire n_28943, n_28944, n_28946, n_28947, n_28948, n_28949, n_28950, n_28951;
wire n_28931, n_28932, n_28934, n_28935, n_28939, n_28940, n_28941, n_28942;
wire n_28923, n_28924, n_28925, n_28926, n_28927, n_28928, n_28929, n_28930;
wire n_28915, n_28916, n_28917, n_28918, n_28919, n_28920, n_28921, n_28922;
wire n_28907, n_28908, n_28909, n_28910, n_28911, n_28912, n_28913, n_28914;
wire n_28896, n_28898, n_28899, n_28900, n_28901, n_28903, n_28905, n_28906;
wire n_28888, n_28889, n_28890, n_28891, n_28892, n_28893, n_28894, n_28895;
wire n_28880, n_28881, n_28882, n_28883, n_28884, n_28885, n_28886, n_28887;
wire n_28870, n_28871, n_28872, n_28874, n_28875, n_28876, n_28877, n_28879;
wire n_28860, n_28861, n_28862, n_28863, n_28864, n_28866, n_28867, n_28869;
wire n_28852, n_28853, n_28854, n_28855, n_28856, n_28857, n_28858, n_28859;
wire n_28840, n_28841, n_28843, n_28844, n_28845, n_28846, n_28849, n_28850;
wire n_28832, n_28833, n_28834, n_28835, n_28836, n_28837, n_28838, n_28839;
wire n_28824, n_28825, n_28826, n_28827, n_28828, n_28829, n_28830, n_28831;
wire n_28809, n_28813, n_28814, n_28816, n_28817, n_28818, n_28820, n_28822;
wire n_28798, n_28799, n_28802, n_28803, n_28804, n_28806, n_28807, n_28808;
wire n_28786, n_28787, n_28789, n_28790, n_28791, n_28793, n_28794, n_28796;
wire n_28778, n_28779, n_28780, n_28781, n_28782, n_28783, n_28784, n_28785;
wire n_28770, n_28771, n_28772, n_28773, n_28774, n_28775, n_28776, n_28777;
wire n_28762, n_28763, n_28764, n_28765, n_28766, n_28767, n_28768, n_28769;
wire n_28753, n_28754, n_28755, n_28756, n_28757, n_28759, n_28760, n_28761;
wire n_28744, n_28745, n_28746, n_28747, n_28748, n_28749, n_28750, n_28751;
wire n_28734, n_28736, n_28737, n_28738, n_28739, n_28740, n_28741, n_28743;
wire n_28725, n_28726, n_28728, n_28729, n_28730, n_28731, n_28732, n_28733;
wire n_28712, n_28713, n_28715, n_28718, n_28721, n_28722, n_28723, n_28724;
wire n_28704, n_28705, n_28706, n_28707, n_28708, n_28709, n_28710, n_28711;
wire n_28692, n_28693, n_28694, n_28695, n_28696, n_28698, n_28701, n_28702;
wire n_28683, n_28684, n_28685, n_28687, n_28688, n_28689, n_28690, n_28691;
wire n_28675, n_28676, n_28677, n_28678, n_28679, n_28680, n_28681, n_28682;
wire n_28667, n_28668, n_28669, n_28670, n_28671, n_28672, n_28673, n_28674;
wire n_28657, n_28658, n_28659, n_28661, n_28663, n_28664, n_28665, n_28666;
wire n_28648, n_28650, n_28651, n_28652, n_28653, n_28654, n_28655, n_28656;
wire n_28639, n_28640, n_28641, n_28642, n_28644, n_28645, n_28646, n_28647;
wire n_28630, n_28631, n_28633, n_28634, n_28635, n_28636, n_28637, n_28638;
wire n_28620, n_28622, n_28623, n_28624, n_28625, n_28626, n_28627, n_28628;
wire n_28610, n_28611, n_28612, n_28614, n_28615, n_28616, n_28618, n_28619;
wire n_28602, n_28603, n_28604, n_28605, n_28606, n_28607, n_28608, n_28609;
wire n_28593, n_28594, n_28595, n_28596, n_28597, n_28599, n_28600, n_28601;
wire n_28583, n_28584, n_28587, n_28588, n_28589, n_28590, n_28591, n_28592;
wire n_28575, n_28576, n_28577, n_28578, n_28579, n_28580, n_28581, n_28582;
wire n_28566, n_28567, n_28568, n_28569, n_28570, n_28572, n_28573, n_28574;
wire n_28555, n_28556, n_28557, n_28559, n_28560, n_28562, n_28563, n_28565;
wire n_28547, n_28548, n_28549, n_28550, n_28551, n_28552, n_28553, n_28554;
wire n_28536, n_28537, n_28538, n_28541, n_28542, n_28543, n_28545, n_28546;
wire n_28527, n_28528, n_28529, n_28530, n_28531, n_28532, n_28533, n_28535;
wire n_28518, n_28519, n_28521, n_28522, n_28523, n_28524, n_28525, n_28526;
wire n_28509, n_28510, n_28511, n_28513, n_28514, n_28515, n_28516, n_28517;
wire n_28501, n_28502, n_28503, n_28504, n_28505, n_28506, n_28507, n_28508;
wire n_28492, n_28493, n_28494, n_28495, n_28496, n_28497, n_28498, n_28500;
wire n_28484, n_28485, n_28486, n_28487, n_28488, n_28489, n_28490, n_28491;
wire n_28475, n_28476, n_28477, n_28479, n_28480, n_28481, n_28482, n_28483;
wire n_28465, n_28467, n_28468, n_28469, n_28471, n_28472, n_28473, n_28474;
wire n_28457, n_28458, n_28459, n_28460, n_28461, n_28462, n_28463, n_28464;
wire n_28449, n_28450, n_28451, n_28452, n_28453, n_28454, n_28455, n_28456;
wire n_28440, n_28441, n_28442, n_28443, n_28444, n_28445, n_28446, n_28448;
wire n_28431, n_28432, n_28433, n_28435, n_28436, n_28437, n_28438, n_28439;
wire n_28423, n_28424, n_28425, n_28426, n_28427, n_28428, n_28429, n_28430;
wire n_28415, n_28416, n_28417, n_28418, n_28419, n_28420, n_28421, n_28422;
wire n_28407, n_28408, n_28409, n_28410, n_28411, n_28412, n_28413, n_28414;
wire n_28398, n_28399, n_28400, n_28401, n_28402, n_28404, n_28405, n_28406;
wire n_28390, n_28391, n_28392, n_28393, n_28394, n_28395, n_28396, n_28397;
wire n_28381, n_28382, n_28383, n_28384, n_28385, n_28386, n_28387, n_28389;
wire n_28373, n_28374, n_28375, n_28376, n_28377, n_28378, n_28379, n_28380;
wire n_28364, n_28365, n_28366, n_28367, n_28368, n_28369, n_28371, n_28372;
wire n_28356, n_28357, n_28358, n_28359, n_28360, n_28361, n_28362, n_28363;
wire n_28346, n_28347, n_28348, n_28349, n_28352, n_28353, n_28354, n_28355;
wire n_28337, n_28338, n_28339, n_28341, n_28342, n_28343, n_28344, n_28345;
wire n_28329, n_28330, n_28331, n_28332, n_28333, n_28334, n_28335, n_28336;
wire n_28321, n_28322, n_28323, n_28324, n_28325, n_28326, n_28327, n_28328;
wire n_28312, n_28314, n_28315, n_28316, n_28317, n_28318, n_28319, n_28320;
wire n_28302, n_28304, n_28305, n_28306, n_28307, n_28308, n_28309, n_28310;
wire n_28293, n_28294, n_28295, n_28296, n_28298, n_28299, n_28300, n_28301;
wire n_28285, n_28286, n_28287, n_28288, n_28289, n_28290, n_28291, n_28292;
wire n_28276, n_28277, n_28279, n_28280, n_28281, n_28282, n_28283, n_28284;
wire n_28266, n_28267, n_28268, n_28270, n_28271, n_28273, n_28274, n_28275;
wire n_28255, n_28256, n_28258, n_28259, n_28260, n_28261, n_28263, n_28265;
wire n_28247, n_28248, n_28249, n_28250, n_28251, n_28252, n_28253, n_28254;
wire n_28238, n_28239, n_28240, n_28241, n_28242, n_28244, n_28245, n_28246;
wire n_28229, n_28230, n_28232, n_28233, n_28234, n_28235, n_28236, n_28237;
wire n_28220, n_28221, n_28222, n_28223, n_28224, n_28225, n_28226, n_28228;
wire n_28212, n_28213, n_28214, n_28215, n_28216, n_28217, n_28218, n_28219;
wire n_28204, n_28205, n_28206, n_28207, n_28208, n_28209, n_28210, n_28211;
wire n_28196, n_28197, n_28198, n_28199, n_28200, n_28201, n_28202, n_28203;
wire n_28186, n_28187, n_28190, n_28191, n_28192, n_28193, n_28194, n_28195;
wire n_28177, n_28178, n_28179, n_28180, n_28181, n_28182, n_28184, n_28185;
wire n_28168, n_28169, n_28171, n_28172, n_28173, n_28174, n_28175, n_28176;
wire n_28159, n_28160, n_28161, n_28162, n_28163, n_28165, n_28166, n_28167;
wire n_28151, n_28152, n_28153, n_28154, n_28155, n_28156, n_28157, n_28158;
wire n_28141, n_28142, n_28143, n_28144, n_28146, n_28147, n_28148, n_28150;
wire n_28132, n_28133, n_28134, n_28135, n_28136, n_28137, n_28138, n_28140;
wire n_28124, n_28125, n_28126, n_28127, n_28128, n_28129, n_28130, n_28131;
wire n_28116, n_28117, n_28118, n_28119, n_28120, n_28121, n_28122, n_28123;
wire n_28105, n_28106, n_28107, n_28108, n_28111, n_28113, n_28114, n_28115;
wire n_28094, n_28096, n_28097, n_28098, n_28099, n_28101, n_28103, n_28104;
wire n_28084, n_28086, n_28088, n_28089, n_28090, n_28091, n_28092, n_28093;
wire n_28076, n_28077, n_28078, n_28079, n_28080, n_28081, n_28082, n_28083;
wire n_28066, n_28067, n_28068, n_28069, n_28072, n_28073, n_28074, n_28075;
wire n_28056, n_28057, n_28058, n_28060, n_28061, n_28063, n_28064, n_28065;
wire n_28047, n_28048, n_28049, n_28050, n_28051, n_28052, n_28053, n_28054;
wire n_28039, n_28040, n_28041, n_28042, n_28043, n_28044, n_28045, n_28046;
wire n_28030, n_28031, n_28032, n_28034, n_28035, n_28036, n_28037, n_28038;
wire n_28020, n_28021, n_28023, n_28024, n_28025, n_28026, n_28027, n_28028;
wire n_28009, n_28011, n_28012, n_28013, n_28014, n_28017, n_28018, n_28019;
wire n_27998, n_27999, n_28000, n_28001, n_28003, n_28004, n_28007, n_28008;
wire n_27989, n_27990, n_27991, n_27992, n_27993, n_27994, n_27995, n_27996;
wire n_27981, n_27982, n_27983, n_27984, n_27985, n_27986, n_27987, n_27988;
wire n_27973, n_27974, n_27975, n_27976, n_27977, n_27978, n_27979, n_27980;
wire n_27961, n_27962, n_27963, n_27967, n_27968, n_27970, n_27971, n_27972;
wire n_27952, n_27954, n_27955, n_27956, n_27957, n_27958, n_27959, n_27960;
wire n_27944, n_27945, n_27946, n_27947, n_27948, n_27949, n_27950, n_27951;
wire n_27936, n_27937, n_27938, n_27939, n_27940, n_27941, n_27942, n_27943;
wire n_27927, n_27928, n_27929, n_27930, n_27931, n_27933, n_27934, n_27935;
wire n_27919, n_27920, n_27921, n_27922, n_27923, n_27924, n_27925, n_27926;
wire n_27910, n_27911, n_27912, n_27913, n_27914, n_27915, n_27916, n_27917;
wire n_27902, n_27903, n_27904, n_27905, n_27906, n_27907, n_27908, n_27909;
wire n_27894, n_27895, n_27896, n_27897, n_27898, n_27899, n_27900, n_27901;
wire n_27884, n_27885, n_27886, n_27887, n_27889, n_27890, n_27891, n_27892;
wire n_27875, n_27876, n_27877, n_27878, n_27879, n_27880, n_27882, n_27883;
wire n_27867, n_27868, n_27869, n_27870, n_27871, n_27872, n_27873, n_27874;
wire n_27858, n_27859, n_27861, n_27862, n_27863, n_27864, n_27865, n_27866;
wire n_27850, n_27851, n_27852, n_27853, n_27854, n_27855, n_27856, n_27857;
wire n_27841, n_27842, n_27843, n_27844, n_27845, n_27846, n_27847, n_27849;
wire n_27833, n_27834, n_27835, n_27836, n_27837, n_27838, n_27839, n_27840;
wire n_27824, n_27825, n_27826, n_27827, n_27828, n_27829, n_27831, n_27832;
wire n_27816, n_27817, n_27818, n_27819, n_27820, n_27821, n_27822, n_27823;
wire n_27807, n_27809, n_27810, n_27811, n_27812, n_27813, n_27814, n_27815;
wire n_27798, n_27799, n_27800, n_27801, n_27802, n_27803, n_27804, n_27805;
wire n_27789, n_27790, n_27791, n_27792, n_27793, n_27794, n_27795, n_27797;
wire n_27774, n_27775, n_27777, n_27778, n_27782, n_27783, n_27784, n_27786;
wire n_27766, n_27767, n_27768, n_27769, n_27770, n_27771, n_27772, n_27773;
wire n_27758, n_27759, n_27760, n_27761, n_27762, n_27763, n_27764, n_27765;
wire n_27748, n_27750, n_27751, n_27752, n_27754, n_27755, n_27756, n_27757;
wire n_27739, n_27741, n_27742, n_27743, n_27744, n_27745, n_27746, n_27747;
wire n_27730, n_27731, n_27732, n_27733, n_27734, n_27735, n_27736, n_27738;
wire n_27720, n_27721, n_27722, n_27725, n_27726, n_27727, n_27728, n_27729;
wire n_27711, n_27712, n_27714, n_27715, n_27716, n_27717, n_27718, n_27719;
wire n_27702, n_27704, n_27705, n_27706, n_27707, n_27708, n_27709, n_27710;
wire n_27691, n_27694, n_27695, n_27696, n_27697, n_27698, n_27699, n_27700;
wire n_27680, n_27681, n_27682, n_27683, n_27685, n_27686, n_27687, n_27689;
wire n_27672, n_27673, n_27674, n_27675, n_27676, n_27677, n_27678, n_27679;
wire n_27662, n_27663, n_27664, n_27665, n_27666, n_27667, n_27668, n_27671;
wire n_27654, n_27655, n_27656, n_27657, n_27658, n_27659, n_27660, n_27661;
wire n_27646, n_27647, n_27648, n_27649, n_27650, n_27651, n_27652, n_27653;
wire n_27636, n_27637, n_27638, n_27639, n_27640, n_27641, n_27644, n_27645;
wire n_27628, n_27629, n_27630, n_27631, n_27632, n_27633, n_27634, n_27635;
wire n_27619, n_27620, n_27621, n_27622, n_27623, n_27625, n_27626, n_27627;
wire n_27610, n_27611, n_27612, n_27613, n_27614, n_27615, n_27616, n_27618;
wire n_27601, n_27602, n_27603, n_27604, n_27606, n_27607, n_27608, n_27609;
wire n_27592, n_27593, n_27594, n_27595, n_27596, n_27598, n_27599, n_27600;
wire n_27584, n_27585, n_27586, n_27587, n_27588, n_27589, n_27590, n_27591;
wire n_27576, n_27577, n_27578, n_27579, n_27580, n_27581, n_27582, n_27583;
wire n_27567, n_27568, n_27569, n_27570, n_27571, n_27572, n_27573, n_27575;
wire n_27559, n_27560, n_27561, n_27562, n_27563, n_27564, n_27565, n_27566;
wire n_27550, n_27551, n_27553, n_27554, n_27555, n_27556, n_27557, n_27558;
wire n_27541, n_27542, n_27543, n_27544, n_27545, n_27547, n_27548, n_27549;
wire n_27532, n_27533, n_27534, n_27535, n_27536, n_27537, n_27538, n_27539;
wire n_27524, n_27525, n_27526, n_27527, n_27528, n_27529, n_27530, n_27531;
wire n_27516, n_27517, n_27518, n_27519, n_27520, n_27521, n_27522, n_27523;
wire n_27508, n_27509, n_27510, n_27511, n_27512, n_27513, n_27514, n_27515;
wire n_27499, n_27500, n_27501, n_27503, n_27504, n_27505, n_27506, n_27507;
wire n_27490, n_27491, n_27492, n_27493, n_27494, n_27495, n_27496, n_27498;
wire n_27480, n_27481, n_27483, n_27484, n_27485, n_27486, n_27487, n_27488;
wire n_27471, n_27472, n_27473, n_27475, n_27476, n_27477, n_27478, n_27479;
wire n_27463, n_27464, n_27465, n_27466, n_27467, n_27468, n_27469, n_27470;
wire n_27449, n_27450, n_27451, n_27453, n_27459, n_27460, n_27461, n_27462;
wire n_27440, n_27441, n_27442, n_27444, n_27445, n_27446, n_27447, n_27448;
wire n_27430, n_27431, n_27433, n_27434, n_27435, n_27436, n_27437, n_27438;
wire n_27422, n_27423, n_27424, n_27425, n_27426, n_27427, n_27428, n_27429;
wire n_27414, n_27415, n_27416, n_27417, n_27418, n_27419, n_27420, n_27421;
wire n_27403, n_27404, n_27405, n_27406, n_27407, n_27408, n_27409, n_27410;
wire n_27391, n_27395, n_27396, n_27397, n_27399, n_27400, n_27401, n_27402;
wire n_27382, n_27383, n_27384, n_27386, n_27387, n_27388, n_27389, n_27390;
wire n_27373, n_27374, n_27375, n_27376, n_27377, n_27378, n_27379, n_27380;
wire n_27364, n_27365, n_27366, n_27367, n_27368, n_27369, n_27370, n_27372;
wire n_27356, n_27357, n_27358, n_27359, n_27360, n_27361, n_27362, n_27363;
wire n_27346, n_27347, n_27348, n_27350, n_27351, n_27352, n_27353, n_27355;
wire n_27337, n_27338, n_27339, n_27340, n_27341, n_27342, n_27343, n_27345;
wire n_27329, n_27330, n_27331, n_27332, n_27333, n_27334, n_27335, n_27336;
wire n_27321, n_27322, n_27323, n_27324, n_27325, n_27326, n_27327, n_27328;
wire n_27311, n_27313, n_27315, n_27316, n_27317, n_27318, n_27319, n_27320;
wire n_27302, n_27303, n_27304, n_27306, n_27307, n_27308, n_27309, n_27310;
wire n_27294, n_27295, n_27296, n_27297, n_27298, n_27299, n_27300, n_27301;
wire n_27284, n_27285, n_27286, n_27287, n_27288, n_27289, n_27290, n_27292;
wire n_27274, n_27275, n_27277, n_27278, n_27280, n_27281, n_27282, n_27283;
wire n_27265, n_27266, n_27267, n_27269, n_27270, n_27271, n_27272, n_27273;
wire n_27257, n_27258, n_27259, n_27260, n_27261, n_27262, n_27263, n_27264;
wire n_27249, n_27250, n_27251, n_27252, n_27253, n_27254, n_27255, n_27256;
wire n_27240, n_27241, n_27243, n_27244, n_27245, n_27246, n_27247, n_27248;
wire n_27232, n_27233, n_27234, n_27235, n_27236, n_27237, n_27238, n_27239;
wire n_27221, n_27222, n_27225, n_27226, n_27227, n_27229, n_27230, n_27231;
wire n_27211, n_27212, n_27214, n_27215, n_27216, n_27217, n_27219, n_27220;
wire n_27200, n_27201, n_27203, n_27204, n_27205, n_27206, n_27207, n_27208;
wire n_27192, n_27193, n_27194, n_27195, n_27196, n_27197, n_27198, n_27199;
wire n_27181, n_27182, n_27183, n_27184, n_27185, n_27186, n_27189, n_27190;
wire n_27172, n_27174, n_27175, n_27176, n_27177, n_27178, n_27179, n_27180;
wire n_27163, n_27164, n_27166, n_27167, n_27168, n_27169, n_27170, n_27171;
wire n_27153, n_27154, n_27155, n_27157, n_27158, n_27159, n_27161, n_27162;
wire n_27144, n_27146, n_27147, n_27148, n_27149, n_27150, n_27151, n_27152;
wire n_27135, n_27136, n_27138, n_27139, n_27140, n_27141, n_27142, n_27143;
wire n_27126, n_27127, n_27128, n_27130, n_27131, n_27132, n_27133, n_27134;
wire n_27114, n_27115, n_27116, n_27117, n_27118, n_27119, n_27122, n_27125;
wire n_27103, n_27105, n_27106, n_27108, n_27109, n_27110, n_27111, n_27112;
wire n_27094, n_27095, n_27097, n_27098, n_27099, n_27100, n_27101, n_27102;
wire n_27085, n_27086, n_27088, n_27089, n_27090, n_27091, n_27092, n_27093;
wire n_27076, n_27077, n_27078, n_27079, n_27080, n_27081, n_27082, n_27083;
wire n_27066, n_27068, n_27069, n_27071, n_27072, n_27073, n_27074, n_27075;
wire n_27056, n_27058, n_27059, n_27061, n_27062, n_27063, n_27064, n_27065;
wire n_27047, n_27048, n_27049, n_27050, n_27051, n_27053, n_27054, n_27055;
wire n_27039, n_27040, n_27041, n_27042, n_27043, n_27044, n_27045, n_27046;
wire n_27028, n_27029, n_27031, n_27032, n_27033, n_27035, n_27036, n_27038;
wire n_27018, n_27019, n_27021, n_27022, n_27023, n_27024, n_27025, n_27026;
wire n_27010, n_27011, n_27012, n_27013, n_27014, n_27015, n_27016, n_27017;
wire n_27001, n_27002, n_27004, n_27005, n_27006, n_27007, n_27008, n_27009;
wire n_26991, n_26992, n_26993, n_26995, n_26996, n_26997, n_26998, n_27000;
wire n_26982, n_26983, n_26984, n_26985, n_26986, n_26987, n_26989, n_26990;
wire n_26974, n_26975, n_26976, n_26977, n_26978, n_26979, n_26980, n_26981;
wire n_26966, n_26967, n_26968, n_26969, n_26970, n_26971, n_26972, n_26973;
wire n_26958, n_26959, n_26960, n_26961, n_26962, n_26963, n_26964, n_26965;
wire n_26945, n_26946, n_26947, n_26948, n_26949, n_26950, n_26951, n_26952;
wire n_26936, n_26937, n_26938, n_26939, n_26940, n_26941, n_26942, n_26944;
wire n_26927, n_26928, n_26929, n_26930, n_26931, n_26933, n_26934, n_26935;
wire n_26919, n_26920, n_26921, n_26922, n_26923, n_26924, n_26925, n_26926;
wire n_26911, n_26912, n_26913, n_26914, n_26915, n_26916, n_26917, n_26918;
wire n_26899, n_26901, n_26902, n_26903, n_26904, n_26908, n_26909, n_26910;
wire n_26891, n_26892, n_26893, n_26894, n_26895, n_26896, n_26897, n_26898;
wire n_26883, n_26884, n_26885, n_26886, n_26887, n_26888, n_26889, n_26890;
wire n_26873, n_26875, n_26876, n_26877, n_26878, n_26879, n_26880, n_26881;
wire n_26865, n_26866, n_26867, n_26868, n_26869, n_26870, n_26871, n_26872;
wire n_26856, n_26857, n_26858, n_26860, n_26861, n_26862, n_26863, n_26864;
wire n_26846, n_26847, n_26848, n_26850, n_26852, n_26853, n_26854, n_26855;
wire n_26838, n_26839, n_26840, n_26841, n_26842, n_26843, n_26844, n_26845;
wire n_26830, n_26831, n_26832, n_26833, n_26834, n_26835, n_26836, n_26837;
wire n_26822, n_26823, n_26824, n_26825, n_26826, n_26827, n_26828, n_26829;
wire n_26813, n_26814, n_26815, n_26816, n_26818, n_26819, n_26820, n_26821;
wire n_26804, n_26805, n_26807, n_26808, n_26809, n_26810, n_26811, n_26812;
wire n_26794, n_26796, n_26797, n_26798, n_26799, n_26800, n_26801, n_26802;
wire n_26786, n_26787, n_26788, n_26789, n_26790, n_26791, n_26792, n_26793;
wire n_26778, n_26779, n_26780, n_26781, n_26782, n_26783, n_26784, n_26785;
wire n_26770, n_26771, n_26772, n_26773, n_26774, n_26775, n_26776, n_26777;
wire n_26760, n_26761, n_26762, n_26763, n_26765, n_26766, n_26767, n_26769;
wire n_26752, n_26753, n_26754, n_26755, n_26756, n_26757, n_26758, n_26759;
wire n_26743, n_26744, n_26745, n_26746, n_26747, n_26748, n_26749, n_26751;
wire n_26735, n_26736, n_26737, n_26738, n_26739, n_26740, n_26741, n_26742;
wire n_26727, n_26728, n_26729, n_26730, n_26731, n_26732, n_26733, n_26734;
wire n_26717, n_26718, n_26719, n_26720, n_26721, n_26723, n_26725, n_26726;
wire n_26707, n_26708, n_26710, n_26711, n_26712, n_26713, n_26715, n_26716;
wire n_26698, n_26699, n_26700, n_26702, n_26703, n_26704, n_26705, n_26706;
wire n_26689, n_26690, n_26691, n_26692, n_26694, n_26695, n_26696, n_26697;
wire n_26676, n_26677, n_26678, n_26680, n_26683, n_26684, n_26687, n_26688;
wire n_26665, n_26666, n_26668, n_26670, n_26671, n_26672, n_26673, n_26675;
wire n_26657, n_26658, n_26659, n_26660, n_26661, n_26662, n_26663, n_26664;
wire n_26648, n_26649, n_26650, n_26652, n_26653, n_26654, n_26655, n_26656;
wire n_26638, n_26639, n_26640, n_26641, n_26643, n_26644, n_26646, n_26647;
wire n_26630, n_26631, n_26632, n_26633, n_26634, n_26635, n_26636, n_26637;
wire n_26622, n_26623, n_26624, n_26625, n_26626, n_26627, n_26628, n_26629;
wire n_26612, n_26613, n_26614, n_26615, n_26616, n_26619, n_26620, n_26621;
wire n_26603, n_26605, n_26606, n_26607, n_26608, n_26609, n_26610, n_26611;
wire n_26595, n_26596, n_26597, n_26598, n_26599, n_26600, n_26601, n_26602;
wire n_26584, n_26585, n_26587, n_26588, n_26589, n_26590, n_26591, n_26594;
wire n_26575, n_26576, n_26577, n_26578, n_26580, n_26581, n_26582, n_26583;
wire n_26565, n_26568, n_26569, n_26570, n_26571, n_26572, n_26573, n_26574;
wire n_26553, n_26554, n_26557, n_26558, n_26559, n_26560, n_26562, n_26564;
wire n_26545, n_26546, n_26547, n_26548, n_26549, n_26550, n_26551, n_26552;
wire n_26535, n_26536, n_26538, n_26539, n_26540, n_26541, n_26542, n_26543;
wire n_26525, n_26528, n_26529, n_26530, n_26531, n_26532, n_26533, n_26534;
wire n_26516, n_26517, n_26519, n_26520, n_26521, n_26522, n_26523, n_26524;
wire n_26506, n_26507, n_26508, n_26509, n_26510, n_26511, n_26513, n_26514;
wire n_26497, n_26498, n_26499, n_26500, n_26502, n_26503, n_26504, n_26505;
wire n_26487, n_26488, n_26490, n_26491, n_26492, n_26493, n_26494, n_26496;
wire n_26478, n_26479, n_26480, n_26481, n_26482, n_26483, n_26485, n_26486;
wire n_26470, n_26471, n_26472, n_26473, n_26474, n_26475, n_26476, n_26477;
wire n_26459, n_26460, n_26461, n_26462, n_26463, n_26464, n_26465, n_26466;
wire n_26444, n_26447, n_26449, n_26450, n_26455, n_26456, n_26457, n_26458;
wire n_26435, n_26436, n_26438, n_26439, n_26440, n_26441, n_26442, n_26443;
wire n_26426, n_26427, n_26428, n_26430, n_26431, n_26432, n_26433, n_26434;
wire n_26418, n_26419, n_26420, n_26421, n_26422, n_26423, n_26424, n_26425;
wire n_26407, n_26408, n_26409, n_26411, n_26412, n_26415, n_26416, n_26417;
wire n_26396, n_26397, n_26398, n_26400, n_26401, n_26402, n_26404, n_26405;
wire n_26387, n_26389, n_26390, n_26391, n_26392, n_26393, n_26394, n_26395;
wire n_26377, n_26379, n_26380, n_26381, n_26382, n_26383, n_26385, n_26386;
wire n_26369, n_26370, n_26371, n_26372, n_26373, n_26374, n_26375, n_26376;
wire n_26361, n_26362, n_26363, n_26364, n_26365, n_26366, n_26367, n_26368;
wire n_26353, n_26354, n_26355, n_26356, n_26357, n_26358, n_26359, n_26360;
wire n_26345, n_26346, n_26347, n_26348, n_26349, n_26350, n_26351, n_26352;
wire n_26336, n_26337, n_26338, n_26339, n_26340, n_26341, n_26342, n_26344;
wire n_26327, n_26328, n_26330, n_26331, n_26332, n_26333, n_26334, n_26335;
wire n_26319, n_26320, n_26321, n_26322, n_26323, n_26324, n_26325, n_26326;
wire n_26311, n_26312, n_26313, n_26314, n_26315, n_26316, n_26317, n_26318;
wire n_26303, n_26304, n_26305, n_26306, n_26307, n_26308, n_26309, n_26310;
wire n_26295, n_26296, n_26297, n_26298, n_26299, n_26300, n_26301, n_26302;
wire n_26287, n_26288, n_26289, n_26290, n_26291, n_26292, n_26293, n_26294;
wire n_26279, n_26280, n_26281, n_26282, n_26283, n_26284, n_26285, n_26286;
wire n_26270, n_26271, n_26272, n_26273, n_26274, n_26275, n_26277, n_26278;
wire n_26260, n_26261, n_26262, n_26264, n_26265, n_26266, n_26268, n_26269;
wire n_26252, n_26253, n_26254, n_26255, n_26256, n_26257, n_26258, n_26259;
wire n_26244, n_26245, n_26246, n_26247, n_26248, n_26249, n_26250, n_26251;
wire n_26235, n_26236, n_26238, n_26239, n_26240, n_26241, n_26242, n_26243;
wire n_26225, n_26227, n_26229, n_26230, n_26231, n_26232, n_26233, n_26234;
wire n_26217, n_26218, n_26219, n_26220, n_26221, n_26222, n_26223, n_26224;
wire n_26208, n_26209, n_26210, n_26212, n_26213, n_26214, n_26215, n_26216;
wire n_26197, n_26199, n_26200, n_26202, n_26203, n_26204, n_26205, n_26207;
wire n_26186, n_26187, n_26189, n_26190, n_26192, n_26193, n_26194, n_26195;
wire n_26177, n_26178, n_26180, n_26181, n_26182, n_26183, n_26184, n_26185;
wire n_26169, n_26170, n_26171, n_26172, n_26173, n_26174, n_26175, n_26176;
wire n_26161, n_26162, n_26163, n_26164, n_26165, n_26166, n_26167, n_26168;
wire n_26152, n_26154, n_26155, n_26156, n_26157, n_26158, n_26159, n_26160;
wire n_26143, n_26144, n_26145, n_26146, n_26147, n_26148, n_26150, n_26151;
wire n_26133, n_26136, n_26137, n_26138, n_26139, n_26140, n_26141, n_26142;
wire n_26124, n_26125, n_26126, n_26128, n_26129, n_26130, n_26131, n_26132;
wire n_26115, n_26117, n_26118, n_26119, n_26120, n_26121, n_26122, n_26123;
wire n_26107, n_26108, n_26109, n_26110, n_26111, n_26112, n_26113, n_26114;
wire n_26099, n_26100, n_26101, n_26102, n_26103, n_26104, n_26105, n_26106;
wire n_26090, n_26091, n_26092, n_26094, n_26095, n_26096, n_26097, n_26098;
wire n_26077, n_26080, n_26082, n_26083, n_26084, n_26085, n_26087, n_26088;
wire n_26069, n_26070, n_26071, n_26072, n_26073, n_26074, n_26075, n_26076;
wire n_26059, n_26060, n_26061, n_26062, n_26063, n_26064, n_26067, n_26068;
wire n_26051, n_26052, n_26053, n_26054, n_26055, n_26056, n_26057, n_26058;
wire n_26040, n_26042, n_26043, n_26045, n_26046, n_26048, n_26049, n_26050;
wire n_26029, n_26030, n_26032, n_26033, n_26034, n_26036, n_26038, n_26039;
wire n_26021, n_26022, n_26023, n_26024, n_26025, n_26026, n_26027, n_26028;
wire n_26012, n_26013, n_26014, n_26015, n_26016, n_26017, n_26018, n_26020;
wire n_26004, n_26005, n_26006, n_26007, n_26008, n_26009, n_26010, n_26011;
wire n_25996, n_25997, n_25998, n_25999, n_26000, n_26001, n_26002, n_26003;
wire n_25988, n_25989, n_25990, n_25991, n_25992, n_25993, n_25994, n_25995;
wire n_25980, n_25981, n_25982, n_25983, n_25984, n_25985, n_25986, n_25987;
wire n_25972, n_25973, n_25974, n_25975, n_25976, n_25977, n_25978, n_25979;
wire n_25962, n_25964, n_25965, n_25966, n_25967, n_25968, n_25969, n_25970;
wire n_25954, n_25955, n_25956, n_25957, n_25958, n_25959, n_25960, n_25961;
wire n_25943, n_25945, n_25947, n_25948, n_25949, n_25951, n_25952, n_25953;
wire n_25926, n_25927, n_25928, n_25929, n_25937, n_25940, n_25941, n_25942;
wire n_25918, n_25919, n_25920, n_25921, n_25922, n_25923, n_25924, n_25925;
wire n_25909, n_25910, n_25911, n_25913, n_25914, n_25915, n_25916, n_25917;
wire n_25901, n_25902, n_25903, n_25904, n_25905, n_25906, n_25907, n_25908;
wire n_25891, n_25893, n_25894, n_25895, n_25896, n_25898, n_25899, n_25900;
wire n_25882, n_25883, n_25885, n_25886, n_25887, n_25888, n_25889, n_25890;
wire n_25873, n_25874, n_25875, n_25876, n_25877, n_25879, n_25880, n_25881;
wire n_25863, n_25865, n_25866, n_25867, n_25868, n_25870, n_25871, n_25872;
wire n_25855, n_25856, n_25857, n_25858, n_25859, n_25860, n_25861, n_25862;
wire n_25844, n_25845, n_25846, n_25847, n_25848, n_25849, n_25850, n_25852;
wire n_25835, n_25836, n_25837, n_25838, n_25839, n_25841, n_25842, n_25843;
wire n_25826, n_25827, n_25828, n_25829, n_25830, n_25832, n_25833, n_25834;
wire n_25817, n_25818, n_25820, n_25821, n_25822, n_25823, n_25824, n_25825;
wire n_25807, n_25808, n_25810, n_25811, n_25812, n_25813, n_25814, n_25815;
wire n_25795, n_25797, n_25798, n_25801, n_25802, n_25803, n_25805, n_25806;
wire n_25787, n_25788, n_25789, n_25790, n_25791, n_25792, n_25793, n_25794;
wire n_25779, n_25780, n_25781, n_25782, n_25783, n_25784, n_25785, n_25786;
wire n_25770, n_25771, n_25772, n_25774, n_25775, n_25776, n_25777, n_25778;
wire n_25762, n_25763, n_25764, n_25765, n_25766, n_25767, n_25768, n_25769;
wire n_25752, n_25753, n_25755, n_25756, n_25757, n_25758, n_25759, n_25761;
wire n_25744, n_25745, n_25746, n_25747, n_25748, n_25749, n_25750, n_25751;
wire n_25734, n_25735, n_25736, n_25737, n_25738, n_25739, n_25740, n_25742;
wire n_25723, n_25724, n_25725, n_25727, n_25728, n_25729, n_25730, n_25732;
wire n_25713, n_25715, n_25716, n_25717, n_25719, n_25720, n_25721, n_25722;
wire n_25704, n_25705, n_25706, n_25707, n_25708, n_25709, n_25710, n_25712;
wire n_25694, n_25695, n_25696, n_25698, n_25699, n_25701, n_25702, n_25703;
wire n_25686, n_25687, n_25688, n_25689, n_25690, n_25691, n_25692, n_25693;
wire n_25677, n_25678, n_25679, n_25680, n_25681, n_25682, n_25683, n_25684;
wire n_25667, n_25668, n_25669, n_25670, n_25671, n_25672, n_25673, n_25675;
wire n_25657, n_25658, n_25659, n_25660, n_25661, n_25662, n_25664, n_25666;
wire n_25648, n_25649, n_25651, n_25652, n_25653, n_25654, n_25655, n_25656;
wire n_25640, n_25641, n_25642, n_25643, n_25644, n_25645, n_25646, n_25647;
wire n_25631, n_25632, n_25633, n_25634, n_25635, n_25636, n_25637, n_25638;
wire n_25623, n_25624, n_25625, n_25626, n_25627, n_25628, n_25629, n_25630;
wire n_25615, n_25616, n_25617, n_25618, n_25619, n_25620, n_25621, n_25622;
wire n_25606, n_25607, n_25608, n_25609, n_25610, n_25611, n_25612, n_25613;
wire n_25596, n_25598, n_25599, n_25600, n_25602, n_25603, n_25604, n_25605;
wire n_25587, n_25589, n_25590, n_25591, n_25592, n_25593, n_25594, n_25595;
wire n_25578, n_25579, n_25580, n_25581, n_25582, n_25583, n_25584, n_25586;
wire n_25570, n_25571, n_25572, n_25573, n_25574, n_25575, n_25576, n_25577;
wire n_25562, n_25563, n_25564, n_25565, n_25566, n_25567, n_25568, n_25569;
wire n_25554, n_25555, n_25556, n_25557, n_25558, n_25559, n_25560, n_25561;
wire n_25544, n_25545, n_25546, n_25547, n_25548, n_25550, n_25552, n_25553;
wire n_25535, n_25536, n_25537, n_25538, n_25539, n_25540, n_25541, n_25543;
wire n_25527, n_25528, n_25529, n_25530, n_25531, n_25532, n_25533, n_25534;
wire n_25517, n_25519, n_25520, n_25521, n_25522, n_25523, n_25525, n_25526;
wire n_25505, n_25506, n_25507, n_25508, n_25513, n_25514, n_25515, n_25516;
wire n_25497, n_25498, n_25499, n_25500, n_25501, n_25502, n_25503, n_25504;
wire n_25489, n_25490, n_25491, n_25492, n_25493, n_25494, n_25495, n_25496;
wire n_25481, n_25482, n_25483, n_25484, n_25485, n_25486, n_25487, n_25488;
wire n_25473, n_25474, n_25475, n_25476, n_25477, n_25478, n_25479, n_25480;
wire n_25464, n_25465, n_25466, n_25467, n_25469, n_25470, n_25471, n_25472;
wire n_25454, n_25455, n_25456, n_25457, n_25460, n_25461, n_25462, n_25463;
wire n_25446, n_25447, n_25448, n_25449, n_25450, n_25451, n_25452, n_25453;
wire n_25436, n_25437, n_25438, n_25439, n_25441, n_25442, n_25443, n_25444;
wire n_25427, n_25429, n_25430, n_25431, n_25432, n_25433, n_25434, n_25435;
wire n_25417, n_25419, n_25421, n_25422, n_25423, n_25424, n_25425, n_25426;
wire n_25409, n_25410, n_25411, n_25412, n_25413, n_25414, n_25415, n_25416;
wire n_25400, n_25402, n_25403, n_25404, n_25405, n_25406, n_25407, n_25408;
wire n_25390, n_25391, n_25392, n_25393, n_25394, n_25395, n_25396, n_25399;
wire n_25382, n_25383, n_25384, n_25385, n_25386, n_25387, n_25388, n_25389;
wire n_25374, n_25375, n_25376, n_25377, n_25378, n_25379, n_25380, n_25381;
wire n_25365, n_25366, n_25367, n_25368, n_25369, n_25371, n_25372, n_25373;
wire n_25355, n_25357, n_25359, n_25360, n_25361, n_25362, n_25363, n_25364;
wire n_25346, n_25347, n_25348, n_25350, n_25351, n_25352, n_25353, n_25354;
wire n_25338, n_25339, n_25340, n_25341, n_25342, n_25343, n_25344, n_25345;
wire n_25326, n_25327, n_25328, n_25329, n_25331, n_25335, n_25336, n_25337;
wire n_25318, n_25319, n_25320, n_25321, n_25322, n_25323, n_25324, n_25325;
wire n_25308, n_25309, n_25311, n_25312, n_25313, n_25315, n_25316, n_25317;
wire n_25299, n_25301, n_25302, n_25303, n_25304, n_25305, n_25306, n_25307;
wire n_25290, n_25292, n_25293, n_25294, n_25295, n_25296, n_25297, n_25298;
wire n_25279, n_25283, n_25284, n_25285, n_25286, n_25287, n_25288, n_25289;
wire n_25270, n_25271, n_25272, n_25274, n_25275, n_25276, n_25277, n_25278;
wire n_25260, n_25261, n_25262, n_25263, n_25264, n_25266, n_25268, n_25269;
wire n_25251, n_25252, n_25253, n_25255, n_25256, n_25257, n_25258, n_25259;
wire n_25243, n_25244, n_25245, n_25246, n_25247, n_25248, n_25249, n_25250;
wire n_25235, n_25236, n_25237, n_25238, n_25239, n_25240, n_25241, n_25242;
wire n_25226, n_25228, n_25229, n_25230, n_25231, n_25232, n_25233, n_25234;
wire n_25217, n_25219, n_25220, n_25221, n_25222, n_25223, n_25224, n_25225;
wire n_25209, n_25210, n_25211, n_25212, n_25213, n_25214, n_25215, n_25216;
wire n_25201, n_25202, n_25203, n_25204, n_25205, n_25206, n_25207, n_25208;
wire n_25193, n_25194, n_25195, n_25196, n_25197, n_25198, n_25199, n_25200;
wire n_25177, n_25178, n_25179, n_25180, n_25181, n_25182, n_25183, n_25185;
wire n_25168, n_25169, n_25170, n_25171, n_25172, n_25173, n_25175, n_25176;
wire n_25160, n_25161, n_25162, n_25163, n_25164, n_25165, n_25166, n_25167;
wire n_25151, n_25152, n_25153, n_25154, n_25155, n_25157, n_25158, n_25159;
wire n_25143, n_25144, n_25145, n_25146, n_25147, n_25148, n_25149, n_25150;
wire n_25135, n_25136, n_25137, n_25138, n_25139, n_25140, n_25141, n_25142;
wire n_25127, n_25128, n_25129, n_25130, n_25131, n_25132, n_25133, n_25134;
wire n_25119, n_25120, n_25121, n_25122, n_25123, n_25124, n_25125, n_25126;
wire n_25109, n_25110, n_25111, n_25112, n_25113, n_25115, n_25116, n_25118;
wire n_25099, n_25100, n_25101, n_25102, n_25103, n_25105, n_25106, n_25107;
wire n_25088, n_25089, n_25092, n_25094, n_25095, n_25096, n_25097, n_25098;
wire n_25079, n_25080, n_25081, n_25082, n_25083, n_25084, n_25085, n_25086;
wire n_25070, n_25071, n_25072, n_25073, n_25074, n_25075, n_25076, n_25078;
wire n_25062, n_25063, n_25064, n_25065, n_25066, n_25067, n_25068, n_25069;
wire n_25053, n_25054, n_25055, n_25056, n_25057, n_25058, n_25059, n_25061;
wire n_25043, n_25046, n_25047, n_25048, n_25049, n_25050, n_25051, n_25052;
wire n_25032, n_25033, n_25034, n_25035, n_25037, n_25038, n_25039, n_25041;
wire n_25022, n_25023, n_25024, n_25025, n_25027, n_25028, n_25029, n_25030;
wire n_25014, n_25015, n_25016, n_25017, n_25018, n_25019, n_25020, n_25021;
wire n_25004, n_25005, n_25006, n_25007, n_25008, n_25009, n_25010, n_25011;
wire n_24993, n_24994, n_24995, n_24997, n_24998, n_24999, n_25001, n_25003;
wire n_24985, n_24986, n_24987, n_24988, n_24989, n_24990, n_24991, n_24992;
wire n_24977, n_24978, n_24979, n_24980, n_24981, n_24982, n_24983, n_24984;
wire n_24965, n_24966, n_24970, n_24971, n_24972, n_24973, n_24975, n_24976;
wire n_24950, n_24951, n_24955, n_24959, n_24960, n_24962, n_24963, n_24964;
wire n_24941, n_24942, n_24943, n_24944, n_24945, n_24946, n_24947, n_24949;
wire n_24932, n_24933, n_24934, n_24935, n_24936, n_24937, n_24938, n_24940;
wire n_24924, n_24925, n_24926, n_24927, n_24928, n_24929, n_24930, n_24931;
wire n_24914, n_24915, n_24917, n_24918, n_24919, n_24920, n_24922, n_24923;
wire n_24904, n_24905, n_24907, n_24908, n_24909, n_24911, n_24912, n_24913;
wire n_24895, n_24896, n_24897, n_24898, n_24899, n_24900, n_24901, n_24903;
wire n_24887, n_24888, n_24889, n_24890, n_24891, n_24892, n_24893, n_24894;
wire n_24879, n_24880, n_24881, n_24882, n_24883, n_24884, n_24885, n_24886;
wire n_24869, n_24871, n_24872, n_24873, n_24874, n_24875, n_24876, n_24877;
wire n_24860, n_24861, n_24863, n_24864, n_24865, n_24866, n_24867, n_24868;
wire n_24847, n_24848, n_24850, n_24852, n_24853, n_24857, n_24858, n_24859;
wire n_24838, n_24839, n_24840, n_24841, n_24842, n_24843, n_24844, n_24845;
wire n_24829, n_24830, n_24831, n_24832, n_24833, n_24835, n_24836, n_24837;
wire n_24821, n_24822, n_24823, n_24824, n_24825, n_24826, n_24827, n_24828;
wire n_24812, n_24814, n_24815, n_24816, n_24817, n_24818, n_24819, n_24820;
wire n_24804, n_24805, n_24806, n_24807, n_24808, n_24809, n_24810, n_24811;
wire n_24795, n_24796, n_24797, n_24798, n_24799, n_24801, n_24802, n_24803;
wire n_24787, n_24788, n_24789, n_24790, n_24791, n_24792, n_24793, n_24794;
wire n_24777, n_24779, n_24780, n_24781, n_24782, n_24783, n_24785, n_24786;
wire n_24769, n_24770, n_24771, n_24772, n_24773, n_24774, n_24775, n_24776;
wire n_24760, n_24761, n_24762, n_24763, n_24764, n_24765, n_24766, n_24767;
wire n_24752, n_24753, n_24754, n_24755, n_24756, n_24757, n_24758, n_24759;
wire n_24744, n_24745, n_24746, n_24747, n_24748, n_24749, n_24750, n_24751;
wire n_24734, n_24735, n_24737, n_24738, n_24739, n_24741, n_24742, n_24743;
wire n_24725, n_24726, n_24727, n_24728, n_24729, n_24731, n_24732, n_24733;
wire n_24716, n_24717, n_24718, n_24719, n_24721, n_24722, n_24723, n_24724;
wire n_24706, n_24708, n_24709, n_24710, n_24711, n_24712, n_24713, n_24715;
wire n_24698, n_24699, n_24700, n_24701, n_24702, n_24703, n_24704, n_24705;
wire n_24688, n_24689, n_24692, n_24693, n_24694, n_24695, n_24696, n_24697;
wire n_24679, n_24680, n_24681, n_24682, n_24684, n_24685, n_24686, n_24687;
wire n_24671, n_24672, n_24673, n_24674, n_24675, n_24676, n_24677, n_24678;
wire n_24663, n_24664, n_24665, n_24666, n_24667, n_24668, n_24669, n_24670;
wire n_24655, n_24656, n_24657, n_24658, n_24659, n_24660, n_24661, n_24662;
wire n_24647, n_24648, n_24649, n_24650, n_24651, n_24652, n_24653, n_24654;
wire n_24639, n_24640, n_24641, n_24642, n_24643, n_24644, n_24645, n_24646;
wire n_24627, n_24628, n_24629, n_24630, n_24631, n_24632, n_24633, n_24638;
wire n_24619, n_24620, n_24621, n_24622, n_24623, n_24624, n_24625, n_24626;
wire n_24611, n_24612, n_24613, n_24614, n_24615, n_24616, n_24617, n_24618;
wire n_24603, n_24604, n_24605, n_24606, n_24607, n_24608, n_24609, n_24610;
wire n_24593, n_24594, n_24595, n_24597, n_24599, n_24600, n_24601, n_24602;
wire n_24583, n_24584, n_24585, n_24586, n_24588, n_24589, n_24590, n_24592;
wire n_24575, n_24576, n_24577, n_24578, n_24579, n_24580, n_24581, n_24582;
wire n_24565, n_24566, n_24567, n_24569, n_24571, n_24572, n_24573, n_24574;
wire n_24557, n_24558, n_24559, n_24560, n_24561, n_24562, n_24563, n_24564;
wire n_24548, n_24549, n_24550, n_24552, n_24553, n_24554, n_24555, n_24556;
wire n_24538, n_24539, n_24540, n_24542, n_24543, n_24545, n_24546, n_24547;
wire n_24528, n_24529, n_24530, n_24531, n_24532, n_24534, n_24535, n_24537;
wire n_24518, n_24519, n_24521, n_24523, n_24524, n_24525, n_24526, n_24527;
wire n_24509, n_24510, n_24511, n_24512, n_24513, n_24514, n_24516, n_24517;
wire n_24500, n_24501, n_24502, n_24503, n_24505, n_24506, n_24507, n_24508;
wire n_24491, n_24492, n_24493, n_24494, n_24495, n_24497, n_24498, n_24499;
wire n_24483, n_24484, n_24485, n_24486, n_24487, n_24488, n_24489, n_24490;
wire n_24474, n_24476, n_24477, n_24478, n_24479, n_24480, n_24481, n_24482;
wire n_24466, n_24467, n_24468, n_24469, n_24470, n_24471, n_24472, n_24473;
wire n_24458, n_24459, n_24460, n_24461, n_24462, n_24463, n_24464, n_24465;
wire n_24448, n_24449, n_24451, n_24452, n_24453, n_24454, n_24455, n_24457;
wire n_24440, n_24441, n_24442, n_24443, n_24444, n_24445, n_24446, n_24447;
wire n_24432, n_24433, n_24434, n_24435, n_24436, n_24437, n_24438, n_24439;
wire n_24424, n_24425, n_24426, n_24427, n_24428, n_24429, n_24430, n_24431;
wire n_24415, n_24416, n_24417, n_24418, n_24419, n_24420, n_24421, n_24422;
wire n_24404, n_24405, n_24407, n_24409, n_24410, n_24411, n_24412, n_24413;
wire n_24395, n_24396, n_24397, n_24398, n_24399, n_24400, n_24401, n_24402;
wire n_24386, n_24387, n_24388, n_24389, n_24390, n_24391, n_24393, n_24394;
wire n_24378, n_24379, n_24380, n_24381, n_24382, n_24383, n_24384, n_24385;
wire n_24369, n_24370, n_24372, n_24373, n_24374, n_24375, n_24376, n_24377;
wire n_24361, n_24362, n_24363, n_24364, n_24365, n_24366, n_24367, n_24368;
wire n_24351, n_24352, n_24353, n_24354, n_24357, n_24358, n_24359, n_24360;
wire n_24343, n_24344, n_24345, n_24346, n_24347, n_24348, n_24349, n_24350;
wire n_24335, n_24336, n_24337, n_24338, n_24339, n_24340, n_24341, n_24342;
wire n_24325, n_24326, n_24329, n_24330, n_24331, n_24332, n_24333, n_24334;
wire n_24311, n_24312, n_24313, n_24314, n_24318, n_24321, n_24323, n_24324;
wire n_24302, n_24303, n_24304, n_24305, n_24306, n_24307, n_24308, n_24309;
wire n_24294, n_24295, n_24296, n_24297, n_24298, n_24299, n_24300, n_24301;
wire n_24286, n_24287, n_24288, n_24289, n_24290, n_24291, n_24292, n_24293;
wire n_24278, n_24279, n_24280, n_24281, n_24282, n_24283, n_24284, n_24285;
wire n_24270, n_24271, n_24272, n_24273, n_24274, n_24275, n_24276, n_24277;
wire n_24262, n_24263, n_24264, n_24265, n_24266, n_24267, n_24268, n_24269;
wire n_24252, n_24254, n_24255, n_24257, n_24258, n_24259, n_24260, n_24261;
wire n_24243, n_24245, n_24246, n_24247, n_24248, n_24249, n_24250, n_24251;
wire n_24234, n_24235, n_24237, n_24238, n_24239, n_24240, n_24241, n_24242;
wire n_24225, n_24226, n_24227, n_24228, n_24229, n_24230, n_24232, n_24233;
wire n_24216, n_24217, n_24219, n_24220, n_24221, n_24222, n_24223, n_24224;
wire n_24207, n_24208, n_24209, n_24210, n_24211, n_24213, n_24214, n_24215;
wire n_24197, n_24198, n_24199, n_24200, n_24202, n_24204, n_24205, n_24206;
wire n_24188, n_24189, n_24190, n_24191, n_24192, n_24194, n_24195, n_24196;
wire n_24177, n_24178, n_24179, n_24182, n_24184, n_24185, n_24186, n_24187;
wire n_24167, n_24168, n_24169, n_24170, n_24172, n_24173, n_24174, n_24175;
wire n_24159, n_24160, n_24161, n_24162, n_24163, n_24164, n_24165, n_24166;
wire n_24151, n_24152, n_24153, n_24154, n_24155, n_24156, n_24157, n_24158;
wire n_24143, n_24144, n_24145, n_24146, n_24147, n_24148, n_24149, n_24150;
wire n_24135, n_24136, n_24137, n_24138, n_24139, n_24140, n_24141, n_24142;
wire n_24126, n_24127, n_24128, n_24129, n_24130, n_24131, n_24133, n_24134;
wire n_24117, n_24118, n_24120, n_24121, n_24122, n_24123, n_24124, n_24125;
wire n_24108, n_24109, n_24110, n_24111, n_24112, n_24113, n_24114, n_24116;
wire n_24100, n_24101, n_24102, n_24103, n_24104, n_24105, n_24106, n_24107;
wire n_24091, n_24092, n_24093, n_24094, n_24095, n_24096, n_24098, n_24099;
wire n_24082, n_24083, n_24084, n_24085, n_24086, n_24088, n_24089, n_24090;
wire n_24074, n_24075, n_24076, n_24077, n_24078, n_24079, n_24080, n_24081;
wire n_24065, n_24067, n_24068, n_24069, n_24070, n_24071, n_24072, n_24073;
wire n_24054, n_24055, n_24056, n_24057, n_24059, n_24060, n_24062, n_24063;
wire n_24046, n_24047, n_24048, n_24049, n_24050, n_24051, n_24052, n_24053;
wire n_24038, n_24039, n_24040, n_24041, n_24042, n_24043, n_24044, n_24045;
wire n_24030, n_24031, n_24032, n_24033, n_24034, n_24035, n_24036, n_24037;
wire n_24021, n_24022, n_24023, n_24024, n_24025, n_24027, n_24028, n_24029;
wire n_24013, n_24014, n_24015, n_24016, n_24017, n_24018, n_24019, n_24020;
wire n_24003, n_24005, n_24006, n_24007, n_24008, n_24009, n_24011, n_24012;
wire n_23995, n_23996, n_23997, n_23998, n_23999, n_24000, n_24001, n_24002;
wire n_23986, n_23987, n_23988, n_23989, n_23990, n_23991, n_23992, n_23993;
wire n_23977, n_23978, n_23980, n_23981, n_23982, n_23983, n_23984, n_23985;
wire n_23969, n_23970, n_23971, n_23972, n_23973, n_23974, n_23975, n_23976;
wire n_23958, n_23960, n_23963, n_23964, n_23965, n_23966, n_23967, n_23968;
wire n_23950, n_23951, n_23952, n_23953, n_23954, n_23955, n_23956, n_23957;
wire n_23940, n_23941, n_23943, n_23944, n_23946, n_23947, n_23948, n_23949;
wire n_23931, n_23932, n_23933, n_23934, n_23935, n_23936, n_23937, n_23939;
wire n_23922, n_23923, n_23924, n_23925, n_23926, n_23927, n_23929, n_23930;
wire n_23911, n_23912, n_23913, n_23914, n_23918, n_23919, n_23920, n_23921;
wire n_23901, n_23902, n_23903, n_23904, n_23905, n_23907, n_23909, n_23910;
wire n_23892, n_23893, n_23894, n_23896, n_23897, n_23898, n_23899, n_23900;
wire n_23884, n_23885, n_23886, n_23887, n_23888, n_23889, n_23890, n_23891;
wire n_23875, n_23876, n_23878, n_23879, n_23880, n_23881, n_23882, n_23883;
wire n_23867, n_23868, n_23869, n_23870, n_23871, n_23872, n_23873, n_23874;
wire n_23859, n_23860, n_23861, n_23862, n_23863, n_23864, n_23865, n_23866;
wire n_23850, n_23851, n_23852, n_23853, n_23854, n_23855, n_23856, n_23858;
wire n_23839, n_23840, n_23843, n_23844, n_23846, n_23847, n_23848, n_23849;
wire n_23830, n_23831, n_23832, n_23834, n_23835, n_23836, n_23837, n_23838;
wire n_23822, n_23823, n_23824, n_23825, n_23826, n_23827, n_23828, n_23829;
wire n_23813, n_23814, n_23816, n_23817, n_23818, n_23819, n_23820, n_23821;
wire n_23805, n_23806, n_23807, n_23808, n_23809, n_23810, n_23811, n_23812;
wire n_23797, n_23798, n_23799, n_23800, n_23801, n_23802, n_23803, n_23804;
wire n_23788, n_23790, n_23791, n_23792, n_23793, n_23794, n_23795, n_23796;
wire n_23779, n_23780, n_23781, n_23782, n_23783, n_23784, n_23785, n_23786;
wire n_23771, n_23772, n_23773, n_23774, n_23775, n_23776, n_23777, n_23778;
wire n_23762, n_23763, n_23764, n_23765, n_23767, n_23768, n_23769, n_23770;
wire n_23754, n_23755, n_23756, n_23757, n_23758, n_23759, n_23760, n_23761;
wire n_23745, n_23746, n_23747, n_23748, n_23749, n_23750, n_23751, n_23752;
wire n_23736, n_23737, n_23738, n_23739, n_23740, n_23742, n_23743, n_23744;
wire n_23728, n_23729, n_23730, n_23731, n_23732, n_23733, n_23734, n_23735;
wire n_23720, n_23721, n_23722, n_23723, n_23724, n_23725, n_23726, n_23727;
wire n_23711, n_23713, n_23714, n_23715, n_23716, n_23717, n_23718, n_23719;
wire n_23702, n_23703, n_23704, n_23705, n_23706, n_23708, n_23709, n_23710;
wire n_23694, n_23695, n_23696, n_23697, n_23698, n_23699, n_23700, n_23701;
wire n_23686, n_23687, n_23688, n_23689, n_23690, n_23691, n_23692, n_23693;
wire n_23678, n_23679, n_23680, n_23681, n_23682, n_23683, n_23684, n_23685;
wire n_23667, n_23668, n_23669, n_23670, n_23672, n_23674, n_23676, n_23677;
wire n_23659, n_23660, n_23661, n_23662, n_23663, n_23664, n_23665, n_23666;
wire n_23649, n_23650, n_23651, n_23652, n_23655, n_23656, n_23657, n_23658;
wire n_23640, n_23641, n_23642, n_23643, n_23644, n_23645, n_23647, n_23648;
wire n_23632, n_23633, n_23634, n_23635, n_23636, n_23637, n_23638, n_23639;
wire n_23623, n_23624, n_23625, n_23626, n_23627, n_23628, n_23629, n_23630;
wire n_23615, n_23616, n_23617, n_23618, n_23619, n_23620, n_23621, n_23622;
wire n_23606, n_23607, n_23609, n_23610, n_23611, n_23612, n_23613, n_23614;
wire n_23597, n_23598, n_23599, n_23600, n_23602, n_23603, n_23604, n_23605;
wire n_23588, n_23589, n_23590, n_23591, n_23592, n_23593, n_23594, n_23596;
wire n_23579, n_23580, n_23581, n_23582, n_23584, n_23585, n_23586, n_23587;
wire n_23571, n_23572, n_23573, n_23574, n_23575, n_23576, n_23577, n_23578;
wire n_23562, n_23563, n_23564, n_23565, n_23566, n_23567, n_23568, n_23569;
wire n_23554, n_23555, n_23556, n_23557, n_23558, n_23559, n_23560, n_23561;
wire n_23543, n_23544, n_23545, n_23546, n_23548, n_23550, n_23551, n_23552;
wire n_23533, n_23534, n_23535, n_23536, n_23538, n_23539, n_23541, n_23542;
wire n_23523, n_23524, n_23526, n_23527, n_23528, n_23530, n_23531, n_23532;
wire n_23514, n_23515, n_23517, n_23518, n_23519, n_23520, n_23521, n_23522;
wire n_23505, n_23506, n_23507, n_23509, n_23510, n_23511, n_23512, n_23513;
wire n_23496, n_23497, n_23498, n_23499, n_23500, n_23501, n_23502, n_23504;
wire n_23487, n_23488, n_23489, n_23490, n_23491, n_23493, n_23494, n_23495;
wire n_23477, n_23478, n_23480, n_23481, n_23483, n_23484, n_23485, n_23486;
wire n_23468, n_23470, n_23471, n_23472, n_23473, n_23474, n_23475, n_23476;
wire n_23460, n_23461, n_23462, n_23463, n_23464, n_23465, n_23466, n_23467;
wire n_23452, n_23453, n_23454, n_23455, n_23456, n_23457, n_23458, n_23459;
wire n_23444, n_23445, n_23446, n_23447, n_23448, n_23449, n_23450, n_23451;
wire n_23436, n_23437, n_23438, n_23439, n_23440, n_23441, n_23442, n_23443;
wire n_23428, n_23429, n_23430, n_23431, n_23432, n_23433, n_23434, n_23435;
wire n_23420, n_23421, n_23422, n_23423, n_23424, n_23425, n_23426, n_23427;
wire n_23412, n_23413, n_23414, n_23415, n_23416, n_23417, n_23418, n_23419;
wire n_23404, n_23405, n_23406, n_23407, n_23408, n_23409, n_23410, n_23411;
wire n_23396, n_23397, n_23398, n_23399, n_23400, n_23401, n_23402, n_23403;
wire n_23385, n_23386, n_23387, n_23389, n_23390, n_23392, n_23393, n_23395;
wire n_23377, n_23378, n_23379, n_23380, n_23381, n_23382, n_23383, n_23384;
wire n_23367, n_23368, n_23369, n_23370, n_23371, n_23372, n_23373, n_23376;
wire n_23358, n_23359, n_23360, n_23361, n_23363, n_23364, n_23365, n_23366;
wire n_23347, n_23348, n_23349, n_23350, n_23351, n_23355, n_23356, n_23357;
wire n_23339, n_23340, n_23341, n_23342, n_23343, n_23344, n_23345, n_23346;
wire n_23330, n_23331, n_23332, n_23333, n_23334, n_23335, n_23337, n_23338;
wire n_23322, n_23323, n_23324, n_23325, n_23326, n_23327, n_23328, n_23329;
wire n_23312, n_23313, n_23314, n_23315, n_23317, n_23318, n_23319, n_23321;
wire n_23303, n_23304, n_23305, n_23306, n_23308, n_23309, n_23310, n_23311;
wire n_23295, n_23296, n_23297, n_23298, n_23299, n_23300, n_23301, n_23302;
wire n_23286, n_23287, n_23288, n_23290, n_23291, n_23292, n_23293, n_23294;
wire n_23278, n_23279, n_23280, n_23281, n_23282, n_23283, n_23284, n_23285;
wire n_23269, n_23270, n_23271, n_23272, n_23273, n_23274, n_23275, n_23277;
wire n_23259, n_23260, n_23261, n_23262, n_23263, n_23264, n_23266, n_23267;
wire n_23251, n_23252, n_23253, n_23254, n_23255, n_23256, n_23257, n_23258;
wire n_23243, n_23244, n_23245, n_23246, n_23247, n_23248, n_23249, n_23250;
wire n_23235, n_23236, n_23237, n_23238, n_23239, n_23240, n_23241, n_23242;
wire n_23227, n_23228, n_23229, n_23230, n_23231, n_23232, n_23233, n_23234;
wire n_23218, n_23219, n_23220, n_23222, n_23223, n_23224, n_23225, n_23226;
wire n_23210, n_23211, n_23212, n_23213, n_23214, n_23215, n_23216, n_23217;
wire n_23201, n_23202, n_23203, n_23204, n_23205, n_23206, n_23207, n_23208;
wire n_23191, n_23192, n_23193, n_23195, n_23196, n_23198, n_23199, n_23200;
wire n_23183, n_23184, n_23185, n_23186, n_23187, n_23188, n_23189, n_23190;
wire n_23175, n_23176, n_23177, n_23178, n_23179, n_23180, n_23181, n_23182;
wire n_23167, n_23168, n_23169, n_23170, n_23171, n_23172, n_23173, n_23174;
wire n_23158, n_23159, n_23160, n_23161, n_23162, n_23164, n_23165, n_23166;
wire n_23150, n_23151, n_23152, n_23153, n_23154, n_23155, n_23156, n_23157;
wire n_23141, n_23142, n_23143, n_23145, n_23146, n_23147, n_23148, n_23149;
wire n_23131, n_23132, n_23133, n_23135, n_23136, n_23137, n_23138, n_23139;
wire n_23120, n_23121, n_23123, n_23124, n_23125, n_23128, n_23129, n_23130;
wire n_23111, n_23112, n_23113, n_23114, n_23115, n_23116, n_23117, n_23119;
wire n_23100, n_23101, n_23102, n_23103, n_23104, n_23108, n_23109, n_23110;
wire n_23092, n_23093, n_23094, n_23095, n_23096, n_23097, n_23098, n_23099;
wire n_23084, n_23085, n_23086, n_23087, n_23088, n_23089, n_23090, n_23091;
wire n_23075, n_23076, n_23077, n_23079, n_23080, n_23081, n_23082, n_23083;
wire n_23067, n_23068, n_23069, n_23070, n_23071, n_23072, n_23073, n_23074;
wire n_23059, n_23060, n_23061, n_23062, n_23063, n_23064, n_23065, n_23066;
wire n_23051, n_23052, n_23053, n_23054, n_23055, n_23056, n_23057, n_23058;
wire n_23042, n_23043, n_23044, n_23045, n_23046, n_23047, n_23049, n_23050;
wire n_23034, n_23035, n_23036, n_23037, n_23038, n_23039, n_23040, n_23041;
wire n_23026, n_23027, n_23028, n_23029, n_23030, n_23031, n_23032, n_23033;
wire n_23016, n_23017, n_23018, n_23019, n_23020, n_23022, n_23023, n_23024;
wire n_23007, n_23008, n_23009, n_23010, n_23011, n_23012, n_23013, n_23014;
wire n_22999, n_23000, n_23001, n_23002, n_23003, n_23004, n_23005, n_23006;
wire n_22991, n_22992, n_22993, n_22994, n_22995, n_22996, n_22997, n_22998;
wire n_22981, n_22982, n_22985, n_22986, n_22987, n_22988, n_22989, n_22990;
wire n_22972, n_22973, n_22974, n_22976, n_22977, n_22978, n_22979, n_22980;
wire n_22963, n_22964, n_22965, n_22966, n_22967, n_22969, n_22970, n_22971;
wire n_22955, n_22956, n_22957, n_22958, n_22959, n_22960, n_22961, n_22962;
wire n_22947, n_22948, n_22949, n_22950, n_22951, n_22952, n_22953, n_22954;
wire n_22939, n_22940, n_22941, n_22942, n_22943, n_22944, n_22945, n_22946;
wire n_22931, n_22932, n_22933, n_22934, n_22935, n_22936, n_22937, n_22938;
wire n_22922, n_22924, n_22925, n_22926, n_22927, n_22928, n_22929, n_22930;
wire n_22914, n_22915, n_22916, n_22917, n_22918, n_22919, n_22920, n_22921;
wire n_22906, n_22907, n_22908, n_22909, n_22910, n_22911, n_22912, n_22913;
wire n_22898, n_22899, n_22900, n_22901, n_22902, n_22903, n_22904, n_22905;
wire n_22886, n_22887, n_22888, n_22889, n_22894, n_22895, n_22896, n_22897;
wire n_22875, n_22876, n_22877, n_22878, n_22879, n_22880, n_22883, n_22884;
wire n_22866, n_22867, n_22868, n_22869, n_22870, n_22871, n_22873, n_22874;
wire n_22857, n_22858, n_22859, n_22861, n_22862, n_22863, n_22864, n_22865;
wire n_22849, n_22850, n_22851, n_22852, n_22853, n_22854, n_22855, n_22856;
wire n_22840, n_22841, n_22842, n_22843, n_22844, n_22845, n_22846, n_22848;
wire n_22831, n_22832, n_22833, n_22835, n_22836, n_22837, n_22838, n_22839;
wire n_22820, n_22821, n_22822, n_22823, n_22825, n_22826, n_22828, n_22829;
wire n_22810, n_22811, n_22812, n_22813, n_22814, n_22815, n_22818, n_22819;
wire n_22802, n_22803, n_22804, n_22805, n_22806, n_22807, n_22808, n_22809;
wire n_22793, n_22794, n_22795, n_22796, n_22797, n_22798, n_22800, n_22801;
wire n_22785, n_22786, n_22787, n_22788, n_22789, n_22790, n_22791, n_22792;
wire n_22777, n_22778, n_22779, n_22780, n_22781, n_22782, n_22783, n_22784;
wire n_22769, n_22770, n_22771, n_22772, n_22773, n_22774, n_22775, n_22776;
wire n_22760, n_22761, n_22762, n_22763, n_22764, n_22765, n_22766, n_22768;
wire n_22751, n_22752, n_22753, n_22754, n_22756, n_22757, n_22758, n_22759;
wire n_22741, n_22743, n_22745, n_22746, n_22747, n_22748, n_22749, n_22750;
wire n_22731, n_22733, n_22734, n_22735, n_22736, n_22737, n_22738, n_22740;
wire n_22723, n_22724, n_22725, n_22726, n_22727, n_22728, n_22729, n_22730;
wire n_22715, n_22716, n_22717, n_22718, n_22719, n_22720, n_22721, n_22722;
wire n_22706, n_22708, n_22709, n_22710, n_22711, n_22712, n_22713, n_22714;
wire n_22697, n_22698, n_22700, n_22701, n_22702, n_22703, n_22704, n_22705;
wire n_22687, n_22688, n_22689, n_22690, n_22691, n_22692, n_22694, n_22696;
wire n_22677, n_22678, n_22679, n_22680, n_22681, n_22682, n_22683, n_22685;
wire n_22669, n_22670, n_22671, n_22672, n_22673, n_22674, n_22675, n_22676;
wire n_22660, n_22661, n_22662, n_22663, n_22664, n_22666, n_22667, n_22668;
wire n_22651, n_22652, n_22653, n_22654, n_22656, n_22657, n_22658, n_22659;
wire n_22642, n_22643, n_22644, n_22645, n_22646, n_22647, n_22648, n_22650;
wire n_22630, n_22631, n_22632, n_22634, n_22635, n_22637, n_22638, n_22641;
wire n_22622, n_22623, n_22624, n_22625, n_22626, n_22627, n_22628, n_22629;
wire n_22613, n_22614, n_22615, n_22616, n_22617, n_22618, n_22619, n_22620;
wire n_22604, n_22605, n_22607, n_22608, n_22609, n_22610, n_22611, n_22612;
wire n_22596, n_22597, n_22598, n_22599, n_22600, n_22601, n_22602, n_22603;
wire n_22587, n_22588, n_22589, n_22591, n_22592, n_22593, n_22594, n_22595;
wire n_22577, n_22578, n_22579, n_22580, n_22581, n_22584, n_22585, n_22586;
wire n_22565, n_22567, n_22569, n_22571, n_22572, n_22573, n_22575, n_22576;
wire n_22557, n_22558, n_22559, n_22560, n_22561, n_22562, n_22563, n_22564;
wire n_22548, n_22549, n_22550, n_22551, n_22552, n_22554, n_22555, n_22556;
wire n_22539, n_22540, n_22541, n_22542, n_22543, n_22544, n_22545, n_22546;
wire n_22530, n_22532, n_22533, n_22534, n_22535, n_22536, n_22537, n_22538;
wire n_22522, n_22523, n_22524, n_22525, n_22526, n_22527, n_22528, n_22529;
wire n_22514, n_22515, n_22516, n_22517, n_22518, n_22519, n_22520, n_22521;
wire n_22506, n_22507, n_22508, n_22509, n_22510, n_22511, n_22512, n_22513;
wire n_22498, n_22499, n_22500, n_22501, n_22502, n_22503, n_22504, n_22505;
wire n_22487, n_22488, n_22489, n_22490, n_22491, n_22492, n_22494, n_22497;
wire n_22478, n_22479, n_22480, n_22481, n_22482, n_22483, n_22484, n_22485;
wire n_22470, n_22471, n_22472, n_22473, n_22474, n_22475, n_22476, n_22477;
wire n_22462, n_22463, n_22464, n_22465, n_22466, n_22467, n_22468, n_22469;
wire n_22454, n_22455, n_22456, n_22457, n_22458, n_22459, n_22460, n_22461;
wire n_22445, n_22446, n_22447, n_22448, n_22449, n_22450, n_22451, n_22453;
wire n_22436, n_22437, n_22438, n_22440, n_22441, n_22442, n_22443, n_22444;
wire n_22425, n_22428, n_22429, n_22430, n_22431, n_22432, n_22434, n_22435;
wire n_22417, n_22418, n_22419, n_22420, n_22421, n_22422, n_22423, n_22424;
wire n_22409, n_22410, n_22411, n_22412, n_22413, n_22414, n_22415, n_22416;
wire n_22401, n_22402, n_22403, n_22404, n_22405, n_22406, n_22407, n_22408;
wire n_22389, n_22390, n_22392, n_22395, n_22396, n_22397, n_22399, n_22400;
wire n_22381, n_22382, n_22383, n_22384, n_22385, n_22386, n_22387, n_22388;
wire n_22373, n_22374, n_22375, n_22376, n_22377, n_22378, n_22379, n_22380;
wire n_22365, n_22366, n_22367, n_22368, n_22369, n_22370, n_22371, n_22372;
wire n_22356, n_22357, n_22358, n_22359, n_22361, n_22362, n_22363, n_22364;
wire n_22348, n_22349, n_22350, n_22351, n_22352, n_22353, n_22354, n_22355;
wire n_22339, n_22340, n_22341, n_22342, n_22344, n_22345, n_22346, n_22347;
wire n_22328, n_22329, n_22330, n_22332, n_22333, n_22335, n_22336, n_22338;
wire n_22319, n_22320, n_22322, n_22323, n_22324, n_22325, n_22326, n_22327;
wire n_22310, n_22311, n_22312, n_22313, n_22314, n_22315, n_22316, n_22318;
wire n_22302, n_22303, n_22304, n_22305, n_22306, n_22307, n_22308, n_22309;
wire n_22292, n_22293, n_22294, n_22295, n_22296, n_22297, n_22300, n_22301;
wire n_22283, n_22284, n_22286, n_22287, n_22288, n_22289, n_22290, n_22291;
wire n_22272, n_22273, n_22274, n_22275, n_22276, n_22277, n_22278, n_22279;
wire n_22264, n_22265, n_22266, n_22267, n_22268, n_22269, n_22270, n_22271;
wire n_22255, n_22256, n_22257, n_22258, n_22259, n_22260, n_22262, n_22263;
wire n_22246, n_22247, n_22248, n_22249, n_22250, n_22251, n_22252, n_22254;
wire n_22238, n_22239, n_22240, n_22241, n_22242, n_22243, n_22244, n_22245;
wire n_22229, n_22230, n_22231, n_22232, n_22233, n_22234, n_22236, n_22237;
wire n_22220, n_22221, n_22222, n_22223, n_22224, n_22225, n_22226, n_22228;
wire n_22211, n_22212, n_22213, n_22214, n_22215, n_22216, n_22218, n_22219;
wire n_22202, n_22203, n_22204, n_22205, n_22206, n_22207, n_22208, n_22210;
wire n_22194, n_22195, n_22196, n_22197, n_22198, n_22199, n_22200, n_22201;
wire n_22186, n_22187, n_22188, n_22189, n_22190, n_22191, n_22192, n_22193;
wire n_22176, n_22177, n_22179, n_22180, n_22181, n_22182, n_22183, n_22184;
wire n_22164, n_22165, n_22166, n_22167, n_22168, n_22169, n_22170, n_22171;
wire n_22155, n_22156, n_22157, n_22158, n_22160, n_22161, n_22162, n_22163;
wire n_22146, n_22147, n_22148, n_22149, n_22150, n_22152, n_22153, n_22154;
wire n_22137, n_22139, n_22140, n_22141, n_22142, n_22143, n_22144, n_22145;
wire n_22129, n_22130, n_22131, n_22132, n_22133, n_22134, n_22135, n_22136;
wire n_22115, n_22117, n_22119, n_22121, n_22122, n_22123, n_22124, n_22128;
wire n_22106, n_22107, n_22108, n_22109, n_22110, n_22111, n_22113, n_22114;
wire n_22098, n_22099, n_22100, n_22101, n_22102, n_22103, n_22104, n_22105;
wire n_22090, n_22091, n_22092, n_22093, n_22094, n_22095, n_22096, n_22097;
wire n_22082, n_22083, n_22084, n_22085, n_22086, n_22087, n_22088, n_22089;
wire n_22074, n_22075, n_22076, n_22077, n_22078, n_22079, n_22080, n_22081;
wire n_22065, n_22066, n_22067, n_22068, n_22070, n_22071, n_22072, n_22073;
wire n_22056, n_22057, n_22058, n_22059, n_22061, n_22062, n_22063, n_22064;
wire n_22047, n_22048, n_22049, n_22050, n_22051, n_22052, n_22053, n_22054;
wire n_22038, n_22039, n_22041, n_22042, n_22043, n_22044, n_22045, n_22046;
wire n_22030, n_22031, n_22032, n_22033, n_22034, n_22035, n_22036, n_22037;
wire n_22022, n_22023, n_22024, n_22025, n_22026, n_22027, n_22028, n_22029;
wire n_22012, n_22013, n_22015, n_22016, n_22017, n_22018, n_22020, n_22021;
wire n_22002, n_22003, n_22004, n_22005, n_22006, n_22008, n_22010, n_22011;
wire n_21993, n_21995, n_21996, n_21997, n_21998, n_21999, n_22000, n_22001;
wire n_21984, n_21985, n_21986, n_21987, n_21988, n_21989, n_21990, n_21992;
wire n_21976, n_21977, n_21978, n_21979, n_21980, n_21981, n_21982, n_21983;
wire n_21968, n_21969, n_21970, n_21971, n_21972, n_21973, n_21974, n_21975;
wire n_21960, n_21961, n_21962, n_21963, n_21964, n_21965, n_21966, n_21967;
wire n_21951, n_21953, n_21954, n_21955, n_21956, n_21957, n_21958, n_21959;
wire n_21943, n_21944, n_21945, n_21946, n_21947, n_21948, n_21949, n_21950;
wire n_21935, n_21936, n_21937, n_21938, n_21939, n_21940, n_21941, n_21942;
wire n_21927, n_21928, n_21929, n_21930, n_21931, n_21932, n_21933, n_21934;
wire n_21919, n_21920, n_21921, n_21922, n_21923, n_21924, n_21925, n_21926;
wire n_21911, n_21912, n_21913, n_21914, n_21915, n_21916, n_21917, n_21918;
wire n_21903, n_21904, n_21905, n_21906, n_21907, n_21908, n_21909, n_21910;
wire n_21895, n_21896, n_21897, n_21898, n_21899, n_21900, n_21901, n_21902;
wire n_21886, n_21887, n_21888, n_21889, n_21890, n_21891, n_21892, n_21894;
wire n_21878, n_21879, n_21880, n_21881, n_21882, n_21883, n_21884, n_21885;
wire n_21870, n_21871, n_21872, n_21873, n_21874, n_21875, n_21876, n_21877;
wire n_21862, n_21863, n_21864, n_21865, n_21866, n_21867, n_21868, n_21869;
wire n_21854, n_21855, n_21856, n_21857, n_21858, n_21859, n_21860, n_21861;
wire n_21846, n_21847, n_21848, n_21849, n_21850, n_21851, n_21852, n_21853;
wire n_21836, n_21837, n_21838, n_21839, n_21841, n_21842, n_21844, n_21845;
wire n_21827, n_21828, n_21829, n_21830, n_21831, n_21832, n_21833, n_21835;
wire n_21819, n_21820, n_21821, n_21822, n_21823, n_21824, n_21825, n_21826;
wire n_21810, n_21811, n_21812, n_21813, n_21814, n_21815, n_21816, n_21818;
wire n_21801, n_21802, n_21803, n_21804, n_21805, n_21806, n_21807, n_21809;
wire n_21790, n_21792, n_21793, n_21794, n_21795, n_21796, n_21797, n_21798;
wire n_21782, n_21783, n_21784, n_21785, n_21786, n_21787, n_21788, n_21789;
wire n_21774, n_21775, n_21776, n_21777, n_21778, n_21779, n_21780, n_21781;
wire n_21766, n_21767, n_21768, n_21769, n_21770, n_21771, n_21772, n_21773;
wire n_21758, n_21759, n_21760, n_21761, n_21762, n_21763, n_21764, n_21765;
wire n_21747, n_21748, n_21749, n_21750, n_21754, n_21755, n_21756, n_21757;
wire n_21739, n_21740, n_21741, n_21742, n_21743, n_21744, n_21745, n_21746;
wire n_21730, n_21731, n_21733, n_21734, n_21735, n_21736, n_21737, n_21738;
wire n_21721, n_21722, n_21723, n_21724, n_21726, n_21727, n_21728, n_21729;
wire n_21709, n_21712, n_21714, n_21715, n_21716, n_21717, n_21718, n_21720;
wire n_21700, n_21701, n_21702, n_21703, n_21704, n_21705, n_21706, n_21708;
wire n_21691, n_21692, n_21693, n_21694, n_21695, n_21696, n_21698, n_21699;
wire n_21677, n_21678, n_21682, n_21683, n_21685, n_21687, n_21689, n_21690;
wire n_21666, n_21667, n_21668, n_21669, n_21671, n_21673, n_21674, n_21675;
wire n_21657, n_21658, n_21660, n_21661, n_21662, n_21663, n_21664, n_21665;
wire n_21649, n_21650, n_21651, n_21652, n_21653, n_21654, n_21655, n_21656;
wire n_21640, n_21641, n_21643, n_21644, n_21645, n_21646, n_21647, n_21648;
wire n_21632, n_21633, n_21634, n_21635, n_21636, n_21637, n_21638, n_21639;
wire n_21624, n_21625, n_21626, n_21627, n_21628, n_21629, n_21630, n_21631;
wire n_21616, n_21617, n_21618, n_21619, n_21620, n_21621, n_21622, n_21623;
wire n_21607, n_21608, n_21609, n_21611, n_21612, n_21613, n_21614, n_21615;
wire n_21598, n_21599, n_21600, n_21601, n_21602, n_21603, n_21604, n_21605;
wire n_21589, n_21590, n_21591, n_21592, n_21593, n_21594, n_21595, n_21596;
wire n_21580, n_21581, n_21582, n_21584, n_21585, n_21586, n_21587, n_21588;
wire n_21572, n_21573, n_21574, n_21575, n_21576, n_21577, n_21578, n_21579;
wire n_21563, n_21564, n_21565, n_21567, n_21568, n_21569, n_21570, n_21571;
wire n_21554, n_21555, n_21556, n_21557, n_21558, n_21559, n_21560, n_21561;
wire n_21545, n_21546, n_21547, n_21548, n_21549, n_21550, n_21551, n_21552;
wire n_21537, n_21538, n_21539, n_21540, n_21541, n_21542, n_21543, n_21544;
wire n_21528, n_21529, n_21530, n_21531, n_21532, n_21533, n_21534, n_21536;
wire n_21520, n_21521, n_21522, n_21523, n_21524, n_21525, n_21526, n_21527;
wire n_21512, n_21513, n_21514, n_21515, n_21516, n_21517, n_21518, n_21519;
wire n_21503, n_21504, n_21505, n_21506, n_21507, n_21508, n_21509, n_21511;
wire n_21493, n_21494, n_21495, n_21496, n_21497, n_21498, n_21501, n_21502;
wire n_21485, n_21486, n_21487, n_21488, n_21489, n_21490, n_21491, n_21492;
wire n_21476, n_21477, n_21478, n_21479, n_21480, n_21482, n_21483, n_21484;
wire n_21466, n_21467, n_21468, n_21469, n_21470, n_21471, n_21472, n_21475;
wire n_21458, n_21459, n_21460, n_21461, n_21462, n_21463, n_21464, n_21465;
wire n_21450, n_21451, n_21452, n_21453, n_21454, n_21455, n_21456, n_21457;
wire n_21442, n_21443, n_21444, n_21445, n_21446, n_21447, n_21448, n_21449;
wire n_21431, n_21432, n_21433, n_21437, n_21438, n_21439, n_21440, n_21441;
wire n_21423, n_21424, n_21425, n_21426, n_21427, n_21428, n_21429, n_21430;
wire n_21413, n_21414, n_21415, n_21416, n_21418, n_21419, n_21421, n_21422;
wire n_21405, n_21406, n_21407, n_21408, n_21409, n_21410, n_21411, n_21412;
wire n_21395, n_21396, n_21397, n_21398, n_21399, n_21402, n_21403, n_21404;
wire n_21387, n_21388, n_21389, n_21390, n_21391, n_21392, n_21393, n_21394;
wire n_21379, n_21380, n_21381, n_21382, n_21383, n_21384, n_21385, n_21386;
wire n_21369, n_21371, n_21373, n_21374, n_21375, n_21376, n_21377, n_21378;
wire n_21361, n_21362, n_21363, n_21364, n_21365, n_21366, n_21367, n_21368;
wire n_21348, n_21349, n_21353, n_21354, n_21355, n_21357, n_21358, n_21360;
wire n_21337, n_21338, n_21341, n_21343, n_21344, n_21345, n_21346, n_21347;
wire n_21329, n_21330, n_21331, n_21332, n_21333, n_21334, n_21335, n_21336;
wire n_21318, n_21320, n_21322, n_21324, n_21325, n_21326, n_21327, n_21328;
wire n_21308, n_21309, n_21310, n_21311, n_21312, n_21313, n_21314, n_21315;
wire n_21299, n_21300, n_21301, n_21302, n_21303, n_21304, n_21306, n_21307;
wire n_21288, n_21289, n_21290, n_21291, n_21293, n_21294, n_21295, n_21297;
wire n_21274, n_21276, n_21278, n_21279, n_21281, n_21282, n_21286, n_21287;
wire n_21265, n_21266, n_21267, n_21268, n_21269, n_21270, n_21271, n_21272;
wire n_21257, n_21258, n_21259, n_21260, n_21261, n_21262, n_21263, n_21264;
wire n_21249, n_21250, n_21251, n_21252, n_21253, n_21254, n_21255, n_21256;
wire n_21241, n_21242, n_21243, n_21244, n_21245, n_21246, n_21247, n_21248;
wire n_21231, n_21232, n_21233, n_21234, n_21235, n_21237, n_21239, n_21240;
wire n_21221, n_21222, n_21223, n_21224, n_21225, n_21227, n_21228, n_21230;
wire n_21210, n_21211, n_21212, n_21214, n_21215, n_21216, n_21217, n_21219;
wire n_21201, n_21202, n_21203, n_21204, n_21205, n_21206, n_21207, n_21208;
wire n_21192, n_21193, n_21194, n_21195, n_21196, n_21197, n_21199, n_21200;
wire n_21184, n_21185, n_21186, n_21187, n_21188, n_21189, n_21190, n_21191;
wire n_21176, n_21177, n_21178, n_21179, n_21180, n_21181, n_21182, n_21183;
wire n_21167, n_21168, n_21169, n_21170, n_21171, n_21172, n_21173, n_21174;
wire n_21157, n_21158, n_21159, n_21160, n_21161, n_21162, n_21164, n_21165;
wire n_21147, n_21148, n_21149, n_21151, n_21152, n_21153, n_21154, n_21156;
wire n_21139, n_21140, n_21141, n_21142, n_21143, n_21144, n_21145, n_21146;
wire n_21131, n_21132, n_21133, n_21134, n_21135, n_21136, n_21137, n_21138;
wire n_21123, n_21124, n_21125, n_21126, n_21127, n_21128, n_21129, n_21130;
wire n_21114, n_21115, n_21116, n_21117, n_21118, n_21120, n_21121, n_21122;
wire n_21106, n_21107, n_21108, n_21109, n_21110, n_21111, n_21112, n_21113;
wire n_21098, n_21099, n_21100, n_21101, n_21102, n_21103, n_21104, n_21105;
wire n_21090, n_21091, n_21092, n_21093, n_21094, n_21095, n_21096, n_21097;
wire n_21081, n_21082, n_21083, n_21084, n_21085, n_21087, n_21088, n_21089;
wire n_21072, n_21073, n_21074, n_21075, n_21076, n_21078, n_21079, n_21080;
wire n_21064, n_21065, n_21066, n_21067, n_21068, n_21069, n_21070, n_21071;
wire n_21054, n_21056, n_21058, n_21059, n_21060, n_21061, n_21062, n_21063;
wire n_21046, n_21047, n_21048, n_21049, n_21050, n_21051, n_21052, n_21053;
wire n_21038, n_21039, n_21040, n_21041, n_21042, n_21043, n_21044, n_21045;
wire n_21029, n_21030, n_21031, n_21032, n_21033, n_21034, n_21036, n_21037;
wire n_21020, n_21021, n_21022, n_21023, n_21024, n_21025, n_21026, n_21027;
wire n_21012, n_21013, n_21014, n_21015, n_21016, n_21017, n_21018, n_21019;
wire n_21004, n_21005, n_21006, n_21007, n_21008, n_21009, n_21010, n_21011;
wire n_20995, n_20996, n_20998, n_20999, n_21000, n_21001, n_21002, n_21003;
wire n_20985, n_20986, n_20987, n_20988, n_20989, n_20990, n_20992, n_20993;
wire n_20977, n_20978, n_20979, n_20980, n_20981, n_20982, n_20983, n_20984;
wire n_20969, n_20970, n_20971, n_20972, n_20973, n_20974, n_20975, n_20976;
wire n_20960, n_20961, n_20962, n_20964, n_20965, n_20966, n_20967, n_20968;
wire n_20951, n_20953, n_20954, n_20955, n_20956, n_20957, n_20958, n_20959;
wire n_20938, n_20940, n_20944, n_20945, n_20946, n_20947, n_20948, n_20950;
wire n_20929, n_20930, n_20931, n_20932, n_20933, n_20934, n_20935, n_20937;
wire n_20921, n_20922, n_20923, n_20924, n_20925, n_20926, n_20927, n_20928;
wire n_20913, n_20914, n_20915, n_20916, n_20917, n_20918, n_20919, n_20920;
wire n_20899, n_20901, n_20902, n_20904, n_20906, n_20908, n_20909, n_20912;
wire n_20889, n_20890, n_20891, n_20892, n_20893, n_20894, n_20895, n_20898;
wire n_20879, n_20880, n_20882, n_20883, n_20884, n_20886, n_20887, n_20888;
wire n_20867, n_20868, n_20871, n_20872, n_20874, n_20875, n_20876, n_20877;
wire n_20858, n_20859, n_20861, n_20862, n_20863, n_20864, n_20865, n_20866;
wire n_20850, n_20851, n_20852, n_20853, n_20854, n_20855, n_20856, n_20857;
wire n_20838, n_20839, n_20840, n_20843, n_20844, n_20845, n_20847, n_20848;
wire n_20830, n_20831, n_20832, n_20833, n_20834, n_20835, n_20836, n_20837;
wire n_20818, n_20819, n_20822, n_20823, n_20825, n_20826, n_20827, n_20829;
wire n_20809, n_20810, n_20812, n_20813, n_20814, n_20815, n_20816, n_20817;
wire n_20796, n_20797, n_20798, n_20802, n_20803, n_20804, n_20805, n_20808;
wire n_20785, n_20787, n_20788, n_20790, n_20791, n_20792, n_20794, n_20795;
wire n_20775, n_20776, n_20777, n_20778, n_20781, n_20782, n_20783, n_20784;
wire n_20766, n_20767, n_20769, n_20770, n_20771, n_20772, n_20773, n_20774;
wire n_20757, n_20759, n_20760, n_20761, n_20762, n_20763, n_20764, n_20765;
wire n_20747, n_20748, n_20749, n_20750, n_20752, n_20754, n_20755, n_20756;
wire n_20736, n_20737, n_20739, n_20740, n_20741, n_20743, n_20744, n_20746;
wire n_20726, n_20727, n_20728, n_20729, n_20730, n_20732, n_20733, n_20734;
wire n_20718, n_20719, n_20720, n_20721, n_20722, n_20723, n_20724, n_20725;
wire n_20710, n_20711, n_20712, n_20713, n_20714, n_20715, n_20716, n_20717;
wire n_20700, n_20701, n_20702, n_20703, n_20704, n_20706, n_20707, n_20708;
wire n_20689, n_20690, n_20692, n_20694, n_20695, n_20697, n_20698, n_20699;
wire n_20679, n_20681, n_20682, n_20683, n_20684, n_20685, n_20687, n_20688;
wire n_20668, n_20670, n_20671, n_20672, n_20673, n_20674, n_20675, n_20676;
wire n_20660, n_20661, n_20662, n_20663, n_20664, n_20665, n_20666, n_20667;
wire n_20650, n_20651, n_20652, n_20655, n_20656, n_20657, n_20658, n_20659;
wire n_20641, n_20642, n_20643, n_20645, n_20646, n_20647, n_20648, n_20649;
wire n_20631, n_20632, n_20633, n_20635, n_20637, n_20638, n_20639, n_20640;
wire n_20622, n_20624, n_20625, n_20626, n_20627, n_20628, n_20629, n_20630;
wire n_20613, n_20614, n_20615, n_20616, n_20618, n_20619, n_20620, n_20621;
wire n_20604, n_20605, n_20606, n_20607, n_20609, n_20610, n_20611, n_20612;
wire n_20596, n_20597, n_20598, n_20599, n_20600, n_20601, n_20602, n_20603;
wire n_20586, n_20588, n_20589, n_20591, n_20592, n_20593, n_20594, n_20595;
wire n_20577, n_20578, n_20579, n_20580, n_20581, n_20582, n_20583, n_20584;
wire n_20569, n_20570, n_20571, n_20572, n_20573, n_20574, n_20575, n_20576;
wire n_20561, n_20562, n_20563, n_20564, n_20565, n_20566, n_20567, n_20568;
wire n_20551, n_20552, n_20554, n_20555, n_20556, n_20557, n_20558, n_20559;
wire n_20543, n_20544, n_20545, n_20546, n_20547, n_20548, n_20549, n_20550;
wire n_20532, n_20535, n_20537, n_20538, n_20539, n_20540, n_20541, n_20542;
wire n_20523, n_20524, n_20525, n_20527, n_20528, n_20529, n_20530, n_20531;
wire n_20515, n_20516, n_20517, n_20518, n_20519, n_20520, n_20521, n_20522;
wire n_20507, n_20508, n_20509, n_20510, n_20511, n_20512, n_20513, n_20514;
wire n_20497, n_20499, n_20500, n_20501, n_20502, n_20503, n_20504, n_20505;
wire n_20488, n_20490, n_20491, n_20492, n_20493, n_20494, n_20495, n_20496;
wire n_20480, n_20481, n_20482, n_20483, n_20484, n_20485, n_20486, n_20487;
wire n_20472, n_20473, n_20474, n_20475, n_20476, n_20477, n_20478, n_20479;
wire n_20464, n_20465, n_20466, n_20467, n_20468, n_20469, n_20470, n_20471;
wire n_20455, n_20456, n_20458, n_20459, n_20460, n_20461, n_20462, n_20463;
wire n_20444, n_20445, n_20446, n_20447, n_20448, n_20450, n_20451, n_20454;
wire n_20436, n_20437, n_20438, n_20439, n_20440, n_20441, n_20442, n_20443;
wire n_20427, n_20428, n_20429, n_20431, n_20432, n_20433, n_20434, n_20435;
wire n_20411, n_20412, n_20414, n_20418, n_20419, n_20422, n_20424, n_20425;
wire n_20402, n_20404, n_20405, n_20406, n_20407, n_20408, n_20409, n_20410;
wire n_20394, n_20395, n_20396, n_20397, n_20398, n_20399, n_20400, n_20401;
wire n_20385, n_20386, n_20387, n_20388, n_20389, n_20390, n_20392, n_20393;
wire n_20377, n_20378, n_20379, n_20380, n_20381, n_20382, n_20383, n_20384;
wire n_20368, n_20370, n_20371, n_20372, n_20373, n_20374, n_20375, n_20376;
wire n_20358, n_20359, n_20360, n_20361, n_20362, n_20363, n_20364, n_20365;
wire n_20347, n_20349, n_20350, n_20352, n_20354, n_20355, n_20356, n_20357;
wire n_20337, n_20338, n_20339, n_20340, n_20341, n_20342, n_20343, n_20346;
wire n_20326, n_20327, n_20328, n_20329, n_20330, n_20332, n_20335, n_20336;
wire n_20316, n_20317, n_20318, n_20319, n_20322, n_20323, n_20324, n_20325;
wire n_20302, n_20303, n_20304, n_20305, n_20307, n_20311, n_20312, n_20315;
wire n_20293, n_20294, n_20295, n_20297, n_20298, n_20299, n_20300, n_20301;
wire n_20284, n_20285, n_20286, n_20287, n_20288, n_20290, n_20291, n_20292;
wire n_20275, n_20277, n_20278, n_20279, n_20280, n_20281, n_20282, n_20283;
wire n_20266, n_20267, n_20268, n_20269, n_20270, n_20271, n_20272, n_20274;
wire n_20255, n_20257, n_20258, n_20261, n_20262, n_20263, n_20264, n_20265;
wire n_20246, n_20247, n_20248, n_20249, n_20250, n_20251, n_20253, n_20254;
wire n_20238, n_20239, n_20240, n_20241, n_20242, n_20243, n_20244, n_20245;
wire n_20230, n_20231, n_20232, n_20233, n_20234, n_20235, n_20236, n_20237;
wire n_20221, n_20223, n_20224, n_20225, n_20226, n_20227, n_20228, n_20229;
wire n_20210, n_20211, n_20212, n_20213, n_20215, n_20217, n_20218, n_20220;
wire n_20200, n_20201, n_20202, n_20203, n_20204, n_20207, n_20208, n_20209;
wire n_20191, n_20193, n_20194, n_20195, n_20196, n_20197, n_20198, n_20199;
wire n_20182, n_20183, n_20184, n_20185, n_20186, n_20187, n_20188, n_20189;
wire n_20172, n_20173, n_20174, n_20175, n_20177, n_20178, n_20179, n_20181;
wire n_20161, n_20163, n_20164, n_20165, n_20167, n_20168, n_20170, n_20171;
wire n_20153, n_20154, n_20155, n_20156, n_20157, n_20158, n_20159, n_20160;
wire n_20144, n_20145, n_20146, n_20147, n_20148, n_20149, n_20150, n_20151;
wire n_20134, n_20135, n_20136, n_20137, n_20138, n_20139, n_20141, n_20143;
wire n_20124, n_20125, n_20127, n_20128, n_20129, n_20130, n_20131, n_20133;
wire n_20116, n_20117, n_20118, n_20119, n_20120, n_20121, n_20122, n_20123;
wire n_20108, n_20109, n_20110, n_20111, n_20112, n_20113, n_20114, n_20115;
wire n_20099, n_20101, n_20102, n_20103, n_20104, n_20105, n_20106, n_20107;
wire n_20091, n_20092, n_20093, n_20094, n_20095, n_20096, n_20097, n_20098;
wire n_20083, n_20084, n_20085, n_20086, n_20087, n_20088, n_20089, n_20090;
wire n_20075, n_20076, n_20077, n_20078, n_20079, n_20080, n_20081, n_20082;
wire n_20067, n_20068, n_20069, n_20070, n_20071, n_20072, n_20073, n_20074;
wire n_20058, n_20059, n_20060, n_20061, n_20062, n_20063, n_20064, n_20065;
wire n_20050, n_20051, n_20052, n_20053, n_20054, n_20055, n_20056, n_20057;
wire n_20041, n_20042, n_20044, n_20045, n_20046, n_20047, n_20048, n_20049;
wire n_20032, n_20033, n_20034, n_20035, n_20036, n_20037, n_20038, n_20040;
wire n_20023, n_20024, n_20025, n_20026, n_20027, n_20028, n_20029, n_20031;
wire n_20015, n_20016, n_20017, n_20018, n_20019, n_20020, n_20021, n_20022;
wire n_20007, n_20008, n_20009, n_20010, n_20011, n_20012, n_20013, n_20014;
wire n_19998, n_19999, n_20000, n_20001, n_20003, n_20004, n_20005, n_20006;
wire n_19989, n_19990, n_19991, n_19992, n_19993, n_19994, n_19995, n_19996;
wire n_19979, n_19980, n_19982, n_19983, n_19984, n_19986, n_19987, n_19988;
wire n_19971, n_19972, n_19973, n_19974, n_19975, n_19976, n_19977, n_19978;
wire n_19962, n_19963, n_19964, n_19965, n_19966, n_19967, n_19968, n_19969;
wire n_19952, n_19953, n_19955, n_19957, n_19958, n_19959, n_19960, n_19961;
wire n_19944, n_19945, n_19946, n_19947, n_19948, n_19949, n_19950, n_19951;
wire n_19936, n_19937, n_19938, n_19939, n_19940, n_19941, n_19942, n_19943;
wire n_19926, n_19928, n_19930, n_19931, n_19932, n_19933, n_19934, n_19935;
wire n_19917, n_19918, n_19919, n_19921, n_19922, n_19923, n_19924, n_19925;
wire n_19909, n_19910, n_19911, n_19912, n_19913, n_19914, n_19915, n_19916;
wire n_19897, n_19898, n_19900, n_19902, n_19903, n_19904, n_19905, n_19906;
wire n_19888, n_19889, n_19890, n_19891, n_19892, n_19893, n_19894, n_19895;
wire n_19880, n_19881, n_19882, n_19883, n_19884, n_19885, n_19886, n_19887;
wire n_19868, n_19870, n_19871, n_19873, n_19874, n_19875, n_19876, n_19878;
wire n_19859, n_19860, n_19861, n_19862, n_19863, n_19864, n_19866, n_19867;
wire n_19849, n_19850, n_19851, n_19852, n_19853, n_19856, n_19857, n_19858;
wire n_19841, n_19842, n_19843, n_19844, n_19845, n_19846, n_19847, n_19848;
wire n_19833, n_19834, n_19835, n_19836, n_19837, n_19838, n_19839, n_19840;
wire n_19821, n_19822, n_19825, n_19827, n_19828, n_19830, n_19831, n_19832;
wire n_19813, n_19814, n_19815, n_19816, n_19817, n_19818, n_19819, n_19820;
wire n_19805, n_19806, n_19807, n_19808, n_19809, n_19810, n_19811, n_19812;
wire n_19797, n_19798, n_19799, n_19800, n_19801, n_19802, n_19803, n_19804;
wire n_19789, n_19790, n_19791, n_19792, n_19793, n_19794, n_19795, n_19796;
wire n_19781, n_19782, n_19783, n_19784, n_19785, n_19786, n_19787, n_19788;
wire n_19772, n_19773, n_19774, n_19776, n_19777, n_19778, n_19779, n_19780;
wire n_19761, n_19763, n_19766, n_19767, n_19768, n_19769, n_19770, n_19771;
wire n_19746, n_19748, n_19750, n_19753, n_19755, n_19757, n_19758, n_19759;
wire n_19737, n_19738, n_19739, n_19740, n_19741, n_19742, n_19743, n_19744;
wire n_19729, n_19730, n_19731, n_19732, n_19733, n_19734, n_19735, n_19736;
wire n_19720, n_19721, n_19722, n_19723, n_19724, n_19725, n_19726, n_19728;
wire n_19709, n_19710, n_19711, n_19712, n_19713, n_19715, n_19717, n_19719;
wire n_19695, n_19696, n_19702, n_19703, n_19704, n_19706, n_19707, n_19708;
wire n_19686, n_19687, n_19688, n_19689, n_19690, n_19691, n_19693, n_19694;
wire n_19678, n_19679, n_19680, n_19681, n_19682, n_19683, n_19684, n_19685;
wire n_19670, n_19671, n_19672, n_19673, n_19674, n_19675, n_19676, n_19677;
wire n_19662, n_19663, n_19664, n_19665, n_19666, n_19667, n_19668, n_19669;
wire n_19652, n_19653, n_19654, n_19655, n_19658, n_19659, n_19660, n_19661;
wire n_19642, n_19643, n_19645, n_19646, n_19647, n_19649, n_19650, n_19651;
wire n_19630, n_19631, n_19632, n_19633, n_19634, n_19637, n_19639, n_19641;
wire n_19621, n_19622, n_19623, n_19624, n_19625, n_19626, n_19627, n_19629;
wire n_19611, n_19613, n_19614, n_19615, n_19616, n_19617, n_19619, n_19620;
wire n_19602, n_19603, n_19604, n_19605, n_19606, n_19607, n_19608, n_19610;
wire n_19591, n_19593, n_19595, n_19596, n_19597, n_19598, n_19600, n_19601;
wire n_19580, n_19581, n_19582, n_19583, n_19584, n_19587, n_19589, n_19590;
wire n_19570, n_19571, n_19572, n_19573, n_19575, n_19576, n_19577, n_19578;
wire n_19562, n_19563, n_19564, n_19565, n_19566, n_19567, n_19568, n_19569;
wire n_19553, n_19554, n_19555, n_19557, n_19558, n_19559, n_19560, n_19561;
wire n_19544, n_19545, n_19546, n_19548, n_19549, n_19550, n_19551, n_19552;
wire n_19536, n_19537, n_19538, n_19539, n_19540, n_19541, n_19542, n_19543;
wire n_19527, n_19528, n_19529, n_19530, n_19531, n_19532, n_19533, n_19534;
wire n_19516, n_19519, n_19520, n_19522, n_19523, n_19524, n_19525, n_19526;
wire n_19504, n_19505, n_19506, n_19507, n_19508, n_19510, n_19511, n_19513;
wire n_19494, n_19495, n_19496, n_19498, n_19500, n_19501, n_19502, n_19503;
wire n_19483, n_19484, n_19485, n_19489, n_19490, n_19491, n_19492, n_19493;
wire n_19475, n_19476, n_19477, n_19478, n_19479, n_19480, n_19481, n_19482;
wire n_19462, n_19463, n_19467, n_19468, n_19469, n_19471, n_19473, n_19474;
wire n_19454, n_19455, n_19456, n_19457, n_19458, n_19459, n_19460, n_19461;
wire n_19443, n_19445, n_19446, n_19447, n_19448, n_19451, n_19452, n_19453;
wire n_19435, n_19436, n_19437, n_19438, n_19439, n_19440, n_19441, n_19442;
wire n_19427, n_19428, n_19429, n_19430, n_19431, n_19432, n_19433, n_19434;
wire n_19419, n_19420, n_19421, n_19422, n_19423, n_19424, n_19425, n_19426;
wire n_19411, n_19412, n_19413, n_19414, n_19415, n_19416, n_19417, n_19418;
wire n_19403, n_19404, n_19405, n_19406, n_19407, n_19408, n_19409, n_19410;
wire n_19390, n_19391, n_19397, n_19398, n_19399, n_19400, n_19401, n_19402;
wire n_19381, n_19382, n_19383, n_19384, n_19385, n_19387, n_19388, n_19389;
wire n_19373, n_19374, n_19375, n_19376, n_19377, n_19378, n_19379, n_19380;
wire n_19365, n_19366, n_19367, n_19368, n_19369, n_19370, n_19371, n_19372;
wire n_19357, n_19358, n_19359, n_19360, n_19361, n_19362, n_19363, n_19364;
wire n_19348, n_19350, n_19351, n_19352, n_19353, n_19354, n_19355, n_19356;
wire n_19339, n_19341, n_19342, n_19343, n_19344, n_19345, n_19346, n_19347;
wire n_19331, n_19332, n_19333, n_19334, n_19335, n_19336, n_19337, n_19338;
wire n_19323, n_19324, n_19325, n_19326, n_19327, n_19328, n_19329, n_19330;
wire n_19313, n_19314, n_19316, n_19318, n_19319, n_19320, n_19321, n_19322;
wire n_19304, n_19305, n_19306, n_19307, n_19308, n_19309, n_19311, n_19312;
wire n_19294, n_19295, n_19296, n_19297, n_19298, n_19299, n_19300, n_19302;
wire n_19282, n_19284, n_19285, n_19286, n_19287, n_19288, n_19290, n_19291;
wire n_19272, n_19273, n_19274, n_19276, n_19277, n_19278, n_19279, n_19280;
wire n_19262, n_19263, n_19264, n_19266, n_19267, n_19268, n_19270, n_19271;
wire n_19252, n_19253, n_19255, n_19256, n_19258, n_19259, n_19260, n_19261;
wire n_19243, n_19244, n_19245, n_19246, n_19247, n_19248, n_19249, n_19250;
wire n_19235, n_19236, n_19237, n_19238, n_19239, n_19240, n_19241, n_19242;
wire n_19227, n_19228, n_19229, n_19230, n_19231, n_19232, n_19233, n_19234;
wire n_19215, n_19217, n_19218, n_19219, n_19220, n_19221, n_19222, n_19225;
wire n_19207, n_19208, n_19209, n_19210, n_19211, n_19212, n_19213, n_19214;
wire n_19198, n_19200, n_19201, n_19202, n_19203, n_19204, n_19205, n_19206;
wire n_19187, n_19189, n_19190, n_19191, n_19192, n_19193, n_19195, n_19196;
wire n_19177, n_19178, n_19179, n_19180, n_19182, n_19183, n_19184, n_19186;
wire n_19168, n_19169, n_19170, n_19171, n_19172, n_19173, n_19174, n_19175;
wire n_19159, n_19160, n_19161, n_19162, n_19164, n_19165, n_19166, n_19167;
wire n_19151, n_19152, n_19153, n_19154, n_19155, n_19156, n_19157, n_19158;
wire n_19142, n_19143, n_19144, n_19146, n_19147, n_19148, n_19149, n_19150;
wire n_19134, n_19135, n_19136, n_19137, n_19138, n_19139, n_19140, n_19141;
wire n_19125, n_19127, n_19128, n_19129, n_19130, n_19131, n_19132, n_19133;
wire n_19116, n_19117, n_19119, n_19120, n_19121, n_19122, n_19123, n_19124;
wire n_19107, n_19108, n_19109, n_19110, n_19111, n_19113, n_19114, n_19115;
wire n_19097, n_19098, n_19099, n_19101, n_19102, n_19103, n_19104, n_19105;
wire n_19085, n_19086, n_19088, n_19090, n_19091, n_19093, n_19094, n_19095;
wire n_19076, n_19077, n_19079, n_19080, n_19081, n_19082, n_19083, n_19084;
wire n_19064, n_19065, n_19068, n_19071, n_19072, n_19073, n_19074, n_19075;
wire n_19056, n_19057, n_19058, n_19059, n_19060, n_19061, n_19062, n_19063;
wire n_19047, n_19048, n_19049, n_19050, n_19051, n_19052, n_19053, n_19055;
wire n_19039, n_19040, n_19041, n_19042, n_19043, n_19044, n_19045, n_19046;
wire n_19030, n_19031, n_19032, n_19033, n_19035, n_19036, n_19037, n_19038;
wire n_19021, n_19022, n_19023, n_19024, n_19026, n_19027, n_19028, n_19029;
wire n_19011, n_19012, n_19013, n_19014, n_19016, n_19017, n_19019, n_19020;
wire n_19001, n_19003, n_19004, n_19005, n_19006, n_19007, n_19008, n_19010;
wire n_18989, n_18993, n_18994, n_18996, n_18997, n_18998, n_18999, n_19000;
wire n_18977, n_18978, n_18979, n_18980, n_18981, n_18982, n_18984, n_18987;
wire n_18964, n_18965, n_18967, n_18968, n_18969, n_18971, n_18974, n_18976;
wire n_18953, n_18954, n_18956, n_18957, n_18958, n_18959, n_18960, n_18961;
wire n_18943, n_18944, n_18945, n_18946, n_18947, n_18948, n_18950, n_18952;
wire n_18935, n_18936, n_18937, n_18938, n_18939, n_18940, n_18941, n_18942;
wire n_18923, n_18924, n_18926, n_18927, n_18929, n_18930, n_18931, n_18933;
wire n_18914, n_18916, n_18917, n_18918, n_18919, n_18920, n_18921, n_18922;
wire n_18904, n_18906, n_18907, n_18908, n_18909, n_18910, n_18911, n_18912;
wire n_18894, n_18895, n_18896, n_18897, n_18898, n_18899, n_18900, n_18902;
wire n_18886, n_18887, n_18888, n_18889, n_18890, n_18891, n_18892, n_18893;
wire n_18877, n_18878, n_18880, n_18881, n_18882, n_18883, n_18884, n_18885;
wire n_18865, n_18868, n_18870, n_18871, n_18872, n_18873, n_18875, n_18876;
wire n_18856, n_18857, n_18858, n_18859, n_18860, n_18861, n_18862, n_18864;
wire n_18848, n_18849, n_18850, n_18851, n_18852, n_18853, n_18854, n_18855;
wire n_18840, n_18841, n_18842, n_18843, n_18844, n_18845, n_18846, n_18847;
wire n_18830, n_18832, n_18833, n_18834, n_18835, n_18836, n_18838, n_18839;
wire n_18819, n_18820, n_18821, n_18823, n_18824, n_18826, n_18828, n_18829;
wire n_18809, n_18810, n_18811, n_18812, n_18813, n_18814, n_18815, n_18816;
wire n_18801, n_18802, n_18803, n_18804, n_18805, n_18806, n_18807, n_18808;
wire n_18791, n_18792, n_18793, n_18794, n_18795, n_18798, n_18799, n_18800;
wire n_18781, n_18782, n_18784, n_18786, n_18787, n_18788, n_18789, n_18790;
wire n_18771, n_18772, n_18773, n_18774, n_18775, n_18776, n_18778, n_18779;
wire n_18763, n_18764, n_18765, n_18766, n_18767, n_18768, n_18769, n_18770;
wire n_18754, n_18755, n_18756, n_18757, n_18758, n_18759, n_18760, n_18761;
wire n_18745, n_18746, n_18747, n_18748, n_18749, n_18750, n_18751, n_18753;
wire n_18735, n_18736, n_18737, n_18738, n_18739, n_18742, n_18743, n_18744;
wire n_18724, n_18726, n_18727, n_18728, n_18729, n_18730, n_18732, n_18734;
wire n_18713, n_18714, n_18715, n_18716, n_18717, n_18720, n_18721, n_18722;
wire n_18704, n_18705, n_18706, n_18708, n_18709, n_18710, n_18711, n_18712;
wire n_18695, n_18696, n_18697, n_18698, n_18700, n_18701, n_18702, n_18703;
wire n_18684, n_18685, n_18687, n_18689, n_18690, n_18691, n_18692, n_18694;
wire n_18675, n_18676, n_18677, n_18679, n_18680, n_18681, n_18682, n_18683;
wire n_18666, n_18667, n_18668, n_18669, n_18670, n_18671, n_18672, n_18674;
wire n_18655, n_18656, n_18658, n_18659, n_18660, n_18661, n_18662, n_18663;
wire n_18643, n_18644, n_18645, n_18646, n_18648, n_18650, n_18652, n_18653;
wire n_18635, n_18636, n_18637, n_18638, n_18639, n_18640, n_18641, n_18642;
wire n_18625, n_18626, n_18627, n_18628, n_18631, n_18632, n_18633, n_18634;
wire n_18616, n_18617, n_18618, n_18619, n_18620, n_18621, n_18622, n_18623;
wire n_18608, n_18609, n_18610, n_18611, n_18612, n_18613, n_18614, n_18615;
wire n_18600, n_18601, n_18602, n_18603, n_18604, n_18605, n_18606, n_18607;
wire n_18591, n_18592, n_18593, n_18594, n_18595, n_18596, n_18597, n_18599;
wire n_18583, n_18584, n_18585, n_18586, n_18587, n_18588, n_18589, n_18590;
wire n_18575, n_18576, n_18577, n_18578, n_18579, n_18580, n_18581, n_18582;
wire n_18564, n_18565, n_18567, n_18568, n_18569, n_18572, n_18573, n_18574;
wire n_18553, n_18554, n_18557, n_18559, n_18560, n_18561, n_18562, n_18563;
wire n_18536, n_18541, n_18542, n_18543, n_18545, n_18546, n_18547, n_18550;
wire n_18527, n_18529, n_18530, n_18531, n_18532, n_18533, n_18534, n_18535;
wire n_18517, n_18518, n_18519, n_18520, n_18521, n_18523, n_18524, n_18526;
wire n_18505, n_18506, n_18507, n_18509, n_18511, n_18512, n_18515, n_18516;
wire n_18495, n_18496, n_18497, n_18498, n_18499, n_18500, n_18501, n_18504;
wire n_18479, n_18480, n_18482, n_18484, n_18486, n_18487, n_18492, n_18493;
wire n_18467, n_18468, n_18470, n_18471, n_18474, n_18475, n_18476, n_18478;
wire n_18457, n_18458, n_18459, n_18460, n_18461, n_18464, n_18465, n_18466;
wire n_18444, n_18447, n_18448, n_18449, n_18450, n_18454, n_18455, n_18456;
wire n_18435, n_18437, n_18438, n_18439, n_18440, n_18441, n_18442, n_18443;
wire n_18426, n_18427, n_18428, n_18429, n_18430, n_18432, n_18433, n_18434;
wire n_18416, n_18417, n_18418, n_18419, n_18420, n_18421, n_18424, n_18425;
wire n_18403, n_18405, n_18406, n_18407, n_18408, n_18410, n_18412, n_18414;
wire n_18394, n_18395, n_18396, n_18397, n_18399, n_18400, n_18401, n_18402;
wire n_18383, n_18384, n_18386, n_18387, n_18388, n_18389, n_18390, n_18391;
wire n_18373, n_18374, n_18375, n_18376, n_18377, n_18378, n_18379, n_18380;
wire n_18355, n_18356, n_18360, n_18362, n_18365, n_18368, n_18371, n_18372;
wire n_18346, n_18347, n_18348, n_18349, n_18351, n_18352, n_18353, n_18354;
wire n_18337, n_18338, n_18339, n_18340, n_18341, n_18342, n_18344, n_18345;
wire n_18329, n_18330, n_18331, n_18332, n_18333, n_18334, n_18335, n_18336;
wire n_18320, n_18321, n_18322, n_18323, n_18324, n_18325, n_18326, n_18328;
wire n_18306, n_18307, n_18309, n_18310, n_18311, n_18316, n_18317, n_18319;
wire n_18294, n_18295, n_18296, n_18298, n_18300, n_18302, n_18303, n_18304;
wire n_18283, n_18284, n_18285, n_18287, n_18288, n_18289, n_18290, n_18291;
wire n_18270, n_18271, n_18272, n_18274, n_18275, n_18276, n_18279, n_18281;
wire n_18258, n_18260, n_18261, n_18262, n_18263, n_18264, n_18265, n_18268;
wire n_18249, n_18250, n_18251, n_18252, n_18253, n_18254, n_18255, n_18256;
wire n_18229, n_18230, n_18231, n_18232, n_18234, n_18235, n_18236, n_18237;
wire n_18221, n_18222, n_18223, n_18224, n_18225, n_18226, n_18227, n_18228;
wire n_18211, n_18212, n_18213, n_18214, n_18217, n_18218, n_18219, n_18220;
wire n_18202, n_18203, n_18204, n_18205, n_18206, n_18207, n_18208, n_18209;
wire n_18194, n_18195, n_18196, n_18197, n_18198, n_18199, n_18200, n_18201;
wire n_18186, n_18187, n_18188, n_18189, n_18190, n_18191, n_18192, n_18193;
wire n_18178, n_18179, n_18180, n_18181, n_18182, n_18183, n_18184, n_18185;
wire n_18168, n_18169, n_18170, n_18171, n_18172, n_18173, n_18174, n_18176;
wire n_18159, n_18160, n_18161, n_18162, n_18163, n_18164, n_18165, n_18166;
wire n_18151, n_18152, n_18153, n_18154, n_18155, n_18156, n_18157, n_18158;
wire n_18142, n_18143, n_18144, n_18145, n_18146, n_18147, n_18149, n_18150;
wire n_18131, n_18134, n_18135, n_18136, n_18137, n_18138, n_18139, n_18140;
wire n_18122, n_18124, n_18125, n_18126, n_18127, n_18128, n_18129, n_18130;
wire n_18112, n_18113, n_18114, n_18115, n_18117, n_18118, n_18120, n_18121;
wire n_18101, n_18102, n_18103, n_18104, n_18106, n_18107, n_18108, n_18110;
wire n_18092, n_18093, n_18095, n_18096, n_18097, n_18098, n_18099, n_18100;
wire n_18080, n_18083, n_18085, n_18086, n_18087, n_18088, n_18089, n_18091;
wire n_18070, n_18071, n_18072, n_18073, n_18074, n_18077, n_18078, n_18079;
wire n_18061, n_18062, n_18063, n_18064, n_18065, n_18066, n_18068, n_18069;
wire n_18050, n_18051, n_18052, n_18055, n_18056, n_18057, n_18059, n_18060;
wire n_18042, n_18043, n_18044, n_18045, n_18046, n_18047, n_18048, n_18049;
wire n_18033, n_18034, n_18035, n_18036, n_18038, n_18039, n_18040, n_18041;
wire n_18024, n_18025, n_18026, n_18028, n_18029, n_18030, n_18031, n_18032;
wire n_18015, n_18016, n_18017, n_18018, n_18019, n_18020, n_18021, n_18023;
wire n_18006, n_18007, n_18008, n_18009, n_18010, n_18011, n_18012, n_18013;
wire n_17993, n_17994, n_17997, n_17999, n_18000, n_18001, n_18004, n_18005;
wire n_17982, n_17983, n_17984, n_17986, n_17987, n_17989, n_17990, n_17991;
wire n_17971, n_17972, n_17973, n_17974, n_17975, n_17977, n_17978, n_17980;
wire n_17958, n_17961, n_17962, n_17963, n_17967, n_17968, n_17969, n_17970;
wire n_17944, n_17945, n_17947, n_17948, n_17950, n_17951, n_17955, n_17956;
wire n_17933, n_17935, n_17937, n_17938, n_17939, n_17940, n_17942, n_17943;
wire n_17925, n_17926, n_17927, n_17928, n_17929, n_17930, n_17931, n_17932;
wire n_17916, n_17917, n_17918, n_17919, n_17920, n_17921, n_17922, n_17923;
wire n_17903, n_17904, n_17906, n_17907, n_17908, n_17909, n_17912, n_17915;
wire n_17894, n_17895, n_17896, n_17897, n_17898, n_17900, n_17901, n_17902;
wire n_17883, n_17884, n_17885, n_17886, n_17887, n_17888, n_17889, n_17892;
wire n_17873, n_17874, n_17876, n_17878, n_17879, n_17880, n_17881, n_17882;
wire n_17864, n_17865, n_17866, n_17867, n_17868, n_17870, n_17871, n_17872;
wire n_17855, n_17856, n_17858, n_17859, n_17860, n_17861, n_17862, n_17863;
wire n_17846, n_17847, n_17848, n_17849, n_17851, n_17852, n_17853, n_17854;
wire n_17836, n_17837, n_17839, n_17841, n_17842, n_17843, n_17844, n_17845;
wire n_17827, n_17828, n_17829, n_17830, n_17831, n_17832, n_17833, n_17835;
wire n_17815, n_17816, n_17817, n_17818, n_17820, n_17822, n_17824, n_17826;
wire n_17804, n_17806, n_17808, n_17809, n_17810, n_17812, n_17813, n_17814;
wire n_17796, n_17797, n_17798, n_17799, n_17800, n_17801, n_17802, n_17803;
wire n_17785, n_17786, n_17787, n_17788, n_17789, n_17793, n_17794, n_17795;
wire n_17776, n_17777, n_17778, n_17780, n_17781, n_17782, n_17783, n_17784;
wire n_17766, n_17767, n_17768, n_17770, n_17772, n_17773, n_17774, n_17775;
wire n_17755, n_17756, n_17758, n_17759, n_17760, n_17763, n_17764, n_17765;
wire n_17742, n_17743, n_17745, n_17747, n_17748, n_17750, n_17752, n_17754;
wire n_17725, n_17727, n_17729, n_17731, n_17732, n_17735, n_17739, n_17740;
wire n_17716, n_17717, n_17718, n_17719, n_17720, n_17721, n_17723, n_17724;
wire n_17707, n_17709, n_17710, n_17711, n_17712, n_17713, n_17714, n_17715;
wire n_17692, n_17698, n_17699, n_17701, n_17703, n_17704, n_17705, n_17706;
wire n_17684, n_17685, n_17686, n_17687, n_17688, n_17689, n_17690, n_17691;
wire n_17675, n_17677, n_17678, n_17679, n_17680, n_17681, n_17682, n_17683;
wire n_17665, n_17666, n_17668, n_17669, n_17670, n_17672, n_17673, n_17674;
wire n_17655, n_17656, n_17657, n_17659, n_17660, n_17661, n_17662, n_17664;
wire n_17635, n_17636, n_17637, n_17639, n_17647, n_17649, n_17652, n_17653;
wire n_17624, n_17625, n_17627, n_17628, n_17630, n_17631, n_17632, n_17634;
wire n_17616, n_17617, n_17618, n_17619, n_17620, n_17621, n_17622, n_17623;
wire n_17608, n_17609, n_17610, n_17611, n_17612, n_17613, n_17614, n_17615;
wire n_17598, n_17599, n_17602, n_17603, n_17604, n_17605, n_17606, n_17607;
wire n_17588, n_17589, n_17590, n_17591, n_17592, n_17595, n_17596, n_17597;
wire n_17580, n_17581, n_17582, n_17583, n_17584, n_17585, n_17586, n_17587;
wire n_17569, n_17570, n_17571, n_17573, n_17574, n_17576, n_17578, n_17579;
wire n_17557, n_17559, n_17560, n_17561, n_17562, n_17564, n_17565, n_17568;
wire n_17546, n_17549, n_17550, n_17551, n_17552, n_17553, n_17555, n_17556;
wire n_17535, n_17536, n_17537, n_17539, n_17540, n_17542, n_17543, n_17545;
wire n_17524, n_17525, n_17526, n_17527, n_17529, n_17532, n_17533, n_17534;
wire n_17513, n_17515, n_17516, n_17517, n_17518, n_17520, n_17521, n_17523;
wire n_17505, n_17506, n_17507, n_17508, n_17509, n_17510, n_17511, n_17512;
wire n_17497, n_17498, n_17499, n_17500, n_17501, n_17502, n_17503, n_17504;
wire n_17487, n_17488, n_17489, n_17491, n_17492, n_17493, n_17494, n_17495;
wire n_17475, n_17476, n_17479, n_17480, n_17481, n_17482, n_17483, n_17486;
wire n_17467, n_17468, n_17469, n_17470, n_17471, n_17472, n_17473, n_17474;
wire n_17453, n_17455, n_17458, n_17461, n_17463, n_17464, n_17465, n_17466;
wire n_17443, n_17444, n_17446, n_17447, n_17448, n_17450, n_17451, n_17452;
wire n_17429, n_17430, n_17431, n_17432, n_17433, n_17439, n_17441, n_17442;
wire n_17416, n_17418, n_17419, n_17424, n_17425, n_17426, n_17427, n_17428;
wire n_17407, n_17409, n_17410, n_17411, n_17412, n_17413, n_17414, n_17415;
wire n_17399, n_17400, n_17401, n_17402, n_17403, n_17404, n_17405, n_17406;
wire n_17389, n_17390, n_17391, n_17392, n_17395, n_17396, n_17397, n_17398;
wire n_17372, n_17374, n_17378, n_17380, n_17384, n_17386, n_17387, n_17388;
wire n_17361, n_17363, n_17364, n_17365, n_17366, n_17369, n_17370, n_17371;
wire n_17349, n_17351, n_17352, n_17356, n_17357, n_17358, n_17359, n_17360;
wire n_17340, n_17341, n_17342, n_17343, n_17344, n_17345, n_17346, n_17348;
wire n_17329, n_17330, n_17331, n_17334, n_17335, n_17337, n_17338, n_17339;
wire n_17316, n_17317, n_17318, n_17320, n_17322, n_17325, n_17326, n_17328;
wire n_17305, n_17307, n_17308, n_17309, n_17311, n_17312, n_17314, n_17315;
wire n_17297, n_17298, n_17299, n_17300, n_17301, n_17302, n_17303, n_17304;
wire n_17286, n_17287, n_17288, n_17289, n_17292, n_17293, n_17295, n_17296;
wire n_17277, n_17278, n_17279, n_17280, n_17282, n_17283, n_17284, n_17285;
wire n_17264, n_17267, n_17268, n_17270, n_17271, n_17273, n_17274, n_17276;
wire n_17255, n_17256, n_17257, n_17259, n_17260, n_17261, n_17262, n_17263;
wire n_17246, n_17247, n_17248, n_17249, n_17250, n_17251, n_17252, n_17253;
wire n_17234, n_17235, n_17236, n_17239, n_17240, n_17241, n_17242, n_17243;
wire n_17223, n_17224, n_17226, n_17228, n_17230, n_17231, n_17232, n_17233;
wire n_17204, n_17206, n_17207, n_17218, n_17219, n_17220, n_17221, n_17222;
wire n_17179, n_17181, n_17182, n_17183, n_17185, n_17186, n_17188, n_17203;
wire n_17166, n_17168, n_17172, n_17173, n_17174, n_17175, n_17177, n_17178;
wire n_17150, n_17155, n_17158, n_17161, n_17162, n_17163, n_17164, n_17165;
wire n_17139, n_17140, n_17142, n_17143, n_17145, n_17146, n_17147, n_17149;
wire n_17129, n_17130, n_17131, n_17132, n_17133, n_17136, n_17137, n_17138;
wire n_17090, n_17092, n_17112, n_17116, n_17117, n_17123, n_17125, n_17128;
wire n_17082, n_17083, n_17084, n_17085, n_17086, n_17087, n_17088, n_17089;
wire n_17073, n_17074, n_17075, n_17076, n_17077, n_17079, n_17080, n_17081;
wire n_17065, n_17066, n_17067, n_17068, n_17069, n_17070, n_17071, n_17072;
wire n_17057, n_17058, n_17059, n_17060, n_17061, n_17062, n_17063, n_17064;
wire n_17048, n_17049, n_17051, n_17052, n_17053, n_17054, n_17055, n_17056;
wire n_17036, n_17037, n_17038, n_17039, n_17040, n_17045, n_17046, n_17047;
wire n_17027, n_17028, n_17029, n_17030, n_17032, n_17033, n_17034, n_17035;
wire n_17018, n_17020, n_17021, n_17022, n_17023, n_17024, n_17025, n_17026;
wire n_17009, n_17010, n_17012, n_17013, n_17014, n_17015, n_17016, n_17017;
wire n_16999, n_17000, n_17001, n_17002, n_17003, n_17004, n_17007, n_17008;
wire n_16987, n_16988, n_16989, n_16991, n_16993, n_16994, n_16997, n_16998;
wire n_16975, n_16978, n_16980, n_16982, n_16983, n_16984, n_16985, n_16986;
wire n_16965, n_16966, n_16967, n_16968, n_16970, n_16972, n_16973, n_16974;
wire n_16949, n_16950, n_16951, n_16955, n_16958, n_16959, n_16960, n_16963;
wire n_16937, n_16938, n_16939, n_16943, n_16944, n_16945, n_16946, n_16947;
wire n_16922, n_16926, n_16927, n_16929, n_16930, n_16932, n_16934, n_16936;
wire n_16912, n_16914, n_16915, n_16916, n_16917, n_16918, n_16920, n_16921;
wire n_16900, n_16901, n_16902, n_16903, n_16904, n_16905, n_16907, n_16910;
wire n_16891, n_16892, n_16893, n_16894, n_16895, n_16897, n_16898, n_16899;
wire n_16879, n_16880, n_16881, n_16885, n_16886, n_16887, n_16888, n_16890;
wire n_16870, n_16871, n_16872, n_16873, n_16874, n_16875, n_16876, n_16878;
wire n_16857, n_16858, n_16861, n_16862, n_16864, n_16866, n_16867, n_16869;
wire n_16847, n_16848, n_16849, n_16851, n_16853, n_16854, n_16855, n_16856;
wire n_16837, n_16838, n_16840, n_16841, n_16842, n_16843, n_16844, n_16845;
wire n_16829, n_16830, n_16831, n_16832, n_16833, n_16834, n_16835, n_16836;
wire n_16818, n_16819, n_16820, n_16821, n_16823, n_16824, n_16825, n_16826;
wire n_16798, n_16799, n_16800, n_16801, n_16804, n_16808, n_16810, n_16817;
wire n_16786, n_16791, n_16792, n_16793, n_16794, n_16795, n_16796, n_16797;
wire n_16774, n_16776, n_16777, n_16778, n_16779, n_16782, n_16783, n_16785;
wire n_16765, n_16767, n_16768, n_16769, n_16770, n_16771, n_16772, n_16773;
wire n_16750, n_16754, n_16755, n_16757, n_16759, n_16760, n_16761, n_16764;
wire n_16741, n_16742, n_16743, n_16745, n_16746, n_16747, n_16748, n_16749;
wire n_16732, n_16733, n_16734, n_16735, n_16737, n_16738, n_16739, n_16740;
wire n_16696, n_16697, n_16699, n_16701, n_16702, n_16707, n_16728, n_16731;
wire n_16688, n_16689, n_16690, n_16691, n_16692, n_16693, n_16694, n_16695;
wire n_16679, n_16680, n_16682, n_16683, n_16684, n_16685, n_16686, n_16687;
wire n_16671, n_16672, n_16673, n_16674, n_16675, n_16676, n_16677, n_16678;
wire n_16662, n_16663, n_16664, n_16665, n_16666, n_16667, n_16669, n_16670;
wire n_16650, n_16652, n_16653, n_16655, n_16656, n_16658, n_16659, n_16660;
wire n_16637, n_16640, n_16641, n_16643, n_16644, n_16645, n_16646, n_16647;
wire n_16628, n_16629, n_16630, n_16631, n_16632, n_16633, n_16635, n_16636;
wire n_16614, n_16615, n_16616, n_16618, n_16619, n_16621, n_16624, n_16626;
wire n_16605, n_16606, n_16607, n_16609, n_16610, n_16611, n_16612, n_16613;
wire n_16589, n_16590, n_16591, n_16593, n_16594, n_16598, n_16599, n_16602;
wire n_16578, n_16580, n_16582, n_16583, n_16584, n_16585, n_16586, n_16587;
wire n_16570, n_16571, n_16572, n_16573, n_16574, n_16575, n_16576, n_16577;
wire n_16562, n_16563, n_16564, n_16565, n_16566, n_16567, n_16568, n_16569;
wire n_16553, n_16555, n_16556, n_16557, n_16558, n_16559, n_16560, n_16561;
wire n_16544, n_16546, n_16547, n_16548, n_16549, n_16550, n_16551, n_16552;
wire n_16535, n_16537, n_16538, n_16539, n_16540, n_16541, n_16542, n_16543;
wire n_16524, n_16526, n_16528, n_16529, n_16530, n_16531, n_16532, n_16533;
wire n_16511, n_16512, n_16514, n_16517, n_16518, n_16519, n_16521, n_16522;
wire n_16499, n_16500, n_16501, n_16502, n_16504, n_16505, n_16506, n_16510;
wire n_16477, n_16481, n_16486, n_16488, n_16494, n_16495, n_16496, n_16497;
wire n_16459, n_16460, n_16465, n_16468, n_16469, n_16473, n_16474, n_16475;
wire n_16450, n_16451, n_16452, n_16454, n_16455, n_16456, n_16457, n_16458;
wire n_16439, n_16440, n_16442, n_16443, n_16444, n_16445, n_16446, n_16448;
wire n_16428, n_16429, n_16430, n_16433, n_16434, n_16435, n_16436, n_16438;
wire n_16417, n_16419, n_16420, n_16421, n_16423, n_16424, n_16425, n_16427;
wire n_16403, n_16404, n_16406, n_16407, n_16411, n_16414, n_16415, n_16416;
wire n_16388, n_16389, n_16390, n_16391, n_16392, n_16396, n_16400, n_16402;
wire n_16379, n_16380, n_16381, n_16382, n_16383, n_16385, n_16386, n_16387;
wire n_16370, n_16371, n_16373, n_16374, n_16375, n_16376, n_16377, n_16378;
wire n_16361, n_16363, n_16364, n_16365, n_16366, n_16367, n_16368, n_16369;
wire n_16351, n_16353, n_16354, n_16355, n_16357, n_16358, n_16359, n_16360;
wire n_16341, n_16342, n_16344, n_16346, n_16347, n_16348, n_16349, n_16350;
wire n_16327, n_16328, n_16331, n_16334, n_16336, n_16337, n_16338, n_16339;
wire n_16319, n_16320, n_16321, n_16322, n_16323, n_16324, n_16325, n_16326;
wire n_16305, n_16306, n_16309, n_16311, n_16312, n_16315, n_16317, n_16318;
wire n_16293, n_16294, n_16295, n_16296, n_16297, n_16298, n_16299, n_16301;
wire n_16284, n_16285, n_16286, n_16288, n_16289, n_16290, n_16291, n_16292;
wire n_16274, n_16275, n_16276, n_16277, n_16278, n_16279, n_16281, n_16283;
wire n_16263, n_16265, n_16266, n_16267, n_16268, n_16269, n_16272, n_16273;
wire n_16253, n_16254, n_16255, n_16256, n_16257, n_16258, n_16260, n_16261;
wire n_16241, n_16242, n_16243, n_16245, n_16249, n_16250, n_16251, n_16252;
wire n_16228, n_16229, n_16230, n_16231, n_16234, n_16237, n_16238, n_16239;
wire n_16210, n_16212, n_16213, n_16214, n_16218, n_16219, n_16222, n_16225;
wire n_16191, n_16194, n_16196, n_16197, n_16199, n_16202, n_16203, n_16209;
wire n_16180, n_16181, n_16182, n_16183, n_16184, n_16186, n_16187, n_16188;
wire n_16170, n_16171, n_16172, n_16173, n_16174, n_16176, n_16177, n_16178;
wire n_16162, n_16163, n_16164, n_16165, n_16166, n_16167, n_16168, n_16169;
wire n_16149, n_16150, n_16151, n_16152, n_16154, n_16158, n_16160, n_16161;
wire n_16136, n_16137, n_16138, n_16140, n_16145, n_16146, n_16147, n_16148;
wire n_16115, n_16117, n_16120, n_16126, n_16130, n_16131, n_16134, n_16135;
wire n_16102, n_16103, n_16105, n_16107, n_16109, n_16112, n_16113, n_16114;
wire n_16092, n_16095, n_16096, n_16097, n_16098, n_16099, n_16100, n_16101;
wire n_16083, n_16084, n_16085, n_16086, n_16087, n_16089, n_16090, n_16091;
wire n_16072, n_16073, n_16074, n_16075, n_16076, n_16078, n_16079, n_16080;
wire n_16063, n_16064, n_16065, n_16066, n_16067, n_16068, n_16069, n_16071;
wire n_16047, n_16048, n_16051, n_16052, n_16054, n_16060, n_16061, n_16062;
wire n_16036, n_16039, n_16040, n_16041, n_16042, n_16043, n_16044, n_16046;
wire n_16015, n_16016, n_16025, n_16026, n_16027, n_16028, n_16031, n_16034;
wire n_16004, n_16005, n_16007, n_16008, n_16009, n_16010, n_16011, n_16012;
wire n_15989, n_15992, n_15995, n_15996, n_15997, n_15998, n_16002, n_16003;
wire n_15979, n_15980, n_15981, n_15982, n_15983, n_15984, n_15985, n_15988;
wire n_15969, n_15971, n_15972, n_15973, n_15974, n_15975, n_15976, n_15977;
wire n_15958, n_15959, n_15960, n_15962, n_15965, n_15966, n_15967, n_15968;
wire n_15947, n_15948, n_15949, n_15950, n_15951, n_15952, n_15953, n_15955;
wire n_15935, n_15936, n_15937, n_15938, n_15940, n_15943, n_15945, n_15946;
wire n_15924, n_15926, n_15928, n_15929, n_15930, n_15931, n_15932, n_15934;
wire n_15912, n_15913, n_15918, n_15919, n_15920, n_15921, n_15922, n_15923;
wire n_15904, n_15905, n_15906, n_15907, n_15908, n_15909, n_15910, n_15911;
wire n_15893, n_15894, n_15896, n_15897, n_15898, n_15899, n_15900, n_15902;
wire n_15877, n_15878, n_15879, n_15881, n_15884, n_15887, n_15889, n_15891;
wire n_15863, n_15864, n_15865, n_15868, n_15870, n_15872, n_15873, n_15875;
wire n_15854, n_15855, n_15856, n_15858, n_15859, n_15860, n_15861, n_15862;
wire n_15843, n_15844, n_15845, n_15849, n_15850, n_15851, n_15852, n_15853;
wire n_15835, n_15836, n_15837, n_15838, n_15839, n_15840, n_15841, n_15842;
wire n_15825, n_15827, n_15828, n_15829, n_15830, n_15831, n_15832, n_15833;
wire n_15813, n_15814, n_15815, n_15817, n_15819, n_15820, n_15821, n_15824;
wire n_15805, n_15806, n_15807, n_15808, n_15809, n_15810, n_15811, n_15812;
wire n_15793, n_15795, n_15797, n_15798, n_15800, n_15801, n_15802, n_15804;
wire n_15776, n_15778, n_15779, n_15783, n_15784, n_15785, n_15787, n_15791;
wire n_15766, n_15767, n_15768, n_15769, n_15771, n_15772, n_15773, n_15775;
wire n_15752, n_15753, n_15757, n_15761, n_15762, n_15763, n_15764, n_15765;
wire n_15736, n_15737, n_15739, n_15743, n_15745, n_15746, n_15747, n_15749;
wire n_15725, n_15726, n_15727, n_15728, n_15729, n_15731, n_15732, n_15733;
wire n_15715, n_15717, n_15718, n_15720, n_15721, n_15722, n_15723, n_15724;
wire n_15706, n_15707, n_15708, n_15709, n_15710, n_15711, n_15712, n_15714;
wire n_15698, n_15699, n_15700, n_15701, n_15702, n_15703, n_15704, n_15705;
wire n_15687, n_15688, n_15689, n_15690, n_15691, n_15692, n_15693, n_15696;
wire n_15676, n_15677, n_15678, n_15679, n_15680, n_15681, n_15685, n_15686;
wire n_15667, n_15668, n_15670, n_15671, n_15672, n_15673, n_15674, n_15675;
wire n_15656, n_15657, n_15658, n_15659, n_15661, n_15663, n_15665, n_15666;
wire n_15647, n_15649, n_15650, n_15651, n_15652, n_15653, n_15654, n_15655;
wire n_15639, n_15640, n_15641, n_15642, n_15643, n_15644, n_15645, n_15646;
wire n_15631, n_15632, n_15633, n_15634, n_15635, n_15636, n_15637, n_15638;
wire n_15622, n_15623, n_15625, n_15626, n_15627, n_15628, n_15629, n_15630;
wire n_15612, n_15613, n_15614, n_15615, n_15616, n_15619, n_15620, n_15621;
wire n_15598, n_15599, n_15601, n_15602, n_15603, n_15608, n_15609, n_15610;
wire n_15587, n_15588, n_15589, n_15590, n_15591, n_15592, n_15593, n_15596;
wire n_15578, n_15579, n_15580, n_15581, n_15583, n_15584, n_15585, n_15586;
wire n_15570, n_15571, n_15572, n_15573, n_15574, n_15575, n_15576, n_15577;
wire n_15562, n_15563, n_15564, n_15565, n_15566, n_15567, n_15568, n_15569;
wire n_15551, n_15552, n_15556, n_15557, n_15558, n_15559, n_15560, n_15561;
wire n_15541, n_15542, n_15544, n_15545, n_15546, n_15547, n_15548, n_15549;
wire n_15533, n_15534, n_15535, n_15536, n_15537, n_15538, n_15539, n_15540;
wire n_15524, n_15526, n_15527, n_15528, n_15529, n_15530, n_15531, n_15532;
wire n_15516, n_15517, n_15518, n_15519, n_15520, n_15521, n_15522, n_15523;
wire n_15506, n_15508, n_15509, n_15510, n_15511, n_15512, n_15513, n_15514;
wire n_15497, n_15498, n_15499, n_15500, n_15501, n_15502, n_15504, n_15505;
wire n_15484, n_15485, n_15486, n_15487, n_15490, n_15491, n_15492, n_15493;
wire n_15474, n_15476, n_15477, n_15478, n_15479, n_15480, n_15481, n_15482;
wire n_15462, n_15464, n_15465, n_15466, n_15467, n_15470, n_15471, n_15473;
wire n_15453, n_15454, n_15456, n_15457, n_15458, n_15459, n_15460, n_15461;
wire n_15445, n_15446, n_15447, n_15448, n_15449, n_15450, n_15451, n_15452;
wire n_15435, n_15436, n_15437, n_15440, n_15441, n_15442, n_15443, n_15444;
wire n_15427, n_15428, n_15429, n_15430, n_15431, n_15432, n_15433, n_15434;
wire n_15414, n_15415, n_15416, n_15419, n_15421, n_15422, n_15424, n_15426;
wire n_15404, n_15405, n_15406, n_15407, n_15408, n_15409, n_15410, n_15413;
wire n_15394, n_15395, n_15396, n_15397, n_15398, n_15399, n_15400, n_15403;
wire n_15384, n_15385, n_15387, n_15389, n_15390, n_15391, n_15392, n_15393;
wire n_15375, n_15376, n_15377, n_15378, n_15379, n_15380, n_15381, n_15382;
wire n_15366, n_15367, n_15368, n_15369, n_15370, n_15371, n_15372, n_15374;
wire n_15353, n_15356, n_15357, n_15358, n_15360, n_15362, n_15363, n_15365;
wire n_15342, n_15344, n_15345, n_15346, n_15347, n_15348, n_15350, n_15352;
wire n_15334, n_15335, n_15336, n_15337, n_15338, n_15339, n_15340, n_15341;
wire n_15320, n_15322, n_15324, n_15325, n_15327, n_15329, n_15332, n_15333;
wire n_15306, n_15311, n_15313, n_15314, n_15315, n_15316, n_15317, n_15318;
wire n_15298, n_15299, n_15300, n_15301, n_15302, n_15303, n_15304, n_15305;
wire n_15290, n_15291, n_15292, n_15293, n_15294, n_15295, n_15296, n_15297;
wire n_15280, n_15281, n_15282, n_15284, n_15285, n_15287, n_15288, n_15289;
wire n_15269, n_15271, n_15272, n_15273, n_15275, n_15277, n_15278, n_15279;
wire n_15259, n_15260, n_15261, n_15262, n_15263, n_15264, n_15266, n_15267;
wire n_15251, n_15252, n_15253, n_15254, n_15255, n_15256, n_15257, n_15258;
wire n_15238, n_15239, n_15240, n_15244, n_15245, n_15247, n_15249, n_15250;
wire n_15229, n_15230, n_15231, n_15232, n_15234, n_15235, n_15236, n_15237;
wire n_15216, n_15218, n_15220, n_15222, n_15224, n_15226, n_15227, n_15228;
wire n_15206, n_15208, n_15209, n_15210, n_15211, n_15212, n_15213, n_15214;
wire n_15196, n_15197, n_15198, n_15199, n_15201, n_15202, n_15203, n_15205;
wire n_15185, n_15186, n_15187, n_15190, n_15192, n_15193, n_15194, n_15195;
wire n_15177, n_15178, n_15179, n_15180, n_15181, n_15182, n_15183, n_15184;
wire n_15168, n_15169, n_15170, n_15172, n_15173, n_15174, n_15175, n_15176;
wire n_15157, n_15158, n_15160, n_15161, n_15162, n_15163, n_15164, n_15165;
wire n_15148, n_15149, n_15150, n_15151, n_15152, n_15153, n_15154, n_15155;
wire n_15140, n_15141, n_15142, n_15143, n_15144, n_15145, n_15146, n_15147;
wire n_15130, n_15131, n_15132, n_15133, n_15134, n_15136, n_15138, n_15139;
wire n_15121, n_15122, n_15123, n_15125, n_15126, n_15127, n_15128, n_15129;
wire n_15113, n_15114, n_15115, n_15116, n_15117, n_15118, n_15119, n_15120;
wire n_15104, n_15105, n_15106, n_15107, n_15109, n_15110, n_15111, n_15112;
wire n_15092, n_15094, n_15095, n_15096, n_15097, n_15098, n_15101, n_15103;
wire n_15082, n_15083, n_15085, n_15086, n_15087, n_15088, n_15089, n_15090;
wire n_15073, n_15074, n_15075, n_15076, n_15077, n_15078, n_15079, n_15081;
wire n_15059, n_15060, n_15061, n_15066, n_15067, n_15069, n_15071, n_15072;
wire n_15051, n_15052, n_15053, n_15054, n_15055, n_15056, n_15057, n_15058;
wire n_15039, n_15041, n_15043, n_15044, n_15045, n_15046, n_15047, n_15049;
wire n_15029, n_15030, n_15031, n_15032, n_15034, n_15036, n_15037, n_15038;
wire n_15020, n_15021, n_15023, n_15024, n_15025, n_15026, n_15027, n_15028;
wire n_15008, n_15009, n_15010, n_15011, n_15013, n_15016, n_15017, n_15018;
wire n_15000, n_15001, n_15002, n_15003, n_15004, n_15005, n_15006, n_15007;
wire n_14991, n_14993, n_14994, n_14995, n_14996, n_14997, n_14998, n_14999;
wire n_14982, n_14983, n_14984, n_14985, n_14986, n_14987, n_14989, n_14990;
wire n_14972, n_14973, n_14975, n_14976, n_14977, n_14978, n_14979, n_14980;
wire n_14963, n_14964, n_14965, n_14966, n_14967, n_14968, n_14970, n_14971;
wire n_14955, n_14956, n_14957, n_14958, n_14959, n_14960, n_14961, n_14962;
wire n_14946, n_14947, n_14948, n_14949, n_14950, n_14951, n_14952, n_14953;
wire n_14935, n_14936, n_14939, n_14940, n_14941, n_14943, n_14944, n_14945;
wire n_14925, n_14927, n_14928, n_14929, n_14930, n_14931, n_14932, n_14933;
wire n_14917, n_14918, n_14919, n_14920, n_14921, n_14922, n_14923, n_14924;
wire n_14908, n_14909, n_14910, n_14911, n_14912, n_14913, n_14915, n_14916;
wire n_14899, n_14900, n_14901, n_14902, n_14903, n_14904, n_14905, n_14907;
wire n_14887, n_14888, n_14889, n_14891, n_14893, n_14895, n_14896, n_14897;
wire n_14879, n_14880, n_14881, n_14882, n_14883, n_14884, n_14885, n_14886;
wire n_14870, n_14871, n_14872, n_14873, n_14875, n_14876, n_14877, n_14878;
wire n_14862, n_14863, n_14864, n_14865, n_14866, n_14867, n_14868, n_14869;
wire n_14854, n_14855, n_14856, n_14857, n_14858, n_14859, n_14860, n_14861;
wire n_14846, n_14847, n_14848, n_14849, n_14850, n_14851, n_14852, n_14853;
wire n_14834, n_14835, n_14837, n_14838, n_14839, n_14843, n_14844, n_14845;
wire n_14825, n_14826, n_14827, n_14828, n_14829, n_14831, n_14832, n_14833;
wire n_14817, n_14818, n_14819, n_14820, n_14821, n_14822, n_14823, n_14824;
wire n_14809, n_14810, n_14811, n_14812, n_14813, n_14814, n_14815, n_14816;
wire n_14801, n_14802, n_14803, n_14804, n_14805, n_14806, n_14807, n_14808;
wire n_14793, n_14794, n_14795, n_14796, n_14797, n_14798, n_14799, n_14800;
wire n_14785, n_14786, n_14787, n_14788, n_14789, n_14790, n_14791, n_14792;
wire n_14777, n_14778, n_14779, n_14780, n_14781, n_14782, n_14783, n_14784;
wire n_14768, n_14769, n_14771, n_14772, n_14773, n_14774, n_14775, n_14776;
wire n_14756, n_14757, n_14758, n_14759, n_14761, n_14763, n_14764, n_14765;
wire n_14745, n_14747, n_14748, n_14749, n_14750, n_14752, n_14753, n_14755;
wire n_14736, n_14737, n_14738, n_14740, n_14741, n_14742, n_14743, n_14744;
wire n_14727, n_14728, n_14729, n_14731, n_14732, n_14733, n_14734, n_14735;
wire n_14719, n_14720, n_14721, n_14722, n_14723, n_14724, n_14725, n_14726;
wire n_14709, n_14711, n_14712, n_14714, n_14715, n_14716, n_14717, n_14718;
wire n_14701, n_14702, n_14703, n_14704, n_14705, n_14706, n_14707, n_14708;
wire n_14692, n_14693, n_14694, n_14695, n_14696, n_14697, n_14698, n_14700;
wire n_14684, n_14685, n_14686, n_14687, n_14688, n_14689, n_14690, n_14691;
wire n_14675, n_14676, n_14677, n_14678, n_14679, n_14680, n_14682, n_14683;
wire n_14666, n_14667, n_14668, n_14669, n_14670, n_14672, n_14673, n_14674;
wire n_14658, n_14659, n_14660, n_14661, n_14662, n_14663, n_14664, n_14665;
wire n_14649, n_14650, n_14652, n_14653, n_14654, n_14655, n_14656, n_14657;
wire n_14641, n_14642, n_14643, n_14644, n_14645, n_14646, n_14647, n_14648;
wire n_14633, n_14634, n_14635, n_14636, n_14637, n_14638, n_14639, n_14640;
wire n_14625, n_14626, n_14627, n_14628, n_14629, n_14630, n_14631, n_14632;
wire n_14615, n_14616, n_14617, n_14618, n_14621, n_14622, n_14623, n_14624;
wire n_14606, n_14608, n_14609, n_14610, n_14611, n_14612, n_14613, n_14614;
wire n_14598, n_14599, n_14600, n_14601, n_14602, n_14603, n_14604, n_14605;
wire n_14589, n_14590, n_14592, n_14593, n_14594, n_14595, n_14596, n_14597;
wire n_14580, n_14581, n_14582, n_14583, n_14584, n_14585, n_14586, n_14587;
wire n_14572, n_14573, n_14574, n_14575, n_14576, n_14577, n_14578, n_14579;
wire n_14564, n_14565, n_14566, n_14567, n_14568, n_14569, n_14570, n_14571;
wire n_14556, n_14557, n_14558, n_14559, n_14560, n_14561, n_14562, n_14563;
wire n_14547, n_14548, n_14549, n_14550, n_14551, n_14552, n_14554, n_14555;
wire n_14537, n_14538, n_14539, n_14540, n_14542, n_14543, n_14544, n_14545;
wire n_14528, n_14529, n_14531, n_14532, n_14533, n_14534, n_14535, n_14536;
wire n_14520, n_14521, n_14522, n_14523, n_14524, n_14525, n_14526, n_14527;
wire n_14510, n_14511, n_14512, n_14513, n_14514, n_14516, n_14517, n_14518;
wire n_14498, n_14499, n_14503, n_14504, n_14505, n_14506, n_14508, n_14509;
wire n_14486, n_14490, n_14491, n_14492, n_14494, n_14495, n_14496, n_14497;
wire n_14478, n_14479, n_14480, n_14481, n_14482, n_14483, n_14484, n_14485;
wire n_14468, n_14469, n_14470, n_14471, n_14473, n_14474, n_14476, n_14477;
wire n_14460, n_14461, n_14462, n_14463, n_14464, n_14465, n_14466, n_14467;
wire n_14452, n_14453, n_14454, n_14455, n_14456, n_14457, n_14458, n_14459;
wire n_14440, n_14442, n_14444, n_14445, n_14446, n_14448, n_14449, n_14450;
wire n_14431, n_14432, n_14433, n_14434, n_14435, n_14436, n_14437, n_14439;
wire n_14422, n_14423, n_14424, n_14425, n_14426, n_14428, n_14429, n_14430;
wire n_14414, n_14415, n_14416, n_14417, n_14418, n_14419, n_14420, n_14421;
wire n_14406, n_14407, n_14408, n_14409, n_14410, n_14411, n_14412, n_14413;
wire n_14397, n_14398, n_14399, n_14400, n_14401, n_14403, n_14404, n_14405;
wire n_14386, n_14387, n_14388, n_14389, n_14390, n_14391, n_14394, n_14395;
wire n_14377, n_14379, n_14380, n_14381, n_14382, n_14383, n_14384, n_14385;
wire n_14369, n_14370, n_14371, n_14372, n_14373, n_14374, n_14375, n_14376;
wire n_14360, n_14361, n_14362, n_14363, n_14365, n_14366, n_14367, n_14368;
wire n_14352, n_14353, n_14354, n_14355, n_14356, n_14357, n_14358, n_14359;
wire n_14344, n_14345, n_14346, n_14347, n_14348, n_14349, n_14350, n_14351;
wire n_14335, n_14336, n_14337, n_14339, n_14340, n_14341, n_14342, n_14343;
wire n_14327, n_14328, n_14329, n_14330, n_14331, n_14332, n_14333, n_14334;
wire n_14318, n_14319, n_14320, n_14321, n_14322, n_14323, n_14325, n_14326;
wire n_14305, n_14306, n_14307, n_14309, n_14311, n_14313, n_14316, n_14317;
wire n_14291, n_14292, n_14295, n_14297, n_14298, n_14299, n_14303, n_14304;
wire n_14272, n_14274, n_14275, n_14276, n_14279, n_14282, n_14286, n_14287;
wire n_14263, n_14264, n_14266, n_14267, n_14268, n_14269, n_14270, n_14271;
wire n_14252, n_14254, n_14256, n_14257, n_14258, n_14259, n_14260, n_14261;
wire n_14241, n_14242, n_14243, n_14244, n_14246, n_14247, n_14248, n_14249;
wire n_14233, n_14234, n_14235, n_14236, n_14237, n_14238, n_14239, n_14240;
wire n_14223, n_14224, n_14225, n_14226, n_14227, n_14229, n_14230, n_14232;
wire n_14213, n_14214, n_14217, n_14218, n_14219, n_14220, n_14221, n_14222;
wire n_14204, n_14206, n_14207, n_14208, n_14209, n_14210, n_14211, n_14212;
wire n_14196, n_14197, n_14198, n_14199, n_14200, n_14201, n_14202, n_14203;
wire n_14187, n_14188, n_14189, n_14190, n_14191, n_14192, n_14193, n_14194;
wire n_14178, n_14179, n_14180, n_14181, n_14182, n_14184, n_14185, n_14186;
wire n_14163, n_14164, n_14168, n_14169, n_14172, n_14173, n_14176, n_14177;
wire n_14154, n_14155, n_14157, n_14158, n_14159, n_14160, n_14161, n_14162;
wire n_14141, n_14143, n_14147, n_14148, n_14150, n_14151, n_14152, n_14153;
wire n_14126, n_14128, n_14129, n_14131, n_14133, n_14134, n_14135, n_14139;
wire n_14112, n_14116, n_14117, n_14118, n_14121, n_14123, n_14124, n_14125;
wire n_14097, n_14100, n_14101, n_14102, n_14104, n_14107, n_14108, n_14109;
wire n_14080, n_14084, n_14086, n_14087, n_14089, n_14090, n_14094, n_14096;
wire n_14058, n_14059, n_14071, n_14072, n_14074, n_14076, n_14078, n_14079;
wire n_14045, n_14049, n_14051, n_14053, n_14054, n_14055, n_14056, n_14057;
wire n_14023, n_14024, n_14025, n_14026, n_14027, n_14032, n_14036, n_14042;
wire n_14011, n_14012, n_14014, n_14016, n_14017, n_14018, n_14019, n_14022;
wire n_14002, n_14003, n_14005, n_14006, n_14007, n_14008, n_14009, n_14010;
wire n_13991, n_13992, n_13993, n_13994, n_13996, n_13998, n_13999, n_14001;
wire n_13983, n_13984, n_13985, n_13986, n_13987, n_13988, n_13989, n_13990;
wire n_13970, n_13973, n_13974, n_13976, n_13977, n_13978, n_13979, n_13981;
wire n_13961, n_13962, n_13963, n_13964, n_13965, n_13966, n_13967, n_13968;
wire n_13953, n_13954, n_13955, n_13956, n_13957, n_13958, n_13959, n_13960;
wire n_13944, n_13945, n_13946, n_13948, n_13949, n_13950, n_13951, n_13952;
wire n_13936, n_13937, n_13938, n_13939, n_13940, n_13941, n_13942, n_13943;
wire n_13927, n_13928, n_13929, n_13930, n_13931, n_13932, n_13933, n_13935;
wire n_13918, n_13919, n_13920, n_13921, n_13922, n_13923, n_13924, n_13925;
wire n_13908, n_13909, n_13911, n_13912, n_13913, n_13914, n_13915, n_13917;
wire n_13899, n_13900, n_13901, n_13902, n_13903, n_13904, n_13905, n_13907;
wire n_13891, n_13892, n_13893, n_13894, n_13895, n_13896, n_13897, n_13898;
wire n_13877, n_13878, n_13880, n_13881, n_13883, n_13885, n_13888, n_13890;
wire n_13862, n_13863, n_13864, n_13866, n_13868, n_13871, n_13873, n_13875;
wire n_13839, n_13840, n_13842, n_13843, n_13845, n_13850, n_13852, n_13854;
wire n_13813, n_13817, n_13820, n_13821, n_13822, n_13823, n_13826, n_13838;
wire n_13803, n_13804, n_13805, n_13806, n_13807, n_13809, n_13810, n_13811;
wire n_13791, n_13793, n_13796, n_13798, n_13799, n_13800, n_13801, n_13802;
wire n_13783, n_13784, n_13785, n_13786, n_13787, n_13788, n_13789, n_13790;
wire n_13775, n_13776, n_13777, n_13778, n_13779, n_13780, n_13781, n_13782;
wire n_13766, n_13767, n_13768, n_13769, n_13770, n_13771, n_13773, n_13774;
wire n_13758, n_13759, n_13760, n_13761, n_13762, n_13763, n_13764, n_13765;
wire n_13744, n_13745, n_13746, n_13747, n_13748, n_13749, n_13755, n_13757;
wire n_13735, n_13736, n_13737, n_13738, n_13739, n_13741, n_13742, n_13743;
wire n_13720, n_13721, n_13723, n_13724, n_13727, n_13728, n_13732, n_13734;
wire n_13699, n_13701, n_13709, n_13711, n_13712, n_13714, n_13716, n_13717;
wire n_13687, n_13689, n_13690, n_13692, n_13695, n_13696, n_13697, n_13698;
wire n_13675, n_13677, n_13678, n_13679, n_13680, n_13681, n_13683, n_13686;
wire n_13663, n_13664, n_13665, n_13667, n_13668, n_13669, n_13670, n_13673;
wire n_13653, n_13654, n_13655, n_13657, n_13659, n_13660, n_13661, n_13662;
wire n_13644, n_13645, n_13646, n_13647, n_13648, n_13650, n_13651, n_13652;
wire n_13633, n_13634, n_13635, n_13637, n_13638, n_13639, n_13640, n_13641;
wire n_13616, n_13620, n_13622, n_13624, n_13627, n_13628, n_13629, n_13632;
wire n_13582, n_13584, n_13588, n_13600, n_13601, n_13602, n_13604, n_13613;
wire n_13564, n_13569, n_13571, n_13572, n_13573, n_13574, n_13579, n_13581;
wire n_13551, n_13552, n_13553, n_13554, n_13555, n_13557, n_13558, n_13559;
wire n_13540, n_13541, n_13542, n_13544, n_13545, n_13546, n_13548, n_13549;
wire n_13528, n_13529, n_13530, n_13531, n_13533, n_13536, n_13537, n_13538;
wire n_13519, n_13520, n_13521, n_13523, n_13524, n_13525, n_13526, n_13527;
wire n_13504, n_13507, n_13509, n_13510, n_13511, n_13515, n_13516, n_13518;
wire n_13492, n_13493, n_13494, n_13496, n_13497, n_13498, n_13499, n_13502;
wire n_13482, n_13484, n_13485, n_13487, n_13488, n_13489, n_13490, n_13491;
wire n_13458, n_13461, n_13464, n_13466, n_13467, n_13469, n_13470, n_13478;
wire n_13435, n_13437, n_13444, n_13448, n_13452, n_13454, n_13455, n_13457;
wire n_13421, n_13425, n_13426, n_13427, n_13428, n_13429, n_13432, n_13434;
wire n_13411, n_13412, n_13413, n_13415, n_13416, n_13417, n_13418, n_13419;
wire n_13402, n_13403, n_13404, n_13406, n_13407, n_13408, n_13409, n_13410;
wire n_13388, n_13389, n_13393, n_13394, n_13396, n_13399, n_13400, n_13401;
wire n_13378, n_13379, n_13380, n_13381, n_13383, n_13385, n_13386, n_13387;
wire n_13368, n_13370, n_13372, n_13373, n_13374, n_13375, n_13376, n_13377;
wire n_13355, n_13357, n_13358, n_13359, n_13361, n_13365, n_13366, n_13367;
wire n_13346, n_13347, n_13348, n_13350, n_13351, n_13352, n_13353, n_13354;
wire n_13336, n_13337, n_13338, n_13340, n_13341, n_13342, n_13343, n_13344;
wire n_13325, n_13327, n_13329, n_13330, n_13332, n_13333, n_13334, n_13335;
wire n_13313, n_13316, n_13317, n_13318, n_13320, n_13321, n_13322, n_13323;
wire n_13287, n_13296, n_13297, n_13299, n_13301, n_13304, n_13311, n_13312;
wire n_13274, n_13277, n_13279, n_13280, n_13281, n_13283, n_13284, n_13285;
wire n_13243, n_13245, n_13248, n_13251, n_13252, n_13264, n_13268, n_13273;
wire n_13234, n_13235, n_13236, n_13237, n_13238, n_13239, n_13240, n_13242;
wire n_13223, n_13225, n_13227, n_13228, n_13230, n_13231, n_13232, n_13233;
wire n_13214, n_13215, n_13216, n_13217, n_13219, n_13220, n_13221, n_13222;
wire n_13205, n_13206, n_13207, n_13208, n_13209, n_13211, n_13212, n_13213;
wire n_13197, n_13198, n_13199, n_13200, n_13201, n_13202, n_13203, n_13204;
wire n_13188, n_13189, n_13191, n_13192, n_13193, n_13194, n_13195, n_13196;
wire n_13179, n_13180, n_13181, n_13183, n_13184, n_13185, n_13186, n_13187;
wire n_13166, n_13167, n_13169, n_13170, n_13171, n_13173, n_13174, n_13175;
wire n_13145, n_13147, n_13150, n_13151, n_13152, n_13154, n_13156, n_13163;
wire n_13125, n_13126, n_13128, n_13130, n_13131, n_13134, n_13137, n_13143;
wire n_13114, n_13117, n_13119, n_13120, n_13121, n_13122, n_13123, n_13124;
wire n_13102, n_13103, n_13104, n_13105, n_13106, n_13108, n_13111, n_13112;
wire n_13093, n_13094, n_13095, n_13096, n_13097, n_13098, n_13100, n_13101;
wire n_13084, n_13085, n_13086, n_13087, n_13088, n_13090, n_13091, n_13092;
wire n_13071, n_13072, n_13075, n_13076, n_13078, n_13080, n_13081, n_13082;
wire n_13059, n_13060, n_13062, n_13064, n_13065, n_13066, n_13067, n_13068;
wire n_13046, n_13049, n_13051, n_13053, n_13054, n_13055, n_13056, n_13058;
wire n_13033, n_13034, n_13035, n_13038, n_13039, n_13040, n_13042, n_13045;
wire n_13023, n_13024, n_13025, n_13026, n_13027, n_13028, n_13031, n_13032;
wire n_13014, n_13015, n_13016, n_13017, n_13018, n_13019, n_13020, n_13022;
wire n_13006, n_13007, n_13008, n_13009, n_13010, n_13011, n_13012, n_13013;
wire n_12998, n_12999, n_13000, n_13001, n_13002, n_13003, n_13004, n_13005;
wire n_12989, n_12991, n_12992, n_12993, n_12994, n_12995, n_12996, n_12997;
wire n_12976, n_12977, n_12978, n_12979, n_12981, n_12985, n_12986, n_12987;
wire n_12968, n_12969, n_12970, n_12971, n_12972, n_12973, n_12974, n_12975;
wire n_12960, n_12961, n_12962, n_12963, n_12964, n_12965, n_12966, n_12967;
wire n_12950, n_12951, n_12952, n_12953, n_12954, n_12955, n_12956, n_12959;
wire n_12941, n_12942, n_12943, n_12944, n_12945, n_12947, n_12948, n_12949;
wire n_12931, n_12933, n_12934, n_12936, n_12937, n_12938, n_12939, n_12940;
wire n_12918, n_12920, n_12921, n_12923, n_12925, n_12926, n_12927, n_12930;
wire n_12908, n_12910, n_12911, n_12912, n_12913, n_12915, n_12916, n_12917;
wire n_12897, n_12899, n_12900, n_12901, n_12902, n_12905, n_12906, n_12907;
wire n_12889, n_12890, n_12891, n_12892, n_12893, n_12894, n_12895, n_12896;
wire n_12880, n_12881, n_12882, n_12883, n_12885, n_12886, n_12887, n_12888;
wire n_12872, n_12873, n_12874, n_12875, n_12876, n_12877, n_12878, n_12879;
wire n_12861, n_12862, n_12863, n_12865, n_12866, n_12867, n_12869, n_12871;
wire n_12850, n_12851, n_12852, n_12853, n_12856, n_12857, n_12858, n_12860;
wire n_12839, n_12840, n_12841, n_12843, n_12844, n_12845, n_12846, n_12848;
wire n_12829, n_12830, n_12831, n_12832, n_12834, n_12835, n_12836, n_12838;
wire n_12820, n_12821, n_12822, n_12823, n_12824, n_12825, n_12826, n_12827;
wire n_12812, n_12813, n_12814, n_12815, n_12816, n_12817, n_12818, n_12819;
wire n_12804, n_12805, n_12806, n_12807, n_12808, n_12809, n_12810, n_12811;
wire n_12795, n_12796, n_12798, n_12799, n_12800, n_12801, n_12802, n_12803;
wire n_12786, n_12787, n_12788, n_12789, n_12790, n_12791, n_12792, n_12793;
wire n_12778, n_12779, n_12780, n_12781, n_12782, n_12783, n_12784, n_12785;
wire n_12769, n_12770, n_12771, n_12772, n_12774, n_12775, n_12776, n_12777;
wire n_12761, n_12762, n_12763, n_12764, n_12765, n_12766, n_12767, n_12768;
wire n_12752, n_12753, n_12754, n_12755, n_12756, n_12757, n_12759, n_12760;
wire n_12740, n_12741, n_12742, n_12744, n_12746, n_12749, n_12750, n_12751;
wire n_12732, n_12733, n_12734, n_12735, n_12736, n_12737, n_12738, n_12739;
wire n_12723, n_12724, n_12725, n_12726, n_12728, n_12729, n_12730, n_12731;
wire n_12715, n_12716, n_12717, n_12718, n_12719, n_12720, n_12721, n_12722;
wire n_12705, n_12706, n_12707, n_12709, n_12711, n_12712, n_12713, n_12714;
wire n_12696, n_12697, n_12698, n_12700, n_12701, n_12702, n_12703, n_12704;
wire n_12688, n_12689, n_12690, n_12691, n_12692, n_12693, n_12694, n_12695;
wire n_12680, n_12681, n_12682, n_12683, n_12684, n_12685, n_12686, n_12687;
wire n_12671, n_12672, n_12673, n_12674, n_12675, n_12676, n_12677, n_12678;
wire n_12662, n_12663, n_12664, n_12665, n_12667, n_12668, n_12669, n_12670;
wire n_12653, n_12654, n_12655, n_12656, n_12657, n_12658, n_12659, n_12661;
wire n_12644, n_12645, n_12646, n_12647, n_12648, n_12649, n_12650, n_12651;
wire n_12635, n_12636, n_12638, n_12639, n_12640, n_12641, n_12642, n_12643;
wire n_12626, n_12627, n_12628, n_12629, n_12630, n_12631, n_12632, n_12633;
wire n_12617, n_12618, n_12619, n_12621, n_12622, n_12623, n_12624, n_12625;
wire n_12607, n_12609, n_12611, n_12612, n_12613, n_12614, n_12615, n_12616;
wire n_12598, n_12599, n_12600, n_12601, n_12602, n_12603, n_12605, n_12606;
wire n_12589, n_12591, n_12592, n_12593, n_12594, n_12595, n_12596, n_12597;
wire n_12579, n_12580, n_12581, n_12582, n_12585, n_12586, n_12587, n_12588;
wire n_12568, n_12570, n_12572, n_12574, n_12575, n_12576, n_12577, n_12578;
wire n_12557, n_12559, n_12561, n_12562, n_12563, n_12564, n_12565, n_12566;
wire n_12545, n_12546, n_12547, n_12549, n_12551, n_12553, n_12555, n_12556;
wire n_12536, n_12537, n_12538, n_12539, n_12540, n_12542, n_12543, n_12544;
wire n_12525, n_12526, n_12527, n_12528, n_12530, n_12531, n_12532, n_12535;
wire n_12516, n_12517, n_12518, n_12519, n_12520, n_12521, n_12522, n_12523;
wire n_12505, n_12507, n_12508, n_12510, n_12511, n_12512, n_12514, n_12515;
wire n_12494, n_12495, n_12496, n_12498, n_12500, n_12502, n_12503, n_12504;
wire n_12484, n_12486, n_12487, n_12488, n_12489, n_12491, n_12492, n_12493;
wire n_12475, n_12476, n_12477, n_12479, n_12480, n_12481, n_12482, n_12483;
wire n_12464, n_12466, n_12467, n_12468, n_12469, n_12470, n_12471, n_12473;
wire n_12455, n_12456, n_12457, n_12458, n_12459, n_12460, n_12461, n_12462;
wire n_12443, n_12445, n_12446, n_12449, n_12450, n_12451, n_12452, n_12454;
wire n_12431, n_12432, n_12433, n_12434, n_12435, n_12436, n_12437, n_12442;
wire n_12423, n_12424, n_12425, n_12426, n_12427, n_12428, n_12429, n_12430;
wire n_12410, n_12412, n_12414, n_12415, n_12417, n_12418, n_12419, n_12422;
wire n_12398, n_12400, n_12402, n_12403, n_12404, n_12405, n_12407, n_12408;
wire n_12389, n_12390, n_12391, n_12393, n_12394, n_12395, n_12396, n_12397;
wire n_12379, n_12380, n_12381, n_12383, n_12384, n_12385, n_12386, n_12388;
wire n_12366, n_12367, n_12368, n_12369, n_12373, n_12374, n_12376, n_12378;
wire n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364, n_12365;
wire n_12350, n_12351, n_12352, n_12353, n_12354, n_12355, n_12356, n_12357;
wire n_12341, n_12342, n_12343, n_12344, n_12345, n_12347, n_12348, n_12349;
wire n_12333, n_12334, n_12335, n_12336, n_12337, n_12338, n_12339, n_12340;
wire n_12323, n_12325, n_12326, n_12328, n_12329, n_12330, n_12331, n_12332;
wire n_12312, n_12313, n_12314, n_12318, n_12319, n_12320, n_12321, n_12322;
wire n_12301, n_12302, n_12304, n_12305, n_12308, n_12309, n_12310, n_12311;
wire n_12288, n_12289, n_12290, n_12291, n_12292, n_12294, n_12297, n_12299;
wire n_12279, n_12280, n_12281, n_12283, n_12284, n_12285, n_12286, n_12287;
wire n_12269, n_12270, n_12271, n_12272, n_12273, n_12274, n_12276, n_12278;
wire n_12258, n_12260, n_12261, n_12262, n_12263, n_12264, n_12266, n_12267;
wire n_12248, n_12249, n_12250, n_12251, n_12253, n_12255, n_12256, n_12257;
wire n_12239, n_12240, n_12241, n_12242, n_12243, n_12245, n_12246, n_12247;
wire n_12227, n_12228, n_12232, n_12233, n_12234, n_12235, n_12236, n_12237;
wire n_12218, n_12220, n_12221, n_12222, n_12223, n_12224, n_12225, n_12226;
wire n_12210, n_12211, n_12212, n_12213, n_12214, n_12215, n_12216, n_12217;
wire n_12198, n_12200, n_12203, n_12204, n_12206, n_12207, n_12208, n_12209;
wire n_12190, n_12191, n_12192, n_12193, n_12194, n_12195, n_12196, n_12197;
wire n_12181, n_12183, n_12184, n_12185, n_12186, n_12187, n_12188, n_12189;
wire n_12169, n_12171, n_12173, n_12174, n_12175, n_12176, n_12178, n_12180;
wire n_12157, n_12159, n_12160, n_12161, n_12163, n_12166, n_12167, n_12168;
wire n_12141, n_12142, n_12143, n_12144, n_12147, n_12151, n_12154, n_12156;
wire n_12130, n_12131, n_12133, n_12135, n_12136, n_12137, n_12138, n_12139;
wire n_12119, n_12120, n_12121, n_12122, n_12124, n_12126, n_12127, n_12128;
wire n_12111, n_12112, n_12113, n_12114, n_12115, n_12116, n_12117, n_12118;
wire n_12103, n_12104, n_12105, n_12106, n_12107, n_12108, n_12109, n_12110;
wire n_12093, n_12094, n_12096, n_12097, n_12098, n_12099, n_12100, n_12101;
wire n_12082, n_12083, n_12084, n_12086, n_12087, n_12089, n_12090, n_12091;
wire n_12070, n_12071, n_12073, n_12075, n_12077, n_12078, n_12079, n_12081;
wire n_12060, n_12061, n_12062, n_12063, n_12064, n_12066, n_12068, n_12069;
wire n_12050, n_12051, n_12052, n_12053, n_12054, n_12055, n_12056, n_12057;
wire n_12042, n_12043, n_12044, n_12045, n_12046, n_12047, n_12048, n_12049;
wire n_12033, n_12034, n_12035, n_12036, n_12037, n_12038, n_12039, n_12041;
wire n_12023, n_12025, n_12026, n_12027, n_12028, n_12029, n_12030, n_12031;
wire n_12013, n_12014, n_12015, n_12016, n_12018, n_12020, n_12021, n_12022;
wire n_12002, n_12003, n_12004, n_12005, n_12006, n_12007, n_12008, n_12009;
wire n_11993, n_11994, n_11995, n_11996, n_11997, n_11999, n_12000, n_12001;
wire n_11982, n_11985, n_11987, n_11988, n_11989, n_11990, n_11991, n_11992;
wire n_11968, n_11970, n_11971, n_11973, n_11976, n_11977, n_11978, n_11981;
wire n_11954, n_11955, n_11957, n_11958, n_11961, n_11962, n_11965, n_11966;
wire n_11936, n_11937, n_11938, n_11939, n_11940, n_11941, n_11952, n_11953;
wire n_11928, n_11929, n_11930, n_11931, n_11932, n_11933, n_11934, n_11935;
wire n_11918, n_11919, n_11920, n_11921, n_11922, n_11923, n_11925, n_11926;
wire n_11909, n_11911, n_11912, n_11913, n_11914, n_11915, n_11916, n_11917;
wire n_11899, n_11900, n_11901, n_11903, n_11904, n_11905, n_11906, n_11908;
wire n_11890, n_11891, n_11892, n_11893, n_11894, n_11896, n_11897, n_11898;
wire n_11882, n_11883, n_11884, n_11885, n_11886, n_11887, n_11888, n_11889;
wire n_11870, n_11871, n_11873, n_11874, n_11875, n_11876, n_11877, n_11880;
wire n_11862, n_11863, n_11864, n_11865, n_11866, n_11867, n_11868, n_11869;
wire n_11854, n_11855, n_11856, n_11857, n_11858, n_11859, n_11860, n_11861;
wire n_11846, n_11847, n_11848, n_11849, n_11850, n_11851, n_11852, n_11853;
wire n_11837, n_11839, n_11840, n_11841, n_11842, n_11843, n_11844, n_11845;
wire n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835, n_11836;
wire n_11820, n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827;
wire n_11812, n_11813, n_11814, n_11815, n_11816, n_11817, n_11818, n_11819;
wire n_11804, n_11805, n_11806, n_11807, n_11808, n_11809, n_11810, n_11811;
wire n_11792, n_11793, n_11797, n_11799, n_11800, n_11801, n_11802, n_11803;
wire n_11784, n_11785, n_11786, n_11787, n_11788, n_11789, n_11790, n_11791;
wire n_11776, n_11777, n_11778, n_11779, n_11780, n_11781, n_11782, n_11783;
wire n_11766, n_11769, n_11770, n_11771, n_11772, n_11773, n_11774, n_11775;
wire n_11751, n_11752, n_11756, n_11759, n_11760, n_11762, n_11763, n_11764;
wire n_11736, n_11737, n_11738, n_11740, n_11742, n_11747, n_11748, n_11750;
wire n_11720, n_11725, n_11727, n_11730, n_11731, n_11732, n_11733, n_11734;
wire n_11704, n_11705, n_11708, n_11709, n_11710, n_11712, n_11713, n_11716;
wire n_11696, n_11697, n_11698, n_11699, n_11700, n_11701, n_11702, n_11703;
wire n_11688, n_11689, n_11690, n_11691, n_11692, n_11693, n_11694, n_11695;
wire n_11677, n_11679, n_11680, n_11682, n_11683, n_11685, n_11686, n_11687;
wire n_11667, n_11668, n_11670, n_11671, n_11672, n_11674, n_11675, n_11676;
wire n_11658, n_11659, n_11660, n_11661, n_11662, n_11664, n_11665, n_11666;
wire n_11648, n_11649, n_11650, n_11651, n_11652, n_11654, n_11655, n_11657;
wire n_11640, n_11641, n_11642, n_11643, n_11644, n_11645, n_11646, n_11647;
wire n_11632, n_11633, n_11634, n_11635, n_11636, n_11637, n_11638, n_11639;
wire n_11624, n_11625, n_11626, n_11627, n_11628, n_11629, n_11630, n_11631;
wire n_11615, n_11616, n_11617, n_11619, n_11620, n_11621, n_11622, n_11623;
wire n_11607, n_11608, n_11609, n_11610, n_11611, n_11612, n_11613, n_11614;
wire n_11598, n_11599, n_11600, n_11601, n_11602, n_11604, n_11605, n_11606;
wire n_11590, n_11591, n_11592, n_11593, n_11594, n_11595, n_11596, n_11597;
wire n_11582, n_11583, n_11584, n_11585, n_11586, n_11587, n_11588, n_11589;
wire n_11574, n_11575, n_11576, n_11577, n_11578, n_11579, n_11580, n_11581;
wire n_11566, n_11567, n_11568, n_11569, n_11570, n_11571, n_11572, n_11573;
wire n_11555, n_11556, n_11558, n_11559, n_11561, n_11563, n_11564, n_11565;
wire n_11545, n_11546, n_11548, n_11549, n_11550, n_11551, n_11552, n_11553;
wire n_11536, n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544;
wire n_11526, n_11527, n_11528, n_11529, n_11530, n_11533, n_11534, n_11535;
wire n_11513, n_11515, n_11518, n_11519, n_11520, n_11521, n_11523, n_11525;
wire n_11500, n_11501, n_11503, n_11504, n_11506, n_11507, n_11508, n_11512;
wire n_11490, n_11491, n_11492, n_11493, n_11495, n_11496, n_11497, n_11498;
wire n_11481, n_11482, n_11483, n_11485, n_11486, n_11487, n_11488, n_11489;
wire n_11464, n_11468, n_11470, n_11476, n_11477, n_11478, n_11479, n_11480;
wire n_11450, n_11451, n_11452, n_11453, n_11454, n_11456, n_11457, n_11458;
wire n_11441, n_11442, n_11443, n_11445, n_11446, n_11447, n_11448, n_11449;
wire n_11433, n_11434, n_11435, n_11436, n_11437, n_11438, n_11439, n_11440;
wire n_11425, n_11426, n_11427, n_11428, n_11429, n_11430, n_11431, n_11432;
wire n_11417, n_11418, n_11419, n_11420, n_11421, n_11422, n_11423, n_11424;
wire n_11407, n_11410, n_11411, n_11412, n_11413, n_11414, n_11415, n_11416;
wire n_11396, n_11397, n_11399, n_11401, n_11402, n_11403, n_11404, n_11405;
wire n_11388, n_11389, n_11390, n_11391, n_11392, n_11393, n_11394, n_11395;
wire n_11380, n_11381, n_11382, n_11383, n_11384, n_11385, n_11386, n_11387;
wire n_11372, n_11373, n_11374, n_11375, n_11376, n_11377, n_11378, n_11379;
wire n_11364, n_11365, n_11366, n_11367, n_11368, n_11369, n_11370, n_11371;
wire n_11356, n_11357, n_11358, n_11359, n_11360, n_11361, n_11362, n_11363;
wire n_11348, n_11349, n_11350, n_11351, n_11352, n_11353, n_11354, n_11355;
wire n_11340, n_11341, n_11342, n_11343, n_11344, n_11345, n_11346, n_11347;
wire n_11327, n_11328, n_11329, n_11330, n_11333, n_11334, n_11338, n_11339;
wire n_11318, n_11319, n_11320, n_11321, n_11322, n_11324, n_11325, n_11326;
wire n_11309, n_11310, n_11311, n_11312, n_11313, n_11314, n_11315, n_11317;
wire n_11301, n_11302, n_11303, n_11304, n_11305, n_11306, n_11307, n_11308;
wire n_11290, n_11293, n_11294, n_11295, n_11296, n_11297, n_11299, n_11300;
wire n_11277, n_11278, n_11280, n_11281, n_11283, n_11285, n_11286, n_11288;
wire n_11266, n_11267, n_11268, n_11269, n_11272, n_11274, n_11275, n_11276;
wire n_11253, n_11254, n_11256, n_11258, n_11260, n_11261, n_11264, n_11265;
wire n_11222, n_11226, n_11227, n_11245, n_11246, n_11247, n_11249, n_11250;
wire n_11207, n_11208, n_11209, n_11210, n_11211, n_11213, n_11215, n_11218;
wire n_11198, n_11199, n_11200, n_11201, n_11202, n_11203, n_11205, n_11206;
wire n_11188, n_11190, n_11191, n_11192, n_11194, n_11195, n_11196, n_11197;
wire n_11179, n_11181, n_11182, n_11183, n_11184, n_11185, n_11186, n_11187;
wire n_11171, n_11172, n_11173, n_11174, n_11175, n_11176, n_11177, n_11178;
wire n_11163, n_11164, n_11165, n_11166, n_11167, n_11168, n_11169, n_11170;
wire n_11155, n_11156, n_11157, n_11158, n_11159, n_11160, n_11161, n_11162;
wire n_11147, n_11148, n_11149, n_11150, n_11151, n_11152, n_11153, n_11154;
wire n_11137, n_11138, n_11139, n_11140, n_11141, n_11143, n_11144, n_11146;
wire n_11121, n_11122, n_11124, n_11129, n_11130, n_11134, n_11135, n_11136;
wire n_11110, n_11111, n_11112, n_11113, n_11116, n_11117, n_11118, n_11120;
wire n_11097, n_11098, n_11099, n_11101, n_11104, n_11105, n_11107, n_11109;
wire n_11079, n_11080, n_11086, n_11087, n_11088, n_11089, n_11092, n_11096;
wire n_11069, n_11070, n_11072, n_11074, n_11075, n_11076, n_11077, n_11078;
wire n_11058, n_11060, n_11061, n_11062, n_11063, n_11064, n_11065, n_11066;
wire n_11047, n_11048, n_11050, n_11051, n_11052, n_11053, n_11055, n_11057;
wire n_11036, n_11037, n_11040, n_11042, n_11043, n_11044, n_11045, n_11046;
wire n_11008, n_11009, n_11010, n_11012, n_11022, n_11030, n_11033, n_11034;
wire n_10990, n_10991, n_10998, n_10999, n_11002, n_11003, n_11006, n_11007;
wire n_10982, n_10983, n_10984, n_10985, n_10986, n_10987, n_10988, n_10989;
wire n_10974, n_10975, n_10976, n_10977, n_10978, n_10979, n_10980, n_10981;
wire n_10966, n_10967, n_10968, n_10969, n_10970, n_10971, n_10972, n_10973;
wire n_10958, n_10959, n_10960, n_10961, n_10962, n_10963, n_10964, n_10965;
wire n_10950, n_10951, n_10952, n_10953, n_10954, n_10955, n_10956, n_10957;
wire n_10942, n_10943, n_10944, n_10945, n_10946, n_10947, n_10948, n_10949;
wire n_10934, n_10935, n_10936, n_10937, n_10938, n_10939, n_10940, n_10941;
wire n_10925, n_10926, n_10927, n_10929, n_10930, n_10931, n_10932, n_10933;
wire n_10917, n_10918, n_10919, n_10920, n_10921, n_10922, n_10923, n_10924;
wire n_10909, n_10910, n_10911, n_10912, n_10913, n_10914, n_10915, n_10916;
wire n_10898, n_10899, n_10901, n_10903, n_10905, n_10906, n_10907, n_10908;
wire n_10884, n_10885, n_10886, n_10887, n_10889, n_10890, n_10893, n_10897;
wire n_10871, n_10872, n_10873, n_10874, n_10875, n_10879, n_10880, n_10882;
wire n_10854, n_10856, n_10858, n_10859, n_10860, n_10862, n_10865, n_10868;
wire n_10840, n_10841, n_10843, n_10847, n_10848, n_10851, n_10852, n_10853;
wire n_10829, n_10831, n_10833, n_10834, n_10836, n_10837, n_10838, n_10839;
wire n_10800, n_10808, n_10819, n_10821, n_10822, n_10823, n_10825, n_10826;
wire n_10790, n_10792, n_10793, n_10794, n_10795, n_10796, n_10797, n_10799;
wire n_10768, n_10769, n_10770, n_10771, n_10774, n_10776, n_10779, n_10785;
wire n_10758, n_10759, n_10760, n_10761, n_10763, n_10764, n_10765, n_10767;
wire n_10746, n_10747, n_10752, n_10753, n_10754, n_10755, n_10756, n_10757;
wire n_10736, n_10737, n_10739, n_10740, n_10741, n_10743, n_10744, n_10745;
wire n_10710, n_10711, n_10712, n_10713, n_10716, n_10717, n_10718, n_10734;
wire n_10691, n_10693, n_10696, n_10697, n_10699, n_10706, n_10708, n_10709;
wire n_10676, n_10678, n_10680, n_10682, n_10684, n_10686, n_10688, n_10689;
wire n_10658, n_10665, n_10666, n_10667, n_10669, n_10671, n_10672, n_10675;
wire n_10645, n_10646, n_10647, n_10648, n_10653, n_10655, n_10656, n_10657;
wire n_10637, n_10638, n_10639, n_10640, n_10641, n_10642, n_10643, n_10644;
wire n_10626, n_10627, n_10628, n_10629, n_10630, n_10631, n_10634, n_10635;
wire n_10616, n_10617, n_10619, n_10621, n_10622, n_10623, n_10624, n_10625;
wire n_10606, n_10607, n_10608, n_10610, n_10611, n_10612, n_10613, n_10615;
wire n_10594, n_10596, n_10597, n_10600, n_10601, n_10602, n_10603, n_10604;
wire n_10582, n_10583, n_10586, n_10587, n_10588, n_10589, n_10590, n_10593;
wire n_10573, n_10574, n_10575, n_10576, n_10577, n_10578, n_10580, n_10581;
wire n_10561, n_10562, n_10563, n_10565, n_10566, n_10569, n_10570, n_10571;
wire n_10550, n_10551, n_10552, n_10553, n_10554, n_10555, n_10556, n_10557;
wire n_10517, n_10525, n_10540, n_10542, n_10543, n_10545, n_10546, n_10548;
wire n_10487, n_10489, n_10490, n_10491, n_10497, n_10504, n_10505, n_10514;
wire n_10476, n_10477, n_10478, n_10480, n_10481, n_10482, n_10484, n_10485;
wire n_10465, n_10466, n_10467, n_10468, n_10470, n_10472, n_10474, n_10475;
wire n_10456, n_10457, n_10458, n_10459, n_10460, n_10461, n_10463, n_10464;
wire n_10447, n_10448, n_10449, n_10450, n_10451, n_10452, n_10453, n_10455;
wire n_10433, n_10435, n_10436, n_10440, n_10441, n_10443, n_10444, n_10445;
wire n_10418, n_10420, n_10423, n_10426, n_10427, n_10429, n_10431, n_10432;
wire n_10405, n_10406, n_10407, n_10409, n_10413, n_10414, n_10415, n_10416;
wire n_10395, n_10397, n_10398, n_10399, n_10400, n_10401, n_10402, n_10403;
wire n_10383, n_10384, n_10385, n_10389, n_10390, n_10392, n_10393, n_10394;
wire n_10370, n_10372, n_10373, n_10375, n_10376, n_10378, n_10379, n_10381;
wire n_10361, n_10362, n_10363, n_10364, n_10366, n_10367, n_10368, n_10369;
wire n_10351, n_10352, n_10354, n_10355, n_10356, n_10357, n_10358, n_10360;
wire n_10334, n_10335, n_10342, n_10343, n_10345, n_10346, n_10348, n_10349;
wire n_10322, n_10324, n_10325, n_10326, n_10329, n_10330, n_10331, n_10333;
wire n_10312, n_10314, n_10315, n_10316, n_10317, n_10318, n_10319, n_10320;
wire n_10283, n_10286, n_10287, n_10289, n_10292, n_10299, n_10303, n_10309;
wire n_10272, n_10273, n_10274, n_10275, n_10276, n_10277, n_10278, n_10279;
wire n_10261, n_10262, n_10263, n_10264, n_10267, n_10268, n_10270, n_10271;
wire n_10251, n_10253, n_10254, n_10256, n_10257, n_10258, n_10259, n_10260;
wire n_10240, n_10242, n_10244, n_10245, n_10246, n_10247, n_10248, n_10249;
wire n_10224, n_10225, n_10228, n_10230, n_10232, n_10234, n_10236, n_10238;
wire n_10215, n_10217, n_10218, n_10219, n_10220, n_10221, n_10222, n_10223;
wire n_10204, n_10205, n_10206, n_10208, n_10210, n_10211, n_10212, n_10214;
wire n_10192, n_10196, n_10197, n_10198, n_10200, n_10201, n_10202, n_10203;
wire n_10181, n_10182, n_10183, n_10187, n_10188, n_10189, n_10190, n_10191;
wire n_10173, n_10174, n_10175, n_10176, n_10177, n_10178, n_10179, n_10180;
wire n_10165, n_10166, n_10167, n_10168, n_10169, n_10170, n_10171, n_10172;
wire n_10157, n_10158, n_10159, n_10160, n_10161, n_10162, n_10163, n_10164;
wire n_10149, n_10150, n_10151, n_10152, n_10153, n_10154, n_10155, n_10156;
wire n_10139, n_10140, n_10141, n_10143, n_10144, n_10145, n_10147, n_10148;
wire n_10129, n_10131, n_10133, n_10134, n_10135, n_10136, n_10137, n_10138;
wire n_10119, n_10120, n_10122, n_10123, n_10124, n_10126, n_10127, n_10128;
wire n_10110, n_10111, n_10112, n_10113, n_10114, n_10115, n_10116, n_10117;
wire n_10097, n_10098, n_10100, n_10102, n_10103, n_10104, n_10105, n_10108;
wire n_10088, n_10089, n_10090, n_10092, n_10093, n_10094, n_10095, n_10096;
wire n_10074, n_10076, n_10079, n_10080, n_10081, n_10082, n_10083, n_10084;
wire n_10059, n_10061, n_10063, n_10064, n_10066, n_10067, n_10069, n_10071;
wire n_10047, n_10048, n_10049, n_10050, n_10052, n_10053, n_10056, n_10057;
wire n_10037, n_10038, n_10040, n_10041, n_10042, n_10043, n_10044, n_10046;
wire n_10023, n_10030, n_10031, n_10032, n_10033, n_10034, n_10035, n_10036;
wire n_9997, n_9998, n_10002, n_10003, n_10006, n_10014, n_10020, n_10021;
wire n_9962, n_9963, n_9964, n_9971, n_9978, n_9983, n_9994, n_9995;
wire n_9947, n_9953, n_9955, n_9956, n_9958, n_9959, n_9960, n_9961;
wire n_9938, n_9939, n_9940, n_9942, n_9943, n_9944, n_9945, n_9946;
wire n_9930, n_9931, n_9932, n_9933, n_9934, n_9935, n_9936, n_9937;
wire n_9921, n_9922, n_9923, n_9924, n_9925, n_9927, n_9928, n_9929;
wire n_9909, n_9910, n_9911, n_9912, n_9916, n_9917, n_9919, n_9920;
wire n_9899, n_9900, n_9902, n_9903, n_9905, n_9906, n_9907, n_9908;
wire n_9890, n_9891, n_9893, n_9894, n_9895, n_9896, n_9897, n_9898;
wire n_9879, n_9880, n_9881, n_9882, n_9883, n_9887, n_9888, n_9889;
wire n_9867, n_9868, n_9869, n_9871, n_9873, n_9875, n_9876, n_9878;
wire n_9858, n_9859, n_9860, n_9861, n_9862, n_9863, n_9864, n_9866;
wire n_9850, n_9851, n_9852, n_9853, n_9854, n_9855, n_9856, n_9857;
wire n_9842, n_9843, n_9844, n_9845, n_9846, n_9847, n_9848, n_9849;
wire n_9834, n_9835, n_9836, n_9837, n_9838, n_9839, n_9840, n_9841;
wire n_9823, n_9825, n_9826, n_9827, n_9828, n_9830, n_9832, n_9833;
wire n_9813, n_9814, n_9815, n_9816, n_9818, n_9819, n_9820, n_9822;
wire n_9803, n_9804, n_9806, n_9807, n_9809, n_9810, n_9811, n_9812;
wire n_9793, n_9794, n_9795, n_9797, n_9798, n_9800, n_9801, n_9802;
wire n_9778, n_9780, n_9783, n_9785, n_9788, n_9789, n_9791, n_9792;
wire n_9769, n_9770, n_9771, n_9772, n_9773, n_9774, n_9775, n_9776;
wire n_9755, n_9758, n_9760, n_9761, n_9763, n_9765, n_9766, n_9767;
wire n_9742, n_9744, n_9745, n_9746, n_9748, n_9749, n_9752, n_9754;
wire n_9722, n_9725, n_9726, n_9729, n_9730, n_9733, n_9738, n_9741;
wire n_9709, n_9710, n_9711, n_9713, n_9714, n_9718, n_9719, n_9720;
wire n_9698, n_9699, n_9700, n_9701, n_9703, n_9704, n_9706, n_9708;
wire n_9684, n_9687, n_9688, n_9689, n_9691, n_9692, n_9693, n_9695;
wire n_9673, n_9674, n_9675, n_9676, n_9677, n_9679, n_9682, n_9683;
wire n_9665, n_9666, n_9667, n_9668, n_9669, n_9670, n_9671, n_9672;
wire n_9653, n_9654, n_9655, n_9657, n_9658, n_9659, n_9662, n_9663;
wire n_9644, n_9645, n_9646, n_9647, n_9648, n_9650, n_9651, n_9652;
wire n_9635, n_9637, n_9638, n_9639, n_9640, n_9641, n_9642, n_9643;
wire n_9625, n_9626, n_9627, n_9628, n_9629, n_9631, n_9632, n_9634;
wire n_9615, n_9616, n_9617, n_9618, n_9621, n_9622, n_9623, n_9624;
wire n_9606, n_9607, n_9608, n_9609, n_9610, n_9612, n_9613, n_9614;
wire n_9597, n_9598, n_9599, n_9601, n_9602, n_9603, n_9604, n_9605;
wire n_9587, n_9589, n_9590, n_9591, n_9592, n_9594, n_9595, n_9596;
wire n_9575, n_9577, n_9578, n_9580, n_9581, n_9583, n_9585, n_9586;
wire n_9562, n_9563, n_9565, n_9566, n_9567, n_9569, n_9571, n_9573;
wire n_9553, n_9554, n_9555, n_9556, n_9557, n_9558, n_9559, n_9561;
wire n_9544, n_9546, n_9547, n_9548, n_9549, n_9550, n_9551, n_9552;
wire n_9529, n_9530, n_9531, n_9532, n_9534, n_9538, n_9541, n_9542;
wire n_9520, n_9521, n_9522, n_9523, n_9524, n_9525, n_9527, n_9528;
wire n_9511, n_9512, n_9513, n_9514, n_9515, n_9516, n_9517, n_9519;
wire n_9502, n_9503, n_9505, n_9506, n_9507, n_9508, n_9509, n_9510;
wire n_9475, n_9476, n_9482, n_9483, n_9490, n_9493, n_9495, n_9498;
wire n_9431, n_9435, n_9436, n_9441, n_9455, n_9458, n_9473, n_9474;
wire n_9421, n_9422, n_9424, n_9425, n_9426, n_9428, n_9429, n_9430;
wire n_9392, n_9404, n_9413, n_9415, n_9416, n_9418, n_9419, n_9420;
wire n_9383, n_9384, n_9385, n_9386, n_9387, n_9388, n_9390, n_9391;
wire n_9374, n_9375, n_9377, n_9378, n_9379, n_9380, n_9381, n_9382;
wire n_9363, n_9364, n_9366, n_9368, n_9369, n_9371, n_9372, n_9373;
wire n_9354, n_9355, n_9356, n_9357, n_9358, n_9360, n_9361, n_9362;
wire n_9346, n_9347, n_9348, n_9349, n_9350, n_9351, n_9352, n_9353;
wire n_9336, n_9337, n_9338, n_9340, n_9341, n_9342, n_9343, n_9345;
wire n_9322, n_9327, n_9329, n_9331, n_9332, n_9333, n_9334, n_9335;
wire n_9309, n_9310, n_9311, n_9313, n_9314, n_9318, n_9320, n_9321;
wire n_9297, n_9298, n_9299, n_9300, n_9302, n_9303, n_9307, n_9308;
wire n_9285, n_9286, n_9288, n_9290, n_9291, n_9292, n_9294, n_9295;
wire n_9274, n_9276, n_9277, n_9278, n_9279, n_9280, n_9281, n_9284;
wire n_9257, n_9260, n_9262, n_9263, n_9264, n_9268, n_9269, n_9272;
wire n_9239, n_9240, n_9242, n_9243, n_9247, n_9249, n_9252, n_9253;
wire n_9230, n_9231, n_9232, n_9234, n_9235, n_9236, n_9237, n_9238;
wire n_9211, n_9212, n_9219, n_9223, n_9225, n_9226, n_9227, n_9228;
wire n_9201, n_9203, n_9204, n_9205, n_9206, n_9207, n_9209, n_9210;
wire n_9186, n_9188, n_9190, n_9194, n_9195, n_9197, n_9198, n_9199;
wire n_9177, n_9178, n_9179, n_9180, n_9181, n_9182, n_9184, n_9185;
wire n_9165, n_9166, n_9167, n_9169, n_9171, n_9172, n_9173, n_9176;
wire n_9146, n_9149, n_9152, n_9154, n_9159, n_9161, n_9162, n_9163;
wire n_9135, n_9136, n_9137, n_9139, n_9141, n_9142, n_9143, n_9145;
wire n_9125, n_9126, n_9127, n_9128, n_9130, n_9131, n_9132, n_9133;
wire n_9114, n_9117, n_9119, n_9120, n_9121, n_9122, n_9123, n_9124;
wire n_9103, n_9104, n_9105, n_9106, n_9108, n_9109, n_9110, n_9111;
wire n_9094, n_9095, n_9096, n_9097, n_9099, n_9100, n_9101, n_9102;
wire n_9086, n_9087, n_9088, n_9089, n_9090, n_9091, n_9092, n_9093;
wire n_9077, n_9078, n_9079, n_9080, n_9081, n_9082, n_9083, n_9085;
wire n_9066, n_9067, n_9068, n_9071, n_9072, n_9073, n_9074, n_9076;
wire n_9058, n_9059, n_9060, n_9061, n_9062, n_9063, n_9064, n_9065;
wire n_9050, n_9051, n_9052, n_9053, n_9054, n_9055, n_9056, n_9057;
wire n_9042, n_9043, n_9044, n_9045, n_9046, n_9047, n_9048, n_9049;
wire n_9032, n_9034, n_9035, n_9036, n_9038, n_9039, n_9040, n_9041;
wire n_9023, n_9024, n_9025, n_9026, n_9027, n_9028, n_9030, n_9031;
wire n_9014, n_9015, n_9016, n_9017, n_9018, n_9019, n_9020, n_9021;
wire n_8996, n_8998, n_9001, n_9003, n_9009, n_9010, n_9011, n_9013;
wire n_8965, n_8966, n_8977, n_8979, n_8980, n_8981, n_8989, n_8990;
wire n_8942, n_8945, n_8946, n_8947, n_8948, n_8949, n_8954, n_8958;
wire n_8922, n_8925, n_8927, n_8933, n_8934, n_8935, n_8936, n_8940;
wire n_8909, n_8910, n_8911, n_8912, n_8914, n_8915, n_8916, n_8917;
wire n_8897, n_8898, n_8899, n_8900, n_8901, n_8903, n_8905, n_8906;
wire n_8889, n_8890, n_8891, n_8892, n_8893, n_8894, n_8895, n_8896;
wire n_8881, n_8882, n_8883, n_8884, n_8885, n_8886, n_8887, n_8888;
wire n_8872, n_8873, n_8874, n_8875, n_8876, n_8877, n_8878, n_8880;
wire n_8862, n_8864, n_8865, n_8867, n_8868, n_8869, n_8870, n_8871;
wire n_8851, n_8853, n_8856, n_8857, n_8858, n_8859, n_8860, n_8861;
wire n_8842, n_8843, n_8844, n_8845, n_8846, n_8847, n_8849, n_8850;
wire n_8832, n_8833, n_8835, n_8837, n_8838, n_8839, n_8840, n_8841;
wire n_8824, n_8825, n_8826, n_8827, n_8828, n_8829, n_8830, n_8831;
wire n_8816, n_8817, n_8818, n_8819, n_8820, n_8821, n_8822, n_8823;
wire n_8803, n_8809, n_8810, n_8811, n_8812, n_8813, n_8814, n_8815;
wire n_8794, n_8795, n_8796, n_8797, n_8798, n_8799, n_8801, n_8802;
wire n_8784, n_8785, n_8787, n_8788, n_8790, n_8791, n_8792, n_8793;
wire n_8776, n_8777, n_8778, n_8779, n_8780, n_8781, n_8782, n_8783;
wire n_8754, n_8755, n_8756, n_8757, n_8758, n_8759, n_8761, n_8762;
wire n_8744, n_8745, n_8746, n_8747, n_8749, n_8750, n_8752, n_8753;
wire n_8736, n_8737, n_8738, n_8739, n_8740, n_8741, n_8742, n_8743;
wire n_8718, n_8719, n_8721, n_8726, n_8729, n_8732, n_8734, n_8735;
wire n_8705, n_8709, n_8710, n_8711, n_8713, n_8714, n_8715, n_8716;
wire n_8692, n_8693, n_8695, n_8696, n_8697, n_8699, n_8703, n_8704;
wire n_8672, n_8677, n_8678, n_8679, n_8680, n_8682, n_8686, n_8687;
wire n_8641, n_8642, n_8643, n_8644, n_8661, n_8664, n_8668, n_8671;
wire n_8616, n_8618, n_8619, n_8622, n_8623, n_8625, n_8633, n_8635;
wire n_8606, n_8609, n_8610, n_8611, n_8612, n_8613, n_8614, n_8615;
wire n_8598, n_8599, n_8600, n_8601, n_8602, n_8603, n_8604, n_8605;
wire n_8588, n_8589, n_8591, n_8592, n_8593, n_8595, n_8596, n_8597;
wire n_8579, n_8580, n_8581, n_8582, n_8584, n_8585, n_8586, n_8587;
wire n_8571, n_8572, n_8573, n_8574, n_8575, n_8576, n_8577, n_8578;
wire n_8561, n_8562, n_8564, n_8565, n_8566, n_8567, n_8568, n_8569;
wire n_8553, n_8554, n_8555, n_8556, n_8557, n_8558, n_8559, n_8560;
wire n_8542, n_8544, n_8545, n_8547, n_8549, n_8550, n_8551, n_8552;
wire n_8526, n_8527, n_8528, n_8534, n_8535, n_8537, n_8540, n_8541;
wire n_8515, n_8516, n_8517, n_8518, n_8522, n_8523, n_8524, n_8525;
wire n_8485, n_8486, n_8492, n_8493, n_8505, n_8511, n_8512, n_8513;
wire n_8469, n_8470, n_8471, n_8472, n_8473, n_8474, n_8479, n_8484;
wire n_8457, n_8458, n_8460, n_8462, n_8464, n_8465, n_8467, n_8468;
wire n_8447, n_8448, n_8449, n_8451, n_8452, n_8453, n_8454, n_8455;
wire n_8438, n_8440, n_8441, n_8442, n_8443, n_8444, n_8445, n_8446;
wire n_8429, n_8430, n_8431, n_8432, n_8433, n_8434, n_8435, n_8436;
wire n_8420, n_8421, n_8422, n_8424, n_8425, n_8426, n_8427, n_8428;
wire n_8408, n_8409, n_8410, n_8412, n_8413, n_8416, n_8417, n_8418;
wire n_8393, n_8394, n_8395, n_8397, n_8399, n_8400, n_8401, n_8407;
wire n_8379, n_8380, n_8381, n_8382, n_8384, n_8387, n_8390, n_8392;
wire n_8370, n_8371, n_8372, n_8374, n_8375, n_8376, n_8377, n_8378;
wire n_8360, n_8361, n_8363, n_8364, n_8365, n_8366, n_8367, n_8369;
wire n_8350, n_8351, n_8352, n_8354, n_8355, n_8356, n_8357, n_8358;
wire n_8336, n_8337, n_8340, n_8343, n_8344, n_8345, n_8346, n_8347;
wire n_8326, n_8329, n_8330, n_8331, n_8332, n_8333, n_8334, n_8335;
wire n_8314, n_8316, n_8319, n_8320, n_8321, n_8322, n_8324, n_8325;
wire n_8293, n_8295, n_8303, n_8304, n_8305, n_8306, n_8309, n_8313;
wire n_8279, n_8280, n_8281, n_8283, n_8284, n_8285, n_8286, n_8291;
wire n_8267, n_8269, n_8270, n_8272, n_8273, n_8274, n_8275, n_8277;
wire n_8258, n_8259, n_8260, n_8261, n_8262, n_8263, n_8264, n_8266;
wire n_8249, n_8250, n_8251, n_8252, n_8254, n_8255, n_8256, n_8257;
wire n_8241, n_8242, n_8243, n_8244, n_8245, n_8246, n_8247, n_8248;
wire n_8232, n_8233, n_8234, n_8235, n_8236, n_8238, n_8239, n_8240;
wire n_8214, n_8224, n_8225, n_8226, n_8228, n_8229, n_8230, n_8231;
wire n_8205, n_8206, n_8207, n_8208, n_8209, n_8210, n_8212, n_8213;
wire n_8196, n_8197, n_8198, n_8199, n_8200, n_8202, n_8203, n_8204;
wire n_8188, n_8189, n_8190, n_8191, n_8192, n_8193, n_8194, n_8195;
wire n_8178, n_8179, n_8181, n_8182, n_8183, n_8185, n_8186, n_8187;
wire n_8169, n_8170, n_8172, n_8173, n_8174, n_8175, n_8176, n_8177;
wire n_8157, n_8158, n_8162, n_8163, n_8164, n_8165, n_8166, n_8168;
wire n_8149, n_8150, n_8151, n_8152, n_8153, n_8154, n_8155, n_8156;
wire n_8141, n_8142, n_8143, n_8144, n_8145, n_8146, n_8147, n_8148;
wire n_8132, n_8134, n_8135, n_8136, n_8137, n_8138, n_8139, n_8140;
wire n_8121, n_8122, n_8124, n_8125, n_8128, n_8129, n_8130, n_8131;
wire n_8109, n_8112, n_8113, n_8114, n_8115, n_8116, n_8117, n_8119;
wire n_8090, n_8093, n_8096, n_8099, n_8102, n_8103, n_8105, n_8106;
wire n_8078, n_8079, n_8080, n_8082, n_8083, n_8084, n_8085, n_8086;
wire n_8058, n_8059, n_8060, n_8065, n_8066, n_8070, n_8074, n_8075;
wire n_8048, n_8049, n_8050, n_8051, n_8052, n_8054, n_8055, n_8056;
wire n_8032, n_8033, n_8034, n_8035, n_8036, n_8037, n_8039, n_8047;
wire n_8016, n_8020, n_8022, n_8023, n_8024, n_8027, n_8029, n_8031;
wire n_8007, n_8008, n_8009, n_8010, n_8011, n_8013, n_8014, n_8015;
wire n_7997, n_7998, n_8000, n_8001, n_8002, n_8003, n_8004, n_8005;
wire n_7984, n_7985, n_7986, n_7987, n_7988, n_7992, n_7993, n_7994;
wire n_7972, n_7973, n_7975, n_7976, n_7977, n_7978, n_7981, n_7983;
wire n_7961, n_7962, n_7963, n_7964, n_7966, n_7967, n_7970, n_7971;
wire n_7953, n_7954, n_7955, n_7956, n_7957, n_7958, n_7959, n_7960;
wire n_7939, n_7940, n_7942, n_7943, n_7944, n_7945, n_7949, n_7952;
wire n_7930, n_7932, n_7933, n_7934, n_7935, n_7936, n_7937, n_7938;
wire n_7921, n_7923, n_7924, n_7925, n_7926, n_7927, n_7928, n_7929;
wire n_7912, n_7914, n_7915, n_7916, n_7917, n_7918, n_7919, n_7920;
wire n_7903, n_7904, n_7905, n_7906, n_7907, n_7909, n_7910, n_7911;
wire n_7894, n_7895, n_7896, n_7897, n_7898, n_7900, n_7901, n_7902;
wire n_7885, n_7886, n_7887, n_7888, n_7890, n_7891, n_7892, n_7893;
wire n_7877, n_7878, n_7879, n_7880, n_7881, n_7882, n_7883, n_7884;
wire n_7863, n_7864, n_7865, n_7869, n_7870, n_7871, n_7873, n_7876;
wire n_7850, n_7851, n_7852, n_7856, n_7858, n_7859, n_7860, n_7862;
wire n_7841, n_7842, n_7843, n_7844, n_7845, n_7847, n_7848, n_7849;
wire n_7830, n_7832, n_7833, n_7834, n_7836, n_7838, n_7839, n_7840;
wire n_7819, n_7820, n_7821, n_7822, n_7823, n_7827, n_7828, n_7829;
wire n_7809, n_7810, n_7811, n_7812, n_7813, n_7814, n_7815, n_7816;
wire n_7796, n_7797, n_7798, n_7799, n_7804, n_7805, n_7806, n_7807;
wire n_7785, n_7786, n_7787, n_7788, n_7789, n_7791, n_7793, n_7794;
wire n_7775, n_7776, n_7777, n_7778, n_7779, n_7781, n_7782, n_7783;
wire n_7766, n_7767, n_7769, n_7770, n_7771, n_7772, n_7773, n_7774;
wire n_7756, n_7758, n_7759, n_7760, n_7761, n_7762, n_7763, n_7764;
wire n_7747, n_7748, n_7749, n_7750, n_7752, n_7753, n_7754, n_7755;
wire n_7738, n_7739, n_7740, n_7741, n_7743, n_7744, n_7745, n_7746;
wire n_7730, n_7731, n_7732, n_7733, n_7734, n_7735, n_7736, n_7737;
wire n_7720, n_7721, n_7722, n_7723, n_7724, n_7725, n_7727, n_7728;
wire n_7711, n_7712, n_7713, n_7714, n_7715, n_7716, n_7717, n_7719;
wire n_7699, n_7700, n_7701, n_7702, n_7703, n_7704, n_7705, n_7706;
wire n_7691, n_7692, n_7693, n_7694, n_7695, n_7696, n_7697, n_7698;
wire n_7681, n_7682, n_7683, n_7684, n_7685, n_7686, n_7687, n_7689;
wire n_7673, n_7674, n_7675, n_7676, n_7677, n_7678, n_7679, n_7680;
wire n_7664, n_7665, n_7666, n_7668, n_7669, n_7670, n_7671, n_7672;
wire n_7656, n_7657, n_7658, n_7659, n_7660, n_7661, n_7662, n_7663;
wire n_7646, n_7647, n_7648, n_7649, n_7651, n_7653, n_7654, n_7655;
wire n_7635, n_7636, n_7637, n_7638, n_7639, n_7640, n_7641, n_7644;
wire n_7625, n_7626, n_7628, n_7629, n_7630, n_7631, n_7633, n_7634;
wire n_7616, n_7617, n_7618, n_7619, n_7620, n_7622, n_7623, n_7624;
wire n_7607, n_7608, n_7609, n_7610, n_7612, n_7613, n_7614, n_7615;
wire n_7595, n_7596, n_7597, n_7598, n_7602, n_7603, n_7604, n_7606;
wire n_7584, n_7586, n_7587, n_7590, n_7591, n_7592, n_7593, n_7594;
wire n_7572, n_7573, n_7574, n_7575, n_7578, n_7580, n_7581, n_7582;
wire n_7563, n_7565, n_7566, n_7567, n_7568, n_7569, n_7570, n_7571;
wire n_7552, n_7553, n_7555, n_7556, n_7558, n_7559, n_7561, n_7562;
wire n_7543, n_7544, n_7545, n_7546, n_7547, n_7549, n_7550, n_7551;
wire n_7533, n_7534, n_7535, n_7536, n_7538, n_7539, n_7540, n_7541;
wire n_7524, n_7525, n_7526, n_7527, n_7528, n_7530, n_7531, n_7532;
wire n_7515, n_7516, n_7517, n_7519, n_7520, n_7521, n_7522, n_7523;
wire n_7504, n_7505, n_7507, n_7509, n_7510, n_7512, n_7513, n_7514;
wire n_7496, n_7497, n_7498, n_7499, n_7500, n_7501, n_7502, n_7503;
wire n_7488, n_7489, n_7490, n_7491, n_7492, n_7493, n_7494, n_7495;
wire n_7478, n_7479, n_7480, n_7481, n_7482, n_7483, n_7484, n_7485;
wire n_7470, n_7471, n_7472, n_7473, n_7474, n_7475, n_7476, n_7477;
wire n_7461, n_7462, n_7463, n_7465, n_7466, n_7467, n_7468, n_7469;
wire n_7445, n_7452, n_7454, n_7455, n_7457, n_7458, n_7459, n_7460;
wire n_7436, n_7437, n_7438, n_7440, n_7441, n_7442, n_7443, n_7444;
wire n_7428, n_7429, n_7430, n_7431, n_7432, n_7433, n_7434, n_7435;
wire n_7415, n_7417, n_7418, n_7419, n_7420, n_7422, n_7426, n_7427;
wire n_7403, n_7404, n_7405, n_7406, n_7407, n_7408, n_7411, n_7414;
wire n_7395, n_7396, n_7397, n_7398, n_7399, n_7400, n_7401, n_7402;
wire n_7385, n_7386, n_7387, n_7389, n_7390, n_7391, n_7393, n_7394;
wire n_7374, n_7375, n_7376, n_7378, n_7379, n_7380, n_7381, n_7383;
wire n_7363, n_7364, n_7367, n_7368, n_7369, n_7370, n_7372, n_7373;
wire n_7353, n_7354, n_7355, n_7358, n_7359, n_7360, n_7361, n_7362;
wire n_7344, n_7345, n_7346, n_7347, n_7348, n_7349, n_7351, n_7352;
wire n_7335, n_7337, n_7338, n_7339, n_7340, n_7341, n_7342, n_7343;
wire n_7326, n_7327, n_7328, n_7329, n_7331, n_7332, n_7333, n_7334;
wire n_7317, n_7318, n_7319, n_7320, n_7321, n_7322, n_7323, n_7325;
wire n_7309, n_7310, n_7311, n_7312, n_7313, n_7314, n_7315, n_7316;
wire n_7298, n_7299, n_7301, n_7302, n_7305, n_7306, n_7307, n_7308;
wire n_7286, n_7287, n_7289, n_7290, n_7291, n_7293, n_7295, n_7297;
wire n_7275, n_7276, n_7278, n_7279, n_7280, n_7283, n_7284, n_7285;
wire n_7262, n_7266, n_7267, n_7268, n_7269, n_7270, n_7272, n_7273;
wire n_7252, n_7253, n_7254, n_7255, n_7257, n_7258, n_7259, n_7260;
wire n_7241, n_7242, n_7243, n_7244, n_7245, n_7246, n_7249, n_7250;
wire n_7231, n_7232, n_7233, n_7236, n_7237, n_7238, n_7239, n_7240;
wire n_7219, n_7221, n_7222, n_7224, n_7225, n_7227, n_7228, n_7230;
wire n_7209, n_7210, n_7212, n_7213, n_7214, n_7216, n_7217, n_7218;
wire n_7201, n_7202, n_7203, n_7204, n_7205, n_7206, n_7207, n_7208;
wire n_7193, n_7194, n_7195, n_7196, n_7197, n_7198, n_7199, n_7200;
wire n_7183, n_7186, n_7187, n_7188, n_7189, n_7190, n_7191, n_7192;
wire n_7172, n_7173, n_7175, n_7177, n_7179, n_7180, n_7181, n_7182;
wire n_7162, n_7163, n_7165, n_7166, n_7168, n_7169, n_7170, n_7171;
wire n_7154, n_7155, n_7156, n_7157, n_7158, n_7159, n_7160, n_7161;
wire n_7145, n_7146, n_7148, n_7149, n_7150, n_7151, n_7152, n_7153;
wire n_7135, n_7136, n_7137, n_7139, n_7140, n_7142, n_7143, n_7144;
wire n_7125, n_7126, n_7127, n_7128, n_7131, n_7132, n_7133, n_7134;
wire n_7116, n_7118, n_7119, n_7120, n_7121, n_7122, n_7123, n_7124;
wire n_7106, n_7107, n_7109, n_7110, n_7111, n_7112, n_7113, n_7115;
wire n_7092, n_7094, n_7096, n_7098, n_7102, n_7103, n_7104, n_7105;
wire n_7082, n_7083, n_7084, n_7085, n_7086, n_7088, n_7090, n_7091;
wire n_7073, n_7074, n_7075, n_7076, n_7077, n_7078, n_7079, n_7081;
wire n_7058, n_7059, n_7062, n_7065, n_7066, n_7068, n_7069, n_7071;
wire n_7049, n_7050, n_7051, n_7052, n_7053, n_7054, n_7055, n_7057;
wire n_7034, n_7040, n_7041, n_7042, n_7043, n_7044, n_7046, n_7048;
wire n_7022, n_7024, n_7025, n_7026, n_7027, n_7030, n_7031, n_7033;
wire n_7012, n_7013, n_7014, n_7015, n_7016, n_7017, n_7020, n_7021;
wire n_7003, n_7004, n_7005, n_7007, n_7008, n_7009, n_7010, n_7011;
wire n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999, n_7001;
wire n_6983, n_6984, n_6985, n_6986, n_6987, n_6988, n_6990, n_6992;
wire n_6973, n_6974, n_6975, n_6976, n_6977, n_6979, n_6980, n_6982;
wire n_6962, n_6963, n_6964, n_6965, n_6968, n_6970, n_6971, n_6972;
wire n_6950, n_6951, n_6952, n_6954, n_6956, n_6959, n_6960, n_6961;
wire n_6939, n_6940, n_6942, n_6943, n_6944, n_6945, n_6947, n_6948;
wire n_6928, n_6929, n_6931, n_6932, n_6933, n_6936, n_6937, n_6938;
wire n_6918, n_6919, n_6921, n_6922, n_6923, n_6924, n_6926, n_6927;
wire n_6909, n_6910, n_6911, n_6912, n_6913, n_6914, n_6916, n_6917;
wire n_6899, n_6900, n_6901, n_6902, n_6903, n_6904, n_6906, n_6908;
wire n_6888, n_6891, n_6892, n_6893, n_6894, n_6895, n_6896, n_6897;
wire n_6876, n_6877, n_6878, n_6881, n_6882, n_6883, n_6885, n_6887;
wire n_6865, n_6867, n_6868, n_6869, n_6870, n_6871, n_6874, n_6875;
wire n_6854, n_6855, n_6856, n_6857, n_6858, n_6860, n_6861, n_6863;
wire n_6844, n_6845, n_6847, n_6848, n_6850, n_6851, n_6852, n_6853;
wire n_6834, n_6835, n_6836, n_6837, n_6838, n_6840, n_6841, n_6842;
wire n_6818, n_6822, n_6823, n_6825, n_6829, n_6831, n_6832, n_6833;
wire n_6797, n_6798, n_6800, n_6802, n_6803, n_6806, n_6810, n_6814;
wire n_6779, n_6782, n_6783, n_6785, n_6787, n_6792, n_6793, n_6796;
wire n_6762, n_6763, n_6765, n_6767, n_6769, n_6770, n_6773, n_6774;
wire n_6751, n_6752, n_6753, n_6754, n_6755, n_6756, n_6757, n_6761;
wire n_6740, n_6741, n_6743, n_6744, n_6745, n_6747, n_6748, n_6750;
wire n_6731, n_6732, n_6734, n_6735, n_6736, n_6737, n_6738, n_6739;
wire n_6722, n_6723, n_6724, n_6725, n_6726, n_6727, n_6728, n_6730;
wire n_6708, n_6712, n_6714, n_6715, n_6716, n_6718, n_6720, n_6721;
wire n_6697, n_6698, n_6701, n_6702, n_6703, n_6704, n_6706, n_6707;
wire n_6687, n_6688, n_6689, n_6690, n_6692, n_6693, n_6695, n_6696;
wire n_6675, n_6676, n_6677, n_6680, n_6681, n_6683, n_6684, n_6685;
wire n_6664, n_6665, n_6666, n_6667, n_6668, n_6671, n_6672, n_6674;
wire n_6653, n_6655, n_6656, n_6657, n_6658, n_6659, n_6661, n_6662;
wire n_6644, n_6645, n_6646, n_6647, n_6648, n_6650, n_6651, n_6652;
wire n_6630, n_6631, n_6634, n_6637, n_6638, n_6639, n_6641, n_6643;
wire n_6621, n_6622, n_6623, n_6624, n_6625, n_6626, n_6628, n_6629;
wire n_6612, n_6613, n_6614, n_6615, n_6616, n_6618, n_6619, n_6620;
wire n_6601, n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608;
wire n_6592, n_6593, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600;
wire n_6582, n_6583, n_6584, n_6585, n_6587, n_6588, n_6589, n_6591;
wire n_6571, n_6572, n_6574, n_6575, n_6576, n_6577, n_6579, n_6581;
wire n_6560, n_6562, n_6563, n_6564, n_6565, n_6566, n_6568, n_6570;
wire n_6546, n_6547, n_6548, n_6549, n_6550, n_6551, n_6556, n_6559;
wire n_6534, n_6537, n_6538, n_6539, n_6540, n_6541, n_6544, n_6545;
wire n_6521, n_6522, n_6524, n_6526, n_6527, n_6528, n_6529, n_6532;
wire n_6511, n_6512, n_6514, n_6515, n_6517, n_6518, n_6519, n_6520;
wire n_6499, n_6500, n_6501, n_6502, n_6503, n_6504, n_6506, n_6510;
wire n_6482, n_6483, n_6484, n_6488, n_6491, n_6493, n_6495, n_6496;
wire n_6468, n_6469, n_6471, n_6473, n_6477, n_6478, n_6480, n_6481;
wire n_6454, n_6455, n_6459, n_6460, n_6463, n_6464, n_6466, n_6467;
wire n_6441, n_6443, n_6445, n_6446, n_6447, n_6448, n_6452, n_6453;
wire n_6421, n_6425, n_6429, n_6435, n_6436, n_6437, n_6438, n_6439;
wire n_6405, n_6406, n_6407, n_6408, n_6409, n_6414, n_6416, n_6419;
wire n_6396, n_6398, n_6399, n_6400, n_6401, n_6402, n_6403, n_6404;
wire n_6383, n_6385, n_6387, n_6389, n_6392, n_6393, n_6394, n_6395;
wire n_6372, n_6374, n_6375, n_6376, n_6377, n_6378, n_6379, n_6382;
wire n_6356, n_6357, n_6359, n_6360, n_6362, n_6365, n_6368, n_6371;
wire n_6347, n_6348, n_6349, n_6351, n_6352, n_6353, n_6354, n_6355;
wire n_6338, n_6339, n_6341, n_6342, n_6343, n_6344, n_6345, n_6346;
wire n_6330, n_6331, n_6332, n_6333, n_6334, n_6335, n_6336, n_6337;
wire n_6321, n_6322, n_6323, n_6324, n_6326, n_6327, n_6328, n_6329;
wire n_6306, n_6309, n_6310, n_6311, n_6313, n_6315, n_6316, n_6320;
wire n_6296, n_6297, n_6298, n_6299, n_6301, n_6302, n_6303, n_6304;
wire n_6284, n_6285, n_6286, n_6289, n_6290, n_6291, n_6292, n_6293;
wire n_6276, n_6277, n_6278, n_6279, n_6280, n_6281, n_6282, n_6283;
wire n_6268, n_6269, n_6270, n_6271, n_6272, n_6273, n_6274, n_6275;
wire n_6253, n_6255, n_6256, n_6258, n_6259, n_6262, n_6265, n_6266;
wire n_6244, n_6246, n_6247, n_6248, n_6249, n_6250, n_6251, n_6252;
wire n_6236, n_6237, n_6238, n_6239, n_6240, n_6241, n_6242, n_6243;
wire n_6224, n_6227, n_6230, n_6231, n_6232, n_6233, n_6234, n_6235;
wire n_6212, n_6213, n_6214, n_6215, n_6218, n_6220, n_6221, n_6222;
wire n_6204, n_6205, n_6206, n_6207, n_6208, n_6209, n_6210, n_6211;
wire n_6196, n_6197, n_6198, n_6199, n_6200, n_6201, n_6202, n_6203;
wire n_6188, n_6189, n_6190, n_6191, n_6192, n_6193, n_6194, n_6195;
wire n_6177, n_6178, n_6179, n_6180, n_6182, n_6183, n_6185, n_6186;
wire n_6167, n_6168, n_6169, n_6170, n_6172, n_6173, n_6174, n_6175;
wire n_6155, n_6156, n_6157, n_6158, n_6160, n_6164, n_6165, n_6166;
wire n_6146, n_6147, n_6148, n_6149, n_6150, n_6151, n_6153, n_6154;
wire n_6138, n_6139, n_6140, n_6141, n_6142, n_6143, n_6144, n_6145;
wire n_6130, n_6131, n_6132, n_6133, n_6134, n_6135, n_6136, n_6137;
wire n_6121, n_6122, n_6123, n_6124, n_6125, n_6126, n_6127, n_6128;
wire n_6113, n_6114, n_6115, n_6116, n_6117, n_6118, n_6119, n_6120;
wire n_6103, n_6105, n_6106, n_6107, n_6109, n_6110, n_6111, n_6112;
wire n_6095, n_6096, n_6097, n_6098, n_6099, n_6100, n_6101, n_6102;
wire n_6087, n_6088, n_6089, n_6090, n_6091, n_6092, n_6093, n_6094;
wire n_6077, n_6078, n_6079, n_6080, n_6081, n_6083, n_6085, n_6086;
wire n_6069, n_6070, n_6071, n_6072, n_6073, n_6074, n_6075, n_6076;
wire n_6061, n_6062, n_6063, n_6064, n_6065, n_6066, n_6067, n_6068;
wire n_6053, n_6054, n_6055, n_6056, n_6057, n_6058, n_6059, n_6060;
wire n_6045, n_6046, n_6047, n_6048, n_6049, n_6050, n_6051, n_6052;
wire n_6036, n_6037, n_6038, n_6039, n_6040, n_6042, n_6043, n_6044;
wire n_6028, n_6029, n_6030, n_6031, n_6032, n_6033, n_6034, n_6035;
wire n_6020, n_6021, n_6022, n_6023, n_6024, n_6025, n_6026, n_6027;
wire n_6010, n_6011, n_6012, n_6015, n_6016, n_6017, n_6018, n_6019;
wire n_6002, n_6003, n_6004, n_6005, n_6006, n_6007, n_6008, n_6009;
wire n_5994, n_5995, n_5996, n_5997, n_5998, n_5999, n_6000, n_6001;
wire n_5982, n_5986, n_5988, n_5989, n_5990, n_5991, n_5992, n_5993;
wire n_5974, n_5975, n_5976, n_5977, n_5978, n_5979, n_5980, n_5981;
wire n_5964, n_5965, n_5967, n_5969, n_5970, n_5971, n_5972, n_5973;
wire n_5956, n_5957, n_5958, n_5959, n_5960, n_5961, n_5962, n_5963;
wire n_5948, n_5949, n_5950, n_5951, n_5952, n_5953, n_5954, n_5955;
wire n_5940, n_5941, n_5942, n_5943, n_5944, n_5945, n_5946, n_5947;
wire n_5932, n_5933, n_5934, n_5935, n_5936, n_5937, n_5938, n_5939;
wire n_5924, n_5925, n_5926, n_5927, n_5928, n_5929, n_5930, n_5931;
wire n_5916, n_5917, n_5918, n_5919, n_5920, n_5921, n_5922, n_5923;
wire n_5908, n_5909, n_5910, n_5911, n_5912, n_5913, n_5914, n_5915;
wire n_5898, n_5901, n_5902, n_5903, n_5904, n_5905, n_5906, n_5907;
wire n_5890, n_5891, n_5892, n_5893, n_5894, n_5895, n_5896, n_5897;
wire n_5880, n_5881, n_5882, n_5883, n_5886, n_5887, n_5888, n_5889;
wire n_5871, n_5872, n_5873, n_5874, n_5875, n_5877, n_5878, n_5879;
wire n_5863, n_5864, n_5865, n_5866, n_5867, n_5868, n_5869, n_5870;
wire n_5855, n_5856, n_5857, n_5858, n_5859, n_5860, n_5861, n_5862;
wire n_5847, n_5848, n_5849, n_5850, n_5851, n_5852, n_5853, n_5854;
wire n_5837, n_5839, n_5840, n_5841, n_5842, n_5843, n_5844, n_5845;
wire n_5828, n_5829, n_5830, n_5831, n_5832, n_5833, n_5834, n_5836;
wire n_5820, n_5821, n_5822, n_5823, n_5824, n_5825, n_5826, n_5827;
wire n_5812, n_5813, n_5814, n_5815, n_5816, n_5817, n_5818, n_5819;
wire n_5803, n_5804, n_5805, n_5806, n_5807, n_5808, n_5809, n_5811;
wire n_5795, n_5796, n_5797, n_5798, n_5799, n_5800, n_5801, n_5802;
wire n_5786, n_5787, n_5789, n_5790, n_5791, n_5792, n_5793, n_5794;
wire n_5778, n_5779, n_5780, n_5781, n_5782, n_5783, n_5784, n_5785;
wire n_5770, n_5771, n_5772, n_5773, n_5774, n_5775, n_5776, n_5777;
wire n_5762, n_5763, n_5764, n_5765, n_5766, n_5767, n_5768, n_5769;
wire n_5754, n_5755, n_5756, n_5757, n_5758, n_5759, n_5760, n_5761;
wire n_5746, n_5747, n_5748, n_5749, n_5750, n_5751, n_5752, n_5753;
wire n_5738, n_5739, n_5740, n_5741, n_5742, n_5743, n_5744, n_5745;
wire n_5729, n_5730, n_5731, n_5732, n_5734, n_5735, n_5736, n_5737;
wire n_5720, n_5721, n_5722, n_5723, n_5724, n_5725, n_5726, n_5727;
wire n_5712, n_5713, n_5714, n_5715, n_5716, n_5717, n_5718, n_5719;
wire n_5704, n_5705, n_5706, n_5707, n_5708, n_5709, n_5710, n_5711;
wire n_5696, n_5697, n_5698, n_5699, n_5700, n_5701, n_5702, n_5703;
wire n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5695;
wire n_5678, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686;
wire n_5670, n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677;
wire n_5662, n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669;
wire n_5654, n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661;
wire n_5646, n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653;
wire n_5638, n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645;
wire n_5630, n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637;
wire n_5621, n_5623, n_5624, n_5625, n_5626, n_5627, n_5628, n_5629;
wire n_5613, n_5614, n_5615, n_5616, n_5617, n_5618, n_5619, n_5620;
wire n_5605, n_5606, n_5607, n_5608, n_5609, n_5610, n_5611, n_5612;
wire n_5597, n_5598, n_5599, n_5600, n_5601, n_5602, n_5603, n_5604;
wire n_5588, n_5589, n_5590, n_5591, n_5592, n_5593, n_5595, n_5596;
wire n_5579, n_5580, n_5581, n_5582, n_5583, n_5585, n_5586, n_5587;
wire n_5569, n_5570, n_5571, n_5573, n_5575, n_5576, n_5577, n_5578;
wire n_5561, n_5562, n_5563, n_5564, n_5565, n_5566, n_5567, n_5568;
wire n_5553, n_5554, n_5555, n_5556, n_5557, n_5558, n_5559, n_5560;
wire n_5545, n_5546, n_5547, n_5548, n_5549, n_5550, n_5551, n_5552;
wire n_5537, n_5538, n_5539, n_5540, n_5541, n_5542, n_5543, n_5544;
wire n_5529, n_5530, n_5531, n_5532, n_5533, n_5534, n_5535, n_5536;
wire n_5518, n_5519, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526;
wire n_5510, n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517;
wire n_5502, n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509;
wire n_5494, n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501;
wire n_5485, n_5486, n_5487, n_5488, n_5489, n_5491, n_5492, n_5493;
wire n_5474, n_5475, n_5478, n_5479, n_5480, n_5481, n_5483, n_5484;
wire n_5465, n_5466, n_5467, n_5468, n_5469, n_5470, n_5471, n_5472;
wire n_5457, n_5458, n_5459, n_5460, n_5461, n_5462, n_5463, n_5464;
wire n_5448, n_5450, n_5451, n_5452, n_5453, n_5454, n_5455, n_5456;
wire n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446, n_5447;
wire n_5431, n_5432, n_5433, n_5435, n_5436, n_5437, n_5438, n_5439;
wire n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429, n_5430;
wire n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421, n_5422;
wire n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413, n_5414;
wire n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405, n_5406;
wire n_5391, n_5392, n_5393, n_5394, n_5395, n_5396, n_5397, n_5398;
wire n_5383, n_5384, n_5385, n_5386, n_5387, n_5388, n_5389, n_5390;
wire n_5375, n_5376, n_5377, n_5378, n_5379, n_5380, n_5381, n_5382;
wire n_5367, n_5368, n_5369, n_5370, n_5371, n_5372, n_5373, n_5374;
wire n_5355, n_5356, n_5357, n_5358, n_5359, n_5361, n_5364, n_5366;
wire n_5347, n_5348, n_5349, n_5350, n_5351, n_5352, n_5353, n_5354;
wire n_5338, n_5340, n_5341, n_5342, n_5343, n_5344, n_5345, n_5346;
wire n_5330, n_5331, n_5332, n_5333, n_5334, n_5335, n_5336, n_5337;
wire n_5320, n_5321, n_5322, n_5325, n_5326, n_5327, n_5328, n_5329;
wire n_5308, n_5310, n_5312, n_5315, n_5316, n_5317, n_5318, n_5319;
wire n_5300, n_5301, n_5302, n_5303, n_5304, n_5305, n_5306, n_5307;
wire n_5292, n_5293, n_5294, n_5295, n_5296, n_5297, n_5298, n_5299;
wire n_5284, n_5285, n_5286, n_5287, n_5288, n_5289, n_5290, n_5291;
wire n_5276, n_5277, n_5278, n_5279, n_5280, n_5281, n_5282, n_5283;
wire n_5266, n_5269, n_5270, n_5271, n_5272, n_5273, n_5274, n_5275;
wire n_5255, n_5257, n_5258, n_5259, n_5260, n_5261, n_5262, n_5263;
wire n_5247, n_5248, n_5249, n_5250, n_5251, n_5252, n_5253, n_5254;
wire n_5238, n_5239, n_5240, n_5241, n_5242, n_5244, n_5245, n_5246;
wire n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236, n_5237;
wire n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228, n_5229;
wire n_5213, n_5214, n_5215, n_5216, n_5218, n_5219, n_5220, n_5221;
wire n_5203, n_5204, n_5205, n_5206, n_5207, n_5208, n_5210, n_5211;
wire n_5194, n_5195, n_5196, n_5197, n_5198, n_5199, n_5200, n_5202;
wire n_5186, n_5187, n_5188, n_5189, n_5190, n_5191, n_5192, n_5193;
wire n_5177, n_5178, n_5179, n_5180, n_5181, n_5182, n_5183, n_5185;
wire n_5169, n_5170, n_5171, n_5172, n_5173, n_5174, n_5175, n_5176;
wire n_5158, n_5159, n_5160, n_5161, n_5163, n_5164, n_5167, n_5168;
wire n_5148, n_5149, n_5150, n_5151, n_5152, n_5155, n_5156, n_5157;
wire n_5140, n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147;
wire n_5132, n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139;
wire n_5123, n_5124, n_5125, n_5126, n_5127, n_5129, n_5130, n_5131;
wire n_5115, n_5116, n_5117, n_5118, n_5119, n_5120, n_5121, n_5122;
wire n_5107, n_5108, n_5109, n_5110, n_5111, n_5112, n_5113, n_5114;
wire n_5096, n_5098, n_5099, n_5100, n_5101, n_5104, n_5105, n_5106;
wire n_5088, n_5089, n_5090, n_5091, n_5092, n_5093, n_5094, n_5095;
wire n_5080, n_5081, n_5082, n_5083, n_5084, n_5085, n_5086, n_5087;
wire n_5072, n_5073, n_5074, n_5075, n_5076, n_5077, n_5078, n_5079;
wire n_5061, n_5062, n_5063, n_5064, n_5065, n_5067, n_5070, n_5071;
wire n_5051, n_5052, n_5053, n_5054, n_5055, n_5056, n_5059, n_5060;
wire n_5043, n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050;
wire n_5033, n_5034, n_5035, n_5037, n_5038, n_5039, n_5041, n_5042;
wire n_5023, n_5024, n_5027, n_5028, n_5029, n_5030, n_5031, n_5032;
wire n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5021, n_5022;
wire n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011;
wire n_4993, n_4994, n_4997, n_4998, n_5000, n_5001, n_5002, n_5003;
wire n_4985, n_4986, n_4987, n_4988, n_4989, n_4990, n_4991, n_4992;
wire n_4976, n_4977, n_4978, n_4980, n_4981, n_4982, n_4983, n_4984;
wire n_4968, n_4969, n_4970, n_4971, n_4972, n_4973, n_4974, n_4975;
wire n_4959, n_4960, n_4961, n_4962, n_4963, n_4965, n_4966, n_4967;
wire n_4947, n_4948, n_4949, n_4953, n_4954, n_4955, n_4956, n_4957;
wire n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946;
wire n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938;
wire n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930;
wire n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922;
wire n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914;
wire n_4899, n_4900, n_4901, n_4902, n_4903, n_4904, n_4905, n_4906;
wire n_4888, n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895;
wire n_4880, n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887;
wire n_4867, n_4868, n_4870, n_4871, n_4872, n_4873, n_4874, n_4877;
wire n_4859, n_4860, n_4861, n_4862, n_4863, n_4864, n_4865, n_4866;
wire n_4848, n_4851, n_4852, n_4853, n_4854, n_4855, n_4856, n_4857;
wire n_4839, n_4840, n_4841, n_4842, n_4844, n_4845, n_4846, n_4847;
wire n_4828, n_4829, n_4830, n_4832, n_4833, n_4834, n_4835, n_4836;
wire n_4818, n_4820, n_4821, n_4822, n_4823, n_4824, n_4825, n_4826;
wire n_4808, n_4810, n_4811, n_4812, n_4813, n_4814, n_4815, n_4817;
wire n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806, n_4807;
wire n_4791, n_4792, n_4793, n_4794, n_4796, n_4797, n_4798, n_4799;
wire n_4782, n_4783, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790;
wire n_4772, n_4774, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781;
wire n_4762, n_4764, n_4766, n_4767, n_4768, n_4769, n_4770, n_4771;
wire n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4759;
wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
wire n_4734, n_4735, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742;
wire n_4725, n_4726, n_4727, n_4728, n_4730, n_4731, n_4732, n_4733;
wire n_4714, n_4718, n_4719, n_4720, n_4721, n_4722, n_4723, n_4724;
wire n_4703, n_4706, n_4707, n_4708, n_4710, n_4711, n_4712, n_4713;
wire n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701;
wire n_4682, n_4684, n_4685, n_4688, n_4689, n_4690, n_4692, n_4693;
wire n_4668, n_4669, n_4670, n_4671, n_4674, n_4675, n_4677, n_4681;
wire n_4654, n_4655, n_4656, n_4657, n_4658, n_4663, n_4665, n_4666;
wire n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653;
wire n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645;
wire n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637;
wire n_4619, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629;
wire n_4611, n_4612, n_4613, n_4614, n_4615, n_4616, n_4617, n_4618;
wire n_4601, n_4602, n_4605, n_4606, n_4607, n_4608, n_4609, n_4610;
wire n_4593, n_4594, n_4595, n_4596, n_4597, n_4598, n_4599, n_4600;
wire n_4584, n_4585, n_4586, n_4588, n_4589, n_4590, n_4591, n_4592;
wire n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581, n_4582;
wire n_4566, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573, n_4574;
wire n_4556, n_4557, n_4559, n_4560, n_4561, n_4562, n_4563, n_4565;
wire n_4548, n_4549, n_4550, n_4551, n_4552, n_4553, n_4554, n_4555;
wire n_4538, n_4540, n_4541, n_4542, n_4544, n_4545, n_4546, n_4547;
wire n_4530, n_4531, n_4532, n_4533, n_4534, n_4535, n_4536, n_4537;
wire n_4519, n_4520, n_4521, n_4523, n_4524, n_4525, n_4526, n_4528;
wire n_4508, n_4509, n_4511, n_4512, n_4514, n_4515, n_4516, n_4518;
wire n_4497, n_4498, n_4499, n_4502, n_4503, n_4504, n_4505, n_4507;
wire n_4486, n_4487, n_4488, n_4491, n_4493, n_4494, n_4495, n_4496;
wire n_4472, n_4473, n_4474, n_4475, n_4476, n_4477, n_4478, n_4481;
wire n_4464, n_4465, n_4466, n_4467, n_4468, n_4469, n_4470, n_4471;
wire n_4455, n_4456, n_4457, n_4459, n_4460, n_4461, n_4462, n_4463;
wire n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453, n_4454;
wire n_4437, n_4439, n_4441, n_4442, n_4443, n_4444, n_4445, n_4446;
wire n_4426, n_4428, n_4429, n_4430, n_4431, n_4432, n_4433, n_4436;
wire n_4418, n_4419, n_4420, n_4421, n_4422, n_4423, n_4424, n_4425;
wire n_4409, n_4410, n_4411, n_4412, n_4414, n_4415, n_4416, n_4417;
wire n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4408;
wire n_4388, n_4389, n_4391, n_4392, n_4394, n_4395, n_4396, n_4398;
wire n_4378, n_4379, n_4380, n_4381, n_4382, n_4384, n_4385, n_4386;
wire n_4367, n_4368, n_4371, n_4372, n_4373, n_4375, n_4376, n_4377;
wire n_4357, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365;
wire n_4347, n_4349, n_4350, n_4351, n_4353, n_4354, n_4355, n_4356;
wire n_4339, n_4340, n_4341, n_4342, n_4343, n_4344, n_4345, n_4346;
wire n_4323, n_4324, n_4325, n_4326, n_4328, n_4334, n_4335, n_4336;
wire n_4311, n_4313, n_4315, n_4318, n_4319, n_4320, n_4321, n_4322;
wire n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4310;
wire n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301;
wire n_4285, n_4286, n_4287, n_4288, n_4289, n_4290, n_4291, n_4293;
wire n_4277, n_4278, n_4279, n_4280, n_4281, n_4282, n_4283, n_4284;
wire n_4263, n_4264, n_4265, n_4266, n_4267, n_4270, n_4271, n_4274;
wire n_4255, n_4256, n_4257, n_4258, n_4259, n_4260, n_4261, n_4262;
wire n_4247, n_4248, n_4249, n_4250, n_4251, n_4252, n_4253, n_4254;
wire n_4236, n_4237, n_4240, n_4241, n_4242, n_4243, n_4244, n_4246;
wire n_4226, n_4229, n_4230, n_4231, n_4232, n_4233, n_4234, n_4235;
wire n_4215, n_4217, n_4218, n_4219, n_4220, n_4223, n_4224, n_4225;
wire n_4202, n_4205, n_4206, n_4209, n_4210, n_4211, n_4212, n_4213;
wire n_4193, n_4194, n_4195, n_4196, n_4197, n_4198, n_4200, n_4201;
wire n_4185, n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192;
wire n_4175, n_4176, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184;
wire n_4162, n_4164, n_4165, n_4166, n_4167, n_4169, n_4170, n_4174;
wire n_4152, n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160;
wire n_4143, n_4145, n_4146, n_4147, n_4148, n_4149, n_4150, n_4151;
wire n_4134, n_4135, n_4136, n_4137, n_4138, n_4139, n_4141, n_4142;
wire n_4124, n_4125, n_4127, n_4129, n_4130, n_4131, n_4132, n_4133;
wire n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121, n_4122;
wire n_4101, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113, n_4114;
wire n_4091, n_4092, n_4094, n_4095, n_4096, n_4097, n_4099, n_4100;
wire n_4079, n_4080, n_4081, n_4082, n_4083, n_4085, n_4086, n_4087;
wire n_4068, n_4069, n_4070, n_4072, n_4073, n_4075, n_4077, n_4078;
wire n_4056, n_4058, n_4059, n_4060, n_4061, n_4065, n_4066, n_4067;
wire n_4046, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055;
wire n_4037, n_4038, n_4039, n_4040, n_4041, n_4042, n_4043, n_4045;
wire n_4029, n_4030, n_4031, n_4032, n_4033, n_4034, n_4035, n_4036;
wire n_4021, n_4022, n_4023, n_4024, n_4025, n_4026, n_4027, n_4028;
wire n_4011, n_4012, n_4013, n_4014, n_4015, n_4017, n_4019, n_4020;
wire n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4009, n_4010;
wire n_3991, n_3992, n_3993, n_3994, n_3995, n_3996, n_3997, n_3999;
wire n_3982, n_3983, n_3984, n_3985, n_3986, n_3987, n_3989, n_3990;
wire n_3973, n_3974, n_3976, n_3977, n_3978, n_3979, n_3980, n_3981;
wire n_3962, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969, n_3971;
wire n_3953, n_3954, n_3955, n_3957, n_3958, n_3959, n_3960, n_3961;
wire n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952;
wire n_3937, n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944;
wire n_3926, n_3927, n_3928, n_3930, n_3932, n_3933, n_3935, n_3936;
wire n_3916, n_3917, n_3919, n_3920, n_3921, n_3922, n_3923, n_3925;
wire n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, n_3915;
wire n_3897, n_3899, n_3902, n_3903, n_3904, n_3905, n_3906, n_3907;
wire n_3888, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896;
wire n_3879, n_3880, n_3881, n_3883, n_3884, n_3885, n_3886, n_3887;
wire n_3868, n_3869, n_3870, n_3871, n_3873, n_3876, n_3877, n_3878;
wire n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, n_3866;
wire n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856;
wire n_3836, n_3837, n_3838, n_3841, n_3842, n_3845, n_3847, n_3848;
wire n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, n_3834, n_3835;
wire n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825, n_3826;
wire n_3809, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817;
wire n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, n_3808;
wire n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, n_3798, n_3799;
wire n_3784, n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791;
wire n_3775, n_3776, n_3777, n_3778, n_3779, n_3781, n_3782, n_3783;
wire n_3765, n_3766, n_3767, n_3768, n_3770, n_3771, n_3772, n_3774;
wire n_3753, n_3754, n_3758, n_3759, n_3760, n_3761, n_3762, n_3764;
wire n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752;
wire n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744;
wire n_3724, n_3725, n_3726, n_3727, n_3728, n_3730, n_3731, n_3736;
wire n_3709, n_3713, n_3714, n_3715, n_3716, n_3719, n_3720, n_3723;
wire n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3707, n_3708;
wire n_3689, n_3690, n_3691, n_3693, n_3694, n_3695, n_3697, n_3698;
wire n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688;
wire n_3672, n_3673, n_3674, n_3675, n_3676, n_3678, n_3679, n_3680;
wire n_3663, n_3664, n_3665, n_3666, n_3668, n_3669, n_3670, n_3671;
wire n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661;
wire n_3645, n_3646, n_3647, n_3648, n_3650, n_3651, n_3652, n_3653;
wire n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644;
wire n_3627, n_3628, n_3629, n_3630, n_3631, n_3634, n_3635, n_3636;
wire n_3611, n_3612, n_3613, n_3614, n_3615, n_3617, n_3618, n_3621;
wire n_3599, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3609;
wire n_3586, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3596;
wire n_3573, n_3576, n_3577, n_3578, n_3580, n_3582, n_3583, n_3585;
wire n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3570;
wire n_3551, n_3552, n_3553, n_3556, n_3558, n_3559, n_3560, n_3561;
wire n_3541, n_3542, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550;
wire n_3531, n_3532, n_3533, n_3534, n_3536, n_3537, n_3538, n_3540;
wire n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530;
wire n_3514, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522;
wire n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513;
wire n_3496, n_3497, n_3498, n_3500, n_3501, n_3502, n_3504, n_3505;
wire n_3486, n_3487, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495;
wire n_3474, n_3476, n_3477, n_3478, n_3479, n_3481, n_3483, n_3485;
wire n_3464, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472;
wire n_3453, n_3454, n_3455, n_3456, n_3457, n_3460, n_3462, n_3463;
wire n_3443, n_3444, n_3445, n_3447, n_3449, n_3450, n_3451, n_3452;
wire n_3432, n_3433, n_3434, n_3436, n_3438, n_3440, n_3441, n_3442;
wire n_3421, n_3422, n_3423, n_3425, n_3426, n_3427, n_3429, n_3431;
wire n_3410, n_3411, n_3412, n_3413, n_3416, n_3418, n_3419, n_3420;
wire n_3399, n_3402, n_3403, n_3404, n_3405, n_3406, n_3408, n_3409;
wire n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3397;
wire n_3379, n_3380, n_3381, n_3382, n_3385, n_3386, n_3387, n_3388;
wire n_3367, n_3368, n_3370, n_3372, n_3373, n_3374, n_3375, n_3377;
wire n_3357, n_3359, n_3360, n_3361, n_3362, n_3364, n_3365, n_3366;
wire n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356;
wire n_3340, n_3341, n_3342, n_3343, n_3345, n_3346, n_3347, n_3348;
wire n_3329, n_3331, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338;
wire n_3320, n_3321, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328;
wire n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, n_3318;
wire n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309;
wire n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301;
wire n_3282, n_3283, n_3284, n_3285, n_3288, n_3289, n_3292, n_3293;
wire n_3273, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281;
wire n_3263, n_3264, n_3266, n_3268, n_3269, n_3270, n_3271, n_3272;
wire n_3253, n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3262;
wire n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252;
wire n_3234, n_3235, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244;
wire n_3225, n_3226, n_3227, n_3228, n_3230, n_3231, n_3232, n_3233;
wire n_3215, n_3217, n_3218, n_3220, n_3221, n_3222, n_3223, n_3224;
wire n_3203, n_3204, n_3205, n_3206, n_3207, n_3209, n_3210, n_3212;
wire n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202;
wire n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194;
wire n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, n_3186;
wire n_3169, n_3170, n_3171, n_3173, n_3174, n_3176, n_3177, n_3178;
wire n_3159, n_3160, n_3161, n_3162, n_3165, n_3166, n_3167, n_3168;
wire n_3148, n_3150, n_3151, n_3152, n_3153, n_3156, n_3157, n_3158;
wire n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147;
wire n_3126, n_3127, n_3129, n_3133, n_3136, n_3137, n_3138, n_3139;
wire n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3124, n_3125;
wire n_3106, n_3107, n_3108, n_3109, n_3110, n_3112, n_3114, n_3115;
wire n_3097, n_3098, n_3099, n_3100, n_3101, n_3103, n_3104, n_3105;
wire n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, n_3096;
wire n_3079, n_3081, n_3082, n_3084, n_3085, n_3086, n_3087, n_3088;
wire n_3068, n_3069, n_3070, n_3071, n_3072, n_3074, n_3075, n_3078;
wire n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3067;
wire n_3049, n_3050, n_3052, n_3054, n_3055, n_3056, n_3057, n_3058;
wire n_3039, n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048;
wire n_3027, n_3029, n_3032, n_3034, n_3035, n_3036, n_3037, n_3038;
wire n_3018, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026;
wire n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3017;
wire n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005;
wire n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, n_2997;
wire n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, n_2988, n_2989;
wire n_2971, n_2972, n_2974, n_2975, n_2976, n_2977, n_2979, n_2980;
wire n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2969;
wire n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960;
wire n_2944, n_2945, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952;
wire n_2934, n_2936, n_2937, n_2938, n_2939, n_2941, n_2942, n_2943;
wire n_2921, n_2926, n_2927, n_2928, n_2929, n_2931, n_2932, n_2933;
wire n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2920;
wire n_2903, n_2904, n_2905, n_2907, n_2908, n_2909, n_2910, n_2911;
wire n_2892, n_2893, n_2894, n_2895, n_2896, n_2898, n_2899, n_2900;
wire n_2883, n_2884, n_2885, n_2886, n_2887, n_2889, n_2890, n_2891;
wire n_2875, n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882;
wire n_2864, n_2865, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874;
wire n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863;
wire n_2848, n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855;
wire n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847;
wire n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839;
wire n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831;
wire n_2815, n_2816, n_2817, n_2819, n_2820, n_2821, n_2822, n_2823;
wire n_2806, n_2807, n_2808, n_2810, n_2811, n_2812, n_2813, n_2814;
wire n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805;
wire n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797;
wire n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789;
wire n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, n_2781;
wire n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, n_2772, n_2773;
wire n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, n_2763, n_2764;
wire n_2747, n_2748, n_2749, n_2751, n_2752, n_2753, n_2754, n_2755;
wire n_2737, n_2738, n_2739, n_2740, n_2742, n_2743, n_2745, n_2746;
wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
wire n_2712, n_2713, n_2714, n_2715, n_2716, n_2718, n_2719, n_2720;
wire n_2701, n_2704, n_2705, n_2706, n_2707, n_2708, n_2710, n_2711;
wire n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2698, n_2699;
wire n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689;
wire n_2673, n_2674, n_2675, n_2676, n_2678, n_2679, n_2680, n_2681;
wire n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
wire n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664;
wire n_2645, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654;
wire n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644;
wire n_2628, n_2629, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636;
wire n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627;
wire n_2608, n_2609, n_2610, n_2611, n_2612, n_2615, n_2616, n_2618;
wire n_2599, n_2600, n_2601, n_2602, n_2603, n_2605, n_2606, n_2607;
wire n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598;
wire n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590;
wire n_2574, n_2575, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582;
wire n_2565, n_2566, n_2567, n_2569, n_2570, n_2571, n_2572, n_2573;
wire n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564;
wire n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2556;
wire n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, n_2547;
wire n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, n_2538, n_2539;
wire n_2524, n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531;
wire n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, n_2520, n_2523;
wire n_2505, n_2506, n_2507, n_2508, n_2509, n_2511, n_2512, n_2513;
wire n_2497, n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504;
wire n_2488, n_2489, n_2490, n_2491, n_2493, n_2494, n_2495, n_2496;
wire n_2479, n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486;
wire n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478;
wire n_2461, n_2462, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469;
wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
wire n_2443, n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450;
wire n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442;
wire n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434;
wire n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426;
wire n_2409, n_2410, n_2412, n_2413, n_2414, n_2415, n_2417, n_2418;
wire n_2400, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408;
wire n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2399;
wire n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390;
wire n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382;
wire n_2366, n_2367, n_2368, n_2369, n_2370, n_2372, n_2373, n_2374;
wire n_2356, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365;
wire n_2346, n_2347, n_2348, n_2349, n_2351, n_2352, n_2353, n_2355;
wire n_2336, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344;
wire n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334;
wire n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325;
wire n_2306, n_2307, n_2309, n_2310, n_2311, n_2312, n_2313, n_2317;
wire n_2296, n_2297, n_2298, n_2300, n_2301, n_2302, n_2303, n_2305;
wire n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, n_2295;
wire n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2286, n_2287;
wire n_2268, n_2269, n_2270, n_2271, n_2275, n_2276, n_2277, n_2278;
wire n_2259, n_2260, n_2261, n_2263, n_2264, n_2265, n_2266, n_2267;
wire n_2250, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258;
wire n_2241, n_2242, n_2243, n_2244, n_2245, n_2247, n_2248, n_2249;
wire n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240;
wire n_2224, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, n_2232;
wire n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, n_2223;
wire n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215;
wire n_2199, n_2200, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207;
wire n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198;
wire n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190;
wire n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182;
wire n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174;
wire n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165;
wire n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2155, n_2156;
wire n_2135, n_2136, n_2137, n_2138, n_2140, n_2141, n_2145, n_2146;
wire n_2126, n_2127, n_2129, n_2130, n_2131, n_2132, n_2133, n_2134;
wire n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, n_2124, n_2125;
wire n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117;
wire n_2098, n_2099, n_2100, n_2101, n_2105, n_2106, n_2107, n_2109;
wire n_2087, n_2089, n_2090, n_2091, n_2094, n_2095, n_2096, n_2097;
wire n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086;
wire n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078;
wire n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, n_2070;
wire n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062;
wire n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054;
wire n_2037, n_2038, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046;
wire n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036;
wire n_2015, n_2016, n_2017, n_2020, n_2021, n_2024, n_2026, n_2028;
wire n_2003, n_2004, n_2005, n_2009, n_2010, n_2011, n_2012, n_2013;
wire n_1993, n_1994, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001;
wire n_1980, n_1985, n_1986, n_1987, n_1989, n_1990, n_1991, n_1992;
wire n_1971, n_1972, n_1973, n_1974, n_1976, n_1977, n_1978, n_1979;
wire n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970;
wire n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962;
wire n_1943, n_1944, n_1945, n_1947, n_1949, n_1950, n_1951, n_1952;
wire n_1934, n_1935, n_1936, n_1937, n_1939, n_1940, n_1941, n_1942;
wire n_1925, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933;
wire n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924;
wire n_1908, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916;
wire n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1906, n_1907;
wire n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1897, n_1898;
wire n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887;
wire n_1871, n_1872, n_1873, n_1874, n_1875, n_1877, n_1878, n_1879;
wire n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870;
wire n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1860, n_1861;
wire n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852;
wire n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1844;
wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1834;
wire n_1813, n_1814, n_1817, n_1818, n_1821, n_1822, n_1823, n_1824;
wire n_1804, n_1805, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812;
wire n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803;
wire n_1787, n_1788, n_1789, n_1790, n_1791, n_1793, n_1794, n_1795;
wire n_1778, n_1779, n_1780, n_1782, n_1783, n_1784, n_1785, n_1786;
wire n_1768, n_1769, n_1770, n_1771, n_1772, n_1774, n_1775, n_1777;
wire n_1759, n_1760, n_1761, n_1762, n_1763, n_1765, n_1766, n_1767;
wire n_1748, n_1749, n_1750, n_1753, n_1754, n_1756, n_1757, n_1758;
wire n_1737, n_1738, n_1739, n_1740, n_1742, n_1745, n_1746, n_1747;
wire n_1725, n_1727, n_1728, n_1729, n_1731, n_1732, n_1733, n_1735;
wire n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724;
wire n_1705, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1715;
wire n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704;
wire n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696;
wire n_1680, n_1681, n_1682, n_1683, n_1684, n_1686, n_1687, n_1688;
wire n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1675, n_1677;
wire n_1658, n_1659, n_1661, n_1662, n_1663, n_1664, n_1666, n_1667;
wire n_1647, n_1648, n_1651, n_1652, n_1653, n_1654, n_1655, n_1657;
wire n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646;
wire n_1625, n_1626, n_1627, n_1629, n_1630, n_1632, n_1633, n_1634;
wire n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624;
wire n_1608, n_1609, n_1610, n_1611, n_1612, n_1614, n_1615, n_1616;
wire n_1592, n_1593, n_1595, n_1602, n_1603, n_1604, n_1605, n_1607;
wire n_1582, n_1583, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591;
wire n_1573, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581;
wire n_1563, n_1564, n_1565, n_1566, n_1568, n_1569, n_1570, n_1572;
wire n_1554, n_1555, n_1556, n_1558, n_1559, n_1560, n_1561, n_1562;
wire n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553;
wire n_1535, n_1536, n_1537, n_1541, n_1542, n_1543, n_1544, n_1545;
wire n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
wire n_1517, n_1518, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526;
wire n_1503, n_1504, n_1508, n_1509, n_1510, n_1511, n_1512, n_1516;
wire n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502;
wire n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1494;
wire n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1484, n_1485;
wire n_1467, n_1468, n_1469, n_1470, n_1471, n_1473, n_1474, n_1475;
wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1464, n_1465, n_1466;
wire n_1449, n_1450, n_1451, n_1453, n_1454, n_1455, n_1456, n_1457;
wire n_1438, n_1439, n_1440, n_1444, n_1445, n_1446, n_1447, n_1448;
wire n_1429, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437;
wire n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428;
wire n_1412, n_1413, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420;
wire n_1400, n_1401, n_1402, n_1403, n_1405, n_1407, n_1409, n_1411;
wire n_1388, n_1391, n_1393, n_1394, n_1396, n_1397, n_1398, n_1399;
wire n_1379, n_1380, n_1381, n_1382, n_1383, n_1385, n_1386, n_1387;
wire n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1377, n_1378;
wire n_1361, n_1362, n_1363, n_1364, n_1365, n_1367, n_1368, n_1369;
wire n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1359, n_1360;
wire n_1341, n_1343, n_1344, n_1345, n_1346, n_1347, n_1350, n_1351;
wire n_1331, n_1332, n_1333, n_1334, n_1336, n_1338, n_1339, n_1340;
wire n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330;
wire n_1313, n_1314, n_1315, n_1316, n_1317, n_1319, n_1320, n_1321;
wire n_1304, n_1305, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312;
wire n_1294, n_1296, n_1297, n_1298, n_1299, n_1300, n_1302, n_1303;
wire n_1279, n_1282, n_1283, n_1284, n_1287, n_1289, n_1290, n_1292;
wire n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277;
wire n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268;
wire n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260;
wire n_1243, n_1244, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251;
wire n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241;
wire n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233;
wire n_1217, n_1218, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225;
wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
wire n_1198, n_1199, n_1200, n_1202, n_1203, n_1204, n_1206, n_1207;
wire n_1184, n_1185, n_1189, n_1190, n_1193, n_1194, n_1195, n_1197;
wire n_1172, n_1173, n_1175, n_1177, n_1178, n_1179, n_1182, n_1183;
wire n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171;
wire n_1154, n_1156, n_1157, n_1158, n_1159, n_1160, n_1162, n_1163;
wire n_1142, n_1143, n_1144, n_1145, n_1148, n_1149, n_1150, n_1153;
wire n_1133, n_1134, n_1135, n_1136, n_1137, n_1139, n_1140, n_1141;
wire n_1120, n_1121, n_1123, n_1124, n_1125, n_1126, n_1131, n_1132;
wire n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1117, n_1119;
wire n_1099, n_1100, n_1101, n_1102, n_1104, n_1106, n_1107, n_1108;
wire n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098;
wire n_1081, n_1082, n_1083, n_1085, n_1087, n_1088, n_1089, n_1090;
wire n_1072, n_1073, n_1074, n_1075, n_1076, n_1078, n_1079, n_1080;
wire n_1061, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070;
wire n_1045, n_1047, n_1048, n_1049, n_1052, n_1054, n_1056, n_1058;
wire n_1035, n_1036, n_1037, n_1040, n_1041, n_1042, n_1043, n_1044;
wire n_1023, n_1026, n_1027, n_1029, n_1030, n_1031, n_1032, n_1033;
wire n_1013, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1022;
wire n_1002, n_1003, n_1004, n_1006, n_1007, n_1009, n_1011, n_1012;
wire n_991, n_992, n_994, n_997, n_998, n_999, n_1000, n_1001;
wire n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_989;
wire n_963, n_965, n_967, n_969, n_972, n_973, n_978, n_979;
wire n_951, n_953, n_954, n_955, n_956, n_957, n_959, n_962;
wire n_939, n_940, n_943, n_944, n_946, n_947, n_949, n_950;
wire n_925, n_926, n_927, n_928, n_929, n_931, n_934, n_937;
wire n_911, n_912, n_914, n_915, n_917, n_918, n_921, n_922;
wire n_897, n_898, n_900, n_902, n_903, n_905, n_908, n_910;
wire n_880, n_886, n_888, n_889, n_892, n_893, n_895, n_896;
wire n_869, n_870, n_871, n_873, n_874, n_877, n_878, n_879;
wire n_855, n_856, n_858, n_861, n_862, n_863, n_864, n_865;
wire n_846, n_847, n_849, n_850, n_851, n_852, n_853, n_854;
wire n_831, n_832, n_833, n_835, n_840, n_842, n_844, n_845;
wire n_820, n_824, n_825, n_826, n_827, n_828, n_829, n_830;
wire n_806, n_808, n_809, n_810, n_811, n_812, n_814, n_817;
wire n_795, n_796, n_799, n_800, n_801, n_802, n_804, n_805;
wire n_779, n_780, n_781, n_782, n_787, n_788, n_790, n_794;
wire n_761, n_762, n_763, n_764, n_765, n_767, n_773, n_774;
wire n_746, n_747, n_748, n_752, n_753, n_757, n_758, n_760;
wire n_733, n_734, n_735, n_736, n_739, n_741, n_743, n_744;
wire n_721, n_722, n_724, n_725, n_727, n_728, n_731, n_732;
wire n_708, n_710, n_711, n_714, n_715, n_716, n_718, n_720;
wire n_688, n_693, n_696, n_698, n_701, n_704, n_706, n_707;
wire n_680, n_681, n_682, n_683, n_684, n_685, n_686, n_687;
wire n_663, n_664, n_665, n_666, n_667, n_668, n_670, n_679;
wire n_649, n_650, n_651, n_652, n_653, n_654, n_657, n_658;
wire n_635, n_636, n_637, n_638, n_639, n_640, n_641, n_647;
wire n_622, n_625, n_628, n_629, n_630, n_631, n_632, n_634;
wire n_609, n_611, n_612, n_614, n_615, n_618, n_619, n_620;
wire n_600, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
wire n_592, n_593, n_594, n_595, n_596, n_597, n_598, n_599;
wire n_579, n_584, n_585, n_586, n_587, n_588, n_589, n_590;
wire n_562, n_563, n_564, n_565, n_567, n_571, n_572, n_578;
wire n_551, n_552, n_553, n_554, n_555, n_557, n_558, n_561;
wire n_540, n_543, n_544, n_545, n_546, n_547, n_549, n_550;
wire n_525, n_527, n_528, n_529, n_535, n_536, n_538, n_539;
wire n_502, n_513, n_515, n_516, n_521, n_522, n_523, n_524;
wire n_492, n_493, n_494, n_496, n_497, n_498, n_499, n_500;
wire n_477, n_479, n_481, n_482, n_485, n_488, n_489, n_491;
wire n_463, n_464, n_465, n_466, n_472, n_474, n_475, n_476;
wire n_450, n_451, n_452, n_453, n_454, n_455, n_457, n_458;
wire n_435, n_439, n_440, n_441, n_442, n_443, n_447, n_449;
wire n_421, n_424, n_428, n_430, n_431, n_432, n_433, n_434;
wire n_410, n_411, n_412, n_414, n_415, n_416, n_417, n_419;
wire n_396, n_397, n_399, n_400, n_403, n_405, n_406, n_409;
wire n_387, n_388, n_389, n_390, n_392, n_393, n_394, n_395;
wire n_375, n_376, n_377, n_379, n_380, n_381, n_382, n_384;
wire n_362, n_363, n_365, n_366, n_367, n_371, n_372, n_373;
wire n_343, n_345, n_346, n_349, n_352, n_354, n_358, n_361;
wire n_331, n_333, n_334, n_335, n_336, n_338, n_339, n_341;
wire n_319, n_320, n_321, n_322, n_323, n_324, n_327, n_330;
wire n_301, n_303, n_304, n_307, n_309, n_311, n_316, n_318;
wire n_287, n_288, n_289, n_290, n_294, n_295, n_296, n_300;
wire n_273, n_274, n_275, n_277, n_279, n_282, n_284, n_286;
wire n_263, n_265, n_266, n_267, n_268, n_269, n_271, n_272;
wire n_241, n_242, n_243, n_247, n_252, n_259, n_261, n_262;
wire n_228, n_229, n_230, n_231, n_233, n_235, n_237, n_238;
wire n_210, n_211, n_212, n_215, n_216, n_218, n_224, n_225;
wire n_200, n_201, n_202, n_203, n_204, n_205, n_207, n_209;
wire n_185, n_188, n_190, n_191, n_192, n_194, n_196, n_198;
wire n_167, n_168, n_169, n_171, n_172, n_173, n_174, n_182;
wire n_150, n_151, n_153, n_154, n_156, n_158, n_164, n_165;
wire n_141, n_142, n_143, n_144, n_146, n_147, n_148, n_149;
wire n_122, n_125, n_126, n_127, n_130, n_134, n_137, n_138;
wire n_113, n_114, n_115, n_116, n_117, n_118, n_120, n_121;
wire n_95, n_96, n_99, n_100, n_101, n_103, n_109, n_110;
wire n_74, n_75, n_77, n_79, n_83, n_85, n_88, n_94;
wire n_64, n_65, n_66, n_68, n_69, n_70, n_72, n_73;
wire n_49, n_50, n_52, n_54, n_56, n_60, n_61, n_62;
wire n_33, n_34, n_35, n_36, n_40, n_41, n_45, n_46;
wire n_17, n_19, n_21, n_22, n_25, n_28, n_31, n_32;
wire n_3, n_5, n_6, n_7, n_10, n_11, n_13, n_15;
wire datao_2[25], datao_2[26], datao_2[27], datao_2[29], datao_2[31], n_0, n_1, n_2;
wire datao_2[16], datao_2[17], datao_2[18], datao_2[19], datao_2[20], datao_2[21], datao_2[22], datao_2[23] ;
wire datao_2[6], datao_2[7], datao_2[8], datao_2[9], datao_2[10], datao_2[13], datao_2[14], datao_2[15] ;
wire datao_1[30], datao_1[31], datao_2[0], datao_2[1], datao_2[2], datao_2[3], datao_2[4], datao_2[5] ;
wire datao_1[10], datao_1[11], datao_1[19], datao_1[23], datao_1[24], datao_1[27], datao_1[28], datao_1[29] ;
wire addr_496, addr_497, datao_1[0], datao_1[1], datao_1[4], datao_1[5], datao_1[7], datao_1[9] ;
wire addr_487, addr_488, addr_489, addr_490, addr_491, addr_492, addr_494, addr_495;
wire addr_454, addr_455, addr_456, addr_457, addr_461, addr_483, addr_484, addr_485;
wire addr_444, addr_445, addr_446, addr_447, addr_450, addr_451, addr_452, addr_453;
wire addr_435, addr_436, addr_437, addr_438, addr_439, addr_441, addr_442, addr_443;
wire addr_425, addr_426, addr_429, addr_430, addr_431, addr_432, addr_433, addr_434;
wire P3_reg_150, P3_reg_151, P3_reg_152, P3_reg_153, addr_1, addr_2, addr_3, addr_424;
wire P3_reg3[26], P3_reg3[27], P3_reg3[28], P3_reg_145, P3_reg_146, P3_reg_147, P3_reg_148, P3_reg_149;
wire P3_reg3[18], P3_reg3[19], P3_reg3[20], P3_reg3[21], P3_reg3[22], P3_reg3[23], P3_reg3[24], P3_reg3[25] ;
wire P3_reg3[10], P3_reg3[11], P3_reg3[12], P3_reg3[13], P3_reg3[14], P3_reg3[15], P3_reg3[16], P3_reg3[17] ;
wire P3_reg3[2], P3_reg3[3], P3_reg3[4], P3_reg3[5], P3_reg3[6], P3_reg3[7], P3_reg3[8], P3_reg3[9] ;
wire P3_reg2[10], P3_reg2[13], P3_reg2[15], P3_reg2[18], P3_reg2[28], P3_reg2[29], P3_reg2[30], P3_reg3[0] ;
wire P3_reg1[12], P3_reg1[15], P3_reg1[16], P3_reg1[17], P3_reg1[18], P3_reg1[26], P3_reg2[6], P3_reg2[9] ;
wire P3_reg1[1], P3_reg1[3], P3_reg1[4], P3_reg1[5], P3_reg1[6], P3_reg1[7], P3_reg1[9], P3_reg1[11] ;
wire P3_d_400, P3_d_401, P3_d_402, P3_d_403, P3_d_404, P3_d_405, P3_d_406, P3_d_407;
wire P3_d_392, P3_d_393, P3_d_394, P3_d_395, P3_d_396, P3_d_397, P3_d_398, P3_d_399;
wire P3_d_384, P3_d_385, P3_d_386, P3_d_387, P3_d_388, P3_d_389, P3_d_390, P3_d_391;
wire P3_d, P3_d_377, P3_d_378, P3_d_379, P3_d_380, P3_d_381, P3_d_382, P3_d_383;
wire P3_IR[23], P3_IR[24], P3_IR[25], P3_IR[26], P3_IR[27], P3_IR[28], P3_IR[30], P3_IR[31] ;
wire P3_IR[15], P3_IR[16], P3_IR[17], P3_IR[18], P3_IR[19], P3_IR[20], P3_IR[21], P3_IR[22] ;
wire P3_IR[7], P3_IR[8], P3_IR[9], P3_IR[10], P3_IR[11], P3_IR[12], P3_IR[13], P3_IR[14] ;
wire P3_B, P3_IR[0], P3_IR[1], P3_IR[2], P3_IR[3], P3_IR[4], P3_IR[5], P3_IR[6] ;
wire P2_reg_106, P2_reg_107, P2_reg_108, P2_reg_109, P2_reg_110, P2_reg_111, P2_reg_112, P2_reg_113;
wire P2_reg3[23], P2_reg3[24], P2_reg3[25], P2_reg3[26], P2_reg3[27], P2_reg3[28], P2_reg_95, P2_reg_104;
wire P2_reg3[15], P2_reg3[16], P2_reg3[17], P2_reg3[18], P2_reg3[19], P2_reg3[20], P2_reg3[21], P2_reg3[22] ;
wire P2_reg3[5], P2_reg3[6], P2_reg3[7], P2_reg3[10], P2_reg3[11], P2_reg3[12], P2_reg3[13], P2_reg3[14] ;
wire P2_reg2[25], P2_reg2[26], P2_reg2[27], P2_reg2[28], P2_reg2[29], P2_reg3[1], P2_reg3[3], P2_reg3[4] ;
wire P2_reg2[10], P2_reg2[11], P2_reg2[12], P2_reg2[15], P2_reg2[16], P2_reg2[18], P2_reg2[19], P2_reg2[24] ;
wire P2_reg1[28], P2_reg1[29], P2_reg1[31], P2_reg2[1], P2_reg2[2], P2_reg2[3], P2_reg2[8], P2_reg2[9] ;
wire P2_reg1[19], P2_reg1[20], P2_reg1[21], P2_reg1[22], P2_reg1[23], P2_reg1[25], P2_reg1[26], P2_reg1[27] ;
wire P2_reg1[10], P2_reg1[11], P2_reg1[12], P2_reg1[13], P2_reg1[15], P2_reg1[16], P2_reg1[17], P2_reg1[18] ;
wire P2_reg1[1], P2_reg1[2], P2_reg1[3], P2_reg1[4], P2_reg1[5], P2_reg1[6], P2_reg1[8], P2_reg1[9] ;
wire P2_d_402, P2_d_403, P2_d_404, P2_d_405, P2_d_406, P2_d_407, P2_d_408, P2_n_749;
wire P2_d_394, P2_d_395, P2_d_396, P2_d_397, P2_d_398, P2_d_399, P2_d_400, P2_d_401;
wire P2_d_386, P2_d_387, P2_d_388, P2_d_389, P2_d_390, P2_d_391, P2_d_392, P2_d_393;
wire P2_d_378, P2_d_379, P2_d_380, P2_d_381, P2_d_382, P2_d_383, P2_d_384, P2_d_385;
wire P2_IR[25], P2_IR[26], P2_IR[27], P2_IR[28], P2_IR[29], P2_IR[30], P2_IR[31], P2_d;
wire P2_IR[17], P2_IR[18], P2_IR[19], P2_IR[20], P2_IR[21], P2_IR[22], P2_IR[23], P2_IR[24] ;
wire P2_IR[9], P2_IR[10], P2_IR[11], P2_IR[12], P2_IR[13], P2_IR[14], P2_IR[15], P2_IR[16] ;
wire P2_IR[1], P2_IR[2], P2_IR[3], P2_IR[4], P2_IR[5], P2_IR[6], P2_IR[7], P2_IR[8] ;
wire P1_reg_175, P1_reg_176, P1_reg_177, P1_reg_178, P1_reg_179, P1_reg_180, P2_B, P2_IR[0] ;
wire P1_reg3[24], P1_reg3[25], P1_reg3[26], P1_reg3[27], P1_reg3[28], P1_reg_172, P1_reg_173, P1_reg_174;
wire P1_reg3[16], P1_reg3[17], P1_reg3[18], P1_reg3[19], P1_reg3[20], P1_reg3[21], P1_reg3[22], P1_reg3[23] ;
wire P1_reg3[8], P1_reg3[9], P1_reg3[10], P1_reg3[11], P1_reg3[12], P1_reg3[13], P1_reg3[14], P1_reg3[15] ;
wire P1_reg2[28], P1_reg2[29], P1_reg2[30], P1_reg3[3], P1_reg3[4], P1_reg3[5], P1_reg3[6], P1_reg3[7] ;
wire P1_reg2[9], P1_reg2[14], P1_reg2[16], P1_reg2[19], P1_reg2[24], P1_reg2[25], P1_reg2[26], P1_reg2[27] ;
wire P1_reg1[25], P1_reg1[26], P1_reg1[27], P1_reg1[28], P1_reg1[29], P1_reg1[30], P1_reg2[0], P1_reg2[1] ;
wire P1_n_449, P1_reg1[0], P1_reg1[1], P1_reg1[12], P1_reg1[14], P1_reg1[16], P1_reg1[19], P1_reg1[24] ;
wire P1_d_121, P1_d_122, P1_d_123, P1_d_124, P1_d_125, P1_d_126, P1_d_127, P1_d_128;
wire P1_d_113, P1_d_114, P1_d_115, P1_d_116, P1_d_117, P1_d_118, P1_d_119, P1_d_120;
wire P1_d_105, P1_d_106, P1_d_107, P1_d_108, P1_d_109, P1_d_110, P1_d_111, P1_d_112;
wire P1_d, P1_d_98, P1_d_99, P1_d_100, P1_d_101, P1_d_102, P1_d_103, P1_d_104;
wire P1_IR[24], P1_IR[25], P1_IR[26], P1_IR[27], P1_IR[28], P1_IR[29], P1_IR[30], P1_IR[31] ;
wire P1_IR[16], P1_IR[17], P1_IR[18], P1_IR[19], P1_IR[20], P1_IR[21], P1_IR[22], P1_IR[23] ;
wire P1_IR[8], P1_IR[9], P1_IR[10], P1_IR[11], P1_IR[12], P1_IR[13], P1_IR[14], P1_IR[15] ;
wire P1_IR[0], P1_IR[1], P1_IR[2], P1_IR[3], P1_IR[4], P1_IR[5], P1_IR[6], P1_IR[7] ;
wire rd, wr;
wire [19:0] so;
wire [31:0] si;
wire clock, reset;
CLKBUFX1 gbuf_d_1(.A(n_32009), .Y(d_out_1));
CLKBUFX1 gbuf_qn_1(.A(qn_in_1), .Y(P1_reg2[29]));
CLKBUFX1 gbuf_d_2(.A(n_32006), .Y(d_out_2));
CLKBUFX1 gbuf_qn_2(.A(qn_in_2), .Y(P1_reg1[29]));
CLKBUFX1 gbuf_d_3(.A(n_32007), .Y(d_out_3));
CLKBUFX1 gbuf_q_3(.A(q_in_3), .Y(P2_reg2[29]));
CLKBUFX1 gbuf_d_4(.A(n_32008), .Y(d_out_4));
CLKBUFX1 gbuf_q_4(.A(q_in_4), .Y(P3_reg2[28]));
CLKBUFX1 gbuf_d_5(.A(n_32005), .Y(d_out_5));
CLKBUFX1 gbuf_q_5(.A(q_in_5), .Y(P3_reg2[29]));
CLKBUFX1 gbuf_d_6(.A(n_32004), .Y(d_out_6));
CLKBUFX1 gbuf_q_6(.A(q_in_6), .Y(n_12670));
CLKBUFX1 gbuf_d_7(.A(n_32002), .Y(d_out_7));
CLKBUFX1 gbuf_qn_7(.A(qn_in_7), .Y(P2_reg_113));
CLKBUFX1 gbuf_d_8(.A(n_32001), .Y(d_out_8));
CLKBUFX1 gbuf_qn_8(.A(qn_in_8), .Y(P2_reg1[29]));
CLKBUFX1 gbuf_d_9(.A(n_31999), .Y(d_out_9));
CLKBUFX1 gbuf_q_9(.A(q_in_9), .Y(n_13689));
CLKBUFX1 gbuf_d_10(.A(n_32000), .Y(d_out_10));
CLKBUFX1 gbuf_q_10(.A(q_in_10), .Y(n_524));
CLKBUFX1 gbuf_d_11(.A(n_31998), .Y(d_out_11));
CLKBUFX1 gbuf_q_11(.A(q_in_11), .Y(n_13690));
NAND2X1 g105376(.A (n_35640), .B (n_35641), .Y (n_32009));
NAND2X2 g105394(.A (n_32068), .B (n_32069), .Y (n_32008));
CLKBUFX1 gbuf_d_12(.A(n_31993), .Y(d_out_12));
CLKBUFX1 gbuf_q_12(.A(q_in_12), .Y(P3_reg3[28]));
CLKBUFX1 gbuf_d_13(.A(n_31989), .Y(d_out_13));
CLKBUFX1 gbuf_q_13(.A(q_in_13), .Y(n_13330));
CLKBUFX1 gbuf_d_14(.A(n_34704), .Y(d_out_14));
CLKBUFX1 gbuf_q_14(.A(q_in_14), .Y(P2_B));
CLKBUFX1 gbuf_d_15(.A(n_31992), .Y(d_out_15));
CLKBUFX1 gbuf_q_15(.A(q_in_15), .Y(P1_reg3[28]));
CLKBUFX1 gbuf_d_16(.A(n_31990), .Y(d_out_16));
CLKBUFX1 gbuf_q_16(.A(q_in_16), .Y(P2_reg1[27]));
CLKBUFX1 gbuf_d_17(.A(n_31988), .Y(d_out_17));
CLKBUFX1 gbuf_qn_17(.A(qn_in_17), .Y(P1_reg1[25]));
NAND2X2 g105396(.A (n_32281), .B (n_32282), .Y (n_32007));
NAND2X2 g105398(.A (n_32893), .B (n_32894), .Y (n_32006));
NAND2X2 g105434(.A (n_32072), .B (n_32073), .Y (n_32005));
NAND2X1 g105392(.A (n_31975), .B (n_12858), .Y (n_32004));
NAND2X1 g105391(.A (n_31985), .B (n_31201), .Y (n_35640));
CLKBUFX1 gbuf_d_18(.A(n_31980), .Y(d_out_18));
CLKBUFX1 gbuf_q_18(.A(q_in_18), .Y(n_13201));
CLKBUFX1 gbuf_d_19(.A(n_31973), .Y(d_out_19));
CLKBUFX1 gbuf_q_19(.A(q_in_19), .Y(n_13334));
CLKBUFX1 gbuf_d_20(.A(n_31976), .Y(d_out_20));
CLKBUFX1 gbuf_q_20(.A(q_in_20), .Y(n_13344));
CLKBUFX1 gbuf_d_21(.A(n_31969), .Y(d_out_21));
CLKBUFX1 gbuf_qn_21(.A(qn_in_21), .Y(P1_reg_179));
CLKBUFX1 gbuf_d_22(.A(n_31981), .Y(d_out_22));
CLKBUFX1 gbuf_q_22(.A(q_in_22), .Y(P3_reg3[25]));
CLKBUFX1 gbuf_d_23(.A(n_31971), .Y(d_out_23));
CLKBUFX1 gbuf_qn_23(.A(qn_in_23), .Y(P1_reg1[28]));
CLKBUFX1 gbuf_d_24(.A(n_31970), .Y(d_out_24));
CLKBUFX1 gbuf_qn_24(.A(qn_in_24), .Y(P1_reg2[27]));
CLKBUFX1 gbuf_d_25(.A(n_31968), .Y(d_out_25));
CLKBUFX1 gbuf_qn_25(.A(qn_in_25), .Y(P1_reg2[28]));
CLKBUFX1 gbuf_d_26(.A(n_34675), .Y(d_out_26));
CLKBUFX1 gbuf_qn_26(.A(qn_in_26), .Y(P1_reg_178));
CLKBUFX1 gbuf_d_27(.A(n_31972), .Y(d_out_27));
CLKBUFX1 gbuf_q_27(.A(q_in_27), .Y(n_13336));
CLKBUFX1 gbuf_d_28(.A(n_31974), .Y(d_out_28));
CLKBUFX1 gbuf_q_28(.A(q_in_28), .Y(P3_reg3[20]));
CLKBUFX1 gbuf_d_29(.A(n_31984), .Y(d_out_29));
CLKBUFX1 gbuf_q_29(.A(q_in_29), .Y(P1_reg_174));
CLKBUFX1 gbuf_d_30(.A(n_31983), .Y(d_out_30));
CLKBUFX1 gbuf_q_30(.A(q_in_30), .Y(P1_reg1[24]));
NAND2X2 g105429(.A (n_32248), .B (n_32249), .Y (n_32002));
NAND2X2 g105430(.A (n_32263), .B (n_32264), .Y (n_32001));
NAND2X1 g105500(.A (n_6761), .B (n_31987), .Y (n_32000));
NAND2X1 g105433(.A (n_32166), .B (n_32167), .Y (n_31999));
NAND2X1 g105501(.A (n_6732), .B (n_31986), .Y (n_31998));
NAND2X2 g105416(.A (n_917), .B (n_35889), .Y (n_32068));
NAND2X1 g105418(.A (n_31345), .B (n_35614), .Y (n_32281));
NAND2X1 g105419(.A (n_31912), .B (n_35291), .Y (n_32893));
CLKBUFX1 gbuf_d_31(.A(n_31959), .Y(d_out_31));
CLKBUFX1 gbuf_q_31(.A(q_in_31), .Y(P3_reg3[24]));
CLKBUFX1 gbuf_d_32(.A(n_33728), .Y(d_out_32));
CLKBUFX1 gbuf_qn_32(.A(qn_in_32), .Y(P1_reg2[25]));
CLKBUFX1 gbuf_d_33(.A(n_31945), .Y(d_out_33));
CLKBUFX1 gbuf_q_33(.A(q_in_33), .Y(P2_reg3[27]));
CLKBUFX1 gbuf_d_34(.A(n_31942), .Y(d_out_34));
CLKBUFX1 gbuf_q_34(.A(q_in_34), .Y(P3_reg3[27]));
CLKBUFX1 gbuf_d_35(.A(n_31950), .Y(d_out_35));
CLKBUFX1 gbuf_qn_35(.A(qn_in_35), .Y(P1_reg1[27]));
CLKBUFX1 gbuf_d_36(.A(n_31949), .Y(d_out_36));
CLKBUFX1 gbuf_qn_36(.A(qn_in_36), .Y(P2_reg_109));
CLKBUFX1 gbuf_d_37(.A(n_31948), .Y(d_out_37));
CLKBUFX1 gbuf_qn_37(.A(qn_in_37), .Y(P2_reg1[25]));
CLKBUFX1 gbuf_d_38(.A(n_31946), .Y(d_out_38));
CLKBUFX1 gbuf_qn_38(.A(qn_in_38), .Y(P1_reg_177));
CLKBUFX1 gbuf_d_39(.A(n_31954), .Y(d_out_39));
CLKBUFX1 gbuf_q_39(.A(q_in_39), .Y(n_13368));
CLKBUFX1 gbuf_d_40(.A(n_31962), .Y(d_out_40));
CLKBUFX1 gbuf_q_40(.A(q_in_40), .Y(P1_reg3[24]));
CLKBUFX1 gbuf_d_41(.A(n_34307), .Y(d_out_41));
CLKBUFX1 gbuf_q_41(.A(q_in_41), .Y(P2_reg3[24]));
CLKBUFX1 gbuf_d_42(.A(n_31955), .Y(d_out_42));
CLKBUFX1 gbuf_q_42(.A(q_in_42), .Y(P1_reg3[27]));
CLKBUFX1 gbuf_d_43(.A(n_34382), .Y(d_out_43));
CLKBUFX1 gbuf_qn_43(.A(qn_in_43), .Y(P2_reg2[24]));
NAND2X1 g105480(.A (n_31951), .B (n_35609), .Y (n_32072));
OAI21X1 g105397(.A0 (n_31901), .A1 (n_31569), .B0 (n_7604), .Y(n_31993));
NAND2X2 g105426(.A (n_32317), .B (n_32318), .Y (n_31992));
NAND2X2 g105496(.A (n_35145), .B (n_35146), .Y (n_31990));
NAND2X2 g105432(.A (n_32252), .B (n_32253), .Y (n_31989));
NAND2X2 g105503(.A (n_35276), .B (n_35277), .Y (n_31988));
NAND2X1 g105540(.A (n_31932), .B (n_31783), .Y (n_31987));
NAND2X1 g105541(.A (n_31937), .B (n_31850), .Y (n_31986));
OAI21X1 g105417(.A0 (n_8584), .A1 (n_30691), .B0 (n_31910), .Y(n_31985));
NAND2X1 g105716(.A (n_7030), .B (n_31913), .Y (n_31984));
NAND2X1 g105721(.A (n_7119), .B (n_31909), .Y (n_31983));
NAND2X1 g105473(.A (n_31928), .B (n_31922), .Y (n_32166));
OAI21X1 g105421(.A0 (n_31871), .A1 (n_31979), .B0 (n_7402), .Y(n_31981));
OAI21X1 g105395(.A0 (n_31979), .A1 (n_35290), .B0 (n_6471), .Y(n_31980));
CLKBUFX1 gbuf_d_44(.A(n_31914), .Y(d_out_44));
CLKBUFX1 gbuf_q_44(.A(q_in_44), .Y(n_13343));
CLKBUFX1 gbuf_d_45(.A(n_31905), .Y(d_out_45));
CLKBUFX1 gbuf_q_45(.A(q_in_45), .Y(P3_reg3[19]));
CLKBUFX1 gbuf_d_46(.A(n_31911), .Y(d_out_46));
CLKBUFX1 gbuf_qn_46(.A(qn_in_46), .Y(P2_reg_111));
CLKBUFX1 gbuf_d_47(.A(n_33200), .Y(d_out_47));
CLKBUFX1 gbuf_qn_47(.A(qn_in_47), .Y(P2_reg1[28]));
CLKBUFX1 gbuf_d_48(.A(n_33349), .Y(d_out_48));
CLKBUFX1 gbuf_qn_48(.A(qn_in_48), .Y(P2_reg_112));
CLKBUFX1 gbuf_d_49(.A(n_31904), .Y(d_out_49));
CLKBUFX1 gbuf_qn_49(.A(qn_in_49), .Y(P2_reg2[27]));
CLKBUFX1 gbuf_d_50(.A(n_31902), .Y(d_out_50));
CLKBUFX1 gbuf_qn_50(.A(qn_in_50), .Y(P1_reg_175));
CLKBUFX1 gbuf_d_51(.A(n_31903), .Y(d_out_51));
CLKBUFX1 gbuf_qn_51(.A(qn_in_51), .Y(P2_reg2[28]));
CLKBUFX1 gbuf_d_52(.A(n_31900), .Y(d_out_52));
CLKBUFX1 gbuf_q_52(.A(q_in_52), .Y(n_13695));
CLKBUFX1 gbuf_d_53(.A(n_31920), .Y(d_out_53));
CLKBUFX1 gbuf_q_53(.A(q_in_53), .Y(P3_reg3[21]));
CLKBUFX1 gbuf_d_54(.A(n_31915), .Y(d_out_54));
CLKBUFX1 gbuf_q_54(.A(q_in_54), .Y(n_13335));
CLKBUFX1 gbuf_d_55(.A(n_31919), .Y(d_out_55));
CLKBUFX1 gbuf_q_55(.A(q_in_55), .Y(P3_reg3[22]));
CLKBUFX1 gbuf_d_56(.A(n_31916), .Y(d_out_56));
CLKBUFX1 gbuf_q_56(.A(q_in_56), .Y(P2_reg3[28]));
CLKBUFX1 gbuf_d_57(.A(n_31917), .Y(d_out_57));
CLKBUFX1 gbuf_q_57(.A(q_in_57), .Y(P1_reg3[25]));
CLKBUFX1 gbuf_d_58(.A(n_31929), .Y(d_out_58));
CLKBUFX1 gbuf_q_58(.A(q_in_58), .Y(P2_reg_108));
CLKBUFX1 gbuf_d_59(.A(n_31927), .Y(d_out_59));
CLKBUFX1 gbuf_q_59(.A(q_in_59), .Y(P2_reg1[22]));
CLKBUFX1 gbuf_d_60(.A(n_31926), .Y(d_out_60));
CLKBUFX1 gbuf_q_60(.A(q_in_60), .Y(n_9231));
CLKBUFX1 gbuf_d_61(.A(n_31925), .Y(d_out_61));
CLKBUFX1 gbuf_qn_61(.A(qn_in_61), .Y(P1_reg2[24]));
CLKBUFX1 gbuf_d_62(.A(n_31924), .Y(d_out_62));
CLKBUFX1 gbuf_q_62(.A(q_in_62), .Y(n_13687));
NAND2X2 g105481(.A (n_34737), .B (n_31493), .Y (n_32248));
NAND2X1 g105482(.A (n_31930), .B (n_31965), .Y (n_32263));
NAND2X2 g105424(.A (n_6477), .B (n_31923), .Y (n_31976));
NOR2X1 g105425(.A (n_1943), .B (n_31907), .Y (n_31975));
OAI21X1 g105488(.A0 (n_31877), .A1 (n_31958), .B0 (n_7419), .Y(n_31974));
NAND2X2 g105428(.A (n_32157), .B (n_32158), .Y (n_31973));
NAND2X1 g105492(.A (n_6667), .B (n_31939), .Y (n_31972));
NAND2X2 g105494(.A (n_32883), .B (n_32884), .Y (n_31971));
NAND2X2 g105495(.A (n_32271), .B (n_32272), .Y (n_31970));
NAND2X1 g105431(.A (n_6923), .B (n_31921), .Y (n_31969));
NAND2X2 g105497(.A (n_32556), .B (n_32557), .Y (n_31968));
NAND2X2 g105536(.A (n_31965), .B (n_35292), .Y (n_35145));
NAND2X1 g105542(.A (n_31882), .B (n_31891), .Y (n_35276));
OAI21X1 g105549(.A0 (n_31800), .A1 (n_31726), .B0 (n_7249), .Y(n_31962));
OAI21X1 g105551(.A0 (n_31801), .A1 (n_31936), .B0 (n_10440), .Y(n_35609));
NAND2X1 g105469(.A (n_35023), .B (n_35615), .Y (n_32317));
OAI21X1 g105420(.A0 (n_31820), .A1 (n_31958), .B0 (n_7420), .Y(n_31959));
CLKBUFX1 gbuf_d_63(.A(n_31868), .Y(d_out_63));
CLKBUFX1 gbuf_q_63(.A(q_in_63), .Y(P3_reg3[26]));
CLKBUFX1 gbuf_d_64(.A(n_31860), .Y(d_out_64));
CLKBUFX1 gbuf_q_64(.A(q_in_64), .Y(n_13348));
CLKBUFX1 gbuf_d_65(.A(n_31858), .Y(d_out_65));
CLKBUFX1 gbuf_q_65(.A(q_in_65), .Y(n_13692));
CLKBUFX1 gbuf_d_66(.A(n_33458), .Y(d_out_66));
CLKBUFX1 gbuf_q_66(.A(q_in_66), .Y(P1_reg3[26]));
CLKBUFX1 gbuf_d_67(.A(n_31862), .Y(d_out_67));
CLKBUFX1 gbuf_q_67(.A(q_in_67), .Y(n_13353));
CLKBUFX1 gbuf_d_68(.A(n_31861), .Y(d_out_68));
CLKBUFX1 gbuf_q_68(.A(q_in_68), .Y(n_13698));
CLKBUFX1 gbuf_d_69(.A(n_31863), .Y(d_out_69));
CLKBUFX1 gbuf_q_69(.A(q_in_69), .Y(n_13354));
CLKBUFX1 gbuf_d_70(.A(n_31869), .Y(d_out_70));
CLKBUFX1 gbuf_q_70(.A(q_in_70), .Y(n_13329));
CLKBUFX1 gbuf_d_71(.A(n_31867), .Y(d_out_71));
CLKBUFX1 gbuf_q_71(.A(q_in_71), .Y(n_13352));
CLKBUFX1 gbuf_d_72(.A(n_31873), .Y(d_out_72));
CLKBUFX1 gbuf_q_72(.A(q_in_72), .Y(n_13359));
CLKBUFX1 gbuf_d_73(.A(n_35022), .Y(d_out_73));
CLKBUFX1 gbuf_q_73(.A(q_in_73), .Y(P1_reg3[20]));
CLKBUFX1 gbuf_d_74(.A(n_31886), .Y(d_out_74));
CLKBUFX1 gbuf_q_74(.A(q_in_74), .Y(P2_reg3[17]));
CLKBUFX1 gbuf_d_75(.A(n_31885), .Y(d_out_75));
CLKBUFX1 gbuf_q_75(.A(q_in_75), .Y(P2_reg3[19]));
CLKBUFX1 gbuf_d_76(.A(n_31887), .Y(d_out_76));
CLKBUFX1 gbuf_q_76(.A(q_in_76), .Y(P1_reg3[17]));
CLKBUFX1 gbuf_d_77(.A(n_34195), .Y(d_out_77));
CLKBUFX1 gbuf_q_77(.A(q_in_77), .Y(P3_reg3[18]));
CLKBUFX1 gbuf_d_78(.A(n_31857), .Y(d_out_78));
CLKBUFX1 gbuf_q_78(.A(q_in_78), .Y(n_10893));
CLKBUFX1 gbuf_d_79(.A(n_31859), .Y(d_out_79));
CLKBUFX1 gbuf_q_79(.A(q_in_79), .Y(n_11120));
CLKBUFX1 gbuf_d_80(.A(n_31897), .Y(d_out_80));
CLKBUFX1 gbuf_q_80(.A(q_in_80), .Y(n_13673));
CLKBUFX1 gbuf_d_81(.A(n_31896), .Y(d_out_81));
CLKBUFX1 gbuf_q_81(.A(q_in_81), .Y(n_13699));
CLKBUFX1 gbuf_d_82(.A(n_31865), .Y(d_out_82));
CLKBUFX1 gbuf_q_82(.A(q_in_82), .Y(P1_reg3[19]));
OAI21X1 g105476(.A0 (n_9839), .A1 (n_31536), .B0 (n_31879), .Y(n_35889));
OAI21X1 g105477(.A0 (n_9291), .A1 (n_35012), .B0 (n_31875), .Y(n_35614));
NAND2X2 g105564(.A (n_35264), .B (n_35265), .Y (n_31955));
NAND2X1 g105565(.A (n_6549), .B (n_31890), .Y (n_31954));
NAND2X1 g105479(.A (n_31874), .B (n_31951), .Y (n_32252));
NAND2X1 g105571(.A (n_6951), .B (n_31895), .Y (n_31950));
NAND2X2 g105572(.A (n_35101), .B (n_35102), .Y (n_31949));
NAND2X1 g105575(.A (n_6585), .B (n_31888), .Y (n_31948));
OAI21X1 g105486(.A0 (n_8600), .A1 (n_31881), .B0 (n_31872), .Y(n_35291));
NAND2X1 g105582(.A (n_32925), .B (n_32926), .Y (n_31946));
OAI21X1 g105490(.A0 (n_31836), .A1 (n_34300), .B0 (n_6885), .Y(n_31945));
NAND2X1 g105493(.A (n_7391), .B (n_31893), .Y (n_31942));
NAND2X1 g105529(.A (n_31894), .B (n_35899), .Y (n_32883));
NAND2X1 g105532(.A (n_31840), .B (n_31774), .Y (n_31939));
OAI21X1 g105695(.A0 (n_31766), .A1 (n_31936), .B0 (n_10356), .Y(n_31937));
NAND2X2 g105537(.A (n_31933), .B (n_35618), .Y (n_32556));
NAND2X2 g105538(.A (n_31933), .B (n_35890), .Y (n_32271));
OAI21X1 g105700(.A0 (n_31765), .A1 (n_31936), .B0 (n_10368), .Y(n_31932));
OAI21X1 g105545(.A0 (n_9308), .A1 (n_31740), .B0 (n_31827), .Y(n_31930));
NAND2X1 g105709(.A (n_35880), .B (n_35881), .Y (n_31929));
OAI21X1 g105548(.A0 (n_31733), .A1 (n_31936), .B0 (n_10384), .Y(n_31928));
NAND2X2 g105711(.A (n_32056), .B (n_32057), .Y (n_31927));
NAND2X1 g105712(.A (n_6630), .B (n_31813), .Y (n_31926));
NAND2X1 g105714(.A (n_35141), .B (n_35142), .Y (n_31925));
NAND2X1 g105719(.A (n_6601), .B (n_31812), .Y (n_31924));
NAND2X1 g105470(.A (n_31838), .B (n_31922), .Y (n_31923));
OAI21X1 g105472(.A0 (n_31780), .A1 (n_8891), .B0 (n_31845), .Y(n_31921));
OAI21X1 g105555(.A0 (n_31731), .A1 (n_31388), .B0 (n_7253), .Y(n_31920));
NAND2X2 g105556(.A (n_7411), .B (n_31851), .Y (n_31919));
NAND2X1 g105474(.A (n_31835), .B (n_31922), .Y (n_32157));
CLKBUFX1 gbuf_d_83(.A(n_31825), .Y(d_out_83));
CLKBUFX1 gbuf_q_83(.A(q_in_83), .Y(P3_B));
CLKBUFX1 gbuf_d_84(.A(n_31802), .Y(d_out_84));
CLKBUFX1 gbuf_qn_84(.A(qn_in_84), .Y(P1_reg1[26]));
CLKBUFX1 gbuf_d_85(.A(n_31810), .Y(d_out_85));
CLKBUFX1 gbuf_qn_85(.A(qn_in_85), .Y(P1_reg2[26]));
CLKBUFX1 gbuf_d_86(.A(n_31806), .Y(d_out_86));
CLKBUFX1 gbuf_qn_86(.A(qn_in_86), .Y(P1_reg_176));
CLKBUFX1 gbuf_d_87(.A(n_31803), .Y(d_out_87));
CLKBUFX1 gbuf_q_87(.A(q_in_87), .Y(P3_reg1[26]));
CLKBUFX1 gbuf_d_88(.A(n_31824), .Y(d_out_88));
CLKBUFX1 gbuf_qn_88(.A(qn_in_88), .Y(P2_reg2[25]));
CLKBUFX1 gbuf_d_89(.A(n_31826), .Y(d_out_89));
CLKBUFX1 gbuf_q_89(.A(q_in_89), .Y(P2_reg3[25]));
CLKBUFX1 gbuf_d_90(.A(n_34975), .Y(d_out_90));
CLKBUFX1 gbuf_q_90(.A(q_in_90), .Y(P2_reg3[18]));
CLKBUFX1 gbuf_d_91(.A(n_31837), .Y(d_out_91));
CLKBUFX1 gbuf_q_91(.A(q_in_91), .Y(P3_reg3[17]));
CLKBUFX1 gbuf_d_92(.A(n_31853), .Y(d_out_92));
CLKBUFX1 gbuf_q_92(.A(q_in_92), .Y(n_9475));
CLKBUFX1 gbuf_d_93(.A(n_31796), .Y(d_out_93));
CLKBUFX1 gbuf_q_93(.A(q_in_93), .Y(n_9139));
CLKBUFX1 gbuf_d_94(.A(n_31794), .Y(d_out_94));
CLKBUFX1 gbuf_q_94(.A(q_in_94), .Y(P2_reg1[17]));
CLKBUFX1 gbuf_d_95(.A(n_31795), .Y(d_out_95));
CLKBUFX1 gbuf_q_95(.A(q_in_95), .Y(n_11141));
CLKBUFX1 gbuf_d_96(.A(n_31793), .Y(d_out_96));
CLKBUFX1 gbuf_q_96(.A(q_in_96), .Y(P2_reg1[19]));
CLKBUFX1 gbuf_d_97(.A(n_31791), .Y(d_out_97));
CLKBUFX1 gbuf_q_97(.A(q_in_97), .Y(n_13212));
CLKBUFX1 gbuf_d_98(.A(n_31790), .Y(d_out_98));
CLKBUFX1 gbuf_q_98(.A(q_in_98), .Y(n_13203));
CLKBUFX1 gbuf_d_99(.A(n_31856), .Y(d_out_99));
CLKBUFX1 gbuf_q_99(.A(q_in_99), .Y(n_13367));
CLKBUFX1 gbuf_d_100(.A(n_31797), .Y(d_out_100));
CLKBUFX1 gbuf_q_100(.A(q_in_100), .Y(P2_reg2[19]));
CLKBUFX1 gbuf_d_101(.A(n_31792), .Y(d_out_101));
CLKBUFX1 gbuf_q_101(.A(q_in_101), .Y(n_10171));
CLKBUFX1 gbuf_d_102(.A(n_31855), .Y(d_out_102));
CLKBUFX1 gbuf_q_102(.A(q_in_102), .Y(n_13697));
CLKBUFX1 gbuf_d_103(.A(n_31854), .Y(d_out_103));
CLKBUFX1 gbuf_q_103(.A(q_in_103), .Y(n_10167));
CLKBUFX1 gbuf_d_104(.A(n_31799), .Y(d_out_104));
CLKBUFX1 gbuf_q_104(.A(q_in_104), .Y(P2_reg3[21]));
CLKBUFX1 gbuf_d_105(.A(n_31798), .Y(d_out_105));
CLKBUFX1 gbuf_q_105(.A(q_in_105), .Y(P3_reg3[23]));
CLKBUFX1 gbuf_d_106(.A(n_31805), .Y(d_out_106));
CLKBUFX1 gbuf_q_106(.A(q_in_106), .Y(P1_reg3[18]));
CLKBUFX1 gbuf_d_107(.A(n_31804), .Y(d_out_107));
CLKBUFX1 gbuf_q_107(.A(q_in_107), .Y(P3_reg3[16]));
CLKBUFX1 gbuf_d_108(.A(n_31816), .Y(d_out_108));
CLKBUFX1 gbuf_q_108(.A(q_in_108), .Y(P1_reg2[19]));
CLKBUFX1 gbuf_d_109(.A(n_31817), .Y(d_out_109));
CLKBUFX1 gbuf_q_109(.A(q_in_109), .Y(n_4277));
CLKBUFX1 gbuf_d_110(.A(n_31815), .Y(d_out_110));
CLKBUFX1 gbuf_q_110(.A(q_in_110), .Y(n_10217));
CLKBUFX1 gbuf_d_111(.A(n_31829), .Y(d_out_111));
CLKBUFX1 gbuf_q_111(.A(q_in_111), .Y(P3_reg3[13]));
NAND2X1 g105562(.A (n_7414), .B (n_31849), .Y (n_31917));
NAND2X2 g105563(.A (n_35075), .B (n_35076), .Y (n_31916));
NAND2X2 g105567(.A (n_32091), .B (n_32092), .Y (n_31915));
NAND2X1 g105423(.A (n_35906), .B (n_35907), .Y (n_31914));
NAND2X1 g105771(.A (n_31912), .B (n_35932), .Y (n_31913));
NAND2X1 g105573(.A (n_6675), .B (n_31848), .Y (n_31911));
OAI21X1 g105483(.A0 (n_31778), .A1 (n_31090), .B0 (n_31771), .Y(n_31910));
NAND2X1 g105775(.A (n_31822), .B (n_31933), .Y (n_31909));
AOI21X1 g105484(.A0 (n_31768), .A1 (n_31622), .B0 (n_6371), .Y(n_31907));
NAND2X1 g105485(.A (n_31821), .B (n_13003), .Y (n_31905));
NAND2X1 g105578(.A (n_6624), .B (n_31847), .Y (n_31904));
NAND2X2 g105579(.A (n_6629), .B (n_31841), .Y (n_31903));
NAND2X1 g105580(.A (n_6904), .B (n_31846), .Y (n_31902));
AOI22X1 g105489(.A0 (n_31767), .A1 (n_31878), .B0 (n_9167), .B1(n_31876), .Y (n_31901));
NAND2X1 g105587(.A (n_6677), .B (n_31844), .Y (n_31900));
NAND2X1 g105647(.A (n_31714), .B (n_34668), .Y (n_35264));
NAND2X1 g105878(.A (n_6603), .B (n_31777), .Y (n_31897));
NAND2X1 g105880(.A (n_6757), .B (n_31776), .Y (n_31896));
NAND2X1 g105652(.A (n_31742), .B (n_31894), .Y (n_31895));
NAND2X1 g105528(.A (n_31764), .B (n_31694), .Y (n_31893));
NAND2X1 g105658(.A (n_31735), .B (n_31891), .Y (n_32925));
NAND2X1 g105662(.A (n_31748), .B (n_31781), .Y (n_31890));
NAND2X1 g105671(.A (n_31741), .B (n_31965), .Y (n_35101));
NAND2X1 g105672(.A (n_31738), .B (n_31683), .Y (n_31888));
NAND2X1 g105676(.A (n_31728), .B (n_12714), .Y (n_31887));
NAND2X2 g105677(.A (n_31732), .B (n_12883), .Y (n_31886));
NAND2X1 g105679(.A (n_31736), .B (n_12955), .Y (n_31885));
OAI21X1 g105691(.A0 (n_9311), .A1 (n_30731), .B0 (n_31729), .Y(n_35292));
OAI21X1 g105697(.A0 (n_8577), .A1 (n_31881), .B0 (n_31730), .Y(n_31882));
OAI21X1 g105543(.A0 (n_31636), .A1 (n_31016), .B0 (n_31878), .Y(n_31879));
AOI22X1 g105703(.A0 (n_31669), .A1 (n_31878), .B0 (n_9318), .B1(n_31876), .Y (n_31877));
OAI21X1 g105546(.A0 (n_34427), .A1 (n_30909), .B0 (n_31402), .Y(n_31875));
OAI21X1 g105550(.A0 (n_9863), .A1 (n_31834), .B0 (n_31779), .Y(n_31874));
OAI21X1 g105717(.A0 (n_31659), .A1 (n_30792), .B0 (n_6539), .Y(n_31873));
OAI21X1 g105554(.A0 (n_35878), .A1 (n_35879), .B0 (n_31160), .Y(n_31872));
AOI22X1 g105557(.A0 (n_31631), .A1 (n_31878), .B0 (n_9307), .B1(n_31819), .Y (n_31871));
AOI22X1 g105475(.A0 (n_31706), .A1 (n_31878), .B0 (n_9149), .B1(n_31495), .Y (n_35290));
NAND2X1 g105560(.A (n_6607), .B (n_31785), .Y (n_31869));
CLKBUFX1 gbuf_d_112(.A(n_33218), .Y(d_out_112));
CLKBUFX1 gbuf_qn_112(.A(qn_in_112), .Y(P2_reg2[26]));
CLKBUFX1 gbuf_d_113(.A(n_31745), .Y(d_out_113));
CLKBUFX1 gbuf_q_113(.A(q_in_113), .Y(n_13351));
CLKBUFX1 gbuf_d_114(.A(n_31752), .Y(d_out_114));
CLKBUFX1 gbuf_q_114(.A(q_in_114), .Y(P2_reg3[26]));
CLKBUFX1 gbuf_d_115(.A(n_31719), .Y(d_out_115));
CLKBUFX1 gbuf_q_115(.A(q_in_115), .Y(n_9165));
CLKBUFX1 gbuf_d_116(.A(n_31718), .Y(d_out_116));
CLKBUFX1 gbuf_q_116(.A(q_in_116), .Y(P2_reg_106));
CLKBUFX1 gbuf_d_117(.A(n_31717), .Y(d_out_117));
CLKBUFX1 gbuf_q_117(.A(q_in_117), .Y(P2_reg1[18]));
CLKBUFX1 gbuf_d_118(.A(n_31716), .Y(d_out_118));
CLKBUFX1 gbuf_q_118(.A(q_in_118), .Y(n_10897));
CLKBUFX1 gbuf_d_119(.A(n_31712), .Y(d_out_119));
CLKBUFX1 gbuf_q_119(.A(q_in_119), .Y(n_10165));
CLKBUFX1 gbuf_d_120(.A(n_31711), .Y(d_out_120));
CLKBUFX1 gbuf_q_120(.A(q_in_120), .Y(n_13216));
CLKBUFX1 gbuf_d_121(.A(n_31715), .Y(d_out_121));
CLKBUFX1 gbuf_q_121(.A(q_in_121), .Y(n_10610));
CLKBUFX1 gbuf_d_122(.A(n_31720), .Y(d_out_122));
CLKBUFX1 gbuf_q_122(.A(q_in_122), .Y(P2_reg2[18]));
CLKBUFX1 gbuf_d_123(.A(n_31789), .Y(d_out_123));
CLKBUFX1 gbuf_q_123(.A(q_in_123), .Y(n_13355));
CLKBUFX1 gbuf_d_124(.A(n_31788), .Y(d_out_124));
CLKBUFX1 gbuf_q_124(.A(q_in_124), .Y(P3_reg1[18]));
CLKBUFX1 gbuf_d_125(.A(n_31787), .Y(d_out_125));
CLKBUFX1 gbuf_q_125(.A(q_in_125), .Y(n_13724));
CLKBUFX1 gbuf_d_126(.A(n_31786), .Y(d_out_126));
CLKBUFX1 gbuf_q_126(.A(q_in_126), .Y(n_10158));
CLKBUFX1 gbuf_d_127(.A(n_31724), .Y(d_out_127));
CLKBUFX1 gbuf_q_127(.A(q_in_127), .Y(P1_reg3[21]));
CLKBUFX1 gbuf_d_128(.A(n_31722), .Y(d_out_128));
CLKBUFX1 gbuf_q_128(.A(q_in_128), .Y(P1_reg3[23]));
CLKBUFX1 gbuf_d_129(.A(n_31725), .Y(d_out_129));
CLKBUFX1 gbuf_q_129(.A(q_in_129), .Y(P2_reg3[22]));
CLKBUFX1 gbuf_d_130(.A(n_31727), .Y(d_out_130));
CLKBUFX1 gbuf_q_130(.A(q_in_130), .Y(P1_reg3[22]));
CLKBUFX1 gbuf_d_131(.A(n_31761), .Y(d_out_131));
CLKBUFX1 gbuf_q_131(.A(q_in_131), .Y(n_9135));
CLKBUFX1 gbuf_d_132(.A(n_31759), .Y(d_out_132));
CLKBUFX1 gbuf_q_132(.A(q_in_132), .Y(n_10613));
CLKBUFX1 gbuf_d_133(.A(n_31758), .Y(d_out_133));
CLKBUFX1 gbuf_q_133(.A(q_in_133), .Y(n_10175));
CLKBUFX1 gbuf_d_134(.A(n_31756), .Y(d_out_134));
CLKBUFX1 gbuf_q_134(.A(q_in_134), .Y(n_10128));
CLKBUFX1 gbuf_d_135(.A(n_31760), .Y(d_out_135));
CLKBUFX1 gbuf_q_135(.A(q_in_135), .Y(P2_reg1[21]));
CLKBUFX1 gbuf_d_136(.A(n_31753), .Y(d_out_136));
CLKBUFX1 gbuf_q_136(.A(q_in_136), .Y(n_10223));
CLKBUFX1 gbuf_d_137(.A(n_31754), .Y(d_out_137));
CLKBUFX1 gbuf_q_137(.A(q_in_137), .Y(P1_reg1[19]));
CLKBUFX1 gbuf_d_138(.A(n_31762), .Y(d_out_138));
CLKBUFX1 gbuf_q_138(.A(q_in_138), .Y(P2_reg3[23]));
CLKBUFX1 gbuf_d_139(.A(n_31723), .Y(d_out_139));
CLKBUFX1 gbuf_qn_139(.A(qn_in_139), .Y(P3_reg_153));
CLKBUFX1 gbuf_d_140(.A(n_31747), .Y(d_out_140));
CLKBUFX1 gbuf_q_140(.A(q_in_140), .Y(P2_reg3[14]));
CLKBUFX1 gbuf_d_141(.A(n_31746), .Y(d_out_141));
CLKBUFX1 gbuf_q_141(.A(q_in_141), .Y(P2_reg3[15]));
CLKBUFX1 gbuf_d_142(.A(n_31769), .Y(d_out_142));
CLKBUFX1 gbuf_q_142(.A(q_in_142), .Y(P3_reg2[15]));
OAI21X1 g105422(.A0 (n_31650), .A1 (n_13197), .B0 (n_7254), .Y(n_31868));
NAND2X2 g105566(.A (n_35692), .B (n_35693), .Y (n_31867));
OAI21X1 g105570(.A0 (n_8103), .A1 (n_31713), .B0 (n_31772), .Y(n_35615));
NAND2X1 g105791(.A (n_31763), .B (n_12814), .Y (n_31865));
OAI21X1 g105583(.A0 (n_31616), .A1 (n_31273), .B0 (n_6680), .Y(n_31863));
OAI21X1 g105584(.A0 (n_31618), .A1 (n_31605), .B0 (n_6637), .Y(n_31862));
NAND2X1 g105586(.A (n_6626), .B (n_31784), .Y (n_31861));
OAI21X1 g105499(.A0 (n_31671), .A1 (n_31278), .B0 (n_6570), .Y(n_31860));
NAND2X1 g105856(.A (n_35696), .B (n_35697), .Y (n_31859));
NAND2X2 g105502(.A (n_35416), .B (n_35417), .Y (n_31858));
NAND2X1 g105859(.A (n_6936), .B (n_31773), .Y (n_31857));
OAI21X1 g105871(.A0 (n_31505), .A1 (n_30792), .B0 (n_6672), .Y(n_31856));
NAND2X1 g105879(.A (n_6616), .B (n_31695), .Y (n_31855));
NAND2X1 g105886(.A (n_7118), .B (n_31693), .Y (n_31854));
NAND2X2 g105887(.A (n_35137), .B (n_35138), .Y (n_31853));
NAND2X2 g105646(.A (n_31534), .B (n_35150), .Y (n_35075));
NAND2X1 g105649(.A (n_31850), .B (n_35706), .Y (n_31851));
OAI21X1 g105645(.A0 (n_31558), .A1 (n_8935), .B0 (n_31601), .Y(n_31849));
OAI21X1 g105653(.A0 (n_31566), .A1 (n_9942), .B0 (n_31588), .Y(n_31848));
OAI21X1 g105655(.A0 (n_31563), .A1 (n_10415), .B0 (n_31644), .Y(n_31847));
OAI21X1 g105656(.A0 (n_31576), .A1 (n_8892), .B0 (n_31845), .Y(n_31846));
NAND2X1 g105660(.A (n_31621), .B (n_31696), .Y (n_31844));
NAND2X2 g105664(.A (n_31640), .B (n_31850), .Y (n_32091));
NAND2X2 g105667(.A (n_35015), .B (n_31965), .Y (n_31841));
OAI21X1 g105668(.A0 (n_9867), .A1 (n_25823), .B0 (n_31632), .Y(n_31840));
OAI21X1 g105533(.A0 (n_9878), .A1 (n_31680), .B0 (n_31690), .Y(n_31838));
NAND2X1 g105684(.A (n_31610), .B (n_13005), .Y (n_31837));
NOR2X1 g105687(.A (n_10477), .B (n_31623), .Y (n_31836));
OAI21X1 g105535(.A0 (n_9854), .A1 (n_31834), .B0 (n_31691), .Y(n_31835));
OAI21X1 g105690(.A0 (n_31552), .A1 (n_30935), .B0 (n_8623), .Y(n_35899));
OAI21X1 g105701(.A0 (n_8238), .A1 (n_31881), .B0 (n_31629), .Y(n_35890));
OAI21X1 g105702(.A0 (n_8585), .A1 (n_31734), .B0 (n_31630), .Y(n_35618));
NAND2X1 g106025(.A (n_31617), .B (n_13014), .Y (n_31829));
OAI21X1 g105706(.A0 (n_34962), .A1 (n_31170), .B0 (n_30353), .Y(n_31827));
NAND2X1 g105707(.A (n_7098), .B (n_31648), .Y (n_31826));
NAND3X1 g105393(.A (n_32188), .B (n_2247), .C (n_32189), .Y(n_31825));
NAND2X1 g105715(.A (n_6730), .B (n_31645), .Y (n_31824));
OAI21X1 g106051(.A0 (n_31603), .A1 (n_31482), .B0 (n_8603), .Y(n_35932));
OAI21X1 g106054(.A0 (n_31600), .A1 (n_31410), .B0 (n_8602), .Y(n_31822));
NOR2X1 g105552(.A (n_7076), .B (n_31707), .Y (n_31821));
AOI22X1 g105553(.A0 (n_31513), .A1 (n_31878), .B0 (n_9260), .B1(n_31819), .Y (n_31820));
NAND2X1 g105471(.A (n_31681), .B (n_31922), .Y (n_35906));
NAND2X2 g106072(.A (n_35120), .B (n_35121), .Y (n_31817));
NAND2X1 g106073(.A (n_6888), .B (n_31642), .Y (n_31816));
NAND2X1 g106090(.A (n_6917), .B (n_31646), .Y (n_31815));
CLKBUFX1 gbuf_d_143(.A(n_31667), .Y(d_out_143));
CLKBUFX1 gbuf_qn_143(.A(qn_in_143), .Y(P2_reg_110));
CLKBUFX1 gbuf_d_144(.A(n_31664), .Y(d_out_144));
CLKBUFX1 gbuf_qn_144(.A(qn_in_144), .Y(P2_reg1[26]));
CLKBUFX1 gbuf_d_145(.A(n_31609), .Y(d_out_145));
CLKBUFX1 gbuf_q_145(.A(q_in_145), .Y(n_4475));
CLKBUFX1 gbuf_d_146(.A(n_31710), .Y(d_out_146));
CLKBUFX1 gbuf_q_146(.A(q_in_146), .Y(n_13357));
CLKBUFX1 gbuf_d_147(.A(n_31708), .Y(d_out_147));
CLKBUFX1 gbuf_q_147(.A(q_in_147), .Y(P3_reg2[18]));
CLKBUFX1 gbuf_d_148(.A(n_31619), .Y(d_out_148));
CLKBUFX1 gbuf_q_148(.A(q_in_148), .Y(P2_reg3[20]));
CLKBUFX1 gbuf_d_149(.A(n_31656), .Y(d_out_149));
CLKBUFX1 gbuf_q_149(.A(q_in_149), .Y(P2_reg_104));
CLKBUFX1 gbuf_d_150(.A(n_31655), .Y(d_out_150));
CLKBUFX1 gbuf_q_150(.A(q_in_150), .Y(P2_reg1[20]));
CLKBUFX1 gbuf_d_151(.A(n_31654), .Y(d_out_151));
CLKBUFX1 gbuf_q_151(.A(q_in_151), .Y(n_11148));
CLKBUFX1 gbuf_d_152(.A(n_31653), .Y(d_out_152));
CLKBUFX1 gbuf_q_152(.A(q_in_152), .Y(n_10047));
CLKBUFX1 gbuf_d_153(.A(n_31651), .Y(d_out_153));
CLKBUFX1 gbuf_q_153(.A(q_in_153), .Y(P1_reg_173));
CLKBUFX1 gbuf_d_154(.A(n_31652), .Y(d_out_154));
CLKBUFX1 gbuf_q_154(.A(q_in_154), .Y(P1_reg_172));
CLKBUFX1 gbuf_d_155(.A(n_31649), .Y(d_out_155));
CLKBUFX1 gbuf_q_155(.A(q_in_155), .Y(n_10136));
CLKBUFX1 gbuf_d_156(.A(n_31672), .Y(d_out_156));
CLKBUFX1 gbuf_q_156(.A(q_in_156), .Y(P2_reg3[13]));
CLKBUFX1 gbuf_d_157(.A(n_31673), .Y(d_out_157));
CLKBUFX1 gbuf_q_157(.A(q_in_157), .Y(P1_reg3[11]));
CLKBUFX1 gbuf_d_158(.A(n_31670), .Y(d_out_158));
CLKBUFX1 gbuf_q_158(.A(q_in_158), .Y(P3_reg3[11]));
CLKBUFX1 gbuf_d_159(.A(n_31614), .Y(d_out_159));
CLKBUFX1 gbuf_q_159(.A(q_in_159), .Y(P2_reg_107));
CLKBUFX1 gbuf_d_160(.A(n_31613), .Y(d_out_160));
CLKBUFX1 gbuf_q_160(.A(q_in_160), .Y(P2_reg1[23]));
CLKBUFX1 gbuf_d_161(.A(n_31611), .Y(d_out_161));
CLKBUFX1 gbuf_q_161(.A(q_in_161), .Y(n_10043));
CLKBUFX1 gbuf_d_162(.A(n_31637), .Y(d_out_162));
CLKBUFX1 gbuf_q_162(.A(q_in_162), .Y(P2_reg3[16]));
CLKBUFX1 gbuf_d_163(.A(n_31634), .Y(d_out_163));
CLKBUFX1 gbuf_q_163(.A(q_in_163), .Y(P3_reg3[15]));
CLKBUFX1 gbuf_d_164(.A(n_31688), .Y(d_out_164));
CLKBUFX1 gbuf_q_164(.A(q_in_164), .Y(P2_reg1[15]));
CLKBUFX1 gbuf_d_165(.A(n_31685), .Y(d_out_165));
CLKBUFX1 gbuf_q_165(.A(q_in_165), .Y(P2_reg2[15]));
CLKBUFX1 gbuf_d_166(.A(n_31687), .Y(d_out_166));
CLKBUFX1 gbuf_q_166(.A(q_in_166), .Y(n_4367));
CLKBUFX1 gbuf_d_167(.A(n_31676), .Y(d_out_167));
CLKBUFX1 gbuf_q_167(.A(q_in_167), .Y(n_9101));
OAI21X1 g105764(.A0 (n_31525), .A1 (n_10447), .B0 (n_31647), .Y(n_35880));
OAI21X1 g105766(.A0 (n_31524), .A1 (n_10432), .B0 (n_31528), .Y(n_31813));
NAND2X1 g105773(.A (n_31661), .B (n_31951), .Y (n_31812));
NAND2X1 g105577(.A (n_7125), .B (n_31705), .Y (n_31810));
NAND2X2 g105783(.A (n_31666), .B (n_31594), .Y (n_32056));
NAND2X1 g105786(.A (n_31660), .B (n_31933), .Y (n_35141));
NAND2X1 g105581(.A (n_6853), .B (n_31704), .Y (n_31806));
NAND2X1 g105790(.A (n_31657), .B (n_12806), .Y (n_31805));
NAND2X1 g105795(.A (n_31658), .B (n_13007), .Y (n_31804));
NAND2X2 g105588(.A (n_6534), .B (n_31703), .Y (n_31803));
NAND2X1 g105589(.A (n_7102), .B (n_31702), .Y (n_31802));
NOR2X1 g105819(.A (n_31225), .B (n_31668), .Y (n_31801));
AOI22X1 g105825(.A0 (n_31398), .A1 (n_35933), .B0 (n_8516), .B1(n_9387), .Y (n_31800));
OAI21X1 g105832(.A0 (n_31517), .A1 (n_12969), .B0 (n_6903), .Y(n_31799));
OAI21X1 g105842(.A0 (n_31979), .A1 (n_35931), .B0 (n_7364), .Y(n_31798));
NAND2X1 g105844(.A (n_6511), .B (n_31701), .Y (n_31797));
NAND2X1 g105847(.A (n_6683), .B (n_31678), .Y (n_31796));
NAND2X1 g105853(.A (n_7111), .B (n_31692), .Y (n_31795));
NAND2X2 g105854(.A (n_35281), .B (n_35282), .Y (n_31794));
NAND2X1 g105857(.A (n_32205), .B (n_32206), .Y (n_31793));
NAND2X1 g105866(.A (n_6937), .B (n_31700), .Y (n_31792));
NAND2X1 g105869(.A (n_6584), .B (n_31699), .Y (n_31791));
NAND2X1 g105870(.A (n_6599), .B (n_31697), .Y (n_31790));
OAI21X1 g105874(.A0 (n_31404), .A1 (n_31744), .B0 (n_6664), .Y(n_31789));
NAND2X1 g105876(.A (n_6593), .B (n_31582), .Y (n_31788));
NAND2X1 g105877(.A (n_6647), .B (n_31580), .Y (n_31787));
NAND2X1 g105885(.A (n_6882), .B (n_31578), .Y (n_31786));
NAND2X1 g105650(.A (n_31526), .B (n_31850), .Y (n_31785));
NAND2X1 g105659(.A (n_31506), .B (n_31783), .Y (n_31784));
NAND2X1 g105663(.A (n_31522), .B (n_31781), .Y (n_35692));
AOI21X1 g105669(.A0 (n_31489), .A1 (n_31243), .B0 (n_8070), .Y(n_31780));
OAI21X1 g105670(.A0 (n_31454), .A1 (n_31322), .B0 (n_33123), .Y(n_31779));
NAND3X1 g105673(.A (n_32920), .B (n_32921), .C (n_30439), .Y(n_31778));
NAND2X1 g105971(.A (n_31511), .B (n_31698), .Y (n_31777));
NAND2X1 g105973(.A (n_31510), .B (n_31260), .Y (n_31776));
NAND2X1 g105531(.A (n_31561), .B (n_31774), .Y (n_35416));
NAND2X1 g105977(.A (n_31507), .B (n_31933), .Y (n_31773));
OAI21X1 g105680(.A0 (n_34228), .A1 (n_31252), .B0 (n_31771), .Y(n_31772));
NAND2X1 g105994(.A (n_31508), .B (n_31933), .Y (n_35696));
NAND2X1 g106565(.A (n_6650), .B (n_31549), .Y (n_31769));
INVX1 g105688(.A (n_31679), .Y (n_31768));
OR4X1 g105696(.A (n_30600), .B (n_31223), .C (n_18926), .D (n_31314),.Y (n_31767));
NOR2X1 g106018(.A (n_31230), .B (n_31499), .Y (n_31766));
NOR2X1 g106036(.A (n_31315), .B (n_31509), .Y (n_31765));
OAI21X1 g105720(.A0 (n_9766), .A1 (n_31834), .B0 (n_31520), .Y(n_31764));
NOR2X1 g106064(.A (n_6902), .B (n_31533), .Y (n_31763));
NAND2X2 g106067(.A (n_35097), .B (n_35098), .Y (n_31762));
NAND2X1 g106069(.A (n_6652), .B (n_31531), .Y (n_31761));
NAND2X1 g106075(.A (n_6644), .B (n_31530), .Y (n_31760));
NAND2X1 g106077(.A (n_6662), .B (n_31529), .Y (n_31759));
OAI21X1 g106081(.A0 (n_31488), .A1 (n_31541), .B0 (n_6840), .Y(n_31758));
OAI21X1 g106082(.A0 (n_31487), .A1 (P1_n_449), .B0 (n_7175), .Y(n_31756));
NAND2X1 g106088(.A (n_6982), .B (n_31527), .Y (n_31754));
OAI21X1 g106089(.A0 (n_31486), .A1 (n_31541), .B0 (n_6914), .Y(n_31753));
CLKBUFX1 gbuf_d_168(.A(n_31539), .Y(d_out_168));
CLKBUFX1 gbuf_q_168(.A(q_in_168), .Y(n_13640));
CLKBUFX1 gbuf_d_169(.A(n_31583), .Y(d_out_169));
CLKBUFX1 gbuf_q_169(.A(q_in_169), .Y(P1_reg3[16]));
CLKBUFX1 gbuf_d_170(.A(n_31608), .Y(d_out_170));
CLKBUFX1 gbuf_q_170(.A(q_in_170), .Y(P3_reg1[17]));
CLKBUFX1 gbuf_d_171(.A(n_31606), .Y(d_out_171));
CLKBUFX1 gbuf_q_171(.A(q_in_171), .Y(n_13502));
CLKBUFX1 gbuf_d_172(.A(n_31514), .Y(d_out_172));
CLKBUFX1 gbuf_q_172(.A(q_in_172), .Y(P1_reg3[9]));
CLKBUFX1 gbuf_d_173(.A(n_31542), .Y(d_out_173));
CLKBUFX1 gbuf_q_173(.A(q_in_173), .Y(n_10178));
CLKBUFX1 gbuf_d_174(.A(n_31540), .Y(d_out_174));
CLKBUFX1 gbuf_q_174(.A(q_in_174), .Y(n_4477));
CLKBUFX1 gbuf_d_175(.A(n_31562), .Y(d_out_175));
CLKBUFX1 gbuf_q_175(.A(q_in_175), .Y(P1_reg3[13]));
CLKBUFX1 gbuf_d_176(.A(n_31560), .Y(d_out_176));
CLKBUFX1 gbuf_q_176(.A(q_in_176), .Y(P2_reg3[10]));
CLKBUFX1 gbuf_d_177(.A(n_31559), .Y(d_out_177));
CLKBUFX1 gbuf_q_177(.A(q_in_177), .Y(P2_reg3[12]));
CLKBUFX1 gbuf_d_178(.A(n_31554), .Y(d_out_178));
CLKBUFX1 gbuf_q_178(.A(q_in_178), .Y(P3_reg3[12]));
CLKBUFX1 gbuf_d_179(.A(n_31553), .Y(d_out_179));
CLKBUFX1 gbuf_q_179(.A(q_in_179), .Y(P3_reg3[14]));
CLKBUFX1 gbuf_d_180(.A(n_31503), .Y(d_out_180));
CLKBUFX1 gbuf_q_180(.A(q_in_180), .Y(P2_reg1[13]));
CLKBUFX1 gbuf_d_181(.A(n_31504), .Y(d_out_181));
CLKBUFX1 gbuf_q_181(.A(q_in_181), .Y(n_4160));
CLKBUFX1 gbuf_d_182(.A(n_31502), .Y(d_out_182));
CLKBUFX1 gbuf_qn_182(.A(qn_in_182), .Y(P3_reg_151));
CLKBUFX1 gbuf_d_183(.A(n_31501), .Y(d_out_183));
CLKBUFX1 gbuf_q_183(.A(q_in_183), .Y(n_13213));
CLKBUFX1 gbuf_d_184(.A(n_31500), .Y(d_out_184));
CLKBUFX1 gbuf_q_184(.A(q_in_184), .Y(n_13680));
CLKBUFX1 gbuf_d_185(.A(n_31498), .Y(d_out_185));
CLKBUFX1 gbuf_q_185(.A(q_in_185), .Y(P3_reg2[13]));
CLKBUFX1 gbuf_d_186(.A(n_31497), .Y(d_out_186));
CLKBUFX1 gbuf_q_186(.A(q_in_186), .Y(n_9103));
CLKBUFX1 gbuf_d_187(.A(n_31521), .Y(d_out_187));
CLKBUFX1 gbuf_q_187(.A(q_in_187), .Y(P1_reg3[14]));
OAI21X1 g105561(.A0 (n_31418), .A1 (n_31149), .B0 (n_7051), .Y(n_31752));
CLKBUFX1 gbuf_d_188(.A(n_31518), .Y(d_out_188));
CLKBUFX1 gbuf_q_188(.A(q_in_188), .Y(P3_reg3[8]));
CLKBUFX1 gbuf_d_189(.A(n_31575), .Y(d_out_189));
CLKBUFX1 gbuf_q_189(.A(q_in_189), .Y(P1_reg2[14]));
CLKBUFX1 gbuf_d_190(.A(n_31572), .Y(d_out_190));
CLKBUFX1 gbuf_q_190(.A(q_in_190), .Y(P2_reg2[16]));
CLKBUFX1 gbuf_d_191(.A(n_31568), .Y(d_out_191));
CLKBUFX1 gbuf_q_191(.A(q_in_191), .Y(P3_reg1[15]));
CLKBUFX1 gbuf_d_192(.A(n_31570), .Y(d_out_192));
CLKBUFX1 gbuf_q_192(.A(q_in_192), .Y(n_13365));
CLKBUFX1 gbuf_d_193(.A(n_31532), .Y(d_out_193));
CLKBUFX1 gbuf_q_193(.A(q_in_193), .Y(n_9773));
OAI21X1 g105777(.A0 (n_9880), .A1 (n_31639), .B0 (n_31556), .Y(n_31748));
NAND2X1 g106172(.A (n_31579), .B (n_12888), .Y (n_31747));
NAND2X1 g106173(.A (n_31581), .B (n_12879), .Y (n_31746));
OAI21X1 g105585(.A0 (n_31401), .A1 (n_31744), .B0 (n_6755), .Y(n_31745));
OAI21X1 g105804(.A0 (n_8275), .A1 (n_29486), .B0 (n_31577), .Y(n_31742));
OAI21X1 g105806(.A0 (n_9795), .A1 (n_31740), .B0 (n_31545), .Y(n_31741));
OAI21X1 g105808(.A0 (n_8819), .A1 (n_31422), .B0 (n_31543), .Y(n_31738));
NOR2X1 g105812(.A (n_7084), .B (n_31587), .Y (n_31736));
OAI21X1 g105815(.A0 (n_8562), .A1 (n_31734), .B0 (n_31574), .Y(n_31735));
NOR2X1 g105818(.A (n_31229), .B (n_33086), .Y (n_31733));
NOR2X1 g105821(.A (n_6765), .B (n_31596), .Y (n_31732));
AOI22X1 g105827(.A0 (n_31428), .A1 (n_31878), .B0 (n_9335), .B1(n_6891), .Y (n_31731));
OAI21X1 g105829(.A0 (n_33655), .A1 (n_30650), .B0 (n_31628), .Y(n_31730));
OAI21X1 g105830(.A0 (n_31419), .A1 (n_30988), .B0 (n_31544), .Y(n_31729));
NOR2X1 g105831(.A (n_7016), .B (n_31604), .Y (n_31728));
OAI21X1 g105836(.A0 (n_31399), .A1 (n_31726), .B0 (n_7246), .Y(n_31727));
NAND2X1 g105837(.A (n_7094), .B (n_31599), .Y (n_31725));
NAND2X1 g105838(.A (n_7237), .B (n_31602), .Y (n_31724));
NAND2X1 g106284(.A (n_6634), .B (n_31607), .Y (n_31723));
NAND2X1 g105839(.A (n_35923), .B (n_35924), .Y (n_31722));
NAND2X1 g105845(.A (n_6491), .B (n_31591), .Y (n_31720));
NAND2X2 g105846(.A (n_35139), .B (n_35140), .Y (n_31719));
NAND2X1 g105849(.A (n_6681), .B (n_31595), .Y (n_31718));
NAND2X1 g105855(.A (n_6575), .B (n_31567), .Y (n_31717));
NAND2X1 g105858(.A (n_6926), .B (n_31593), .Y (n_31716));
NAND2X1 g105862(.A (n_6735), .B (n_31589), .Y (n_31715));
OAI21X1 g105864(.A0 (n_8234), .A1 (n_31713), .B0 (n_31557), .Y(n_31714));
NAND2X1 g105867(.A (n_6869), .B (n_31585), .Y (n_31712));
NAND2X1 g105868(.A (n_6564), .B (n_31584), .Y (n_31711));
OAI21X1 g105872(.A0 (n_31293), .A1 (n_31273), .B0 (n_6510), .Y(n_31710));
OAI21X1 g105883(.A0 (n_31292), .A1 (n_31744), .B0 (n_6707), .Y(n_31708));
AOI21X1 g105648(.A0 (n_10456), .A1 (n_31338), .B0 (n_31490), .Y(n_31707));
OR4X1 g105651(.A (n_30051), .B (n_30042), .C (n_10589), .D (n_33998),.Y (n_31706));
OAI21X1 g105654(.A0 (n_31361), .A1 (n_8889), .B0 (n_31592), .Y(n_31705));
OAI21X1 g105657(.A0 (n_31357), .A1 (n_8894), .B0 (n_31845), .Y(n_31704));
NAND2X1 g105661(.A (n_31406), .B (n_31783), .Y (n_31703));
OAI21X1 g105665(.A0 (n_31354), .A1 (n_8917), .B0 (n_31845), .Y(n_31702));
NAND2X1 g105958(.A (n_31435), .B (n_31590), .Y (n_31701));
NAND2X1 g105963(.A (n_31415), .B (n_31912), .Y (n_31700));
NAND2X1 g105966(.A (n_31413), .B (n_31698), .Y (n_31699));
NAND2X1 g105967(.A (n_31412), .B (n_31696), .Y (n_31697));
NAND2X1 g105972(.A (n_31407), .B (n_31694), .Y (n_31695));
NAND2X1 g105975(.A (n_31411), .B (n_31205), .Y (n_31693));
NAND2X1 g105980(.A (n_31405), .B (n_31933), .Y (n_31692));
OAI21X1 g105681(.A0 (n_31350), .A1 (n_30770), .B0 (n_31689), .Y(n_31691));
OAI21X1 g105682(.A0 (n_31336), .A1 (n_30769), .B0 (n_31689), .Y(n_31690));
NAND2X1 g106550(.A (n_32874), .B (n_32875), .Y (n_31688));
OAI21X1 g106553(.A0 (n_31295), .A1 (n_33201), .B0 (n_6592), .Y(n_31687));
NAND2X1 g106554(.A (n_6613), .B (n_31462), .Y (n_31685));
NAND2X1 g105990(.A (n_31423), .B (n_31683), .Y (n_35281));
NAND2X1 g105992(.A (n_31408), .B (n_31677), .Y (n_35137));
OAI21X1 g105534(.A0 (n_9847), .A1 (n_31680), .B0 (n_31474), .Y(n_31681));
NAND4X1 g105689(.A (n_30987), .B (n_30356), .C (n_31189), .D(n_30767), .Y (n_31679));
NAND2X1 g105997(.A (n_31424), .B (n_31677), .Y (n_31678));
NAND2X1 g106570(.A (n_6643), .B (n_31460), .Y (n_31676));
NAND2X1 g106001(.A (n_31677), .B (n_35293), .Y (n_32205));
NAND2X1 g106005(.A (n_31417), .B (n_12723), .Y (n_31673));
NAND2X1 g106010(.A (n_31416), .B (n_12881), .Y (n_31672));
NOR2X1 g105698(.A (n_10393), .B (n_31431), .Y (n_31671));
NAND2X1 g106023(.A (n_31400), .B (n_13016), .Y (n_31670));
OR4X1 g106028(.A (n_30141), .B (n_30955), .C (n_18927), .D (n_31181),.Y (n_31669));
NAND2X1 g106039(.A (n_31432), .B (n_31133), .Y (n_31668));
NAND2X1 g105710(.A (n_6696), .B (n_31439), .Y (n_31667));
OAI21X1 g106041(.A0 (n_9752), .A1 (n_31129), .B0 (n_31403), .Y(n_31666));
NAND2X1 g105713(.A (n_6731), .B (n_31436), .Y (n_31664));
OAI21X1 g106055(.A0 (n_31368), .A1 (n_31620), .B0 (n_10379), .Y(n_31661));
OAI21X1 g106058(.A0 (n_8586), .A1 (n_30527), .B0 (n_31426), .Y(n_31660));
NOR2X1 g106061(.A (n_9898), .B (n_31434), .Y (n_31659));
NOR2X1 g106062(.A (n_7026), .B (n_31444), .Y (n_31658));
NOR2X1 g106063(.A (n_6894), .B (n_31443), .Y (n_31657));
NAND2X1 g106068(.A (n_6551), .B (n_31441), .Y (n_31656));
NAND2X1 g106074(.A (n_32159), .B (n_32160), .Y (n_31655));
CLKBUFX1 gbuf_d_194(.A(n_31457), .Y(d_out_194));
CLKBUFX1 gbuf_q_194(.A(q_in_194), .Y(P3_reg3[9]));
NAND2X1 g106076(.A (n_35131), .B (n_35132), .Y (n_31654));
NAND2X1 g106079(.A (n_6532), .B (n_31437), .Y (n_31653));
OAI21X1 g106083(.A0 (n_31371), .A1 (n_31472), .B0 (n_6847), .Y(n_31652));
OAI21X1 g106084(.A0 (n_31370), .A1 (n_31470), .B0 (n_7126), .Y(n_31651));
AOI22X1 g105558(.A0 (n_31306), .A1 (n_31878), .B0 (n_9236), .B1(n_31876), .Y (n_31650));
NAND2X1 g106091(.A (n_35329), .B (n_35330), .Y (n_31649));
CLKBUFX1 gbuf_d_195(.A(n_31452), .Y(d_out_195));
CLKBUFX1 gbuf_q_195(.A(q_in_195), .Y(n_13322));
CLKBUFX1 gbuf_d_196(.A(n_31455), .Y(d_out_196));
CLKBUFX1 gbuf_q_196(.A(q_in_196), .Y(n_13893));
CLKBUFX1 gbuf_d_197(.A(n_31449), .Y(d_out_197));
CLKBUFX1 gbuf_q_197(.A(q_in_197), .Y(n_13635));
CLKBUFX1 gbuf_d_198(.A(n_31391), .Y(d_out_198));
CLKBUFX1 gbuf_q_198(.A(q_in_198), .Y(P1_reg2[16]));
CLKBUFX1 gbuf_d_199(.A(n_31390), .Y(d_out_199));
CLKBUFX1 gbuf_q_199(.A(q_in_199), .Y(n_10180));
CLKBUFX1 gbuf_d_200(.A(n_31492), .Y(d_out_200));
CLKBUFX1 gbuf_q_200(.A(q_in_200), .Y(P1_reg1[16]));
CLKBUFX1 gbuf_d_201(.A(n_31447), .Y(d_out_201));
CLKBUFX1 gbuf_q_201(.A(q_in_201), .Y(n_4011));
CLKBUFX1 gbuf_d_202(.A(n_31446), .Y(d_out_202));
CLKBUFX1 gbuf_q_202(.A(q_in_202), .Y(P1_reg2[9]));
CLKBUFX1 gbuf_d_203(.A(n_31445), .Y(d_out_203));
CLKBUFX1 gbuf_q_203(.A(q_in_203), .Y(n_10154));
CLKBUFX1 gbuf_d_204(.A(n_31463), .Y(d_out_204));
CLKBUFX1 gbuf_q_204(.A(q_in_204), .Y(P1_reg3[15]));
CLKBUFX1 gbuf_d_205(.A(n_31459), .Y(d_out_205));
CLKBUFX1 gbuf_q_205(.A(q_in_205), .Y(n_1319));
CLKBUFX1 gbuf_d_206(.A(n_31397), .Y(d_out_206));
CLKBUFX1 gbuf_q_206(.A(q_in_206), .Y(P2_reg1[10]));
CLKBUFX1 gbuf_d_207(.A(n_31396), .Y(d_out_207));
CLKBUFX1 gbuf_q_207(.A(q_in_207), .Y(n_13377));
CLKBUFX1 gbuf_d_208(.A(n_31395), .Y(d_out_208));
CLKBUFX1 gbuf_q_208(.A(q_in_208), .Y(P3_reg1[16]));
CLKBUFX1 gbuf_d_209(.A(n_31394), .Y(d_out_209));
CLKBUFX1 gbuf_q_209(.A(q_in_209), .Y(n_13342));
CLKBUFX1 gbuf_d_210(.A(n_31393), .Y(d_out_210));
CLKBUFX1 gbuf_q_210(.A(q_in_210), .Y(n_13507));
CLKBUFX1 gbuf_d_211(.A(n_31392), .Y(d_out_211));
CLKBUFX1 gbuf_q_211(.A(q_in_211), .Y(n_9067));
CLKBUFX1 gbuf_d_212(.A(n_31430), .Y(d_out_212));
CLKBUFX1 gbuf_q_212(.A(q_in_212), .Y(P2_reg3[11]));
CLKBUFX1 gbuf_d_213(.A(n_31473), .Y(d_out_213));
CLKBUFX1 gbuf_q_213(.A(q_in_213), .Y(n_10201));
CLKBUFX1 gbuf_d_214(.A(n_31471), .Y(d_out_214));
CLKBUFX1 gbuf_q_214(.A(q_in_214), .Y(n_10189));
CLKBUFX1 gbuf_d_215(.A(n_31467), .Y(d_out_215));
CLKBUFX1 gbuf_q_215(.A(q_in_215), .Y(n_4534));
CLKBUFX1 gbuf_d_216(.A(n_31466), .Y(d_out_216));
CLKBUFX1 gbuf_q_216(.A(q_in_216), .Y(P1_reg1[14]));
OAI21X1 g105761(.A0 (n_31311), .A1 (n_9963), .B0 (n_31647), .Y(n_31648));
NAND2X1 g106141(.A (n_31483), .B (n_31891), .Y (n_31646));
OAI21X1 g105769(.A0 (n_31318), .A1 (n_9900), .B0 (n_31644), .Y(n_31645));
NAND2X1 g106155(.A (n_31481), .B (n_31641), .Y (n_35120));
NAND2X1 g106156(.A (n_31479), .B (n_31641), .Y (n_31642));
OAI21X1 g105779(.A0 (n_9855), .A1 (n_31639), .B0 (n_31458), .Y(n_31640));
OAI21X1 g105780(.A0 (n_31326), .A1 (n_31244), .B0 (n_31573), .Y(n_31638));
NAND2X2 g106174(.A (n_31477), .B (n_12886), .Y (n_31637));
OR4X1 g105787(.A (n_30586), .B (n_9039), .C (n_30998), .D (n_31226),.Y (n_31636));
NAND2X1 g106184(.A (n_31485), .B (n_13009), .Y (n_31634));
OAI21X1 g105794(.A0 (n_31320), .A1 (n_30734), .B0 (n_31555), .Y(n_31632));
OR4X1 g105797(.A (n_30261), .B (n_30813), .C (n_20748), .D (n_31256),.Y (n_31631));
OAI21X1 g105800(.A0 (n_33133), .A1 (n_31253), .B0 (n_30403), .Y(n_31630));
OAI21X1 g105801(.A0 (n_31305), .A1 (n_31046), .B0 (n_31628), .Y(n_31629));
NAND4X1 g105805(.A (n_32132), .B (n_30440), .C (n_32133), .D(n_26973), .Y (n_35879));
AOI21X1 g105813(.A0 (n_31303), .A1 (n_30816), .B0 (n_31564), .Y(n_31623));
NOR2X1 g105814(.A (n_31451), .B (n_30993), .Y (n_31622));
OAI21X1 g105816(.A0 (n_31297), .A1 (n_31620), .B0 (n_10429), .Y(n_31621));
NAND2X1 g105822(.A (n_7096), .B (n_31478), .Y (n_31619));
NOR2X1 g105823(.A (n_9899), .B (n_31475), .Y (n_31618));
NOR2X1 g106257(.A (n_7069), .B (n_31389), .Y (n_31617));
NOR2X1 g105826(.A (n_10370), .B (n_31469), .Y (n_31616));
OAI21X1 g105828(.A0 (n_9765), .A1 (n_24484), .B0 (n_31450), .Y(n_35706));
OAI21X1 g106265(.A0 (n_31333), .A1 (n_29285), .B0 (n_6701), .Y(n_31614));
OAI21X1 g106273(.A0 (n_31331), .A1 (n_33201), .B0 (n_6604), .Y(n_31613));
OAI21X1 g105834(.A0 (n_9154), .A1 (n_31122), .B0 (n_34784), .Y(n_35150));
NAND2X2 g106278(.A (n_35103), .B (n_35104), .Y (n_31611));
NOR2X1 g105840(.A (n_7059), .B (n_31491), .Y (n_31610));
OAI21X1 g105843(.A0 (n_31324), .A1 (n_31328), .B0 (n_6646), .Y(n_31609));
OAI21X1 g105875(.A0 (n_31135), .A1 (n_31273), .B0 (n_6514), .Y(n_31608));
NAND2X1 g106364(.A (n_31330), .B (n_31698), .Y (n_31607));
OAI21X1 g105882(.A0 (n_31128), .A1 (n_31605), .B0 (n_6565), .Y(n_31606));
CLKBUFX1 gbuf_d_217(.A(n_31277), .Y(d_out_217));
CLKBUFX1 gbuf_q_217(.A(q_in_217), .Y(n_13679));
AOI21X1 g105941(.A0 (n_9426), .A1 (n_31242), .B0 (n_34676), .Y(n_31604));
NOR2X1 g106475(.A (n_31056), .B (n_31335), .Y (n_31603));
OAI21X1 g105942(.A0 (n_31234), .A1 (n_8934), .B0 (n_31601), .Y(n_31602));
NOR2X1 g106477(.A (n_31055), .B (n_31334), .Y (n_31600));
OAI21X1 g105943(.A0 (n_31203), .A1 (n_9964), .B0 (n_31644), .Y(n_31599));
NAND2X1 g105944(.A (n_31287), .B (n_35023), .Y (n_35923));
AOI21X1 g105948(.A0 (n_10403), .A1 (n_31209), .B0 (n_31586), .Y(n_31596));
NAND2X1 g105951(.A (n_31309), .B (n_31594), .Y (n_31595));
OAI21X1 g105954(.A0 (n_31255), .A1 (n_8714), .B0 (n_31592), .Y(n_31593));
NAND2X1 g105957(.A (n_31323), .B (n_31590), .Y (n_31591));
OAI21X1 g105959(.A0 (n_31237), .A1 (n_9917), .B0 (n_31588), .Y(n_31589));
AOI21X1 g105961(.A0 (n_10401), .A1 (n_31208), .B0 (n_31586), .Y(n_31587));
OAI21X1 g105964(.A0 (n_31250), .A1 (n_8896), .B0 (n_31592), .Y(n_31585));
NAND2X1 g105965(.A (n_31301), .B (n_31951), .Y (n_31584));
NAND2X1 g105675(.A (n_31283), .B (n_12812), .Y (n_31583));
NAND2X1 g105969(.A (n_31300), .B (n_31781), .Y (n_31582));
NOR2X1 g106525(.A (n_6792), .B (n_31344), .Y (n_31581));
NAND2X1 g105970(.A (n_31298), .B (n_31698), .Y (n_31580));
CLKBUFX1 gbuf_d_218(.A(n_31271), .Y(d_out_218));
CLKBUFX1 gbuf_q_218(.A(q_in_218), .Y(n_4920));
NOR2X1 g106534(.A (n_7085), .B (n_31347), .Y (n_31579));
OAI21X1 g105976(.A0 (n_31247), .A1 (n_8911), .B0 (n_31592), .Y(n_31578));
OAI21X1 g105981(.A0 (n_31112), .A1 (n_33512), .B0 (n_31628), .Y(n_31577));
AOI21X1 g105983(.A0 (n_31264), .A1 (n_30827), .B0 (n_31360), .Y(n_31576));
NAND2X2 g106548(.A (n_32283), .B (n_32284), .Y (n_31575));
OAI21X1 g105985(.A0 (n_31267), .A1 (n_33501), .B0 (n_31573), .Y(n_31574));
NAND2X1 g106555(.A (n_6499), .B (n_31346), .Y (n_31572));
NAND2X2 g105989(.A (n_31310), .B (n_31590), .Y (n_35139));
OAI21X1 g106560(.A0 (n_31119), .A1 (n_31569), .B0 (n_6697), .Y(n_31570));
OAI21X1 g106562(.A0 (n_31118), .A1 (n_31569), .B0 (n_6615), .Y(n_31568));
NAND2X1 g105991(.A (n_31683), .B (n_35610), .Y (n_31567));
AOI21X1 g105999(.A0 (n_31265), .A1 (n_30829), .B0 (n_31523), .Y(n_31566));
AOI21X1 g106003(.A0 (n_31220), .A1 (n_30828), .B0 (n_31236), .Y(n_31563));
NAND2X1 g106006(.A (n_31304), .B (n_12718), .Y (n_31562));
OAI21X1 g105694(.A0 (n_31159), .A1 (n_8505), .B0 (n_10367), .Y(n_31561));
NAND2X1 g106008(.A (n_31291), .B (n_12896), .Y (n_31560));
NAND2X1 g106009(.A (n_31294), .B (n_12873), .Y (n_31559));
AOI21X1 g106012(.A0 (n_31232), .A1 (n_30815), .B0 (n_31233), .Y(n_31558));
OAI21X1 g106013(.A0 (n_33548), .A1 (n_31047), .B0 (n_31771), .Y(n_31557));
OAI21X1 g106019(.A0 (n_31239), .A1 (n_30420), .B0 (n_31555), .Y(n_31556));
NAND2X1 g106024(.A (n_31296), .B (n_13023), .Y (n_31554));
NAND2X1 g106026(.A (n_31290), .B (n_13012), .Y (n_31553));
NOR2X1 g106033(.A (n_31327), .B (n_31313), .Y (n_31552));
NAND2X1 g106668(.A (n_31289), .B (n_31694), .Y (n_31549));
CLKBUFX1 gbuf_d_219(.A(n_31285), .Y(d_out_219));
CLKBUFX1 gbuf_q_219(.A(q_in_219), .Y(n_9121));
NOR2X1 g106049(.A (n_31302), .B (n_29973), .Y (n_31548));
OAI21X1 g106065(.A0 (n_31214), .A1 (n_30324), .B0 (n_31544), .Y(n_31545));
OAI21X1 g106066(.A0 (n_31212), .A1 (n_30314), .B0 (n_30914), .Y(n_31543));
OAI21X1 g106080(.A0 (n_31207), .A1 (n_31541), .B0 (n_6922), .Y(n_31542));
OAI21X1 g106087(.A0 (n_31204), .A1 (n_31538), .B0 (n_6994), .Y(n_31540));
OAI21X1 g105559(.A0 (n_31146), .A1 (n_31538), .B0 (n_6929), .Y(n_31539));
CLKBUFX1 gbuf_d_220(.A(n_31366), .Y(d_out_220));
CLKBUFX1 gbuf_q_220(.A(q_in_220), .Y(P1_reg3[12]));
CLKBUFX1 gbuf_d_221(.A(n_31272), .Y(d_out_221));
CLKBUFX1 gbuf_q_221(.A(q_in_221), .Y(P1_reg1[30]));
CLKBUFX1 gbuf_d_222(.A(n_31270), .Y(d_out_222));
CLKBUFX1 gbuf_q_222(.A(q_in_222), .Y(n_14133));
CLKBUFX1 gbuf_d_223(.A(n_31268), .Y(d_out_223));
CLKBUFX1 gbuf_q_223(.A(q_in_223), .Y(P1_reg2[30]));
CLKBUFX1 gbuf_d_224(.A(n_31269), .Y(d_out_224));
CLKBUFX1 gbuf_q_224(.A(q_in_224), .Y(P2_reg1[31]));
CLKBUFX1 gbuf_d_225(.A(n_31387), .Y(d_out_225));
CLKBUFX1 gbuf_q_225(.A(q_in_225), .Y(P1_reg_180));
CLKBUFX1 gbuf_d_226(.A(n_31340), .Y(d_out_226));
CLKBUFX1 gbuf_q_226(.A(q_in_226), .Y(P3_reg3[10]));
CLKBUFX1 gbuf_d_227(.A(n_31286), .Y(d_out_227));
CLKBUFX1 gbuf_q_227(.A(q_in_227), .Y(n_4213));
CLKBUFX1 gbuf_d_228(.A(n_31284), .Y(d_out_228));
CLKBUFX1 gbuf_q_228(.A(q_in_228), .Y(P2_reg1[9]));
CLKBUFX1 gbuf_d_229(.A(n_31288), .Y(d_out_229));
CLKBUFX1 gbuf_q_229(.A(q_in_229), .Y(P2_reg2[9]));
CLKBUFX1 gbuf_d_230(.A(n_31282), .Y(d_out_230));
CLKBUFX1 gbuf_q_230(.A(q_in_230), .Y(n_10182));
CLKBUFX1 gbuf_d_231(.A(n_31281), .Y(d_out_231));
CLKBUFX1 gbuf_qn_231(.A(qn_in_231), .Y(P3_reg_152));
CLKBUFX1 gbuf_d_232(.A(n_31279), .Y(d_out_232));
CLKBUFX1 gbuf_q_232(.A(q_in_232), .Y(P3_reg1[11]));
CLKBUFX1 gbuf_d_233(.A(n_31280), .Y(d_out_233));
CLKBUFX1 gbuf_qn_233(.A(qn_in_233), .Y(P3_reg_149));
CLKBUFX1 gbuf_d_234(.A(n_31274), .Y(d_out_234));
CLKBUFX1 gbuf_q_234(.A(q_in_234), .Y(n_13338));
CLKBUFX1 gbuf_d_235(.A(n_31276), .Y(d_out_235));
CLKBUFX1 gbuf_q_235(.A(q_in_235), .Y(n_13366));
CLKBUFX1 gbuf_d_236(.A(n_31316), .Y(d_out_236));
CLKBUFX1 gbuf_q_236(.A(q_in_236), .Y(P1_reg3[10]));
CLKBUFX1 gbuf_d_237(.A(n_31359), .Y(d_out_237));
CLKBUFX1 gbuf_q_237(.A(q_in_237), .Y(n_4151));
CLKBUFX1 gbuf_d_238(.A(n_31358), .Y(d_out_238));
CLKBUFX1 gbuf_q_238(.A(q_in_238), .Y(n_4590));
CLKBUFX1 gbuf_d_239(.A(n_31356), .Y(d_out_239));
CLKBUFX1 gbuf_q_239(.A(q_in_239), .Y(P2_reg1[16]));
CLKBUFX1 gbuf_d_240(.A(n_31353), .Y(d_out_240));
CLKBUFX1 gbuf_q_240(.A(q_in_240), .Y(n_10191));
CLKBUFX1 gbuf_d_241(.A(n_31352), .Y(d_out_241));
CLKBUFX1 gbuf_q_241(.A(q_in_241), .Y(n_3958));
CLKBUFX1 gbuf_d_242(.A(n_31348), .Y(d_out_242));
CLKBUFX1 gbuf_q_242(.A(q_in_242), .Y(n_9565));
CLKBUFX1 gbuf_d_243(.A(n_31349), .Y(d_out_243));
CLKBUFX1 gbuf_q_243(.A(q_in_243), .Y(n_9071));
CLKBUFX1 gbuf_d_244(.A(n_31376), .Y(d_out_244));
CLKBUFX1 gbuf_q_244(.A(q_in_244), .Y(P1_reg3[6]));
CLKBUFX1 gbuf_d_245(.A(n_31375), .Y(d_out_245));
CLKBUFX1 gbuf_q_245(.A(q_in_245), .Y(P1_reg3[7]));
CLKBUFX1 gbuf_d_246(.A(n_31329), .Y(d_out_246));
CLKBUFX1 gbuf_q_246(.A(q_in_246), .Y(n_9586));
NAND3X1 g105478(.A (n_35669), .B (n_27232), .C (n_31536), .Y(n_32188));
NAND2X1 g106129(.A (n_31534), .B (n_35900), .Y (n_35097));
AOI21X1 g106132(.A0 (n_9388), .A1 (n_31175), .B0 (n_30702), .Y(n_31533));
NAND2X1 g106828(.A (n_6540), .B (n_31321), .Y (n_31532));
OAI21X1 g106136(.A0 (n_31173), .A1 (n_9947), .B0 (n_31588), .Y(n_31531));
OAI21X1 g106138(.A0 (n_31171), .A1 (n_10433), .B0 (n_31588), .Y(n_31530));
OAI21X1 g106139(.A0 (n_31169), .A1 (n_9920), .B0 (n_31528), .Y(n_31529));
OAI21X1 g106140(.A0 (n_9378), .A1 (n_31176), .B0 (n_31845), .Y(n_31527));
OAI21X1 g105774(.A0 (n_9857), .A1 (n_31834), .B0 (n_31339), .Y(n_31526));
AOI21X1 g106161(.A0 (n_31184), .A1 (n_30787), .B0 (n_8377), .Y(n_31525));
AOI21X1 g106164(.A0 (n_31183), .A1 (n_30786), .B0 (n_31523), .Y(n_31524));
OAI21X1 g105778(.A0 (n_9858), .A1 (n_31639), .B0 (n_31341), .Y(n_31522));
NAND2X1 g106170(.A (n_31362), .B (n_12716), .Y (n_31521));
OAI21X1 g105782(.A0 (n_31139), .A1 (n_30161), .B0 (n_33123), .Y(n_31520));
NAND2X1 g106185(.A (n_31365), .B (n_12997), .Y (n_31518));
AOI22X1 g106189(.A0 (n_31168), .A1 (n_35008), .B0 (n_9347), .B1(n_34706), .Y (n_31517));
NAND2X1 g105793(.A (n_31332), .B (n_12728), .Y (n_31514));
OR4X1 g105796(.A (n_30251), .B (n_30653), .C (n_18929), .D (n_31104),.Y (n_31513));
OAI21X1 g106236(.A0 (n_31156), .A1 (n_31936), .B0 (n_10357), .Y(n_31511));
OAI21X1 g106238(.A0 (n_31155), .A1 (n_31936), .B0 (n_10445), .Y(n_31510));
NAND2X1 g106239(.A (n_31383), .B (n_31369), .Y (n_31509));
OAI21X1 g106242(.A0 (n_8591), .A1 (n_31414), .B0 (n_31372), .Y(n_31508));
OAI21X1 g106243(.A0 (n_8588), .A1 (n_31480), .B0 (n_31382), .Y(n_31507));
OAI21X1 g105820(.A0 (n_31134), .A1 (n_31620), .B0 (n_10372), .Y(n_31506));
NOR2X1 g106245(.A (n_9897), .B (n_31381), .Y (n_31505));
NAND2X1 g106261(.A (n_6726), .B (n_31386), .Y (n_31504));
NAND2X1 g106272(.A (n_6689), .B (n_31379), .Y (n_31503));
NAND2X1 g106282(.A (n_6706), .B (n_31385), .Y (n_31502));
NAND2X1 g106285(.A (n_6600), .B (n_31384), .Y (n_31501));
OAI21X1 g106291(.A0 (n_31157), .A1 (n_31275), .B0 (n_6583), .Y(n_31500));
NAND2X1 g106294(.A (n_31374), .B (n_31367), .Y (n_31499));
OAI21X1 g106299(.A0 (n_31154), .A1 (n_31605), .B0 (n_6504), .Y(n_31498));
NAND2X1 g106305(.A (n_35262), .B (n_35263), .Y (n_31497));
AOI22X1 g106306(.A0 (n_31165), .A1 (n_31878), .B0 (n_9272), .B1(n_31495), .Y (n_35931));
CLKBUFX1 gbuf_d_247(.A(n_31351), .Y(d_out_247));
CLKBUFX1 gbuf_q_247(.A(q_in_247), .Y(n_4215));
NAND2X1 g106372(.A (n_31158), .B (n_31493), .Y (n_35103));
NAND2X1 g105884(.A (n_6906), .B (n_31196), .Y (n_31492));
AOI21X1 g105945(.A0 (n_10491), .A1 (n_31100), .B0 (n_31490), .Y(n_31491));
NOR3X1 g105949(.A (n_30720), .B (n_26455), .C (n_31070), .Y(n_31489));
NOR2X1 g106496(.A (n_9380), .B (n_31180), .Y (n_31488));
NOR2X1 g106497(.A (n_8897), .B (n_31179), .Y (n_31487));
NOR2X1 g106509(.A (n_8912), .B (n_31177), .Y (n_31486));
NOR2X1 g106510(.A (n_7021), .B (n_31167), .Y (n_31485));
OAI21X1 g106512(.A0 (n_30983), .A1 (n_31482), .B0 (n_9887), .Y(n_31483));
OAI21X1 g106521(.A0 (n_8263), .A1 (n_31480), .B0 (n_31162), .Y(n_31481));
OAI21X1 g106522(.A0 (n_8599), .A1 (n_31199), .B0 (n_31161), .Y(n_31479));
NAND2X1 g105978(.A (n_31137), .B (n_31534), .Y (n_31478));
AOI22X1 g106540(.A0 (n_30975), .A1 (n_31528), .B0 (n_3647), .B1(n_35007), .Y (n_31477));
AOI21X1 g105986(.A0 (n_31083), .A1 (n_30903), .B0 (n_33125), .Y(n_31475));
OAI21X1 g105683(.A0 (n_31034), .A1 (n_30263), .B0 (n_31555), .Y(n_31474));
OAI21X1 g106557(.A0 (n_30981), .A1 (n_31472), .B0 (n_7113), .Y(n_31473));
OAI21X1 g106559(.A0 (n_30980), .A1 (n_31470), .B0 (n_7116), .Y(n_31471));
AOI21X1 g105993(.A0 (n_31084), .A1 (n_30870), .B0 (n_33125), .Y(n_31469));
NAND2X1 g106566(.A (n_7115), .B (n_31182), .Y (n_31467));
OAI21X1 g106568(.A0 (n_30977), .A1 (P1_n_449), .B0 (n_6918), .Y(n_31466));
NAND2X1 g106595(.A (n_31132), .B (n_31683), .Y (n_32874));
NAND2X1 g106007(.A (n_31125), .B (n_12818), .Y (n_31463));
NAND2X1 g106597(.A (n_31130), .B (n_31097), .Y (n_31462));
NAND2X1 g106606(.A (n_31123), .B (n_31677), .Y (n_31460));
NAND2X1 g106014(.A (n_31127), .B (n_12871), .Y (n_31459));
OAI21X1 g106021(.A0 (n_31091), .A1 (n_30105), .B0 (n_31689), .Y(n_31458));
NAND2X2 g106027(.A (n_31126), .B (n_13026), .Y (n_31457));
NAND2X1 g105704(.A (n_6656), .B (n_31145), .Y (n_31455));
CLKBUFX1 gbuf_d_248(.A(n_31120), .Y(d_out_248));
CLKBUFX1 gbuf_q_248(.A(q_in_248), .Y(P2_reg2[12]));
NAND4X1 g106031(.A (n_31068), .B (n_15247), .C (n_30840), .D(n_30635), .Y (n_31454));
INVX1 g106034(.A (n_31337), .Y (n_31453));
NAND2X1 g105708(.A (n_6909), .B (n_31148), .Y (n_31452));
NAND4X1 g106050(.A (n_30216), .B (n_11087), .C (n_30898), .D(n_30158), .Y (n_31451));
OAI21X1 g106053(.A0 (n_33637), .A1 (n_29005), .B0 (n_24695), .Y(n_31450));
NAND2X1 g105718(.A (n_6911), .B (n_31144), .Y (n_31449));
NOR2X1 g106057(.A (n_26462), .B (n_35050), .Y (n_32920));
NAND2X1 g106070(.A (n_6944), .B (n_31143), .Y (n_31447));
NAND2X1 g106078(.A (n_7121), .B (n_31147), .Y (n_31446));
NAND2X1 g106085(.A (n_6912), .B (n_31141), .Y (n_31445));
CLKBUFX1 gbuf_d_249(.A(n_31115), .Y(d_out_249));
CLKBUFX1 gbuf_q_249(.A(q_in_249), .Y(n_4445));
CLKBUFX1 gbuf_d_250(.A(n_31114), .Y(d_out_250));
CLKBUFX1 gbuf_q_250(.A(q_in_250), .Y(n_10156));
CLKBUFX1 gbuf_d_251(.A(n_31257), .Y(d_out_251));
CLKBUFX1 gbuf_q_251(.A(q_in_251), .Y(P1_reg1[12]));
CLKBUFX1 gbuf_d_252(.A(n_31121), .Y(d_out_252));
CLKBUFX1 gbuf_q_252(.A(q_in_252), .Y(n_4824));
CLKBUFX1 gbuf_d_253(.A(n_31124), .Y(d_out_253));
CLKBUFX1 gbuf_q_253(.A(q_in_253), .Y(P2_reg2[10]));
CLKBUFX1 gbuf_d_254(.A(n_31117), .Y(d_out_254));
CLKBUFX1 gbuf_qn_254(.A(qn_in_254), .Y(P3_reg_150));
CLKBUFX1 gbuf_d_255(.A(n_31116), .Y(d_out_255));
CLKBUFX1 gbuf_q_255(.A(q_in_255), .Y(P3_reg1[12]));
CLKBUFX1 gbuf_d_256(.A(n_31187), .Y(d_out_256));
CLKBUFX1 gbuf_q_256(.A(q_in_256), .Y(P2_reg2[11]));
CLKBUFX1 gbuf_d_257(.A(n_31188), .Y(d_out_257));
CLKBUFX1 gbuf_q_257(.A(q_in_257), .Y(n_10205));
CLKBUFX1 gbuf_d_258(.A(n_31222), .Y(d_out_258));
CLKBUFX1 gbuf_q_258(.A(q_in_258), .Y(P3_reg3[5]));
CLKBUFX1 gbuf_d_259(.A(n_31221), .Y(d_out_259));
CLKBUFX1 gbuf_q_259(.A(q_in_259), .Y(P3_reg3[6]));
CLKBUFX1 gbuf_d_260(.A(n_31153), .Y(d_out_260));
CLKBUFX1 gbuf_q_260(.A(q_in_260), .Y(P2_reg1[11]));
CLKBUFX1 gbuf_d_261(.A(n_31152), .Y(d_out_261));
CLKBUFX1 gbuf_q_261(.A(q_in_261), .Y(n_3416));
CLKBUFX1 gbuf_d_262(.A(n_31151), .Y(d_out_262));
CLKBUFX1 gbuf_q_262(.A(q_in_262), .Y(n_4561));
CLKBUFX1 gbuf_d_263(.A(n_31150), .Y(d_out_263));
CLKBUFX1 gbuf_q_263(.A(q_in_263), .Y(P2_reg_95));
AOI21X1 g106130(.A0 (n_10458), .A1 (n_31035), .B0 (n_31490), .Y(n_31444));
AOI21X1 g106131(.A0 (n_9386), .A1 (n_31036), .B0 (n_30702), .Y(n_31443));
NAND2X1 g106135(.A (n_31215), .B (n_31677), .Y (n_31441));
NAND2X1 g106137(.A (n_31213), .B (n_31677), .Y (n_32159));
OAI21X1 g105765(.A0 (n_30996), .A1 (n_9944), .B0 (n_31528), .Y(n_31439));
OAI21X1 g106142(.A0 (n_35694), .A1 (n_35695), .B0 (n_31845), .Y(n_35329));
NAND2X1 g106143(.A (n_31210), .B (n_31677), .Y (n_31437));
OAI21X1 g105767(.A0 (n_30995), .A1 (n_9895), .B0 (n_31644), .Y(n_31436));
OAI21X1 g106151(.A0 (n_8813), .A1 (n_31420), .B0 (n_31211), .Y(n_31435));
AOI21X1 g106152(.A0 (n_31032), .A1 (n_30799), .B0 (n_33125), .Y(n_31434));
NAND2X1 g106154(.A (n_31200), .B (n_31641), .Y (n_35131));
AOI21X1 g106158(.A0 (n_15039), .A1 (n_15413), .B0 (n_31190), .Y(n_31432));
AOI21X1 g105781(.A0 (n_30991), .A1 (n_30942), .B0 (n_8397), .Y(n_31431));
NAND2X1 g106171(.A (n_31198), .B (n_12892), .Y (n_31430));
OR4X1 g106186(.A (n_29762), .B (n_30471), .C (n_18284), .D (n_30826),.Y (n_31428));
OAI21X1 g106192(.A0 (n_31028), .A1 (n_30825), .B0 (n_31240), .Y(n_31426));
OAI21X1 g106198(.A0 (n_8865), .A1 (n_31307), .B0 (n_31193), .Y(n_31424));
OAI21X1 g106201(.A0 (n_8812), .A1 (n_31422), .B0 (n_31197), .Y(n_31423));
OAI21X1 g106203(.A0 (n_9783), .A1 (n_31420), .B0 (n_31192), .Y(n_35293));
NAND4X1 g106204(.A (n_32260), .B (n_29970), .C (n_32261), .D(n_26040), .Y (n_31419));
NOR2X1 g105799(.A (n_10466), .B (n_31164), .Y (n_31418));
NOR2X1 g106208(.A (n_6897), .B (n_31259), .Y (n_31417));
NOR2X1 g106211(.A (n_7091), .B (n_31263), .Y (n_31416));
OAI21X1 g106219(.A0 (n_8264), .A1 (n_31414), .B0 (n_31251), .Y(n_31415));
OAI21X1 g106221(.A0 (n_9868), .A1 (n_31299), .B0 (n_31249), .Y(n_31413));
OAI21X1 g106222(.A0 (n_31012), .A1 (n_8505), .B0 (n_10431), .Y(n_31412));
OAI21X1 g106233(.A0 (n_31027), .A1 (n_31410), .B0 (n_9910), .Y(n_31411));
OAI21X1 g106235(.A0 (n_8776), .A1 (n_31740), .B0 (n_31195), .Y(n_31408));
OAI21X1 g106237(.A0 (n_31017), .A1 (n_31936), .B0 (n_10352), .Y(n_31407));
OAI21X1 g105817(.A0 (n_30984), .A1 (n_31620), .B0 (n_10346), .Y(n_31406));
OAI21X1 g106241(.A0 (n_8592), .A1 (n_31414), .B0 (n_31241), .Y(n_31405));
NOR2X1 g106247(.A (n_9896), .B (n_31246), .Y (n_31404));
OAI21X1 g106250(.A0 (n_31024), .A1 (n_30485), .B0 (n_31402), .Y(n_31403));
NOR2X1 g105824(.A (n_10369), .B (n_31186), .Y (n_31401));
NOR2X1 g106256(.A (n_7001), .B (n_31113), .Y (n_31400));
AOI22X1 g106263(.A0 (n_31031), .A1 (n_31398), .B0 (n_8512), .B1(n_30881), .Y (n_31399));
NAND2X1 g106271(.A (n_6483), .B (n_31238), .Y (n_31397));
NAND2X1 g106286(.A (n_6728), .B (n_31262), .Y (n_31396));
NAND2X1 g106293(.A (n_6484), .B (n_31261), .Y (n_31395));
NAND2X1 g106298(.A (n_6515), .B (n_31228), .Y (n_31394));
NAND2X1 g106301(.A (n_6582), .B (n_31227), .Y (n_31393));
NAND2X1 g106303(.A (n_6708), .B (n_31224), .Y (n_31392));
NAND2X1 g105852(.A (n_6939), .B (n_31206), .Y (n_31391));
NAND2X1 g105865(.A (n_6870), .B (n_31202), .Y (n_31390));
AOI21X1 g106343(.A0 (n_10457), .A1 (n_30992), .B0 (n_31388), .Y(n_31389));
NAND2X1 g105873(.A (n_7048), .B (n_31066), .Y (n_31387));
NAND2X1 g106356(.A (n_31040), .B (n_31965), .Y (n_31386));
NAND2X1 g106363(.A (n_31021), .B (n_31698), .Y (n_31385));
NAND2X1 g106365(.A (n_31020), .B (n_31694), .Y (n_31384));
NOR2X1 g106373(.A (n_29985), .B (n_31004), .Y (n_31383));
CLKBUFX1 gbuf_d_264(.A(n_31060), .Y(d_out_264));
CLKBUFX1 gbuf_q_264(.A(q_in_264), .Y(P2_reg1[12]));
OAI21X1 g106399(.A0 (n_30810), .A1 (n_30492), .B0 (n_31628), .Y(n_31382));
AOI21X1 g106400(.A0 (n_30814), .A1 (n_30764), .B0 (n_31245), .Y(n_31381));
NAND3X1 g106414(.A (n_33806), .B (n_30095), .C (n_30820), .Y(n_35878));
NAND2X1 g106418(.A (n_31025), .B (n_31493), .Y (n_31379));
NOR3X1 g106421(.A (n_30117), .B (n_25176), .C (n_30794), .Y(n_31378));
NOR3X1 g106427(.A (n_30113), .B (n_25163), .C (n_30795), .Y(n_31377));
NAND2X1 g106436(.A (n_31009), .B (n_12822), .Y (n_31376));
NAND2X1 g106437(.A (n_31008), .B (n_12820), .Y (n_31375));
NOR2X1 g106446(.A (n_31010), .B (n_31006), .Y (n_31374));
NAND2X1 g106454(.A (n_31015), .B (n_31683), .Y (n_35262));
OAI21X1 g106467(.A0 (n_30809), .A1 (n_30576), .B0 (n_31628), .Y(n_31372));
NOR2X1 g106499(.A (n_8895), .B (n_31045), .Y (n_31371));
NOR2X1 g106500(.A (n_9381), .B (n_31043), .Y (n_31370));
NOR2X1 g106502(.A (n_9558), .B (n_31003), .Y (n_31369));
NOR2X1 g106504(.A (n_30543), .B (n_31014), .Y (n_31368));
NOR2X1 g106505(.A (n_9051), .B (n_31007), .Y (n_31367));
CLKBUFX1 gbuf_d_265(.A(n_30970), .Y(d_out_265));
CLKBUFX1 gbuf_q_265(.A(q_in_265), .Y(P3_reg2[9]));
NAND2X1 g105674(.A (n_30974), .B (n_12808), .Y (n_31366));
NOR2X1 g106518(.A (n_6854), .B (n_31054), .Y (n_31365));
OAI21X1 g106535(.A0 (n_9343), .A1 (n_31420), .B0 (n_34819), .Y(n_35900));
NOR2X1 g106539(.A (n_6997), .B (n_31058), .Y (n_31362));
AOI21X1 g105982(.A0 (n_30940), .A1 (n_30415), .B0 (n_31360), .Y(n_31361));
NAND2X1 g106546(.A (n_6942), .B (n_31037), .Y (n_31359));
NAND2X1 g106547(.A (n_6874), .B (n_31038), .Y (n_31358));
AOI21X1 g105984(.A0 (n_30966), .A1 (n_30414), .B0 (n_31360), .Y(n_31357));
OAI21X1 g106551(.A0 (n_30807), .A1 (n_33350), .B0 (n_6687), .Y(n_31356));
AOI21X1 g105988(.A0 (n_30965), .A1 (n_30416), .B0 (n_31360), .Y(n_31354));
NAND2X1 g106558(.A (n_7110), .B (n_31052), .Y (n_31353));
NAND2X1 g106564(.A (n_7107), .B (n_31051), .Y (n_31352));
OAI21X1 g106567(.A0 (n_30804), .A1 (P1_n_449), .B0 (n_7180), .Y(n_31351));
OR4X1 g105996(.A (n_30243), .B (n_10104), .C (n_29953), .D (n_30740),.Y (n_31350));
NAND2X1 g106569(.A (n_35429), .B (n_35430), .Y (n_31349));
OAI21X1 g106571(.A0 (n_30803), .A1 (n_33201), .B0 (n_6562), .Y(n_31348));
AOI21X1 g106587(.A0 (n_10398), .A1 (n_30959), .B0 (n_31586), .Y(n_31347));
NAND2X1 g106598(.A (n_30982), .B (n_31345), .Y (n_31346));
AOI21X1 g106600(.A0 (n_10405), .A1 (n_30957), .B0 (n_31343), .Y(n_31344));
NAND2X1 g106608(.A (n_31894), .B (n_35611), .Y (n_32283));
OAI21X1 g106020(.A0 (n_30948), .A1 (n_29781), .B0 (n_31689), .Y(n_31341));
NAND2X1 g106022(.A (n_30978), .B (n_13018), .Y (n_31340));
OAI21X1 g106030(.A0 (n_30933), .A1 (n_29383), .B0 (n_31555), .Y(n_31339));
OAI21X1 g106032(.A0 (n_30932), .A1 (n_28559), .B0 (n_31099), .Y(n_31338));
NAND4X1 g106035(.A (n_30239), .B (n_30139), .C (n_30584), .D(n_29504), .Y (n_31337));
OR4X1 g106037(.A (n_35300), .B (n_10113), .C (n_35299), .D (n_30739),.Y (n_31336));
NAND2X1 g106677(.A (n_30979), .B (n_30939), .Y (n_31335));
NAND2X1 g106678(.A (n_30976), .B (n_30937), .Y (n_31334));
NOR2X1 g106692(.A (n_9945), .B (n_30990), .Y (n_31333));
AOI22X1 g106060(.A0 (n_30949), .A1 (n_31601), .B0 (n_3205), .B1(n_9382), .Y (n_31332));
NOR2X1 g106701(.A (n_9931), .B (n_30989), .Y (n_31331));
OAI21X1 g106715(.A0 (n_9864), .A1 (n_31019), .B0 (n_30994), .Y(n_31330));
CLKBUFX1 gbuf_d_266(.A(n_31048), .Y(d_out_266));
CLKBUFX1 gbuf_q_266(.A(q_in_266), .Y(P1_reg3[8]));
CLKBUFX1 gbuf_d_267(.A(n_31018), .Y(d_out_267));
CLKBUFX1 gbuf_q_267(.A(q_in_267), .Y(n_4231));
CLKBUFX1 gbuf_d_268(.A(n_31013), .Y(d_out_268));
CLKBUFX1 gbuf_q_268(.A(q_in_268), .Y(n_10150));
CLKBUFX1 gbuf_d_269(.A(n_30972), .Y(d_out_269));
CLKBUFX1 gbuf_q_269(.A(q_in_269), .Y(P3_reg1[9]));
CLKBUFX1 gbuf_d_270(.A(n_31061), .Y(d_out_270));
CLKBUFX1 gbuf_q_270(.A(q_in_270), .Y(n_3716));
CLKBUFX1 gbuf_d_271(.A(n_31059), .Y(d_out_271));
CLKBUFX1 gbuf_q_271(.A(q_in_271), .Y(n_10221));
CLKBUFX1 gbuf_d_272(.A(n_31085), .Y(d_out_272));
CLKBUFX1 gbuf_q_272(.A(q_in_272), .Y(P1_reg3[5]));
CLKBUFX1 gbuf_d_273(.A(n_31002), .Y(d_out_273));
CLKBUFX1 gbuf_qn_273(.A(qn_in_273), .Y(P3_reg_145));
CLKBUFX1 gbuf_d_274(.A(n_31001), .Y(d_out_274));
CLKBUFX1 gbuf_qn_274(.A(qn_in_274), .Y(P3_reg_146));
CLKBUFX1 gbuf_d_275(.A(n_31000), .Y(d_out_275));
CLKBUFX1 gbuf_qn_275(.A(qn_in_275), .Y(P3_reg_148));
CLKBUFX1 gbuf_d_276(.A(n_30999), .Y(d_out_276));
CLKBUFX1 gbuf_q_276(.A(q_in_276), .Y(n_13681));
CLKBUFX1 gbuf_d_277(.A(n_31033), .Y(d_out_277));
CLKBUFX1 gbuf_q_277(.A(q_in_277), .Y(P2_reg3[7]));
OAI21X1 g106802(.A0 (n_30947), .A1 (n_31328), .B0 (n_6577), .Y(n_31329));
NAND4X1 g106133(.A (n_30755), .B (n_10170), .C (n_30676), .D(n_29913), .Y (n_31327));
NAND4X1 g106134(.A (n_30754), .B (n_10153), .C (n_30660), .D(n_29907), .Y (n_31326));
OAI21X1 g106148(.A0 (n_30904), .A1 (n_30334), .B0 (n_30403), .Y(n_31325));
NOR2X1 g106149(.A (n_9912), .B (n_31075), .Y (n_31324));
OAI21X1 g106150(.A0 (n_8693), .A1 (n_31420), .B0 (n_31074), .Y(n_31323));
NAND4X1 g106153(.A (n_30851), .B (n_30656), .C (n_19562), .D(n_30681), .Y (n_31322));
NAND2X1 g106875(.A (n_31094), .B (n_31677), .Y (n_31321));
OR4X1 g106157(.A (n_30135), .B (n_10120), .C (n_30133), .D (n_33721),.Y (n_31320));
NOR3X1 g106166(.A (n_30194), .B (n_26576), .C (n_33448), .Y(n_31319));
AOI21X1 g106168(.A0 (n_30901), .A1 (n_30331), .B0 (n_8377), .Y(n_31318));
NAND2X1 g106169(.A (n_31062), .B (n_12712), .Y (n_31316));
CLKBUFX1 gbuf_d_278(.A(n_31079), .Y(d_out_278));
CLKBUFX1 gbuf_q_278(.A(q_in_278), .Y(P3_reg3[7]));
NAND4X1 g106180(.A (n_30347), .B (n_30856), .C (n_30637), .D(n_30304), .Y (n_31315));
NAND4X1 g106188(.A (n_32066), .B (n_32067), .C (n_30651), .D(n_30292), .Y (n_31314));
NAND4X1 g106191(.A (n_30853), .B (n_30674), .C (n_30673), .D(n_21660), .Y (n_31313));
AOI21X1 g106194(.A0 (n_30908), .A1 (n_30552), .B0 (n_8377), .Y(n_31311));
OAI21X1 g106197(.A0 (n_8792), .A1 (n_31420), .B0 (n_31065), .Y(n_31310));
OAI21X1 g106199(.A0 (n_30899), .A1 (n_27557), .B0 (n_10450), .Y(n_31309));
OAI21X1 g106202(.A0 (n_9708), .A1 (n_31307), .B0 (n_31063), .Y(n_35610));
OR4X1 g105798(.A (n_29670), .B (n_29738), .C (n_21224), .D (n_30781),.Y (n_31306));
NAND4X1 g106205(.A (n_32028), .B (n_30590), .C (n_32029), .D(n_30554), .Y (n_31305));
NOR2X1 g106210(.A (n_6851), .B (n_31106), .Y (n_31304));
NOR3X1 g106215(.A (n_30188), .B (n_26909), .C (n_33382), .Y(n_31303));
NAND4X1 g106218(.A (n_28678), .B (n_9508), .C (n_30776), .D(n_29339), .Y (n_31302));
OAI21X1 g106220(.A0 (n_9860), .A1 (n_31639), .B0 (n_31103), .Y(n_31301));
OAI21X1 g106224(.A0 (n_9844), .A1 (n_31299), .B0 (n_31102), .Y(n_31300));
OAI21X1 g106225(.A0 (n_30867), .A1 (n_31936), .B0 (n_10739), .Y(n_31298));
NOR2X1 g106227(.A (n_30407), .B (n_33671), .Y (n_31297));
NOR2X1 g106232(.A (n_6893), .B (n_31082), .Y (n_31296));
NOR2X1 g107071(.A (n_9924), .B (n_31108), .Y (n_31295));
NOR2X1 g106244(.A (n_6783), .B (n_31109), .Y (n_31294));
NOR2X1 g106246(.A (n_9639), .B (n_31095), .Y (n_31293));
NOR2X1 g106249(.A (n_10400), .B (n_31101), .Y (n_31292));
NOR2X1 g106252(.A (n_7086), .B (n_30969), .Y (n_31291));
NOR2X1 g106254(.A (n_6855), .B (n_31111), .Y (n_31290));
OAI21X1 g107096(.A0 (n_9840), .A1 (n_30886), .B0 (n_33124), .Y(n_31289));
NAND2X1 g106262(.A (n_6529), .B (n_31110), .Y (n_31288));
OAI21X1 g106264(.A0 (n_8225), .A1 (n_31713), .B0 (n_31089), .Y(n_31287));
NAND2X1 g106268(.A (n_6921), .B (n_31093), .Y (n_31286));
NAND2X1 g106270(.A (n_35412), .B (n_35413), .Y (n_31285));
NAND2X1 g106275(.A (n_6753), .B (n_31096), .Y (n_31284));
NOR2X1 g105835(.A (n_6899), .B (n_31076), .Y (n_31283));
OAI21X1 g106280(.A0 (n_30891), .A1 (n_31726), .B0 (n_7109), .Y(n_31282));
OAI21X1 g106283(.A0 (n_30866), .A1 (n_31569), .B0 (n_6622), .Y(n_31281));
NAND2X1 g106287(.A (n_6612), .B (n_31107), .Y (n_31280));
OAI21X1 g106288(.A0 (n_30889), .A1 (n_31278), .B0 (n_6747), .Y(n_31279));
OAI21X1 g106292(.A0 (n_30888), .A1 (n_31278), .B0 (n_6688), .Y(n_31277));
OAI21X1 g106296(.A0 (n_30865), .A1 (n_31275), .B0 (n_6581), .Y(n_31276));
OAI21X1 g106300(.A0 (n_30864), .A1 (n_31273), .B0 (n_6521), .Y(n_31274));
NAND2X1 g105848(.A (n_7128), .B (n_31072), .Y (n_31272));
OAI21X1 g106302(.A0 (n_30882), .A1 (n_31726), .B0 (n_7103), .Y(n_31271));
NAND2X1 g105851(.A (n_6741), .B (n_31071), .Y (n_31270));
NAND2X1 g105860(.A (n_6745), .B (n_31069), .Y (n_31269));
NAND2X1 g105861(.A (n_7112), .B (n_31067), .Y (n_31268));
NAND4X1 g106346(.A (n_30489), .B (n_10220), .C (n_30548), .D(n_29453), .Y (n_31267));
NOR2X1 g106349(.A (n_30280), .B (n_30896), .Y (n_31266));
NOR2X1 g106350(.A (n_30921), .B (n_30257), .Y (n_31265));
NOR2X1 g106351(.A (n_33790), .B (n_30256), .Y (n_31264));
AOI21X1 g106361(.A0 (n_10406), .A1 (n_30621), .B0 (n_30968), .Y(n_31263));
NAND2X1 g106366(.A (n_30890), .B (n_31850), .Y (n_31262));
NAND2X1 g106368(.A (n_30887), .B (n_31260), .Y (n_31261));
AOI21X1 g106369(.A0 (n_9391), .A1 (n_30649), .B0 (n_31105), .Y(n_31259));
NOR2X1 g107305(.A (n_30913), .B (n_30895), .Y (n_31258));
OAI21X1 g105881(.A0 (n_30632), .A1 (n_31472), .B0 (n_6948), .Y(n_31257));
NAND4X1 g106374(.A (n_32147), .B (n_14622), .C (n_32148), .D(n_30168), .Y (n_31256));
AOI21X1 g106376(.A0 (n_30640), .A1 (n_30214), .B0 (n_8070), .Y(n_31255));
NAND3X1 g106377(.A (n_11146), .B (n_30488), .C (n_30669), .Y(n_31253));
NAND2X1 g106380(.A (n_30875), .B (n_21196), .Y (n_31252));
OAI21X1 g106383(.A0 (n_30700), .A1 (n_30328), .B0 (n_31573), .Y(n_31251));
AOI21X1 g106384(.A0 (n_30698), .A1 (n_30213), .B0 (n_8070), .Y(n_31250));
OAI21X1 g106386(.A0 (n_30662), .A1 (n_30177), .B0 (n_33123), .Y(n_31249));
NAND2X1 g106396(.A (n_30878), .B (n_26002), .Y (n_31248));
AOI21X1 g106391(.A0 (n_30697), .A1 (n_30211), .B0 (n_8070), .Y(n_31247));
AOI21X1 g106402(.A0 (n_30658), .A1 (n_30512), .B0 (n_31245), .Y(n_31246));
NAND2X1 g106404(.A (n_30844), .B (n_30869), .Y (n_31244));
NOR2X1 g106405(.A (n_30841), .B (n_30868), .Y (n_31243));
OAI21X1 g106406(.A0 (n_30648), .A1 (n_29653), .B0 (n_31174), .Y(n_31242));
OAI21X1 g106408(.A0 (n_30629), .A1 (n_29642), .B0 (n_31240), .Y(n_31241));
OR4X1 g106410(.A (n_29749), .B (n_10117), .C (n_29324), .D (n_30562),.Y (n_31239));
NAND2X1 g106417(.A (n_30894), .B (n_31493), .Y (n_31238));
AOI21X1 g106420(.A0 (n_30225), .A1 (n_30639), .B0 (n_31236), .Y(n_31237));
AOI21X1 g106426(.A0 (n_30664), .A1 (n_30191), .B0 (n_31233), .Y(n_31234));
NOR2X1 g106430(.A (n_25843), .B (n_30876), .Y (n_31232));
NAND2X1 g106445(.A (n_30873), .B (n_30341), .Y (n_31230));
NAND2X1 g106447(.A (n_30885), .B (n_30838), .Y (n_31229));
NAND2X1 g106448(.A (n_30884), .B (n_31698), .Y (n_31228));
NAND2X1 g106449(.A (n_30883), .B (n_31260), .Y (n_31227));
NAND2X1 g106450(.A (n_30858), .B (n_30835), .Y (n_31226));
NAND2X1 g106451(.A (n_30880), .B (n_30850), .Y (n_31225));
NAND2X1 g106452(.A (n_30879), .B (n_31683), .Y (n_31224));
NAND3X1 g106456(.A (n_32200), .B (n_32201), .C (n_30679), .Y(n_31223));
NAND2X1 g106457(.A (n_30859), .B (n_13001), .Y (n_31222));
NAND2X1 g106458(.A (n_30862), .B (n_12995), .Y (n_31221));
NOR2X1 g106470(.A (n_26440), .B (n_30854), .Y (n_31220));
NOR2X1 g106473(.A (n_30900), .B (n_30591), .Y (n_31218));
NOR2X1 g106478(.A (n_10246), .B (n_30857), .Y (n_32132));
OAI21X1 g106479(.A0 (n_8861), .A1 (n_31740), .B0 (n_30915), .Y(n_31215));
NAND3X1 g106480(.A (n_32265), .B (n_32266), .C (n_29491), .Y(n_31214));
OAI21X1 g106483(.A0 (n_8795), .A1 (n_31307), .B0 (n_30912), .Y(n_31213));
NAND3X1 g106484(.A (n_35080), .B (n_35081), .C (n_29489), .Y(n_31212));
OAI21X1 g106489(.A0 (n_30667), .A1 (n_29797), .B0 (n_34731), .Y(n_31211));
OAI21X1 g106490(.A0 (n_8811), .A1 (n_31307), .B0 (n_30910), .Y(n_31210));
OAI21X1 g106491(.A0 (n_30631), .A1 (n_29437), .B0 (n_27485), .Y(n_31209));
OAI21X1 g106493(.A0 (n_30666), .A1 (n_29795), .B0 (n_30958), .Y(n_31208));
NOR2X1 g106495(.A (n_8898), .B (n_30917), .Y (n_31207));
NAND2X1 g105953(.A (n_30818), .B (n_31205), .Y (n_31206));
NOR2X1 g106508(.A (n_8726), .B (n_30916), .Y (n_31204));
AOI21X1 g106513(.A0 (n_30190), .A1 (n_30647), .B0 (n_31236), .Y(n_31203));
NAND2X1 g105962(.A (n_30812), .B (n_31201), .Y (n_31202));
OAI21X1 g106523(.A0 (n_8587), .A1 (n_31199), .B0 (n_30902), .Y(n_31200));
NOR2X1 g106524(.A (n_6782), .B (n_30924), .Y (n_31198));
OAI21X1 g106530(.A0 (n_30628), .A1 (n_30119), .B0 (n_30958), .Y(n_31197));
NAND2X1 g105974(.A (n_30808), .B (n_31891), .Y (n_31196));
OAI21X1 g106533(.A0 (n_30614), .A1 (n_30120), .B0 (n_30958), .Y(n_31195));
OAI21X1 g106536(.A0 (n_30630), .A1 (n_29801), .B0 (n_31544), .Y(n_31193));
OAI21X1 g106537(.A0 (n_30627), .A1 (n_29798), .B0 (n_34731), .Y(n_31192));
NAND3X1 g106541(.A (n_32145), .B (n_30072), .C (n_32146), .Y(n_31190));
NAND4X1 g106543(.A (n_7427), .B (n_30897), .C (n_29944), .D(n_30333), .Y (n_31189));
OAI21X1 g106544(.A0 (n_30622), .A1 (n_31472), .B0 (n_6850), .Y(n_31188));
OAI21X1 g106552(.A0 (n_30624), .A1 (n_33201), .B0 (n_6655), .Y(n_31187));
AOI21X1 g105987(.A0 (n_30759), .A1 (n_30456), .B0 (n_33125), .Y(n_31186));
NAND3X1 g105686(.A (n_30905), .B (n_30721), .C (n_29669), .Y(n_35669));
CLKBUFX1 gbuf_d_279(.A(n_30793), .Y(d_out_279));
CLKBUFX1 gbuf_q_279(.A(q_in_279), .Y(n_13721));
NOR2X1 g106590(.A (n_30831), .B (n_29493), .Y (n_31184));
NOR2X1 g106592(.A (n_30830), .B (n_29490), .Y (n_31183));
NAND2X1 g106604(.A (n_30805), .B (n_31205), .Y (n_31182));
NAND4X1 g106615(.A (n_30451), .B (n_14704), .C (n_30455), .D(n_30110), .Y (n_31181));
AOI21X1 g106620(.A0 (n_30582), .A1 (n_30496), .B0 (n_31178), .Y(n_31180));
AOI21X1 g106621(.A0 (n_30581), .A1 (n_30495), .B0 (n_31178), .Y(n_31179));
AOI21X1 g106625(.A0 (n_30580), .A1 (n_30494), .B0 (n_8070), .Y(n_31177));
AOI21X1 g106626(.A0 (n_30579), .A1 (n_30493), .B0 (n_31041), .Y(n_31176));
OAI21X1 g106633(.A0 (n_30782), .A1 (n_30227), .B0 (n_31174), .Y(n_31175));
AOI21X1 g106647(.A0 (n_30578), .A1 (n_30127), .B0 (n_8377), .Y(n_31173));
AOI21X1 g106652(.A0 (n_30577), .A1 (n_30727), .B0 (n_31236), .Y(n_31171));
NAND3X1 g106653(.A (n_30061), .B (n_30565), .C (n_30010), .Y(n_31170));
AOI21X1 g106655(.A0 (n_30777), .A1 (n_30125), .B0 (n_31236), .Y(n_31169));
NAND4X1 g106657(.A (n_35078), .B (n_29247), .C (n_35079), .D(n_25328), .Y (n_31168));
AOI21X1 g106669(.A0 (n_10743), .A1 (n_30766), .B0 (n_7058), .Y(n_31167));
NAND3X1 g106673(.A (n_30215), .B (n_30571), .C (n_30531), .Y(n_31165));
AOI21X1 g106046(.A0 (n_30750), .A1 (n_30002), .B0 (n_31523), .Y(n_31164));
OAI21X1 g106682(.A0 (n_30780), .A1 (n_30223), .B0 (n_31628), .Y(n_31162));
OAI21X1 g106683(.A0 (n_30779), .A1 (n_30222), .B0 (n_31160), .Y(n_31161));
NOR2X1 g106052(.A (n_30467), .B (n_30819), .Y (n_31159));
OAI21X1 g106707(.A0 (n_9772), .A1 (n_31131), .B0 (n_30817), .Y(n_31158));
NOR2X1 g106722(.A (n_10360), .B (n_30824), .Y (n_31157));
NOR2X1 g106725(.A (n_30473), .B (n_30801), .Y (n_31156));
NOR2X1 g106727(.A (n_30174), .B (n_30800), .Y (n_31155));
NOR2X1 g106766(.A (n_9890), .B (n_30823), .Y (n_31154));
CLKBUFX1 gbuf_d_280(.A(n_30791), .Y(d_out_280));
CLKBUFX1 gbuf_q_280(.A(q_in_280), .Y(P3_reg2[10]));
CLKBUFX1 gbuf_d_281(.A(n_30944), .Y(d_out_281));
CLKBUFX1 gbuf_q_281(.A(q_in_281), .Y(P2_reg3[5]));
CLKBUFX1 gbuf_d_282(.A(n_30848), .Y(d_out_282));
CLKBUFX1 gbuf_q_282(.A(q_in_282), .Y(n_4554));
CLKBUFX1 gbuf_d_283(.A(n_30846), .Y(d_out_283));
CLKBUFX1 gbuf_q_283(.A(q_in_283), .Y(n_10138));
CLKBUFX1 gbuf_d_284(.A(n_30907), .Y(d_out_284));
CLKBUFX1 gbuf_q_284(.A(q_in_284), .Y(P2_reg3[6]));
CLKBUFX1 gbuf_d_285(.A(n_30906), .Y(d_out_285));
CLKBUFX1 gbuf_q_285(.A(q_in_285), .Y(P3_reg3[4]));
CLKBUFX1 gbuf_d_286(.A(n_30790), .Y(d_out_286));
CLKBUFX1 gbuf_q_286(.A(q_in_286), .Y(n_3402));
CLKBUFX1 gbuf_d_287(.A(n_30789), .Y(d_out_287));
CLKBUFX1 gbuf_q_287(.A(q_in_287), .Y(n_4344));
CLKBUFX1 gbuf_d_288(.A(n_30788), .Y(d_out_288));
CLKBUFX1 gbuf_q_288(.A(q_in_288), .Y(n_10140));
OAI21X1 g106801(.A0 (n_30775), .A1 (n_31328), .B0 (n_6659), .Y(n_31153));
NAND2X1 g106806(.A (n_6919), .B (n_30833), .Y (n_31152));
NAND2X1 g106807(.A (n_7122), .B (n_30832), .Y (n_31151));
OAI21X1 g106827(.A0 (n_30768), .A1 (n_31149), .B0 (n_6526), .Y(n_31150));
NAND2X1 g105763(.A (n_30927), .B (n_31201), .Y (n_31148));
NAND2X1 g106145(.A (n_30931), .B (n_31092), .Y (n_31147));
NOR2X1 g105768(.A (n_8905), .B (n_30926), .Y (n_31146));
NAND2X1 g105770(.A (n_30929), .B (n_31594), .Y (n_31145));
NAND2X1 g105772(.A (n_30919), .B (n_31912), .Y (n_31144));
CLKBUFX1 gbuf_d_289(.A(n_30847), .Y(d_out_289));
CLKBUFX1 gbuf_qn_289(.A(qn_in_289), .Y(P3_reg_147));
NAND2X1 g106163(.A (n_30936), .B (n_31641), .Y (n_31143));
NAND2X1 g106182(.A (n_30934), .B (n_31201), .Y (n_31141));
NAND2X1 g106187(.A (n_30952), .B (n_30938), .Y (n_31139));
NOR2X1 g106953(.A (n_30946), .B (n_30941), .Y (n_31138));
OAI21X1 g106212(.A0 (n_9290), .A1 (n_31420), .B0 (n_30945), .Y(n_31137));
NOR2X1 g106223(.A (n_9902), .B (n_30953), .Y (n_31135));
NOR2X1 g106226(.A (n_30382), .B (n_30930), .Y (n_31134));
NOR3X1 g106230(.A (n_8686), .B (n_8013), .C (n_30709), .Y (n_31133));
OAI21X1 g107056(.A0 (n_8842), .A1 (n_31131), .B0 (n_30964), .Y(n_31132));
OAI21X1 g107072(.A0 (n_9778), .A1 (n_31129), .B0 (n_30961), .Y(n_31130));
NOR2X1 g106248(.A (n_9889), .B (n_30951), .Y (n_31128));
NOR2X1 g106251(.A (n_7065), .B (n_30785), .Y (n_31127));
NOR2X1 g106253(.A (n_7082), .B (n_30967), .Y (n_31126));
NOR2X1 g106258(.A (n_6900), .B (n_30784), .Y (n_31125));
OAI21X1 g106260(.A0 (n_30744), .A1 (n_31149), .B0 (n_6645), .Y(n_31124));
OAI21X1 g107103(.A0 (n_8810), .A1 (n_31122), .B0 (n_30954), .Y(n_31123));
OAI21X1 g106269(.A0 (n_30722), .A1 (n_31726), .B0 (n_7123), .Y(n_31121));
OAI21X1 g106276(.A0 (n_30729), .A1 (n_33201), .B0 (n_6628), .Y(n_31120));
AOI22X1 g107132(.A0 (n_30737), .A1 (n_31878), .B0 (n_9360), .B1(n_31876), .Y (n_31119));
AOI22X1 g107133(.A0 (n_30736), .A1 (n_31878), .B0 (n_9351), .B1(n_31495), .Y (n_31118));
NAND2X1 g106281(.A (n_6591), .B (n_30962), .Y (n_31117));
OAI21X1 g106290(.A0 (n_30719), .A1 (n_31958), .B0 (n_6740), .Y(n_31116));
NAND2X1 g105850(.A (n_35644), .B (n_35645), .Y (n_31115));
OAI21X1 g105863(.A0 (n_30652), .A1 (n_31541), .B0 (n_6924), .Y(n_31114));
AOI21X1 g106342(.A0 (n_10463), .A1 (n_30684), .B0 (n_31388), .Y(n_31113));
NAND4X1 g106344(.A (n_30491), .B (n_10248), .C (n_30561), .D(n_29457), .Y (n_31112));
AOI21X1 g106347(.A0 (n_10734), .A1 (n_30408), .B0 (n_31081), .Y(n_31111));
NAND2X1 g106359(.A (n_30743), .B (n_31493), .Y (n_31110));
AOI21X1 g106360(.A0 (n_10407), .A1 (n_30393), .B0 (n_16415), .Y(n_31109));
AOI21X1 g107289(.A0 (n_30429), .A1 (n_30009), .B0 (n_30537), .Y(n_31108));
NAND2X1 g106367(.A (n_30728), .B (n_31781), .Y (n_31107));
AOI21X1 g106370(.A0 (n_8610), .A1 (n_30381), .B0 (n_31105), .Y(n_31106));
NAND4X1 g106371(.A (n_32564), .B (n_14965), .C (n_32565), .D(n_29881), .Y (n_31104));
OAI21X1 g106385(.A0 (n_30389), .A1 (n_29886), .B0 (n_33123), .Y(n_31103));
OAI21X1 g106388(.A0 (n_30384), .A1 (n_29651), .B0 (n_33123), .Y(n_31102));
AOI21X1 g106394(.A0 (n_30362), .A1 (n_29883), .B0 (n_33125), .Y(n_31101));
OAI21X1 g106395(.A0 (n_30339), .A1 (n_29222), .B0 (n_31099), .Y(n_31100));
NAND2X1 g106397(.A (n_30732), .B (n_31097), .Y (n_35412));
NAND2X1 g106398(.A (n_30730), .B (n_31097), .Y (n_31096));
AOI21X1 g106401(.A0 (n_30388), .A1 (n_30259), .B0 (n_31245), .Y(n_31095));
OAI21X1 g107388(.A0 (n_9774), .A1 (n_31131), .B0 (n_30746), .Y(n_31094));
NAND2X1 g106407(.A (n_30723), .B (n_31092), .Y (n_31093));
OR4X1 g106412(.A (n_29325), .B (n_10115), .C (n_29323), .D (n_30326),.Y (n_31091));
CLKBUFX1 gbuf_d_290(.A(n_30685), .Y(d_out_290));
CLKBUFX1 gbuf_q_290(.A(q_in_290), .Y(P1_reg3[4]));
NAND3X1 g106419(.A (n_30726), .B (n_30093), .C (n_30397), .Y(n_31090));
OAI21X1 g106428(.A0 (n_30379), .A1 (n_29935), .B0 (n_30403), .Y(n_31089));
NAND2X1 g106435(.A (n_30717), .B (n_12824), .Y (n_31085));
NOR2X1 g106441(.A (n_30244), .B (n_30742), .Y (n_31084));
NOR2X1 g106442(.A (n_30233), .B (n_30741), .Y (n_31083));
AOI21X1 g106453(.A0 (n_10737), .A1 (n_30364), .B0 (n_31081), .Y(n_31082));
NAND2X1 g106459(.A (n_30718), .B (n_12999), .Y (n_31079));
AOI21X1 g105940(.A0 (n_9955), .A1 (n_30517), .B0 (n_30783), .Y(n_31076));
AOI21X1 g106487(.A0 (n_30395), .A1 (n_29444), .B0 (n_31523), .Y(n_31075));
OAI21X1 g106488(.A0 (n_30394), .A1 (n_29443), .B0 (n_31064), .Y(n_31074));
OAI21X1 g106492(.A0 (n_30392), .A1 (n_29436), .B0 (n_30956), .Y(n_31073));
NAND2X1 g105950(.A (n_30692), .B (n_31912), .Y (n_31072));
NAND2X1 g105952(.A (n_30665), .B (n_31683), .Y (n_31071));
NAND3X1 g106501(.A (n_10212), .B (n_30088), .C (n_30387), .Y(n_31070));
NAND2X1 g105955(.A (n_30659), .B (n_31590), .Y (n_31069));
NOR2X1 g106503(.A (n_9188), .B (n_30713), .Y (n_31068));
NAND2X1 g105956(.A (n_30657), .B (n_31205), .Y (n_31067));
NAND2X1 g105968(.A (n_30682), .B (n_31891), .Y (n_31066));
OAI21X1 g106529(.A0 (n_30375), .A1 (n_29802), .B0 (n_31064), .Y(n_31065));
OAI21X1 g106531(.A0 (n_30373), .A1 (n_29799), .B0 (n_30958), .Y(n_31063));
NOR2X1 g106538(.A (n_6999), .B (n_30747), .Y (n_31062));
NAND2X1 g106545(.A (n_6992), .B (n_30738), .Y (n_31061));
OAI21X1 g106549(.A0 (n_30374), .A1 (n_31328), .B0 (n_6614), .Y(n_31060));
NAND2X1 g106563(.A (n_6881), .B (n_30735), .Y (n_31059));
AOI21X1 g106586(.A0 (n_9015), .A1 (n_30330), .B0 (n_34676), .Y(n_31058));
NAND4X1 g106588(.A (n_30076), .B (n_10160), .C (n_30185), .D(n_29909), .Y (n_31056));
NAND4X1 g106589(.A (n_30075), .B (n_10177), .C (n_30167), .D(n_29905), .Y (n_31055));
AOI21X1 g106594(.A0 (n_10455), .A1 (n_30516), .B0 (n_7058), .Y(n_31054));
NAND2X1 g106601(.A (n_30620), .B (n_31205), .Y (n_31052));
NAND2X1 g106603(.A (n_30617), .B (n_31205), .Y (n_31051));
NAND2X1 g106605(.A (n_30615), .B (n_31683), .Y (n_35429));
NOR2X1 g106611(.A (n_30583), .B (n_30626), .Y (n_31049));
NAND2X1 g106015(.A (n_30616), .B (n_12730), .Y (n_31048));
NAND3X1 g106613(.A (n_20750), .B (n_29454), .C (n_30549), .Y(n_31047));
NAND2X1 g106617(.A (n_30595), .B (n_11328), .Y (n_31046));
AOI21X1 g106622(.A0 (n_30338), .A1 (n_30534), .B0 (n_31233), .Y(n_31045));
AOI21X1 g106623(.A0 (n_30337), .A1 (n_30212), .B0 (n_31233), .Y(n_31043));
AOI21X1 g106627(.A0 (n_30336), .A1 (n_30210), .B0 (n_31041), .Y(n_35694));
OAI21X1 g106631(.A0 (n_8862), .A1 (n_35012), .B0 (n_30623), .Y(n_31040));
NAND2X1 g106634(.A (n_30611), .B (n_31894), .Y (n_31038));
NAND2X1 g106635(.A (n_31641), .B (n_35648), .Y (n_31037));
OAI21X1 g106636(.A0 (n_30553), .A1 (n_30228), .B0 (n_7827), .Y(n_31036));
OAI21X1 g106637(.A0 (n_30540), .A1 (n_29113), .B0 (n_29633), .Y(n_31035));
OR4X1 g106038(.A (n_29655), .B (n_10111), .C (n_29657), .D (n_33663),.Y (n_31034));
NAND2X1 g106660(.A (n_30598), .B (n_12890), .Y (n_31033));
NOR2X1 g106665(.A (n_30136), .B (n_30678), .Y (n_31032));
NAND4X1 g106674(.A (n_30224), .B (n_29057), .C (n_29777), .D(n_30189), .Y (n_31031));
CLKBUFX1 gbuf_d_291(.A(n_30610), .Y(d_out_291));
CLKBUFX1 gbuf_q_291(.A(q_in_291), .Y(n_13645));
NAND4X1 g106685(.A (n_35646), .B (n_35647), .C (n_30221), .D(n_29927), .Y (n_31028));
NOR2X1 g106691(.A (n_30699), .B (n_30643), .Y (n_31027));
NOR2X1 g106695(.A (n_9089), .B (n_30605), .Y (n_32571));
OAI21X1 g106699(.A0 (n_8845), .A1 (n_30893), .B0 (n_30599), .Y(n_31025));
NAND4X1 g106700(.A (n_32290), .B (n_29026), .C (n_32291), .D(n_25296), .Y (n_31024));
NOR2X1 g106702(.A (n_9082), .B (n_30596), .Y (n_31023));
OAI21X1 g106714(.A0 (n_9845), .A1 (n_30447), .B0 (n_30687), .Y(n_31021));
OAI21X1 g106716(.A0 (n_9852), .A1 (n_31019), .B0 (n_30686), .Y(n_31020));
NAND2X1 g106071(.A (n_6932), .B (n_30705), .Y (n_31018));
NOR2X1 g106726(.A (n_29884), .B (n_30613), .Y (n_31017));
OAI21X1 g106734(.A0 (n_30050), .A1 (n_29833), .B0 (n_30601), .Y(n_31016));
OAI21X1 g106738(.A0 (n_8793), .A1 (n_35012), .B0 (n_30597), .Y(n_31015));
NAND4X1 g106744(.A (n_30771), .B (n_15072), .C (n_29827), .D(n_29415), .Y (n_31014));
NAND2X1 g106086(.A (n_6933), .B (n_30704), .Y (n_31013));
NOR2X1 g106751(.A (n_30176), .B (n_30661), .Y (n_31012));
CLKBUFX1 gbuf_d_292(.A(n_30706), .Y(d_out_292));
CLKBUFX1 gbuf_q_292(.A(q_in_292), .Y(n_13515));
CLKBUFX1 gbuf_d_293(.A(n_30612), .Y(d_out_293));
CLKBUFX1 gbuf_q_293(.A(q_in_293), .Y(n_14135));
CLKBUFX1 gbuf_d_294(.A(n_30608), .Y(d_out_294));
CLKBUFX1 gbuf_q_294(.A(q_in_294), .Y(n_4230));
CLKBUFX1 gbuf_d_295(.A(n_30606), .Y(d_out_295));
CLKBUFX1 gbuf_q_295(.A(q_in_295), .Y(n_14096));
CLKBUFX1 gbuf_d_296(.A(n_30765), .Y(d_out_296));
CLKBUFX1 gbuf_q_296(.A(q_in_296), .Y(P1_reg3[3]));
CLKBUFX1 gbuf_d_297(.A(n_30716), .Y(d_out_297));
CLKBUFX1 gbuf_q_297(.A(q_in_297), .Y(n_10443));
CLKBUFX1 gbuf_d_298(.A(n_30715), .Y(d_out_298));
CLKBUFX1 gbuf_q_298(.A(q_in_298), .Y(P2_reg1[5]));
CLKBUFX1 gbuf_d_299(.A(n_30714), .Y(d_out_299));
CLKBUFX1 gbuf_q_299(.A(q_in_299), .Y(n_3709));
CLKBUFX1 gbuf_d_300(.A(n_30712), .Y(d_out_300));
CLKBUFX1 gbuf_q_300(.A(q_in_300), .Y(P3_reg1[5]));
CLKBUFX1 gbuf_d_301(.A(n_30708), .Y(d_out_301));
CLKBUFX1 gbuf_q_301(.A(q_in_301), .Y(n_13498));
CLKBUFX1 gbuf_d_302(.A(n_30707), .Y(d_out_302));
CLKBUFX1 gbuf_q_302(.A(q_in_302), .Y(P3_reg2[6]));
CLKBUFX1 gbuf_d_303(.A(n_30585), .Y(d_out_303));
CLKBUFX1 gbuf_q_303(.A(q_in_303), .Y(n_3724));
NAND2X1 g106778(.A (n_30644), .B (n_15491), .Y (n_31010));
NOR2X1 g106781(.A (n_6998), .B (n_30703), .Y (n_31009));
NOR2X1 g106782(.A (n_6896), .B (n_30701), .Y (n_31008));
NAND2X1 g106790(.A (n_30655), .B (n_20124), .Y (n_31007));
NAND2X1 g106792(.A (n_30646), .B (n_30299), .Y (n_31006));
NAND2X1 g106794(.A (n_30302), .B (n_30642), .Y (n_31004));
OAI21X1 g106809(.A0 (n_20114), .A1 (n_25540), .B0 (n_30638), .Y(n_31003));
NAND2X1 g106812(.A (n_6587), .B (n_30696), .Y (n_31002));
NAND2X1 g106813(.A (n_6695), .B (n_30695), .Y (n_31001));
NAND2X1 g106815(.A (n_6579), .B (n_30689), .Y (n_31000));
NAND2X1 g106820(.A (n_6736), .B (n_30694), .Y (n_30999));
NAND2X1 g106821(.A (n_30634), .B (n_20107), .Y (n_30998));
CLKBUFX1 gbuf_d_304(.A(n_30711), .Y(d_out_304));
CLKBUFX1 gbuf_q_304(.A(q_in_304), .Y(P3_reg1[6]));
AOI21X1 g106162(.A0 (n_30475), .A1 (n_29711), .B0 (n_31523), .Y(n_30996));
AOI21X1 g106165(.A0 (n_30474), .A1 (n_29710), .B0 (n_31523), .Y(n_30995));
OAI21X1 g106900(.A0 (n_30476), .A1 (n_28887), .B0 (n_33123), .Y(n_30994));
NAND3X1 g106177(.A (n_27548), .B (n_28516), .C (n_30463), .Y(n_30993));
OAI21X1 g106921(.A0 (n_30457), .A1 (n_26472), .B0 (n_30683), .Y(n_30992));
NOR2X1 g106179(.A (n_30043), .B (n_30773), .Y (n_30991));
AOI21X1 g106948(.A0 (n_30498), .A1 (n_30160), .B0 (n_31564), .Y(n_30990));
AOI21X1 g106951(.A0 (n_30497), .A1 (n_30126), .B0 (n_31564), .Y(n_30989));
NAND3X1 g106952(.A (n_30774), .B (n_29624), .C (n_30481), .Y(n_30988));
NOR2X1 g105802(.A (n_30748), .B (n_30745), .Y (n_30987));
NOR3X1 g106216(.A (n_29591), .B (n_26373), .C (n_30441), .Y(n_30986));
NOR2X1 g106228(.A (n_29766), .B (n_30757), .Y (n_30984));
NOR2X1 g107047(.A (n_30040), .B (n_30778), .Y (n_30983));
OAI21X1 g107073(.A0 (n_30468), .A1 (n_29681), .B0 (n_10420), .Y(n_30982));
NOR2X1 g107078(.A (n_8721), .B (n_30575), .Y (n_30981));
NOR2X1 g107083(.A (n_9383), .B (n_30573), .Y (n_30980));
NOR2X1 g107084(.A (n_30183), .B (n_30762), .Y (n_30979));
NOR2X1 g106255(.A (n_7075), .B (n_30568), .Y (n_30978));
NOR2X1 g107099(.A (n_9385), .B (n_30572), .Y (n_30977));
NOR2X1 g107105(.A (n_30166), .B (n_30761), .Y (n_30976));
OAI21X1 g107120(.A0 (n_30466), .A1 (n_34336), .B0 (n_10480), .Y(n_30975));
NOR2X1 g105833(.A (n_6852), .B (n_30751), .Y (n_30974));
OAI21X1 g107129(.A0 (n_8593), .A1 (n_31713), .B0 (n_30570), .Y(n_35611));
OAI21X1 g106295(.A0 (n_30442), .A1 (n_30792), .B0 (n_6571), .Y(n_30972));
OAI21X1 g106304(.A0 (n_30437), .A1 (n_31273), .B0 (n_6756), .Y(n_30970));
AOI21X1 g106338(.A0 (n_10283), .A1 (n_30361), .B0 (n_30968), .Y(n_30969));
AOI21X1 g106348(.A0 (n_10355), .A1 (n_30100), .B0 (n_31081), .Y(n_30967));
NOR2X1 g106352(.A (n_30470), .B (n_29969), .Y (n_30966));
NOR2X1 g106353(.A (n_30469), .B (n_29971), .Y (n_30965));
OAI21X1 g107282(.A0 (n_30129), .A1 (n_29293), .B0 (n_31544), .Y(n_30964));
NAND2X1 g106362(.A (n_30448), .B (n_31781), .Y (n_30962));
OAI21X1 g107291(.A0 (n_30108), .A1 (n_30008), .B0 (n_31402), .Y(n_30961));
NOR2X1 g107293(.A (n_30460), .B (n_30450), .Y (n_30960));
OAI21X1 g107301(.A0 (n_30116), .A1 (n_28832), .B0 (n_30958), .Y(n_30959));
OAI21X1 g107302(.A0 (n_30115), .A1 (n_29261), .B0 (n_30956), .Y(n_30957));
CLKBUFX1 gbuf_d_305(.A(n_30482), .Y(d_out_305));
CLKBUFX1 gbuf_q_305(.A(q_in_305), .Y(n_3668));
NAND3X1 g107339(.A (n_32171), .B (n_29441), .C (n_32172), .Y(n_30955));
OAI21X1 g107347(.A0 (n_30128), .A1 (n_29291), .B0 (n_31544), .Y(n_30954));
AOI21X1 g106387(.A0 (n_30083), .A1 (n_29652), .B0 (n_8397), .Y(n_30953));
NOR2X1 g106392(.A (n_30047), .B (n_30459), .Y (n_30952));
AOI21X1 g106393(.A0 (n_30048), .A1 (n_29561), .B0 (n_33125), .Y(n_30951));
OAI21X1 g106409(.A0 (n_30084), .A1 (n_31360), .B0 (n_9420), .Y(n_30949));
OR4X1 g106411(.A (n_28979), .B (n_10105), .C (n_33737), .D (n_30022),.Y (n_30948));
NOR2X1 g107399(.A (n_9933), .B (n_30487), .Y (n_30947));
OAI21X1 g107403(.A0 (n_29771), .A1 (n_29388), .B0 (n_22480), .Y(n_30946));
OAI21X1 g106425(.A0 (n_30055), .A1 (n_29648), .B0 (n_35008), .Y(n_30945));
NAND2X1 g106432(.A (n_30436), .B (n_12877), .Y (n_30944));
NOR2X1 g106466(.A (n_30472), .B (n_30132), .Y (n_30942));
OAI21X1 g107523(.A0 (n_29020), .A1 (n_10790), .B0 (n_30480), .Y(n_30941));
NOR2X1 g106469(.A (n_26391), .B (n_30435), .Y (n_30940));
INVX1 g107524(.A (n_30753), .Y (n_30939));
AOI21X1 g106471(.A0 (n_15296), .A1 (n_30530), .B0 (n_30453), .Y(n_30938));
INVX1 g107528(.A (n_30752), .Y (n_30937));
OAI21X1 g106481(.A0 (n_30086), .A1 (n_30935), .B0 (n_8616), .Y(n_30936));
OAI21X1 g106506(.A0 (n_30082), .A1 (n_30935), .B0 (n_8611), .Y(n_30934));
OR4X1 g106507(.A (n_28537), .B (n_10268), .C (n_28976), .D (n_30023),.Y (n_30933));
OR4X1 g106511(.A (n_29004), .B (n_20754), .C (n_29006), .D (n_29998),.Y (n_30932));
OAI21X1 g106514(.A0 (n_30085), .A1 (n_31482), .B0 (n_9916), .Y(n_30931));
NAND4X1 g106517(.A (n_32908), .B (n_32909), .C (n_29957), .D(n_29166), .Y (n_30930));
OAI21X1 g105979(.A0 (n_9769), .A1 (n_31129), .B0 (n_30385), .Y(n_30929));
NAND2X1 g105995(.A (n_31933), .B (n_35619), .Y (n_35644));
OAI21X1 g105998(.A0 (n_8567), .A1 (n_31734), .B0 (n_30419), .Y(n_30927));
AOI21X1 g106002(.A0 (n_30232), .A1 (n_21313), .B0 (n_8070), .Y(n_30926));
CLKBUFX1 gbuf_d_306(.A(n_30428), .Y(d_out_306));
CLKBUFX1 gbuf_q_306(.A(q_in_306), .Y(n_13361));
AOI21X1 g106599(.A0 (n_10394), .A1 (n_30311), .B0 (n_16415), .Y(n_30924));
NAND4X1 g106610(.A (n_35088), .B (n_9133), .C (n_29904), .D(n_35089), .Y (n_30921));
OAI21X1 g106017(.A0 (n_8565), .A1 (n_31734), .B0 (n_30404), .Y(n_30919));
AOI21X1 g106619(.A0 (n_30037), .A1 (n_30274), .B0 (n_31233), .Y(n_30917));
AOI21X1 g106624(.A0 (n_30036), .A1 (n_30273), .B0 (n_31233), .Y(n_30916));
OAI21X1 g106646(.A0 (n_30039), .A1 (n_29942), .B0 (n_30914), .Y(n_30915));
OAI21X1 g107951(.A0 (n_29712), .A1 (n_30523), .B0 (n_21205), .Y(n_30913));
OAI21X1 g106651(.A0 (n_30038), .A1 (n_29940), .B0 (n_35008), .Y(n_30912));
OAI21X1 g106654(.A0 (n_30286), .A1 (n_29641), .B0 (n_31064), .Y(n_30910));
NAND3X1 g106656(.A (n_30057), .B (n_30028), .C (n_30003), .Y(n_30909));
NOR2X1 g106658(.A (n_25672), .B (n_30363), .Y (n_30908));
NAND2X1 g106659(.A (n_30352), .B (n_12875), .Y (n_30907));
NAND2X1 g106671(.A (n_30349), .B (n_13187), .Y (n_30906));
INVX1 g106047(.A (n_30733), .Y (n_30905));
NAND4X1 g106676(.A (n_30282), .B (n_29840), .C (n_29849), .D(n_29435), .Y (n_30904));
NOR2X1 g106679(.A (n_30417), .B (n_30368), .Y (n_30903));
OAI21X1 g106681(.A0 (n_30277), .A1 (n_29938), .B0 (n_30569), .Y(n_30902));
NOR2X1 g106684(.A (n_25719), .B (n_30348), .Y (n_30901));
NAND3X1 g106687(.A (n_30322), .B (n_22089), .C (n_30318), .Y(n_30900));
NOR2X1 g106688(.A (n_29941), .B (n_30424), .Y (n_30899));
NAND3X1 g106690(.A (n_8947), .B (n_30307), .C (n_30897), .Y(n_30898));
NAND3X1 g106694(.A (n_9604), .B (n_29612), .C (n_30323), .Y(n_30896));
OAI21X1 g108055(.A0 (n_27847), .A1 (n_8664), .B0 (n_30433), .Y(n_30895));
OAI21X1 g106698(.A0 (n_8821), .A1 (n_30893), .B0 (n_30354), .Y(n_30894));
NOR2X1 g106711(.A (n_9186), .B (n_30413), .Y (n_30891));
OAI21X1 g106717(.A0 (n_30267), .A1 (n_31620), .B0 (n_10441), .Y(n_30890));
NOR2X1 g106721(.A (n_10427), .B (n_30411), .Y (n_30889));
NOR2X1 g106723(.A (n_9893), .B (n_30410), .Y (n_30888));
OAI21X1 g106724(.A0 (n_9851), .A1 (n_30886), .B0 (n_30409), .Y(n_30887));
AOI21X1 g106729(.A0 (n_30171), .A1 (n_30837), .B0 (n_29723), .Y(n_30885));
OAI21X1 g106731(.A0 (n_9873), .A1 (n_30886), .B0 (n_30366), .Y(n_30884));
OAI21X1 g106732(.A0 (n_9876), .A1 (n_31299), .B0 (n_30365), .Y(n_30883));
AOI22X1 g106733(.A0 (n_30272), .A1 (n_31398), .B0 (n_8246), .B1(n_30881), .Y (n_30882));
AOI21X1 g106735(.A0 (n_30171), .A1 (n_35307), .B0 (n_29726), .Y(n_30880));
OAI21X1 g106736(.A0 (n_8823), .A1 (n_30893), .B0 (n_30350), .Y(n_30879));
NAND4X1 g106737(.A (n_32213), .B (n_32214), .C (n_28560), .D(n_28541), .Y (n_30878));
NAND4X1 g106741(.A (n_35408), .B (n_22090), .C (n_29894), .D(n_35409), .Y (n_30876));
AOI22X1 g106743(.A0 (n_30874), .A1 (n_30668), .B0 (n_32340), .B1(n_33785), .Y (n_30875));
NOR2X1 g106745(.A (n_30542), .B (n_30351), .Y (n_30873));
NOR2X1 g106750(.A (n_30418), .B (n_30054), .Y (n_30870));
AOI22X1 g106754(.A0 (n_30842), .A1 (n_30180), .B0 (n_20692), .B1(n_22123), .Y (n_30869));
OAI21X1 g106755(.A0 (n_30253), .A1 (n_29388), .B0 (n_20734), .Y(n_30868));
NOR2X1 g106756(.A (n_29650), .B (n_30383), .Y (n_30867));
AOI22X1 g106761(.A0 (n_30268), .A1 (n_31878), .B0 (n_9371), .B1(n_31819), .Y (n_30866));
NOR2X1 g106765(.A (n_9906), .B (n_30406), .Y (n_30865));
NOR2X1 g106767(.A (n_10354), .B (n_30405), .Y (n_30864));
AOI22X1 g106770(.A0 (n_30860), .A1 (n_33738), .B0 (n_20136), .B1(n_30505), .Y (n_32067));
NOR2X1 g106771(.A (n_7083), .B (n_30425), .Y (n_30862));
AOI21X1 g106773(.A0 (n_30860), .A1 (n_28158), .B0 (n_15408), .Y(n_32066));
NOR2X1 g106774(.A (n_7191), .B (n_30427), .Y (n_30859));
AOI21X1 g106775(.A0 (n_30834), .A1 (n_29155), .B0 (n_15410), .Y(n_30858));
OAI21X1 g106776(.A0 (n_33800), .A1 (n_9493), .B0 (n_30090), .Y(n_30857));
AOI21X1 g106777(.A0 (n_30641), .A1 (n_28158), .B0 (n_15416), .Y(n_30856));
CLKBUFX1 gbuf_d_307(.A(n_30432), .Y(d_out_307));
CLKBUFX1 gbuf_q_307(.A(q_in_307), .Y(n_3470));
CLKBUFX1 gbuf_d_308(.A(n_30430), .Y(d_out_308));
CLKBUFX1 gbuf_q_308(.A(q_in_308), .Y(P3_reg1[7]));
CLKBUFX1 gbuf_d_309(.A(n_30345), .Y(d_out_309));
CLKBUFX1 gbuf_q_309(.A(q_in_309), .Y(n_4237));
CLKBUFX1 gbuf_d_310(.A(n_30346), .Y(d_out_310));
CLKBUFX1 gbuf_q_310(.A(q_in_310), .Y(n_9595));
CLKBUFX1 gbuf_d_311(.A(n_30390), .Y(d_out_311));
CLKBUFX1 gbuf_q_311(.A(q_in_311), .Y(n_10854));
NAND4X1 g106786(.A (n_29630), .B (n_10603), .C (n_29901), .D(n_29605), .Y (n_30854));
AOI22X1 g106787(.A0 (n_30675), .A1 (n_33494), .B0 (n_34774), .B1(n_28926), .Y (n_30853));
AOI21X1 g106795(.A0 (n_30839), .A1 (n_29341), .B0 (n_30378), .Y(n_30851));
AOI21X1 g106797(.A0 (n_35307), .A1 (n_30836), .B0 (n_20105), .Y(n_30850));
NAND2X1 g106799(.A (n_6945), .B (n_30423), .Y (n_30848));
NAND2X1 g106814(.A (n_6537), .B (n_30422), .Y (n_30847));
OAI21X1 g106816(.A0 (n_30264), .A1 (n_31541), .B0 (n_6927), .Y(n_30846));
AOI22X1 g106830(.A0 (n_33546), .A1 (n_30842), .B0 (n_29906), .B1(n_28926), .Y (n_30844));
OAI21X1 g106831(.A0 (n_29972), .A1 (n_10790), .B0 (n_30412), .Y(n_30841));
AOI21X1 g106832(.A0 (n_30839), .A1 (n_29430), .B0 (n_30376), .Y(n_30840));
AOI21X1 g106833(.A0 (n_30837), .A1 (n_30836), .B0 (n_20130), .Y(n_30838));
AOI21X1 g106834(.A0 (n_30834), .A1 (n_29253), .B0 (n_30541), .Y(n_30835));
NAND2X1 g106869(.A (n_30528), .B (n_31205), .Y (n_30833));
NAND2X1 g106870(.A (n_30526), .B (n_31912), .Y (n_30832));
NAND4X1 g106876(.A (n_35107), .B (n_9176), .C (n_35108), .D(n_28654), .Y (n_30831));
NAND4X1 g106879(.A (n_32119), .B (n_9105), .C (n_32120), .D(n_28652), .Y (n_30830));
NOR2X1 g106889(.A (n_30502), .B (n_30529), .Y (n_30829));
NOR2X1 g106891(.A (n_30501), .B (n_30525), .Y (n_30828));
NOR2X1 g106892(.A (n_30500), .B (n_30520), .Y (n_30827));
NAND4X1 g106894(.A (n_29759), .B (n_14812), .C (n_35147), .D(n_35148), .Y (n_30826));
NAND3X1 g106895(.A (n_10859), .B (n_29911), .C (n_30195), .Y(n_30825));
AOI21X1 g106906(.A0 (n_30175), .A1 (n_29314), .B0 (n_8340), .Y(n_30824));
AOI21X1 g106916(.A0 (n_30143), .A1 (n_27935), .B0 (n_33125), .Y(n_30823));
CLKBUFX1 gbuf_d_312(.A(n_30431), .Y(d_out_312));
CLKBUFX1 gbuf_q_312(.A(q_in_312), .Y(n_3693));
NAND2X1 g106945(.A (n_33801), .B (n_30399), .Y (n_32133));
NAND2X1 g106946(.A (n_33801), .B (n_33513), .Y (n_30820));
NAND4X1 g106190(.A (n_30443), .B (n_15414), .C (n_29718), .D(n_29252), .Y (n_30819));
OAI21X1 g106195(.A0 (n_8568), .A1 (n_30811), .B0 (n_30521), .Y(n_30818));
OAI21X1 g106967(.A0 (n_30162), .A1 (n_29461), .B0 (n_31544), .Y(n_30817));
NOR2X1 g106975(.A (n_30524), .B (n_30515), .Y (n_30816));
NOR2X1 g106976(.A (n_30507), .B (n_30522), .Y (n_30815));
NOR2X1 g106992(.A (n_29750), .B (n_30327), .Y (n_30814));
NAND3X1 g107007(.A (n_32598), .B (n_32599), .C (n_32144), .Y(n_30813));
OAI21X1 g106217(.A0 (n_8256), .A1 (n_30811), .B0 (n_30539), .Y(n_30812));
NAND3X1 g107025(.A (n_32913), .B (n_32914), .C (n_29758), .Y(n_30810));
NAND3X1 g107034(.A (n_35449), .B (n_35450), .C (n_29851), .Y(n_30809));
OAI21X1 g106231(.A0 (n_8572), .A1 (n_30811), .B0 (n_30535), .Y(n_30808));
NOR2X1 g107057(.A (n_9932), .B (n_30555), .Y (n_30807));
NOR2X1 g107061(.A (n_9096), .B (n_30504), .Y (n_32260));
OAI21X1 g107095(.A0 (n_30149), .A1 (n_30619), .B0 (n_8601), .Y(n_30805));
NOR2X1 g107098(.A (n_8887), .B (n_30329), .Y (n_30804));
NOR2X1 g107104(.A (n_9903), .B (n_30538), .Y (n_30803));
NAND4X1 g107110(.A (n_30452), .B (n_15003), .C (n_28990), .D(n_9047), .Y (n_30801));
NAND3X1 g107112(.A (n_30150), .B (n_30142), .C (n_15112), .Y(n_30800));
NOR2X1 g107117(.A (n_30332), .B (n_30518), .Y (n_30799));
AOI21X1 g107126(.A0 (n_30566), .A1 (n_34952), .B0 (n_15490), .Y(n_32570));
NAND4X1 g107145(.A (n_28661), .B (n_19475), .C (n_29794), .D(n_28648), .Y (n_30795));
NAND4X1 g107156(.A (n_28663), .B (n_10083), .C (n_29796), .D(n_28650), .Y (n_30794));
OAI21X1 g106289(.A0 (n_30130), .A1 (n_30792), .B0 (n_6566), .Y(n_30793));
OAI21X1 g106297(.A0 (n_30121), .A1 (n_31273), .B0 (n_6598), .Y(n_30791));
OAI21X1 g107172(.A0 (n_30159), .A1 (n_31538), .B0 (n_6987), .Y(n_30790));
NAND2X1 g107178(.A (n_6651), .B (n_30335), .Y (n_30789));
OAI21X1 g107182(.A0 (n_30151), .A1 (n_31538), .B0 (n_6842), .Y(n_30788));
NOR2X1 g107233(.A (n_30446), .B (n_30465), .Y (n_30787));
NOR2X1 g107235(.A (n_30444), .B (n_30461), .Y (n_30786));
AOI21X1 g106339(.A0 (n_10489), .A1 (n_30046), .B0 (n_31586), .Y(n_30785));
AOI21X1 g106345(.A0 (n_9390), .A1 (n_30097), .B0 (n_30783), .Y(n_30784));
NAND3X1 g107303(.A (n_29458), .B (n_29755), .C (n_29391), .Y(n_30782));
NAND4X1 g106375(.A (n_30071), .B (n_15263), .C (n_28739), .D(n_22111), .Y (n_30781));
NAND3X1 g107353(.A (n_35927), .B (n_29746), .C (n_35928), .Y(n_30780));
NAND3X1 g107354(.A (n_32611), .B (n_29745), .C (n_32612), .Y(n_30779));
NAND2X1 g107365(.A (n_30146), .B (n_29753), .Y (n_30778));
NOR2X1 g107373(.A (n_25066), .B (n_30140), .Y (n_30777));
NAND3X1 g107386(.A (n_7778), .B (n_29793), .C (n_6878), .Y (n_30776));
NOR2X1 g107398(.A (n_9936), .B (n_30196), .Y (n_30775));
AOI22X1 g107402(.A0 (n_35248), .A1 (n_30063), .B0 (n_9629), .B1(n_21251), .Y (n_30774));
NAND4X1 g106413(.A (n_35703), .B (n_29248), .C (n_35704), .D(n_35298), .Y (n_30773));
NOR3X1 g106422(.A (n_28628), .B (n_25863), .C (n_29722), .Y(n_30772));
NOR2X1 g107431(.A (n_9040), .B (n_30137), .Y (n_30771));
NAND2X1 g107438(.A (n_30173), .B (n_29129), .Y (n_30770));
NAND2X1 g107439(.A (n_30172), .B (n_29484), .Y (n_30769));
NOR2X1 g107442(.A (n_9927), .B (n_30170), .Y (n_30768));
OAI21X1 g106431(.A0 (n_30462), .A1 (n_12670), .B0 (n_30180), .Y(n_30767));
OAI21X1 g107443(.A0 (n_29747), .A1 (n_28397), .B0 (n_31878), .Y(n_30766));
NAND2X1 g106434(.A (n_30118), .B (n_12732), .Y (n_30765));
NOR2X1 g107456(.A (n_30226), .B (n_29861), .Y (n_30764));
OAI21X1 g107462(.A0 (n_18298), .A1 (n_21365), .B0 (n_30181), .Y(n_30762));
OAI21X1 g107463(.A0 (n_18295), .A1 (n_21365), .B0 (n_30164), .Y(n_30761));
NOR2X1 g106443(.A (n_29656), .B (n_30157), .Y (n_30759));
NAND4X1 g106462(.A (n_30052), .B (n_15266), .C (n_29234), .D(n_28707), .Y (n_30757));
NOR2X1 g106463(.A (n_34776), .B (n_28665), .Y (n_30755));
NOR2X1 g106465(.A (n_35326), .B (n_35325), .Y (n_30754));
NAND2X1 g107525(.A (n_29920), .B (n_30179), .Y (n_30753));
NAND2X1 g107529(.A (n_29916), .B (n_30163), .Y (n_30752));
AOI21X1 g105947(.A0 (n_8372), .A1 (n_29997), .B0 (n_30702), .Y(n_30751));
NOR3X1 g106494(.A (n_28619), .B (n_25844), .C (n_33339), .Y(n_30750));
OAI21X1 g106542(.A0 (n_30462), .A1 (n_8940), .B0 (n_28517), .Y(n_30748));
AOI21X1 g106585(.A0 (n_9418), .A1 (n_29709), .B0 (n_30783), .Y(n_30747));
OAI21X1 g107853(.A0 (n_29740), .A1 (n_28867), .B0 (n_31064), .Y(n_30746));
NAND3X1 g106016(.A (n_12426), .B (n_26486), .C (n_29945), .Y(n_30745));
NOR2X1 g106630(.A (n_9911), .B (n_30058), .Y (n_30744));
OAI21X1 g106632(.A0 (n_8820), .A1 (n_35012), .B0 (n_30056), .Y(n_30743));
NAND4X1 g106640(.A (n_15271), .B (n_29161), .C (n_29160), .D(n_29586), .Y (n_30742));
NAND4X1 g106641(.A (n_15175), .B (n_29534), .C (n_29533), .D(n_29580), .Y (n_30741));
NAND4X1 g106643(.A (n_15096), .B (n_29157), .C (n_29560), .D(n_29159), .Y (n_30740));
NAND4X1 g106644(.A (n_15017), .B (n_29527), .C (n_29559), .D(n_29532), .Y (n_30739));
NAND2X1 g106649(.A (n_30065), .B (n_31641), .Y (n_30738));
NAND3X1 g107968(.A (n_29732), .B (n_29733), .C (n_29717), .Y(n_30737));
NAND4X1 g107980(.A (n_29313), .B (n_29716), .C (n_29228), .D(n_28761), .Y (n_30736));
NAND2X1 g106667(.A (n_30053), .B (n_31201), .Y (n_30735));
NAND2X1 g107988(.A (n_30111), .B (n_29344), .Y (n_30734));
NAND4X1 g106048(.A (n_32879), .B (n_29692), .C (n_32880), .D(n_27043), .Y (n_30733));
OAI21X1 g106697(.A0 (n_8798), .A1 (n_30731), .B0 (n_30045), .Y(n_30732));
OAI21X1 g106705(.A0 (n_8832), .A1 (n_35012), .B0 (n_30044), .Y(n_30730));
AOI22X1 g106706(.A0 (n_29991), .A1 (n_35008), .B0 (n_9225), .B1(n_34706), .Y (n_30729));
OAI21X1 g106719(.A0 (n_9861), .A1 (n_30886), .B0 (n_30103), .Y(n_30728));
NOR2X1 g108145(.A (n_30325), .B (n_28859), .Y (n_30727));
AOI22X1 g106753(.A0 (n_35042), .A1 (n_33802), .B0 (n_19496), .B1(n_33803), .Y (n_30726));
OAI21X1 g106758(.A0 (n_8266), .A1 (n_31199), .B0 (n_30070), .Y(n_30723));
AOI22X1 g106759(.A0 (n_29994), .A1 (n_31398), .B0 (n_8024), .B1(n_30881), .Y (n_30722));
NOR2X1 g106092(.A (n_29786), .B (n_30098), .Y (n_30721));
NAND2X1 g106762(.A (n_30096), .B (n_15404), .Y (n_30720));
AOI22X1 g106763(.A0 (n_29983), .A1 (n_31878), .B0 (n_9428), .B1(n_31819), .Y (n_30719));
NOR2X1 g106772(.A (n_7033), .B (n_30106), .Y (n_30718));
CLKBUFX1 gbuf_d_313(.A(n_30049), .Y(d_out_313));
CLKBUFX1 gbuf_q_313(.A(q_in_313), .Y(n_3333));
CLKBUFX1 gbuf_d_314(.A(n_30242), .Y(d_out_314));
CLKBUFX1 gbuf_q_314(.A(q_in_314), .Y(n_3337));
CLKBUFX1 gbuf_d_315(.A(n_30241), .Y(d_out_315));
CLKBUFX1 gbuf_q_315(.A(q_in_315), .Y(n_9597));
CLKBUFX1 gbuf_d_316(.A(n_30240), .Y(d_out_316));
CLKBUFX1 gbuf_q_316(.A(q_in_316), .Y(P2_reg1[6]));
CLKBUFX1 gbuf_d_317(.A(n_30238), .Y(d_out_317));
CLKBUFX1 gbuf_q_317(.A(q_in_317), .Y(n_3259));
CLKBUFX1 gbuf_d_318(.A(n_30237), .Y(d_out_318));
CLKBUFX1 gbuf_q_318(.A(q_in_318), .Y(n_10148));
CLKBUFX1 gbuf_d_319(.A(n_30134), .Y(d_out_319));
CLKBUFX1 gbuf_q_319(.A(q_in_319), .Y(n_13209));
NOR2X1 g106780(.A (n_7079), .B (n_30107), .Y (n_30717));
NAND2X1 g106800(.A (n_6692), .B (n_30062), .Y (n_30716));
NAND2X1 g106803(.A (n_6743), .B (n_30059), .Y (n_30715));
NAND2X1 g106808(.A (n_6641), .B (n_30104), .Y (n_30714));
OAI21X1 g106810(.A0 (n_30377), .A1 (n_28528), .B0 (n_19563), .Y(n_30713));
OAI21X1 g106817(.A0 (n_29982), .A1 (n_31605), .B0 (n_6618), .Y(n_30712));
OAI21X1 g106818(.A0 (n_29981), .A1 (n_31605), .B0 (n_6619), .Y(n_30711));
NAND2X1 g106822(.A (n_30066), .B (n_19551), .Y (n_30709));
OAI21X1 g106823(.A0 (n_29967), .A1 (n_31605), .B0 (n_6568), .Y(n_30708));
OAI21X1 g106824(.A0 (n_29966), .A1 (n_30792), .B0 (n_6605), .Y(n_30707));
NAND2X1 g106826(.A (n_6503), .B (n_30081), .Y (n_30706));
NAND2X1 g106144(.A (n_30219), .B (n_31891), .Y (n_30705));
NAND2X1 g106146(.A (n_30218), .B (n_31092), .Y (n_30704));
AOI21X1 g106854(.A0 (n_9422), .A1 (n_29892), .B0 (n_30702), .Y(n_30703));
AOI21X1 g106855(.A0 (n_9421), .A1 (n_29891), .B0 (n_30702), .Y(n_30701));
NAND4X1 g106861(.A (n_29683), .B (n_10172), .C (n_29433), .D(n_28909), .Y (n_30700));
NAND4X1 g106862(.A (n_30283), .B (n_10168), .C (n_29423), .D(n_28906), .Y (n_30699));
NOR2X1 g106864(.A (n_30034), .B (n_29364), .Y (n_30698));
NOR2X1 g106865(.A (n_30033), .B (n_29363), .Y (n_30697));
NAND2X1 g106871(.A (n_30266), .B (n_31260), .Y (n_30696));
NAND2X1 g106872(.A (n_30265), .B (n_30421), .Y (n_30695));
NAND2X1 g106874(.A (n_30254), .B (n_31781), .Y (n_30694));
NOR2X1 g106877(.A (n_24685), .B (n_30271), .Y (n_32265));
OAI21X1 g106159(.A0 (n_8274), .A1 (n_30691), .B0 (n_30269), .Y(n_30692));
NOR2X1 g106880(.A (n_24674), .B (n_30270), .Y (n_35080));
NAND2X1 g106884(.A (n_30255), .B (n_31850), .Y (n_30689));
OAI21X1 g106899(.A0 (n_29888), .A1 (n_27949), .B0 (n_33123), .Y(n_30687));
OAI21X1 g106901(.A0 (n_29887), .A1 (n_28886), .B0 (n_33123), .Y(n_30686));
NAND2X1 g106175(.A (n_30217), .B (n_13091), .Y (n_30685));
OAI21X1 g106920(.A0 (n_29852), .A1 (n_25572), .B0 (n_30683), .Y(n_30684));
OAI21X1 g106178(.A0 (n_8257), .A1 (n_30691), .B0 (n_30258), .Y(n_30682));
NAND2X1 g106923(.A (n_30839), .B (n_8922), .Y (n_30681));
NAND2X1 g106925(.A (n_35308), .B (n_30291), .Y (n_32145));
NAND2X1 g106928(.A (n_30200), .B (n_30860), .Y (n_30679));
NAND4X1 g106937(.A (n_15250), .B (n_29406), .C (n_29404), .D(n_29431), .Y (n_30678));
NAND2X1 g106942(.A (n_30675), .B (n_30184), .Y (n_30676));
NAND2X1 g106943(.A (n_30675), .B (n_26611), .Y (n_30674));
NAND2X1 g106944(.A (n_30675), .B (n_30180), .Y (n_30673));
NAND2X1 g106956(.A (n_33129), .B (n_30668), .Y (n_30669));
NAND4X1 g106965(.A (n_27298), .B (n_25865), .C (n_29462), .D(n_28829), .Y (n_30667));
NAND4X1 g106973(.A (n_32275), .B (n_32276), .C (n_29465), .D(n_28825), .Y (n_30666));
OAI21X1 g106200(.A0 (n_8716), .A1 (n_31422), .B0 (n_30235), .Y(n_30665));
NOR2X1 g106974(.A (n_25845), .B (n_30281), .Y (n_30664));
NAND3X1 g106987(.A (n_29863), .B (n_29836), .C (n_15186), .Y(n_30662));
NAND3X1 g106990(.A (n_29862), .B (n_29835), .C (n_15273), .Y(n_30661));
NAND2X1 g106991(.A (n_30842), .B (n_30559), .Y (n_30660));
OAI21X1 g106206(.A0 (n_8777), .A1 (n_31422), .B0 (n_30234), .Y(n_30659));
NOR2X1 g106994(.A (n_29326), .B (n_30025), .Y (n_30658));
OAI21X1 g106207(.A0 (n_8582), .A1 (n_30811), .B0 (n_30301), .Y(n_30657));
NAND2X1 g106997(.A (n_30248), .B (n_27522), .Y (n_30656));
NAND2X1 g107002(.A (n_30645), .B (n_8954), .Y (n_30655));
NAND2X1 g107003(.A (n_30837), .B (n_29684), .Y (n_32606));
NAND3X1 g107006(.A (n_32152), .B (n_29569), .C (n_32153), .Y(n_30653));
NOR2X1 g106213(.A (n_8901), .B (n_30300), .Y (n_30652));
NAND2X1 g107009(.A (n_30860), .B (n_26238), .Y (n_30651));
NAND3X1 g107011(.A (n_30262), .B (n_29616), .C (n_29875), .Y(n_30650));
OAI21X1 g107013(.A0 (n_29869), .A1 (n_28044), .B0 (n_30380), .Y(n_30649));
NAND3X1 g107015(.A (n_28079), .B (n_29900), .C (n_29373), .Y(n_30648));
NOR2X1 g107016(.A (n_25323), .B (n_30260), .Y (n_30647));
NAND2X1 g107018(.A (n_30645), .B (n_30636), .Y (n_30646));
NAND2X1 g107019(.A (n_30645), .B (n_29405), .Y (n_30644));
NAND4X1 g107026(.A (n_29829), .B (n_29421), .C (n_29419), .D(n_20733), .Y (n_30643));
NAND2X1 g107028(.A (n_30641), .B (n_28136), .Y (n_30642));
NOR2X1 g107030(.A (n_25868), .B (n_30247), .Y (n_30640));
NOR2X1 g107031(.A (n_25365), .B (n_30246), .Y (n_30639));
NAND2X1 g107033(.A (n_30641), .B (n_8954), .Y (n_30638));
NAND2X1 g107035(.A (n_30641), .B (n_30636), .Y (n_30637));
NAND2X1 g107036(.A (n_29962), .B (n_27902), .Y (n_30635));
NAND2X1 g107043(.A (n_30834), .B (n_33738), .Y (n_30634));
NOR2X1 g106229(.A (n_9377), .B (n_30285), .Y (n_30632));
OAI21X1 g107046(.A0 (n_27069), .A1 (n_8678), .B0 (n_30309), .Y(n_30631));
NAND4X1 g107049(.A (n_35095), .B (n_35096), .C (n_29399), .D(n_25419), .Y (n_30630));
NAND3X1 g107054(.A (n_28080), .B (n_29872), .C (n_29330), .Y(n_30629));
NAND4X1 g107058(.A (n_32070), .B (n_32071), .C (n_29395), .D(n_24246), .Y (n_30628));
NAND4X1 g107060(.A (n_35633), .B (n_35634), .C (n_29394), .D(n_25411), .Y (n_30627));
OAI21X1 g107062(.A0 (n_32409), .A1 (n_8285), .B0 (n_22088), .Y(n_30626));
AOI21X1 g107065(.A0 (n_30594), .A1 (n_30180), .B0 (n_21726), .Y(n_32028));
AOI22X1 g107068(.A0 (n_29870), .A1 (n_35008), .B0 (n_9295), .B1(n_34706), .Y (n_30624));
OAI21X1 g107069(.A0 (n_29902), .A1 (n_28789), .B0 (n_30914), .Y(n_30623));
NOR2X1 g107074(.A (n_8906), .B (n_30030), .Y (n_30622));
OAI21X1 g107079(.A0 (n_29899), .A1 (n_27777), .B0 (n_30360), .Y(n_30621));
OAI21X1 g107082(.A0 (n_29867), .A1 (n_30619), .B0 (n_8392), .Y(n_30620));
OAI21X1 g107093(.A0 (n_29856), .A1 (n_30619), .B0 (n_8606), .Y(n_30617));
NOR2X1 g106259(.A (n_7020), .B (n_30029), .Y (n_30616));
OAI21X1 g107102(.A0 (n_8787), .A1 (n_31131), .B0 (n_30294), .Y(n_30615));
NAND4X1 g107106(.A (n_28786), .B (n_27390), .C (n_29379), .D(n_24202), .Y (n_30614));
NAND3X1 g107111(.A (n_35908), .B (n_35909), .C (n_15071), .Y(n_30613));
NAND2X1 g106267(.A (n_6638), .B (n_30319), .Y (n_30612));
OAI21X1 g107127(.A0 (n_8023), .A1 (n_31199), .B0 (n_30278), .Y(n_30611));
NAND2X1 g106274(.A (n_6625), .B (n_30317), .Y (n_30610));
OAI21X1 g107128(.A0 (n_8597), .A1 (n_31713), .B0 (n_30279), .Y(n_35648));
NAND2X1 g106277(.A (n_6875), .B (n_30316), .Y (n_30608));
NAND2X1 g106279(.A (n_6657), .B (n_30315), .Y (n_30606));
OAI21X1 g107137(.A0 (n_30145), .A1 (n_33340), .B0 (n_30018), .Y(n_30605));
OAI21X1 g107138(.A0 (n_34963), .A1 (n_33340), .B0 (n_30012), .Y(n_30604));
NAND2X1 g107140(.A (n_30296), .B (n_8316), .Y (n_30601));
NAND2X1 g107144(.A (n_30287), .B (n_20137), .Y (n_30600));
OAI21X1 g107147(.A0 (n_29871), .A1 (n_27792), .B0 (n_30353), .Y(n_30599));
NOR2X1 g107149(.A (n_7017), .B (n_30041), .Y (n_30598));
OAI21X1 g107154(.A0 (n_29855), .A1 (n_27746), .B0 (n_30914), .Y(n_30597));
OAI21X1 g107159(.A0 (n_32409), .A1 (n_30138), .B0 (n_29607), .Y(n_30596));
AOI22X1 g107160(.A0 (n_30594), .A1 (n_30668), .B0 (n_30589), .B1(n_33785), .Y (n_30595));
NAND2X1 g107164(.A (n_29625), .B (n_30320), .Y (n_30591));
AOI22X1 g107165(.A0 (n_30594), .A1 (n_33494), .B0 (n_30589), .B1(n_28926), .Y (n_30590));
OAI21X1 g107171(.A0 (n_29832), .A1 (n_8352), .B0 (n_20108), .Y(n_30586));
NAND2X1 g107177(.A (n_6563), .B (n_30035), .Y (n_30585));
NAND4X1 g107180(.A (n_7131), .B (n_6878), .C (n_7552), .D (n_29470),.Y (n_30584));
OAI21X1 g107184(.A0 (n_32409), .A1 (n_30445), .B0 (n_29622), .Y(n_30583));
NOR2X1 g107210(.A (n_29811), .B (n_30153), .Y (n_30582));
NOR2X1 g107211(.A (n_29810), .B (n_30152), .Y (n_30581));
NOR2X1 g107212(.A (n_29809), .B (n_30148), .Y (n_30580));
NOR2X1 g107213(.A (n_29808), .B (n_30147), .Y (n_30579));
CLKBUFX1 gbuf_d_320(.A(n_30192), .Y(d_out_320));
CLKBUFX1 gbuf_q_320(.A(q_in_320), .Y(n_10144));
NOR2X1 g107222(.A (n_30229), .B (n_29278), .Y (n_30578));
NOR3X1 g107223(.A (n_29277), .B (n_24676), .C (n_29787), .Y(n_30577));
NAND3X1 g107238(.A (n_11121), .B (n_29736), .C (n_29446), .Y(n_30576));
AOI21X1 g107241(.A0 (n_29816), .A1 (n_29311), .B0 (n_8070), .Y(n_30575));
AOI21X1 g107242(.A0 (n_29815), .A1 (n_29310), .B0 (n_8070), .Y(n_30573));
AOI21X1 g107245(.A0 (n_29814), .A1 (n_29309), .B0 (n_31178), .Y(n_30572));
NOR2X1 g107247(.A (n_29343), .B (n_30169), .Y (n_30571));
OAI21X1 g107251(.A0 (n_29789), .A1 (n_28953), .B0 (n_30569), .Y(n_30570));
AOI21X1 g106341(.A0 (n_10460), .A1 (n_29763), .B0 (n_31388), .Y(n_30568));
NAND2X1 g107254(.A (n_30566), .B (n_30563), .Y (n_30567));
NAND2X1 g107255(.A (n_34950), .B (n_30563), .Y (n_30565));
NAND4X1 g107266(.A (n_32273), .B (n_28345), .C (n_28875), .D(n_32274), .Y (n_30562));
NAND2X1 g107269(.A (n_33503), .B (n_30559), .Y (n_30561));
AOI21X1 g107283(.A0 (n_29447), .A1 (n_29451), .B0 (n_31236), .Y(n_30555));
NAND2X1 g107288(.A (n_30594), .B (n_26665), .Y (n_30554));
NAND4X1 g107300(.A (n_34717), .B (n_29042), .C (n_25343), .D(n_28949), .Y (n_30553));
NOR2X1 g107306(.A (n_29843), .B (n_29513), .Y (n_30552));
NAND2X1 g107311(.A (n_33541), .B (n_30559), .Y (n_30549));
NAND2X1 g107317(.A (n_33495), .B (n_30559), .Y (n_30548));
NAND2X1 g107325(.A (n_29853), .B (n_29818), .Y (n_30543));
NOR2X1 g107328(.A (n_30050), .B (n_29834), .Y (n_30542));
NOR2X1 g107334(.A (n_10002), .B (n_29833), .Y (n_30541));
NAND2X1 g107337(.A (n_29932), .B (n_28599), .Y (n_30540));
OAI21X1 g106382(.A0 (n_29589), .A1 (n_29337), .B0 (n_31628), .Y(n_30539));
AOI21X1 g107352(.A0 (n_35382), .A1 (n_35383), .B0 (n_30537), .Y(n_30538));
OAI21X1 g106390(.A0 (n_29555), .A1 (n_29331), .B0 (n_31573), .Y(n_30535));
NOR2X1 g107364(.A (n_29866), .B (n_29329), .Y (n_30534));
NOR2X1 g107367(.A (n_29930), .B (n_25562), .Y (n_30533));
AOI21X1 g107381(.A0 (n_14486), .A1 (n_30530), .B0 (n_29873), .Y(n_30531));
OAI21X1 g107394(.A0 (n_29360), .A1 (n_8321), .B0 (n_22136), .Y(n_30529));
OAI21X1 g107409(.A0 (n_8580), .A1 (n_30527), .B0 (n_29937), .Y(n_30528));
OAI21X1 g107410(.A0 (n_8578), .A1 (n_30527), .B0 (n_29936), .Y(n_30526));
OAI21X1 g107411(.A0 (n_29356), .A1 (n_8321), .B0 (n_22131), .Y(n_30525));
OAI21X1 g107412(.A0 (n_30514), .A1 (n_30523), .B0 (n_22129), .Y(n_30524));
OAI21X1 g107413(.A0 (n_29376), .A1 (n_29388), .B0 (n_22478), .Y(n_30522));
OAI21X1 g106416(.A0 (n_29543), .A1 (n_29338), .B0 (n_31628), .Y(n_30521));
OAI21X1 g107418(.A0 (n_29347), .A1 (n_29388), .B0 (n_22476), .Y(n_30520));
NAND3X1 g107422(.A (n_9077), .B (n_20120), .C (n_29409), .Y(n_30518));
OAI21X1 g106424(.A0 (n_29594), .A1 (n_29298), .B0 (n_7827), .Y(n_30517));
OAI21X1 g107445(.A0 (n_29380), .A1 (n_27827), .B0 (n_30099), .Y(n_30516));
OAI21X1 g107451(.A0 (n_30514), .A1 (n_8678), .B0 (n_29618), .Y(n_30515));
NOR2X1 g107458(.A (n_29943), .B (n_29859), .Y (n_30512));
AOI21X1 g107460(.A0 (n_30220), .A1 (n_30180), .B0 (n_19621), .Y(n_35646));
AOI21X1 g107469(.A0 (n_30454), .A1 (n_29547), .B0 (n_29880), .Y(n_32147));
OAI21X1 g107488(.A0 (n_29035), .A1 (n_34719), .B0 (n_29934), .Y(n_30507));
AOI22X1 g107498(.A0 (n_30201), .A1 (n_33738), .B0 (n_21702), .B1(n_30505), .Y (n_32148));
OAI21X1 g107517(.A0 (n_35247), .A1 (n_10276), .B0 (n_29610), .Y(n_30504));
OAI21X1 g107553(.A0 (n_30445), .A1 (n_29360), .B0 (n_29626), .Y(n_30502));
OAI21X1 g107555(.A0 (n_30445), .A1 (n_29356), .B0 (n_29621), .Y(n_30501));
OAI21X1 g107556(.A0 (n_29015), .A1 (n_10790), .B0 (n_29933), .Y(n_30500));
NOR2X1 g107572(.A (n_29290), .B (n_29788), .Y (n_30498));
NOR2X1 g107573(.A (n_29288), .B (n_29785), .Y (n_30497));
NOR2X1 g107600(.A (n_29744), .B (n_29385), .Y (n_30496));
NOR2X1 g107601(.A (n_29743), .B (n_29784), .Y (n_30495));
NOR2X1 g107603(.A (n_29742), .B (n_29382), .Y (n_30494));
NOR2X1 g107604(.A (n_29741), .B (n_29780), .Y (n_30493));
NAND3X1 g107613(.A (n_32560), .B (n_28467), .C (n_32561), .Y(n_30492));
NOR2X1 g107642(.A (n_29807), .B (n_27535), .Y (n_30491));
NOR2X1 g107643(.A (n_29806), .B (n_27532), .Y (n_32029));
NOR2X1 g107644(.A (n_29805), .B (n_27530), .Y (n_30489));
NAND2X1 g107694(.A (n_29768), .B (n_25636), .Y (n_30488));
AOI21X1 g107720(.A0 (n_29315), .A1 (n_29294), .B0 (n_31236), .Y(n_30487));
NAND2X1 g107721(.A (n_32886), .B (n_32887), .Y (n_30485));
NAND2X1 g107724(.A (n_35248), .B (n_25756), .Y (n_32261));
NAND2X1 g106556(.A (n_6980), .B (n_29885), .Y (n_30482));
NAND2X1 g107726(.A (n_35248), .B (n_26528), .Y (n_30481));
NAND2X1 g107728(.A (n_29357), .B (n_33513), .Y (n_30480));
NAND3X1 g107783(.A (n_27869), .B (n_29265), .C (n_15153), .Y(n_30476));
NOR2X1 g106591(.A (n_29782), .B (n_29135), .Y (n_30475));
NOR2X1 g106593(.A (n_29779), .B (n_29134), .Y (n_30474));
NAND4X1 g107816(.A (n_28881), .B (n_28305), .C (n_20719), .D(n_28880), .Y (n_30473));
NAND3X1 g106609(.A (n_35425), .B (n_35426), .C (n_29251), .Y(n_30472));
OAI21X1 g107848(.A0 (n_28787), .A1 (n_8927), .B0 (n_29761), .Y(n_30471));
NAND4X1 g106614(.A (n_25943), .B (n_10135), .C (n_29179), .D(n_29195), .Y (n_30470));
NAND4X1 g106616(.A (n_25886), .B (n_10162), .C (n_29193), .D(n_29200), .Y (n_30469));
NOR2X1 g107878(.A (n_29056), .B (n_29804), .Y (n_30468));
NAND2X1 g106628(.A (n_29730), .B (n_29720), .Y (n_30467));
NOR2X1 g107920(.A (n_29109), .B (n_29775), .Y (n_30466));
OAI21X1 g107921(.A0 (n_29276), .A1 (n_8321), .B0 (n_21221), .Y(n_30465));
NAND2X1 g106639(.A (n_30462), .B (n_8946), .Y (n_30463));
OAI21X1 g107935(.A0 (n_29273), .A1 (n_29150), .B0 (n_21212), .Y(n_30461));
OAI21X1 g107942(.A0 (n_30449), .A1 (n_30523), .B0 (n_20739), .Y(n_30460));
NAND3X1 g106670(.A (n_29688), .B (n_29687), .C (n_28843), .Y(n_30459));
NOR2X1 g108007(.A (n_29260), .B (n_29813), .Y (n_35078));
NAND4X1 g108016(.A (n_29803), .B (n_26011), .C (n_27606), .D(n_27616), .Y (n_30457));
NOR2X1 g106680(.A (n_29778), .B (n_29734), .Y (n_30456));
AOI21X1 g108026(.A0 (n_30454), .A1 (n_29440), .B0 (n_29790), .Y(n_30455));
NAND3X1 g106686(.A (n_29256), .B (n_29685), .C (n_29255), .Y(n_30453));
NOR2X1 g108057(.A (n_28377), .B (n_29751), .Y (n_30452));
AOI22X1 g108061(.A0 (n_30122), .A1 (n_33738), .B0 (n_20185), .B1(n_21328), .Y (n_30451));
OAI21X1 g108087(.A0 (n_30449), .A1 (n_27564), .B0 (n_28656), .Y(n_30450));
OAI21X1 g106713(.A0 (n_9841), .A1 (n_30447), .B0 (n_29776), .Y(n_30448));
OAI21X1 g108108(.A0 (n_30445), .A1 (n_29276), .B0 (n_28658), .Y(n_30446));
OAI21X1 g108111(.A0 (n_30445), .A1 (n_29273), .B0 (n_28657), .Y(n_30444));
NOR2X1 g106728(.A (n_9052), .B (n_29721), .Y (n_30443));
NOR2X1 g106730(.A (n_10351), .B (n_29770), .Y (n_30442));
NAND4X1 g106742(.A (n_29208), .B (n_20752), .C (n_29182), .D(n_29196), .Y (n_30441));
AOI21X1 g106757(.A0 (n_30438), .A1 (n_30094), .B0 (n_15345), .Y(n_30440));
AOI21X1 g106760(.A0 (n_30438), .A1 (n_32850), .B0 (n_15342), .Y(n_30439));
NOR2X1 g106768(.A (n_10348), .B (n_29765), .Y (n_30437));
AOI22X1 g106769(.A0 (n_29267), .A1 (n_31528), .B0 (n_2833), .B1(n_35007), .Y (n_30436));
CLKBUFX1 gbuf_d_321(.A(n_29791), .Y(d_out_321));
CLKBUFX1 gbuf_q_321(.A(q_in_321), .Y(n_10197));
CLKBUFX1 gbuf_d_322(.A(n_29860), .Y(d_out_322));
CLKBUFX1 gbuf_q_322(.A(q_in_322), .Y(n_1976));
CLKBUFX1 gbuf_d_323(.A(n_29737), .Y(d_out_323));
CLKBUFX1 gbuf_q_323(.A(q_in_323), .Y(P3_reg3[3]));
CLKBUFX1 gbuf_d_324(.A(n_30000), .Y(d_out_324));
CLKBUFX1 gbuf_q_324(.A(q_in_324), .Y(P3_reg3[2]));
CLKBUFX1 gbuf_d_325(.A(n_29826), .Y(d_out_325));
CLKBUFX1 gbuf_q_325(.A(q_in_325), .Y(P1_reg2[1]));
CLKBUFX1 gbuf_d_326(.A(n_29954), .Y(d_out_326));
CLKBUFX1 gbuf_q_326(.A(q_in_326), .Y(P3_reg1[4]));
CLKBUFX1 gbuf_d_327(.A(n_29825), .Y(d_out_327));
CLKBUFX1 gbuf_q_327(.A(q_in_327), .Y(n_10173));
CLKBUFX1 gbuf_d_328(.A(n_29823), .Y(d_out_328));
CLKBUFX1 gbuf_q_328(.A(q_in_328), .Y(P1_reg1[1]));
CLKBUFX1 gbuf_d_329(.A(n_29898), .Y(d_out_329));
CLKBUFX1 gbuf_q_329(.A(q_in_329), .Y(n_10566));
NAND4X1 g106785(.A (n_29209), .B (n_10887), .C (n_29189), .D(n_29198), .Y (n_30435));
NAND2X1 g108294(.A (n_29269), .B (n_26528), .Y (n_30433));
NAND2X1 g106804(.A (n_6928), .B (n_29783), .Y (n_30432));
OAI21X1 g106805(.A0 (n_29676), .A1 (n_31726), .B0 (n_7055), .Y(n_30431));
OAI21X1 g106819(.A0 (n_29673), .A1 (n_31605), .B0 (n_6548), .Y(n_30430));
NOR2X1 g108368(.A (n_29724), .B (n_27176), .Y (n_30429));
OAI21X1 g106825(.A0 (n_29664), .A1 (n_30792), .B0 (n_6518), .Y(n_30428));
AOI21X1 g106856(.A0 (n_10459), .A1 (n_29632), .B0 (n_349), .Y(n_30427));
AOI21X1 g106859(.A0 (n_10389), .A1 (n_29634), .B0 (n_7058), .Y(n_30425));
NAND4X1 g106863(.A (n_29028), .B (n_25011), .C (n_28997), .D(n_9607), .Y (n_30424));
NAND2X1 g106867(.A (n_29995), .B (n_31891), .Y (n_30423));
NAND2X1 g106873(.A (n_29984), .B (n_30421), .Y (n_30422));
NAND2X1 g108475(.A (n_29727), .B (n_28320), .Y (n_30420));
OAI21X1 g106160(.A0 (n_29516), .A1 (n_21322), .B0 (n_31771), .Y(n_30419));
NAND3X1 g106885(.A (n_29507), .B (n_29584), .C (n_29164), .Y(n_30418));
NAND3X1 g106886(.A (n_29506), .B (n_29577), .C (n_29539), .Y(n_30417));
NOR2X1 g106888(.A (n_29952), .B (n_29996), .Y (n_30416));
NOR2X1 g106890(.A (n_29951), .B (n_29993), .Y (n_30415));
NOR2X1 g106893(.A (n_29950), .B (n_29986), .Y (n_30414));
AOI21X1 g106896(.A0 (n_29654), .A1 (n_28958), .B0 (n_31041), .Y(n_30413));
NAND2X1 g106902(.A (n_33546), .B (n_30386), .Y (n_30412));
AOI21X1 g106905(.A0 (n_29571), .A1 (n_28519), .B0 (n_29769), .Y(n_30411));
AOI21X1 g106907(.A0 (n_29570), .A1 (n_28518), .B0 (n_33125), .Y(n_30410));
OAI21X1 g106908(.A0 (n_29643), .A1 (n_28671), .B0 (n_24695), .Y(n_30409));
OAI21X1 g106910(.A0 (n_29540), .A1 (n_26946), .B0 (n_30683), .Y(n_30408));
NAND2X1 g106912(.A (n_29978), .B (n_29960), .Y (n_30407));
AOI21X1 g106915(.A0 (n_29496), .A1 (n_26948), .B0 (n_8340), .Y(n_30406));
AOI21X1 g106917(.A0 (n_29495), .A1 (n_28404), .B0 (n_8401), .Y(n_30405));
OAI21X1 g106181(.A0 (n_29503), .A1 (n_21294), .B0 (n_30403), .Y(n_30404));
CLKBUFX1 gbuf_d_330(.A(n_29792), .Y(d_out_330));
CLKBUFX1 gbuf_q_330(.A(q_in_330), .Y(n_3235));
NAND2X1 g106959(.A (n_35042), .B (n_30399), .Y (n_32921));
NAND2X1 g106961(.A (n_35042), .B (n_33513), .Y (n_30397));
NOR3X1 g106963(.A (n_28263), .B (n_24912), .C (n_29477), .Y(n_30395));
NAND4X1 g106964(.A (n_35904), .B (n_24595), .C (n_35905), .D(n_27345), .Y (n_30394));
OAI21X1 g106971(.A0 (n_29593), .A1 (n_28515), .B0 (n_30956), .Y(n_30393));
NAND4X1 g106972(.A (n_28258), .B (n_25262), .C (n_29112), .D(n_27343), .Y (n_30392));
NOR2X1 g106978(.A (n_29990), .B (n_29976), .Y (n_30391));
NAND2X1 g106981(.A (n_29988), .B (n_13093), .Y (n_30390));
NAND3X1 g106986(.A (n_29510), .B (n_29481), .C (n_15158), .Y(n_30389));
NOR2X1 g106993(.A (n_28984), .B (n_29708), .Y (n_30388));
NAND2X1 g106995(.A (n_30386), .B (n_24786), .Y (n_30387));
OAI21X1 g106209(.A0 (n_29475), .A1 (n_22464), .B0 (n_31402), .Y(n_30385));
NAND4X1 g106999(.A (n_35440), .B (n_35441), .C (n_28531), .D(n_9066), .Y (n_30384));
NAND4X1 g107000(.A (n_32615), .B (n_32616), .C (n_28530), .D(n_27903), .Y (n_30383));
NAND2X1 g107001(.A (n_29980), .B (n_29948), .Y (n_30382));
OAI21X1 g107014(.A0 (n_29517), .A1 (n_27509), .B0 (n_30380), .Y(n_30381));
NAND3X1 g107017(.A (n_28594), .B (n_29592), .C (n_29032), .Y(n_30379));
NOR2X1 g107029(.A (n_30377), .B (n_29725), .Y (n_30378));
NOR2X1 g107037(.A (n_30377), .B (n_8661), .Y (n_30376));
NAND4X1 g107048(.A (n_28281), .B (n_27395), .C (n_29052), .D(n_24261), .Y (n_30375));
NOR2X1 g107055(.A (n_9935), .B (n_30015), .Y (n_30374));
NAND4X1 g107059(.A (n_32080), .B (n_32081), .C (n_29048), .D(n_24850), .Y (n_30373));
OAI21X1 g106240(.A0 (n_8595), .A1 (n_31414), .B0 (n_29961), .Y(n_35619));
NAND3X1 g107086(.A (n_9060), .B (n_21683), .C (n_29536), .Y(n_30368));
NOR2X1 g107090(.A (n_9076), .B (n_29958), .Y (n_32909));
OAI21X1 g107094(.A0 (n_29473), .A1 (n_27545), .B0 (n_33123), .Y(n_30366));
OAI21X1 g107097(.A0 (n_29485), .A1 (n_28119), .B0 (n_33123), .Y(n_30365));
OAI21X1 g107101(.A0 (n_29471), .A1 (n_27002), .B0 (n_30683), .Y(n_30364));
NAND4X1 g107108(.A (n_29106), .B (n_21663), .C (n_28620), .D(n_29088), .Y (n_30363));
NOR2X1 g107115(.A (n_29645), .B (n_30024), .Y (n_30362));
OAI21X1 g107118(.A0 (n_29514), .A1 (n_27292), .B0 (n_30360), .Y(n_30361));
MX2X1 g107136(.A (n_30355), .B (n_35043), .S0 (n_33092), .Y(n_30356));
OAI21X1 g107146(.A0 (n_29520), .A1 (n_27307), .B0 (n_30353), .Y(n_30354));
NOR2X1 g107148(.A (n_7078), .B (n_29715), .Y (n_30352));
AOI21X1 g107151(.A0 (n_15347), .A1 (n_30297), .B0 (n_29725), .Y(n_30351));
OAI21X1 g107153(.A0 (n_29502), .A1 (n_27267), .B0 (n_30353), .Y(n_30350));
NOR2X1 g107155(.A (n_7073), .B (n_29714), .Y (n_30349));
NAND4X1 g107157(.A (n_29108), .B (n_10608), .C (n_28630), .D(n_29089), .Y (n_30348));
AOI21X1 g107169(.A0 (n_8922), .A1 (n_30303), .B0 (n_20115), .Y(n_30347));
NAND2X1 g107173(.A (n_35431), .B (n_35432), .Y (n_30346));
OAI21X1 g107175(.A0 (n_29519), .A1 (n_33350), .B0 (n_6541), .Y(n_30345));
AOI21X1 g107187(.A0 (n_30298), .A1 (n_30836), .B0 (n_20724), .Y(n_30341));
NAND3X1 g107190(.A (n_29999), .B (n_28057), .C (n_29029), .Y(n_30339));
NOR2X1 g107214(.A (n_29413), .B (n_29865), .Y (n_30338));
NOR2X1 g107219(.A (n_29060), .B (n_29864), .Y (n_30337));
NOR2X1 g107221(.A (n_29059), .B (n_29854), .Y (n_30336));
NAND2X1 g107226(.A (n_29868), .B (n_31590), .Y (n_30335));
NAND2X1 g107228(.A (n_29842), .B (n_18933), .Y (n_30334));
NAND2X1 g107229(.A (n_32841), .B (n_991), .Y (n_30333));
NAND3X1 g107232(.A (n_29384), .B (n_29428), .C (n_29412), .Y(n_30332));
NOR2X1 g107237(.A (n_29822), .B (n_29518), .Y (n_30331));
OAI21X1 g107240(.A0 (n_29442), .A1 (n_28965), .B0 (n_31174), .Y(n_30330));
AOI21X1 g107244(.A0 (n_29467), .A1 (n_28957), .B0 (n_31178), .Y(n_30329));
NAND2X1 g107253(.A (n_29820), .B (n_29848), .Y (n_30328));
NAND4X1 g107260(.A (n_15152), .B (n_28355), .C (n_28354), .D(n_28884), .Y (n_30327));
NAND4X1 g107268(.A (n_32296), .B (n_28343), .C (n_28400), .D(n_32297), .Y (n_30326));
NAND2X1 g109477(.A (n_29700), .B (n_28288), .Y (n_30325));
NAND3X1 g107273(.A (n_29153), .B (n_29104), .C (n_28640), .Y(n_30324));
NAND2X1 g107274(.A (n_30321), .B (n_34753), .Y (n_30323));
NAND2X1 g107275(.A (n_30321), .B (n_28798), .Y (n_30322));
NAND2X1 g107276(.A (n_30321), .B (n_28785), .Y (n_30320));
NAND2X1 g106354(.A (n_29482), .B (n_31493), .Y (n_30319));
NAND2X1 g107277(.A (n_30321), .B (n_27798), .Y (n_30318));
NAND2X1 g106355(.A (n_29479), .B (n_31493), .Y (n_30317));
NAND2X1 g106357(.A (n_29487), .B (n_31201), .Y (n_30316));
NAND2X1 g106358(.A (n_29476), .B (n_31965), .Y (n_30315));
NAND3X1 g107284(.A (n_29146), .B (n_29101), .C (n_28475), .Y(n_30314));
OAI21X1 g107299(.A0 (n_29080), .A1 (n_27829), .B0 (n_30956), .Y(n_30311));
NOR2X1 g107304(.A (n_24885), .B (n_29494), .Y (n_30309));
NAND2X1 g107316(.A (n_33092), .B (n_991), .Y (n_30307));
NAND2X1 g107323(.A (n_28347), .B (n_30303), .Y (n_30304));
NAND2X1 g107324(.A (n_29695), .B (n_30303), .Y (n_30302));
OAI21X1 g106378(.A0 (n_28975), .A1 (n_22101), .B0 (n_31771), .Y(n_30301));
NAND2X1 g107329(.A (n_29480), .B (n_30295), .Y (n_30645));
AOI21X1 g106379(.A0 (n_29046), .A1 (n_28669), .B0 (n_31233), .Y(n_30300));
NAND2X1 g107330(.A (n_30298), .B (n_27632), .Y (n_30299));
NAND2X1 g107333(.A (n_30297), .B (n_29478), .Y (n_30834));
NAND2X1 g107335(.A (n_30295), .B (n_15409), .Y (n_30296));
OAI21X1 g107338(.A0 (n_29115), .A1 (n_28600), .B0 (n_30353), .Y(n_30294));
NAND2X1 g107346(.A (n_30291), .B (n_30288), .Y (n_30292));
NAND2X1 g107348(.A (n_29573), .B (n_29505), .Y (n_32201));
NAND2X1 g107349(.A (n_29568), .B (n_30288), .Y (n_32200));
NAND2X1 g107350(.A (n_29551), .B (n_30288), .Y (n_30287));
NAND4X1 g107355(.A (n_29062), .B (n_28583), .C (n_28035), .D(n_28489), .Y (n_30286));
AOI21X1 g106389(.A0 (n_29044), .A1 (n_28668), .B0 (n_31233), .Y(n_30285));
NOR2X1 g107358(.A (n_29307), .B (n_26185), .Y (n_35450));
NOR2X1 g107360(.A (n_29305), .B (n_26150), .Y (n_30283));
NOR2X1 g107362(.A (n_29306), .B (n_26120), .Y (n_30282));
NAND4X1 g107363(.A (n_28500), .B (n_19473), .C (n_28433), .D(n_28460), .Y (n_30281));
OAI21X1 g107366(.A0 (n_29023), .A1 (n_9626), .B0 (n_25230), .Y(n_30280));
OAI21X1 g107371(.A0 (n_29071), .A1 (n_28039), .B0 (n_31160), .Y(n_30279));
OAI21X1 g107372(.A0 (n_29070), .A1 (n_28038), .B0 (n_31628), .Y(n_30278));
NAND4X1 g107374(.A (n_35874), .B (n_35875), .C (n_35702), .D(n_28026), .Y (n_30277));
AOI21X1 g107378(.A0 (n_14399), .A1 (n_15029), .B0 (n_29530), .Y(n_32213));
NOR2X1 g107382(.A (n_29528), .B (n_28992), .Y (n_30274));
NOR2X1 g107384(.A (n_29522), .B (n_28991), .Y (n_30273));
NAND3X1 g107387(.A (n_28956), .B (n_28115), .C (n_28852), .Y(n_30272));
NAND3X1 g107391(.A (n_9065), .B (n_29092), .C (n_28641), .Y(n_30271));
NAND3X1 g107400(.A (n_9099), .B (n_29091), .C (n_28637), .Y(n_30270));
OAI21X1 g106415(.A0 (n_28994), .A1 (n_22102), .B0 (n_31771), .Y(n_30269));
NAND3X1 g107419(.A (n_29076), .B (n_29077), .C (n_28580), .Y(n_30268));
NOR2X1 g107421(.A (n_29647), .B (n_28731), .Y (n_30267));
OAI21X1 g107425(.A0 (n_9848), .A1 (n_30447), .B0 (n_29640), .Y(n_30266));
OAI21X1 g107426(.A0 (n_9879), .A1 (n_30447), .B0 (n_29639), .Y(n_30265));
NOR2X1 g107430(.A (n_8890), .B (n_29636), .Y (n_30264));
OAI21X1 g107440(.A0 (n_27543), .A1 (n_23138), .B0 (n_29558), .Y(n_30263));
AOI22X1 g107446(.A0 (n_29878), .A1 (n_33802), .B0 (n_21669), .B1(n_33803), .Y (n_30262));
NAND2X2 g107447(.A (n_29590), .B (n_29034), .Y (n_30874));
NAND2X1 g107453(.A (n_29548), .B (n_21704), .Y (n_30261));
NAND4X1 g107455(.A (n_28498), .B (n_18935), .C (n_27970), .D(n_28458), .Y (n_30260));
NOR2X1 g107457(.A (n_29646), .B (n_29509), .Y (n_30259));
OAI21X1 g106444(.A0 (n_28955), .A1 (n_22098), .B0 (n_30403), .Y(n_30258));
OAI21X1 g107472(.A0 (n_29024), .A1 (n_9625), .B0 (n_15350), .Y(n_30257));
NAND2X1 g107474(.A (n_29627), .B (n_15176), .Y (n_30256));
OAI21X1 g107476(.A0 (n_29036), .A1 (n_8505), .B0 (n_10362), .Y(n_30255));
OAI21X1 g107477(.A0 (n_9850), .A1 (n_28332), .B0 (n_29635), .Y(n_30254));
NAND2X2 g107482(.A (n_29598), .B (n_13493), .Y (n_30675));
NAND2X2 g107489(.A (n_29521), .B (n_29545), .Y (n_30860));
NAND2X1 g107490(.A (n_29588), .B (n_29014), .Y (n_30842));
INVX1 g107491(.A (n_30386), .Y (n_30253));
AOI21X1 g107493(.A0 (n_30454), .A1 (n_29567), .B0 (n_29554), .Y(n_32565));
NAND2X1 g107499(.A (n_29552), .B (n_20167), .Y (n_30251));
AOI22X1 g107500(.A0 (n_29917), .A1 (n_33738), .B0 (n_20165), .B1(n_30505), .Y (n_32564));
NAND2X1 g107501(.A (n_29574), .B (n_29662), .Y (n_30839));
NAND2X1 g107503(.A (n_29575), .B (n_29576), .Y (n_30641));
NAND2X1 g107511(.A (n_29538), .B (n_14885), .Y (n_30248));
NAND2X1 g107513(.A (n_29537), .B (n_29694), .Y (n_30837));
NAND4X1 g107515(.A (n_28503), .B (n_10898), .C (n_28445), .D(n_28472), .Y (n_30247));
NAND4X1 g107516(.A (n_28501), .B (n_10611), .C (n_27980), .D(n_28462), .Y (n_30246));
NAND2X1 g107534(.A (n_29587), .B (n_20118), .Y (n_30244));
OAI21X1 g107535(.A0 (n_29335), .A1 (n_30230), .B0 (n_20111), .Y(n_30243));
NAND2X1 g107536(.A (n_6940), .B (n_29597), .Y (n_30242));
NAND2X1 g107538(.A (n_6500), .B (n_29649), .Y (n_30241));
OAI21X1 g107540(.A0 (n_29047), .A1 (n_27698), .B0 (n_6520), .Y(n_30240));
NOR2X1 g106476(.A (n_29439), .B (n_29312), .Y (n_30239));
NAND2X1 g107541(.A (n_6931), .B (n_29644), .Y (n_30238));
NAND2X1 g107543(.A (n_6916), .B (n_29583), .Y (n_30237));
OAI21X1 g107548(.A0 (n_21228), .A1 (n_25540), .B0 (n_29524), .Y(n_35300));
OAI21X1 g106482(.A0 (n_28986), .A1 (n_22466), .B0 (n_35008), .Y(n_30235));
OAI21X1 g106485(.A0 (n_28980), .A1 (n_22465), .B0 (n_31544), .Y(n_30234));
NAND2X1 g107558(.A (n_29582), .B (n_21685), .Y (n_30233));
NOR2X1 g106486(.A (n_15013), .B (n_29500), .Y (n_30232));
OAI21X1 g107561(.A0 (n_32934), .A1 (n_30230), .B0 (n_21687), .Y(n_35299));
NAND4X1 g107584(.A (n_35268), .B (n_9136), .C (n_28277), .D(n_35269), .Y (n_30229));
NAND3X1 g107585(.A (n_20747), .B (n_28916), .C (n_28435), .Y(n_30228));
NAND3X1 g107586(.A (n_20215), .B (n_28914), .C (n_28894), .Y(n_30227));
NAND3X1 g107589(.A (n_28854), .B (n_28882), .C (n_28363), .Y(n_30226));
NOR2X1 g107598(.A (n_29320), .B (n_29045), .Y (n_30225));
NOR2X1 g107599(.A (n_29374), .B (n_19469), .Y (n_30224));
NAND3X1 g107611(.A (n_11129), .B (n_28919), .C (n_28446), .Y(n_30223));
NAND3X1 g107612(.A (n_11124), .B (n_28917), .C (n_28901), .Y(n_30222));
NAND2X1 g107615(.A (n_33546), .B (n_30220), .Y (n_30221));
OAI21X1 g106515(.A0 (n_28913), .A1 (n_31410), .B0 (n_9943), .Y(n_30219));
OAI21X1 g106516(.A0 (n_28912), .A1 (n_31410), .B0 (n_8619), .Y(n_30218));
NOR2X1 g106526(.A (n_6895), .B (n_29563), .Y (n_30217));
INVX1 g106527(.A (n_29931), .Y (n_30216));
NOR2X1 g107645(.A (n_29340), .B (n_18283), .Y (n_30215));
NOR2X1 g107646(.A (n_29321), .B (n_29371), .Y (n_30214));
NOR2X1 g107647(.A (n_29319), .B (n_29369), .Y (n_30213));
NOR2X1 g107648(.A (n_29318), .B (n_29368), .Y (n_30212));
NOR2X1 g107649(.A (n_29317), .B (n_29367), .Y (n_30211));
NOR2X1 g107650(.A (n_29316), .B (n_29365), .Y (n_30210));
NOR2X1 g107656(.A (n_9172), .B (n_30203), .Y (n_30208));
NOR2X1 g107666(.A (n_9172), .B (n_29346), .Y (n_35325));
NAND2X1 g107681(.A (n_30201), .B (n_30200), .Y (n_32599));
NAND2X1 g107696(.A (n_29353), .B (n_30197), .Y (n_32222));
AOI21X1 g107719(.A0 (n_28964), .A1 (n_28369), .B0 (n_31236), .Y(n_30196));
NAND2X1 g107723(.A (n_30220), .B (n_29445), .Y (n_30195));
NOR2X1 g107725(.A (n_29771), .B (n_8718), .Y (n_30194));
OAI21X1 g106561(.A0 (n_28888), .A1 (n_31538), .B0 (n_7106), .Y(n_30192));
NOR2X1 g107752(.A (n_29352), .B (n_29389), .Y (n_30191));
NOR2X1 g107753(.A (n_29350), .B (n_29039), .Y (n_30190));
NOR2X1 g107754(.A (n_28893), .B (n_29387), .Y (n_30189));
NOR2X1 g107758(.A (n_8382), .B (n_30514), .Y (n_30188));
NAND2X1 g107761(.A (n_29767), .B (n_24786), .Y (n_30187));
NAND2X1 g107775(.A (n_30182), .B (n_30184), .Y (n_30185));
AND2X1 g107776(.A (n_30182), .B (n_30557), .Y (n_30183));
NAND2X1 g107777(.A (n_30182), .B (n_30180), .Y (n_30181));
NAND2X1 g107778(.A (n_30182), .B (n_33513), .Y (n_30179));
NAND3X1 g107788(.A (n_27529), .B (n_28863), .C (n_20428), .Y(n_30177));
NAND3X1 g107790(.A (n_28072), .B (n_28862), .C (n_21708), .Y(n_30176));
NOR2X1 g107814(.A (n_29410), .B (n_27404), .Y (n_30175));
NAND4X1 g107819(.A (n_28408), .B (n_28304), .C (n_19568), .D(n_28407), .Y (n_30174));
NAND2X1 g107835(.A (n_30171), .B (n_28999), .Y (n_30173));
NAND2X1 g107837(.A (n_30171), .B (n_32935), .Y (n_30172));
CLKBUFX1 gbuf_d_331(.A(n_29474), .Y(d_out_331));
CLKBUFX1 gbuf_q_331(.A(q_in_331), .Y(n_13677));
AOI21X1 g107846(.A0 (n_28962), .A1 (n_28368), .B0 (n_31564), .Y(n_30170));
OAI21X1 g107850(.A0 (n_28240), .A1 (n_8927), .B0 (n_29342), .Y(n_30169));
NAND2X1 g107855(.A (n_30201), .B (n_30109), .Y (n_30168));
NAND2X1 g107869(.A (n_30165), .B (n_30184), .Y (n_30167));
AND2X1 g107870(.A (n_30165), .B (n_30557), .Y (n_30166));
NAND2X1 g107871(.A (n_30165), .B (n_30180), .Y (n_30164));
NAND2X1 g107872(.A (n_30165), .B (n_33494), .Y (n_30163));
NAND4X1 g107877(.A (n_29262), .B (n_27877), .C (n_25545), .D(n_28827), .Y (n_30162));
NAND3X1 g106629(.A (n_21225), .B (n_22479), .C (n_28841), .Y(n_30161));
NOR2X1 g107907(.A (n_29055), .B (n_29706), .Y (n_30160));
NOR2X1 g107922(.A (n_8915), .B (n_29464), .Y (n_30159));
NAND2X1 g106638(.A (n_29729), .B (n_28915), .Y (n_30158));
NAND4X1 g106642(.A (n_15269), .B (n_28702), .C (n_28701), .D(n_28728), .Y (n_30157));
NOR2X1 g107933(.A (n_28900), .B (n_29370), .Y (n_32913));
NOR2X1 g107934(.A (n_9095), .B (n_29332), .Y (n_32290));
NAND3X1 g107958(.A (n_10176), .B (n_28911), .C (n_28426), .Y(n_30153));
NAND3X1 g107960(.A (n_10129), .B (n_28910), .C (n_28892), .Y(n_30152));
NOR2X1 g107981(.A (n_8900), .B (n_29460), .Y (n_30151));
NOR2X1 g107985(.A (n_9044), .B (n_29328), .Y (n_30150));
NOR2X1 g107987(.A (n_29468), .B (n_29053), .Y (n_30149));
NAND3X1 g107992(.A (n_10224), .B (n_28908), .C (n_28399), .Y(n_30148));
NAND3X1 g107993(.A (n_10208), .B (n_28907), .C (n_28871), .Y(n_30147));
NOR2X1 g107996(.A (n_28383), .B (n_29366), .Y (n_30146));
INVX1 g107998(.A (n_30145), .Y (n_30566));
NOR2X1 g108011(.A (n_28959), .B (n_29450), .Y (n_30143));
NOR2X1 g108059(.A (n_28373), .B (n_29327), .Y (n_30142));
NAND2X1 g108060(.A (n_29417), .B (n_20186), .Y (n_30141));
NAND4X1 g108082(.A (n_28828), .B (n_10615), .C (n_28261), .D(n_28804), .Y (n_30140));
MX2X1 g108085(.A (n_27564), .B (n_30138), .S0 (n_28007), .Y(n_30139));
NAND2X1 g108090(.A (n_29426), .B (n_20128), .Y (n_30137));
NAND2X1 g108092(.A (n_29432), .B (n_20121), .Y (n_30136));
OAI21X1 g108094(.A0 (n_29263), .A1 (n_8333), .B0 (n_20113), .Y(n_30135));
NAND2X1 g108101(.A (n_6602), .B (n_29466), .Y (n_30134));
OAI21X1 g108104(.A0 (n_19485), .A1 (n_25540), .B0 (n_29400), .Y(n_30133));
OAI21X1 g106718(.A0 (n_9557), .A1 (n_215), .B0 (n_29287), .Y(n_30132));
AOI21X1 g108110(.A0 (n_33546), .A1 (n_29850), .B0 (n_29303), .Y(n_35449));
NOR2X1 g106720(.A (n_10361), .B (n_29361), .Y (n_30130));
NAND2X1 g108127(.A (n_28367), .B (n_29671), .Y (n_30129));
NAND4X1 g108130(.A (n_29663), .B (n_27582), .C (n_15284), .D(n_23803), .Y (n_30128));
NOR2X1 g108143(.A (n_29705), .B (n_28860), .Y (n_30127));
NOR2X1 g108146(.A (n_29704), .B (n_28341), .Y (n_30126));
NOR2X1 g108147(.A (n_29703), .B (n_28858), .Y (n_30125));
NOR2X1 g108164(.A (n_29308), .B (n_25721), .Y (n_35927));
NAND2X1 g108199(.A (n_30122), .B (n_30200), .Y (n_32171));
NOR2X1 g106764(.A (n_10448), .B (n_29348), .Y (n_30121));
NAND4X1 g108228(.A (n_32084), .B (n_28799), .C (n_32085), .D(n_27342), .Y (n_30120));
NAND4X1 g108246(.A (n_32088), .B (n_28794), .C (n_32089), .D(n_27337), .Y (n_30119));
CLKBUFX1 gbuf_d_332(.A(n_29660), .Y(d_out_332));
CLKBUFX1 gbuf_q_332(.A(q_in_332), .Y(n_10363));
CLKBUFX1 gbuf_d_333(.A(n_29282), .Y(d_out_333));
CLKBUFX1 gbuf_q_333(.A(q_in_333), .Y(n_13341));
CLKBUFX1 gbuf_d_334(.A(n_29284), .Y(d_out_334));
CLKBUFX1 gbuf_q_334(.A(q_in_334), .Y(P2_reg1[8]));
CLKBUFX1 gbuf_d_335(.A(n_29286), .Y(d_out_335));
CLKBUFX1 gbuf_q_335(.A(q_in_335), .Y(n_9592));
CLKBUFX1 gbuf_d_336(.A(n_29283), .Y(d_out_336));
CLKBUFX1 gbuf_q_336(.A(q_in_336), .Y(P2_reg2[8]));
CLKBUFX1 gbuf_d_337(.A(n_29659), .Y(d_out_337));
CLKBUFX1 gbuf_q_337(.A(q_in_337), .Y(P2_reg1[4]));
CLKBUFX1 gbuf_d_338(.A(n_29658), .Y(d_out_338));
CLKBUFX1 gbuf_q_338(.A(q_in_338), .Y(n_13202));
CLKBUFX1 gbuf_d_339(.A(n_29472), .Y(d_out_339));
CLKBUFX1 gbuf_q_339(.A(q_in_339), .Y(n_13332));
NOR2X1 g106779(.A (n_7081), .B (n_29398), .Y (n_30118));
NOR2X1 g108267(.A (n_30449), .B (n_8382), .Y (n_30117));
NAND3X1 g108282(.A (n_27082), .B (n_29243), .C (n_28708), .Y(n_30116));
NAND2X1 g108283(.A (n_29300), .B (n_28366), .Y (n_30115));
NOR2X1 g108289(.A (n_28856), .B (n_29279), .Y (n_35079));
NOR2X1 g108291(.A (n_29712), .B (n_8382), .Y (n_30113));
NAND2X1 g108333(.A (n_30171), .B (n_28840), .Y (n_30111));
NAND2X1 g108349(.A (n_30122), .B (n_30109), .Y (n_30110));
NAND4X1 g108369(.A (n_29292), .B (n_28684), .C (n_15290), .D(n_23805), .Y (n_30108));
AOI21X1 g106853(.A0 (n_9424), .A1 (n_29181), .B0 (n_31105), .Y(n_30107));
AOI21X1 g106860(.A0 (n_10345), .A1 (n_29214), .B0 (n_349), .Y(n_30106));
NAND2X1 g108477(.A (n_29297), .B (n_28318), .Y (n_30105));
NAND2X1 g106883(.A (n_29682), .B (n_31594), .Y (n_30104));
OAI21X1 g106903(.A0 (n_29175), .A1 (n_27449), .B0 (n_33123), .Y(n_30103));
OAI21X1 g106911(.A0 (n_29165), .A1 (n_25568), .B0 (n_30099), .Y(n_30100));
OAI21X1 g106176(.A0 (n_27568), .A1 (n_7971), .B0 (n_29637), .Y(n_30098));
OAI21X1 g106922(.A0 (n_29185), .A1 (n_28043), .B0 (n_31174), .Y(n_30097));
NAND2X1 g106924(.A (n_9503), .B (n_30087), .Y (n_30096));
NAND2X1 g106926(.A (n_30094), .B (n_29925), .Y (n_30095));
NAND2X1 g106927(.A (n_32850), .B (n_29925), .Y (n_30093));
NAND2X1 g106929(.A (n_30094), .B (n_25980), .Y (n_30090));
NAND2X1 g106934(.A (n_30087), .B (n_33785), .Y (n_30088));
NOR2X1 g106949(.A (n_26977), .B (n_29679), .Y (n_30086));
NOR2X1 g106968(.A (n_28012), .B (n_29702), .Y (n_30085));
NOR2X1 g106983(.A (n_26942), .B (n_29701), .Y (n_30084));
NOR2X1 g106998(.A (n_29680), .B (n_29139), .Y (n_30083));
NOR2X1 g107004(.A (n_26976), .B (n_29674), .Y (n_30082));
NAND2X1 g107005(.A (n_29672), .B (n_31850), .Y (n_30081));
NAND2X1 g107021(.A (n_30079), .B (n_26238), .Y (n_32607));
AOI21X1 g107022(.A0 (n_28597), .A1 (n_29926), .B0 (n_25552), .Y(n_35647));
AOI21X1 g107023(.A0 (n_29065), .A1 (n_29919), .B0 (n_25550), .Y(n_30076));
AOI21X1 g107024(.A0 (n_28948), .A1 (n_29915), .B0 (n_25546), .Y(n_30075));
NAND2X1 g107038(.A (n_30068), .B (n_28374), .Y (n_30072));
NOR2X1 g107039(.A (n_29167), .B (n_29665), .Y (n_30071));
OAI21X1 g107041(.A0 (n_29149), .A1 (n_27507), .B0 (n_31240), .Y(n_30070));
NAND2X1 g107044(.A (n_30068), .B (n_29405), .Y (n_32146));
NAND2X1 g107045(.A (n_30068), .B (n_33738), .Y (n_30066));
OAI21X1 g107050(.A0 (n_29190), .A1 (n_28588), .B0 (n_8618), .Y(n_30065));
AOI22X1 g107051(.A0 (n_30020), .A1 (n_30063), .B0 (n_9629), .B1(n_20080), .Y (n_30064));
NAND2X1 g107053(.A (n_29678), .B (n_31594), .Y (n_30062));
AOI22X1 g107063(.A0 (n_30013), .A1 (n_30063), .B0 (n_9629), .B1(n_20077), .Y (n_30061));
NAND2X1 g107066(.A (n_29677), .B (n_31594), .Y (n_30059));
AOI21X1 g107067(.A0 (n_29186), .A1 (n_28790), .B0 (n_31564), .Y(n_30058));
AOI22X1 g107076(.A0 (n_30005), .A1 (n_30063), .B0 (n_20304), .B1(n_20076), .Y (n_30057));
OAI21X1 g107077(.A0 (n_29184), .A1 (n_26872), .B0 (n_30353), .Y(n_30056));
NAND3X1 g107080(.A (n_29058), .B (n_29183), .C (n_29010), .Y(n_30055));
NAND3X1 g107085(.A (n_9124), .B (n_20117), .C (n_29163), .Y(n_30054));
OAI21X1 g107089(.A0 (n_29174), .A1 (n_30619), .B0 (n_8612), .Y(n_30053));
NOR2X1 g107092(.A (n_9581), .B (n_29661), .Y (n_30052));
OAI21X1 g107100(.A0 (n_30050), .A1 (n_29127), .B0 (n_29238), .Y(n_30051));
OAI21X1 g106266(.A0 (n_29131), .A1 (n_31726), .B0 (n_7157), .Y(n_30049));
NOR2X1 g107114(.A (n_29223), .B (n_29707), .Y (n_30048));
NAND2X1 g107116(.A (n_29689), .B (n_22473), .Y (n_30047));
OAI21X1 g107119(.A0 (n_29141), .A1 (n_26862), .B0 (n_30360), .Y(n_30046));
OAI21X1 g107142(.A0 (n_29147), .A1 (n_26884), .B0 (n_31544), .Y(n_30045));
OAI21X1 g107143(.A0 (n_29144), .A1 (n_26878), .B0 (n_30353), .Y(n_30044));
NAND2X1 g107186(.A (n_29699), .B (n_22470), .Y (n_30043));
OAI21X1 g107188(.A0 (n_29127), .A1 (n_8352), .B0 (n_22471), .Y(n_30042));
AOI21X1 g107206(.A0 (n_10464), .A1 (n_29038), .B0 (n_30968), .Y(n_30041));
NAND4X1 g107215(.A (n_29066), .B (n_10218), .C (n_28385), .D(n_28450), .Y (n_30040));
NAND4X1 g107216(.A (n_29064), .B (n_9608), .C (n_28004), .D(n_28473), .Y (n_30039));
NAND4X1 g107217(.A (n_29063), .B (n_9583), .C (n_27991), .D(n_28469), .Y (n_30038));
NOR2X1 g107218(.A (n_28596), .B (n_29511), .Y (n_30037));
NOR2X1 g107220(.A (n_28595), .B (n_29501), .Y (n_30036));
NAND2X1 g107225(.A (n_29515), .B (n_31965), .Y (n_30035));
NAND4X1 g107230(.A (n_25744), .B (n_10166), .C (n_28424), .D(n_28456), .Y (n_30034));
NAND4X1 g107231(.A (n_25730), .B (n_10159), .C (n_28391), .D(n_28454), .Y (n_30033));
AOI21X1 g107239(.A0 (n_29118), .A1 (n_28514), .B0 (n_8070), .Y(n_30030));
AOI21X1 g106340(.A0 (n_9961), .A1 (n_28961), .B0 (n_30702), .Y(n_30029));
NAND2X1 g107256(.A (n_30027), .B (n_28492), .Y (n_30028));
NAND2X1 g107258(.A (n_30027), .B (n_10063), .Y (n_30026));
NAND4X1 g107262(.A (n_15285), .B (n_28353), .C (n_28352), .D(n_28412), .Y (n_30025));
NAND4X1 g107264(.A (n_15034), .B (n_27887), .C (n_27931), .D(n_27890), .Y (n_30024));
NAND4X1 g107265(.A (n_14742), .B (n_27884), .C (n_27434), .D(n_27889), .Y (n_30023));
NAND4X1 g107267(.A (n_32230), .B (n_27882), .C (n_27930), .D(n_32231), .Y (n_30022));
NAND2X1 g107278(.A (n_30020), .B (n_25756), .Y (n_32112));
NAND2X1 g107279(.A (n_34753), .B (n_30020), .Y (n_30018));
NAND2X1 g107280(.A (n_30020), .B (n_26528), .Y (n_30017));
AOI21X1 g107281(.A0 (n_28672), .A1 (n_28601), .B0 (n_31236), .Y(n_30015));
NAND2X2 g107286(.A (n_30013), .B (n_34753), .Y (n_30012));
NAND2X1 g107287(.A (n_30013), .B (n_26528), .Y (n_30010));
NOR2X1 g109515(.A (n_29140), .B (n_11117), .Y (n_30009));
NAND3X1 g109516(.A (n_10847), .B (n_28682), .C (n_25775), .Y(n_30008));
NOR2X1 g107294(.A (n_29143), .B (n_29123), .Y (n_30007));
NAND2X1 g107297(.A (n_30005), .B (n_10808), .Y (n_30004));
NAND2X1 g107298(.A (n_30005), .B (n_26528), .Y (n_30003));
NOR2X1 g107307(.A (n_29142), .B (n_29138), .Y (n_30002));
NAND2X1 g107351(.A (n_29136), .B (n_13194), .Y (n_30000));
AOI21X1 g107377(.A0 (n_14336), .A1 (n_15029), .B0 (n_29158), .Y(n_29999));
NAND4X1 g107379(.A (n_14735), .B (n_27929), .C (n_27917), .D(n_27426), .Y (n_29998));
OAI21X1 g106403(.A0 (n_28521), .A1 (n_28120), .B0 (n_31174), .Y(n_29997));
OAI21X1 g107389(.A0 (n_28557), .A1 (n_29388), .B0 (n_22140), .Y(n_29996));
OAI21X1 g107392(.A0 (n_8270), .A1 (n_31480), .B0 (n_29220), .Y(n_29995));
NAND4X1 g107397(.A (n_32315), .B (n_28116), .C (n_32316), .D(n_27666), .Y (n_29994));
OAI21X1 g107404(.A0 (n_28552), .A1 (n_29388), .B0 (n_22134), .Y(n_29993));
NAND4X1 g107406(.A (n_28036), .B (n_27812), .C (n_27678), .D(n_27878), .Y (n_29991));
OAI21X1 g107414(.A0 (n_29975), .A1 (n_29388), .B0 (n_22128), .Y(n_29990));
AOI22X1 g107416(.A0 (n_28566), .A1 (n_15723), .B0 (n_1721), .B1(n_9382), .Y (n_29988));
OAI21X1 g107420(.A0 (n_28546), .A1 (n_29388), .B0 (n_22121), .Y(n_29986));
AOI21X1 g107424(.A0 (n_15415), .A1 (n_29544), .B0 (n_8927), .Y(n_29985));
OAI21X1 g107428(.A0 (n_9846), .A1 (n_31019), .B0 (n_29217), .Y(n_29984));
NAND4X1 g107429(.A (n_29114), .B (n_28576), .C (n_28296), .D(n_26916), .Y (n_29983));
NOR2X1 g107434(.A (n_9891), .B (n_29216), .Y (n_29982));
NOR2X1 g107435(.A (n_10279), .B (n_29215), .Y (n_29981));
AOI21X1 g107448(.A0 (n_30171), .A1 (n_29947), .B0 (n_28677), .Y(n_29980));
AOI21X1 g107449(.A0 (n_30171), .A1 (n_29959), .B0 (n_29128), .Y(n_29978));
OAI21X1 g107452(.A0 (n_29975), .A1 (n_25119), .B0 (n_29202), .Y(n_29976));
NOR2X1 g106438(.A (n_29082), .B (n_27550), .Y (n_32880));
NAND4X1 g106440(.A (n_29002), .B (n_26960), .C (n_25252), .D(n_25246), .Y (n_29973));
INVX1 g107467(.A (n_30087), .Y (n_29972));
OAI21X1 g107471(.A0 (n_14933), .A1 (n_29968), .B0 (n_29211), .Y(n_29971));
AOI21X1 g107473(.A0 (n_29623), .A1 (n_34952), .B0 (n_15304), .Y(n_29970));
OAI21X1 g107475(.A0 (n_14925), .A1 (n_29968), .B0 (n_29206), .Y(n_29969));
NOR2X1 g107478(.A (n_9923), .B (n_29213), .Y (n_29967));
NOR2X1 g107479(.A (n_10390), .B (n_29212), .Y (n_29966));
NAND2X1 g107492(.A (n_29177), .B (n_29666), .Y (n_30386));
INVX2 g107506(.A (n_29962), .Y (n_30377));
OAI21X1 g106468(.A0 (n_28502), .A1 (n_28118), .B0 (n_31240), .Y(n_29961));
AOI21X1 g107526(.A0 (n_29959), .A1 (n_13952), .B0 (n_22119), .Y(n_29960));
NAND2X1 g107530(.A (n_29171), .B (n_20125), .Y (n_29958));
AOI21X1 g107531(.A0 (n_29170), .A1 (n_29955), .B0 (n_29173), .Y(n_29957));
NAND2X1 g107546(.A (n_6684), .B (n_29225), .Y (n_29954));
NAND2X1 g107547(.A (n_29154), .B (n_20110), .Y (n_29953));
NAND2X1 g107552(.A (n_29204), .B (n_29221), .Y (n_29952));
OAI21X1 g107554(.A0 (n_28553), .A1 (n_10790), .B0 (n_29219), .Y(n_29951));
OAI21X1 g107557(.A0 (n_28547), .A1 (n_10790), .B0 (n_29218), .Y(n_29950));
AOI21X1 g107560(.A0 (n_29947), .A1 (n_13952), .B0 (n_20725), .Y(n_29948));
NAND3X1 g106498(.A (n_7559), .B (n_28562), .C (n_29944), .Y(n_29945));
NAND3X1 g107591(.A (n_28334), .B (n_28410), .C (n_28362), .Y(n_29943));
NAND4X1 g107594(.A (n_28494), .B (n_28040), .C (n_28001), .D(n_21222), .Y (n_29942));
NAND2X1 g107595(.A (n_28972), .B (n_28587), .Y (n_29941));
NAND4X1 g107596(.A (n_28491), .B (n_28037), .C (n_27989), .D(n_21214), .Y (n_29940));
NOR2X1 g107606(.A (n_29007), .B (n_19117), .Y (n_32214));
NAND3X1 g107614(.A (n_11149), .B (n_28443), .C (n_28014), .Y(n_29938));
OAI21X1 g107619(.A0 (n_28439), .A1 (n_27183), .B0 (n_30569), .Y(n_29937));
OAI21X1 g107620(.A0 (n_28438), .A1 (n_27182), .B0 (n_30569), .Y(n_29936));
NAND3X1 g107622(.A (n_18287), .B (n_28429), .C (n_28011), .Y(n_29935));
NAND2X1 g107623(.A (n_33546), .B (n_29893), .Y (n_29934));
NAND2X1 g107624(.A (n_33546), .B (n_29889), .Y (n_29933));
NOR2X1 g107635(.A (n_28328), .B (n_29072), .Y (n_29932));
NAND2X1 g106528(.A (n_29121), .B (n_27022), .Y (n_29931));
NOR2X1 g107653(.A (n_29019), .B (n_9626), .Y (n_29930));
NAND2X1 g107670(.A (n_29926), .B (n_29925), .Y (n_29927));
NOR2X1 g107675(.A (n_29923), .B (n_8668), .Y (n_29924));
NAND2X1 g107679(.A (n_29919), .B (n_29925), .Y (n_29920));
NAND2X1 g107680(.A (n_29917), .B (n_30200), .Y (n_32152));
NAND2X1 g107683(.A (n_29915), .B (n_29925), .Y (n_29916));
NAND2X1 g107686(.A (n_34774), .B (n_29908), .Y (n_29913));
NAND2X1 g107689(.A (n_29926), .B (n_28013), .Y (n_29911));
NAND2X1 g107698(.A (n_35058), .B (n_33785), .Y (n_29910));
NAND2X1 g107702(.A (n_29919), .B (n_29908), .Y (n_29909));
NAND2X1 g107705(.A (n_29906), .B (n_29455), .Y (n_29907));
NAND2X1 g107707(.A (n_29908), .B (n_29915), .Y (n_29905));
NAND2X1 g107715(.A (n_29359), .B (n_34753), .Y (n_29904));
NAND4X1 g107736(.A (n_25783), .B (n_24597), .C (n_28286), .D(n_27036), .Y (n_29902));
NAND2X1 g107737(.A (n_29355), .B (n_10808), .Y (n_29901));
NOR2X1 g107744(.A (n_27976), .B (n_29043), .Y (n_29900));
NAND4X1 g107746(.A (n_25764), .B (n_24577), .C (n_28291), .D(n_26163), .Y (n_29899));
NAND2X1 g107747(.A (n_29025), .B (n_12810), .Y (n_29898));
NAND2X1 g107763(.A (n_29893), .B (n_28431), .Y (n_29894));
OAI21X1 g107770(.A0 (n_28338), .A1 (n_27185), .B0 (n_31398), .Y(n_29892));
OAI21X1 g107771(.A0 (n_28337), .A1 (n_27184), .B0 (n_30380), .Y(n_29891));
NAND3X1 g107782(.A (n_26935), .B (n_28309), .C (n_15267), .Y(n_29888));
NAND3X1 g107784(.A (n_28335), .B (n_28308), .C (n_15253), .Y(n_29887));
NAND3X1 g107786(.A (n_28073), .B (n_28365), .C (n_21343), .Y(n_29886));
NAND2X1 g106596(.A (n_28896), .B (n_31092), .Y (n_29885));
NAND4X1 g107817(.A (n_27940), .B (n_27839), .C (n_20726), .D(n_27939), .Y (n_29884));
NOR2X1 g107833(.A (n_28977), .B (n_10622), .Y (n_29883));
NAND2X1 g107851(.A (n_29917), .B (n_30109), .Y (n_29881));
NOR2X1 g107856(.A (n_29345), .B (n_29553), .Y (n_29880));
NAND2X1 g107875(.A (n_29878), .B (n_33513), .Y (n_29875));
NAND3X1 g107906(.A (n_28389), .B (n_28387), .C (n_28386), .Y(n_29873));
NOR2X1 g107908(.A (n_27998), .B (n_29051), .Y (n_29872));
NAND4X1 g107931(.A (n_32161), .B (n_32162), .C (n_28236), .D(n_24248), .Y (n_29871));
NAND4X1 g107941(.A (n_28287), .B (n_27258), .C (n_27587), .D(n_28235), .Y (n_29870));
NAND3X1 g107945(.A (n_28031), .B (n_28436), .C (n_28190), .Y(n_29869));
OAI21X1 g107948(.A0 (n_8822), .A1 (n_31122), .B0 (n_29081), .Y(n_29868));
NOR2X1 g107954(.A (n_29117), .B (n_28078), .Y (n_29867));
NAND3X1 g107965(.A (n_28421), .B (n_19584), .C (n_28419), .Y(n_29866));
NAND3X1 g107966(.A (n_10164), .B (n_28455), .C (n_28422), .Y(n_29865));
NAND3X1 g107967(.A (n_10163), .B (n_28417), .C (n_28009), .Y(n_29864));
NOR2X1 g107971(.A (n_9064), .B (n_28983), .Y (n_29863));
NOR2X1 g107972(.A (n_9078), .B (n_28982), .Y (n_29862));
NAND3X1 g107973(.A (n_9063), .B (n_20715), .C (n_28361), .Y(n_29861));
NAND2X1 g106661(.A (n_28866), .B (n_12894), .Y (n_29860));
NAND3X1 g107975(.A (n_9061), .B (n_19565), .C (n_28359), .Y(n_29859));
NOR2X1 g107983(.A (n_9053), .B (n_28996), .Y (n_32616));
NOR2X1 g107984(.A (n_9058), .B (n_28988), .Y (n_35909));
NOR2X1 g107986(.A (n_29116), .B (n_29054), .Y (n_29856));
NAND4X1 g107995(.A (n_32113), .B (n_32114), .C (n_28223), .D(n_24228), .Y (n_29855));
NAND3X1 g107997(.A (n_10137), .B (n_28381), .C (n_28008), .Y(n_29854));
INVX1 g107999(.A (n_29498), .Y (n_30145));
AOI21X1 g108008(.A0 (n_30171), .A1 (n_29817), .B0 (n_29001), .Y(n_29853));
NAND4X1 g108015(.A (n_29086), .B (n_25212), .C (n_26574), .D(n_26605), .Y (n_29852));
AOI21X1 g108020(.A0 (n_29850), .A1 (n_30180), .B0 (n_20187), .Y(n_29851));
AOI21X1 g108021(.A0 (n_29841), .A1 (n_30180), .B0 (n_20159), .Y(n_29849));
AOI22X1 g108023(.A0 (n_29819), .A1 (n_30180), .B0 (n_19493), .B1(n_33803), .Y (n_29848));
NAND2X2 g108041(.A (n_29084), .B (n_28325), .Y (n_30594));
OAI21X1 g108045(.A0 (n_30445), .A1 (n_27862), .B0 (n_29097), .Y(n_29843));
AOI22X1 g108051(.A0 (n_29841), .A1 (n_30668), .B0 (n_29839), .B1(n_33785), .Y (n_29842));
AOI22X1 g108054(.A0 (n_29841), .A1 (n_33494), .B0 (n_29839), .B1(n_34709), .Y (n_29840));
NOR2X1 g108056(.A (n_27906), .B (n_28987), .Y (n_35440));
NOR2X1 g108058(.A (n_27901), .B (n_28985), .Y (n_35908));
NOR2X1 g108064(.A (n_28357), .B (n_28970), .Y (n_29836));
NOR2X1 g108065(.A (n_28356), .B (n_28967), .Y (n_29835));
INVX1 g108071(.A (n_30298), .Y (n_29834));
INVX2 g108077(.A (n_29831), .Y (n_29833));
INVX1 g108078(.A (n_29831), .Y (n_29832));
AOI22X1 g108089(.A0 (n_29422), .A1 (n_33494), .B0 (n_28905), .B1(n_28926), .Y (n_29829));
AOI21X1 g108091(.A0 (n_29425), .A1 (n_30636), .B0 (n_29074), .Y(n_29827));
NAND2X1 g108096(.A (n_6863), .B (n_29111), .Y (n_29826));
NAND2X1 g108100(.A (n_6910), .B (n_29078), .Y (n_29825));
NAND2X1 g108251(.A (n_29272), .B (n_34753), .Y (n_32119));
NAND2X1 g108107(.A (n_6908), .B (n_29073), .Y (n_29823));
OAI21X1 g108113(.A0 (n_30445), .A1 (n_27850), .B0 (n_29099), .Y(n_29822));
AOI21X1 g108114(.A0 (n_33546), .A1 (n_29819), .B0 (n_28928), .Y(n_29820));
AOI21X1 g108115(.A0 (n_29817), .A1 (n_13952), .B0 (n_20728), .Y(n_29818));
NOR2X1 g108121(.A (n_27505), .B (n_28857), .Y (n_29816));
NOR2X1 g108128(.A (n_28784), .B (n_28855), .Y (n_29815));
NOR2X1 g108129(.A (n_28783), .B (n_28853), .Y (n_29814));
NAND3X1 g108148(.A (n_18290), .B (n_28802), .C (n_28256), .Y(n_29813));
NAND3X1 g108167(.A (n_28947), .B (n_24980), .C (n_14877), .Y(n_29811));
NAND3X1 g108168(.A (n_28946), .B (n_25947), .C (n_14967), .Y(n_29810));
NAND3X1 g108170(.A (n_28944), .B (n_14434), .C (n_24929), .Y(n_29809));
NAND3X1 g108171(.A (n_28943), .B (n_25893), .C (n_14966), .Y(n_29808));
NOR2X1 g108175(.A (n_9172), .B (n_28846), .Y (n_29807));
NOR2X1 g108178(.A (n_9502), .B (n_28845), .Y (n_29806));
NOR2X1 g108186(.A (n_9172), .B (n_28844), .Y (n_29805));
OAI21X1 g108216(.A0 (n_15079), .A1 (n_8614), .B0 (n_28861), .Y(n_29804));
NOR2X1 g108224(.A (n_28849), .B (n_14376), .Y (n_29803));
NAND4X1 g108229(.A (n_35091), .B (n_28280), .C (n_35092), .D(n_27339), .Y (n_29802));
NAND3X1 g108231(.A (n_27373), .B (n_28824), .C (n_27310), .Y(n_29801));
NAND2X1 g108233(.A (n_29275), .B (n_34753), .Y (n_35107));
NAND4X1 g108247(.A (n_35093), .B (n_28271), .C (n_35094), .D(n_27334), .Y (n_29799));
NAND3X1 g108249(.A (n_27372), .B (n_28820), .C (n_27302), .Y(n_29798));
CLKBUFX1 gbuf_d_340(.A(n_28963), .Y(d_out_340));
CLKBUFX1 gbuf_q_340(.A(q_in_340), .Y(P2_reg3[3]));
CLKBUFX1 gbuf_d_341(.A(n_29232), .Y(d_out_341));
CLKBUFX1 gbuf_q_341(.A(q_in_341), .Y(n_13511));
CLKBUFX1 gbuf_d_342(.A(n_29168), .Y(d_out_342));
CLKBUFX1 gbuf_q_342(.A(q_in_342), .Y(n_13675));
CLKBUFX1 gbuf_d_343(.A(n_28978), .Y(d_out_343));
CLKBUFX1 gbuf_q_343(.A(q_in_343), .Y(n_13211));
NAND3X1 g108266(.A (n_27370), .B (n_28816), .C (n_27295), .Y(n_29797));
NAND2X1 g108268(.A (n_29270), .B (n_34753), .Y (n_29796));
NAND3X1 g108287(.A (n_27369), .B (n_34695), .C (n_27288), .Y(n_29795));
NAND2X1 g108293(.A (n_29269), .B (n_34753), .Y (n_29794));
NAND2X1 g108307(.A (n_28007), .B (n_7967), .Y (n_29793));
NAND2X1 g106798(.A (n_6947), .B (n_29037), .Y (n_29792));
OAI21X1 g106811(.A0 (n_28782), .A1 (n_31541), .B0 (n_6943), .Y(n_29791));
NOR2X1 g108350(.A (n_29268), .B (n_29553), .Y (n_29790));
NAND3X1 g108361(.A (n_28239), .B (n_28754), .C (n_27254), .Y(n_29789));
NAND3X1 g108418(.A (n_9606), .B (n_28807), .C (n_27802), .Y(n_29788));
NAND3X1 g108429(.A (n_9042), .B (n_28806), .C (n_28268), .Y(n_29787));
NAND3X1 g106147(.A (n_12142), .B (n_27005), .C (n_28687), .Y(n_29786));
NAND3X1 g108431(.A (n_35111), .B (n_35112), .C (n_27790), .Y(n_29785));
NAND2X1 g108453(.A (n_21712), .B (n_28889), .Y (n_29784));
NAND2X1 g106868(.A (n_29244), .B (n_31205), .Y (n_29783));
NAND4X1 g106878(.A (n_25123), .B (n_9179), .C (n_28093), .D(n_28098), .Y (n_29782));
NAND2X1 g108476(.A (n_28872), .B (n_27843), .Y (n_29781));
OAI21X1 g108479(.A0 (n_28767), .A1 (n_8718), .B0 (n_21709), .Y(n_29780));
NAND4X1 g106881(.A (n_32115), .B (n_9143), .C (n_32116), .D(n_28097), .Y (n_29779));
NAND3X1 g106887(.A (n_28685), .B (n_28725), .C (n_28706), .Y(n_29778));
INVX1 g108506(.A (n_29372), .Y (n_29777));
OAI21X1 g106898(.A0 (n_28732), .A1 (n_27464), .B0 (n_33123), .Y(n_29776));
OAI21X1 g108525(.A0 (n_14701), .A1 (n_8614), .B0 (n_28895), .Y(n_29775));
AOI21X1 g108526(.A0 (n_30454), .A1 (n_29760), .B0 (n_28869), .Y(n_35148));
AOI21X1 g106909(.A0 (n_28718), .A1 (n_27510), .B0 (n_29769), .Y(n_29770));
INVX1 g108566(.A (n_30203), .Y (n_29768));
INVX1 g108578(.A (n_29767), .Y (n_30478));
NAND2X1 g106913(.A (n_29242), .B (n_29235), .Y (n_29766));
AOI21X1 g106918(.A0 (n_28680), .A1 (n_26947), .B0 (n_33125), .Y(n_29765));
OAI21X1 g106919(.A0 (n_28679), .A1 (n_25573), .B0 (n_30099), .Y(n_29763));
NAND2X1 g108614(.A (n_28876), .B (n_19602), .Y (n_29762));
AOI21X1 g108620(.A0 (n_29427), .A1 (n_29760), .B0 (n_28921), .Y(n_29761));
AOI21X1 g108623(.A0 (n_29295), .A1 (n_29523), .B0 (n_20143), .Y(n_29759));
AOI21X1 g108660(.A0 (n_29067), .A1 (n_25988), .B0 (n_28898), .Y(n_29758));
AOI21X1 g108661(.A0 (n_29392), .A1 (n_26528), .B0 (n_28939), .Y(n_32886));
AOI21X1 g108663(.A0 (n_34712), .A1 (n_29390), .B0 (n_28935), .Y(n_29755));
AOI21X1 g108664(.A0 (n_28384), .A1 (n_33513), .B0 (n_28920), .Y(n_29753));
NAND2X1 g108673(.A (n_28375), .B (n_28877), .Y (n_29751));
NAND2X1 g108676(.A (n_28885), .B (n_20716), .Y (n_29750));
OAI21X1 g108682(.A0 (n_29230), .A1 (n_8333), .B0 (n_19560), .Y(n_29749));
NAND4X1 g108697(.A (n_27659), .B (n_28224), .C (n_28171), .D(n_28216), .Y (n_29747));
AOI21X1 g108699(.A0 (n_34712), .A1 (n_29049), .B0 (n_28942), .Y(n_29746));
AOI21X1 g108700(.A0 (n_34712), .A1 (n_29396), .B0 (n_28941), .Y(n_29745));
NAND2X1 g108703(.A (n_28932), .B (n_28509), .Y (n_29744));
NAND2X1 g108704(.A (n_28930), .B (n_28951), .Y (n_29743));
NAND2X1 g108710(.A (n_28925), .B (n_28506), .Y (n_29742));
NAND2X1 g108711(.A (n_28923), .B (n_28950), .Y (n_29741));
NAND2X1 g108727(.A (n_27175), .B (n_29239), .Y (n_29740));
NAND3X1 g107008(.A (n_28713), .B (n_28730), .C (n_28740), .Y(n_29738));
NAND2X1 g107010(.A (n_29236), .B (n_13192), .Y (n_29737));
NAND2X1 g108861(.A (n_28214), .B (n_28013), .Y (n_29736));
NAND3X1 g107087(.A (n_9073), .B (n_22104), .C (n_28705), .Y(n_29734));
NOR2X1 g109027(.A (n_29233), .B (n_29224), .Y (n_29733));
NOR2X1 g109028(.A (n_29227), .B (n_28778), .Y (n_29732));
AOI21X1 g107113(.A0 (n_30171), .A1 (n_29719), .B0 (n_28773), .Y(n_29730));
NAND2X1 g109102(.A (n_30171), .B (n_28759), .Y (n_29727));
AOI21X1 g107141(.A0 (n_29693), .A1 (n_15038), .B0 (n_29725), .Y(n_29726));
NAND2X1 g109172(.A (n_29241), .B (n_28690), .Y (n_29724));
AOI21X1 g107152(.A0 (n_14678), .A1 (n_34220), .B0 (n_29725), .Y(n_29723));
NAND4X1 g107158(.A (n_32890), .B (n_10606), .C (n_32891), .D(n_28096), .Y (n_29722));
NAND2X1 g107162(.A (n_29258), .B (n_22474), .Y (n_29721));
AOI21X1 g107167(.A0 (n_29719), .A1 (n_13952), .B0 (n_22846), .Y(n_29720));
AOI21X1 g107168(.A0 (n_29257), .A1 (n_30636), .B0 (n_29259), .Y(n_29718));
NOR2X1 g109274(.A (n_9120), .B (n_29226), .Y (n_29717));
NOR2X1 g109287(.A (n_9079), .B (n_29229), .Y (n_29716));
AOI21X1 g107205(.A0 (n_10277), .A1 (n_28581), .B0 (n_16415), .Y(n_29715));
AOI21X1 g107209(.A0 (n_10746), .A1 (n_28602), .B0 (n_31081), .Y(n_29714));
NAND2X1 g107224(.A (n_29148), .B (n_31965), .Y (n_35431));
NOR2X1 g107234(.A (n_29120), .B (n_29151), .Y (n_29711));
NOR2X1 g107236(.A (n_29119), .B (n_29145), .Y (n_29710));
OAI21X1 g107252(.A0 (n_28627), .A1 (n_28045), .B0 (n_31174), .Y(n_29709));
NAND4X1 g107261(.A (n_15249), .B (n_27892), .C (n_27891), .D(n_27946), .Y (n_29708));
NAND4X1 g107263(.A (n_15005), .B (n_27410), .C (n_27435), .D(n_27416), .Y (n_29707));
OAI21X1 g109464(.A0 (n_28141), .A1 (n_8664), .B0 (n_27797), .Y(n_29706));
NAND2X1 g109475(.A (n_28822), .B (n_28289), .Y (n_29705));
NAND2X1 g109478(.A (n_28818), .B (n_27824), .Y (n_29704));
NAND2X1 g109479(.A (n_28814), .B (n_28285), .Y (n_29703));
NAND4X1 g107292(.A (n_20477), .B (n_24594), .C (n_27506), .D(n_25998), .Y (n_29702));
NAND4X1 g107313(.A (n_20463), .B (n_24571), .C (n_27512), .D(n_25997), .Y (n_29701));
NAND2X1 g109563(.A (n_28138), .B (n_28485), .Y (n_29700));
NAND2X1 g107320(.A (n_30836), .B (n_29697), .Y (n_29699));
NAND2X1 g107321(.A (n_27632), .B (n_29697), .Y (n_35703));
NAND2X1 g107322(.A (n_29695), .B (n_29697), .Y (n_35425));
NAND2X1 g107331(.A (n_29694), .B (n_29693), .Y (n_30079));
NOR2X1 g106381(.A (n_28667), .B (n_11197), .Y (n_29692));
NAND2X1 g107336(.A (n_34220), .B (n_29690), .Y (n_30068));
NAND2X1 g107340(.A (n_8284), .B (n_29686), .Y (n_29689));
NAND2X1 g107341(.A (n_28710), .B (n_27109), .Y (n_29688));
NAND2X1 g107342(.A (n_29341), .B (n_29686), .Y (n_29687));
NAND2X1 g107344(.A (n_29684), .B (n_29686), .Y (n_29685));
AOI21X1 g107359(.A0 (n_34770), .A1 (n_28927), .B0 (n_25449), .Y(n_29683));
OAI21X1 g107361(.A0 (n_28117), .A1 (n_29681), .B0 (n_10383), .Y(n_29682));
NAND4X1 g107370(.A (n_14825), .B (n_27421), .C (n_27448), .D(n_27419), .Y (n_29680));
NAND4X1 g107395(.A (n_20491), .B (n_26380), .C (n_27409), .D(n_24252), .Y (n_29679));
OAI21X1 g107396(.A0 (n_28090), .A1 (n_29681), .B0 (n_10444), .Y(n_29678));
OAI21X1 g107405(.A0 (n_28088), .A1 (n_29681), .B0 (n_10381), .Y(n_29677));
NOR2X1 g107408(.A (n_9392), .B (n_28745), .Y (n_29676));
NAND2X1 g107423(.A (n_28724), .B (n_29505), .Y (n_35426));
NAND4X1 g107433(.A (n_20393), .B (n_26379), .C (n_27403), .D(n_24209), .Y (n_29674));
NOR2X1 g107436(.A (n_10373), .B (n_28744), .Y (n_29673));
OAI21X1 g107441(.A0 (n_9881), .A1 (n_31019), .B0 (n_28683), .Y(n_29672));
NOR2X1 g109894(.A (n_9117), .B (n_28693), .Y (n_29671));
NAND2X1 g107454(.A (n_28712), .B (n_22133), .Y (n_29670));
NOR2X1 g106439(.A (n_28348), .B (n_28622), .Y (n_29669));
NAND2X1 g107464(.A (n_28737), .B (n_33792), .Y (n_30094));
NAND2X1 g107465(.A (n_28736), .B (n_29667), .Y (n_32851));
OAI21X1 g107468(.A0 (n_28049), .A1 (n_13434), .B0 (n_29666), .Y(n_30087));
NAND2X1 g107470(.A (n_32313), .B (n_32314), .Y (n_29665));
NOR2X1 g107480(.A (n_10385), .B (n_28743), .Y (n_29664));
NOR2X1 g109958(.A (n_9102), .B (n_28692), .Y (n_29663));
NAND2X1 g107507(.A (n_28723), .B (n_29662), .Y (n_29962));
NAND2X1 g107519(.A (n_28722), .B (n_22117), .Y (n_29661));
NAND2X1 g107521(.A (n_6693), .B (n_28756), .Y (n_29660));
NAND2X1 g107522(.A (n_6606), .B (n_28755), .Y (n_29659));
NAND2X1 g107544(.A (n_6595), .B (n_28753), .Y (n_29658));
NAND2X1 g107549(.A (n_28695), .B (n_22107), .Y (n_29657));
NAND2X1 g107559(.A (n_28729), .B (n_22105), .Y (n_29656));
OAI21X1 g107562(.A0 (n_28533), .A1 (n_8333), .B0 (n_22109), .Y(n_29655));
NOR2X1 g107570(.A (n_27555), .B (n_28336), .Y (n_29654));
NAND4X1 g107571(.A (n_27494), .B (n_27972), .C (n_20207), .D(n_10823), .Y (n_29653));
NOR2X1 g107574(.A (n_28545), .B (n_28565), .Y (n_29652));
NAND2X1 g107575(.A (n_27524), .B (n_28563), .Y (n_29651));
NAND4X1 g107576(.A (n_27444), .B (n_27840), .C (n_21728), .D(n_27442), .Y (n_29650));
NAND2X1 g107579(.A (n_28584), .B (n_31590), .Y (n_29649));
NAND4X1 g107587(.A (n_28461), .B (n_27971), .C (n_10042), .D(n_18910), .Y (n_29648));
NAND2X1 g107588(.A (n_28579), .B (n_28578), .Y (n_29647));
NAND3X1 g107590(.A (n_27868), .B (n_27944), .C (n_27897), .Y(n_29646));
NAND3X1 g107593(.A (n_28573), .B (n_27934), .C (n_20386), .Y(n_29645));
NAND2X1 g107597(.A (n_28567), .B (n_31912), .Y (n_29644));
NAND4X1 g107602(.A (n_28575), .B (n_26845), .C (n_15336), .D(n_26821), .Y (n_29643));
NAND3X1 g107610(.A (n_11143), .B (n_27496), .C (n_27992), .Y(n_29642));
NAND4X1 g107621(.A (n_28463), .B (n_27981), .C (n_10048), .D(n_9505), .Y (n_29641));
OAI21X1 g107627(.A0 (n_27943), .A1 (n_26265), .B0 (n_33123), .Y(n_29640));
OAI21X1 g107628(.A0 (n_27898), .A1 (n_26623), .B0 (n_24695), .Y(n_29639));
NAND4X1 g106520(.A (n_6556), .B (n_7165), .C (n_27567), .D (n_27809),.Y (n_29637));
AOI21X1 g107630(.A0 (n_28048), .A1 (n_28242), .B0 (n_31041), .Y(n_29636));
OAI21X1 g107634(.A0 (n_27880), .A1 (n_27272), .B0 (n_33123), .Y(n_29635));
OAI21X1 g107636(.A0 (n_27899), .A1 (n_25182), .B0 (n_29633), .Y(n_29634));
OAI21X1 g107641(.A0 (n_27857), .A1 (n_24822), .B0 (n_29633), .Y(n_29632));
NAND2X1 g107657(.A (n_29620), .B (n_28864), .Y (n_29630));
NAND2X1 g107661(.A (n_9503), .B (n_29601), .Y (n_35409));
NAND2X1 g107664(.A (n_9503), .B (n_33783), .Y (n_29627));
NAND2X1 g107668(.A (n_29613), .B (n_29619), .Y (n_29626));
NAND2X1 g107669(.A (n_29611), .B (n_30563), .Y (n_29625));
NAND2X1 g107671(.A (n_29623), .B (n_30563), .Y (n_29624));
NAND2X1 g107672(.A (n_29606), .B (n_29008), .Y (n_29622));
NAND2X1 g107674(.A (n_29620), .B (n_29619), .Y (n_29621));
NAND2X1 g107676(.A (n_33377), .B (n_28485), .Y (n_29618));
NAND2X1 g107684(.A (n_29615), .B (n_34709), .Y (n_29616));
NAND2X1 g107687(.A (n_29613), .B (n_28808), .Y (n_35088));
NAND2X1 g107688(.A (n_29611), .B (n_30197), .Y (n_29612));
NAND2X2 g107690(.A (n_29623), .B (n_27326), .Y (n_29610));
NAND2X1 g107692(.A (n_29606), .B (n_29604), .Y (n_29607));
NAND2X1 g107695(.A (n_29620), .B (n_29604), .Y (n_29605));
NAND2X1 g107700(.A (n_29601), .B (n_33785), .Y (n_35408));
NAND2X1 g107711(.A (n_29595), .B (n_27747), .Y (n_29598));
NAND2X1 g107713(.A (n_28589), .B (n_31912), .Y (n_29597));
NAND2X1 g107731(.A (n_29595), .B (n_28441), .Y (n_29596));
NAND4X1 g107742(.A (n_26981), .B (n_27875), .C (n_27823), .D(n_26897), .Y (n_29594));
NAND3X1 g107745(.A (n_27810), .B (n_27874), .C (n_27694), .Y(n_29593));
NOR2X1 g107755(.A (n_27472), .B (n_28582), .Y (n_29592));
NOR2X1 g107764(.A (n_29975), .B (n_8718), .Y (n_29591));
NAND2X2 g107766(.A (n_29595), .B (n_27770), .Y (n_29590));
NAND4X1 g107772(.A (n_26913), .B (n_27872), .C (n_27821), .D(n_26895), .Y (n_29589));
NAND2X1 g107791(.A (n_29595), .B (n_13274), .Y (n_29588));
NAND2X1 g107793(.A (n_8284), .B (n_29585), .Y (n_29587));
NAND2X1 g107794(.A (n_26255), .B (n_29585), .Y (n_29586));
NAND2X1 g107795(.A (n_29695), .B (n_29585), .Y (n_29584));
NAND2X1 g107796(.A (n_28577), .B (n_31641), .Y (n_29583));
NAND2X1 g107797(.A (n_8284), .B (n_29578), .Y (n_29582));
NAND2X1 g107798(.A (n_26255), .B (n_29578), .Y (n_29580));
NAND2X1 g107799(.A (n_29427), .B (n_29578), .Y (n_29577));
NAND2X1 g107805(.A (n_29576), .B (n_29572), .Y (n_30303));
NAND2X1 g107806(.A (n_29562), .B (n_17968), .Y (n_29575));
NAND2X1 g107808(.A (n_29556), .B (n_14439), .Y (n_29574));
NAND2X1 g107809(.A (n_29572), .B (n_15407), .Y (n_29573));
NOR2X1 g107813(.A (n_28592), .B (n_26435), .Y (n_29571));
NOR2X1 g107815(.A (n_28591), .B (n_27867), .Y (n_29570));
NAND2X1 g107818(.A (n_29568), .B (n_29567), .Y (n_29569));
NAND2X1 g107823(.A (n_29565), .B (n_33738), .Y (n_29566));
AOI21X1 g106602(.A0 (n_9384), .A1 (n_28282), .B0 (n_34676), .Y(n_29563));
NAND2X1 g107829(.A (n_29562), .B (n_35736), .Y (n_30297));
NOR2X1 g107832(.A (n_28527), .B (n_10588), .Y (n_29561));
NAND2X1 g107834(.A (n_28999), .B (n_28874), .Y (n_29560));
NAND2X2 g107836(.A (n_30454), .B (n_32935), .Y (n_29559));
NAND2X1 g107839(.A (n_30171), .B (n_28052), .Y (n_29558));
NAND2X1 g107842(.A (n_29556), .B (n_35816), .Y (n_29557));
NAND4X1 g107843(.A (n_26912), .B (n_27865), .C (n_27818), .D(n_26893), .Y (n_29555));
NOR2X1 g107852(.A (n_29553), .B (n_29011), .Y (n_29554));
NAND2X1 g107854(.A (n_29551), .B (n_29567), .Y (n_29552));
NAND2X1 g107857(.A (n_28624), .B (n_29505), .Y (n_32144));
NAND2X1 g107858(.A (n_29551), .B (n_29547), .Y (n_29548));
NAND2X1 g107859(.A (n_29568), .B (n_29547), .Y (n_32598));
NAND2X1 g107867(.A (n_29544), .B (n_29545), .Y (n_30288));
NAND4X1 g107876(.A (n_26979), .B (n_27879), .C (n_27826), .D(n_26899), .Y (n_29543));
NAND2X1 g107882(.A (n_28604), .B (n_29505), .Y (n_32153));
NAND4X1 g107884(.A (n_28644), .B (n_26360), .C (n_26217), .D(n_26250), .Y (n_29540));
NAND2X1 g107887(.A (n_29535), .B (n_29411), .Y (n_29539));
NAND2X1 g107889(.A (n_29556), .B (n_35473), .Y (n_29538));
NAND2X1 g107890(.A (n_29556), .B (n_26234), .Y (n_29537));
NAND2X1 g107892(.A (n_29535), .B (n_8954), .Y (n_29536));
NAND2X1 g107896(.A (n_29535), .B (n_29405), .Y (n_29534));
NAND2X1 g107897(.A (n_29535), .B (n_30636), .Y (n_29533));
NAND2X1 g107901(.A (n_29526), .B (n_33991), .Y (n_29532));
NAND3X1 g107904(.A (n_27921), .B (n_26963), .C (n_27919), .Y(n_29530));
NAND3X1 g107909(.A (n_27955), .B (n_22124), .C (n_27958), .Y(n_29528));
NAND2X1 g107910(.A (n_29562), .B (n_28053), .Y (n_30295));
NAND2X1 g107914(.A (n_29526), .B (n_28158), .Y (n_29527));
NAND2X1 g107915(.A (n_29526), .B (n_29523), .Y (n_29524));
NAND3X1 g107918(.A (n_27927), .B (n_22114), .C (n_27925), .Y(n_29522));
NAND2X1 g107919(.A (n_29562), .B (n_35500), .Y (n_29521));
NAND4X1 g107930(.A (n_32163), .B (n_32164), .C (n_27736), .D(n_23156), .Y (n_29520));
NOR2X1 g107938(.A (n_9907), .B (n_28631), .Y (n_29519));
OAI21X1 g107943(.A0 (n_27850), .A1 (n_8321), .B0 (n_22849), .Y(n_29518));
NAND3X1 g107946(.A (n_27348), .B (n_27978), .C (n_27695), .Y(n_29517));
NAND4X1 g106648(.A (n_14180), .B (n_13743), .C (n_28993), .D(n_27562), .Y (n_29516));
OAI21X1 g107947(.A0 (n_8778), .A1 (n_35012), .B0 (n_28623), .Y(n_29515));
NAND4X1 g107950(.A (n_25768), .B (n_23433), .C (n_27816), .D(n_25144), .Y (n_29514));
OAI21X1 g107952(.A0 (n_27862), .A1 (n_8321), .B0 (n_22848), .Y(n_29513));
NAND3X1 g107957(.A (n_10179), .B (n_27492), .C (n_27959), .Y(n_29511));
NOR2X1 g107969(.A (n_9080), .B (n_28529), .Y (n_29510));
NAND3X1 g107974(.A (n_9062), .B (n_20712), .C (n_27896), .Y(n_29509));
NAND3X1 g106662(.A (n_7772), .B (n_27855), .C (n_7165), .Y (n_32879));
NAND2X1 g107976(.A (n_28616), .B (n_29505), .Y (n_29507));
NAND2X1 g107977(.A (n_28614), .B (n_29505), .Y (n_29506));
OAI21X1 g106664(.A0 (n_29438), .A1 (n_8687), .B0 (n_30063), .Y(n_29504));
NAND4X1 g106666(.A (n_14551), .B (n_14158), .C (n_28954), .D(n_27560), .Y (n_29503));
NAND4X1 g107989(.A (n_32138), .B (n_32139), .C (n_27729), .D(n_23148), .Y (n_29502));
NAND3X1 g107991(.A (n_10127), .B (n_27491), .C (n_27928), .Y(n_29501));
NAND4X1 g106672(.A (n_35046), .B (n_14320), .C (n_28974), .D(n_27561), .Y (n_29500));
NAND2X1 g108000(.A (n_28638), .B (n_29133), .Y (n_29498));
NAND2X1 g108004(.A (n_28625), .B (n_26570), .Y (n_30027));
NOR2X1 g108010(.A (n_28042), .B (n_28646), .Y (n_29496));
NOR2X1 g108012(.A (n_28041), .B (n_28645), .Y (n_29495));
NAND4X1 g108018(.A (n_32103), .B (n_18405), .C (n_32104), .D(n_27321), .Y (n_29494));
OAI21X1 g108027(.A0 (n_27852), .A1 (n_9625), .B0 (n_15337), .Y(n_29493));
AOI21X1 g108028(.A0 (n_29103), .A1 (n_29061), .B0 (n_15027), .Y(n_29491));
OAI21X1 g108030(.A0 (n_27851), .A1 (n_9625), .B0 (n_15378), .Y(n_29490));
AOI21X1 g108031(.A0 (n_29100), .A1 (n_29061), .B0 (n_15024), .Y(n_29489));
NAND2X1 g108034(.A (n_28639), .B (n_13662), .Y (n_30321));
OAI21X1 g106689(.A0 (n_8228), .A1 (n_29486), .B0 (n_28526), .Y(n_29487));
NAND2X1 g108039(.A (n_28635), .B (n_28554), .Y (n_29845));
NAND2X1 g108042(.A (n_28626), .B (n_28549), .Y (n_30342));
NAND3X1 g108049(.A (n_28574), .B (n_26915), .C (n_26930), .Y(n_29485));
NAND2X1 g108053(.A (n_28609), .B (n_8316), .Y (n_29484));
OAI21X1 g106696(.A0 (n_8856), .A1 (n_30731), .B0 (n_28448), .Y(n_29482));
NOR2X1 g108063(.A (n_27894), .B (n_28525), .Y (n_29481));
NAND2X1 g108072(.A (n_28590), .B (n_29480), .Y (n_30298));
OAI21X1 g106704(.A0 (n_8699), .A1 (n_35012), .B0 (n_28440), .Y(n_29479));
NAND2X2 g108080(.A (n_28607), .B (n_29478), .Y (n_29831));
NAND4X1 g108081(.A (n_27346), .B (n_10586), .C (n_27784), .D(n_27324), .Y (n_29477));
OAI21X1 g106708(.A0 (n_9770), .A1 (n_30893), .B0 (n_28522), .Y(n_29476));
NAND4X1 g106709(.A (n_15306), .B (n_34423), .C (n_27636), .D(n_14521), .Y (n_29475));
OAI21X1 g108102(.A0 (n_27866), .A1 (n_30792), .B0 (n_6506), .Y(n_29474));
NAND2X1 g108103(.A (n_28670), .B (n_28611), .Y (n_29473));
OAI21X1 g108105(.A0 (n_27853), .A1 (n_30792), .B0 (n_6488), .Y(n_29472));
CLKBUFX1 gbuf_d_344(.A(n_28674), .Y(d_out_344));
CLKBUFX1 gbuf_q_344(.A(q_in_344), .Y(P2_reg1[2]));
NAND4X1 g108106(.A (n_35918), .B (n_27400), .C (n_35919), .D(n_26432), .Y (n_29471));
NAND2X1 g108118(.A (n_28903), .B (n_7967), .Y (n_29470));
NAND2X1 g108124(.A (n_28032), .B (n_28331), .Y (n_29468));
NOR2X1 g108125(.A (n_27813), .B (n_28330), .Y (n_29467));
NAND2X1 g108136(.A (n_28333), .B (n_30421), .Y (n_29466));
NOR2X1 g108140(.A (n_19526), .B (n_28321), .Y (n_29465));
AOI21X1 g108153(.A0 (n_28293), .A1 (n_28273), .B0 (n_31041), .Y(n_29464));
NOR2X1 g108156(.A (n_10084), .B (n_28836), .Y (n_29462));
NAND4X1 g108157(.A (n_28803), .B (n_27783), .C (n_10044), .D(n_9622), .Y (n_29461));
AOI21X1 g108159(.A0 (n_28292), .A1 (n_28244), .B0 (n_31041), .Y(n_29460));
AOI21X1 g108165(.A0 (n_29068), .A1 (n_28940), .B0 (n_26802), .Y(n_32612));
AOI21X1 g108173(.A0 (n_9003), .A1 (n_28934), .B0 (n_26784), .Y(n_29458));
NAND2X1 g108200(.A (n_33509), .B (n_29455), .Y (n_29457));
NAND2X1 g108213(.A (n_28329), .B (n_25980), .Y (n_29454));
NAND2X1 g108214(.A (n_33498), .B (n_29455), .Y (n_29453));
AOI21X1 g108215(.A0 (n_15254), .A1 (n_22821), .B0 (n_28349), .Y(n_29451));
NAND4X1 g108219(.A (n_15006), .B (n_26233), .C (n_27618), .D(n_26239), .Y (n_29450));
AOI21X1 g108226(.A0 (n_15256), .A1 (n_22821), .B0 (n_28346), .Y(n_35382));
NOR2X1 g108245(.A (n_28185), .B (n_28307), .Y (n_29447));
CLKBUFX1 gbuf_d_345(.A(n_28763), .Y(d_out_345));
CLKBUFX1 gbuf_q_345(.A(q_in_345), .Y(P3_reg1[3]));
NAND2X1 g108250(.A (n_29850), .B (n_29445), .Y (n_29446));
CLKBUFX1 gbuf_d_346(.A(n_28764), .Y(d_out_346));
CLKBUFX1 gbuf_q_346(.A(q_in_346), .Y(P2_reg2[3]));
CLKBUFX1 gbuf_d_347(.A(n_28760), .Y(d_out_347));
CLKBUFX1 gbuf_q_347(.A(q_in_347), .Y(n_13358));
CLKBUFX1 gbuf_d_348(.A(n_28830), .Y(d_out_348));
CLKBUFX1 gbuf_q_348(.A(q_in_348), .Y(P2_reg3[4]));
CLKBUFX1 gbuf_d_349(.A(n_28675), .Y(d_out_349));
CLKBUFX1 gbuf_q_349(.A(q_in_349), .Y(n_10435));
CLKBUFX1 gbuf_d_350(.A(n_28673), .Y(d_out_350));
CLKBUFX1 gbuf_q_350(.A(q_in_350), .Y(P2_reg2[2]));
CLKBUFX1 gbuf_d_351(.A(n_28733), .Y(d_out_351));
CLKBUFX1 gbuf_q_351(.A(q_in_351), .Y(n_9634));
NOR2X1 g108264(.A (n_28316), .B (n_28834), .Y (n_29444));
NAND2X1 g108265(.A (n_28314), .B (n_28833), .Y (n_29443));
NAND4X1 g108278(.A (n_28765), .B (n_27248), .C (n_24797), .D(n_27655), .Y (n_29442));
NAND2X1 g108280(.A (n_29568), .B (n_29440), .Y (n_29441));
OAI21X1 g106789(.A0 (n_29438), .A1 (n_26052), .B0 (n_26457), .Y(n_29439));
NAND4X1 g108284(.A (n_20278), .B (n_27775), .C (n_27773), .D(n_27330), .Y (n_29437));
NAND2X1 g108285(.A (n_28312), .B (n_28317), .Y (n_29436));
NAND2X1 g108286(.A (n_29841), .B (n_30557), .Y (n_29435));
NAND2X1 g108304(.A (n_29819), .B (n_30559), .Y (n_29433));
NAND2X1 g108309(.A (n_8284), .B (n_29429), .Y (n_29432));
NAND2X1 g108310(.A (n_29430), .B (n_29429), .Y (n_29431));
NAND2X1 g108311(.A (n_29427), .B (n_29429), .Y (n_29428));
NAND2X1 g108324(.A (n_29425), .B (n_33738), .Y (n_29426));
NAND2X1 g108346(.A (n_29422), .B (n_30184), .Y (n_29423));
NAND2X1 g108347(.A (n_29422), .B (n_26665), .Y (n_29421));
NAND2X1 g108348(.A (n_29422), .B (n_30180), .Y (n_29419));
NAND2X1 g108351(.A (n_28395), .B (n_29505), .Y (n_32172));
NAND2X1 g108352(.A (n_29551), .B (n_29440), .Y (n_29417));
NOR2X1 g108358(.A (n_28180), .B (n_28301), .Y (n_35383));
NAND2X1 g108365(.A (n_29425), .B (n_29405), .Y (n_29415));
NAND3X1 g108371(.A (n_28496), .B (n_25100), .C (n_14923), .Y(n_29413));
NAND2X1 g108387(.A (n_29408), .B (n_29411), .Y (n_29412));
NAND4X1 g108390(.A (n_14820), .B (n_26245), .C (n_27627), .D(n_26243), .Y (n_29410));
NAND2X1 g108393(.A (n_29408), .B (n_8954), .Y (n_29409));
NAND2X1 g108394(.A (n_29408), .B (n_29405), .Y (n_29406));
NAND2X1 g108395(.A (n_29408), .B (n_29955), .Y (n_29404));
NAND2X1 g108411(.A (n_29401), .B (n_29523), .Y (n_29400));
NOR2X1 g108415(.A (n_9141), .B (n_28839), .Y (n_29399));
AOI21X1 g106852(.A0 (n_9425), .A1 (n_28167), .B0 (n_30702), .Y(n_29398));
AOI21X1 g108425(.A0 (n_29396), .A1 (n_30557), .B0 (n_21371), .Y(n_32611));
NOR2X1 g108426(.A (n_9114), .B (n_28838), .Y (n_29395));
NOR2X1 g108428(.A (n_9108), .B (n_28837), .Y (n_29394));
AOI22X1 g108430(.A0 (n_29392), .A1 (n_26288), .B0 (n_20304), .B1(n_19501), .Y (n_32887));
AOI21X1 g108441(.A0 (n_29390), .A1 (n_29040), .B0 (n_21366), .Y(n_29391));
OAI21X1 g108443(.A0 (n_28221), .A1 (n_29388), .B0 (n_20737), .Y(n_29389));
OAI21X1 g108445(.A0 (n_28218), .A1 (n_33807), .B0 (n_19603), .Y(n_29387));
OAI21X1 g108452(.A0 (n_28203), .A1 (n_29381), .B0 (n_22122), .Y(n_29385));
NAND2X1 g108461(.A (n_28414), .B (n_29505), .Y (n_29384));
NAND2X1 g108473(.A (n_28402), .B (n_27844), .Y (n_29383));
OAI21X1 g108478(.A0 (n_28197), .A1 (n_29381), .B0 (n_22113), .Y(n_29382));
NAND2X1 g108480(.A (n_28378), .B (n_26396), .Y (n_29380));
NOR2X1 g108481(.A (n_9476), .B (n_28835), .Y (n_29379));
INVX2 g108483(.A (n_29378), .Y (n_30514));
INVX1 g108491(.A (n_29893), .Y (n_29376));
NAND2X1 g108501(.A (n_28457), .B (n_28430), .Y (n_29374));
INVX1 g108504(.A (n_29033), .Y (n_29373));
OAI21X1 g108507(.A0 (n_28220), .A1 (n_30355), .B0 (n_28482), .Y(n_29372));
OAI21X1 g108510(.A0 (n_28210), .A1 (n_29388), .B0 (n_21215), .Y(n_29371));
OAI21X1 g108511(.A0 (n_28899), .A1 (n_33807), .B0 (n_19623), .Y(n_29370));
OAI21X1 g108513(.A0 (n_28201), .A1 (n_29388), .B0 (n_21200), .Y(n_29369));
OAI21X1 g108514(.A0 (n_28200), .A1 (n_29388), .B0 (n_20146), .Y(n_29368));
OAI21X1 g108515(.A0 (n_28193), .A1 (n_29388), .B0 (n_21208), .Y(n_29367));
OAI21X1 g108516(.A0 (n_18947), .A1 (n_21365), .B0 (n_28382), .Y(n_29366));
OAI21X1 g108517(.A0 (n_28191), .A1 (n_33807), .B0 (n_20135), .Y(n_29365));
NAND2X1 g108532(.A (n_28497), .B (n_14828), .Y (n_29364));
NAND2X1 g108534(.A (n_28495), .B (n_14602), .Y (n_29363));
AOI21X1 g106904(.A0 (n_28162), .A1 (n_26984), .B0 (n_8355), .Y(n_29361));
INVX1 g108542(.A (n_29359), .Y (n_29360));
NAND2X1 g108549(.A (n_28442), .B (n_13628), .Y (n_30220));
INVX1 g108555(.A (n_29357), .Y (n_29771));
INVX2 g108567(.A (n_29018), .Y (n_30203));
INVX1 g108570(.A (n_29355), .Y (n_29356));
INVX1 g108573(.A (n_29923), .Y (n_29353));
OAI21X1 g108576(.A0 (n_28222), .A1 (n_34719), .B0 (n_28510), .Y(n_29352));
OAI21X1 g108577(.A0 (n_30445), .A1 (n_27726), .B0 (n_28484), .Y(n_29350));
NAND2X1 g108579(.A (n_28428), .B (n_35057), .Y (n_29767));
AOI21X1 g106914(.A0 (n_28128), .A1 (n_26949), .B0 (n_33125), .Y(n_29348));
NAND2X2 g108585(.A (n_28415), .B (n_13487), .Y (n_30182));
INVX1 g108588(.A (n_29889), .Y (n_29347));
INVX1 g108594(.A (n_29906), .Y (n_29346));
NAND2X2 g108603(.A (n_28379), .B (n_13181), .Y (n_30165));
NAND2X1 g108610(.A (n_28437), .B (n_8316), .Y (n_29344));
NAND2X1 g108616(.A (n_28393), .B (n_19582), .Y (n_29343));
AOI21X1 g108622(.A0 (n_29341), .A1 (n_28392), .B0 (n_28474), .Y(n_29342));
NAND2X1 g108625(.A (n_19572), .B (n_28452), .Y (n_29340));
NAND2X1 g106932(.A (n_28774), .B (n_26142), .Y (n_29339));
NAND4X1 g106935(.A (n_15107), .B (n_25959), .C (n_26883), .D(n_27793), .Y (n_29338));
NAND4X1 g106936(.A (n_15103), .B (n_25915), .C (n_26860), .D(n_27769), .Y (n_29337));
OAI21X1 g108650(.A0 (n_28207), .A1 (n_10276), .B0 (n_28465), .Y(n_29332));
NAND4X1 g106939(.A (n_15109), .B (n_25870), .C (n_26831), .D(n_27752), .Y (n_29331));
INVX1 g108658(.A (n_28995), .Y (n_29330));
NAND2X1 g108666(.A (n_28477), .B (n_28418), .Y (n_29329));
OAI21X1 g108670(.A0 (n_18938), .A1 (n_25540), .B0 (n_28405), .Y(n_29328));
OAI21X1 g108675(.A0 (n_28184), .A1 (n_8677), .B0 (n_28371), .Y(n_29327));
NAND2X1 g108678(.A (n_28413), .B (n_19566), .Y (n_29326));
OAI21X1 g108684(.A0 (n_28757), .A1 (n_8352), .B0 (n_19554), .Y(n_29325));
OAI21X1 g108694(.A0 (n_28241), .A1 (n_33734), .B0 (n_19559), .Y(n_29324));
OAI21X1 g108696(.A0 (n_28245), .A1 (n_33734), .B0 (n_19553), .Y(n_29323));
OAI21X1 g108701(.A0 (n_28212), .A1 (n_10790), .B0 (n_28513), .Y(n_29321));
OAI21X1 g108702(.A0 (n_30445), .A1 (n_27715), .B0 (n_28487), .Y(n_29320));
NAND2X1 g108705(.A (n_28480), .B (n_28508), .Y (n_29319));
NAND2X1 g108706(.A (n_28024), .B (n_28507), .Y (n_29318));
OAI21X1 g108712(.A0 (n_28194), .A1 (n_10790), .B0 (n_28505), .Y(n_29317));
NAND2X1 g108713(.A (n_28019), .B (n_28504), .Y (n_29316));
NOR2X1 g108726(.A (n_27177), .B (n_28781), .Y (n_29315));
NOR2X1 g108738(.A (n_28769), .B (n_28777), .Y (n_29314));
NOR2X1 g108740(.A (n_28768), .B (n_28776), .Y (n_29313));
NAND3X1 g106989(.A (n_12380), .B (n_25253), .C (n_28130), .Y(n_29312));
NOR2X1 g108758(.A (n_28751), .B (n_28779), .Y (n_29311));
NOR2X1 g108759(.A (n_28750), .B (n_27731), .Y (n_29310));
NOR2X1 g108762(.A (n_28746), .B (n_27730), .Y (n_29309));
NOR2X1 g108801(.A (n_9172), .B (n_28775), .Y (n_29308));
NOR2X1 g108802(.A (n_14162), .B (n_29302), .Y (n_29307));
NOR2X1 g108807(.A (n_9172), .B (n_28771), .Y (n_29306));
NOR2X1 g108819(.A (n_34771), .B (n_28766), .Y (n_29305));
NOR2X1 g108826(.A (n_29302), .B (n_27158), .Y (n_29303));
NAND2X1 g108929(.A (n_28772), .B (n_30559), .Y (n_32560));
NOR2X1 g108970(.A (n_27245), .B (n_28694), .Y (n_29300));
INVX1 g107123(.A (n_30462), .Y (n_29729));
NAND4X1 g107125(.A (n_15094), .B (n_25941), .C (n_26871), .D(n_27778), .Y (n_29298));
NAND2X1 g109106(.A (n_30171), .B (n_28181), .Y (n_29297));
NAND2X1 g109135(.A (n_29295), .B (n_30109), .Y (n_35147));
NOR2X1 g109170(.A (n_28780), .B (n_28131), .Y (n_29294));
NAND3X1 g109171(.A (n_28691), .B (n_26529), .C (n_27054), .Y(n_29293));
NOR2X1 g109173(.A (n_27250), .B (n_28689), .Y (n_29292));
NAND3X1 g109177(.A (n_28688), .B (n_25727), .C (n_26182), .Y(n_29291));
OAI21X1 g109182(.A0 (n_28141), .A1 (n_9626), .B0 (n_25547), .Y(n_29290));
NAND3X1 g109184(.A (n_28831), .B (n_25204), .C (n_15344), .Y(n_29288));
AOI22X1 g107170(.A0 (n_29250), .A1 (n_8954), .B0 (n_22469), .B1(n_21328), .Y (n_29287));
OAI21X1 g107174(.A0 (n_28135), .A1 (n_29285), .B0 (n_6727), .Y(n_29286));
OAI21X1 g107176(.A0 (n_28133), .A1 (n_33350), .B0 (n_6671), .Y(n_29284));
NAND2X1 g107179(.A (n_6496), .B (n_28326), .Y (n_29283));
OAI21X1 g107181(.A0 (n_28129), .A1 (n_31958), .B0 (n_6620), .Y(n_29282));
OAI21X1 g109322(.A0 (n_28147), .A1 (n_8668), .B0 (n_28255), .Y(n_29279));
OAI21X1 g109332(.A0 (n_28142), .A1 (n_9625), .B0 (n_15164), .Y(n_29278));
OAI21X1 g109336(.A0 (n_28698), .A1 (n_26748), .B0 (n_15157), .Y(n_29277));
INVX1 g109345(.A (n_29275), .Y (n_29276));
INVX1 g109357(.A (n_29272), .Y (n_29273));
INVX1 g109368(.A (n_29270), .Y (n_30449));
INVX1 g109381(.A (n_29269), .Y (n_29712));
INVX2 g109391(.A (n_29268), .Y (n_30122));
OAI21X1 g107246(.A0 (n_28077), .A1 (n_34336), .B0 (n_10478), .Y(n_29267));
NOR2X1 g109422(.A (n_26591), .B (n_28749), .Y (n_29265));
AOI21X1 g109480(.A0 (n_28826), .A1 (n_34694), .B0 (n_28284), .Y(n_29262));
NAND3X1 g109503(.A (n_20697), .B (n_27572), .C (n_25753), .Y(n_29261));
NOR2X1 g109554(.A (n_28147), .B (n_26748), .Y (n_29260));
NOR2X1 g107326(.A (n_28676), .B (n_29172), .Y (n_29259));
NAND2X1 g107327(.A (n_29257), .B (n_33738), .Y (n_29258));
NAND2X1 g107343(.A (n_29254), .B (n_28158), .Y (n_29256));
NAND2X1 g107345(.A (n_29254), .B (n_29253), .Y (n_29255));
NAND2X1 g107357(.A (n_29257), .B (n_29405), .Y (n_29252));
NAND2X1 g107369(.A (n_29250), .B (n_8966), .Y (n_29251));
NAND2X1 g107376(.A (n_29250), .B (n_29955), .Y (n_35298));
NAND2X1 g107375(.A (n_29250), .B (n_29405), .Y (n_29248));
NAND2X1 g109713(.A (n_28254), .B (n_25756), .Y (n_29247));
OAI21X1 g107407(.A0 (n_8581), .A1 (n_30527), .B0 (n_28169), .Y(n_29244));
NOR2X1 g109857(.A (n_27028), .B (n_28143), .Y (n_29243));
NOR2X1 g107450(.A (n_28157), .B (n_28123), .Y (n_29242));
NOR2X1 g109899(.A (n_27566), .B (n_28134), .Y (n_29241));
NAND2X1 g109945(.A (n_27101), .B (n_28137), .Y (n_29240));
NOR2X1 g109957(.A (n_9094), .B (n_28132), .Y (n_29239));
NAND2X1 g107496(.A (n_28152), .B (n_8966), .Y (n_29238));
NOR2X1 g107514(.A (n_7071), .B (n_28175), .Y (n_29236));
AOI21X1 g107527(.A0 (n_27520), .A1 (n_30836), .B0 (n_22475), .Y(n_29235));
AOI21X1 g107533(.A0 (n_28721), .A1 (n_29955), .B0 (n_28156), .Y(n_29234));
NAND2X1 g110132(.A (n_28160), .B (n_15287), .Y (n_29233));
NAND2X1 g107551(.A (n_6739), .B (n_28150), .Y (n_29232));
NAND2X1 g110174(.A (n_28166), .B (n_19862), .Y (n_29229));
AND2X1 g110190(.A (n_28163), .B (n_27623), .Y (n_29228));
NAND2X1 g110194(.A (n_28161), .B (n_19882), .Y (n_29227));
OAI21X1 g110199(.A0 (n_27553), .A1 (n_33734), .B0 (n_19883), .Y(n_29226));
NAND2X1 g107583(.A (n_28068), .B (n_30421), .Y (n_29225));
OAI21X1 g110224(.A0 (n_27553), .A1 (n_28747), .B0 (n_27633), .Y(n_29224));
NAND3X1 g107592(.A (n_28067), .B (n_27437), .C (n_21331), .Y(n_29223));
NAND3X1 g107605(.A (n_19658), .B (n_21361), .C (n_27490), .Y(n_29222));
NAND2X1 g107607(.A (n_33546), .B (n_29192), .Y (n_29221));
OAI21X1 g107609(.A0 (n_27513), .A1 (n_27795), .B0 (n_31771), .Y(n_29220));
NAND2X1 g107616(.A (n_33546), .B (n_29188), .Y (n_29219));
NAND2X1 g107625(.A (n_33546), .B (n_29178), .Y (n_29218));
OAI21X1 g107629(.A0 (n_27450), .A1 (n_25929), .B0 (n_33123), .Y(n_29217));
AOI21X1 g107631(.A0 (n_27438), .A1 (n_26762), .B0 (n_8355), .Y(n_29216));
AOI21X1 g107632(.A0 (n_27418), .A1 (n_26759), .B0 (n_29769), .Y(n_29215));
OAI21X1 g107637(.A0 (n_27417), .A1 (n_24470), .B0 (n_31099), .Y(n_29214));
AOI21X1 g107638(.A0 (n_27397), .A1 (n_25902), .B0 (n_33125), .Y(n_29213));
AOI21X1 g107639(.A0 (n_27396), .A1 (n_26251), .B0 (n_8355), .Y(n_29212));
NAND2X1 g107651(.A (n_9503), .B (n_35917), .Y (n_29211));
NAND2X1 g107655(.A (n_34770), .B (n_29197), .Y (n_29209));
NAND2X1 g107662(.A (n_34770), .B (n_29201), .Y (n_29208));
NAND2X1 g107665(.A (n_9503), .B (n_29194), .Y (n_29206));
NAND2X1 g107667(.A (n_35917), .B (n_34709), .Y (n_29204));
NAND2X1 g107678(.A (n_29201), .B (n_29925), .Y (n_29202));
NAND2X1 g107685(.A (n_35917), .B (n_29199), .Y (n_29200));
NAND2X1 g107693(.A (n_29197), .B (n_28013), .Y (n_29198));
NAND2X1 g107701(.A (n_29201), .B (n_29199), .Y (n_29196));
NAND2X1 g107704(.A (n_29194), .B (n_33785), .Y (n_29195));
NAND2X1 g107709(.A (n_29192), .B (n_29191), .Y (n_29193));
NOR2X1 g107714(.A (n_25985), .B (n_28076), .Y (n_29190));
NAND2X1 g107729(.A (n_29188), .B (n_28890), .Y (n_29189));
NAND2X1 g107733(.A (n_33808), .B (n_28734), .Y (n_29187));
NOR3X1 g107735(.A (n_26124), .B (n_23754), .C (n_27359), .Y(n_29186));
NAND3X1 g107740(.A (n_28114), .B (n_27677), .C (n_27733), .Y(n_29185));
NAND4X1 g107741(.A (n_24772), .B (n_23661), .C (n_27353), .D(n_25441), .Y (n_29184));
NOR2X1 g107751(.A (n_27476), .B (n_28075), .Y (n_29183));
NAND2X1 g107765(.A (n_28568), .B (n_25968), .Y (n_29182));
OAI21X1 g107769(.A0 (n_27405), .A1 (n_26010), .B0 (n_31398), .Y(n_29181));
NAND2X1 g107781(.A (n_29178), .B (n_29191), .Y (n_29179));
NAND2X1 g107792(.A (n_33808), .B (n_27950), .Y (n_29177));
NAND3X1 g107810(.A (n_26931), .B (n_27366), .C (n_15149), .Y(n_29175));
NOR2X1 g107811(.A (n_25976), .B (n_28069), .Y (n_29174));
NOR2X1 g107820(.A (n_28536), .B (n_29172), .Y (n_29173));
NAND2X1 g107821(.A (n_29170), .B (n_33738), .Y (n_29171));
NOR2X1 g107822(.A (n_28535), .B (n_29172), .Y (n_29169));
NAND2X1 g107847(.A (n_28065), .B (n_13196), .Y (n_29168));
NOR2X1 g107860(.A (n_22528), .B (n_32299), .Y (n_29167));
NAND2X1 g107879(.A (n_29170), .B (n_29405), .Y (n_29166));
NAND4X1 g107883(.A (n_28094), .B (n_25211), .C (n_25857), .D(n_25888), .Y (n_29165));
NAND2X1 g107886(.A (n_29162), .B (n_29411), .Y (n_29164));
NAND2X1 g107891(.A (n_29162), .B (n_8954), .Y (n_29163));
NAND2X1 g107894(.A (n_29162), .B (n_29405), .Y (n_29161));
NAND2X1 g107895(.A (n_29162), .B (n_29955), .Y (n_29160));
NAND2X1 g107900(.A (n_29156), .B (n_33991), .Y (n_29159));
NAND3X1 g107903(.A (n_27430), .B (n_27429), .C (n_27428), .Y(n_29158));
NAND2X1 g107912(.A (n_29156), .B (n_29155), .Y (n_29157));
NAND2X1 g107913(.A (n_29156), .B (n_33738), .Y (n_29154));
AOI22X1 g107923(.A0 (n_28642), .A1 (n_30063), .B0 (n_9629), .B1(n_22095), .Y (n_29153));
OAI21X1 g107924(.A0 (n_27387), .A1 (n_29150), .B0 (n_22137), .Y(n_29151));
NAND4X1 g107926(.A (n_26427), .B (n_27679), .C (n_26804), .D(n_26321), .Y (n_29149));
OAI21X1 g107927(.A0 (n_8781), .A1 (n_35012), .B0 (n_28089), .Y(n_29148));
NAND4X1 g107929(.A (n_32134), .B (n_32135), .C (n_27252), .D(n_23348), .Y (n_29147));
AOI22X1 g107936(.A0 (n_28741), .A1 (n_30063), .B0 (n_9629), .B1(n_22094), .Y (n_29146));
OAI21X1 g107937(.A0 (n_27383), .A1 (n_29150), .B0 (n_22135), .Y(n_29145));
NAND4X1 g107940(.A (n_32149), .B (n_32150), .C (n_27251), .D(n_23879), .Y (n_29144));
OAI21X1 g107944(.A0 (n_29122), .A1 (n_30523), .B0 (n_22132), .Y(n_29143));
OAI21X1 g107953(.A0 (n_35627), .A1 (n_30523), .B0 (n_22130), .Y(n_29142));
NAND4X1 g107955(.A (n_32082), .B (n_24184), .C (n_32083), .D(n_25439), .Y (n_29141));
OAI21X1 g111065(.A0 (n_25587), .A1 (n_33340), .B0 (n_28127), .Y(n_29140));
NAND3X1 g107982(.A (n_9045), .B (n_27447), .C (n_21337), .Y(n_29139));
CLKBUFX1 gbuf_d_352(.A(n_28050), .Y(d_out_352));
CLKBUFX1 gbuf_q_352(.A(q_in_352), .Y(n_13337));
OAI21X1 g108017(.A0 (n_35626), .A1 (n_8678), .B0 (n_28101), .Y(n_29138));
NOR2X1 g108019(.A (n_7015), .B (n_28121), .Y (n_29136));
OAI21X1 g108029(.A0 (n_15085), .A1 (n_8614), .B0 (n_28113), .Y(n_29135));
OAI21X1 g108032(.A0 (n_15060), .A1 (n_8614), .B0 (n_28111), .Y(n_29134));
NAND2X2 g108035(.A (n_28092), .B (n_29133), .Y (n_30020));
NAND2X2 g108040(.A (n_28099), .B (n_29132), .Y (n_30013));
NAND2X2 g108043(.A (n_28086), .B (n_26570), .Y (n_30005));
AOI22X1 g106693(.A0 (n_27834), .A1 (n_30380), .B0 (n_8273), .B1(n_9387), .Y (n_29131));
NAND2X1 g108052(.A (n_28082), .B (n_8316), .Y (n_29129));
AOI21X1 g108067(.A0 (n_14610), .A1 (n_28610), .B0 (n_29000), .Y(n_29128));
INVX1 g108073(.A (n_29125), .Y (n_29127));
OAI21X1 g108088(.A0 (n_29122), .A1 (n_8678), .B0 (n_28104), .Y(n_29123));
OAI21X1 g106712(.A0 (n_33319), .A1 (n_12670), .B0 (n_14956), .Y(n_29121));
OAI21X1 g108109(.A0 (n_30445), .A1 (n_27387), .B0 (n_28108), .Y(n_29120));
OAI21X1 g108112(.A0 (n_30445), .A1 (n_27383), .B0 (n_28106), .Y(n_29119));
NOR2X1 g108120(.A (n_27814), .B (n_27876), .Y (n_29118));
NAND2X1 g108122(.A (n_26426), .B (n_27873), .Y (n_29117));
NAND4X1 g108123(.A (n_28283), .B (n_10147), .C (n_25497), .D(n_26707), .Y (n_29116));
CLKBUFX1 gbuf_d_353(.A(n_28122), .Y(d_out_353));
CLKBUFX1 gbuf_q_353(.A(q_in_353), .Y(n_3565));
NAND2X1 g108126(.A (n_27811), .B (n_27863), .Y (n_29115));
NOR2X1 g108131(.A (n_27846), .B (n_27858), .Y (n_29114));
NAND3X1 g108133(.A (n_20221), .B (n_27750), .C (n_20945), .Y(n_29113));
NOR2X1 g108139(.A (n_20090), .B (n_27845), .Y (n_29112));
NAND2X1 g108144(.A (n_27859), .B (n_31641), .Y (n_29111));
NOR2X1 g108155(.A (n_10557), .B (n_28298), .Y (n_35904));
NAND4X1 g108174(.A (n_27744), .B (n_26754), .C (n_27161), .D(n_20788), .Y (n_29109));
NAND2X1 g108180(.A (n_29098), .B (n_28864), .Y (n_29108));
NAND2X1 g108183(.A (n_29096), .B (n_28864), .Y (n_29106));
NOR2X1 g108185(.A (n_9172), .B (n_29093), .Y (n_29105));
NAND2X1 g108188(.A (n_29103), .B (n_34694), .Y (n_29104));
NAND2X1 g108191(.A (n_29100), .B (n_34694), .Y (n_29101));
NAND2X1 g108194(.A (n_29098), .B (n_29619), .Y (n_29099));
NAND2X1 g108196(.A (n_29096), .B (n_29619), .Y (n_29097));
NAND2X1 g108202(.A (n_29103), .B (n_29090), .Y (n_29092));
NAND2X1 g108205(.A (n_29100), .B (n_29090), .Y (n_29091));
NAND2X1 g108208(.A (n_29098), .B (n_29604), .Y (n_29089));
NAND2X1 g108211(.A (n_29096), .B (n_29604), .Y (n_29088));
NOR2X1 g108223(.A (n_27854), .B (n_14741), .Y (n_29086));
NAND2X1 g108230(.A (n_29083), .B (n_27089), .Y (n_29085));
CLKBUFX1 gbuf_d_354(.A(n_28168), .Y(d_out_354));
CLKBUFX1 gbuf_q_354(.A(q_in_354), .Y(P2_reg3[1]));
CLKBUFX1 gbuf_d_355(.A(n_28051), .Y(d_out_355));
CLKBUFX1 gbuf_q_355(.A(q_in_355), .Y(P3_reg1[1]));
CLKBUFX1 gbuf_d_356(.A(n_27923), .Y(d_out_356));
CLKBUFX1 gbuf_q_356(.A(q_in_356), .Y(P3_reg3[0]));
NAND2X1 g108259(.A (n_29083), .B (n_25554), .Y (n_29084));
NAND2X1 g106783(.A (n_28056), .B (n_27006), .Y (n_29082));
OAI21X1 g108279(.A0 (n_27828), .A1 (n_26166), .B0 (n_30353), .Y(n_29081));
NAND4X1 g108281(.A (n_28234), .B (n_27595), .C (n_23801), .D(n_25822), .Y (n_29080));
NAND2X1 g108299(.A (n_29083), .B (n_35054), .Y (n_29079));
NAND2X1 g108301(.A (n_27871), .B (n_31201), .Y (n_29078));
NOR2X1 g108305(.A (n_27365), .B (n_28294), .Y (n_29077));
NOR2X1 g108306(.A (n_27836), .B (n_27870), .Y (n_29076));
NAND2X1 g108308(.A (n_29083), .B (n_23578), .Y (n_29075));
NOR2X1 g108323(.A (n_28306), .B (n_29172), .Y (n_29074));
NAND2X1 g108343(.A (n_27864), .B (n_31201), .Y (n_29073));
OAI21X1 g108344(.A0 (n_26266), .A1 (n_9616), .B0 (n_28295), .Y(n_29072));
NAND3X1 g108359(.A (n_32592), .B (n_32593), .C (n_26393), .Y(n_29071));
NAND3X1 g108360(.A (n_35133), .B (n_35134), .C (n_27738), .Y(n_29070));
AOI21X1 g108367(.A0 (n_29068), .A1 (n_29067), .B0 (n_25866), .Y(n_32914));
AOI21X1 g108370(.A0 (n_29065), .A1 (n_28449), .B0 (n_25871), .Y(n_29066));
AOI21X1 g108374(.A0 (n_28493), .A1 (n_29061), .B0 (n_25070), .Y(n_29064));
AOI21X1 g108376(.A0 (n_28490), .A1 (n_29027), .B0 (n_25069), .Y(n_29063));
AOI21X1 g108378(.A0 (n_28488), .A1 (n_29061), .B0 (n_25068), .Y(n_29062));
NAND3X1 g108380(.A (n_28030), .B (n_26033), .C (n_14980), .Y(n_29060));
NAND3X1 g108382(.A (n_28028), .B (n_26030), .C (n_14982), .Y(n_29059));
AOI21X1 g108384(.A0 (n_29009), .A1 (n_28864), .B0 (n_25046), .Y(n_29058));
AOI21X1 g108385(.A0 (n_29068), .A1 (n_28481), .B0 (n_25833), .Y(n_29057));
NAND4X1 g108398(.A (n_27815), .B (n_26757), .C (n_27163), .D(n_20791), .Y (n_29056));
NAND3X1 g108401(.A (n_27801), .B (n_20198), .C (n_27799), .Y(n_29055));
NAND3X1 g108408(.A (n_28177), .B (n_25496), .C (n_26018), .Y(n_29054));
NAND3X1 g108409(.A (n_28176), .B (n_26612), .C (n_27236), .Y(n_29053));
NOR2X1 g108413(.A (n_9166), .B (n_28300), .Y (n_29052));
OAI21X1 g108423(.A0 (n_20772), .A1 (n_21365), .B0 (n_27996), .Y(n_29051));
AOI21X1 g108424(.A0 (n_29049), .A1 (n_30557), .B0 (n_21729), .Y(n_35928));
NOR2X1 g108427(.A (n_9109), .B (n_28299), .Y (n_29048));
NOR2X1 g108435(.A (n_9929), .B (n_27982), .Y (n_29047));
NOR2X1 g106857(.A (n_26919), .B (n_28074), .Y (n_29046));
OAI21X1 g108437(.A0 (n_27715), .A1 (n_8321), .B0 (n_20172), .Y(n_29045));
NOR2X1 g106858(.A (n_26917), .B (n_28066), .Y (n_29044));
OAI21X1 g108439(.A0 (n_10525), .A1 (n_20770), .B0 (n_27975), .Y(n_29043));
AOI21X1 g108440(.A0 (n_34714), .A1 (n_29040), .B0 (n_21720), .Y(n_29042));
OAI21X1 g108444(.A0 (n_27726), .A1 (n_8321), .B0 (n_20736), .Y(n_29039));
OAI21X1 g108449(.A0 (n_27732), .A1 (n_26108), .B0 (n_30958), .Y(n_29038));
NAND2X1 g106866(.A (n_28249), .B (n_31891), .Y (n_29037));
NOR2X1 g108464(.A (n_27900), .B (n_26952), .Y (n_29036));
NAND2X1 g108484(.A (n_27963), .B (n_28572), .Y (n_29378));
INVX1 g108489(.A (n_29601), .Y (n_29035));
NAND2X1 g108492(.A (n_27962), .B (n_28569), .Y (n_29893));
NAND2X2 g108497(.A (n_27960), .B (n_29034), .Y (n_32340));
OAI21X1 g108505(.A0 (n_27231), .A1 (n_27696), .B0 (n_27973), .Y(n_29033));
AOI21X1 g108508(.A0 (n_28593), .A1 (n_25988), .B0 (n_27968), .Y(n_29032));
AOI21X1 g108512(.A0 (n_28511), .A1 (n_30180), .B0 (n_19622), .Y(n_35874));
NOR2X1 g108521(.A (n_27922), .B (n_26945), .Y (n_29029));
AOI21X1 g108527(.A0 (n_27720), .A1 (n_29027), .B0 (n_15086), .Y(n_29028));
AOI21X1 g108528(.A0 (n_28464), .A1 (n_34952), .B0 (n_15082), .Y(n_29026));
NOR2X1 g108529(.A (n_7068), .B (n_28047), .Y (n_29025));
INVX1 g108540(.A (n_29613), .Y (n_29024));
NAND2X1 g108544(.A (n_28000), .B (n_28556), .Y (n_29359));
INVX1 g108545(.A (n_29611), .Y (n_29023));
NAND2X1 g108548(.A (n_27988), .B (n_13628), .Y (n_29926));
NAND2X2 g108552(.A (n_27987), .B (n_25151), .Y (n_35248));
NAND2X1 g108556(.A (n_27985), .B (n_28555), .Y (n_29357));
INVX1 g108558(.A (n_33444), .Y (n_29020));
INVX1 g108560(.A (n_29606), .Y (n_29019));
NAND2X1 g108568(.A (n_27984), .B (n_26985), .Y (n_29018));
NAND2X1 g108572(.A (n_27979), .B (n_28551), .Y (n_29355));
INVX2 g108574(.A (n_28550), .Y (n_29923));
NAND2X1 g108584(.A (n_27952), .B (n_13487), .Y (n_29919));
INVX1 g108586(.A (n_33783), .Y (n_29015));
NAND2X1 g108589(.A (n_27951), .B (n_28548), .Y (n_29889));
NAND2X1 g108595(.A (n_27948), .B (n_29014), .Y (n_29906));
INVX1 g108600(.A (n_30201), .Y (n_29345));
NAND2X1 g108602(.A (n_27910), .B (n_13181), .Y (n_29915));
NAND2X1 g108604(.A (n_27909), .B (n_28542), .Y (n_29878));
INVX1 g108605(.A (n_29615), .Y (n_29012));
INVX2 g108607(.A (n_29011), .Y (n_29917));
AOI21X1 g108611(.A0 (n_29009), .A1 (n_29008), .B0 (n_27473), .Y(n_29010));
OAI21X1 g108612(.A0 (n_27719), .A1 (n_28528), .B0 (n_20383), .Y(n_29007));
OAI21X1 g108613(.A0 (n_27704), .A1 (n_33734), .B0 (n_21723), .Y(n_29006));
OAI21X1 g108615(.A0 (n_10021), .A1 (n_20160), .B0 (n_27911), .Y(n_29005));
OAI21X1 g108619(.A0 (n_27704), .A1 (n_29000), .B0 (n_21693), .Y(n_29004));
NAND2X1 g108621(.A (n_27977), .B (n_28021), .Y (n_29003));
NAND2X1 g106933(.A (n_29438), .B (n_18909), .Y (n_29002));
AOI21X1 g108631(.A0 (n_14665), .A1 (n_28401), .B0 (n_29000), .Y(n_29001));
INVX1 g108639(.A (n_28999), .Y (n_29335));
AOI21X1 g108648(.A0 (n_28971), .A1 (n_28275), .B0 (n_28017), .Y(n_28997));
NAND2X1 g108657(.A (n_27942), .B (n_21731), .Y (n_28996));
OAI21X1 g108659(.A0 (n_27226), .A1 (n_27696), .B0 (n_27994), .Y(n_28995));
NAND4X1 g106947(.A (n_14181), .B (n_13747), .C (n_28993), .D(n_26993), .Y (n_28994));
NAND2X1 g108665(.A (n_27501), .B (n_27954), .Y (n_28992));
NAND2X1 g108667(.A (n_27499), .B (n_27924), .Y (n_28991));
AOI21X1 g108668(.A0 (n_28376), .A1 (n_8954), .B0 (n_20127), .Y(n_28990));
NAND2X1 g108669(.A (n_27936), .B (n_20718), .Y (n_28988));
NAND2X1 g108671(.A (n_27904), .B (n_26951), .Y (n_28987));
NAND4X1 g106950(.A (n_14989), .B (n_14527), .C (n_27134), .D(n_26992), .Y (n_28986));
NAND2X1 g108674(.A (n_27908), .B (n_27937), .Y (n_28985));
NAND2X1 g108677(.A (n_27947), .B (n_20713), .Y (n_28984));
OAI21X1 g108680(.A0 (n_28969), .A1 (n_27192), .B0 (n_20429), .Y(n_28983));
OAI21X1 g108681(.A0 (n_28966), .A1 (n_33734), .B0 (n_21706), .Y(n_28982));
NAND4X1 g106954(.A (n_14775), .B (n_14768), .C (n_27118), .D(n_26991), .Y (n_28980));
OAI21X1 g108683(.A0 (n_28182), .A1 (n_8333), .B0 (n_19557), .Y(n_28979));
NAND2X1 g108687(.A (n_6572), .B (n_28046), .Y (n_28978));
NAND2X1 g108691(.A (n_27885), .B (n_20385), .Y (n_28977));
OAI21X1 g108692(.A0 (n_27759), .A1 (n_28528), .B0 (n_21699), .Y(n_28976));
NAND4X1 g106962(.A (n_15165), .B (n_14522), .C (n_28974), .D(n_26990), .Y (n_28975));
AOI21X1 g108698(.A0 (n_34312), .A1 (n_28971), .B0 (n_28027), .Y(n_28972));
OAI21X1 g108708(.A0 (n_28969), .A1 (n_8661), .B0 (n_26959), .Y(n_28970));
OAI21X1 g108709(.A0 (n_28966), .A1 (n_28523), .B0 (n_27460), .Y(n_28967));
NAND3X1 g108728(.A (n_20220), .B (n_27641), .C (n_26659), .Y(n_28965));
NOR2X1 g108731(.A (n_27742), .B (n_28237), .Y (n_28964));
NAND2X1 g106977(.A (n_28211), .B (n_12962), .Y (n_28963));
NOR2X1 g108734(.A (n_27741), .B (n_28225), .Y (n_28962));
OAI21X1 g106982(.A0 (n_27466), .A1 (n_27569), .B0 (n_7827), .Y(n_28961));
NAND3X1 g108753(.A (n_28229), .B (n_27620), .C (n_20865), .Y(n_28959));
NOR2X1 g108760(.A (n_28173), .B (n_28232), .Y (n_28958));
NOR2X1 g108761(.A (n_28172), .B (n_28228), .Y (n_28957));
NOR2X1 g108763(.A (n_28174), .B (n_28226), .Y (n_28956));
NAND4X1 g106996(.A (n_14552), .B (n_14163), .C (n_28954), .D(n_26987), .Y (n_28955));
NAND3X1 g108768(.A (n_10865), .B (n_27644), .C (n_26700), .Y(n_28953));
NOR2X1 g108769(.A (n_28179), .B (n_11130), .Y (n_32316));
NAND2X1 g108779(.A (n_34712), .B (n_28891), .Y (n_28951));
NAND2X1 g108787(.A (n_34712), .B (n_28870), .Y (n_28950));
NAND2X1 g108806(.A (n_28948), .B (n_34718), .Y (n_28949));
NAND2X1 g108811(.A (n_34770), .B (n_28931), .Y (n_28947));
NAND2X1 g108812(.A (n_34770), .B (n_28929), .Y (n_28946));
NAND2X1 g108817(.A (n_34770), .B (n_28924), .Y (n_28944));
NAND2X1 g108818(.A (n_29065), .B (n_28922), .Y (n_28943));
AND2X1 g108824(.A (n_28918), .B (n_28926), .Y (n_28942));
AND2X1 g108825(.A (n_28940), .B (n_28926), .Y (n_28941));
NOR2X1 g108828(.A (n_28206), .B (n_8319), .Y (n_28939));
AND2X1 g108833(.A (n_28934), .B (n_34708), .Y (n_28935));
NAND2X1 g108837(.A (n_28931), .B (n_29925), .Y (n_28932));
NAND2X1 g108838(.A (n_28929), .B (n_29925), .Y (n_28930));
AND2X1 g108839(.A (n_28927), .B (n_28926), .Y (n_28928));
NAND2X1 g108844(.A (n_28924), .B (n_29925), .Y (n_28925));
NAND2X1 g108845(.A (n_28922), .B (n_29925), .Y (n_28923));
NOR2X1 g108846(.A (n_28770), .B (n_29000), .Y (n_28921));
NOR2X1 g108849(.A (n_28192), .B (n_10790), .Y (n_28920));
NAND2X1 g108859(.A (n_28918), .B (n_28013), .Y (n_28919));
NAND2X1 g108860(.A (n_28940), .B (n_28013), .Y (n_28917));
NAND2X1 g108872(.A (n_34718), .B (n_28915), .Y (n_28916));
NAND2X1 g108873(.A (n_28934), .B (n_28013), .Y (n_28914));
NOR2X1 g107040(.A (n_26027), .B (n_28248), .Y (n_28913));
NOR2X1 g107042(.A (n_26026), .B (n_28238), .Y (n_28912));
NAND2X1 g108880(.A (n_28931), .B (n_28013), .Y (n_28911));
NAND2X1 g108881(.A (n_28929), .B (n_29455), .Y (n_28910));
NAND2X1 g108882(.A (n_28927), .B (n_29455), .Y (n_28909));
NAND2X1 g108888(.A (n_28924), .B (n_29455), .Y (n_28908));
NAND2X1 g108889(.A (n_28922), .B (n_29908), .Y (n_28907));
NAND2X1 g108891(.A (n_28905), .B (n_29908), .Y (n_28906));
NAND2X1 g108922(.A (n_29396), .B (n_30559), .Y (n_28901));
NOR2X1 g108926(.A (n_28899), .B (n_8718), .Y (n_28900));
NOR2X1 g108927(.A (n_28209), .B (n_30355), .Y (n_28898));
NAND2X1 g108928(.A (n_29392), .B (n_25756), .Y (n_32291));
OAI21X1 g107070(.A0 (n_8261), .A1 (n_30691), .B0 (n_28290), .Y(n_28896));
AOI21X1 g108971(.A0 (n_23166), .A1 (n_8303), .B0 (n_28233), .Y(n_28895));
NAND2X1 g108972(.A (n_29390), .B (n_28431), .Y (n_28894));
NOR2X1 g108977(.A (n_28217), .B (n_8718), .Y (n_28893));
NAND2X1 g109006(.A (n_28891), .B (n_28890), .Y (n_28892));
NAND2X1 g109007(.A (n_28891), .B (n_26665), .Y (n_28889));
NOR2X1 g107088(.A (n_8903), .B (n_27841), .Y (n_28888));
NAND3X1 g109024(.A (n_28230), .B (n_27081), .C (n_20895), .Y(n_28887));
NAND3X1 g109026(.A (n_26796), .B (n_27612), .C (n_20908), .Y(n_28886));
NAND2X1 g109039(.A (n_8284), .B (n_28883), .Y (n_28885));
NAND2X1 g109041(.A (n_26255), .B (n_28883), .Y (n_28884));
NAND2X1 g109042(.A (n_29427), .B (n_28883), .Y (n_28882));
NAND2X1 g109071(.A (n_30171), .B (n_28879), .Y (n_28881));
NAND2X1 g109072(.A (n_28879), .B (n_8922), .Y (n_28880));
NAND2X1 g109073(.A (n_28879), .B (n_29684), .Y (n_28877));
NAND2X1 g109074(.A (n_8284), .B (n_29760), .Y (n_28876));
NAND2X1 g109101(.A (n_28759), .B (n_28874), .Y (n_28875));
NAND3X1 g107124(.A (n_21633), .B (n_24842), .C (n_27590), .Y(n_30462));
NAND2X1 g109104(.A (n_30171), .B (n_27682), .Y (n_28872));
NAND2X1 g109118(.A (n_28870), .B (n_29191), .Y (n_28871));
NOR2X1 g109136(.A (n_28199), .B (n_29553), .Y (n_28869));
NAND3X1 g109174(.A (n_27585), .B (n_27015), .C (n_27593), .Y(n_28867));
NOR2X1 g107150(.A (n_6779), .B (n_27856), .Y (n_28866));
NAND2X1 g109189(.A (n_27691), .B (n_28364), .Y (n_28863));
NAND2X1 g109190(.A (n_27689), .B (n_28319), .Y (n_28862));
AOI21X1 g109214(.A0 (n_23165), .A1 (n_8303), .B0 (n_28187), .Y(n_28861));
OAI21X1 g109234(.A0 (n_27603), .A1 (n_8321), .B0 (n_20199), .Y(n_28860));
OAI21X1 g109242(.A0 (n_27600), .A1 (n_29150), .B0 (n_20184), .Y(n_28859));
OAI21X1 g109247(.A0 (n_27598), .A1 (n_29150), .B0 (n_19617), .Y(n_28858));
NAND3X1 g109254(.A (n_10202), .B (n_27638), .C (n_26710), .Y(n_28857));
OAI21X1 g109255(.A0 (n_28148), .A1 (n_8285), .B0 (n_20158), .Y(n_28856));
NAND3X1 g109264(.A (n_10190), .B (n_27640), .C (n_26640), .Y(n_28855));
NAND2X1 g109278(.A (n_28247), .B (n_29505), .Y (n_28854));
NAND3X1 g109296(.A (n_10133), .B (n_27639), .C (n_26608), .Y(n_28853));
NOR2X1 g109298(.A (n_10131), .B (n_28178), .Y (n_28852));
NAND3X1 g109328(.A (n_25526), .B (n_27615), .C (n_25491), .Y(n_28849));
AOI21X1 g109331(.A0 (n_26565), .A1 (n_34952), .B0 (n_15279), .Y(n_35095));
AOI21X1 g109335(.A0 (n_26562), .A1 (n_34952), .B0 (n_15106), .Y(n_35633));
INVX1 g109341(.A (n_33509), .Y (n_28846));
NAND2X1 g109347(.A (n_28274), .B (n_27389), .Y (n_29275));
NAND2X1 g109359(.A (n_28266), .B (n_27384), .Y (n_29272));
INVX1 g109366(.A (n_30589), .Y (n_28845));
NAND2X1 g109369(.A (n_28259), .B (n_27380), .Y (n_29270));
NAND2X1 g109382(.A (n_28250), .B (n_27377), .Y (n_29269));
INVX1 g109386(.A (n_33498), .Y (n_28844));
INVX1 g109392(.A (n_28323), .Y (n_29268));
NAND2X1 g107257(.A (n_29254), .B (n_8966), .Y (n_28843));
NAND2X1 g107259(.A (n_29254), .B (n_33738), .Y (n_28841));
INVX1 g109445(.A (n_28840), .Y (n_29263));
OAI21X1 g109453(.A0 (n_27604), .A1 (n_33340), .B0 (n_27311), .Y(n_28839));
OAI21X1 g109454(.A0 (n_27602), .A1 (n_10276), .B0 (n_27327), .Y(n_28838));
OAI21X1 g109456(.A0 (n_27601), .A1 (n_33340), .B0 (n_27303), .Y(n_28837));
OAI21X1 g109458(.A0 (n_27599), .A1 (n_27045), .B0 (n_27296), .Y(n_28836));
OAI21X1 g109462(.A0 (n_27596), .A1 (n_10276), .B0 (n_27317), .Y(n_28835));
OAI21X1 g109465(.A0 (n_28315), .A1 (n_8285), .B0 (n_27332), .Y(n_28834));
AOI21X1 g109466(.A0 (n_30369), .A1 (n_35201), .B0 (n_27807), .Y(n_28833));
NAND3X1 g109505(.A (n_19001), .B (n_26139), .C (n_27023), .Y(n_28832));
NAND2X1 g109545(.A (n_28817), .B (n_28864), .Y (n_28831));
NAND2X1 g107309(.A (n_27570), .B (n_12966), .Y (n_28830));
NAND2X1 g109548(.A (n_26559), .B (n_29061), .Y (n_28829));
NAND2X1 g109549(.A (n_28813), .B (n_28864), .Y (n_28828));
NAND2X1 g109550(.A (n_28826), .B (n_29061), .Y (n_28827));
NAND2X1 g109553(.A (n_34692), .B (n_29061), .Y (n_28825));
NAND2X1 g109557(.A (n_26565), .B (n_30563), .Y (n_28824));
NAND2X1 g109558(.A (n_28809), .B (n_28485), .Y (n_28822));
NAND2X1 g109562(.A (n_26562), .B (n_30563), .Y (n_28820));
NAND2X1 g109564(.A (n_28817), .B (n_28485), .Y (n_28818));
NAND2X1 g109567(.A (n_26559), .B (n_30563), .Y (n_28816));
NAND2X1 g109568(.A (n_28813), .B (n_28485), .Y (n_28814));
NAND2X1 g109576(.A (n_28809), .B (n_28808), .Y (n_35268));
NAND2X1 g109577(.A (n_28140), .B (n_30197), .Y (n_28807));
NAND2X1 g109581(.A (n_28138), .B (n_29604), .Y (n_28806));
NAND2X1 g109582(.A (n_28817), .B (n_30197), .Y (n_35111));
NAND2X1 g109586(.A (n_28813), .B (n_29604), .Y (n_28804));
NAND2X1 g109587(.A (n_28826), .B (n_30197), .Y (n_28803));
NAND2X1 g109590(.A (n_28146), .B (n_33378), .Y (n_28802));
NAND2X1 g109591(.A (n_28850), .B (n_30197), .Y (n_32187));
NAND2X1 g109605(.A (n_28796), .B (n_28798), .Y (n_28799));
NAND2X1 g109606(.A (n_28796), .B (n_28791), .Y (n_32084));
NAND2X1 g109644(.A (n_28793), .B (n_28785), .Y (n_32071));
NAND2X1 g109645(.A (n_28793), .B (n_28798), .Y (n_28794));
NAND2X1 g109646(.A (n_28793), .B (n_28791), .Y (n_32088));
NOR2X1 g109672(.A (n_27594), .B (n_27588), .Y (n_28790));
NAND3X1 g109674(.A (n_26187), .B (n_27035), .C (n_25780), .Y(n_28789));
NAND2X1 g109718(.A (n_27066), .B (n_34753), .Y (n_35073));
NOR2X1 g109795(.A (n_27629), .B (n_13519), .Y (n_28787));
NAND2X1 g109834(.A (n_28796), .B (n_28785), .Y (n_28786));
NAND3X1 g109846(.A (n_27654), .B (n_24439), .C (n_15077), .Y(n_28784));
NAND3X1 g109849(.A (n_27653), .B (n_24455), .C (n_15061), .Y(n_28783));
NOR2X1 g107427(.A (n_8888), .B (n_27656), .Y (n_28782));
NAND3X1 g109890(.A (n_9587), .B (n_26145), .C (n_27033), .Y(n_28781));
NAND3X1 g109892(.A (n_27032), .B (n_20292), .C (n_27029), .Y(n_28780));
OAI21X1 g109913(.A0 (n_27013), .A1 (n_33807), .B0 (n_20471), .Y(n_28779));
NAND2X1 g109928(.A (n_27631), .B (n_26575), .Y (n_28778));
OAI21X1 g109982(.A0 (n_26382), .A1 (n_27010), .B0 (n_26173), .Y(n_28777));
OAI21X1 g109984(.A0 (n_26382), .A1 (n_27011), .B0 (n_27592), .Y(n_28776));
INVX1 g110004(.A (n_28918), .Y (n_28775));
INVX1 g107508(.A (n_29438), .Y (n_28774));
INVX1 g110010(.A (n_28214), .Y (n_29302));
AOI21X1 g107512(.A0 (n_15299), .A1 (n_28154), .B0 (n_29000), .Y(n_28773));
INVX1 g110020(.A (n_28899), .Y (n_28772));
INVX1 g110046(.A (n_29839), .Y (n_28771));
INVX1 g110071(.A (n_28770), .Y (n_29295));
NAND2X1 g110076(.A (n_27626), .B (n_20886), .Y (n_28769));
NAND2X1 g110078(.A (n_27622), .B (n_19842), .Y (n_28768));
INVX1 g110085(.A (n_28870), .Y (n_28767));
INVX1 g110091(.A (n_28905), .Y (n_28766));
AOI21X1 g110101(.A0 (n_34712), .A1 (n_27247), .B0 (n_27650), .Y(n_28765));
NAND2X1 g107542(.A (n_6481), .B (n_27667), .Y (n_28764));
OAI21X1 g107545(.A0 (n_26998), .A1 (n_31275), .B0 (n_6512), .Y(n_28763));
NAND2X1 g110129(.A (n_27610), .B (n_15111), .Y (n_28762));
AOI21X1 g110133(.A0 (n_28165), .A1 (n_29405), .B0 (n_14979), .Y(n_28761));
OAI21X1 g107550(.A0 (n_26995), .A1 (n_31278), .B0 (n_6574), .Y(n_28760));
INVX1 g110156(.A (n_28759), .Y (n_29230));
NAND2X1 g107578(.A (n_27558), .B (n_31097), .Y (n_28756));
NAND2X1 g107580(.A (n_27556), .B (n_31594), .Y (n_28755));
AOI21X1 g110212(.A0 (n_34712), .A1 (n_27253), .B0 (n_27652), .Y(n_28754));
NAND2X1 g107582(.A (n_27528), .B (n_917), .Y (n_28753));
NAND2X1 g110217(.A (n_26731), .B (n_27657), .Y (n_28751));
NAND2X1 g110218(.A (n_27648), .B (n_26752), .Y (n_28750));
OAI21X1 g110222(.A0 (n_27193), .A1 (n_27662), .B0 (n_27635), .Y(n_28749));
OAI21X1 g110227(.A0 (n_27017), .A1 (n_28747), .B0 (n_27098), .Y(n_28748));
NAND2X1 g110228(.A (n_27646), .B (n_26751), .Y (n_28746));
AOI21X1 g107618(.A0 (n_26968), .A1 (n_26354), .B0 (n_31041), .Y(n_28745));
AOI21X1 g107633(.A0 (n_26950), .A1 (n_26357), .B0 (n_8340), .Y(n_28744));
AOI21X1 g107640(.A0 (n_26928), .A1 (n_25495), .B0 (n_8340), .Y(n_28743));
NAND2X1 g108252(.A (n_28741), .B (n_25756), .Y (n_35081));
NAND2X1 g107682(.A (n_28738), .B (n_30200), .Y (n_28740));
NAND2X1 g107706(.A (n_28738), .B (n_33738), .Y (n_28739));
NAND2X1 g107712(.A (n_33626), .B (n_23356), .Y (n_28737));
NAND2X1 g107734(.A (n_33626), .B (n_28734), .Y (n_28736));
NAND2X1 g107762(.A (n_27526), .B (n_12960), .Y (n_28733));
NAND3X1 g107780(.A (n_26936), .B (n_26918), .C (n_15187), .Y(n_28732));
NAND4X1 g107785(.A (n_27358), .B (n_26794), .C (n_26816), .D(n_26856), .Y (n_28731));
NAND2X1 g107789(.A (n_29568), .B (n_28715), .Y (n_28730));
NAND2X1 g107800(.A (n_8284), .B (n_28726), .Y (n_28729));
NAND2X1 g107801(.A (n_27632), .B (n_28726), .Y (n_28728));
NAND2X1 g107802(.A (n_29427), .B (n_28726), .Y (n_28725));
NAND2X1 g107803(.A (n_28709), .B (n_28124), .Y (n_29697));
NAND2X1 g107804(.A (n_15302), .B (n_28711), .Y (n_28724));
NAND2X1 g107807(.A (n_34215), .B (n_18262), .Y (n_28723));
NAND2X1 g107826(.A (n_28721), .B (n_33738), .Y (n_28722));
NOR2X1 g107831(.A (n_27536), .B (n_26434), .Y (n_28718));
NAND2X1 g107861(.A (n_28874), .B (n_28715), .Y (n_32314));
NAND2X1 g107862(.A (n_28738), .B (n_26238), .Y (n_32313));
NAND2X1 g107863(.A (n_27538), .B (n_29505), .Y (n_28713));
NAND2X1 g107864(.A (n_29551), .B (n_28715), .Y (n_28712));
NAND2X1 g107865(.A (n_28125), .B (n_28711), .Y (n_29686));
NAND2X1 g107866(.A (n_28709), .B (n_15295), .Y (n_28710));
INVX1 g110877(.A (n_28144), .Y (n_28708));
NAND2X1 g107881(.A (n_28721), .B (n_29405), .Y (n_28707));
NAND2X1 g107888(.A (n_28704), .B (n_29411), .Y (n_28706));
NAND2X1 g107893(.A (n_28704), .B (n_8954), .Y (n_28705));
NAND2X1 g107898(.A (n_28704), .B (n_29405), .Y (n_28702));
NAND2X1 g107899(.A (n_28704), .B (n_30636), .Y (n_28701));
NAND2X1 g107911(.A (n_34215), .B (n_26584), .Y (n_29693));
NAND2X1 g107917(.A (n_28696), .B (n_33738), .Y (n_28695));
NAND2X1 g110989(.A (n_27578), .B (n_25755), .Y (n_28694));
OAI21X1 g111061(.A0 (n_26067), .A1 (n_30138), .B0 (n_27573), .Y(n_28693));
NAND2X1 g111074(.A (n_27571), .B (n_25728), .Y (n_28692));
AOI21X1 g111078(.A0 (n_27053), .A1 (n_28791), .B0 (n_27580), .Y(n_28691));
AOI21X1 g111081(.A0 (n_28126), .A1 (n_30369), .B0 (n_26540), .Y(n_28690));
OAI21X1 g111082(.A0 (n_27527), .A1 (n_8319), .B0 (n_25776), .Y(n_28689));
AOI21X1 g111086(.A0 (n_26181), .A1 (n_28791), .B0 (n_27576), .Y(n_28688));
OAI21X1 g106663(.A0 (n_28666), .A1 (n_27042), .B0 (n_8284), .Y(n_28687));
NAND2X1 g107978(.A (n_27547), .B (n_29505), .Y (n_28685));
NAND2X1 g111133(.A (n_28681), .B (n_26160), .Y (n_28684));
OAI21X1 g107990(.A0 (n_26922), .A1 (n_26830), .B0 (n_33123), .Y(n_28683));
NAND2X1 g111179(.A (n_28681), .B (n_30197), .Y (n_28682));
NOR2X1 g108013(.A (n_26982), .B (n_27554), .Y (n_28680));
NAND4X1 g108014(.A (n_27551), .B (n_25213), .C (n_25462), .D(n_25494), .Y (n_28679));
CLKBUFX1 gbuf_d_357(.A(n_27516), .Y(d_out_357));
CLKBUFX1 gbuf_q_357(.A(q_in_357), .Y(n_10452));
AOI21X1 g108046(.A0 (n_25247), .A1 (n_26213), .B0 (n_27531), .Y(n_28678));
AOI21X1 g108066(.A0 (n_14719), .A1 (n_28084), .B0 (n_29000), .Y(n_28677));
INVX1 g108069(.A (n_28676), .Y (n_29719));
NAND2X1 g108076(.A (n_27541), .B (n_28153), .Y (n_29125));
NAND2X1 g108095(.A (n_6546), .B (n_27534), .Y (n_28675));
NAND2X1 g108097(.A (n_6597), .B (n_27533), .Y (n_28674));
NAND2X1 g108098(.A (n_6576), .B (n_27559), .Y (n_28673));
NOR2X1 g108119(.A (n_27347), .B (n_27408), .Y (n_28672));
NAND3X1 g108132(.A (n_27376), .B (n_26843), .C (n_26778), .Y(n_28671));
NOR2X1 g108142(.A (n_27363), .B (n_27402), .Y (n_28670));
NOR2X1 g108150(.A (n_27833), .B (n_27406), .Y (n_28669));
NOR2X1 g108152(.A (n_27831), .B (n_27401), .Y (n_28668));
OAI21X1 g106739(.A0 (n_28666), .A1 (n_28528), .B0 (n_27563), .Y(n_28667));
OAI21X1 g106746(.A0 (n_15130), .A1 (n_29968), .B0 (n_27518), .Y(n_28665));
OAI21X1 g106747(.A0 (n_15141), .A1 (n_28659), .B0 (n_27514), .Y(n_28664));
NAND2X1 g108179(.A (n_28655), .B (n_34952), .Y (n_28663));
NAND2X1 g108182(.A (n_28647), .B (n_34952), .Y (n_28661));
OAI21X1 g106749(.A0 (n_15281), .A1 (n_28659), .B0 (n_27508), .Y(n_35326));
NAND2X1 g108187(.A (n_28653), .B (n_29619), .Y (n_28658));
NAND2X1 g108190(.A (n_28651), .B (n_29619), .Y (n_28657));
NAND2X1 g108193(.A (n_28655), .B (n_28485), .Y (n_28656));
NAND2X1 g108201(.A (n_28653), .B (n_28808), .Y (n_28654));
NAND2X1 g108204(.A (n_28651), .B (n_28808), .Y (n_28652));
NAND2X1 g108207(.A (n_28655), .B (n_26142), .Y (n_28650));
NAND2X1 g108210(.A (n_28647), .B (n_26142), .Y (n_28648));
NAND4X1 g108218(.A (n_15098), .B (n_25470), .C (n_26614), .D(n_25479), .Y (n_28646));
NAND4X1 g108220(.A (n_15067), .B (n_26589), .C (n_26256), .D(n_26590), .Y (n_28645));
NOR2X1 g108225(.A (n_27360), .B (n_14921), .Y (n_28644));
NAND2X1 g108234(.A (n_28642), .B (n_25756), .Y (n_32266));
NAND2X1 g108235(.A (n_28642), .B (n_28636), .Y (n_28641));
NAND2X1 g108236(.A (n_28642), .B (n_26528), .Y (n_28640));
NAND2X1 g108238(.A (n_28634), .B (n_27999), .Y (n_28639));
NAND2X1 g108240(.A (n_24652), .B (n_33368), .Y (n_28638));
CLKBUFX1 gbuf_d_358(.A(n_27699), .Y(d_out_358));
CLKBUFX1 gbuf_q_358(.A(q_in_358), .Y(P2_reg1[3]));
NAND2X1 g108253(.A (n_28741), .B (n_28636), .Y (n_28637));
NAND2X1 g108256(.A (n_28634), .B (n_23270), .Y (n_28635));
CLKBUFX1 gbuf_d_359(.A(n_27700), .Y(d_out_359));
CLKBUFX1 gbuf_q_359(.A(q_in_359), .Y(n_9599));
CLKBUFX1 gbuf_d_360(.A(n_27515), .Y(d_out_360));
CLKBUFX1 gbuf_q_360(.A(q_in_360), .Y(P2_reg1[1]));
CLKBUFX1 gbuf_d_361(.A(n_27674), .Y(d_out_361));
CLKBUFX1 gbuf_q_361(.A(q_in_361), .Y(n_13215));
CLKBUFX1 gbuf_d_362(.A(n_27672), .Y(d_out_362));
CLKBUFX1 gbuf_q_362(.A(q_in_362), .Y(n_2718));
NAND2X1 g108258(.A (n_33368), .B (n_18384), .Y (n_28633));
AOI21X1 g108261(.A0 (n_27355), .A1 (n_27140), .B0 (n_30537), .Y(n_28631));
NAND2X1 g108269(.A (n_27849), .B (n_10808), .Y (n_28630));
NOR2X1 g108270(.A (n_8382), .B (n_29122), .Y (n_28628));
NAND4X1 g108272(.A (n_27712), .B (n_26800), .C (n_24089), .D(n_26747), .Y (n_28627));
NAND2X1 g108273(.A (n_28634), .B (n_32664), .Y (n_28626));
NAND2X1 g108275(.A (n_33368), .B (n_32798), .Y (n_28625));
NAND2X1 g108276(.A (n_28615), .B (n_14207), .Y (n_28624));
OAI21X1 g108277(.A0 (n_27350), .A1 (n_25825), .B0 (n_34731), .Y(n_28623));
OAI21X1 g106788(.A0 (n_28666), .A1 (n_25540), .B0 (n_26487), .Y(n_28622));
NAND2X1 g108295(.A (n_27861), .B (n_10808), .Y (n_28620));
NOR2X1 g108296(.A (n_8382), .B (n_35629), .Y (n_28619));
NAND2X1 g108298(.A (n_28634), .B (n_34688), .Y (n_28618));
NAND2X1 g108312(.A (n_28054), .B (n_28603), .Y (n_29585));
NAND2X1 g108313(.A (n_14946), .B (n_28605), .Y (n_28616));
NAND2X1 g108314(.A (n_28538), .B (n_28615), .Y (n_29578));
NAND2X1 g108315(.A (n_14838), .B (n_28612), .Y (n_28614));
NAND2X1 g108320(.A (n_28606), .B (n_17968), .Y (n_29572));
NAND2X1 g108322(.A (n_28543), .B (n_28612), .Y (n_29547));
NAND2X1 g108326(.A (n_20755), .B (n_28608), .Y (n_29565));
NOR2X1 g108329(.A (n_27368), .B (n_27832), .Y (n_28611));
NAND2X2 g108336(.A (n_28532), .B (n_28610), .Y (n_29526));
NAND2X1 g108337(.A (n_28608), .B (n_14608), .Y (n_28609));
NAND2X2 g108340(.A (n_28606), .B (n_35842), .Y (n_28607));
NAND2X1 g108353(.A (n_28605), .B (n_28058), .Y (n_29567));
NAND2X1 g108354(.A (n_28603), .B (n_14478), .Y (n_28604));
OAI21X1 g108357(.A0 (n_27259), .A1 (n_25443), .B0 (n_30099), .Y(n_28602));
NOR2X1 g108366(.A (n_27407), .B (n_27197), .Y (n_28601));
NAND3X1 g108372(.A (n_27675), .B (n_26247), .C (n_26782), .Y(n_28600));
NOR2X1 g108373(.A (n_27318), .B (n_27391), .Y (n_28599));
AOI21X1 g108377(.A0 (n_28597), .A1 (n_28025), .B0 (n_26442), .Y(n_35702));
NAND3X1 g108379(.A (n_27504), .B (n_14829), .C (n_25287), .Y(n_28596));
NAND3X1 g108381(.A (n_27503), .B (n_25276), .C (n_14377), .Y(n_28595));
AOI21X1 g108386(.A0 (n_34770), .A1 (n_28593), .B0 (n_26910), .Y(n_28594));
NAND4X1 g108389(.A (n_15101), .B (n_25487), .C (n_26622), .D(n_25485), .Y (n_28592));
NAND4X1 g108391(.A (n_15074), .B (n_26595), .C (n_35607), .D(n_35608), .Y (n_28591));
NAND2X1 g108404(.A (n_28606), .B (n_35508), .Y (n_29544));
NAND2X1 g108407(.A (n_28606), .B (n_25596), .Y (n_28590));
OAI21X1 g108416(.A0 (n_27309), .A1 (n_28588), .B0 (n_8622), .Y(n_28589));
AOI22X1 g108417(.A0 (n_28971), .A1 (n_26288), .B0 (n_20304), .B1(n_19502), .Y (n_28587));
OAI21X1 g108422(.A0 (n_8783), .A1 (n_30731), .B0 (n_27486), .Y(n_28584));
AOI21X1 g108436(.A0 (n_28034), .A1 (n_30369), .B0 (n_20740), .Y(n_28583));
OAI21X1 g108446(.A0 (n_27967), .A1 (n_33807), .B0 (n_20156), .Y(n_28582));
OAI21X1 g108448(.A0 (n_27244), .A1 (n_25826), .B0 (n_30958), .Y(n_28581));
NOR2X1 g108454(.A (n_9553), .B (n_27835), .Y (n_28580));
NOR2X1 g108456(.A (n_27257), .B (n_27364), .Y (n_28579));
NOR2X1 g108457(.A (n_9043), .B (n_27837), .Y (n_28578));
OAI21X1 g108462(.A0 (n_27281), .A1 (n_28588), .B0 (n_8605), .Y(n_28577));
NOR2X1 g108465(.A (n_9184), .B (n_27838), .Y (n_28576));
NOR2X1 g108467(.A (n_9083), .B (n_27375), .Y (n_28575));
NOR2X1 g108470(.A (n_27255), .B (n_27367), .Y (n_28574));
AOI21X1 g108472(.A0 (n_27100), .A1 (n_27933), .B0 (n_27374), .Y(n_28573));
NAND2X1 g108490(.A (n_27468), .B (n_28569), .Y (n_29601));
INVX1 g108493(.A (n_28568), .Y (n_29975));
OAI21X1 g108499(.A0 (n_27299), .A1 (n_28588), .B0 (n_8613), .Y(n_28567));
OAI21X1 g108500(.A0 (n_27286), .A1 (n_31360), .B0 (n_8394), .Y(n_28566));
OAI21X1 g108502(.A0 (n_26382), .A1 (n_27206), .B0 (n_27362), .Y(n_28565));
AOI21X1 g108503(.A0 (n_24925), .A1 (n_27523), .B0 (n_27361), .Y(n_28563));
NAND2X1 g106897(.A (n_33319), .B (n_991), .Y (n_28562));
NOR2X1 g108522(.A (n_27427), .B (n_26449), .Y (n_28560));
OAI21X1 g108523(.A0 (n_27263), .A1 (n_8927), .B0 (n_27425), .Y(n_28559));
INVX1 g108536(.A (n_29192), .Y (n_28557));
NAND2X1 g108541(.A (n_27488), .B (n_28556), .Y (n_29613));
NAND2X1 g108546(.A (n_27487), .B (n_13662), .Y (n_29611));
NAND2X2 g108557(.A (n_27484), .B (n_25151), .Y (n_29623));
NAND2X1 g108561(.A (n_27480), .B (n_28554), .Y (n_29606));
INVX1 g108562(.A (n_29197), .Y (n_28553));
INVX1 g108564(.A (n_29188), .Y (n_28552));
NAND2X1 g108569(.A (n_27478), .B (n_28551), .Y (n_29620));
NAND2X1 g108575(.A (n_27477), .B (n_28549), .Y (n_28550));
INVX1 g108590(.A (n_29194), .Y (n_28547));
INVX1 g108592(.A (n_29178), .Y (n_28546));
NAND2X1 g108596(.A (n_27446), .B (n_21336), .Y (n_28545));
OAI21X1 g108601(.A0 (n_32845), .A1 (n_35538), .B0 (n_28543), .Y(n_30201));
NAND2X1 g108606(.A (n_27423), .B (n_28542), .Y (n_29615));
INVX2 g108608(.A (n_28060), .Y (n_29011));
AOI21X1 g108618(.A0 (n_27920), .A1 (n_8966), .B0 (n_20935), .Y(n_28541));
OAI21X1 g108627(.A0 (n_32843), .A1 (n_13736), .B0 (n_28538), .Y(n_29535));
OAI21X1 g108629(.A0 (n_27683), .A1 (n_8927), .B0 (n_21700), .Y(n_28537));
INVX1 g108632(.A (n_28536), .Y (n_29947));
INVX1 g108634(.A (n_28535), .Y (n_29959));
NAND2X1 g108640(.A (n_27433), .B (n_28083), .Y (n_28999));
NAND2X1 g108646(.A (n_27431), .B (n_28532), .Y (n_32935));
AOI21X1 g108656(.A0 (n_27905), .A1 (n_8954), .B0 (n_20875), .Y(n_28531));
AOI21X1 g108672(.A0 (n_27941), .A1 (n_29955), .B0 (n_27440), .Y(n_28530));
OAI21X1 g108679(.A0 (n_28524), .A1 (n_28528), .B0 (n_21347), .Y(n_28529));
NAND2X1 g108690(.A (n_27415), .B (n_21330), .Y (n_28527));
OAI21X1 g106966(.A0 (n_26944), .A1 (n_27139), .B0 (n_31628), .Y(n_28526));
OAI21X1 g108707(.A0 (n_28524), .A1 (n_28523), .B0 (n_27463), .Y(n_28525));
OAI21X1 g106969(.A0 (n_27111), .A1 (n_22100), .B0 (n_31064), .Y(n_28522));
NAND4X1 g106970(.A (n_27357), .B (n_26939), .C (n_25113), .D(n_26348), .Y (n_28521));
OAI21X1 g108714(.A0 (n_33917), .A1 (n_27451), .B0 (n_27453), .Y(n_29556));
NAND2X2 g108715(.A (n_32058), .B (n_32059), .Y (n_29595));
NAND2X2 g108718(.A (n_32918), .B (n_32919), .Y (n_29562));
NOR2X1 g108737(.A (n_27706), .B (n_27722), .Y (n_28519));
NOR2X1 g108739(.A (n_27216), .B (n_27721), .Y (n_28518));
NAND2X1 g106984(.A (n_33319), .B (n_26870), .Y (n_28517));
OR2X1 g106985(.A (n_33319), .B (n_10067), .Y (n_28516));
NAND3X1 g108750(.A (n_18406), .B (n_26330), .C (n_27132), .Y(n_28515));
NOR2X1 g108757(.A (n_27664), .B (n_27246), .Y (n_28514));
NAND2X1 g108770(.A (n_33546), .B (n_28444), .Y (n_28513));
NAND2X1 g108772(.A (n_33546), .B (n_28511), .Y (n_35875));
NAND2X1 g108777(.A (n_33546), .B (n_28432), .Y (n_28510));
NAND2X1 g108778(.A (n_34712), .B (n_28425), .Y (n_28509));
NAND2X1 g108780(.A (n_33546), .B (n_28423), .Y (n_28508));
NAND2X1 g108781(.A (n_33546), .B (n_28416), .Y (n_28507));
NAND2X1 g108786(.A (n_34712), .B (n_28398), .Y (n_28506));
NAND2X1 g108788(.A (n_33546), .B (n_28390), .Y (n_28505));
NAND2X1 g108789(.A (n_33546), .B (n_28380), .Y (n_28504));
NAND2X1 g108803(.A (n_29068), .B (n_28471), .Y (n_28503));
NAND3X1 g107012(.A (n_26431), .B (n_27356), .C (n_26941), .Y(n_28502));
NAND2X1 g108804(.A (n_28486), .B (n_28864), .Y (n_28501));
NAND2X1 g108808(.A (n_34770), .B (n_28459), .Y (n_28500));
NAND2X1 g108809(.A (n_28483), .B (n_28864), .Y (n_28498));
NAND2X1 g108813(.A (n_9503), .B (n_28479), .Y (n_28497));
NAND2X1 g108814(.A (n_34770), .B (n_28476), .Y (n_28496));
NAND2X1 g108820(.A (n_9503), .B (n_28453), .Y (n_28495));
NAND2X1 g108822(.A (n_28493), .B (n_28492), .Y (n_28494));
NAND2X1 g108827(.A (n_28490), .B (n_28492), .Y (n_28491));
NAND2X1 g108830(.A (n_28488), .B (n_34694), .Y (n_28489));
NAND2X1 g108831(.A (n_28486), .B (n_28485), .Y (n_28487));
NAND2X1 g108834(.A (n_28483), .B (n_28485), .Y (n_28484));
NAND2X1 g108835(.A (n_28481), .B (n_28926), .Y (n_28482));
NAND2X1 g108840(.A (n_28479), .B (n_34709), .Y (n_28480));
NAND2X1 g108841(.A (n_28476), .B (n_34709), .Y (n_28477));
NAND2X1 g108254(.A (n_28741), .B (n_26528), .Y (n_28475));
AND2X1 g108848(.A (n_28451), .B (n_8966), .Y (n_28474));
NAND2X1 g108855(.A (n_28493), .B (n_28468), .Y (n_28473));
NAND2X1 g108863(.A (n_28471), .B (n_28013), .Y (n_28472));
NAND2X1 g108864(.A (n_28490), .B (n_28468), .Y (n_28469));
NAND2X1 g108865(.A (n_29067), .B (n_25980), .Y (n_28467));
NAND2X1 g108866(.A (n_28464), .B (n_29090), .Y (n_28465));
NAND2X1 g108868(.A (n_28488), .B (n_30197), .Y (n_28463));
NAND2X1 g108869(.A (n_28486), .B (n_28808), .Y (n_28462));
NAND2X1 g108874(.A (n_29009), .B (n_26535), .Y (n_28461));
NAND2X1 g108875(.A (n_28459), .B (n_28013), .Y (n_28460));
NAND2X1 g108876(.A (n_28483), .B (n_28808), .Y (n_28458));
NAND2X1 g108877(.A (n_28481), .B (n_33785), .Y (n_28457));
NAND2X1 g108883(.A (n_28479), .B (n_33785), .Y (n_28456));
NAND2X1 g108884(.A (n_28476), .B (n_29455), .Y (n_28455));
NAND2X1 g108892(.A (n_28453), .B (n_33785), .Y (n_28454));
NAND2X1 g108893(.A (n_28451), .B (n_8954), .Y (n_28452));
NAND2X1 g108894(.A (n_28449), .B (n_33784), .Y (n_28450));
INVX1 g108898(.A (n_28007), .Y (n_28903));
OAI21X1 g107052(.A0 (n_27135), .A1 (n_21315), .B0 (n_34731), .Y(n_28448));
NAND2X1 g108921(.A (n_29049), .B (n_30559), .Y (n_28446));
NAND2X1 g108923(.A (n_28444), .B (n_28890), .Y (n_28445));
NAND2X1 g108930(.A (n_28511), .B (n_30559), .Y (n_28443));
NAND2X1 g108932(.A (n_28427), .B (n_28441), .Y (n_28442));
OAI21X1 g107064(.A0 (n_27119), .A1 (n_21314), .B0 (n_34731), .Y(n_28440));
NAND4X1 g108950(.A (n_35135), .B (n_35136), .C (n_23168), .D(n_25656), .Y (n_28439));
NAND4X1 g108951(.A (n_35122), .B (n_35123), .C (n_24469), .D(n_25655), .Y (n_28438));
NAND2X1 g108957(.A (n_28409), .B (n_14670), .Y (n_28437));
NOR2X1 g108959(.A (n_26666), .B (n_27734), .Y (n_28436));
NAND2X1 g108969(.A (n_34714), .B (n_28431), .Y (n_28435));
NAND2X1 g108976(.A (n_28432), .B (n_28431), .Y (n_28433));
NAND2X1 g108979(.A (n_28219), .B (n_24786), .Y (n_28430));
NAND2X1 g108982(.A (n_27229), .B (n_30668), .Y (n_28429));
NAND2X1 g108983(.A (n_28427), .B (n_26965), .Y (n_28428));
NAND2X1 g109003(.A (n_28425), .B (n_28890), .Y (n_28426));
NAND2X1 g109009(.A (n_28423), .B (n_29191), .Y (n_28424));
NAND2X1 g109010(.A (n_28420), .B (n_28890), .Y (n_28422));
NAND2X1 g109011(.A (n_28420), .B (n_30557), .Y (n_28421));
NAND2X1 g109012(.A (n_28420), .B (n_27993), .Y (n_28419));
NAND2X1 g109013(.A (n_28420), .B (n_33513), .Y (n_28418));
NAND2X1 g109014(.A (n_28416), .B (n_30559), .Y (n_28417));
NAND2X1 g109017(.A (n_28427), .B (n_23578), .Y (n_28415));
NAND2X1 g109037(.A (n_28310), .B (n_28394), .Y (n_29429));
NAND2X1 g109038(.A (n_14889), .B (n_28396), .Y (n_28414));
NAND2X1 g109047(.A (n_8284), .B (n_28411), .Y (n_28413));
NAND2X1 g109048(.A (n_27632), .B (n_28411), .Y (n_28412));
NAND2X1 g109049(.A (n_29427), .B (n_28411), .Y (n_28410));
NAND2X1 g109070(.A (n_18939), .B (n_28409), .Y (n_29425));
NAND2X1 g109079(.A (n_30171), .B (n_28406), .Y (n_28408));
NAND2X1 g109080(.A (n_28406), .B (n_8922), .Y (n_28407));
NAND2X1 g109081(.A (n_28372), .B (n_33738), .Y (n_28405));
NOR2X1 g109091(.A (n_27671), .B (n_10571), .Y (n_28404));
NAND2X1 g109099(.A (n_24925), .B (n_27203), .Y (n_28402));
NAND2X1 g109100(.A (n_28401), .B (n_28302), .Y (n_29401));
NAND2X1 g109105(.A (n_28181), .B (n_30454), .Y (n_28400));
NAND2X1 g109117(.A (n_28398), .B (n_26660), .Y (n_28399));
NAND3X1 g109120(.A (n_18007), .B (n_19835), .C (n_27083), .Y(n_28397));
NAND2X1 g109133(.A (n_28396), .B (n_28322), .Y (n_29440));
NAND2X1 g109134(.A (n_28394), .B (n_14247), .Y (n_28395));
NAND2X1 g109141(.A (n_8922), .B (n_28392), .Y (n_28393));
NAND2X1 g109142(.A (n_28390), .B (n_29191), .Y (n_28391));
NAND2X1 g109143(.A (n_28451), .B (n_28158), .Y (n_28389));
NAND2X1 g109144(.A (n_30291), .B (n_28392), .Y (n_28387));
NAND2X1 g109145(.A (n_28451), .B (n_29253), .Y (n_28386));
NAND2X1 g109146(.A (n_28384), .B (n_26660), .Y (n_28385));
AND2X1 g109147(.A (n_28384), .B (n_29040), .Y (n_28383));
NAND2X1 g109148(.A (n_28384), .B (n_30180), .Y (n_28382));
NAND2X1 g109149(.A (n_28380), .B (n_28890), .Y (n_28381));
NAND2X1 g109152(.A (n_28427), .B (n_25734), .Y (n_28379));
NOR2X1 g109153(.A (n_27049), .B (n_27745), .Y (n_28378));
AND2X1 g109164(.A (n_28376), .B (n_28158), .Y (n_28377));
NAND2X1 g109165(.A (n_28376), .B (n_28374), .Y (n_28375));
AND2X1 g109167(.A (n_28372), .B (n_28158), .Y (n_28373));
NAND2X1 g109168(.A (n_28372), .B (n_26238), .Y (n_28371));
NOR2X1 g109169(.A (n_27735), .B (n_27589), .Y (n_28369));
NOR2X1 g109176(.A (n_27728), .B (n_27586), .Y (n_28368));
NOR2X1 g109183(.A (n_27583), .B (n_24477), .Y (n_28367));
NOR2X1 g109185(.A (n_27581), .B (n_24476), .Y (n_28366));
NAND2X1 g109188(.A (n_27208), .B (n_28364), .Y (n_28365));
NAND2X1 g109191(.A (n_28360), .B (n_29411), .Y (n_28363));
NAND2X1 g109193(.A (n_28358), .B (n_29411), .Y (n_28362));
NAND2X1 g109194(.A (n_28360), .B (n_8954), .Y (n_28361));
NAND2X1 g109196(.A (n_28358), .B (n_8954), .Y (n_28359));
NOR2X1 g109198(.A (n_28969), .B (n_25881), .Y (n_28357));
NOR2X1 g109199(.A (n_28966), .B (n_25881), .Y (n_28356));
NAND2X1 g109200(.A (n_28360), .B (n_29405), .Y (n_28355));
NAND2X1 g109201(.A (n_28360), .B (n_30636), .Y (n_28354));
NAND2X1 g109204(.A (n_28358), .B (n_29405), .Y (n_28353));
NAND2X1 g109205(.A (n_28358), .B (n_30636), .Y (n_28352));
NAND2X1 g109209(.A (n_28344), .B (n_33991), .Y (n_32273));
NAND2X1 g109211(.A (n_28342), .B (n_33991), .Y (n_32296));
NAND3X1 g109213(.A (n_24452), .B (n_27142), .C (n_26696), .Y(n_28349));
MX2X1 g107161(.A (n_29695), .B (n_28347), .S0 (n_27041), .Y(n_28348));
NAND3X1 g109216(.A (n_32060), .B (n_32061), .C (n_26597), .Y(n_28346));
NAND2X1 g109228(.A (n_28344), .B (n_29155), .Y (n_28345));
NAND2X1 g109230(.A (n_28342), .B (n_28158), .Y (n_28343));
OAI21X1 g109243(.A0 (n_27062), .A1 (n_8285), .B0 (n_20183), .Y(n_28341));
OAI21X1 g109256(.A0 (n_28252), .A1 (n_29150), .B0 (n_20157), .Y(n_28339));
NAND4X1 g109263(.A (n_27608), .B (n_21357), .C (n_23161), .D(n_25654), .Y (n_28338));
NAND4X1 g109265(.A (n_27607), .B (n_19909), .C (n_24459), .D(n_25653), .Y (n_28337));
NAND3X1 g109266(.A (n_10183), .B (n_27117), .C (n_26708), .Y(n_28336));
NOR2X1 g109273(.A (n_9131), .B (n_27673), .Y (n_28335));
NAND2X1 g109280(.A (n_27765), .B (n_29505), .Y (n_28334));
OAI21X1 g109281(.A0 (n_9842), .A1 (n_28332), .B0 (n_27819), .Y(n_28333));
NOR2X1 g109292(.A (n_10214), .B (n_27680), .Y (n_28331));
NAND3X1 g109295(.A (n_10242), .B (n_26705), .C (n_27106), .Y(n_28330));
INVX1 g109311(.A (n_29093), .Y (n_28329));
NAND2X1 g109329(.A (n_27751), .B (n_20855), .Y (n_28328));
NAND2X1 g109354(.A (n_27791), .B (n_28213), .Y (n_29850));
NAND2X1 g107227(.A (n_27591), .B (n_31097), .Y (n_28326));
NAND2X2 g109367(.A (n_27786), .B (n_28325), .Y (n_30589));
NAND2X1 g109378(.A (n_27772), .B (n_28204), .Y (n_29841));
NAND2X1 g109385(.A (n_27768), .B (n_19492), .Y (n_29819));
NAND2X1 g109390(.A (n_27748), .B (n_28195), .Y (n_29422));
OAI21X1 g109393(.A0 (n_27038), .A1 (n_35520), .B0 (n_28322), .Y(n_28323));
OAI21X1 g109397(.A0 (n_34691), .A1 (n_9455), .B0 (n_27289), .Y(n_28321));
NAND2X1 g109402(.A (n_27755), .B (n_28319), .Y (n_28320));
OAI21X1 g109404(.A0 (n_27077), .A1 (n_13912), .B0 (n_27842), .Y(n_28318));
AOI21X1 g109409(.A0 (n_35197), .A1 (n_30063), .B0 (n_27805), .Y(n_28317));
OAI21X1 g109412(.A0 (n_28315), .A1 (n_8382), .B0 (n_20283), .Y(n_28316));
AOI22X1 g109413(.A0 (n_35201), .A1 (n_25756), .B0 (n_20304), .B1(n_20093), .Y (n_28314));
AOI22X1 g109415(.A0 (n_35197), .A1 (n_26213), .B0 (n_9629), .B1(n_20091), .Y (n_28312));
OAI21X1 g109417(.A0 (n_27038), .A1 (n_13214), .B0 (n_28310), .Y(n_29408));
NOR2X1 g109421(.A (n_25880), .B (n_27663), .Y (n_28309));
NOR2X1 g109423(.A (n_27080), .B (n_27661), .Y (n_28308));
NAND3X1 g109431(.A (n_26758), .B (n_20794), .C (n_27164), .Y(n_28307));
INVX1 g109438(.A (n_28306), .Y (n_29817));
NAND2X1 g109440(.A (n_27763), .B (n_26548), .Y (n_28305));
NAND2X1 g109442(.A (n_27761), .B (n_26548), .Y (n_28304));
NAND2X1 g109446(.A (n_27758), .B (n_28302), .Y (n_28840));
NAND3X1 g109449(.A (n_32117), .B (n_20782), .C (n_32118), .Y(n_28301));
OAI21X1 g109452(.A0 (n_27065), .A1 (n_30138), .B0 (n_27328), .Y(n_28300));
OAI21X1 g109455(.A0 (n_27063), .A1 (n_10276), .B0 (n_27325), .Y(n_28299));
OAI21X1 g109457(.A0 (n_35199), .A1 (n_30138), .B0 (n_27323), .Y(n_28298));
AND2X1 g109469(.A (n_26822), .B (n_27278), .Y (n_28296));
AOI21X1 g109470(.A0 (n_26827), .A1 (n_26553), .B0 (n_27266), .Y(n_28295));
OAI21X1 g109482(.A0 (n_26180), .A1 (n_28747), .B0 (n_27285), .Y(n_28294));
MX2X1 g109489(.A (n_19691), .B (n_19690), .S0 (n_26625), .Y(n_29083));
NOR2X1 g109498(.A (n_26507), .B (n_27075), .Y (n_28293));
NOR2X1 g109499(.A (n_26506), .B (n_27073), .Y (n_28292));
NOR2X1 g109502(.A (n_19528), .B (n_27056), .Y (n_28291));
OAI21X1 g107290(.A0 (n_26877), .A1 (n_25623), .B0 (n_31628), .Y(n_28290));
NAND2X1 g109508(.A (n_34312), .B (n_28276), .Y (n_28289));
NAND2X1 g109511(.A (n_34312), .B (n_28267), .Y (n_28288));
NOR2X1 g109513(.A (n_27047), .B (n_10853), .Y (n_28287));
NOR2X1 g109514(.A (n_10089), .B (n_27046), .Y (n_28286));
NAND2X1 g109517(.A (n_34312), .B (n_28260), .Y (n_28285));
NOR2X1 g109518(.A (n_30445), .B (n_27058), .Y (n_28284));
NOR2X1 g109537(.A (n_27168), .B (n_24427), .Y (n_28283));
OAI21X1 g107312(.A0 (n_26861), .A1 (n_25619), .B0 (n_30569), .Y(n_28282));
NAND2X1 g109607(.A (n_28279), .B (n_28785), .Y (n_28281));
NAND2X1 g109609(.A (n_28279), .B (n_28798), .Y (n_28280));
NAND2X1 g109610(.A (n_28279), .B (n_28791), .Y (n_35091));
NAND2X1 g109615(.A (n_28276), .B (n_28275), .Y (n_28277));
NAND2X1 g109622(.A (n_28265), .B (n_18399), .Y (n_28274));
AOI21X1 g109625(.A0 (n_21245), .A1 (n_22139), .B0 (n_27155), .Y(n_28273));
NAND2X1 g109643(.A (n_28246), .B (n_27707), .Y (n_29760));
NAND2X1 g109647(.A (n_28270), .B (n_28785), .Y (n_32081));
NAND2X1 g109650(.A (n_28270), .B (n_28798), .Y (n_28271));
NAND2X1 g109651(.A (n_28270), .B (n_28791), .Y (n_35093));
NAND2X1 g109656(.A (n_28267), .B (n_28275), .Y (n_28268));
NAND2X1 g109660(.A (n_28265), .B (n_23270), .Y (n_28266));
NOR2X1 g109677(.A (n_28315), .B (n_8678), .Y (n_28263));
NAND2X1 g109679(.A (n_35201), .B (n_28785), .Y (n_35905));
NAND2X1 g109684(.A (n_28260), .B (n_10808), .Y (n_28261));
NAND2X1 g109686(.A (n_28265), .B (n_32728), .Y (n_28259));
NAND2X1 g109706(.A (n_35197), .B (n_28785), .Y (n_28258));
NAND2X1 g109714(.A (n_28254), .B (n_34753), .Y (n_28256));
NAND2X1 g109715(.A (n_28254), .B (n_28785), .Y (n_28255));
NOR2X1 g109716(.A (n_28252), .B (n_8382), .Y (n_28253));
NOR2X1 g109717(.A (n_28252), .B (n_8678), .Y (n_28251));
NAND2X1 g109720(.A (n_28265), .B (n_26866), .Y (n_28250));
OAI21X1 g107390(.A0 (n_8589), .A1 (n_31480), .B0 (n_27186), .Y(n_28249));
NAND2X1 g107393(.A (n_27136), .B (n_25830), .Y (n_28248));
NAND2X1 g109754(.A (n_27687), .B (n_27628), .Y (n_28883));
NAND2X1 g109755(.A (n_14799), .B (n_28246), .Y (n_28247));
INVX1 g109760(.A (n_28342), .Y (n_28245));
AOI21X1 g109782(.A0 (n_21244), .A1 (n_22139), .B0 (n_27152), .Y(n_28244));
AOI21X1 g109789(.A0 (n_18595), .A1 (n_22139), .B0 (n_27151), .Y(n_28242));
INVX1 g109804(.A (n_28344), .Y (n_28241));
NOR2X1 g109829(.A (n_27103), .B (n_13764), .Y (n_28240));
AOI21X1 g109843(.A0 (n_29068), .A1 (n_27651), .B0 (n_25179), .Y(n_28239));
NAND2X1 g107432(.A (n_27079), .B (n_25450), .Y (n_28238));
NAND3X1 g109887(.A (n_9571), .B (n_26536), .C (n_26131), .Y(n_28237));
NOR2X1 g109889(.A (n_9130), .B (n_27048), .Y (n_28236));
NOR2X1 g109898(.A (n_26524), .B (n_27051), .Y (n_28235));
NOR2X1 g109910(.A (n_26115), .B (n_27050), .Y (n_28234));
NAND2X1 g109912(.A (n_34803), .B (n_26654), .Y (n_28233));
OAI21X1 g109920(.A0 (n_26498), .A1 (n_8718), .B0 (n_21715), .Y(n_28232));
AOI21X1 g109926(.A0 (n_24925), .A1 (n_27634), .B0 (n_27074), .Y(n_28230));
AOI21X1 g109941(.A0 (n_27100), .A1 (n_27619), .B0 (n_25848), .Y(n_28229));
OAI21X1 g109946(.A0 (n_26497), .A1 (n_33807), .B0 (n_21696), .Y(n_28228));
OAI21X1 g109948(.A0 (n_26496), .A1 (n_8718), .B0 (n_21724), .Y(n_28226));
NAND3X1 g109953(.A (n_9605), .B (n_26533), .C (n_26107), .Y(n_28225));
NOR2X1 g109954(.A (n_27088), .B (n_27071), .Y (n_28224));
NOR2X1 g109956(.A (n_9104), .B (n_27044), .Y (n_28223));
INVX1 g109962(.A (n_28459), .Y (n_28222));
INVX1 g109964(.A (n_28432), .Y (n_28221));
INVX1 g109970(.A (n_28219), .Y (n_28220));
INVX1 g109971(.A (n_28219), .Y (n_28218));
INVX1 g109972(.A (n_28219), .Y (n_28217));
NOR2X1 g109992(.A (n_27086), .B (n_14984), .Y (n_28216));
NAND2X1 g110005(.A (n_27146), .B (n_27718), .Y (n_28918));
NAND2X1 g110007(.A (n_27144), .B (n_28215), .Y (n_28940));
NAND2X1 g110008(.A (n_27143), .B (n_28215), .Y (n_29396));
NAND3X1 g107509(.A (n_21631), .B (n_24829), .C (n_26478), .Y(n_29438));
NAND2X1 g110011(.A (n_27141), .B (n_28213), .Y (n_28214));
INVX1 g110013(.A (n_28471), .Y (n_28212));
NOR2X1 g107510(.A (n_6814), .B (n_27195), .Y (n_28211));
INVX1 g110015(.A (n_28444), .Y (n_28210));
INVX1 g110019(.A (n_28208), .Y (n_28209));
INVX2 g110021(.A (n_28208), .Y (n_28899));
INVX1 g110027(.A (n_28464), .Y (n_28206));
NAND2X1 g110044(.A (n_27128), .B (n_28205), .Y (n_28934));
NAND2X1 g110045(.A (n_27126), .B (n_28205), .Y (n_29390));
NAND2X1 g110047(.A (n_27122), .B (n_28204), .Y (n_29839));
NAND2X1 g110053(.A (n_27093), .B (n_27705), .Y (n_28924));
NAND2X1 g110056(.A (n_27115), .B (n_27709), .Y (n_28931));
INVX1 g110057(.A (n_28425), .Y (n_28203));
NAND2X1 g110059(.A (n_27114), .B (n_28202), .Y (n_28929));
NAND2X1 g110060(.A (n_27112), .B (n_28202), .Y (n_28891));
NAND2X1 g110061(.A (n_27108), .B (n_19492), .Y (n_28927));
INVX1 g110063(.A (n_28423), .Y (n_28201));
INVX1 g110068(.A (n_28416), .Y (n_28200));
INVX1 g110070(.A (n_28198), .Y (n_28199));
INVX1 g110072(.A (n_28198), .Y (n_28770));
INVX1 g110082(.A (n_28398), .Y (n_28197));
NAND2X1 g110084(.A (n_27092), .B (n_28196), .Y (n_28922));
NAND2X1 g110086(.A (n_27090), .B (n_28196), .Y (n_28870));
NAND2X1 g110092(.A (n_27085), .B (n_28195), .Y (n_28905));
INVX1 g110093(.A (n_28453), .Y (n_28194));
INVX1 g110095(.A (n_28390), .Y (n_28193));
INVX1 g110097(.A (n_28449), .Y (n_28192));
INVX1 g110099(.A (n_28380), .Y (n_28191));
INVX1 g110105(.A (n_27697), .Y (n_28190));
NAND2X1 g110130(.A (n_27138), .B (n_26673), .Y (n_28187));
NAND2X1 g110134(.A (n_27110), .B (n_19850), .Y (n_28186));
NAND2X1 g110136(.A (n_27154), .B (n_9585), .Y (n_28185));
NAND2X1 g110146(.A (n_27078), .B (n_27762), .Y (n_28879));
INVX1 g110148(.A (n_28406), .Y (n_28184));
NAND2X1 g110157(.A (n_27097), .B (n_27756), .Y (n_28759));
INVX1 g110162(.A (n_28181), .Y (n_28757));
NAND2X1 g110164(.A (n_27150), .B (n_9566), .Y (n_28180));
NAND2X1 g110167(.A (n_27147), .B (n_26718), .Y (n_28179));
NAND2X1 g110177(.A (n_27095), .B (n_26704), .Y (n_28178));
AOI21X1 g110186(.A0 (n_26017), .A1 (n_33494), .B0 (n_27159), .Y(n_28177));
AOI21X1 g110187(.A0 (n_27235), .A1 (n_33494), .B0 (n_27157), .Y(n_28176));
AOI21X1 g107569(.A0 (n_10763), .A1 (n_26471), .B0 (n_349), .Y(n_28175));
NAND2X1 g110214(.A (n_26725), .B (n_27179), .Y (n_28174));
NAND2X1 g110219(.A (n_26729), .B (n_27181), .Y (n_28173));
NAND2X1 g110226(.A (n_26727), .B (n_27180), .Y (n_28172));
AOI21X1 g110231(.A0 (n_27658), .A1 (n_26238), .B0 (n_27178), .Y(n_28171));
OAI21X1 g107617(.A0 (n_26461), .A1 (n_25312), .B0 (n_31160), .Y(n_28169));
NAND2X2 g107750(.A (n_26996), .B (n_12968), .Y (n_28168));
OAI21X1 g107768(.A0 (n_26439), .A1 (n_25313), .B0 (n_31398), .Y(n_28167));
NAND2X1 g110634(.A (n_28165), .B (n_8954), .Y (n_28166));
NAND2X1 g110732(.A (n_28165), .B (n_30636), .Y (n_28163));
NOR2X1 g107812(.A (n_27001), .B (n_26436), .Y (n_28162));
NAND2X1 g110742(.A (n_28159), .B (n_28136), .Y (n_28161));
NAND2X1 g110748(.A (n_28159), .B (n_28158), .Y (n_28160));
NOR2X1 g107824(.A (n_30050), .B (n_28155), .Y (n_28157));
NOR2X1 g107825(.A (n_28155), .B (n_29172), .Y (n_28156));
NAND2X1 g107828(.A (n_21666), .B (n_28151), .Y (n_29257));
NAND2X1 g107841(.A (n_28151), .B (n_15297), .Y (n_28152));
NAND2X1 g107845(.A (n_26997), .B (n_31696), .Y (n_28150));
INVX1 g110865(.A (n_28146), .Y (n_28147));
OAI21X1 g110878(.A0 (n_25592), .A1 (n_8319), .B0 (n_27024), .Y(n_28144));
NAND2X1 g110884(.A (n_20279), .B (n_27026), .Y (n_28143));
INVX1 g110903(.A (n_28809), .Y (n_28142));
INVX1 g110907(.A (n_28140), .Y (n_28141));
INVX1 g110927(.A (n_28138), .Y (n_28698));
NAND2X1 g110984(.A (n_27019), .B (n_28136), .Y (n_28137));
NOR2X1 g107928(.A (n_9939), .B (n_27009), .Y (n_28135));
OAI21X1 g110999(.A0 (n_27565), .A1 (n_8322), .B0 (n_20284), .Y(n_28134));
NOR2X1 g107939(.A (n_9925), .B (n_27007), .Y (n_28133));
NAND2X1 g111073(.A (n_26137), .B (n_27016), .Y (n_28132));
OAI21X1 g111077(.A0 (n_26480), .A1 (n_8285), .B0 (n_26156), .Y(n_28131));
NAND3X1 g107970(.A (n_7533), .B (n_26474), .C (n_7552), .Y (n_28130));
AOI22X1 g107979(.A0 (n_26470), .A1 (n_31878), .B0 (n_9353), .B1(n_31495), .Y (n_28129));
NOR2X1 g108009(.A (n_26475), .B (n_27012), .Y (n_28128));
NAND2X1 g111287(.A (n_28126), .B (n_24526), .Y (n_28127));
NAND2X1 g108048(.A (n_27000), .B (n_28125), .Y (n_29254));
NAND2X1 g108062(.A (n_27004), .B (n_28124), .Y (n_29250));
AOI21X1 g108068(.A0 (n_14939), .A1 (n_27544), .B0 (n_29725), .Y(n_28123));
AOI21X1 g108070(.A0 (n_32869), .A1 (n_28053), .B0 (n_13929), .Y(n_28676));
NAND2X1 g108093(.A (n_6653), .B (n_27014), .Y (n_28122));
AOI21X1 g108137(.A0 (n_10392), .A1 (n_26902), .B0 (n_7058), .Y(n_28121));
NAND3X1 g108138(.A (n_19654), .B (n_26331), .C (n_26873), .Y(n_28120));
NAND3X1 g108151(.A (n_10096), .B (n_21689), .C (n_26835), .Y(n_28119));
NAND3X1 g108154(.A (n_11134), .B (n_26335), .C (n_26885), .Y(n_28118));
NOR2X1 g108162(.A (n_25130), .B (n_26967), .Y (n_28117));
NOR2X1 g108163(.A (n_27172), .B (n_25566), .Y (n_28116));
NOR2X1 g108169(.A (n_27166), .B (n_25564), .Y (n_28115));
NOR2X1 g108172(.A (n_27170), .B (n_25560), .Y (n_28114));
NAND2X1 g108176(.A (n_28107), .B (n_26160), .Y (n_28113));
NAND2X1 g108177(.A (n_28105), .B (n_26160), .Y (n_28111));
NAND2X1 g108181(.A (n_28103), .B (n_34952), .Y (n_32891));
NAND2X1 g108189(.A (n_28107), .B (n_29619), .Y (n_28108));
NAND2X1 g108192(.A (n_28105), .B (n_29619), .Y (n_28106));
NAND2X1 g108195(.A (n_28103), .B (n_28485), .Y (n_28104));
NAND2X1 g108197(.A (n_33335), .B (n_28485), .Y (n_28101));
NAND2X1 g108257(.A (n_28091), .B (n_22406), .Y (n_28099));
NAND2X1 g108203(.A (n_28107), .B (n_28808), .Y (n_28098));
NAND2X1 g108206(.A (n_28105), .B (n_28808), .Y (n_28097));
NAND2X1 g108209(.A (n_28103), .B (n_33378), .Y (n_28096));
NOR2X1 g108227(.A (n_26911), .B (n_14601), .Y (n_28094));
NAND2X1 g108237(.A (n_27386), .B (n_34753), .Y (n_28093));
NAND2X1 g108239(.A (n_17719), .B (n_28091), .Y (n_28092));
NOR2X1 g108242(.A (n_25135), .B (n_26927), .Y (n_28090));
OAI21X1 g108243(.A0 (n_26908), .A1 (n_26699), .B0 (n_27485), .Y(n_28089));
CLKBUFX1 gbuf_d_363(.A(n_27190), .Y(d_out_363));
CLKBUFX1 gbuf_q_363(.A(q_in_363), .Y(n_565));
NOR2X1 g108260(.A (n_25133), .B (n_26926), .Y (n_28088));
NAND2X1 g108271(.A (n_27378), .B (n_34753), .Y (n_32890));
NAND2X1 g108274(.A (n_28091), .B (n_32764), .Y (n_28086));
NAND2X1 g108325(.A (n_18936), .B (n_28081), .Y (n_29170));
NAND2X1 g108334(.A (n_28084), .B (n_28083), .Y (n_29156));
NAND2X1 g108335(.A (n_28081), .B (n_14725), .Y (n_28082));
AOI21X1 g108375(.A0 (n_29068), .A1 (n_27495), .B0 (n_26098), .Y(n_28080));
AOI21X1 g108383(.A0 (n_30438), .A1 (n_27493), .B0 (n_26075), .Y(n_28079));
NAND3X1 g108402(.A (n_26770), .B (n_26279), .C (n_26798), .Y(n_28078));
NOR2X1 g108412(.A (n_25071), .B (n_26937), .Y (n_28077));
NAND4X1 g108419(.A (n_19946), .B (n_24726), .C (n_26223), .D(n_23355), .Y (n_28076));
OAI21X1 g108442(.A0 (n_27475), .A1 (n_29150), .B0 (n_21206), .Y(n_28075));
NAND3X1 g108447(.A (n_10157), .B (n_26328), .C (n_26864), .Y(n_28074));
AOI21X1 g108458(.A0 (n_24925), .A1 (n_27461), .B0 (n_26934), .Y(n_28073));
AOI21X1 g108460(.A0 (n_24925), .A1 (n_27459), .B0 (n_26933), .Y(n_28072));
NAND2X1 g108255(.A (n_27382), .B (n_34753), .Y (n_32115));
NAND4X1 g108466(.A (n_19863), .B (n_24723), .C (n_26218), .D(n_23571), .Y (n_28069));
OAI21X1 g108469(.A0 (n_9843), .A1 (n_31680), .B0 (n_26980), .Y(n_28068));
AOI21X1 g108471(.A0 (n_27100), .A1 (n_27436), .B0 (n_26921), .Y(n_28067));
NAND3X1 g108474(.A (n_10210), .B (n_26326), .C (n_26833), .Y(n_28066));
NAND2X1 g108494(.A (n_26966), .B (n_13171), .Y (n_28568));
NAND2X1 g108495(.A (n_26964), .B (n_13171), .Y (n_29201));
NOR2X1 g108509(.A (n_7088), .B (n_26983), .Y (n_28065));
NAND2X1 g108535(.A (n_26975), .B (n_28064), .Y (n_35917));
NAND2X1 g108537(.A (n_26974), .B (n_28064), .Y (n_29192));
NAND2X1 g108563(.A (n_26972), .B (n_28063), .Y (n_29197));
NAND2X1 g108565(.A (n_26970), .B (n_28063), .Y (n_29188));
INVX1 g108581(.A (n_28738), .Y (n_32299));
NAND2X1 g108591(.A (n_26962), .B (n_28061), .Y (n_29194));
NAND2X1 g108593(.A (n_26961), .B (n_28061), .Y (n_29178));
OAI21X1 g108609(.A0 (n_26765), .A1 (n_35546), .B0 (n_28058), .Y(n_28060));
AOI21X1 g108617(.A0 (n_35688), .A1 (n_28136), .B0 (n_20853), .Y(n_28057));
NAND2X1 g106931(.A (n_7988), .B (n_28666), .Y (n_28056));
OAI21X1 g108626(.A0 (n_26765), .A1 (n_13736), .B0 (n_28054), .Y(n_29162));
AOI21X1 g108633(.A0 (n_33644), .A1 (n_28053), .B0 (n_13921), .Y(n_28536));
AOI21X1 g108635(.A0 (n_35649), .A1 (n_28053), .B0 (n_13920), .Y(n_28535));
INVX1 g108642(.A (n_28052), .Y (n_28533));
OAI21X1 g108688(.A0 (n_26793), .A1 (n_31275), .B0 (n_6588), .Y(n_28051));
OAI21X1 g108693(.A0 (n_26788), .A1 (n_31273), .B0 (n_6560), .Y(n_28050));
INVX1 g108721(.A (n_33626), .Y (n_28049));
NOR2X1 g108733(.A (n_26819), .B (n_27072), .Y (n_28048));
AOI21X1 g108742(.A0 (n_8609), .A1 (n_26753), .B0 (n_34676), .Y(n_28047));
NAND2X1 g108744(.A (n_27241), .B (n_31698), .Y (n_28046));
NAND3X1 g108746(.A (n_18025), .B (n_26716), .C (n_26298), .Y(n_28045));
NAND3X1 g108747(.A (n_18569), .B (n_26661), .C (n_26715), .Y(n_28044));
NAND4X1 g108749(.A (n_27133), .B (n_26712), .C (n_19642), .D(n_10825), .Y (n_28043));
NAND3X1 g108752(.A (n_27238), .B (n_26616), .C (n_20866), .Y(n_28042));
NAND3X1 g108754(.A (n_27237), .B (n_26258), .C (n_20861), .Y(n_28041));
NAND2X1 g108764(.A (n_34312), .B (n_28003), .Y (n_28040));
NAND3X1 g108765(.A (n_10998), .B (n_26721), .C (n_25965), .Y(n_28039));
NAND4X1 g108766(.A (n_27148), .B (n_26720), .C (n_10833), .D(n_10040), .Y (n_28038));
NAND2X1 g108771(.A (n_34312), .B (n_27990), .Y (n_28037));
NOR2X1 g108773(.A (n_27201), .B (n_10852), .Y (n_28036));
NAND2X1 g108774(.A (n_34312), .B (n_28034), .Y (n_28035));
NOR2X1 g108796(.A (n_27174), .B (n_25216), .Y (n_35134));
NOR2X1 g108798(.A (n_27167), .B (n_25215), .Y (n_28032));
NOR2X1 g108799(.A (n_27171), .B (n_24824), .Y (n_28031));
NAND2X1 g108815(.A (n_34770), .B (n_28023), .Y (n_28030));
NAND2X1 g108821(.A (n_29065), .B (n_28018), .Y (n_28028));
NOR2X1 g108823(.A (n_34501), .B (n_8668), .Y (n_28027));
NAND2X1 g108829(.A (n_28025), .B (n_29925), .Y (n_28026));
NAND2X1 g108842(.A (n_28023), .B (n_34709), .Y (n_28024));
NAND2X1 g108847(.A (n_8966), .B (n_28020), .Y (n_28021));
NAND2X1 g108850(.A (n_28018), .B (n_29925), .Y (n_28019));
NOR2X1 g108856(.A (n_34501), .B (n_33340), .Y (n_28017));
NAND2X1 g108867(.A (n_28025), .B (n_28013), .Y (n_28014));
NAND3X1 g108870(.A (n_26668), .B (n_25994), .C (n_26755), .Y(n_28012));
NAND2X1 g108878(.A (n_28593), .B (n_28013), .Y (n_28011));
NAND2X1 g108885(.A (n_28023), .B (n_28013), .Y (n_28009));
NAND2X1 g108895(.A (n_28018), .B (n_28013), .Y (n_28008));
NAND3X1 g108899(.A (n_24832), .B (n_26624), .C (n_24491), .Y(n_28007));
NAND2X1 g108906(.A (n_28003), .B (n_24526), .Y (n_28004));
NAND2X1 g108907(.A (n_28003), .B (n_28791), .Y (n_28001));
NAND2X1 g108910(.A (n_27986), .B (n_27999), .Y (n_28000));
AND2X1 g108917(.A (n_27995), .B (n_33494), .Y (n_27998));
NAND2X1 g108918(.A (n_27995), .B (n_27956), .Y (n_27996));
NAND2X1 g108919(.A (n_27995), .B (n_27993), .Y (n_27994));
NAND2X1 g108920(.A (n_27995), .B (n_29445), .Y (n_27992));
NAND2X1 g108924(.A (n_27990), .B (n_24526), .Y (n_27991));
NAND2X1 g108925(.A (n_27990), .B (n_28791), .Y (n_27989));
NAND2X1 g108931(.A (n_35055), .B (n_22831), .Y (n_27988));
NAND2X1 g108934(.A (n_27986), .B (n_22406), .Y (n_27987));
NAND2X1 g108935(.A (n_27961), .B (n_26315), .Y (n_27985));
NAND2X1 g108944(.A (n_27983), .B (n_25554), .Y (n_27984));
AOI21X1 g108945(.A0 (n_26763), .A1 (n_26680), .B0 (n_27008), .Y(n_27982));
NAND2X1 g108952(.A (n_28034), .B (n_34753), .Y (n_27981));
NAND2X1 g108954(.A (n_27714), .B (n_10808), .Y (n_27980));
NAND2X1 g108956(.A (n_27986), .B (n_32685), .Y (n_27979));
NOR2X1 g108961(.A (n_26297), .B (n_27249), .Y (n_27978));
NAND2X1 g108964(.A (n_29341), .B (n_27912), .Y (n_27977));
AND2X1 g108965(.A (n_27974), .B (n_26662), .Y (n_27976));
NAND2X1 g108966(.A (n_27974), .B (n_26665), .Y (n_27975));
NAND2X1 g108967(.A (n_27974), .B (n_27993), .Y (n_27973));
NAND2X1 g108968(.A (n_27974), .B (n_28431), .Y (n_27972));
NAND2X1 g108975(.A (n_26377), .B (n_10808), .Y (n_27971));
NAND2X1 g108978(.A (n_27725), .B (n_10808), .Y (n_27970));
NOR2X1 g108981(.A (n_27967), .B (n_14159), .Y (n_27968));
NAND2X1 g108985(.A (n_27986), .B (n_27470), .Y (n_27963));
NAND2X1 g108990(.A (n_27961), .B (n_35054), .Y (n_27962));
NAND2X1 g108994(.A (n_27983), .B (n_23192), .Y (n_27960));
NAND2X1 g108999(.A (n_27957), .B (n_28890), .Y (n_27959));
NAND2X1 g109000(.A (n_27957), .B (n_27956), .Y (n_27958));
NAND2X1 g109001(.A (n_27957), .B (n_33513), .Y (n_27955));
NAND2X1 g109002(.A (n_27957), .B (n_30180), .Y (n_27954));
NAND2X1 g109015(.A (n_35055), .B (n_25193), .Y (n_27952));
NAND2X1 g109019(.A (n_27961), .B (n_27950), .Y (n_27951));
NAND3X1 g109023(.A (n_27243), .B (n_26241), .C (n_20934), .Y(n_27949));
NAND2X1 g109030(.A (n_27983), .B (n_26631), .Y (n_27948));
NAND2X1 g109043(.A (n_8284), .B (n_27945), .Y (n_27947));
NAND2X1 g109044(.A (n_26255), .B (n_27945), .Y (n_27946));
NAND2X1 g109046(.A (n_29427), .B (n_27945), .Y (n_27944));
NAND3X1 g109058(.A (n_25860), .B (n_26552), .C (n_15150), .Y(n_27943));
NAND2X1 g109069(.A (n_27941), .B (n_33738), .Y (n_27942));
NAND2X1 g109075(.A (n_30171), .B (n_27938), .Y (n_27940));
NAND2X1 g109076(.A (n_27938), .B (n_8922), .Y (n_27939));
NAND2X1 g109077(.A (n_27938), .B (n_29684), .Y (n_27937));
NAND2X1 g109078(.A (n_27907), .B (n_8954), .Y (n_27936));
NOR2X1 g109090(.A (n_27189), .B (n_10874), .Y (n_27935));
NAND2X1 g109096(.A (n_27933), .B (n_29505), .Y (n_27934));
NAND2X1 g109097(.A (n_27933), .B (n_26132), .Y (n_27931));
NAND2X1 g109103(.A (n_27682), .B (n_30454), .Y (n_27930));
NAND2X1 g109110(.A (n_27916), .B (n_28158), .Y (n_27929));
NAND2X1 g109111(.A (n_27926), .B (n_28890), .Y (n_27928));
NAND2X1 g109112(.A (n_27926), .B (n_33513), .Y (n_27927));
NAND2X1 g109113(.A (n_27926), .B (n_27956), .Y (n_27925));
NAND2X1 g109114(.A (n_27926), .B (n_30180), .Y (n_27924));
NAND2X1 g109116(.A (n_27233), .B (n_13189), .Y (n_27923));
NOR2X1 g109121(.A (n_26382), .B (n_27265), .Y (n_27922));
NAND2X1 g109128(.A (n_27920), .B (n_28158), .Y (n_27921));
NAND2X1 g109129(.A (n_27920), .B (n_26238), .Y (n_27919));
NAND2X1 g109131(.A (n_27916), .B (n_26238), .Y (n_27917));
NAND2X1 g109137(.A (n_28020), .B (n_27902), .Y (n_27915));
NAND2X1 g109138(.A (n_28020), .B (n_26238), .Y (n_27914));
NAND2X1 g109139(.A (n_27614), .B (n_27912), .Y (n_27913));
NAND2X1 g109140(.A (n_8284), .B (n_27912), .Y (n_27911));
NAND2X1 g109150(.A (n_35055), .B (n_27091), .Y (n_27910));
NAND2X1 g109154(.A (n_27961), .B (n_27422), .Y (n_27909));
NAND2X1 g109158(.A (n_27907), .B (n_26238), .Y (n_27908));
AND2X1 g109161(.A (n_27905), .B (n_29405), .Y (n_27906));
NAND2X1 g109162(.A (n_27905), .B (n_26238), .Y (n_27904));
NAND2X1 g109163(.A (n_27941), .B (n_27902), .Y (n_27903));
AND2X1 g109166(.A (n_27907), .B (n_29405), .Y (n_27901));
NAND2X1 g109179(.A (n_26387), .B (n_27240), .Y (n_27900));
NAND4X1 g109180(.A (n_27315), .B (n_24419), .C (n_24907), .D(n_24926), .Y (n_27899));
NAND3X1 g109187(.A (n_26219), .B (n_26551), .C (n_15172), .Y(n_27898));
NAND2X1 g109192(.A (n_27895), .B (n_29411), .Y (n_27897));
NAND2X1 g109195(.A (n_27895), .B (n_8954), .Y (n_27896));
NOR2X1 g109197(.A (n_28524), .B (n_25881), .Y (n_27894));
NAND2X1 g109202(.A (n_27895), .B (n_29405), .Y (n_27892));
NAND2X1 g109203(.A (n_27895), .B (n_30636), .Y (n_27891));
NAND2X1 g109207(.A (n_27886), .B (n_30636), .Y (n_27890));
NAND2X1 g109208(.A (n_27883), .B (n_33991), .Y (n_27889));
NAND2X1 g109210(.A (n_33732), .B (n_33991), .Y (n_32230));
NAND2X1 g109225(.A (n_27886), .B (n_29405), .Y (n_27887));
NAND2X1 g109226(.A (n_27886), .B (n_33738), .Y (n_27885));
NAND2X1 g109227(.A (n_27883), .B (n_28158), .Y (n_27884));
NAND2X1 g109229(.A (n_33732), .B (n_29155), .Y (n_27882));
NAND4X1 g109233(.A (n_27239), .B (n_24753), .C (n_14878), .D(n_24742), .Y (n_27880));
AOI21X1 g109239(.A0 (n_27825), .A1 (n_30557), .B0 (n_21730), .Y(n_27879));
NOR2X1 g109246(.A (n_26675), .B (n_27212), .Y (n_27878));
AOI21X1 g109248(.A0 (n_27782), .A1 (n_28791), .B0 (n_19616), .Y(n_27877));
NAND3X1 g109250(.A (n_10206), .B (n_26713), .C (n_26293), .Y(n_27876));
AOI21X1 g109252(.A0 (n_27822), .A1 (n_29040), .B0 (n_21721), .Y(n_27875));
NOR2X1 g109253(.A (n_26658), .B (n_27211), .Y (n_27874));
NOR2X1 g109260(.A (n_10192), .B (n_27200), .Y (n_27873));
AOI21X1 g109267(.A0 (n_27820), .A1 (n_30557), .B0 (n_21714), .Y(n_27872));
OAI21X1 g109268(.A0 (n_26636), .A1 (n_31410), .B0 (n_8604), .Y(n_27871));
NAND2X1 g109271(.A (n_27284), .B (n_26390), .Y (n_27870));
NOR2X1 g109272(.A (n_9554), .B (n_27194), .Y (n_27869));
NAND2X1 g109279(.A (n_27282), .B (n_29505), .Y (n_27868));
NAND3X1 g109286(.A (n_9054), .B (n_26619), .C (n_20883), .Y(n_27867));
NOR2X1 g109288(.A (n_9921), .B (n_27352), .Y (n_27866));
AOI21X1 g109299(.A0 (n_27817), .A1 (n_30557), .B0 (n_21722), .Y(n_27865));
OAI21X1 g109302(.A0 (n_26601), .A1 (n_31482), .B0 (n_9919), .Y(n_27864));
NOR2X1 g109303(.A (n_9072), .B (n_27199), .Y (n_27863));
NAND2X1 g109304(.A (n_27287), .B (n_27399), .Y (n_29096));
INVX1 g109305(.A (n_27861), .Y (n_27862));
AOI21X1 g109312(.A0 (n_27803), .A1 (n_27770), .B0 (n_15119), .Y(n_29093));
OAI21X1 g109313(.A0 (n_26697), .A1 (n_30935), .B0 (n_8615), .Y(n_27859));
OAI21X1 g109314(.A0 (n_26382), .A1 (n_26550), .B0 (n_26779), .Y(n_27858));
NAND4X1 g109315(.A (n_27316), .B (n_24085), .C (n_24908), .D(n_24928), .Y (n_27857));
AOI21X1 g107207(.A0 (n_10759), .A1 (n_26488), .B0 (n_31343), .Y(n_27856));
NAND2X1 g107208(.A (n_27039), .B (n_1054), .Y (n_27855));
NAND3X1 g109327(.A (n_24807), .B (n_26603), .C (n_24808), .Y(n_27854));
NOR2X1 g109337(.A (n_10395), .B (n_27351), .Y (n_27853));
INVX1 g109343(.A (n_28653), .Y (n_27852));
NAND2X1 g109349(.A (n_27308), .B (n_27388), .Y (n_29103));
INVX1 g109355(.A (n_28651), .Y (n_27851));
NAND2X1 g109361(.A (n_27301), .B (n_24673), .Y (n_29100));
NAND2X1 g109371(.A (n_27294), .B (n_27379), .Y (n_29098));
INVX1 g109372(.A (n_27849), .Y (n_27850));
INVX1 g109383(.A (n_28647), .Y (n_27847));
NAND2X1 g109388(.A (n_27280), .B (n_19866), .Y (n_27846));
OAI21X1 g109396(.A0 (n_35196), .A1 (n_10276), .B0 (n_27320), .Y(n_27845));
NAND2X1 g109398(.A (n_27270), .B (n_28319), .Y (n_27844));
OAI21X1 g109403(.A0 (n_26583), .A1 (n_13903), .B0 (n_27842), .Y(n_27843));
AOI21X1 g107243(.A0 (n_26848), .A1 (n_26071), .B0 (n_8070), .Y(n_27841));
NAND2X1 g109437(.A (n_27274), .B (n_26548), .Y (n_27840));
AOI21X1 g109439(.A0 (n_27766), .A1 (n_28053), .B0 (n_13923), .Y(n_28306));
NAND2X1 g109441(.A (n_27273), .B (n_26548), .Y (n_27839));
NAND2X1 g109461(.A (n_26847), .B (n_19867), .Y (n_27838));
NAND2X1 g109468(.A (n_26858), .B (n_20962), .Y (n_27837));
NAND2X1 g109471(.A (n_26818), .B (n_19887), .Y (n_27836));
OAI21X1 g109472(.A0 (n_26180), .A1 (n_33734), .B0 (n_19888), .Y(n_27835));
NAND4X1 g107272(.A (n_25818), .B (n_20954), .C (n_25567), .D(n_25725), .Y (n_27834));
NAND2X1 g109481(.A (n_26339), .B (n_26904), .Y (n_27833));
OAI21X1 g109484(.A0 (n_26282), .A1 (n_28747), .B0 (n_26836), .Y(n_27832));
NAND2X1 g109485(.A (n_26337), .B (n_26903), .Y (n_27831));
AOI21X1 g109486(.A0 (n_26428), .A1 (n_26238), .B0 (n_26901), .Y(n_35918));
NAND2X2 g109487(.A (n_26418), .B (n_26886), .Y (n_28634));
NAND2X2 g109492(.A (n_35929), .B (n_35930), .Y (n_28606));
NAND3X1 g109501(.A (n_19003), .B (n_25815), .C (n_26110), .Y(n_27829));
NAND4X1 g109504(.A (n_26534), .B (n_18729), .C (n_23184), .D(n_24872), .Y (n_27828));
NAND3X1 g109507(.A (n_17278), .B (n_26133), .C (n_19215), .Y(n_27827));
NAND2X1 g109510(.A (n_34712), .B (n_27825), .Y (n_27826));
NAND2X1 g109512(.A (n_34312), .B (n_27789), .Y (n_27824));
NAND2X1 g109520(.A (n_34712), .B (n_27822), .Y (n_27823));
NAND2X1 g109522(.A (n_34712), .B (n_27820), .Y (n_27821));
OAI21X1 g109523(.A0 (n_26100), .A1 (n_25245), .B0 (n_24695), .Y(n_27819));
NAND2X1 g109526(.A (n_34712), .B (n_27817), .Y (n_27818));
NOR2X1 g109528(.A (n_19004), .B (n_26568), .Y (n_27816));
AOI21X1 g109531(.A0 (n_27743), .A1 (n_27162), .B0 (n_10616), .Y(n_27815));
NAND3X1 g109535(.A (n_26746), .B (n_14876), .C (n_23762), .Y(n_27814));
NAND3X1 g109538(.A (n_26741), .B (n_14380), .C (n_24619), .Y(n_27813));
NOR2X1 g109541(.A (n_26749), .B (n_24094), .Y (n_27812));
NOR2X1 g109542(.A (n_26743), .B (n_24092), .Y (n_27811));
NOR2X1 g109543(.A (n_26744), .B (n_24091), .Y (n_27810));
NAND2X1 g107315(.A (n_27040), .B (n_1054), .Y (n_27809));
NOR2X1 g109566(.A (n_26560), .B (n_8319), .Y (n_27807));
NOR2X1 g109571(.A (n_26557), .B (n_8319), .Y (n_27805));
NAND2X1 g109608(.A (n_27803), .B (n_26676), .Y (n_27804));
NAND2X1 g109617(.A (n_27800), .B (n_10808), .Y (n_27802));
NAND2X1 g109618(.A (n_27800), .B (n_28798), .Y (n_27801));
NAND2X1 g109619(.A (n_27800), .B (n_27798), .Y (n_27799));
NAND2X1 g109620(.A (n_27800), .B (n_26528), .Y (n_27797));
NAND4X1 g109628(.A (n_19943), .B (n_25625), .C (n_25660), .D(n_25648), .Y (n_27795));
NAND2X1 g109633(.A (n_26573), .B (n_24451), .Y (n_27794));
NAND2X1 g109639(.A (n_27825), .B (n_28431), .Y (n_27793));
NAND3X1 g109642(.A (n_26189), .B (n_26158), .C (n_25795), .Y(n_27792));
NAND2X1 g109649(.A (n_27771), .B (n_28441), .Y (n_27791));
NAND2X1 g109657(.A (n_27789), .B (n_10808), .Y (n_27790));
NAND2X1 g109668(.A (n_27803), .B (n_25554), .Y (n_27786));
NAND2X1 g109678(.A (n_27061), .B (n_34753), .Y (n_27784));
NAND2X1 g109685(.A (n_27782), .B (n_10808), .Y (n_27783));
NAND2X1 g109699(.A (n_27822), .B (n_24786), .Y (n_27778));
NAND3X1 g109702(.A (n_26186), .B (n_26152), .C (n_25761), .Y(n_27777));
NAND2X1 g109703(.A (n_27774), .B (n_28636), .Y (n_32103));
NAND2X1 g109704(.A (n_27774), .B (n_26213), .Y (n_27775));
NAND2X1 g109705(.A (n_27774), .B (n_27798), .Y (n_27773));
NAND2X1 g109708(.A (n_27771), .B (n_27770), .Y (n_27772));
NAND2X1 g109735(.A (n_27820), .B (n_28431), .Y (n_27769));
NAND2X1 g109741(.A (n_27771), .B (n_13274), .Y (n_27768));
NAND2X1 g109745(.A (n_27803), .B (n_24348), .Y (n_27767));
NAND2X1 g109751(.A (n_27766), .B (n_18546), .Y (n_28394));
NAND2X1 g109758(.A (n_27686), .B (n_27102), .Y (n_28411));
NAND2X1 g109759(.A (n_14973), .B (n_27764), .Y (n_27765));
NAND2X1 g109761(.A (n_27760), .B (n_27681), .Y (n_28342));
NAND2X1 g109778(.A (n_27764), .B (n_27711), .Y (n_28392));
NAND2X1 g109783(.A (n_27739), .B (n_35744), .Y (n_28401));
NAND2X1 g109784(.A (n_14577), .B (n_27757), .Y (n_27763));
NAND2X1 g109785(.A (n_27762), .B (n_27754), .Y (n_28376));
NAND2X1 g109787(.A (n_14745), .B (n_27760), .Y (n_27761));
NAND2X1 g109788(.A (n_27685), .B (n_27076), .Y (n_28372));
INVX1 g109800(.A (n_27883), .Y (n_27759));
NAND2X1 g109803(.A (n_27766), .B (n_35816), .Y (n_27758));
NAND2X2 g109805(.A (n_27757), .B (n_27756), .Y (n_28344));
NAND2X1 g109806(.A (n_27754), .B (n_14194), .Y (n_27755));
NAND2X1 g109810(.A (n_27817), .B (n_28431), .Y (n_27752));
NAND2X1 g109816(.A (n_29551), .B (n_25874), .Y (n_27751));
NAND2X1 g109819(.A (n_28347), .B (n_25874), .Y (n_27750));
NAND2X1 g109826(.A (n_27771), .B (n_27747), .Y (n_27748));
NAND3X1 g109830(.A (n_26183), .B (n_26154), .C (n_25806), .Y(n_27746));
OAI21X1 g109833(.A0 (n_24959), .A1 (n_25376), .B0 (n_26554), .Y(n_27745));
AOI21X1 g109836(.A0 (n_27743), .A1 (n_34801), .B0 (n_19527), .Y(n_27744));
NAND3X1 g109844(.A (n_26545), .B (n_23448), .C (n_15278), .Y(n_27742));
NAND3X1 g109850(.A (n_26543), .B (n_23446), .C (n_15264), .Y(n_27741));
NAND2X1 g109862(.A (n_27766), .B (n_35479), .Y (n_28396));
NAND2X1 g109868(.A (n_27739), .B (n_22021), .Y (n_28409));
AOI21X1 g109881(.A0 (n_27668), .A1 (n_27234), .B0 (n_19940), .Y(n_27738));
AOI21X1 g109884(.A0 (n_27665), .A1 (n_26665), .B0 (n_21373), .Y(n_32315));
NOR2X1 g109886(.A (n_9119), .B (n_26547), .Y (n_27736));
NAND3X1 g109888(.A (n_26130), .B (n_20295), .C (n_26128), .Y(n_27735));
OAI21X1 g109904(.A0 (n_26094), .A1 (n_33807), .B0 (n_19924), .Y(n_27734));
AOI21X1 g109908(.A0 (n_27676), .A1 (n_29040), .B0 (n_21367), .Y(n_27733));
NAND4X1 g109916(.A (n_26504), .B (n_18716), .C (n_23177), .D(n_24871), .Y (n_27732));
OAI21X1 g109918(.A0 (n_26088), .A1 (n_29381), .B0 (n_21716), .Y(n_27731));
OAI21X1 g109947(.A0 (n_26080), .A1 (n_29381), .B0 (n_21695), .Y(n_27730));
NOR2X1 g109949(.A (n_9068), .B (n_26546), .Y (n_27729));
NAND3X1 g109955(.A (n_26104), .B (n_20305), .C (n_26102), .Y(n_27728));
NAND2X1 g109963(.A (n_26650), .B (n_27727), .Y (n_28459));
NAND2X1 g109965(.A (n_26649), .B (n_27727), .Y (n_28432));
NAND2X1 g109966(.A (n_26647), .B (n_27230), .Y (n_28483));
INVX1 g109967(.A (n_27725), .Y (n_27726));
NAND2X2 g109973(.A (n_26646), .B (n_13175), .Y (n_28219));
NAND2X1 g109974(.A (n_26644), .B (n_13175), .Y (n_28481));
OAI21X1 g109981(.A0 (n_26382), .A1 (n_26076), .B0 (n_25452), .Y(n_27722));
OAI21X1 g109983(.A0 (n_26382), .A1 (n_25671), .B0 (n_26549), .Y(n_27721));
NAND2X1 g109993(.A (n_26702), .B (n_13667), .Y (n_28493));
INVX1 g109996(.A (n_34501), .Y (n_27720));
INVX1 g109999(.A (n_27920), .Y (n_27719));
NAND2X1 g110006(.A (n_26698), .B (n_27718), .Y (n_29049));
NAND2X1 g110014(.A (n_26694), .B (n_27717), .Y (n_28471));
NAND2X1 g110016(.A (n_26692), .B (n_27717), .Y (n_28444));
NAND2X1 g110017(.A (n_26691), .B (n_13650), .Y (n_28490));
NAND2X1 g110022(.A (n_26689), .B (n_27716), .Y (n_28208));
NAND2X1 g110023(.A (n_26688), .B (n_27716), .Y (n_29067));
INVX1 g110025(.A (n_29392), .Y (n_28207));
NAND2X1 g110028(.A (n_26687), .B (n_27222), .Y (n_28464));
NAND2X1 g110030(.A (n_26684), .B (n_27221), .Y (n_28511));
NAND2X1 g110031(.A (n_26671), .B (n_27220), .Y (n_28488));
INVX1 g110033(.A (n_27714), .Y (n_27715));
NAND2X1 g110036(.A (n_26670), .B (n_27219), .Y (n_28486));
AOI21X1 g110037(.A0 (n_33546), .A1 (n_26799), .B0 (n_26736), .Y(n_27712));
NAND2X1 g110039(.A (n_26683), .B (n_13180), .Y (n_28384));
NAND2X2 g110040(.A (n_26587), .B (n_27711), .Y (n_28451));
NAND2X1 g110051(.A (n_26652), .B (n_26376), .Y (n_29009));
NAND2X1 g110058(.A (n_26638), .B (n_27709), .Y (n_28425));
NAND2X1 g110062(.A (n_26635), .B (n_27708), .Y (n_28479));
NAND2X1 g110064(.A (n_26634), .B (n_27708), .Y (n_28423));
NAND2X1 g110065(.A (n_26633), .B (n_24299), .Y (n_28476));
NAND2X1 g110066(.A (n_26632), .B (n_24299), .Y (n_28420));
NAND2X1 g110069(.A (n_26630), .B (n_27217), .Y (n_28416));
NAND2X2 g110073(.A (n_26577), .B (n_27707), .Y (n_28198));
NAND2X1 g110075(.A (n_26621), .B (n_20923), .Y (n_27706));
NAND2X1 g110083(.A (n_26606), .B (n_27705), .Y (n_28398));
INVX2 g110088(.A (n_27916), .Y (n_27704));
NAND2X1 g110094(.A (n_26678), .B (n_27702), .Y (n_28453));
NAND2X1 g110096(.A (n_26600), .B (n_27702), .Y (n_28390));
NAND2X1 g110098(.A (n_26599), .B (n_13180), .Y (n_28449));
NAND2X1 g110100(.A (n_26598), .B (n_27227), .Y (n_28380));
NAND2X1 g107537(.A (n_6517), .B (n_26767), .Y (n_27700));
OAI21X1 g107539(.A0 (n_26068), .A1 (n_27698), .B0 (n_6750), .Y(n_27699));
OAI21X1 g110106(.A0 (n_26091), .A1 (n_27696), .B0 (n_26664), .Y(n_27697));
INVX1 g110107(.A (n_27215), .Y (n_27695));
INVX1 g110109(.A (n_27214), .Y (n_27694));
INVX1 g110119(.A (n_27691), .Y (n_28969));
INVX1 g110123(.A (n_27689), .Y (n_28966));
OAI21X1 g110126(.A0 (n_26073), .A1 (n_13214), .B0 (n_27687), .Y(n_28360));
OAI21X1 g110128(.A0 (n_26072), .A1 (n_13736), .B0 (n_27686), .Y(n_28358));
NAND2X1 g110149(.A (n_26581), .B (n_27685), .Y (n_28406));
INVX1 g110159(.A (n_27682), .Y (n_28182));
NAND2X1 g110163(.A (n_26610), .B (n_27681), .Y (n_28181));
NAND2X1 g110176(.A (n_26613), .B (n_26706), .Y (n_27680));
INVX1 g110179(.A (n_27198), .Y (n_27679));
INVX1 g110182(.A (n_27196), .Y (n_27678));
AOI21X1 g110184(.A0 (n_34712), .A1 (n_27676), .B0 (n_26734), .Y(n_27677));
AOI21X1 g110188(.A0 (n_26781), .A1 (n_28791), .B0 (n_26723), .Y(n_27675));
NAND2X1 g110189(.A (n_6685), .B (n_26761), .Y (n_27674));
OAI21X1 g110198(.A0 (n_27660), .A1 (n_33734), .B0 (n_20909), .Y(n_27673));
NAND2X1 g110203(.A (n_6674), .B (n_26760), .Y (n_27672));
OAI21X1 g110208(.A0 (n_20231), .A1 (n_25540), .B0 (n_26580), .Y(n_27671));
AOI21X1 g110210(.A0 (n_33546), .A1 (n_26392), .B0 (n_26740), .Y(n_32592));
AOI21X1 g110211(.A0 (n_33546), .A1 (n_27668), .B0 (n_26738), .Y(n_35133));
NAND2X1 g107581(.A (n_26481), .B (n_31590), .Y (n_27667));
AOI21X1 g110213(.A0 (n_34712), .A1 (n_27665), .B0 (n_26737), .Y(n_27666));
NAND2X1 g110216(.A (n_26733), .B (n_26353), .Y (n_27664));
OAI21X1 g110221(.A0 (n_26368), .A1 (n_27662), .B0 (n_26627), .Y(n_27663));
OAI21X1 g110223(.A0 (n_27660), .A1 (n_28523), .B0 (n_26274), .Y(n_27661));
AOI21X1 g110230(.A0 (n_27658), .A1 (n_28136), .B0 (n_20378), .Y(n_27659));
NAND2X2 g110238(.A (n_26277), .B (n_26628), .Y (n_28427));
NAND2X1 g110290(.A (n_33546), .B (n_27637), .Y (n_27657));
AOI21X1 g107626(.A0 (n_26061), .A1 (n_26105), .B0 (n_31041), .Y(n_27656));
NAND2X1 g110325(.A (n_29065), .B (n_27649), .Y (n_27655));
NAND2X1 g110331(.A (n_34770), .B (n_27647), .Y (n_27654));
NAND2X1 g110338(.A (n_34770), .B (n_27645), .Y (n_27653));
AND2X1 g110344(.A (n_27651), .B (n_28926), .Y (n_27652));
AND2X1 g110352(.A (n_27649), .B (n_34709), .Y (n_27650));
NAND2X1 g110359(.A (n_27647), .B (n_29925), .Y (n_27648));
NAND2X1 g110367(.A (n_27645), .B (n_34709), .Y (n_27646));
NAND2X1 g110378(.A (n_27651), .B (n_28013), .Y (n_27644));
NOR2X1 g110383(.A (n_24379), .B (n_26492), .Y (n_35136));
NOR2X1 g110384(.A (n_25622), .B (n_26491), .Y (n_35123));
NAND2X1 g110391(.A (n_27649), .B (n_28915), .Y (n_27641));
NAND2X1 g110397(.A (n_27647), .B (n_28013), .Y (n_27640));
NAND2X1 g110409(.A (n_27645), .B (n_29455), .Y (n_27639));
NAND2X1 g110526(.A (n_27637), .B (n_30559), .Y (n_27638));
NOR2X1 g107739(.A (n_26477), .B (n_15257), .Y (n_27636));
NAND2X1 g110579(.A (n_29430), .B (n_27634), .Y (n_27635));
NAND2X1 g110582(.A (n_27632), .B (n_27630), .Y (n_27633));
NAND2X1 g110583(.A (n_24925), .B (n_27630), .Y (n_27631));
INVX1 g110596(.A (n_27628), .Y (n_27629));
NAND2X1 g110626(.A (n_27625), .B (n_27462), .Y (n_27627));
NAND2X1 g110628(.A (n_27625), .B (n_27522), .Y (n_27626));
NAND2X1 g110633(.A (n_27621), .B (n_8990), .Y (n_27623));
NAND2X1 g110635(.A (n_27621), .B (n_29505), .Y (n_27622));
NAND2X1 g110658(.A (n_27619), .B (n_29505), .Y (n_27620));
NAND2X1 g110659(.A (n_27619), .B (n_26132), .Y (n_27618));
NAND2X1 g110694(.A (n_27100), .B (n_27613), .Y (n_27616));
NAND2X1 g110696(.A (n_27614), .B (n_27613), .Y (n_27615));
NAND2X1 g110741(.A (n_26077), .B (n_28364), .Y (n_27612));
NAND2X1 g110757(.A (n_27609), .B (n_33738), .Y (n_27611));
NAND2X1 g110787(.A (n_27609), .B (n_29405), .Y (n_27610));
NOR2X1 g110801(.A (n_24366), .B (n_26500), .Y (n_27608));
NOR2X1 g110802(.A (n_25613), .B (n_26499), .Y (n_27607));
NAND2X1 g110847(.A (n_26509), .B (n_29505), .Y (n_27606));
INVX1 g110863(.A (n_28254), .Y (n_28148));
NAND2X1 g110867(.A (n_26517), .B (n_27068), .Y (n_28146));
NAND2X1 g110872(.A (n_26516), .B (n_26569), .Y (n_28850));
NAND2X1 g110904(.A (n_26532), .B (n_27064), .Y (n_28809));
INVX1 g110905(.A (n_28276), .Y (n_27603));
NAND2X1 g110909(.A (n_26531), .B (n_26564), .Y (n_28140));
OAI21X1 g110928(.A0 (n_26062), .A1 (n_13843), .B0 (n_24675), .Y(n_28138));
INVX1 g110929(.A (n_28267), .Y (n_27600));
NAND2X1 g110931(.A (n_14128), .B (n_32121), .Y (n_28817));
NAND2X1 g110946(.A (n_26521), .B (n_27059), .Y (n_28813));
INVX1 g110947(.A (n_28260), .Y (n_27598));
NAND2X1 g110949(.A (n_26519), .B (n_26558), .Y (n_28826));
INVX1 g110987(.A (n_27055), .Y (n_27595));
OAI21X1 g110996(.A0 (n_25589), .A1 (n_8382), .B0 (n_20287), .Y(n_27594));
AOI21X1 g111005(.A0 (n_27584), .A1 (n_26213), .B0 (n_19713), .Y(n_27593));
NAND2X1 g111045(.A (n_26511), .B (n_29411), .Y (n_27592));
OAI21X1 g107949(.A0 (n_9767), .A1 (n_35012), .B0 (n_26482), .Y(n_27591));
NAND4X1 g107956(.A (n_21784), .B (n_24841), .C (n_21675), .D(n_26025), .Y (n_27590));
OAI21X1 g111076(.A0 (n_25591), .A1 (n_8285), .B0 (n_26542), .Y(n_27589));
OAI21X1 g111079(.A0 (n_24578), .A1 (n_8664), .B0 (n_26525), .Y(n_27588));
AOI21X1 g111080(.A0 (n_25268), .A1 (n_29619), .B0 (n_26523), .Y(n_27587));
NAND2X1 g111084(.A (n_26539), .B (n_26101), .Y (n_27586));
AOI21X1 g111085(.A0 (n_27584), .A1 (n_28791), .B0 (n_26148), .Y(n_27585));
AND2X1 g111128(.A (n_27579), .B (n_34952), .Y (n_27583));
NAND2X1 g111129(.A (n_27575), .B (n_26160), .Y (n_27582));
AND2X1 g111139(.A (n_27577), .B (n_34952), .Y (n_27581));
AND2X1 g111148(.A (n_27579), .B (n_34693), .Y (n_27580));
NAND2X1 g111157(.A (n_27577), .B (n_27340), .Y (n_27578));
AND2X1 g111160(.A (n_27575), .B (n_34693), .Y (n_27576));
NAND2X1 g111172(.A (n_27579), .B (n_28808), .Y (n_27573));
NAND2X1 g111189(.A (n_27577), .B (n_26535), .Y (n_27572));
NAND2X1 g111196(.A (n_27575), .B (n_26142), .Y (n_27571));
NOR2X1 g108022(.A (n_6774), .B (n_26503), .Y (n_27570));
NAND4X1 g108024(.A (n_14428), .B (n_24124), .C (n_25747), .D(n_24763), .Y (n_27569));
NAND2X1 g108025(.A (n_26502), .B (n_27567), .Y (n_27568));
NOR2X1 g111286(.A (n_27565), .B (n_27564), .Y (n_27566));
OAI21X1 g111370(.A0 (n_27549), .A1 (n_27042), .B0 (n_29505), .Y(n_27563));
NOR2X1 g108083(.A (n_13742), .B (n_26494), .Y (n_27562));
NOR2X1 g108084(.A (n_14173), .B (n_26490), .Y (n_27561));
NOR2X1 g108086(.A (n_14157), .B (n_26485), .Y (n_27560));
NAND2X1 g108141(.A (n_26447), .B (n_31097), .Y (n_27559));
OAI21X1 g108160(.A0 (n_26425), .A1 (n_27557), .B0 (n_10364), .Y(n_27558));
OAI21X1 g108161(.A0 (n_26424), .A1 (n_27557), .B0 (n_10426), .Y(n_27556));
NAND3X1 g108166(.A (n_26742), .B (n_25221), .C (n_15289), .Y(n_27555));
NAND4X1 g108221(.A (n_15009), .B (n_25467), .C (n_25899), .D(n_25478), .Y (n_27554));
INVX1 g111700(.A (n_28159), .Y (n_27553));
NOR2X1 g108222(.A (n_26433), .B (n_14661), .Y (n_27551));
MX2X1 g111783(.A (n_18227), .B (n_18218), .S0 (n_27549), .Y(n_27550));
AOI21X1 g111784(.A0 (n_27021), .A1 (n_8037), .B0 (n_26483), .Y(n_27548));
NAND2X1 g108316(.A (n_27521), .B (n_27537), .Y (n_28726));
NAND2X1 g108317(.A (n_14944), .B (n_27539), .Y (n_27547));
NAND2X1 g108318(.A (n_32869), .B (n_17968), .Y (n_28709));
NAND2X1 g108327(.A (n_13904), .B (n_27542), .Y (n_28721));
NAND4X1 g108330(.A (n_26808), .B (n_19852), .C (n_9529), .D (n_9021),.Y (n_27545));
NAND2X1 g108338(.A (n_27544), .B (n_27519), .Y (n_28696));
AND2X1 g108339(.A (n_27542), .B (n_14936), .Y (n_27543));
NAND2X1 g108342(.A (n_32870), .B (n_35736), .Y (n_27541));
NAND2X1 g108355(.A (n_27539), .B (n_27525), .Y (n_28715));
NAND2X1 g108356(.A (n_27537), .B (n_14930), .Y (n_27538));
NAND4X1 g108392(.A (n_15007), .B (n_25484), .C (n_25913), .D(n_25482), .Y (n_27536));
NAND2X1 g108403(.A (n_32870), .B (n_35500), .Y (n_28711));
OAI21X1 g108414(.A0 (n_15129), .A1 (n_28659), .B0 (n_26464), .Y(n_27535));
NAND2X1 g108420(.A (n_26443), .B (n_31097), .Y (n_27534));
NAND2X1 g108432(.A (n_26441), .B (n_31345), .Y (n_27533));
OAI21X1 g108433(.A0 (n_15127), .A1 (n_26801), .B0 (n_26463), .Y(n_27532));
AOI21X1 g108451(.A0 (n_26402), .A1 (n_7967), .B0 (n_8614), .Y(n_27531));
OAI21X1 g108455(.A0 (n_15123), .A1 (n_28659), .B0 (n_26459), .Y(n_27530));
AOI21X1 g108459(.A0 (n_27100), .A1 (n_26958), .B0 (n_26438), .Y(n_27529));
OAI21X1 g108463(.A0 (n_9849), .A1 (n_28332), .B0 (n_26473), .Y(n_27528));
INVX1 g112360(.A (n_27527), .Y (n_28681));
NOR2X1 g108531(.A (n_7090), .B (n_26476), .Y (n_27526));
NAND2X2 g108582(.A (n_26444), .B (n_27525), .Y (n_28738));
AOI21X1 g108597(.A0 (n_27523), .A1 (n_27522), .B0 (n_20874), .Y(n_27524));
OAI21X1 g108628(.A0 (n_26359), .A1 (n_13214), .B0 (n_27521), .Y(n_28704));
INVX1 g108636(.A (n_28155), .Y (n_27520));
NAND2X1 g108643(.A (n_26450), .B (n_27519), .Y (n_28052));
INVX1 g106940(.A (n_26989), .Y (n_27518));
OAI21X1 g108654(.A0 (n_15120), .A1 (n_28659), .B0 (n_26460), .Y(n_27517));
NAND2X1 g108685(.A (n_6704), .B (n_26466), .Y (n_27516));
NAND2X1 g108686(.A (n_6550), .B (n_26465), .Y (n_27515));
INVX1 g106957(.A (n_26986), .Y (n_27514));
NAND4X1 g108730(.A (n_26395), .B (n_10232), .C (n_25640), .D(n_25627), .Y (n_27513));
NOR2X1 g108735(.A (n_19125), .B (n_26790), .Y (n_27512));
NAND2X1 g106980(.A (n_26825), .B (n_25942), .Y (n_27511));
NOR2X1 g108741(.A (n_26786), .B (n_26789), .Y (n_27510));
NAND3X1 g108748(.A (n_20217), .B (n_26294), .C (n_25979), .Y(n_27509));
NAND2X1 g106988(.A (n_26797), .B (n_8641), .Y (n_27508));
NAND3X1 g108767(.A (n_10868), .B (n_25983), .C (n_26318), .Y(n_27507));
NOR2X1 g108775(.A (n_11147), .B (n_26772), .Y (n_27506));
NAND3X1 g108797(.A (n_26745), .B (n_24472), .C (n_14968), .Y(n_27505));
NAND2X1 g108810(.A (n_34770), .B (n_27500), .Y (n_27504));
NAND2X1 g108816(.A (n_34770), .B (n_27498), .Y (n_27503));
NAND2X1 g108836(.A (n_27500), .B (n_34709), .Y (n_27501));
NAND2X1 g108843(.A (n_27498), .B (n_34709), .Y (n_27499));
NAND2X1 g108858(.A (n_27495), .B (n_25980), .Y (n_27496));
NAND2X1 g108871(.A (n_27493), .B (n_28013), .Y (n_27494));
NAND2X1 g108879(.A (n_27500), .B (n_29455), .Y (n_27492));
NAND2X1 g108887(.A (n_27498), .B (n_29455), .Y (n_27491));
NAND2X1 g108890(.A (n_35688), .B (n_8954), .Y (n_27490));
NAND2X1 g108909(.A (n_27483), .B (n_27999), .Y (n_27488));
NAND2X1 g108912(.A (n_27479), .B (n_26530), .Y (n_27487));
OAI21X1 g108915(.A0 (n_26358), .A1 (n_26317), .B0 (n_27485), .Y(n_27486));
NAND2X1 g108936(.A (n_27483), .B (n_22406), .Y (n_27484));
NAND2X1 g108937(.A (n_27467), .B (n_21919), .Y (n_27481));
NAND2X1 g108938(.A (n_27479), .B (n_22064), .Y (n_27480));
NAND2X1 g108955(.A (n_27483), .B (n_32685), .Y (n_27478));
NAND2X1 g108958(.A (n_27479), .B (n_32739), .Y (n_27477));
NOR2X1 g108973(.A (n_27475), .B (n_8382), .Y (n_27476));
NOR2X1 g108974(.A (n_27475), .B (n_8678), .Y (n_27473));
AND2X1 g108980(.A (n_27229), .B (n_27956), .Y (n_27472));
NAND2X1 g108986(.A (n_27483), .B (n_27470), .Y (n_27471));
NAND2X1 g108988(.A (n_27479), .B (n_25290), .Y (n_27469));
NAND2X1 g108989(.A (n_24361), .B (n_27467), .Y (n_27468));
NAND4X1 g108996(.A (n_26350), .B (n_25173), .C (n_24792), .D(n_25821), .Y (n_27466));
NAND2X1 g109018(.A (n_27467), .B (n_23578), .Y (n_27465));
NAND3X1 g109021(.A (n_26022), .B (n_26242), .C (n_20434), .Y(n_27464));
NAND2X1 g109029(.A (n_27462), .B (n_27461), .Y (n_27463));
NAND2X1 g109034(.A (n_27462), .B (n_27459), .Y (n_27460));
NAND2X1 g109036(.A (n_26853), .B (n_18335), .Y (n_32058));
NAND2X1 g109050(.A (n_33644), .B (n_18546), .Y (n_28603));
NAND2X1 g109051(.A (n_35649), .B (n_18546), .Y (n_28615));
NAND2X1 g109055(.A (n_26850), .B (n_18349), .Y (n_32918));
NAND2X1 g109057(.A (n_33917), .B (n_27451), .Y (n_27453));
NAND3X1 g109059(.A (n_25465), .B (n_26177), .C (n_15245), .Y(n_27450));
NAND3X1 g109061(.A (n_26386), .B (n_26240), .C (n_20892), .Y(n_27449));
NAND2X1 g109062(.A (n_27445), .B (n_27462), .Y (n_27448));
NAND2X1 g109063(.A (n_27420), .B (n_33738), .Y (n_27447));
NAND2X1 g109064(.A (n_27445), .B (n_27522), .Y (n_27446));
NAND2X1 g109066(.A (n_24925), .B (n_27441), .Y (n_27444));
NAND2X1 g109067(.A (n_27441), .B (n_29505), .Y (n_27442));
AND2X1 g109068(.A (n_27441), .B (n_30291), .Y (n_27440));
NAND2X1 g109083(.A (n_33648), .B (n_35816), .Y (n_28610));
NOR2X1 g109086(.A (n_26815), .B (n_25463), .Y (n_27438));
NAND2X1 g109094(.A (n_27436), .B (n_29505), .Y (n_27437));
NAND2X1 g109095(.A (n_27436), .B (n_26132), .Y (n_27435));
NAND2X1 g109098(.A (n_27203), .B (n_28874), .Y (n_27434));
NAND2X1 g109107(.A (n_33644), .B (n_35744), .Y (n_27433));
NAND2X1 g109108(.A (n_35650), .B (n_35822), .Y (n_27431));
NAND2X1 g109123(.A (n_35689), .B (n_28158), .Y (n_27430));
NAND2X1 g109124(.A (n_30454), .B (n_27264), .Y (n_27429));
NAND2X1 g109125(.A (n_33991), .B (n_35689), .Y (n_27428));
NOR2X1 g109126(.A (n_26382), .B (n_26824), .Y (n_27427));
NAND2X1 g109130(.A (n_8989), .B (n_27424), .Y (n_27426));
NAND2X1 g109132(.A (n_24925), .B (n_27424), .Y (n_27425));
NAND2X1 g109155(.A (n_27467), .B (n_27422), .Y (n_27423));
NAND2X1 g109159(.A (n_27420), .B (n_28158), .Y (n_27421));
NAND2X1 g109160(.A (n_27420), .B (n_28374), .Y (n_27419));
NOR2X1 g109175(.A (n_26814), .B (n_25859), .Y (n_27418));
NAND4X1 g109181(.A (n_26889), .B (n_23781), .C (n_24588), .D(n_24615), .Y (n_27417));
NAND2X1 g109206(.A (n_27414), .B (n_26238), .Y (n_27416));
NAND2X1 g109217(.A (n_27414), .B (n_33738), .Y (n_27415));
NAND2X1 g109218(.A (n_33644), .B (n_35479), .Y (n_28605));
NAND2X1 g109219(.A (n_35650), .B (n_35473), .Y (n_28612));
NAND2X1 g109222(.A (n_32844), .B (n_25877), .Y (n_28608));
NAND2X1 g109224(.A (n_27414), .B (n_29405), .Y (n_27410));
NOR2X1 g109235(.A (n_10228), .B (n_26773), .Y (n_27409));
NAND3X1 g109240(.A (n_9589), .B (n_26334), .C (n_26314), .Y(n_27408));
NAND3X1 g109241(.A (n_26313), .B (n_20294), .C (n_26311), .Y(n_27407));
OAI21X1 g109257(.A0 (n_26195), .A1 (n_29388), .B0 (n_21362), .Y(n_27406));
NAND3X1 g109262(.A (n_25855), .B (n_26225), .C (n_19910), .Y(n_27405));
NAND3X1 g109285(.A (n_9055), .B (n_26264), .C (n_20888), .Y(n_27404));
NOR2X1 g109289(.A (n_10155), .B (n_26771), .Y (n_27403));
NAND2X1 g109291(.A (n_26838), .B (n_26783), .Y (n_27402));
OAI21X1 g109294(.A0 (n_26194), .A1 (n_33807), .B0 (n_21338), .Y(n_27401));
NOR2X1 g109301(.A (n_26829), .B (n_26792), .Y (n_27400));
NAND2X1 g109307(.A (n_26865), .B (n_27399), .Y (n_27861));
NOR2X1 g109316(.A (n_26355), .B (n_26891), .Y (n_27397));
NOR2X1 g109317(.A (n_26327), .B (n_26890), .Y (n_27396));
AOI21X1 g109330(.A0 (n_27338), .A1 (n_26162), .B0 (n_15037), .Y(n_27395));
AOI21X1 g109333(.A0 (n_27336), .A1 (n_26162), .B0 (n_15160), .Y(n_32070));
AOI21X1 g109334(.A0 (n_27333), .A1 (n_26162), .B0 (n_15193), .Y(n_32080));
OAI21X1 g109339(.A0 (n_14953), .A1 (n_8949), .B0 (n_26828), .Y(n_27391));
AOI21X1 g109340(.A0 (n_27341), .A1 (n_26162), .B0 (n_15146), .Y(n_27390));
NAND2X1 g109344(.A (n_26888), .B (n_27389), .Y (n_28653));
NAND2X2 g109348(.A (n_26887), .B (n_27388), .Y (n_28642));
INVX1 g109351(.A (n_27386), .Y (n_27387));
NAND2X1 g109356(.A (n_35260), .B (n_27384), .Y (n_28651));
NAND2X2 g109360(.A (n_26880), .B (n_14126), .Y (n_28741));
INVX1 g109363(.A (n_27382), .Y (n_27383));
NAND2X1 g109370(.A (n_26876), .B (n_27380), .Y (n_28655));
NAND2X1 g109374(.A (n_26875), .B (n_27379), .Y (n_27849));
INVX1 g109375(.A (n_27378), .Y (n_29122));
NAND2X1 g109384(.A (n_26867), .B (n_27377), .Y (n_28647));
AND2X1 g109389(.A (n_26844), .B (n_20852), .Y (n_27376));
OAI21X1 g109399(.A0 (n_26172), .A1 (n_10517), .B0 (n_20879), .Y(n_27375));
AOI21X1 g109401(.A0 (n_27275), .A1 (n_14634), .B0 (n_26920), .Y(n_27374));
AOI22X1 g109410(.A0 (n_27313), .A1 (n_26213), .B0 (n_9629), .B1(n_19541), .Y (n_27373));
AOI22X1 g109411(.A0 (n_27304), .A1 (n_26213), .B0 (n_9629), .B1(n_19539), .Y (n_27372));
AOI22X1 g109414(.A0 (n_27297), .A1 (n_26213), .B0 (n_9629), .B1(n_19536), .Y (n_27370));
AOI22X1 g109416(.A0 (n_27290), .A1 (n_26213), .B0 (n_9629), .B1(n_19533), .Y (n_27369));
NAND2X1 g109418(.A (n_26809), .B (n_15069), .Y (n_27368));
NAND2X1 g109419(.A (n_26805), .B (n_15097), .Y (n_27367));
NOR2X1 g109424(.A (n_25879), .B (n_26766), .Y (n_27366));
NAND2X1 g109425(.A (n_26813), .B (n_15251), .Y (n_27365));
NAND2X1 g109426(.A (n_26811), .B (n_15275), .Y (n_27364));
NAND2X1 g109428(.A (n_26839), .B (n_19853), .Y (n_27363));
NAND2X1 g109435(.A (n_26840), .B (n_26548), .Y (n_27362));
AOI21X1 g109436(.A0 (n_14632), .A1 (n_27306), .B0 (n_29725), .Y(n_27361));
NAND3X1 g109448(.A (n_25891), .B (n_26349), .C (n_25889), .Y(n_27360));
NAND4X1 g109451(.A (n_25145), .B (n_10619), .C (n_25784), .D(n_25132), .Y (n_27359));
AOI21X1 g109463(.A0 (n_8922), .A1 (n_26857), .B0 (n_21348), .Y(n_27358));
AOI21X1 g109467(.A0 (n_33546), .A1 (n_26938), .B0 (n_26341), .Y(n_27357));
AOI21X1 g109476(.A0 (n_33546), .A1 (n_26940), .B0 (n_26344), .Y(n_27356));
OAI21X1 g109488(.A0 (n_26416), .A1 (n_26415), .B0 (n_26417), .Y(n_28091));
NOR2X1 g109497(.A (n_25999), .B (n_26097), .Y (n_27355));
NOR2X1 g109506(.A (n_19525), .B (n_26215), .Y (n_32082));
NOR2X1 g109519(.A (n_10590), .B (n_26167), .Y (n_27353));
AOI21X1 g109524(.A0 (n_25724), .A1 (n_24877), .B0 (n_8340), .Y(n_27352));
AOI21X1 g109529(.A0 (n_25709), .A1 (n_24848), .B0 (n_8340), .Y(n_27351));
NAND4X1 g109532(.A (n_26141), .B (n_18730), .C (n_22820), .D(n_24287), .Y (n_27350));
AOI21X1 g109533(.A0 (n_29068), .A1 (n_26739), .B0 (n_24432), .Y(n_32593));
NOR2X1 g109539(.A (n_26347), .B (n_25346), .Y (n_27348));
OAI21X1 g109540(.A0 (n_25703), .A1 (n_9626), .B0 (n_23786), .Y(n_27347));
NAND2X1 g109546(.A (n_27331), .B (n_34952), .Y (n_27346));
NAND2X1 g109547(.A (n_27322), .B (n_28864), .Y (n_27345));
NAND2X1 g109551(.A (n_27329), .B (n_26160), .Y (n_32104));
NAND2X1 g109552(.A (n_27319), .B (n_26162), .Y (n_27343));
NAND2X1 g109555(.A (n_27341), .B (n_27340), .Y (n_27342));
NAND2X1 g109556(.A (n_27338), .B (n_27335), .Y (n_27339));
NAND2X1 g109560(.A (n_27336), .B (n_27335), .Y (n_27337));
NAND2X1 g109561(.A (n_27333), .B (n_27335), .Y (n_27334));
NAND2X1 g109565(.A (n_27331), .B (n_28485), .Y (n_27332));
NAND2X1 g109570(.A (n_27329), .B (n_27340), .Y (n_27330));
NAND2X1 g109575(.A (n_27338), .B (n_29090), .Y (n_27328));
NAND2X1 g109579(.A (n_27336), .B (n_27326), .Y (n_27327));
NAND2X1 g109580(.A (n_27333), .B (n_27326), .Y (n_27325));
NAND2X1 g109584(.A (n_27331), .B (n_33378), .Y (n_27324));
NAND2X1 g109585(.A (n_27322), .B (n_29090), .Y (n_27323));
NAND2X1 g109588(.A (n_27329), .B (n_28468), .Y (n_27321));
NAND2X1 g109589(.A (n_27319), .B (n_27326), .Y (n_27320));
NOR2X1 g109592(.A (n_27256), .B (n_26175), .Y (n_27318));
NAND2X1 g109593(.A (n_27341), .B (n_27326), .Y (n_27317));
NOR2X1 g109595(.A (n_26212), .B (n_14604), .Y (n_27316));
NOR2X1 g109603(.A (n_26176), .B (n_14625), .Y (n_27315));
NAND2X1 g109611(.A (n_27313), .B (n_28785), .Y (n_35096));
NAND2X1 g109612(.A (n_27313), .B (n_34753), .Y (n_27311));
NAND2X1 g109613(.A (n_27313), .B (n_30369), .Y (n_27310));
NOR2X1 g109614(.A (n_24276), .B (n_26224), .Y (n_27309));
NAND2X1 g109624(.A (n_27300), .B (n_23725), .Y (n_27308));
NAND3X1 g109641(.A (n_26190), .B (n_25143), .C (n_25801), .Y(n_27307));
NAND2X1 g109648(.A (n_27306), .B (n_27204), .Y (n_27886));
NAND2X1 g109653(.A (n_27304), .B (n_28785), .Y (n_35634));
NAND2X1 g109654(.A (n_27304), .B (n_34753), .Y (n_27303));
NAND2X1 g109655(.A (n_27304), .B (n_30369), .Y (n_27302));
NAND2X1 g109662(.A (n_27300), .B (n_18384), .Y (n_27301));
NOR2X1 g109671(.A (n_24270), .B (n_26304), .Y (n_27299));
NAND2X1 g109681(.A (n_27297), .B (n_28785), .Y (n_27298));
NAND2X1 g109682(.A (n_27297), .B (n_34753), .Y (n_27296));
NAND2X1 g109683(.A (n_27297), .B (n_30369), .Y (n_27295));
NAND2X1 g109688(.A (n_27300), .B (n_32664), .Y (n_27294));
NAND3X1 g109701(.A (n_26214), .B (n_25141), .C (n_25765), .Y(n_27292));
NAND2X1 g109707(.A (n_27290), .B (n_26528), .Y (n_32276));
NAND2X1 g109709(.A (n_27290), .B (n_28636), .Y (n_27289));
NAND2X1 g109710(.A (n_27290), .B (n_30063), .Y (n_27288));
NAND3X1 g107385(.A (n_22170), .B (n_23876), .C (n_25594), .Y(n_28666));
NAND2X1 g109723(.A (n_27300), .B (n_34688), .Y (n_27287));
NOR2X1 g109731(.A (n_24266), .B (n_26280), .Y (n_27286));
NAND2X1 g109743(.A (n_27632), .B (n_27283), .Y (n_27285));
NAND2X1 g109744(.A (n_24925), .B (n_27283), .Y (n_27284));
NAND2X1 g109756(.A (n_27207), .B (n_27260), .Y (n_27945));
NAND2X1 g109757(.A (n_14887), .B (n_27262), .Y (n_27282));
NOR2X1 g109762(.A (n_24264), .B (n_26220), .Y (n_27281));
NAND2X1 g109768(.A (n_26582), .B (n_27205), .Y (n_27907));
NAND2X1 g109770(.A (n_27277), .B (n_29505), .Y (n_27280));
NAND2X1 g109772(.A (n_27277), .B (n_8990), .Y (n_27278));
NAND2X1 g109779(.A (n_26371), .B (n_27275), .Y (n_27905));
NAND2X1 g109780(.A (n_14721), .B (n_27271), .Y (n_27274));
NAND2X1 g109781(.A (n_26776), .B (n_27269), .Y (n_27941));
NAND2X1 g109786(.A (n_14680), .B (n_33730), .Y (n_27273));
NAND3X1 g109790(.A (n_26170), .B (n_25382), .C (n_24710), .Y(n_27272));
NAND2X1 g109801(.A (n_27271), .B (n_26774), .Y (n_27883));
NAND2X1 g109802(.A (n_27269), .B (n_14266), .Y (n_27270));
NAND3X1 g109813(.A (n_26184), .B (n_25139), .C (n_25786), .Y(n_27267));
NOR2X1 g109817(.A (n_25748), .B (n_26578), .Y (n_27266));
INVX1 g109820(.A (n_27264), .Y (n_27265));
NOR2X1 g109825(.A (n_26270), .B (n_13521), .Y (n_27263));
NAND2X1 g109827(.A (n_27225), .B (n_27262), .Y (n_27912));
NAND2X1 g109828(.A (n_27260), .B (n_14437), .Y (n_27261));
NAND2X1 g109832(.A (n_26351), .B (n_24729), .Y (n_27259));
NOR2X1 g109845(.A (n_26164), .B (n_24098), .Y (n_27258));
NOR2X1 g109856(.A (n_27256), .B (n_26178), .Y (n_27257));
NOR2X1 g109866(.A (n_27256), .B (n_26287), .Y (n_27255));
AOI21X1 g109883(.A0 (n_27253), .A1 (n_30557), .B0 (n_21375), .Y(n_27254));
NOR2X1 g109885(.A (n_9123), .B (n_26169), .Y (n_27252));
NOR2X1 g109897(.A (n_9085), .B (n_26168), .Y (n_27251));
NAND3X1 g109900(.A (n_25779), .B (n_20792), .C (n_25778), .Y(n_27250));
OAI21X1 g109906(.A0 (n_25692), .A1 (n_33807), .B0 (n_21369), .Y(n_27249));
AOI21X1 g109907(.A0 (n_27247), .A1 (n_29040), .B0 (n_21368), .Y(n_27248));
OAI21X1 g109909(.A0 (n_25691), .A1 (n_29388), .B0 (n_19918), .Y(n_27246));
NAND3X1 g109911(.A (n_25759), .B (n_20790), .C (n_25758), .Y(n_27245));
NAND4X1 g109915(.A (n_26099), .B (n_18720), .C (n_22812), .D(n_24286), .Y (n_27244));
AOI21X1 g109923(.A0 (n_24925), .A1 (n_26626), .B0 (n_26222), .Y(n_27243));
OAI21X1 g109931(.A0 (n_9856), .A1 (n_31299), .B0 (n_26352), .Y(n_27241));
NOR2X1 g109933(.A (n_9559), .B (n_26174), .Y (n_27240));
NOR2X1 g109937(.A (n_9074), .B (n_26171), .Y (n_27239));
AOI21X1 g109939(.A0 (n_27100), .A1 (n_26615), .B0 (n_25161), .Y(n_27238));
AOI21X1 g109942(.A0 (n_27100), .A1 (n_26257), .B0 (n_26192), .Y(n_27237));
AOI21X1 g109944(.A0 (n_27235), .A1 (n_27234), .B0 (n_19847), .Y(n_27236));
AOI22X1 g109951(.A0 (n_25707), .A1 (n_27232), .B0 (n_1153), .B1(n_12926), .Y (n_27233));
NAND2X1 g109959(.A (n_26291), .B (n_26791), .Y (n_27974));
INVX1 g109960(.A (n_27493), .Y (n_27231));
NAND2X1 g109969(.A (n_26285), .B (n_27230), .Y (n_27725));
INVX1 g109976(.A (n_27229), .Y (n_27967));
NAND2X1 g109978(.A (n_26284), .B (n_13174), .Y (n_28593));
NAND2X1 g109994(.A (n_26324), .B (n_13667), .Y (n_28003));
NAND2X1 g109995(.A (n_26246), .B (n_27227), .Y (n_28018));
NAND2X1 g109998(.A (n_26323), .B (n_24190), .Y (n_28971));
NAND2X1 g110000(.A (n_26230), .B (n_26398), .Y (n_27920));
NAND2X1 g110001(.A (n_26316), .B (n_24508), .Y (n_27995));
INVX1 g110002(.A (n_27495), .Y (n_27226));
NAND2X2 g110012(.A (n_26227), .B (n_27225), .Y (n_28020));
NAND2X1 g110018(.A (n_26309), .B (n_13650), .Y (n_27990));
NAND2X2 g110026(.A (n_26307), .B (n_27222), .Y (n_29392));
NAND2X1 g110029(.A (n_26305), .B (n_27221), .Y (n_28025));
NAND2X1 g110032(.A (n_26300), .B (n_27220), .Y (n_28034));
NAND2X1 g110035(.A (n_26299), .B (n_27219), .Y (n_27714));
OAI21X1 g110055(.A0 (n_25664), .A1 (n_13273), .B0 (n_26787), .Y(n_27957));
NAND2X1 g110067(.A (n_26278), .B (n_27217), .Y (n_28023));
NAND2X1 g110077(.A (n_26262), .B (n_20882), .Y (n_27216));
OAI21X1 g110081(.A0 (n_25664), .A1 (n_13781), .B0 (n_24505), .Y(n_27926));
NAND2X2 g110090(.A (n_26229), .B (n_26869), .Y (n_27916));
OAI21X1 g110108(.A0 (n_25347), .A1 (n_27696), .B0 (n_26296), .Y(n_27215));
OAI21X1 g110110(.A0 (n_25687), .A1 (n_8319), .B0 (n_26289), .Y(n_27214));
OAI21X1 g110111(.A0 (n_25701), .A1 (n_8382), .B0 (n_20285), .Y(n_27212));
OAI21X1 g110112(.A0 (n_26657), .A1 (n_8382), .B0 (n_20281), .Y(n_27211));
INVX1 g110115(.A (n_27208), .Y (n_28524));
NAND2X1 g110121(.A (n_26272), .B (n_26401), .Y (n_27691));
NAND2X1 g110125(.A (n_26268), .B (n_26854), .Y (n_27689));
OAI21X1 g110127(.A0 (n_25661), .A1 (n_13214), .B0 (n_27207), .Y(n_27895));
INVX1 g110142(.A (n_27445), .Y (n_27206));
NAND2X1 g110147(.A (n_26235), .B (n_27205), .Y (n_27938));
NAND2X1 g110151(.A (n_26254), .B (n_27204), .Y (n_27933));
INVX1 g110153(.A (n_27203), .Y (n_27683));
NAND2X1 g110160(.A (n_26253), .B (n_33731), .Y (n_27682));
NAND2X1 g110169(.A (n_26332), .B (n_26302), .Y (n_27201));
NAND2X1 g110173(.A (n_26281), .B (n_25978), .Y (n_27200));
NAND2X1 g110178(.A (n_26325), .B (n_26248), .Y (n_27199));
OAI21X1 g110180(.A0 (n_25352), .A1 (n_27696), .B0 (n_26319), .Y(n_27198));
NAND2X1 g110181(.A (n_26342), .B (n_26310), .Y (n_27197));
OAI21X1 g110183(.A0 (n_25699), .A1 (n_8319), .B0 (n_26303), .Y(n_27196));
AOI21X1 g107568(.A0 (n_10476), .A1 (n_25565), .B0 (n_31586), .Y(n_27195));
OAI21X1 g110197(.A0 (n_27193), .A1 (n_27192), .B0 (n_20877), .Y(n_27194));
NAND2X1 g110204(.A (n_6482), .B (n_26356), .Y (n_27190));
NAND2X1 g110207(.A (n_26231), .B (n_20863), .Y (n_27189));
NAND2X2 g110233(.A (n_25974), .B (n_26322), .Y (n_27986));
NAND2X2 g110240(.A (n_32307), .B (n_32308), .Y (n_27961));
NAND2X2 g110243(.A (n_26271), .B (n_25937), .Y (n_27983));
OAI21X1 g107608(.A0 (n_25577), .A1 (n_25811), .B0 (n_31628), .Y(n_27186));
NAND3X1 g110274(.A (n_20749), .B (n_25633), .C (n_24364), .Y(n_27185));
NAND3X1 g110277(.A (n_18023), .B (n_25611), .C (n_25631), .Y(n_27184));
NAND3X1 g110284(.A (n_10882), .B (n_25638), .C (n_24377), .Y(n_27183));
NAND3X1 g110285(.A (n_10879), .B (n_25620), .C (n_25635), .Y(n_27182));
NAND2X1 g110293(.A (n_34712), .B (n_27116), .Y (n_27181));
NAND2X1 g110297(.A (n_33546), .B (n_27105), .Y (n_27180));
NAND2X1 g110299(.A (n_34712), .B (n_27094), .Y (n_27179));
NOR2X1 g110306(.A (n_8677), .B (n_26126), .Y (n_27178));
NAND3X1 g110311(.A (n_26165), .B (n_23772), .C (n_15255), .Y(n_27177));
OAI21X1 g110313(.A0 (n_25587), .A1 (n_9626), .B0 (n_24093), .Y(n_27176));
NOR2X1 g110314(.A (n_26159), .B (n_24426), .Y (n_27175));
NOR2X1 g110316(.A (n_9172), .B (n_26096), .Y (n_27174));
NOR2X1 g110317(.A (n_9172), .B (n_26095), .Y (n_27172));
NOR2X1 g110321(.A (n_27169), .B (n_26091), .Y (n_27171));
NOR2X1 g110326(.A (n_27169), .B (n_26090), .Y (n_27170));
NOR2X1 g110334(.A (n_34771), .B (n_26084), .Y (n_27168));
NOR2X1 g110335(.A (n_9172), .B (n_26083), .Y (n_27167));
NOR2X1 g110339(.A (n_9172), .B (n_26087), .Y (n_27166));
NAND2X1 g110347(.A (n_27153), .B (n_34694), .Y (n_27164));
NAND2X1 g110348(.A (n_27162), .B (n_29008), .Y (n_27163));
NAND2X1 g110355(.A (n_34801), .B (n_27340), .Y (n_27161));
NOR2X1 g110363(.A (n_26084), .B (n_27158), .Y (n_27159));
NOR2X1 g110364(.A (n_26083), .B (n_27158), .Y (n_27157));
NAND2X1 g110370(.A (n_27149), .B (n_34694), .Y (n_32117));
NAND3X1 g110372(.A (n_24389), .B (n_25649), .C (n_24413), .Y(n_27155));
NAND2X1 g110381(.A (n_27743), .B (n_27153), .Y (n_27154));
NAND3X1 g110402(.A (n_24353), .B (n_25646), .C (n_24410), .Y(n_27152));
NAND3X1 g110403(.A (n_25607), .B (n_25644), .C (n_25657), .Y(n_27151));
NAND2X1 g110415(.A (n_27743), .B (n_27149), .Y (n_27150));
NAND2X1 g110436(.A (n_27668), .B (n_30668), .Y (n_27148));
NAND2X1 g110444(.A (n_27665), .B (n_29191), .Y (n_27147));
NAND2X1 g110447(.A (n_25554), .B (n_27130), .Y (n_27146));
NAND2X1 g110453(.A (n_27127), .B (n_25554), .Y (n_27144));
NAND2X1 g110454(.A (n_27125), .B (n_28441), .Y (n_27143));
NAND2X1 g110458(.A (n_27153), .B (n_34802), .Y (n_27142));
NAND2X1 g110460(.A (n_35040), .B (n_25302), .Y (n_27141));
AOI21X1 g110480(.A0 (n_9629), .A1 (n_17296), .B0 (n_26144), .Y(n_27140));
NAND4X1 g107708(.A (n_14879), .B (n_24133), .C (n_25406), .D(n_24774), .Y (n_27139));
NAND2X1 g110488(.A (n_27162), .B (n_34802), .Y (n_27138));
NOR2X1 g107716(.A (n_26423), .B (n_26070), .Y (n_27136));
NAND4X1 g107717(.A (n_14990), .B (n_14532), .C (n_27134), .D(n_25536), .Y (n_27135));
NAND2X1 g110508(.A (n_27676), .B (n_30184), .Y (n_27133));
NAND2X1 g110514(.A (n_25688), .B (n_10808), .Y (n_27132));
NAND2X1 g110515(.A (n_27130), .B (n_27770), .Y (n_27131));
NAND2X1 g110519(.A (n_27127), .B (n_25956), .Y (n_27128));
NAND2X1 g110520(.A (n_27125), .B (n_24361), .Y (n_27126));
NAND2X1 g110527(.A (n_35040), .B (n_23192), .Y (n_27122));
NAND4X1 g107730(.A (n_14776), .B (n_14771), .C (n_27118), .D(n_25535), .Y (n_27119));
NAND2X1 g110550(.A (n_27116), .B (n_30559), .Y (n_27117));
NAND2X1 g110553(.A (n_27130), .B (n_18137), .Y (n_27115));
NAND2X1 g110555(.A (n_27127), .B (n_13274), .Y (n_27114));
NAND2X1 g110557(.A (n_27125), .B (n_26637), .Y (n_27112));
NAND4X1 g107738(.A (n_15419), .B (n_15131), .C (n_15258), .D(n_25534), .Y (n_27111));
NAND2X1 g110559(.A (n_27099), .B (n_27109), .Y (n_27110));
NAND2X1 g110560(.A (n_35040), .B (n_23578), .Y (n_27108));
NAND2X1 g110577(.A (n_27105), .B (n_26660), .Y (n_27106));
NAND2X1 g110597(.A (n_35233), .B (n_18546), .Y (n_27628));
INVX1 g110600(.A (n_27102), .Y (n_27103));
NAND2X1 g110664(.A (n_27100), .B (n_27099), .Y (n_27101));
NAND2X1 g110666(.A (n_27099), .B (n_27632), .Y (n_27098));
NAND2X1 g110671(.A (n_35233), .B (n_35744), .Y (n_27097));
NAND2X1 g110675(.A (n_27094), .B (n_29191), .Y (n_27095));
NAND2X1 g110681(.A (n_27130), .B (n_25605), .Y (n_27093));
NAND2X1 g110689(.A (n_27127), .B (n_27091), .Y (n_27092));
NAND2X1 g110695(.A (n_27125), .B (n_27089), .Y (n_27090));
NOR2X1 g110702(.A (n_26382), .B (n_26126), .Y (n_27088));
AND2X1 g110703(.A (n_27658), .B (n_28158), .Y (n_27086));
NAND2X1 g110704(.A (n_35040), .B (n_24386), .Y (n_27085));
NAND2X1 g110715(.A (n_27149), .B (n_34802), .Y (n_32060));
NAND2X1 g110722(.A (n_27658), .B (n_8954), .Y (n_27083));
NOR2X1 g110737(.A (n_26161), .B (n_24420), .Y (n_27082));
NAND2X1 g110740(.A (n_25673), .B (n_28364), .Y (n_27081));
NOR2X1 g110747(.A (n_27660), .B (n_25881), .Y (n_27080));
NAND2X1 g110764(.A (n_35519), .B (n_35233), .Y (n_28246));
NOR2X1 g107827(.A (n_26421), .B (n_26069), .Y (n_27079));
NAND2X1 g110773(.A (n_35233), .B (n_28053), .Y (n_27078));
INVX1 g110778(.A (n_27076), .Y (n_27077));
NAND3X1 g110807(.A (n_10234), .B (n_25642), .C (n_24391), .Y(n_27075));
AOI21X1 g110827(.A0 (n_14797), .A1 (n_26505), .B0 (n_8927), .Y(n_27074));
NAND3X1 g110838(.A (n_10141), .B (n_25629), .C (n_24351), .Y(n_27073));
NAND3X1 g110840(.A (n_10139), .B (n_25609), .C (n_25628), .Y(n_27072));
AOI21X1 g110849(.A0 (n_26513), .A1 (n_14983), .B0 (n_8927), .Y(n_27071));
INVX1 g110859(.A (n_27774), .Y (n_27069));
NAND2X1 g110864(.A (n_26109), .B (n_27068), .Y (n_28254));
INVX2 g110870(.A (n_27066), .Y (n_28252));
INVX1 g110901(.A (n_26565), .Y (n_27604));
NAND2X1 g110906(.A (n_26136), .B (n_27064), .Y (n_28276));
INVX1 g110915(.A (n_28793), .Y (n_27602));
INVX1 g110924(.A (n_26562), .Y (n_27601));
OAI21X1 g110930(.A0 (n_25582), .A1 (n_13647), .B0 (n_24675), .Y(n_28267));
INVX1 g110932(.A (n_27789), .Y (n_27062));
INVX1 g110934(.A (n_27061), .Y (n_28315));
INVX1 g110944(.A (n_26559), .Y (n_27599));
NAND2X1 g110948(.A (n_26119), .B (n_27059), .Y (n_28260));
INVX1 g110950(.A (n_27782), .Y (n_27058));
INVX1 g110974(.A (n_28796), .Y (n_27596));
NAND2X1 g110978(.A (n_26140), .B (n_25762), .Y (n_27056));
OAI21X1 g110988(.A0 (n_25263), .A1 (n_8977), .B0 (n_26111), .Y(n_27055));
AOI21X1 g110994(.A0 (n_27053), .A1 (n_26213), .B0 (n_21281), .Y(n_27054));
OAI21X1 g110997(.A0 (n_26522), .A1 (n_8382), .B0 (n_20286), .Y(n_27051));
NAND2X1 g111001(.A (n_20282), .B (n_26114), .Y (n_27050));
NAND2X1 g111057(.A (n_26117), .B (n_19307), .Y (n_27049));
NAND2X1 g111060(.A (n_26146), .B (n_25797), .Y (n_27048));
OAI21X1 g111063(.A0 (n_25269), .A1 (n_33340), .B0 (n_26122), .Y(n_27047));
OAI21X1 g111064(.A0 (n_26064), .A1 (n_27045), .B0 (n_25781), .Y(n_27046));
NAND2X1 g111072(.A (n_26143), .B (n_25729), .Y (n_27044));
OAI21X1 g107959(.A0 (n_35455), .A1 (n_27042), .B0 (n_15110), .Y(n_27043));
CLKBUFX1 gbuf_d_364(.A(n_26430), .Y(d_out_364));
CLKBUFX1 gbuf_q_364(.A(q_in_364), .Y(P2_reg2[1]));
INVX1 g107961(.A (n_27040), .Y (n_27041));
INVX1 g107962(.A (n_27040), .Y (n_27039));
NAND2X1 g111091(.A (n_32045), .B (n_32046), .Y (n_28265));
INVX2 g111099(.A (n_27739), .Y (n_27038));
NAND2X1 g111132(.A (n_25266), .B (n_29061), .Y (n_27036));
NAND2X1 g111151(.A (n_25266), .B (n_30563), .Y (n_27035));
NAND2X1 g111247(.A (n_27031), .B (n_10808), .Y (n_27033));
NAND2X1 g111248(.A (n_27031), .B (n_26528), .Y (n_27032));
NAND2X1 g111249(.A (n_27031), .B (n_26213), .Y (n_27029));
AND2X1 g111329(.A (n_27025), .B (n_28785), .Y (n_27028));
NAND2X1 g111330(.A (n_27025), .B (n_26112), .Y (n_27026));
NAND2X1 g111331(.A (n_27025), .B (n_26288), .Y (n_27024));
NAND2X1 g111332(.A (n_27025), .B (n_24526), .Y (n_27023));
OAI21X1 g111374(.A0 (n_27021), .A1 (n_12670), .B0 (n_27956), .Y(n_27022));
NAND2X1 g111416(.A (n_26493), .B (n_27018), .Y (n_28165));
NAND2X1 g111431(.A (n_27018), .B (n_14748), .Y (n_27019));
INVX1 g111432(.A (n_27609), .Y (n_27017));
NAND2X1 g111451(.A (n_27584), .B (n_28275), .Y (n_27016));
NAND2X1 g111452(.A (n_27584), .B (n_26528), .Y (n_27015));
NAND2X1 g108134(.A (n_26056), .B (n_31594), .Y (n_27014));
INVX1 g111635(.A (n_27637), .Y (n_27013));
NAND4X1 g108217(.A (n_15030), .B (n_25473), .C (n_25498), .D(n_25480), .Y (n_27012));
OAI21X1 g111702(.A0 (n_25571), .A1 (n_13163), .B0 (n_26514), .Y(n_28159));
INVX1 g111731(.A (n_27621), .Y (n_27011));
INVX1 g111735(.A (n_27625), .Y (n_27010));
AOI21X1 g108244(.A0 (n_26043), .A1 (n_26046), .B0 (n_27008), .Y(n_27009));
CLKBUFX1 gbuf_d_365(.A(n_26058), .Y(d_out_365));
CLKBUFX1 gbuf_q_365(.A(q_in_365), .Y(n_13727));
CLKBUFX1 gbuf_d_366(.A(n_26057), .Y(d_out_366));
CLKBUFX1 gbuf_q_366(.A(q_in_366), .Y(n_13732));
AOI21X1 g108262(.A0 (n_26039), .A1 (n_26045), .B0 (n_27008), .Y(n_27007));
NAND2X1 g108302(.A (n_26050), .B (n_33991), .Y (n_27006));
OR2X1 g111886(.A (n_27549), .B (n_29725), .Y (n_27005));
NAND2X1 g108319(.A (n_35341), .B (n_13130), .Y (n_27004));
NAND2X2 g108328(.A (n_35761), .B (n_35342), .Y (n_28154));
NAND3X1 g108341(.A (n_17991), .B (n_19836), .C (n_26029), .Y(n_27002));
NAND4X1 g108388(.A (n_14881), .B (n_25490), .C (n_25507), .D(n_25488), .Y (n_27001));
NAND2X1 g108405(.A (n_35341), .B (n_35515), .Y (n_27000));
NAND2X1 g108406(.A (n_35342), .B (n_22021), .Y (n_28151));
NOR2X1 g108468(.A (n_10416), .B (n_26060), .Y (n_26998));
OAI21X1 g108498(.A0 (n_9866), .A1 (n_28332), .B0 (n_26048), .Y(n_26997));
INVX1 g112352(.A (n_27565), .Y (n_28126));
INVX1 g112361(.A (n_26479), .Y (n_27527));
AOI22X1 g108530(.A0 (n_26028), .A1 (n_31528), .B0 (n_1485), .B1(n_35007), .Y (n_26996));
NOR2X1 g108533(.A (n_9940), .B (n_26059), .Y (n_26995));
AOI21X1 g108637(.A0 (n_33755), .A1 (n_28053), .B0 (n_13905), .Y(n_28155));
NOR2X1 g108647(.A (n_13746), .B (n_26055), .Y (n_26993));
NOR2X1 g108649(.A (n_14526), .B (n_26054), .Y (n_26992));
NOR2X1 g108651(.A (n_14523), .B (n_26053), .Y (n_26991));
AOI21X1 g108652(.A0 (n_21240), .A1 (n_15288), .B0 (n_26051), .Y(n_26990));
AOI21X1 g106941(.A0 (n_25961), .A1 (n_34773), .B0 (n_9430), .Y(n_26989));
NOR2X1 g108655(.A (n_14161), .B (n_26049), .Y (n_26987));
AOI21X1 g106958(.A0 (n_25954), .A1 (n_26985), .B0 (n_8942), .Y(n_26986));
NOR2X1 g108736(.A (n_26375), .B (n_26383), .Y (n_26984));
AOI21X1 g108745(.A0 (n_10376), .A1 (n_26003), .B0 (n_7058), .Y(n_26983));
NAND3X1 g108756(.A (n_26385), .B (n_25901), .C (n_20859), .Y(n_26982));
AOI21X1 g108776(.A0 (n_26978), .A1 (n_26896), .B0 (n_21232), .Y(n_26981));
OAI21X1 g108785(.A0 (n_26008), .A1 (n_25147), .B0 (n_33123), .Y(n_26980));
AOI21X1 g108791(.A0 (n_26978), .A1 (n_26898), .B0 (n_11325), .Y(n_26979));
NAND3X1 g108857(.A (n_25973), .B (n_25996), .C (n_26007), .Y(n_26977));
NAND3X1 g108886(.A (n_25917), .B (n_25987), .C (n_26004), .Y(n_26976));
NAND2X1 g108900(.A (n_26971), .B (n_26676), .Y (n_26975));
NAND2X1 g108901(.A (n_26969), .B (n_24101), .Y (n_26974));
NAND2X1 g108905(.A (n_26381), .B (n_25942), .Y (n_26973));
NAND2X1 g108939(.A (n_26971), .B (n_25554), .Y (n_26972));
NAND2X1 g108940(.A (n_26969), .B (n_28441), .Y (n_26970));
NOR2X1 g108949(.A (n_25531), .B (n_26409), .Y (n_26968));
NAND4X1 g108962(.A (n_19282), .B (n_23313), .C (n_25442), .D(n_23983), .Y (n_26967));
NAND2X1 g108991(.A (n_26969), .B (n_26965), .Y (n_26966));
NAND2X1 g108992(.A (n_26971), .B (n_22994), .Y (n_26964));
NAND2X1 g108995(.A (n_28874), .B (n_26823), .Y (n_26963));
NAND2X1 g109020(.A (n_26971), .B (n_23578), .Y (n_26962));
NAND2X1 g109022(.A (n_26969), .B (n_18137), .Y (n_26961));
NAND2X1 g109031(.A (n_26402), .B (n_10196), .Y (n_26960));
NAND2X1 g109032(.A (n_29430), .B (n_26958), .Y (n_26959));
NAND2X1 g109035(.A (n_18334), .B (n_26852), .Y (n_32059));
NAND2X1 g109054(.A (n_34859), .B (n_18348), .Y (n_32919));
NAND4X1 g109060(.A (n_25841), .B (n_25361), .C (n_24739), .D(n_25389), .Y (n_26952));
NAND2X1 g109065(.A (n_27523), .B (n_29684), .Y (n_26951));
NAND2X1 g109082(.A (n_34209), .B (n_35816), .Y (n_28084));
NOR2X1 g109087(.A (n_26394), .B (n_25171), .Y (n_26950));
NOR2X1 g109088(.A (n_26365), .B (n_10587), .Y (n_26949));
NOR2X1 g109089(.A (n_26364), .B (n_10581), .Y (n_26948));
NOR2X1 g109115(.A (n_26363), .B (n_10837), .Y (n_26947));
NAND3X1 g109119(.A (n_19109), .B (n_20901), .C (n_25885), .Y(n_26946));
AOI21X1 g109122(.A0 (n_26855), .A1 (n_14335), .B0 (n_8927), .Y(n_26945));
NAND4X1 g109157(.A (n_25883), .B (n_25177), .C (n_24794), .D(n_25434), .Y (n_26944));
NAND2X1 g109221(.A (n_34209), .B (n_22021), .Y (n_28081));
NAND3X1 g109232(.A (n_25952), .B (n_25990), .C (n_26006), .Y(n_26942));
AOI21X1 g109237(.A0 (n_26940), .A1 (n_27234), .B0 (n_20953), .Y(n_26941));
AOI21X1 g109251(.A0 (n_26938), .A1 (n_30180), .B0 (n_20937), .Y(n_26939));
NAND4X1 g109259(.A (n_19748), .B (n_23302), .C (n_25444), .D(n_23982), .Y (n_26937));
NOR2X1 g109269(.A (n_9567), .B (n_26370), .Y (n_26936));
NOR2X1 g109270(.A (n_9562), .B (n_26369), .Y (n_26935));
AOI21X1 g109275(.A0 (n_14803), .A1 (n_26826), .B0 (n_8927), .Y(n_26934));
AOI21X1 g109277(.A0 (n_14948), .A1 (n_26868), .B0 (n_8927), .Y(n_26933));
NOR2X1 g109282(.A (n_9555), .B (n_26367), .Y (n_26931));
AOI21X1 g109293(.A0 (n_24925), .A1 (n_26914), .B0 (n_26374), .Y(n_26930));
NAND2X2 g109309(.A (n_26405), .B (n_26929), .Y (n_35630));
NOR2X1 g109318(.A (n_26009), .B (n_26422), .Y (n_26928));
NAND4X1 g109324(.A (n_32136), .B (n_32137), .C (n_25367), .D(n_23014), .Y (n_26927));
NAND4X1 g109325(.A (n_32063), .B (n_32064), .C (n_25366), .D(n_23010), .Y (n_26926));
NAND2X1 g109350(.A (n_26420), .B (n_26925), .Y (n_28107));
NAND2X1 g109353(.A (n_26419), .B (n_26925), .Y (n_27386));
NAND2X1 g109362(.A (n_35109), .B (n_26924), .Y (n_28105));
NAND2X1 g109365(.A (n_26411), .B (n_26924), .Y (n_27382));
NAND2X1 g109376(.A (n_26408), .B (n_26923), .Y (n_27378));
NAND2X1 g109377(.A (n_26407), .B (n_26923), .Y (n_28103));
NAND4X1 g109394(.A (n_25836), .B (n_25858), .C (n_25155), .D(n_24734), .Y (n_26922));
AOI21X1 g109400(.A0 (n_26841), .A1 (n_14583), .B0 (n_26920), .Y(n_26921));
NAND3X1 g107249(.A (n_26346), .B (n_24700), .C (n_15078), .Y(n_26919));
NOR2X1 g109420(.A (n_25882), .B (n_26362), .Y (n_26918));
NAND3X1 g107250(.A (n_26345), .B (n_24689), .C (n_15066), .Y(n_26917));
AOI21X1 g109427(.A0 (n_26846), .A1 (n_29405), .B0 (n_14715), .Y(n_26916));
AOI21X1 g109429(.A0 (n_26914), .A1 (n_27522), .B0 (n_21332), .Y(n_26915));
AOI21X1 g109434(.A0 (n_26978), .A1 (n_26894), .B0 (n_10181), .Y(n_26913));
AOI21X1 g109447(.A0 (n_26978), .A1 (n_26892), .B0 (n_10143), .Y(n_26912));
NAND3X1 g109450(.A (n_24805), .B (n_26000), .C (n_24803), .Y(n_26911));
OAI21X1 g109459(.A0 (n_14275), .A1 (n_28659), .B0 (n_26036), .Y(n_26910));
OAI21X1 g109460(.A0 (n_15122), .A1 (n_25862), .B0 (n_26034), .Y(n_26909));
MX2X1 g109490(.A (n_19738), .B (n_21392), .S0 (n_25481), .Y(n_32870));
NAND4X1 g109496(.A (n_25532), .B (n_9596), .C (n_23721), .D(n_24861), .Y (n_26908));
NAND2X1 g109521(.A (n_33546), .B (n_26863), .Y (n_26904));
NAND2X1 g109525(.A (n_33546), .B (n_26832), .Y (n_26903));
OAI21X1 g109527(.A0 (n_25372), .A1 (n_23930), .B0 (n_31099), .Y(n_26902));
NOR2X1 g109530(.A (n_8677), .B (n_25895), .Y (n_26901));
NAND2X1 g109559(.A (n_26898), .B (n_29925), .Y (n_26899));
NAND2X1 g109569(.A (n_26896), .B (n_29925), .Y (n_26897));
NAND2X1 g109573(.A (n_26894), .B (n_29925), .Y (n_26895));
NAND2X1 g109574(.A (n_26892), .B (n_29925), .Y (n_26893));
NAND4X1 g109601(.A (n_15001), .B (n_24332), .C (n_24931), .D(n_24338), .Y (n_26891));
NAND4X1 g109602(.A (n_15018), .B (n_24601), .C (n_24930), .D(n_24603), .Y (n_26890));
NOR2X1 g109604(.A (n_25834), .B (n_14707), .Y (n_26889));
NAND2X1 g109621(.A (n_26881), .B (n_27999), .Y (n_26888));
NAND2X1 g109623(.A (n_26879), .B (n_13574), .Y (n_26887));
NAND2X1 g109631(.A (n_25967), .B (n_20084), .Y (n_26886));
NAND2X1 g109635(.A (n_26940), .B (n_29445), .Y (n_26885));
NAND3X1 g109638(.A (n_25159), .B (n_25438), .C (n_24781), .Y(n_26884));
NAND2X1 g109640(.A (n_26898), .B (n_26870), .Y (n_26883));
NAND2X1 g109659(.A (n_26881), .B (n_26412), .Y (n_35260));
NAND2X1 g109661(.A (n_26879), .B (n_13604), .Y (n_26880));
NAND3X1 g109670(.A (n_25158), .B (n_25436), .C (n_24775), .Y(n_26878));
NAND4X1 g109675(.A (n_35127), .B (n_35128), .C (n_11116), .D(n_24269), .Y (n_26877));
NAND2X1 g109687(.A (n_26881), .B (n_32739), .Y (n_26876));
NAND2X1 g109689(.A (n_26879), .B (n_32798), .Y (n_26875));
NAND2X1 g109696(.A (n_26938), .B (n_28431), .Y (n_26873));
NAND3X1 g109698(.A (n_25157), .B (n_25432), .C (n_24769), .Y(n_26872));
NAND2X1 g109700(.A (n_26896), .B (n_26870), .Y (n_26871));
NAND2X1 g109712(.A (n_26869), .B (n_26868), .Y (n_27424));
NAND2X1 g109721(.A (n_26881), .B (n_26866), .Y (n_26867));
NAND2X1 g109724(.A (n_26879), .B (n_23791), .Y (n_26865));
NAND2X1 g109729(.A (n_26863), .B (n_26660), .Y (n_26864));
NAND3X1 g109730(.A (n_25169), .B (n_25430), .C (n_24765), .Y(n_26862));
NAND4X1 g109732(.A (n_25813), .B (n_20932), .C (n_19113), .D(n_24265), .Y (n_26861));
NAND2X1 g109736(.A (n_26894), .B (n_26870), .Y (n_26860));
NAND2X1 g109746(.A (n_27632), .B (n_26857), .Y (n_26858));
NAND2X1 g109747(.A (n_29695), .B (n_26857), .Y (n_26856));
NAND2X1 g109748(.A (n_26780), .B (n_26855), .Y (n_27461));
NAND2X1 g109750(.A (n_26854), .B (n_26269), .Y (n_27459));
INVX1 g109752(.A (n_26852), .Y (n_26853));
NAND2X1 g109763(.A (n_25832), .B (n_18325), .Y (n_35929));
INVX1 g109765(.A (n_34859), .Y (n_26850));
NOR2X1 g109769(.A (n_24884), .B (n_25926), .Y (n_26848));
NAND2X1 g109773(.A (n_26846), .B (n_8954), .Y (n_26847));
NAND2X1 g109774(.A (n_24752), .B (n_26820), .Y (n_26845));
NAND2X1 g109775(.A (n_26842), .B (n_27109), .Y (n_26844));
NAND2X1 g109776(.A (n_24925), .B (n_26842), .Y (n_26843));
NAND2X1 g109777(.A (n_26777), .B (n_26841), .Y (n_27420));
NAND2X1 g109791(.A (n_14360), .B (n_26834), .Y (n_26840));
NAND2X1 g109792(.A (n_26837), .B (n_27109), .Y (n_26839));
NAND2X1 g109793(.A (n_27100), .B (n_26837), .Y (n_26838));
NAND2X1 g109794(.A (n_26837), .B (n_27632), .Y (n_26836));
NAND2X1 g109796(.A (n_26914), .B (n_26132), .Y (n_26835));
NAND2X1 g109797(.A (n_26834), .B (n_26775), .Y (n_27414));
NAND2X1 g109799(.A (n_26832), .B (n_26660), .Y (n_26833));
NAND2X1 g109811(.A (n_26892), .B (n_26870), .Y (n_26831));
NAND3X1 g109812(.A (n_10108), .B (n_19222), .C (n_25380), .Y(n_26830));
NOR2X1 g109814(.A (n_26382), .B (n_25896), .Y (n_26829));
NAND2X1 g109818(.A (n_26827), .B (n_28158), .Y (n_26828));
NAND2X1 g109821(.A (n_26785), .B (n_26826), .Y (n_27264));
NAND2X1 g107415(.A (n_25922), .B (n_29034), .Y (n_26825));
INVX1 g109822(.A (n_26823), .Y (n_26824));
NAND2X1 g109838(.A (n_26846), .B (n_30636), .Y (n_26822));
NAND2X1 g109839(.A (n_26820), .B (n_27902), .Y (n_26821));
NAND2X1 g109848(.A (n_25651), .B (n_24467), .Y (n_26819));
NAND2X1 g109851(.A (n_26812), .B (n_28136), .Y (n_26818));
NAND2X1 g109852(.A (n_26810), .B (n_28136), .Y (n_26816));
NAND4X1 g109853(.A (n_14822), .B (n_24342), .C (n_24946), .D(n_24340), .Y (n_26815));
NAND4X1 g109854(.A (n_14845), .B (n_24609), .C (n_24943), .D(n_24611), .Y (n_26814));
NAND2X1 g109858(.A (n_26812), .B (n_28158), .Y (n_26813));
NAND2X1 g109859(.A (n_26810), .B (n_28158), .Y (n_26811));
NAND2X1 g109864(.A (n_26807), .B (n_29405), .Y (n_26809));
NAND2X1 g109865(.A (n_26807), .B (n_33738), .Y (n_26808));
NAND2X1 g109867(.A (n_26286), .B (n_29405), .Y (n_26805));
AOI21X1 g109882(.A0 (n_26320), .A1 (n_30180), .B0 (n_21376), .Y(n_26804));
OAI21X1 g109891(.A0 (n_14469), .A1 (n_26801), .B0 (n_25962), .Y(n_26802));
AOI21X1 g109903(.A0 (n_26799), .A1 (n_30180), .B0 (n_19376), .Y(n_26800));
AOI21X1 g109917(.A0 (n_26769), .A1 (n_33802), .B0 (n_21360), .Y(n_26798));
NAND2X1 g107466(.A (n_25898), .B (n_29014), .Y (n_26797));
AOI21X1 g109927(.A0 (n_24925), .A1 (n_26273), .B0 (n_25861), .Y(n_26796));
INVX1 g109929(.A (n_26389), .Y (n_26794));
NOR2X1 g109935(.A (n_10358), .B (n_26005), .Y (n_26793));
AOI21X1 g109952(.A0 (n_26275), .A1 (n_14473), .B0 (n_8927), .Y(n_26792));
NAND2X1 g109961(.A (n_25958), .B (n_26791), .Y (n_27493));
OAI21X1 g109977(.A0 (n_25662), .A1 (n_25694), .B0 (n_13174), .Y(n_27229));
NAND2X1 g109979(.A (n_25977), .B (n_25949), .Y (n_26790));
OAI21X1 g109985(.A0 (n_26382), .A1 (n_25326), .B0 (n_25451), .Y(n_26789));
NOR2X1 g109991(.A (n_10343), .B (n_26001), .Y (n_26788));
NAND2X1 g110003(.A (n_25964), .B (n_24508), .Y (n_27495));
INVX1 g110049(.A (n_26377), .Y (n_27475));
NAND2X1 g110054(.A (n_25948), .B (n_26787), .Y (n_27500));
NAND2X1 g110079(.A (n_25911), .B (n_20868), .Y (n_26786));
OAI21X1 g110080(.A0 (n_25316), .A1 (n_13316), .B0 (n_24505), .Y(n_27498));
NAND2X1 g110087(.A (n_25872), .B (n_26785), .Y (n_35689));
OAI21X1 g110102(.A0 (n_14461), .A1 (n_14658), .B0 (n_25955), .Y(n_26784));
NAND2X1 g110103(.A (n_25909), .B (n_28136), .Y (n_26783));
AOI21X1 g110113(.A0 (n_26781), .A1 (n_26213), .B0 (n_19715), .Y(n_26782));
NAND2X1 g110117(.A (n_25940), .B (n_26780), .Y (n_27208));
NAND2X1 g110140(.A (n_25924), .B (n_29411), .Y (n_26779));
NAND2X1 g110141(.A (n_25920), .B (n_28136), .Y (n_26778));
NAND2X1 g110143(.A (n_25876), .B (n_26777), .Y (n_27445));
NAND2X1 g110145(.A (n_25875), .B (n_26776), .Y (n_27441));
NAND2X1 g110150(.A (n_25907), .B (n_26775), .Y (n_27436));
NAND2X1 g110154(.A (n_25904), .B (n_26774), .Y (n_27203));
NAND2X1 g110165(.A (n_25984), .B (n_25969), .Y (n_26773));
OAI21X1 g110170(.A0 (n_25695), .A1 (n_23487), .B0 (n_25981), .Y(n_26772));
NAND2X1 g110175(.A (n_25975), .B (n_25914), .Y (n_26771));
AOI21X1 g110185(.A0 (n_26769), .A1 (n_33513), .B0 (n_25992), .Y(n_26770));
NAND2X1 g107577(.A (n_25604), .B (n_31590), .Y (n_26767));
OAI21X1 g110225(.A0 (n_26366), .A1 (n_27662), .B0 (n_25928), .Y(n_26766));
MX2X1 g110232(.A (n_20783), .B (n_22512), .S0 (n_25373), .Y(n_27483));
NAND2X2 g110234(.A (n_25970), .B (n_25528), .Y (n_27479));
NAND2X1 g110239(.A (n_25517), .B (n_25945), .Y (n_27467));
INVX2 g110245(.A (n_34209), .Y (n_26765));
NOR2X1 g110265(.A (n_24922), .B (n_25720), .Y (n_26763));
NOR2X1 g110267(.A (n_25708), .B (n_25712), .Y (n_26762));
NAND2X1 g110269(.A (n_25824), .B (n_31781), .Y (n_26761));
NAND2X1 g110271(.A (n_25716), .B (n_31696), .Y (n_26760));
NOR2X1 g110279(.A (n_25670), .B (n_25710), .Y (n_26759));
NAND2X1 g110281(.A (n_26756), .B (n_26695), .Y (n_26758));
NAND2X1 g110282(.A (n_26756), .B (n_26672), .Y (n_26757));
NAND2X1 g110286(.A (n_33546), .B (n_25052), .Y (n_26755));
NAND2X1 g110288(.A (n_26756), .B (n_26653), .Y (n_26754));
OAI21X1 g110289(.A0 (n_25289), .A1 (n_24492), .B0 (n_30380), .Y(n_26753));
NAND2X1 g110291(.A (n_34712), .B (n_26639), .Y (n_26752));
NAND2X1 g110298(.A (n_34712), .B (n_26607), .Y (n_26751));
NAND2X1 g110302(.A (n_26756), .B (n_26596), .Y (n_32118));
NOR2X1 g110318(.A (n_25699), .B (n_26748), .Y (n_26749));
NAND2X1 g110320(.A (n_28948), .B (n_26735), .Y (n_26747));
NAND2X1 g110322(.A (n_28597), .B (n_26732), .Y (n_26746));
NAND2X1 g110327(.A (n_34770), .B (n_26730), .Y (n_26745));
NOR2X1 g110328(.A (n_25687), .B (n_26748), .Y (n_26744));
NOR2X1 g110329(.A (n_25678), .B (n_26748), .Y (n_26743));
NAND2X1 g110332(.A (n_34770), .B (n_26728), .Y (n_26742));
NAND2X1 g110337(.A (n_34770), .B (n_26726), .Y (n_26741));
AND2X1 g110341(.A (n_26739), .B (n_28926), .Y (n_26740));
AND2X1 g110342(.A (n_26719), .B (n_28926), .Y (n_26738));
AND2X1 g110345(.A (n_26717), .B (n_28926), .Y (n_26737));
AND2X1 g110350(.A (n_26735), .B (n_34709), .Y (n_26736));
AND2X1 g110353(.A (n_26711), .B (n_34708), .Y (n_26734));
NAND2X1 g110354(.A (n_26732), .B (n_34709), .Y (n_26733));
NAND2X1 g110356(.A (n_26730), .B (n_34709), .Y (n_26731));
NAND2X1 g110361(.A (n_26728), .B (n_29925), .Y (n_26729));
NAND2X1 g110366(.A (n_26726), .B (n_29925), .Y (n_26727));
NAND2X1 g110368(.A (n_26703), .B (n_25988), .Y (n_26725));
NOR2X1 g110369(.A (n_25678), .B (n_8319), .Y (n_26723));
NAND2X1 g110374(.A (n_26739), .B (n_28013), .Y (n_26721));
NAND2X1 g110375(.A (n_26719), .B (n_28013), .Y (n_26720));
NAND2X1 g110379(.A (n_26717), .B (n_33785), .Y (n_26718));
NAND2X1 g110386(.A (n_26735), .B (n_28915), .Y (n_26716));
NAND2X1 g110387(.A (n_26092), .B (n_33784), .Y (n_26715));
NAND2X1 g110390(.A (n_26732), .B (n_29455), .Y (n_26713));
NAND2X1 g110392(.A (n_26711), .B (n_28013), .Y (n_26712));
NAND2X1 g110394(.A (n_26730), .B (n_28013), .Y (n_26710));
NAND2X1 g110399(.A (n_26728), .B (n_28013), .Y (n_26708));
NAND2X1 g110405(.A (n_26085), .B (n_33784), .Y (n_26707));
NAND2X1 g110406(.A (n_26082), .B (n_33785), .Y (n_26706));
NAND2X1 g110408(.A (n_26726), .B (n_28013), .Y (n_26705));
NAND2X1 g110410(.A (n_26703), .B (n_33785), .Y (n_26704));
NAND2X1 g110417(.A (n_26690), .B (n_25309), .Y (n_26702));
NAND2X1 g110441(.A (n_27253), .B (n_29445), .Y (n_26700));
NAND4X1 g110443(.A (n_18764), .B (n_23719), .C (n_23738), .D(n_24869), .Y (n_26699));
NAND2X1 g110448(.A (n_26655), .B (n_25554), .Y (n_26698));
NOR2X1 g110457(.A (n_23883), .B (n_25794), .Y (n_26697));
NAND2X1 g110459(.A (n_26695), .B (n_10808), .Y (n_26696));
NAND2X1 g110461(.A (n_26677), .B (n_25554), .Y (n_26694));
NAND2X1 g110462(.A (n_26648), .B (n_28441), .Y (n_26692));
NAND2X1 g110463(.A (n_26690), .B (n_25297), .Y (n_26691));
NAND2X1 g110465(.A (n_17713), .B (n_34838), .Y (n_26689));
NAND2X1 g110466(.A (n_26643), .B (n_28441), .Y (n_26688));
NAND2X1 g110468(.A (n_34496), .B (n_18384), .Y (n_26687));
NAND2X1 g110471(.A (n_26629), .B (n_28441), .Y (n_26684));
NAND2X1 g110477(.A (n_34838), .B (n_24101), .Y (n_26683));
AOI21X1 g110478(.A0 (n_9629), .A1 (n_17305), .B0 (n_25817), .Y(n_26680));
NAND2X1 g110483(.A (n_26677), .B (n_26676), .Y (n_26678));
NOR2X1 g110484(.A (n_25701), .B (n_8678), .Y (n_26675));
NAND2X1 g110489(.A (n_26672), .B (n_34753), .Y (n_26673));
NAND2X1 g110490(.A (n_26690), .B (n_32815), .Y (n_26671));
NAND2X1 g110492(.A (n_34496), .B (n_32786), .Y (n_26670));
NAND2X1 g110495(.A (n_25052), .B (n_24629), .Y (n_26668));
AND2X1 g110499(.A (n_26663), .B (n_26665), .Y (n_26666));
NAND2X1 g110500(.A (n_26663), .B (n_26662), .Y (n_26664));
NAND2X1 g110501(.A (n_26663), .B (n_26660), .Y (n_26661));
NAND2X1 g110507(.A (n_27247), .B (n_28431), .Y (n_26659));
NOR2X1 g110512(.A (n_26657), .B (n_27564), .Y (n_26658));
NAND2X1 g110516(.A (n_26655), .B (n_24361), .Y (n_26656));
NAND2X1 g110523(.A (n_26653), .B (n_34753), .Y (n_26654));
NAND2X1 g110528(.A (n_26690), .B (n_34688), .Y (n_26652));
NAND2X1 g110529(.A (n_26677), .B (n_35054), .Y (n_26650));
NAND2X1 g110530(.A (n_26648), .B (n_35054), .Y (n_26649));
NAND2X1 g110531(.A (n_34496), .B (n_24984), .Y (n_26647));
NAND2X1 g110533(.A (n_34838), .B (n_22994), .Y (n_26646));
NAND2X1 g110534(.A (n_26643), .B (n_24361), .Y (n_26644));
NAND2X1 g110546(.A (n_26639), .B (n_26660), .Y (n_26640));
NAND2X1 g110554(.A (n_26655), .B (n_26637), .Y (n_26638));
NOR2X1 g110558(.A (n_23882), .B (n_25717), .Y (n_26636));
NAND2X1 g110561(.A (n_26677), .B (n_23578), .Y (n_26635));
NAND2X1 g110562(.A (n_26648), .B (n_27950), .Y (n_26634));
NAND2X1 g110563(.A (n_26643), .B (n_26637), .Y (n_26633));
NAND2X1 g110564(.A (n_34838), .B (n_26631), .Y (n_26632));
NAND2X1 g110567(.A (n_26629), .B (n_13274), .Y (n_26630));
NAND2X1 g110569(.A (n_25829), .B (n_18329), .Y (n_26628));
NAND2X1 g110576(.A (n_27462), .B (n_26626), .Y (n_26627));
NAND3X1 g110584(.A (n_32237), .B (n_20335), .C (n_23220), .Y(n_26625));
NAND3X1 g110586(.A (n_25722), .B (n_25258), .C (n_25259), .Y(n_26624));
NAND2X1 g110601(.A (n_26609), .B (n_18546), .Y (n_27102));
NAND3X1 g110614(.A (n_25362), .B (n_25274), .C (n_19341), .Y(n_26623));
NAND2X1 g110621(.A (n_26620), .B (n_8990), .Y (n_26622));
NAND2X1 g110623(.A (n_26620), .B (n_27522), .Y (n_26621));
NAND2X1 g110631(.A (n_26594), .B (n_33738), .Y (n_26619));
NAND2X1 g110641(.A (n_26585), .B (n_35744), .Y (n_27757));
NAND2X1 g110643(.A (n_35816), .B (n_33812), .Y (n_27760));
NAND2X1 g110654(.A (n_26615), .B (n_29505), .Y (n_26616));
NAND2X1 g110655(.A (n_26615), .B (n_26255), .Y (n_26614));
NAND2X1 g110663(.A (n_27235), .B (n_29191), .Y (n_26613));
NAND2X1 g110665(.A (n_27235), .B (n_26611), .Y (n_26612));
NAND2X1 g110673(.A (n_26609), .B (n_35736), .Y (n_26610));
NAND2X1 g110674(.A (n_26607), .B (n_28890), .Y (n_26608));
NAND2X1 g110682(.A (n_26655), .B (n_25098), .Y (n_26606));
NAND2X1 g110685(.A (n_27100), .B (n_26602), .Y (n_26605));
NAND2X1 g110686(.A (n_27614), .B (n_26602), .Y (n_26603));
NOR2X1 g110701(.A (n_23881), .B (n_25715), .Y (n_26601));
NAND2X1 g110709(.A (n_26648), .B (n_24101), .Y (n_26600));
NAND2X1 g110710(.A (n_26643), .B (n_24101), .Y (n_26599));
NAND2X1 g110713(.A (n_26629), .B (n_27091), .Y (n_26598));
NAND2X1 g110716(.A (n_26596), .B (n_10808), .Y (n_26597));
NAND2X1 g110730(.A (n_26594), .B (n_28158), .Y (n_26595));
NAND2X1 g110731(.A (n_26594), .B (n_28374), .Y (n_35607));
NOR2X1 g110746(.A (n_27193), .B (n_25881), .Y (n_26591));
NAND2X1 g110752(.A (n_26588), .B (n_30636), .Y (n_26590));
NAND2X1 g110758(.A (n_26588), .B (n_29405), .Y (n_26589));
NAND2X1 g110759(.A (n_33812), .B (n_35578), .Y (n_26587));
CLKBUFX1 gbuf_d_367(.A(n_25576), .Y(d_out_367));
CLKBUFX1 gbuf_q_367(.A(q_in_367), .Y(n_14168));
NAND2X1 g110766(.A (n_26609), .B (n_35500), .Y (n_27764));
NAND2X1 g110774(.A (n_26585), .B (n_26584), .Y (n_27754));
INVX1 g110775(.A (n_26582), .Y (n_26583));
NAND2X1 g110777(.A (n_26609), .B (n_28053), .Y (n_26581));
NAND2X1 g110779(.A (n_33812), .B (n_26584), .Y (n_27076));
NAND2X1 g110786(.A (n_26588), .B (n_33738), .Y (n_26580));
NAND2X2 g110795(.A (n_26585), .B (n_35578), .Y (n_26577));
OAI21X1 g110812(.A0 (n_14832), .A1 (n_26372), .B0 (n_25789), .Y(n_26576));
INVX1 g110829(.A (n_26221), .Y (n_26575));
NAND2X1 g110846(.A (n_25812), .B (n_29505), .Y (n_26574));
NAND2X1 g110852(.A (n_25808), .B (n_29133), .Y (n_26573));
NAND2X1 g110854(.A (n_25788), .B (n_29132), .Y (n_26572));
NAND2X1 g110856(.A (n_25771), .B (n_26570), .Y (n_26571));
NAND2X1 g110858(.A (n_25770), .B (n_25856), .Y (n_27822));
NAND2X1 g110860(.A (n_25752), .B (n_26216), .Y (n_27774));
NAND2X1 g110871(.A (n_25750), .B (n_26569), .Y (n_27066));
NAND2X1 g110874(.A (n_25129), .B (n_25766), .Y (n_26568));
AOI21X1 g110890(.A0 (n_26157), .A1 (n_34952), .B0 (n_15161), .Y(n_32161));
AOI21X1 g110893(.A0 (n_35359), .A1 (n_29061), .B0 (n_15154), .Y(n_32113));
INVX1 g110896(.A (n_28279), .Y (n_27065));
OAI21X1 g110902(.A0 (n_34696), .A1 (n_13817), .B0 (n_26208), .Y(n_26565));
NAND2X1 g110910(.A (n_25810), .B (n_26564), .Y (n_27800));
NAND2X1 g110913(.A (n_25807), .B (n_25852), .Y (n_27825));
OAI21X1 g110916(.A0 (n_25255), .A1 (n_26204), .B0 (n_26207), .Y(n_28793));
INVX1 g110919(.A (n_28270), .Y (n_27063));
OAI21X1 g110925(.A0 (n_34696), .A1 (n_14116), .B0 (n_26203), .Y(n_26562));
NAND2X1 g110933(.A (n_25791), .B (n_14128), .Y (n_27789));
NAND2X1 g110935(.A (n_25774), .B (n_26202), .Y (n_27061));
INVX1 g110940(.A (n_27322), .Y (n_26560));
OAI21X1 g110945(.A0 (n_34696), .A1 (n_32707), .B0 (n_26199), .Y(n_26559));
NAND2X1 g110951(.A (n_25772), .B (n_26558), .Y (n_27782));
INVX1 g110957(.A (n_27319), .Y (n_26557));
NAND2X1 g110968(.A (n_25746), .B (n_25850), .Y (n_27820));
NAND2X1 g110972(.A (n_25735), .B (n_25849), .Y (n_27817));
OAI21X1 g110975(.A0 (n_25255), .A1 (n_26210), .B0 (n_26193), .Y(n_28796));
AOI21X1 g110990(.A0 (n_24743), .A1 (n_26553), .B0 (n_25749), .Y(n_26554));
NOR2X1 g111014(.A (n_24605), .B (n_25667), .Y (n_26552));
NOR2X1 g111015(.A (n_24918), .B (n_25666), .Y (n_26551));
INVX1 g111041(.A (n_27277), .Y (n_26550));
NAND2X1 g111044(.A (n_25737), .B (n_26548), .Y (n_26549));
NAND2X1 g111059(.A (n_25134), .B (n_25802), .Y (n_26547));
NAND2X1 g111071(.A (n_25126), .B (n_25732), .Y (n_26546));
AOI21X1 g107963(.A0 (n_25593), .A1 (n_25235), .B0 (n_24975), .Y(n_27040));
NAND2X1 g111096(.A (n_25745), .B (n_25399), .Y (n_27771));
NAND2X2 g111097(.A (n_32596), .B (n_32597), .Y (n_27803));
NAND2X1 g111098(.A (n_25740), .B (n_25393), .Y (n_27766));
NAND2X1 g111101(.A (n_25739), .B (n_25392), .Y (n_27739));
NAND2X1 g111126(.A (n_26541), .B (n_28864), .Y (n_26545));
NAND2X1 g111141(.A (n_26538), .B (n_28864), .Y (n_26543));
NAND2X1 g111145(.A (n_26541), .B (n_28485), .Y (n_26542));
NOR2X1 g111152(.A (n_25587), .B (n_8319), .Y (n_26540));
NAND2X1 g111162(.A (n_26538), .B (n_30563), .Y (n_26539));
NAND2X1 g111169(.A (n_26541), .B (n_26535), .Y (n_26536));
NOR2X1 g111183(.A (n_23701), .B (n_25583), .Y (n_26534));
NAND2X1 g111190(.A (n_26538), .B (n_26535), .Y (n_26533));
NAND2X1 g111203(.A (n_26520), .B (n_27999), .Y (n_26532));
NAND2X1 g111206(.A (n_33233), .B (n_26530), .Y (n_26531));
NAND2X1 g111250(.A (n_27053), .B (n_26528), .Y (n_26529));
NAND2X1 g111262(.A (n_25003), .B (n_33233), .Y (n_32121));
NAND2X1 g111277(.A (n_25270), .B (n_26288), .Y (n_26525));
INVX1 g111278(.A (n_26123), .Y (n_26524));
NOR2X1 g111280(.A (n_26522), .B (n_8285), .Y (n_26523));
NAND2X1 g111298(.A (n_26520), .B (n_32664), .Y (n_26521));
NAND2X1 g111302(.A (n_33233), .B (n_32815), .Y (n_26519));
NAND2X1 g111342(.A (n_26520), .B (n_26866), .Y (n_26517));
NAND2X1 g111345(.A (n_33233), .B (n_34688), .Y (n_26516));
NAND2X1 g111385(.A (n_25331), .B (n_26508), .Y (n_27634));
NAND2X1 g111389(.A (n_26514), .B (n_26513), .Y (n_27630));
NAND2X1 g111417(.A (n_14978), .B (n_26510), .Y (n_26511));
NAND2X1 g111433(.A (n_26510), .B (n_26074), .Y (n_27609));
NAND2X1 g111442(.A (n_26508), .B (n_14375), .Y (n_26509));
OAI21X1 g111474(.A0 (n_9172), .A1 (n_25242), .B0 (n_23169), .Y(n_26507));
NAND2X1 g111477(.A (n_25652), .B (n_23167), .Y (n_26506));
NAND2X1 g111495(.A (n_24709), .B (n_26505), .Y (n_27613));
NOR2X1 g111500(.A (n_23688), .B (n_25584), .Y (n_26504));
AOI21X1 g108135(.A0 (n_10397), .A1 (n_25543), .B0 (n_31343), .Y(n_26503));
NAND2X1 g108158(.A (n_35455), .B (n_1054), .Y (n_26502));
NAND2X1 g111555(.A (n_25618), .B (n_25713), .Y (n_27649));
NAND2X1 g111586(.A (n_25624), .B (n_25705), .Y (n_27651));
NAND2X1 g111636(.A (n_25616), .B (n_25689), .Y (n_27637));
NAND2X1 g111637(.A (n_25606), .B (n_25679), .Y (n_27645));
NAND2X1 g111642(.A (n_25615), .B (n_25684), .Y (n_27647));
OAI21X1 g111644(.A0 (n_25244), .A1 (n_27696), .B0 (n_24411), .Y(n_26500));
OAI21X1 g111647(.A0 (n_25243), .A1 (n_27696), .B0 (n_25658), .Y(n_26499));
INVX1 g111649(.A (n_27116), .Y (n_26498));
INVX1 g111668(.A (n_27105), .Y (n_26497));
INVX1 g111672(.A (n_27094), .Y (n_26496));
AOI21X1 g108232(.A0 (n_25557), .A1 (n_18303), .B0 (n_8942), .Y(n_26494));
NAND2X1 g111732(.A (n_25598), .B (n_26493), .Y (n_27621));
NAND2X1 g111736(.A (n_25600), .B (n_25387), .Y (n_27625));
NAND2X1 g111744(.A (n_25603), .B (n_25400), .Y (n_27619));
OAI21X1 g111776(.A0 (n_25241), .A1 (n_34719), .B0 (n_24412), .Y(n_26492));
OAI21X1 g111777(.A0 (n_25240), .A1 (n_34719), .B0 (n_25659), .Y(n_26491));
CLKBUFX1 gbuf_d_368(.A(n_25960), .Y(d_out_368));
CLKBUFX1 gbuf_q_368(.A(q_in_368), .Y(n_10562));
CLKBUFX1 gbuf_d_369(.A(n_25668), .Y(d_out_369));
CLKBUFX1 gbuf_q_369(.A(q_in_369), .Y(P1_reg1[0]));
CLKBUFX1 gbuf_d_370(.A(n_25669), .Y(d_out_370));
CLKBUFX1 gbuf_q_370(.A(q_in_370), .Y(n_10187));
CLKBUFX1 gbuf_d_371(.A(n_25575), .Y(d_out_371));
CLKBUFX1 gbuf_q_371(.A(q_in_371), .Y(n_14513));
CLKBUFX1 gbuf_d_372(.A(n_25574), .Y(d_out_372));
CLKBUFX1 gbuf_q_372(.A(q_in_372), .Y(P3_reg2[30]));
AOI21X1 g108263(.A0 (n_25556), .A1 (n_14172), .B0 (n_8942), .Y(n_26490));
OAI21X1 g108300(.A0 (n_25559), .A1 (n_25537), .B0 (n_30956), .Y(n_26488));
NAND2X1 g108303(.A (n_35456), .B (n_29405), .Y (n_26487));
OR2X1 g111885(.A (n_27021), .B (n_10790), .Y (n_26486));
AOI21X1 g108321(.A0 (n_25553), .A1 (n_21293), .B0 (n_8942), .Y(n_26485));
NOR2X1 g111904(.A (n_27021), .B (n_8679), .Y (n_26483));
OAI21X1 g108399(.A0 (n_25548), .A1 (n_25558), .B0 (n_35008), .Y(n_26482));
OAI21X1 g108438(.A0 (n_8864), .A1 (n_35012), .B0 (n_25569), .Y(n_26481));
INVX1 g112329(.A (n_27031), .Y (n_26480));
NAND2X1 g112331(.A (n_25581), .B (n_25590), .Y (n_27579));
INVX2 g112353(.A (n_26063), .Y (n_27565));
OAI21X1 g112362(.A0 (n_25232), .A1 (n_32662), .B0 (n_23181), .Y(n_26479));
NAND2X1 g112375(.A (n_25580), .B (n_24892), .Y (n_27577));
NAND2X1 g112380(.A (n_25578), .B (n_24890), .Y (n_27575));
NAND4X1 g108630(.A (n_23475), .B (n_21760), .C (n_21271), .D(n_25210), .Y (n_26478));
OAI21X1 g108653(.A0 (n_25538), .A1 (n_26052), .B0 (n_14520), .Y(n_26477));
AOI21X1 g108743(.A0 (n_10423), .A1 (n_25520), .B0 (n_30968), .Y(n_26476));
NAND3X1 g108751(.A (n_26020), .B (n_25500), .C (n_20390), .Y(n_26475));
NAND2X1 g108782(.A (n_26456), .B (n_7967), .Y (n_26474));
OAI21X1 g108783(.A0 (n_25508), .A1 (n_24354), .B0 (n_33123), .Y(n_26473));
NAND3X1 g108794(.A (n_19119), .B (n_20933), .C (n_25530), .Y(n_26472));
OAI21X1 g108795(.A0 (n_25455), .A1 (n_23175), .B0 (n_29633), .Y(n_26471));
NAND4X1 g108800(.A (n_24040), .B (n_25065), .C (n_25146), .D(n_23990), .Y (n_26470));
NAND2X1 g108854(.A (n_26024), .B (n_31097), .Y (n_26466));
NAND2X1 g108862(.A (n_26023), .B (n_31534), .Y (n_26465));
NAND2X1 g108903(.A (n_26015), .B (n_26458), .Y (n_26464));
NAND2X1 g108942(.A (n_26014), .B (n_9431), .Y (n_26463));
AOI21X1 g108946(.A0 (n_25522), .A1 (n_29667), .B0 (n_8940), .Y(n_26462));
NAND4X1 g108948(.A (n_35124), .B (n_35125), .C (n_23452), .D(n_24169), .Y (n_26461));
NAND2X1 g108993(.A (n_26016), .B (n_8641), .Y (n_26460));
NAND2X1 g109025(.A (n_26013), .B (n_26458), .Y (n_26459));
NAND2X1 g109033(.A (n_26456), .B (n_34802), .Y (n_26457));
AOI21X1 g109040(.A0 (n_25514), .A1 (n_29666), .B0 (n_25867), .Y(n_26455));
NAND2X1 g109052(.A (n_33755), .B (n_18546), .Y (n_27537));
NAND2X1 g109084(.A (n_34187), .B (n_35790), .Y (n_27544));
NAND2X1 g109109(.A (n_33754), .B (n_35744), .Y (n_26450));
AOI21X1 g109127(.A0 (n_26400), .A1 (n_14398), .B0 (n_8927), .Y(n_26449));
OAI21X1 g109178(.A0 (n_25533), .A1 (n_29681), .B0 (n_10413), .Y(n_26447));
NAND2X1 g109220(.A (n_35528), .B (n_33754), .Y (n_27539));
NAND2X1 g109223(.A (n_34187), .B (n_25877), .Y (n_27542));
NAND2X2 g109231(.A (n_35528), .B (n_34187), .Y (n_26444));
OAI21X1 g109236(.A0 (n_25527), .A1 (n_29681), .B0 (n_10436), .Y(n_26443));
OAI21X1 g109244(.A0 (n_14485), .A1 (n_14916), .B0 (n_26042), .Y(n_26442));
OAI21X1 g109245(.A0 (n_25523), .A1 (n_29681), .B0 (n_10378), .Y(n_26441));
OAI21X1 g109249(.A0 (n_15125), .A1 (n_8614), .B0 (n_26038), .Y(n_26440));
NAND4X1 g109261(.A (n_25595), .B (n_19911), .C (n_23450), .D(n_24168), .Y (n_26439));
AOI21X1 g109276(.A0 (n_14858), .A1 (n_26397), .B0 (n_8927), .Y(n_26438));
NAND3X1 g109283(.A (n_9185), .B (n_25506), .C (n_20398), .Y(n_26436));
NAND3X1 g109284(.A (n_9056), .B (n_25503), .C (n_20890), .Y(n_26435));
NAND3X1 g109290(.A (n_9050), .B (n_25501), .C (n_20871), .Y(n_26434));
NAND3X1 g109326(.A (n_24806), .B (n_25502), .C (n_24809), .Y(n_26433));
NOR2X1 g109338(.A (n_26032), .B (n_14474), .Y (n_26432));
AOI21X1 g107248(.A0 (n_29068), .A1 (n_32532), .B0 (n_25456), .Y(n_26431));
OAI21X1 g109474(.A0 (n_25178), .A1 (n_34300), .B0 (n_6734), .Y(n_26430));
AOI21X1 g109483(.A0 (n_26428), .A1 (n_28136), .B0 (n_20380), .Y(n_35919));
AOI21X1 g109534(.A0 (n_28597), .A1 (n_25982), .B0 (n_25369), .Y(n_26427));
AOI21X1 g109536(.A0 (n_9503), .A1 (n_25991), .B0 (n_25364), .Y(n_26426));
NOR2X1 g109578(.A (n_23629), .B (n_25461), .Y (n_26425));
NOR2X1 g109583(.A (n_23628), .B (n_25460), .Y (n_26424));
NAND3X1 g109594(.A (n_14249), .B (n_25137), .C (n_10230), .Y(n_26423));
NAND4X1 g109599(.A (n_15081), .B (n_24018), .C (n_24616), .D(n_24021), .Y (n_26422));
NAND3X1 g109600(.A (n_14654), .B (n_25128), .C (n_10151), .Y(n_26421));
NAND2X1 g109626(.A (n_35163), .B (n_18399), .Y (n_26420));
NAND2X1 g109627(.A (n_35151), .B (n_27999), .Y (n_26419));
NAND2X1 g109630(.A (n_20083), .B (n_25966), .Y (n_26418));
NAND2X1 g109632(.A (n_26416), .B (n_26415), .Y (n_26417));
NAND2X1 g109663(.A (n_35163), .B (n_26412), .Y (n_35109));
NAND2X1 g109664(.A (n_35151), .B (n_23270), .Y (n_26411));
NAND4X1 g109680(.A (n_19928), .B (n_24669), .C (n_24699), .D(n_24402), .Y (n_26409));
NAND2X1 g109690(.A (n_35152), .B (n_32794), .Y (n_26408));
NAND2X1 g109691(.A (n_35164), .B (n_32739), .Y (n_26407));
NAND2X1 g109725(.A (n_35152), .B (n_27470), .Y (n_26405));
NAND2X2 g109726(.A (n_35164), .B (n_27470), .Y (n_26404));
INVX1 g109738(.A (n_26456), .Y (n_26402));
NAND2X1 g109749(.A (n_26401), .B (n_26400), .Y (n_26958));
NAND3X1 g109753(.A (n_32217), .B (n_21431), .C (n_32218), .Y(n_26852));
NAND2X1 g109764(.A (n_18965), .B (n_34514), .Y (n_35930));
NAND2X1 g109823(.A (n_26398), .B (n_26397), .Y (n_26823));
NOR2X1 g109840(.A (n_25125), .B (n_25457), .Y (n_26396));
AOI21X1 g109842(.A0 (n_28597), .A1 (n_25647), .B0 (n_24801), .Y(n_26395));
NAND4X1 g109855(.A (n_15058), .B (n_24025), .C (n_24625), .D(n_24023), .Y (n_26394));
AOI21X1 g109879(.A0 (n_26392), .A1 (n_27234), .B0 (n_19379), .Y(n_26393));
OAI21X1 g109896(.A0 (n_14929), .A1 (n_29968), .B0 (n_25525), .Y(n_26391));
INVX1 g109924(.A (n_26021), .Y (n_26390));
AOI21X1 g109930(.A0 (n_14950), .A1 (n_25873), .B0 (n_8927), .Y(n_26389));
NOR2X1 g109932(.A (n_25076), .B (n_25454), .Y (n_26387));
AOI21X1 g109934(.A0 (n_27100), .A1 (n_25927), .B0 (n_25464), .Y(n_26386));
AOI21X1 g109950(.A0 (n_27100), .A1 (n_25900), .B0 (n_25160), .Y(n_26385));
OAI21X1 g109980(.A0 (n_26382), .A1 (n_25030), .B0 (n_25453), .Y(n_26383));
OAI21X1 g109986(.A0 (n_25020), .A1 (n_24312), .B0 (n_33792), .Y(n_26381));
AOI21X1 g109989(.A0 (n_34770), .A1 (n_25995), .B0 (n_14341), .Y(n_26380));
AOI21X1 g109990(.A0 (n_34770), .A1 (n_25986), .B0 (n_14785), .Y(n_26379));
OAI21X1 g110050(.A0 (n_25317), .A1 (n_13579), .B0 (n_26376), .Y(n_26377));
NAND2X1 g110074(.A (n_25505), .B (n_20397), .Y (n_26375));
AOI21X1 g110104(.A0 (n_25921), .A1 (n_14716), .B0 (n_29725), .Y(n_26374));
OAI21X1 g110138(.A0 (n_14698), .A1 (n_26372), .B0 (n_25519), .Y(n_26373));
NAND2X1 g110144(.A (n_25474), .B (n_26371), .Y (n_27523));
OAI21X1 g110195(.A0 (n_26361), .A1 (n_28528), .B0 (n_20435), .Y(n_26370));
OAI21X1 g110196(.A0 (n_26368), .A1 (n_27192), .B0 (n_20915), .Y(n_26369));
OAI21X1 g110200(.A0 (n_26366), .A1 (n_27192), .B0 (n_20893), .Y(n_26367));
NAND2X1 g110205(.A (n_25471), .B (n_20492), .Y (n_26365));
OAI21X1 g110206(.A0 (n_20229), .A1 (n_25540), .B0 (n_25466), .Y(n_26364));
NAND2X1 g110209(.A (n_25477), .B (n_20858), .Y (n_26363));
OAI21X1 g110220(.A0 (n_26361), .A1 (n_27662), .B0 (n_25516), .Y(n_26362));
AOI21X1 g110229(.A0 (n_25890), .A1 (n_28136), .B0 (n_20400), .Y(n_26360));
MX2X1 g110241(.A (n_19732), .B (n_21387), .S0 (n_25078), .Y(n_26971));
MX2X1 g110242(.A (n_21259), .B (n_21258), .S0 (n_25075), .Y(n_26969));
INVX1 g110253(.A (n_34187), .Y (n_26359));
NAND4X1 g110263(.A (n_24608), .B (n_9598), .C (n_24556), .D(n_24273), .Y (n_26358));
NOR2X1 g110268(.A (n_25337), .B (n_25354), .Y (n_26357));
NAND2X1 g110272(.A (n_25360), .B (n_31698), .Y (n_26356));
NAND3X1 g110275(.A (n_25359), .B (n_24933), .C (n_19839), .Y(n_26355));
NOR2X1 g110283(.A (n_25324), .B (n_11567), .Y (n_26354));
NAND2X1 g110287(.A (n_33546), .B (n_26292), .Y (n_26353));
OAI21X1 g110294(.A0 (n_24962), .A1 (n_24136), .B0 (n_24695), .Y(n_26352));
NOR2X1 g110301(.A (n_24909), .B (n_25377), .Y (n_26351));
AOI21X1 g110303(.A0 (n_26978), .A1 (n_25820), .B0 (n_20223), .Y(n_26350));
NAND2X1 g110305(.A (n_27614), .B (n_26249), .Y (n_26349));
NAND2X1 g110323(.A (n_29065), .B (n_26340), .Y (n_26348));
NOR2X1 g110324(.A (n_27169), .B (n_25347), .Y (n_26347));
NAND2X1 g110330(.A (n_34770), .B (n_26338), .Y (n_26346));
NAND2X1 g110336(.A (n_34770), .B (n_26336), .Y (n_26345));
AND2X1 g110343(.A (n_32532), .B (n_28926), .Y (n_26344));
NAND2X1 g110346(.A (n_26333), .B (n_30563), .Y (n_26342));
AND2X1 g110351(.A (n_26340), .B (n_34709), .Y (n_26341));
NAND2X1 g110357(.A (n_26338), .B (n_34709), .Y (n_26339));
NAND2X1 g110365(.A (n_26336), .B (n_34709), .Y (n_26337));
NAND2X1 g110376(.A (n_32532), .B (n_28013), .Y (n_26335));
NAND2X1 g110380(.A (n_26333), .B (n_30197), .Y (n_26334));
NAND2X1 g110382(.A (n_25698), .B (n_29604), .Y (n_26332));
NAND2X1 g110388(.A (n_26340), .B (n_28915), .Y (n_26331));
NAND2X1 g110393(.A (n_25686), .B (n_26535), .Y (n_26330));
NAND2X1 g110395(.A (n_26338), .B (n_28013), .Y (n_26328));
NAND3X1 g110400(.A (n_25357), .B (n_24990), .C (n_19357), .Y(n_26327));
NAND2X1 g110407(.A (n_26336), .B (n_28013), .Y (n_26326));
NAND2X1 g110414(.A (n_25677), .B (n_28808), .Y (n_26325));
NAND2X1 g110418(.A (n_26308), .B (n_22412), .Y (n_26324));
NAND2X1 g110420(.A (n_26306), .B (n_27999), .Y (n_26323));
NAND2X2 g110423(.A (n_25446), .B (n_20773), .Y (n_26322));
NAND2X1 g110437(.A (n_26320), .B (n_26665), .Y (n_26321));
NAND2X1 g110438(.A (n_26320), .B (n_33494), .Y (n_26319));
NAND2X1 g110439(.A (n_26320), .B (n_29445), .Y (n_26318));
NAND4X1 g110440(.A (n_18767), .B (n_24554), .C (n_24565), .D(n_24284), .Y (n_26317));
NAND2X1 g110445(.A (n_26290), .B (n_26315), .Y (n_26316));
NAND2X1 g110449(.A (n_26312), .B (n_10808), .Y (n_26314));
NAND2X1 g110450(.A (n_26312), .B (n_26528), .Y (n_26313));
NAND2X1 g110451(.A (n_26312), .B (n_26213), .Y (n_26311));
NAND2X1 g110452(.A (n_26312), .B (n_26288), .Y (n_26310));
NAND2X1 g110464(.A (n_26308), .B (n_23270), .Y (n_26309));
NAND2X1 g110467(.A (n_26306), .B (n_18384), .Y (n_26307));
NAND2X1 g110470(.A (n_26283), .B (n_25198), .Y (n_26305));
NAND4X1 g110481(.A (n_20479), .B (n_22072), .C (n_24562), .D(n_23290), .Y (n_26304));
NAND2X1 g110485(.A (n_26301), .B (n_27798), .Y (n_26303));
NAND2X1 g110486(.A (n_26301), .B (n_10808), .Y (n_26302));
NAND2X1 g110491(.A (n_26308), .B (n_32764), .Y (n_26300));
NAND2X1 g110493(.A (n_26306), .B (n_32664), .Y (n_26299));
NAND2X1 g110498(.A (n_26799), .B (n_28890), .Y (n_26298));
AND2X1 g110503(.A (n_26295), .B (n_26665), .Y (n_26297));
NAND2X1 g110504(.A (n_26295), .B (n_26662), .Y (n_26296));
NAND2X1 g110505(.A (n_26295), .B (n_26660), .Y (n_26294));
NAND2X1 g110506(.A (n_26292), .B (n_28890), .Y (n_26293));
NAND2X1 g110510(.A (n_26290), .B (n_27770), .Y (n_26291));
NAND2X1 g110513(.A (n_25688), .B (n_26288), .Y (n_26289));
INVX1 g110524(.A (n_26286), .Y (n_26287));
NAND2X1 g110532(.A (n_26306), .B (n_34688), .Y (n_26285));
NAND2X1 g110537(.A (n_26283), .B (n_23457), .Y (n_26284));
INVX1 g110538(.A (n_26807), .Y (n_26282));
NAND2X1 g110543(.A (n_26769), .B (n_29191), .Y (n_26281));
NAND4X1 g110544(.A (n_20466), .B (n_22071), .C (n_24559), .D(n_23288), .Y (n_26280));
NAND2X1 g110545(.A (n_26769), .B (n_30399), .Y (n_26279));
NAND2X1 g110565(.A (n_26283), .B (n_26637), .Y (n_26278));
NAND2X1 g110568(.A (n_25828), .B (n_18328), .Y (n_26277));
NAND2X1 g110573(.A (n_25448), .B (n_20244), .Y (n_32307));
NAND2X1 g110578(.A (n_25847), .B (n_26275), .Y (n_27283));
NAND2X1 g110580(.A (n_29430), .B (n_26273), .Y (n_26274));
NAND2X1 g110589(.A (n_26260), .B (n_18262), .Y (n_26272));
NAND2X1 g110591(.A (n_25339), .B (n_17782), .Y (n_26271));
INVX1 g110593(.A (n_26269), .Y (n_26270));
NAND2X1 g110595(.A (n_26259), .B (n_17968), .Y (n_26268));
NAND2X1 g110599(.A (n_26252), .B (n_18546), .Y (n_27260));
NOR2X1 g110611(.A (n_25395), .B (n_14952), .Y (n_26266));
NAND3X1 g110613(.A (n_25363), .B (n_24920), .C (n_19939), .Y(n_26265));
NAND2X1 g110627(.A (n_26244), .B (n_33738), .Y (n_26264));
NAND2X1 g110630(.A (n_26261), .B (n_8990), .Y (n_35608));
NAND2X1 g110632(.A (n_26261), .B (n_27522), .Y (n_26262));
NAND2X1 g110639(.A (n_26260), .B (n_35736), .Y (n_27306));
NAND2X1 g110640(.A (n_26259), .B (n_35816), .Y (n_27271));
NAND2X1 g110661(.A (n_26257), .B (n_29505), .Y (n_26258));
NAND2X1 g110662(.A (n_26257), .B (n_26255), .Y (n_26256));
INVX1 g110668(.A (n_25905), .Y (n_26254));
NAND2X1 g110672(.A (n_26252), .B (n_35744), .Y (n_26253));
NOR2X1 g110677(.A (n_25541), .B (n_10548), .Y (n_26251));
NAND2X1 g110698(.A (n_27100), .B (n_26249), .Y (n_26250));
NAND2X1 g110705(.A (n_26781), .B (n_28275), .Y (n_26248));
NAND2X1 g110706(.A (n_26781), .B (n_26528), .Y (n_26247));
NAND2X1 g110711(.A (n_26283), .B (n_27089), .Y (n_26246));
NAND2X1 g110728(.A (n_26244), .B (n_28158), .Y (n_26245));
NAND2X1 g110729(.A (n_26244), .B (n_28374), .Y (n_26243));
NAND2X1 g110738(.A (n_25043), .B (n_28364), .Y (n_26242));
NAND2X1 g110739(.A (n_25041), .B (n_28364), .Y (n_26241));
NAND2X1 g110743(.A (n_25039), .B (n_28364), .Y (n_26240));
NAND2X1 g110754(.A (n_26232), .B (n_26238), .Y (n_26239));
NAND2X1 g110765(.A (n_26252), .B (n_35578), .Y (n_27262));
NAND2X1 g110769(.A (n_26260), .B (n_26584), .Y (n_27275));
NAND2X1 g110772(.A (n_26259), .B (n_22021), .Y (n_27269));
NAND2X1 g110776(.A (n_26236), .B (n_25877), .Y (n_26582));
NAND2X1 g110780(.A (n_26252), .B (n_26234), .Y (n_26235));
NAND2X1 g110784(.A (n_26232), .B (n_29405), .Y (n_26233));
NAND2X1 g110785(.A (n_26232), .B (n_33738), .Y (n_26231));
INVX1 g110790(.A (n_25874), .Y (n_26578));
NAND2X1 g110793(.A (n_26260), .B (n_35515), .Y (n_26230));
NAND2X1 g110794(.A (n_26259), .B (n_35528), .Y (n_26229));
NAND2X1 g110797(.A (n_26236), .B (n_35540), .Y (n_26227));
NOR2X1 g110800(.A (n_24648), .B (n_25340), .Y (n_26225));
NAND4X1 g110804(.A (n_20504), .B (n_23632), .C (n_24517), .D(n_14381), .Y (n_26224));
NOR2X1 g110806(.A (n_10236), .B (n_25325), .Y (n_26223));
AOI21X1 g110826(.A0 (n_14941), .A1 (n_25723), .B0 (n_8927), .Y(n_26222));
AOI21X1 g110830(.A0 (n_14976), .A1 (n_25792), .B0 (n_8927), .Y(n_26221));
NAND4X1 g110831(.A (n_20409), .B (n_23630), .C (n_24514), .D(n_14826), .Y (n_26220));
NOR2X1 g110834(.A (n_9569), .B (n_25321), .Y (n_26219));
NOR2X1 g110837(.A (n_10222), .B (n_25322), .Y (n_26218));
NAND2X1 g110848(.A (n_25379), .B (n_29505), .Y (n_26217));
NAND2X1 g110861(.A (n_25405), .B (n_26216), .Y (n_27329));
NAND2X1 g110875(.A (n_25423), .B (n_24766), .Y (n_26215));
AOI21X1 g110879(.A0 (n_25767), .A1 (n_26213), .B0 (n_19753), .Y(n_26214));
NAND3X1 g110887(.A (n_23765), .B (n_24936), .C (n_23756), .Y(n_26212));
OAI21X1 g110897(.A0 (n_26205), .A1 (n_26210), .B0 (n_26209), .Y(n_28279));
NAND2X1 g110898(.A (n_25422), .B (n_26209), .Y (n_27338));
NAND2X1 g110899(.A (n_25421), .B (n_26208), .Y (n_27313));
CLKBUFX1 gbuf_d_373(.A(n_25320), .Y(d_out_373));
CLKBUFX1 gbuf_q_373(.A(q_in_373), .Y(P1_reg2[0]));
NAND2X1 g110917(.A (n_25416), .B (n_26207), .Y (n_27336));
OAI21X1 g110920(.A0 (n_26205), .A1 (n_26204), .B0 (n_24121), .Y(n_28270));
NAND2X1 g110921(.A (n_25415), .B (n_24121), .Y (n_27333));
NAND2X1 g110922(.A (n_25413), .B (n_26203), .Y (n_27304));
NAND2X1 g110936(.A (n_25410), .B (n_26202), .Y (n_27331));
OAI21X1 g110939(.A0 (n_26205), .A1 (n_32690), .B0 (n_26200), .Y(n_35201));
NAND2X1 g110941(.A (n_25408), .B (n_26200), .Y (n_27322));
NAND2X1 g110942(.A (n_25407), .B (n_26199), .Y (n_27297));
OAI21X1 g110956(.A0 (n_26205), .A1 (n_13579), .B0 (n_26197), .Y(n_35198));
NAND2X1 g110958(.A (n_25403), .B (n_26197), .Y (n_27319));
NAND2X1 g110959(.A (n_35920), .B (n_34690), .Y (n_27290));
INVX1 g110964(.A (n_26863), .Y (n_26195));
INVX1 g110969(.A (n_26832), .Y (n_26194));
NAND2X1 g110976(.A (n_25375), .B (n_26193), .Y (n_27341));
AOI21X1 g110983(.A0 (n_25738), .A1 (n_14672), .B0 (n_29725), .Y(n_26192));
AOI21X1 g110992(.A0 (n_25803), .A1 (n_26213), .B0 (n_19755), .Y(n_26190));
AOI21X1 g110993(.A0 (n_25798), .A1 (n_26213), .B0 (n_20293), .Y(n_26189));
AOI22X1 g110998(.A0 (n_25782), .A1 (n_26213), .B0 (n_9629), .B1(n_18416), .Y (n_26187));
AOI21X1 g111002(.A0 (n_25763), .A1 (n_26213), .B0 (n_20280), .Y(n_26186));
OAI21X1 g107932(.A0 (n_14647), .A1 (n_8945), .B0 (n_25319), .Y(n_26185));
AOI21X1 g111003(.A0 (n_25785), .A1 (n_26213), .B0 (n_19717), .Y(n_26184));
AOI21X1 g111004(.A0 (n_25805), .A1 (n_26213), .B0 (n_20298), .Y(n_26183));
AOI21X1 g111006(.A0 (n_26181), .A1 (n_26213), .B0 (n_21279), .Y(n_26182));
INVX1 g111007(.A (n_26812), .Y (n_26180));
INVX1 g111010(.A (n_26810), .Y (n_26178));
NOR2X1 g111016(.A (n_24337), .B (n_25318), .Y (n_26177));
NAND3X1 g111027(.A (n_24059), .B (n_25017), .C (n_24057), .Y(n_26176));
INVX1 g111035(.A (n_26827), .Y (n_26175));
NAND2X1 g111037(.A (n_25391), .B (n_19227), .Y (n_26174));
NAND2X1 g111042(.A (n_25371), .B (n_25925), .Y (n_27277));
NAND2X1 g111043(.A (n_25385), .B (n_28364), .Y (n_26173));
INVX1 g111046(.A (n_26842), .Y (n_26172));
OAI21X1 g111048(.A0 (n_24883), .A1 (n_10517), .B0 (n_19221), .Y(n_26171));
AND2X1 g111049(.A (n_25383), .B (n_19308), .Y (n_26170));
NAND2X1 g111058(.A (n_25427), .B (n_24782), .Y (n_26169));
NAND2X1 g111062(.A (n_25426), .B (n_24776), .Y (n_26168));
NAND2X1 g111066(.A (n_25425), .B (n_24770), .Y (n_26167));
NAND2X2 g111093(.A (n_25124), .B (n_25417), .Y (n_27300));
NAND3X1 g111123(.A (n_10593), .B (n_24858), .C (n_23699), .Y(n_26166));
NAND2X1 g111127(.A (n_26155), .B (n_28864), .Y (n_26165));
NOR2X1 g111131(.A (n_25269), .B (n_26748), .Y (n_26164));
NAND2X1 g111137(.A (n_26151), .B (n_26162), .Y (n_26163));
AND2X1 g111138(.A (n_26138), .B (n_26160), .Y (n_26161));
AND2X1 g111142(.A (n_26147), .B (n_34952), .Y (n_26159));
NAND2X1 g111146(.A (n_26157), .B (n_34694), .Y (n_26158));
NAND2X1 g111147(.A (n_26155), .B (n_28485), .Y (n_26156));
NAND2X1 g111149(.A (n_35359), .B (n_34694), .Y (n_26154));
NAND2X1 g111156(.A (n_26151), .B (n_28492), .Y (n_26152));
OAI21X1 g107994(.A0 (n_14432), .A1 (n_29968), .B0 (n_25304), .Y(n_26150));
AND2X1 g111163(.A (n_26147), .B (n_34693), .Y (n_26148));
NAND2X1 g111170(.A (n_26157), .B (n_26142), .Y (n_26146));
NAND2X1 g111171(.A (n_26155), .B (n_30197), .Y (n_26145));
NAND3X1 g111175(.A (n_23708), .B (n_24867), .C (n_23736), .Y(n_26144));
NAND2X1 g111180(.A (n_35359), .B (n_26142), .Y (n_26143));
NOR2X1 g111182(.A (n_24538), .B (n_25256), .Y (n_26141));
NAND2X1 g111187(.A (n_26151), .B (n_29090), .Y (n_26140));
NAND2X1 g111188(.A (n_26138), .B (n_26535), .Y (n_26139));
NAND2X1 g111195(.A (n_26147), .B (n_29604), .Y (n_26137));
NAND2X1 g111204(.A (n_26118), .B (n_18399), .Y (n_26136));
NAND2X1 g111212(.A (n_25308), .B (n_20085), .Y (n_32045));
NAND2X1 g111226(.A (n_26132), .B (n_24613), .Y (n_26133));
NAND2X1 g111241(.A (n_26129), .B (n_26106), .Y (n_26131));
NAND2X1 g111242(.A (n_26129), .B (n_26528), .Y (n_26130));
NAND2X1 g111243(.A (n_26129), .B (n_26213), .Y (n_26128));
INVX1 g111259(.A (n_26125), .Y (n_26126));
NOR2X1 g111275(.A (n_25589), .B (n_8678), .Y (n_26124));
NAND2X1 g111279(.A (n_26121), .B (n_28785), .Y (n_26123));
NAND2X1 g111282(.A (n_26121), .B (n_34753), .Y (n_26122));
OAI21X1 g108050(.A0 (n_14426), .A1 (n_28659), .B0 (n_25315), .Y(n_26120));
NAND2X1 g111299(.A (n_26118), .B (n_32685), .Y (n_26119));
NAND2X1 g111307(.A (n_29551), .B (n_24613), .Y (n_26117));
AND2X1 g111321(.A (n_26113), .B (n_28785), .Y (n_26115));
NAND2X1 g111322(.A (n_26112), .B (n_26113), .Y (n_26114));
NAND2X1 g111323(.A (n_26288), .B (n_26113), .Y (n_26111));
NAND2X1 g111325(.A (n_26113), .B (n_10808), .Y (n_26110));
NAND2X1 g111341(.A (n_26118), .B (n_25402), .Y (n_26109));
NAND3X1 g111353(.A (n_17268), .B (n_24857), .C (n_23686), .Y(n_26108));
NAND2X1 g111363(.A (n_26103), .B (n_26106), .Y (n_26107));
AOI21X1 g111402(.A0 (n_18596), .A1 (n_22139), .B0 (n_25311), .Y(n_26105));
NAND2X1 g111444(.A (n_26103), .B (n_26528), .Y (n_26104));
NAND2X1 g111445(.A (n_26103), .B (n_26213), .Y (n_26102));
NAND2X1 g111446(.A (n_26103), .B (n_26288), .Y (n_26101));
NAND3X1 g111479(.A (n_24844), .B (n_24836), .C (n_15151), .Y(n_26100));
NOR2X1 g111499(.A (n_24529), .B (n_25261), .Y (n_26099));
OAI21X1 g111508(.A0 (n_14340), .A1 (n_26801), .B0 (n_25301), .Y(n_26098));
NAND3X1 g111515(.A (n_9575), .B (n_24860), .C (n_23710), .Y(n_26097));
INVX1 g111579(.A (n_26719), .Y (n_26096));
NAND2X1 g111581(.A (n_25306), .B (n_25706), .Y (n_27668));
INVX1 g111588(.A (n_26717), .Y (n_26095));
NAND2X1 g111590(.A (n_25303), .B (n_25704), .Y (n_27665));
NAND2X1 g111594(.A (n_25299), .B (n_25702), .Y (n_27153));
NAND2X1 g111603(.A (n_25295), .B (n_25696), .Y (n_27162));
INVX1 g111608(.A (n_26663), .Y (n_26094));
INVX1 g111611(.A (n_26092), .Y (n_26091));
INVX1 g111623(.A (n_26711), .Y (n_26090));
NAND2X1 g111625(.A (n_25294), .B (n_25690), .Y (n_27676));
INVX1 g111645(.A (n_26639), .Y (n_26088));
NAND2X1 g111650(.A (n_25288), .B (n_25683), .Y (n_27116));
INVX1 g111654(.A (n_26703), .Y (n_26087));
INVX1 g111660(.A (n_26085), .Y (n_26084));
INVX1 g111663(.A (n_26082), .Y (n_26083));
NAND2X1 g111669(.A (n_25278), .B (n_25682), .Y (n_27105));
INVX1 g111670(.A (n_26607), .Y (n_26080));
NAND2X1 g111673(.A (n_25277), .B (n_25681), .Y (n_27094));
NAND2X1 g111678(.A (n_25675), .B (n_32022), .Y (n_27149));
INVX1 g111697(.A (n_26077), .Y (n_27660));
INVX1 g111716(.A (n_26620), .Y (n_26076));
OAI21X1 g111721(.A0 (n_14184), .A1 (n_8945), .B0 (n_25292), .Y(n_26075));
NAND2X1 g111745(.A (n_25279), .B (n_26074), .Y (n_27099));
OAI21X1 g111749(.A0 (n_25610), .A1 (n_35494), .B0 (n_25793), .Y(n_27658));
CLKBUFX1 gbuf_d_374(.A(n_25521), .Y(d_out_374));
CLKBUFX1 gbuf_q_374(.A(q_in_374), .Y(n_11135));
CLKBUFX1 gbuf_d_375(.A(n_25233), .Y(d_out_375));
CLKBUFX1 gbuf_q_375(.A(q_in_375), .Y(n_14317));
OAI21X1 g111795(.A0 (n_25285), .A1 (n_25284), .B0 (n_25286), .Y(n_27130));
NAND2X1 g111797(.A (n_24976), .B (n_25283), .Y (n_27127));
MX2X1 g111798(.A (n_21268), .B (n_21269), .S0 (n_24875), .Y(n_27125));
NAND2X2 g111814(.A (n_35876), .B (n_35877), .Y (n_35233));
INVX1 g111815(.A (n_26585), .Y (n_26073));
INVX1 g111821(.A (n_33812), .Y (n_26072));
AOI21X1 g108364(.A0 (n_14595), .A1 (n_14956), .B0 (n_25231), .Y(n_26071));
NAND3X1 g108397(.A (n_24143), .B (n_24787), .C (n_25121), .Y(n_26070));
NAND3X1 g108400(.A (n_24111), .B (n_24755), .C (n_25089), .Y(n_26069));
NOR2X1 g108434(.A (n_9930), .B (n_25237), .Y (n_26068));
NAND2X1 g112224(.A (n_25570), .B (n_28053), .Y (n_27018));
NAND2X1 g112291(.A (n_25249), .B (n_25271), .Y (n_27025));
NAND2X1 g112330(.A (n_25250), .B (n_23136), .Y (n_27031));
INVX1 g112332(.A (n_27053), .Y (n_26067));
OAI21X1 g112354(.A0 (n_24827), .A1 (n_32745), .B0 (n_25264), .Y(n_26063));
OAI21X1 g112393(.A0 (n_24828), .A1 (n_13817), .B0 (n_25260), .Y(n_27584));
INVX1 g112453(.A (n_26520), .Y (n_26062));
NAND4X1 g112815(.A (n_25236), .B (n_24137), .C (n_24173), .D(n_23892), .Y (n_27549));
NOR2X1 g108732(.A (n_25217), .B (n_25272), .Y (n_26061));
AOI21X1 g108784(.A0 (n_25183), .A1 (n_24418), .B0 (n_29769), .Y(n_26060));
AOI21X1 g108790(.A0 (n_25170), .A1 (n_24031), .B0 (n_8340), .Y(n_26059));
NAND2X1 g112965(.A (n_6751), .B (n_25239), .Y (n_26058));
NAND2X1 g112966(.A (n_6589), .B (n_25238), .Y (n_26057));
OAI21X1 g108805(.A0 (n_9748), .A1 (n_31129), .B0 (n_25544), .Y(n_26056));
AOI21X1 g108908(.A0 (n_25208), .A1 (n_34417), .B0 (n_8942), .Y(n_26055));
AOI21X1 g108913(.A0 (n_25206), .A1 (n_20072), .B0 (n_26052), .Y(n_26054));
AOI21X1 g108941(.A0 (n_25203), .A1 (n_13622), .B0 (n_26052), .Y(n_26053));
AOI21X1 g108947(.A0 (n_25200), .A1 (n_20173), .B0 (n_8942), .Y(n_26051));
INVX1 g109004(.A (n_35456), .Y (n_26050));
AOI21X1 g109053(.A0 (n_25185), .A1 (n_22097), .B0 (n_8942), .Y(n_26049));
OAI21X1 g109300(.A0 (n_25164), .A1 (n_24795), .B0 (n_33123), .Y(n_26048));
AOI21X1 g109596(.A0 (n_15182), .A1 (n_22821), .B0 (n_25181), .Y(n_26046));
AOI21X1 g109597(.A0 (n_15180), .A1 (n_22821), .B0 (n_25180), .Y(n_26045));
NAND2X1 g109629(.A (n_25154), .B (n_25122), .Y (n_35089));
NOR2X1 g109636(.A (n_24716), .B (n_25153), .Y (n_26043));
NAND2X1 g109658(.A (n_25168), .B (n_8641), .Y (n_26042));
NAND2X1 g109665(.A (n_25152), .B (n_8303), .Y (n_26040));
NOR2X1 g109669(.A (n_24712), .B (n_25150), .Y (n_26039));
NAND2X1 g109692(.A (n_25149), .B (n_8303), .Y (n_26038));
NAND2X1 g109722(.A (n_25175), .B (n_8641), .Y (n_26036));
NAND2X1 g109727(.A (n_25165), .B (n_8303), .Y (n_26034));
NAND2X1 g109739(.A (n_24703), .B (n_25195), .Y (n_26456));
NAND2X1 g109742(.A (n_25167), .B (n_9431), .Y (n_26033));
AND2X1 g109815(.A (n_26428), .B (n_27902), .Y (n_26032));
NAND2X1 g109831(.A (n_25166), .B (n_25942), .Y (n_26030));
NAND2X1 g109835(.A (n_26428), .B (n_8954), .Y (n_26029));
OAI21X1 g109837(.A0 (n_24796), .A1 (n_34336), .B0 (n_10375), .Y(n_26028));
NAND3X1 g109861(.A (n_24790), .B (n_21377), .C (n_24789), .Y(n_26027));
NAND3X1 g109863(.A (n_24758), .B (n_21334), .C (n_24757), .Y(n_26026));
NAND4X1 g109869(.A (n_22492), .B (n_22340), .C (n_24326), .D(n_22287), .Y (n_26025));
OAI21X1 g109876(.A0 (n_24732), .A1 (n_29681), .B0 (n_10453), .Y(n_26024));
OAI21X1 g109895(.A0 (n_24731), .A1 (n_27557), .B0 (n_10418), .Y(n_26023));
AOI21X1 g109922(.A0 (n_24925), .A1 (n_25515), .B0 (n_25172), .Y(n_26022));
AOI21X1 g109925(.A0 (n_14905), .A1 (n_25492), .B0 (n_8927), .Y(n_26021));
AOI21X1 g109938(.A0 (n_27100), .A1 (n_25499), .B0 (n_25162), .Y(n_26020));
AOI21X1 g109940(.A0 (n_26017), .A1 (n_27234), .B0 (n_19360), .Y(n_26018));
NAND2X1 g110052(.A (n_25196), .B (n_13170), .Y (n_26016));
NAND2X1 g110135(.A (n_25209), .B (n_28327), .Y (n_26015));
NAND2X1 g110137(.A (n_25202), .B (n_28325), .Y (n_26014));
NAND2X1 g110139(.A (n_25194), .B (n_28324), .Y (n_26013));
OAI21X1 g110172(.A0 (n_14734), .A1 (n_8614), .B0 (n_25197), .Y(n_26012));
AOI21X1 g110193(.A0 (n_25529), .A1 (n_29411), .B0 (n_20379), .Y(n_26011));
NAND3X1 g110273(.A (n_18010), .B (n_24396), .C (n_24646), .Y(n_26010));
NAND3X1 g110276(.A (n_25061), .B (n_24618), .C (n_20382), .Y(n_26009));
NAND4X1 g110278(.A (n_25062), .B (n_23402), .C (n_14846), .D(n_23396), .Y (n_26008));
NAND2X1 g110280(.A (n_33546), .B (n_25972), .Y (n_26007));
NAND2X1 g110292(.A (n_33546), .B (n_25951), .Y (n_26006));
AOI21X1 g110295(.A0 (n_24627), .A1 (n_23891), .B0 (n_8355), .Y(n_26005));
NAND2X1 g110296(.A (n_33546), .B (n_25916), .Y (n_26004));
NAND2X1 g110300(.A (n_25059), .B (n_26002), .Y (n_26003));
AOI21X1 g110304(.A0 (n_24586), .A1 (n_23868), .B0 (n_33125), .Y(n_26001));
NAND2X1 g110307(.A (n_27614), .B (n_25887), .Y (n_26000));
OAI21X1 g110312(.A0 (n_24489), .A1 (n_9626), .B0 (n_23185), .Y(n_25999));
NAND2X1 g110319(.A (n_34770), .B (n_25993), .Y (n_25998));
NAND2X1 g110333(.A (n_34770), .B (n_25989), .Y (n_25997));
NAND2X1 g110340(.A (n_25995), .B (n_34709), .Y (n_25996));
NAND2X1 g110349(.A (n_25993), .B (n_34709), .Y (n_25994));
AND2X1 g110358(.A (n_25991), .B (n_28926), .Y (n_25992));
NAND2X1 g110360(.A (n_25989), .B (n_25988), .Y (n_25990));
NAND2X1 g110362(.A (n_25986), .B (n_34709), .Y (n_25987));
NAND3X1 g110371(.A (n_24688), .B (n_24405), .C (n_24701), .Y(n_25985));
NAND2X1 g110373(.A (n_25995), .B (n_29199), .Y (n_25984));
NAND2X1 g110377(.A (n_25982), .B (n_28013), .Y (n_25983));
NAND2X1 g110385(.A (n_25993), .B (n_25980), .Y (n_25981));
NAND2X1 g110389(.A (n_25348), .B (n_33784), .Y (n_25979));
NAND2X1 g110396(.A (n_25991), .B (n_33785), .Y (n_25978));
NAND2X1 g110398(.A (n_25989), .B (n_25980), .Y (n_25977));
NAND3X1 g110401(.A (n_24630), .B (n_24400), .C (n_24697), .Y(n_25976));
NAND2X1 g110404(.A (n_25986), .B (n_29199), .Y (n_25975));
NAND2X1 g110421(.A (n_34521), .B (n_20774), .Y (n_25974));
NAND2X1 g110424(.A (n_25972), .B (n_24629), .Y (n_25973));
NAND2X2 g110425(.A (n_25025), .B (n_24490), .Y (n_25970));
NAND2X1 g110427(.A (n_25972), .B (n_25968), .Y (n_25969));
INVX1 g110428(.A (n_25966), .Y (n_25967));
NAND2X1 g110432(.A (n_26392), .B (n_30559), .Y (n_25965));
NAND2X1 g110446(.A (n_25957), .B (n_25554), .Y (n_25964));
NAND2X1 g110455(.A (n_25037), .B (n_26458), .Y (n_25962));
NAND2X1 g107710(.A (n_25953), .B (n_26676), .Y (n_25961));
NAND2X1 g110509(.A (n_25057), .B (n_12964), .Y (n_25960));
NAND2X1 g107718(.A (n_24880), .B (n_9431), .Y (n_25959));
NAND2X1 g110511(.A (n_25957), .B (n_25956), .Y (n_25958));
NAND2X1 g110521(.A (n_25034), .B (n_8641), .Y (n_25955));
NAND2X1 g110525(.A (n_25919), .B (n_25837), .Y (n_26286));
NAND2X1 g110539(.A (n_25923), .B (n_25838), .Y (n_26807));
NAND2X1 g107732(.A (n_25953), .B (n_25554), .Y (n_25954));
NAND2X1 g110548(.A (n_25951), .B (n_30180), .Y (n_25952));
NAND2X1 g110549(.A (n_25951), .B (n_26660), .Y (n_25949));
NAND2X1 g110552(.A (n_25957), .B (n_26637), .Y (n_25948));
NAND2X1 g110556(.A (n_25033), .B (n_9431), .Y (n_25947));
NAND2X1 g110571(.A (n_25097), .B (n_19731), .Y (n_25945));
NAND2X1 g110572(.A (n_25447), .B (n_20245), .Y (n_32308));
NAND2X1 g110574(.A (n_25032), .B (n_25942), .Y (n_25943));
NAND2X1 g107743(.A (n_24898), .B (n_9431), .Y (n_25941));
NAND2X1 g110585(.A (n_25846), .B (n_25394), .Y (n_26857));
NAND2X1 g110587(.A (n_25918), .B (n_18262), .Y (n_25940));
NAND2X1 g110588(.A (n_25906), .B (n_18262), .Y (n_26855));
NAND2X1 g110592(.A (n_25338), .B (n_18365), .Y (n_25937));
NAND2X1 g110594(.A (n_25903), .B (n_18546), .Y (n_26269));
NAND2X1 g110605(.A (n_25092), .B (n_19739), .Y (n_32196));
NAND3X1 g110615(.A (n_25064), .B (n_24607), .C (n_20377), .Y(n_25929));
NAND2X1 g110616(.A (n_27462), .B (n_25927), .Y (n_25928));
NAND4X1 g110618(.A (n_20894), .B (n_23405), .C (n_23426), .D(n_24277), .Y (n_25926));
NAND2X1 g110624(.A (n_25925), .B (n_25908), .Y (n_26846));
NAND2X1 g110625(.A (n_14714), .B (n_25923), .Y (n_25924));
NAND2X1 g107767(.A (n_25953), .B (n_35054), .Y (n_25922));
NAND2X1 g110636(.A (n_25839), .B (n_25921), .Y (n_26820));
NAND2X1 g110637(.A (n_15087), .B (n_25919), .Y (n_25920));
NAND2X1 g110638(.A (n_25918), .B (n_35736), .Y (n_26834));
NAND2X1 g110645(.A (n_25916), .B (n_24629), .Y (n_25917));
NAND2X1 g107773(.A (n_24876), .B (n_9431), .Y (n_25915));
NAND2X1 g110647(.A (n_25916), .B (n_25968), .Y (n_25914));
NAND2X1 g110648(.A (n_25910), .B (n_8990), .Y (n_25913));
NAND2X1 g110650(.A (n_25910), .B (n_27522), .Y (n_25911));
NAND2X1 g110657(.A (n_25908), .B (n_14674), .Y (n_25909));
NAND2X1 g110667(.A (n_25906), .B (n_35794), .Y (n_25907));
NOR2X1 g110669(.A (n_25021), .B (n_35766), .Y (n_25905));
NAND2X1 g110670(.A (n_25903), .B (n_35744), .Y (n_25904));
NOR2X1 g110676(.A (n_24826), .B (n_10873), .Y (n_25902));
NAND2X1 g110679(.A (n_25900), .B (n_29505), .Y (n_25901));
NAND2X1 g110680(.A (n_25900), .B (n_26255), .Y (n_25899));
NAND2X1 g107787(.A (n_25953), .B (n_23578), .Y (n_25898));
INVX1 g110690(.A (n_25894), .Y (n_25896));
INVX1 g110691(.A (n_25894), .Y (n_25895));
NAND2X1 g110693(.A (n_25038), .B (n_25942), .Y (n_25893));
NAND2X1 g110699(.A (n_25890), .B (n_28158), .Y (n_25891));
NAND2X1 g110700(.A (n_25890), .B (n_26238), .Y (n_25889));
NAND2X1 g110717(.A (n_27100), .B (n_25887), .Y (n_25888));
NAND2X1 g110720(.A (n_25029), .B (n_25942), .Y (n_25886));
NAND2X1 g110721(.A (n_25890), .B (n_8954), .Y (n_25885));
AOI21X1 g110735(.A0 (n_26978), .A1 (n_25433), .B0 (n_11326), .Y(n_25883));
NOR2X1 g110744(.A (n_26361), .B (n_25881), .Y (n_25882));
NOR2X1 g110745(.A (n_26368), .B (n_25881), .Y (n_25880));
NOR2X1 g110749(.A (n_26366), .B (n_25881), .Y (n_25879));
NAND2X1 g110761(.A (n_25906), .B (n_35540), .Y (n_26826));
NAND2X1 g110763(.A (n_25903), .B (n_35528), .Y (n_26868));
NAND2X1 g110767(.A (n_25918), .B (n_25877), .Y (n_26841));
NAND2X1 g110768(.A (n_25906), .B (n_25599), .Y (n_25876));
NAND2X1 g110771(.A (n_25903), .B (n_25072), .Y (n_25875));
NAND2X2 g110791(.A (n_25873), .B (n_25842), .Y (n_25874));
NAND2X1 g110792(.A (n_25918), .B (n_35457), .Y (n_25872));
OAI21X1 g110803(.A0 (n_14246), .A1 (n_26372), .B0 (n_25083), .Y(n_25871));
NAND2X1 g107844(.A (n_24873), .B (n_9431), .Y (n_25870));
OAI21X1 g110810(.A0 (n_24580), .A1 (n_25867), .B0 (n_14833), .Y(n_25868));
OAI21X1 g110811(.A0 (n_14433), .A1 (n_28659), .B0 (n_25115), .Y(n_25866));
AOI21X1 g110815(.A0 (n_24582), .A1 (n_8303), .B0 (n_15277), .Y(n_25865));
OAI21X1 g110820(.A0 (n_14927), .A1 (n_25862), .B0 (n_25112), .Y(n_25863));
AOI21X1 g110828(.A0 (n_14902), .A1 (n_25388), .B0 (n_8927), .Y(n_25861));
NOR2X1 g110833(.A (n_9556), .B (n_25027), .Y (n_25860));
NAND3X1 g110842(.A (n_9100), .B (n_24626), .C (n_19363), .Y(n_25859));
AOI21X1 g110844(.A0 (n_27100), .A1 (n_25835), .B0 (n_24421), .Y(n_25858));
NAND2X1 g110850(.A (n_25080), .B (n_29505), .Y (n_25857));
NAND2X1 g110857(.A (n_25107), .B (n_25856), .Y (n_26896));
AOI21X1 g110873(.A0 (n_22656), .A1 (n_25942), .B0 (n_25028), .Y(n_25855));
AOI21X1 g110888(.A0 (n_25437), .A1 (n_29061), .B0 (n_15136), .Y(n_32134));
AOI21X1 g110891(.A0 (n_25435), .A1 (n_34952), .B0 (n_15132), .Y(n_32149));
NAND2X1 g110911(.A (n_25118), .B (n_25353), .Y (n_26940));
NAND2X1 g110912(.A (n_25116), .B (n_25852), .Y (n_26898));
NAND2X1 g110952(.A (n_25110), .B (n_25350), .Y (n_26938));
AOI21X1 g110960(.A0 (n_24581), .A1 (n_25111), .B0 (n_15104), .Y(n_32275));
NAND2X1 g110965(.A (n_25102), .B (n_25342), .Y (n_26863));
NAND2X1 g110967(.A (n_25101), .B (n_25850), .Y (n_26894));
NAND2X1 g110970(.A (n_25099), .B (n_25336), .Y (n_26832));
NAND2X1 g110971(.A (n_25084), .B (n_25849), .Y (n_26892));
AOI21X1 g110982(.A0 (n_25386), .A1 (n_14570), .B0 (n_29725), .Y(n_25848));
OAI21X1 g111009(.A0 (n_24292), .A1 (n_13163), .B0 (n_25847), .Y(n_26812));
NAND2X1 g111011(.A (n_25095), .B (n_25846), .Y (n_26810));
OAI21X1 g111030(.A0 (n_24593), .A1 (n_25867), .B0 (n_14594), .Y(n_25845));
OAI21X1 g111031(.A0 (n_15056), .A1 (n_9458), .B0 (n_25103), .Y(n_25844));
OAI21X1 g111032(.A0 (n_24592), .A1 (n_25867), .B0 (n_15168), .Y(n_25843));
NAND2X1 g111036(.A (n_25074), .B (n_25842), .Y (n_26827));
AOI21X1 g111038(.A0 (n_8922), .A1 (n_25390), .B0 (n_19773), .Y(n_25841));
OAI21X1 g111047(.A0 (n_24566), .A1 (n_13739), .B0 (n_25839), .Y(n_26842));
NAND2X1 g111051(.A (n_25088), .B (n_25838), .Y (n_26837));
NAND2X1 g111052(.A (n_25086), .B (n_25837), .Y (n_26914));
AOI21X1 g111054(.A0 (n_25835), .A1 (n_29505), .B0 (n_18781), .Y(n_25836));
NAND3X1 g111056(.A (n_23444), .B (n_24694), .C (n_23440), .Y(n_25834));
OAI21X1 g111067(.A0 (n_14243), .A1 (n_9971), .B0 (n_25105), .Y(n_25833));
INVX1 g111069(.A (n_34514), .Y (n_25832));
AOI21X1 g111075(.A0 (n_25136), .A1 (n_34709), .B0 (n_25120), .Y(n_25830));
MX2X1 g111090(.A (n_21302), .B (n_18984), .S0 (n_24702), .Y(n_26881));
NAND2X2 g111092(.A (n_32078), .B (n_32079), .Y (n_26879));
INVX1 g111103(.A (n_25828), .Y (n_25829));
NAND3X1 g111108(.A (n_35638), .B (n_35639), .C (n_23030), .Y(n_25827));
NAND3X1 g111118(.A (n_17270), .B (n_24267), .C (n_24527), .Y(n_25826));
NAND3X1 g111122(.A (n_10596), .B (n_24268), .C (n_24535), .Y(n_25825));
OAI21X1 g111125(.A0 (n_9853), .A1 (n_25823), .B0 (n_24966), .Y(n_25824));
NAND2X1 g111136(.A (n_25814), .B (n_26162), .Y (n_25822));
NAND2X1 g111159(.A (n_25820), .B (n_29925), .Y (n_25821));
NOR2X1 g111164(.A (n_23727), .B (n_24882), .Y (n_25818));
NAND3X1 g111174(.A (n_24545), .B (n_24282), .C (n_24564), .Y(n_25817));
NOR2X1 g111178(.A (n_23421), .B (n_24881), .Y (n_35128));
NAND2X1 g111186(.A (n_25814), .B (n_26535), .Y (n_25815));
NOR2X1 g111192(.A (n_23416), .B (n_24879), .Y (n_25813));
NAND2X1 g111205(.A (n_25742), .B (n_14740), .Y (n_25812));
NAND4X1 g111207(.A (n_19947), .B (n_23602), .C (n_23618), .D(n_24165), .Y (n_25811));
NAND2X1 g111208(.A (n_25790), .B (n_18399), .Y (n_25810));
NAND2X1 g111211(.A (n_25307), .B (n_20086), .Y (n_32046));
NAND2X1 g111227(.A (n_18340), .B (n_25787), .Y (n_25808));
NAND2X1 g111233(.A (n_25769), .B (n_25554), .Y (n_25807));
NAND2X1 g111236(.A (n_25805), .B (n_26288), .Y (n_25806));
NAND2X1 g111237(.A (n_25803), .B (n_28785), .Y (n_32164));
NAND2X1 g111238(.A (n_25803), .B (n_24526), .Y (n_25802));
NAND2X1 g111239(.A (n_25803), .B (n_26288), .Y (n_25801));
NAND2X1 g111244(.A (n_25798), .B (n_28785), .Y (n_32162));
NAND2X1 g111245(.A (n_25798), .B (n_24526), .Y (n_25797));
NAND2X1 g111246(.A (n_25798), .B (n_26288), .Y (n_25795));
NAND4X1 g111251(.A (n_20484), .B (n_21613), .C (n_24172), .D(n_22936), .Y (n_25794));
NAND2X1 g111260(.A (n_25793), .B (n_25792), .Y (n_26125));
NAND2X1 g111263(.A (n_25790), .B (n_22792), .Y (n_25791));
NAND2X1 g111268(.A (n_24905), .B (n_25942), .Y (n_25789));
NAND2X1 g111270(.A (n_25787), .B (n_24446), .Y (n_25788));
NAND2X1 g111271(.A (n_25785), .B (n_26288), .Y (n_25786));
NAND2X1 g111276(.A (n_25270), .B (n_34753), .Y (n_25784));
NAND2X1 g111283(.A (n_25782), .B (n_28785), .Y (n_25783));
NAND2X1 g111284(.A (n_25782), .B (n_34753), .Y (n_25781));
NAND2X1 g111285(.A (n_25782), .B (n_26288), .Y (n_25780));
NAND2X1 g111288(.A (n_25777), .B (n_26528), .Y (n_25779));
NAND2X1 g111289(.A (n_25777), .B (n_25756), .Y (n_25778));
NAND2X1 g111290(.A (n_25777), .B (n_26288), .Y (n_25776));
NAND2X1 g111291(.A (n_25777), .B (n_10808), .Y (n_25775));
NAND2X1 g111293(.A (n_25751), .B (n_32815), .Y (n_25774));
NAND2X1 g111303(.A (n_25790), .B (n_32652), .Y (n_25772));
NAND2X1 g111308(.A (n_25787), .B (n_32685), .Y (n_25771));
NAND2X1 g111317(.A (n_25769), .B (n_27770), .Y (n_25770));
NAND2X1 g111318(.A (n_25767), .B (n_28785), .Y (n_25768));
NAND2X1 g111319(.A (n_25767), .B (n_34753), .Y (n_25766));
NAND2X1 g111320(.A (n_25767), .B (n_26288), .Y (n_25765));
NAND2X1 g111326(.A (n_25763), .B (n_28785), .Y (n_25764));
NAND2X1 g111327(.A (n_25763), .B (n_34753), .Y (n_25762));
NAND2X1 g111328(.A (n_25763), .B (n_26288), .Y (n_25761));
NAND2X1 g111333(.A (n_25757), .B (n_28785), .Y (n_25759));
NAND2X1 g111334(.A (n_25757), .B (n_25756), .Y (n_25758));
NAND2X1 g111335(.A (n_25757), .B (n_30063), .Y (n_25755));
NAND2X1 g111336(.A (n_25757), .B (n_10808), .Y (n_25753));
NAND2X1 g111337(.A (n_25751), .B (n_25404), .Y (n_25752));
NAND2X1 g111343(.A (n_25790), .B (n_25290), .Y (n_25750));
NOR2X1 g111351(.A (n_25748), .B (n_25275), .Y (n_25749));
NAND2X1 g111361(.A (n_25820), .B (n_26870), .Y (n_25747));
NAND2X1 g111366(.A (n_25769), .B (n_23578), .Y (n_25746));
NAND2X1 g111371(.A (n_24973), .B (n_19510), .Y (n_25745));
NAND2X1 g111373(.A (n_24900), .B (n_25942), .Y (n_25744));
NAND2X1 g111383(.A (n_24718), .B (n_25742), .Y (n_26626));
NAND2X1 g111388(.A (n_24911), .B (n_19244), .Y (n_32597));
NAND2X1 g111393(.A (n_34515), .B (n_18968), .Y (n_25740));
NAND2X1 g111396(.A (n_34860), .B (n_18346), .Y (n_25739));
NAND2X1 g111414(.A (n_25327), .B (n_25738), .Y (n_26594));
NAND2X1 g111415(.A (n_14685), .B (n_25736), .Y (n_25737));
NAND2X1 g111430(.A (n_25329), .B (n_25736), .Y (n_26588));
NAND2X1 g111437(.A (n_25769), .B (n_25734), .Y (n_25735));
NAND2X1 g111438(.A (n_25785), .B (n_28785), .Y (n_32139));
NAND2X1 g111440(.A (n_25785), .B (n_24526), .Y (n_25732));
NAND2X1 g111447(.A (n_25805), .B (n_28785), .Y (n_32114));
NAND2X1 g111448(.A (n_24899), .B (n_25942), .Y (n_25730));
NAND2X1 g111449(.A (n_25805), .B (n_24526), .Y (n_25729));
NAND2X1 g111454(.A (n_26181), .B (n_34753), .Y (n_25728));
NAND2X1 g111456(.A (n_26181), .B (n_26528), .Y (n_25727));
AOI21X1 g111463(.A0 (n_13978), .A1 (n_9436), .B0 (n_24886), .Y(n_25725));
NOR2X1 g111471(.A (n_24919), .B (n_24513), .Y (n_25724));
NAND2X1 g111487(.A (n_25723), .B (n_24086), .Y (n_26602));
NOR2X1 g111501(.A (n_21761), .B (n_25019), .Y (n_25722));
OAI21X1 g111510(.A0 (n_14406), .A1 (n_25563), .B0 (n_25005), .Y(n_25721));
NAND3X1 g111513(.A (n_9577), .B (n_24272), .C (n_24547), .Y(n_25720));
OAI21X1 g111521(.A0 (n_15011), .A1 (n_8614), .B0 (n_25001), .Y(n_25719));
NAND4X1 g111527(.A (n_20445), .B (n_23246), .C (n_24128), .D(n_21571), .Y (n_25717));
OAI21X1 g111535(.A0 (n_9862), .A1 (n_31680), .B0 (n_25018), .Y(n_25716));
NAND4X1 g111542(.A (n_20376), .B (n_23245), .C (n_24129), .D(n_21565), .Y (n_25715));
NAND2X1 g111548(.A (n_24999), .B (n_25355), .Y (n_26735));
NAND2X1 g111550(.A (n_24986), .B (n_34800), .Y (n_26653));
NAND2X1 g111556(.A (n_24994), .B (n_25713), .Y (n_27247));
OAI21X1 g111558(.A0 (n_26382), .A1 (n_24501), .B0 (n_24295), .Y(n_25712));
OAI21X1 g111559(.A0 (n_26382), .A1 (n_24502), .B0 (n_24575), .Y(n_25710));
NOR2X1 g111561(.A (n_24558), .B (n_25015), .Y (n_25709));
NAND2X1 g111568(.A (n_24945), .B (n_19870), .Y (n_25708));
OAI21X1 g111574(.A0 (n_24511), .A1 (n_8397), .B0 (n_10349), .Y(n_25707));
NAND2X1 g111577(.A (n_25009), .B (n_25055), .Y (n_26739));
NAND2X1 g111580(.A (n_25008), .B (n_25706), .Y (n_26719));
NAND2X1 g111587(.A (n_25007), .B (n_25705), .Y (n_27253));
NAND2X1 g111589(.A (n_25006), .B (n_25704), .Y (n_26717));
INVX1 g111591(.A (n_26333), .Y (n_25703));
NAND2X1 g111595(.A (n_25004), .B (n_25702), .Y (n_26695));
INVX1 g111596(.A (n_26301), .Y (n_25701));
INVX1 g111599(.A (n_25698), .Y (n_25699));
OAI21X1 g111602(.A0 (n_24493), .A1 (n_32748), .B0 (n_25696), .Y(n_26672));
NAND2X1 g111609(.A (n_24997), .B (n_25693), .Y (n_26663));
OAI21X1 g111612(.A0 (n_24498), .A1 (n_25694), .B0 (n_25693), .Y(n_26092));
NAND2X1 g111613(.A (n_24995), .B (n_25345), .Y (n_26732));
INVX1 g111615(.A (n_26295), .Y (n_25692));
INVX1 g111621(.A (n_26292), .Y (n_25691));
NAND2X1 g111624(.A (n_24992), .B (n_25690), .Y (n_26711));
NAND2X1 g111626(.A (n_24988), .B (n_25689), .Y (n_26730));
INVX1 g111628(.A (n_25688), .Y (n_26657));
INVX1 g111630(.A (n_25686), .Y (n_25687));
NAND2X1 g111646(.A (n_24982), .B (n_25684), .Y (n_26639));
NAND2X1 g111648(.A (n_24981), .B (n_25683), .Y (n_26728));
NAND2X1 g111651(.A (n_24937), .B (n_25682), .Y (n_26726));
NAND2X1 g111655(.A (n_24934), .B (n_25681), .Y (n_26703));
OAI21X1 g111661(.A0 (n_24499), .A1 (n_24312), .B0 (n_24721), .Y(n_26085));
NAND2X1 g111665(.A (n_24938), .B (n_25680), .Y (n_26082));
OAI21X1 g111666(.A0 (n_25305), .A1 (n_24312), .B0 (n_25680), .Y(n_27235));
NAND2X1 g111671(.A (n_24935), .B (n_25679), .Y (n_26607));
INVX1 g111674(.A (n_25677), .Y (n_25678));
NAND2X1 g111679(.A (n_24923), .B (n_25675), .Y (n_26596));
INVX1 g111693(.A (n_25673), .Y (n_27193));
NAND2X1 g111699(.A (n_24964), .B (n_25396), .Y (n_26077));
NAND2X1 g111717(.A (n_24913), .B (n_24760), .Y (n_26620));
OAI21X1 g111726(.A0 (n_14592), .A1 (n_8614), .B0 (n_24983), .Y(n_25672));
INVX1 g111737(.A (n_26261), .Y (n_25671));
NAND2X1 g111743(.A (n_24941), .B (n_24785), .Y (n_26615));
NAND2X1 g111751(.A (n_25010), .B (n_19362), .Y (n_25670));
OAI21X1 g111769(.A0 (n_24516), .A1 (n_31470), .B0 (n_7105), .Y(n_25669));
OAI21X1 g111770(.A0 (n_24512), .A1 (n_31470), .B0 (n_6913), .Y(n_25668));
CLKBUFX1 gbuf_d_376(.A(n_25023), .Y(d_out_376));
CLKBUFX1 gbuf_q_376(.A(q_in_376), .Y(n_9590));
CLKBUFX1 gbuf_d_377(.A(n_25022), .Y(d_out_377));
CLKBUFX1 gbuf_q_377(.A(q_in_377), .Y(n_9549));
OAI21X1 g111779(.A0 (n_24604), .A1 (n_27662), .B0 (n_24951), .Y(n_25667));
OAI21X1 g111780(.A0 (n_24917), .A1 (n_27662), .B0 (n_24949), .Y(n_25666));
NAND2X1 g111785(.A (n_25014), .B (n_24692), .Y (n_26690));
INVX1 g111792(.A (n_26290), .Y (n_25664));
OAI21X1 g111796(.A0 (n_24978), .A1 (n_24977), .B0 (n_24979), .Y(n_26655));
NAND2X1 g111800(.A (n_24971), .B (n_24642), .Y (n_26677));
NAND2X1 g111801(.A (n_24641), .B (n_24970), .Y (n_26648));
MX2X1 g111802(.A (n_17780), .B (n_19651), .S0 (n_24500), .Y(n_26643));
INVX1 g111805(.A (n_25662), .Y (n_26629));
NAND2X2 g111816(.A (n_32243), .B (n_32244), .Y (n_26585));
INVX1 g111818(.A (n_26236), .Y (n_25661));
NAND2X2 g111820(.A (n_24633), .B (n_24955), .Y (n_26609));
NAND2X1 g111849(.A (n_33546), .B (n_25626), .Y (n_25660));
NAND2X1 g111855(.A (n_33546), .B (n_25621), .Y (n_25659));
NAND2X1 g111860(.A (n_33546), .B (n_25612), .Y (n_25658));
NAND2X1 g111864(.A (n_33546), .B (n_25608), .Y (n_25657));
NAND2X1 g111870(.A (n_28597), .B (n_25637), .Y (n_25656));
NAND2X1 g111871(.A (n_28597), .B (n_25634), .Y (n_25655));
NAND2X1 g111873(.A (n_29065), .B (n_25632), .Y (n_25654));
NAND2X1 g111874(.A (n_29065), .B (n_25630), .Y (n_25653));
NAND2X1 g111875(.A (n_34770), .B (n_25645), .Y (n_25652));
NAND2X1 g111876(.A (n_34770), .B (n_25643), .Y (n_25651));
NAND2X1 g111878(.A (n_25641), .B (n_25988), .Y (n_25649));
NAND2X1 g111879(.A (n_25647), .B (n_28926), .Y (n_25648));
NAND2X1 g111888(.A (n_25645), .B (n_25988), .Y (n_25646));
NAND2X1 g111889(.A (n_25643), .B (n_25988), .Y (n_25644));
NAND2X1 g111892(.A (n_25641), .B (n_29455), .Y (n_25642));
NAND2X1 g111893(.A (n_25647), .B (n_25980), .Y (n_25640));
NOR2X1 g111897(.A (n_23592), .B (n_24835), .Y (n_35125));
NAND2X1 g111899(.A (n_25637), .B (n_25636), .Y (n_25638));
NAND2X1 g111900(.A (n_25634), .B (n_29455), .Y (n_25635));
NAND2X1 g111902(.A (n_25632), .B (n_28915), .Y (n_25633));
NAND2X1 g111903(.A (n_25630), .B (n_33784), .Y (n_25631));
NAND2X1 g111907(.A (n_25645), .B (n_29455), .Y (n_25629));
NAND2X1 g111908(.A (n_25643), .B (n_28013), .Y (n_25628));
NAND2X1 g111936(.A (n_25626), .B (n_30559), .Y (n_25627));
NAND2X1 g111937(.A (n_25626), .B (n_30180), .Y (n_25625));
NAND2X1 g111951(.A (n_25617), .B (n_25554), .Y (n_25624));
NAND4X1 g108362(.A (n_14851), .B (n_23460), .C (n_24234), .D(n_23419), .Y (n_25623));
AND2X1 g111990(.A (n_25621), .B (n_27993), .Y (n_25622));
NAND2X1 g111992(.A (n_25621), .B (n_30559), .Y (n_25620));
NAND4X1 g108363(.A (n_14401), .B (n_22850), .C (n_24226), .D(n_23414), .Y (n_25619));
NAND2X1 g112008(.A (n_25617), .B (n_23192), .Y (n_25618));
NAND2X1 g112030(.A (n_24497), .B (n_13274), .Y (n_25616));
NAND2X1 g112047(.A (n_25617), .B (n_18137), .Y (n_25615));
AND2X1 g112053(.A (n_25612), .B (n_27993), .Y (n_25613));
NAND2X1 g112054(.A (n_25612), .B (n_26660), .Y (n_25611));
NAND2X1 g112089(.A (n_25602), .B (n_24965), .Y (n_26508));
NAND2X1 g112092(.A (n_24494), .B (n_17968), .Y (n_26513));
OR2X1 g112126(.A (n_25610), .B (n_35771), .Y (n_26510));
NAND2X1 g112130(.A (n_25608), .B (n_30559), .Y (n_25609));
NAND2X1 g112131(.A (n_25608), .B (n_30180), .Y (n_25607));
NAND2X1 g112156(.A (n_25617), .B (n_25605), .Y (n_25606));
OAI21X1 g108421(.A0 (n_8704), .A1 (n_31122), .B0 (n_24831), .Y(n_25604));
NAND2X1 g112171(.A (n_25602), .B (n_35736), .Y (n_25603));
NAND2X1 g112214(.A (n_25602), .B (n_35457), .Y (n_26505));
NAND2X1 g112221(.A (n_25602), .B (n_25599), .Y (n_25600));
NAND2X1 g112225(.A (n_24494), .B (n_25596), .Y (n_25598));
NOR2X1 g112235(.A (n_23582), .B (n_24838), .Y (n_25595));
NAND3X1 g108450(.A (n_25593), .B (n_25234), .C (n_23874), .Y(n_25594));
INVX1 g112292(.A (n_26138), .Y (n_25592));
NAND2X1 g112323(.A (n_24853), .B (n_22839), .Y (n_26541));
INVX1 g112324(.A (n_26129), .Y (n_25591));
NAND2X1 g112333(.A (n_24852), .B (n_25590), .Y (n_27053));
INVX1 g112343(.A (n_26121), .Y (n_26522));
INVX1 g112350(.A (n_25266), .Y (n_26064));
INVX1 g112356(.A (n_25586), .Y (n_25587));
NAND2X1 g112378(.A (n_24864), .B (n_23731), .Y (n_25584));
NAND2X1 g112388(.A (n_24847), .B (n_22836), .Y (n_26538));
NAND2X1 g112442(.A (n_24866), .B (n_23733), .Y (n_25583));
NAND2X1 g112454(.A (n_24845), .B (n_24518), .Y (n_26520));
INVX1 g112455(.A (n_26118), .Y (n_25582));
NAND2X1 g112607(.A (n_25579), .B (n_18918), .Y (n_25581));
NAND2X1 g112667(.A (n_25579), .B (n_24984), .Y (n_25580));
NAND2X1 g112685(.A (n_25579), .B (n_21627), .Y (n_25578));
AOI21X1 g111774(.A0 (n_16615), .A1 (n_17958), .B0 (n_25016), .Y(n_26641));
NAND4X1 g112799(.A (n_24830), .B (n_24177), .C (n_23625), .D(n_23296), .Y (n_27021));
NAND4X1 g108729(.A (n_24825), .B (n_10240), .C (n_23604), .D(n_24161), .Y (n_25577));
OAI21X1 g112959(.A0 (n_24487), .A1 (n_31605), .B0 (n_6665), .Y(n_25576));
OAI21X1 g112961(.A0 (n_24486), .A1 (n_31744), .B0 (n_6502), .Y(n_25575));
OAI21X1 g112967(.A0 (n_24481), .A1 (n_31273), .B0 (n_6648), .Y(n_25574));
NAND3X1 g108792(.A (n_18573), .B (n_20387), .C (n_24821), .Y(n_25573));
NAND3X1 g108793(.A (n_19128), .B (n_20856), .C (n_24819), .Y(n_25572));
INVX1 g113012(.A (n_25570), .Y (n_25571));
OAI21X1 g108960(.A0 (n_24823), .A1 (n_23735), .B0 (n_31064), .Y(n_25569));
NAND3X1 g109156(.A (n_19107), .B (n_20944), .C (n_24802), .Y(n_25568));
AOI21X1 g109212(.A0 (n_22087), .A1 (n_25082), .B0 (n_24887), .Y(n_25567));
OAI21X1 g109238(.A0 (n_14738), .A1 (n_25563), .B0 (n_25226), .Y(n_25566));
OAI21X1 g109258(.A0 (n_24799), .A1 (n_23692), .B0 (n_30360), .Y(n_25565));
OAI21X1 g109297(.A0 (n_14737), .A1 (n_25563), .B0 (n_25219), .Y(n_25564));
OAI21X1 g109320(.A0 (n_15293), .A1 (n_8614), .B0 (n_25225), .Y(n_25562));
OAI21X1 g109321(.A0 (n_15291), .A1 (n_15026), .B0 (n_25224), .Y(n_25561));
OAI21X1 g109395(.A0 (n_14732), .A1 (n_25368), .B0 (n_25223), .Y(n_25560));
NAND4X1 g109544(.A (n_24422), .B (n_24077), .C (n_24072), .D(n_21274), .Y (n_25559));
NAND4X1 g109598(.A (n_35635), .B (n_35636), .C (n_24052), .D(n_24053), .Y (n_25558));
NAND2X1 g109616(.A (n_25555), .B (n_25207), .Y (n_25557));
NAND2X1 g109673(.A (n_25555), .B (n_25554), .Y (n_25556));
NAND2X1 g109767(.A (n_25555), .B (n_13274), .Y (n_25553));
OAI21X1 g107401(.A0 (n_14468), .A1 (n_14916), .B0 (n_24812), .Y(n_25552));
OAI21X1 g107417(.A0 (n_14467), .A1 (n_26372), .B0 (n_24810), .Y(n_25550));
NAND4X1 g109860(.A (n_24434), .B (n_24078), .C (n_24074), .D(n_21276), .Y (n_25548));
AOI22X1 g109877(.A0 (n_14963), .A1 (n_25229), .B0 (n_24425), .B1(n_25228), .Y (n_25547));
OAI21X1 g107444(.A0 (n_14463), .A1 (n_26372), .B0 (n_24798), .Y(n_25546));
NOR2X1 g109902(.A (n_24815), .B (n_15341), .Y (n_25545));
OAI21X1 g109905(.A0 (n_24431), .A1 (n_24436), .B0 (n_34731), .Y(n_25544));
OAI21X1 g109914(.A0 (n_24429), .A1 (n_24435), .B0 (n_27485), .Y(n_25543));
OAI21X1 g111772(.A0 (n_18575), .A1 (n_25540), .B0 (n_24599), .Y(n_25541));
OAI21X1 g107494(.A0 (n_14460), .A1 (n_9971), .B0 (n_24811), .Y(n_25539));
AOI21X1 g109987(.A0 (n_25205), .A1 (n_32777), .B0 (n_19494), .Y(n_25538));
NAND4X1 g109988(.A (n_15183), .B (n_22828), .C (n_24048), .D(n_24049), .Y (n_25537));
NOR2X1 g110166(.A (n_14531), .B (n_24817), .Y (n_25536));
NOR2X1 g110168(.A (n_14524), .B (n_24816), .Y (n_25535));
AOI21X1 g110171(.A0 (n_14496), .A1 (n_8313), .B0 (n_24814), .Y(n_25534));
NOR2X1 g110308(.A (n_23113), .B (n_24773), .Y (n_25533));
AOI21X1 g110310(.A0 (n_24868), .A1 (n_29027), .B0 (n_22841), .Y(n_25532));
NAND2X1 g110315(.A (n_24725), .B (n_23346), .Y (n_25531));
NAND2X1 g110413(.A (n_25529), .B (n_8954), .Y (n_25530));
NAND2X1 g110426(.A (n_25024), .B (n_19519), .Y (n_25528));
NAND3X1 g110429(.A (n_32039), .B (n_21790), .C (n_32040), .Y(n_25966));
NOR2X1 g110431(.A (n_23115), .B (n_24728), .Y (n_25527));
NAND2X1 g110442(.A (n_25529), .B (n_28158), .Y (n_25526));
NAND2X1 g110472(.A (n_24715), .B (n_25082), .Y (n_25525));
NOR2X1 g110473(.A (n_23114), .B (n_24727), .Y (n_25523));
NAND2X1 g110479(.A (n_25513), .B (n_17713), .Y (n_25522));
NAND2X1 g110497(.A (n_24724), .B (n_12816), .Y (n_25521));
OAI21X1 g110540(.A0 (n_24409), .A1 (n_23120), .B0 (n_27485), .Y(n_25520));
NAND2X1 g110541(.A (n_24722), .B (n_25942), .Y (n_25519));
NAND2X1 g110570(.A (n_25096), .B (n_21389), .Y (n_25517));
NAND2X1 g110575(.A (n_27462), .B (n_25515), .Y (n_25516));
NAND2X1 g110590(.A (n_25475), .B (n_18262), .Y (n_26400));
NAND2X1 g110598(.A (n_25513), .B (n_17340), .Y (n_25514));
NAND2X1 g110604(.A (n_34493), .B (n_21393), .Y (n_32197));
NAND3X1 g110612(.A (n_24015), .B (n_24296), .C (n_15184), .Y(n_25508));
NAND2X1 g110617(.A (n_25504), .B (n_8990), .Y (n_25507));
NAND2X1 g110619(.A (n_25489), .B (n_33738), .Y (n_25506));
NAND2X1 g110620(.A (n_25504), .B (n_27522), .Y (n_25505));
NAND2X1 g110622(.A (n_25486), .B (n_33738), .Y (n_25503));
NAND2X1 g110629(.A (n_28874), .B (n_25493), .Y (n_25502));
NAND2X1 g110649(.A (n_25483), .B (n_33738), .Y (n_25501));
NAND2X1 g110651(.A (n_25499), .B (n_29505), .Y (n_25500));
NAND2X1 g110652(.A (n_25499), .B (n_26255), .Y (n_25498));
NAND2X1 g110653(.A (n_26017), .B (n_26660), .Y (n_25497));
NAND2X1 g110656(.A (n_26017), .B (n_26611), .Y (n_25496));
NOR2X1 g110678(.A (n_24704), .B (n_10577), .Y (n_25495));
NAND2X1 g110683(.A (n_27100), .B (n_25493), .Y (n_25494));
NAND2X1 g110692(.A (n_25148), .B (n_25492), .Y (n_25894));
NAND2X1 g110697(.A (n_25529), .B (n_26238), .Y (n_25491));
NAND2X1 g110724(.A (n_25489), .B (n_28158), .Y (n_25490));
NAND2X1 g110725(.A (n_25489), .B (n_28374), .Y (n_25488));
NAND2X1 g110726(.A (n_25486), .B (n_28158), .Y (n_25487));
NAND2X1 g110727(.A (n_25486), .B (n_28374), .Y (n_25485));
NAND2X1 g110733(.A (n_25483), .B (n_28158), .Y (n_25484));
NAND2X1 g110734(.A (n_25483), .B (n_28374), .Y (n_25482));
NAND3X1 g110736(.A (n_32239), .B (n_32240), .C (n_22575), .Y(n_25481));
NAND2X1 g110750(.A (n_25472), .B (n_26238), .Y (n_25480));
NAND2X1 g110751(.A (n_25469), .B (n_30636), .Y (n_25479));
NAND2X1 g110753(.A (n_25476), .B (n_30636), .Y (n_25478));
NAND2X1 g110760(.A (n_25476), .B (n_33738), .Y (n_25477));
NAND2X1 g110762(.A (n_25475), .B (n_35508), .Y (n_26397));
NAND2X1 g110770(.A (n_25475), .B (n_28053), .Y (n_25474));
NAND2X1 g110781(.A (n_25472), .B (n_29405), .Y (n_25473));
NAND2X1 g110782(.A (n_25472), .B (n_33738), .Y (n_25471));
NAND2X1 g110783(.A (n_25469), .B (n_29405), .Y (n_25470));
NAND2X1 g110788(.A (n_25476), .B (n_29405), .Y (n_25467));
NAND2X1 g110796(.A (n_25469), .B (n_33738), .Y (n_25466));
NAND3X1 g110798(.A (n_32881), .B (n_32882), .C (n_22208), .Y(n_26416));
NOR2X1 g110835(.A (n_9547), .B (n_24706), .Y (n_25465));
AOI21X1 g110836(.A0 (n_14807), .A1 (n_25081), .B0 (n_8927), .Y(n_25464));
CLKBUFX1 gbuf_d_378(.A(n_24705), .Y(d_out_378));
CLKBUFX1 gbuf_q_378(.A(q_in_378), .Y(n_10563));
NAND3X1 g110841(.A (n_9086), .B (n_24347), .C (n_19857), .Y(n_25463));
NAND2X1 g110845(.A (n_24746), .B (n_29505), .Y (n_25462));
NAND3X1 g110881(.A (n_19295), .B (n_24030), .C (n_24335), .Y(n_25461));
NAND3X1 g110882(.A (n_19291), .B (n_24029), .C (n_24334), .Y(n_25460));
AOI21X1 g110889(.A0 (n_25142), .A1 (n_34952), .B0 (n_15194), .Y(n_32163));
AOI21X1 g110892(.A0 (n_25138), .A1 (n_29061), .B0 (n_15192), .Y(n_32138));
OAI21X1 g110894(.A0 (n_14222), .A1 (n_33713), .B0 (n_24744), .Y(n_25457));
OAI21X1 g107925(.A0 (n_14663), .A1 (n_26372), .B0 (n_24708), .Y(n_25456));
NAND4X1 g110986(.A (n_35885), .B (n_35886), .C (n_23065), .D(n_23064), .Y (n_25455));
NAND2X1 g111020(.A (n_24738), .B (n_15185), .Y (n_25454));
NAND2X1 g111039(.A (n_24761), .B (n_28364), .Y (n_25453));
NAND2X1 g111040(.A (n_24780), .B (n_26548), .Y (n_25452));
NAND2X1 g111050(.A (n_24749), .B (n_26548), .Y (n_25451));
AOI21X1 g111083(.A0 (n_25127), .A1 (n_34709), .B0 (n_24754), .Y(n_25450));
OAI21X1 g107964(.A0 (n_24107), .A1 (n_8940), .B0 (n_15075), .Y(n_25449));
NAND3X1 g111104(.A (n_21307), .B (n_24220), .C (n_23312), .Y(n_25828));
INVX1 g111109(.A (n_25447), .Y (n_25448));
INVX1 g111115(.A (n_34521), .Y (n_25446));
NOR2X1 g111117(.A (n_18403), .B (n_24585), .Y (n_25444));
NAND3X1 g111119(.A (n_17489), .B (n_24245), .C (n_18191), .Y(n_25443));
NOR2X1 g111121(.A (n_10597), .B (n_24572), .Y (n_25442));
NAND2X1 g111134(.A (n_25431), .B (n_28864), .Y (n_25441));
NAND2X1 g111140(.A (n_25429), .B (n_26162), .Y (n_25439));
NAND2X1 g111143(.A (n_25437), .B (n_34694), .Y (n_25438));
NAND2X1 g111150(.A (n_25435), .B (n_34694), .Y (n_25436));
NAND2X1 g111153(.A (n_25433), .B (n_29925), .Y (n_25434));
NAND2X1 g111154(.A (n_25431), .B (n_28492), .Y (n_25432));
NAND2X1 g111158(.A (n_25429), .B (n_28492), .Y (n_25430));
NAND2X1 g111167(.A (n_25437), .B (n_25424), .Y (n_25427));
NAND2X1 g111176(.A (n_25435), .B (n_26142), .Y (n_25426));
NAND2X1 g111184(.A (n_25431), .B (n_25424), .Y (n_25425));
NAND2X1 g111191(.A (n_25429), .B (n_29090), .Y (n_25423));
NAND2X1 g111200(.A (n_25414), .B (n_25374), .Y (n_25422));
NAND2X1 g111201(.A (n_25412), .B (n_17719), .Y (n_25421));
NAND2X1 g111202(.A (n_24584), .B (n_8303), .Y (n_25419));
NAND2X1 g111215(.A (n_24684), .B (n_20784), .Y (n_25417));
NAND2X1 g111253(.A (n_25409), .B (n_22406), .Y (n_25416));
NAND2X1 g111254(.A (n_25414), .B (n_22406), .Y (n_25415));
NAND2X1 g111256(.A (n_25412), .B (n_22406), .Y (n_25413));
NAND2X1 g111257(.A (n_24583), .B (n_8303), .Y (n_25411));
NAND2X1 g111294(.A (n_25409), .B (n_32794), .Y (n_25410));
NAND2X1 g111295(.A (n_25414), .B (n_32664), .Y (n_25408));
NAND2X1 g111296(.A (n_25412), .B (n_32777), .Y (n_25407));
NAND2X1 g111301(.A (n_25433), .B (n_26870), .Y (n_25406));
NAND2X1 g111338(.A (n_25409), .B (n_25404), .Y (n_25405));
NAND2X1 g111339(.A (n_25414), .B (n_25402), .Y (n_25403));
NAND2X1 g111340(.A (n_25412), .B (n_25404), .Y (n_35920));
NAND2X1 g111357(.A (n_25384), .B (n_25400), .Y (n_26232));
NAND2X1 g111372(.A (n_24972), .B (n_19511), .Y (n_25399));
NAND2X1 g111384(.A (n_24291), .B (n_14439), .Y (n_26275));
NAND2X1 g111386(.A (n_34834), .B (n_21388), .Y (n_32596));
NAND2X1 g111387(.A (n_25396), .B (n_25378), .Y (n_26273));
INVX1 g111391(.A (n_25394), .Y (n_25395));
NAND2X1 g111394(.A (n_24901), .B (n_19508), .Y (n_25393));
NAND2X1 g111397(.A (n_24960), .B (n_18347), .Y (n_25392));
NAND2X1 g111403(.A (n_27632), .B (n_25390), .Y (n_25391));
NAND2X1 g111404(.A (n_29695), .B (n_25390), .Y (n_25389));
NAND2X1 g111409(.A (n_25388), .B (n_25035), .Y (n_26249));
NAND2X1 g111412(.A (n_25387), .B (n_25386), .Y (n_26244));
NAND2X1 g111413(.A (n_14362), .B (n_25384), .Y (n_25385));
NAND2X1 g111424(.A (n_25381), .B (n_27109), .Y (n_25383));
NAND2X1 g111425(.A (n_24925), .B (n_25381), .Y (n_25382));
NAND2X1 g111439(.A (n_25835), .B (n_26132), .Y (n_25380));
NAND2X1 g111443(.A (n_25378), .B (n_14920), .Y (n_25379));
OAI21X1 g111455(.A0 (n_23322), .A1 (n_25376), .B0 (n_24576), .Y(n_25377));
NAND2X1 g111462(.A (n_25409), .B (n_25374), .Y (n_25375));
NAND3X1 g111464(.A (n_32568), .B (n_32569), .C (n_22858), .Y(n_25373));
NAND4X1 g111473(.A (n_24693), .B (n_23300), .C (n_22372), .D(n_22377), .Y (n_25372));
NAND2X1 g111491(.A (n_24291), .B (n_25596), .Y (n_25371));
OAI21X1 g111505(.A0 (n_14189), .A1 (n_25368), .B0 (n_24680), .Y(n_25369));
NOR2X1 g111506(.A (n_9126), .B (n_24574), .Y (n_25367));
NOR2X1 g111512(.A (n_9087), .B (n_24573), .Y (n_25366));
OAI21X1 g111520(.A0 (n_14869), .A1 (n_8614), .B0 (n_24666), .Y(n_25365));
OAI21X1 g111526(.A0 (n_14188), .A1 (n_25563), .B0 (n_24649), .Y(n_25364));
AOI21X1 g111530(.A0 (n_24925), .A1 (n_24950), .B0 (n_24590), .Y(n_25363));
AOI21X1 g111531(.A0 (n_27100), .A1 (n_24947), .B0 (n_24589), .Y(n_25362));
INVX1 g111533(.A (n_25063), .Y (n_25361));
OAI21X1 g111537(.A0 (n_9875), .A1 (n_25823), .B0 (n_24696), .Y(n_25360));
AOI21X1 g111539(.A0 (n_27100), .A1 (n_24932), .B0 (n_24000), .Y(n_25359));
AOI21X1 g111540(.A0 (n_27100), .A1 (n_24989), .B0 (n_24303), .Y(n_25357));
NAND2X1 g111549(.A (n_24665), .B (n_25355), .Y (n_26799));
OAI21X1 g111560(.A0 (n_26382), .A1 (n_24186), .B0 (n_23991), .Y(n_25354));
NAND2X1 g111582(.A (n_24681), .B (n_25353), .Y (n_32532));
OAI21X1 g111583(.A0 (n_25341), .A1 (n_13758), .B0 (n_25053), .Y(n_26320));
INVX1 g111584(.A (n_25982), .Y (n_25352));
NAND2X1 g111592(.A (n_24679), .B (n_25351), .Y (n_26333));
NAND2X1 g111593(.A (n_24678), .B (n_25351), .Y (n_26312));
NAND2X1 g111598(.A (n_24672), .B (n_13639), .Y (n_26301));
NAND2X1 g111601(.A (n_24671), .B (n_13639), .Y (n_25698));
INVX1 g111605(.A (n_25052), .Y (n_25695));
NAND2X1 g111614(.A (n_24664), .B (n_25350), .Y (n_26340));
NAND2X1 g111616(.A (n_24660), .B (n_25049), .Y (n_26295));
INVX1 g111618(.A (n_25348), .Y (n_25347));
OAI21X1 g111620(.A0 (n_13944), .A1 (n_25368), .B0 (n_24659), .Y(n_25346));
NAND2X1 g111622(.A (n_24658), .B (n_25345), .Y (n_26292));
NAND2X1 g111629(.A (n_24656), .B (n_25344), .Y (n_25688));
NAND2X1 g111632(.A (n_24655), .B (n_25344), .Y (n_25686));
AOI21X1 g111634(.A0 (n_24188), .A1 (n_25220), .B0 (n_14436), .Y(n_25343));
NAND2X1 g111638(.A (n_24651), .B (n_25342), .Y (n_26338));
OAI21X1 g111641(.A0 (n_25341), .A1 (n_13273), .B0 (n_25048), .Y(n_26769));
OAI21X1 g111643(.A0 (n_23910), .A1 (n_27696), .B0 (n_24698), .Y(n_25340));
INVX1 g111652(.A (n_25338), .Y (n_25339));
NAND2X1 g111658(.A (n_24624), .B (n_20374), .Y (n_25337));
NAND2X1 g111667(.A (n_24620), .B (n_25336), .Y (n_26336));
NAND2X1 g111676(.A (n_24653), .B (n_25335), .Y (n_25677));
NAND2X1 g111677(.A (n_24682), .B (n_25335), .Y (n_26781));
NAND2X1 g111695(.A (n_24639), .B (n_25331), .Y (n_25673));
NAND2X1 g111720(.A (n_24622), .B (n_25329), .Y (n_26257));
AOI21X1 g111725(.A0 (n_14557), .A1 (n_14490), .B0 (n_24654), .Y(n_25328));
NAND2X1 g111738(.A (n_24602), .B (n_25327), .Y (n_26261));
INVX1 g111741(.A (n_25910), .Y (n_25326));
NAND2X1 g111752(.A (n_24398), .B (n_24686), .Y (n_25325));
NAND2X1 g111753(.A (n_24397), .B (n_24667), .Y (n_25324));
OAI21X1 g111754(.A0 (n_14866), .A1 (n_8614), .B0 (n_24650), .Y(n_25323));
NAND2X1 g111757(.A (n_24394), .B (n_24662), .Y (n_25322));
OAI21X1 g111761(.A0 (n_18577), .A1 (n_25540), .B0 (n_24606), .Y(n_25321));
OAI21X1 g111765(.A0 (n_24197), .A1 (n_31541), .B0 (n_7104), .Y(n_25320));
NAND2X1 g108248(.A (n_24480), .B (n_25942), .Y (n_25319));
OAI21X1 g111781(.A0 (n_24336), .A1 (n_27662), .B0 (n_24632), .Y(n_25318));
INVX1 g111786(.A (n_25317), .Y (n_26308));
NAND2X2 g111789(.A (n_35279), .B (n_35280), .Y (n_26306));
INVX1 g111790(.A (n_25957), .Y (n_25316));
NAND2X1 g111794(.A (n_24645), .B (n_24644), .Y (n_26290));
MX2X1 g111804(.A (n_17247), .B (n_19652), .S0 (n_24179), .Y(n_26283));
MX2X1 g111806(.A (n_18330), .B (n_18331), .S0 (n_24288), .Y(n_25662));
NAND2X2 g111809(.A (n_32277), .B (n_32278), .Y (n_26260));
NAND2X2 g111813(.A (n_24638), .B (n_24357), .Y (n_26259));
NAND2X1 g111817(.A (n_32922), .B (n_32923), .Y (n_26252));
NAND2X2 g111819(.A (n_35921), .B (n_35922), .Y (n_26236));
NAND2X1 g108288(.A (n_24479), .B (n_25942), .Y (n_25315));
NAND3X1 g111844(.A (n_18024), .B (n_24157), .C (n_23580), .Y(n_25313));
NAND3X1 g111852(.A (n_10884), .B (n_23590), .C (n_24160), .Y(n_25312));
NAND3X1 g111905(.A (n_23572), .B (n_24163), .C (n_23613), .Y(n_25311));
NAND2X1 g111912(.A (n_25298), .B (n_25309), .Y (n_32022));
INVX1 g111924(.A (n_25307), .Y (n_25308));
OR2X1 g111946(.A (n_25305), .B (n_25054), .Y (n_25306));
NAND2X1 g108345(.A (n_24478), .B (n_8641), .Y (n_25304));
NAND2X1 g111954(.A (n_25293), .B (n_25302), .Y (n_25303));
NAND2X1 g111957(.A (n_24509), .B (n_9431), .Y (n_25301));
NAND2X1 g111965(.A (n_25298), .B (n_25297), .Y (n_25299));
NAND2X1 g111970(.A (n_24503), .B (n_24247), .Y (n_25296));
NAND2X1 g111984(.A (n_25298), .B (n_32746), .Y (n_25295));
NAND2X1 g112016(.A (n_25293), .B (n_24361), .Y (n_25294));
NAND2X1 g112022(.A (n_24510), .B (n_8641), .Y (n_25292));
NAND3X1 g112029(.A (n_24154), .B (n_24158), .C (n_20474), .Y(n_25289));
NAND2X1 g112058(.A (n_25293), .B (n_18137), .Y (n_25288));
NAND2X1 g112059(.A (n_24507), .B (n_25942), .Y (n_25287));
NAND2X1 g112062(.A (n_25285), .B (n_25284), .Y (n_25286));
NAND2X1 g112066(.A (n_24525), .B (n_20785), .Y (n_25283));
NAND3X1 g112093(.A (n_24874), .B (n_23523), .C (n_23218), .Y(n_32237));
NAND2X1 g112104(.A (n_24519), .B (n_18967), .Y (n_35876));
OR2X1 g112150(.A (n_24833), .B (n_35719), .Y (n_25279));
NAND2X1 g112155(.A (n_24175), .B (n_18065), .Y (n_25278));
NAND2X1 g112159(.A (n_25293), .B (n_27089), .Y (n_25277));
NAND2X1 g112163(.A (n_24506), .B (n_25220), .Y (n_25276));
NAND2X1 g112194(.A (n_24192), .B (n_28136), .Y (n_25274));
NAND3X1 g112260(.A (n_10198), .B (n_24155), .C (n_23574), .Y(n_25272));
NAND2X1 g112293(.A (n_24531), .B (n_25271), .Y (n_26138));
NAND2X1 g112325(.A (n_24553), .B (n_22839), .Y (n_26129));
NAND2X1 g112327(.A (n_24552), .B (n_23542), .Y (n_26157));
NAND2X1 g112328(.A (n_24550), .B (n_23136), .Y (n_26155));
INVX1 g112339(.A (n_25270), .Y (n_25589));
NAND2X1 g112344(.A (n_24543), .B (n_24897), .Y (n_26121));
INVX1 g112345(.A (n_25268), .Y (n_25269));
OAI21X1 g112351(.A0 (n_24116), .A1 (n_32669), .B0 (n_24896), .Y(n_25266));
NAND2X1 g112358(.A (n_24540), .B (n_25264), .Y (n_25586));
NAND2X1 g112368(.A (n_24534), .B (n_24895), .Y (n_26113));
INVX1 g112369(.A (n_25814), .Y (n_25263));
NAND2X1 g112373(.A (n_24532), .B (n_24894), .Y (n_26151));
AOI21X1 g112376(.A0 (n_14394), .A1 (n_25229), .B0 (n_24530), .Y(n_25262));
NAND2X1 g112377(.A (n_24279), .B (n_24560), .Y (n_25261));
OAI21X1 g112389(.A0 (n_24113), .A1 (n_13661), .B0 (n_22836), .Y(n_26103));
NAND2X1 g112391(.A (n_24549), .B (n_24888), .Y (n_35359));
NAND2X1 g112392(.A (n_24523), .B (n_25260), .Y (n_26147));
NAND3X1 g112404(.A (n_18077), .B (n_23053), .C (n_25257), .Y(n_25259));
NAND3X1 g112436(.A (n_20562), .B (n_25257), .C (n_17345), .Y(n_25258));
NAND2X1 g112441(.A (n_24281), .B (n_24561), .Y (n_25256));
NAND2X1 g112456(.A (n_24557), .B (n_24258), .Y (n_26118));
INVX2 g112459(.A (n_25751), .Y (n_25255));
OR2X1 g112531(.A (n_25251), .B (n_8668), .Y (n_25253));
OR2X1 g112554(.A (n_25251), .B (n_7776), .Y (n_25252));
NAND2X1 g112606(.A (n_25248), .B (n_26412), .Y (n_25250));
NAND2X1 g112664(.A (n_25248), .B (n_13582), .Y (n_25249));
OR2X1 g112714(.A (n_25251), .B (n_8687), .Y (n_25247));
NAND2X1 g112724(.A (n_25251), .B (n_8680), .Y (n_25246));
NAND3X1 g112738(.A (n_22764), .B (n_24109), .C (n_19831), .Y(n_25245));
INVX1 g112851(.A (n_25632), .Y (n_25244));
INVX1 g112854(.A (n_25630), .Y (n_25243));
INVX1 g112866(.A (n_25641), .Y (n_25242));
INVX1 g112879(.A (n_25637), .Y (n_25241));
INVX1 g112882(.A (n_25634), .Y (n_25240));
INVX1 g113013(.A (n_25610), .Y (n_25570));
NAND2X1 g113036(.A (n_24485), .B (n_31850), .Y (n_25239));
NAND2X1 g113037(.A (n_24483), .B (n_31783), .Y (n_25238));
AOI21X1 g108943(.A0 (n_24474), .A1 (n_24380), .B0 (n_27008), .Y(n_25237));
NOR2X1 g113322(.A (n_21503), .B (n_24482), .Y (n_25236));
AND2X1 g109008(.A (n_25234), .B (n_33748), .Y (n_25235));
NAND2X1 g113441(.A (n_6501), .B (n_24488), .Y (n_25233));
INVX1 g113483(.A (n_25579), .Y (n_25232));
NAND3X1 g109215(.A (n_23455), .B (n_23403), .C (n_24230), .Y(n_25231));
AOI22X1 g109319(.A0 (n_15346), .A1 (n_25229), .B0 (n_24466), .B1(n_25228), .Y (n_25230));
NAND2X1 g109637(.A (n_24463), .B (n_25942), .Y (n_25226));
NAND2X1 g109666(.A (n_24465), .B (n_23771), .Y (n_25225));
NAND2X1 g109693(.A (n_24464), .B (n_8303), .Y (n_25224));
NAND2X1 g109697(.A (n_24462), .B (n_25082), .Y (n_25223));
NAND2X1 g109728(.A (n_24468), .B (n_25228), .Y (n_25222));
NAND2X1 g109734(.A (n_24461), .B (n_25220), .Y (n_25221));
NAND2X1 g109809(.A (n_24460), .B (n_9431), .Y (n_25219));
NAND2X1 g109847(.A (n_24166), .B (n_23451), .Y (n_25217));
OAI21X1 g109880(.A0 (n_14477), .A1 (n_9971), .B0 (n_24473), .Y(n_25216));
OAI21X1 g109943(.A0 (n_14470), .A1 (n_25563), .B0 (n_24471), .Y(n_25215));
NAND4X1 g110131(.A (n_24458), .B (n_21531), .C (n_19590), .D(n_22906), .Y (n_25214));
AOI21X1 g110191(.A0 (n_24820), .A1 (n_28136), .B0 (n_19919), .Y(n_25213));
AOI21X1 g110192(.A0 (n_24818), .A1 (n_28136), .B0 (n_20381), .Y(n_25212));
AOI21X1 g110215(.A0 (n_24804), .A1 (n_28136), .B0 (n_20410), .Y(n_25211));
NAND2X1 g110270(.A (n_24428), .B (n_23623), .Y (n_25210));
NAND2X1 g110416(.A (n_25201), .B (n_27091), .Y (n_25209));
NAND2X1 g110419(.A (n_25199), .B (n_25207), .Y (n_25208));
NAND2X1 g110435(.A (n_25205), .B (n_26530), .Y (n_25206));
NAND2X1 g110469(.A (n_24424), .B (n_23771), .Y (n_25204));
NAND2X1 g110475(.A (n_25205), .B (n_18918), .Y (n_25203));
NAND2X1 g110476(.A (n_25201), .B (n_28441), .Y (n_25202));
NAND2X1 g110482(.A (n_25199), .B (n_25198), .Y (n_25200));
NAND2X1 g110535(.A (n_24430), .B (n_25228), .Y (n_25197));
NAND2X1 g110542(.A (n_25201), .B (n_35054), .Y (n_25196));
NAND4X1 g110566(.A (n_24416), .B (n_21014), .C (n_22867), .D(n_23839), .Y (n_25195));
NAND2X1 g110581(.A (n_25201), .B (n_25193), .Y (n_25194));
NAND2X1 g110610(.A (n_25199), .B (n_13274), .Y (n_25185));
NOR2X1 g110646(.A (n_24433), .B (n_23752), .Y (n_25183));
NAND3X1 g110714(.A (n_17476), .B (n_19345), .C (n_24027), .Y(n_25182));
NAND3X1 g110755(.A (n_32099), .B (n_32100), .C (n_24063), .Y(n_25181));
NAND3X1 g110756(.A (n_23423), .B (n_24056), .C (n_24055), .Y(n_25180));
OAI21X1 g110809(.A0 (n_14662), .A1 (n_26372), .B0 (n_24453), .Y(n_25179));
NOR2X1 g110816(.A (n_9922), .B (n_24445), .Y (n_25178));
AOI21X1 g110818(.A0 (n_24793), .A1 (n_30180), .B0 (n_20940), .Y(n_25177));
OAI21X1 g110819(.A0 (n_14919), .A1 (n_25862), .B0 (n_24444), .Y(n_25176));
NAND2X1 g110821(.A (n_24442), .B (n_13174), .Y (n_25175));
AOI21X1 g110824(.A0 (n_24791), .A1 (n_30180), .B0 (n_20930), .Y(n_25173));
AOI21X1 g110825(.A0 (n_14860), .A1 (n_24735), .B0 (n_8927), .Y(n_25172));
NAND3X1 g110843(.A (n_9125), .B (n_24037), .C (n_20392), .Y(n_25171));
NOR2X1 g110876(.A (n_24081), .B (n_24457), .Y (n_25170));
AOI21X1 g110880(.A0 (n_24767), .A1 (n_26213), .B0 (n_20277), .Y(n_25169));
NAND2X1 g110883(.A (n_24449), .B (n_27221), .Y (n_25168));
NAND2X1 g110885(.A (n_24438), .B (n_27217), .Y (n_25167));
NAND2X1 g110886(.A (n_24437), .B (n_27227), .Y (n_25166));
NAND2X1 g110966(.A (n_24440), .B (n_28572), .Y (n_25165));
NAND4X1 g110977(.A (n_23993), .B (n_24014), .C (n_23740), .D(n_23392), .Y (n_25164));
OAI21X1 g110979(.A0 (n_15055), .A1 (n_8614), .B0 (n_24443), .Y(n_25163));
AOI21X1 g110980(.A0 (n_24762), .A1 (n_14630), .B0 (n_26920), .Y(n_25162));
AOI21X1 g110981(.A0 (n_24759), .A1 (n_14727), .B0 (n_29725), .Y(n_25161));
AOI21X1 g110985(.A0 (n_24750), .A1 (n_14561), .B0 (n_29725), .Y(n_25160));
AOI21X1 g110991(.A0 (n_24783), .A1 (n_26213), .B0 (n_20297), .Y(n_25159));
AOI21X1 g110995(.A0 (n_24777), .A1 (n_26213), .B0 (n_20288), .Y(n_25158));
AOI22X1 g111000(.A0 (n_24771), .A1 (n_26213), .B0 (n_20304), .B1(n_18414), .Y (n_25157));
AOI21X1 g111012(.A0 (n_24733), .A1 (n_28158), .B0 (n_15032), .Y(n_25155));
NAND2X1 g111022(.A (n_24454), .B (n_28556), .Y (n_25154));
NAND3X1 g111024(.A (n_24080), .B (n_21282), .C (n_24076), .Y(n_25153));
NAND2X1 g111025(.A (n_24448), .B (n_25151), .Y (n_25152));
NAND3X1 g111026(.A (n_24079), .B (n_21278), .C (n_24075), .Y(n_25150));
OAI21X1 g111028(.A0 (n_23987), .A1 (n_32765), .B0 (n_28551), .Y(n_25149));
OAI21X1 g111055(.A0 (n_24292), .A1 (n_35555), .B0 (n_25148), .Y(n_26428));
NAND3X1 g111106(.A (n_24318), .B (n_23668), .C (n_23376), .Y(n_25147));
NAND3X1 g111110(.A (n_33015), .B (n_33016), .C (n_23639), .Y(n_25447));
NOR2X1 g111113(.A (n_23384), .B (n_24293), .Y (n_25146));
NAND2X1 g111130(.A (n_25131), .B (n_34952), .Y (n_25145));
NAND2X1 g111135(.A (n_25140), .B (n_26162), .Y (n_25144));
NAND2X1 g111144(.A (n_25142), .B (n_34694), .Y (n_25143));
NAND2X1 g111155(.A (n_25140), .B (n_28492), .Y (n_25141));
NAND2X1 g111161(.A (n_25138), .B (n_28492), .Y (n_25139));
NAND2X1 g111165(.A (n_26978), .B (n_25136), .Y (n_25137));
NAND3X1 g111166(.A (n_23724), .B (n_23981), .C (n_23739), .Y(n_25135));
NAND2X1 g111168(.A (n_25142), .B (n_26142), .Y (n_25134));
NAND3X1 g111173(.A (n_23714), .B (n_23978), .C (n_23737), .Y(n_25133));
NAND2X1 g111177(.A (n_25131), .B (n_26142), .Y (n_25132));
NAND3X1 g111181(.A (n_23704), .B (n_23976), .C (n_23734), .Y(n_25130));
NAND2X1 g111185(.A (n_25140), .B (n_29090), .Y (n_25129));
NAND2X1 g111193(.A (n_26978), .B (n_25127), .Y (n_25128));
NAND2X1 g111194(.A (n_25138), .B (n_26142), .Y (n_25126));
NOR2X1 g111197(.A (n_27256), .B (n_24304), .Y (n_25125));
NAND2X1 g111214(.A (n_34810), .B (n_21272), .Y (n_25124));
NAND2X1 g111216(.A (n_24314), .B (n_25122), .Y (n_25123));
NAND2X1 g111222(.A (n_25136), .B (n_26870), .Y (n_25121));
NOR2X1 g111223(.A (n_24313), .B (n_25119), .Y (n_25120));
NAND2X1 g111228(.A (n_25109), .B (n_25554), .Y (n_25118));
NAND2X1 g111232(.A (n_25106), .B (n_28441), .Y (n_25116));
NAND2X1 g111261(.A (n_24302), .B (n_8641), .Y (n_25115));
NAND2X1 g111266(.A (n_24311), .B (n_25122), .Y (n_32116));
AOI21X1 g108044(.A0 (n_23818), .A1 (n_26458), .B0 (n_14924), .Y(n_25113));
NAND2X1 g111305(.A (n_24308), .B (n_25111), .Y (n_25112));
NAND2X1 g111310(.A (n_25109), .B (n_24361), .Y (n_25110));
NAND2X1 g111316(.A (n_25106), .B (n_27770), .Y (n_25107));
NAND2X1 g111344(.A (n_24321), .B (n_25220), .Y (n_25105));
NAND2X1 g111348(.A (n_24323), .B (n_8303), .Y (n_25103));
NAND2X1 g111349(.A (n_25109), .B (n_26637), .Y (n_25102));
NAND2X1 g111362(.A (n_25094), .B (n_35736), .Y (n_25919));
NAND2X1 g111365(.A (n_25106), .B (n_25193), .Y (n_25101));
NAND2X1 g111375(.A (n_24300), .B (n_25220), .Y (n_25100));
NAND2X1 g111377(.A (n_25109), .B (n_25098), .Y (n_25099));
INVX1 g111380(.A (n_25096), .Y (n_25097));
NAND2X1 g111390(.A (n_25094), .B (n_14439), .Y (n_25095));
NAND2X1 g111392(.A (n_25085), .B (n_24965), .Y (n_25394));
NAND2X1 g111395(.A (n_21429), .B (n_24643), .Y (n_32217));
INVX1 g111399(.A (n_34493), .Y (n_25092));
NAND2X1 g111406(.A (n_24717), .B (n_25079), .Y (n_25927));
NAND2X1 g111411(.A (n_25073), .B (n_35816), .Y (n_25923));
NAND2X1 g111421(.A (n_25127), .B (n_26870), .Y (n_25089));
OR2X1 g111429(.A (n_24567), .B (n_35775), .Y (n_25088));
NAND2X1 g111434(.A (n_25085), .B (n_35822), .Y (n_25086));
NAND2X1 g111436(.A (n_25106), .B (n_27091), .Y (n_25084));
NAND2X1 g111450(.A (n_24298), .B (n_25082), .Y (n_25083));
NAND2X1 g111460(.A (n_24090), .B (n_25081), .Y (n_25887));
NAND2X1 g111461(.A (n_25079), .B (n_14600), .Y (n_25080));
NAND4X1 g111467(.A (n_24217), .B (n_23562), .C (n_22559), .D(n_19889), .Y (n_25078));
NAND2X1 g111470(.A (n_24415), .B (n_20778), .Y (n_32078));
NOR2X1 g111483(.A (n_27256), .B (n_24297), .Y (n_25076));
NAND4X1 g111485(.A (n_32876), .B (n_32877), .C (n_22557), .D(n_20432), .Y (n_25075));
NAND2X1 g111486(.A (n_25094), .B (n_35479), .Y (n_25074));
NAND2X1 g111489(.A (n_25085), .B (n_35576), .Y (n_25873));
NAND2X1 g111490(.A (n_25073), .B (n_25072), .Y (n_25908));
NAND2X1 g111493(.A (n_25094), .B (n_22021), .Y (n_25921));
NAND3X1 g111498(.A (n_23691), .B (n_23974), .C (n_23732), .Y(n_25071));
OAI21X1 g111503(.A0 (n_14650), .A1 (n_8614), .B0 (n_24393), .Y(n_25070));
OAI21X1 g111511(.A0 (n_14646), .A1 (n_25067), .B0 (n_24381), .Y(n_25069));
OAI21X1 g111518(.A0 (n_14870), .A1 (n_25067), .B0 (n_24376), .Y(n_25068));
OAI21X1 g111519(.A0 (n_23911), .A1 (n_8065), .B0 (n_15353), .Y(n_25066));
NOR2X1 g111529(.A (n_9046), .B (n_24294), .Y (n_25065));
AOI21X1 g111532(.A0 (n_24925), .A1 (n_24631), .B0 (n_24325), .Y(n_25064));
AOI21X1 g111534(.A0 (n_14854), .A1 (n_24612), .B0 (n_8927), .Y(n_25063));
NOR2X1 g111536(.A (n_9059), .B (n_24306), .Y (n_25062));
AOI21X1 g111541(.A0 (n_27100), .A1 (n_24617), .B0 (n_23742), .Y(n_25061));
NAND4X1 g111544(.A (n_23323), .B (n_23964), .C (n_23250), .D(n_22950), .Y (n_25059));
NAND2X1 g111552(.A (n_24363), .B (n_25058), .Y (n_25951));
NAND2X1 g111553(.A (n_24362), .B (n_25058), .Y (n_25989));
NOR2X1 g111572(.A (n_6773), .B (n_24417), .Y (n_25057));
NAND2X1 g111575(.A (n_24387), .B (n_25056), .Y (n_25972));
NAND2X1 g111576(.A (n_24385), .B (n_25056), .Y (n_25995));
NAND2X1 g111578(.A (n_24384), .B (n_25055), .Y (n_26392));
OAI21X1 g111585(.A0 (n_25050), .A1 (n_25054), .B0 (n_25053), .Y(n_25982));
NAND2X1 g111606(.A (n_24375), .B (n_25051), .Y (n_25052));
NAND2X1 g111607(.A (n_24373), .B (n_25051), .Y (n_25993));
OAI21X1 g111619(.A0 (n_25050), .A1 (n_25694), .B0 (n_25049), .Y(n_25348));
NAND2X1 g111640(.A (n_24367), .B (n_25048), .Y (n_25991));
AOI21X1 g111653(.A0 (n_21467), .A1 (n_35035), .B0 (n_22609), .Y(n_25338));
NAND2X1 g111656(.A (n_24350), .B (n_25047), .Y (n_25916));
NAND2X1 g111657(.A (n_24349), .B (n_25047), .Y (n_25986));
OAI21X1 g111682(.A0 (n_14640), .A1 (n_8614), .B0 (n_24368), .Y(n_25046));
INVX1 g111685(.A (n_25043), .Y (n_26361));
INVX1 g111689(.A (n_25041), .Y (n_26368));
INVX1 g111704(.A (n_25039), .Y (n_26366));
NAND2X1 g111709(.A (n_24344), .B (n_28196), .Y (n_25038));
NAND2X1 g111710(.A (n_24382), .B (n_28215), .Y (n_25037));
OAI21X1 g111711(.A0 (n_24174), .A1 (n_35570), .B0 (n_25035), .Y(n_25890));
NAND2X1 g111724(.A (n_24370), .B (n_28205), .Y (n_25034));
NAND2X1 g111728(.A (n_24360), .B (n_28202), .Y (n_25033));
NAND2X1 g111729(.A (n_24359), .B (n_28061), .Y (n_25032));
NAND3X1 g111730(.A (n_24640), .B (n_33017), .C (n_21482), .Y(n_32141));
INVX1 g111733(.A (n_25504), .Y (n_25030));
NAND2X1 g111742(.A (n_24333), .B (n_24751), .Y (n_25910));
NAND2X1 g111746(.A (n_24346), .B (n_24764), .Y (n_25900));
NAND2X1 g111750(.A (n_24343), .B (n_28064), .Y (n_25029));
NAND2X1 g111756(.A (n_14329), .B (n_24407), .Y (n_25028));
OAI21X1 g111760(.A0 (n_19139), .A1 (n_25540), .B0 (n_24339), .Y(n_25027));
INVX1 g111763(.A (n_25024), .Y (n_25025));
OAI21X1 g111767(.A0 (n_23922), .A1 (n_31149), .B0 (n_6737), .Y(n_25023));
OAI21X1 g111771(.A0 (n_23914), .A1 (n_33201), .B0 (n_6623), .Y(n_25022));
MX2X1 g111787(.A (n_18323), .B (n_18322), .S0 (n_23913), .Y(n_25317));
MX2X1 g111791(.A (n_19730), .B (n_21735), .S0 (n_23947), .Y(n_25957));
NAND2X1 g111807(.A (n_24043), .B (n_24358), .Y (n_25918));
MX2X1 g111808(.A (n_20269), .B (n_22144), .S0 (n_23944), .Y(n_25906));
INVX1 g111810(.A (n_25475), .Y (n_25021));
MX2X1 g111812(.A (n_22143), .B (n_20787), .S0 (n_23927), .Y(n_25903));
INVX1 g111824(.A (n_25513), .Y (n_25020));
NAND3X1 g111843(.A (n_23814), .B (n_23888), .C (n_23212), .Y(n_25019));
OAI21X1 g111861(.A0 (n_23863), .A1 (n_22526), .B0 (n_33123), .Y(n_25018));
NAND2X1 g111866(.A (n_27614), .B (n_24924), .Y (n_25017));
NAND2X1 g111894(.A (n_22962), .B (n_24914), .Y (n_25016));
NAND4X1 g111910(.A (n_15002), .B (n_23497), .C (n_22382), .D(n_23498), .Y (n_25015));
NAND2X1 g111913(.A (n_24260), .B (n_18354), .Y (n_25014));
NAND2X1 g111916(.A (n_24195), .B (n_8303), .Y (n_35269));
NAND2X1 g111921(.A (n_24191), .B (n_8303), .Y (n_25011));
NAND3X1 g111925(.A (n_32107), .B (n_23862), .C (n_32108), .Y(n_25307));
NAND2X1 g111933(.A (n_24942), .B (n_27522), .Y (n_25010));
NAND2X1 g111940(.A (n_24998), .B (n_25554), .Y (n_25009));
NAND2X1 g111944(.A (n_24987), .B (n_25554), .Y (n_25008));
NAND2X1 g111952(.A (n_24993), .B (n_25554), .Y (n_25007));
NAND2X1 g111953(.A (n_24991), .B (n_25554), .Y (n_25006));
NAND2X1 g111959(.A (n_24189), .B (n_25942), .Y (n_25005));
NAND2X1 g111966(.A (n_24985), .B (n_25003), .Y (n_25004));
NAND2X1 g111980(.A (n_24963), .B (n_35736), .Y (n_25736));
OR2X1 g111997(.A (n_24194), .B (n_8065), .Y (n_25001));
NAND2X1 g111998(.A (n_24998), .B (n_27770), .Y (n_24999));
NAND2X1 g112000(.A (n_24497), .B (n_27770), .Y (n_24997));
NAND2X1 g112002(.A (n_24998), .B (n_13274), .Y (n_24995));
NAND2X1 g112009(.A (n_24993), .B (n_24361), .Y (n_24994));
NAND2X1 g112015(.A (n_24991), .B (n_23192), .Y (n_24992));
NAND2X1 g112017(.A (n_24989), .B (n_29505), .Y (n_24990));
NAND2X1 g112018(.A (n_24987), .B (n_18137), .Y (n_24988));
NAND2X1 g112026(.A (n_24985), .B (n_24984), .Y (n_24986));
NAND2X1 g112040(.A (n_24196), .B (n_8303), .Y (n_24983));
NAND2X1 g112052(.A (n_24993), .B (n_26637), .Y (n_24982));
NAND2X1 g112055(.A (n_24991), .B (n_26637), .Y (n_24981));
NAND2X1 g112063(.A (n_24187), .B (n_9431), .Y (n_24980));
NAND2X1 g112064(.A (n_24978), .B (n_24977), .Y (n_24979));
NAND2X1 g112065(.A (n_24524), .B (n_20267), .Y (n_24976));
NAND2X1 g112069(.A (n_24182), .B (n_21740), .Y (n_24975));
INVX1 g112074(.A (n_24972), .Y (n_24973));
NAND2X1 g112077(.A (n_24200), .B (n_18362), .Y (n_24971));
NAND2X1 g112080(.A (n_24221), .B (n_18333), .Y (n_24970));
OAI21X1 g112082(.A0 (n_23864), .A1 (n_22527), .B0 (n_31878), .Y(n_24966));
NAND2X1 g112087(.A (n_24940), .B (n_24965), .Y (n_25742));
NAND2X1 g112090(.A (n_24963), .B (n_18262), .Y (n_24964));
NAND3X1 g112098(.A (n_23860), .B (n_23852), .C (n_15163), .Y(n_24962));
NOR2X1 g112102(.A (n_24211), .B (n_14221), .Y (n_24959));
NAND2X1 g112103(.A (n_33911), .B (n_20212), .Y (n_35877));
NAND2X1 g112105(.A (n_24215), .B (n_18978), .Y (n_32244));
NAND2X1 g112112(.A (n_24213), .B (n_18326), .Y (n_24955));
NAND2X1 g112117(.A (n_8990), .B (n_24950), .Y (n_24951));
NAND2X1 g112118(.A (n_8990), .B (n_24947), .Y (n_24949));
NAND2X1 g112134(.A (n_24944), .B (n_27462), .Y (n_24946));
NAND2X1 g112136(.A (n_24944), .B (n_27522), .Y (n_24945));
NAND2X1 g112137(.A (n_24942), .B (n_27462), .Y (n_24943));
NAND2X1 g112146(.A (n_24940), .B (n_35794), .Y (n_24941));
NAND2X1 g112147(.A (n_24987), .B (n_26676), .Y (n_24938));
NAND2X1 g112153(.A (n_23894), .B (n_25605), .Y (n_24937));
NAND2X1 g112154(.A (n_27614), .B (n_24927), .Y (n_24936));
NAND2X1 g112157(.A (n_24993), .B (n_25098), .Y (n_24935));
NAND2X1 g112158(.A (n_24991), .B (n_24101), .Y (n_24934));
NAND2X1 g112161(.A (n_24932), .B (n_29505), .Y (n_24933));
NAND2X1 g112162(.A (n_24932), .B (n_26132), .Y (n_24931));
NAND2X1 g112164(.A (n_24989), .B (n_29430), .Y (n_24930));
NAND2X1 g112168(.A (n_24185), .B (n_25220), .Y (n_24929));
NAND2X1 g112172(.A (n_24925), .B (n_24927), .Y (n_24928));
NAND2X1 g112174(.A (n_24925), .B (n_24924), .Y (n_24926));
NAND2X1 g112175(.A (n_24985), .B (n_26530), .Y (n_24923));
INVX1 g112178(.A (n_24613), .Y (n_25275));
OAI21X1 g112192(.A0 (n_23855), .A1 (n_9626), .B0 (n_22822), .Y(n_24922));
NAND2X1 g112193(.A (n_23905), .B (n_28136), .Y (n_24920));
NAND4X1 g112196(.A (n_14823), .B (n_23502), .C (n_22387), .D(n_23500), .Y (n_24919));
NOR2X1 g112202(.A (n_24917), .B (n_25881), .Y (n_24918));
NAND2X1 g112211(.A (n_22278), .B (n_24914), .Y (n_24915));
NAND2X1 g112213(.A (n_24940), .B (n_35540), .Y (n_25723));
NAND2X1 g112216(.A (n_24494), .B (n_35528), .Y (n_25792));
NAND2X1 g112220(.A (n_24940), .B (n_25599), .Y (n_24913));
NAND2X1 g112222(.A (n_24963), .B (n_25877), .Y (n_25738));
OAI21X1 g112246(.A0 (n_14791), .A1 (n_25862), .B0 (n_24232), .Y(n_24912));
INVX1 g112257(.A (n_34834), .Y (n_24911));
NAND2X1 g112268(.A (n_24254), .B (n_18225), .Y (n_24909));
NAND2X1 g112269(.A (n_24208), .B (n_27522), .Y (n_24908));
NAND2X1 g112270(.A (n_24205), .B (n_27522), .Y (n_24907));
NAND2X1 g112274(.A (n_24243), .B (n_28555), .Y (n_24905));
NAND2X1 g112275(.A (n_24241), .B (n_28542), .Y (n_24904));
OAI21X1 g112277(.A0 (n_23846), .A1 (n_24013), .B0 (n_24324), .Y(n_25767));
NAND2X1 g112283(.A (n_24224), .B (n_24011), .Y (n_25820));
NAND2X1 g112285(.A (n_24219), .B (n_28548), .Y (n_24903));
NAND2X1 g112306(.A (n_24222), .B (n_27708), .Y (n_24900));
NAND2X1 g112307(.A (n_24206), .B (n_27702), .Y (n_24899));
NAND2X1 g108482(.A (n_24131), .B (n_25856), .Y (n_24898));
NAND2X1 g112321(.A (n_24251), .B (n_22441), .Y (n_25803));
NAND2X1 g112326(.A (n_24250), .B (n_23542), .Y (n_25798));
NAND2X1 g112340(.A (n_24240), .B (n_24309), .Y (n_25270));
OAI21X1 g112347(.A0 (n_24114), .A1 (n_32654), .B0 (n_24897), .Y(n_25268));
NAND2X1 g112348(.A (n_24238), .B (n_24896), .Y (n_25782));
NAND2X1 g112359(.A (n_24235), .B (n_13638), .Y (n_25777));
NAND2X1 g112370(.A (n_24229), .B (n_24895), .Y (n_25814));
OAI21X1 g112371(.A0 (n_23843), .A1 (n_24893), .B0 (n_24894), .Y(n_25763));
OAI21X1 g112374(.A0 (n_24891), .A1 (n_24893), .B0 (n_24892), .Y(n_25757));
OAI21X1 g112381(.A0 (n_24891), .A1 (n_26210), .B0 (n_24890), .Y(n_26181));
OAI21X1 g112386(.A0 (n_23846), .A1 (n_24889), .B0 (n_24305), .Y(n_25785));
OAI21X1 g112390(.A0 (n_23843), .A1 (n_24889), .B0 (n_24888), .Y(n_25805));
OAI21X1 g112412(.A0 (n_23856), .A1 (n_8305), .B0 (n_23425), .Y(n_24887));
NAND2X1 g112414(.A (n_24275), .B (n_10238), .Y (n_24886));
NAND2X1 g112416(.A (n_15000), .B (n_24227), .Y (n_24885));
NAND2X1 g112418(.A (n_24263), .B (n_10145), .Y (n_24884));
INVX1 g112423(.A (n_25381), .Y (n_24883));
NAND2X1 g112437(.A (n_24285), .B (n_23431), .Y (n_24882));
OAI21X1 g112440(.A0 (n_23854), .A1 (n_10785), .B0 (n_23430), .Y(n_24881));
NAND2X1 g108547(.A (n_24142), .B (n_25852), .Y (n_24880));
OAI21X1 g112443(.A0 (n_23853), .A1 (n_27696), .B0 (n_23429), .Y(n_24879));
INVX2 g112447(.A (n_24569), .Y (n_26205));
NAND2X2 g112458(.A (n_23960), .B (n_24255), .Y (n_25790));
NAND2X2 g112461(.A (n_32916), .B (n_32917), .Y (n_25751));
NAND2X1 g112464(.A (n_23948), .B (n_24223), .Y (n_25769));
NAND2X1 g112477(.A (n_24290), .B (n_23984), .Y (n_25787));
NOR2X1 g112483(.A (n_23033), .B (n_24127), .Y (n_24877));
NAND2X1 g108583(.A (n_24123), .B (n_25850), .Y (n_24876));
INVX1 g112504(.A (n_24874), .Y (n_24875));
OAI21X1 g108598(.A0 (n_24100), .A1 (n_13317), .B0 (n_25849), .Y(n_24873));
NAND2X1 g112514(.A (n_24865), .B (n_28864), .Y (n_24872));
NAND2X1 g112517(.A (n_24863), .B (n_29061), .Y (n_24871));
NAND2X1 g112521(.A (n_24868), .B (n_27335), .Y (n_24869));
NAND2X1 g112524(.A (n_24859), .B (n_30563), .Y (n_24867));
NAND2X1 g112527(.A (n_24865), .B (n_28485), .Y (n_24866));
NAND2X1 g112530(.A (n_24863), .B (n_28485), .Y (n_24864));
NAND2X1 g112537(.A (n_24868), .B (n_29604), .Y (n_24861));
NAND2X1 g112541(.A (n_24859), .B (n_26535), .Y (n_24860));
NAND2X1 g112547(.A (n_24865), .B (n_30197), .Y (n_24858));
NAND2X1 g112551(.A (n_24863), .B (n_28468), .Y (n_24857));
NAND2X1 g112599(.A (n_23844), .B (n_25003), .Y (n_24853));
NAND2X1 g112608(.A (n_23847), .B (n_18918), .Y (n_24852));
NAND2X1 g112611(.A (n_24122), .B (n_8303), .Y (n_24850));
NOR2X1 g112762(.A (n_24118), .B (n_10556), .Y (n_24848));
NAND2X1 g112765(.A (n_23844), .B (n_26530), .Y (n_24847));
NAND2X1 g112787(.A (n_24126), .B (n_23226), .Y (n_24845));
NAND2X1 g108720(.A (n_23884), .B (n_24167), .Y (n_25953));
NOR2X1 g112827(.A (n_9111), .B (n_24120), .Y (n_24844));
NAND2X1 g112852(.A (n_24141), .B (n_23647), .Y (n_25632));
NAND2X1 g112853(.A (n_24140), .B (n_24843), .Y (n_25612));
NAND2X1 g112855(.A (n_24139), .B (n_24843), .Y (n_25630));
AOI22X1 g112860(.A0 (n_23832), .A1 (n_24841), .B0 (n_20629), .B1(n_22883), .Y (n_24842));
NAND2X1 g112867(.A (n_24153), .B (n_23642), .Y (n_25641));
NAND2X1 g112869(.A (n_24152), .B (n_24840), .Y (n_25647));
NAND2X1 g112870(.A (n_24151), .B (n_24840), .Y (n_25626));
NAND2X1 g112880(.A (n_24148), .B (n_23640), .Y (n_25637));
NAND2X1 g112881(.A (n_24147), .B (n_24839), .Y (n_25621));
NAND2X1 g112883(.A (n_24145), .B (n_24839), .Y (n_25634));
OAI21X1 g112888(.A0 (n_23829), .A1 (n_27696), .B0 (n_23615), .Y(n_24838));
NAND2X1 g112891(.A (n_24135), .B (n_24837), .Y (n_25608));
NAND2X1 g112896(.A (n_24150), .B (n_23637), .Y (n_25645));
NAND2X1 g112898(.A (n_24134), .B (n_24837), .Y (n_25643));
NOR2X1 g112921(.A (n_23835), .B (n_24117), .Y (n_24836));
OAI21X1 g112971(.A0 (n_23828), .A1 (n_10785), .B0 (n_23616), .Y(n_24835));
XOR2X1 g112998(.A (n_22193), .B (n_23831), .Y (n_25617));
NAND2X1 g113008(.A (n_24138), .B (n_23869), .Y (n_25602));
INVX1 g113014(.A (n_24495), .Y (n_25610));
NAND2X1 g113032(.A (n_23465), .B (n_24112), .Y (n_24832));
OAI21X1 g108914(.A0 (n_24099), .A1 (n_24065), .B0 (n_27485), .Y(n_24831));
NOR2X1 g113207(.A (n_22198), .B (n_24108), .Y (n_24830));
AOI22X1 g113371(.A0 (n_23820), .A1 (n_23474), .B0 (n_20622), .B1(n_23215), .Y (n_24829));
NAND2X1 g113484(.A (n_24110), .B (n_23836), .Y (n_25579));
INVX1 g113485(.A (n_25248), .Y (n_24828));
INVX1 g113486(.A (n_25248), .Y (n_24827));
NAND2X1 g111766(.A (n_24330), .B (n_19938), .Y (n_24826));
AOI21X1 g109841(.A0 (n_28597), .A1 (n_24164), .B0 (n_23802), .Y(n_24825));
OAI21X1 g109921(.A0 (n_23800), .A1 (n_22239), .B0 (n_23896), .Y(n_25234));
OAI21X1 g110038(.A0 (n_23784), .A1 (n_8940), .B0 (n_14744), .Y(n_24824));
NAND4X1 g110266(.A (n_23970), .B (n_19189), .C (n_22077), .D(n_22731), .Y (n_24823));
NAND3X1 g110309(.A (n_18013), .B (n_19930), .C (n_23777), .Y(n_24822));
NAND2X1 g110411(.A (n_24820), .B (n_8954), .Y (n_24821));
NAND2X1 g110412(.A (n_24818), .B (n_8954), .Y (n_24819));
AOI21X1 g110433(.A0 (n_23773), .A1 (n_18310), .B0 (n_26052), .Y(n_24817));
AOI21X1 g110474(.A0 (n_23768), .A1 (n_13646), .B0 (n_26052), .Y(n_24816));
AOI21X1 g110496(.A0 (n_23764), .A1 (n_26558), .B0 (n_26052), .Y(n_24815));
AOI21X1 g110502(.A0 (n_23763), .A1 (n_14097), .B0 (n_26052), .Y(n_24814));
NAND2X1 g107722(.A (n_24001), .B (n_8641), .Y (n_24812));
NAND2X1 g107759(.A (n_23999), .B (n_26458), .Y (n_24811));
NAND2X1 g107774(.A (n_23998), .B (n_8641), .Y (n_24810));
NAND2X1 g110684(.A (n_24820), .B (n_26238), .Y (n_24809));
NAND2X1 g110687(.A (n_24818), .B (n_26238), .Y (n_24808));
NAND2X1 g110688(.A (n_24818), .B (n_28158), .Y (n_24807));
NAND2X1 g110707(.A (n_24820), .B (n_28158), .Y (n_24806));
NAND2X1 g110718(.A (n_24804), .B (n_28158), .Y (n_24805));
NAND2X1 g110719(.A (n_24804), .B (n_26238), .Y (n_24803));
NAND2X1 g110723(.A (n_24804), .B (n_8954), .Y (n_24802));
OAI21X1 g110808(.A0 (n_14017), .A1 (n_14658), .B0 (n_24096), .Y(n_24801));
NAND4X1 g110823(.A (n_23923), .B (n_19276), .C (n_22076), .D(n_22730), .Y (n_24799));
NAND2X1 g107868(.A (n_23997), .B (n_8641), .Y (n_24798));
AOI21X1 g111013(.A0 (n_23747), .A1 (n_26458), .B0 (n_14917), .Y(n_24797));
XOR2X1 g111102(.A (n_16777), .B (n_23755), .Y (n_25555));
NOR2X1 g111105(.A (n_22420), .B (n_24050), .Y (n_24796));
NAND3X1 g111114(.A (n_10122), .B (n_19358), .C (n_23664), .Y(n_24795));
NAND2X1 g111120(.A (n_33546), .B (n_24793), .Y (n_24794));
NAND2X1 g111124(.A (n_33546), .B (n_24791), .Y (n_24792));
NAND2X1 g111218(.A (n_24788), .B (n_26611), .Y (n_24790));
NAND2X1 g111220(.A (n_24788), .B (n_30180), .Y (n_24789));
NAND2X1 g111221(.A (n_24788), .B (n_24786), .Y (n_24787));
NAND2X1 g111225(.A (n_24785), .B (n_24779), .Y (n_25469));
NAND2X1 g111231(.A (n_24783), .B (n_28785), .Y (n_32135));
NAND2X1 g111234(.A (n_24783), .B (n_24526), .Y (n_24782));
NAND2X1 g111235(.A (n_24783), .B (n_26288), .Y (n_24781));
NAND2X1 g111255(.A (n_14723), .B (n_24779), .Y (n_24780));
NAND2X1 g111272(.A (n_24777), .B (n_28785), .Y (n_32150));
NAND2X1 g111273(.A (n_24777), .B (n_24526), .Y (n_24776));
NAND2X1 g111274(.A (n_24777), .B (n_26288), .Y (n_24775));
NAND2X1 g111300(.A (n_24793), .B (n_28431), .Y (n_24774));
NAND4X1 g111309(.A (n_18742), .B (n_20689), .C (n_23365), .D(n_21987), .Y (n_24773));
NAND2X1 g111312(.A (n_24771), .B (n_28785), .Y (n_24772));
NAND2X1 g111314(.A (n_24771), .B (n_24526), .Y (n_24770));
NAND2X1 g111315(.A (n_24771), .B (n_30063), .Y (n_24769));
NAND2X1 g111354(.A (n_24767), .B (n_28785), .Y (n_32083));
NAND2X1 g111355(.A (n_24767), .B (n_34753), .Y (n_24766));
NAND2X1 g111356(.A (n_24767), .B (n_26288), .Y (n_24765));
NAND2X1 g111359(.A (n_24748), .B (n_24764), .Y (n_25476));
NAND2X1 g111360(.A (n_24791), .B (n_24786), .Y (n_24763));
NAND3X1 g111381(.A (n_20826), .B (n_23660), .C (n_23682), .Y(n_25096));
NAND2X1 g111382(.A (n_24719), .B (n_24745), .Y (n_25515));
NAND2X1 g111407(.A (n_24711), .B (n_24762), .Y (n_25489));
NAND2X1 g111408(.A (n_14414), .B (n_24747), .Y (n_24761));
NAND2X1 g111410(.A (n_24760), .B (n_24759), .Y (n_25486));
NAND2X1 g111418(.A (n_24756), .B (n_26611), .Y (n_24758));
NAND2X1 g111419(.A (n_24756), .B (n_30180), .Y (n_24757));
NAND2X1 g111420(.A (n_24756), .B (n_24786), .Y (n_24755));
AND2X1 g111422(.A (n_24756), .B (n_33513), .Y (n_24754));
NAND2X1 g111423(.A (n_24752), .B (n_24741), .Y (n_24753));
NAND2X1 g111426(.A (n_24751), .B (n_24750), .Y (n_25483));
NAND2X1 g111427(.A (n_14572), .B (n_24748), .Y (n_24749));
NAND2X1 g111428(.A (n_24747), .B (n_24713), .Y (n_25472));
NAND2X1 g111441(.A (n_24745), .B (n_14660), .Y (n_24746));
NAND2X1 g111458(.A (n_24743), .B (n_29405), .Y (n_24744));
NAND2X1 g111468(.A (n_24741), .B (n_27902), .Y (n_24742));
NAND2X1 g111469(.A (n_34604), .B (n_20777), .Y (n_32079));
NAND2X1 g111481(.A (n_24737), .B (n_28136), .Y (n_24739));
NAND2X1 g111484(.A (n_24737), .B (n_29405), .Y (n_24738));
NAND2X1 g111488(.A (n_24291), .B (n_35479), .Y (n_25492));
NAND2X1 g111492(.A (n_24088), .B (n_24735), .Y (n_25493));
NAND2X1 g111494(.A (n_24752), .B (n_24733), .Y (n_24734));
NOR2X1 g111496(.A (n_22422), .B (n_23989), .Y (n_24732));
NOR2X1 g111497(.A (n_22421), .B (n_23988), .Y (n_24731));
NOR2X1 g111502(.A (n_24020), .B (n_14643), .Y (n_35885));
NOR2X1 g111554(.A (n_23728), .B (n_23995), .Y (n_24729));
NAND4X1 g111566(.A (n_19296), .B (n_22436), .C (n_23315), .D(n_15162), .Y (n_24728));
NAND4X1 g111567(.A (n_32871), .B (n_22435), .C (n_23314), .D(n_32872), .Y (n_24727));
AOI21X1 g111569(.A0 (n_34770), .A1 (n_24404), .B0 (n_14342), .Y(n_24726));
AOI21X1 g111570(.A0 (n_28948), .A1 (n_24401), .B0 (n_14560), .Y(n_24725));
NOR2X1 g111571(.A (n_6995), .B (n_24083), .Y (n_24724));
AOI21X1 g111573(.A0 (n_34770), .A1 (n_24399), .B0 (n_14787), .Y(n_24723));
OAI21X1 g111639(.A0 (n_33555), .A1 (n_13183), .B0 (n_13171), .Y(n_24722));
OAI21X1 g111662(.A0 (n_24383), .A1 (n_13184), .B0 (n_24721), .Y(n_26017));
NAND2X1 g111687(.A (n_24046), .B (n_24719), .Y (n_25043));
NAND2X1 g111691(.A (n_24044), .B (n_24718), .Y (n_25041));
NAND2X1 g111706(.A (n_24039), .B (n_24717), .Y (n_25039));
NAND2X1 g111708(.A (n_24070), .B (n_9594), .Y (n_24716));
OAI21X1 g111712(.A0 (n_33555), .A1 (n_13990), .B0 (n_28063), .Y(n_24715));
NAND2X1 g111713(.A (n_24033), .B (n_24713), .Y (n_25499));
NAND2X1 g111715(.A (n_24068), .B (n_9573), .Y (n_24712));
NAND2X1 g111734(.A (n_24019), .B (n_24711), .Y (n_25504));
NAND2X1 g111740(.A (n_24036), .B (n_28136), .Y (n_24710));
OAI21X1 g111748(.A0 (n_23893), .A1 (n_35520), .B0 (n_24709), .Y(n_25529));
NAND2X1 g108241(.A (n_23819), .B (n_8641), .Y (n_24708));
NAND3X1 g111758(.A (n_35389), .B (n_32151), .C (n_21480), .Y(n_32019));
OAI21X1 g111762(.A0 (n_19664), .A1 (n_25540), .B0 (n_24022), .Y(n_24706));
AOI21X1 g111764(.A0 (n_23963), .A1 (n_32095), .B0 (n_22617), .Y(n_25024));
NAND2X1 g111768(.A (n_6639), .B (n_24084), .Y (n_24705));
OAI21X1 g111773(.A0 (n_19672), .A1 (n_25540), .B0 (n_24016), .Y(n_24704));
MX2X1 g111811(.A (n_19273), .B (n_22142), .S0 (n_23677), .Y(n_25475));
XOR2X1 g111825(.A (n_16740), .B (n_23674), .Y (n_25513));
AOI21X1 g111837(.A0 (n_22612), .A1 (n_23298), .B0 (n_23840), .Y(n_24703));
NAND3X1 g111846(.A (n_35272), .B (n_35273), .C (n_22666), .Y(n_24702));
NAND2X1 g111847(.A (n_33546), .B (n_24687), .Y (n_24701));
NAND2X1 g108292(.A (n_23817), .B (n_9431), .Y (n_24700));
NAND2X1 g111853(.A (n_33546), .B (n_24668), .Y (n_24699));
NAND2X1 g111858(.A (n_33546), .B (n_24647), .Y (n_24698));
NAND2X1 g111862(.A (n_33546), .B (n_24661), .Y (n_24697));
OAI21X1 g111865(.A0 (n_23622), .A1 (n_22637), .B0 (n_24695), .Y(n_24696));
NAND2X1 g111867(.A (n_27614), .B (n_24614), .Y (n_24694));
NOR2X1 g111911(.A (n_23897), .B (n_14598), .Y (n_24693));
NAND2X1 g111914(.A (n_24259), .B (n_18982), .Y (n_24692));
NAND2X1 g111920(.A (n_32358), .B (n_18960), .Y (n_35280));
NAND2X1 g108331(.A (n_23816), .B (n_9431), .Y (n_24689));
NAND2X1 g111926(.A (n_24687), .B (n_24629), .Y (n_24688));
NAND2X1 g111927(.A (n_24687), .B (n_25968), .Y (n_24686));
AOI21X1 g111928(.A0 (n_23598), .A1 (n_27388), .B0 (n_8065), .Y(n_24685));
INVX1 g111929(.A (n_34810), .Y (n_24684));
NAND2X1 g111943(.A (n_24677), .B (n_18399), .Y (n_24682));
NAND2X1 g111948(.A (n_24663), .B (n_25554), .Y (n_24681));
NAND2X1 g111950(.A (n_23903), .B (n_8641), .Y (n_24680));
NAND2X1 g111958(.A (n_24670), .B (n_18918), .Y (n_24679));
NAND2X1 g111960(.A (n_24677), .B (n_26412), .Y (n_24678));
AOI21X1 g111969(.A0 (n_23596), .A1 (n_24675), .B0 (n_8065), .Y(n_24676));
AOI21X1 g111972(.A0 (n_23594), .A1 (n_24673), .B0 (n_8065), .Y(n_24674));
NAND2X1 g111981(.A (n_24677), .B (n_32798), .Y (n_24672));
NAND2X1 g111982(.A (n_24670), .B (n_32764), .Y (n_24671));
NAND2X1 g111985(.A (n_24668), .B (n_30180), .Y (n_24669));
NAND2X1 g111986(.A (n_24668), .B (n_30668), .Y (n_24667));
NAND2X1 g111993(.A (n_23902), .B (n_8303), .Y (n_24666));
NAND2X1 g111999(.A (n_24657), .B (n_24361), .Y (n_24665));
NAND2X1 g112004(.A (n_24663), .B (n_23192), .Y (n_24664));
NAND2X1 g112005(.A (n_24661), .B (n_25968), .Y (n_24662));
NAND2X1 g112006(.A (n_24175), .B (n_27770), .Y (n_24660));
NAND2X1 g112007(.A (n_23900), .B (n_8641), .Y (n_24659));
NAND2X1 g112012(.A (n_24657), .B (n_26637), .Y (n_24658));
NAND2X1 g112019(.A (n_24677), .B (n_25402), .Y (n_24656));
NAND2X1 g112020(.A (n_24670), .B (n_26866), .Y (n_24655));
AOI21X1 g112033(.A0 (n_23585), .A1 (n_27068), .B0 (n_8065), .Y(n_24654));
NAND2X1 g112034(.A (n_24670), .B (n_24652), .Y (n_24653));
NAND2X1 g112035(.A (n_24663), .B (n_18137), .Y (n_24651));
NAND2X1 g112036(.A (n_23907), .B (n_8303), .Y (n_24650));
NAND2X1 g112044(.A (n_23899), .B (n_25942), .Y (n_24649));
AND2X1 g112048(.A (n_24647), .B (n_24629), .Y (n_24648));
NAND2X1 g112049(.A (n_24647), .B (n_28431), .Y (n_24646));
NAND2X1 g112060(.A (n_23921), .B (n_20257), .Y (n_24645));
NAND2X1 g112061(.A (n_23920), .B (n_20258), .Y (n_24644));
INVX1 g112075(.A (n_24643), .Y (n_24972));
NAND2X1 g112078(.A (n_24199), .B (n_18987), .Y (n_24642));
NAND2X1 g112079(.A (n_24640), .B (n_18332), .Y (n_24641));
NAND2X1 g112088(.A (n_24628), .B (n_18262), .Y (n_24639));
NAND2X1 g112091(.A (n_24621), .B (n_24965), .Y (n_25378));
NAND2X1 g112096(.A (n_23967), .B (n_20290), .Y (n_24638));
INVX1 g112100(.A (n_34860), .Y (n_24960));
NAND2X1 g112106(.A (n_24214), .B (n_18979), .Y (n_32243));
NAND2X1 g112108(.A (n_23941), .B (n_17748), .Y (n_32922));
NAND2X1 g112110(.A (n_23986), .B (n_18977), .Y (n_35921));
NAND2X1 g112111(.A (n_33615), .B (n_17747), .Y (n_24633));
NAND2X1 g112119(.A (n_8990), .B (n_24631), .Y (n_24632));
NAND2X1 g112120(.A (n_23996), .B (n_24210), .Y (n_25390));
NAND2X1 g112123(.A (n_24661), .B (n_24629), .Y (n_24630));
NAND2X1 g112125(.A (n_24628), .B (n_35744), .Y (n_25384));
NOR2X1 g112129(.A (n_23924), .B (n_23551), .Y (n_24627));
NAND2X1 g112138(.A (n_24610), .B (n_33738), .Y (n_24626));
NAND2X1 g112139(.A (n_24623), .B (n_8990), .Y (n_24625));
NAND2X1 g112141(.A (n_24623), .B (n_27522), .Y (n_24624));
NAND2X1 g112148(.A (n_24621), .B (n_35790), .Y (n_24622));
NAND2X1 g112151(.A (n_24663), .B (n_25605), .Y (n_24620));
NAND2X1 g112152(.A (n_23898), .B (n_25220), .Y (n_24619));
NAND2X1 g112165(.A (n_24617), .B (n_29505), .Y (n_24618));
NAND2X1 g112166(.A (n_24617), .B (n_29430), .Y (n_24616));
NAND2X1 g112176(.A (n_24925), .B (n_24614), .Y (n_24615));
NAND2X2 g112179(.A (n_24612), .B (n_24002), .Y (n_24613));
NAND2X1 g112185(.A (n_24610), .B (n_28374), .Y (n_24611));
NAND2X1 g112188(.A (n_24610), .B (n_28158), .Y (n_24609));
AOI21X1 g112191(.A0 (n_24283), .A1 (n_29027), .B0 (n_22453), .Y(n_24608));
NAND2X1 g112195(.A (n_23636), .B (n_28136), .Y (n_24607));
NAND2X1 g112199(.A (n_24192), .B (n_33738), .Y (n_24606));
NOR2X1 g112201(.A (n_24604), .B (n_25881), .Y (n_24605));
NAND2X1 g112204(.A (n_24600), .B (n_30636), .Y (n_24603));
NAND2X1 g112215(.A (n_24621), .B (n_35528), .Y (n_25388));
NAND2X1 g112223(.A (n_24621), .B (n_25599), .Y (n_24602));
NAND2X1 g112229(.A (n_24628), .B (n_25877), .Y (n_25386));
NAND2X1 g112230(.A (n_24600), .B (n_29405), .Y (n_24601));
NAND2X1 g112233(.A (n_24600), .B (n_33738), .Y (n_24599));
NAND2X1 g112237(.A (n_23909), .B (n_19721), .Y (n_32277));
AOI21X1 g112245(.A0 (n_23541), .A1 (n_23771), .B0 (n_15155), .Y(n_24597));
AOI21X1 g112247(.A0 (n_23528), .A1 (n_23771), .B0 (n_15190), .Y(n_24595));
AOI21X1 g112250(.A0 (n_23546), .A1 (n_25942), .B0 (n_14789), .Y(n_24594));
AOI21X1 g112252(.A0 (n_24579), .A1 (n_24361), .B0 (n_14593), .Y(n_24593));
AOI21X1 g112253(.A0 (n_24242), .A1 (n_24361), .B0 (n_22477), .Y(n_24592));
AOI21X1 g112261(.A0 (n_14805), .A1 (n_24198), .B0 (n_8927), .Y(n_24590));
AOI21X1 g112262(.A0 (n_14835), .A1 (n_24216), .B0 (n_8927), .Y(n_24589));
NAND2X1 g112271(.A (n_23943), .B (n_27522), .Y (n_24588));
NAND2X1 g112282(.A (n_23949), .B (n_24012), .Y (n_25429));
INVX1 g112287(.A (n_34515), .Y (n_24901));
NOR2X1 g112295(.A (n_23619), .B (n_23965), .Y (n_24586));
NAND2X1 g112296(.A (n_23968), .B (n_23689), .Y (n_24585));
OAI21X1 g112297(.A0 (n_23517), .A1 (n_23178), .B0 (n_26208), .Y(n_24584));
NAND2X1 g112299(.A (n_23957), .B (n_26203), .Y (n_24583));
OAI21X1 g112301(.A0 (n_23517), .A1 (n_32654), .B0 (n_26199), .Y(n_24582));
NAND2X1 g112303(.A (n_23951), .B (n_34690), .Y (n_24581));
AOI21X1 g112305(.A0 (n_24579), .A1 (n_20178), .B0 (n_13883), .Y(n_24580));
NAND2X1 g112320(.A (n_23958), .B (n_24007), .Y (n_25437));
NAND2X1 g112336(.A (n_23956), .B (n_23242), .Y (n_25435));
INVX1 g112341(.A (n_25131), .Y (n_24578));
NAND2X1 g112363(.A (n_23954), .B (n_24006), .Y (n_25433));
NAND2X1 g112367(.A (n_23953), .B (n_24005), .Y (n_25431));
AOI21X1 g112372(.A0 (n_14327), .A1 (n_22821), .B0 (n_23952), .Y(n_24577));
AOI21X1 g112406(.A0 (n_23407), .A1 (n_26553), .B0 (n_23936), .Y(n_24576));
NAND2X1 g112420(.A (n_23933), .B (n_27842), .Y (n_24575));
NAND2X1 g112422(.A (n_23946), .B (n_24060), .Y (n_25835));
OAI21X1 g112424(.A0 (n_23034), .A1 (n_23519), .B0 (n_24042), .Y(n_25381));
NAND2X1 g112426(.A (n_23972), .B (n_23722), .Y (n_24574));
NAND2X1 g112427(.A (n_23971), .B (n_23711), .Y (n_24573));
NAND2X1 g112428(.A (n_23969), .B (n_23702), .Y (n_24572));
AOI21X1 g112430(.A0 (n_23555), .A1 (n_25220), .B0 (n_14328), .Y(n_24571));
NAND3X1 g112435(.A (n_23858), .B (n_32304), .C (n_21787), .Y(n_32210));
MX2X1 g112448(.A (n_19094), .B (n_19093), .S0 (n_23610), .Y(n_24569));
MX2X1 g112449(.A (n_20242), .B (n_19549), .S0 (n_23538), .Y(n_25414));
MX2X1 g112450(.A (n_20200), .B (n_20201), .S0 (n_23550), .Y(n_25412));
INVX1 g112472(.A (n_25085), .Y (n_24566));
MX2X1 g112474(.A (n_19050), .B (n_21742), .S0 (n_23611), .Y(n_25409));
NAND2X1 g112488(.A (n_24563), .B (n_24555), .Y (n_24565));
NAND2X1 g112491(.A (n_24563), .B (n_24546), .Y (n_24564));
NOR2X1 g112493(.A (n_11118), .B (n_23850), .Y (n_24562));
NAND2X1 g112497(.A (n_24563), .B (n_24537), .Y (n_24561));
NAND2X1 g112500(.A (n_24563), .B (n_24528), .Y (n_24560));
NOR2X1 g112502(.A (n_19114), .B (n_23849), .Y (n_24559));
NAND2X1 g112505(.A (n_22593), .B (n_23871), .Y (n_24874));
NAND3X1 g112548(.A (n_23859), .B (n_22384), .C (n_19843), .Y(n_24558));
NAND2X1 g112567(.A (n_23866), .B (n_19506), .Y (n_24557));
NAND2X1 g112588(.A (n_24555), .B (n_24526), .Y (n_24556));
NAND2X1 g112590(.A (n_24555), .B (n_28798), .Y (n_24554));
NAND2X1 g112601(.A (n_24542), .B (n_26412), .Y (n_24553));
NAND2X1 g112604(.A (n_24548), .B (n_18384), .Y (n_24552));
NAND2X1 g112605(.A (n_24539), .B (n_25003), .Y (n_24550));
NAND2X1 g112616(.A (n_24548), .B (n_24652), .Y (n_24549));
NAND2X1 g112622(.A (n_24546), .B (n_26106), .Y (n_24547));
NAND2X1 g112623(.A (n_24546), .B (n_25756), .Y (n_24545));
NAND2X1 g112632(.A (n_24542), .B (n_32764), .Y (n_24543));
NAND2X1 g112635(.A (n_24539), .B (n_32685), .Y (n_24540));
AND2X1 g112649(.A (n_24537), .B (n_26213), .Y (n_24538));
NAND2X1 g112650(.A (n_24537), .B (n_34753), .Y (n_24535));
NAND2X1 g112659(.A (n_24542), .B (n_13582), .Y (n_24534));
NAND2X1 g112663(.A (n_24548), .B (n_13582), .Y (n_24532));
NAND2X1 g112665(.A (n_24539), .B (n_26866), .Y (n_24531));
AOI21X1 g112669(.A0 (n_23507), .A1 (n_26197), .B0 (n_8065), .Y(n_24530));
AND2X1 g112681(.A (n_24528), .B (n_26213), .Y (n_24529));
NAND2X1 g112682(.A (n_24528), .B (n_24526), .Y (n_24527));
NAND3X1 g112700(.A (n_23463), .B (n_23505), .C (n_22942), .Y(n_25285));
INVX1 g112702(.A (n_24524), .Y (n_24525));
NAND2X1 g112768(.A (n_24539), .B (n_34499), .Y (n_24523));
INVX1 g112776(.A (n_35036), .Y (n_24521));
INVX1 g112785(.A (n_33911), .Y (n_24519));
NAND2X1 g112788(.A (n_24125), .B (n_18374), .Y (n_24518));
NOR2X1 g112800(.A (n_10244), .B (n_23851), .Y (n_24517));
NOR2X1 g112808(.A (n_8715), .B (n_23886), .Y (n_24516));
NAND2X1 g112816(.A (n_23861), .B (n_23029), .Y (n_35638));
NOR2X1 g112825(.A (n_10149), .B (n_23848), .Y (n_24514));
NAND3X1 g112830(.A (n_9049), .B (n_23504), .C (n_19861), .Y(n_24513));
NOR2X1 g112831(.A (n_8909), .B (n_23885), .Y (n_24512));
NOR2X1 g112834(.A (n_23887), .B (n_23293), .Y (n_24511));
NAND2X1 g112843(.A (n_23878), .B (n_26791), .Y (n_24510));
OAI21X1 g112873(.A0 (n_23480), .A1 (n_19330), .B0 (n_24508), .Y(n_24509));
NAND2X1 g112889(.A (n_23873), .B (n_26787), .Y (n_24507));
OAI21X1 g112899(.A0 (n_23480), .A1 (n_13317), .B0 (n_24505), .Y(n_24506));
NAND2X1 g112928(.A (n_23880), .B (n_27222), .Y (n_24503));
INVX1 g112938(.A (n_24942), .Y (n_24502));
INVX1 g112942(.A (n_24944), .Y (n_24501));
NAND4X1 g112976(.A (n_23838), .B (n_22558), .C (n_22919), .D(n_22876), .Y (n_24500));
NAND2X2 g112978(.A (n_23867), .B (n_23565), .Y (n_25298));
INVX1 g112981(.A (n_24998), .Y (n_24499));
INVX1 g112986(.A (n_24987), .Y (n_24498));
INVX1 g112989(.A (n_24497), .Y (n_25305));
XOR2X1 g113001(.A (n_19710), .B (n_23515), .Y (n_25293));
MX2X1 g113015(.A (n_19288), .B (n_19287), .S0 (n_23514), .Y(n_24495));
INVX1 g113017(.A (n_24494), .Y (n_24833));
INVX1 g113025(.A (n_24985), .Y (n_24493));
NAND3X1 g113056(.A (n_18568), .B (n_23473), .C (n_22333), .Y(n_24492));
NAND3X1 g113282(.A (n_22865), .B (n_23468), .C (n_23467), .Y(n_24491));
NAND4X1 g113328(.A (n_23837), .B (n_33365), .C (n_24490), .D(n_18924), .Y (n_25251));
INVX1 g113387(.A (n_24859), .Y (n_24489));
NAND2X2 g113487(.A (n_32279), .B (n_32280), .Y (n_25248));
NAND2X1 g113503(.A (n_23821), .B (n_31781), .Y (n_24488));
NOR2X1 g113541(.A (n_10366), .B (n_23826), .Y (n_24487));
NOR2X1 g113553(.A (n_9894), .B (n_23827), .Y (n_24486));
OAI21X1 g113694(.A0 (n_9882), .A1 (n_24484), .B0 (n_23825), .Y(n_24485));
OAI21X1 g113695(.A0 (n_9838), .A1 (n_24484), .B0 (n_23824), .Y(n_24483));
NAND4X1 g113759(.A (n_23822), .B (n_22949), .C (n_22638), .D(n_22947), .Y (n_24482));
NOR2X1 g113766(.A (n_9905), .B (n_23823), .Y (n_24481));
NAND2X1 g109405(.A (n_24106), .B (n_28213), .Y (n_24480));
NAND2X1 g109406(.A (n_24104), .B (n_28204), .Y (n_24479));
NAND2X1 g109408(.A (n_24102), .B (n_28195), .Y (n_24478));
OAI21X1 g109893(.A0 (n_14972), .A1 (n_9458), .B0 (n_23806), .Y(n_24477));
OAI21X1 g110043(.A0 (n_15092), .A1 (n_9458), .B0 (n_23804), .Y(n_24476));
NOR2X1 g110264(.A (n_23445), .B (n_23662), .Y (n_24474));
NAND2X1 g110434(.A (n_23785), .B (n_25942), .Y (n_24473));
NAND2X1 g110517(.A (n_23783), .B (n_9431), .Y (n_24472));
NAND2X1 g110660(.A (n_23782), .B (n_9431), .Y (n_24471));
NAND3X1 g110708(.A (n_18564), .B (n_20472), .C (n_23438), .Y(n_24470));
AOI21X1 g110817(.A0 (n_23436), .A1 (n_25942), .B0 (n_14711), .Y(n_24469));
NAND2X1 g110822(.A (n_23792), .B (n_28570), .Y (n_24468));
AOI21X1 g110839(.A0 (n_23434), .A1 (n_25220), .B0 (n_14471), .Y(n_24467));
NAND2X1 g110851(.A (n_23799), .B (n_13662), .Y (n_24466));
NAND2X1 g110853(.A (n_23797), .B (n_28554), .Y (n_24465));
NAND2X1 g110855(.A (n_23795), .B (n_28549), .Y (n_24464));
NAND2X1 g111023(.A (n_23798), .B (n_25704), .Y (n_24463));
NAND2X1 g111029(.A (n_23794), .B (n_25690), .Y (n_24462));
NAND2X1 g111034(.A (n_23790), .B (n_25683), .Y (n_24461));
NAND2X1 g111053(.A (n_23788), .B (n_25681), .Y (n_24460));
AOI21X1 g111068(.A0 (n_23435), .A1 (n_25220), .B0 (n_14462), .Y(n_24459));
NAND2X1 g111107(.A (n_23759), .B (n_23624), .Y (n_24458));
NAND4X1 g111199(.A (n_15028), .B (n_22769), .C (n_23068), .D(n_22770), .Y (n_24457));
NAND2X1 g111210(.A (n_23751), .B (n_25122), .Y (n_35108));
NAND2X1 g111213(.A (n_23744), .B (n_9431), .Y (n_24455));
NAND2X1 g111219(.A (n_24447), .B (n_23725), .Y (n_24454));
NAND2X1 g111229(.A (n_23746), .B (n_26458), .Y (n_24453));
NAND2X1 g111252(.A (n_23743), .B (n_24451), .Y (n_24452));
NAND2X1 g111264(.A (n_23750), .B (n_25122), .Y (n_32120));
NAND2X1 g111265(.A (n_24441), .B (n_25554), .Y (n_24449));
NAND2X1 g111267(.A (n_24447), .B (n_24446), .Y (n_24448));
AOI21X1 g111297(.A0 (n_23432), .A1 (n_22749), .B0 (n_31523), .Y(n_24445));
NAND2X1 g111304(.A (n_23749), .B (n_25111), .Y (n_24444));
NAND2X1 g111346(.A (n_23748), .B (n_25111), .Y (n_24443));
NAND2X1 g111347(.A (n_24441), .B (n_35054), .Y (n_24442));
NAND2X1 g111350(.A (n_24447), .B (n_23696), .Y (n_24440));
NAND2X1 g111358(.A (n_23745), .B (n_9431), .Y (n_24439));
NAND2X1 g111376(.A (n_24441), .B (n_23578), .Y (n_24438));
NAND2X1 g111453(.A (n_24441), .B (n_25207), .Y (n_24437));
NAND4X1 g111465(.A (n_15178), .B (n_22062), .C (n_23092), .D(n_22789), .Y (n_24436));
NAND4X1 g111466(.A (n_15177), .B (n_22057), .C (n_23087), .D(n_22788), .Y (n_24435));
AOI21X1 g111472(.A0 (n_27743), .A1 (n_24073), .B0 (n_10875), .Y(n_24434));
NAND4X1 g111482(.A (n_14875), .B (n_22774), .C (n_23075), .D(n_22772), .Y (n_24433));
OAI21X1 g111504(.A0 (n_14408), .A1 (n_26801), .B0 (n_23774), .Y(n_24432));
NAND4X1 g111522(.A (n_23160), .B (n_18734), .C (n_23121), .D(n_22808), .Y (n_24431));
NAND2X1 g111524(.A (n_23760), .B (n_26569), .Y (n_24430));
NAND4X1 g111525(.A (n_23159), .B (n_19274), .C (n_23119), .D(n_22806), .Y (n_24429));
NAND4X1 g111528(.A (n_21444), .B (n_21823), .C (n_20487), .D(n_23054), .Y (n_24428));
OAI21X1 g111538(.A0 (n_13801), .A1 (n_29968), .B0 (n_23758), .Y(n_24427));
OAI21X1 g111545(.A0 (n_14867), .A1 (n_8614), .B0 (n_23757), .Y(n_24426));
NAND2X1 g111546(.A (n_23775), .B (n_26564), .Y (n_24425));
NAND2X1 g111547(.A (n_23770), .B (n_14128), .Y (n_24424));
AOI21X1 g111557(.A0 (n_27743), .A1 (n_24071), .B0 (n_20089), .Y(n_24422));
AOI21X1 g111683(.A0 (n_24041), .A1 (n_15031), .B0 (n_23138), .Y(n_24421));
OAI21X1 g111722(.A0 (n_14863), .A1 (n_8614), .B0 (n_23761), .Y(n_24420));
XOR2X1 g111778(.A (n_20175), .B (n_23428), .Y (n_25201));
AOI21X1 g111782(.A0 (n_33288), .A1 (n_29411), .B0 (n_18835), .Y(n_24419));
OAI21X1 g111823(.A0 (n_23779), .A1 (n_23778), .B0 (n_23780), .Y(n_25205));
XOR2X1 g111826(.A (n_16400), .B (n_23386), .Y (n_25199));
NOR2X1 g111833(.A (n_23644), .B (n_23645), .Y (n_24418));
AOI21X1 g111836(.A0 (n_10409), .A1 (n_23341), .B0 (n_16415), .Y(n_24417));
NAND2X1 g111838(.A (n_23683), .B (n_23020), .Y (n_24416));
INVX1 g111839(.A (n_34604), .Y (n_24415));
NAND2X1 g111848(.A (n_33546), .B (n_24390), .Y (n_24413));
NAND2X1 g111854(.A (n_33546), .B (n_24378), .Y (n_24412));
NAND2X1 g111859(.A (n_33546), .B (n_24365), .Y (n_24411));
NAND2X1 g111863(.A (n_33546), .B (n_24352), .Y (n_24410));
NAND3X1 g111868(.A (n_23366), .B (n_23359), .C (n_19278), .Y(n_24409));
NAND3X1 g111869(.A (n_23926), .B (n_22552), .C (n_22573), .Y(n_32239));
NAND2X1 g111872(.A (n_9503), .B (n_24395), .Y (n_24407));
NAND2X1 g111877(.A (n_24404), .B (n_34709), .Y (n_24405));
NAND2X1 g111882(.A (n_24401), .B (n_28926), .Y (n_24402));
NAND2X1 g111887(.A (n_24399), .B (n_34709), .Y (n_24400));
NAND2X1 g111891(.A (n_24404), .B (n_29199), .Y (n_24398));
NAND2X1 g111898(.A (n_24401), .B (n_25980), .Y (n_24397));
NAND2X1 g111901(.A (n_24395), .B (n_28013), .Y (n_24396));
NAND2X1 g111906(.A (n_24399), .B (n_29199), .Y (n_24394));
NAND2X1 g111915(.A (n_23652), .B (n_25228), .Y (n_24393));
NAND2X1 g111919(.A (n_32359), .B (n_18961), .Y (n_35279));
NAND2X1 g111931(.A (n_24390), .B (n_28890), .Y (n_24391));
NAND2X1 g111932(.A (n_24390), .B (n_30180), .Y (n_24389));
NAND3X1 g111935(.A (n_22859), .B (n_23351), .C (n_22753), .Y(n_24388));
NAND2X1 g111938(.A (n_24374), .B (n_24386), .Y (n_24387));
NAND2X1 g111939(.A (n_24372), .B (n_24386), .Y (n_24385));
OR2X1 g111941(.A (n_24383), .B (n_25054), .Y (n_24384));
NAND2X1 g111963(.A (n_24369), .B (n_28441), .Y (n_24382));
NAND2X1 g111968(.A (n_23651), .B (n_25228), .Y (n_24381));
AOI21X1 g111976(.A0 (n_9629), .A1 (n_19007), .B0 (n_23730), .Y(n_24380));
AND2X1 g111987(.A (n_24378), .B (n_27993), .Y (n_24379));
NAND2X1 g111989(.A (n_24378), .B (n_30668), .Y (n_24377));
NAND2X1 g111991(.A (n_23650), .B (n_25228), .Y (n_24376));
NAND2X1 g111994(.A (n_24374), .B (n_26315), .Y (n_24375));
NAND2X1 g111996(.A (n_24372), .B (n_17713), .Y (n_24373));
NAND2X1 g112027(.A (n_24369), .B (n_24361), .Y (n_24370));
NAND2X1 g112032(.A (n_23649), .B (n_25228), .Y (n_24368));
NAND2X1 g112041(.A (n_23894), .B (n_27950), .Y (n_24367));
AND2X1 g112050(.A (n_24365), .B (n_27993), .Y (n_24366));
NAND2X1 g112051(.A (n_24365), .B (n_28431), .Y (n_24364));
NAND2X1 g112056(.A (n_24374), .B (n_24361), .Y (n_24363));
NAND2X1 g112057(.A (n_24372), .B (n_24361), .Y (n_24362));
NAND2X1 g112067(.A (n_24369), .B (n_23578), .Y (n_24360));
NAND2X1 g112076(.A (n_23684), .B (n_22894), .Y (n_24643));
OR2X1 g112083(.A (n_33555), .B (n_13432), .Y (n_24359));
NAND2X1 g112095(.A (n_23658), .B (n_19770), .Y (n_24358));
NAND2X1 g112097(.A (n_23966), .B (n_20291), .Y (n_24357));
NAND2X1 g112107(.A (n_23940), .B (n_20211), .Y (n_32923));
NAND2X1 g112109(.A (n_23985), .B (n_18976), .Y (n_35922));
NAND3X1 g112115(.A (n_23385), .B (n_23318), .C (n_19935), .Y(n_24354));
NAND2X1 g112122(.A (n_24345), .B (n_24965), .Y (n_25079));
NAND2X1 g112127(.A (n_24352), .B (n_30180), .Y (n_24353));
NAND2X1 g112128(.A (n_24352), .B (n_28890), .Y (n_24351));
NAND2X1 g112132(.A (n_24374), .B (n_23329), .Y (n_24350));
NAND2X1 g112133(.A (n_24372), .B (n_24348), .Y (n_24349));
NAND2X1 g112135(.A (n_24341), .B (n_33738), .Y (n_24347));
NAND2X1 g112167(.A (n_24345), .B (n_35794), .Y (n_24346));
NAND2X1 g112169(.A (n_24369), .B (n_25605), .Y (n_24344));
OR2X1 g112180(.A (n_33555), .B (n_17287), .Y (n_24343));
NAND2X1 g112186(.A (n_24341), .B (n_28158), .Y (n_24342));
NAND2X1 g112187(.A (n_24341), .B (n_28374), .Y (n_24340));
NAND2X1 g112197(.A (n_23905), .B (n_33738), .Y (n_24339));
NAND2X1 g112200(.A (n_24331), .B (n_26238), .Y (n_24338));
NOR2X1 g112203(.A (n_24336), .B (n_25881), .Y (n_24337));
AOI21X1 g112206(.A0 (n_21174), .A1 (n_23771), .B0 (n_23634), .Y(n_24335));
AOI21X1 g112207(.A0 (n_21172), .A1 (n_25122), .B0 (n_23633), .Y(n_24334));
NAND2X1 g112209(.A (n_24345), .B (n_35457), .Y (n_25081));
NAND2X1 g112226(.A (n_24345), .B (n_25599), .Y (n_24333));
NAND2X1 g112227(.A (n_24331), .B (n_29405), .Y (n_24332));
NAND2X1 g112228(.A (n_24331), .B (n_33738), .Y (n_24330));
NAND3X1 g112234(.A (n_22242), .B (n_23032), .C (n_23247), .Y(n_24329));
NAND2X1 g112236(.A (n_33710), .B (n_19722), .Y (n_32278));
NAND2X1 g112241(.A (n_21746), .B (n_23912), .Y (n_32039));
NAND4X1 g112256(.A (n_21021), .B (n_22286), .C (n_22491), .D(n_22963), .Y (n_24326));
AOI21X1 g112263(.A0 (n_14883), .A1 (n_23929), .B0 (n_22762), .Y(n_24325));
NAND2X1 g112278(.A (n_23698), .B (n_24324), .Y (n_25140));
NAND2X1 g112280(.A (n_23697), .B (n_26929), .Y (n_24323));
NAND3X1 g112289(.A (n_20365), .B (n_23560), .C (n_19694), .Y(n_32881));
OAI21X1 g112304(.A0 (n_24301), .A1 (n_13183), .B0 (n_13175), .Y(n_24321));
AND2X1 g112308(.A (n_23685), .B (n_18222), .Y (n_24318));
AOI21X1 g112310(.A0 (n_23980), .A1 (n_34952), .B0 (n_15138), .Y(n_32136));
AOI21X1 g112311(.A0 (n_23977), .A1 (n_26162), .B0 (n_15133), .Y(n_32063));
NAND2X1 g112314(.A (n_23726), .B (n_26925), .Y (n_24314));
INVX1 g112315(.A (n_24788), .Y (n_24313));
OAI21X1 g112317(.A0 (n_24307), .A1 (n_24312), .B0 (n_24009), .Y(n_25136));
NAND2X1 g112322(.A (n_23717), .B (n_22441), .Y (n_25142));
NAND2X1 g112334(.A (n_23716), .B (n_26924), .Y (n_24311));
OAI21X1 g112342(.A0 (n_23294), .A1 (n_32748), .B0 (n_24309), .Y(n_25131));
OAI21X1 g112365(.A0 (n_23297), .A1 (n_32812), .B0 (n_26923), .Y(n_24308));
OAI21X1 g112383(.A0 (n_24307), .A1 (n_13653), .B0 (n_24003), .Y(n_25127));
OAI21X1 g112384(.A0 (n_23304), .A1 (n_10517), .B0 (n_18206), .Y(n_24306));
NAND2X1 g112387(.A (n_23706), .B (n_24305), .Y (n_25138));
INVX1 g112397(.A (n_24743), .Y (n_24304));
AOI21X1 g112400(.A0 (n_23934), .A1 (n_14612), .B0 (n_29725), .Y(n_24303));
OAI21X1 g112402(.A0 (n_24301), .A1 (n_19330), .B0 (n_27716), .Y(n_24302));
OAI21X1 g112403(.A0 (n_24301), .A1 (n_14430), .B0 (n_24299), .Y(n_24300));
NAND2X1 g112405(.A (n_23663), .B (n_13180), .Y (n_24298));
INVX1 g112407(.A (n_24737), .Y (n_24297));
NOR2X1 g112413(.A (n_23056), .B (n_23627), .Y (n_24296));
NAND2X1 g112419(.A (n_23681), .B (n_26548), .Y (n_24295));
OAI21X1 g112431(.A0 (n_18213), .A1 (n_25540), .B0 (n_23669), .Y(n_24294));
OAI21X1 g112432(.A0 (n_23035), .A1 (n_29725), .B0 (n_23672), .Y(n_24293));
OAI21X1 g112462(.A0 (n_23694), .A1 (n_23693), .B0 (n_23695), .Y(n_25109));
MX2X1 g112463(.A (n_21736), .B (n_20268), .S0 (n_23358), .Y(n_25106));
INVX1 g112466(.A (n_24292), .Y (n_25073));
INVX1 g112469(.A (n_24291), .Y (n_24567));
NAND2X1 g112471(.A (n_23679), .B (n_23411), .Y (n_25094));
NAND2X2 g112473(.A (n_23678), .B (n_23410), .Y (n_25085));
NAND2X1 g112485(.A (n_23559), .B (n_17150), .Y (n_24290));
OAI21X1 g112510(.A0 (n_21461), .A1 (n_22879), .B0 (n_23561), .Y(n_24289));
NAND2X1 g112511(.A (n_23524), .B (n_23260), .Y (n_24288));
NAND2X1 g112513(.A (n_24280), .B (n_28864), .Y (n_24287));
NAND2X1 g112516(.A (n_24278), .B (n_29061), .Y (n_24286));
NAND2X1 g112518(.A (n_24274), .B (n_25988), .Y (n_24285));
NAND2X1 g112520(.A (n_24283), .B (n_27340), .Y (n_24284));
NAND2X1 g112523(.A (n_24271), .B (n_30563), .Y (n_24282));
NAND2X1 g112526(.A (n_24280), .B (n_28485), .Y (n_24281));
NAND2X1 g112529(.A (n_24278), .B (n_28485), .Y (n_24279));
NAND2X1 g112532(.A (n_24262), .B (n_28926), .Y (n_24277));
NAND3X1 g112533(.A (n_22712), .B (n_23287), .C (n_22752), .Y(n_24276));
NAND2X1 g112534(.A (n_26978), .B (n_24274), .Y (n_24275));
NAND2X1 g112536(.A (n_24283), .B (n_29604), .Y (n_24273));
NAND2X1 g112540(.A (n_24271), .B (n_26535), .Y (n_24272));
NAND3X1 g112542(.A (n_22703), .B (n_23285), .C (n_22750), .Y(n_24270));
NAND2X1 g112543(.A (n_26978), .B (n_24233), .Y (n_24269));
NAND2X1 g112546(.A (n_24280), .B (n_30197), .Y (n_24268));
NAND2X1 g112550(.A (n_24278), .B (n_26535), .Y (n_24267));
NAND3X1 g112552(.A (n_22692), .B (n_23283), .C (n_22747), .Y(n_24266));
NAND2X1 g112553(.A (n_26978), .B (n_24225), .Y (n_24265));
NAND3X1 g112558(.A (n_22677), .B (n_23281), .C (n_22751), .Y(n_24264));
NAND2X1 g112559(.A (n_26978), .B (n_24262), .Y (n_24263));
NAND2X1 g112563(.A (n_23532), .B (n_8303), .Y (n_24261));
INVX1 g112564(.A (n_24259), .Y (n_24260));
NAND2X1 g112568(.A (n_23865), .B (n_19507), .Y (n_24258));
INVX1 g112569(.A (n_34765), .Y (n_24257));
NAND2X1 g112576(.A (n_23600), .B (n_20088), .Y (n_24255));
NAND2X1 g112580(.A (n_29551), .B (n_23061), .Y (n_24254));
NAND3X1 g112583(.A (n_23889), .B (n_34725), .C (n_22857), .Y(n_32568));
NAND2X1 g112585(.A (n_23548), .B (n_25942), .Y (n_24252));
NAND2X1 g112596(.A (n_24239), .B (n_24249), .Y (n_24251));
NAND2X1 g112602(.A (n_24237), .B (n_24249), .Y (n_24250));
NAND2X1 g112603(.A (n_23543), .B (n_24247), .Y (n_24248));
NAND2X1 g112610(.A (n_23531), .B (n_8303), .Y (n_24246));
NAND2X1 g112615(.A (n_26132), .B (n_23061), .Y (n_24245));
NAND2X1 g112617(.A (n_24242), .B (n_24105), .Y (n_24243));
NAND2X1 g112621(.A (n_24242), .B (n_34418), .Y (n_24241));
NAND2X1 g112630(.A (n_24239), .B (n_32728), .Y (n_24240));
NAND2X1 g112633(.A (n_24237), .B (n_32685), .Y (n_24238));
NAND2X1 g112637(.A (n_23847), .B (n_32777), .Y (n_24235));
NAND2X1 g112639(.A (n_24233), .B (n_26870), .Y (n_24234));
NAND2X1 g112641(.A (n_23530), .B (n_8303), .Y (n_24232));
NAND2X1 g112645(.A (n_24262), .B (n_26870), .Y (n_24230));
NAND2X1 g112660(.A (n_23844), .B (n_27470), .Y (n_24229));
NAND2X1 g112666(.A (n_23539), .B (n_24247), .Y (n_24228));
NAND2X1 g112668(.A (n_23536), .B (n_25228), .Y (n_24227));
NAND2X1 g112691(.A (n_24225), .B (n_26870), .Y (n_24226));
NAND2X1 g112695(.A (n_23518), .B (n_27770), .Y (n_24224));
NAND2X1 g112698(.A (n_23621), .B (n_19708), .Y (n_24223));
NAND3X1 g112701(.A (n_23210), .B (n_22746), .C (n_23234), .Y(n_24978));
NAND2X1 g112703(.A (n_23614), .B (n_22940), .Y (n_24524));
NAND2X1 g112705(.A (n_24579), .B (n_23578), .Y (n_24222));
INVX1 g112706(.A (n_24640), .Y (n_24221));
NAND2X1 g112711(.A (n_23554), .B (n_21769), .Y (n_24220));
NAND2X1 g112712(.A (n_24242), .B (n_23578), .Y (n_24219));
NAND3X1 g112715(.A (n_22510), .B (n_24178), .C (n_22875), .Y(n_24217));
NAND2X1 g112722(.A (n_24216), .B (n_33287), .Y (n_24924));
INVX1 g112728(.A (n_24214), .Y (n_24215));
INVX1 g112733(.A (n_33615), .Y (n_24213));
NAND2X1 g112742(.A (n_23635), .B (n_24207), .Y (n_24950));
NAND2X1 g112743(.A (n_23904), .B (n_24204), .Y (n_24947));
INVX1 g112746(.A (n_24210), .Y (n_24211));
NAND2X1 g112751(.A (n_23544), .B (n_25942), .Y (n_24209));
NAND2X1 g112766(.A (n_24207), .B (n_14603), .Y (n_24208));
NAND2X1 g112767(.A (n_24579), .B (n_23356), .Y (n_24206));
NAND2X1 g112771(.A (n_24204), .B (n_14624), .Y (n_24205));
NAND2X1 g112774(.A (n_23576), .B (n_18459), .Y (n_32916));
NAND2X1 g112775(.A (n_23526), .B (n_8303), .Y (n_24202));
INVX1 g112782(.A (n_24199), .Y (n_24200));
NAND2X1 g112792(.A (n_23130), .B (n_24198), .Y (n_24927));
NOR2X1 g112801(.A (n_8914), .B (n_23617), .Y (n_24197));
OAI21X1 g112811(.A0 (n_23237), .A1 (n_18441), .B0 (n_27399), .Y(n_24196));
NAND2X1 g112838(.A (n_23607), .B (n_27064), .Y (n_24195));
AND2X1 g112842(.A (n_23588), .B (n_27379), .Y (n_24194));
NAND2X1 g112861(.A (n_23273), .B (n_23589), .Y (n_24914));
INVX1 g112909(.A (n_24192), .Y (n_24917));
NAND2X1 g112922(.A (n_23605), .B (n_24190), .Y (n_24191));
NAND2X1 g112926(.A (n_23597), .B (n_27718), .Y (n_24189));
NAND2X1 g112934(.A (n_23587), .B (n_27710), .Y (n_24188));
NAND2X1 g112936(.A (n_23579), .B (n_27709), .Y (n_24187));
NAND2X1 g112939(.A (n_23556), .B (n_23935), .Y (n_24942));
INVX1 g112940(.A (n_24623), .Y (n_24186));
NAND2X1 g112943(.A (n_23557), .B (n_23666), .Y (n_24944));
NAND2X1 g112945(.A (n_23609), .B (n_23932), .Y (n_24989));
NAND2X1 g112947(.A (n_23566), .B (n_27705), .Y (n_24185));
NAND2X1 g112951(.A (n_23568), .B (n_23718), .Y (n_24932));
AOI21X1 g112954(.A0 (n_14512), .A1 (n_22821), .B0 (n_23584), .Y(n_24184));
AOI21X1 g112958(.A0 (n_23875), .A1 (n_33748), .B0 (n_17656), .Y(n_24182));
NAND4X1 g112977(.A (n_22991), .B (n_22497), .C (n_22916), .D(n_21908), .Y (n_24179));
XOR2X1 g112982(.A (n_22197), .B (n_24178), .Y (n_24998));
XOR2X1 g112987(.A (n_24177), .B (n_23261), .Y (n_24987));
XOR2X1 g112990(.A (n_19711), .B (n_23870), .Y (n_24497));
INVX1 g112996(.A (n_24175), .Y (n_25341));
XOR2X1 g112999(.A (n_19209), .B (n_23256), .Y (n_24993));
XOR2X1 g113000(.A (n_22194), .B (n_23253), .Y (n_24991));
NAND2X1 g113005(.A (n_23577), .B (n_23335), .Y (n_24940));
INVX1 g113009(.A (n_24174), .Y (n_24963));
MX2X1 g113018(.A (n_18689), .B (n_24173), .S0 (n_23251), .Y(n_24494));
NAND2X1 g113026(.A (n_23563), .B (n_23321), .Y (n_24985));
NOR2X1 g113049(.A (n_10860), .B (n_23488), .Y (n_24172));
NOR2X1 g113066(.A (n_22306), .B (n_23491), .Y (n_25257));
NAND2X1 g113078(.A (n_28597), .B (n_24159), .Y (n_24169));
NAND2X1 g113079(.A (n_29065), .B (n_24156), .Y (n_24168));
NAND2X1 g108852(.A (n_23812), .B (n_17639), .Y (n_24167));
NAND2X1 g113080(.A (n_34770), .B (n_24162), .Y (n_24166));
NAND2X1 g113081(.A (n_24164), .B (n_28926), .Y (n_24165));
NAND2X1 g113085(.A (n_24162), .B (n_25988), .Y (n_24163));
NAND2X1 g113086(.A (n_24164), .B (n_28013), .Y (n_24161));
NAND2X1 g113092(.A (n_24159), .B (n_29455), .Y (n_24160));
NOR2X1 g113094(.A (n_22336), .B (n_23481), .Y (n_24158));
NAND2X1 g113096(.A (n_24156), .B (n_28915), .Y (n_24157));
NAND2X1 g113101(.A (n_24162), .B (n_29455), .Y (n_24155));
AOI21X1 g113104(.A0 (n_13670), .A1 (n_14956), .B0 (n_23486), .Y(n_24154));
NAND2X1 g113123(.A (n_24149), .B (n_27091), .Y (n_24153));
NAND2X1 g113127(.A (n_24144), .B (n_25734), .Y (n_24152));
NAND2X1 g113129(.A (n_24146), .B (n_27091), .Y (n_24151));
NAND2X1 g113147(.A (n_24149), .B (n_26637), .Y (n_24150));
NAND2X1 g113162(.A (n_24149), .B (n_25554), .Y (n_24148));
NAND2X1 g113164(.A (n_24146), .B (n_18498), .Y (n_24147));
NAND2X1 g113165(.A (n_24144), .B (n_25554), .Y (n_24145));
NAND2X1 g108911(.A (n_23810), .B (n_25942), .Y (n_24143));
NAND2X1 g108916(.A (n_24130), .B (n_21919), .Y (n_24142));
NAND2X1 g113201(.A (n_24149), .B (n_22994), .Y (n_24141));
NAND2X1 g113202(.A (n_24146), .B (n_25956), .Y (n_24140));
NAND2X1 g113203(.A (n_24144), .B (n_22994), .Y (n_24139));
NAND2X1 g113217(.A (n_23494), .B (n_24137), .Y (n_24138));
NAND3X1 g113222(.A (n_22663), .B (n_23232), .C (n_18224), .Y(n_24136));
NAND2X1 g113241(.A (n_24146), .B (n_25193), .Y (n_24135));
NAND2X1 g113266(.A (n_24144), .B (n_26637), .Y (n_24134));
NAND2X1 g108953(.A (n_23809), .B (n_9431), .Y (n_24133));
NAND2X1 g108963(.A (n_24130), .B (n_23192), .Y (n_24131));
NOR2X1 g113319(.A (n_10126), .B (n_23484), .Y (n_24129));
NOR2X1 g113323(.A (n_10174), .B (n_23485), .Y (n_24128));
NAND2X1 g113349(.A (n_23506), .B (n_23045), .Y (n_24863));
OAI21X1 g113356(.A0 (n_26382), .A1 (n_21938), .B0 (n_23489), .Y(n_24127));
INVX1 g113363(.A (n_24125), .Y (n_24126));
NAND2X1 g108997(.A (n_23808), .B (n_9431), .Y (n_24124));
NAND2X1 g108998(.A (n_24130), .B (n_19597), .Y (n_24123));
NAND2X1 g113380(.A (n_23513), .B (n_23042), .Y (n_24868));
NAND2X1 g113388(.A (n_23511), .B (n_23040), .Y (n_24859));
NAND2X1 g113398(.A (n_23509), .B (n_23038), .Y (n_24865));
NAND2X1 g113415(.A (n_23512), .B (n_24121), .Y (n_24122));
OAI21X1 g113436(.A0 (n_19123), .A1 (n_25540), .B0 (n_23499), .Y(n_24120));
OAI21X1 g113440(.A0 (n_19121), .A1 (n_25540), .B0 (n_23495), .Y(n_24118));
OAI21X1 g113443(.A0 (n_23834), .A1 (n_28523), .B0 (n_22390), .Y(n_24117));
INVX1 g113455(.A (n_24548), .Y (n_24116));
INVX1 g113478(.A (n_24542), .Y (n_24113));
NOR2X1 g113500(.A (n_23231), .B (n_23199), .Y (n_24112));
NAND2X1 g109085(.A (n_23807), .B (n_25942), .Y (n_24111));
NAND2X1 g113727(.A (n_23472), .B (n_20323), .Y (n_24110));
NAND2X1 g113732(.A (n_23222), .B (n_28136), .Y (n_24109));
NAND4X1 g113760(.A (n_23470), .B (n_22361), .C (n_23476), .D(n_23477), .Y (n_24108));
NOR2X1 g109407(.A (n_23813), .B (n_14084), .Y (n_24107));
NAND2X1 g109652(.A (n_24103), .B (n_24105), .Y (n_24106));
NAND2X1 g109711(.A (n_24103), .B (n_35054), .Y (n_24104));
NAND2X1 g109824(.A (n_24103), .B (n_24101), .Y (n_24102));
INVX1 g110235(.A (n_24130), .Y (n_24100));
NAND4X1 g110262(.A (n_23186), .B (n_9601), .C (n_22418), .D(n_22718), .Y (n_24099));
OAI21X1 g110813(.A0 (n_14928), .A1 (n_9458), .B0 (n_23447), .Y(n_24098));
NAND2X1 g111217(.A (n_23437), .B (n_25082), .Y (n_24096));
NAND3X1 g111369(.A (n_18701), .B (n_23128), .C (n_21806), .Y(n_24095));
OAI21X1 g111516(.A0 (n_14880), .A1 (n_8614), .B0 (n_23442), .Y(n_24094));
AOI22X1 g111517(.A0 (n_14871), .A1 (n_14490), .B0 (n_23135), .B1(n_25111), .Y (n_24093));
OAI21X1 g111543(.A0 (n_14656), .A1 (n_9458), .B0 (n_23439), .Y(n_24092));
OAI21X1 g111633(.A0 (n_14644), .A1 (n_8614), .B0 (n_23441), .Y(n_24091));
OAI21X1 g111714(.A0 (n_23367), .A1 (n_35520), .B0 (n_24090), .Y(n_24804));
AOI21X1 g111718(.A0 (n_23142), .A1 (n_25220), .B0 (n_14429), .Y(n_24089));
OAI21X1 g111727(.A0 (n_23369), .A1 (n_35520), .B0 (n_24088), .Y(n_24820));
OAI21X1 g111747(.A0 (n_23370), .A1 (n_35520), .B0 (n_24086), .Y(n_24818));
AOI21X1 g111759(.A0 (n_23776), .A1 (n_29411), .B0 (n_19346), .Y(n_24085));
NAND2X1 g111834(.A (n_23387), .B (n_31345), .Y (n_24084));
AOI21X1 g111835(.A0 (n_9379), .A1 (n_23123), .B0 (n_30702), .Y(n_24083));
AOI21X1 g111841(.A0 (n_21850), .A1 (n_22907), .B0 (n_23372), .Y(n_24082));
NAND3X1 g111842(.A (n_23383), .B (n_23070), .C (n_19840), .Y(n_24081));
NAND2X1 g111850(.A (n_26756), .B (n_24062), .Y (n_24080));
NAND2X1 g111851(.A (n_26756), .B (n_24054), .Y (n_24079));
NAND2X1 g111856(.A (n_26756), .B (n_24051), .Y (n_24078));
NAND2X1 g111857(.A (n_26756), .B (n_24047), .Y (n_24077));
NAND2X1 g111880(.A (n_24069), .B (n_34694), .Y (n_24076));
NAND2X1 g111881(.A (n_24067), .B (n_34694), .Y (n_24075));
NAND2X1 g111883(.A (n_24073), .B (n_30563), .Y (n_24074));
NAND2X1 g111884(.A (n_24071), .B (n_34694), .Y (n_24072));
NAND2X1 g111895(.A (n_27743), .B (n_24069), .Y (n_24070));
NAND2X1 g111896(.A (n_27743), .B (n_24067), .Y (n_24068));
NAND2X1 g111934(.A (n_24045), .B (n_35744), .Y (n_24747));
NAND4X1 g111949(.A (n_19190), .B (n_22416), .C (n_22431), .D(n_22727), .Y (n_24065));
NAND2X1 g111955(.A (n_24069), .B (n_34802), .Y (n_32099));
NAND2X1 g111956(.A (n_24062), .B (n_10808), .Y (n_24063));
NAND2X1 g111967(.A (n_24035), .B (n_24060), .Y (n_24733));
NAND2X1 g111973(.A (n_33288), .B (n_28158), .Y (n_24059));
NAND2X1 g111974(.A (n_33288), .B (n_26238), .Y (n_24057));
NAND2X1 g111978(.A (n_24067), .B (n_34802), .Y (n_24056));
NAND2X1 g111979(.A (n_24054), .B (n_10808), .Y (n_24055));
NAND2X1 g112013(.A (n_24073), .B (n_34802), .Y (n_24053));
NAND2X1 g112014(.A (n_24051), .B (n_10808), .Y (n_24052));
NAND4X1 g112031(.A (n_18622), .B (n_20650), .C (n_22748), .D(n_21141), .Y (n_24050));
NAND2X1 g112045(.A (n_24071), .B (n_34802), .Y (n_24049));
NAND2X1 g112046(.A (n_24047), .B (n_10808), .Y (n_24048));
NAND2X1 g112084(.A (n_24045), .B (n_18262), .Y (n_24046));
NAND2X1 g112085(.A (n_24032), .B (n_24965), .Y (n_24745));
NAND2X1 g112086(.A (n_24038), .B (n_18262), .Y (n_24044));
NAND2X1 g112094(.A (n_23657), .B (n_19769), .Y (n_24043));
NAND2X1 g112114(.A (n_24042), .B (n_24041), .Y (n_24741));
AOI21X1 g112116(.A0 (n_9546), .A1 (n_23036), .B0 (n_15174), .Y(n_24040));
NAND2X1 g112121(.A (n_24034), .B (n_18262), .Y (n_24039));
NAND2X1 g112124(.A (n_24038), .B (n_35816), .Y (n_24779));
NAND2X1 g112140(.A (n_24024), .B (n_33738), .Y (n_24037));
NAND2X1 g112142(.A (n_14410), .B (n_24035), .Y (n_24036));
NAND2X1 g112143(.A (n_24034), .B (n_35736), .Y (n_24748));
NAND2X1 g112145(.A (n_24032), .B (n_35790), .Y (n_24033));
NOR2X1 g112160(.A (n_23371), .B (n_10621), .Y (n_24031));
AOI21X1 g112181(.A0 (n_14819), .A1 (n_24028), .B0 (n_23378), .Y(n_24030));
AOI21X1 g112182(.A0 (n_14818), .A1 (n_24028), .B0 (n_23377), .Y(n_24029));
NAND2X1 g112183(.A (n_33288), .B (n_8954), .Y (n_24027));
NAND2X1 g112189(.A (n_24024), .B (n_28158), .Y (n_24025));
NAND2X1 g112190(.A (n_24024), .B (n_28374), .Y (n_24023));
NAND2X1 g112198(.A (n_23636), .B (n_33738), .Y (n_24022));
NAND2X1 g112205(.A (n_24017), .B (n_26238), .Y (n_24021));
NAND3X1 g112208(.A (n_22054), .B (n_23063), .C (n_22051), .Y(n_24020));
NAND2X1 g112210(.A (n_24032), .B (n_25599), .Y (n_24019));
NAND2X1 g112212(.A (n_24032), .B (n_35519), .Y (n_24735));
NAND2X1 g112217(.A (n_24034), .B (n_25877), .Y (n_24750));
NAND2X1 g112218(.A (n_24045), .B (n_25877), .Y (n_24762));
NAND2X1 g112219(.A (n_24038), .B (n_26584), .Y (n_24759));
NAND2X1 g112231(.A (n_24017), .B (n_29405), .Y (n_24018));
NAND2X1 g112232(.A (n_24017), .B (n_33738), .Y (n_24016));
NOR2X1 g112259(.A (n_9057), .B (n_23373), .Y (n_24015));
AOI21X1 g112267(.A0 (n_27100), .A1 (n_23992), .B0 (n_23139), .Y(n_24014));
OAI21X1 g112281(.A0 (n_24008), .A1 (n_24013), .B0 (n_24012), .Y(n_24767));
NAND2X1 g112284(.A (n_23413), .B (n_24011), .Y (n_24791));
OAI21X1 g112316(.A0 (n_23026), .A1 (n_24312), .B0 (n_24009), .Y(n_24788));
OAI21X1 g112319(.A0 (n_24008), .A1 (n_24889), .B0 (n_24007), .Y(n_24783));
NAND2X1 g112335(.A (n_23422), .B (n_23242), .Y (n_24777));
NAND2X1 g112364(.A (n_23417), .B (n_24006), .Y (n_24793));
OAI21X1 g112366(.A0 (n_24008), .A1 (n_32791), .B0 (n_24005), .Y(n_24771));
OAI21X1 g112382(.A0 (n_23026), .A1 (n_13653), .B0 (n_24003), .Y(n_24756));
NAND2X1 g112398(.A (n_23389), .B (n_24002), .Y (n_24743));
NAND2X1 g108518(.A (n_23331), .B (n_13628), .Y (n_24001));
AOI21X1 g112399(.A0 (n_23665), .A1 (n_14563), .B0 (n_26920), .Y(n_24000));
NAND2X1 g108519(.A (n_23309), .B (n_35057), .Y (n_23999));
NAND2X1 g108520(.A (n_23305), .B (n_13487), .Y (n_23998));
NAND2X1 g108524(.A (n_23264), .B (n_13181), .Y (n_23997));
NAND2X1 g112408(.A (n_23406), .B (n_23996), .Y (n_24737));
OAI21X1 g112409(.A0 (n_14210), .A1 (n_33713), .B0 (n_23408), .Y(n_23995));
AOI21X1 g112410(.A0 (n_23992), .A1 (n_27522), .B0 (n_18839), .Y(n_23993));
NAND2X1 g112421(.A (n_23399), .B (n_28364), .Y (n_23991));
AOI21X1 g112425(.A0 (n_8922), .A1 (n_23670), .B0 (n_18214), .Y(n_23990));
NAND4X1 g112433(.A (n_18625), .B (n_21599), .C (n_22667), .D(n_15139), .Y (n_23989));
NAND4X1 g112434(.A (n_32093), .B (n_32094), .C (n_22664), .D(n_20037), .Y (n_23988));
INVX1 g112438(.A (n_24447), .Y (n_23987));
MX2X1 g112467(.A (n_17536), .B (n_17537), .S0 (n_23655), .Y(n_24292));
MX2X1 g112470(.A (n_17557), .B (n_21502), .S0 (n_35170), .Y(n_24291));
INVX1 g112480(.A (n_23985), .Y (n_23986));
NAND2X1 g112486(.A (n_23558), .B (n_16411), .Y (n_23984));
NAND2X1 g112512(.A (n_23975), .B (n_28864), .Y (n_23983));
NAND2X1 g112515(.A (n_23973), .B (n_34952), .Y (n_23982));
NAND2X1 g112519(.A (n_23980), .B (n_28485), .Y (n_23981));
NAND2X1 g112522(.A (n_23977), .B (n_28485), .Y (n_23978));
NAND2X1 g112525(.A (n_23975), .B (n_28485), .Y (n_23976));
NAND2X1 g112528(.A (n_23973), .B (n_28492), .Y (n_23974));
NAND2X1 g112535(.A (n_23980), .B (n_25424), .Y (n_23972));
NAND2X1 g112539(.A (n_23977), .B (n_25424), .Y (n_23971));
NOR2X1 g112544(.A (n_22403), .B (n_23301), .Y (n_23970));
NAND2X1 g112545(.A (n_23975), .B (n_25424), .Y (n_23969));
NAND2X1 g112549(.A (n_23973), .B (n_29090), .Y (n_23968));
INVX1 g112555(.A (n_23966), .Y (n_23967));
NAND4X1 g112561(.A (n_15004), .B (n_22597), .C (n_22311), .D(n_22598), .Y (n_23965));
NOR2X1 g112562(.A (n_23303), .B (n_14606), .Y (n_23964));
INVX1 g112565(.A (n_23963), .Y (n_24259));
NAND2X1 g112575(.A (n_20087), .B (n_23599), .Y (n_23960));
NAND2X1 g112595(.A (n_23955), .B (n_24652), .Y (n_23958));
NAND2X1 g112612(.A (n_23950), .B (n_24446), .Y (n_23957));
NAND2X1 g112629(.A (n_23955), .B (n_18384), .Y (n_23956));
OR2X1 g112643(.A (n_24307), .B (n_25054), .Y (n_23954));
NAND2X1 g112656(.A (n_23955), .B (n_32664), .Y (n_23953));
AOI21X1 g112662(.A0 (n_23003), .A1 (n_24894), .B0 (n_26052), .Y(n_23952));
NAND2X1 g112670(.A (n_23950), .B (n_18378), .Y (n_23951));
NAND2X1 g112687(.A (n_23955), .B (n_13582), .Y (n_23949));
NAND2X1 g112697(.A (n_23620), .B (n_19707), .Y (n_23948));
NAND2X1 g112699(.A (n_23364), .B (n_23050), .Y (n_23947));
NAND2X2 g112707(.A (n_23338), .B (n_22588), .Y (n_24640));
NAND2X1 g112708(.A (n_35794), .B (n_23937), .Y (n_23946));
NAND2X1 g112721(.A (n_23361), .B (n_23047), .Y (n_23944));
NAND2X1 g112723(.A (n_23939), .B (n_14706), .Y (n_23943));
INVX1 g112729(.A (n_35388), .Y (n_24214));
INVX1 g112731(.A (n_23940), .Y (n_23941));
NAND2X1 g112744(.A (n_23379), .B (n_23939), .Y (n_24631));
NAND2X1 g112747(.A (n_18546), .B (n_23937), .Y (n_24210));
NOR2X1 g112750(.A (n_25748), .B (n_23564), .Y (n_23936));
NAND2X1 g112755(.A (n_23935), .B (n_23934), .Y (n_24610));
NAND2X1 g112756(.A (n_14387), .B (n_23931), .Y (n_23933));
NAND2X1 g112763(.A (n_23932), .B (n_23931), .Y (n_24600));
NAND3X1 g112770(.A (n_18008), .B (n_19925), .C (n_22974), .Y(n_23930));
NAND2X1 g112772(.A (n_23929), .B (n_22813), .Y (n_24614));
NAND2X1 g112773(.A (n_23575), .B (n_18458), .Y (n_32917));
INVX1 g112779(.A (n_23926), .Y (n_23927));
INVX1 g112783(.A (n_23925), .Y (n_24199));
NAND4X1 g112789(.A (n_14824), .B (n_22605), .C (n_22316), .D(n_22603), .Y (n_23924));
NAND2X1 g112793(.A (n_35540), .B (n_23937), .Y (n_24612));
NOR2X1 g112798(.A (n_22397), .B (n_23306), .Y (n_23923));
NOR2X1 g112803(.A (n_9938), .B (n_23347), .Y (n_23922));
NAND2X1 g112813(.A (n_23919), .B (n_23918), .Y (n_23921));
AND2X1 g112814(.A (n_23919), .B (n_23918), .Y (n_23920));
NAND2X1 g112818(.A (n_23337), .B (n_20412), .Y (n_33015));
NAND2X2 g112822(.A (n_23311), .B (n_19059), .Y (n_32096));
NAND2X1 g112824(.A (n_23334), .B (n_20904), .Y (n_32575));
NOR2X1 g112832(.A (n_9888), .B (n_23327), .Y (n_23914));
INVX1 g112836(.A (n_23912), .Y (n_23913));
AOI21X1 g112841(.A0 (n_23606), .A1 (n_32644), .B0 (n_15352), .Y(n_23911));
INVX1 g112847(.A (n_24395), .Y (n_23910));
NAND2X1 g112849(.A (n_23339), .B (n_23648), .Y (n_24647));
INVX1 g112856(.A (n_33710), .Y (n_23909));
NAND2X1 g112864(.A (n_23357), .B (n_23643), .Y (n_24687));
NAND2X1 g112877(.A (n_23345), .B (n_23641), .Y (n_24668));
OAI21X1 g112887(.A0 (n_23901), .A1 (n_17848), .B0 (n_27230), .Y(n_23907));
NAND2X1 g112894(.A (n_23330), .B (n_23638), .Y (n_24661));
INVX1 g112906(.A (n_23905), .Y (n_24604));
NAND2X1 g112910(.A (n_23333), .B (n_23904), .Y (n_24192));
NAND2X1 g112925(.A (n_23349), .B (n_25053), .Y (n_23903));
OAI21X1 g112930(.A0 (n_23901), .A1 (n_32698), .B0 (n_27219), .Y(n_23902));
NAND2X1 g112933(.A (n_23343), .B (n_25049), .Y (n_23900));
NAND2X1 g112935(.A (n_23340), .B (n_25048), .Y (n_23899));
NAND2X1 g112941(.A (n_23317), .B (n_23401), .Y (n_24623));
NAND2X1 g112944(.A (n_23328), .B (n_25682), .Y (n_23898));
NAND2X1 g112946(.A (n_23326), .B (n_23418), .Y (n_24617));
NAND3X1 g112948(.A (n_22988), .B (n_22423), .C (n_22982), .Y(n_23897));
AOI21X1 g112957(.A0 (n_22955), .A1 (n_22237), .B0 (n_21851), .Y(n_23896));
INVX1 g112983(.A (n_24383), .Y (n_24657));
NAND2X1 g112985(.A (n_23059), .B (n_23319), .Y (n_24670));
XOR2X1 g112991(.A (n_20832), .B (n_22973), .Y (n_24663));
INVX1 g112993(.A (n_23894), .Y (n_25050));
XOR2X1 g112997(.A (n_19211), .B (n_22997), .Y (n_24175));
INVX1 g113006(.A (n_23893), .Y (n_24628));
MX2X1 g113010(.A (n_19740), .B (n_19741), .S0 (n_23022), .Y(n_24174));
MX2X1 g113011(.A (n_19253), .B (n_23892), .S0 (n_22964), .Y(n_24621));
NAND2X1 g113024(.A (n_23067), .B (n_23324), .Y (n_24677));
NOR2X1 g113033(.A (n_22957), .B (n_23248), .Y (n_23891));
INVX1 g113043(.A (n_23889), .Y (n_23890));
NAND2X1 g113069(.A (n_21824), .B (n_23490), .Y (n_23888));
NAND3X1 g113073(.A (n_22252), .B (n_22895), .C (n_14599), .Y(n_23887));
AOI21X1 g113075(.A0 (n_22938), .A1 (n_22247), .B0 (n_8070), .Y(n_23886));
AOI21X1 g113076(.A0 (n_22937), .A1 (n_22245), .B0 (n_31041), .Y(n_23885));
NAND2X1 g108851(.A (n_23811), .B (n_16173), .Y (n_23884));
NAND3X1 g113089(.A (n_22924), .B (n_22934), .C (n_22945), .Y(n_23883));
NAND3X1 g113098(.A (n_22328), .B (n_22932), .C (n_22357), .Y(n_23882));
NAND3X1 g113102(.A (n_22309), .B (n_22930), .C (n_22350), .Y(n_23881));
NAND2X1 g113144(.A (n_23239), .B (n_18384), .Y (n_23880));
NAND2X1 g113154(.A (n_23243), .B (n_24247), .Y (n_23879));
NAND2X1 g113179(.A (n_23872), .B (n_24361), .Y (n_23878));
NAND2X1 g113204(.A (n_23875), .B (n_23874), .Y (n_23876));
NAND2X1 g113205(.A (n_23872), .B (n_13274), .Y (n_23873));
NAND2X1 g113208(.A (n_21454), .B (n_23870), .Y (n_23871));
NAND2X1 g113218(.A (n_23493), .B (n_19252), .Y (n_23869));
NOR2X1 g113250(.A (n_23240), .B (n_10554), .Y (n_23868));
NAND2X1 g113275(.A (n_23263), .B (n_21741), .Y (n_23867));
INVX1 g113283(.A (n_23865), .Y (n_23866));
NAND2X1 g113308(.A (n_23023), .B (n_23266), .Y (n_23864));
NAND3X1 g113312(.A (n_22946), .B (n_22905), .C (n_15008), .Y(n_23863));
NAND2X1 g113313(.A (n_23257), .B (n_21745), .Y (n_23862));
NAND2X1 g113324(.A (n_23292), .B (n_22499), .Y (n_23861));
NOR2X1 g113330(.A (n_9110), .B (n_23241), .Y (n_23860));
AOI21X1 g113338(.A0 (n_27100), .A1 (n_22383), .B0 (n_23244), .Y(n_23859));
NAND2X1 g113346(.A (n_23545), .B (n_32220), .Y (n_24528));
INVX1 g113364(.A (n_23858), .Y (n_24125));
AOI21X1 g113368(.A0 (n_21768), .A1 (n_23233), .B0 (n_21430), .Y(n_32876));
INVX1 g113374(.A (n_24274), .Y (n_23856));
NAND2X1 g113379(.A (n_23274), .B (n_23535), .Y (n_24555));
INVX1 g113384(.A (n_24271), .Y (n_23855));
NAND2X1 g113386(.A (n_23272), .B (n_23534), .Y (n_24546));
INVX1 g113391(.A (n_24233), .Y (n_23854));
NAND2X1 g113395(.A (n_23269), .B (n_23533), .Y (n_24537));
INVX1 g113401(.A (n_24225), .Y (n_23853));
NOR2X1 g113419(.A (n_22903), .B (n_23238), .Y (n_23852));
NAND2X1 g113428(.A (n_22710), .B (n_23279), .Y (n_23851));
NAND2X1 g113431(.A (n_22701), .B (n_23278), .Y (n_23850));
NAND2X1 g113433(.A (n_22690), .B (n_23277), .Y (n_23849));
NAND2X1 g113434(.A (n_22675), .B (n_23275), .Y (n_23848));
NAND2X1 g113456(.A (n_22971), .B (n_23259), .Y (n_24548));
MX2X1 g113457(.A (n_18447), .B (n_20322), .S0 (n_22901), .Y(n_24539));
INVX1 g113459(.A (n_23847), .Y (n_24891));
INVX1 g113461(.A (n_24239), .Y (n_23846));
INVX1 g113476(.A (n_23844), .Y (n_24114));
NAND2X1 g113479(.A (n_23258), .B (n_22967), .Y (n_24542));
INVX1 g113480(.A (n_24237), .Y (n_23843));
NAND2X1 g113614(.A (n_23224), .B (n_17921), .Y (n_32279));
AND2X1 g113653(.A (n_23235), .B (n_23839), .Y (n_23840));
NAND2X1 g113654(.A (n_23830), .B (n_22917), .Y (n_23838));
NOR2X1 g113667(.A (n_22513), .B (n_23227), .Y (n_23837));
NAND2X1 g113726(.A (n_23471), .B (n_17870), .Y (n_23836));
NOR2X1 g113737(.A (n_23834), .B (n_25881), .Y (n_23835));
NAND4X1 g113744(.A (n_23228), .B (n_21748), .C (n_21747), .D(n_18493), .Y (n_23832));
AOI21X1 g113753(.A0 (n_23478), .A1 (n_22918), .B0 (n_23830), .Y(n_23831));
INVX1 g113773(.A (n_24156), .Y (n_23829));
INVX1 g113805(.A (n_24159), .Y (n_23828));
AOI21X1 g114047(.A0 (n_23205), .A1 (n_13968), .B0 (n_31245), .Y(n_23827));
AOI21X1 g114048(.A0 (n_23204), .A1 (n_14204), .B0 (n_33125), .Y(n_23826));
OAI21X1 g114062(.A0 (n_23203), .A1 (n_14998), .B0 (n_24695), .Y(n_23825));
OAI21X1 g114063(.A0 (n_23202), .A1 (n_15145), .B0 (n_24695), .Y(n_23824));
AOI21X1 g114070(.A0 (n_23200), .A1 (n_14639), .B0 (n_8401), .Y(n_23823));
NOR2X1 g114123(.A (n_20606), .B (n_23466), .Y (n_23822));
OAI21X1 g114168(.A0 (n_9869), .A1 (n_24484), .B0 (n_23217), .Y(n_23821));
AOI21X1 g114195(.A0 (n_22854), .A1 (n_21270), .B0 (n_23464), .Y(n_23820));
NAND2X1 g109430(.A (n_23461), .B (n_25353), .Y (n_23819));
NAND2X1 g109432(.A (n_23459), .B (n_25350), .Y (n_23818));
NAND2X1 g109433(.A (n_23456), .B (n_25342), .Y (n_23817));
NAND2X1 g109443(.A (n_23454), .B (n_25336), .Y (n_23816));
NOR2X1 g109740(.A (n_23449), .B (n_14218), .Y (n_23813));
INVX1 g109870(.A (n_23811), .Y (n_23812));
NAND2X1 g109878(.A (n_23198), .B (n_24009), .Y (n_23810));
NAND2X1 g109901(.A (n_23196), .B (n_24006), .Y (n_23809));
NAND2X1 g109919(.A (n_23193), .B (n_24011), .Y (n_23808));
NAND2X1 g109936(.A (n_23189), .B (n_24003), .Y (n_23807));
OAI21X1 g110236(.A0 (n_23190), .A1 (n_23453), .B0 (n_23191), .Y(n_24130));
NAND2X1 g110456(.A (n_23183), .B (n_25111), .Y (n_23806));
NAND2X1 g110487(.A (n_23182), .B (n_24247), .Y (n_23805));
NAND2X1 g110518(.A (n_23180), .B (n_25111), .Y (n_23804));
NAND2X1 g110712(.A (n_23179), .B (n_8303), .Y (n_23803));
OAI21X1 g110805(.A0 (n_14003), .A1 (n_25368), .B0 (n_23188), .Y(n_23802));
NOR2X1 g110953(.A (n_23187), .B (n_15105), .Y (n_23801));
AOI21X1 g111198(.A0 (n_21896), .A1 (n_22823), .B0 (n_23031), .Y(n_23800));
NAND2X1 g111224(.A (n_23796), .B (n_18399), .Y (n_23799));
NAND2X1 g111230(.A (n_23793), .B (n_25198), .Y (n_23798));
NAND2X1 g111269(.A (n_23796), .B (n_20050), .Y (n_23797));
NAND2X1 g111306(.A (n_23796), .B (n_32723), .Y (n_23795));
NAND2X1 g111313(.A (n_23793), .B (n_35054), .Y (n_23794));
NAND2X1 g111352(.A (n_23796), .B (n_23791), .Y (n_23792));
NAND2X1 g111364(.A (n_23793), .B (n_23578), .Y (n_23790));
NAND2X1 g111435(.A (n_23793), .B (n_25207), .Y (n_23788));
NAND2X1 g111457(.A (n_23162), .B (n_24451), .Y (n_32061));
AOI22X1 g111509(.A0 (n_14882), .A1 (n_8313), .B0 (n_22819), .B1(n_25228), .Y (n_23786));
NAND2X1 g111707(.A (n_23174), .B (n_25706), .Y (n_23785));
NOR2X1 g111719(.A (n_23173), .B (n_13304), .Y (n_23784));
NAND2X1 g111723(.A (n_23171), .B (n_25689), .Y (n_23783));
NAND2X1 g111739(.A (n_23170), .B (n_25680), .Y (n_23782));
AOI21X1 g111775(.A0 (n_23443), .A1 (n_29411), .B0 (n_19833), .Y(n_23781));
NAND2X1 g111890(.A (n_23779), .B (n_23778), .Y (n_23780));
NAND2X1 g111909(.A (n_23776), .B (n_8954), .Y (n_23777));
NAND2X1 g111923(.A (n_23769), .B (n_18399), .Y (n_23775));
NAND2X1 g111942(.A (n_23132), .B (n_26458), .Y (n_23774));
NAND2X1 g111945(.A (n_23767), .B (n_22052), .Y (n_23773));
NAND2X1 g111961(.A (n_23137), .B (n_23771), .Y (n_23772));
NAND2X1 g111971(.A (n_23769), .B (n_24446), .Y (n_23770));
NAND2X1 g111975(.A (n_23767), .B (n_18918), .Y (n_23768));
NAND2X1 g111988(.A (n_23776), .B (n_28158), .Y (n_23765));
NAND2X1 g111995(.A (n_23769), .B (n_32652), .Y (n_23764));
NAND2X1 g112003(.A (n_23767), .B (n_32728), .Y (n_23763));
NAND2X1 g112011(.A (n_23129), .B (n_25220), .Y (n_23762));
NAND2X1 g112023(.A (n_23143), .B (n_25228), .Y (n_23761));
NAND2X1 g112037(.A (n_23769), .B (n_17797), .Y (n_23760));
NAND4X1 g112068(.A (n_21048), .B (n_22761), .C (n_20541), .D(n_20974), .Y (n_23759));
NAND2X1 g112144(.A (n_23131), .B (n_8641), .Y (n_23758));
NAND2X1 g112170(.A (n_23133), .B (n_8303), .Y (n_23757));
NAND2X1 g112173(.A (n_23776), .B (n_26238), .Y (n_23756));
NAND3X1 g112238(.A (n_22884), .B (n_18465), .C (n_23427), .Y(n_23755));
OAI21X1 g112244(.A0 (n_14852), .A1 (n_8614), .B0 (n_23152), .Y(n_23754));
NAND3X1 g112266(.A (n_9041), .B (n_22780), .C (n_19859), .Y(n_23752));
NAND2X1 g112272(.A (n_23158), .B (n_27389), .Y (n_23751));
NAND2X1 g112273(.A (n_23154), .B (n_27384), .Y (n_23750));
OAI21X1 g112276(.A0 (n_22754), .A1 (n_32707), .B0 (n_27380), .Y(n_23749));
NAND2X1 g112279(.A (n_23147), .B (n_27377), .Y (n_23748));
NAND2X1 g112290(.A (n_23151), .B (n_25713), .Y (n_23747));
NAND2X1 g112318(.A (n_23157), .B (n_25705), .Y (n_23746));
NAND2X1 g112379(.A (n_23146), .B (n_25684), .Y (n_23745));
NAND2X1 g112385(.A (n_23145), .B (n_25679), .Y (n_23744));
NAND2X1 g112394(.A (n_23155), .B (n_25702), .Y (n_23743));
AOI21X1 g112396(.A0 (n_23400), .A1 (n_14667), .B0 (n_29725), .Y(n_23742));
AOI21X1 g112411(.A0 (n_23390), .A1 (n_28158), .B0 (n_15021), .Y(n_23740));
XOR2X1 g112439(.A (n_21344), .B (n_22811), .Y (n_24447));
XOR2X1 g112475(.A (n_17712), .B (n_22784), .Y (n_24441));
NAND3X1 g112481(.A (n_22679), .B (n_22554), .C (n_22680), .Y(n_23985));
NAND2X1 g112487(.A (n_24563), .B (n_23723), .Y (n_23739));
NAND2X1 g112489(.A (n_24563), .B (n_23720), .Y (n_23738));
NAND2X1 g112490(.A (n_24563), .B (n_23713), .Y (n_23737));
NAND2X1 g112492(.A (n_24563), .B (n_23709), .Y (n_23736));
NAND3X1 g112495(.A (n_10600), .B (n_22715), .C (n_22401), .Y(n_23735));
NAND2X1 g112496(.A (n_24563), .B (n_23703), .Y (n_23734));
NAND2X1 g112498(.A (n_24563), .B (n_23700), .Y (n_23733));
NAND2X1 g112499(.A (n_24563), .B (n_23690), .Y (n_23732));
NAND2X1 g112501(.A (n_24563), .B (n_23687), .Y (n_23731));
NAND3X1 g112538(.A (n_22409), .B (n_22725), .C (n_22430), .Y(n_23730));
INVX1 g112556(.A (n_23729), .Y (n_23966));
NOR2X1 g112560(.A (n_27256), .B (n_23037), .Y (n_23728));
NAND2X1 g112566(.A (n_23058), .B (n_22546), .Y (n_23963));
NAND4X1 g112572(.A (n_22153), .B (n_22279), .C (n_22346), .D(n_21864), .Y (n_32359));
NOR2X1 g112577(.A (n_23044), .B (n_33807), .Y (n_23727));
NAND2X1 g112581(.A (n_23715), .B (n_23725), .Y (n_23726));
NAND2X1 g112586(.A (n_23723), .B (n_25756), .Y (n_23724));
NAND2X1 g112587(.A (n_23723), .B (n_34753), .Y (n_23722));
NAND2X1 g112591(.A (n_23720), .B (n_24526), .Y (n_23721));
NAND2X1 g112592(.A (n_23720), .B (n_28798), .Y (n_23719));
NAND2X1 g112593(.A (n_23680), .B (n_23718), .Y (n_24331));
NAND2X1 g112598(.A (n_23705), .B (n_18384), .Y (n_23717));
NAND2X1 g112614(.A (n_23715), .B (n_24446), .Y (n_23716));
NAND2X1 g112619(.A (n_23713), .B (n_25756), .Y (n_23714));
NAND2X1 g112620(.A (n_23713), .B (n_34753), .Y (n_23711));
NAND2X1 g112624(.A (n_23709), .B (n_26106), .Y (n_23710));
NAND2X1 g112625(.A (n_23709), .B (n_26213), .Y (n_23708));
NAND2X1 g112626(.A (n_23705), .B (n_24652), .Y (n_23706));
NAND2X1 g112647(.A (n_23703), .B (n_25756), .Y (n_23704));
NAND2X1 g112648(.A (n_23703), .B (n_34753), .Y (n_23702));
AND2X1 g112651(.A (n_23700), .B (n_26213), .Y (n_23701));
NAND2X1 g112653(.A (n_23700), .B (n_34753), .Y (n_23699));
NAND2X1 g112658(.A (n_23705), .B (n_13582), .Y (n_23698));
NAND2X1 g112675(.A (n_23715), .B (n_23696), .Y (n_23697));
NAND2X1 g112676(.A (n_23694), .B (n_23693), .Y (n_23695));
NAND3X1 g112678(.A (n_18408), .B (n_22714), .C (n_22395), .Y(n_23692));
NAND2X1 g112679(.A (n_23690), .B (n_25756), .Y (n_23691));
NAND2X1 g112680(.A (n_23690), .B (n_28636), .Y (n_23689));
AND2X1 g112683(.A (n_23687), .B (n_26112), .Y (n_23688));
NAND2X1 g112684(.A (n_23687), .B (n_24526), .Y (n_23686));
NAND2X1 g112693(.A (n_23667), .B (n_27109), .Y (n_23685));
NAND2X1 g112704(.A (n_23694), .B (n_21775), .Y (n_23684));
NAND3X1 g112710(.A (n_20436), .B (n_22687), .C (n_21015), .Y(n_23683));
NAND3X1 g112713(.A (n_23363), .B (n_23659), .C (n_20920), .Y(n_23682));
NAND2X1 g112716(.A (n_14347), .B (n_23680), .Y (n_23681));
NAND2X1 g112717(.A (n_23083), .B (n_19298), .Y (n_23679));
NAND2X1 g112719(.A (n_23112), .B (n_22145), .Y (n_23678));
NAND3X1 g112725(.A (n_22240), .B (n_22683), .C (n_22630), .Y(n_23677));
NAND2X1 g112726(.A (n_35170), .B (n_21427), .Y (n_23676));
NAND3X1 g112727(.A (n_23052), .B (n_21779), .C (n_22576), .Y(n_23674));
NAND3X1 g112732(.A (n_22986), .B (n_21918), .C (n_22681), .Y(n_23940));
NAND2X1 g112740(.A (n_29341), .B (n_23670), .Y (n_23672));
NAND2X1 g112741(.A (n_8990), .B (n_23670), .Y (n_23669));
NAND2X1 g112753(.A (n_24925), .B (n_23667), .Y (n_23668));
NAND2X1 g112754(.A (n_23666), .B (n_23665), .Y (n_24341));
NAND2X1 g112764(.A (n_23992), .B (n_26132), .Y (n_23664));
NAND2X1 g112769(.A (n_23299), .B (n_22036), .Y (n_23663));
NAND2X1 g112780(.A (n_22353), .B (n_23117), .Y (n_23926));
NAND2X1 g112784(.A (n_23116), .B (n_22356), .Y (n_23925));
NAND3X1 g112804(.A (n_9580), .B (n_22717), .C (n_22411), .Y(n_23662));
AOI22X1 g112810(.A0 (n_22653), .A1 (n_25122), .B0 (n_14758), .B1(n_8313), .Y (n_23661));
NAND2X1 g112817(.A (n_23051), .B (n_23659), .Y (n_23660));
INVX1 g112819(.A (n_23657), .Y (n_23658));
NAND2X2 g112821(.A (n_23655), .B (n_21002), .Y (n_23656));
NAND2X1 g112835(.A (n_23110), .B (n_13667), .Y (n_23652));
NAND2X2 g112837(.A (n_23109), .B (n_21596), .Y (n_23912));
NAND2X1 g112839(.A (n_23101), .B (n_13650), .Y (n_23651));
NAND2X1 g112840(.A (n_23093), .B (n_27220), .Y (n_23650));
NAND2X1 g112844(.A (n_23088), .B (n_26376), .Y (n_23649));
NAND2X1 g112848(.A (n_23085), .B (n_23648), .Y (n_24395));
NAND2X1 g112850(.A (n_23084), .B (n_23647), .Y (n_24365));
NAND2X1 g112858(.A (n_23049), .B (n_21416), .Y (n_33058));
OAI21X1 g112859(.A0 (n_26382), .A1 (n_22647), .B0 (n_22756), .Y(n_23645));
NAND2X1 g112862(.A (n_23074), .B (n_19933), .Y (n_23644));
NAND2X1 g112865(.A (n_23108), .B (n_23643), .Y (n_24404));
NAND2X1 g112868(.A (n_23104), .B (n_23642), .Y (n_24390));
NAND2X1 g112876(.A (n_23097), .B (n_23641), .Y (n_24401));
NAND2X1 g112878(.A (n_23095), .B (n_23640), .Y (n_24378));
NAND3X1 g112890(.A (n_22219), .B (n_23626), .C (n_21349), .Y(n_23639));
NAND2X1 g112895(.A (n_23077), .B (n_23638), .Y (n_24399));
NAND2X1 g112897(.A (n_23076), .B (n_23637), .Y (n_24352));
INVX1 g112903(.A (n_23636), .Y (n_24336));
NAND2X1 g112907(.A (n_23079), .B (n_23635), .Y (n_23905));
NAND2X1 g112919(.A (n_22801), .B (n_23103), .Y (n_23634));
NAND2X1 g112920(.A (n_22797), .B (n_23099), .Y (n_23633));
AOI21X1 g112952(.A0 (n_34770), .A1 (n_23286), .B0 (n_21644), .Y(n_23632));
AOI21X1 g112955(.A0 (n_34770), .A1 (n_23280), .B0 (n_21184), .Y(n_23630));
OAI21X1 g112969(.A0 (n_22371), .A1 (n_8664), .B0 (n_23125), .Y(n_23629));
NAND2X1 g112970(.A (n_22809), .B (n_23124), .Y (n_23628));
XOR2X1 g112973(.A (n_19624), .B (n_22720), .Y (n_24369));
OAI21X1 g112975(.A0 (n_23055), .A1 (n_27662), .B0 (n_23081), .Y(n_23627));
MX2X1 g112984(.A (n_18051), .B (n_18050), .S0 (n_22729), .Y(n_24383));
XOR2X1 g112994(.A (n_20831), .B (n_22662), .Y (n_23894));
MX2X1 g113007(.A (n_18056), .B (n_18055), .S0 (n_22685), .Y(n_23893));
OAI21X1 g113021(.A0 (n_32968), .A1 (n_23089), .B0 (n_23090), .Y(n_24345));
XOR2X1 g113022(.A (n_18047), .B (n_23626), .Y (n_24374));
XOR2X1 g113023(.A (n_23625), .B (n_22660), .Y (n_24372));
OAI21X1 g113034(.A0 (n_20543), .A1 (n_22269), .B0 (n_22992), .Y(n_23624));
OAI21X1 g113035(.A0 (n_22610), .A1 (n_16892), .B0 (n_22544), .Y(n_23623));
NAND4X1 g113038(.A (n_22904), .B (n_15148), .C (n_10074), .D(n_21827), .Y (n_23622));
INVX1 g113039(.A (n_23620), .Y (n_23621));
NAND3X1 g113042(.A (n_22961), .B (n_22313), .C (n_18202), .Y(n_23619));
NAND2X2 g113044(.A (n_32620), .B (n_32621), .Y (n_23889));
NAND2X1 g113045(.A (n_33546), .B (n_23603), .Y (n_23618));
AOI21X1 g113047(.A0 (n_22625), .A1 (n_22565), .B0 (n_31233), .Y(n_23617));
NAND2X1 g113051(.A (n_33546), .B (n_23591), .Y (n_23616));
NAND2X1 g113059(.A (n_33546), .B (n_23581), .Y (n_23615));
NAND2X1 g113064(.A (n_23552), .B (n_22165), .Y (n_23614));
NAND2X1 g113070(.A (n_33546), .B (n_23573), .Y (n_23613));
NAND2X1 g113074(.A (n_23249), .B (n_21426), .Y (n_23612));
NAND2X1 g113077(.A (n_22969), .B (n_34683), .Y (n_23611));
NAND3X1 g113105(.A (n_35690), .B (n_35691), .C (n_21932), .Y(n_23610));
NAND2X1 g113107(.A (n_35744), .B (n_23569), .Y (n_23609));
NAND2X1 g113109(.A (n_23606), .B (n_23725), .Y (n_23607));
OR2X1 g113111(.A (n_23901), .B (n_17288), .Y (n_23605));
NAND2X1 g113113(.A (n_23603), .B (n_30668), .Y (n_23604));
NAND2X1 g113114(.A (n_23603), .B (n_30180), .Y (n_23602));
INVX1 g113115(.A (n_23599), .Y (n_23600));
NAND2X1 g113122(.A (n_23593), .B (n_17719), .Y (n_23598));
NAND2X1 g113140(.A (n_23586), .B (n_24105), .Y (n_23597));
NAND2X1 g113143(.A (n_23606), .B (n_18384), .Y (n_23596));
NAND2X1 g113145(.A (n_23593), .B (n_18384), .Y (n_23594));
AND2X1 g113156(.A (n_23591), .B (n_27993), .Y (n_23592));
NAND2X1 g113157(.A (n_23591), .B (n_30559), .Y (n_23590));
NAND2X1 g113167(.A (n_21530), .B (n_22965), .Y (n_23589));
NAND2X1 g113168(.A (n_23593), .B (n_32764), .Y (n_23588));
NAND2X1 g113181(.A (n_23586), .B (n_23149), .Y (n_23587));
NAND2X1 g113184(.A (n_23606), .B (n_20154), .Y (n_23585));
AOI21X1 g113194(.A0 (n_22613), .A1 (n_24012), .B0 (n_26052), .Y(n_23584));
AND2X1 g113195(.A (n_23581), .B (n_27993), .Y (n_23582));
NAND2X1 g113196(.A (n_23581), .B (n_28431), .Y (n_23580));
NAND2X1 g113206(.A (n_23586), .B (n_23578), .Y (n_23579));
NAND2X1 g113213(.A (n_22959), .B (n_19258), .Y (n_23577));
INVX1 g113225(.A (n_23575), .Y (n_23576));
NAND2X1 g113230(.A (n_13957), .B (n_23567), .Y (n_24207));
NAND2X1 g113231(.A (n_23573), .B (n_28890), .Y (n_23574));
NAND2X1 g113233(.A (n_23573), .B (n_30180), .Y (n_23572));
NAND2X1 g113238(.A (n_22951), .B (n_25942), .Y (n_23571));
NAND2X1 g113251(.A (n_13957), .B (n_23569), .Y (n_24204));
NAND2X1 g113258(.A (n_35790), .B (n_23567), .Y (n_23568));
NAND2X1 g113260(.A (n_23586), .B (n_25207), .Y (n_23566));
NAND2X1 g113262(.A (n_23262), .B (n_19550), .Y (n_23565));
NAND2X1 g113276(.A (n_23019), .B (n_19614), .Y (n_23563));
AOI21X1 g113278(.A0 (n_21012), .A1 (n_22941), .B0 (n_21801), .Y(n_23562));
NAND4X1 g113279(.A (n_19903), .B (n_18702), .C (n_22878), .D(n_19968), .Y (n_23561));
INVX1 g113284(.A (n_23560), .Y (n_23865));
INVX1 g113295(.A (n_23558), .Y (n_23559));
NAND2X1 g113297(.A (n_35528), .B (n_23567), .Y (n_24198));
NAND2X1 g113300(.A (n_35540), .B (n_23569), .Y (n_24216));
NAND2X1 g113303(.A (n_25596), .B (n_23567), .Y (n_23557));
NAND2X1 g113305(.A (n_25596), .B (n_23569), .Y (n_23556));
NAND2X1 g113321(.A (n_22993), .B (n_25058), .Y (n_23555));
NAND2X1 g113325(.A (n_22989), .B (n_22192), .Y (n_23554));
NAND3X1 g113337(.A (n_9048), .B (n_22608), .C (n_18209), .Y(n_23551));
INVX1 g113339(.A (n_34522), .Y (n_23550));
OAI21X1 g113341(.A0 (n_22567), .A1 (n_24312), .B0 (n_25056), .Y(n_23548));
OAI21X1 g113343(.A0 (n_22567), .A1 (n_19330), .B0 (n_25051), .Y(n_23546));
NAND2X1 g113347(.A (n_22998), .B (n_23545), .Y (n_24278));
NAND2X1 g113351(.A (n_22981), .B (n_25047), .Y (n_23544));
NAND2X1 g113358(.A (n_23012), .B (n_23542), .Y (n_23543));
OAI21X1 g113360(.A0 (n_22569), .A1 (n_32803), .B0 (n_24896), .Y(n_23541));
OAI21X1 g113362(.A0 (n_22569), .A1 (n_23178), .B0 (n_24888), .Y(n_23539));
NAND2X2 g113365(.A (n_23017), .B (n_22243), .Y (n_23858));
NAND3X1 g113366(.A (n_22520), .B (n_22305), .C (n_22874), .Y(n_23538));
NAND2X1 g113367(.A (n_22966), .B (n_21379), .Y (n_35272));
NAND2X1 g113370(.A (n_23000), .B (n_26216), .Y (n_23536));
NAND2X1 g113375(.A (n_23016), .B (n_22760), .Y (n_24274));
NAND2X1 g113378(.A (n_23013), .B (n_23535), .Y (n_24283));
NAND2X1 g113385(.A (n_23009), .B (n_23534), .Y (n_24271));
NAND2X1 g113392(.A (n_23006), .B (n_22844), .Y (n_24233));
NAND2X1 g113396(.A (n_23004), .B (n_23533), .Y (n_24280));
NAND2X1 g113402(.A (n_22995), .B (n_22759), .Y (n_24225));
NAND2X1 g113405(.A (n_22976), .B (n_22842), .Y (n_24262));
OAI21X1 g113413(.A0 (n_23527), .A1 (n_23178), .B0 (n_26209), .Y(n_23532));
NAND2X1 g113414(.A (n_23011), .B (n_26207), .Y (n_23531));
OAI21X1 g113416(.A0 (n_22571), .A1 (n_32803), .B0 (n_26202), .Y(n_23530));
OAI21X1 g113417(.A0 (n_23527), .A1 (n_32654), .B0 (n_26200), .Y(n_23528));
OAI21X1 g113418(.A0 (n_22571), .A1 (n_23178), .B0 (n_26193), .Y(n_23526));
AOI22X1 g113420(.A0 (n_22898), .A1 (n_22161), .B0 (n_22592), .B1(n_23523), .Y (n_23524));
AOI22X1 g113421(.A0 (n_22896), .A1 (n_21409), .B0 (n_22589), .B1(n_23521), .Y (n_23522));
AOI22X1 g113438(.A0 (n_23254), .A1 (n_22163), .B0 (n_21836), .B1(n_23393), .Y (n_23520));
MX2X1 g113460(.A (n_19064), .B (n_19063), .S0 (n_22594), .Y(n_23847));
OAI21X1 g113463(.A0 (n_23350), .A1 (n_22978), .B0 (n_22979), .Y(n_24239));
INVX1 g113466(.A (n_23937), .Y (n_23519));
INVX1 g113471(.A (n_24307), .Y (n_23518));
MX2X1 g113477(.A (n_20327), .B (n_18444), .S0 (n_22587), .Y(n_23844));
NAND2X1 g113482(.A (n_22671), .B (n_22977), .Y (n_24237));
XOR2X1 g113488(.A (n_19471), .B (n_22591), .Y (n_24579));
INVX1 g113489(.A (n_23950), .Y (n_23517));
XOR2X1 g113497(.A (n_19000), .B (n_22579), .Y (n_24242));
OAI21X1 g113515(.A0 (n_22862), .A1 (n_22514), .B0 (n_22899), .Y(n_23515));
NAND2X1 g113523(.A (n_21953), .B (n_22897), .Y (n_23514));
NAND2X1 g113588(.A (n_23510), .B (n_27999), .Y (n_23513));
NAND2X1 g113594(.A (n_22886), .B (n_24446), .Y (n_23512));
NAND2X1 g113605(.A (n_23510), .B (n_23007), .Y (n_23511));
NAND2X1 g113624(.A (n_23510), .B (n_32652), .Y (n_23509));
NAND2X1 g113629(.A (n_22886), .B (n_23001), .Y (n_23507));
NAND2X1 g113641(.A (n_23510), .B (n_25290), .Y (n_23506));
NAND2X1 g113651(.A (n_22944), .B (n_23462), .Y (n_23505));
NAND2X1 g113692(.A (n_23501), .B (n_33738), .Y (n_23504));
NAND2X1 g113707(.A (n_23223), .B (n_17920), .Y (n_32280));
NAND2X1 g113722(.A (n_23501), .B (n_28158), .Y (n_23502));
NAND2X1 g113723(.A (n_23501), .B (n_28374), .Y (n_23500));
NAND2X1 g113733(.A (n_23222), .B (n_33738), .Y (n_23499));
NAND2X1 g113736(.A (n_23496), .B (n_26238), .Y (n_23498));
NAND2X1 g113741(.A (n_23496), .B (n_29405), .Y (n_23497));
NAND2X1 g113742(.A (n_23496), .B (n_33738), .Y (n_23495));
NAND2X1 g113774(.A (n_22920), .B (n_22960), .Y (n_24156));
INVX1 g113780(.A (n_23493), .Y (n_23494));
NAND2X1 g113797(.A (n_22925), .B (n_22954), .Y (n_24164));
NAND2X1 g113806(.A (n_22922), .B (n_22953), .Y (n_24159));
NAND2X1 g113811(.A (n_22913), .B (n_22952), .Y (n_24162));
INVX1 g113832(.A (n_23490), .Y (n_23491));
NAND2X1 g113834(.A (n_22909), .B (n_26548), .Y (n_23489));
OAI21X1 g113837(.A0 (n_22536), .A1 (n_23487), .B0 (n_22928), .Y(n_23488));
NAND2X1 g113840(.A (n_21120), .B (n_22935), .Y (n_23486));
NAND2X1 g113841(.A (n_22927), .B (n_22326), .Y (n_23485));
NAND2X1 g113842(.A (n_22307), .B (n_22926), .Y (n_23484));
AOI22X1 g113843(.A0 (n_23229), .A1 (n_21384), .B0 (n_22871), .B1(n_34725), .Y (n_23483));
OAI21X1 g113850(.A0 (n_23208), .A1 (n_10790), .B0 (n_22358), .Y(n_23481));
INVX1 g113870(.A (n_23872), .Y (n_23480));
OAI21X1 g113882(.A0 (n_23478), .A1 (n_23477), .B0 (n_22912), .Y(n_24149));
OAI21X1 g113884(.A0 (n_23252), .A1 (n_23476), .B0 (n_22911), .Y(n_24144));
XOR2X1 g113885(.A (n_19207), .B (n_22863), .Y (n_24146));
AND2X1 g113891(.A (n_21759), .B (n_23474), .Y (n_23475));
NAND2X1 g113969(.A (n_22861), .B (n_28915), .Y (n_23473));
INVX1 g114107(.A (n_23471), .Y (n_23472));
NOR2X1 g114125(.A (n_22196), .B (n_23216), .Y (n_23470));
NAND2X1 g114213(.A (n_23214), .B (n_21346), .Y (n_23468));
NAND3X1 g114214(.A (n_23207), .B (n_22864), .C (n_21345), .Y(n_23467));
OR4X1 g114364(.A (n_21394), .B (n_20213), .C (n_22146), .D (n_20330),.Y (n_23466));
INVX1 g114435(.A (n_23213), .Y (n_23465));
NOR2X1 g114444(.A (n_22855), .B (n_23230), .Y (n_23464));
NAND4X1 g114523(.A (n_21858), .B (n_21857), .C (n_21856), .D(n_23462), .Y (n_23463));
NAND2X1 g109634(.A (n_23458), .B (n_25554), .Y (n_23461));
NAND2X1 g109676(.A (n_22845), .B (n_9431), .Y (n_23460));
INVX1 g114852(.A (n_23199), .Y (n_23814));
NAND2X1 g109695(.A (n_23458), .B (n_23457), .Y (n_23459));
NAND2X1 g109719(.A (n_23458), .B (n_23578), .Y (n_23456));
NAND2X1 g109771(.A (n_22843), .B (n_9431), .Y (n_23455));
NAND2X1 g109798(.A (n_23458), .B (n_27422), .Y (n_23454));
NAND3X1 g109871(.A (n_21300), .B (n_23453), .C (n_21654), .Y(n_23811));
AOI21X1 g110814(.A0 (n_22455), .A1 (n_25942), .B0 (n_14659), .Y(n_23452));
AOI21X1 g110832(.A0 (n_22454), .A1 (n_25220), .B0 (n_14435), .Y(n_23451));
AOI21X1 g111033(.A0 (n_22457), .A1 (n_25220), .B0 (n_14244), .Y(n_23450));
INVX1 g111088(.A (n_23449), .Y (n_24103));
NAND2X1 g111240(.A (n_22840), .B (n_23771), .Y (n_23448));
NAND2X1 g111281(.A (n_22838), .B (n_25111), .Y (n_23447));
NAND2X1 g111311(.A (n_22837), .B (n_23771), .Y (n_23446));
OAI21X1 g111476(.A0 (n_22291), .A1 (n_9626), .B0 (n_22078), .Y(n_23445));
NAND2X1 g111922(.A (n_23443), .B (n_28158), .Y (n_23444));
NAND2X1 g111983(.A (n_22818), .B (n_8303), .Y (n_23442));
NAND2X1 g112021(.A (n_22815), .B (n_25228), .Y (n_23441));
NAND2X1 g112042(.A (n_23443), .B (n_26238), .Y (n_23440));
NAND2X1 g112070(.A (n_22814), .B (n_25111), .Y (n_23439));
NAND2X1 g112184(.A (n_23443), .B (n_8954), .Y (n_23438));
NAND2X1 g112240(.A (n_22835), .B (n_24840), .Y (n_23437));
NAND2X1 g112249(.A (n_22833), .B (n_24839), .Y (n_23436));
NAND2X1 g112255(.A (n_22826), .B (n_24843), .Y (n_23435));
NAND2X1 g112265(.A (n_22825), .B (n_24837), .Y (n_23434));
AOI21X1 g112415(.A0 (n_14395), .A1 (n_22821), .B0 (n_22829), .Y(n_23433));
NOR2X1 g112479(.A (n_22432), .B (n_22790), .Y (n_23432));
NAND2X1 g112484(.A (n_33546), .B (n_23424), .Y (n_23431));
NAND2X1 g112494(.A (n_33546), .B (n_23420), .Y (n_23430));
NAND2X1 g112503(.A (n_33546), .B (n_23415), .Y (n_23429));
NAND2X1 g112506(.A (n_22853), .B (n_23427), .Y (n_23428));
NAND2X1 g112507(.A (n_33546), .B (n_23404), .Y (n_23426));
NAND2X2 g112557(.A (n_32235), .B (n_32236), .Y (n_23729));
NAND2X1 g112579(.A (n_23424), .B (n_24786), .Y (n_23425));
NAND2X1 g112627(.A (n_22757), .B (n_24451), .Y (n_23423));
NAND2X1 g112628(.A (n_23027), .B (n_24249), .Y (n_23422));
AND2X1 g112636(.A (n_23420), .B (n_27993), .Y (n_23421));
NAND2X1 g112638(.A (n_23420), .B (n_28431), .Y (n_23419));
NAND2X1 g112640(.A (n_23418), .B (n_23398), .Y (n_24017));
NAND2X1 g112644(.A (n_23412), .B (n_25554), .Y (n_23417));
AND2X1 g112689(.A (n_23415), .B (n_27993), .Y (n_23416));
NAND2X1 g112690(.A (n_23415), .B (n_24786), .Y (n_23414));
NAND2X1 g112696(.A (n_23412), .B (n_27770), .Y (n_23413));
NAND2X1 g112718(.A (n_23082), .B (n_19299), .Y (n_23411));
NAND2X1 g112720(.A (n_23111), .B (n_19737), .Y (n_23410));
NAND3X1 g112736(.A (n_21519), .B (n_23368), .C (n_21917), .Y(n_23409));
NAND2X1 g112737(.A (n_23407), .B (n_29405), .Y (n_23408));
NAND2X1 g112745(.A (n_14439), .B (n_23397), .Y (n_23406));
NAND2X1 g112748(.A (n_23404), .B (n_30180), .Y (n_23405));
NAND2X1 g112749(.A (n_23404), .B (n_28890), .Y (n_23403));
NAND2X1 g112752(.A (n_24752), .B (n_23395), .Y (n_23402));
NAND2X1 g112757(.A (n_23401), .B (n_23400), .Y (n_24024));
NAND2X1 g112758(.A (n_14676), .B (n_23398), .Y (n_23399));
NAND2X1 g112759(.A (n_35744), .B (n_23397), .Y (n_24035));
NAND2X1 g112781(.A (n_23395), .B (n_27902), .Y (n_23396));
NAND3X1 g112791(.A (n_22507), .B (n_22728), .C (n_23393), .Y(n_32877));
NAND2X1 g112794(.A (n_24752), .B (n_23390), .Y (n_23392));
NAND2X1 g112795(.A (n_13311), .B (n_23397), .Y (n_24041));
NAND2X1 g112796(.A (n_35576), .B (n_23397), .Y (n_23389));
OAI21X1 g112807(.A0 (n_8831), .A1 (n_35012), .B0 (n_22791), .Y(n_23387));
NAND2X1 g112820(.A (n_22783), .B (n_22301), .Y (n_23657));
NAND4X1 g112826(.A (n_22022), .B (n_22487), .C (n_18344), .D(n_19580), .Y (n_23386));
AOI21X1 g112828(.A0 (n_24925), .A1 (n_23080), .B0 (n_22763), .Y(n_23385));
AOI21X1 g112829(.A0 (n_15173), .A1 (n_23060), .B0 (n_8927), .Y(n_23384));
AOI21X1 g112833(.A0 (n_27100), .A1 (n_23069), .B0 (n_22437), .Y(n_23383));
NAND2X1 g112845(.A (n_22787), .B (n_14049), .Y (n_24047));
NAND2X1 g112846(.A (n_22785), .B (n_14049), .Y (n_24071));
NAND2X1 g112871(.A (n_23382), .B (n_32062), .Y (n_24069));
NAND2X1 g112872(.A (n_22798), .B (n_23382), .Y (n_24062));
NAND2X1 g112874(.A (n_22796), .B (n_23381), .Y (n_24067));
NAND2X1 g112875(.A (n_22794), .B (n_23381), .Y (n_24054));
OAI21X1 g112885(.A0 (n_22363), .A1 (n_32673), .B0 (n_23380), .Y(n_24051));
OAI21X1 g112886(.A0 (n_22364), .A1 (n_32720), .B0 (n_23380), .Y(n_24073));
NAND2X1 g112904(.A (n_22782), .B (n_23379), .Y (n_23636));
NAND2X1 g112924(.A (n_22804), .B (n_9127), .Y (n_23378));
NAND2X1 g112929(.A (n_22803), .B (n_9090), .Y (n_23377));
NAND2X1 g112937(.A (n_22777), .B (n_26548), .Y (n_23376));
OAI21X1 g112960(.A0 (n_19137), .A1 (n_25540), .B0 (n_22771), .Y(n_23373));
AOI22X1 g112964(.A0 (n_22370), .A1 (n_17912), .B0 (n_21607), .B1(n_21521), .Y (n_23372));
OAI21X1 g112968(.A0 (n_19148), .A1 (n_25540), .B0 (n_22765), .Y(n_23371));
INVX1 g112979(.A (n_23370), .Y (n_24038));
INVX1 g113002(.A (n_23369), .Y (n_24045));
MX2X1 g113004(.A (n_19821), .B (n_18694), .S0 (n_23368), .Y(n_24032));
INVX1 g113019(.A (n_23367), .Y (n_24034));
NAND2X1 g113040(.A (n_22689), .B (n_22601), .Y (n_23620));
AOI21X1 g113041(.A0 (n_18899), .A1 (n_24247), .B0 (n_22657), .Y(n_23366));
NOR2X1 g113053(.A (n_10090), .B (n_22644), .Y (n_23365));
INVX1 g113061(.A (n_23363), .Y (n_23364));
NAND2X1 g113063(.A (n_23626), .B (n_21778), .Y (n_23919));
NAND2X1 g113065(.A (n_22972), .B (n_23028), .Y (n_32903));
INVX1 g113067(.A (n_23360), .Y (n_23361));
NOR2X1 g113095(.A (n_21957), .B (n_22643), .Y (n_23359));
AOI21X1 g113097(.A0 (n_21782), .A1 (n_23295), .B0 (n_23291), .Y(n_23358));
NAND3X1 g113116(.A (n_22622), .B (n_22223), .C (n_22341), .Y(n_23599));
NAND2X1 g113117(.A (n_23344), .B (n_23356), .Y (n_23357));
NAND2X1 g113119(.A (n_22651), .B (n_25942), .Y (n_23355));
NAND3X1 g113128(.A (n_21477), .B (n_23350), .C (n_19300), .Y(n_23351));
NAND2X1 g113133(.A (n_23342), .B (n_25302), .Y (n_23349));
NAND2X1 g113137(.A (n_22654), .B (n_24247), .Y (n_23348));
AOI21X1 g113138(.A0 (n_22348), .A1 (n_21884), .B0 (n_30537), .Y(n_23347));
NAND2X1 g113158(.A (n_22648), .B (n_25082), .Y (n_23346));
NAND2X1 g113160(.A (n_23344), .B (n_25554), .Y (n_23345));
NAND2X1 g113173(.A (n_23342), .B (n_35054), .Y (n_23343));
OAI21X1 g113177(.A0 (n_22304), .A1 (n_21586), .B0 (n_30956), .Y(n_23341));
NAND2X1 g113192(.A (n_23342), .B (n_26637), .Y (n_23340));
NAND2X1 g113199(.A (n_23344), .B (n_22994), .Y (n_23339));
NAND2X1 g113209(.A (n_22996), .B (n_21774), .Y (n_23338));
OAI21X1 g113211(.A0 (n_23918), .A1 (n_20919), .B0 (n_22522), .Y(n_23337));
NAND2X1 g113212(.A (n_35816), .B (n_23332), .Y (n_23931));
NAND2X1 g113214(.A (n_22958), .B (n_19820), .Y (n_23335));
NAND2X1 g113223(.A (n_22736), .B (n_22225), .Y (n_23334));
NAND2X1 g113226(.A (n_22740), .B (n_22373), .Y (n_23575));
NAND2X1 g113232(.A (n_18546), .B (n_23332), .Y (n_23333));
NAND2X1 g108933(.A (n_23308), .B (n_25554), .Y (n_23331));
NAND2X1 g113235(.A (n_13957), .B (n_23325), .Y (n_23939));
NAND2X1 g113236(.A (n_23344), .B (n_23329), .Y (n_23330));
NAND2X1 g113252(.A (n_23342), .B (n_25207), .Y (n_23328));
AOI21X1 g113254(.A0 (n_22347), .A1 (n_21882), .B0 (n_30537), .Y(n_23327));
NAND2X1 g113259(.A (n_35790), .B (n_23325), .Y (n_23326));
NAND2X1 g113264(.A (n_22672), .B (n_17396), .Y (n_23324));
NOR2X1 g113265(.A (n_22641), .B (n_17002), .Y (n_23323));
INVX1 g113272(.A (n_23061), .Y (n_23564));
NOR2X1 g113274(.A (n_22674), .B (n_14209), .Y (n_23322));
NAND2X1 g113277(.A (n_23018), .B (n_19615), .Y (n_23321));
NAND2X1 g113285(.A (n_22735), .B (n_21594), .Y (n_23560));
AOI21X1 g113286(.A0 (n_22629), .A1 (n_32924), .B0 (n_21488), .Y(n_32173));
NAND2X1 g113288(.A (n_22734), .B (n_18448), .Y (n_23319));
NAND2X1 g113290(.A (n_22368), .B (n_28136), .Y (n_23318));
NOR3X1 g113296(.A (n_20798), .B (n_20311), .C (n_22292), .Y(n_23558));
NAND2X1 g113301(.A (n_35528), .B (n_23325), .Y (n_23929));
NAND2X1 g113304(.A (n_25877), .B (n_23332), .Y (n_23934));
NAND2X1 g113306(.A (n_25596), .B (n_23325), .Y (n_23317));
NAND3X1 g113311(.A (n_32203), .B (n_32204), .C (n_21030), .Y(n_33059));
NOR2X1 g113315(.A (n_9128), .B (n_22646), .Y (n_23315));
NOR2X1 g113316(.A (n_9091), .B (n_22645), .Y (n_23314));
AOI21X1 g113318(.A0 (n_14759), .A1 (n_20688), .B0 (n_22698), .Y(n_23313));
NAND3X1 g113326(.A (n_22697), .B (n_21770), .C (n_21354), .Y(n_23312));
NAND2X1 g113331(.A (n_22738), .B (n_22187), .Y (n_23311));
NAND3X1 g113332(.A (n_32904), .B (n_32905), .C (n_19900), .Y(n_23310));
NAND2X1 g113345(.A (n_23046), .B (n_32076), .Y (n_23973));
NAND2X1 g108987(.A (n_23308), .B (n_24361), .Y (n_23309));
NAND2X1 g113377(.A (n_22709), .B (n_23043), .Y (n_23980));
NAND2X1 g113383(.A (n_22705), .B (n_23041), .Y (n_23977));
NAND2X1 g113394(.A (n_22700), .B (n_23039), .Y (n_23975));
NAND2X1 g113399(.A (n_22722), .B (n_22428), .Y (n_23306));
NAND2X1 g109016(.A (n_23308), .B (n_23578), .Y (n_23305));
INVX1 g113423(.A (n_23667), .Y (n_23304));
NAND3X1 g113426(.A (n_21963), .B (n_22349), .C (n_21964), .Y(n_23303));
AOI21X1 g113432(.A0 (n_14985), .A1 (n_23176), .B0 (n_22694), .Y(n_23302));
NAND2X1 g113442(.A (n_22724), .B (n_22429), .Y (n_23301));
AOI21X1 g113444(.A0 (n_22987), .A1 (n_29411), .B0 (n_19350), .Y(n_23300));
INVX1 g113445(.A (n_23299), .Y (n_24301));
NAND4X1 g113447(.A (n_20764), .B (n_18474), .C (n_22611), .D(n_21449), .Y (n_23298));
INVX1 g113450(.A (n_23715), .Y (n_23297));
OAI21X1 g113454(.A0 (n_32433), .A1 (n_22706), .B0 (n_22708), .Y(n_23955));
NAND2X1 g113467(.A (n_22388), .B (n_22682), .Y (n_23937));
XOR2X1 g113472(.A (n_23296), .B (n_23295), .Y (n_24307));
INVX1 g113473(.A (n_23705), .Y (n_23294));
XOR2X1 g113491(.A (n_17831), .B (n_22359), .Y (n_23950));
NAND4X1 g113504(.A (n_22856), .B (n_18228), .C (n_20601), .D(n_20618), .Y (n_23293));
NAND2X1 g113517(.A (n_23291), .B (n_22632), .Y (n_23292));
NAND2X1 g113537(.A (n_34770), .B (n_23284), .Y (n_23290));
NAND2X1 g113540(.A (n_34770), .B (n_23282), .Y (n_23288));
NAND2X1 g113544(.A (n_23286), .B (n_34709), .Y (n_23287));
NAND2X1 g113547(.A (n_23284), .B (n_34709), .Y (n_23285));
NAND2X1 g113550(.A (n_23282), .B (n_25988), .Y (n_23283));
NAND2X1 g113552(.A (n_23280), .B (n_34709), .Y (n_23281));
NAND2X1 g113555(.A (n_23286), .B (n_29199), .Y (n_23279));
NAND2X1 g113559(.A (n_23284), .B (n_29199), .Y (n_23278));
NAND2X1 g113560(.A (n_21859), .B (n_22943), .Y (n_24178));
NAND2X1 g113564(.A (n_23282), .B (n_28013), .Y (n_23277));
NAND2X1 g113567(.A (n_23280), .B (n_29199), .Y (n_23275));
NAND2X1 g113587(.A (n_23271), .B (n_22412), .Y (n_23274));
NAND2X1 g113595(.A (n_22616), .B (n_21867), .Y (n_23273));
NAND2X1 g113604(.A (n_23271), .B (n_23270), .Y (n_23272));
NAND2X1 g113621(.A (n_23271), .B (n_32798), .Y (n_23269));
NAND2X1 g113638(.A (n_23271), .B (n_26866), .Y (n_32220));
AOI21X1 g113655(.A0 (n_22516), .A1 (n_23255), .B0 (n_22556), .Y(n_23267));
AOI21X1 g113662(.A0 (n_14780), .A1 (n_15147), .B0 (n_22631), .Y(n_23266));
NAND2X1 g109151(.A (n_23308), .B (n_26676), .Y (n_23264));
INVX1 g113712(.A (n_23262), .Y (n_23263));
INVX1 g113716(.A (n_23552), .Y (n_23261));
NAND2X2 g113724(.A (n_22624), .B (n_21540), .Y (n_23870));
AOI21X1 g113725(.A0 (n_22515), .A1 (n_22623), .B0 (n_23219), .Y(n_23260));
NAND2X1 g113728(.A (n_22602), .B (n_17871), .Y (n_23259));
NAND2X1 g113734(.A (n_22581), .B (n_18500), .Y (n_23258));
NAND2X1 g113748(.A (n_22635), .B (n_20982), .Y (n_23257));
AOI21X1 g113754(.A0 (n_23255), .A1 (n_21786), .B0 (n_23254), .Y(n_23256));
AOI21X1 g113755(.A0 (n_23252), .A1 (n_22915), .B0 (n_22990), .Y(n_23253));
AOI21X1 g113758(.A0 (n_20460), .A1 (n_22535), .B0 (n_22249), .Y(n_23875));
NAND2X1 g113762(.A (n_22324), .B (n_22627), .Y (n_23251));
NOR2X1 g113767(.A (n_22607), .B (n_21945), .Y (n_23250));
INVX1 g113781(.A (n_23249), .Y (n_23493));
OAI21X1 g113783(.A0 (n_26382), .A1 (n_22241), .B0 (n_22572), .Y(n_23248));
AOI21X1 g113790(.A0 (n_21034), .A1 (n_22873), .B0 (n_21804), .Y(n_23247));
AOI21X1 g113795(.A0 (n_34770), .A1 (n_22931), .B0 (n_14788), .Y(n_23246));
AOI21X1 g113796(.A0 (n_34770), .A1 (n_22929), .B0 (n_14333), .Y(n_23245));
AOI21X1 g113815(.A0 (n_22910), .A1 (n_14565), .B0 (n_29725), .Y(n_23244));
NAND2X1 g113821(.A (n_22614), .B (n_23242), .Y (n_23243));
NAND2X1 g113833(.A (n_22585), .B (n_22555), .Y (n_23490));
OAI21X1 g113844(.A0 (n_17492), .A1 (n_25540), .B0 (n_22599), .Y(n_23241));
NAND2X1 g113846(.A (n_22595), .B (n_18207), .Y (n_23240));
INVX1 g113847(.A (n_23901), .Y (n_23239));
OAI21X1 g113856(.A0 (n_22902), .A1 (n_8661), .B0 (n_22323), .Y(n_23238));
XOR2X1 g113872(.A (n_20830), .B (n_22562), .Y (n_23872));
INVX1 g113889(.A (n_23593), .Y (n_23237));
OAI21X1 g113909(.A0 (n_22504), .A1 (n_22169), .B0 (n_21818), .Y(n_23830));
NAND4X1 g114033(.A (n_22157), .B (n_22177), .C (n_19720), .D(n_22231), .Y (n_23236));
NAND3X1 g114034(.A (n_22868), .B (n_21286), .C (n_21733), .Y(n_23235));
INVX1 g114082(.A (n_23233), .Y (n_23234));
NAND2X1 g114094(.A (n_22534), .B (n_28136), .Y (n_23232));
NOR3X1 g114103(.A (n_23230), .B (n_20913), .C (n_23211), .Y(n_23231));
AOI21X1 g114108(.A0 (n_22619), .A1 (n_20845), .B0 (n_23229), .Y(n_23471));
INVX1 g114116(.A (n_22900), .Y (n_23228));
NAND4X1 g114129(.A (n_22866), .B (n_23226), .C (n_33230), .D(n_23225), .Y (n_23227));
INVX1 g114152(.A (n_23223), .Y (n_23224));
INVX1 g114190(.A (n_23222), .Y (n_23834));
AOI22X1 g114196(.A0 (n_33008), .A1 (n_22985), .B0 (n_18420), .B1(n_20411), .Y (n_32174));
AOI22X1 g114210(.A0 (n_23219), .A1 (n_23218), .B0 (n_19028), .B1(n_20499), .Y (n_23220));
OAI21X1 g114296(.A0 (n_22490), .A1 (n_15406), .B0 (n_33123), .Y(n_23217));
OR4X1 g114369(.A (n_19779), .B (n_21391), .C (n_21737), .D (n_19653),.Y (n_23216));
NAND3X1 g114377(.A (n_19689), .B (n_21364), .C (n_22489), .Y(n_23215));
NOR2X1 g114393(.A (n_23206), .B (n_22188), .Y (n_23214));
AOI21X1 g114436(.A0 (n_21758), .A1 (n_23212), .B0 (n_23211), .Y(n_23213));
NAND4X1 g114466(.A (n_21507), .B (n_21636), .C (n_21506), .D(n_22745), .Y (n_23210));
NOR2X1 g114529(.A (n_22494), .B (n_22158), .Y (n_23474));
NOR2X1 g114672(.A (n_23206), .B (n_11716), .Y (n_23207));
NOR2X1 g114730(.A (n_22141), .B (n_22483), .Y (n_23205));
NOR2X1 g114731(.A (n_22488), .B (n_22484), .Y (n_23204));
NAND4X1 g114732(.A (n_22468), .B (n_14352), .C (n_23201), .D(n_21230), .Y (n_23203));
NAND4X1 g114733(.A (n_22467), .B (n_14574), .C (n_23201), .D(n_21231), .Y (n_23202));
NOR2X1 g114734(.A (n_22115), .B (n_22481), .Y (n_23200));
NAND3X1 g114853(.A (n_22485), .B (n_22171), .C (n_20510), .Y(n_23199));
NAND2X1 g110422(.A (n_23195), .B (n_25605), .Y (n_23198));
NAND2X1 g110494(.A (n_23195), .B (n_21919), .Y (n_23196));
NAND2X1 g110547(.A (n_23195), .B (n_23192), .Y (n_23193));
NAND2X1 g110551(.A (n_23190), .B (n_23453), .Y (n_23191));
NAND2X1 g110644(.A (n_23195), .B (n_18137), .Y (n_23189));
XOR2X1 g111089(.A (n_18275), .B (n_22079), .Y (n_23449));
NAND2X1 g111209(.A (n_22456), .B (n_25082), .Y (n_23188));
AOI21X1 g111324(.A0 (n_22074), .A1 (n_24895), .B0 (n_26052), .Y(n_23187));
AOI21X1 g111475(.A0 (n_22726), .A1 (n_29027), .B0 (n_21651), .Y(n_23186));
AOI21X1 g111514(.A0 (n_14872), .A1 (n_22821), .B0 (n_22462), .Y(n_23185));
AOI21X1 g111523(.A0 (n_14868), .A1 (n_22821), .B0 (n_22461), .Y(n_23184));
NAND2X1 g111562(.A (n_22463), .B (n_25590), .Y (n_23183));
OAI21X1 g111563(.A0 (n_22070), .A1 (n_32646), .B0 (n_23181), .Y(n_23182));
NAND2X1 g111564(.A (n_22460), .B (n_24892), .Y (n_23180));
OAI21X1 g111565(.A0 (n_22070), .A1 (n_23178), .B0 (n_24890), .Y(n_23179));
AOI21X1 g111755(.A0 (n_14864), .A1 (n_23176), .B0 (n_22458), .Y(n_23177));
NAND3X1 g111845(.A (n_18015), .B (n_19834), .C (n_22067), .Y(n_23175));
NAND2X1 g111947(.A (n_23172), .B (n_24105), .Y (n_23174));
AND2X1 g112001(.A (n_23172), .B (n_27770), .Y (n_23173));
NAND2X1 g112024(.A (n_23172), .B (n_23578), .Y (n_23171));
NAND2X1 g112149(.A (n_23172), .B (n_25605), .Y (n_23170));
AOI21X1 g112239(.A0 (n_22048), .A1 (n_25942), .B0 (n_14409), .Y(n_23169));
AOI21X1 g112248(.A0 (n_22047), .A1 (n_25942), .B0 (n_14849), .Y(n_23168));
AOI21X1 g112264(.A0 (n_22046), .A1 (n_9431), .B0 (n_14400), .Y(n_23167));
OAI21X1 g112294(.A0 (n_23164), .A1 (n_19037), .B0 (n_34800), .Y(n_23166));
OAI21X1 g112395(.A0 (n_23164), .A1 (n_32765), .B0 (n_25696), .Y(n_23165));
OAI21X1 g112401(.A0 (n_23164), .A1 (n_22042), .B0 (n_25675), .Y(n_23162));
AOI21X1 g112429(.A0 (n_22049), .A1 (n_25220), .B0 (n_14397), .Y(n_23161));
XOR2X1 g112444(.A (n_19098), .B (n_23427), .Y (n_23793));
MX2X1 g112476(.A (n_20741), .B (n_16420), .S0 (n_22050), .Y(n_23796));
AOI21X1 g112508(.A0 (n_27743), .A1 (n_22807), .B0 (n_10555), .Y(n_23160));
AOI21X1 g112509(.A0 (n_27743), .A1 (n_22805), .B0 (n_17833), .Y(n_23159));
NAND2X1 g112578(.A (n_23153), .B (n_23725), .Y (n_23158));
NAND2X1 g112589(.A (n_23150), .B (n_25554), .Y (n_23157));
NAND2X1 g112597(.A (n_22442), .B (n_8303), .Y (n_23156));
NAND2X1 g112609(.A (n_22434), .B (n_18384), .Y (n_23155));
NAND2X1 g112613(.A (n_23153), .B (n_24446), .Y (n_23154));
NAND2X1 g112631(.A (n_22440), .B (n_25111), .Y (n_23152));
NAND2X1 g112652(.A (n_23150), .B (n_23149), .Y (n_23151));
NAND2X1 g112654(.A (n_22438), .B (n_8303), .Y (n_23148));
NAND2X1 g112671(.A (n_23153), .B (n_22786), .Y (n_23147));
NAND2X1 g112692(.A (n_23150), .B (n_23578), .Y (n_23146));
NAND2X1 g112760(.A (n_23150), .B (n_27422), .Y (n_23145));
NAND3X1 g112797(.A (n_22523), .B (n_19633), .C (n_22810), .Y(n_23779));
NAND2X1 g112863(.A (n_22444), .B (n_25271), .Y (n_23143));
NAND2X1 g112884(.A (n_22447), .B (n_25355), .Y (n_23142));
NAND3X1 g112892(.A (n_21079), .B (n_35324), .C (n_35414), .Y(n_23141));
AOI21X1 g112900(.A0 (n_22778), .A1 (n_15020), .B0 (n_23138), .Y(n_23139));
NAND2X1 g112913(.A (n_22450), .B (n_23136), .Y (n_23137));
OAI21X1 g112915(.A0 (n_22010), .A1 (n_32765), .B0 (n_25264), .Y(n_23135));
NAND2X1 g112918(.A (n_22449), .B (n_25260), .Y (n_23133));
NAND2X1 g112923(.A (n_22451), .B (n_25055), .Y (n_23132));
NAND2X1 g112927(.A (n_22443), .B (n_24721), .Y (n_23131));
OAI21X1 g112931(.A0 (n_35532), .A1 (n_22362), .B0 (n_23130), .Y(n_23776));
NAND2X1 g112932(.A (n_22445), .B (n_25345), .Y (n_23129));
NAND4X1 g112956(.A (n_17511), .B (n_17958), .C (n_20008), .D(n_21598), .Y (n_23128));
MX2X1 g112980(.A (n_18674), .B (n_18675), .S0 (n_22766), .Y(n_23370));
MX2X1 g113003(.A (n_18085), .B (n_18086), .S0 (n_34290), .Y(n_23369));
MX2X1 g113020(.A (n_18120), .B (n_18121), .S0 (n_35324), .Y(n_23367));
XOR2X1 g113030(.A (n_17715), .B (n_22038), .Y (n_23769));
XOR2X1 g113031(.A (n_16423), .B (n_22011), .Y (n_23767));
NAND2X1 g113048(.A (n_26756), .B (n_23102), .Y (n_23125));
NAND2X1 g113050(.A (n_26756), .B (n_23098), .Y (n_23124));
OAI21X1 g113052(.A0 (n_21961), .A1 (n_21922), .B0 (n_7827), .Y(n_23123));
NAND2X1 g113054(.A (n_26756), .B (n_23091), .Y (n_23121));
NAND3X1 g113057(.A (n_17276), .B (n_21976), .C (n_21955), .Y(n_23120));
NAND2X1 g113058(.A (n_26756), .B (n_23086), .Y (n_23119));
AND2X1 g113062(.A (n_22659), .B (n_21460), .Y (n_23363));
AND2X1 g113068(.A (n_32969), .B (n_21006), .Y (n_23360));
NAND2X1 g113071(.A (n_21005), .B (n_22658), .Y (n_23117));
NAND2X1 g113072(.A (n_22661), .B (n_21448), .Y (n_23116));
NAND3X1 g113087(.A (n_21971), .B (n_21986), .C (n_22005), .Y(n_23115));
NAND3X1 g113090(.A (n_21968), .B (n_21984), .C (n_22004), .Y(n_23114));
NAND3X1 g113093(.A (n_21960), .B (n_21982), .C (n_22003), .Y(n_23113));
INVX1 g113099(.A (n_23111), .Y (n_23112));
NAND2X1 g113106(.A (n_23100), .B (n_27999), .Y (n_23110));
NAND2X1 g113108(.A (n_23066), .B (n_20961), .Y (n_23109));
NAND2X1 g113118(.A (n_23096), .B (n_24386), .Y (n_23108));
NAND2X1 g113126(.A (n_23094), .B (n_27747), .Y (n_23104));
NAND2X1 g113132(.A (n_23102), .B (n_34753), .Y (n_23103));
NAND2X1 g113142(.A (n_23100), .B (n_23270), .Y (n_23101));
NAND2X1 g113149(.A (n_23098), .B (n_34753), .Y (n_23099));
NAND2X1 g113159(.A (n_23096), .B (n_25554), .Y (n_23097));
NAND2X1 g113161(.A (n_23094), .B (n_22032), .Y (n_23095));
NAND2X1 g113166(.A (n_23100), .B (n_32786), .Y (n_23093));
NAND2X1 g113171(.A (n_23091), .B (n_10808), .Y (n_23092));
NAND2X1 g113180(.A (n_32968), .B (n_23089), .Y (n_23090));
NAND2X1 g113183(.A (n_23100), .B (n_34688), .Y (n_23088));
NAND2X2 g113185(.A (n_22696), .B (n_21492), .Y (n_23694));
NAND2X1 g113187(.A (n_23086), .B (n_10808), .Y (n_23087));
NAND2X1 g113198(.A (n_23096), .B (n_22994), .Y (n_23085));
NAND2X1 g113200(.A (n_23094), .B (n_25956), .Y (n_23084));
NAND2X2 g113215(.A (n_22743), .B (n_20600), .Y (n_23655));
NAND2X2 g113216(.A (n_22741), .B (n_21053), .Y (n_35170));
INVX1 g113219(.A (n_23082), .Y (n_23083));
NAND2X1 g113227(.A (n_8990), .B (n_23080), .Y (n_23081));
NAND2X1 g113228(.A (n_13504), .B (n_22673), .Y (n_23670));
NAND2X1 g113229(.A (n_24965), .B (n_23071), .Y (n_23079));
NAND2X1 g113237(.A (n_23096), .B (n_23329), .Y (n_23077));
NAND2X1 g113239(.A (n_23094), .B (n_25193), .Y (n_23076));
NAND2X1 g113242(.A (n_23073), .B (n_8990), .Y (n_23075));
NAND2X1 g113244(.A (n_23073), .B (n_27522), .Y (n_23074));
NAND2X2 g113247(.A (n_33781), .B (n_21001), .Y (n_23072));
NAND2X1 g113248(.A (n_35736), .B (n_23071), .Y (n_23680));
NAND2X1 g113255(.A (n_23069), .B (n_29505), .Y (n_23070));
NAND2X1 g113256(.A (n_23069), .B (n_26255), .Y (n_23068));
NAND2X1 g113263(.A (n_23066), .B (n_17395), .Y (n_23067));
NAND2X1 g113267(.A (n_22379), .B (n_27522), .Y (n_23065));
NAND2X1 g113268(.A (n_24925), .B (n_23062), .Y (n_23064));
NAND2X1 g113269(.A (n_27614), .B (n_23062), .Y (n_23063));
NAND2X2 g113273(.A (n_23060), .B (n_22758), .Y (n_23061));
NAND2X1 g113287(.A (n_23057), .B (n_20325), .Y (n_23059));
NAND2X1 g113289(.A (n_23057), .B (n_20847), .Y (n_23058));
NOR2X1 g113292(.A (n_23055), .B (n_25881), .Y (n_23056));
NAND2X1 g113302(.A (n_25877), .B (n_23071), .Y (n_23665));
NAND4X1 g113309(.A (n_23053), .B (n_33768), .C (n_33770), .D(n_21904), .Y (n_23054));
NOR2X1 g113310(.A (n_22367), .B (n_21312), .Y (n_23052));
OAI21X1 g113327(.A0 (n_23050), .A1 (n_20440), .B0 (n_22190), .Y(n_23051));
NAND2X1 g113333(.A (n_22425), .B (n_21809), .Y (n_23049));
NAND2X1 g113344(.A (n_35261), .B (n_23046), .Y (n_23690));
NAND2X1 g113348(.A (n_23045), .B (n_32212), .Y (n_23687));
INVX1 g113372(.A (n_23424), .Y (n_23044));
NAND2X1 g113376(.A (n_22415), .B (n_23043), .Y (n_23723));
NAND2X1 g113381(.A (n_22413), .B (n_23042), .Y (n_23720));
NAND2X1 g113382(.A (n_22408), .B (n_23041), .Y (n_23713));
NAND2X1 g113389(.A (n_22405), .B (n_23040), .Y (n_23709));
NAND2X1 g113393(.A (n_22400), .B (n_23039), .Y (n_23703));
NAND2X1 g113397(.A (n_22399), .B (n_23038), .Y (n_23700));
INVX1 g113403(.A (n_23407), .Y (n_23037));
INVX1 g113411(.A (n_23035), .Y (n_23036));
OAI21X1 g113424(.A0 (n_23034), .A1 (n_21933), .B0 (n_22779), .Y(n_23667));
NAND2X1 g113425(.A (n_22381), .B (n_22776), .Y (n_23992));
NAND2X1 g113427(.A (n_22386), .B (n_19936), .Y (n_23033));
NAND3X1 g113435(.A (n_21792), .B (n_23024), .C (n_20307), .Y(n_23032));
NAND2X1 g113437(.A (n_22419), .B (n_22329), .Y (n_23031));
NAND4X1 g113439(.A (n_23295), .B (n_21999), .C (n_23029), .D(n_23028), .Y (n_23030));
XOR2X1 g113446(.A (n_16126), .B (n_21995), .Y (n_23299));
XOR2X1 g113451(.A (n_20195), .B (n_21974), .Y (n_23715));
INVX1 g113452(.A (n_23027), .Y (n_24008));
INVX1 g113468(.A (n_23412), .Y (n_23026));
MX2X1 g113474(.A (n_17868), .B (n_20328), .S0 (n_23024), .Y(n_23705));
NOR2X1 g113499(.A (n_21629), .B (n_22533), .Y (n_23023));
NAND2X1 g113526(.A (n_21954), .B (n_22303), .Y (n_23022));
NAND2X1 g113535(.A (n_22586), .B (n_35119), .Y (n_32620));
OAI21X1 g113565(.A0 (n_22268), .A1 (n_21396), .B0 (n_22256), .Y(n_23020));
INVX1 g113568(.A (n_23018), .Y (n_23019));
NAND2X1 g113574(.A (n_22970), .B (n_20503), .Y (n_23017));
NAND2X1 g113577(.A (n_23005), .B (n_26676), .Y (n_23016));
NAND2X1 g113585(.A (n_22290), .B (n_24247), .Y (n_23014));
NAND2X1 g113586(.A (n_23008), .B (n_27999), .Y (n_23013));
NAND2X1 g113592(.A (n_23002), .B (n_24446), .Y (n_23012));
NAND2X1 g113593(.A (n_22999), .B (n_24446), .Y (n_23011));
NAND2X1 g113602(.A (n_22289), .B (n_8303), .Y (n_23010));
NAND2X1 g113603(.A (n_23008), .B (n_23007), .Y (n_23009));
NAND2X1 g113611(.A (n_23005), .B (n_25302), .Y (n_23006));
NAND2X1 g113622(.A (n_23008), .B (n_32652), .Y (n_23004));
NAND2X1 g113626(.A (n_23002), .B (n_23001), .Y (n_23003));
NAND2X1 g113628(.A (n_22999), .B (n_34688), .Y (n_23000));
NAND2X1 g113639(.A (n_23008), .B (n_25290), .Y (n_22998));
INVX1 g113643(.A (n_22996), .Y (n_22997));
NAND2X1 g113647(.A (n_23005), .B (n_22994), .Y (n_22995));
NAND2X1 g113649(.A (n_22980), .B (n_23149), .Y (n_22993));
NAND3X1 g113652(.A (n_21049), .B (n_22270), .C (n_16655), .Y(n_22992));
NAND2X1 g113656(.A (n_22990), .B (n_22914), .Y (n_22991));
NAND2X1 g113660(.A (n_22600), .B (n_32847), .Y (n_22989));
NAND2X1 g113673(.A (n_22987), .B (n_28158), .Y (n_22988));
AOI21X1 g113676(.A0 (n_21844), .A1 (n_22948), .B0 (n_22985), .Y(n_22986));
NAND2X1 g113683(.A (n_22987), .B (n_26238), .Y (n_22982));
NAND2X1 g113697(.A (n_22980), .B (n_22080), .Y (n_22981));
NAND2X1 g113703(.A (n_23350), .B (n_22978), .Y (n_22979));
NAND2X1 g113704(.A (n_22295), .B (n_19056), .Y (n_22977));
NAND2X1 g113705(.A (n_23005), .B (n_18137), .Y (n_22976));
AOI21X1 g113713(.A0 (n_20843), .A1 (n_35934), .B0 (n_22539), .Y(n_23262));
NAND2X1 g113715(.A (n_22987), .B (n_8954), .Y (n_22974));
NAND3X1 g113717(.A (n_21871), .B (n_21916), .C (n_20609), .Y(n_23552));
INVX1 g113718(.A (n_22972), .Y (n_22973));
NAND2X1 g113729(.A (n_22970), .B (n_20324), .Y (n_22971));
INVX1 g113730(.A (n_34450), .Y (n_22969));
NAND2X1 g113735(.A (n_22580), .B (n_18501), .Y (n_22967));
OAI21X1 g113746(.A0 (n_22538), .A1 (n_32363), .B0 (n_22150), .Y(n_22966));
NOR2X1 g113752(.A (n_18724), .B (n_22615), .Y (n_22965));
NAND2X1 g113756(.A (n_22325), .B (n_22355), .Y (n_22964));
NAND2X1 g113757(.A (n_21897), .B (n_22962), .Y (n_22963));
AOI21X1 g113765(.A0 (n_27100), .A1 (n_22312), .B0 (n_22288), .Y(n_22961));
NAND2X1 g113772(.A (n_22330), .B (n_22960), .Y (n_23581));
INVX1 g113777(.A (n_22958), .Y (n_22959));
NAND2X1 g113782(.A (n_22310), .B (n_21616), .Y (n_23249));
NAND2X1 g113789(.A (n_22315), .B (n_18221), .Y (n_22957));
AOI21X1 g113793(.A0 (n_34386), .A1 (n_20763), .B0 (n_22294), .Y(n_22956));
AOI21X1 g113794(.A0 (n_22246), .A1 (n_19261), .B0 (n_20272), .Y(n_22955));
NAND2X1 g113798(.A (n_22342), .B (n_22954), .Y (n_23603));
NAND2X1 g113804(.A (n_22339), .B (n_22953), .Y (n_23591));
NAND2X1 g113812(.A (n_22320), .B (n_22952), .Y (n_23573));
NAND2X1 g113829(.A (n_22318), .B (n_23638), .Y (n_22951));
AOI21X1 g113848(.A0 (n_22344), .A1 (n_18948), .B0 (n_22345), .Y(n_23901));
XOR2X1 g113853(.A (n_20188), .B (n_22272), .Y (n_23586));
INVX1 g113854(.A (n_22642), .Y (n_22950));
OAI21X1 g113875(.A0 (n_35402), .A1 (n_22949), .B0 (n_22332), .Y(n_23567));
OAI21X1 g113876(.A0 (n_22948), .A1 (n_22947), .B0 (n_22319), .Y(n_23569));
XOR2X1 g113888(.A (n_18288), .B (n_22259), .Y (n_23606));
XOR2X1 g113890(.A (n_19520), .B (n_22260), .Y (n_23593));
NOR2X1 g113892(.A (n_21552), .B (n_22537), .Y (n_22946));
NAND2X1 g113898(.A (n_33546), .B (n_21891), .Y (n_22945));
INVX1 g113901(.A (n_22943), .Y (n_22944));
INVX1 g113915(.A (n_22941), .Y (n_22942));
INVX1 g113917(.A (n_22939), .Y (n_22940));
NOR2X1 g113950(.A (n_21880), .B (n_22545), .Y (n_22938));
NOR2X1 g113952(.A (n_21878), .B (n_22542), .Y (n_22937));
NAND2X1 g113955(.A (n_34770), .B (n_22933), .Y (n_22936));
NAND2X1 g113957(.A (n_9503), .B (n_22861), .Y (n_22935));
NAND2X1 g113959(.A (n_22933), .B (n_34709), .Y (n_22934));
NAND2X1 g113963(.A (n_22931), .B (n_34709), .Y (n_22932));
NAND2X1 g113964(.A (n_22929), .B (n_34709), .Y (n_22930));
NAND2X1 g113966(.A (n_22933), .B (n_25980), .Y (n_22928));
NAND2X1 g113971(.A (n_22931), .B (n_29199), .Y (n_22927));
NAND2X1 g113973(.A (n_22929), .B (n_29199), .Y (n_22926));
NAND2X1 g113979(.A (n_22921), .B (n_27089), .Y (n_22925));
NAND2X1 g113992(.A (n_21891), .B (n_24629), .Y (n_22924));
NAND2X1 g114005(.A (n_22921), .B (n_25554), .Y (n_22922));
NAND2X1 g114025(.A (n_22921), .B (n_26965), .Y (n_22920));
NAND3X1 g114035(.A (n_23478), .B (n_22918), .C (n_22917), .Y(n_22919));
NAND3X1 g114036(.A (n_23252), .B (n_22915), .C (n_22914), .Y(n_22916));
NAND2X1 g114051(.A (n_22921), .B (n_26637), .Y (n_22913));
NAND2X1 g114055(.A (n_23478), .B (n_23477), .Y (n_22912));
NAND2X1 g114059(.A (n_23252), .B (n_23476), .Y (n_22911));
NAND2X1 g114060(.A (n_21601), .B (n_22910), .Y (n_23501));
NAND2X1 g114061(.A (n_14356), .B (n_22908), .Y (n_22909));
NAND2X1 g114069(.A (n_21600), .B (n_22908), .Y (n_23496));
NAND2X1 g114083(.A (n_22283), .B (n_21835), .Y (n_23233));
AND2X1 g114084(.A (n_22560), .B (n_22906), .Y (n_22907));
AOI21X1 g114086(.A0 (n_20619), .A1 (n_28347), .B0 (n_22525), .Y(n_22905));
NOR2X1 g114087(.A (n_21083), .B (n_22524), .Y (n_22904));
NOR2X1 g114096(.A (n_22902), .B (n_25881), .Y (n_22903));
NAND2X1 g114113(.A (n_22262), .B (n_22541), .Y (n_22901));
AOI21X1 g114117(.A0 (n_22182), .A1 (n_19720), .B0 (n_21674), .Y(n_22900));
INVX1 g114118(.A (n_22898), .Y (n_22899));
INVX1 g114137(.A (n_22896), .Y (n_22897));
NOR2X1 g114148(.A (n_21094), .B (n_22529), .Y (n_22895));
NAND2X1 g114153(.A (n_22550), .B (n_21926), .Y (n_23223));
AOI21X1 g114160(.A0 (n_22181), .A1 (n_32847), .B0 (n_22191), .Y(n_22894));
NAND2X1 g114191(.A (n_22551), .B (n_21622), .Y (n_23222));
NAND2X1 g114211(.A (n_22563), .B (n_21718), .Y (n_22888));
NAND3X1 g114212(.A (n_22222), .B (n_22869), .C (n_21717), .Y(n_22887));
INVX1 g114217(.A (n_23527), .Y (n_22886));
XOR2X1 g114229(.A (n_17873), .B (n_22215), .Y (n_23510));
NOR2X1 g114280(.A (n_17123), .B (n_22852), .Y (n_22884));
NAND2X1 g114347(.A (n_22204), .B (n_34386), .Y (n_22883));
INVX1 g114354(.A (n_22878), .Y (n_22879));
NAND3X1 g114362(.A (n_22179), .B (n_22517), .C (n_20781), .Y(n_22877));
NAND2X1 g114371(.A (n_22200), .B (n_22875), .Y (n_22876));
INVX1 g114428(.A (n_22873), .Y (n_22874));
AOI21X1 g114430(.A0 (n_22147), .A1 (n_20957), .B0 (n_22871), .Y(n_32621));
NAND2X1 g114439(.A (n_20470), .B (n_22869), .Y (n_22870));
NOR2X1 g114440(.A (n_22203), .B (n_21750), .Y (n_24841));
NAND2X1 g114441(.A (n_22232), .B (n_22867), .Y (n_22868));
NOR2X1 g114443(.A (n_21743), .B (n_22218), .Y (n_22866));
NAND2X1 g114446(.A (n_20501), .B (n_22864), .Y (n_22865));
NAND2X1 g114453(.A (n_21532), .B (n_22148), .Y (n_23229));
INVX1 g114457(.A (n_22862), .Y (n_22863));
INVX1 g114482(.A (n_22861), .Y (n_23208));
AOI22X1 g114512(.A0 (n_22152), .A1 (n_20840), .B0 (n_19530), .B1(n_20839), .Y (n_22859));
AOI22X1 g114513(.A0 (n_22618), .A1 (n_22857), .B0 (n_19543), .B1(n_20488), .Y (n_22858));
INVX1 g114520(.A (n_22532), .Y (n_22856));
NAND2X1 g114665(.A (n_20912), .B (n_22854), .Y (n_22855));
INVX1 g114717(.A (n_22505), .Y (n_24170));
INVX1 g114728(.A (n_22852), .Y (n_22853));
INVX1 g114756(.A (n_22502), .Y (n_22851));
NAND2X1 g109733(.A (n_22086), .B (n_9431), .Y (n_22850));
NAND2X1 g115452(.A (n_9629), .B (n_22093), .Y (n_22849));
NAND2X1 g115500(.A (n_9629), .B (n_22096), .Y (n_22848));
NOR2X1 g115755(.A (n_20727), .B (n_22092), .Y (n_22846));
XOR2X1 g110255(.A (n_16172), .B (n_21655), .Y (n_23308));
NAND2X1 g111018(.A (n_22084), .B (n_22844), .Y (n_22845));
NAND2X1 g111021(.A (n_22082), .B (n_22842), .Y (n_22843));
XOR2X1 g111087(.A (n_19085), .B (n_21653), .Y (n_23458));
OAI21X1 g111507(.A0 (n_21645), .A1 (n_26052), .B0 (n_15083), .Y(n_22841));
NAND2X1 g112298(.A (n_22075), .B (n_22839), .Y (n_22840));
OAI21X1 g112300(.A0 (n_21643), .A1 (n_32748), .B0 (n_24897), .Y(n_22838));
OAI21X1 g112302(.A0 (n_21643), .A1 (n_22042), .B0 (n_22836), .Y(n_22837));
NAND2X1 g112582(.A (n_22832), .B (n_25734), .Y (n_22835));
NAND2X1 g112594(.A (n_22044), .B (n_24451), .Y (n_32100));
NAND2X1 g112642(.A (n_22832), .B (n_22831), .Y (n_22833));
NAND2X1 g112655(.A (n_22041), .B (n_23771), .Y (n_35635));
AOI21X1 g112657(.A0 (n_21640), .A1 (n_24324), .B0 (n_26052), .Y(n_22829));
NAND2X1 g112686(.A (n_22045), .B (n_25122), .Y (n_22828));
NAND2X1 g112694(.A (n_22832), .B (n_23457), .Y (n_22826));
NAND2X1 g112761(.A (n_22832), .B (n_13274), .Y (n_22825));
NAND3X1 g112790(.A (n_21107), .B (n_21638), .C (n_18099), .Y(n_22823));
AOI21X1 g112805(.A0 (n_14816), .A1 (n_22821), .B0 (n_22063), .Y(n_22822));
AOI21X1 g112809(.A0 (n_14814), .A1 (n_22821), .B0 (n_22061), .Y(n_22820));
NAND2X1 g112912(.A (n_22065), .B (n_25351), .Y (n_22819));
OAI21X1 g112914(.A0 (n_21637), .A1 (n_32802), .B0 (n_13639), .Y(n_22818));
NAND2X1 g112916(.A (n_22059), .B (n_25344), .Y (n_22815));
NAND2X1 g112917(.A (n_22053), .B (n_25335), .Y (n_22814));
OAI21X1 g112950(.A0 (n_35478), .A1 (n_22006), .B0 (n_22813), .Y(n_23443));
AOI21X1 g112953(.A0 (n_14590), .A1 (n_23176), .B0 (n_22056), .Y(n_22812));
NAND2X1 g113046(.A (n_22155), .B (n_22810), .Y (n_22811));
NAND2X1 g113082(.A (n_22802), .B (n_30563), .Y (n_22809));
NAND2X1 g113083(.A (n_22807), .B (n_34694), .Y (n_22808));
NAND2X1 g113084(.A (n_22805), .B (n_29008), .Y (n_22806));
NAND2X1 g113088(.A (n_27743), .B (n_22800), .Y (n_22804));
NAND2X1 g113091(.A (n_27743), .B (n_22802), .Y (n_22803));
AOI21X1 g113100(.A0 (n_20989), .A1 (n_32932), .B0 (n_22737), .Y(n_23111));
NAND2X1 g113131(.A (n_22800), .B (n_34802), .Y (n_22801));
NAND2X1 g113135(.A (n_22795), .B (n_25309), .Y (n_32062));
NAND2X1 g113136(.A (n_22793), .B (n_26530), .Y (n_22798));
NAND2X1 g113148(.A (n_22802), .B (n_34802), .Y (n_22797));
NAND2X1 g113152(.A (n_22795), .B (n_25297), .Y (n_22796));
NAND2X1 g113153(.A (n_22793), .B (n_22792), .Y (n_22794));
OAI21X1 g113155(.A0 (n_21630), .A1 (n_21587), .B0 (n_34731), .Y(n_22791));
NAND4X1 g113163(.A (n_18623), .B (n_20662), .C (n_20674), .D(n_21136), .Y (n_22790));
NAND2X1 g113170(.A (n_22807), .B (n_34802), .Y (n_22789));
NAND2X1 g113186(.A (n_22805), .B (n_34802), .Y (n_22788));
NAND2X1 g113191(.A (n_22793), .B (n_22786), .Y (n_22787));
NAND2X1 g113193(.A (n_22795), .B (n_24984), .Y (n_22785));
NAND2X1 g113210(.A (n_21178), .B (n_22719), .Y (n_22784));
AOI21X1 g113220(.A0 (n_21032), .A1 (n_35305), .B0 (n_22424), .Y(n_23082));
NAND2X1 g113221(.A (n_35324), .B (n_20566), .Y (n_22783));
NAND2X1 g113234(.A (n_24965), .B (n_22781), .Y (n_22782));
NAND2X1 g113240(.A (n_35816), .B (n_22781), .Y (n_23398));
NAND2X1 g113243(.A (n_22773), .B (n_33738), .Y (n_22780));
NAND2X1 g113245(.A (n_22779), .B (n_22778), .Y (n_23395));
NAND2X1 g113246(.A (n_14382), .B (n_22775), .Y (n_22777));
NAND2X1 g113257(.A (n_22776), .B (n_22775), .Y (n_23390));
NAND2X1 g113280(.A (n_22773), .B (n_28158), .Y (n_22774));
NAND2X1 g113281(.A (n_22773), .B (n_28374), .Y (n_22772));
NAND2X1 g113291(.A (n_22368), .B (n_33738), .Y (n_22771));
NAND2X1 g113293(.A (n_22768), .B (n_30636), .Y (n_22770));
NAND2X1 g113294(.A (n_25877), .B (n_22781), .Y (n_23400));
NAND2X1 g113298(.A (n_22768), .B (n_29405), .Y (n_22769));
NAND2X1 g113299(.A (n_22766), .B (n_32320), .Y (n_32235));
NAND2X1 g113307(.A (n_22768), .B (n_33738), .Y (n_22765));
AOI21X1 g113335(.A0 (n_24925), .A1 (n_22389), .B0 (n_22017), .Y(n_22764));
AOI21X1 g113336(.A0 (n_14856), .A1 (n_22375), .B0 (n_22762), .Y(n_22763));
NAND4X1 g113350(.A (n_22018), .B (n_18100), .C (n_18088), .D(n_19967), .Y (n_22761));
NAND2X1 g113373(.A (n_22037), .B (n_22760), .Y (n_23424));
NAND2X1 g113390(.A (n_22034), .B (n_22844), .Y (n_23420));
NAND2X1 g113400(.A (n_22031), .B (n_22759), .Y (n_23415));
NAND2X1 g113404(.A (n_22020), .B (n_22758), .Y (n_23407));
NAND2X1 g113406(.A (n_22028), .B (n_22842), .Y (n_23404));
NAND2X1 g113408(.A (n_22035), .B (n_23381), .Y (n_22757));
NOR2X1 g113412(.A (n_22029), .B (n_17012), .Y (n_23035));
NAND2X1 g113422(.A (n_22030), .B (n_28364), .Y (n_22756));
MX2X1 g113453(.A (n_17933), .B (n_17932), .S0 (n_34557), .Y(n_23027));
XOR2X1 g113465(.A (n_16891), .B (n_35305), .Y (n_23397));
XOR2X1 g113470(.A (n_19205), .B (n_22688), .Y (n_23412));
INVX1 g113495(.A (n_23153), .Y (n_22754));
AOI21X1 g113502(.A0 (n_21476), .A1 (n_21931), .B0 (n_21789), .Y(n_22753));
NAND2X1 g113505(.A (n_33546), .B (n_22711), .Y (n_22752));
NAND2X1 g113507(.A (n_33546), .B (n_22676), .Y (n_22751));
NAND2X1 g113509(.A (n_33546), .B (n_22702), .Y (n_22750));
NOR2X1 g113510(.A (n_21935), .B (n_11113), .Y (n_22749));
NOR2X1 g113512(.A (n_17282), .B (n_21934), .Y (n_22748));
NAND2X1 g113514(.A (n_33546), .B (n_22691), .Y (n_22747));
NAND2X1 g113516(.A (n_22002), .B (n_22745), .Y (n_22746));
INVX1 g113519(.A (n_22743), .Y (n_32204));
INVX1 g113521(.A (n_22741), .Y (n_32905));
INVX1 g113524(.A (n_34605), .Y (n_22740));
NAND2X1 g113527(.A (n_22737), .B (n_33025), .Y (n_22738));
NAND2X1 g113529(.A (n_22300), .B (n_35414), .Y (n_22736));
NAND2X1 g113532(.A (n_22670), .B (n_20502), .Y (n_22735));
INVX1 g113533(.A (n_23057), .Y (n_22734));
OAI21X1 g113536(.A0 (n_34683), .A1 (n_34445), .B0 (n_21739), .Y(n_22733));
NAND2X1 g113538(.A (n_22723), .B (n_28864), .Y (n_22731));
NAND2X1 g113539(.A (n_22721), .B (n_29061), .Y (n_22730));
INVX1 g113542(.A (n_22728), .Y (n_22729));
NAND2X1 g113545(.A (n_22726), .B (n_27340), .Y (n_22727));
NAND2X1 g113546(.A (n_22716), .B (n_30563), .Y (n_22725));
NAND2X1 g113548(.A (n_22723), .B (n_28485), .Y (n_22724));
NAND2X1 g113549(.A (n_22721), .B (n_28485), .Y (n_22722));
NAND2X1 g113551(.A (n_22719), .B (n_20048), .Y (n_22720));
NAND2X1 g113556(.A (n_22726), .B (n_29604), .Y (n_22718));
NAND2X1 g113558(.A (n_22716), .B (n_26535), .Y (n_22717));
NAND2X1 g113561(.A (n_22723), .B (n_30197), .Y (n_22715));
NAND2X1 g113563(.A (n_22721), .B (n_28468), .Y (n_22714));
AOI21X1 g113569(.A0 (n_20947), .A1 (n_22008), .B0 (n_22634), .Y(n_23018));
NAND2X2 g113571(.A (n_22296), .B (n_32601), .Y (n_22713));
NAND2X1 g113572(.A (n_22711), .B (n_24629), .Y (n_22712));
NAND2X1 g113573(.A (n_22711), .B (n_25968), .Y (n_22710));
NAND2X1 g113584(.A (n_22704), .B (n_22414), .Y (n_22709));
NAND2X1 g113590(.A (n_32433), .B (n_22706), .Y (n_22708));
NAND2X1 g113601(.A (n_22704), .B (n_18384), .Y (n_22705));
NAND2X1 g113608(.A (n_22702), .B (n_24629), .Y (n_22703));
NAND2X1 g113609(.A (n_22702), .B (n_25968), .Y (n_22701));
NAND2X1 g113619(.A (n_22704), .B (n_32815), .Y (n_22700));
AOI21X1 g113620(.A0 (n_21581), .A1 (n_23039), .B0 (n_8065), .Y(n_22698));
INVX1 g113630(.A (n_22696), .Y (n_22697));
NAND2X1 g113636(.A (n_22704), .B (n_25402), .Y (n_32076));
AOI21X1 g113637(.A0 (n_21915), .A1 (n_23046), .B0 (n_26052), .Y(n_22694));
NAND2X1 g113642(.A (n_22691), .B (n_30180), .Y (n_22692));
NAND2X1 g113644(.A (n_21948), .B (n_21947), .Y (n_22996));
NAND2X1 g113645(.A (n_22691), .B (n_35044), .Y (n_22690));
NAND2X1 g113650(.A (n_22168), .B (n_22688), .Y (n_22689));
INVX1 g113657(.A (n_22392), .Y (n_22687));
INVX1 g113665(.A (n_33781), .Y (n_22685));
NAND2X1 g113671(.A (n_21989), .B (n_21037), .Y (n_22683));
NAND2X1 g113672(.A (n_32930), .B (n_17378), .Y (n_22682));
NAND2X1 g113675(.A (n_22354), .B (n_21424), .Y (n_22681));
NAND2X1 g113677(.A (n_22302), .B (n_21413), .Y (n_22680));
AOI21X1 g113678(.A0 (n_21842), .A1 (n_22365), .B0 (n_22678), .Y(n_22679));
NAND2X1 g113681(.A (n_22676), .B (n_24629), .Y (n_22677));
NAND2X1 g113682(.A (n_22676), .B (n_25968), .Y (n_22675));
INVX1 g113686(.A (n_22673), .Y (n_22674));
INVX1 g113708(.A (n_23066), .Y (n_22672));
NAND2X1 g113714(.A (n_22670), .B (n_19055), .Y (n_22671));
NAND2X1 g113719(.A (n_21593), .B (n_22000), .Y (n_22972));
NAND3X1 g113720(.A (n_21575), .B (n_21909), .C (n_21539), .Y(n_23626));
AOI21X1 g113721(.A0 (n_21841), .A1 (n_35230), .B0 (n_22668), .Y(n_22669));
NOR2X1 g113745(.A (n_9137), .B (n_21937), .Y (n_22667));
NAND3X1 g113747(.A (n_21951), .B (n_21380), .C (n_35353), .Y(n_22666));
NAND3X1 g113749(.A (n_32198), .B (n_32199), .C (n_19277), .Y(n_32107));
NOR2X1 g113751(.A (n_9106), .B (n_21936), .Y (n_22664));
AOI21X1 g113763(.A0 (n_27100), .A1 (n_22322), .B0 (n_21943), .Y(n_22663));
INVX1 g113770(.A (n_22661), .Y (n_22662));
INVX1 g113775(.A (n_22659), .Y (n_22660));
INVX1 g113778(.A (n_22658), .Y (n_22958));
OAI21X1 g113791(.A0 (n_21888), .A1 (n_26748), .B0 (n_15010), .Y(n_22657));
OAI21X1 g113792(.A0 (n_22650), .A1 (n_14702), .B0 (n_23648), .Y(n_22656));
OAI21X1 g113820(.A0 (n_22652), .A1 (n_23178), .B0 (n_24007), .Y(n_22654));
OAI21X1 g113822(.A0 (n_22652), .A1 (n_32745), .B0 (n_24005), .Y(n_22653));
OAI21X1 g113824(.A0 (n_22650), .A1 (n_13317), .B0 (n_23643), .Y(n_22651));
OAI21X1 g113826(.A0 (n_22650), .A1 (n_14404), .B0 (n_23641), .Y(n_22648));
INVX1 g113830(.A (n_23073), .Y (n_22647));
NAND2X1 g113836(.A (n_21979), .B (n_21969), .Y (n_22646));
NAND2X1 g113838(.A (n_21978), .B (n_21966), .Y (n_22645));
NAND2X1 g113839(.A (n_21977), .B (n_21958), .Y (n_22644));
NAND2X1 g113851(.A (n_21980), .B (n_21997), .Y (n_22643));
XOR2X1 g113852(.A (n_17398), .B (n_22366), .Y (n_23342));
OAI21X1 g113855(.A0 (n_21873), .A1 (n_8965), .B0 (n_18197), .Y(n_22642));
NAND2X1 g113857(.A (n_18211), .B (n_21949), .Y (n_22641));
INVX1 g113864(.A (n_33286), .Y (n_23332));
OAI21X1 g113879(.A0 (n_33611), .A1 (n_22638), .B0 (n_21965), .Y(n_23325));
XOR2X1 g113880(.A (n_18619), .B (n_21912), .Y (n_23344));
NAND3X1 g113893(.A (n_22254), .B (n_21517), .C (n_18223), .Y(n_22637));
NAND2X1 g113896(.A (n_22634), .B (n_21595), .Y (n_22635));
AOI21X1 g113902(.A0 (n_21821), .A1 (n_21857), .B0 (n_22503), .Y(n_22943));
NAND2X1 g113911(.A (n_22273), .B (n_22202), .Y (n_23291));
OAI21X1 g113916(.A0 (n_21818), .A1 (n_20450), .B0 (n_22199), .Y(n_22941));
NAND2X1 g113918(.A (n_22271), .B (n_21907), .Y (n_22939));
AOI21X1 g113920(.A0 (n_22201), .A1 (n_22632), .B0 (n_22498), .Y(n_32902));
NAND3X1 g113923(.A (n_20626), .B (n_18217), .C (n_21866), .Y(n_22631));
INVX1 g113933(.A (n_22629), .Y (n_22630));
AOI21X1 g113937(.A0 (n_21992), .A1 (n_20948), .B0 (n_22213), .Y(n_22628));
INVX1 g113944(.A (n_22626), .Y (n_22627));
NOR2X1 g113948(.A (n_22248), .B (n_21881), .Y (n_22625));
NAND2X1 g113951(.A (n_22623), .B (n_21463), .Y (n_22624));
NAND2X1 g113954(.A (n_21591), .B (n_22184), .Y (n_23254));
AOI21X1 g113974(.A0 (n_21793), .A1 (n_34646), .B0 (n_22530), .Y(n_22622));
NAND2X1 g113975(.A (n_21928), .B (n_20965), .Y (n_35690));
AOI21X1 g113980(.A0 (n_21794), .A1 (n_22619), .B0 (n_22618), .Y(n_22620));
NAND3X1 g113985(.A (n_35631), .B (n_20265), .C (n_21805), .Y(n_22617));
INVX1 g113995(.A (n_22615), .Y (n_22616));
NAND2X1 g114001(.A (n_22236), .B (n_24446), .Y (n_22614));
NAND2X1 g114021(.A (n_22236), .B (n_23001), .Y (n_22613));
NAND2X1 g114027(.A (n_22611), .B (n_22220), .Y (n_22612));
NAND2X1 g114039(.A (n_21526), .B (n_22584), .Y (n_22610));
NAND3X1 g114042(.A (n_18681), .B (n_21433), .C (n_21802), .Y(n_22609));
NAND2X1 g114057(.A (n_22604), .B (n_33738), .Y (n_22608));
NOR2X1 g114076(.A (n_26382), .B (n_22277), .Y (n_22607));
NAND2X1 g114081(.A (n_22604), .B (n_28158), .Y (n_22605));
NAND2X1 g114085(.A (n_22604), .B (n_28374), .Y (n_22603));
INVX1 g114090(.A (n_22970), .Y (n_22602));
INVX1 g114092(.A (n_22600), .Y (n_22601));
NAND2X1 g114095(.A (n_22534), .B (n_33738), .Y (n_22599));
NAND2X1 g114097(.A (n_22596), .B (n_26238), .Y (n_22598));
NAND2X1 g114099(.A (n_22596), .B (n_29405), .Y (n_22597));
NAND2X1 g114102(.A (n_22596), .B (n_33738), .Y (n_22595));
NAND2X1 g114105(.A (n_21122), .B (n_21924), .Y (n_22594));
NAND2X1 g114119(.A (n_22274), .B (n_22234), .Y (n_22898));
AOI21X1 g114124(.A0 (n_22233), .A1 (n_21771), .B0 (n_22592), .Y(n_22593));
NAND3X1 g114126(.A (n_22578), .B (n_21913), .C (n_22577), .Y(n_22591));
AOI21X1 g114127(.A0 (n_35411), .A1 (n_22229), .B0 (n_22589), .Y(n_32236));
AOI21X1 g114128(.A0 (n_21536), .A1 (n_21349), .B0 (n_22521), .Y(n_22588));
INVX1 g114132(.A (n_22586), .Y (n_22587));
NAND2X1 g114138(.A (n_21903), .B (n_22230), .Y (n_22896));
NAND2X1 g114140(.A (n_21527), .B (n_22584), .Y (n_22585));
INVX1 g114149(.A (n_22580), .Y (n_22581));
NAND2X1 g114170(.A (n_21921), .B (n_21942), .Y (n_23286));
NAND2X1 g114178(.A (n_21920), .B (n_21941), .Y (n_23284));
NAND2X1 g114183(.A (n_22275), .B (n_21939), .Y (n_23282));
NAND2X1 g114184(.A (n_22267), .B (n_21940), .Y (n_23280));
NAND4X1 g114188(.A (n_22577), .B (n_22578), .C (n_22561), .D(n_22576), .Y (n_22579));
AOI21X1 g114198(.A0 (n_33613), .A1 (n_22573), .B0 (n_20899), .Y(n_22575));
NAND2X1 g114200(.A (n_22264), .B (n_26548), .Y (n_22572));
XOR2X1 g114219(.A (n_17830), .B (n_21825), .Y (n_23527));
INVX1 g114220(.A (n_22999), .Y (n_22571));
XOR2X1 g114228(.A (n_16563), .B (n_22549), .Y (n_23271));
INVX1 g114239(.A (n_23002), .Y (n_22569));
INVX1 g114245(.A (n_22980), .Y (n_22567));
NOR2X1 g114282(.A (n_22176), .B (n_11319), .Y (n_22565));
AND2X1 g114334(.A (n_22207), .B (n_22500), .Y (n_22564));
NOR2X1 g114341(.A (n_22221), .B (n_22205), .Y (n_22563));
AND2X1 g114355(.A (n_21807), .B (n_19709), .Y (n_22878));
NAND2X1 g114356(.A (n_22577), .B (n_22561), .Y (n_22562));
NAND3X1 g114365(.A (n_21803), .B (n_21849), .C (n_17983), .Y(n_22560));
OR2X1 g114375(.A (n_22558), .B (n_22509), .Y (n_22559));
NAND2X1 g114376(.A (n_22556), .B (n_22506), .Y (n_22557));
NAND2X1 g114389(.A (n_22543), .B (n_20950), .Y (n_22555));
NAND2X1 g114395(.A (n_21861), .B (n_34282), .Y (n_22554));
NAND2X1 g114400(.A (n_18546), .B (n_22548), .Y (n_22551));
NAND2X1 g114405(.A (n_22549), .B (n_20476), .Y (n_22550));
NAND2X1 g114406(.A (n_35736), .B (n_22548), .Y (n_22908));
NAND2X1 g114415(.A (n_21466), .B (n_21822), .Y (n_23478));
NAND2X1 g114422(.A (n_26584), .B (n_22548), .Y (n_22910));
OAI21X1 g114429(.A0 (n_22251), .A1 (n_19201), .B0 (n_21405), .Y(n_22873));
AOI21X1 g114431(.A0 (n_22250), .A1 (n_32366), .B0 (n_22149), .Y(n_22546));
NAND3X1 g114437(.A (n_10188), .B (n_18745), .C (n_21470), .Y(n_22545));
NAND2X1 g114445(.A (n_19993), .B (n_22543), .Y (n_22544));
NAND3X1 g114447(.A (n_10200), .B (n_18663), .C (n_21411), .Y(n_22542));
INVX1 g114451(.A (n_22540), .Y (n_22541));
INVX1 g114454(.A (n_22538), .Y (n_22539));
INVX1 g114458(.A (n_22623), .Y (n_22862));
OAI21X1 g114462(.A0 (n_26382), .A1 (n_19961), .B0 (n_21798), .Y(n_22537));
NAND2X1 g114475(.A (n_21863), .B (n_21890), .Y (n_22933));
NAND2X1 g114483(.A (n_21855), .B (n_21889), .Y (n_22861));
NAND2X1 g114491(.A (n_21848), .B (n_21885), .Y (n_22931));
NAND2X1 g114492(.A (n_21865), .B (n_21892), .Y (n_22929));
AND2X1 g114507(.A (n_21833), .B (n_22369), .Y (n_22535));
INVX1 g114509(.A (n_22534), .Y (n_22902));
NAND2X1 g114515(.A (n_18220), .B (n_21847), .Y (n_22533));
OAI21X1 g114521(.A0 (n_17503), .A1 (n_7985), .B0 (n_21839), .Y(n_22532));
OAI21X1 g114525(.A0 (n_21402), .A1 (n_22528), .B0 (n_18199), .Y(n_22529));
NAND2X1 g114528(.A (n_21845), .B (n_9561), .Y (n_22527));
NAND2X1 g114530(.A (n_21830), .B (n_9551), .Y (n_22526));
OAI21X1 g114531(.A0 (n_17502), .A1 (n_25540), .B0 (n_21831), .Y(n_22525));
NAND2X1 g114532(.A (n_21828), .B (n_18204), .Y (n_22524));
XOR2X1 g114543(.A (n_21398), .B (n_21407), .Y (n_22921));
NOR2X1 g114556(.A (n_17173), .B (n_22154), .Y (n_22523));
INVX1 g114593(.A (n_22521), .Y (n_22522));
NAND3X1 g114604(.A (n_20508), .B (n_21325), .C (n_20010), .Y(n_22520));
AOI21X1 g114610(.A0 (n_19941), .A1 (n_34805), .B0 (n_18256), .Y(n_22519));
NAND2X1 g114644(.A (n_22517), .B (n_33311), .Y (n_22518));
NOR2X1 g114651(.A (n_21785), .B (n_22162), .Y (n_22516));
NOR2X1 g114653(.A (n_22514), .B (n_22160), .Y (n_22515));
NAND4X1 g114655(.A (n_17181), .B (n_21303), .C (n_22512), .D(n_22511), .Y (n_22513));
NOR2X1 g114662(.A (n_22166), .B (n_22509), .Y (n_22510));
NOR2X1 g114667(.A (n_21767), .B (n_22164), .Y (n_22508));
NAND2X1 g114671(.A (n_21734), .B (n_17155), .Y (n_23211));
AND2X1 g114697(.A (n_22745), .B (n_22506), .Y (n_22507));
NAND3X1 g114718(.A (n_21749), .B (n_20469), .C (n_21386), .Y(n_22505));
NAND3X1 g114729(.A (n_21765), .B (n_19604), .C (n_18324), .Y(n_22852));
NAND2X1 g114743(.A (n_21756), .B (n_18418), .Y (n_22985));
INVX1 g114746(.A (n_22503), .Y (n_22504));
AOI21X1 g114757(.A0 (n_22501), .A1 (n_22500), .B0 (n_22156), .Y(n_22502));
INVX1 g114787(.A (n_22498), .Y (n_22499));
INVX1 g114795(.A (n_34823), .Y (n_22497));
AND2X1 g114816(.A (n_21757), .B (n_21290), .Y (n_32218));
NAND2X1 g114830(.A (n_21691), .B (n_21103), .Y (n_22494));
OAI21X1 g114870(.A0 (n_22226), .A1 (n_20916), .B0 (n_19030), .Y(n_23219));
AND2X1 g114881(.A (n_20795), .B (n_21788), .Y (n_32211));
AOI21X1 g114883(.A0 (n_21542), .A1 (n_22491), .B0 (n_32977), .Y(n_22492));
NAND4X1 g114917(.A (n_21223), .B (n_15181), .C (n_20699), .D(n_13965), .Y (n_22490));
INVX1 g114919(.A (n_22489), .Y (n_23206));
NAND4X1 g115194(.A (n_15144), .B (n_13771), .C (n_20708), .D(n_13774), .Y (n_22488));
INVX1 g115219(.A (n_33557), .Y (n_22487));
AOI21X1 g115228(.A0 (n_21235), .A1 (n_21690), .B0 (n_19170), .Y(n_22485));
NAND4X1 g115298(.A (n_13777), .B (n_22482), .C (n_20707), .D(n_14586), .Y (n_22484));
NAND4X1 g115304(.A (n_13769), .B (n_22482), .C (n_14514), .D(n_20704), .Y (n_22483));
NAND4X1 g115305(.A (n_13961), .B (n_15405), .C (n_14763), .D(n_20701), .Y (n_22481));
NAND2X1 g115430(.A (n_21673), .B (n_21694), .Y (n_22480));
NAND2X1 g115456(.A (n_22472), .B (n_21328), .Y (n_22479));
OAI21X1 g115506(.A0 (n_21203), .A1 (n_22477), .B0 (n_20473), .Y(n_22478));
NAND2X1 g115653(.A (n_21671), .B (n_22139), .Y (n_22476));
NOR2X1 g115752(.A (n_10020), .B (n_21668), .Y (n_22475));
NAND2X1 g115756(.A (n_22091), .B (n_21328), .Y (n_22474));
NAND2X1 g115848(.A (n_20864), .B (n_22472), .Y (n_22473));
NAND2X1 g115875(.A (n_21703), .B (n_21665), .Y (n_22471));
NAND2X1 g115889(.A (n_20112), .B (n_22469), .Y (n_22470));
NOR2X1 g115902(.A (n_15023), .B (n_21662), .Y (n_22468));
NOR2X1 g115903(.A (n_15170), .B (n_21661), .Y (n_22467));
NAND3X1 g115926(.A (n_14548), .B (n_14525), .C (n_21216), .Y(n_22466));
NAND3X1 g115931(.A (n_14772), .B (n_14765), .C (n_21210), .Y(n_22465));
INVX1 g115942(.A (n_22099), .Y (n_22464));
INVX1 g111367(.A (n_22083), .Y (n_23453));
XOR2X1 g111827(.A (n_35679), .B (n_21192), .Y (n_23195));
NAND2X1 g111964(.A (n_22459), .B (n_18918), .Y (n_22463));
AOI21X1 g111977(.A0 (n_21189), .A1 (n_23040), .B0 (n_8065), .Y(n_22462));
AOI21X1 g112010(.A0 (n_21188), .A1 (n_23038), .B0 (n_26052), .Y(n_22461));
NAND2X1 g112025(.A (n_22459), .B (n_22786), .Y (n_22460));
AOI21X1 g112043(.A0 (n_21186), .A1 (n_23045), .B0 (n_8065), .Y(n_22458));
NAND2X1 g112254(.A (n_21647), .B (n_22960), .Y (n_22457));
NAND2X1 g112309(.A (n_21650), .B (n_22954), .Y (n_22456));
NAND2X1 g112312(.A (n_21649), .B (n_22953), .Y (n_22455));
NAND2X1 g112313(.A (n_21646), .B (n_22952), .Y (n_22454));
OAI21X1 g112802(.A0 (n_21173), .A1 (n_26052), .B0 (n_15025), .Y(n_22453));
AOI21X1 g112901(.A0 (n_22066), .A1 (n_29411), .B0 (n_19348), .Y(n_35886));
XOR2X1 g112972(.A (n_17399), .B (n_22068), .Y (n_23172));
NAND2X1 g113130(.A (n_22446), .B (n_28441), .Y (n_22451));
NAND2X1 g113141(.A (n_22448), .B (n_24446), .Y (n_22450));
NAND2X1 g113146(.A (n_22448), .B (n_26530), .Y (n_22449));
NAND2X1 g113169(.A (n_22446), .B (n_23149), .Y (n_22447));
NAND2X1 g113174(.A (n_22446), .B (n_13274), .Y (n_22445));
NAND2X1 g113182(.A (n_22448), .B (n_34688), .Y (n_22444));
NAND2X1 g113249(.A (n_22446), .B (n_24101), .Y (n_22443));
NAND2X1 g113357(.A (n_21641), .B (n_22441), .Y (n_22442));
OAI21X1 g113359(.A0 (n_21151), .A1 (n_32812), .B0 (n_24309), .Y(n_22440));
OAI21X1 g113361(.A0 (n_21151), .A1 (n_23178), .B0 (n_24305), .Y(n_22438));
AOI21X1 g113410(.A0 (n_22026), .A1 (n_14626), .B0 (n_29725), .Y(n_22437));
AOI21X1 g113429(.A0 (n_21985), .A1 (n_26162), .B0 (n_19463), .Y(n_22436));
AOI21X1 g113430(.A0 (n_21983), .A1 (n_34952), .B0 (n_19462), .Y(n_22435));
INVX1 g113448(.A (n_23164), .Y (n_22434));
XOR2X1 g113464(.A (n_19629), .B (n_33558), .Y (n_23150));
XOR2X1 g113496(.A (n_19474), .B (n_21156), .Y (n_23153));
NAND2X1 g113501(.A (n_21605), .B (n_19445), .Y (n_22432));
NAND2X1 g113506(.A (n_24563), .B (n_22417), .Y (n_22431));
NAND2X1 g113508(.A (n_24563), .B (n_22410), .Y (n_22430));
NAND2X1 g113511(.A (n_24563), .B (n_22402), .Y (n_22429));
NAND2X1 g113513(.A (n_24563), .B (n_22396), .Y (n_22428));
NAND2X2 g113520(.A (n_35306), .B (n_21031), .Y (n_22743));
NAND2X2 g113522(.A (n_32933), .B (n_34068), .Y (n_22741));
NAND2X1 g113528(.A (n_22424), .B (n_33857), .Y (n_22425));
NAND2X1 g113531(.A (n_27614), .B (n_22376), .Y (n_22423));
NAND2X2 g113534(.A (n_21950), .B (n_21404), .Y (n_23057));
NAND2X1 g113543(.A (n_21508), .B (n_22001), .Y (n_22728));
NAND3X1 g113554(.A (n_20672), .B (n_21140), .C (n_20676), .Y(n_22422));
NAND3X1 g113557(.A (n_20666), .B (n_21138), .C (n_20675), .Y(n_22421));
NAND3X1 g113562(.A (n_20658), .B (n_21134), .C (n_20673), .Y(n_22420));
NAND2X1 g113566(.A (n_20032), .B (n_21988), .Y (n_23368));
NAND3X1 g113570(.A (n_21557), .B (n_21559), .C (n_21886), .Y(n_22419));
NAND2X1 g113581(.A (n_22417), .B (n_24526), .Y (n_22418));
NAND2X1 g113582(.A (n_22417), .B (n_28798), .Y (n_22416));
NAND2X1 g113583(.A (n_22407), .B (n_22414), .Y (n_22415));
NAND2X1 g113589(.A (n_22404), .B (n_22412), .Y (n_22413));
NAND2X1 g113598(.A (n_22410), .B (n_26106), .Y (n_22411));
NAND2X1 g113599(.A (n_22410), .B (n_26213), .Y (n_22409));
NAND2X1 g113600(.A (n_22407), .B (n_22406), .Y (n_22408));
NAND2X1 g113606(.A (n_22404), .B (n_23007), .Y (n_22405));
AND2X1 g113615(.A (n_22402), .B (n_26213), .Y (n_22403));
NAND2X1 g113617(.A (n_22402), .B (n_34753), .Y (n_22401));
NAND2X1 g113618(.A (n_22407), .B (n_32764), .Y (n_22400));
NAND2X1 g113623(.A (n_22404), .B (n_32728), .Y (n_22399));
NAND2X2 g113631(.A (n_22688), .B (n_22167), .Y (n_22696));
AND2X1 g113632(.A (n_22396), .B (n_26112), .Y (n_22397));
NAND2X1 g113634(.A (n_22396), .B (n_24526), .Y (n_22395));
NAND2X1 g113635(.A (n_22407), .B (n_25404), .Y (n_35261));
NAND2X1 g113640(.A (n_22404), .B (n_26866), .Y (n_32212));
AOI21X1 g113658(.A0 (n_19333), .A1 (n_21143), .B0 (n_20024), .Y(n_22392));
NAND2X1 g113684(.A (n_29430), .B (n_22389), .Y (n_22390));
NAND2X1 g113685(.A (n_22012), .B (n_22378), .Y (n_23080));
NAND2X1 g113687(.A (n_24965), .B (n_22380), .Y (n_22673));
NAND2X1 g113690(.A (n_32932), .B (n_21501), .Y (n_22388));
NAND2X1 g113691(.A (n_22385), .B (n_8990), .Y (n_22387));
NAND2X1 g113693(.A (n_22385), .B (n_27522), .Y (n_22386));
NAND2X1 g113699(.A (n_22383), .B (n_29505), .Y (n_22384));
NAND2X1 g113700(.A (n_22383), .B (n_29430), .Y (n_22382));
NAND2X1 g113702(.A (n_35794), .B (n_22380), .Y (n_22381));
NAND2X1 g113706(.A (n_22378), .B (n_14642), .Y (n_22379));
NAND2X2 g113709(.A (n_21990), .B (n_20976), .Y (n_23066));
NAND2X1 g113710(.A (n_24925), .B (n_22376), .Y (n_22377));
NAND2X1 g113711(.A (n_22375), .B (n_21168), .Y (n_23062));
NAND2X1 g113739(.A (n_35540), .B (n_22380), .Y (n_23060));
OAI21X1 g113750(.A0 (n_22373), .A1 (n_34601), .B0 (n_20978), .Y(n_22374));
NAND2X1 g113768(.A (n_21620), .B (n_27522), .Y (n_22372));
NAND3X1 g113769(.A (n_32590), .B (n_32591), .C (n_32125), .Y(n_32969));
OAI21X1 g113771(.A0 (n_32302), .A1 (n_32325), .B0 (n_21635), .Y(n_22661));
NAND3X1 g113776(.A (n_21578), .B (n_21577), .C (n_21067), .Y(n_22659));
NAND2X1 g113779(.A (n_21632), .B (n_20596), .Y (n_22658));
INVX1 g113799(.A (n_22800), .Y (n_22371));
NAND2X1 g113801(.A (n_21628), .B (n_22016), .Y (n_23102));
NAND2X1 g113803(.A (n_21626), .B (n_22015), .Y (n_23098));
OAI21X1 g113808(.A0 (n_21544), .A1 (n_32662), .B0 (n_22013), .Y(n_23091));
NAND2X1 g113810(.A (n_21624), .B (n_14089), .Y (n_23086));
AOI21X1 g113816(.A0 (n_22369), .A1 (n_17904), .B0 (n_21608), .Y(n_22370));
INVX1 g113818(.A (n_22368), .Y (n_23055));
NAND4X1 g113823(.A (n_22366), .B (n_19084), .C (n_16173), .D(n_19523), .Y (n_22367));
NAND2X1 g113831(.A (n_21614), .B (n_22027), .Y (n_23073));
NAND2X1 g113835(.A (n_21623), .B (n_22024), .Y (n_23069));
INVX1 g113866(.A (n_22795), .Y (n_22364));
INVX1 g113868(.A (n_22793), .Y (n_22363));
INVX1 g113873(.A (n_22362), .Y (n_23071));
XOR2X1 g113881(.A (n_22361), .B (n_32325), .Y (n_23096));
XOR2X1 g113883(.A (n_17505), .B (n_23255), .Y (n_23094));
XOR2X1 g113887(.A (n_18917), .B (n_21556), .Y (n_23100));
NOR2X1 g113894(.A (n_21796), .B (n_20057), .Y (n_22359));
NAND2X1 g113905(.A (n_33546), .B (n_22335), .Y (n_22358));
OAI21X1 g113910(.A0 (n_20609), .A1 (n_21464), .B0 (n_21815), .Y(n_22990));
NAND2X1 g113912(.A (n_21910), .B (n_21505), .Y (n_23295));
NAND2X1 g113919(.A (n_33546), .B (n_22327), .Y (n_22357));
AOI21X1 g113921(.A0 (n_21996), .A1 (n_20920), .B0 (n_22189), .Y(n_22356));
INVX1 g113928(.A (n_22354), .Y (n_22355));
OAI21X1 g113934(.A0 (n_21993), .A1 (n_19871), .B0 (n_21495), .Y(n_22629));
AOI21X1 g113935(.A0 (n_21810), .A1 (n_21421), .B0 (n_22352), .Y(n_22353));
AOI21X1 g113936(.A0 (n_21497), .A1 (n_33027), .B0 (n_22186), .Y(n_22351));
NAND2X1 g113938(.A (n_33546), .B (n_22308), .Y (n_22350));
NAND2X1 g113945(.A (n_21569), .B (n_21811), .Y (n_22626));
NAND2X1 g113946(.A (n_28874), .B (n_22276), .Y (n_22349));
NOR2X1 g113949(.A (n_21547), .B (n_21895), .Y (n_22348));
NOR2X1 g113953(.A (n_21546), .B (n_21894), .Y (n_22347));
NAND2X1 g113972(.A (n_21927), .B (n_35126), .Y (n_23350));
NAND2X1 g113977(.A (n_21925), .B (n_20959), .Y (n_22346));
NOR2X1 g113978(.A (n_22344), .B (n_18948), .Y (n_22345));
NAND2X1 g113981(.A (n_22338), .B (n_25098), .Y (n_22342));
NAND2X1 g113983(.A (n_21923), .B (n_21382), .Y (n_22341));
NAND3X1 g113996(.A (n_32978), .B (n_21543), .C (n_22340), .Y(n_22615));
NAND2X1 g114003(.A (n_22338), .B (n_18498), .Y (n_22339));
AND2X1 g114012(.A (n_22335), .B (n_24629), .Y (n_22336));
NAND2X1 g114013(.A (n_22335), .B (n_28431), .Y (n_22333));
NAND2X1 g114022(.A (n_35402), .B (n_22949), .Y (n_22332));
NAND2X1 g114024(.A (n_22338), .B (n_22994), .Y (n_22330));
AND2X1 g114028(.A (n_21887), .B (n_19880), .Y (n_22329));
NAND2X1 g114031(.A (n_22327), .B (n_24629), .Y (n_22328));
NAND2X1 g114032(.A (n_22327), .B (n_25968), .Y (n_22326));
NAND2X1 g114038(.A (n_22948), .B (n_21024), .Y (n_22325));
NAND2X1 g114041(.A (n_33611), .B (n_21763), .Y (n_22324));
NAND2X1 g114043(.A (n_27462), .B (n_22322), .Y (n_22323));
NAND2X1 g114052(.A (n_22338), .B (n_25193), .Y (n_22320));
NAND2X1 g114053(.A (n_22948), .B (n_22947), .Y (n_22319));
OR2X1 g114054(.A (n_22650), .B (n_13432), .Y (n_22318));
NAND2X1 g114056(.A (n_22314), .B (n_8990), .Y (n_22316));
NAND2X1 g114058(.A (n_22314), .B (n_27522), .Y (n_22315));
NAND2X1 g114066(.A (n_22312), .B (n_29505), .Y (n_22313));
NAND2X1 g114067(.A (n_22312), .B (n_26132), .Y (n_22311));
NAND2X1 g114071(.A (n_35403), .B (n_19984), .Y (n_22310));
NAND2X1 g114072(.A (n_22308), .B (n_24629), .Y (n_22309));
NAND2X1 g114075(.A (n_22308), .B (n_25968), .Y (n_22307));
AOI21X1 g114088(.A0 (n_16583), .A1 (n_17299), .B0 (n_21902), .Y(n_22306));
NAND2X1 g114089(.A (n_21877), .B (n_21325), .Y (n_22305));
NAND2X2 g114091(.A (n_21906), .B (n_21554), .Y (n_22970));
NAND2X1 g114093(.A (n_21589), .B (n_22180), .Y (n_22600));
NAND2X1 g114106(.A (n_21883), .B (n_21879), .Y (n_22304));
INVX1 g114120(.A (n_21946), .Y (n_23918));
OAI21X1 g114133(.A0 (n_21837), .A1 (n_18634), .B0 (n_20523), .Y(n_22586));
INVX1 g114135(.A (n_22302), .Y (n_22303));
INVX1 g114141(.A (n_22300), .Y (n_22301));
AOI21X1 g114147(.A0 (n_35414), .A1 (n_35415), .B0 (n_22224), .Y(n_22297));
INVX1 g114150(.A (n_22296), .Y (n_22580));
INVX1 g114158(.A (n_22670), .Y (n_22295));
OAI21X1 g114167(.A0 (n_19791), .A1 (n_21326), .B0 (n_22293), .Y(n_22294));
NAND3X1 g114171(.A (n_20743), .B (n_22284), .C (n_18515), .Y(n_22292));
INVX1 g114174(.A (n_22716), .Y (n_22291));
NAND2X1 g114185(.A (n_21585), .B (n_23043), .Y (n_22290));
NAND2X1 g114186(.A (n_21582), .B (n_23041), .Y (n_22289));
AOI21X1 g114187(.A0 (n_22265), .A1 (n_14567), .B0 (n_29725), .Y(n_22288));
NAND3X1 g114193(.A (n_21898), .B (n_22491), .C (n_22286), .Y(n_22287));
OAI21X1 g114204(.A0 (n_35478), .A1 (n_21797), .B0 (n_21617), .Y(n_22987));
OAI21X1 g114215(.A0 (n_21509), .A1 (n_18639), .B0 (n_20569), .Y(n_22962));
XOR2X1 g114222(.A (n_19766), .B (n_21494), .Y (n_22999));
XOR2X1 g114227(.A (n_18599), .B (n_34767), .Y (n_23008));
XOR2X1 g114234(.A (n_22195), .B (n_21493), .Y (n_23005));
XOR2X1 g114241(.A (n_16417), .B (n_22284), .Y (n_23002));
XOR2X1 g114247(.A (n_19179), .B (n_22561), .Y (n_22980));
NAND2X1 g114264(.A (n_21854), .B (n_21820), .Y (n_23252));
NAND2X1 g114266(.A (n_22183), .B (n_21773), .Y (n_22283));
NAND2X1 g114302(.A (n_21478), .B (n_22549), .Y (n_22279));
NAND3X1 g114332(.A (n_21868), .B (n_21020), .C (n_20016), .Y(n_22278));
INVX1 g114339(.A (n_22276), .Y (n_22277));
NAND2X1 g114344(.A (n_22266), .B (n_24361), .Y (n_22275));
NAND2X1 g114348(.A (n_21541), .B (n_21462), .Y (n_22274));
NAND2X1 g114350(.A (n_21998), .B (n_21781), .Y (n_22273));
OR2X1 g114361(.A (n_21522), .B (n_21145), .Y (n_22272));
NAND2X1 g114363(.A (n_21814), .B (n_21776), .Y (n_22271));
INVX1 g114367(.A (n_22269), .Y (n_22270));
NAND2X1 g114373(.A (n_22255), .B (n_17928), .Y (n_22268));
NOR2X1 g114384(.A (n_21869), .B (n_21395), .Y (n_22584));
NAND2X1 g114399(.A (n_22266), .B (n_23329), .Y (n_22267));
NAND2X1 g114402(.A (n_21874), .B (n_22265), .Y (n_22604));
NAND2X1 g114403(.A (n_14358), .B (n_22263), .Y (n_22264));
NAND2X1 g114404(.A (n_22263), .B (n_21875), .Y (n_22596));
NAND2X1 g114414(.A (n_34767), .B (n_34769), .Y (n_22262));
NAND4X1 g114423(.A (n_22258), .B (n_22257), .C (n_21872), .D(n_20796), .Y (n_22260));
NAND3X1 g114433(.A (n_22258), .B (n_20986), .C (n_22257), .Y(n_22259));
NAND2X1 g114442(.A (n_20437), .B (n_22255), .Y (n_22256));
AOI21X1 g114448(.A0 (n_24925), .A1 (n_21516), .B0 (n_21490), .Y(n_22254));
AOI21X1 g114450(.A0 (n_24752), .A1 (n_21838), .B0 (n_17003), .Y(n_22252));
NAND2X1 g114452(.A (n_21512), .B (n_22251), .Y (n_22540));
AOI21X1 g114455(.A0 (n_21403), .A1 (n_35355), .B0 (n_22250), .Y(n_22538));
NAND2X2 g114459(.A (n_21524), .B (n_20613), .Y (n_22623));
NOR3X1 g114467(.A (n_21456), .B (n_21832), .C (n_22249), .Y(n_25593));
NAND3X1 g114468(.A (n_21484), .B (n_20584), .C (n_18770), .Y(n_22248));
INVX1 g114473(.A (n_21891), .Y (n_22536));
AOI21X1 g114478(.A0 (n_22244), .A1 (n_21469), .B0 (n_21486), .Y(n_22247));
AOI21X1 g114489(.A0 (n_21525), .A1 (n_22238), .B0 (n_19876), .Y(n_22246));
AOI21X1 g114493(.A0 (n_22244), .A1 (n_21410), .B0 (n_21485), .Y(n_22245));
AOI21X1 g114506(.A0 (n_34682), .A1 (n_34446), .B0 (n_21738), .Y(n_22243));
NAND2X1 g114510(.A (n_21520), .B (n_21900), .Y (n_22534));
AOI22X1 g114511(.A0 (n_34766), .A1 (n_20497), .B0 (n_20099), .B1(n_19945), .Y (n_22242));
INVX1 g114516(.A (n_22314), .Y (n_22241));
NAND3X1 g114526(.A (n_19416), .B (n_21037), .C (n_20031), .Y(n_22240));
NAND4X1 g114527(.A (n_19742), .B (n_22238), .C (n_22237), .D(n_19781), .Y (n_22239));
INVX1 g114534(.A (n_22652), .Y (n_22236));
INVX1 g114566(.A (n_22233), .Y (n_22234));
NAND2X1 g114571(.A (n_21397), .B (n_33032), .Y (n_22232));
OR2X1 g114576(.A (n_22206), .B (n_20363), .Y (n_22231));
INVX1 g114581(.A (n_22229), .Y (n_22230));
NOR2X1 g114590(.A (n_21327), .B (n_22228), .Y (n_22880));
NAND2X1 g114594(.A (n_21447), .B (n_22226), .Y (n_22521));
NOR2X1 g114595(.A (n_21764), .B (n_21455), .Y (n_22719));
INVX1 g114600(.A (n_22224), .Y (n_22225));
NAND2X1 g114609(.A (n_21929), .B (n_35179), .Y (n_22223));
NOR2X1 g114638(.A (n_22221), .B (n_34384), .Y (n_22222));
NOR2X1 g114652(.A (n_21309), .B (n_22220), .Y (n_23839));
NOR2X1 g114654(.A (n_21777), .B (n_19062), .Y (n_22219));
NAND2X1 g114660(.A (n_21446), .B (n_21445), .Y (n_22218));
AOI21X1 g114684(.A0 (n_20405), .A1 (n_21295), .B0 (n_17699), .Y(n_22216));
INVX1 g114692(.A (n_22619), .Y (n_22215));
AOI21X1 g114710(.A0 (n_20371), .A1 (n_21304), .B0 (n_17701), .Y(n_22214));
NAND2X1 g114737(.A (n_22211), .B (n_22210), .Y (n_22213));
AND2X1 g114738(.A (n_22211), .B (n_22210), .Y (n_22212));
AOI21X1 g114739(.A0 (n_21318), .A1 (n_21744), .B0 (n_20805), .Y(n_32040));
AOI21X1 g114740(.A0 (n_20364), .A1 (n_34599), .B0 (n_17777), .Y(n_22208));
NAND2X1 g114747(.A (n_21468), .B (n_19809), .Y (n_22503));
AOI21X1 g114762(.A0 (n_19828), .A1 (n_20928), .B0 (n_22206), .Y(n_22207));
INVX1 g114763(.A (n_22205), .Y (n_22869));
AOI21X1 g114772(.A0 (n_19270), .A1 (n_18496), .B0 (n_22221), .Y(n_22204));
NAND2X1 g114773(.A (n_21355), .B (n_21105), .Y (n_22203));
INVX1 g114777(.A (n_22201), .Y (n_22202));
INVX1 g114780(.A (n_22199), .Y (n_22200));
OR2X1 g114785(.A (n_21399), .B (n_22197), .Y (n_22198));
NAND4X1 g114786(.A (n_22195), .B (n_20833), .C (n_22194), .D(n_22193), .Y (n_22196));
NAND2X1 g114788(.A (n_21453), .B (n_20813), .Y (n_22498));
INVX1 g114789(.A (n_22191), .Y (n_22192));
INVX1 g114791(.A (n_22189), .Y (n_22190));
INVX1 g114813(.A (n_22188), .Y (n_22864));
INVX1 g114817(.A (n_22186), .Y (n_22187));
NAND2X1 g114821(.A (n_21422), .B (n_20822), .Y (n_22678));
INVX1 g114844(.A (n_22183), .Y (n_22184));
NAND2X1 g114868(.A (n_21479), .B (n_20819), .Y (n_22668));
AOI21X1 g114869(.A0 (n_21783), .A1 (n_21513), .B0 (n_19703), .Y(n_22182));
INVX1 g114871(.A (n_22180), .Y (n_22181));
AOI22X1 g114884(.A0 (n_20809), .A1 (n_33313), .B0 (n_22177), .B1(n_17951), .Y (n_22179));
OAI21X1 g114894(.A0 (n_20837), .A1 (n_35043), .B0 (n_18769), .Y(n_22176));
NAND3X1 g114895(.A (n_19949), .B (n_20965), .C (n_20532), .Y(n_35691));
AND2X1 g114896(.A (n_20251), .B (n_21471), .Y (n_32882));
AND2X1 g114900(.A (n_19202), .B (n_21483), .Y (n_32142));
AND2X1 g114901(.A (n_32613), .B (n_32614), .Y (n_32020));
NAND2X1 g114920(.A (n_20337), .B (n_22171), .Y (n_22489));
AND2X1 g114928(.A (n_21288), .B (n_17526), .Y (n_22170));
NOR2X1 g115026(.A (n_20938), .B (n_22169), .Y (n_22918));
AND2X1 g115038(.A (n_22167), .B (n_20925), .Y (n_22168));
INVX1 g115054(.A (n_22166), .Y (n_23462));
INVX1 g115061(.A (n_22164), .Y (n_22165));
INVX1 g115081(.A (n_22162), .Y (n_22163));
INVX1 g115084(.A (n_22160), .Y (n_22161));
AOI21X1 g115099(.A0 (n_18980), .A1 (n_16748), .B0 (n_21301), .Y(n_22854));
NOR2X1 g115153(.A (n_33024), .B (n_34509), .Y (n_32904));
NAND2X1 g115182(.A (n_22171), .B (n_20621), .Y (n_22158));
INVX1 g115190(.A (n_22156), .Y (n_22157));
INVX1 g115195(.A (n_22154), .Y (n_22155));
INVX1 g115203(.A (n_22152), .Y (n_22153));
INVX1 g115264(.A (n_22149), .Y (n_22150));
INVX1 g115267(.A (n_22147), .Y (n_22148));
NAND4X1 g115300(.A (n_22145), .B (n_22144), .C (n_22143), .D(n_22142), .Y (n_22146));
NAND3X1 g115331(.A (n_15311), .B (n_13770), .C (n_20710), .Y(n_22141));
NAND2X1 g115345(.A (n_21256), .B (n_22139), .Y (n_22140));
NAND2X1 g115386(.A (n_9629), .B (n_21254), .Y (n_22137));
NAND2X1 g115391(.A (n_9629), .B (n_21253), .Y (n_22136));
NAND2X1 g115427(.A (n_9629), .B (n_21252), .Y (n_22135));
NAND2X1 g115431(.A (n_21250), .B (n_22139), .Y (n_22134));
NAND2X1 g115446(.A (n_21703), .B (n_22110), .Y (n_22133));
NAND2X1 g115453(.A (n_9629), .B (n_21249), .Y (n_22132));
NAND2X1 g115454(.A (n_9629), .B (n_21248), .Y (n_22131));
NAND2X1 g115501(.A (n_9629), .B (n_21266), .Y (n_22130));
NAND2X1 g115502(.A (n_9629), .B (n_21265), .Y (n_22129));
NAND2X1 g115510(.A (n_21264), .B (n_21694), .Y (n_22128));
NAND2X1 g115571(.A (n_21261), .B (n_22123), .Y (n_22124));
NAND2X1 g115579(.A (n_21260), .B (n_21694), .Y (n_22122));
NAND2X1 g115647(.A (n_21247), .B (n_22139), .Y (n_22121));
NOR2X1 g115748(.A (n_10020), .B (n_21234), .Y (n_22119));
NAND2X1 g115754(.A (n_21667), .B (n_21328), .Y (n_22117));
NAND3X1 g115803(.A (n_15169), .B (n_13950), .C (n_20702), .Y(n_22115));
NAND2X1 g115814(.A (n_21267), .B (n_22123), .Y (n_22114));
NAND2X1 g115833(.A (n_21257), .B (n_21694), .Y (n_22113));
NAND2X1 g115847(.A (n_22110), .B (n_21328), .Y (n_22111));
NAND2X1 g115874(.A (n_20864), .B (n_22106), .Y (n_22109));
NOR2X1 g115884(.A (n_21664), .B (n_25540), .Y (n_22108));
NAND2X1 g115885(.A (n_22106), .B (n_21328), .Y (n_22107));
NAND2X1 g115888(.A (n_20864), .B (n_22103), .Y (n_22105));
NAND2X1 g115891(.A (n_22103), .B (n_21328), .Y (n_22104));
NAND2X1 g115907(.A (n_13763), .B (n_21242), .Y (n_22102));
NAND2X1 g115934(.A (n_14542), .B (n_21241), .Y (n_22101));
INVX1 g115940(.A (n_21678), .Y (n_22100));
AOI21X1 g115943(.A0 (n_21677), .A1 (n_19494), .B0 (n_21239), .Y(n_22099));
OAI21X1 g116011(.A0 (n_13761), .A1 (n_22097), .B0 (n_21237), .Y(n_22098));
NAND2X1 g116952(.A (n_21204), .B (n_27399), .Y (n_22096));
NAND2X1 g117015(.A (n_21219), .B (n_27388), .Y (n_22095));
NAND2X1 g117018(.A (n_21211), .B (n_24673), .Y (n_22094));
NAND2X1 g117025(.A (n_21207), .B (n_27379), .Y (n_22093));
INVX1 g117190(.A (n_22091), .Y (n_22092));
AOI22X1 g117275(.A0 (n_10573), .A1 (n_10889), .B0 (n_19000), .B1(n_8946), .Y (n_22090));
NAND2X1 g117691(.A (n_20304), .B (n_21199), .Y (n_22089));
NAND2X1 g117749(.A (n_9629), .B (n_21197), .Y (n_22088));
OAI21X1 g111017(.A0 (n_22085), .A1 (n_24312), .B0 (n_22760), .Y(n_22087));
OAI21X1 g111019(.A0 (n_22085), .A1 (n_14702), .B0 (n_22759), .Y(n_22086));
NAND2X1 g111292(.A (n_22081), .B (n_21919), .Y (n_22084));
NAND2X1 g111368(.A (n_21652), .B (n_19744), .Y (n_22083));
NAND2X1 g111405(.A (n_22081), .B (n_22080), .Y (n_22082));
NOR2X1 g112073(.A (n_21451), .B (n_21195), .Y (n_22079));
AOI21X1 g112243(.A0 (n_14853), .A1 (n_22821), .B0 (n_21194), .Y(n_22078));
AOI21X1 g112251(.A0 (n_14848), .A1 (n_22821), .B0 (n_21193), .Y(n_22077));
AOI21X1 g112417(.A0 (n_14621), .A1 (n_23176), .B0 (n_21190), .Y(n_22076));
NAND2X1 g112600(.A (n_22073), .B (n_24446), .Y (n_22075));
NAND2X1 g112661(.A (n_22073), .B (n_22786), .Y (n_22074));
AOI21X1 g112806(.A0 (n_20687), .A1 (n_25942), .B0 (n_14831), .Y(n_22072));
AOI21X1 g112812(.A0 (n_20685), .A1 (n_25220), .B0 (n_14379), .Y(n_22071));
INVX1 g113027(.A (n_22459), .Y (n_22070));
NOR2X1 g113060(.A (n_20274), .B (n_22068), .Y (n_23427));
NAND2X1 g113103(.A (n_22066), .B (n_8954), .Y (n_22067));
NAND2X1 g113139(.A (n_22058), .B (n_22064), .Y (n_22065));
AOI21X1 g113150(.A0 (n_20684), .A1 (n_23534), .B0 (n_8065), .Y(n_22063));
NAND2X1 g113172(.A (n_21171), .B (n_23771), .Y (n_22062));
AOI21X1 g113175(.A0 (n_20682), .A1 (n_23533), .B0 (n_26052), .Y(n_22061));
NAND2X1 g113178(.A (n_22058), .B (n_34688), .Y (n_22059));
NAND2X1 g113188(.A (n_21170), .B (n_25122), .Y (n_22057));
AOI21X1 g113189(.A0 (n_20679), .A1 (n_23545), .B0 (n_8065), .Y(n_22056));
NAND2X1 g113253(.A (n_22066), .B (n_28158), .Y (n_22054));
NAND2X1 g113261(.A (n_22058), .B (n_22052), .Y (n_22053));
NAND2X1 g113270(.A (n_22066), .B (n_26238), .Y (n_22051));
NAND4X1 g113314(.A (n_22039), .B (n_21555), .C (n_21153), .D(n_20300), .Y (n_22050));
NAND2X1 g113320(.A (n_21179), .B (n_23647), .Y (n_22049));
NAND2X1 g113352(.A (n_21183), .B (n_23642), .Y (n_22048));
NAND2X1 g113353(.A (n_21182), .B (n_23640), .Y (n_22047));
NAND2X1 g113354(.A (n_21176), .B (n_23637), .Y (n_22046));
OAI21X1 g113355(.A0 (n_22043), .A1 (n_21169), .B0 (n_14049), .Y(n_22045));
OAI21X1 g113407(.A0 (n_22043), .A1 (n_22042), .B0 (n_23382), .Y(n_22044));
OAI21X1 g113409(.A0 (n_22043), .A1 (n_32646), .B0 (n_23380), .Y(n_22041));
XOR2X1 g113449(.A (n_18561), .B (n_22039), .Y (n_23164));
XOR2X1 g113498(.A (n_17411), .B (n_20049), .Y (n_22832));
NAND2X1 g113575(.A (n_20058), .B (n_21795), .Y (n_22038));
NAND2X1 g113576(.A (n_22033), .B (n_22036), .Y (n_22037));
NAND2X1 g113607(.A (n_21152), .B (n_18384), .Y (n_22035));
NAND2X1 g113610(.A (n_22033), .B (n_22032), .Y (n_22034));
NAND2X1 g113646(.A (n_22033), .B (n_25956), .Y (n_22031));
NAND2X1 g113661(.A (n_14412), .B (n_22023), .Y (n_22030));
NAND2X2 g113664(.A (n_21167), .B (n_21095), .Y (n_22766));
NAND3X1 g113669(.A (n_20045), .B (n_21111), .C (n_21058), .Y(n_35324));
AND2X1 g113688(.A (n_18546), .B (n_22025), .Y (n_22029));
NAND2X1 g113689(.A (n_22033), .B (n_23578), .Y (n_22028));
NAND2X1 g113696(.A (n_22027), .B (n_22026), .Y (n_22773));
NAND2X1 g113698(.A (n_35736), .B (n_22025), .Y (n_22775));
NAND2X1 g113701(.A (n_22024), .B (n_22023), .Y (n_22768));
NOR2X1 g113738(.A (n_16740), .B (n_33558), .Y (n_22022));
NAND2X1 g113740(.A (n_22021), .B (n_22025), .Y (n_22778));
NAND2X1 g113743(.A (n_35578), .B (n_22025), .Y (n_22020));
NAND3X1 g113761(.A (n_21160), .B (n_18200), .C (n_19966), .Y(n_22018));
AOI21X1 g113764(.A0 (n_14795), .A1 (n_21618), .B0 (n_22762), .Y(n_22017));
NAND2X1 g113800(.A (n_22016), .B (n_35252), .Y (n_22800));
NAND2X1 g113802(.A (n_21165), .B (n_22015), .Y (n_22802));
OAI21X1 g113807(.A0 (n_21102), .A1 (n_32803), .B0 (n_22013), .Y(n_22807));
NAND2X1 g113809(.A (n_21162), .B (n_14089), .Y (n_22805));
NAND2X1 g113819(.A (n_21159), .B (n_22012), .Y (n_22368));
NAND4X1 g113845(.A (n_21973), .B (n_17689), .C (n_18515), .D(n_21972), .Y (n_22011));
INVX1 g113862(.A (n_22448), .Y (n_22010));
XOR2X1 g113867(.A (n_18450), .B (n_35934), .Y (n_22795));
XOR2X1 g113869(.A (n_16947), .B (n_22008), .Y (n_22793));
XOR2X1 g113874(.A (n_17037), .B (n_33782), .Y (n_22362));
INVX1 g113877(.A (n_22006), .Y (n_22781));
NAND2X1 g113897(.A (n_24563), .B (n_21970), .Y (n_22005));
NAND2X1 g113899(.A (n_24563), .B (n_21967), .Y (n_22004));
NAND2X1 g113900(.A (n_24563), .B (n_21959), .Y (n_22003));
INVX1 g113903(.A (n_22001), .Y (n_22002));
AOI21X1 g113906(.A0 (n_21504), .A1 (n_21999), .B0 (n_21998), .Y(n_22000));
NAND2X1 g113907(.A (n_24563), .B (n_21956), .Y (n_21997));
AOI21X1 g113914(.A0 (n_21634), .A1 (n_20454), .B0 (n_21996), .Y(n_23050));
NOR2X1 g113922(.A (n_21310), .B (n_21146), .Y (n_21995));
NAND2X1 g113929(.A (n_21113), .B (n_21993), .Y (n_22354));
NAND2X1 g113931(.A (n_21568), .B (n_21498), .Y (n_22737));
AOI21X1 g113932(.A0 (n_21615), .A1 (n_19921), .B0 (n_21992), .Y(n_23047));
INVX1 g113939(.A (n_21990), .Y (n_32199));
INVX1 g113942(.A (n_21988), .Y (n_21989));
NAND2X1 g113956(.A (n_21981), .B (n_28864), .Y (n_21987));
NAND2X1 g113958(.A (n_21985), .B (n_28485), .Y (n_21986));
NAND2X1 g113960(.A (n_21983), .B (n_28485), .Y (n_21984));
NAND2X1 g113961(.A (n_21981), .B (n_28485), .Y (n_21982));
NAND2X1 g113962(.A (n_21975), .B (n_28485), .Y (n_21980));
NAND2X1 g113965(.A (n_21985), .B (n_25424), .Y (n_21979));
NAND2X1 g113967(.A (n_21983), .B (n_25424), .Y (n_21978));
NAND2X1 g113968(.A (n_21981), .B (n_29090), .Y (n_21977));
NAND2X1 g113970(.A (n_21975), .B (n_28468), .Y (n_21976));
NAND2X1 g113984(.A (n_21973), .B (n_21972), .Y (n_21974));
NAND2X1 g113986(.A (n_21970), .B (n_25756), .Y (n_21971));
NAND2X1 g113987(.A (n_21970), .B (n_34753), .Y (n_21969));
NAND2X1 g113993(.A (n_21967), .B (n_25756), .Y (n_21968));
NAND2X1 g113994(.A (n_21967), .B (n_34753), .Y (n_21966));
NAND2X1 g114002(.A (n_33611), .B (n_22638), .Y (n_21965));
NAND2X1 g114004(.A (n_21962), .B (n_26238), .Y (n_21964));
NAND2X1 g114006(.A (n_21962), .B (n_28158), .Y (n_21963));
NAND4X1 g114007(.A (n_21089), .B (n_21043), .C (n_18750), .D(n_20583), .Y (n_21961));
NAND2X1 g114009(.A (n_21959), .B (n_25756), .Y (n_21960));
NAND2X1 g114010(.A (n_21959), .B (n_34753), .Y (n_21958));
AND2X1 g114016(.A (n_21956), .B (n_26112), .Y (n_21957));
NAND2X1 g114017(.A (n_21956), .B (n_24526), .Y (n_21955));
NAND2X1 g114037(.A (n_22365), .B (n_21438), .Y (n_21954));
NAND2X1 g114040(.A (n_35230), .B (n_21442), .Y (n_21953));
INVX1 g114073(.A (n_21950), .Y (n_21951));
NAND2X1 g114080(.A (n_21962), .B (n_33738), .Y (n_21949));
NAND2X1 g114114(.A (n_21911), .B (n_20551), .Y (n_21948));
AOI21X1 g114115(.A0 (n_21538), .A1 (n_21459), .B0 (n_21572), .Y(n_21947));
NAND2X1 g114121(.A (n_21573), .B (n_21537), .Y (n_21946));
AOI21X1 g114122(.A0 (n_21899), .A1 (n_14605), .B0 (n_25376), .Y(n_21945));
NAND2X1 g114136(.A (n_21570), .B (n_21944), .Y (n_22302));
NAND2X1 g114142(.A (n_21567), .B (n_21534), .Y (n_22300));
AOI21X1 g114145(.A0 (n_14801), .A1 (n_21914), .B0 (n_22762), .Y(n_21943));
NAND2X2 g114151(.A (n_21147), .B (n_19972), .Y (n_22296));
NAND2X1 g114155(.A (n_21580), .B (n_21609), .Y (n_22721));
NAND2X2 g114159(.A (n_21561), .B (n_20047), .Y (n_22670));
NAND2X1 g114161(.A (n_20013), .B (n_21876), .Y (n_23024));
NAND2X1 g114169(.A (n_21127), .B (n_21942), .Y (n_22711));
NAND2X1 g114172(.A (n_21126), .B (n_21604), .Y (n_22726));
NAND2X1 g114175(.A (n_21124), .B (n_21603), .Y (n_22716));
NAND2X1 g114177(.A (n_21123), .B (n_21941), .Y (n_22702));
NAND2X1 g114179(.A (n_21564), .B (n_21940), .Y (n_22676));
NAND2X1 g114181(.A (n_21121), .B (n_21602), .Y (n_22723));
NAND2X1 g114182(.A (n_21579), .B (n_21939), .Y (n_22691));
INVX1 g114201(.A (n_22385), .Y (n_21938));
NAND2X1 g114205(.A (n_21131), .B (n_20670), .Y (n_21937));
NAND2X1 g114207(.A (n_20664), .B (n_21130), .Y (n_21936));
OAI21X1 g114208(.A0 (n_20598), .A1 (n_10276), .B0 (n_21129), .Y(n_21935));
NAND2X1 g114209(.A (n_21128), .B (n_20656), .Y (n_21934));
XOR2X1 g114226(.A (n_18601), .B (n_21905), .Y (n_22704));
INVX1 g114231(.A (n_22380), .Y (n_21933));
INVX1 g114248(.A (n_21931), .Y (n_21932));
AOI21X1 g114250(.A0 (n_20983), .A1 (n_20955), .B0 (n_21929), .Y(n_21930));
INVX1 g114270(.A (n_21927), .Y (n_21928));
INVX1 g114272(.A (n_21925), .Y (n_21926));
INVX1 g114274(.A (n_21923), .Y (n_21924));
NAND2X1 g114276(.A (n_21515), .B (n_20525), .Y (n_22634));
NAND3X1 g114286(.A (n_17837), .B (n_18747), .C (n_21026), .Y(n_21922));
NOR2X1 g114295(.A (n_21487), .B (n_18149), .Y (n_22611));
NAND2X1 g114300(.A (n_22266), .B (n_23356), .Y (n_21921));
NAND2X1 g114316(.A (n_22266), .B (n_21919), .Y (n_21920));
NAND2X1 g114326(.A (n_21496), .B (n_21917), .Y (n_21918));
NAND2X1 g114327(.A (n_21819), .B (n_21870), .Y (n_21916));
NAND2X1 g114338(.A (n_21584), .B (n_21185), .Y (n_21915));
NAND2X1 g114340(.A (n_21545), .B (n_21914), .Y (n_22276));
AND2X1 g114342(.A (n_21780), .B (n_21913), .Y (n_22366));
INVX1 g114345(.A (n_21911), .Y (n_21912));
NAND2X1 g114349(.A (n_21592), .B (n_19914), .Y (n_21910));
NAND2X1 g114359(.A (n_21099), .B (n_21574), .Y (n_21909));
NAND2X1 g114368(.A (n_21051), .B (n_35912), .Y (n_22269));
OR2X1 g114372(.A (n_21907), .B (n_21772), .Y (n_21908));
NAND2X1 g114374(.A (n_21905), .B (n_19352), .Y (n_21906));
NAND2X1 g114380(.A (n_19398), .B (n_21901), .Y (n_21904));
NAND2X1 g114385(.A (n_21096), .B (n_21010), .Y (n_21903));
NAND2X1 g114388(.A (n_21901), .B (n_19397), .Y (n_21902));
NAND2X1 g114394(.A (n_21900), .B (n_21899), .Y (n_22322));
NAND3X1 g114416(.A (n_21528), .B (n_19904), .C (n_21529), .Y(n_21898));
NOR2X1 g114424(.A (n_21065), .B (n_19206), .Y (n_21897));
INVX1 g114425(.A (n_21558), .Y (n_21896));
NAND2X1 g114427(.A (n_19418), .B (n_21064), .Y (n_22948));
NAND3X1 g114434(.A (n_9591), .B (n_18763), .C (n_20568), .Y(n_21895));
NAND3X1 g114449(.A (n_9550), .B (n_18656), .C (n_20529), .Y(n_21894));
NAND2X1 g114471(.A (n_21093), .B (n_21892), .Y (n_22308));
NAND2X1 g114474(.A (n_21091), .B (n_21890), .Y (n_21891));
NAND2X1 g114484(.A (n_21088), .B (n_21889), .Y (n_22335));
INVX1 g114485(.A (n_21975), .Y (n_21888));
AOI21X1 g114488(.A0 (n_18185), .A1 (n_21886), .B0 (n_18097), .Y(n_21887));
NAND2X1 g114490(.A (n_21081), .B (n_21885), .Y (n_22327));
AOI21X1 g114494(.A0 (n_26756), .A1 (n_20567), .B0 (n_21046), .Y(n_21884));
AOI21X1 g114495(.A0 (n_26756), .A1 (n_20557), .B0 (n_21045), .Y(n_21883));
AOI21X1 g114497(.A0 (n_26756), .A1 (n_20528), .B0 (n_21044), .Y(n_21882));
NAND3X1 g114498(.A (n_20580), .B (n_20570), .C (n_14587), .Y(n_21881));
NAND3X1 g114500(.A (n_20578), .B (n_20561), .C (n_14809), .Y(n_21880));
NOR2X1 g114501(.A (n_20576), .B (n_21050), .Y (n_21879));
NAND3X1 g114502(.A (n_20575), .B (n_20531), .C (n_14346), .Y(n_21878));
INVX1 g114504(.A (n_21876), .Y (n_21877));
NAND2X1 g114514(.A (n_21076), .B (n_21875), .Y (n_22312));
NAND2X1 g114517(.A (n_21070), .B (n_21874), .Y (n_22314));
INVX1 g114518(.A (n_21962), .Y (n_21873));
AOI21X1 g114533(.A0 (n_17413), .A1 (n_21082), .B0 (n_21078), .Y(n_22650));
XOR2X1 g114536(.A (n_16728), .B (n_21872), .Y (n_22652));
XOR2X1 g114544(.A (n_18640), .B (n_21523), .Y (n_22338));
NAND3X1 g114558(.A (n_21853), .B (n_21870), .C (n_21852), .Y(n_21871));
NAND2X1 g114567(.A (n_21022), .B (n_19337), .Y (n_22233));
OAI21X1 g114570(.A0 (n_21097), .A1 (n_17580), .B0 (n_20835), .Y(n_22592));
INVX1 g114579(.A (n_21869), .Y (n_22543));
NAND2X1 g114582(.A (n_21009), .B (n_19819), .Y (n_22229));
INVX1 g114587(.A (n_21867), .Y (n_21868));
NAND2X1 g114598(.A (n_21846), .B (n_30109), .Y (n_21866));
NAND2X1 g114601(.A (n_21000), .B (n_20803), .Y (n_22224));
NAND2X1 g114605(.A (n_21862), .B (n_23356), .Y (n_21865));
NAND2X1 g114608(.A (n_20980), .B (n_19300), .Y (n_21864));
NAND2X1 g114614(.A (n_21862), .B (n_26315), .Y (n_21863));
INVX1 g114620(.A (n_21860), .Y (n_21861));
NAND3X1 g114627(.A (n_21858), .B (n_21857), .C (n_21856), .Y(n_21859));
NAND2X1 g114629(.A (n_21862), .B (n_22994), .Y (n_21855));
NAND2X1 g114642(.A (n_21853), .B (n_21852), .Y (n_21854));
NAND3X1 g114646(.A (n_18487), .B (n_20448), .C (n_33051), .Y(n_21851));
NAND2X1 g114647(.A (n_21849), .B (n_19589), .Y (n_21850));
NAND2X1 g114650(.A (n_21862), .B (n_24348), .Y (n_21848));
NAND2X1 g114657(.A (n_21846), .B (n_29411), .Y (n_21847));
NAND2X1 g114659(.A (n_24752), .B (n_21846), .Y (n_21845));
NOR2X1 g114675(.A (n_21023), .B (n_21423), .Y (n_21844));
NOR2X1 g114677(.A (n_21437), .B (n_21412), .Y (n_21842));
NOR2X1 g114679(.A (n_21441), .B (n_21408), .Y (n_21841));
NAND2X1 g114691(.A (n_21838), .B (n_8966), .Y (n_21839));
INVX1 g114693(.A (n_21837), .Y (n_22619));
INVX1 g114706(.A (n_21835), .Y (n_21836));
OR2X1 g114712(.A (n_19782), .B (n_21832), .Y (n_21833));
NAND2X1 g114720(.A (n_21829), .B (n_30109), .Y (n_21831));
NAND2X1 g114721(.A (n_24752), .B (n_21829), .Y (n_21830));
NAND2X1 g114723(.A (n_21826), .B (n_29405), .Y (n_21828));
NAND2X1 g114724(.A (n_24752), .B (n_21826), .Y (n_21827));
OR2X1 g114735(.A (n_21039), .B (n_21100), .Y (n_21825));
NAND3X1 g114736(.A (n_20951), .B (n_21823), .C (n_21443), .Y(n_21824));
INVX1 g114744(.A (n_21821), .Y (n_21822));
INVX1 g114751(.A (n_21819), .Y (n_21820));
NAND3X1 g114764(.A (n_16782), .B (n_20468), .C (n_18443), .Y(n_22205));
INVX1 g114769(.A (n_21816), .Y (n_21818));
INVX1 g114774(.A (n_21814), .Y (n_21815));
NAND2X1 g114778(.A (n_21019), .B (n_20815), .Y (n_22201));
AOI21X1 g114781(.A0 (n_20814), .A1 (n_19897), .B0 (n_21452), .Y(n_22199));
NAND2X1 g114790(.A (n_21018), .B (n_21812), .Y (n_22191));
NAND2X1 g114792(.A (n_21017), .B (n_21813), .Y (n_22189));
AOI21X1 g114793(.A0 (n_20812), .A1 (n_19891), .B0 (n_19239), .Y(n_22558));
OAI21X1 g114794(.A0 (n_21812), .A1 (n_18356), .B0 (n_19040), .Y(n_22556));
INVX1 g114807(.A (n_21810), .Y (n_21811));
NAND3X1 g114814(.A (n_17686), .B (n_20512), .C (n_19053), .Y(n_22188));
NAND2X1 g114815(.A (n_20537), .B (n_20817), .Y (n_22352));
NAND2X1 g114818(.A (n_21004), .B (n_20810), .Y (n_22186));
INVX1 g114819(.A (n_33858), .Y (n_21809));
NAND2X1 g114840(.A (n_19351), .B (n_20973), .Y (n_22549));
NAND2X1 g114845(.A (n_21042), .B (n_21040), .Y (n_22183));
NOR2X1 g114872(.A (n_21041), .B (n_21514), .Y (n_22180));
AOI22X1 g114878(.A0 (n_19313), .A1 (n_21806), .B0 (n_22340), .B1(n_16974), .Y (n_21807));
AOI22X1 g114880(.A0 (n_21804), .A1 (n_19942), .B0 (n_20264), .B1(n_18467), .Y (n_21805));
AOI21X1 g114885(.A0 (n_20347), .A1 (n_20318), .B0 (n_19250), .Y(n_21803));
AOI22X1 g114886(.A0 (n_21801), .A1 (n_20395), .B0 (n_19247), .B1(n_18680), .Y (n_21802));
NAND2X1 g114890(.A (n_21029), .B (n_8966), .Y (n_21798));
INVX1 g114910(.A (n_21797), .Y (n_22548));
INVX1 g114923(.A (n_21795), .Y (n_21796));
NOR2X1 g114938(.A (n_20804), .B (n_17240), .Y (n_22517));
NOR2X1 g114964(.A (n_20844), .B (n_21383), .Y (n_21794));
NOR2X1 g114965(.A (n_20480), .B (n_21381), .Y (n_21793));
NOR2X1 g114970(.A (n_21324), .B (n_21033), .Y (n_21792));
NAND2X1 g114978(.A (n_21320), .B (n_21027), .Y (n_35631));
NAND2X1 g114979(.A (n_21789), .B (n_20838), .Y (n_21790));
NAND2X1 g114983(.A (n_21291), .B (n_21787), .Y (n_21788));
INVX1 g115028(.A (n_21785), .Y (n_21786));
AND2X1 g115030(.A (n_21783), .B (n_20929), .Y (n_21784));
AND2X1 g115036(.A (n_21999), .B (n_21781), .Y (n_21782));
AND2X1 g115046(.A (n_21780), .B (n_21779), .Y (n_22577));
INVX1 g115049(.A (n_21777), .Y (n_21778));
NAND2X1 g115055(.A (n_21358), .B (n_20451), .Y (n_22166));
INVX1 g115058(.A (n_21457), .Y (n_22745));
NAND2X1 g115062(.A (n_20927), .B (n_21776), .Y (n_22164));
NOR2X1 g115072(.A (n_21353), .B (n_20921), .Y (n_21775));
NOR2X1 g115078(.A (n_20919), .B (n_20924), .Y (n_21774));
NAND2X1 g115082(.A (n_20918), .B (n_21773), .Y (n_22162));
NOR2X1 g115083(.A (n_21772), .B (n_20922), .Y (n_22914));
NAND2X1 g115085(.A (n_23523), .B (n_21771), .Y (n_22160));
AND2X1 g115087(.A (n_32847), .B (n_21769), .Y (n_21770));
AND2X1 g115096(.A (n_23393), .B (n_22506), .Y (n_21768));
INVX1 g115107(.A (n_21766), .Y (n_21767));
NOR2X1 g115112(.A (n_21177), .B (n_21764), .Y (n_21765));
INVX1 g115116(.A (n_21762), .Y (n_21763));
NAND3X1 g115122(.A (n_21760), .B (n_21759), .C (n_21758), .Y(n_21761));
NAND2X1 g115136(.A (n_21306), .B (n_21428), .Y (n_21757));
NAND2X1 g115147(.A (n_19794), .B (n_18466), .Y (n_21756));
INVX1 g115150(.A (n_21754), .Y (n_21755));
NOR2X1 g115154(.A (n_35396), .B (n_19581), .Y (n_32203));
INVX1 g115162(.A (n_21749), .Y (n_21750));
NAND3X1 g115191(.A (n_21748), .B (n_17239), .C (n_21747), .Y(n_22156));
NAND3X1 g115196(.A (n_20496), .B (n_20194), .C (n_19524), .Y(n_22154));
NAND2X2 g115204(.A (n_20850), .B (n_35708), .Y (n_22152));
NAND2X1 g115205(.A (n_20956), .B (n_19545), .Y (n_22618));
AND2X1 g115206(.A (n_21745), .B (n_21744), .Y (n_21746));
NAND4X1 g115207(.A (n_18354), .B (n_20243), .C (n_21742), .D(n_21741), .Y (n_21743));
AOI21X1 g115218(.A0 (n_33748), .A1 (n_21287), .B0 (n_18930), .Y(n_21740));
NAND2X1 g115265(.A (n_20968), .B (n_20970), .Y (n_22149));
NAND2X1 g115268(.A (n_20966), .B (n_18579), .Y (n_22147));
INVX1 g115287(.A (n_21738), .Y (n_21739));
NAND4X1 g115302(.A (n_21736), .B (n_21735), .C (n_20267), .D(n_25284), .Y (n_21737));
AOI22X1 g115303(.A0 (n_20316), .A1 (n_23212), .B0 (n_18321), .B1(n_21733), .Y (n_21734));
NOR2X1 g115376(.A (n_19548), .B (n_20312), .Y (n_32198));
NAND2X1 g115384(.A (n_21727), .B (n_21328), .Y (n_21731));
AOI21X1 g115409(.A0 (n_20191), .A1 (n_25852), .B0 (n_21374), .Y(n_21730));
AOI21X1 g115411(.A0 (n_20189), .A1 (n_27718), .B0 (n_21374), .Y(n_21729));
NAND2X1 g115424(.A (n_21703), .B (n_21727), .Y (n_21728));
AOI21X1 g115432(.A0 (n_20177), .A1 (n_28325), .B0 (n_10525), .Y(n_21726));
NAND2X1 g115440(.A (n_20771), .B (n_21694), .Y (n_21724));
NAND2X1 g115444(.A (n_21692), .B (n_21328), .Y (n_21723));
AOI21X1 g115466(.A0 (n_20141), .A1 (n_25849), .B0 (n_21374), .Y(n_21722));
AOI21X1 g115473(.A0 (n_20164), .A1 (n_25856), .B0 (n_21374), .Y(n_21721));
AOI21X1 g115483(.A0 (n_20163), .A1 (n_27710), .B0 (n_21374), .Y(n_21720));
AND2X1 g115515(.A (n_21717), .B (n_20175), .Y (n_21718));
NAND2X1 g115534(.A (n_20767), .B (n_21694), .Y (n_21716));
NAND2X1 g115546(.A (n_20766), .B (n_21333), .Y (n_21715));
AOI21X1 g115557(.A0 (n_20149), .A1 (n_25850), .B0 (n_21374), .Y(n_21714));
NAND2X1 g115591(.A (n_20765), .B (n_22139), .Y (n_21712));
NAND2X1 g115615(.A (n_20760), .B (n_21658), .Y (n_21709));
NAND2X1 g115674(.A (n_20864), .B (n_21705), .Y (n_21708));
NAND2X1 g115675(.A (n_21705), .B (n_21328), .Y (n_21706));
NAND2X1 g115730(.A (n_21703), .B (n_21702), .Y (n_21704));
NAND2X1 g115749(.A (n_21233), .B (n_21328), .Y (n_21701));
NAND2X1 g115792(.A (n_20112), .B (n_21698), .Y (n_21700));
NAND2X1 g115793(.A (n_21698), .B (n_21328), .Y (n_21699));
NAND2X1 g115799(.A (n_20762), .B (n_21694), .Y (n_21696));
NAND2X1 g115801(.A (n_20761), .B (n_21694), .Y (n_21695));
NAND2X1 g115832(.A (n_20864), .B (n_21692), .Y (n_21693));
NAND4X1 g115861(.A (n_12174), .B (n_21690), .C (n_20138), .D(n_17677), .Y (n_21691));
NAND2X1 g115863(.A (n_20757), .B (n_21328), .Y (n_21689));
NAND2X1 g115873(.A (n_20864), .B (n_21227), .Y (n_21687));
NAND2X1 g115887(.A (n_20112), .B (n_21682), .Y (n_21685));
NAND2X1 g115890(.A (n_21682), .B (n_21328), .Y (n_21683));
AOI21X1 g115941(.A0 (n_21677), .A1 (n_14496), .B0 (n_20759), .Y(n_21678));
INVX1 g116480(.A (n_21674), .Y (n_21675));
OAI21X1 g117021(.A0 (n_13990), .A1 (n_19523), .B0 (n_28555), .Y(n_21673));
OAI21X1 g117029(.A0 (n_21243), .A1 (n_19523), .B0 (n_28548), .Y(n_21671));
NAND2X1 g117041(.A (n_20732), .B (n_28542), .Y (n_21669));
NAND2X1 g117085(.A (n_20729), .B (n_28125), .Y (n_22472));
INVX1 g117188(.A (n_21667), .Y (n_21668));
NAND2X1 g117191(.A (n_20730), .B (n_21666), .Y (n_22091));
NAND2X1 g117233(.A (n_20746), .B (n_28124), .Y (n_22469));
INVX1 g117243(.A (n_21664), .Y (n_21665));
AOI21X1 g117272(.A0 (n_21217), .A1 (n_10848), .B0 (n_9513), .Y(n_21663));
NAND2X1 g117328(.A (n_14354), .B (n_20723), .Y (n_21662));
NAND2X1 g117329(.A (n_14582), .B (n_20721), .Y (n_21661));
NAND2X1 g117656(.A (n_20695), .B (n_21694), .Y (n_21660));
AOI21X1 g117798(.A0 (n_20065), .A1 (n_28549), .B0 (n_10023), .Y(n_21657));
AOI21X1 g117874(.A0 (n_20064), .A1 (n_28570), .B0 (n_10023), .Y(n_21656));
NAND4X1 g111378(.A (n_21191), .B (n_21450), .C (n_21299), .D(n_21654), .Y (n_21655));
INVX1 g112038(.A (n_21652), .Y (n_21653));
OAI21X1 g112242(.A0 (n_20062), .A1 (n_26052), .B0 (n_15036), .Y(n_21651));
NAND2X1 g112574(.A (n_21648), .B (n_25734), .Y (n_21650));
NAND2X1 g112634(.A (n_21648), .B (n_22831), .Y (n_21649));
NAND2X1 g112688(.A (n_21648), .B (n_23457), .Y (n_21647));
NAND2X1 g112739(.A (n_21648), .B (n_13274), .Y (n_21646));
NOR2X1 g112911(.A (n_20690), .B (n_14309), .Y (n_21645));
XOR2X1 g113029(.A (n_17116), .B (n_22810), .Y (n_22459));
AOI21X1 g113110(.A0 (n_20059), .A1 (n_21942), .B0 (n_8942), .Y(n_21644));
INVX1 g113492(.A (n_22073), .Y (n_21643));
NAND2X1 g113591(.A (n_21639), .B (n_24446), .Y (n_21641));
NAND2X1 g113625(.A (n_21639), .B (n_23001), .Y (n_21640));
OAI21X1 g113814(.A0 (n_20651), .A1 (n_17552), .B0 (n_20615), .Y(n_21638));
XOR2X1 g113849(.A (n_17409), .B (n_21161), .Y (n_22446));
INVX1 g113860(.A (n_22058), .Y (n_21637));
XOR2X1 g113863(.A (n_17259), .B (n_21972), .Y (n_22448));
XOR2X1 g113878(.A (n_18089), .B (n_35230), .Y (n_22006));
AOI21X1 g113904(.A0 (n_20610), .A1 (n_21636), .B0 (n_21590), .Y(n_22001));
AOI21X1 g113908(.A0 (n_21066), .A1 (n_20552), .B0 (n_21634), .Y(n_21635));
AND2X1 g113913(.A (n_21106), .B (n_16268), .Y (n_21633));
NAND2X1 g113925(.A (n_33610), .B (n_21440), .Y (n_21632));
NAND2X2 g113927(.A (n_21114), .B (n_18895), .Y (n_32933));
AND2X1 g113930(.A (n_21104), .B (n_18108), .Y (n_21631));
NAND2X2 g113940(.A (n_22008), .B (n_20946), .Y (n_21990));
NAND4X1 g113941(.A (n_20638), .B (n_20588), .C (n_18756), .D(n_20005), .Y (n_21630));
AOI21X1 g113943(.A0 (n_21063), .A1 (n_20550), .B0 (n_21112), .Y(n_21988));
NAND3X1 g113947(.A (n_18226), .B (n_20627), .C (n_20604), .Y(n_21629));
NAND2X1 g113989(.A (n_21625), .B (n_21627), .Y (n_21628));
NAND2X1 g113998(.A (n_21625), .B (n_14045), .Y (n_21626));
NAND2X2 g114015(.A (n_20655), .B (n_20027), .Y (n_22688));
NAND2X1 g114019(.A (n_21625), .B (n_22786), .Y (n_21624));
NAND2X1 g114029(.A (n_35790), .B (n_21621), .Y (n_21623));
NAND2X1 g114046(.A (n_21622), .B (n_21619), .Y (n_22389));
NAND2X1 g114050(.A (n_13957), .B (n_21621), .Y (n_22378));
NAND2X1 g114065(.A (n_21619), .B (n_14597), .Y (n_21620));
NAND2X1 g114068(.A (n_21618), .B (n_21617), .Y (n_22376));
NAND2X2 g114074(.A (n_35935), .B (n_34745), .Y (n_21950));
AOI21X1 g114079(.A0 (n_21054), .A1 (n_19845), .B0 (n_21615), .Y(n_21616));
NAND2X1 g114098(.A (n_35500), .B (n_21621), .Y (n_22375));
NAND2X1 g114101(.A (n_25596), .B (n_21621), .Y (n_21614));
AOI21X1 g114104(.A0 (n_20595), .A1 (n_25942), .B0 (n_14792), .Y(n_21613));
INVX1 g114130(.A (n_21611), .Y (n_21612));
NAND2X1 g114139(.A (n_33851), .B (n_32180), .Y (n_22424));
NAND2X1 g114154(.A (n_21118), .B (n_21609), .Y (n_22396));
NAND2X1 g114162(.A (n_20544), .B (n_21607), .Y (n_21608));
AOI21X1 g114165(.A0 (n_21137), .A1 (n_26162), .B0 (n_15134), .Y(n_32093));
AOI21X1 g114166(.A0 (n_21135), .A1 (n_34952), .B0 (n_14790), .Y(n_21605));
NAND2X1 g114173(.A (n_20668), .B (n_21604), .Y (n_22417));
NAND2X1 g114176(.A (n_20663), .B (n_21603), .Y (n_22410));
NAND2X1 g114180(.A (n_20659), .B (n_21602), .Y (n_22402));
NAND2X1 g114202(.A (n_21108), .B (n_21601), .Y (n_22385));
NAND2X1 g114203(.A (n_20660), .B (n_21600), .Y (n_22383));
AOI21X1 g114206(.A0 (n_21139), .A1 (n_34952), .B0 (n_19446), .Y(n_21599));
NAND3X1 g114216(.A (n_21117), .B (n_17516), .C (n_17508), .Y(n_21598));
XOR2X1 g114225(.A (n_16879), .B (n_21560), .Y (n_22407));
XOR2X1 g114230(.A (n_16949), .B (n_34646), .Y (n_22404));
XOR2X1 g114232(.A (n_20605), .B (n_20603), .Y (n_22380));
OAI21X1 g114249(.A0 (n_21588), .A1 (n_19772), .B0 (n_20979), .Y(n_21931));
AOI21X1 g114252(.A0 (n_21595), .A1 (n_32303), .B0 (n_20981), .Y(n_21596));
AOI21X1 g114253(.A0 (n_21142), .A1 (n_34606), .B0 (n_20977), .Y(n_21594));
NOR2X1 g114254(.A (n_21378), .B (n_21101), .Y (n_22344));
NAND2X1 g114259(.A (n_21592), .B (n_20555), .Y (n_21593));
NAND2X1 g114262(.A (n_21590), .B (n_21465), .Y (n_21591));
NAND2X1 g114265(.A (n_21491), .B (n_20925), .Y (n_21589));
AOI21X1 g114271(.A0 (n_34845), .A1 (n_20972), .B0 (n_21073), .Y(n_21927));
NAND2X1 g114273(.A (n_21074), .B (n_21588), .Y (n_21925));
NAND2X1 g114275(.A (n_21072), .B (n_20984), .Y (n_21923));
NAND3X1 g114284(.A (n_10565), .B (n_18755), .C (n_20564), .Y(n_21587));
NAND3X1 g114287(.A (n_17835), .B (n_18727), .C (n_20558), .Y(n_21586));
INVX1 g114289(.A (n_21132), .Y (n_22293));
NAND2X1 g114307(.A (n_21584), .B (n_18340), .Y (n_21585));
NAND2X1 g114314(.A (n_21584), .B (n_24446), .Y (n_21582));
NAND2X1 g114324(.A (n_21584), .B (n_32697), .Y (n_21581));
NAND2X1 g114337(.A (n_21125), .B (n_25290), .Y (n_21580));
NAND2X1 g114343(.A (n_21563), .B (n_24361), .Y (n_21579));
NAND2X1 g114346(.A (n_20631), .B (n_21098), .Y (n_21911));
NAND3X1 g114352(.A (n_21149), .B (n_19971), .C (n_21576), .Y(n_21578));
NAND2X1 g114353(.A (n_21148), .B (n_21576), .Y (n_21577));
NAND3X1 g114357(.A (n_19957), .B (n_20630), .C (n_21574), .Y(n_21575));
NAND2X1 g114360(.A (n_21572), .B (n_21458), .Y (n_21573));
NAND2X1 g114370(.A (n_20591), .B (n_25942), .Y (n_21571));
NAND2X1 g114381(.A (n_19438), .B (n_20647), .Y (n_22365));
NAND2X1 g114382(.A (n_21157), .B (n_21007), .Y (n_21570));
NAND2X1 g114386(.A (n_20597), .B (n_21439), .Y (n_21569));
NAND2X1 g114387(.A (n_21052), .B (n_19900), .Y (n_21568));
NAND2X1 g114391(.A (n_35939), .B (n_19996), .Y (n_21567));
NAND2X1 g114396(.A (n_20593), .B (n_25942), .Y (n_21565));
NAND2X1 g114398(.A (n_21563), .B (n_24348), .Y (n_21564));
NAND2X1 g114411(.A (n_21560), .B (n_18858), .Y (n_21561));
NAND3X1 g114418(.A (n_21047), .B (n_20015), .C (n_17559), .Y(n_21559));
NAND4X1 g114426(.A (n_21886), .B (n_21557), .C (n_20014), .D(n_18851), .Y (n_21558));
NAND3X1 g114432(.A (n_19440), .B (n_21154), .C (n_21555), .Y(n_21556));
AOI21X1 g114464(.A0 (n_19196), .A1 (n_20521), .B0 (n_34678), .Y(n_21554));
NAND2X1 g114465(.A (n_20620), .B (n_18212), .Y (n_21552));
NAND2X1 g114469(.A (n_20645), .B (n_21551), .Y (n_21970));
NAND2X1 g114470(.A (n_20643), .B (n_21551), .Y (n_21985));
NAND2X1 g114476(.A (n_20642), .B (n_21550), .Y (n_21967));
NAND2X1 g114477(.A (n_20640), .B (n_21550), .Y (n_21983));
NAND2X1 g114479(.A (n_20637), .B (n_21549), .Y (n_21959));
NAND2X1 g114480(.A (n_20635), .B (n_21549), .Y (n_21981));
NAND2X1 g114486(.A (n_20633), .B (n_21548), .Y (n_21975));
NAND2X1 g114487(.A (n_20632), .B (n_21548), .Y (n_21956));
NAND3X1 g114499(.A (n_20001), .B (n_19998), .C (n_15143), .Y(n_21547));
NAND3X1 g114503(.A (n_19999), .B (n_19980), .C (n_15140), .Y(n_21546));
AOI21X1 g114505(.A0 (n_20518), .A1 (n_20011), .B0 (n_21511), .Y(n_21876));
OAI21X1 g114519(.A0 (n_35538), .A1 (n_20516), .B0 (n_21545), .Y(n_21962));
INVX1 g114539(.A (n_21625), .Y (n_21544));
NAND2X1 g114557(.A (n_21542), .B (n_21533), .Y (n_21543));
INVX1 g114559(.A (n_21540), .Y (n_21541));
INVX1 g114563(.A (n_21538), .Y (n_21539));
INVX1 g114568(.A (n_21536), .Y (n_21537));
NOR3X1 g114572(.A (n_17231), .B (n_17349), .C (n_19953), .Y(n_22255));
NAND3X1 g114580(.A (n_18708), .B (n_19885), .C (n_18709), .Y(n_21869));
INVX1 g114583(.A (n_21534), .Y (n_35415));
NAND2X1 g114585(.A (n_19982), .B (n_20358), .Y (n_22589));
NAND2X1 g114588(.A (n_19793), .B (n_21533), .Y (n_21867));
NAND2X1 g114592(.A (n_20524), .B (n_20368), .Y (n_21532));
AOI21X1 g114597(.A0 (n_17888), .A1 (n_19309), .B0 (n_20319), .Y(n_21531));
AND2X1 g114599(.A (n_21529), .B (n_21528), .Y (n_21530));
AND2X1 g114616(.A (n_21526), .B (n_17346), .Y (n_21527));
AOI21X1 g114621(.A0 (n_35902), .A1 (n_21059), .B0 (n_21525), .Y(n_21860));
NAND2X1 g114631(.A (n_21523), .B (n_19832), .Y (n_21524));
AND2X1 g114643(.A (n_17289), .B (n_20546), .Y (n_22561));
OR2X1 g114645(.A (n_21144), .B (n_20829), .Y (n_21522));
NOR2X1 g114648(.A (n_20447), .B (n_21521), .Y (n_22906));
INVX1 g114669(.A (n_21080), .Y (n_21944));
NAND2X1 g114673(.A (n_18546), .B (n_21518), .Y (n_21520));
NOR2X1 g114681(.A (n_21036), .B (n_21419), .Y (n_21519));
NAND2X1 g114683(.A (n_35736), .B (n_21518), .Y (n_22263));
NAND2X1 g114687(.A (n_21516), .B (n_27522), .Y (n_21517));
AOI21X1 g114694(.A0 (n_32379), .A1 (n_18059), .B0 (n_20520), .Y(n_21837));
NOR2X1 g114698(.A (n_19217), .B (n_20985), .Y (n_22284));
NAND2X1 g114702(.A (n_20975), .B (n_19277), .Y (n_21515));
AOI21X1 g114707(.A0 (n_20442), .A1 (n_21514), .B0 (n_21513), .Y(n_21835));
NAND2X1 g114716(.A (n_21511), .B (n_20848), .Y (n_21512));
NAND2X1 g114722(.A (n_26584), .B (n_21518), .Y (n_22265));
INVX1 g114741(.A (n_21069), .Y (n_21509));
NAND2X1 g114745(.A (n_20559), .B (n_18808), .Y (n_21821));
NAND3X1 g114748(.A (n_21507), .B (n_21636), .C (n_21506), .Y(n_21508));
NAND2X1 g114752(.A (n_20556), .B (n_18804), .Y (n_21819));
INVX1 g114758(.A (n_21504), .Y (n_21505));
NAND2X1 g114760(.A (n_20554), .B (n_18802), .Y (n_21998));
NAND2X1 g114771(.A (n_20549), .B (n_20349), .Y (n_21816));
NAND2X1 g114775(.A (n_20548), .B (n_19805), .Y (n_21814));
NAND2X1 g114779(.A (n_20547), .B (n_19803), .Y (n_21996));
NAND4X1 g114782(.A (n_21502), .B (n_19822), .C (n_23089), .D(n_21501), .Y (n_21503));
INVX1 g114805(.A (n_21060), .Y (n_21993));
NAND2X1 g114808(.A (n_20539), .B (n_19798), .Y (n_21810));
INVX1 g114811(.A (n_21497), .Y (n_21498));
INVX1 g114823(.A (n_21495), .Y (n_21496));
NAND2X2 g114831(.A (n_20538), .B (n_19807), .Y (n_21992));
NAND4X1 g114832(.A (n_19218), .B (n_20572), .C (n_20571), .D(n_20797), .Y (n_21494));
INVX1 g114833(.A (n_21592), .Y (n_21493));
INVX1 g114842(.A (n_21491), .Y (n_21492));
AOI21X1 g114882(.A0 (n_20990), .A1 (n_14781), .B0 (n_23138), .Y(n_21490));
AOI22X1 g114888(.A0 (n_21488), .A1 (n_20408), .B0 (n_19255), .B1(n_18504), .Y (n_21489));
NAND2X1 g114891(.A (n_19366), .B (n_20589), .Y (n_21487));
NAND2X1 g114898(.A (n_20581), .B (n_18744), .Y (n_21486));
OAI21X1 g114902(.A0 (n_19812), .A1 (n_10790), .B0 (n_18662), .Y(n_21485));
XOR2X1 g114909(.A (n_19735), .B (n_21858), .Y (n_22266));
XOR2X1 g114911(.A (n_18043), .B (n_19335), .Y (n_21797));
NAND2X1 g114914(.A (n_22244), .B (n_20836), .Y (n_21484));
AND2X1 g114922(.A (n_20340), .B (n_21414), .Y (n_22221));
NOR2X1 g114924(.A (n_20495), .B (n_20505), .Y (n_21795));
AND2X1 g114931(.A (n_20359), .B (n_20931), .Y (n_22206));
NAND2X1 g114940(.A (n_20336), .B (n_21482), .Y (n_21483));
NAND2X1 g114942(.A (n_34098), .B (n_21480), .Y (n_32613));
NAND2X1 g114959(.A (n_20802), .B (n_19079), .Y (n_21479));
NOR2X1 g114963(.A (n_20475), .B (n_20958), .Y (n_21478));
NOR2X1 g114972(.A (n_20964), .B (n_21475), .Y (n_21477));
NOR2X1 g114973(.A (n_19761), .B (n_21475), .Y (n_21476));
NAND2X1 g114980(.A (n_33184), .B (n_19694), .Y (n_21471));
NAND2X1 g114996(.A (n_21469), .B (n_28890), .Y (n_21470));
NAND2X1 g114998(.A (n_19323), .B (n_18857), .Y (n_21468));
AND2X1 g114999(.A (n_23029), .B (n_21432), .Y (n_21467));
NAND2X1 g115025(.A (n_21858), .B (n_21856), .Y (n_21466));
NAND2X1 g115029(.A (n_21636), .B (n_21465), .Y (n_21785));
NOR2X1 g115031(.A (n_19917), .B (n_21464), .Y (n_22915));
NAND2X1 g115033(.A (n_21463), .B (n_21462), .Y (n_22514));
AND2X1 g115041(.A (n_21806), .B (n_18113), .Y (n_21461));
NOR2X1 g115042(.A (n_18854), .B (n_20455), .Y (n_21460));
NAND2X1 g115050(.A (n_21459), .B (n_21458), .Y (n_21777));
NAND2X1 g115059(.A (n_21465), .B (n_21773), .Y (n_21457));
NOR2X1 g115060(.A (n_20370), .B (n_10470), .Y (n_21456));
NAND2X1 g115063(.A (n_21180), .B (n_20275), .Y (n_21455));
AND2X1 g115066(.A (n_21462), .B (n_21771), .Y (n_21454));
NOR2X1 g115069(.A (n_20926), .B (n_20444), .Y (n_23028));
NAND2X1 g115070(.A (n_21452), .B (n_19894), .Y (n_21453));
NAND2X1 g115071(.A (n_21450), .B (n_21654), .Y (n_21451));
OR2X1 g115074(.A (n_20339), .B (n_21308), .Y (n_21449));
NOR2X1 g115076(.A (n_20440), .B (n_20455), .Y (n_21448));
NAND2X1 g115079(.A (n_20834), .B (n_20439), .Y (n_21447));
AND2X1 g115080(.A (n_22875), .B (n_20451), .Y (n_22917));
NOR2X1 g115091(.A (n_19789), .B (n_20329), .Y (n_21446));
NOR2X1 g115094(.A (n_20326), .B (n_19778), .Y (n_21445));
NOR2X1 g115108(.A (n_21772), .B (n_34825), .Y (n_21766));
AND2X1 g115111(.A (n_19992), .B (n_21443), .Y (n_21444));
INVX1 g115113(.A (n_21441), .Y (n_21442));
NAND2X1 g115117(.A (n_21440), .B (n_21439), .Y (n_21762));
INVX1 g115119(.A (n_21437), .Y (n_21438));
NAND2X1 g115128(.A (n_20827), .B (n_21432), .Y (n_21433));
NAND2X1 g115134(.A (n_21430), .B (n_20372), .Y (n_21431));
AND2X1 g115135(.A (n_21769), .B (n_21428), .Y (n_21429));
NOR2X1 g115137(.A (n_20456), .B (n_33026), .Y (n_21427));
NOR2X1 g115141(.A (n_21425), .B (n_19922), .Y (n_21426));
NAND2X1 g115142(.A (n_20816), .B (n_20486), .Y (n_22211));
INVX1 g115145(.A (n_21423), .Y (n_21424));
NAND2X1 g115148(.A (n_20425), .B (n_19061), .Y (n_21422));
NAND2X1 g115151(.A (n_21421), .B (n_22552), .Y (n_21754));
NOR2X1 g115155(.A (n_20902), .B (n_21419), .Y (n_32924));
NAND2X1 g115158(.A (n_20823), .B (n_34511), .Y (n_21418));
AND2X1 g115163(.A (n_21414), .B (n_20628), .Y (n_21749));
INVX1 g115166(.A (n_21412), .Y (n_21413));
NAND2X1 g115170(.A (n_21410), .B (n_28890), .Y (n_21411));
INVX1 g115174(.A (n_21408), .Y (n_21409));
INVX1 g115188(.A (n_21853), .Y (n_21407));
NAND2X1 g115198(.A (n_20507), .B (n_18589), .Y (n_21929));
INVX1 g115259(.A (n_21405), .Y (n_21406));
INVX1 g115261(.A (n_21403), .Y (n_21404));
INVX1 g115272(.A (n_20971), .Y (n_22251));
INVX1 g115277(.A (n_21838), .Y (n_21402));
NAND2X1 g115279(.A (n_35114), .B (n_35115), .Y (n_22530));
NAND4X1 g115285(.A (n_18748), .B (n_20969), .C (n_21398), .D(n_19734), .Y (n_21399));
NAND2X1 g115288(.A (n_20515), .B (n_19661), .Y (n_21738));
AOI22X1 g115290(.A0 (n_19688), .A1 (n_21013), .B0 (n_17774), .B1(n_17243), .Y (n_21397));
OAI21X1 g115291(.A0 (n_21395), .A1 (n_16955), .B0 (n_20514), .Y(n_21396));
NAND4X1 g115299(.A (n_21392), .B (n_21393), .C (n_33638), .D(n_33752), .Y (n_21394));
NAND4X1 g115301(.A (n_21390), .B (n_21389), .C (n_21388), .D(n_21387), .Y (n_21391));
OR2X1 g115316(.A (n_20225), .B (n_21385), .Y (n_21386));
INVX1 g115366(.A (n_21383), .Y (n_21384));
INVX1 g115370(.A (n_21381), .Y (n_21382));
AND2X1 g115375(.A (n_21379), .B (n_32364), .Y (n_21380));
NOR2X1 g115378(.A (n_21378), .B (n_20302), .Y (n_21973));
NAND2X1 g115388(.A (n_20253), .B (n_21333), .Y (n_21377));
AOI21X1 g115401(.A0 (n_19632), .A1 (n_25053), .B0 (n_21201), .Y(n_21376));
AOI21X1 g115402(.A0 (n_19630), .A1 (n_25705), .B0 (n_21374), .Y(n_21375));
AOI21X1 g115403(.A0 (n_19627), .A1 (n_25704), .B0 (n_21365), .Y(n_21373));
NAND3X1 g115413(.A (n_20210), .B (n_34612), .C (n_20299), .Y(n_22171));
AOI21X1 g115414(.A0 (n_19625), .A1 (n_28215), .B0 (n_21374), .Y(n_21371));
NAND2X1 g115445(.A (n_20236), .B (n_33803), .Y (n_35135));
NAND2X1 g115465(.A (n_33803), .B (n_20250), .Y (n_21369));
AOI21X1 g115467(.A0 (n_19610), .A1 (n_25713), .B0 (n_21365), .Y(n_21368));
AOI21X1 g115469(.A0 (n_19607), .A1 (n_25690), .B0 (n_21365), .Y(n_21367));
AOI21X1 g115485(.A0 (n_19605), .A1 (n_28205), .B0 (n_21365), .Y(n_21366));
NAND2X1 g115487(.A (n_20263), .B (n_11747), .Y (n_21364));
NOR2X1 g115505(.A (n_18118), .B (n_35216), .Y (n_21363));
NAND2X1 g115507(.A (n_20249), .B (n_21694), .Y (n_21362));
NAND2X1 g115516(.A (n_20238), .B (n_21328), .Y (n_21361));
AOI21X1 g115524(.A0 (n_19598), .A1 (n_25048), .B0 (n_21374), .Y(n_21360));
INVX1 g115526(.A (n_21358), .Y (n_22169));
NAND2X1 g115529(.A (n_21333), .B (n_20248), .Y (n_21357));
NAND4X1 g115533(.A (n_11544), .B (n_19088), .C (n_20224), .D(n_16443), .Y (n_21355));
NAND4X1 g115542(.A (n_11301), .B (n_33976), .C (n_20586), .D(n_19099), .Y (n_22491));
INVX1 g115552(.A (n_21353), .Y (n_21354));
NOR2X1 g115663(.A (n_10021), .B (n_20227), .Y (n_21348));
NAND2X1 g115665(.A (n_21341), .B (n_21328), .Y (n_21347));
AND2X1 g115666(.A (n_21345), .B (n_21344), .Y (n_21346));
NAND2X1 g115667(.A (n_21703), .B (n_21341), .Y (n_21343));
NAND2X1 g115735(.A (n_20239), .B (n_21694), .Y (n_21338));
NAND2X1 g115742(.A (n_21335), .B (n_21328), .Y (n_21337));
NAND2X1 g115743(.A (n_21703), .B (n_21335), .Y (n_21336));
NAND2X1 g115753(.A (n_20240), .B (n_21333), .Y (n_21334));
NOR2X1 g115785(.A (n_10021), .B (n_20756), .Y (n_21332));
NAND2X1 g115788(.A (n_20864), .B (n_21329), .Y (n_21331));
NAND2X1 g115789(.A (n_21329), .B (n_21328), .Y (n_21330));
OR2X1 g115880(.A (n_21326), .B (n_19204), .Y (n_21327));
INVX1 g115893(.A (n_21324), .Y (n_21325));
NAND2X1 g115908(.A (n_13762), .B (n_20234), .Y (n_21322));
INVX1 g115909(.A (n_21320), .Y (n_35273));
INVX1 g115911(.A (n_21318), .Y (n_32108));
NAND3X1 g115925(.A (n_14549), .B (n_14517), .C (n_19634), .Y(n_21315));
NAND3X1 g115930(.A (n_14773), .B (n_14769), .C (n_19620), .Y(n_21314));
AOI21X1 g115935(.A0 (n_11356), .A1 (n_14319), .B0 (n_20233), .Y(n_21313));
INVX1 g115978(.A (n_22578), .Y (n_21312));
INVX1 g115980(.A (n_21310), .Y (n_21311));
OR2X1 g115982(.A (n_21308), .B (n_20247), .Y (n_21309));
INVX1 g115986(.A (n_21306), .Y (n_21307));
INVX1 g115991(.A (n_21304), .Y (n_33016));
NOR2X1 g115993(.A (n_21302), .B (n_20784), .Y (n_21303));
NAND2X1 g115996(.A (n_20317), .B (n_17155), .Y (n_21301));
AND2X1 g116000(.A (n_20262), .B (n_21299), .Y (n_21300));
INVX1 g116005(.A (n_21297), .Y (n_33055));
INVX1 g116009(.A (n_21295), .Y (n_32576));
OAI21X1 g116012(.A0 (n_13761), .A1 (n_21293), .B0 (n_20232), .Y(n_21294));
INVX1 g116046(.A (n_21291), .Y (n_32569));
INVX1 g116151(.A (n_20808), .Y (n_22226));
NAND2X1 g116176(.A (n_19168), .B (n_21326), .Y (n_21290));
AOI21X1 g116183(.A0 (n_18536), .A1 (n_23190), .B0 (n_20271), .Y(n_21289));
AOI22X1 g116185(.A0 (n_23874), .A1 (n_21287), .B0 (n_18402), .B1(n_16548), .Y (n_21288));
AOI22X1 g116190(.A0 (n_19529), .A1 (n_19044), .B0 (n_17155), .B1(n_18320), .Y (n_21286));
NAND2X1 g116226(.A (n_9629), .B (n_20097), .Y (n_35092));
NAND2X1 g116287(.A (n_20304), .B (n_20096), .Y (n_21282));
AOI21X1 g116300(.A0 (n_19522), .A1 (n_25590), .B0 (n_10023), .Y(n_21281));
NAND2X1 g116305(.A (n_9629), .B (n_20095), .Y (n_35094));
AOI21X1 g116310(.A0 (n_19516), .A1 (n_24890), .B0 (n_10023), .Y(n_21279));
NAND2X1 g116323(.A (n_20304), .B (n_20094), .Y (n_21278));
NAND2X1 g116388(.A (n_9629), .B (n_20092), .Y (n_21276));
NAND2X1 g116462(.A (n_9629), .B (n_20101), .Y (n_21274));
NAND2X1 g116481(.A (n_20104), .B (n_22501), .Y (n_21674));
INVX1 g116678(.A (n_21270), .Y (n_21271));
INVX1 g116835(.A (n_21268), .Y (n_21269));
NAND2X1 g116939(.A (n_20197), .B (n_24505), .Y (n_21267));
NAND2X1 g116953(.A (n_20155), .B (n_26929), .Y (n_21266));
NAND2X1 g116954(.A (n_20150), .B (n_28572), .Y (n_21265));
INVX1 g116956(.A (n_20769), .Y (n_21264));
OAI21X1 g116958(.A0 (n_18344), .A1 (n_25694), .B0 (n_21262), .Y(n_21263));
NAND2X1 g116968(.A (n_20148), .B (n_26787), .Y (n_21261));
NAND2X1 g116969(.A (n_20147), .B (n_27709), .Y (n_21260));
INVX1 g116990(.A (n_21258), .Y (n_21259));
NAND2X1 g117006(.A (n_20171), .B (n_27705), .Y (n_21257));
NAND2X1 g117013(.A (n_20202), .B (n_28064), .Y (n_21256));
OAI21X1 g117014(.A0 (n_13317), .A1 (n_18344), .B0 (n_28327), .Y(n_21255));
NAND2X1 g117016(.A (n_20196), .B (n_26925), .Y (n_21254));
NAND2X1 g117017(.A (n_20193), .B (n_28556), .Y (n_21253));
NAND2X1 g117019(.A (n_20182), .B (n_26924), .Y (n_21252));
NAND2X1 g117020(.A (n_20181), .B (n_25151), .Y (n_21251));
NAND2X1 g117022(.A (n_20179), .B (n_28063), .Y (n_21250));
NAND2X1 g117026(.A (n_20170), .B (n_26923), .Y (n_21249));
NAND2X1 g117027(.A (n_20168), .B (n_28551), .Y (n_21248));
NAND2X1 g117030(.A (n_20145), .B (n_28061), .Y (n_21247));
NAND2X1 g117031(.A (n_20144), .B (n_28324), .Y (n_21246));
OAI21X1 g117045(.A0 (n_20235), .A1 (n_13425), .B0 (n_23642), .Y(n_21245));
OAI21X1 g117054(.A0 (n_20235), .A1 (n_21243), .B0 (n_23637), .Y(n_21244));
NAND2X1 g117089(.A (n_20129), .B (n_27525), .Y (n_22110));
AOI21X1 g117090(.A0 (n_20473), .A1 (n_19498), .B0 (n_13745), .Y(n_21242));
AOI21X1 g117092(.A0 (n_33513), .A1 (n_21240), .B0 (n_20174), .Y(n_21241));
OAI21X1 g117094(.A0 (n_10023), .A1 (n_19495), .B0 (n_14518), .Y(n_21239));
AOI21X1 g117095(.A0 (n_20473), .A1 (n_19490), .B0 (n_14160), .Y(n_21237));
AOI21X1 g117104(.A0 (n_34609), .A1 (n_19186), .B0 (n_20139), .Y(n_21235));
INVX1 g117186(.A (n_21233), .Y (n_21234));
NAND2X1 g117189(.A (n_20134), .B (n_13904), .Y (n_21667));
OAI21X1 g117213(.A0 (n_8981), .A1 (n_3157), .B0 (n_20208), .Y(n_21232));
AOI21X1 g117216(.A0 (n_20720), .A1 (n_21328), .B0 (n_13931), .Y(n_21231));
NAND2X1 g117217(.A (n_20203), .B (n_27519), .Y (n_22106));
NAND2X1 g117232(.A (n_20209), .B (n_27521), .Y (n_22103));
AOI21X1 g117242(.A0 (n_20722), .A1 (n_21328), .B0 (n_13915), .Y(n_21230));
NOR2X1 g117244(.A (n_20204), .B (n_13333), .Y (n_21664));
INVX1 g117245(.A (n_21227), .Y (n_21228));
AOI21X1 g117280(.A0 (n_20744), .A1 (n_19108), .B0 (n_9519), .Y(n_21225));
OAI21X1 g117282(.A0 (n_9520), .A1 (n_10110), .B0 (n_20131), .Y(n_21224));
AOI21X1 g117283(.A0 (n_20698), .A1 (n_21328), .B0 (n_14190), .Y(n_21223));
NAND2X1 g117661(.A (n_9629), .B (n_20082), .Y (n_21222));
NAND2X1 g117680(.A (n_9629), .B (n_20081), .Y (n_21221));
NAND2X1 g117683(.A (n_22412), .B (n_21217), .Y (n_21219));
NAND2X1 g117707(.A (n_9629), .B (n_20073), .Y (n_21216));
NAND2X1 g117732(.A (n_20071), .B (n_22139), .Y (n_21215));
NAND2X1 g117734(.A (n_9629), .B (n_20079), .Y (n_21214));
NAND2X1 g117739(.A (n_9629), .B (n_20078), .Y (n_21212));
NAND2X1 g117745(.A (n_22064), .B (n_21217), .Y (n_21211));
NAND2X1 g117760(.A (n_9629), .B (n_20070), .Y (n_21210));
NAND2X1 g117776(.A (n_20068), .B (n_22139), .Y (n_21208));
NAND2X1 g117790(.A (n_32794), .B (n_21217), .Y (n_21207));
NAND2X1 g117833(.A (n_20304), .B (n_20075), .Y (n_21206));
NAND2X1 g117850(.A (n_9629), .B (n_20074), .Y (n_21205));
NAND2X1 g117855(.A (n_21217), .B (n_18375), .Y (n_21204));
NOR2X1 g117876(.A (n_19523), .B (n_13147), .Y (n_21203));
AOI21X1 g117891(.A0 (n_19468), .A1 (n_29034), .B0 (n_21201), .Y(n_21202));
NAND2X1 g118127(.A (n_20069), .B (n_22139), .Y (n_21200));
OAI21X1 g119430(.A0 (n_22042), .A1 (n_16420), .B0 (n_13662), .Y(n_21199));
NAND2X1 g119438(.A (n_20067), .B (n_28554), .Y (n_21197));
AOI22X1 g119698(.A0 (n_20218), .A1 (n_13301), .B0 (n_17639), .B1(n_8946), .Y (n_21196));
NOR2X1 g112039(.A (n_21195), .B (n_20443), .Y (n_21652));
INVX1 g112445(.A (n_22085), .Y (n_22081));
AOI21X1 g112618(.A0 (n_19461), .A1 (n_21603), .B0 (n_8065), .Y(n_21194));
AOI21X1 g112646(.A0 (n_19459), .A1 (n_21602), .B0 (n_26052), .Y(n_21193));
INVX1 g112672(.A (n_21191), .Y (n_21192));
AOI21X1 g112677(.A0 (n_19457), .A1 (n_21609), .B0 (n_8065), .Y(n_21190));
NAND2X1 g113151(.A (n_21187), .B (n_22792), .Y (n_21189));
NAND2X1 g113176(.A (n_21187), .B (n_32739), .Y (n_21188));
NAND2X1 g113190(.A (n_21187), .B (n_21185), .Y (n_21186));
AOI21X1 g113224(.A0 (n_19455), .A1 (n_21940), .B0 (n_8940), .Y(n_21184));
XOR2X1 g113494(.A (n_16836), .B (n_19453), .Y (n_22073));
NAND2X1 g113578(.A (n_21181), .B (n_25207), .Y (n_21183));
NAND2X1 g113612(.A (n_21181), .B (n_22831), .Y (n_21182));
NAND2X1 g113627(.A (n_20048), .B (n_21180), .Y (n_22068));
NAND2X1 g113648(.A (n_21181), .B (n_23457), .Y (n_21179));
NOR2X1 g113659(.A (n_20049), .B (n_21177), .Y (n_21178));
NAND2X1 g113674(.A (n_21181), .B (n_13274), .Y (n_21176));
NAND2X1 g113784(.A (n_20053), .B (n_22016), .Y (n_21174));
NOR2X1 g113785(.A (n_20055), .B (n_14506), .Y (n_21173));
NAND2X1 g113786(.A (n_20052), .B (n_22015), .Y (n_21172));
OAI21X1 g113787(.A0 (n_20040), .A1 (n_32745), .B0 (n_22013), .Y(n_21171));
OAI21X1 g113788(.A0 (n_20040), .A1 (n_21169), .B0 (n_14089), .Y(n_21170));
OAI21X1 g113813(.A0 (n_35532), .A1 (n_20648), .B0 (n_21168), .Y(n_22066));
XOR2X1 g113861(.A (n_17814), .B (n_20683), .Y (n_22058));
NAND2X1 g113924(.A (n_35231), .B (n_21011), .Y (n_21167));
NAND2X1 g113988(.A (n_21164), .B (n_34499), .Y (n_35252));
NAND2X1 g113997(.A (n_21164), .B (n_18384), .Y (n_21165));
NAND2X1 g114018(.A (n_21164), .B (n_24984), .Y (n_21162));
NAND2X1 g114030(.A (n_20649), .B (n_16677), .Y (n_21160));
NAND2X1 g114049(.A (n_24965), .B (n_21158), .Y (n_21159));
NAND2X1 g114064(.A (n_35816), .B (n_21158), .Y (n_22023));
NAND2X1 g114100(.A (n_25877), .B (n_21158), .Y (n_22026));
AOI21X1 g114131(.A0 (n_20646), .A1 (n_21008), .B0 (n_21157), .Y(n_21611));
NAND4X1 g114192(.A (n_19440), .B (n_21154), .C (n_21153), .D(n_21555), .Y (n_21156));
INVX1 g114223(.A (n_22043), .Y (n_21152));
XOR2X1 g114233(.A (n_17027), .B (n_21115), .Y (n_22025));
XOR2X1 g114235(.A (n_17506), .B (n_32970), .Y (n_22033));
INVX1 g114236(.A (n_21639), .Y (n_21151));
AOI21X1 g114260(.A0 (n_19971), .A1 (n_21149), .B0 (n_21148), .Y(n_32325));
NAND2X1 g114261(.A (n_20007), .B (n_20611), .Y (n_23255));
NAND2X1 g114263(.A (n_34645), .B (n_19932), .Y (n_21147));
OR2X1 g114267(.A (n_21145), .B (n_21144), .Y (n_21146));
NAND3X1 g114268(.A (n_16950), .B (n_16898), .C (n_19965), .Y(n_21143));
AOI21X1 g114277(.A0 (n_35217), .A1 (n_20046), .B0 (n_21142), .Y(n_22373));
NAND2X1 g114279(.A (n_21133), .B (n_26162), .Y (n_21141));
NAND2X1 g114281(.A (n_21139), .B (n_28485), .Y (n_21140));
NAND2X1 g114283(.A (n_21137), .B (n_28485), .Y (n_21138));
NAND2X1 g114285(.A (n_21135), .B (n_27335), .Y (n_21136));
NAND2X1 g114288(.A (n_21133), .B (n_28492), .Y (n_21134));
NAND2X1 g114290(.A (n_20592), .B (n_18163), .Y (n_21132));
NAND2X1 g114291(.A (n_21139), .B (n_25424), .Y (n_21131));
NAND2X1 g114292(.A (n_21137), .B (n_29090), .Y (n_21130));
NAND2X1 g114293(.A (n_21135), .B (n_30197), .Y (n_21129));
NAND2X1 g114294(.A (n_21133), .B (n_29090), .Y (n_21128));
NAND2X1 g114299(.A (n_21563), .B (n_24386), .Y (n_21127));
NAND2X1 g114305(.A (n_21125), .B (n_27999), .Y (n_21126));
NAND2X1 g114312(.A (n_21125), .B (n_23007), .Y (n_21124));
NAND2X1 g114315(.A (n_21563), .B (n_26315), .Y (n_21123));
NAND2X1 g114317(.A (n_34646), .B (n_20481), .Y (n_21122));
NAND2X1 g114323(.A (n_21125), .B (n_32739), .Y (n_21121));
NAND2X1 g114328(.A (n_20594), .B (n_25082), .Y (n_21120));
NAND2X1 g114331(.A (n_21061), .B (n_20652), .Y (n_32591));
NAND2X1 g114336(.A (n_20667), .B (n_26866), .Y (n_21118));
NAND3X1 g114358(.A (n_21068), .B (n_18643), .C (n_19436), .Y(n_21117));
NOR3X1 g114366(.A (n_18401), .B (n_18847), .C (n_19425), .Y(n_21607));
NAND2X1 g114378(.A (n_21115), .B (n_17613), .Y (n_21116));
NAND2X1 g114379(.A (n_20602), .B (n_17087), .Y (n_21114));
NAND2X1 g114383(.A (n_21112), .B (n_20574), .Y (n_21113));
NAND2X1 g114390(.A (n_21110), .B (n_35665), .Y (n_21111));
NAND2X1 g114401(.A (n_13957), .B (n_21109), .Y (n_21619));
NAND2X1 g114419(.A (n_35519), .B (n_21109), .Y (n_21618));
NAND2X1 g114421(.A (n_25596), .B (n_21109), .Y (n_21108));
AOI21X1 g114461(.A0 (n_18820), .A1 (n_20614), .B0 (n_17060), .Y(n_21107));
AOI22X1 g114463(.A0 (n_20467), .A1 (n_21105), .B0 (n_18114), .B1(n_18164), .Y (n_21106));
AOI22X1 g114496(.A0 (n_20511), .A1 (n_21103), .B0 (n_18150), .B1(n_18159), .Y (n_21104));
INVX1 g114537(.A (n_21164), .Y (n_21102));
XOR2X1 g114540(.A (n_16075), .B (n_19391), .Y (n_21625));
XOR2X1 g114545(.A (n_17556), .B (n_19400), .Y (n_21621));
OR2X1 g114555(.A (n_21100), .B (n_21038), .Y (n_21101));
AOI21X1 g114560(.A0 (n_19339), .A1 (n_18853), .B0 (n_18885), .Y(n_21540));
INVX1 g114561(.A (n_21098), .Y (n_21099));
NAND2X1 g114564(.A (n_19989), .B (n_19338), .Y (n_21538));
NAND2X1 g114569(.A (n_19986), .B (n_21097), .Y (n_21536));
INVX1 g114574(.A (n_21095), .Y (n_21096));
AOI21X1 g114584(.A0 (n_19365), .A1 (n_19818), .B0 (n_34111), .Y(n_21534));
NOR2X1 g114589(.A (n_10003), .B (n_19978), .Y (n_21094));
NAND2X1 g114606(.A (n_21090), .B (n_21092), .Y (n_21093));
NAND2X1 g114613(.A (n_21090), .B (n_26315), .Y (n_21091));
AOI21X1 g114624(.A0 (n_10901), .A1 (n_20582), .B0 (n_14198), .Y(n_21089));
NAND2X1 g114630(.A (n_21090), .B (n_22994), .Y (n_21088));
AND2X1 g114633(.A (n_21084), .B (n_17411), .Y (n_21087));
AND2X1 g114634(.A (n_21084), .B (n_9788), .Y (n_21085));
NOR2X1 g114637(.A (n_20517), .B (n_10517), .Y (n_21083));
AND2X1 g114639(.A (n_21082), .B (n_19271), .Y (n_21913));
NAND2X1 g114649(.A (n_21090), .B (n_23329), .Y (n_21081));
NAND3X1 g114668(.A (n_17075), .B (n_19342), .C (n_17076), .Y(n_21901));
NAND2X1 g114670(.A (n_19983), .B (n_18826), .Y (n_21080));
NAND2X1 g114674(.A (n_24965), .B (n_21075), .Y (n_21899));
NOR2X1 g114680(.A (n_20565), .B (n_19611), .Y (n_21079));
NOR2X1 g114686(.A (n_17413), .B (n_21082), .Y (n_21078));
NAND2X1 g114688(.A (n_35744), .B (n_21075), .Y (n_21076));
NAND2X1 g114699(.A (n_21073), .B (n_20509), .Y (n_21074));
NAND2X1 g114701(.A (n_19973), .B (n_19931), .Y (n_21072));
NAND2X1 g114705(.A (n_19960), .B (n_18659), .Y (n_21071));
NAND2X1 g114719(.A (n_35457), .B (n_21075), .Y (n_21914));
NAND2X1 g114725(.A (n_25596), .B (n_21075), .Y (n_21070));
AOI22X1 g114742(.A0 (n_19378), .A1 (n_18888), .B0 (n_18620), .B1(n_21068), .Y (n_21069));
NAND2X1 g114759(.A (n_19428), .B (n_20352), .Y (n_21504));
INVX1 g114766(.A (n_21066), .Y (n_21067));
NAND2X1 g114776(.A (n_19902), .B (n_21084), .Y (n_21065));
AOI21X1 g114784(.A0 (n_19802), .A1 (n_19892), .B0 (n_21016), .Y(n_21907));
INVX1 g114798(.A (n_21063), .Y (n_21064));
INVX1 g114803(.A (n_21061), .Y (n_21062));
NAND2X1 g114806(.A (n_19990), .B (n_18795), .Y (n_21060));
NAND2X2 g114812(.A (n_19417), .B (n_19796), .Y (n_21497));
AOI21X1 g114824(.A0 (n_19795), .A1 (n_18670), .B0 (n_21003), .Y(n_21495));
NAND2X1 g114828(.A (n_19415), .B (n_19801), .Y (n_21615));
NAND2X2 g114834(.A (n_19991), .B (n_19811), .Y (n_21592));
INVX1 g114838(.A (n_33777), .Y (n_21058));
OAI21X1 g114843(.A0 (n_21056), .A1 (n_20465), .B0 (n_19813), .Y(n_21491));
NAND2X2 g114846(.A (n_19976), .B (n_19959), .Y (n_21905));
OAI21X1 g114847(.A0 (n_18169), .A1 (n_19923), .B0 (n_21056), .Y(n_21590));
INVX1 g114861(.A (n_21054), .Y (n_32590));
INVX1 g114866(.A (n_21052), .Y (n_21053));
AOI21X1 g114879(.A0 (n_18798), .A1 (n_20542), .B0 (n_18098), .Y(n_21051));
NAND2X1 g114892(.A (n_19995), .B (n_14995), .Y (n_21050));
AOI22X1 g114893(.A0 (n_18162), .A1 (n_21048), .B0 (n_21047), .B1(n_16641), .Y (n_21049));
NAND2X1 g114897(.A (n_20006), .B (n_18761), .Y (n_21046));
NAND2X1 g114899(.A (n_20003), .B (n_18728), .Y (n_21045));
OAI21X1 g114903(.A0 (n_19324), .A1 (n_8319), .B0 (n_18714), .Y(n_21044));
XOR2X1 g114905(.A (n_16518), .B (n_20527), .Y (n_21584));
NAND2X1 g114915(.A (n_22244), .B (n_21025), .Y (n_21043));
NOR2X1 g114930(.A (n_19780), .B (n_18435), .Y (n_21849));
NAND2X1 g114943(.A (n_19814), .B (n_19746), .Y (n_21042));
NOR2X1 g114944(.A (n_21040), .B (n_20458), .Y (n_21041));
OR2X1 g114960(.A (n_21038), .B (n_18520), .Y (n_21039));
INVX1 g114966(.A (n_21036), .Y (n_21037));
NOR2X1 g114971(.A (n_20960), .B (n_21033), .Y (n_21034));
AND2X1 g114974(.A (n_21031), .B (n_21030), .Y (n_21032));
NAND2X1 g114975(.A (n_14555), .B (n_20987), .Y (n_21029));
AND2X1 g114977(.A (n_21379), .B (n_21027), .Y (n_32095));
NAND2X1 g114994(.A (n_21025), .B (n_28431), .Y (n_21026));
INVX1 g115022(.A (n_21023), .Y (n_21024));
NAND2X1 g115034(.A (n_18821), .B (n_32947), .Y (n_21022));
AND2X1 g115035(.A (n_19906), .B (n_21020), .Y (n_21021));
NAND2X1 g115037(.A (n_35718), .B (n_20461), .Y (n_21019));
NOR2X1 g115040(.A (n_12337), .B (n_32175), .Y (n_21832));
NAND3X1 g115056(.A (n_11772), .B (n_19072), .C (n_19105), .Y(n_22238));
NAND2X1 g115075(.A (n_21513), .B (n_20441), .Y (n_21018));
NAND2X1 g115077(.A (n_21016), .B (n_19893), .Y (n_21017));
AND2X1 g115086(.A (n_19785), .B (n_20513), .Y (n_21015));
AND2X1 g115088(.A (n_19815), .B (n_21013), .Y (n_21014));
NOR2X1 g115095(.A (n_20438), .B (n_22509), .Y (n_21012));
NAND2X1 g115114(.A (n_21011), .B (n_21010), .Y (n_21441));
NAND2X1 g115115(.A (n_19817), .B (n_19377), .Y (n_21009));
NAND2X1 g115120(.A (n_21008), .B (n_21007), .Y (n_21437));
NOR2X1 g115123(.A (n_19846), .B (n_19922), .Y (n_21006));
NOR2X1 g115131(.A (n_20482), .B (n_20483), .Y (n_21005));
NAND2X1 g115138(.A (n_21003), .B (n_19219), .Y (n_21004));
NOR2X1 g115139(.A (n_19944), .B (n_35397), .Y (n_21002));
NOR2X1 g115143(.A (n_20422), .B (n_19385), .Y (n_21001));
NAND2X1 g115144(.A (n_20357), .B (n_19875), .Y (n_21000));
NAND2X1 g115146(.A (n_20419), .B (n_20573), .Y (n_21423));
NAND2X1 g115149(.A (n_34828), .B (n_20998), .Y (n_20999));
NAND2X1 g115152(.A (n_19787), .B (n_17756), .Y (n_32589));
NOR2X1 g115156(.A (n_34283), .B (n_20995), .Y (n_20996));
NAND2X1 g115161(.A (n_33912), .B (n_20350), .Y (n_20992));
NAND2X1 g115164(.A (n_19389), .B (n_20990), .Y (n_21829));
NOR2X1 g115165(.A (n_34067), .B (n_20456), .Y (n_20989));
NAND2X1 g115167(.A (n_34282), .B (n_20988), .Y (n_21412));
NAND2X1 g115171(.A (n_20987), .B (n_13510), .Y (n_21826));
NAND2X1 g115175(.A (n_23521), .B (n_35411), .Y (n_21408));
INVX1 g115184(.A (n_20985), .Y (n_20986));
NAND2X1 g115189(.A (n_19916), .B (n_18806), .Y (n_21853));
NAND2X1 g115193(.A (n_19844), .B (n_19422), .Y (n_21846));
INVX1 g115199(.A (n_20983), .Y (n_20984));
INVX1 g115201(.A (n_20981), .Y (n_20982));
INVX1 g115239(.A (n_20979), .Y (n_20980));
INVX1 g115241(.A (n_20977), .Y (n_20978));
INVX1 g115249(.A (n_20975), .Y (n_20976));
AOI21X1 g115255(.A0 (n_18006), .A1 (n_18011), .B0 (n_19895), .Y(n_20974));
INVX1 g115257(.A (n_20972), .Y (n_20973));
AOI21X1 g115260(.A0 (n_19115), .A1 (n_17880), .B0 (n_20967), .Y(n_21405));
NAND2X1 g115262(.A (n_19952), .B (n_19130), .Y (n_21403));
NAND2X1 g115263(.A (n_19387), .B (n_19660), .Y (n_22871));
NAND2X1 g115266(.A (n_19951), .B (n_19116), .Y (n_22250));
NAND2X1 g115273(.A (n_19950), .B (n_19132), .Y (n_20971));
NAND2X1 g115278(.A (n_19837), .B (n_19410), .Y (n_21838));
OAI21X1 g115310(.A0 (n_20969), .A1 (n_21149), .B0 (n_19830), .Y(n_21862));
NAND2X1 g115328(.A (n_20967), .B (n_19763), .Y (n_20968));
NAND2X1 g115334(.A (n_18572), .B (n_18631), .Y (n_20966));
INVX1 g115341(.A (n_20964), .Y (n_20965));
NAND2X1 g115347(.A (n_20226), .B (n_21328), .Y (n_20962));
NOR2X1 g115355(.A (n_19750), .B (n_20312), .Y (n_20961));
INVX1 g115363(.A (n_20958), .Y (n_20959));
NAND2X2 g115367(.A (n_34725), .B (n_20957), .Y (n_21383));
NAND2X1 g115368(.A (n_19662), .B (n_34723), .Y (n_20956));
NAND2X1 g115371(.A (n_35179), .B (n_20955), .Y (n_21381));
NAND2X1 g115373(.A (n_19684), .B (n_20490), .Y (n_20954));
AOI21X1 g115400(.A0 (n_19086), .A1 (n_25353), .B0 (n_21374), .Y(n_20953));
INVX1 g115404(.A (n_20950), .Y (n_20951));
INVX1 g115407(.A (n_21425), .Y (n_20948));
AND2X1 g115428(.A (n_20946), .B (n_19277), .Y (n_20947));
NAND2X1 g115429(.A (n_20854), .B (n_21328), .Y (n_20945));
NAND2X1 g115437(.A (n_19680), .B (n_21328), .Y (n_20944));
NAND2X1 g115442(.A (n_19683), .B (n_33803), .Y (n_35127));
AOI21X1 g115448(.A0 (n_19082), .A1 (n_24006), .B0 (n_21374), .Y(n_20940));
AOI21X1 g115464(.A0 (n_19081), .A1 (n_25350), .B0 (n_21365), .Y(n_20937));
NOR2X1 g115486(.A (n_10020), .B (n_19686), .Y (n_20935));
NAND2X1 g115489(.A (n_21703), .B (n_20914), .Y (n_20934));
NAND2X1 g115494(.A (n_19678), .B (n_21328), .Y (n_20933));
NAND2X1 g115525(.A (n_21333), .B (n_19682), .Y (n_20932));
NOR2X1 g115527(.A (n_17065), .B (n_18713), .Y (n_21358));
NAND3X1 g115530(.A (n_19670), .B (n_11773), .C (n_20931), .Y(n_21783));
AOI21X1 g115535(.A0 (n_19074), .A1 (n_24011), .B0 (n_21374), .Y(n_20930));
NAND3X1 g115536(.A (n_19667), .B (n_11774), .C (n_20928), .Y(n_20929));
INVX1 g115539(.A (n_21464), .Y (n_20927));
INVX1 g115549(.A (n_20926), .Y (n_21781));
INVX1 g115554(.A (n_20925), .Y (n_21353));
INVX1 g115569(.A (n_21458), .Y (n_20924));
NAND2X1 g115577(.A (n_20112), .B (n_20889), .Y (n_20923));
INVX1 g115581(.A (n_21776), .Y (n_20922));
INVX1 g115605(.A (n_20919), .Y (n_21349));
INVX1 g115609(.A (n_20917), .Y (n_23393));
INVX1 g115610(.A (n_20917), .Y (n_20918));
NOR2X1 g115614(.A (n_18642), .B (n_20916), .Y (n_23523));
NAND2X1 g115637(.A (n_20914), .B (n_21328), .Y (n_20915));
INVX1 g115644(.A (n_20912), .Y (n_20913));
NAND2X1 g115656(.A (n_20906), .B (n_21328), .Y (n_20909));
NAND2X1 g115657(.A (n_21703), .B (n_20906), .Y (n_20908));
AND2X1 g115668(.A (n_20904), .B (n_20404), .Y (n_32151));
INVX1 g115687(.A (n_20902), .Y (n_21917));
NAND2X1 g115696(.A (n_19676), .B (n_21328), .Y (n_20901));
INVX1 g115700(.A (n_21419), .Y (n_33008));
NOR2X1 g115703(.A (n_20355), .B (n_19280), .Y (n_20899));
NOR2X1 g115708(.A (n_20818), .B (n_19191), .Y (n_20898));
NAND2X1 g115715(.A (n_21703), .B (n_20876), .Y (n_20895));
NAND2X1 g115720(.A (n_19681), .B (n_21658), .Y (n_20894));
NAND2X1 g115721(.A (n_20891), .B (n_21328), .Y (n_20893));
NAND2X1 g115722(.A (n_21703), .B (n_20891), .Y (n_20892));
NAND2X1 g115728(.A (n_20889), .B (n_20887), .Y (n_20890));
NAND2X1 g115733(.A (n_20884), .B (n_20887), .Y (n_20888));
NAND2X1 g115734(.A (n_21703), .B (n_20884), .Y (n_20886));
NAND2X1 g115736(.A (n_20880), .B (n_20887), .Y (n_20883));
NAND2X1 g115737(.A (n_20112), .B (n_20880), .Y (n_20882));
NAND2X1 g115740(.A (n_20851), .B (n_21328), .Y (n_20879));
NAND2X1 g115741(.A (n_20876), .B (n_21328), .Y (n_20877));
NOR2X1 g115744(.A (n_20872), .B (n_25540), .Y (n_20875));
NOR2X1 g115745(.A (n_10021), .B (n_20872), .Y (n_20874));
NAND2X1 g115757(.A (n_20867), .B (n_21328), .Y (n_20871));
NAND2X1 g115771(.A (n_21703), .B (n_20867), .Y (n_20868));
NAND2X1 g115775(.A (n_20864), .B (n_20228), .Y (n_20866));
NAND2X1 g115779(.A (n_20864), .B (n_20862), .Y (n_20865));
NAND2X1 g115780(.A (n_20862), .B (n_21328), .Y (n_20863));
NAND2X1 g115781(.A (n_20864), .B (n_20230), .Y (n_20861));
NAND2X1 g115815(.A (n_20864), .B (n_20857), .Y (n_20859));
NAND2X1 g115816(.A (n_20857), .B (n_21328), .Y (n_20858));
NAND2X1 g115821(.A (n_19674), .B (n_21328), .Y (n_20856));
NAND2X1 g115828(.A (n_21703), .B (n_20854), .Y (n_20855));
NOR2X1 g115830(.A (n_10021), .B (n_20237), .Y (n_20853));
NAND2X1 g115839(.A (n_20864), .B (n_20851), .Y (n_20852));
NAND2X1 g115864(.A (n_23230), .B (n_19049), .Y (n_20850));
NOR2X1 g115871(.A (n_19777), .B (n_19629), .Y (n_21779));
OR2X1 g115872(.A (n_19776), .B (n_20830), .Y (n_21764));
NAND2X1 g115895(.A (n_20848), .B (n_19200), .Y (n_21324));
NOR2X1 g115897(.A (n_35354), .B (n_32365), .Y (n_20847));
INVX1 g115898(.A (n_20844), .Y (n_20845));
AND2X1 g115900(.A (n_34745), .B (n_35353), .Y (n_20843));
NAND2X1 g115910(.A (n_19759), .B (n_20098), .Y (n_21320));
OAI21X1 g115912(.A0 (n_35707), .A1 (n_18319), .B0 (n_19531), .Y(n_21318));
INVX1 g115917(.A (n_21475), .Y (n_20840));
AND2X1 g115920(.A (n_20839), .B (n_20838), .Y (n_21744));
INVX1 g115922(.A (n_20836), .Y (n_20837));
INVX1 g115973(.A (n_20834), .Y (n_20835));
AND2X1 g115976(.A (n_20832), .B (n_20831), .Y (n_20833));
NOR2X1 g115979(.A (n_19728), .B (n_20830), .Y (n_22578));
OR2X1 g115981(.A (n_20829), .B (n_19726), .Y (n_21310));
INVX1 g115984(.A (n_20827), .Y (n_35639));
INVX1 g115987(.A (n_20362), .Y (n_21306));
INVX1 g115989(.A (n_20825), .Y (n_20826));
NAND2X1 g115992(.A (n_19725), .B (n_19027), .Y (n_21304));
INVX1 g116003(.A (n_20823), .Y (n_32097));
OAI21X1 g116006(.A0 (n_20822), .A1 (n_17257), .B0 (n_19042), .Y(n_21297));
OAI21X1 g116010(.A0 (n_20819), .A1 (n_18352), .B0 (n_20818), .Y(n_21295));
OAI21X1 g116047(.A0 (n_18468), .A1 (n_20354), .B0 (n_19723), .Y(n_21291));
INVX1 g116048(.A (n_20816), .Y (n_20817));
INVX1 g116081(.A (n_20814), .Y (n_20815));
INVX1 g116090(.A (n_20812), .Y (n_20813));
INVX1 g116092(.A (n_20346), .Y (n_21813));
OAI21X1 g116141(.A0 (n_20270), .A1 (n_19208), .B0 (n_19827), .Y(n_20809));
NAND2X1 g116152(.A (n_19704), .B (n_18969), .Y (n_20808));
AOI21X1 g116153(.A0 (n_20341), .A1 (n_20338), .B0 (n_20246), .Y(n_21789));
AND2X1 g116156(.A (n_19696), .B (n_21308), .Y (n_20805));
OAI21X1 g116162(.A0 (n_19045), .A1 (n_19073), .B0 (n_17787), .Y(n_20804));
INVX1 g116180(.A (n_20802), .Y (n_20803));
NAND3X1 g116217(.A (n_20102), .B (n_18989), .C (n_20103), .Y(n_22500));
NAND2X1 g116275(.A (n_20797), .B (n_20796), .Y (n_20798));
NAND2X1 g116278(.A (n_18981), .B (n_19583), .Y (n_20795));
NAND2X1 g116301(.A (n_9629), .B (n_19540), .Y (n_20794));
NAND2X1 g116336(.A (n_9629), .B (n_19538), .Y (n_20792));
NAND2X1 g116337(.A (n_9629), .B (n_19537), .Y (n_20791));
NAND2X1 g116419(.A (n_9629), .B (n_19534), .Y (n_20790));
NAND2X1 g116421(.A (n_9629), .B (n_19546), .Y (n_20788));
INVX1 g116569(.A (n_22143), .Y (n_20787));
INVX1 g116638(.A (n_20784), .Y (n_21272));
INVX1 g116642(.A (n_22512), .Y (n_20783));
NAND2X1 g116679(.A (n_20315), .B (n_21758), .Y (n_21270));
NAND2X1 g116766(.A (n_9629), .B (n_19532), .Y (n_20782));
NAND2X1 g116836(.A (n_22177), .B (n_20781), .Y (n_21268));
INVX1 g116914(.A (n_20777), .Y (n_20778));
INVX1 g116917(.A (n_20775), .Y (n_20776));
INVX1 g116922(.A (n_20773), .Y (n_20774));
NAND2X1 g116933(.A (n_19641), .B (n_26869), .Y (n_21692));
AOI21X1 g116934(.A0 (n_20830), .A1 (n_22831), .B0 (n_13655), .Y(n_20772));
NAND2X1 g116942(.A (n_19576), .B (n_25681), .Y (n_20771));
NOR2X1 g116946(.A (n_19606), .B (n_14182), .Y (n_20770));
AOI21X1 g116957(.A0 (n_33556), .A1 (n_23192), .B0 (n_13464), .Y(n_20769));
NAND2X1 g116959(.A (n_19601), .B (n_17390), .Y (n_21717));
NAND2X1 g116964(.A (n_19596), .B (n_25684), .Y (n_20767));
NAND2X1 g116966(.A (n_19593), .B (n_25683), .Y (n_20766));
NAND2X1 g116972(.A (n_19575), .B (n_28202), .Y (n_20765));
NAND2X1 g116976(.A (n_19689), .B (n_20342), .Y (n_20764));
OR2X1 g116991(.A (n_19601), .B (n_20763), .Y (n_21258));
NAND2X1 g117003(.A (n_19578), .B (n_25682), .Y (n_20762));
NAND2X1 g117004(.A (n_19573), .B (n_25679), .Y (n_20761));
NAND2X1 g117005(.A (n_19619), .B (n_28196), .Y (n_20760));
OAI21X1 g117028(.A0 (n_8678), .A1 (n_14097), .B0 (n_19613), .Y(n_20759));
NAND2X1 g117076(.A (n_19643), .B (n_26776), .Y (n_21727));
NAND2X1 g117086(.A (n_19569), .B (n_28543), .Y (n_21702));
INVX1 g117137(.A (n_20756), .Y (n_20757));
NAND2X1 g117140(.A (n_19649), .B (n_26774), .Y (n_21698));
NAND2X1 g117180(.A (n_19650), .B (n_26854), .Y (n_21705));
NAND2X1 g117187(.A (n_19570), .B (n_20755), .Y (n_21233));
OAI21X1 g117210(.A0 (n_9520), .A1 (n_9313), .B0 (n_19645), .Y(n_20754));
NAND2X1 g117231(.A (n_19646), .B (n_28538), .Y (n_21682));
NAND2X1 g117246(.A (n_19639), .B (n_28532), .Y (n_21227));
AOI22X1 g117276(.A0 (n_20218), .A1 (n_10885), .B0 (n_33556), .B1(n_8946), .Y (n_20752));
AOI22X1 g117277(.A0 (n_10573), .A1 (n_13169), .B0 (n_20175), .B1(n_8946), .Y (n_20750));
AOI22X1 g117279(.A0 (n_16798), .A1 (n_8946), .B0 (n_20218), .B1(n_10880), .Y (n_20749));
OAI21X1 g117281(.A0 (n_9520), .A1 (n_10112), .B0 (n_19567), .Y(n_20748));
AOI22X1 g117291(.A0 (n_20188), .A1 (n_8946), .B0 (n_10573), .B1(n_7819), .Y (n_20747));
NAND2X1 g117595(.A (n_18546), .B (n_20744), .Y (n_20746));
NOR2X1 g117695(.A (n_19520), .B (n_20741), .Y (n_20743));
AOI21X1 g117781(.A0 (n_18911), .A1 (n_27220), .B0 (n_10023), .Y(n_20740));
OR2X1 g117789(.A (n_10023), .B (n_19500), .Y (n_20739));
OR2X1 g117835(.A (n_21374), .B (n_19504), .Y (n_20737));
NAND2X1 g117837(.A (n_9629), .B (n_19503), .Y (n_20736));
NAND2X1 g118189(.A (n_19491), .B (n_22139), .Y (n_20734));
NAND2X1 g118256(.A (n_19489), .B (n_21694), .Y (n_20733));
NAND2X1 g118277(.A (n_27747), .B (n_19000), .Y (n_20732));
NAND2X1 g118291(.A (n_20133), .B (n_20744), .Y (n_20730));
NAND2X1 g118295(.A (n_35473), .B (n_20744), .Y (n_20729));
NOR2X1 g118298(.A (n_20727), .B (n_19483), .Y (n_20728));
NAND2X1 g118299(.A (n_21703), .B (n_20717), .Y (n_20726));
NOR2X1 g118300(.A (n_20727), .B (n_19479), .Y (n_20725));
NOR2X1 g118301(.A (n_10020), .B (n_19477), .Y (n_20724));
NAND2X1 g118303(.A (n_20864), .B (n_20722), .Y (n_20723));
NAND2X1 g118304(.A (n_20864), .B (n_20720), .Y (n_20721));
NAND2X1 g118305(.A (n_21703), .B (n_19481), .Y (n_20719));
NAND2X1 g118311(.A (n_20717), .B (n_21328), .Y (n_20718));
NAND2X1 g118317(.A (n_20112), .B (n_20714), .Y (n_20716));
NAND2X1 g118318(.A (n_20714), .B (n_21328), .Y (n_20715));
NAND2X1 g118319(.A (n_20112), .B (n_20711), .Y (n_20713));
NAND2X1 g118320(.A (n_20711), .B (n_21328), .Y (n_20712));
NAND2X1 g118328(.A (n_20864), .B (n_20703), .Y (n_20710));
NAND2X1 g118329(.A (n_20864), .B (n_20706), .Y (n_20708));
NAND2X1 g118330(.A (n_20706), .B (n_21328), .Y (n_20707));
NAND2X1 g118331(.A (n_20703), .B (n_21328), .Y (n_20704));
NAND2X1 g118379(.A (n_20864), .B (n_20700), .Y (n_20702));
NAND2X1 g118380(.A (n_20700), .B (n_21328), .Y (n_20701));
NAND2X1 g118381(.A (n_20112), .B (n_20698), .Y (n_20699));
AOI21X1 g118586(.A0 (n_18289), .A1 (n_8467), .B0 (n_19513), .Y(n_20697));
OAI21X1 g119550(.A0 (n_13781), .A1 (n_16173), .B0 (n_13493), .Y(n_20695));
OAI21X1 g119559(.A0 (n_13990), .A1 (n_16173), .B0 (n_14117), .Y(n_20694));
NAND2X1 g119572(.A (n_19467), .B (n_29014), .Y (n_20692));
AOI22X1 g119683(.A0 (n_18289), .A1 (n_8447), .B0 (n_20741), .B1(n_18909), .Y (n_32226));
XOR2X1 g112446(.A (n_18511), .B (n_20063), .Y (n_22085));
INVX1 g112673(.A (n_21195), .Y (n_21191));
NOR2X1 g113134(.A (n_20060), .B (n_20054), .Y (n_20690));
AOI21X1 g113317(.A0 (n_14993), .A1 (n_20688), .B0 (n_19460), .Y(n_20689));
OAI21X1 g113825(.A0 (n_19451), .A1 (n_19330), .B0 (n_21941), .Y(n_20687));
NAND2X1 g113827(.A (n_19456), .B (n_21939), .Y (n_20685));
XOR2X1 g113886(.A (n_17418), .B (n_18898), .Y (n_21648));
NAND2X1 g114000(.A (n_20681), .B (n_25003), .Y (n_20684));
NOR2X1 g114008(.A (n_20683), .B (n_19768), .Y (n_22039));
NAND2X1 g114011(.A (n_20681), .B (n_32794), .Y (n_20682));
NAND2X1 g114020(.A (n_20681), .B (n_23696), .Y (n_20679));
XOR2X1 g114224(.A (n_18997), .B (n_19440), .Y (n_22043));
XOR2X1 g114238(.A (n_16837), .B (n_20042), .Y (n_21639));
NAND2X1 g114251(.A (n_24563), .B (n_20671), .Y (n_20676));
NAND2X1 g114255(.A (n_24563), .B (n_20665), .Y (n_20675));
NAND2X1 g114256(.A (n_24563), .B (n_20661), .Y (n_20674));
NAND2X1 g114258(.A (n_24563), .B (n_20657), .Y (n_20673));
NAND2X2 g114278(.A (n_20029), .B (n_33772), .Y (n_22008));
NAND2X1 g114297(.A (n_20671), .B (n_25756), .Y (n_20672));
NAND2X1 g114298(.A (n_20671), .B (n_34753), .Y (n_20670));
NAND2X1 g114303(.A (n_20599), .B (n_19381), .Y (n_32180));
NAND2X1 g114306(.A (n_20667), .B (n_22412), .Y (n_20668));
NAND2X1 g114308(.A (n_20665), .B (n_25756), .Y (n_20666));
NAND2X1 g114309(.A (n_20665), .B (n_34753), .Y (n_20664));
NAND2X1 g114313(.A (n_20667), .B (n_23270), .Y (n_20663));
NAND2X1 g114319(.A (n_20661), .B (n_28798), .Y (n_20662));
NAND2X1 g114320(.A (n_35790), .B (n_21109), .Y (n_20660));
NAND2X1 g114322(.A (n_20667), .B (n_32728), .Y (n_20659));
NAND2X1 g114329(.A (n_20657), .B (n_25756), .Y (n_20658));
NAND2X1 g114330(.A (n_20657), .B (n_24526), .Y (n_20656));
NAND2X1 g114333(.A (n_32971), .B (n_18830), .Y (n_20655));
NAND3X1 g114392(.A (n_20033), .B (n_18870), .C (n_20652), .Y(n_32125));
OAI21X1 g114417(.A0 (n_19335), .A1 (n_18883), .B0 (n_16684), .Y(n_20651));
AOI21X1 g114438(.A0 (n_14986), .A1 (n_23176), .B0 (n_19443), .Y(n_20650));
NAND2X1 g114460(.A (n_19442), .B (n_19447), .Y (n_35231));
AOI21X1 g114524(.A0 (n_18862), .A1 (n_18179), .B0 (n_17553), .Y(n_20649));
XOR2X1 g114538(.A (n_18602), .B (n_20035), .Y (n_21164));
INVX1 g114541(.A (n_20648), .Y (n_21158));
AOI21X1 g114562(.A0 (n_19314), .A1 (n_18646), .B0 (n_20612), .Y(n_21098));
NAND2X1 g114565(.A (n_18886), .B (n_19825), .Y (n_21572));
AOI21X1 g114575(.A0 (n_33774), .A1 (n_35716), .B0 (n_18873), .Y(n_21095));
NAND2X2 g114586(.A (n_19408), .B (n_34551), .Y (n_21560));
INVX1 g114602(.A (n_20646), .Y (n_20647));
NAND2X1 g114611(.A (n_20641), .B (n_23725), .Y (n_20645));
NAND2X1 g114612(.A (n_20639), .B (n_22414), .Y (n_20643));
NAND2X1 g114617(.A (n_20641), .B (n_22406), .Y (n_20642));
NAND2X1 g114618(.A (n_20639), .B (n_22406), .Y (n_20640));
AOI21X1 g114619(.A0 (n_10124), .A1 (n_20004), .B0 (n_15142), .Y(n_20638));
NAND2X1 g114625(.A (n_20641), .B (n_32664), .Y (n_20637));
NAND2X1 g114626(.A (n_20639), .B (n_32685), .Y (n_20635));
NAND2X1 g114635(.A (n_20639), .B (n_26866), .Y (n_20633));
NAND2X1 g114636(.A (n_20641), .B (n_26866), .Y (n_20632));
NAND2X1 g114640(.A (n_20630), .B (n_18824), .Y (n_20631));
AND2X1 g114641(.A (n_21105), .B (n_20628), .Y (n_20629));
NAND2X1 g114656(.A (n_27100), .B (n_20625), .Y (n_20627));
NAND2X1 g114658(.A (n_8990), .B (n_20625), .Y (n_20626));
NAND3X1 g114661(.A (n_19437), .B (n_21008), .C (n_33705), .Y(n_20624));
AND2X1 g114664(.A (n_21103), .B (n_20621), .Y (n_20622));
NAND2X1 g114685(.A (n_20619), .B (n_29505), .Y (n_20620));
NAND2X1 g114690(.A (n_27100), .B (n_19977), .Y (n_20618));
NAND3X1 g114704(.A (n_19974), .B (n_19975), .C (n_18659), .Y(n_20616));
AND2X1 g114709(.A (n_20614), .B (n_18884), .Y (n_20615));
AOI21X1 g114713(.A0 (n_20612), .A1 (n_19368), .B0 (n_19988), .Y(n_20613));
INVX1 g114749(.A (n_20610), .Y (n_20611));
INVX1 g114753(.A (n_20607), .Y (n_20609));
NAND2X1 g114765(.A (n_19427), .B (n_19321), .Y (n_21148));
NAND2X1 g114767(.A (n_19426), .B (n_20028), .Y (n_21066));
NAND4X1 g114783(.A (n_20605), .B (n_18181), .C (n_19958), .D(n_18604), .Y (n_20606));
NAND2X1 g114797(.A (n_19421), .B (n_29505), .Y (n_20604));
NAND2X1 g114799(.A (n_19420), .B (n_17083), .Y (n_21063));
NAND2X1 g114804(.A (n_19419), .B (n_35356), .Y (n_21061));
INVX1 g114826(.A (n_20602), .Y (n_20603));
NAND2X1 g114829(.A (n_19412), .B (n_29505), .Y (n_20601));
INVX1 g114835(.A (n_20599), .Y (n_20600));
NAND2X1 g114848(.A (n_19404), .B (n_18812), .Y (n_21157));
NAND2X1 g114850(.A (n_19434), .B (n_20022), .Y (n_21139));
NAND2X1 g114855(.A (n_19433), .B (n_20021), .Y (n_21137));
NAND2X1 g114856(.A (n_19431), .B (n_20020), .Y (n_21135));
INVX1 g114857(.A (n_20661), .Y (n_20598));
NAND2X1 g114860(.A (n_19429), .B (n_20019), .Y (n_21133));
NAND2X1 g114862(.A (n_19406), .B (n_18811), .Y (n_21054));
INVX1 g114864(.A (n_20596), .Y (n_20597));
NAND2X1 g114867(.A (n_19435), .B (n_19319), .Y (n_21052));
OAI21X1 g114873(.A0 (n_18786), .A1 (n_19330), .B0 (n_21890), .Y(n_20595));
NAND2X1 g114874(.A (n_19430), .B (n_21889), .Y (n_20594));
OAI21X1 g114875(.A0 (n_18786), .A1 (n_24312), .B0 (n_21892), .Y(n_20593));
AOI21X1 g114876(.A0 (n_18439), .A1 (n_19987), .B0 (n_18230), .Y(n_20592));
NAND2X1 g114877(.A (n_19424), .B (n_21885), .Y (n_20591));
XOR2X1 g114906(.A (n_18614), .B (n_32378), .Y (n_21125));
XOR2X1 g114908(.A (n_21507), .B (n_18621), .Y (n_21563));
OAI21X1 g114916(.A0 (n_18737), .A1 (n_18792), .B0 (n_21020), .Y(n_21529));
NAND2X1 g114918(.A (n_18438), .B (n_20540), .Y (n_20589));
NAND2X1 g114925(.A (n_26756), .B (n_20563), .Y (n_20588));
NAND3X1 g114926(.A (n_33976), .B (n_18751), .C (n_20586), .Y(n_21533));
NAND2X1 g114945(.A (n_20579), .B (n_25988), .Y (n_20584));
NAND2X1 g114948(.A (n_20582), .B (n_25988), .Y (n_20583));
NAND2X1 g114949(.A (n_20577), .B (n_34709), .Y (n_20581));
NAND2X1 g114951(.A (n_26978), .B (n_20579), .Y (n_20580));
NAND2X1 g114953(.A (n_26978), .B (n_20577), .Y (n_20578));
NOR2X1 g114954(.A (n_8682), .B (n_19326), .Y (n_20576));
NAND2X1 g114956(.A (n_26978), .B (n_20530), .Y (n_20575));
NAND2X1 g114968(.A (n_20574), .B (n_20573), .Y (n_21036));
AND2X1 g114969(.A (n_20572), .B (n_20571), .Y (n_21872));
NAND2X1 g114981(.A (n_20579), .B (n_26870), .Y (n_20570));
AND2X1 g114982(.A (n_19380), .B (n_20017), .Y (n_20569));
NAND2X1 g114985(.A (n_20567), .B (n_34753), .Y (n_20568));
INVX1 g114986(.A (n_20565), .Y (n_20566));
NAND2X1 g114990(.A (n_20563), .B (n_34753), .Y (n_20564));
AND2X1 g114991(.A (n_23053), .B (n_9730), .Y (n_20562));
NAND2X1 g114993(.A (n_21823), .B (n_18586), .Y (n_21526));
NAND2X1 g114995(.A (n_20577), .B (n_26870), .Y (n_20561));
NAND2X1 g114997(.A (n_19810), .B (n_19373), .Y (n_20559));
NAND2X1 g115001(.A (n_20557), .B (n_10808), .Y (n_20558));
NAND2X1 g115002(.A (n_19322), .B (n_18124), .Y (n_20556));
NAND2X1 g115006(.A (n_35869), .B (n_35870), .Y (n_21523));
NOR2X1 g115010(.A (n_19374), .B (n_19913), .Y (n_20555));
NAND2X1 g115012(.A (n_19808), .B (n_18856), .Y (n_20554));
NAND2X1 g115016(.A (n_20552), .B (n_21576), .Y (n_32302));
NOR2X1 g115019(.A (n_19369), .B (n_19912), .Y (n_20551));
NAND2X1 g115023(.A (n_20550), .B (n_20574), .Y (n_21023));
NAND2X1 g115027(.A (n_18801), .B (n_20462), .Y (n_20549));
NAND2X1 g115032(.A (n_18800), .B (n_20464), .Y (n_20548));
NAND2X1 g115043(.A (n_19804), .B (n_19264), .Y (n_20547));
NAND3X1 g115045(.A (n_11782), .B (n_17907), .C (n_18563), .Y(n_21886));
NOR2X1 g115047(.A (n_20009), .B (n_19272), .Y (n_20546));
OR2X1 g115057(.A (n_20041), .B (n_20545), .Y (n_21144));
OR2X1 g115065(.A (n_19332), .B (n_20446), .Y (n_20544));
AND2X1 g115067(.A (n_20542), .B (n_20541), .Y (n_20543));
NAND2X1 g115073(.A (n_17778), .B (n_20540), .Y (n_22220));
NAND2X1 g115118(.A (n_19800), .B (n_19934), .Y (n_20539));
NAND2X1 g115124(.A (n_19797), .B (n_19937), .Y (n_20538));
NAND2X1 g115130(.A (n_19806), .B (n_20485), .Y (n_20537));
NOR2X1 g115133(.A (n_19926), .B (n_19878), .Y (n_32320));
NAND2X1 g115140(.A (n_21525), .B (n_33853), .Y (n_20535));
NAND3X1 g115168(.A (n_19948), .B (n_34845), .C (n_20532), .Y(n_35126));
NAND2X1 g115169(.A (n_20530), .B (n_26870), .Y (n_20531));
NAND2X1 g115178(.A (n_20528), .B (n_26106), .Y (n_20529));
NAND2X1 g115185(.A (n_20527), .B (n_17882), .Y (n_20985));
NAND2X1 g115200(.A (n_19347), .B (n_18032), .Y (n_20983));
NAND2X1 g115202(.A (n_19384), .B (n_19146), .Y (n_20981));
NAND2X1 g115237(.A (n_19343), .B (n_19142), .Y (n_21142));
AOI21X1 g115240(.A0 (n_19767), .A1 (n_19962), .B0 (n_20431), .Y(n_20979));
NAND2X1 g115242(.A (n_19382), .B (n_19133), .Y (n_20977));
INVX1 g115244(.A (n_19964), .Y (n_21588));
NAND2X1 g115250(.A (n_19353), .B (n_19963), .Y (n_20975));
INVX1 g115251(.A (n_20525), .Y (n_32303));
NAND2X1 g115258(.A (n_19356), .B (n_18026), .Y (n_20972));
INVX1 g115269(.A (n_20523), .Y (n_20524));
INVX1 g115275(.A (n_20521), .Y (n_20522));
NAND2X1 g115280(.A (n_19355), .B (n_18036), .Y (n_20520));
INVX1 g115283(.A (n_20518), .Y (n_20519));
NAND2X1 g115286(.A (n_18829), .B (n_19127), .Y (n_21511));
INVX1 g115294(.A (n_20517), .Y (n_21516));
INVX1 g115311(.A (n_20516), .Y (n_21518));
AND2X1 g115315(.A (n_19218), .B (n_20797), .Y (n_22257));
NAND2X1 g115323(.A (n_19659), .B (n_34724), .Y (n_20515));
OAI21X1 g115326(.A0 (n_16584), .A1 (n_16512), .B0 (n_20513), .Y(n_20514));
NAND2X1 g115340(.A (n_20511), .B (n_20510), .Y (n_20512));
NAND2X1 g115343(.A (n_20509), .B (n_20500), .Y (n_20964));
AND2X1 g115346(.A (n_20012), .B (n_20011), .Y (n_20508));
NAND2X1 g115349(.A (n_19143), .B (n_19306), .Y (n_20507));
NOR2X1 g115350(.A (n_18757), .B (n_19771), .Y (n_32601));
OR2X1 g115351(.A (n_18900), .B (n_20061), .Y (n_20505));
NAND2X1 g115357(.A (n_19161), .B (n_20478), .Y (n_20504));
NOR2X1 g115358(.A (n_34445), .B (n_18628), .Y (n_20503));
NOR2X1 g115359(.A (n_34601), .B (n_35216), .Y (n_20502));
NAND2X1 g115361(.A (n_20510), .B (n_20621), .Y (n_20501));
NAND2X1 g115364(.A (n_19300), .B (n_20500), .Y (n_20958));
AND2X1 g115365(.A (n_20499), .B (n_19724), .Y (n_23218));
NAND2X1 g115372(.A (n_19134), .B (n_19047), .Y (n_35115));
INVX1 g115379(.A (n_21033), .Y (n_20497));
NOR2X1 g115387(.A (n_20056), .B (n_20495), .Y (n_20496));
NOR2X1 g115389(.A (n_19297), .B (n_19091), .Y (n_22857));
NOR2X1 g115390(.A (n_20493), .B (n_34997), .Y (n_20494));
NAND2X1 g115393(.A (n_20389), .B (n_21328), .Y (n_20492));
NAND2X1 g115394(.A (n_19184), .B (n_20490), .Y (n_20491));
AND2X1 g115395(.A (n_34441), .B (n_20488), .Y (n_32304));
NAND2X1 g115405(.A (n_19178), .B (n_20487), .Y (n_20950));
NAND2X1 g115408(.A (n_20486), .B (n_20485), .Y (n_21425));
NAND2X1 g115417(.A (n_19182), .B (n_22139), .Y (n_20484));
INVX1 g115418(.A (n_20483), .Y (n_21421));
INVX1 g115425(.A (n_20482), .Y (n_21439));
INVX1 g115434(.A (n_20480), .Y (n_20481));
NAND2X1 g115438(.A (n_19160), .B (n_20478), .Y (n_20479));
NAND2X1 g115451(.A (n_19180), .B (n_22139), .Y (n_20477));
INVX1 g115461(.A (n_21857), .Y (n_20938));
NOR2X1 g115463(.A (n_19285), .B (n_17581), .Y (n_21856));
INVX1 g115481(.A (n_20475), .Y (n_20476));
NAND2X1 g115488(.A (n_19177), .B (n_20473), .Y (n_20474));
NAND2X1 g115492(.A (n_19156), .B (n_21328), .Y (n_20472));
NAND2X1 g115493(.A (n_19175), .B (n_21694), .Y (n_20471));
NAND2X1 g115508(.A (n_20628), .B (n_20469), .Y (n_20470));
NAND2X1 g115509(.A (n_20467), .B (n_20469), .Y (n_20468));
NAND2X1 g115517(.A (n_19158), .B (n_20473), .Y (n_20466));
NOR2X1 g115531(.A (n_20465), .B (n_20459), .Y (n_21465));
NAND2X1 g115540(.A (n_17565), .B (n_20464), .Y (n_21464));
NAND2X1 g115541(.A (n_21333), .B (n_19174), .Y (n_20463));
NAND3X1 g115543(.A (n_19141), .B (n_11300), .C (n_19792), .Y(n_22286));
NOR2X1 g115545(.A (n_17061), .B (n_32949), .Y (n_21462));
NAND2X1 g115550(.A (n_20462), .B (n_20461), .Y (n_20926));
NAND2X1 g115551(.A (n_19267), .B (n_12561), .Y (n_20460));
NOR2X1 g115555(.A (n_20459), .B (n_20458), .Y (n_20925));
NAND2X1 g115559(.A (n_19124), .B (n_19111), .Y (n_21806));
INVX1 g115566(.A (n_20454), .Y (n_20455));
NOR2X1 g115570(.A (n_32949), .B (n_17561), .Y (n_21458));
INVX1 g115574(.A (n_20450), .Y (n_20451));
NAND2X1 g115580(.A (n_18427), .B (n_19742), .Y (n_20448));
NOR2X1 g115582(.A (n_18103), .B (n_18703), .Y (n_21776));
OR2X1 g115583(.A (n_20446), .B (n_19783), .Y (n_20447));
NAND2X1 g115592(.A (n_19173), .B (n_20490), .Y (n_20445));
INVX1 g115593(.A (n_20444), .Y (n_22632));
NOR2X1 g115595(.A (n_20443), .B (n_19743), .Y (n_21450));
NAND2X1 g115597(.A (n_20442), .B (n_20441), .Y (n_20921));
NOR2X1 g115598(.A (n_19703), .B (n_19719), .Y (n_21812));
INVX1 g115601(.A (n_20440), .Y (n_20920));
NAND2X1 g115606(.A (n_20439), .B (n_18732), .Y (n_20919));
INVX1 g115607(.A (n_20438), .Y (n_22875));
NAND2X1 g115611(.A (n_20441), .B (n_19065), .Y (n_20917));
NAND2X1 g115616(.A (n_20436), .B (n_19195), .Y (n_20437));
NAND2X1 g115627(.A (n_20433), .B (n_21328), .Y (n_20435));
NAND2X1 g115628(.A (n_21703), .B (n_20433), .Y (n_20434));
NAND2X1 g115636(.A (n_20360), .B (n_20388), .Y (n_20432));
NAND2X1 g115645(.A (n_21760), .B (n_20431), .Y (n_20912));
NAND3X1 g115655(.A (n_17884), .B (n_11748), .C (n_18407), .Y(n_21443));
NAND2X1 g115669(.A (n_20427), .B (n_21328), .Y (n_20429));
NAND2X1 g115670(.A (n_21703), .B (n_20427), .Y (n_20428));
INVX1 g115681(.A (n_20424), .Y (n_20425));
INVX2 g115684(.A (n_20422), .Y (n_35414));
INVX1 g115688(.A (n_20419), .Y (n_20902));
AND2X1 g115690(.A (n_23659), .B (n_34824), .Y (n_20418));
AND2X1 g115695(.A (n_20998), .B (n_34824), .Y (n_20414));
AND2X1 g115697(.A (n_20412), .B (n_20499), .Y (n_33017));
NAND2X2 g115701(.A (n_20411), .B (n_19230), .Y (n_21419));
NOR2X1 g115702(.A (n_20399), .B (n_19679), .Y (n_20410));
NAND2X1 g115706(.A (n_19157), .B (n_20478), .Y (n_20409));
AND2X1 g115711(.A (n_20407), .B (n_20406), .Y (n_21415));
AND2X1 g115712(.A (n_21480), .B (n_20404), .Y (n_20405));
AND2X1 g115714(.A (n_33912), .B (n_20401), .Y (n_20402));
NOR2X1 g115717(.A (n_20399), .B (n_19675), .Y (n_20400));
NAND3X1 g115719(.A (n_19104), .B (n_13095), .C (n_20261), .Y(n_21414));
NAND2X1 g115726(.A (n_20396), .B (n_20887), .Y (n_20398));
NAND2X1 g115727(.A (n_21703), .B (n_20396), .Y (n_20397));
AND2X1 g115729(.A (n_19890), .B (n_20395), .Y (n_21432));
INVX1 g115750(.A (n_20988), .Y (n_20394));
NAND2X1 g115764(.A (n_19166), .B (n_20478), .Y (n_20393));
NAND2X1 g115767(.A (n_20373), .B (n_20887), .Y (n_20392));
NAND2X1 g115774(.A (n_20864), .B (n_20389), .Y (n_20390));
AND2X1 g115786(.A (n_20361), .B (n_20388), .Y (n_22506));
NAND2X1 g115787(.A (n_19154), .B (n_21328), .Y (n_20387));
NAND2X1 g115790(.A (n_20864), .B (n_20384), .Y (n_20386));
NAND2X1 g115791(.A (n_20384), .B (n_21328), .Y (n_20385));
NAND2X1 g115795(.A (n_19685), .B (n_21328), .Y (n_20383));
NAND2X1 g115812(.A (n_20864), .B (n_19671), .Y (n_20382));
NOR2X1 g115819(.A (n_20399), .B (n_19673), .Y (n_20381));
NOR2X1 g115822(.A (n_10021), .B (n_19152), .Y (n_20380));
NOR2X1 g115825(.A (n_20399), .B (n_19677), .Y (n_20379));
NOR2X1 g115826(.A (n_10021), .B (n_19150), .Y (n_20378));
NAND2X1 g115829(.A (n_21703), .B (n_19663), .Y (n_20377));
NAND2X1 g115831(.A (n_19164), .B (n_20490), .Y (n_20376));
INVX1 g115837(.A (n_20995), .Y (n_20375));
NAND2X1 g115842(.A (n_21703), .B (n_20373), .Y (n_20374));
AND2X1 g115881(.A (n_20388), .B (n_20372), .Y (n_21428));
AND2X1 g115882(.A (n_21482), .B (n_20499), .Y (n_20371));
OAI21X1 g115892(.A0 (n_17251), .A1 (n_16134), .B0 (n_19110), .Y(n_20370));
NOR2X1 g115896(.A (n_19193), .B (n_19702), .Y (n_35119));
NAND2X1 g115899(.A (n_18635), .B (n_20368), .Y (n_20844));
NAND2X2 g115918(.A (n_19048), .B (n_20839), .Y (n_21475));
NOR2X1 g115919(.A (n_34997), .B (n_17739), .Y (n_21472));
NOR2X1 g115921(.A (n_34596), .B (n_34997), .Y (n_20365));
OAI21X1 g115923(.A0 (n_18748), .A1 (n_19330), .B0 (n_19329), .Y(n_20836));
NOR2X1 g115924(.A (n_19693), .B (n_34997), .Y (n_20364));
INVX1 g115928(.A (n_21513), .Y (n_20363));
NAND2X1 g115933(.A (n_19290), .B (n_19210), .Y (n_21542));
NAND2X1 g115939(.A (n_19286), .B (n_19328), .Y (n_21469));
NAND2X1 g115974(.A (n_19248), .B (n_19229), .Y (n_20834));
NAND2X1 g115985(.A (n_19240), .B (n_17845), .Y (n_20827));
AOI21X1 g115988(.A0 (n_19039), .A1 (n_20361), .B0 (n_20360), .Y(n_20362));
NAND2X1 g115990(.A (n_19237), .B (n_34830), .Y (n_20825));
AOI21X1 g115995(.A0 (n_11559), .A1 (n_20781), .B0 (n_19668), .Y(n_20359));
INVX1 g116001(.A (n_20357), .Y (n_20358));
NAND2X1 g116004(.A (n_19231), .B (n_18419), .Y (n_20823));
OAI21X1 g116014(.A0 (n_18748), .A1 (n_13316), .B0 (n_19325), .Y(n_21410));
OAI21X1 g116045(.A0 (n_18470), .A1 (n_18355), .B0 (n_20354), .Y(n_21804));
NAND2X1 g116049(.A (n_19234), .B (n_16598), .Y (n_20816));
INVX1 g116060(.A (n_20350), .Y (n_32240));
INVX1 g116077(.A (n_35717), .Y (n_20349));
NAND2X1 g116082(.A (n_19266), .B (n_19320), .Y (n_20814));
NAND2X1 g116085(.A (n_19263), .B (n_19243), .Y (n_21452));
NAND2X1 g116087(.A (n_19249), .B (n_19304), .Y (n_20347));
NAND2X1 g116091(.A (n_19246), .B (n_19729), .Y (n_20812));
NAND2X1 g116093(.A (n_19241), .B (n_17847), .Y (n_20346));
OAI21X1 g116100(.A0 (n_17843), .A1 (n_17902), .B0 (n_19799), .Y(n_21801));
INVX1 g116124(.A (n_19794), .Y (n_20810));
AOI21X1 g116143(.A0 (n_19077), .A1 (n_18667), .B0 (n_35895), .Y(n_22210));
AND2X1 g116146(.A (n_19192), .B (n_20446), .Y (n_20343));
OAI21X1 g116159(.A0 (n_18638), .A1 (n_19169), .B0 (n_20332), .Y(n_20340));
AOI21X1 g116166(.A0 (n_19505), .A1 (n_20341), .B0 (n_20338), .Y(n_20339));
OAI21X1 g116173(.A0 (n_19687), .A1 (n_20338), .B0 (n_20341), .Y(n_20337));
INVX1 g116174(.A (n_20335), .Y (n_20336));
AOI21X1 g116179(.A0 (n_20332), .A1 (n_19169), .B0 (n_19203), .Y(n_21430));
NAND2X1 g116181(.A (n_19232), .B (n_18426), .Y (n_20802));
NAND4X1 g116186(.A (n_18325), .B (n_17631), .C (n_27451), .D(n_17179), .Y (n_20330));
NAND4X1 g116187(.A (n_20328), .B (n_20327), .C (n_22706), .D(n_18449), .Y (n_20329));
NAND4X1 g116188(.A (n_20325), .B (n_20324), .C (n_20323), .D(n_20322), .Y (n_20326));
INVX1 g116199(.A (n_20318), .Y (n_20319));
NAND2X1 g116210(.A (n_20316), .B (n_20315), .Y (n_20317));
NAND2X1 g116212(.A (n_19035), .B (n_20301), .Y (n_23212));
NAND2X1 g116222(.A (n_9629), .B (n_19026), .Y (n_32085));
INVX2 g116234(.A (n_20312), .Y (n_21595));
INVX1 g116236(.A (n_22258), .Y (n_20311));
INVX1 g116246(.A (n_20960), .Y (n_20307));
NAND2X1 g116254(.A (n_20304), .B (n_19019), .Y (n_20305));
NAND2X1 g116265(.A (n_19544), .B (n_18394), .Y (n_20303));
OR2X1 g116266(.A (n_20301), .B (n_21690), .Y (n_20302));
NOR2X1 g116272(.A (n_20299), .B (n_21690), .Y (n_20300));
AOI21X1 g116274(.A0 (n_18368), .A1 (n_24888), .B0 (n_10023), .Y(n_20298));
AOI21X1 g116288(.A0 (n_18391), .A1 (n_24007), .B0 (n_10023), .Y(n_20297));
NAND2X1 g116294(.A (n_20304), .B (n_19023), .Y (n_20295));
NAND2X1 g116295(.A (n_20304), .B (n_19022), .Y (n_20294));
AOI21X1 g116296(.A0 (n_18390), .A1 (n_23542), .B0 (n_10023), .Y(n_20293));
NAND2X1 g116297(.A (n_20304), .B (n_19021), .Y (n_20292));
INVX1 g116302(.A (n_20290), .Y (n_20291));
NAND2X1 g116304(.A (n_9629), .B (n_19020), .Y (n_32089));
AOI21X1 g116324(.A0 (n_18386), .A1 (n_23242), .B0 (n_10023), .Y(n_20288));
NAND2X1 g116329(.A (n_20304), .B (n_19017), .Y (n_20287));
NAND2X1 g116330(.A (n_20304), .B (n_19016), .Y (n_20286));
NAND2X1 g116331(.A (n_9629), .B (n_19014), .Y (n_20285));
NAND2X1 g116332(.A (n_20304), .B (n_19013), .Y (n_20284));
NAND2X1 g116338(.A (n_20304), .B (n_19012), .Y (n_20283));
NAND2X1 g116399(.A (n_20304), .B (n_19011), .Y (n_20282));
NAND2X1 g116400(.A (n_20304), .B (n_19010), .Y (n_20281));
AOI21X1 g116410(.A0 (n_18380), .A1 (n_24894), .B0 (n_10023), .Y(n_20280));
NAND2X1 g116411(.A (n_20304), .B (n_19036), .Y (n_20279));
NAND2X1 g116422(.A (n_9629), .B (n_19038), .Y (n_20278));
AOI21X1 g116465(.A0 (n_18372), .A1 (n_24012), .B0 (n_10023), .Y(n_20277));
INVX1 g116484(.A (n_20274), .Y (n_20275));
NOR2X1 g116535(.A (n_19666), .B (n_20270), .Y (n_20271));
INVX1 g116567(.A (n_22144), .Y (n_20269));
NAND2X1 g116570(.A (n_19786), .B (n_18668), .Y (n_22143));
INVX1 g116611(.A (n_21736), .Y (n_20268));
INVX1 g116617(.A (n_20267), .Y (n_20785));
NAND2X1 g116634(.A (n_17842), .B (n_22501), .Y (n_21747));
AND2X1 g116639(.A (n_20354), .B (n_18471), .Y (n_20784));
INVX1 g116640(.A (n_22511), .Y (n_20266));
NAND2X1 g116643(.A (n_20265), .B (n_20264), .Y (n_22512));
NOR2X1 g116675(.A (n_19695), .B (n_34998), .Y (n_20263));
NAND3X1 g116694(.A (n_19006), .B (n_11788), .C (n_18517), .Y(n_21759));
NOR2X1 g116709(.A (n_19088), .B (n_20261), .Y (n_20262));
INVX1 g116828(.A (n_20257), .Y (n_20258));
INVX1 g116868(.A (n_20848), .Y (n_20255));
NAND2X1 g116915(.A (n_20341), .B (n_19068), .Y (n_20777));
NAND2X1 g116918(.A (n_20254), .B (n_34995), .Y (n_20775));
NAND2X1 g116920(.A (n_19090), .B (n_24009), .Y (n_20253));
NOR2X1 g116923(.A (n_19587), .B (n_19695), .Y (n_20773));
NAND2X1 g116930(.A (n_19587), .B (n_19183), .Y (n_20251));
NAND2X1 g116944(.A (n_19080), .B (n_25049), .Y (n_20250));
NAND2X1 g116955(.A (n_19076), .B (n_25342), .Y (n_20249));
OAI21X1 g116962(.A0 (n_20235), .A1 (n_25694), .B0 (n_23647), .Y(n_20248));
NAND2X1 g116967(.A (n_19600), .B (n_34386), .Y (n_21326));
INVX1 g116979(.A (n_20246), .Y (n_20247));
INVX1 g116982(.A (n_20244), .Y (n_20245));
NOR2X1 g116985(.A (n_20242), .B (n_20241), .Y (n_20243));
OR2X1 g116994(.A (n_20254), .B (n_19695), .Y (n_21345));
NAND2X1 g117000(.A (n_19058), .B (n_24003), .Y (n_20240));
NAND2X1 g117002(.A (n_19057), .B (n_25336), .Y (n_20239));
INVX1 g117007(.A (n_20237), .Y (n_20238));
OAI21X1 g117049(.A0 (n_20235), .A1 (n_13990), .B0 (n_23640), .Y(n_20236));
NAND2X1 g117075(.A (n_19095), .B (n_26777), .Y (n_21335));
AOI21X1 g117091(.A0 (n_20473), .A1 (n_18304), .B0 (n_13741), .Y(n_20234));
OAI21X1 g117093(.A0 (n_25119), .A1 (n_14172), .B0 (n_19083), .Y(n_20233));
AOI21X1 g117096(.A0 (n_20473), .A1 (n_18296), .B0 (n_14155), .Y(n_20232));
INVX1 g117114(.A (n_20230), .Y (n_20231));
INVX1 g117133(.A (n_20228), .Y (n_20229));
NOR2X1 g117138(.A (n_19102), .B (n_13714), .Y (n_20756));
NAND2X1 g117139(.A (n_19101), .B (n_26775), .Y (n_21329));
INVX1 g117176(.A (n_20226), .Y (n_20227));
NAND2X1 g117178(.A (n_19103), .B (n_26780), .Y (n_21341));
OAI21X1 g117196(.A0 (n_16442), .A1 (n_19790), .B0 (n_20224), .Y(n_20225));
OAI21X1 g117220(.A0 (n_8981), .A1 (n_2553), .B0 (n_19097), .Y(n_20223));
AOI21X1 g117259(.A0 (n_18306), .A1 (n_7988), .B0 (n_9510), .Y(n_20221));
AOI22X1 g117270(.A0 (n_19629), .A1 (n_8946), .B0 (n_20218), .B1(n_7575), .Y (n_20220));
AOI22X1 g117290(.A0 (n_19631), .A1 (n_8946), .B0 (n_10573), .B1(n_7706), .Y (n_20217));
AOI22X1 g117292(.A0 (n_19624), .A1 (n_8946), .B0 (n_10573), .B1(n_11122), .Y (n_20215));
NAND4X1 g117302(.A (n_20212), .B (n_18968), .C (n_17747), .D(n_20211), .Y (n_20213));
AOI21X1 g117326(.A0 (n_11747), .A1 (n_17775), .B0 (n_18509), .Y(n_20210));
NAND2X1 g117594(.A (n_14439), .B (n_33000), .Y (n_20209));
NAND2X1 g117611(.A (n_23190), .B (n_8946), .Y (n_20208));
NAND2X1 g117612(.A (n_20830), .B (n_8946), .Y (n_20207));
NOR2X1 g117639(.A (n_35830), .B (n_18371), .Y (n_20204));
NAND2X1 g117641(.A (n_35790), .B (n_33000), .Y (n_20203));
NAND2X1 g117646(.A (n_24101), .B (n_33556), .Y (n_20202));
INVX1 g117654(.A (n_20200), .Y (n_20201));
NAND2X1 g117672(.A (n_9629), .B (n_18954), .Y (n_20199));
NAND2X1 g117674(.A (n_20304), .B (n_18953), .Y (n_20198));
NAND2X1 g117684(.A (n_20830), .B (n_25207), .Y (n_20197));
NAND2X1 g117686(.A (n_18399), .B (n_20195), .Y (n_20196));
NOR2X1 g117688(.A (n_34998), .B (n_19520), .Y (n_20194));
NAND2X1 g117690(.A (n_18399), .B (n_21344), .Y (n_20193));
NAND2X1 g117718(.A (n_23190), .B (n_21919), .Y (n_20191));
NAND2X1 g117721(.A (n_20188), .B (n_17713), .Y (n_20189));
AOI21X1 g117725(.A0 (n_18276), .A1 (n_28213), .B0 (n_21374), .Y(n_20187));
NAND2X1 g117731(.A (n_21703), .B (n_20185), .Y (n_20186));
NAND2X1 g117736(.A (n_9629), .B (n_18952), .Y (n_20184));
NAND2X1 g117738(.A (n_32209), .B (n_9629), .Y (n_20183));
NAND2X1 g117747(.A (n_15089), .B (n_20195), .Y (n_20182));
NAND2X1 g117748(.A (n_22064), .B (n_21344), .Y (n_20181));
NAND2X1 g117757(.A (n_20178), .B (n_33556), .Y (n_20179));
NAND2X1 g117759(.A (n_21919), .B (n_20175), .Y (n_20177));
AOI21X1 g117767(.A0 (n_18270), .A1 (n_20173), .B0 (n_21374), .Y(n_20174));
OR2X1 g117784(.A (n_10023), .B (n_18950), .Y (n_20172));
NAND2X1 g117788(.A (n_20188), .B (n_19577), .Y (n_20171));
NAND2X1 g117793(.A (n_32685), .B (n_20195), .Y (n_20170));
NAND2X1 g117796(.A (n_32685), .B (n_21344), .Y (n_20168));
NAND2X1 g117813(.A (n_21703), .B (n_20165), .Y (n_20167));
NAND2X1 g117814(.A (n_23190), .B (n_27770), .Y (n_20164));
NAND2X1 g117821(.A (n_20188), .B (n_27770), .Y (n_20163));
NOR2X1 g117827(.A (n_20160), .B (n_25540), .Y (n_20161));
AOI21X1 g117830(.A0 (n_18265), .A1 (n_28204), .B0 (n_21201), .Y(n_20159));
NAND2X1 g117836(.A (n_9629), .B (n_18959), .Y (n_20158));
NAND2X1 g117844(.A (n_20304), .B (n_18956), .Y (n_20157));
NAND2X1 g117851(.A (n_18957), .B (n_20490), .Y (n_20156));
NAND2X1 g117866(.A (n_20195), .B (n_20154), .Y (n_20155));
NAND2X1 g117867(.A (n_18946), .B (n_20490), .Y (n_20153));
NAND2X1 g117869(.A (n_21344), .B (n_10848), .Y (n_20151));
NAND2X1 g117870(.A (n_21344), .B (n_18907), .Y (n_20150));
NAND2X1 g117922(.A (n_23190), .B (n_23578), .Y (n_20149));
NAND2X1 g117946(.A (n_20830), .B (n_13274), .Y (n_20148));
NAND2X1 g117954(.A (n_20188), .B (n_19595), .Y (n_20147));
NAND2X1 g118138(.A (n_18945), .B (n_21694), .Y (n_20146));
NAND2X1 g118166(.A (n_17340), .B (n_33556), .Y (n_20145));
NAND2X1 g118181(.A (n_23578), .B (n_20175), .Y (n_20144));
NOR2X1 g118182(.A (n_18943), .B (n_25540), .Y (n_20143));
NAND2X1 g118209(.A (n_23190), .B (n_23356), .Y (n_20141));
INVX1 g118224(.A (n_20138), .Y (n_20139));
NAND2X1 g118264(.A (n_21703), .B (n_20136), .Y (n_20137));
NAND2X1 g118266(.A (n_18944), .B (n_21658), .Y (n_20135));
NAND2X1 g118294(.A (n_20133), .B (n_33000), .Y (n_20134));
NAND2X1 g118297(.A (n_33000), .B (n_19108), .Y (n_20131));
NOR2X1 g118302(.A (n_10020), .B (n_20122), .Y (n_20130));
NAND2X1 g118307(.A (n_35540), .B (n_33000), .Y (n_20129));
NAND2X1 g118309(.A (n_19482), .B (n_21328), .Y (n_20128));
NOR2X1 g118310(.A (n_19480), .B (n_25540), .Y (n_20127));
NAND2X1 g118312(.A (n_19478), .B (n_21328), .Y (n_20125));
NAND2X1 g118313(.A (n_19476), .B (n_21328), .Y (n_20124));
NOR2X1 g118314(.A (n_20122), .B (n_25540), .Y (n_20123));
NAND2X1 g118315(.A (n_20864), .B (n_20119), .Y (n_20121));
NAND2X1 g118316(.A (n_20119), .B (n_21328), .Y (n_20120));
NAND2X1 g118323(.A (n_20112), .B (n_20116), .Y (n_20118));
NAND2X1 g118324(.A (n_20116), .B (n_21328), .Y (n_20117));
NOR2X1 g118325(.A (n_10021), .B (n_20114), .Y (n_20115));
NAND2X1 g118366(.A (n_20112), .B (n_19484), .Y (n_20113));
NAND2X1 g118373(.A (n_20112), .B (n_20109), .Y (n_20111));
NAND2X1 g118374(.A (n_20109), .B (n_21328), .Y (n_20110));
NAND2X1 g118375(.A (n_20112), .B (n_20106), .Y (n_20108));
NAND2X1 g118376(.A (n_20106), .B (n_21328), .Y (n_20107));
NOR2X1 g118377(.A (n_20727), .B (n_18941), .Y (n_20105));
NAND4X1 g118382(.A (n_17163), .B (n_20103), .C (n_20102), .D(n_11775), .Y (n_20104));
NAND2X1 g118422(.A (n_18964), .B (n_19669), .Y (n_21177));
NAND2X1 g118443(.A (n_18993), .B (n_14049), .Y (n_20101));
INVX1 g118465(.A (n_20098), .Y (n_20099));
OAI21X1 g118494(.A0 (n_17830), .A1 (n_19024), .B0 (n_26209), .Y(n_20097));
NAND2X1 g118497(.A (n_18999), .B (n_23382), .Y (n_20096));
OAI21X1 g118503(.A0 (n_17830), .A1 (n_13843), .B0 (n_24121), .Y(n_20095));
NAND2X1 g118507(.A (n_18998), .B (n_23381), .Y (n_20094));
OAI21X1 g118516(.A0 (n_17830), .A1 (n_32673), .B0 (n_26200), .Y(n_20093));
NAND2X1 g118519(.A (n_18996), .B (n_23380), .Y (n_20092));
NAND2X1 g118524(.A (n_18994), .B (n_26197), .Y (n_20091));
NAND2X1 g118589(.A (n_9515), .B (n_18974), .Y (n_20090));
OAI21X1 g118594(.A0 (n_8325), .A1 (n_2979), .B0 (n_18971), .Y(n_20089));
CLKBUFX1 g118898(.A (n_19520), .Y (n_21217));
INVX1 g119282(.A (n_20087), .Y (n_20088));
INVX1 g119286(.A (n_20085), .Y (n_20086));
INVX1 g119290(.A (n_20083), .Y (n_20084));
NAND2X1 g119425(.A (n_18923), .B (n_13667), .Y (n_20082));
NAND2X1 g119429(.A (n_18922), .B (n_27389), .Y (n_20081));
NAND2X1 g119431(.A (n_18921), .B (n_29133), .Y (n_20080));
NAND2X1 g119433(.A (n_18919), .B (n_13650), .Y (n_20079));
NAND2X1 g119437(.A (n_18916), .B (n_27384), .Y (n_20078));
NAND2X1 g119439(.A (n_18914), .B (n_29132), .Y (n_20077));
OAI21X1 g119444(.A0 (n_17150), .A1 (n_32718), .B0 (n_26570), .Y(n_20076));
NAND2X1 g119445(.A (n_18906), .B (n_26376), .Y (n_20075));
NAND2X1 g119446(.A (n_18908), .B (n_27377), .Y (n_20074));
OAI21X1 g119555(.A0 (n_14279), .A1 (n_23778), .B0 (n_20072), .Y(n_20073));
NAND2X1 g119556(.A (n_18920), .B (n_27717), .Y (n_20071));
OAI21X1 g119558(.A0 (n_18429), .A1 (n_23778), .B0 (n_13622), .Y(n_20070));
NAND2X1 g119565(.A (n_18904), .B (n_27708), .Y (n_20069));
NAND2X1 g119576(.A (n_18912), .B (n_27702), .Y (n_20068));
NAND2X1 g119776(.A (n_18384), .B (n_20741), .Y (n_20067));
NAND2X1 g119795(.A (n_32777), .B (n_20741), .Y (n_20065));
NAND2X1 g119812(.A (n_20741), .B (n_18907), .Y (n_20064));
NAND3X1 g112674(.A (n_20063), .B (n_18897), .C (n_17407), .Y(n_21195));
NOR2X1 g113342(.A (n_18902), .B (n_14311), .Y (n_20062));
NOR2X1 g113530(.A (n_20061), .B (n_19452), .Y (n_22810));
INVX1 g113858(.A (n_20060), .Y (n_21187));
OR2X1 g113976(.A (n_19451), .B (n_13663), .Y (n_20059));
NOR2X1 g113982(.A (n_20057), .B (n_20056), .Y (n_20058));
NOR2X1 g113991(.A (n_20038), .B (n_20054), .Y (n_20055));
NAND2X1 g113990(.A (n_20051), .B (n_14690), .Y (n_20053));
NAND2X1 g113999(.A (n_20051), .B (n_20050), .Y (n_20052));
INVX1 g114111(.A (n_20049), .Y (n_20048));
XOR2X1 g114242(.A (n_16798), .B (n_21145), .Y (n_21181));
AOI21X1 g114257(.A0 (n_34554), .A1 (n_18722), .B0 (n_20046), .Y(n_20047));
NAND3X1 g114310(.A (n_17089), .B (n_20044), .C (n_35665), .Y(n_20045));
AND2X1 g114318(.A (n_20042), .B (n_19955), .Y (n_21972));
OR2X1 g114325(.A (n_21145), .B (n_20041), .Y (n_21161));
NAND2X1 g114413(.A (n_19440), .B (n_18460), .Y (n_20683));
XOR2X1 g114542(.A (n_17038), .B (n_19441), .Y (n_20648));
INVX1 g114546(.A (n_20051), .Y (n_20040));
INVX1 g114549(.A (n_20038), .Y (n_20681));
NAND2X1 g114577(.A (n_18877), .B (n_18187), .Y (n_21110));
NAND2X1 g114603(.A (n_18882), .B (n_18819), .Y (n_20646));
NAND2X1 g114615(.A (n_18864), .B (n_8303), .Y (n_20037));
NAND2X1 g114623(.A (n_20035), .B (n_17029), .Y (n_20036));
NAND2X1 g114666(.A (n_18870), .B (n_20033), .Y (n_20034));
NAND3X1 g114695(.A (n_20018), .B (n_20550), .C (n_20031), .Y(n_20032));
NAND2X2 g114708(.A (n_19390), .B (n_17586), .Y (n_20029));
NAND2X1 g114726(.A (n_18881), .B (n_17619), .Y (n_21115));
OAI21X1 g114750(.A0 (n_20023), .A1 (n_33983), .B0 (n_18791), .Y(n_20610));
OAI21X1 g114755(.A0 (n_20028), .A1 (n_19375), .B0 (n_17599), .Y(n_20607));
AOI21X1 g114761(.A0 (n_18790), .A1 (n_18648), .B0 (n_19316), .Y(n_20027));
NAND2X1 g114768(.A (n_18887), .B (n_18799), .Y (n_21634));
NAND2X1 g114800(.A (n_19399), .B (n_17088), .Y (n_20026));
AOI21X1 g114801(.A0 (n_35357), .A1 (n_17030), .B0 (n_19405), .Y(n_20025));
NAND2X1 g114827(.A (n_18173), .B (n_32123), .Y (n_20602));
NAND2X1 g114836(.A (n_18880), .B (n_18844), .Y (n_20599));
NAND3X1 g114837(.A (n_16899), .B (n_18232), .C (n_35850), .Y(n_20024));
NAND2X1 g114841(.A (n_18889), .B (n_20023), .Y (n_32971));
NAND2X1 g114849(.A (n_18893), .B (n_20022), .Y (n_20671));
NAND2X1 g114854(.A (n_18892), .B (n_20021), .Y (n_20665));
OAI21X1 g114858(.A0 (n_18158), .A1 (n_32698), .B0 (n_20020), .Y(n_20661));
NAND2X1 g114859(.A (n_18890), .B (n_20019), .Y (n_20657));
NAND2X1 g114863(.A (n_18872), .B (n_18788), .Y (n_21112));
AOI21X1 g114865(.A0 (n_18810), .A1 (n_17540), .B0 (n_19414), .Y(n_20596));
XOR2X1 g114907(.A (n_16951), .B (n_18178), .Y (n_20667));
XOR2X1 g114912(.A (n_18180), .B (n_20018), .Y (n_21109));
NAND2X1 g114921(.A (n_18168), .B (n_20017), .Y (n_21084));
NAND2X1 g114927(.A (n_18823), .B (n_19905), .Y (n_20016));
NAND2X1 g114929(.A (n_20014), .B (n_18813), .Y (n_20015));
NAND3X1 g114933(.A (n_20012), .B (n_20011), .C (n_20010), .Y(n_20013));
NOR2X1 g114936(.A (n_20009), .B (n_15943), .Y (n_21082));
OAI21X1 g114937(.A0 (n_18044), .A1 (n_18166), .B0 (n_17516), .Y(n_20008));
NAND2X1 g114941(.A (n_21507), .B (n_21506), .Y (n_20007));
NAND2X1 g114946(.A (n_20000), .B (n_30563), .Y (n_20006));
NAND2X1 g114947(.A (n_20004), .B (n_34694), .Y (n_20005));
NAND2X1 g114950(.A (n_19994), .B (n_27340), .Y (n_20003));
NAND2X1 g114952(.A (n_27743), .B (n_20000), .Y (n_20001));
NAND2X1 g114957(.A (n_27743), .B (n_19979), .Y (n_19999));
NAND2X1 g114984(.A (n_20000), .B (n_34802), .Y (n_19998));
NAND2X1 g114987(.A (n_33778), .B (n_19996), .Y (n_20565));
NAND2X1 g115000(.A (n_19994), .B (n_34802), .Y (n_19995));
NAND2X1 g115004(.A (n_20487), .B (n_19992), .Y (n_19993));
NAND2X1 g115009(.A (n_19312), .B (n_19284), .Y (n_19991));
NAND2X1 g115014(.A (n_19318), .B (n_18849), .Y (n_19990));
NAND2X1 g115020(.A (n_19988), .B (n_19367), .Y (n_19989));
NAND3X1 g115039(.A (n_19987), .B (n_18421), .C (n_17165), .Y(n_22228));
NAND2X1 g115052(.A (n_19336), .B (n_18698), .Y (n_19986));
NOR2X1 g115106(.A (n_19359), .B (n_18842), .Y (n_19984));
NAND2X1 g115109(.A (n_18845), .B (n_18672), .Y (n_19983));
NAND2X1 g115132(.A (n_34111), .B (n_19874), .Y (n_19982));
NAND2X1 g115177(.A (n_19979), .B (n_34802), .Y (n_19980));
INVX1 g115179(.A (n_19977), .Y (n_19978));
NAND2X1 g115183(.A (n_19975), .B (n_19974), .Y (n_19976));
INVX1 g115208(.A (n_19972), .Y (n_19973));
INVX1 g115210(.A (n_19969), .Y (n_19971));
NAND2X1 g115214(.A (n_18793), .B (n_18701), .Y (n_19968));
NAND2X1 g115217(.A (n_17079), .B (n_19966), .Y (n_19967));
NAND3X1 g115238(.A (n_18789), .B (n_16288), .C (n_16663), .Y(n_19965));
NAND2X1 g115243(.A (n_18838), .B (n_19144), .Y (n_21073));
OAI21X1 g115245(.A0 (n_19963), .A1 (n_18774), .B0 (n_18587), .Y(n_19964));
AOI21X1 g115252(.A0 (n_19884), .A1 (n_17881), .B0 (n_19962), .Y(n_20525));
AOI21X1 g115270(.A0 (n_18017), .A1 (n_18046), .B0 (n_18859), .Y(n_20523));
NAND2X1 g115276(.A (n_18836), .B (n_18016), .Y (n_20521));
NAND2X1 g115284(.A (n_18861), .B (n_17498), .Y (n_20518));
INVX1 g115292(.A (n_20619), .Y (n_19961));
NOR2X1 g115295(.A (n_18840), .B (n_13509), .Y (n_20517));
INVX1 g115296(.A (n_19959), .Y (n_19960));
OAI21X1 g115308(.A0 (n_19958), .A1 (n_20033), .B0 (n_18841), .Y(n_21075));
XOR2X1 g115309(.A (n_19957), .B (n_18048), .Y (n_21090));
XOR2X1 g115312(.A (n_17089), .B (n_18072), .Y (n_20516));
NAND2X1 g115314(.A (n_18759), .B (n_19955), .Y (n_21038));
OAI21X1 g115324(.A0 (n_20744), .A1 (n_33000), .B0 (n_18565), .Y(n_32175));
NOR2X1 g115325(.A (n_18042), .B (n_19784), .Y (n_19953));
NAND2X1 g115329(.A (n_35062), .B (n_34742), .Y (n_19952));
NAND2X1 g115330(.A (n_19131), .B (n_17876), .Y (n_19951));
NAND2X1 g115333(.A (n_19129), .B (n_17874), .Y (n_19950));
AND2X1 g115344(.A (n_19948), .B (n_34845), .Y (n_19949));
NAND2X1 g115369(.A (n_18618), .B (n_21694), .Y (n_19947));
NAND2X1 g115377(.A (n_18592), .B (n_20490), .Y (n_19946));
NAND2X2 g115380(.A (n_19945), .B (n_19758), .Y (n_21033));
INVX1 g115381(.A (n_19944), .Y (n_21030));
NAND2X1 g115385(.A (n_18617), .B (n_21694), .Y (n_19943));
AND2X1 g115392(.A (n_19945), .B (n_19942), .Y (n_21027));
AND2X1 g115396(.A (n_21787), .B (n_20488), .Y (n_19941));
AOI21X1 g115399(.A0 (n_17935), .A1 (n_25706), .B0 (n_21374), .Y(n_19940));
NAND2X1 g115410(.A (n_21703), .B (n_19138), .Y (n_19939));
NAND2X1 g115416(.A (n_19838), .B (n_21328), .Y (n_19938));
NAND2X2 g115419(.A (n_19937), .B (n_20485), .Y (n_20483));
NAND2X1 g115421(.A (n_21703), .B (n_19860), .Y (n_19936));
NAND2X1 g115423(.A (n_21703), .B (n_19136), .Y (n_19935));
NAND2X1 g115426(.A (n_19413), .B (n_19934), .Y (n_20482));
NAND2X1 g115433(.A (n_21703), .B (n_19858), .Y (n_19933));
NAND2X1 g115435(.A (n_19932), .B (n_19931), .Y (n_20480));
NAND2X1 g115436(.A (n_18594), .B (n_21328), .Y (n_19930));
NAND2X1 g115441(.A (n_18613), .B (n_33803), .Y (n_35124));
NAND2X1 g115443(.A (n_18591), .B (n_21694), .Y (n_19928));
NAND2X1 g115447(.A (n_18612), .B (n_33803), .Y (n_35122));
INVX1 g115449(.A (n_19926), .Y (n_21010));
NAND2X1 g115458(.A (n_18582), .B (n_21328), .Y (n_19925));
NAND2X1 g115459(.A (n_18611), .B (n_33803), .Y (n_19924));
NOR2X1 g115462(.A (n_18131), .B (n_17582), .Y (n_21857));
NOR2X1 g115468(.A (n_19923), .B (n_18052), .Y (n_21636));
INVX1 g115470(.A (n_19921), .Y (n_19922));
NOR2X1 g115474(.A (n_20399), .B (n_19153), .Y (n_19919));
NAND2X1 g115475(.A (n_18610), .B (n_21694), .Y (n_19918));
INVX1 g115476(.A (n_21870), .Y (n_19917));
NAND3X1 g115478(.A (n_21149), .B (n_16915), .C (n_17365), .Y(n_19916));
NOR2X1 g115479(.A (n_19280), .B (n_19915), .Y (n_22573));
NAND2X1 g115482(.A (n_34845), .B (n_20509), .Y (n_20475));
NOR2X1 g115491(.A (n_16689), .B (n_17571), .Y (n_21463));
INVX1 g115497(.A (n_19913), .Y (n_19914));
INVX1 g115520(.A (n_19912), .Y (n_21574));
NAND2X1 g115523(.A (n_18607), .B (n_21658), .Y (n_19911));
NAND2X1 g115528(.A (n_21333), .B (n_18606), .Y (n_19910));
NAND2X1 g115532(.A (n_21333), .B (n_18605), .Y (n_19909));
NAND3X1 g115544(.A (n_18585), .B (n_11304), .C (n_19905), .Y(n_19906));
NAND3X1 g115547(.A (n_9725), .B (n_16616), .C (n_19903), .Y(n_19904));
NAND2X1 g115548(.A (n_18650), .B (n_11022), .Y (n_19902));
NAND2X1 g115556(.A (n_22340), .B (n_32979), .Y (n_21514));
INVX1 g115561(.A (n_19900), .Y (n_20456));
NOR2X1 g115568(.A (n_19268), .B (n_18703), .Y (n_20454));
NAND2X1 g115572(.A (n_18697), .B (n_18113), .Y (n_19898));
NAND2X1 g115576(.A (n_19897), .B (n_20461), .Y (n_20450));
NOR2X1 g115578(.A (n_19262), .B (n_20458), .Y (n_21773));
NOR2X1 g115586(.A (n_17561), .B (n_17580), .Y (n_21771));
INVX1 g115587(.A (n_20542), .Y (n_19895));
NAND2X1 g115594(.A (n_19897), .B (n_19894), .Y (n_20444));
NAND2X1 g115602(.A (n_19893), .B (n_19892), .Y (n_20440));
NAND2X1 g115608(.A (n_19894), .B (n_19891), .Y (n_20438));
NAND2X1 g115613(.A (n_19893), .B (n_17892), .Y (n_21772));
NAND2X1 g115626(.A (n_19238), .B (n_19890), .Y (n_22509));
NAND2X1 g115629(.A (n_17844), .B (n_19890), .Y (n_19889));
NAND2X1 g115643(.A (n_19886), .B (n_21328), .Y (n_19888));
NAND2X1 g115646(.A (n_20864), .B (n_19886), .Y (n_19887));
NAND2X1 g115658(.A (n_19884), .B (n_20487), .Y (n_19885));
NAND2X1 g115659(.A (n_19881), .B (n_21328), .Y (n_19883));
NAND2X1 g115660(.A (n_20864), .B (n_19881), .Y (n_19882));
NAND2X2 g115661(.A (n_34112), .B (n_19880), .Y (n_21059));
NOR2X1 g115662(.A (n_18846), .B (n_18080), .Y (n_21007));
INVX1 g115671(.A (n_19878), .Y (n_35411));
NOR2X1 g115680(.A (n_19364), .B (n_19873), .Y (n_33027));
NOR2X1 g115682(.A (n_19876), .B (n_19260), .Y (n_20424));
NAND2X2 g115686(.A (n_19875), .B (n_19874), .Y (n_20422));
NOR2X1 g115689(.A (n_19873), .B (n_17228), .Y (n_20419));
NOR2X1 g115698(.A (n_19233), .B (n_17224), .Y (n_22552));
INVX1 g115704(.A (n_20573), .Y (n_19871));
NOR2X1 g115707(.A (n_19191), .B (n_18352), .Y (n_22889));
NAND2X1 g115718(.A (n_21703), .B (n_19856), .Y (n_19870));
NAND2X1 g115724(.A (n_35736), .B (n_19868), .Y (n_20987));
NAND2X1 g115725(.A (n_25877), .B (n_19868), .Y (n_20990));
NAND2X1 g115731(.A (n_19864), .B (n_21328), .Y (n_19867));
NAND2X1 g115732(.A (n_20864), .B (n_19864), .Y (n_19866));
NAND2X1 g115738(.A (n_18590), .B (n_20478), .Y (n_19863));
NAND2X1 g115739(.A (n_19841), .B (n_21328), .Y (n_19862));
NOR2X1 g115751(.A (n_35901), .B (n_18776), .Y (n_20988));
NAND2X1 g115759(.A (n_19860), .B (n_21328), .Y (n_19861));
NAND2X1 g115760(.A (n_19858), .B (n_20887), .Y (n_19859));
NAND2X1 g115763(.A (n_19856), .B (n_20887), .Y (n_19857));
NAND2X1 g115777(.A (n_20864), .B (n_19851), .Y (n_19853));
NAND2X1 g115778(.A (n_19851), .B (n_21328), .Y (n_19852));
NAND2X1 g115782(.A (n_20864), .B (n_19848), .Y (n_19850));
NAND2X1 g115783(.A (n_19848), .B (n_21328), .Y (n_19849));
AOI21X1 g115784(.A0 (n_17915), .A1 (n_25680), .B0 (n_21374), .Y(n_19847));
INVX1 g115796(.A (n_19845), .Y (n_19846));
NAND2X1 g115800(.A (n_17968), .B (n_19868), .Y (n_19844));
NAND2X1 g115802(.A (n_20864), .B (n_19120), .Y (n_19843));
NAND2X1 g115804(.A (n_20864), .B (n_19841), .Y (n_19842));
NAND2X1 g115805(.A (n_20864), .B (n_19147), .Y (n_19840));
NAND2X1 g115809(.A (n_20864), .B (n_19838), .Y (n_19839));
NAND2X1 g115817(.A (n_35479), .B (n_19868), .Y (n_19837));
NAND2X1 g115823(.A (n_19151), .B (n_21328), .Y (n_19836));
NAND2X1 g115827(.A (n_19149), .B (n_21328), .Y (n_19835));
NAND2X1 g115838(.A (n_19060), .B (n_20407), .Y (n_20995));
NAND2X1 g115852(.A (n_18609), .B (n_21328), .Y (n_19834));
NOR2X1 g115859(.A (n_20399), .B (n_19155), .Y (n_19833));
AND2X1 g115868(.A (n_18784), .B (n_16353), .Y (n_21180));
NOR2X1 g115878(.A (n_18045), .B (n_18049), .Y (n_19832));
NAND2X1 g115883(.A (n_21703), .B (n_19122), .Y (n_19831));
NAND2X1 g115904(.A (n_20969), .B (n_21149), .Y (n_19830));
NAND2X2 g115929(.A (n_18779), .B (n_19706), .Y (n_21513));
NAND2X1 g115938(.A (n_18749), .B (n_19327), .Y (n_21025));
AOI21X1 g115954(.A0 (n_19666), .A1 (n_19827), .B0 (n_19665), .Y(n_19828));
NOR2X1 g115971(.A (n_19821), .B (n_19820), .Y (n_19822));
INVX1 g115997(.A (n_19818), .Y (n_19819));
NAND2X1 g116002(.A (n_18753), .B (n_18695), .Y (n_20357));
INVX1 g116016(.A (n_19816), .Y (n_19817));
NAND2X1 g116023(.A (n_17770), .B (n_18562), .Y (n_19815));
INVX1 g116033(.A (n_19813), .Y (n_19814));
NAND2X1 g116035(.A (n_18712), .B (n_18112), .Y (n_21040));
INVX1 g116041(.A (n_20530), .Y (n_19812));
NAND2X1 g116050(.A (n_18653), .B (n_19736), .Y (n_21003));
INVX1 g116051(.A (n_19810), .Y (n_19811));
INVX1 g116056(.A (n_19323), .Y (n_20352));
INVX1 g116058(.A (n_19808), .Y (n_19809));
OAI21X1 g116061(.A0 (n_17374), .A1 (n_19788), .B0 (n_18505), .Y(n_20350));
INVX1 g116073(.A (n_19806), .Y (n_19807));
INVX1 g116079(.A (n_19804), .Y (n_19805));
INVX1 g116083(.A (n_19802), .Y (n_19803));
NAND2X1 g116086(.A (n_18692), .B (n_18677), .Y (n_21016));
INVX1 g116112(.A (n_19800), .Y (n_19801));
INVX1 g116118(.A (n_19797), .Y (n_19798));
INVX1 g116120(.A (n_19795), .Y (n_19796));
NAND2X1 g116125(.A (n_18669), .B (n_19786), .Y (n_19794));
NAND3X1 g116128(.A (n_18739), .B (n_19140), .C (n_19792), .Y(n_19793));
AOI21X1 g116136(.A0 (n_19790), .A1 (n_20332), .B0 (n_19169), .Y(n_19791));
NAND3X1 g116137(.A (n_18616), .B (n_16876), .C (n_18157), .Y(n_19789));
OAI21X1 g116138(.A0 (n_17925), .A1 (n_17222), .B0 (n_19788), .Y(n_21488));
OAI21X1 g116142(.A0 (n_19786), .A1 (n_16774), .B0 (n_35896), .Y(n_19787));
AOI21X1 g116144(.A0 (n_17829), .A1 (n_17828), .B0 (n_19784), .Y(n_19785));
AND2X1 g116145(.A (n_18627), .B (n_19783), .Y (n_20993));
AND2X1 g116161(.A (n_18706), .B (n_19331), .Y (n_19782));
NAND3X1 g116163(.A (n_17590), .B (n_17977), .C (n_11778), .Y(n_19781));
OAI21X1 g116164(.A0 (n_17867), .A1 (n_16855), .B0 (n_17785), .Y(n_19780));
NOR2X1 g116175(.A (n_19075), .B (n_35381), .Y (n_20335));
NAND4X1 g116184(.A (n_17782), .B (n_16795), .C (n_33621), .D(n_16794), .Y (n_19779));
NAND2X1 g116189(.A (n_18603), .B (n_18600), .Y (n_19778));
AOI21X1 g116200(.A0 (n_12986), .A1 (n_17732), .B0 (n_17984), .Y(n_20318));
NAND2X1 g116215(.A (n_17398), .B (n_19774), .Y (n_19777));
NAND2X1 g116216(.A (n_17219), .B (n_19774), .Y (n_19776));
NOR2X1 g116218(.A (n_10021), .B (n_18507), .Y (n_19773));
INVX1 g116224(.A (n_20500), .Y (n_19772));
INVX1 g116227(.A (n_19771), .Y (n_20955));
INVX1 g116230(.A (n_19769), .Y (n_19770));
NOR2X1 g116232(.A (n_18461), .B (n_19768), .Y (n_21154));
NAND2X2 g116235(.A (n_19767), .B (n_19383), .Y (n_20312));
NOR2X1 g116237(.A (n_18516), .B (n_19766), .Y (n_22258));
NAND2X2 g116248(.A (n_19763), .B (n_17824), .Y (n_20960));
NAND3X1 g116253(.A (n_18519), .B (n_17802), .C (n_17147), .Y(n_21378));
NAND2X1 g116263(.A (n_19032), .B (n_19758), .Y (n_19759));
NAND2X1 g116264(.A (n_19008), .B (n_19046), .Y (n_19757));
NAND2X1 g116282(.A (n_9629), .B (n_18432), .Y (n_32137));
AOI21X1 g116293(.A0 (n_17817), .A1 (n_22441), .B0 (n_10023), .Y(n_19755));
NAND2X1 g116303(.A (n_17973), .B (n_17983), .Y (n_20290));
NAND2X1 g116322(.A (n_9629), .B (n_18430), .Y (n_32064));
AOI21X1 g116398(.A0 (n_17801), .A1 (n_24324), .B0 (n_10023), .Y(n_19753));
NAND2X1 g116457(.A (n_9629), .B (n_18442), .Y (n_19748));
INVX1 g116477(.A (n_20459), .Y (n_19746));
NAND2X1 g116485(.A (n_18492), .B (n_17386), .Y (n_20274));
INVX1 g116496(.A (n_19743), .Y (n_19744));
NOR2X1 g116499(.A (n_18440), .B (n_13232), .Y (n_22249));
INVX1 g116532(.A (n_19742), .Y (n_20272));
NAND3X1 g116539(.A (n_35404), .B (n_17132), .C (n_17724), .Y(n_22237));
INVX1 g116543(.A (n_19740), .Y (n_19741));
INVX1 g116559(.A (n_21393), .Y (n_19739));
INVX1 g116563(.A (n_21392), .Y (n_19738));
INVX1 g116565(.A (n_22145), .Y (n_19737));
NAND2X1 g116568(.A (n_19736), .B (n_18652), .Y (n_22144));
INVX1 g116580(.A (n_19734), .Y (n_19735));
NAND2X1 g116595(.A (n_19733), .B (n_18710), .Y (n_20831));
NAND2X1 g116596(.A (n_17903), .B (n_18711), .Y (n_22193));
INVX1 g116598(.A (n_21387), .Y (n_19732));
INVX1 g116602(.A (n_21389), .Y (n_19731));
NOR2X1 g116607(.A (n_20931), .B (n_20928), .Y (n_21654));
NAND2X1 g116612(.A (n_17895), .B (n_18106), .Y (n_21736));
INVX1 g116613(.A (n_21735), .Y (n_19730));
NAND2X1 g116618(.A (n_19729), .B (n_19245), .Y (n_20267));
OR2X1 g116619(.A (n_20931), .B (n_18275), .Y (n_19728));
OR2X1 g116629(.A (n_20931), .B (n_20102), .Y (n_19726));
NAND2X1 g116636(.A (n_19029), .B (n_19724), .Y (n_19725));
NAND2X1 g116641(.A (n_18771), .B (n_19723), .Y (n_22511));
INVX1 g116705(.A (n_19721), .Y (n_19722));
INVX1 g116726(.A (n_19719), .Y (n_19720));
AOI21X1 g116780(.A0 (n_17758), .A1 (n_24305), .B0 (n_10023), .Y(n_19717));
AOI21X1 g116792(.A0 (n_17809), .A1 (n_25335), .B0 (n_10023), .Y(n_19715));
AOI21X1 g116800(.A0 (n_17755), .A1 (n_25260), .B0 (n_10023), .Y(n_19713));
NOR2X1 g116818(.A (n_16978), .B (n_16975), .Y (n_19711));
AND2X1 g116822(.A (n_22340), .B (n_19709), .Y (n_19710));
INVX1 g116823(.A (n_19707), .Y (n_19708));
NAND2X1 g116829(.A (n_19706), .B (n_19827), .Y (n_20257));
NAND2X1 g116840(.A (n_19703), .B (n_16785), .Y (n_19704));
INVX1 g116854(.A (n_19702), .Y (n_20957));
NOR2X1 g116869(.A (n_34743), .B (n_17315), .Y (n_20848));
NOR2X1 g116925(.A (n_19695), .B (n_20342), .Y (n_20838));
NAND2X1 g116926(.A (n_19689), .B (n_19695), .Y (n_19696));
INVX1 g116927(.A (n_19693), .Y (n_19694));
INVX1 g116931(.A (n_19690), .Y (n_19691));
NAND2X1 g116975(.A (n_20254), .B (n_19689), .Y (n_21308));
INVX1 g116977(.A (n_19171), .Y (n_19688));
AND2X1 g116980(.A (n_19687), .B (n_20341), .Y (n_20246));
NOR2X1 g116983(.A (n_18497), .B (n_19169), .Y (n_20244));
NOR2X1 g117008(.A (n_18531), .B (n_13940), .Y (n_20237));
INVX1 g117010(.A (n_19685), .Y (n_19686));
NAND2X1 g117043(.A (n_18512), .B (n_22760), .Y (n_19684));
NAND2X1 g117047(.A (n_18499), .B (n_22844), .Y (n_19683));
NAND2X1 g117051(.A (n_18495), .B (n_22759), .Y (n_19682));
NAND2X1 g117053(.A (n_18464), .B (n_22842), .Y (n_19681));
INVX1 g117056(.A (n_19679), .Y (n_19680));
INVX1 g117058(.A (n_19677), .Y (n_19678));
NOR2X1 g117066(.A (n_18527), .B (n_14154), .Y (n_20872));
INVX1 g117067(.A (n_19675), .Y (n_19676));
NAND2X1 g117069(.A (n_18526), .B (n_24751), .Y (n_20867));
NAND2X1 g117071(.A (n_18524), .B (n_24760), .Y (n_20889));
NAND2X1 g117072(.A (n_18530), .B (n_25327), .Y (n_20880));
NAND2X1 g117074(.A (n_18534), .B (n_25839), .Y (n_20851));
NAND2X1 g117077(.A (n_18529), .B (n_25387), .Y (n_20884));
INVX1 g117078(.A (n_19673), .Y (n_19674));
NAND2X1 g117084(.A (n_18523), .B (n_25842), .Y (n_20854));
NAND2X1 g117115(.A (n_18557), .B (n_25329), .Y (n_20230));
INVX1 g117120(.A (n_19671), .Y (n_19672));
NAND2X2 g117123(.A (n_35176), .B (n_17774), .Y (n_23230));
NAND2X1 g117132(.A (n_18545), .B (n_24764), .Y (n_20857));
NAND2X1 g117134(.A (n_18559), .B (n_24785), .Y (n_20228));
NAND2X1 g117136(.A (n_18550), .B (n_25400), .Y (n_20862));
AOI21X1 g117149(.A0 (n_11559), .A1 (n_19669), .B0 (n_19668), .Y(n_19670));
AOI21X1 g117150(.A0 (n_19666), .A1 (n_16808), .B0 (n_19665), .Y(n_19667));
NAND2X1 g117170(.A (n_18543), .B (n_24717), .Y (n_20891));
NAND2X1 g117171(.A (n_18547), .B (n_25396), .Y (n_20906));
NAND2X1 g117173(.A (n_18553), .B (n_24718), .Y (n_20914));
NAND2X1 g117175(.A (n_18542), .B (n_25331), .Y (n_20876));
NAND2X1 g117177(.A (n_18554), .B (n_25846), .Y (n_20226));
INVX1 g117182(.A (n_19663), .Y (n_19664));
INVX1 g117197(.A (n_19661), .Y (n_19662));
NAND2X1 g117199(.A (n_18455), .B (n_16497), .Y (n_20967));
INVX1 g117200(.A (n_19659), .Y (n_19660));
AOI21X1 g117241(.A0 (n_17975), .A1 (n_7988), .B0 (n_9521), .Y(n_19658));
AOI22X1 g117289(.A0 (n_19085), .A1 (n_8946), .B0 (n_20218), .B1(n_7730), .Y (n_19654));
NAND4X1 g117308(.A (n_35041), .B (n_18362), .C (n_19652), .D(n_19651), .Y (n_19653));
NAND2X1 g117452(.A (n_14439), .B (n_19647), .Y (n_19650));
NAND2X1 g117466(.A (n_35790), .B (n_19647), .Y (n_19649));
INVX1 g117577(.A (n_19703), .Y (n_22177));
NAND2X1 g117593(.A (n_14439), .B (n_19637), .Y (n_19646));
NAND2X1 g117598(.A (n_19647), .B (n_7988), .Y (n_19645));
NAND2X1 g117600(.A (n_18533), .B (n_19647), .Y (n_19643));
NAND2X1 g117610(.A (n_19626), .B (n_8946), .Y (n_19642));
NAND2X1 g117617(.A (n_35528), .B (n_19647), .Y (n_19641));
NAND2X1 g117640(.A (n_35822), .B (n_19637), .Y (n_19639));
NAND2X1 g117655(.A (n_17774), .B (n_33032), .Y (n_20200));
NAND2X1 g117705(.A (n_9629), .B (n_18311), .Y (n_19634));
NOR2X1 g117706(.A (n_21344), .B (n_20741), .Y (n_19633));
NAND2X1 g117710(.A (n_19631), .B (n_17727), .Y (n_19632));
NAND2X1 g117711(.A (n_19629), .B (n_17713), .Y (n_19630));
NAND2X1 g117713(.A (n_19626), .B (n_18498), .Y (n_19627));
NAND2X1 g117722(.A (n_19624), .B (n_17713), .Y (n_19625));
NAND2X1 g117735(.A (n_18302), .B (n_33803), .Y (n_19623));
AOI21X1 g117737(.A0 (n_17714), .A1 (n_27221), .B0 (n_21374), .Y(n_19622));
AOI21X1 g117746(.A0 (n_17711), .A1 (n_13628), .B0 (n_21374), .Y(n_19621));
NAND2X1 g117758(.A (n_9629), .B (n_18309), .Y (n_19620));
NAND2X1 g117766(.A (n_19624), .B (n_34418), .Y (n_19619));
OR2X1 g117782(.A (n_10023), .B (n_18307), .Y (n_19617));
AOI21X1 g117785(.A0 (n_17709), .A1 (n_26558), .B0 (n_10023), .Y(n_19616));
INVX1 g117786(.A (n_19614), .Y (n_19615));
OAI21X1 g117801(.A0 (n_17707), .A1 (n_14496), .B0 (n_20304), .Y(n_19613));
INVX1 g117806(.A (n_19611), .Y (n_20904));
NAND2X1 g117808(.A (n_19629), .B (n_23192), .Y (n_19610));
NAND2X1 g117810(.A (n_23190), .B (n_20830), .Y (n_19608));
NAND2X1 g117812(.A (n_19626), .B (n_27770), .Y (n_19607));
NOR2X1 g117820(.A (n_16808), .B (n_14261), .Y (n_19606));
NAND2X1 g117823(.A (n_19624), .B (n_27770), .Y (n_19605));
NOR2X1 g117828(.A (n_33556), .B (n_19000), .Y (n_19604));
NAND2X1 g117838(.A (n_18317), .B (n_20490), .Y (n_19603));
NAND2X1 g117843(.A (n_21703), .B (n_18942), .Y (n_19602));
INVX1 g117887(.A (n_19600), .Y (n_19601));
NAND2X1 g117896(.A (n_19631), .B (n_19597), .Y (n_19598));
NAND2X1 g117905(.A (n_19629), .B (n_19595), .Y (n_19596));
NAND3X1 g117913(.A (n_18291), .B (n_11816), .C (n_33749), .Y(n_23874));
NAND2X1 g117914(.A (n_19626), .B (n_26631), .Y (n_19593));
INVX1 g118023(.A (n_19589), .Y (n_19590));
NAND2X1 g118136(.A (n_18300), .B (n_22123), .Y (n_19584));
INVX1 g118159(.A (n_20265), .Y (n_19583));
NAND2X1 g118168(.A (n_20864), .B (n_19571), .Y (n_19582));
INVX1 g118184(.A (n_19581), .Y (n_21416));
NOR2X1 g118191(.A (n_33556), .B (n_17639), .Y (n_19580));
NAND2X1 g118192(.A (n_19631), .B (n_19577), .Y (n_19578));
NAND2X1 g118201(.A (n_19626), .B (n_27422), .Y (n_19576));
NAND3X1 g118214(.A (n_18285), .B (n_11990), .C (n_17822), .Y(n_21758));
NAND2X1 g118215(.A (n_19624), .B (n_17340), .Y (n_19575));
NAND2X1 g118225(.A (n_11732), .B (n_17776), .Y (n_20138));
NAND2X1 g118226(.A (n_19629), .B (n_19577), .Y (n_19573));
NAND2X1 g118260(.A (n_19571), .B (n_21328), .Y (n_19572));
NAND2X1 g118292(.A (n_20133), .B (n_19637), .Y (n_19570));
NAND2X1 g118293(.A (n_35479), .B (n_19637), .Y (n_19569));
NAND2X1 g118296(.A (n_21703), .B (n_18937), .Y (n_19568));
NAND2X1 g118306(.A (n_19637), .B (n_7988), .Y (n_19567));
NAND2X1 g118321(.A (n_20864), .B (n_19564), .Y (n_19566));
NAND2X1 g118322(.A (n_19564), .B (n_21328), .Y (n_19565));
NAND2X1 g118326(.A (n_19561), .B (n_21328), .Y (n_19563));
NAND2X1 g118327(.A (n_20864), .B (n_19561), .Y (n_19562));
NAND2X1 g118367(.A (n_20864), .B (n_19558), .Y (n_19560));
NAND2X1 g118368(.A (n_19558), .B (n_21328), .Y (n_19559));
NAND2X1 g118369(.A (n_20112), .B (n_19555), .Y (n_19557));
NAND2X1 g118371(.A (n_20112), .B (n_19552), .Y (n_19554));
NAND2X1 g118372(.A (n_19552), .B (n_21328), .Y (n_19553));
NAND2X1 g118378(.A (n_18940), .B (n_21328), .Y (n_19551));
INVX1 g118383(.A (n_21741), .Y (n_19550));
INVX1 g118390(.A (n_20242), .Y (n_19549));
INVX1 g118409(.A (n_19548), .Y (n_21745));
NAND2X1 g118440(.A (n_18342), .B (n_34800), .Y (n_19546));
INVX1 g118463(.A (n_19544), .Y (n_19545));
NOR2X1 g118466(.A (n_18396), .B (n_19031), .Y (n_20098));
INVX1 g118467(.A (n_19542), .Y (n_19543));
OAI21X1 g118470(.A0 (n_17863), .A1 (n_17161), .B0 (n_17864), .Y(n_21287));
NAND2X1 g118495(.A (n_18400), .B (n_26208), .Y (n_19541));
NAND2X1 g118501(.A (n_18389), .B (n_25702), .Y (n_19540));
NAND2X1 g118504(.A (n_18388), .B (n_26203), .Y (n_19539));
OAI21X1 g118513(.A0 (n_17116), .A1 (n_32720), .B0 (n_23181), .Y(n_19538));
NAND2X1 g118514(.A (n_18383), .B (n_25696), .Y (n_19537));
OAI21X1 g118517(.A0 (n_17637), .A1 (n_32774), .B0 (n_26199), .Y(n_19536));
NAND2X1 g118523(.A (n_18377), .B (n_24892), .Y (n_19534));
NAND2X1 g118525(.A (n_18376), .B (n_34690), .Y (n_19533));
NAND2X1 g118526(.A (n_18341), .B (n_25675), .Y (n_19532));
INVX1 g118540(.A (n_19530), .Y (n_19531));
NAND2X1 g118558(.A (n_18316), .B (n_32361), .Y (n_19529));
NAND2X1 g118584(.A (n_9516), .B (n_18339), .Y (n_19528));
OR2X1 g118587(.A (n_9163), .B (n_18338), .Y (n_19527));
NAND2X1 g118590(.A (n_9514), .B (n_18337), .Y (n_19526));
OAI21X1 g118595(.A0 (n_8325), .A1 (n_2693), .B0 (n_18336), .Y(n_19525));
AND2X1 g118729(.A (n_19052), .B (n_19524), .Y (n_20796));
NAND2X1 g118760(.A (n_17647), .B (n_25297), .Y (n_19522));
INVX1 g119068(.A (n_24490), .Y (n_19519));
NAND2X1 g119164(.A (n_17647), .B (n_25309), .Y (n_19516));
AND2X1 g119190(.A (n_17647), .B (n_18909), .Y (n_19513));
INVX1 g119199(.A (n_19510), .Y (n_19511));
INVX1 g119273(.A (n_19506), .Y (n_19507));
NAND2X1 g119283(.A (n_17155), .B (n_21733), .Y (n_20087));
NOR2X1 g119287(.A (n_19505), .B (n_17692), .Y (n_20085));
OAI22X1 g119291(.A0 (n_11961), .A1 (n_20741), .B0 (n_16796), .B1(n_16420), .Y (n_20083));
AOI21X1 g119384(.A0 (n_19471), .A1 (n_13268), .B0 (n_14593), .Y(n_19504));
INVX1 g119386(.A (n_18958), .Y (n_19503));
NAND2X1 g119427(.A (n_18279), .B (n_24190), .Y (n_19502));
NAND2X1 g119435(.A (n_18272), .B (n_27222), .Y (n_19501));
AOI21X1 g119443(.A0 (n_32739), .A1 (n_19474), .B0 (n_14104), .Y(n_19500));
OAI21X1 g119552(.A0 (n_13781), .A1 (n_16734), .B0 (n_34417), .Y(n_19498));
NAND2X1 g119560(.A (n_18271), .B (n_29667), .Y (n_19496));
AOI21X1 g119562(.A0 (n_16731), .A1 (n_32764), .B0 (n_19494), .Y(n_19495));
NAND2X1 g119564(.A (n_18268), .B (n_19492), .Y (n_19493));
NAND2X1 g119569(.A (n_18264), .B (n_29666), .Y (n_19491));
OAI21X1 g119570(.A0 (n_13588), .A1 (n_16734), .B0 (n_22097), .Y(n_19490));
NAND2X1 g119574(.A (n_18254), .B (n_28195), .Y (n_19489));
NAND2X1 g119648(.A (n_18274), .B (n_27687), .Y (n_20714));
NAND2X1 g119649(.A (n_18253), .B (n_27207), .Y (n_20711));
NAND2X1 g119654(.A (n_18261), .B (n_13347), .Y (n_20703));
NAND2X1 g119655(.A (n_18263), .B (n_13346), .Y (n_20706));
NAND2X1 g119659(.A (n_18258), .B (n_13499), .Y (n_20700));
INVX1 g119660(.A (n_19484), .Y (n_19485));
NAND2X1 g119662(.A (n_18260), .B (n_13372), .Y (n_20698));
INVX1 g119668(.A (n_19482), .Y (n_19483));
INVX1 g119671(.A (n_19480), .Y (n_19481));
NAND2X1 g119673(.A (n_18250), .B (n_27205), .Y (n_20717));
INVX1 g119676(.A (n_19478), .Y (n_19479));
INVX1 g119678(.A (n_19476), .Y (n_19477));
NAND2X1 g119681(.A (n_18252), .B (n_13917), .Y (n_20722));
NAND2X1 g119682(.A (n_18251), .B (n_14150), .Y (n_20720));
AOI22X1 g119687(.A0 (n_18289), .A1 (n_10081), .B0 (n_19474), .B1(n_18909), .Y (n_19475));
AOI22X1 g119695(.A0 (n_10573), .A1 (n_8207), .B0 (n_19471), .B1(n_8946), .Y (n_19473));
OAI21X1 g119696(.A0 (n_8981), .A1 (n_8511), .B0 (n_18249), .Y(n_19469));
NAND2X1 g119819(.A (n_17639), .B (n_27770), .Y (n_19468));
NAND2X1 g119959(.A (n_26637), .B (n_17639), .Y (n_19467));
AOI21X1 g113579(.A0 (n_17636), .A1 (n_21551), .B0 (n_8065), .Y(n_19463));
AOI21X1 g113596(.A0 (n_17634), .A1 (n_21550), .B0 (n_8065), .Y(n_19462));
NAND2X1 g113597(.A (n_19458), .B (n_22792), .Y (n_19461));
AOI21X1 g113613(.A0 (n_17632), .A1 (n_21549), .B0 (n_8065), .Y(n_19460));
NAND2X1 g113616(.A (n_19458), .B (n_32739), .Y (n_19459));
NAND2X1 g113633(.A (n_19458), .B (n_23696), .Y (n_19457));
XOR2X1 g113859(.A (n_16275), .B (n_20057), .Y (n_20060));
NAND2X1 g114023(.A (n_19454), .B (n_23149), .Y (n_19456));
NAND2X1 g114044(.A (n_19454), .B (n_23578), .Y (n_19455));
INVX1 g114077(.A (n_19452), .Y (n_19453));
NAND3X1 g114112(.A (n_19448), .B (n_18715), .C (n_18832), .Y(n_20049));
XOR2X1 g114548(.A (n_17273), .B (n_18896), .Y (n_20051));
XOR2X1 g114550(.A (n_16273), .B (n_21100), .Y (n_20038));
INVX1 g114551(.A (n_19454), .Y (n_19451));
AOI21X1 g114573(.A0 (n_18186), .A1 (n_16673), .B0 (n_18875), .Y(n_19447));
AOI21X1 g114607(.A0 (n_17624), .A1 (n_20022), .B0 (n_8065), .Y(n_19446));
OR2X1 g114622(.A (n_18234), .B (n_8065), .Y (n_19445));
AOI21X1 g114632(.A0 (n_17621), .A1 (n_20019), .B0 (n_8065), .Y(n_19443));
NAND2X1 g114663(.A (n_19441), .B (n_17618), .Y (n_19442));
NOR2X1 g114689(.A (n_21100), .B (n_18758), .Y (n_20042));
AOI21X1 g114727(.A0 (n_17546), .A1 (n_18183), .B0 (n_19403), .Y(n_19439));
NAND2X1 g114932(.A (n_19437), .B (n_33705), .Y (n_19438));
NAND2X1 g114939(.A (n_18160), .B (n_19187), .Y (n_21103));
NAND3X1 g114955(.A (n_15935), .B (n_17560), .C (n_17513), .Y(n_19436));
NAND2X1 g114958(.A (n_18787), .B (n_34066), .Y (n_19435));
NAND2X1 g114962(.A (n_19432), .B (n_22414), .Y (n_19434));
NAND2X1 g114989(.A (n_19432), .B (n_22406), .Y (n_19433));
NAND2X1 g114992(.A (n_19432), .B (n_32715), .Y (n_19431));
NAND2X1 g115005(.A (n_19423), .B (n_35054), .Y (n_19430));
NAND2X1 g115008(.A (n_19432), .B (n_25402), .Y (n_19429));
NAND2X1 g115011(.A (n_18807), .B (n_19372), .Y (n_19428));
NAND2X1 g115015(.A (n_18805), .B (n_19402), .Y (n_19427));
NAND2X1 g115017(.A (n_18803), .B (n_18125), .Y (n_19426));
NAND2X1 g115024(.A (n_18165), .B (n_19162), .Y (n_21105));
NAND3X1 g115044(.A (n_11781), .B (n_16937), .C (n_17466), .Y(n_21557));
NAND4X1 g115048(.A (n_11296), .B (n_16605), .C (n_16092), .D(n_16997), .Y (n_20614));
NOR2X1 g115064(.A (n_17865), .B (n_19401), .Y (n_19425));
NAND2X1 g115068(.A (n_19423), .B (n_22080), .Y (n_19424));
NAND2X1 g115089(.A (n_19422), .B (n_19411), .Y (n_20625));
NAND2X1 g115090(.A (n_14778), .B (n_19409), .Y (n_19421));
NAND2X1 g115093(.A (n_18174), .B (n_16675), .Y (n_19420));
NAND2X1 g115105(.A (n_18172), .B (n_18235), .Y (n_19419));
NAND2X1 g115110(.A (n_18878), .B (n_20031), .Y (n_19418));
NAND2X1 g115121(.A (n_18794), .B (n_18848), .Y (n_19417));
AND2X1 g115129(.A (n_20018), .B (n_20550), .Y (n_19416));
NAND2X1 g115173(.A (n_19414), .B (n_19413), .Y (n_19415));
NAND2X1 g115176(.A (n_19411), .B (n_14185), .Y (n_19412));
NAND2X1 g115180(.A (n_19410), .B (n_19409), .Y (n_19977));
NAND2X2 g115181(.A (n_19407), .B (n_16042), .Y (n_19408));
NAND2X1 g115187(.A (n_19405), .B (n_17524), .Y (n_19406));
NAND2X1 g115197(.A (n_18087), .B (n_19403), .Y (n_19404));
AOI21X1 g115209(.A0 (n_17500), .A1 (n_17568), .B0 (n_18194), .Y(n_19972));
NAND3X1 g115212(.A (n_19402), .B (n_16915), .C (n_17365), .Y(n_19969));
NOR3X1 g115213(.A (n_35360), .B (n_16635), .C (n_18049), .Y(n_20630));
OR2X1 g115216(.A (n_17783), .B (n_19401), .Y (n_21521));
INVX1 g115221(.A (n_19399), .Y (n_19400));
AND2X1 g115227(.A (n_19397), .B (n_18229), .Y (n_19398));
NAND2X1 g115236(.A (n_18195), .B (n_18033), .Y (n_20046));
INVX1 g115247(.A (n_19390), .Y (n_19391));
NAND2X1 g115293(.A (n_18188), .B (n_19389), .Y (n_20619));
AOI21X1 g115297(.A0 (n_17483), .A1 (n_18192), .B0 (n_19354), .Y(n_19959));
XOR2X1 g115306(.A (n_16564), .B (n_19948), .Y (n_20641));
XOR2X1 g115307(.A (n_18615), .B (n_20012), .Y (n_20639));
NOR2X1 g115320(.A (n_19388), .B (n_16552), .Y (n_20527));
NOR2X1 g115322(.A (n_19388), .B (n_17883), .Y (n_20571));
NAND2X1 g115327(.A (n_34680), .B (n_19302), .Y (n_19387));
INVX1 g115352(.A (n_19996), .Y (n_19385));
NAND2X1 g115356(.A (n_20431), .B (n_19383), .Y (n_19384));
NAND2X1 g115360(.A (n_18588), .B (n_35001), .Y (n_19382));
INVX1 g115382(.A (n_19381), .Y (n_19944));
NAND2X1 g115397(.A (n_18155), .B (n_18009), .Y (n_19380));
AOI21X1 g115398(.A0 (n_17410), .A1 (n_25055), .B0 (n_21374), .Y(n_19379));
NAND2X1 g115439(.A (n_18147), .B (n_17990), .Y (n_19378));
NAND2X1 g115450(.A (n_35671), .B (n_19377), .Y (n_19926));
AOI21X1 g115455(.A0 (n_17401), .A1 (n_25355), .B0 (n_21374), .Y(n_19376));
NOR2X1 g115472(.A (n_18671), .B (n_18153), .Y (n_19921));
NOR2X1 g115477(.A (n_19375), .B (n_19370), .Y (n_21870));
NOR2X1 g115480(.A (n_19371), .B (n_17068), .Y (n_21852));
NAND3X1 g115484(.A (n_17989), .B (n_11303), .C (n_19279), .Y(n_21020));
INVX2 g115495(.A (n_19374), .Y (n_21999));
NAND2X1 g115498(.A (n_19373), .B (n_19372), .Y (n_19913));
NOR2X1 g115503(.A (n_19923), .B (n_20465), .Y (n_22167));
NOR2X1 g115504(.A (n_18083), .B (n_18079), .Y (n_20574));
NOR2X1 g115513(.A (n_19371), .B (n_19370), .Y (n_21576));
INVX1 g115518(.A (n_19369), .Y (n_21459));
NAND2X1 g115521(.A (n_19368), .B (n_19367), .Y (n_19912));
INVX1 g115563(.A (n_18850), .Y (n_19900));
OR2X1 g115573(.A (n_19334), .B (n_18159), .Y (n_19366));
NAND2X1 g115588(.A (n_18004), .B (n_18021), .Y (n_20542));
NAND2X1 g115589(.A (n_18020), .B (n_17999), .Y (n_20541));
NAND2X1 g115590(.A (n_17994), .B (n_18019), .Y (n_21048));
NAND2X1 g115654(.A (n_19397), .B (n_33767), .Y (n_23053));
NAND2X1 g115673(.A (n_19874), .B (n_19365), .Y (n_19878));
NOR2X1 g115699(.A (n_18660), .B (n_17759), .Y (n_23521));
NOR2X1 g115705(.A (n_19364), .B (n_18078), .Y (n_20573));
NAND2X1 g115765(.A (n_19361), .B (n_20887), .Y (n_19363));
NAND2X1 g115766(.A (n_20112), .B (n_19361), .Y (n_19362));
AOI21X1 g115776(.A0 (n_17338), .A1 (n_24721), .B0 (n_21374), .Y(n_19360));
INVX1 g115797(.A (n_19359), .Y (n_19845));
NAND2X1 g115808(.A (n_18040), .B (n_21328), .Y (n_19358));
NAND2X1 g115810(.A (n_20864), .B (n_18574), .Y (n_19357));
NAND2X1 g115811(.A (n_17077), .B (n_16888), .Y (n_19356));
NAND2X1 g115820(.A (n_19354), .B (n_32878), .Y (n_19355));
NAND2X1 g115835(.A (n_18586), .B (n_17416), .Y (n_19353));
NOR2X1 g115845(.A (n_18636), .B (n_18658), .Y (n_19352));
NAND2X1 g115849(.A (n_19948), .B (n_20532), .Y (n_19351));
NOR2X1 g115850(.A (n_20399), .B (n_18581), .Y (n_19350));
NOR2X1 g115851(.A (n_20399), .B (n_18608), .Y (n_19348));
NAND2X1 g115853(.A (n_18034), .B (n_19213), .Y (n_19347));
NOR2X1 g115855(.A (n_20399), .B (n_18593), .Y (n_19346));
NAND2X1 g115858(.A (n_18029), .B (n_21328), .Y (n_19345));
NAND2X1 g115860(.A (n_17625), .B (n_20010), .Y (n_19344));
NAND2X1 g115862(.A (n_18031), .B (n_19212), .Y (n_19343));
NAND2X1 g115866(.A (n_18068), .B (n_17610), .Y (n_19342));
NAND2X1 g115877(.A (n_21703), .B (n_18576), .Y (n_19341));
NAND2X1 g115927(.A (n_18154), .B (n_17292), .Y (n_20567));
NAND2X1 g115932(.A (n_18143), .B (n_18815), .Y (n_20563));
NAND3X1 g115944(.A (n_16353), .B (n_20235), .C (n_18782), .Y(n_20041));
NAND2X1 g115945(.A (n_18126), .B (n_18814), .Y (n_20557));
INVX1 g115950(.A (n_19338), .Y (n_19339));
INVX1 g115956(.A (n_18821), .Y (n_19825));
INVX1 g115958(.A (n_19336), .Y (n_19337));
AOI21X1 g115964(.A0 (n_19208), .A1 (n_17963), .B0 (n_18778), .Y(n_21097));
NAND2X2 g115970(.A (n_19305), .B (n_35410), .Y (n_21525));
NAND2X1 g115977(.A (n_17550), .B (n_19334), .Y (n_20540));
AOI21X1 g115983(.A0 (n_17267), .A1 (n_17277), .B0 (n_18231), .Y(n_19333));
OAI21X1 g115998(.A0 (n_16991), .A1 (n_17605), .B0 (n_19259), .Y(n_19818));
NAND2X1 g116013(.A (n_18063), .B (n_18809), .Y (n_20528));
INVX1 g116017(.A (n_18816), .Y (n_19816));
AOI21X1 g116024(.A0 (n_17803), .A1 (n_19331), .B0 (n_18704), .Y(n_19332));
OAI21X1 g116025(.A0 (n_19330), .A1 (n_17402), .B0 (n_19329), .Y(n_20579));
NAND2X1 g116028(.A (n_18138), .B (n_19328), .Y (n_20577));
NAND2X1 g116029(.A (n_18136), .B (n_19327), .Y (n_20582));
INVX1 g116030(.A (n_19994), .Y (n_19326));
NAND2X1 g116032(.A (n_17070), .B (n_18696), .Y (n_21056));
NAND2X1 g116034(.A (n_18117), .B (n_18700), .Y (n_19813));
NAND2X1 g116042(.A (n_18066), .B (n_19325), .Y (n_20530));
INVX1 g116043(.A (n_19979), .Y (n_19324));
NAND2X1 g116052(.A (n_18130), .B (n_16589), .Y (n_19810));
NAND2X1 g116057(.A (n_18129), .B (n_16301), .Y (n_19323));
NAND2X1 g116059(.A (n_18128), .B (n_17084), .Y (n_19808));
INVX1 g116064(.A (n_19321), .Y (n_19322));
NAND2X1 g116074(.A (n_16938), .B (n_35700), .Y (n_19806));
OAI21X1 g116080(.A0 (n_17359), .A1 (n_19733), .B0 (n_17903), .Y(n_19804));
OAI21X1 g116084(.A0 (n_17898), .A1 (n_19320), .B0 (n_17895), .Y(n_19802));
INVX1 g116110(.A (n_19318), .Y (n_19319));
NAND2X1 g116113(.A (n_18064), .B (n_18170), .Y (n_19800));
NAND2X1 g116119(.A (n_18152), .B (n_18690), .Y (n_19797));
NAND2X2 g116121(.A (n_18122), .B (n_18102), .Y (n_19795));
INVX1 g116133(.A (n_19314), .Y (n_35869));
NAND2X1 g116139(.A (n_18110), .B (n_17446), .Y (n_19313));
CLKBUFX1 g116149(.A (n_19312), .Y (n_21858));
INVX1 g116170(.A (n_35715), .Y (n_19311));
AOI22X1 g116182(.A0 (n_11227), .A1 (n_34110), .B0 (n_35861), .B1(n_17975), .Y (n_19309));
NAND2X1 g116220(.A (n_20864), .B (n_19220), .Y (n_19308));
NAND2X1 g116221(.A (n_21703), .B (n_19214), .Y (n_19307));
NOR2X1 g116225(.A (n_18521), .B (n_18721), .Y (n_20500));
NAND2X1 g116228(.A (n_19212), .B (n_19306), .Y (n_19771));
NAND3X1 g116229(.A (n_19005), .B (n_17830), .C (n_18456), .Y(n_20495));
NAND2X1 g116231(.A (n_19305), .B (n_19304), .Y (n_19769));
INVX1 g116251(.A (n_19300), .Y (n_19761));
INVX1 g116261(.A (n_19298), .Y (n_19299));
INVX1 g116269(.A (n_20488), .Y (n_19297));
NAND2X1 g116280(.A (n_9629), .B (n_17858), .Y (n_19296));
NAND2X1 g116281(.A (n_9629), .B (n_17855), .Y (n_19295));
INVX2 g116284(.A (n_18766), .Y (n_20411));
NOR2X1 g116306(.A (n_17900), .B (n_19294), .Y (n_20395));
NAND2X1 g116319(.A (n_9629), .B (n_17854), .Y (n_32872));
NAND2X1 g116320(.A (n_9629), .B (n_17853), .Y (n_19291));
NAND2X1 g116328(.A (n_16633), .B (n_17446), .Y (n_19290));
INVX1 g116342(.A (n_19287), .Y (n_19288));
NAND2X1 g116356(.A (n_18410), .B (n_13274), .Y (n_19286));
INVX1 g116367(.A (n_19284), .Y (n_19285));
OR2X1 g116385(.A (n_10023), .B (n_17852), .Y (n_19282));
INVX1 g116433(.A (n_19280), .Y (n_20401));
OR2X1 g116440(.A (n_19279), .B (n_19905), .Y (n_20443));
NAND2X1 g116446(.A (n_20304), .B (n_17859), .Y (n_19278));
INVX1 g116449(.A (n_19277), .Y (n_19750));
NAND2X1 g116451(.A (n_20304), .B (n_17849), .Y (n_19276));
NAND2X1 g116452(.A (n_20304), .B (n_17851), .Y (n_19274));
INVX1 g116459(.A (n_22142), .Y (n_19273));
INVX1 g116463(.A (n_19271), .Y (n_19272));
INVX1 g116473(.A (n_18713), .Y (n_20462));
NOR2X1 g116475(.A (n_19167), .B (n_33556), .Y (n_19270));
NAND2X1 g116478(.A (n_16982), .B (n_17446), .Y (n_20459));
INVX1 g116482(.A (n_19268), .Y (n_20464));
NAND2X1 g116487(.A (n_16973), .B (n_17446), .Y (n_32949));
NOR2X1 g116492(.A (n_19228), .B (n_33000), .Y (n_19267));
NAND2X1 g116493(.A (n_18484), .B (n_18683), .Y (n_19266));
OR2X1 g116497(.A (n_19792), .B (n_33976), .Y (n_19743));
NAND3X1 g116533(.A (n_11210), .B (n_16739), .C (n_17185), .Y(n_19742));
NAND2X1 g116534(.A (n_18476), .B (n_19242), .Y (n_19263));
OR2X1 g116536(.A (n_33976), .B (n_20928), .Y (n_20829));
INVX1 g116537(.A (n_19262), .Y (n_20442));
INVX1 g116541(.A (n_19260), .Y (n_19261));
NAND2X1 g116544(.A (n_19259), .B (n_18096), .Y (n_19740));
INVX1 g116547(.A (n_19820), .Y (n_19258));
NAND2X1 g116560(.A (n_19788), .B (n_18765), .Y (n_21393));
NAND2X1 g116564(.A (n_19256), .B (n_19255), .Y (n_21392));
NAND2X1 g116566(.A (n_16938), .B (n_18074), .Y (n_22145));
INVX1 g116573(.A (n_23892), .Y (n_19253));
INVX1 g116577(.A (n_24137), .Y (n_19252));
NAND2X1 g116581(.A (n_16912), .B (n_17365), .Y (n_19734));
NOR2X1 g116582(.A (n_19876), .B (n_19235), .Y (n_19250));
NAND2X1 g116583(.A (n_19305), .B (n_16640), .Y (n_19249));
NAND2X1 g116588(.A (n_18541), .B (n_16972), .Y (n_19248));
OR2X1 g116599(.A (n_19247), .B (n_19294), .Y (n_21387));
NAND2X1 g116603(.A (n_19799), .B (n_18480), .Y (n_21389));
NAND2X1 g116604(.A (n_17896), .B (n_19245), .Y (n_19246));
INVX1 g116605(.A (n_21388), .Y (n_19244));
INVX1 g116609(.A (n_18679), .Y (n_20441));
NAND2X1 g116614(.A (n_19243), .B (n_19242), .Y (n_21735));
NAND2X1 g116625(.A (n_18478), .B (n_18091), .Y (n_19241));
NAND3X1 g116632(.A (n_16836), .B (n_16505), .C (n_18457), .Y(n_20061));
NAND2X1 g116633(.A (n_19239), .B (n_19238), .Y (n_19240));
NAND2X1 g116635(.A (n_18424), .B (n_19236), .Y (n_19237));
NAND3X1 g116685(.A (n_17832), .B (n_11989), .C (n_18518), .Y(n_21760));
AND2X1 g116706(.A (n_18695), .B (n_19235), .Y (n_19721));
NAND2X1 g116713(.A (n_18486), .B (n_18717), .Y (n_19234));
INVX1 g116718(.A (n_19233), .Y (n_20486));
NAND2X1 g116720(.A (n_17974), .B (n_18061), .Y (n_19232));
NAND2X1 g116722(.A (n_18417), .B (n_19230), .Y (n_19231));
NOR2X1 g116728(.A (n_19229), .B (n_18535), .Y (n_19719));
NOR2X1 g116729(.A (n_19228), .B (n_19225), .Y (n_21480));
NAND2X1 g116734(.A (n_18506), .B (n_21328), .Y (n_19227));
OR2X1 g116739(.A (n_22369), .B (n_19225), .Y (n_32614));
NAND2X1 g116744(.A (n_17930), .B (n_21328), .Y (n_19222));
NAND2X1 g116747(.A (n_19220), .B (n_21328), .Y (n_19221));
INVX1 g116761(.A (n_19873), .Y (n_19219));
INVX1 g116793(.A (n_19217), .Y (n_19218));
NAND2X1 g116801(.A (n_19214), .B (n_21328), .Y (n_19215));
NAND2X1 g116804(.A (n_19213), .B (n_19212), .Y (n_19712));
NAND2X1 g116820(.A (n_19210), .B (n_17446), .Y (n_19211));
NAND2X1 g116821(.A (n_17962), .B (n_16973), .Y (n_19209));
NAND2X1 g116824(.A (n_16970), .B (n_19208), .Y (n_19707));
NAND2X1 g116834(.A (n_19229), .B (n_16972), .Y (n_24977));
INVX1 g116838(.A (n_18642), .Y (n_20439));
NOR2X1 g116843(.A (n_19206), .B (n_17439), .Y (n_19207));
AND2X1 g116844(.A (n_17441), .B (n_17570), .Y (n_19205));
INVX1 g116846(.A (n_19203), .Y (n_19204));
NOR2X1 g116848(.A (n_19790), .B (n_19169), .Y (n_20388));
OR2X1 g116849(.A (n_34386), .B (n_17861), .Y (n_19202));
INVX1 g116851(.A (n_19200), .Y (n_19201));
NAND2X1 g116855(.A (n_19198), .B (n_19302), .Y (n_19702));
NOR2X1 g116858(.A (n_18454), .B (n_18637), .Y (n_32366));
INVX1 g116862(.A (n_19784), .Y (n_19195));
NAND2X1 g116864(.A (n_17827), .B (n_17826), .Y (n_20513));
INVX1 g116874(.A (n_19193), .Y (n_20368));
NAND2X1 g116879(.A (n_22369), .B (n_19228), .Y (n_19192));
NOR2X1 g116880(.A (n_17363), .B (n_19228), .Y (n_20406));
NAND2X1 g116881(.A (n_22369), .B (n_17886), .Y (n_20446));
INVX1 g116884(.A (n_19191), .Y (n_20404));
NAND2X1 g116887(.A (n_9629), .B (n_17839), .Y (n_19190));
NAND2X1 g116890(.A (n_9629), .B (n_17836), .Y (n_19189));
NAND4X1 g116913(.A (n_19187), .B (n_12350), .C (n_16793), .D(n_16733), .Y (n_20510));
AND2X1 g116916(.A (n_19186), .B (n_34996), .Y (n_20839));
OAI21X1 g116924(.A0 (n_19179), .A1 (n_13318), .B0 (n_25056), .Y(n_19184));
NAND2X1 g116929(.A (n_18474), .B (n_19183), .Y (n_19693));
NAND2X1 g116932(.A (n_34386), .B (n_17390), .Y (n_19690));
OAI21X1 g116936(.A0 (n_19172), .A1 (n_13990), .B0 (n_21890), .Y(n_19182));
OAI21X1 g116941(.A0 (n_19179), .A1 (n_13990), .B0 (n_25051), .Y(n_19180));
NAND2X1 g116947(.A (n_17919), .B (n_18855), .Y (n_19178));
OAI21X1 g116948(.A0 (n_19172), .A1 (n_25694), .B0 (n_21889), .Y(n_19177));
NAND2X1 g116951(.A (n_17917), .B (n_25689), .Y (n_19175));
OAI21X1 g116965(.A0 (n_19179), .A1 (n_13147), .B0 (n_25058), .Y(n_19174));
OAI21X1 g116974(.A0 (n_19172), .A1 (n_19165), .B0 (n_21885), .Y(n_19173));
AOI21X1 g116978(.A0 (n_18560), .A1 (n_17772), .B0 (n_16847), .Y(n_19171));
INVX1 g116988(.A (n_20621), .Y (n_19170));
NOR2X1 g116992(.A (n_20763), .B (n_19169), .Y (n_20499));
NAND2X1 g116996(.A (n_34386), .B (n_19167), .Y (n_19168));
OAI21X1 g117001(.A0 (n_19179), .A1 (n_19165), .B0 (n_25047), .Y(n_19166));
OAI21X1 g117009(.A0 (n_19172), .A1 (n_13318), .B0 (n_21892), .Y(n_19164));
NAND2X1 g117011(.A (n_17939), .B (n_26398), .Y (n_19685));
NAND4X1 g117012(.A (n_32888), .B (n_12054), .C (n_16455), .D(n_19162), .Y (n_20469));
OAI21X1 g117042(.A0 (n_19159), .A1 (n_13318), .B0 (n_21942), .Y(n_19161));
OAI21X1 g117046(.A0 (n_19159), .A1 (n_13990), .B0 (n_21941), .Y(n_19160));
OAI21X1 g117050(.A0 (n_19159), .A1 (n_25694), .B0 (n_21939), .Y(n_19158));
OAI21X1 g117052(.A0 (n_19159), .A1 (n_19165), .B0 (n_21940), .Y(n_19157));
NOR2X1 g117057(.A (n_17947), .B (n_13933), .Y (n_19679));
NOR2X1 g117059(.A (n_17940), .B (n_13899), .Y (n_19677));
NAND2X1 g117061(.A (n_17943), .B (n_23401), .Y (n_20373));
INVX1 g117062(.A (n_19155), .Y (n_19156));
INVX1 g117064(.A (n_19153), .Y (n_19154));
NOR2X1 g117068(.A (n_17942), .B (n_13937), .Y (n_19675));
NAND2X1 g117070(.A (n_17948), .B (n_24711), .Y (n_20396));
NOR2X1 g117079(.A (n_17945), .B (n_13900), .Y (n_19673));
INVX1 g117080(.A (n_19151), .Y (n_19152));
INVX1 g117082(.A (n_19149), .Y (n_19150));
INVX1 g117102(.A (n_19147), .Y (n_19148));
NAND2X1 g117107(.A (n_17967), .B (n_24713), .Y (n_20389));
NAND2X1 g117108(.A (n_17986), .B (n_27204), .Y (n_20384));
NAND2X1 g117121(.A (n_17980), .B (n_23418), .Y (n_19671));
NOR2X1 g117124(.A (n_18580), .B (n_35303), .Y (n_19146));
INVX1 g117146(.A (n_19142), .Y (n_19143));
AND2X1 g117151(.A (n_17956), .B (n_19140), .Y (n_19141));
INVX1 g117156(.A (n_19138), .Y (n_19139));
INVX1 g117160(.A (n_19136), .Y (n_19137));
NAND2X1 g117172(.A (n_17987), .B (n_24719), .Y (n_20433));
NAND2X1 g117179(.A (n_17971), .B (n_26401), .Y (n_20427));
NAND2X1 g117183(.A (n_17969), .B (n_23379), .Y (n_19663));
AOI21X1 g117198(.A0 (n_19135), .A1 (n_17767), .B0 (n_16746), .Y(n_19661));
NAND2X1 g117201(.A (n_17879), .B (n_17230), .Y (n_19659));
AOI21X1 g117203(.A0 (n_32837), .A1 (n_17768), .B0 (n_19135), .Y(n_20970));
INVX1 g117204(.A (n_19133), .Y (n_19134));
INVX1 g117206(.A (n_19131), .Y (n_19132));
INVX1 g117208(.A (n_19129), .Y (n_19130));
AOI21X1 g117212(.A0 (n_17993), .A1 (n_7988), .B0 (n_9010), .Y(n_19128));
INVX1 g117214(.A (n_35062), .Y (n_19127));
OAI21X1 g117221(.A0 (n_8981), .A1 (n_2837), .B0 (n_17944), .Y(n_19125));
AOI21X1 g117222(.A0 (n_19626), .A1 (n_33967), .B0 (n_10667), .Y(n_19124));
INVX1 g117236(.A (n_19122), .Y (n_19123));
INVX1 g117247(.A (n_19120), .Y (n_19121));
AOI21X1 g117258(.A0 (n_17997), .A1 (n_7988), .B0 (n_9011), .Y(n_19119));
OAI21X1 g117260(.A0 (n_9520), .A1 (n_3493), .B0 (n_17938), .Y(n_19117));
INVX1 g117262(.A (n_18572), .Y (n_19655));
INVX1 g117266(.A (n_19115), .Y (n_19116));
INVX1 g117295(.A (n_18567), .Y (n_19114));
AOI22X1 g117297(.A0 (n_18511), .A1 (n_8946), .B0 (n_20218), .B1(n_1003), .Y (n_19113));
AOI22X1 g117300(.A0 (n_11055), .A1 (n_19629), .B0 (n_9776), .B1(n_19626), .Y (n_19111));
AOI22X1 g117301(.A0 (n_17906), .A1 (n_16403), .B0 (n_16419), .B1(n_17384), .Y (n_19110));
AOI22X1 g117313(.A0 (n_32984), .A1 (n_19108), .B0 (n_11138), .B1(n_13327), .Y (n_19109));
AOI22X1 g117316(.A0 (n_18005), .A1 (n_19108), .B0 (n_11138), .B1(n_13370), .Y (n_19107));
AOI22X1 g117324(.A0 (n_17916), .A1 (n_19071), .B0 (n_12703), .B1(n_17732), .Y (n_19105));
AOI22X1 g117327(.A0 (n_34384), .A1 (n_33551), .B0 (n_18496), .B1(n_34385), .Y (n_19104));
AOI21X1 g117332(.A0 (n_11987), .A1 (n_17830), .B0 (n_18580), .Y(n_21013));
NAND2X1 g117357(.A (n_17968), .B (n_17975), .Y (n_19103));
NOR2X1 g117454(.A (n_35719), .B (n_16800), .Y (n_19102));
NAND2X1 g117463(.A (n_35776), .B (n_17975), .Y (n_19101));
INVX1 g117475(.A (n_19706), .Y (n_20270));
NAND2X1 g117555(.A (n_10754), .B (n_19098), .Y (n_19099));
NAND2X1 g117615(.A (n_35679), .B (n_8946), .Y (n_19097));
NAND2X1 g117636(.A (n_18533), .B (n_17975), .Y (n_19095));
NAND2X1 g117643(.A (n_10270), .B (n_19523), .Y (n_20224));
INVX1 g117647(.A (n_19093), .Y (n_19094));
NOR2X1 g117679(.A (n_16869), .B (n_18397), .Y (n_21379));
NAND2X1 g117689(.A (n_35679), .B (n_19577), .Y (n_19090));
INVX1 g117692(.A (n_21385), .Y (n_19088));
NAND2X1 g117708(.A (n_19085), .B (n_17713), .Y (n_19086));
INVX1 g117761(.A (n_20261), .Y (n_19084));
OR2X1 g117768(.A (n_21201), .B (n_17729), .Y (n_19083));
NAND2X1 g117783(.A (n_35679), .B (n_21919), .Y (n_19082));
NAND2X1 g117787(.A (n_16238), .B (n_17773), .Y (n_19614));
NAND2X1 g117802(.A (n_19085), .B (n_27770), .Y (n_19081));
NAND2X1 g117805(.A (n_19631), .B (n_27770), .Y (n_19080));
NAND2X1 g117807(.A (n_19079), .B (n_18351), .Y (n_19611));
NAND2X1 g117839(.A (n_17793), .B (n_17183), .Y (n_22501));
NAND2X1 g117877(.A (n_19085), .B (n_19595), .Y (n_19076));
INVX1 g117889(.A (n_19075), .Y (n_19600));
NAND2X1 g117907(.A (n_35679), .B (n_27770), .Y (n_19074));
NOR2X1 g117927(.A (n_19073), .B (n_17789), .Y (n_19591));
NAND2X1 g117953(.A (n_19071), .B (n_17732), .Y (n_19072));
OR2X1 g118024(.A (n_16855), .B (n_19043), .Y (n_19589));
INVX1 g118100(.A (n_20338), .Y (n_19068));
INVX1 g118120(.A (n_19689), .Y (n_19587));
AND2X1 g118142(.A (n_19065), .B (n_20361), .Y (n_21769));
INVX1 g118143(.A (n_19063), .Y (n_19064));
INVX1 g118146(.A (n_20412), .Y (n_19062));
NAND2X1 g118150(.A (n_19520), .B (n_34608), .Y (n_20354));
NAND2X1 g118160(.A (n_18475), .B (n_21344), .Y (n_20265));
NAND4X1 g118165(.A (n_12175), .B (n_20301), .C (n_17136), .D(n_16749), .Y (n_20315));
NAND2X1 g118185(.A (n_19061), .B (n_19060), .Y (n_19581));
INVX1 g118187(.A (n_34509), .Y (n_19059));
NAND2X1 g118210(.A (n_35679), .B (n_19595), .Y (n_19058));
NAND2X1 g118221(.A (n_19085), .B (n_19577), .Y (n_19057));
NAND2X1 g118222(.A (n_17725), .B (n_17723), .Y (n_20628));
INVX1 g118262(.A (n_19055), .Y (n_19056));
OR2X1 g118265(.A (n_19474), .B (n_19520), .Y (n_21690));
NAND3X1 g118280(.A (n_17172), .B (n_17146), .C (n_16732), .Y(n_19053));
NAND3X1 g118290(.A (n_17831), .B (n_19052), .C (n_16407), .Y(n_20056));
NAND2X1 g118384(.A (n_17256), .B (n_17330), .Y (n_21741));
AND2X1 g118391(.A (n_17230), .B (n_17878), .Y (n_20242));
INVX1 g118400(.A (n_20241), .Y (n_19051));
INVX1 g118402(.A (n_21742), .Y (n_19050));
NAND2X1 g118410(.A (n_19049), .B (n_19048), .Y (n_19548));
AOI21X1 g118418(.A0 (n_17710), .A1 (n_18434), .B0 (n_18433), .Y(n_19045));
AND2X1 g118421(.A (n_19044), .B (n_18412), .Y (n_22867));
NAND2X1 g118433(.A (n_17813), .B (n_19043), .Y (n_20822));
INVX1 g118434(.A (n_19041), .Y (n_19042));
INVX1 g118436(.A (n_19039), .Y (n_19040));
OAI21X1 g118441(.A0 (n_19005), .A1 (n_19037), .B0 (n_26216), .Y(n_19038));
NAND2X1 g118458(.A (n_17795), .B (n_25271), .Y (n_19036));
AOI21X1 g118460(.A0 (n_16748), .A1 (n_21733), .B0 (n_17137), .Y(n_19035));
INVX1 g118461(.A (n_19032), .Y (n_19033));
OAI21X1 g118464(.A0 (n_17166), .A1 (n_18428), .B0 (n_18395), .Y(n_19544));
AOI21X1 g118468(.A0 (n_18773), .A1 (n_19031), .B0 (n_17690), .Y(n_19542));
AND2X1 g118478(.A (n_17804), .B (n_18705), .Y (n_20818));
NOR2X1 g118479(.A (n_17764), .B (n_16783), .Y (n_20819));
INVX1 g118482(.A (n_19029), .Y (n_19030));
INVX1 g118485(.A (n_19027), .Y (n_19028));
OAI21X1 g118493(.A0 (n_19005), .A1 (n_19024), .B0 (n_26193), .Y(n_19026));
NAND2X1 g118498(.A (n_17816), .B (n_22839), .Y (n_19023));
NAND2X1 g118499(.A (n_17815), .B (n_25351), .Y (n_19022));
NAND2X1 g118500(.A (n_17812), .B (n_23136), .Y (n_19021));
OAI21X1 g118502(.A0 (n_19005), .A1 (n_13843), .B0 (n_26207), .Y(n_19020));
OAI21X1 g118505(.A0 (n_16836), .A1 (n_22042), .B0 (n_22836), .Y(n_19019));
OAI21X1 g118508(.A0 (n_16837), .A1 (n_32784), .B0 (n_24309), .Y(n_19017));
OAI21X1 g118509(.A0 (n_16836), .A1 (n_32718), .B0 (n_24897), .Y(n_19016));
OAI21X1 g118510(.A0 (n_17112), .A1 (n_32698), .B0 (n_13639), .Y(n_19014));
NAND2X1 g118512(.A (n_17806), .B (n_25264), .Y (n_19013));
OAI21X1 g118515(.A0 (n_19005), .A1 (n_32784), .B0 (n_26202), .Y(n_19012));
NAND2X1 g118521(.A (n_17799), .B (n_24895), .Y (n_19011));
NAND2X1 g118522(.A (n_17796), .B (n_25344), .Y (n_19010));
INVX1 g118538(.A (n_19008), .Y (n_35114));
AOI21X1 g118541(.A0 (n_17155), .A1 (n_17740), .B0 (n_19044), .Y(n_19530));
OR2X1 g118546(.A (n_17765), .B (n_18437), .Y (n_20511));
OAI21X1 g118547(.A0 (n_32417), .A1 (n_17304), .B0 (n_21603), .Y(n_19007));
AOI21X1 g118580(.A0 (n_11278), .A1 (n_19005), .B0 (n_17808), .Y(n_19006));
OR2X1 g118581(.A (n_9018), .B (n_17752), .Y (n_19004));
AOI21X1 g118582(.A0 (n_18289), .A1 (n_7664), .B0 (n_17750), .Y(n_19003));
AOI21X1 g118585(.A0 (n_18289), .A1 (n_3100), .B0 (n_17754), .Y(n_19001));
NAND2X1 g118750(.A (n_18997), .B (n_18340), .Y (n_18999));
NAND2X1 g118780(.A (n_18997), .B (n_18384), .Y (n_18998));
NAND2X1 g118802(.A (n_18997), .B (n_32777), .Y (n_18996));
NAND2X1 g118821(.A (n_17092), .B (n_34688), .Y (n_18994));
NAND2X1 g118835(.A (n_18997), .B (n_18907), .Y (n_18993));
NAND2X1 g118870(.A (n_17162), .B (n_16785), .Y (n_18989));
INVX4 g118900(.A (n_17776), .Y (n_19520));
INVX1 g119040(.A (n_21302), .Y (n_18984));
NAND2X1 g119069(.A (n_18981), .B (n_18255), .Y (n_24490));
NOR2X1 g119070(.A (n_17740), .B (n_17174), .Y (n_18980));
INVX1 g119098(.A (n_18978), .Y (n_18979));
INVX1 g119102(.A (n_18976), .Y (n_18977));
NAND2X1 g119192(.A (n_17092), .B (n_10848), .Y (n_18974));
NAND2X1 g119195(.A (n_18997), .B (n_18909), .Y (n_18971));
NAND2X1 g119200(.A (n_16785), .B (n_18969), .Y (n_19510));
INVX1 g119211(.A (n_18968), .Y (n_19508));
INVX1 g119213(.A (n_20212), .Y (n_18967));
NOR2X1 g119225(.A (n_17653), .B (n_18275), .Y (n_18964));
NAND2X1 g119274(.A (n_16430), .B (n_32361), .Y (n_19506));
INVX1 g119277(.A (n_18960), .Y (n_18961));
NAND2X1 g119385(.A (n_17706), .B (n_27068), .Y (n_18959));
AOI21X1 g119387(.A0 (n_18948), .A1 (n_20154), .B0 (n_14286), .Y(n_18958));
NAND2X1 g119389(.A (n_17704), .B (n_13174), .Y (n_18957));
NAND2X1 g119401(.A (n_17705), .B (n_26569), .Y (n_18956));
NAND2X1 g119426(.A (n_17721), .B (n_27064), .Y (n_18954));
NAND2X1 g119428(.A (n_17720), .B (n_26564), .Y (n_18953));
NAND2X1 g119434(.A (n_17717), .B (n_24675), .Y (n_18952));
NAND2X1 g119436(.A (n_17716), .B (n_14128), .Y (n_32209));
AOI21X1 g119442(.A0 (n_32715), .A1 (n_18948), .B0 (n_14297), .Y(n_18950));
AOI21X1 g119554(.A0 (n_18294), .A1 (n_16396), .B0 (n_13482), .Y(n_18947));
NAND2X1 g119563(.A (n_17703), .B (n_35057), .Y (n_18946));
NAND2X1 g119567(.A (n_17691), .B (n_27217), .Y (n_18945));
NAND2X1 g119573(.A (n_17675), .B (n_27227), .Y (n_18944));
INVX1 g119619(.A (n_18942), .Y (n_18943));
NAND2X1 g119624(.A (n_17672), .B (n_28322), .Y (n_20185));
NOR2X1 g119625(.A (n_17673), .B (n_13941), .Y (n_20160));
NAND2X1 g119626(.A (n_17659), .B (n_29545), .Y (n_20136));
NAND2X1 g119644(.A (n_17661), .B (n_28058), .Y (n_20165));
NAND2X1 g119651(.A (n_17684), .B (n_28054), .Y (n_20116));
NOR2X1 g119652(.A (n_17718), .B (n_13350), .Y (n_20114));
NAND2X1 g119656(.A (n_17685), .B (n_28310), .Y (n_20119));
INVX1 g119657(.A (n_18940), .Y (n_18941));
NAND2X1 g119661(.A (n_17683), .B (n_28302), .Y (n_19484));
NAND2X1 g119666(.A (n_17681), .B (n_28083), .Y (n_20109));
NAND2X1 g119667(.A (n_17679), .B (n_29478), .Y (n_20106));
NAND2X1 g119669(.A (n_17670), .B (n_18939), .Y (n_19482));
NOR2X1 g119672(.A (n_17664), .B (n_13922), .Y (n_19480));
INVX1 g119674(.A (n_18937), .Y (n_18938));
NAND2X1 g119677(.A (n_17669), .B (n_18936), .Y (n_19478));
NAND2X1 g119679(.A (n_17668), .B (n_29480), .Y (n_19476));
NOR2X1 g119680(.A (n_17666), .B (n_14151), .Y (n_20122));
AOI22X1 g119685(.A0 (n_18289), .A1 (n_9209), .B0 (n_18948), .B1(n_10848), .Y (n_18935));
AOI22X1 g119694(.A0 (n_10573), .A1 (n_7957), .B0 (n_18275), .B1(n_8946), .Y (n_18933));
OAI21X1 g119697(.A0 (n_8981), .A1 (n_8515), .B0 (n_17649), .Y(n_18931));
AOI21X1 g119699(.A0 (n_17655), .A1 (n_17592), .B0 (n_17687), .Y(n_18930));
OAI21X1 g119702(.A0 (n_9520), .A1 (n_10103), .B0 (n_17660), .Y(n_18929));
OAI21X1 g119704(.A0 (n_9520), .A1 (n_10119), .B0 (n_17662), .Y(n_18927));
OAI22X1 g119706(.A0 (n_9520), .A1 (n_3601), .B0 (n_17186), .B1(n_8309), .Y (n_18926));
XOR2X1 g119713(.A (n_16452), .B (n_23778), .Y (n_18924));
NAND2X1 g119741(.A (n_26530), .B (n_18917), .Y (n_18923));
NAND2X1 g119747(.A (n_18399), .B (n_19474), .Y (n_18922));
NAND2X1 g119753(.A (n_18399), .B (n_16411), .Y (n_18921));
NAND2X1 g119767(.A (n_20178), .B (n_19471), .Y (n_18920));
NAND2X1 g119768(.A (n_18918), .B (n_18917), .Y (n_18919));
NAND2X1 g119773(.A (n_15089), .B (n_19474), .Y (n_18916));
NAND2X1 g119777(.A (n_22064), .B (n_16411), .Y (n_18914));
NAND2X1 g119784(.A (n_19577), .B (n_19471), .Y (n_18912));
NAND2X1 g119790(.A (n_32739), .B (n_18917), .Y (n_18911));
NAND2X1 g119803(.A (n_18917), .B (n_18909), .Y (n_18910));
NAND2X1 g119808(.A (n_19474), .B (n_18907), .Y (n_18908));
NAND2X1 g119810(.A (n_18917), .B (n_24984), .Y (n_18906));
NAND2X1 g119887(.A (n_17340), .B (n_19471), .Y (n_18904));
NOR2X1 g113580(.A (n_18237), .B (n_20054), .Y (n_18902));
NOR2X1 g114014(.A (n_17418), .B (n_18898), .Y (n_20063));
OR2X1 g114078(.A (n_20057), .B (n_18900), .Y (n_19452));
NAND2X1 g114164(.A (n_18236), .B (n_21548), .Y (n_18899));
INVX1 g114554(.A (n_18898), .Y (n_19448));
NAND3X1 g114628(.A (n_18146), .B (n_18894), .C (n_18897), .Y(n_21145));
NOR2X1 g114715(.A (n_16561), .B (n_18896), .Y (n_19440));
AOI21X1 g114802(.A0 (n_17082), .A1 (n_16670), .B0 (n_18871), .Y(n_18895));
XOR2X1 g114904(.A (n_18833), .B (n_18894), .Y (n_19454));
NAND2X2 g114934(.A (n_17493), .B (n_35258), .Y (n_20035));
NAND2X1 g114961(.A (n_18891), .B (n_22414), .Y (n_18893));
NAND2X1 g114988(.A (n_18891), .B (n_18384), .Y (n_18892));
NAND2X1 g115007(.A (n_18891), .B (n_25404), .Y (n_18890));
NAND2X1 g115013(.A (n_18888), .B (n_17520), .Y (n_18889));
NAND2X1 g115018(.A (n_17598), .B (n_17565), .Y (n_18887));
NAND2X1 g115021(.A (n_18885), .B (n_18852), .Y (n_18886));
NAND3X1 g115051(.A (n_11295), .B (n_16323), .C (n_17001), .Y(n_18884));
NOR2X1 g115053(.A (n_17627), .B (n_10475), .Y (n_18883));
NAND2X1 g115092(.A (n_17620), .B (n_16389), .Y (n_18882));
NAND2X1 g115097(.A (n_18182), .B (n_16696), .Y (n_18881));
NAND2X1 g115098(.A (n_18176), .B (n_17587), .Y (n_18880));
NAND2X1 g115100(.A (n_18878), .B (n_17049), .Y (n_32123));
NAND2X1 g115101(.A (n_17597), .B (n_17048), .Y (n_18877));
NAND2X1 g115103(.A (n_18875), .B (n_17574), .Y (n_18876));
NAND2X1 g115104(.A (n_18873), .B (n_35672), .Y (n_32293));
NAND2X1 g115186(.A (n_18871), .B (n_34063), .Y (n_18872));
NAND2X1 g115222(.A (n_17616), .B (n_18171), .Y (n_19399));
INVX1 g115224(.A (n_18868), .Y (n_18870));
AOI21X1 g115246(.A0 (n_17497), .A1 (n_16886), .B0 (n_18828), .Y(n_18865));
NAND2X2 g115248(.A (n_17611), .B (n_18140), .Y (n_19390));
NAND2X1 g115253(.A (n_17622), .B (n_20021), .Y (n_18864));
NAND3X1 g115289(.A (n_16578), .B (n_16645), .C (n_17009), .Y(n_18862));
NAND2X1 g115318(.A (n_17494), .B (n_16283), .Y (n_18861));
NAND2X1 g115332(.A (n_18859), .B (n_18632), .Y (n_18860));
NOR2X1 g115353(.A (n_18139), .B (n_17532), .Y (n_19996));
NOR2X1 g115374(.A (n_18118), .B (n_34552), .Y (n_18858));
NOR2X1 g115383(.A (n_18080), .B (n_18156), .Y (n_19381));
NAND3X1 g115415(.A (n_17470), .B (n_11063), .C (n_17406), .Y(n_20017));
NAND2X1 g115496(.A (n_18857), .B (n_18856), .Y (n_19374));
NAND3X1 g115499(.A (n_17923), .B (n_18855), .C (n_17918), .Y(n_19992));
INVX1 g115511(.A (n_20552), .Y (n_18854));
NAND2X1 g115519(.A (n_18853), .B (n_18852), .Y (n_19369));
NAND2X1 g115558(.A (n_17475), .B (n_17488), .Y (n_18851));
NAND2X1 g115564(.A (n_18849), .B (n_18848), .Y (n_18850));
NAND2X1 g115565(.A (n_17469), .B (n_17487), .Y (n_20014));
NOR2X1 g115584(.A (n_17527), .B (n_11333), .Y (n_18847));
NAND2X1 g115585(.A (n_17481), .B (n_17486), .Y (n_19966));
NOR2X1 g115632(.A (n_18843), .B (n_17573), .Y (n_21011));
NOR2X1 g115635(.A (n_17539), .B (n_17525), .Y (n_21440));
NOR2X1 g115639(.A (n_18834), .B (n_18846), .Y (n_21031));
INVX1 g115640(.A (n_18844), .Y (n_18845));
INVX1 g115649(.A (n_20652), .Y (n_18842));
NAND2X1 g115676(.A (n_19958), .B (n_20033), .Y (n_18841));
NAND3X1 g115762(.A (n_17885), .B (n_16890), .C (n_16502), .Y(n_21823));
NOR2X1 g115772(.A (n_35719), .B (n_17583), .Y (n_18840));
NAND2X1 g115798(.A (n_17540), .B (n_19413), .Y (n_19359));
NOR2X1 g115806(.A (n_10021), .B (n_18039), .Y (n_18839));
NAND2X1 g115813(.A (n_16943), .B (n_33771), .Y (n_18838));
INVX1 g115843(.A (n_18193), .Y (n_19975));
NAND2X1 g115846(.A (n_18035), .B (n_18060), .Y (n_18836));
NOR2X1 g115857(.A (n_20399), .B (n_18028), .Y (n_18835));
NOR2X1 g115867(.A (n_17053), .B (n_18834), .Y (n_21008));
AND2X1 g115869(.A (n_17589), .B (n_16353), .Y (n_21780));
NAND3X1 g115870(.A (n_18833), .B (n_16590), .C (n_18832), .Y(n_20009));
NOR2X1 g115876(.A (n_17521), .B (n_33983), .Y (n_21506));
NOR2X1 g115879(.A (n_33983), .B (n_18052), .Y (n_18830));
NAND2X1 g115886(.A (n_18828), .B (n_17316), .Y (n_18829));
NAND3X1 g115949(.A (n_18824), .B (n_35364), .C (n_16636), .Y(n_35870));
AOI21X1 g115951(.A0 (n_19206), .A1 (n_17570), .B0 (n_18736), .Y(n_19338));
AOI21X1 g115953(.A0 (n_18584), .A1 (n_17570), .B0 (n_18583), .Y(n_18823));
NAND2X1 g115957(.A (n_17562), .B (n_18644), .Y (n_18821));
OAI21X1 g115959(.A0 (n_16974), .A1 (n_19210), .B0 (n_17443), .Y(n_19336));
INVX1 g115961(.A (n_18819), .Y (n_18820));
INVX1 g115967(.A (n_19437), .Y (n_19335));
NAND2X1 g116015(.A (n_32577), .B (n_32578), .Y (n_32379));
NAND2X1 g116018(.A (n_17535), .B (n_17606), .Y (n_18816));
NAND2X1 g116026(.A (n_17588), .B (n_17292), .Y (n_20000));
OAI21X1 g116027(.A0 (n_32802), .A1 (n_16939), .B0 (n_18815), .Y(n_20004));
NAND2X1 g116031(.A (n_17579), .B (n_18814), .Y (n_19994));
INVX1 g116036(.A (n_18812), .Y (n_18813));
INVX1 g116039(.A (n_18810), .Y (n_18811));
NAND2X1 g116044(.A (n_17523), .B (n_18809), .Y (n_19979));
INVX1 g116053(.A (n_18807), .Y (n_18808));
INVX1 g116062(.A (n_18805), .Y (n_18806));
AOI21X1 g116065(.A0 (n_17364), .A1 (n_18682), .B0 (n_17357), .Y(n_19321));
INVX1 g116066(.A (n_18803), .Y (n_18804));
INVX1 g116071(.A (n_18801), .Y (n_18802));
INVX1 g116075(.A (n_18799), .Y (n_18800));
OR2X1 g116088(.A (n_17551), .B (n_17607), .Y (n_18798));
NAND2X1 g116111(.A (n_17040), .B (n_35310), .Y (n_19318));
INVX1 g116116(.A (n_18794), .Y (n_18795));
INVX1 g116131(.A (n_18169), .Y (n_19316));
NAND2X1 g116134(.A (n_17518), .B (n_17021), .Y (n_19314));
NAND2X1 g116135(.A (n_17517), .B (n_16612), .Y (n_20612));
OAI21X1 g116140(.A0 (n_17570), .A1 (n_18792), .B0 (n_18735), .Y(n_18793));
INVX1 g116147(.A (n_18790), .Y (n_18791));
OAI21X1 g116150(.A0 (n_17366), .A1 (n_16252), .B0 (n_18687), .Y(n_19312));
NAND2X1 g116157(.A (n_17509), .B (n_17504), .Y (n_19988));
NAND3X1 g116167(.A (n_11258), .B (n_16547), .C (n_16873), .Y(n_18789));
INVX1 g116168(.A (n_18787), .Y (n_18788));
INVX1 g116194(.A (n_19423), .Y (n_18786));
AND2X1 g116213(.A (n_16616), .B (n_18782), .Y (n_18784));
NOR2X1 g116219(.A (n_10021), .B (n_17929), .Y (n_18781));
NAND2X1 g116223(.A (n_18778), .B (n_19827), .Y (n_18779));
NOR2X1 g116252(.A (n_17937), .B (n_17742), .Y (n_19300));
INVX1 g116256(.A (n_18775), .Y (n_18776));
NOR2X1 g116260(.A (n_18774), .B (n_32873), .Y (n_20509));
NAND2X1 g116262(.A (n_34110), .B (n_34107), .Y (n_19298));
AND2X1 g116267(.A (n_18773), .B (n_18772), .Y (n_19945));
NOR2X1 g116268(.A (n_34843), .B (n_17415), .Y (n_20946));
AND2X1 g116270(.A (n_18771), .B (n_18772), .Y (n_20488));
AND2X1 g116271(.A (n_18771), .B (n_20264), .Y (n_19942));
NAND2X1 g116273(.A (n_21694), .B (n_18768), .Y (n_18770));
NAND2X1 g116276(.A (n_18768), .B (n_9431), .Y (n_18769));
AND2X1 g116277(.A (n_18981), .B (n_20264), .Y (n_21787));
NAND2X1 g116283(.A (n_9629), .B (n_17307), .Y (n_18767));
NAND2X2 g116285(.A (n_16445), .B (n_18765), .Y (n_18766));
NAND2X1 g116286(.A (n_9629), .B (n_17297), .Y (n_18764));
NAND2X1 g116290(.A (n_18760), .B (n_8303), .Y (n_18763));
NAND2X1 g116292(.A (n_9629), .B (n_18760), .Y (n_18761));
INVX1 g116314(.A (n_18758), .Y (n_18759));
INVX1 g116317(.A (n_18757), .Y (n_19931));
NAND2X1 g116325(.A (n_9629), .B (n_18754), .Y (n_18756));
NAND2X1 g116327(.A (n_18754), .B (n_8303), .Y (n_18755));
NAND2X1 g116341(.A (n_17972), .B (n_19235), .Y (n_18753));
NAND2X1 g116343(.A (n_34112), .B (n_35912), .Y (n_19287));
NAND2X1 g116344(.A (n_10754), .B (n_19709), .Y (n_18751));
NAND2X1 g116349(.A (n_21694), .B (n_18746), .Y (n_18750));
OR2X1 g116350(.A (n_18748), .B (n_14261), .Y (n_18749));
NAND2X1 g116351(.A (n_18746), .B (n_9431), .Y (n_18747));
NAND2X1 g116355(.A (n_18743), .B (n_9431), .Y (n_18745));
NAND2X1 g116357(.A (n_33803), .B (n_18743), .Y (n_18744));
OR2X1 g116360(.A (n_10023), .B (n_17303), .Y (n_18742));
NOR2X1 g116368(.A (n_16910), .B (n_16914), .Y (n_19284));
NAND2X1 g116372(.A (n_17955), .B (n_18645), .Y (n_18739));
OR2X1 g116373(.A (n_32382), .B (n_19256), .Y (n_18738));
NAND2X1 g116376(.A (n_17961), .B (n_16986), .Y (n_32979));
AND2X1 g116379(.A (n_18736), .B (n_18735), .Y (n_18737));
OR2X1 g116380(.A (n_10023), .B (n_17302), .Y (n_18734));
OR2X1 g116386(.A (n_10023), .B (n_17301), .Y (n_18730));
NAND2X1 g116387(.A (n_9629), .B (n_17295), .Y (n_18729));
NAND2X1 g116392(.A (n_9629), .B (n_18726), .Y (n_18728));
NAND2X1 g116396(.A (n_18726), .B (n_8303), .Y (n_18727));
NOR2X1 g116414(.A (n_17374), .B (n_17927), .Y (n_20408));
NAND2X1 g116434(.A (n_18691), .B (n_18765), .Y (n_19280));
NOR2X1 g116435(.A (n_32862), .B (n_16975), .Y (n_18724));
NOR2X1 g116450(.A (n_18774), .B (n_18721), .Y (n_19277));
NAND2X1 g116458(.A (n_9629), .B (n_17309), .Y (n_18720));
NAND2X1 g116460(.A (n_16598), .B (n_18717), .Y (n_22142));
NAND2X1 g116461(.A (n_9629), .B (n_17308), .Y (n_18716));
AND2X1 g116464(.A (n_18782), .B (n_18715), .Y (n_19271));
NAND2X1 g116470(.A (n_16927), .B (n_17271), .Y (n_20487));
NAND2X1 g116471(.A (n_9629), .B (n_18655), .Y (n_18714));
NAND2X1 g116474(.A (n_18685), .B (n_18710), .Y (n_18713));
OR2X1 g116476(.A (n_19279), .B (n_19792), .Y (n_20545));
NAND2X1 g116479(.A (n_19210), .B (n_17447), .Y (n_18712));
NAND2X1 g116483(.A (n_18711), .B (n_18710), .Y (n_19268));
NAND2X1 g116488(.A (n_18708), .B (n_18709), .Y (n_19962));
INVX1 g116489(.A (n_18115), .Y (n_20461));
NAND2X2 g116494(.A (n_19709), .B (n_16973), .Y (n_20458));
OR2X1 g116495(.A (n_18705), .B (n_18704), .Y (n_18706));
INVX1 g116502(.A (n_18703), .Y (n_19264));
NAND2X1 g116508(.A (n_21528), .B (n_17604), .Y (n_18702));
INVX1 g116509(.A (n_18700), .Y (n_18701));
INVX1 g116520(.A (n_18696), .Y (n_18697));
INVX1 g116525(.A (n_18107), .Y (n_19897));
NAND2X1 g116530(.A (n_17978), .B (n_35912), .Y (n_19880));
NAND2X1 g116538(.A (n_19827), .B (n_19208), .Y (n_19262));
NOR2X1 g116542(.A (n_18695), .B (n_17982), .Y (n_19260));
INVX1 g116545(.A (n_19821), .Y (n_18694));
AND2X1 g116548(.A (n_35310), .B (n_34065), .Y (n_19820));
INVX1 g116554(.A (n_18103), .Y (n_19892));
NAND2X1 g116561(.A (n_17897), .B (n_18676), .Y (n_18692));
NAND2X1 g116574(.A (n_18690), .B (n_18151), .Y (n_23892));
INVX1 g116575(.A (n_24173), .Y (n_18689));
OR2X1 g116578(.A (n_16917), .B (n_16916), .Y (n_24137));
NAND2X1 g116579(.A (n_16915), .B (n_18687), .Y (n_20969));
NAND2X1 g116584(.A (n_18705), .B (n_19331), .Y (n_19783));
NAND2X1 g116589(.A (n_16589), .B (n_17067), .Y (n_21398));
NAND2X1 g116590(.A (n_18685), .B (n_18684), .Y (n_20832));
NAND2X1 g116594(.A (n_19320), .B (n_18683), .Y (n_22194));
NAND2X1 g116597(.A (n_17358), .B (n_18682), .Y (n_22195));
INVX1 g116600(.A (n_18095), .Y (n_19894));
NAND2X1 g116606(.A (n_18681), .B (n_18680), .Y (n_21388));
NAND2X1 g116610(.A (n_18641), .B (n_16972), .Y (n_18679));
NAND2X1 g116615(.A (n_18677), .B (n_18676), .Y (n_25284));
INVX1 g116623(.A (n_18092), .Y (n_19893));
NAND2X1 g116626(.A (n_16586), .B (n_35950), .Y (n_23296));
NOR2X1 g116661(.A (n_17902), .B (n_16835), .Y (n_19890));
INVX1 g116668(.A (n_18674), .Y (n_18675));
INVX1 g116695(.A (n_18671), .Y (n_19934));
INVX1 g116707(.A (n_19364), .Y (n_18670));
INVX1 g116711(.A (n_18073), .Y (n_20485));
NAND2X1 g116717(.A (n_17370), .B (n_18668), .Y (n_18669));
NAND2X1 g116719(.A (n_18668), .B (n_18667), .Y (n_19233));
OR2X1 g116721(.A (n_17249), .B (n_18681), .Y (n_18666));
INVX1 g116723(.A (n_18070), .Y (n_20407));
NAND2X1 g116748(.A (n_18661), .B (n_9431), .Y (n_18663));
NAND2X1 g116749(.A (n_21333), .B (n_18661), .Y (n_18662));
AND2X1 g116757(.A (n_16767), .B (n_18680), .Y (n_20998));
NAND2X1 g116762(.A (n_18668), .B (n_18717), .Y (n_19873));
INVX1 g116764(.A (n_18660), .Y (n_19875));
INVX1 g116767(.A (n_18658), .Y (n_18659));
NAND2X1 g116771(.A (n_18655), .B (n_8303), .Y (n_18656));
NAND2X1 g116784(.A (n_17926), .B (n_18652), .Y (n_18653));
NAND3X1 g116795(.A (n_18145), .B (n_16505), .C (n_16821), .Y(n_19217));
NOR2X1 g116805(.A (n_16798), .B (n_17439), .Y (n_18650));
NAND2X1 g116819(.A (n_18645), .B (n_18644), .Y (n_23693));
NAND2X1 g116830(.A (n_17448), .B (n_35361), .Y (n_18643));
NAND2X1 g116839(.A (n_18641), .B (n_16785), .Y (n_18642));
NOR2X1 g116842(.A (n_18639), .B (n_17024), .Y (n_18640));
AND2X1 g116847(.A (n_18638), .B (n_18597), .Y (n_19203));
NOR2X1 g116853(.A (n_18637), .B (n_18633), .Y (n_19200));
INVX1 g116860(.A (n_18636), .Y (n_19196));
NOR2X1 g116863(.A (n_17264), .B (n_17263), .Y (n_19784));
INVX1 g116866(.A (n_18634), .Y (n_18635));
NOR2X1 g116873(.A (n_17315), .B (n_18633), .Y (n_35355));
NAND2X1 g116875(.A (n_18632), .B (n_18631), .Y (n_19193));
INVX1 g116877(.A (n_34677), .Y (n_18628));
NAND2X1 g116882(.A (n_19331), .B (n_18704), .Y (n_18627));
NAND2X2 g116885(.A (n_18626), .B (n_18069), .Y (n_19191));
NAND2X1 g116886(.A (n_9629), .B (n_17286), .Y (n_18625));
NAND2X1 g116888(.A (n_9629), .B (n_17285), .Y (n_32094));
NAND2X1 g116889(.A (n_9629), .B (n_17283), .Y (n_18623));
NAND2X1 g116891(.A (n_20304), .B (n_17280), .Y (n_18622));
NOR2X1 g116906(.A (n_18620), .B (n_35361), .Y (n_18621));
NAND2X1 g116909(.A (n_16930), .B (n_16611), .Y (n_18619));
NAND2X1 g116912(.A (n_17419), .B (n_22954), .Y (n_18618));
NAND2X1 g116919(.A (n_17412), .B (n_24840), .Y (n_18617));
NOR2X1 g116935(.A (n_18615), .B (n_18614), .Y (n_18616));
NAND2X1 g116938(.A (n_17405), .B (n_22953), .Y (n_18613));
NAND2X1 g116940(.A (n_17403), .B (n_24839), .Y (n_18612));
CLKBUFX1 gbuf_d_379(.A(n_17279), .Y(d_out_379));
CLKBUFX1 gbuf_q_379(.A(q_in_379), .Y(P1_IR[26]));
NAND2X1 g116943(.A (n_17400), .B (n_25693), .Y (n_18611));
NAND2X1 g116945(.A (n_17397), .B (n_25345), .Y (n_18610));
INVX1 g116949(.A (n_18608), .Y (n_18609));
NAND2X1 g116960(.A (n_17389), .B (n_22960), .Y (n_18607));
NAND2X1 g116961(.A (n_17388), .B (n_23648), .Y (n_18606));
NAND2X1 g116963(.A (n_17387), .B (n_24843), .Y (n_18605));
INVX1 g116970(.A (n_18604), .Y (n_19868));
NOR2X1 g116986(.A (n_18602), .B (n_18601), .Y (n_18603));
NOR2X1 g116987(.A (n_18599), .B (n_17872), .Y (n_18600));
NAND3X1 g116989(.A (n_17688), .B (n_11533), .C (n_16797), .Y(n_20621));
NOR2X1 g116993(.A (n_20763), .B (n_18597), .Y (n_35381));
NOR2X1 g116995(.A (n_19167), .B (n_20763), .Y (n_20372));
NAND2X1 g116997(.A (n_17342), .B (n_22952), .Y (n_18596));
NAND2X1 g116998(.A (n_17339), .B (n_24837), .Y (n_18595));
INVX1 g117023(.A (n_18593), .Y (n_18594));
NAND2X1 g117037(.A (n_17430), .B (n_22027), .Y (n_19858));
NAND2X1 g117039(.A (n_17427), .B (n_23666), .Y (n_19856));
NAND2X1 g117044(.A (n_17414), .B (n_23643), .Y (n_18592));
NAND2X1 g117048(.A (n_17404), .B (n_23641), .Y (n_18591));
NAND2X1 g117055(.A (n_17341), .B (n_23638), .Y (n_18590));
NAND2X1 g117060(.A (n_17429), .B (n_25925), .Y (n_19864));
NOR2X1 g117063(.A (n_17426), .B (n_13936), .Y (n_19155));
NOR2X1 g117065(.A (n_17425), .B (n_13898), .Y (n_19153));
NAND2X1 g117073(.A (n_17428), .B (n_26493), .Y (n_19841));
NAND2X1 g117081(.A (n_17431), .B (n_25148), .Y (n_19151));
NAND2X1 g117083(.A (n_17432), .B (n_25793), .Y (n_19149));
NAND2X1 g117101(.A (n_17463), .B (n_23718), .Y (n_19838));
NAND2X1 g117103(.A (n_17461), .B (n_22024), .Y (n_19147));
INVX1 g117105(.A (n_18588), .Y (n_18589));
NAND2X1 g117109(.A (n_17450), .B (n_26074), .Y (n_19848));
INVX1 g117110(.A (n_19884), .Y (n_18587));
INVX1 g117130(.A (n_18586), .Y (n_19144));
NAND2X1 g117135(.A (n_17458), .B (n_25838), .Y (n_19851));
INVX1 g117147(.A (n_18030), .Y (n_19142));
AOI21X1 g117152(.A0 (n_18584), .A1 (n_35686), .B0 (n_18583), .Y(n_18585));
NAND2X1 g117157(.A (n_17464), .B (n_23635), .Y (n_19138));
NAND2X1 g117161(.A (n_17465), .B (n_22012), .Y (n_19136));
NAND2X1 g117163(.A (n_17331), .B (n_21601), .Y (n_19860));
INVX1 g117165(.A (n_18581), .Y (n_18582));
NAND2X1 g117169(.A (n_17452), .B (n_26514), .Y (n_19881));
NAND2X1 g117174(.A (n_17455), .B (n_25847), .Y (n_19886));
AOI21X1 g117205(.A0 (n_18580), .A1 (n_35000), .B0 (n_17207), .Y(n_19133));
NAND2X1 g117207(.A (n_17325), .B (n_18018), .Y (n_19131));
NAND2X1 g117209(.A (n_17328), .B (n_16231), .Y (n_19129));
INVX1 g117234(.A (n_18578), .Y (n_18579));
NAND2X1 g117237(.A (n_17433), .B (n_21622), .Y (n_19122));
INVX1 g117238(.A (n_18576), .Y (n_18577));
NAND2X1 g117248(.A (n_17424), .B (n_21600), .Y (n_19120));
INVX1 g117249(.A (n_18574), .Y (n_18575));
AOI21X1 g117252(.A0 (n_16209), .A1 (n_7988), .B0 (n_9013), .Y(n_18573));
NAND2X1 g117263(.A (n_17318), .B (n_16510), .Y (n_18572));
NAND2X1 g117267(.A (n_17322), .B (n_18012), .Y (n_19115));
AOI22X1 g117288(.A0 (n_17399), .A1 (n_8946), .B0 (n_20218), .B1(n_7724), .Y (n_18569));
AOI22X1 g117293(.A0 (n_16486), .A1 (n_8946), .B0 (n_20218), .B1(n_10566), .Y (n_18568));
AOI22X1 g117296(.A0 (n_16465), .A1 (n_8946), .B0 (n_20218), .B1(n_10854), .Y (n_18567));
AOI22X1 g117298(.A0 (n_17909), .A1 (n_33004), .B0 (n_17337), .B1(n_17908), .Y (n_18565));
AOI22X1 g117309(.A0 (n_16202), .A1 (n_7988), .B0 (n_11138), .B1(n_13711), .Y (n_18564));
NOR2X1 g117322(.A (n_16998), .B (n_17453), .Y (n_18563));
AOI22X1 g117325(.A0 (n_32349), .A1 (n_18561), .B0 (n_11498), .B1(n_18560), .Y (n_18562));
NAND2X1 g117348(.A (n_35816), .B (n_17993), .Y (n_18559));
NAND2X1 g117349(.A (n_35736), .B (n_32984), .Y (n_18557));
NAND2X1 g117356(.A (n_18262), .B (n_18532), .Y (n_18554));
NAND2X1 g117381(.A (n_17968), .B (n_17993), .Y (n_18553));
NAND2X1 g117448(.A (n_35776), .B (n_17997), .Y (n_18550));
NAND2X1 g117449(.A (n_18546), .B (n_32984), .Y (n_18547));
NAND2X1 g117453(.A (n_35776), .B (n_18005), .Y (n_18545));
NAND2X1 g117459(.A (n_18546), .B (n_18005), .Y (n_18543));
NAND2X1 g117460(.A (n_18546), .B (n_17997), .Y (n_18542));
NOR2X1 g117468(.A (n_11058), .B (n_20188), .Y (n_19668));
NOR2X1 g117554(.A (n_18536), .B (n_23190), .Y (n_19665));
INVX1 g117579(.A (n_17950), .Y (n_19703));
INVX1 g117584(.A (n_18535), .Y (n_20781));
NAND2X1 g117602(.A (n_18533), .B (n_18532), .Y (n_18534));
NOR2X1 g117605(.A (n_35600), .B (n_17731), .Y (n_18531));
NAND2X1 g117609(.A (n_22021), .B (n_32984), .Y (n_18530));
NAND2X1 g117620(.A (n_22021), .B (n_17997), .Y (n_18529));
NOR2X1 g117621(.A (n_17665), .B (n_19071), .Y (n_18527));
NAND2X1 g117625(.A (n_18533), .B (n_18005), .Y (n_18526));
NAND2X1 g117634(.A (n_18533), .B (n_17993), .Y (n_18524));
NAND2X1 g117635(.A (n_35479), .B (n_18532), .Y (n_18523));
INVX1 g117644(.A (n_18521), .Y (n_19767));
NAND2X1 g117648(.A (n_18038), .B (n_16958), .Y (n_19093));
INVX1 g117649(.A (n_18519), .Y (n_18520));
NOR2X1 g117658(.A (n_18518), .B (n_18517), .Y (n_21555));
OR2X1 g117662(.A (n_18518), .B (n_18917), .Y (n_18516));
INVX1 g117663(.A (n_20299), .Y (n_18515));
NAND2X1 g117675(.A (n_18511), .B (n_24101), .Y (n_18512));
NOR2X1 g117694(.A (n_16172), .B (n_19000), .Y (n_21385));
NOR2X1 g117704(.A (n_11468), .B (n_34998), .Y (n_18509));
INVX1 g117719(.A (n_18506), .Y (n_18507));
INVX1 g117728(.A (n_18504), .Y (n_18505));
NAND2X1 g117762(.A (n_34385), .B (n_33551), .Y (n_20261));
INVX1 g117764(.A (n_18500), .Y (n_18501));
NAND2X1 g117775(.A (n_18511), .B (n_18498), .Y (n_18499));
INVX1 g117841(.A (n_19786), .Y (n_19077));
INVX1 g117879(.A (n_20332), .Y (n_18497));
AND2X1 g117890(.A (n_18496), .B (n_33551), .Y (n_19075));
NAND2X1 g117897(.A (n_18511), .B (n_13268), .Y (n_18495));
NAND2X1 g117906(.A (n_17252), .B (n_17182), .Y (n_18493));
NOR2X1 g117911(.A (n_19629), .B (n_19631), .Y (n_18492));
NOR2X1 g117933(.A (n_19626), .B (n_23190), .Y (n_19774));
NAND2X1 g117955(.A (n_17255), .B (n_35318), .Y (n_18487));
INVX1 g117992(.A (n_18486), .Y (n_19736));
INVX1 g118070(.A (n_19247), .Y (n_18479));
NAND2X2 g118084(.A (n_11226), .B (n_17776), .Y (n_20341));
INVX1 g118088(.A (n_18478), .Y (n_19729));
INVX1 g118101(.A (n_34996), .Y (n_20338));
NAND2X1 g118104(.A (n_34991), .B (n_18360), .Y (n_20254));
NAND2X1 g118122(.A (n_18475), .B (n_17775), .Y (n_19689));
INVX2 g118130(.A (n_18474), .Y (n_19695));
INVX1 g118133(.A (n_34995), .Y (n_20342));
NAND2X1 g118144(.A (n_18709), .B (n_17232), .Y (n_19063));
NOR2X1 g118147(.A (n_20916), .B (n_17235), .Y (n_20412));
INVX1 g118151(.A (n_18470), .Y (n_18471));
INVX1 g118157(.A (n_19723), .Y (n_18467));
NAND2X1 g118186(.A (n_17219), .B (n_19669), .Y (n_20931));
NOR2X1 g118196(.A (n_20175), .B (n_17639), .Y (n_18465));
NAND2X1 g118200(.A (n_18511), .B (n_22080), .Y (n_18464));
INVX1 g118252(.A (n_18460), .Y (n_18461));
NAND2X1 g118263(.A (n_16517), .B (n_35173), .Y (n_19055));
INVX1 g118274(.A (n_18458), .Y (n_18459));
AND2X1 g118276(.A (n_18457), .B (n_18456), .Y (n_20797));
NAND2X1 g118334(.A (n_17810), .B (n_16499), .Y (n_18455));
INVX1 g118338(.A (n_18454), .Y (n_19763));
INVX1 g118388(.A (n_18449), .Y (n_18450));
INVX1 g118392(.A (n_20325), .Y (n_18448));
INVX1 g118396(.A (n_20322), .Y (n_18447));
NOR2X1 g118401(.A (n_19135), .B (n_32836), .Y (n_20241));
NAND2X1 g118403(.A (n_16497), .B (n_16499), .Y (n_21742));
INVX1 g118404(.A (n_20327), .Y (n_18444));
NAND3X1 g118408(.A (n_16734), .B (n_16779), .C (n_16735), .Y(n_18443));
OAI21X1 g118415(.A0 (n_16518), .A1 (n_18441), .B0 (n_23046), .Y(n_18442));
OAI21X1 g118417(.A0 (n_16457), .A1 (n_17678), .B0 (n_17188), .Y(n_18440));
INVX1 g118423(.A (n_17862), .Y (n_18439));
OAI21X1 g118432(.A0 (n_18437), .A1 (n_19183), .B0 (n_17818), .Y(n_18438));
AOI21X1 g118435(.A0 (n_33051), .A1 (n_18435), .B0 (n_17784), .Y(n_19041));
AOI21X1 g118437(.A0 (n_18434), .A1 (n_18433), .B0 (n_17788), .Y(n_19039));
OAI21X1 g118447(.A0 (n_16518), .A1 (n_17856), .B0 (n_23043), .Y(n_18432));
OAI21X1 g118451(.A0 (n_16518), .A1 (n_18429), .B0 (n_23041), .Y(n_18430));
OAI21X1 g118462(.A0 (n_16743), .A1 (n_17766), .B0 (n_18428), .Y(n_19032));
OAI21X1 g118469(.A0 (n_18426), .A1 (n_17866), .B0 (n_18353), .Y(n_18427));
INVX1 g118472(.A (n_18424), .Y (n_18425));
OAI21X1 g118481(.A0 (n_17860), .A1 (n_17165), .B0 (n_18421), .Y(n_20467));
OAI21X1 g118483(.A0 (n_17786), .A1 (n_16425), .B0 (n_35949), .Y(n_19029));
AND2X1 g118486(.A (n_17234), .B (n_18638), .Y (n_19027));
AOI21X1 g118487(.A0 (n_17158), .A1 (n_17221), .B0 (n_17841), .Y(n_20356));
INVX1 g118488(.A (n_18419), .Y (n_18420));
AOI21X1 g118490(.A0 (n_16445), .A1 (n_32959), .B0 (n_16742), .Y(n_20355));
INVX1 g118491(.A (n_18417), .Y (n_18418));
OAI21X1 g118511(.A0 (n_16417), .A1 (n_32698), .B0 (n_24896), .Y(n_18416));
OAI21X1 g118520(.A0 (n_18145), .A1 (n_32748), .B0 (n_24005), .Y(n_18414));
OAI21X1 g118539(.A0 (n_16760), .A1 (n_16430), .B0 (n_17735), .Y(n_19008));
AOI21X1 g118542(.A0 (n_16764), .A1 (n_19186), .B0 (n_17692), .Y(n_20493));
NAND2X1 g118560(.A (n_17204), .B (n_16430), .Y (n_20316));
AOI21X1 g118564(.A0 (n_32428), .A1 (n_18909), .B0 (n_10030), .Y(n_18408));
AOI22X1 g118579(.A0 (n_11791), .A1 (n_17117), .B0 (n_11797), .B1(n_18145), .Y (n_18407));
AOI22X1 g118583(.A0 (n_17814), .A1 (n_18909), .B0 (n_18289), .B1(n_8185), .Y (n_18406));
AOI22X1 g118588(.A0 (n_19766), .A1 (n_18909), .B0 (n_18289), .B1(n_8458), .Y (n_18405));
OAI21X1 g118591(.A0 (n_8325), .A1 (n_2379), .B0 (n_17220), .Y(n_18403));
INVX1 g118612(.A (n_18401), .Y (n_18402));
NAND2X1 g118717(.A (n_18387), .B (n_18399), .Y (n_18400));
INVX1 g118726(.A (n_18397), .Y (n_19758));
NOR2X1 g118728(.A (n_18395), .B (n_18373), .Y (n_18396));
INVX1 g118730(.A (n_19091), .Y (n_18394));
NAND2X1 g118751(.A (n_16728), .B (n_17719), .Y (n_18391));
NAND2X1 g118757(.A (n_18379), .B (n_18384), .Y (n_18390));
NAND2X1 g118761(.A (n_18561), .B (n_18384), .Y (n_18389));
NAND2X1 g118766(.A (n_18387), .B (n_23270), .Y (n_18388));
NAND2X1 g118781(.A (n_16728), .B (n_18384), .Y (n_18386));
NAND2X1 g118788(.A (n_18561), .B (n_32739), .Y (n_18383));
NAND2X1 g118817(.A (n_18379), .B (n_18378), .Y (n_18380));
NAND2X1 g118819(.A (n_17647), .B (n_18375), .Y (n_18377));
NAND2X1 g118823(.A (n_18387), .B (n_18375), .Y (n_18376));
INVX1 g118826(.A (n_23226), .Y (n_18374));
NAND2X1 g118836(.A (n_16728), .B (n_18378), .Y (n_18372));
CLKBUFX1 g118856(.A (n_17251), .Y (n_19637));
NAND2X1 g118881(.A (n_18379), .B (n_17719), .Y (n_18368));
INVX1 g118893(.A (n_18362), .Y (n_18987));
INVX1 g118907(.A (n_18360), .Y (n_20195));
INVX1 g118945(.A (n_19065), .Y (n_18356));
AND2X1 g119041(.A (n_18773), .B (n_18355), .Y (n_21302));
INVX1 g119050(.A (n_18354), .Y (n_18982));
NAND2X1 g119099(.A (n_18353), .B (n_17226), .Y (n_18978));
NAND2X1 g119103(.A (n_16444), .B (n_35399), .Y (n_18976));
INVX1 g119110(.A (n_18351), .Y (n_18352));
INVX1 g119114(.A (n_18348), .Y (n_18349));
INVX1 g119116(.A (n_18346), .Y (n_18347));
INVX1 g119122(.A (n_23225), .Y (n_18345));
NAND2X1 g119147(.A (n_18561), .B (n_22786), .Y (n_18342));
NAND2X1 g119183(.A (n_18561), .B (n_18340), .Y (n_18341));
NAND2X1 g119189(.A (n_18379), .B (n_10848), .Y (n_18339));
AND2X1 g119191(.A (n_18561), .B (n_10848), .Y (n_18338));
NAND2X1 g119193(.A (n_18387), .B (n_10848), .Y (n_18337));
NAND2X1 g119196(.A (n_16728), .B (n_10848), .Y (n_18336));
INVX1 g119197(.A (n_18334), .Y (n_18335));
INVX1 g119201(.A (n_18332), .Y (n_18333));
INVX1 g119204(.A (n_18330), .Y (n_18331));
INVX1 g119206(.A (n_18328), .Y (n_18329));
NAND2X1 g119212(.A (n_18667), .B (n_35896), .Y (n_18968));
NAND2X1 g119214(.A (n_16773), .B (n_16820), .Y (n_20212));
INVX1 g119221(.A (n_18325), .Y (n_18965));
NOR2X1 g119223(.A (n_20102), .B (n_17657), .Y (n_21299));
AND2X1 g119224(.A (n_17652), .B (n_18324), .Y (n_22576));
INVX1 g119271(.A (n_18322), .Y (n_18323));
NOR2X1 g119278(.A (n_18321), .B (n_18320), .Y (n_18960));
INVX1 g119284(.A (n_19048), .Y (n_18319));
OAI21X1 g119388(.A0 (n_16126), .A1 (n_14261), .B0 (n_13175), .Y(n_18317));
OR2X1 g119392(.A (n_17743), .B (n_17206), .Y (n_18316));
OAI21X1 g119432(.A0 (n_14279), .A1 (n_17172), .B0 (n_18310), .Y(n_18311));
OAI21X1 g119440(.A0 (n_13843), .A1 (n_17172), .B0 (n_13646), .Y(n_18309));
AOI21X1 g119441(.A0 (n_32777), .A1 (n_18288), .B0 (n_15352), .Y(n_18307));
INVX2 g119522(.A (n_17732), .Y (n_19647));
INVX1 g119537(.A (n_16800), .Y (n_18306));
NAND2X1 g119553(.A (n_17175), .B (n_18303), .Y (n_18304));
OAI21X1 g119557(.A0 (n_17293), .A1 (n_16126), .B0 (n_27716), .Y(n_18302));
OAI21X1 g119566(.A0 (n_14430), .A1 (n_16126), .B0 (n_24299), .Y(n_18300));
AOI21X1 g119568(.A0 (n_26631), .A1 (n_16172), .B0 (n_13866), .Y(n_18298));
NAND2X1 g119571(.A (n_17143), .B (n_21293), .Y (n_18296));
AOI21X1 g119575(.A0 (n_18294), .A1 (n_16172), .B0 (n_13485), .Y(n_18295));
NAND2X1 g119620(.A (n_17128), .B (n_27707), .Y (n_18942));
OAI21X1 g119623(.A0 (n_35555), .A1 (n_16738), .B0 (n_27711), .Y(n_19571));
NAND2X1 g119650(.A (n_17142), .B (n_27686), .Y (n_19564));
NAND2X1 g119653(.A (n_17145), .B (n_29662), .Y (n_19561));
NAND2X1 g119658(.A (n_17138), .B (n_29690), .Y (n_18940));
NAND2X1 g119663(.A (n_17168), .B (n_27756), .Y (n_19558));
NAND2X1 g119664(.A (n_17140), .B (n_33731), .Y (n_19555));
NAND2X1 g119665(.A (n_17164), .B (n_27681), .Y (n_19552));
AOI21X1 g119670(.A0 (n_11333), .A1 (n_17133), .B0 (n_17177), .Y(n_18291));
NAND2X1 g119675(.A (n_17129), .B (n_27685), .Y (n_18937));
AOI22X1 g119684(.A0 (n_18289), .A1 (n_10612), .B0 (n_18288), .B1(n_18909), .Y (n_18290));
AOI22X1 g119700(.A0 (n_10573), .A1 (n_13173), .B0 (n_17712), .B1(n_8946), .Y (n_18287));
AOI21X1 g119701(.A0 (n_11988), .A1 (n_16407), .B0 (n_17149), .Y(n_18285));
OAI22X1 g119707(.A0 (n_9520), .A1 (n_10116), .B0 (n_17131), .B1(n_8309), .Y (n_18284));
OAI22X1 g119709(.A0 (n_9520), .A1 (n_10114), .B0 (n_16738), .B1(n_8309), .Y (n_18283));
NAND2X1 g119736(.A (n_27747), .B (n_16740), .Y (n_18281));
NAND2X1 g119743(.A (n_26530), .B (n_18948), .Y (n_18279));
NOR2X1 g119748(.A (n_17715), .B (n_19474), .Y (n_19524));
NAND2X1 g119765(.A (n_21919), .B (n_18275), .Y (n_18276));
NAND2X1 g119766(.A (n_14439), .B (n_16130), .Y (n_18274));
NAND2X1 g119770(.A (n_25297), .B (n_18948), .Y (n_18272));
NAND2X1 g119778(.A (n_16740), .B (n_25554), .Y (n_18271));
NAND2X1 g119783(.A (n_16400), .B (n_21919), .Y (n_18270));
NAND2X1 g119886(.A (n_26637), .B (n_18275), .Y (n_18268));
INVX1 g119911(.A (n_17740), .Y (n_21733));
OR2X1 g119920(.A (n_9722), .B (n_19471), .Y (n_20103));
NAND2X1 g119960(.A (n_18275), .B (n_27770), .Y (n_18265));
NAND2X1 g119963(.A (n_17340), .B (n_16740), .Y (n_18264));
NAND2X1 g119967(.A (n_18262), .B (n_17133), .Y (n_18263));
NAND2X1 g119975(.A (n_18262), .B (n_17178), .Y (n_18261));
NAND2X1 g119982(.A (n_35736), .B (n_17133), .Y (n_18260));
NAND2X1 g119983(.A (n_35794), .B (n_17178), .Y (n_18258));
INVX1 g119987(.A (n_18255), .Y (n_18256));
NAND2X1 g119992(.A (n_17674), .B (n_18275), .Y (n_18254));
NAND2X1 g119999(.A (n_14439), .B (n_17139), .Y (n_18253));
NAND2X1 g120011(.A (n_18533), .B (n_17178), .Y (n_18252));
NAND2X1 g120012(.A (n_18533), .B (n_17133), .Y (n_18251));
NAND2X1 g120013(.A (n_22021), .B (n_17139), .Y (n_18250));
NAND2X1 g120033(.A (n_16396), .B (n_8946), .Y (n_18249));
INVX1 g114243(.A (n_18237), .Y (n_19458));
NAND2X1 g114335(.A (n_17635), .B (n_18907), .Y (n_18236));
NAND3X1 g114408(.A (n_16701), .B (n_17335), .C (n_18041), .Y(n_20057));
NAND2X1 g115003(.A (n_18833), .B (n_18894), .Y (n_18898));
NAND2X1 g115172(.A (n_17090), .B (n_17596), .Y (n_19441));
NOR3X1 g115223(.A (n_16621), .B (n_16650), .C (n_17617), .Y(n_20044));
NAND3X1 g115226(.A (n_17615), .B (n_18235), .C (n_17614), .Y(n_18868));
AOI21X1 g115254(.A0 (n_17623), .A1 (n_32786), .B0 (n_14298), .Y(n_18234));
OR2X1 g115317(.A (n_16665), .B (n_18231), .Y (n_18232));
NOR2X1 g115321(.A (n_18184), .B (n_18164), .Y (n_18230));
NAND3X1 g115336(.A (n_16582), .B (n_16580), .C (n_17298), .Y(n_18229));
NAND2X1 g115338(.A (n_18198), .B (n_18227), .Y (n_18228));
NAND2X1 g115339(.A (n_18219), .B (n_18227), .Y (n_18226));
NAND2X1 g115412(.A (n_21703), .B (n_18190), .Y (n_18225));
NAND2X1 g115422(.A (n_21703), .B (n_17491), .Y (n_18224));
NAND2X1 g115457(.A (n_20112), .B (n_18203), .Y (n_18223));
NOR2X1 g115512(.A (n_17564), .B (n_19375), .Y (n_20552));
NAND2X1 g115522(.A (n_20864), .B (n_18205), .Y (n_18222));
NAND2X1 g115612(.A (n_20112), .B (n_18208), .Y (n_18221));
NAND2X1 g115617(.A (n_18546), .B (n_18189), .Y (n_19411));
NAND2X1 g115618(.A (n_18219), .B (n_18218), .Y (n_18220));
NAND2X1 g115619(.A (n_18219), .B (n_21328), .Y (n_18217));
NOR2X1 g115624(.A (n_34062), .B (n_17085), .Y (n_20550));
NOR2X1 g115625(.A (n_16388), .B (n_17086), .Y (n_20031));
NOR2X1 g115641(.A (n_17534), .B (n_35346), .Y (n_18844));
NOR2X1 g115650(.A (n_17035), .B (n_16671), .Y (n_20652));
NOR2X1 g115716(.A (n_10021), .B (n_18213), .Y (n_18214));
NAND2X1 g115723(.A (n_20864), .B (n_17501), .Y (n_18212));
NAND2X1 g115746(.A (n_18196), .B (n_21328), .Y (n_18211));
NAND2X1 g115747(.A (n_18208), .B (n_21328), .Y (n_18209));
NAND2X1 g115758(.A (n_18201), .B (n_21328), .Y (n_18207));
NAND2X1 g115761(.A (n_18205), .B (n_21328), .Y (n_18206));
NAND2X1 g115773(.A (n_18203), .B (n_21328), .Y (n_18204));
NAND2X1 g115794(.A (n_20864), .B (n_18201), .Y (n_18202));
NAND2X1 g115807(.A (n_17010), .B (n_17008), .Y (n_18200));
NAND2X1 g115818(.A (n_18198), .B (n_30505), .Y (n_18199));
NAND2X1 g115836(.A (n_20864), .B (n_18196), .Y (n_18197));
NAND2X1 g115841(.A (n_18194), .B (n_18144), .Y (n_18195));
NAND3X1 g115844(.A (n_17018), .B (n_18192), .C (n_17017), .Y(n_18193));
NAND2X1 g115854(.A (n_18190), .B (n_21328), .Y (n_18191));
NAND2X1 g115905(.A (n_35479), .B (n_18189), .Y (n_19409));
NAND2X1 g115906(.A (n_26234), .B (n_18189), .Y (n_18188));
INVX1 g115936(.A (n_18186), .Y (n_18187));
INVX1 g115947(.A (n_18185), .Y (n_18826));
NAND2X1 g115960(.A (n_16688), .B (n_18184), .Y (n_19987));
INVX1 g115962(.A (n_18183), .Y (n_18819));
CLKBUFX1 g115968(.A (n_18182), .Y (n_19437));
NOR2X1 g115972(.A (n_18180), .B (n_17555), .Y (n_18181));
AOI21X1 g115975(.A0 (n_16363), .A1 (n_18071), .B0 (n_16370), .Y(n_18179));
INVX2 g116019(.A (n_17602), .Y (n_19407));
INVX1 g116021(.A (n_34641), .Y (n_18178));
INVX1 g116037(.A (n_18176), .Y (n_18812));
NAND2X2 g116040(.A (n_17046), .B (n_16922), .Y (n_18810));
OAI21X1 g116054(.A0 (n_16295), .A1 (n_16907), .B0 (n_15924), .Y(n_18807));
OAI21X1 g116063(.A0 (n_16914), .A1 (n_18687), .B0 (n_16912), .Y(n_18805));
NAND2X1 g116067(.A (n_17066), .B (n_17549), .Y (n_18803));
AOI21X1 g116068(.A0 (n_16901), .A1 (n_35950), .B0 (n_18127), .Y(n_20028));
NAND2X1 g116072(.A (n_17062), .B (n_16292), .Y (n_18801));
AOI21X1 g116076(.A0 (n_16900), .A1 (n_18685), .B0 (n_17360), .Y(n_18799));
CLKBUFX1 g116094(.A (n_18878), .Y (n_20018));
INVX1 g116096(.A (n_18173), .Y (n_18174));
INVX1 g116104(.A (n_18171), .Y (n_18172));
NAND2X2 g116107(.A (n_17047), .B (n_16699), .Y (n_35357));
NAND2X1 g116108(.A (n_17034), .B (n_15926), .Y (n_19405));
OAI21X1 g116109(.A0 (n_18104), .A1 (n_18161), .B0 (n_16090), .Y(n_19414));
OAI21X1 g116117(.A0 (n_16916), .A1 (n_18170), .B0 (n_16918), .Y(n_18794));
CLKBUFX1 g116126(.A (n_18888), .Y (n_21507));
NAND2X1 g116129(.A (n_17072), .B (n_17512), .Y (n_20023));
NAND2X1 g116132(.A (n_17071), .B (n_17515), .Y (n_18169));
AND2X1 g116148(.A (n_16667), .B (n_17507), .Y (n_18790));
OAI21X1 g116158(.A0 (n_16612), .A1 (n_18166), .B0 (n_16930), .Y(n_18168));
AOI21X1 g116160(.A0 (n_18164), .A1 (n_18163), .B0 (n_16776), .Y(n_18165));
NAND2X1 g116165(.A (n_17054), .B (n_17569), .Y (n_18162));
NAND2X1 g116169(.A (n_17052), .B (n_18161), .Y (n_18787));
AOI21X1 g116172(.A0 (n_18159), .A1 (n_16872), .B0 (n_16424), .Y(n_18160));
INVX1 g116191(.A (n_18891), .Y (n_18158));
OAI21X1 g116193(.A0 (n_18157), .A1 (n_19974), .B0 (n_17020), .Y(n_19432));
INVX1 g116257(.A (n_18156), .Y (n_18775));
NOR2X1 g116279(.A (n_18897), .B (n_11534), .Y (n_18155));
NAND2X1 g116291(.A (n_18142), .B (n_18918), .Y (n_18154));
INVX1 g116307(.A (n_18153), .Y (n_19937));
NAND2X1 g116309(.A (n_18151), .B (n_16917), .Y (n_18152));
NOR2X1 g116312(.A (n_18149), .B (n_16423), .Y (n_18150));
NOR2X1 g116313(.A (n_18146), .B (n_10765), .Y (n_18147));
NAND3X1 g116315(.A (n_18145), .B (n_16273), .C (n_18057), .Y(n_18758));
NAND2X1 g116318(.A (n_18144), .B (n_19213), .Y (n_18757));
NAND2X1 g116326(.A (n_18142), .B (n_32739), .Y (n_18143));
INVX1 g116339(.A (n_18139), .Y (n_19377));
NAND2X1 g116345(.A (n_18137), .B (n_18135), .Y (n_18138));
NAND2X1 g116348(.A (n_18135), .B (n_14235), .Y (n_18136));
INVX1 g116352(.A (n_34552), .Y (n_18134));
INVX1 g116361(.A (n_18857), .Y (n_18131));
INVX1 g116365(.A (n_17582), .Y (n_19372));
INVX1 g116370(.A (n_17581), .Y (n_19373));
NAND2X1 g116374(.A (n_17067), .B (n_17361), .Y (n_18130));
NAND2X1 g116377(.A (n_16902), .B (n_18093), .Y (n_18129));
NAND2X1 g116378(.A (n_18127), .B (n_17073), .Y (n_18128));
INVX1 g116383(.A (n_17580), .Y (n_18732));
NAND2X1 g116389(.A (n_17570), .B (n_18735), .Y (n_19923));
NAND2X1 g116393(.A (n_18142), .B (n_21185), .Y (n_18126));
INVX1 g116402(.A (n_18125), .Y (n_19370));
INVX1 g116405(.A (n_19371), .Y (n_18124));
NAND2X1 g116423(.A (n_17369), .B (n_18101), .Y (n_18122));
INVX1 g116428(.A (n_17571), .Y (n_19367));
INVX1 g116430(.A (n_18120), .Y (n_18121));
INVX1 g116442(.A (n_18118), .Y (n_18722));
NAND2X1 g116444(.A (n_16626), .B (n_16351), .Y (n_20465));
NAND2X1 g116445(.A (n_21528), .B (n_16975), .Y (n_18117));
NAND2X1 g116490(.A (n_18683), .B (n_18711), .Y (n_18115));
NOR2X1 g116491(.A (n_16870), .B (n_16400), .Y (n_18114));
NAND2X1 g116503(.A (n_18106), .B (n_18683), .Y (n_18703));
INVX1 g116504(.A (n_18112), .Y (n_18113));
NAND2X1 g116507(.A (n_17442), .B (n_19210), .Y (n_18110));
NAND2X1 g116511(.A (n_32862), .B (n_21528), .Y (n_18700));
INVX1 g116514(.A (n_17561), .Y (n_18698));
NAND2X1 g116521(.A (n_17441), .B (n_17603), .Y (n_18696));
NAND2X1 g116522(.A (n_18108), .B (n_16423), .Y (n_19334));
NAND2X1 g116526(.A (n_19242), .B (n_18106), .Y (n_18107));
NAND2X1 g116540(.A (n_34109), .B (n_19304), .Y (n_35410));
NOR2X1 g116546(.A (n_16602), .B (n_18104), .Y (n_19821));
NAND2X1 g116555(.A (n_19242), .B (n_18676), .Y (n_18103));
NAND2X1 g116576(.A (n_18102), .B (n_18101), .Y (n_24173));
NAND2X1 g116586(.A (n_18099), .B (n_15923), .Y (n_18100));
NOR2X1 g116591(.A (n_18097), .B (n_18096), .Y (n_18098));
NAND2X1 g116601(.A (n_19245), .B (n_18676), .Y (n_18095));
NAND2X1 g116621(.A (n_16301), .B (n_18093), .Y (n_23476));
NAND2X1 g116624(.A (n_19245), .B (n_18091), .Y (n_18092));
NAND2X1 g116628(.A (n_16292), .B (n_17064), .Y (n_24177));
NAND2X1 g116630(.A (n_18099), .B (n_18088), .Y (n_18089));
INVX1 g116647(.A (n_18834), .Y (n_18087));
INVX1 g116651(.A (n_18085), .Y (n_18086));
NAND2X1 g116669(.A (n_21047), .B (n_16655), .Y (n_18674));
INVX1 g116680(.A (n_34066), .Y (n_18083));
INVX1 g116689(.A (n_18080), .Y (n_18672));
INVX1 g116691(.A (n_18849), .Y (n_18079));
NAND2X1 g116696(.A (n_18151), .B (n_16591), .Y (n_18671));
INVX1 g116697(.A (n_18848), .Y (n_18078));
NOR2X1 g116701(.A (n_16275), .B (n_17344), .Y (n_18077));
NAND2X1 g116708(.A (n_18074), .B (n_18652), .Y (n_19364));
NAND2X1 g116712(.A (n_18652), .B (n_18717), .Y (n_18073));
INVX2 g116714(.A (n_17529), .Y (n_19874));
NAND2X1 g116716(.A (n_15936), .B (n_18071), .Y (n_18072));
NAND2X1 g116724(.A (n_16771), .B (n_18069), .Y (n_18070));
NAND4X1 g116725(.A (n_16543), .B (n_11051), .C (n_16237), .D(n_15904), .Y (n_18068));
NOR2X1 g116742(.A (n_34744), .B (n_16887), .Y (n_20011));
NAND2X1 g116746(.A (n_18065), .B (n_18135), .Y (n_18066));
NAND2X1 g116756(.A (n_35309), .B (n_17057), .Y (n_18064));
NAND2X1 g116763(.A (n_18142), .B (n_26530), .Y (n_18063));
NAND2X1 g116765(.A (n_18062), .B (n_18061), .Y (n_18660));
NAND2X2 g116769(.A (n_18060), .B (n_32878), .Y (n_18658));
NOR2X1 g116775(.A (n_16573), .B (n_16571), .Y (n_20532));
NOR2X1 g116779(.A (n_16885), .B (n_17028), .Y (n_20010));
NOR2X1 g116781(.A (n_16281), .B (n_16338), .Y (n_18059));
NAND3X1 g116785(.A (n_18145), .B (n_16837), .C (n_18057), .Y(n_18900));
NOR2X1 g116786(.A (n_16278), .B (n_16328), .Y (n_19932));
INVX1 g116787(.A (n_18055), .Y (n_18056));
INVX1 g116807(.A (n_18052), .Y (n_18648));
INVX1 g116811(.A (n_18050), .Y (n_18051));
INVX1 g116814(.A (n_18049), .Y (n_18646));
NOR2X1 g116841(.A (n_16358), .B (n_16989), .Y (n_18048));
NOR2X1 g116845(.A (n_16629), .B (n_18792), .Y (n_18047));
AND2X1 g116850(.A (n_17390), .B (n_16438), .Y (n_21482));
NAND2X2 g116861(.A (n_18046), .B (n_18632), .Y (n_18636));
NAND2X1 g116867(.A (n_18046), .B (n_18060), .Y (n_18634));
INVX1 g116900(.A (n_18045), .Y (n_19368));
NOR2X1 g116905(.A (n_16610), .B (n_33982), .Y (n_18044));
NOR2X1 g116910(.A (n_17080), .B (n_16621), .Y (n_18043));
NOR2X1 g116950(.A (n_16966), .B (n_13942), .Y (n_18608));
OAI21X1 g116971(.A0 (n_12437), .A1 (n_16381), .B0 (n_16599), .Y(n_18604));
AOI21X1 g116984(.A0 (n_32864), .A1 (n_16517), .B0 (n_35171), .Y(n_18042));
NAND3X1 g116999(.A (n_17630), .B (n_17284), .C (n_18041), .Y(n_19388));
NOR2X1 g117024(.A (n_16965), .B (n_13897), .Y (n_18593));
INVX1 g117099(.A (n_18039), .Y (n_18040));
NAND2X1 g117106(.A (n_16959), .B (n_18038), .Y (n_18588));
NAND2X2 g117111(.A (n_16894), .B (n_16517), .Y (n_19884));
INVX1 g117118(.A (n_18035), .Y (n_18036));
NAND2X1 g117122(.A (n_16897), .B (n_18560), .Y (n_20431));
NAND2X2 g117131(.A (n_16893), .B (n_32411), .Y (n_18586));
INVX1 g117142(.A (n_18033), .Y (n_18034));
INVX1 g117144(.A (n_18031), .Y (n_18032));
OAI21X1 g117148(.A0 (n_16849), .A1 (n_18709), .B0 (n_16238), .Y(n_18030));
NAND2X1 g117155(.A (n_16880), .B (n_23935), .Y (n_19361));
NOR2X1 g117166(.A (n_16881), .B (n_13928), .Y (n_18581));
INVX1 g117167(.A (n_18028), .Y (n_18029));
AOI22X1 g117211(.A0 (n_17409), .A1 (n_8946), .B0 (n_10573), .B1(n_7737), .Y (n_18025));
AOI21X1 g117218(.A0 (n_17418), .A1 (n_8946), .B0 (n_10543), .Y(n_18024));
AOI22X1 g117219(.A0 (n_17411), .A1 (n_8946), .B0 (n_10573), .B1(n_7546), .Y (n_18023));
AOI22X1 g117228(.A0 (n_35206), .A1 (n_18001), .B0 (n_32984), .B1(n_18000), .Y (n_18021));
AOI22X1 g117229(.A0 (n_10699), .A1 (n_10314), .B0 (n_32496), .B1(n_17997), .Y (n_18020));
AOI21X1 g117230(.A0 (n_16209), .A1 (n_17993), .B0 (n_11264), .Y(n_18019));
OAI21X1 g117235(.A0 (n_18018), .A1 (n_16538), .B0 (n_16539), .Y(n_18578));
NAND2X1 g117239(.A (n_16967), .B (n_23904), .Y (n_18576));
NAND2X1 g117250(.A (n_16963), .B (n_23932), .Y (n_18574));
NAND2X1 g117255(.A (n_16945), .B (n_17013), .Y (n_19354));
INVX1 g117256(.A (n_18016), .Y (n_18017));
AOI21X1 g117264(.A0 (n_16643), .A1 (n_19108), .B0 (n_9506), .Y(n_18015));
AOI21X1 g117265(.A0 (n_17004), .A1 (n_7988), .B0 (n_9020), .Y(n_18013));
AOI21X1 g117271(.A0 (n_10316), .A1 (n_18005), .B0 (n_16062), .Y(n_18011));
AOI22X1 g117278(.A0 (n_17413), .A1 (n_8946), .B0 (n_10573), .B1(n_13167), .Y (n_18010));
AOI22X1 g117286(.A0 (n_10333), .A1 (n_16799), .B0 (n_16331), .B1(n_16196), .Y (n_18009));
AOI22X1 g117287(.A0 (n_16576), .A1 (n_7988), .B0 (n_11138), .B1(P3_reg3[2] ), .Y (n_18008));
AOI22X1 g117294(.A0 (n_17451), .A1 (n_19108), .B0 (n_11138), .B1(n_13375), .Y (n_18007));
AOI21X1 g117304(.A0 (n_16857), .A1 (n_18005), .B0 (n_11043), .Y(n_18006));
AOI22X1 g117305(.A0 (n_35206), .A1 (n_32984), .B0 (n_18001), .B1(n_18000), .Y (n_18004));
AOI22X1 g117306(.A0 (n_10699), .A1 (n_17997), .B0 (n_10314), .B1(n_32496), .Y (n_17999));
AOI22X1 g117307(.A0 (n_10315), .A1 (n_17993), .B0 (n_11036), .B1(n_16209), .Y (n_17994));
AOI22X1 g117312(.A0 (n_32496), .A1 (n_19108), .B0 (n_11138), .B1(n_13378), .Y (n_17991));
AOI21X1 g117318(.A0 (n_10485), .A1 (n_18833), .B0 (n_16637), .Y(n_17990));
AOI21X1 g117319(.A0 (n_11092), .A1 (n_16616), .B0 (n_16980), .Y(n_17989));
XOR2X1 g117330(.A (n_19172), .B (n_17289), .Y (n_19423));
AOI21X1 g117333(.A0 (n_16895), .A1 (n_16505), .B0 (n_17236), .Y(n_20436));
NAND2X1 g117351(.A (n_17968), .B (n_16209), .Y (n_17987));
NAND2X1 g117352(.A (n_35776), .B (n_17970), .Y (n_17986));
INVX1 g117358(.A (n_17982), .Y (n_17983));
NAND2X1 g117373(.A (n_35776), .B (n_16202), .Y (n_17980));
INVX1 g117424(.A (n_17978), .Y (n_19259));
OR2X1 g117427(.A (n_35861), .B (n_17975), .Y (n_17977));
INVX1 g117430(.A (n_17973), .Y (n_19876));
INVX1 g117431(.A (n_17973), .Y (n_17974));
INVX2 g117433(.A (n_17972), .Y (n_19305));
NAND2X1 g117451(.A (n_18546), .B (n_17970), .Y (n_17971));
NAND2X1 g117458(.A (n_17968), .B (n_16202), .Y (n_17969));
NAND2X1 g117461(.A (n_35776), .B (n_16209), .Y (n_17967));
INVX1 g117477(.A (n_19706), .Y (n_18541));
INVX2 g117505(.A (n_17963), .Y (n_22340));
INVX1 g117508(.A (n_17961), .Y (n_17962));
NAND2X1 g117512(.A (n_10755), .B (n_33968), .Y (n_20586));
INVX1 g117546(.A (n_16975), .Y (n_19903));
NAND2X1 g117556(.A (n_17955), .B (n_16031), .Y (n_17956));
NAND2X1 g117580(.A (n_17351), .B (n_16477), .Y (n_17950));
INVX1 g117585(.A (n_18641), .Y (n_18535));
NAND2X1 g117597(.A (n_22021), .B (n_16209), .Y (n_17948));
NOR2X1 g117604(.A (n_35602), .B (n_17473), .Y (n_17947));
NOR2X1 g117606(.A (n_35596), .B (n_16474), .Y (n_17945));
NAND2X1 g117616(.A (n_16481), .B (n_8946), .Y (n_17944));
NAND2X1 g117624(.A (n_18533), .B (n_16202), .Y (n_17943));
NOR2X1 g117626(.A (n_35596), .B (n_32992), .Y (n_17942));
NOR2X1 g117630(.A (n_35529), .B (n_16473), .Y (n_17940));
NAND2X1 g117631(.A (n_35576), .B (n_17970), .Y (n_17939));
NAND2X1 g117632(.A (n_17970), .B (n_7988), .Y (n_17938));
NAND2X1 g117645(.A (n_16249), .B (n_17242), .Y (n_18521));
NOR2X1 g117650(.A (n_17922), .B (n_18517), .Y (n_18519));
INVX1 g117659(.A (n_17937), .Y (n_19383));
OR2X1 g117665(.A (n_17894), .B (n_34998), .Y (n_20299));
NAND2X1 g117703(.A (n_17399), .B (n_17713), .Y (n_17935));
INVX1 g117716(.A (n_17932), .Y (n_17933));
NAND2X1 g117720(.A (n_16858), .B (n_23996), .Y (n_18506));
INVX1 g117729(.A (n_17931), .Y (n_18504));
INVX1 g117743(.A (n_17929), .Y (n_17930));
NAND2X1 g117765(.A (n_16830), .B (n_17928), .Y (n_18500));
INVX1 g117769(.A (n_17927), .Y (n_19255));
INVX1 g117778(.A (n_18765), .Y (n_17925));
OR2X1 g117803(.A (n_17923), .B (n_17922), .Y (n_19768));
INVX1 g117818(.A (n_17920), .Y (n_17921));
AND2X1 g117826(.A (n_17918), .B (n_17923), .Y (n_17919));
NAND2X1 g117834(.A (n_17399), .B (n_19595), .Y (n_17917));
NAND2X2 g117842(.A (n_19647), .B (n_17916), .Y (n_19786));
NAND2X1 g117875(.A (n_16353), .B (n_35686), .Y (n_19905));
NAND2X1 g117878(.A (n_17203), .B (n_16808), .Y (n_20928));
CLKBUFX1 g117880(.A (n_18597), .Y (n_20332));
INVX2 g117883(.A (n_17391), .Y (n_19169));
NAND2X1 g117886(.A (n_17399), .B (n_23356), .Y (n_17915));
INVX2 g117916(.A (n_17912), .Y (n_19228));
NAND2X1 g117930(.A (n_17908), .B (n_17909), .Y (n_22369));
NAND2X1 g117932(.A (n_32992), .B (n_16203), .Y (n_17907));
NAND2X1 g117987(.A (n_17906), .B (n_17251), .Y (n_19788));
INVX1 g117993(.A (n_17371), .Y (n_18486));
INVX1 g118035(.A (n_18626), .Y (n_17904));
INVX1 g118052(.A (n_17903), .Y (n_18484));
INVX1 g118055(.A (n_18710), .Y (n_18482));
OR2X1 g118065(.A (n_17392), .B (n_19523), .Y (n_19799));
INVX1 g118067(.A (n_17902), .Y (n_18480));
AND2X1 g118071(.A (n_17380), .B (n_33550), .Y (n_19247));
INVX1 g118072(.A (n_17901), .Y (n_19294));
INVX1 g118075(.A (n_18680), .Y (n_17900));
INVX1 g118080(.A (n_17897), .Y (n_19243));
INVX1 g118085(.A (n_18677), .Y (n_17896));
INVX1 g118089(.A (n_17352), .Y (n_18478));
INVX1 g118093(.A (n_17895), .Y (n_18476));
NAND2X1 g118131(.A (n_17348), .B (n_17894), .Y (n_18474));
AND2X1 g118140(.A (n_19891), .B (n_19238), .Y (n_23029));
AND2X1 g118145(.A (n_17892), .B (n_19236), .Y (n_23659));
INVX1 g118152(.A (n_18772), .Y (n_18470));
INVX1 g118155(.A (n_18771), .Y (n_18468));
NAND2X1 g118158(.A (n_34991), .B (n_34998), .Y (n_19723));
INVX1 g118193(.A (n_17889), .Y (n_19212));
NAND2X1 g118211(.A (n_18532), .B (n_17975), .Y (n_17888));
NAND2X1 g118213(.A (n_16819), .B (n_24042), .Y (n_19220));
INVX1 g118227(.A (n_17886), .Y (n_17887));
NOR2X1 g118253(.A (n_17885), .B (n_17884), .Y (n_18460));
INVX1 g118258(.A (n_17882), .Y (n_17883));
NOR2X1 g118261(.A (n_17885), .B (n_17923), .Y (n_19955));
INVX1 g118267(.A (n_18721), .Y (n_17881));
NAND2X1 g118275(.A (n_18560), .B (n_16848), .Y (n_18458));
INVX1 g118332(.A (n_18637), .Y (n_17880));
INVX1 g118335(.A (n_17329), .Y (n_19302));
NAND2X1 g118337(.A (n_17223), .B (n_17878), .Y (n_17879));
NAND2X1 g118339(.A (n_32838), .B (n_17878), .Y (n_18454));
INVX1 g118354(.A (n_18633), .Y (n_17876));
INVX1 g118385(.A (n_17872), .Y (n_17873));
NAND2X1 g118389(.A (n_16844), .B (n_17482), .Y (n_18449));
NAND2X1 g118393(.A (n_17317), .B (n_16510), .Y (n_20325));
INVX1 g118394(.A (n_20324), .Y (n_17871));
NAND2X1 g118397(.A (n_16539), .B (n_16265), .Y (n_20322));
INVX1 g118398(.A (n_20323), .Y (n_17870));
NAND2X1 g118405(.A (n_16231), .B (n_34741), .Y (n_20327));
INVX1 g118406(.A (n_20328), .Y (n_17868));
AOI21X1 g118419(.A0 (n_16178), .A1 (n_18353), .B0 (n_17866), .Y(n_17867));
AOI21X1 g118420(.A0 (n_17864), .A1 (n_19225), .B0 (n_17863), .Y(n_17865));
AOI21X1 g118424(.A0 (n_18421), .A1 (n_17861), .B0 (n_17860), .Y(n_17862));
NAND2X1 g118431(.A (n_16818), .B (n_24002), .Y (n_19214));
AOI21X1 g118438(.A0 (n_17233), .A1 (n_17240), .B0 (n_17250), .Y(n_20360));
OAI21X1 g118444(.A0 (n_17630), .A1 (n_18441), .B0 (n_21548), .Y(n_17859));
OAI21X1 g118445(.A0 (n_17630), .A1 (n_17856), .B0 (n_21551), .Y(n_17858));
NAND2X1 g118446(.A (n_16866), .B (n_22016), .Y (n_17855));
OAI21X1 g118449(.A0 (n_17630), .A1 (n_18429), .B0 (n_21550), .Y(n_17854));
NAND2X1 g118450(.A (n_16862), .B (n_22015), .Y (n_17853));
AND2X1 g118455(.A (n_16861), .B (n_23039), .Y (n_17852));
NAND2X1 g118457(.A (n_16831), .B (n_14089), .Y (n_17851));
OAI21X1 g118459(.A0 (n_32417), .A1 (n_17848), .B0 (n_21609), .Y(n_17849));
OAI21X1 g118471(.A0 (n_17847), .A1 (n_16765), .B0 (n_17846), .Y(n_19239));
OAI21X1 g118473(.A0 (n_17846), .A1 (n_16841), .B0 (n_17300), .Y(n_18424));
INVX1 g118474(.A (n_17844), .Y (n_17845));
OAI21X1 g118484(.A0 (n_18969), .A1 (n_18433), .B0 (n_18434), .Y(n_17842));
AOI21X1 g118489(.A0 (n_17841), .A1 (n_17253), .B0 (n_32959), .Y(n_18419));
OAI21X1 g118492(.A0 (n_16786), .A1 (n_35896), .B0 (n_16773), .Y(n_18417));
OAI21X1 g118543(.A0 (n_32417), .A1 (n_19024), .B0 (n_21604), .Y(n_17839));
AOI22X1 g118549(.A0 (n_15943), .A1 (n_8946), .B0 (n_20218), .B1(n_11135), .Y (n_17837));
OAI21X1 g118550(.A0 (n_32417), .A1 (n_32698), .B0 (n_21602), .Y(n_17836));
AOI22X1 g118551(.A0 (n_16552), .A1 (n_18909), .B0 (n_18289), .B1(n_10562), .Y (n_17835));
INVX1 g118555(.A (n_18748), .Y (n_18410));
INVX1 g118573(.A (n_17274), .Y (n_17833));
AOI22X1 g118575(.A0 (n_16829), .A1 (n_17831), .B0 (n_35244), .B1(n_17830), .Y (n_17832));
AOI21X1 g118600(.A0 (n_9720), .A1 (n_16728), .B0 (n_16840), .Y(n_17829));
AOI21X1 g118601(.A0 (n_16728), .A1 (n_18997), .B0 (n_11274), .Y(n_17828));
NOR2X1 g118604(.A (n_16838), .B (n_11485), .Y (n_17827));
NOR2X1 g118605(.A (n_16833), .B (n_16834), .Y (n_17826));
NOR2X1 g118725(.A (n_17822), .B (n_20301), .Y (n_21153));
NAND2X1 g118727(.A (n_17820), .B (n_34721), .Y (n_18397));
NAND2X1 g118731(.A (n_18773), .B (n_17820), .Y (n_19091));
NAND2X1 g118745(.A (n_17818), .B (n_16792), .Y (n_26415));
INVX1 g118747(.A (n_17257), .Y (n_19060));
NAND2X1 g118752(.A (n_17800), .B (n_18384), .Y (n_17817));
NAND2X1 g118753(.A (n_17798), .B (n_20050), .Y (n_17816));
NAND2X1 g118756(.A (n_17814), .B (n_20050), .Y (n_17815));
NAND2X1 g118758(.A (n_18353), .B (n_17866), .Y (n_17813));
NAND2X1 g118759(.A (n_17794), .B (n_20050), .Y (n_17812));
NAND2X1 g118770(.A (n_17814), .B (n_25309), .Y (n_17809));
NOR2X1 g118777(.A (n_32349), .B (n_18561), .Y (n_17808));
NAND2X1 g118782(.A (n_18426), .B (n_18353), .Y (n_19043));
NAND2X1 g118787(.A (n_17794), .B (n_32794), .Y (n_17806));
OR2X1 g118796(.A (n_33051), .B (n_17803), .Y (n_17804));
INVX1 g118797(.A (n_18518), .Y (n_17802));
NAND2X1 g118809(.A (n_17800), .B (n_18378), .Y (n_17801));
NAND2X1 g118810(.A (n_17798), .B (n_17797), .Y (n_17799));
NAND2X1 g118811(.A (n_17814), .B (n_24984), .Y (n_17796));
NAND2X1 g118818(.A (n_17794), .B (n_17797), .Y (n_17795));
NOR2X1 g118822(.A (n_11254), .B (n_17125), .Y (n_17793));
NAND2X1 g118827(.A (n_18428), .B (n_34720), .Y (n_23226));
INVX1 g118841(.A (n_20744), .Y (n_18371));
INVX1 g118863(.A (n_17788), .Y (n_17789));
NAND2X1 g118869(.A (n_17233), .B (n_17786), .Y (n_17787));
NAND2X1 g118875(.A (n_33051), .B (n_17763), .Y (n_17785));
NAND2X1 g118879(.A (n_17864), .B (n_17161), .Y (n_17783));
INVX1 g118883(.A (n_17782), .Y (n_18365));
INVX1 g118885(.A (n_21390), .Y (n_17781));
INVX1 g118887(.A (n_19651), .Y (n_17780));
NAND2X1 g118894(.A (n_17846), .B (n_16845), .Y (n_18362));
NOR2X1 g118895(.A (n_18437), .B (n_17777), .Y (n_17778));
INVX1 g118909(.A (n_34998), .Y (n_18360));
INVX2 g118917(.A (n_17775), .Y (n_21344));
INVX1 g118933(.A (n_17772), .Y (n_17773));
AND2X1 g118946(.A (n_16785), .B (n_16843), .Y (n_19065));
NAND2X1 g119039(.A (n_18561), .B (n_19766), .Y (n_17770));
NAND2X1 g119051(.A (n_17767), .B (n_17766), .Y (n_18354));
AND2X1 g119089(.A (n_17818), .B (n_17777), .Y (n_17765));
NOR2X1 g119106(.A (n_17763), .B (n_18353), .Y (n_17764));
NOR2X1 g119112(.A (n_18435), .B (n_17803), .Y (n_18351));
OAI22X1 g119115(.A0 (n_9198), .A1 (n_17678), .B0 (n_16435), .B1(n_17186), .Y (n_18348));
NAND2X1 g119117(.A (n_18061), .B (n_18426), .Y (n_18346));
NAND2X1 g119123(.A (n_18395), .B (n_34721), .Y (n_23225));
INVX1 g119135(.A (n_20175), .Y (n_18344));
INVX1 g119142(.A (n_17760), .Y (n_19061));
INVX1 g119155(.A (n_17759), .Y (n_19079));
NAND2X1 g119167(.A (n_17800), .B (n_17719), .Y (n_17758));
NAND2X1 g119181(.A (n_17794), .B (n_25309), .Y (n_17755));
AND2X1 g119186(.A (n_17794), .B (n_18909), .Y (n_17754));
AND2X1 g119187(.A (n_17800), .B (n_10848), .Y (n_17752));
AND2X1 g119188(.A (n_17798), .B (n_18909), .Y (n_17750));
OAI22X1 g119198(.A0 (n_16174), .A1 (n_17639), .B0 (n_11730), .B1(n_16173), .Y (n_18334));
NAND2X1 g119202(.A (n_18434), .B (n_16843), .Y (n_18332));
NAND2X1 g119205(.A (n_21748), .B (n_16164), .Y (n_18330));
NAND2X1 g119207(.A (n_16448), .B (n_18638), .Y (n_18328));
INVX1 g119215(.A (n_20211), .Y (n_17748));
INVX1 g119218(.A (n_17747), .Y (n_18326));
OR2X1 g119222(.A (n_32382), .B (n_17745), .Y (n_18325));
NAND2X1 g119272(.A (n_17743), .B (n_16166), .Y (n_18322));
INVX1 g119275(.A (n_17742), .Y (n_19049));
INVX1 g119280(.A (n_35003), .Y (n_19047));
NOR2X1 g119285(.A (n_17740), .B (n_18320), .Y (n_19048));
INVX1 g119288(.A (n_19046), .Y (n_17739));
INVX1 g119336(.A (n_19626), .Y (n_19098));
AND2X1 g119390(.A (n_17735), .B (n_16168), .Y (n_19044));
INVX1 g119395(.A (n_19669), .Y (n_19624));
AOI21X1 g119561(.A0 (n_16777), .A1 (n_17727), .B0 (n_14319), .Y(n_17729));
AOI21X1 g119686(.A0 (n_16182), .A1 (n_16768), .B0 (n_16737), .Y(n_17725));
AOI22X1 g119692(.A0 (n_12992), .A1 (n_17130), .B0 (n_13071), .B1(n_17131), .Y (n_17724));
AOI21X1 g119693(.A0 (n_16768), .A1 (n_16173), .B0 (n_16741), .Y(n_17723));
NAND2X1 g119742(.A (n_18399), .B (n_18288), .Y (n_17721));
NAND2X1 g119746(.A (n_17719), .B (n_17715), .Y (n_17720));
AND2X1 g119760(.A (n_17968), .B (n_17678), .Y (n_17718));
NAND2X1 g119769(.A (n_15089), .B (n_18288), .Y (n_17717));
NAND2X1 g119771(.A (n_15089), .B (n_17715), .Y (n_17716));
NAND2X1 g119772(.A (n_17713), .B (n_17712), .Y (n_17714));
NAND2X1 g119774(.A (n_17713), .B (n_16172), .Y (n_17711));
NAND2X1 g119791(.A (n_32739), .B (n_17715), .Y (n_17709));
NOR2X1 g119797(.A (n_17172), .B (n_32770), .Y (n_17707));
NAND2X1 g119804(.A (n_18288), .B (n_23696), .Y (n_17706));
NAND2X1 g119807(.A (n_17715), .B (n_17797), .Y (n_17705));
NAND2X1 g119809(.A (n_17712), .B (n_35054), .Y (n_17704));
NAND2X1 g119811(.A (n_16172), .B (n_35054), .Y (n_17703));
NAND2X1 g119860(.A (n_17715), .B (n_18909), .Y (n_17698));
INVX1 g119917(.A (n_17692), .Y (n_19687));
NAND2X1 g119919(.A (n_19595), .B (n_17712), .Y (n_17691));
INVX1 g119940(.A (n_18355), .Y (n_17690));
INVX1 g119945(.A (n_17688), .Y (n_17689));
NAND2X1 g119949(.A (n_33750), .B (n_15962), .Y (n_17687));
NAND2X1 g119956(.A (n_12349), .B (n_16731), .Y (n_17686));
NAND2X1 g119958(.A (n_14439), .B (n_17682), .Y (n_17685));
NAND2X1 g119962(.A (n_14439), .B (n_17680), .Y (n_17684));
NAND2X1 g119974(.A (n_35790), .B (n_17682), .Y (n_17683));
NAND2X1 g119976(.A (n_35736), .B (n_17680), .Y (n_17681));
NAND2X1 g119978(.A (n_35822), .B (n_17678), .Y (n_17679));
NAND2X1 g119988(.A (n_16796), .B (n_20741), .Y (n_18255));
NAND2X1 g119995(.A (n_34609), .B (n_15852), .Y (n_17677));
NAND2X1 g119998(.A (n_17674), .B (n_17712), .Y (n_17675));
NOR2X1 g120003(.A (n_35596), .B (n_16402), .Y (n_17673));
NAND2X1 g120004(.A (n_35515), .B (n_17682), .Y (n_17672));
NAND2X1 g120007(.A (n_20133), .B (n_17682), .Y (n_17670));
NAND2X1 g120008(.A (n_20133), .B (n_17680), .Y (n_17669));
NAND2X1 g120009(.A (n_13311), .B (n_17678), .Y (n_17668));
NOR2X1 g120010(.A (n_17665), .B (n_16404), .Y (n_17666));
NOR2X1 g120014(.A (n_17665), .B (n_17131), .Y (n_17664));
NAND2X1 g120015(.A (n_17682), .B (n_7988), .Y (n_17662));
NAND2X1 g120016(.A (n_35508), .B (n_17680), .Y (n_17661));
NAND2X1 g120017(.A (n_17680), .B (n_7988), .Y (n_17660));
NAND2X1 g120018(.A (n_35540), .B (n_17678), .Y (n_17659));
NOR2X1 g120023(.A (n_17655), .B (n_17592), .Y (n_17656));
INVX1 g120024(.A (n_17652), .Y (n_17653));
NAND2X1 g120034(.A (n_16172), .B (n_8946), .Y (n_17649));
CLKBUFX1 gbuf_d_380(.A(n_16875), .Y(d_out_380));
CLKBUFX1 gbuf_q_380(.A(q_in_380), .Y(P3_IR[27]));
INVX1 g120141(.A (n_18387), .Y (n_17637));
XOR2X1 g114244(.A (n_32417), .B (n_16702), .Y (n_18237));
NAND2X1 g114304(.A (n_17635), .B (n_17719), .Y (n_17636));
NAND2X1 g114311(.A (n_17635), .B (n_18384), .Y (n_17634));
NAND2X1 g114321(.A (n_17635), .B (n_32777), .Y (n_17632));
XOR2X1 g118613(.A (n_8737), .B (n_17592), .Y (n_17631));
AND2X1 g118613_and(.A (n_8737), .B (n_17592), .Y (n_18401));
NAND3X1 g115192(.A (n_16544), .B (n_17628), .C (n_16225), .Y(n_21100));
NAND3X1 g115231(.A (n_17630), .B (n_32426), .C (n_17628), .Y(n_18896));
NAND3X1 g115319(.A (n_16321), .B (n_16369), .C (n_16319), .Y(n_17627));
NAND2X2 g115337(.A (n_17625), .B (n_35943), .Y (n_35258));
NAND2X1 g115354(.A (n_17623), .B (n_17719), .Y (n_17624));
NAND2X1 g115420(.A (n_17623), .B (n_24446), .Y (n_17622));
NAND2X1 g115490(.A (n_17623), .B (n_21185), .Y (n_17621));
INVX1 g115621(.A (n_17619), .Y (n_17620));
NAND2X1 g115623(.A (n_17059), .B (n_16653), .Y (n_19403));
NOR2X1 g115631(.A (n_16385), .B (n_17617), .Y (n_17618));
NAND3X1 g115633(.A (n_20033), .B (n_17615), .C (n_17614), .Y(n_17616));
NOR2X1 g115638(.A (n_17612), .B (n_17053), .Y (n_17613));
CLKBUFX1 gbuf_d_381(.A(n_16549), .Y(d_out_381));
CLKBUFX1 gbuf_q_381(.A(q_in_381), .Y(P1_IR[25]));
NAND2X1 g115834(.A (n_17610), .B (n_16572), .Y (n_17611));
NAND2X1 g115840(.A (n_17608), .B (n_17584), .Y (n_17609));
NAND2X1 g115937(.A (n_16676), .B (n_17026), .Y (n_18186));
OAI21X1 g115948(.A0 (n_17606), .A1 (n_17607), .B0 (n_17605), .Y(n_18185));
OAI21X1 g115952(.A0 (n_17603), .A1 (n_17604), .B0 (n_32862), .Y(n_18885));
NAND2X1 g115963(.A (n_16687), .B (n_34171), .Y (n_18183));
NAND2X1 g115969(.A (n_16686), .B (n_15936), .Y (n_18182));
OAI21X1 g115994(.A0 (n_16641), .A1 (n_32503), .B0 (n_17545), .Y(n_18873));
NAND3X1 g116020(.A (n_16694), .B (n_34546), .C (n_16693), .Y(n_17602));
NAND2X1 g116038(.A (n_16682), .B (n_32503), .Y (n_18176));
INVX1 g116069(.A (n_17598), .Y (n_17599));
NAND2X1 g116089(.A (n_16679), .B (n_16095), .Y (n_18871));
NAND2X1 g116095(.A (n_16680), .B (n_16325), .Y (n_18878));
AOI21X1 g116097(.A0 (n_17595), .A1 (n_16387), .B0 (n_17056), .Y(n_18173));
INVX1 g116101(.A (n_17596), .Y (n_17597));
NAND2X1 g116103(.A (n_16691), .B (n_17015), .Y (n_18875));
AOI21X1 g116105(.A0 (n_16607), .A1 (n_17614), .B0 (n_17595), .Y(n_18171));
NAND2X1 g116127(.A (n_15935), .B (n_32915), .Y (n_18888));
XOR2X1 g116192(.A (n_16042), .B (n_16341), .Y (n_18891));
AOI22X1 g116197(.A0 (n_17591), .A1 (n_17592), .B0 (n_8737), .B1(n_17591), .Y (n_19401));
NAND2X1 g116211(.A (n_16800), .B (n_19304), .Y (n_17590));
NOR2X1 g116214(.A (n_19085), .B (n_19279), .Y (n_17589));
NAND2X1 g116258(.A (n_35913), .B (n_18096), .Y (n_18156));
NAND2X1 g116289(.A (n_17578), .B (n_22792), .Y (n_17588));
INVX1 g116298(.A (n_17587), .Y (n_18846));
NAND2X1 g116308(.A (n_18074), .B (n_18101), .Y (n_18153));
NOR2X1 g116311(.A (n_16571), .B (n_34842), .Y (n_17586));
INVX1 g116334(.A (n_17077), .Y (n_18140));
NAND2X1 g116340(.A (n_18096), .B (n_17533), .Y (n_18139));
CLKBUFX1 gbuf_d_382(.A(n_16555), .Y(d_out_382));
CLKBUFX1 gbuf_q_382(.A(q_in_382), .Y(P2_IR[26]));
INVX1 g116358(.A (n_18189), .Y (n_17583));
INVX1 g116362(.A (n_17074), .Y (n_18857));
NAND2X1 g116366(.A (n_16587), .B (n_18093), .Y (n_17582));
NAND2X1 g116371(.A (n_17576), .B (n_18682), .Y (n_17581));
NAND2X1 g116384(.A (n_19827), .B (n_16972), .Y (n_17580));
NAND2X1 g116391(.A (n_17578), .B (n_18375), .Y (n_17579));
INVX1 g116403(.A (n_17069), .Y (n_18125));
NAND2X1 g116406(.A (n_16587), .B (n_17576), .Y (n_19371));
INVX1 g116408(.A (n_17068), .Y (n_19402));
INVX1 g116416(.A (n_17574), .Y (n_17573));
NAND2X1 g116429(.A (n_16099), .B (n_17570), .Y (n_17571));
NAND2X1 g116431(.A (n_17569), .B (n_32503), .Y (n_18120));
INVX1 g116437(.A (n_17065), .Y (n_18856));
NAND2X2 g116443(.A (n_17568), .B (n_18144), .Y (n_18118));
INVX1 g116454(.A (n_17564), .Y (n_17565));
INVX1 g116467(.A (n_17061), .Y (n_18852));
NAND2X1 g116469(.A (n_16978), .B (n_16632), .Y (n_17562));
NAND2X1 g116506(.A (n_18644), .B (n_19210), .Y (n_18112));
NAND2X1 g116515(.A (n_19208), .B (n_16986), .Y (n_17561));
NAND2X1 g116518(.A (n_16228), .B (n_16988), .Y (n_17560));
INVX1 g116528(.A (n_35345), .Y (n_17559));
NAND2X1 g116549(.A (n_17051), .B (n_18161), .Y (n_23089));
INVX1 g116550(.A (n_21502), .Y (n_17557));
NAND2X1 g116552(.A (n_17615), .B (n_16325), .Y (n_19958));
INVX1 g116556(.A (n_17555), .Y (n_17556));
NAND2X1 g116571(.A (n_16095), .B (n_16678), .Y (n_22638));
NAND2X1 g116572(.A (n_35915), .B (n_16386), .Y (n_22949));
NOR2X1 g116587(.A (n_17552), .B (n_17081), .Y (n_17553));
AND2X1 g116592(.A (n_35349), .B (n_17605), .Y (n_17551));
OR2X1 g116608(.A (n_18159), .B (n_16871), .Y (n_17550));
NAND2X1 g116620(.A (n_17549), .B (n_16587), .Y (n_23477));
NAND2X1 g116622(.A (n_15924), .B (n_17576), .Y (n_22361));
NAND2X1 g116648(.A (n_35632), .B (n_35221), .Y (n_18834));
NAND2X1 g116652(.A (n_17545), .B (n_17543), .Y (n_18085));
NAND2X2 g116666(.A (n_17569), .B (n_17543), .Y (n_18843));
NAND2X1 g116667(.A (n_35221), .B (n_16999), .Y (n_17542));
INVX1 g116671(.A (n_17539), .Y (n_17540));
INVX1 g116676(.A (n_17536), .Y (n_17537));
NAND2X1 g116686(.A (n_35352), .B (n_17534), .Y (n_17535));
NAND2X2 g116690(.A (n_35351), .B (n_17533), .Y (n_18080));
INVX1 g116692(.A (n_17039), .Y (n_18849));
NOR2X1 g116698(.A (n_16566), .B (n_16921), .Y (n_18848));
INVX1 g116699(.A (n_17532), .Y (n_19365));
NAND2X1 g116702(.A (n_18074), .B (n_16920), .Y (n_35700));
NAND2X1 g116715(.A (n_19304), .B (n_19235), .Y (n_17529));
NAND2X1 g116745(.A (n_17526), .B (n_17178), .Y (n_17527));
INVX1 g116753(.A (n_17524), .Y (n_17525));
INVX1 g116759(.A (n_17032), .Y (n_19413));
NAND2X1 g116770(.A (n_25309), .B (n_17578), .Y (n_17523));
NAND2X1 g116788(.A (n_17605), .B (n_17533), .Y (n_18055));
NOR2X1 g116791(.A (n_21395), .B (n_16892), .Y (n_19963));
NAND2X1 g116808(.A (n_17510), .B (n_16099), .Y (n_18052));
INVX1 g116809(.A (n_17520), .Y (n_17521));
NAND2X1 g116812(.A (n_32862), .B (n_16351), .Y (n_18050));
NAND2X2 g116815(.A (n_21068), .B (n_33982), .Y (n_18049));
NAND2X1 g116816(.A (n_16358), .B (n_35366), .Y (n_17518));
NAND2X1 g116817(.A (n_16987), .B (n_33982), .Y (n_17517));
INVX1 g116825(.A (n_17515), .Y (n_17516));
INVX1 g116831(.A (n_17512), .Y (n_17513));
OR2X1 g116833(.A (n_19206), .B (n_17510), .Y (n_17511));
NAND2X1 g116901(.A (n_16611), .B (n_17510), .Y (n_18045));
NAND2X1 g116902(.A (n_16610), .B (n_17510), .Y (n_17509));
INVX1 g116903(.A (n_17507), .Y (n_17508));
AND2X1 g116908(.A (n_16612), .B (n_33982), .Y (n_17506));
AND2X1 g116911(.A (n_17504), .B (n_17510), .Y (n_17505));
INVX1 g117032(.A (n_18198), .Y (n_17503));
INVX1 g117034(.A (n_17501), .Y (n_17502));
NOR2X1 g117100(.A (n_16658), .B (n_13723), .Y (n_18039));
INVX1 g117112(.A (n_17499), .Y (n_17500));
INVX1 g117116(.A (n_17497), .Y (n_17498));
NAND2X1 g117119(.A (n_16575), .B (n_15921), .Y (n_18035));
INVX1 g117125(.A (n_17495), .Y (n_19948));
AOI21X1 g117143(.A0 (n_16514), .A1 (n_32867), .B0 (n_16932), .Y(n_18033));
OAI21X1 g117145(.A0 (n_16051), .A1 (n_16517), .B0 (n_16261), .Y(n_18031));
INVX1 g117153(.A (n_17493), .Y (n_17494));
INVX1 g117158(.A (n_17491), .Y (n_17492));
NOR2X1 g117168(.A (n_16565), .B (n_13938), .Y (n_18028));
INVX1 g117193(.A (n_33767), .Y (n_18026));
AOI21X1 g117202(.A0 (n_16349), .A1 (n_19108), .B0 (n_9522), .Y(n_17489));
AOI22X1 g117223(.A0 (n_17474), .A1 (n_17472), .B0 (n_17471), .B1(n_17473), .Y (n_17488));
AOI21X1 g117224(.A0 (n_17468), .A1 (n_17467), .B0 (n_16606), .Y(n_17487));
AOI22X1 g117225(.A0 (n_17480), .A1 (n_9286), .B0 (n_17479), .B1(n_16202), .Y (n_17486));
OAI21X1 g117240(.A0 (n_35061), .A1 (n_34746), .B0 (n_17311), .Y(n_18859));
NAND2X1 g117251(.A (n_16614), .B (n_16041), .Y (n_18828));
INVX1 g117253(.A (n_17483), .Y (n_32577));
AOI21X1 g117257(.A0 (n_16504), .A1 (n_17482), .B0 (n_35063), .Y(n_18016));
AOI22X1 g117284(.A0 (n_17480), .A1 (n_17479), .B0 (n_9286), .B1(n_16202), .Y (n_17481));
AOI22X1 g117285(.A0 (n_17479), .A1 (n_7988), .B0 (n_11138), .B1(n_13735), .Y (n_17476));
AOI22X1 g117299(.A0 (n_17474), .A1 (n_17473), .B0 (n_17472), .B1(n_17471), .Y (n_17475));
AOI22X1 g117317(.A0 (n_10767), .A1 (n_16299), .B0 (n_9322), .B1(n_20235), .Y (n_17470));
AOI22X1 g117320(.A0 (n_17468), .A1 (n_16474), .B0 (n_17467), .B1(n_16026), .Y (n_17469));
NOR2X1 g117321(.A (n_16373), .B (n_16652), .Y (n_17466));
NAND2X1 g117335(.A (n_17968), .B (n_16643), .Y (n_17465));
NAND2X1 g117336(.A (n_17968), .B (n_17004), .Y (n_17464));
NAND2X1 g117340(.A (n_35816), .B (n_17004), .Y (n_17463));
NAND2X1 g117341(.A (n_35776), .B (n_16643), .Y (n_17461));
NAND2X1 g117350(.A (n_35736), .B (n_32496), .Y (n_17458));
INVX1 g117354(.A (n_18695), .Y (n_17984));
INVX1 g117360(.A (n_18062), .Y (n_17982));
NAND2X1 g117380(.A (n_14439), .B (n_32496), .Y (n_17455));
NOR2X1 g117385(.A (n_35206), .B (n_32984), .Y (n_17453));
INVX1 g117425(.A (n_16994), .Y (n_17978));
NAND2X2 g117432(.A (n_17916), .B (n_17732), .Y (n_17973));
INVX1 g117434(.A (n_16993), .Y (n_17972));
NAND2X1 g117450(.A (n_14439), .B (n_17451), .Y (n_17452));
NAND2X1 g117462(.A (n_35794), .B (n_17451), .Y (n_17450));
NAND2X2 g117478(.A (n_16904), .B (n_16475), .Y (n_19706));
INVX1 g117488(.A (n_17448), .Y (n_18639));
INVX1 g117494(.A (n_17446), .Y (n_17447));
INVX1 g117501(.A (n_17444), .Y (n_19709));
INVX1 g117506(.A (n_16985), .Y (n_17963));
INVX1 g117509(.A (n_17443), .Y (n_17961));
NAND2X1 g117511(.A (n_11089), .B (n_17398), .Y (n_19140));
INVX1 g117513(.A (n_17442), .Y (n_18645));
INVX1 g117520(.A (n_17441), .Y (n_18736));
INVX1 g117539(.A (n_17439), .Y (n_17958));
INVX1 g117570(.A (n_16972), .Y (n_17951));
INVX1 g117582(.A (n_16970), .Y (n_18778));
NAND2X1 g117586(.A (n_16903), .B (n_16028), .Y (n_18641));
NAND2X1 g117592(.A (n_17968), .B (n_16576), .Y (n_17433));
NAND2X1 g117603(.A (n_35540), .B (n_17451), .Y (n_17432));
NAND2X1 g117607(.A (n_35528), .B (n_32496), .Y (n_17431));
NAND2X1 g117608(.A (n_22021), .B (n_16643), .Y (n_17430));
NAND2X1 g117619(.A (n_13311), .B (n_32496), .Y (n_17429));
NAND2X1 g117622(.A (n_13311), .B (n_17451), .Y (n_17428));
NAND2X1 g117623(.A (n_18533), .B (n_17004), .Y (n_17427));
NOR2X1 g117627(.A (n_35529), .B (n_16804), .Y (n_17426));
NOR2X1 g117629(.A (n_35596), .B (n_16026), .Y (n_17425));
NAND2X1 g117642(.A (n_35776), .B (n_16576), .Y (n_17424));
INVX1 g117651(.A (n_16960), .Y (n_19306));
NAND2X1 g117660(.A (n_16958), .B (n_33032), .Y (n_17937));
NAND2X1 g117673(.A (n_17418), .B (n_18294), .Y (n_17419));
INVX1 g117676(.A (n_17416), .Y (n_32873));
INVX1 g117677(.A (n_17416), .Y (n_17415));
NAND2X1 g117681(.A (n_17413), .B (n_24101), .Y (n_17414));
NAND2X1 g117685(.A (n_17411), .B (n_18294), .Y (n_17412));
NAND2X1 g117702(.A (n_17409), .B (n_17713), .Y (n_17410));
NAND2X1 g117717(.A (n_16619), .B (n_32411), .Y (n_17932));
INVX1 g117726(.A (n_17406), .Y (n_17407));
NAND2X1 g117730(.A (n_10319), .B (n_33006), .Y (n_17931));
NOR2X1 g117744(.A (n_16537), .B (n_13738), .Y (n_17929));
NOR2X1 g117770(.A (n_17909), .B (n_17372), .Y (n_17927));
NAND2X1 g117771(.A (n_17418), .B (n_18498), .Y (n_17405));
INVX1 g117773(.A (n_16938), .Y (n_17926));
NAND2X1 g117777(.A (n_17413), .B (n_21919), .Y (n_17404));
NAND2X2 g117779(.A (n_16926), .B (n_17384), .Y (n_18765));
NAND2X1 g117780(.A (n_17411), .B (n_18498), .Y (n_17403));
INVX1 g117794(.A (n_18135), .Y (n_17402));
NAND2X1 g117797(.A (n_17409), .B (n_27770), .Y (n_17401));
NAND2X1 g117800(.A (n_17399), .B (n_27770), .Y (n_17400));
NAND2X1 g117804(.A (n_17398), .B (n_16031), .Y (n_19792));
NOR2X1 g117809(.A (n_35679), .B (n_15897), .Y (n_18782));
NAND2X1 g117815(.A (n_17409), .B (n_19595), .Y (n_17397));
NAND2X1 g117819(.A (n_16261), .B (n_17334), .Y (n_17920));
NOR2X1 g117825(.A (n_17413), .B (n_16798), .Y (n_18715));
INVX1 g117846(.A (n_17395), .Y (n_17396));
OR2X1 g117881(.A (n_17392), .B (n_16867), .Y (n_18597));
NAND2X1 g117884(.A (n_10334), .B (n_16541), .Y (n_17391));
INVX1 g117893(.A (n_17390), .Y (n_19167));
NAND2X1 g117895(.A (n_17418), .B (n_13268), .Y (n_17389));
NAND2X1 g117898(.A (n_17413), .B (n_13268), .Y (n_17388));
NAND2X1 g117904(.A (n_17411), .B (n_13268), .Y (n_17387));
NOR2X1 g117912(.A (n_17399), .B (n_19085), .Y (n_17386));
NAND2X2 g117918(.A (n_10320), .B (n_17372), .Y (n_17912));
INVX1 g117924(.A (n_18069), .Y (n_18704));
NAND2X2 g117929(.A (n_17384), .B (n_17906), .Y (n_19331));
NOR2X1 g117956(.A (n_17380), .B (n_33551), .Y (n_20763));
INVX1 g117965(.A (n_21501), .Y (n_17378));
INVX1 g117988(.A (n_18691), .Y (n_17374));
NAND2X1 g117991(.A (n_17909), .B (n_17372), .Y (n_19256));
NAND2X1 g117994(.A (n_10325), .B (n_16801), .Y (n_17371));
NAND2X1 g117999(.A (n_32602), .B (n_17000), .Y (n_18668));
INVX1 g118007(.A (n_17369), .Y (n_18690));
INVX1 g118036(.A (n_17363), .Y (n_18626));
NAND2X1 g118053(.A (n_16983), .B (n_33967), .Y (n_17903));
NAND2X1 g118056(.A (n_8830), .B (n_16218), .Y (n_18710));
INVX1 g118057(.A (n_18711), .Y (n_17359));
NAND2X1 g118059(.A (n_16984), .B (n_19626), .Y (n_19320));
INVX1 g118061(.A (n_17357), .Y (n_17358));
INVX1 g118068(.A (n_17356), .Y (n_17902));
NAND2X1 g118073(.A (n_10299), .B (n_33551), .Y (n_17901));
NAND2X1 g118074(.A (n_34383), .B (n_34387), .Y (n_18681));
OR2X1 g118076(.A (n_34383), .B (n_34387), .Y (n_18680));
INVX1 g118078(.A (n_18106), .Y (n_17898));
INVX1 g118081(.A (n_16905), .Y (n_17897));
NAND2X1 g118086(.A (n_16968), .B (n_16817), .Y (n_18677));
NAND2X1 g118090(.A (n_17351), .B (n_16810), .Y (n_17352));
NAND2X1 g118094(.A (n_10756), .B (n_16213), .Y (n_17895));
AND2X1 g118148(.A (n_18709), .B (n_16051), .Y (n_17349));
NAND2X1 g118153(.A (n_34617), .B (n_16853), .Y (n_18772));
NAND2X1 g118156(.A (n_34992), .B (n_34993), .Y (n_18771));
NAND2X1 g118161(.A (n_17348), .B (n_16851), .Y (n_20264));
NOR2X1 g118163(.A (n_16239), .B (n_17014), .Y (n_18601));
NAND2X1 g118172(.A (n_16533), .B (n_17343), .Y (n_18708));
INVX1 g118177(.A (n_17344), .Y (n_17345));
NAND2X1 g118195(.A (n_16521), .B (n_17343), .Y (n_17889));
NAND2X1 g118204(.A (n_17418), .B (n_17340), .Y (n_17342));
NAND2X1 g118205(.A (n_17413), .B (n_17340), .Y (n_17341));
NOR2X1 g118207(.A (n_16531), .B (n_16569), .Y (n_18615));
NAND2X1 g118208(.A (n_17411), .B (n_17340), .Y (n_17339));
NAND2X1 g118216(.A (n_17409), .B (n_23356), .Y (n_17338));
NAND2X1 g118228(.A (n_33007), .B (n_17337), .Y (n_17886));
AND2X1 g118259(.A (n_18057), .B (n_17335), .Y (n_17882));
NAND2X1 g118268(.A (n_17343), .B (n_17334), .Y (n_18721));
NAND2X1 g118279(.A (n_18533), .B (n_16576), .Y (n_17331));
NAND2X1 g118333(.A (n_16499), .B (n_17330), .Y (n_18637));
NAND2X1 g118336(.A (n_16499), .B (n_17878), .Y (n_17329));
NAND2X1 g118340(.A (n_16500), .B (n_34741), .Y (n_17328));
INVX1 g118341(.A (n_17326), .Y (n_18631));
NAND2X1 g118343(.A (n_17312), .B (n_16826), .Y (n_17325));
NAND2X1 g118347(.A (n_16864), .B (n_17320), .Y (n_17322));
NAND2X1 g118355(.A (n_17320), .B (n_16265), .Y (n_18633));
NAND2X1 g118356(.A (n_16824), .B (n_17317), .Y (n_17318));
INVX1 g118357(.A (n_34744), .Y (n_17316));
INVX1 g118360(.A (n_17315), .Y (n_17874));
INVX1 g118364(.A (n_17314), .Y (n_19198));
AND2X1 g118386(.A (n_16041), .B (n_16613), .Y (n_17872));
NAND2X1 g118395(.A (n_18018), .B (n_17312), .Y (n_20324));
NAND2X1 g118399(.A (n_18012), .B (n_17320), .Y (n_20323));
NAND2X1 g118407(.A (n_17311), .B (n_34740), .Y (n_20328));
OAI21X1 g118416(.A0 (n_16273), .A1 (n_17848), .B0 (n_23545), .Y(n_17309));
OAI21X1 g118442(.A0 (n_16275), .A1 (n_17848), .B0 (n_23045), .Y(n_17308));
OAI21X1 g118448(.A0 (n_16273), .A1 (n_14279), .B0 (n_23535), .Y(n_17307));
OAI21X1 g118452(.A0 (n_16273), .A1 (n_17304), .B0 (n_23534), .Y(n_17305));
AOI21X1 g118453(.A0 (n_16546), .A1 (n_32715), .B0 (n_14497), .Y(n_17303));
AOI21X1 g118454(.A0 (n_17273), .A1 (n_32786), .B0 (n_14094), .Y(n_17302));
AND2X1 g118456(.A (n_16532), .B (n_23533), .Y (n_17301));
OAI21X1 g118475(.A0 (n_17300), .A1 (n_16842), .B0 (n_16854), .Y(n_17844));
AND2X1 g118480(.A (n_16535), .B (n_17298), .Y (n_17299));
OAI21X1 g118496(.A0 (n_16327), .A1 (n_19024), .B0 (n_23042), .Y(n_17297));
OAI21X1 g118506(.A0 (n_16327), .A1 (n_17304), .B0 (n_23040), .Y(n_17296));
OAI21X1 g118518(.A0 (n_16275), .A1 (n_32677), .B0 (n_23038), .Y(n_17295));
OAI21X1 g118527(.A0 (n_17289), .A1 (n_17293), .B0 (n_19329), .Y(n_18768));
OAI21X1 g118528(.A0 (n_20572), .A1 (n_14042), .B0 (n_17292), .Y(n_18760));
OAI21X1 g118529(.A0 (n_20572), .A1 (n_32646), .B0 (n_18815), .Y(n_18754));
OAI21X1 g118530(.A0 (n_17289), .A1 (n_13183), .B0 (n_19327), .Y(n_18746));
OAI21X1 g118531(.A0 (n_17289), .A1 (n_13434), .B0 (n_19328), .Y(n_18743));
NAND2X1 g118532(.A (n_16529), .B (n_18814), .Y (n_18726));
OAI21X1 g118533(.A0 (n_20572), .A1 (n_17288), .B0 (n_18809), .Y(n_18655));
OAI21X1 g118534(.A0 (n_17289), .A1 (n_17287), .B0 (n_19325), .Y(n_18661));
OAI21X1 g118536(.A0 (n_17284), .A1 (n_17856), .B0 (n_20022), .Y(n_17286));
OAI21X1 g118545(.A0 (n_17284), .A1 (n_18429), .B0 (n_20021), .Y(n_17285));
OAI21X1 g118548(.A0 (n_17284), .A1 (n_32698), .B0 (n_20020), .Y(n_17283));
NAND2X1 g118552(.A (n_9530), .B (n_16528), .Y (n_17282));
OAI21X1 g118556(.A0 (n_12532), .A1 (n_15943), .B0 (n_16856), .Y(n_18748));
OAI21X1 g118557(.A0 (n_17284), .A1 (n_18441), .B0 (n_20019), .Y(n_17280));
OAI22X1 g118565(.A0 (n_16149), .A1 (n_15723), .B0 (n_6303), .B1(n_15722), .Y (n_17279));
AOI22X1 g118566(.A0 (n_16857), .A1 (n_19108), .B0 (n_11138), .B1(n_7755), .Y (n_17278));
AOI21X1 g118571(.A0 (n_10317), .A1 (n_9292), .B0 (n_16495), .Y(n_17277));
AOI22X1 g118572(.A0 (n_16546), .A1 (n_18909), .B0 (n_18289), .B1(n_9634), .Y (n_17276));
AOI22X1 g118574(.A0 (n_17273), .A1 (n_10848), .B0 (n_18289), .B1(n_1183), .Y (n_17274));
INVX1 g118577(.A (n_16874), .Y (n_17271));
AOI21X1 g118592(.A0 (n_18289), .A1 (n_10594), .B0 (n_16494), .Y(n_17270));
AOI21X1 g118593(.A0 (n_18289), .A1 (n_8193), .B0 (n_16496), .Y(n_17268));
AOI21X1 g118598(.A0 (n_9292), .A1 (n_17273), .B0 (n_16519), .Y(n_17267));
OAI22X1 g118602(.A0 (n_17262), .A1 (n_17259), .B0 (n_17261), .B1(n_17260), .Y (n_17264));
OAI22X1 g118603(.A0 (n_17262), .A1 (n_17261), .B0 (n_17260), .B1(n_17259), .Y (n_17263));
INVX1 g118721(.A (n_16869), .Y (n_17824));
INVX1 g118738(.A (n_19523), .Y (n_19000));
NAND2X1 g118748(.A (n_16180), .B (n_35398), .Y (n_17257));
INVX1 g118763(.A (n_17256), .Y (n_17810));
NAND2X1 g118798(.A (n_17831), .B (n_17830), .Y (n_18518));
NOR2X1 g118801(.A (n_18435), .B (n_17139), .Y (n_17255));
NAND2X1 g118824(.A (n_16445), .B (n_17253), .Y (n_19915));
NOR2X1 g118837(.A (n_17240), .B (n_16396), .Y (n_17252));
INVX2 g118842(.A (n_17908), .Y (n_20744));
AND2X1 g118864(.A (n_18969), .B (n_16425), .Y (n_17788));
INVX1 g118865(.A (n_17250), .Y (n_19073));
INVX1 g118877(.A (n_16855), .Y (n_17784));
OR2X1 g118884(.A (n_17249), .B (n_17248), .Y (n_17782));
NAND2X1 g118886(.A (n_17843), .B (n_16433), .Y (n_21390));
NAND2X1 g118888(.A (n_17300), .B (n_16170), .Y (n_19651));
INVX1 g118896(.A (n_19652), .Y (n_17247));
INVX2 g118903(.A (n_17246), .Y (n_17776));
INVX1 g118918(.A (n_17894), .Y (n_17775));
INVX1 g118923(.A (n_18580), .Y (n_17774));
INVX1 g118934(.A (n_17242), .Y (n_17772));
INVX1 g118947(.A (n_17892), .Y (n_17241));
NOR2X1 g118992(.A (n_17240), .B (n_17786), .Y (n_20361));
OR2X1 g118993(.A (n_35949), .B (n_17240), .Y (n_17239));
INVX1 g119003(.A (n_19724), .Y (n_17235));
OR2X1 g119005(.A (n_17233), .B (n_19790), .Y (n_17234));
INVX1 g119014(.A (n_17231), .Y (n_17232));
INVX1 g119043(.A (n_17230), .Y (n_17768));
INVX1 g119100(.A (n_17228), .Y (n_18466));
INVX1 g119108(.A (n_16825), .Y (n_19230));
INVX1 g119136(.A (n_34385), .Y (n_20175));
INVX1 g119140(.A (n_16823), .Y (n_19135));
NAND2X1 g119143(.A (n_18061), .B (n_17226), .Y (n_17760));
NOR2X1 g119145(.A (n_17794), .B (n_18379), .Y (n_18457));
NAND2X1 g119156(.A (n_35398), .B (n_17226), .Y (n_17759));
INVX1 g119171(.A (n_17224), .Y (n_17756));
NOR2X1 g119185(.A (n_17647), .B (n_18561), .Y (n_18456));
NAND2X1 g119216(.A (n_16436), .B (n_17221), .Y (n_20211));
NAND2X1 g119219(.A (n_16772), .B (n_17253), .Y (n_17747));
NAND2X1 g119230(.A (n_15797), .B (n_18909), .Y (n_17220));
INVX1 g119265(.A (n_17219), .Y (n_20188));
NAND2X1 g119276(.A (n_17743), .B (n_32362), .Y (n_17742));
NOR2X1 g119279(.A (n_17206), .B (n_32361), .Y (n_17218));
AND2X1 g119289(.A (n_16759), .B (n_19186), .Y (n_19046));
INVX1 g119306(.A (n_16486), .Y (n_19172));
INVX4 g119337(.A (n_33973), .Y (n_19626));
INVX1 g119346(.A (n_33968), .Y (n_19629));
NOR2X1 g119391(.A (n_17207), .B (n_17206), .Y (n_18412));
CLKBUFX1 g119396(.A (n_16477), .Y (n_19669));
NAND2X1 g119402(.A (n_17207), .B (n_32361), .Y (n_17204));
INVX2 g119407(.A (n_17203), .Y (n_23190));
INVX1 g119531(.A (n_17975), .Y (n_17731));
INVX1 g119607(.A (n_16465), .Y (n_19159));
AOI22X1 g119689(.A0 (n_16435), .A1 (n_16404), .B0 (n_16184), .B1(n_17186), .Y (n_17188));
AOI21X1 g119690(.A0 (n_35318), .A1 (n_16738), .B0 (n_16439), .Y(n_17185));
AOI22X1 g119691(.A0 (n_17182), .A1 (n_15952), .B0 (n_10717), .B1(n_16126), .Y (n_17183));
XOR2X1 g119705(.A (n_18159), .B (n_17172), .Y (n_17181));
NAND2X1 g119714(.A (n_16458), .B (n_16459), .Y (n_27451));
OAI21X1 g119715(.A0 (n_11333), .A1 (n_17178), .B0 (n_16456), .Y(n_17179));
NOR2X1 g119724(.A (n_8737), .B (n_17178), .Y (n_17177));
NAND2X1 g119744(.A (n_17674), .B (n_16777), .Y (n_17175));
NOR2X1 g119745(.A (n_17174), .B (n_16421), .Y (n_19052));
NAND2X1 g119754(.A (n_17172), .B (n_17150), .Y (n_17173));
NAND2X1 g119775(.A (n_35744), .B (n_16130), .Y (n_17168));
INVX1 g119780(.A (n_16785), .Y (n_17710));
INVX1 g119798(.A (n_34721), .Y (n_17166));
INVX1 g119805(.A (n_17820), .Y (n_18373));
INVX1 g119815(.A (n_17165), .Y (n_17701));
NAND2X1 g119820(.A (n_35816), .B (n_16137), .Y (n_17164));
NAND2X1 g119822(.A (n_17162), .B (n_16707), .Y (n_17163));
INVX1 g119828(.A (n_17161), .Y (n_17699));
INVX1 g119888(.A (n_17735), .Y (n_18321));
NOR2X1 g119918(.A (n_16754), .B (n_19474), .Y (n_17692));
NAND2X1 g119941(.A (n_11037), .B (n_19474), .Y (n_18355));
NAND2X1 g119946(.A (n_17150), .B (n_16420), .Y (n_17688));
NOR2X1 g119948(.A (n_11222), .B (n_18288), .Y (n_17149));
INVX1 g119954(.A (n_17822), .Y (n_17147));
NAND2X1 g119957(.A (n_12345), .B (n_23778), .Y (n_17146));
NAND2X1 g119965(.A (n_17968), .B (n_16457), .Y (n_17145));
NAND2X1 g119966(.A (n_22080), .B (n_16777), .Y (n_17143));
NAND2X1 g119977(.A (n_14439), .B (n_16137), .Y (n_17142));
NAND2X1 g119979(.A (n_35816), .B (n_17139), .Y (n_17140));
NAND2X1 g119981(.A (n_35736), .B (n_16457), .Y (n_17138));
INVX1 g119984(.A (n_17136), .Y (n_17137));
NAND2X1 g120002(.A (n_17131), .B (n_17130), .Y (n_17132));
NAND2X1 g120005(.A (n_18533), .B (n_16137), .Y (n_17129));
NAND2X1 g120006(.A (n_35473), .B (n_16130), .Y (n_17128));
INVX1 g120020(.A (n_17125), .Y (n_17657));
NOR2X1 g120025(.A (n_16171), .B (n_19471), .Y (n_17652));
NOR2X1 g120027(.A (n_17712), .B (n_16172), .Y (n_18324));
NAND2X1 g120028(.A (n_16734), .B (n_16454), .Y (n_17123));
CLKBUFX1 gbuf_d_383(.A(n_16556), .Y(d_out_383));
CLKBUFX1 gbuf_q_383(.A(q_in_383), .Y(P2_IR[27]));
CLKBUFX1 gbuf_d_384(.A(n_16553), .Y(d_out_384));
CLKBUFX1 gbuf_q_384(.A(q_in_384), .Y(P2_IR[25]));
CLKBUFX1 gbuf_d_385(.A(n_16550), .Y(d_out_385));
CLKBUFX1 gbuf_q_385(.A(q_in_385), .Y(P3_IR[26]));
CLKBUFX1 gbuf_d_386(.A(n_16551), .Y(d_out_386));
CLKBUFX1 gbuf_q_386(.A(q_in_386), .Y(P3_IR[25]));
CLKBUFX1 gbuf_d_387(.A(n_16416), .Y(d_out_387));
CLKBUFX1 gbuf_q_387(.A(q_in_387), .Y(P2_IR[29]));
CLKBUFX1 gbuf_d_388(.A(n_16414), .Y(d_out_388));
CLKBUFX1 gbuf_q_388(.A(q_in_388), .Y(P3_IR[31]));
INVX1 g120266(.A (n_17814), .Y (n_17112));
INVX1 g120142(.A (n_17831), .Y (n_18387));
XOR2X1 g115313(.A (n_17628), .B (n_17630), .Y (n_17635));
NOR2X1 g115622(.A (n_16683), .B (n_17552), .Y (n_17619));
NAND3X1 g115630(.A (n_17089), .B (n_17081), .C (n_16685), .Y(n_17090));
NOR2X1 g115634(.A (n_16671), .B (n_16672), .Y (n_17088));
NOR2X1 g115642(.A (n_17086), .B (n_17085), .Y (n_17087));
OAI21X1 g116070(.A0 (n_17055), .A1 (n_17084), .B0 (n_16305), .Y(n_17598));
INVX1 g116098(.A (n_17082), .Y (n_17083));
AOI21X1 g116102(.A0 (n_16370), .A1 (n_17081), .B0 (n_17080), .Y(n_17596));
OAI21X1 g116122(.A0 (n_16371), .A1 (n_17025), .B0 (n_17036), .Y(n_17079));
INVX1 g116196(.A (n_16630), .Y (n_18894));
NOR2X1 g116299(.A (n_16641), .B (n_17058), .Y (n_17587));
NAND2X1 g116321(.A (n_15926), .B (n_17033), .Y (n_22947));
NAND2X2 g116335(.A (n_17076), .B (n_17075), .Y (n_17077));
NAND2X1 g116359(.A (n_16364), .B (n_17089), .Y (n_18189));
NAND2X1 g116363(.A (n_35951), .B (n_17073), .Y (n_17074));
NAND2X1 g116390(.A (n_17022), .B (n_17024), .Y (n_17072));
NAND2X1 g116395(.A (n_17023), .B (n_16628), .Y (n_17071));
NAND2X1 g116397(.A (n_16629), .B (n_17603), .Y (n_17070));
NAND2X1 g116401(.A (n_17063), .B (n_17073), .Y (n_19375));
NAND2X1 g116404(.A (n_18093), .B (n_35951), .Y (n_17069));
NAND2X1 g116409(.A (n_18682), .B (n_17067), .Y (n_17068));
NAND2X1 g116412(.A (n_16298), .B (n_16587), .Y (n_17066));
NOR2X1 g116413(.A (n_17595), .B (n_16326), .Y (n_18180));
INVX1 g116417(.A (n_16692), .Y (n_17574));
CLKBUFX1 gbuf_d_389(.A(n_16277), .Y(d_out_389));
CLKBUFX1 gbuf_q_389(.A(q_in_389), .Y(P1_IR[27]));
INVX1 g116425(.A (n_16689), .Y (n_18853));
NAND2X2 g116438(.A (n_17064), .B (n_17063), .Y (n_17065));
NAND2X1 g116439(.A (n_16306), .B (n_17064), .Y (n_17062));
NAND2X1 g116456(.A (n_17064), .B (n_18685), .Y (n_17564));
NAND2X1 g116468(.A (n_16626), .B (n_16355), .Y (n_17061));
NAND2X1 g116498(.A (n_16268), .B (n_15953), .Y (n_18184));
INVX1 g116516(.A (n_17059), .Y (n_17060));
NAND2X1 g116551(.A (n_17057), .B (n_18170), .Y (n_21502));
NOR2X1 g116557(.A (n_17056), .B (n_16097), .Y (n_17555));
NOR2X1 g116585(.A (n_16306), .B (n_17055), .Y (n_22197));
NAND2X1 g116593(.A (n_35218), .B (n_32503), .Y (n_17054));
NAND2X1 g116627(.A (n_17073), .B (n_17084), .Y (n_23625));
NOR2X1 g116631(.A (n_16274), .B (n_16272), .Y (n_18231));
INVX1 g116645(.A (n_17053), .Y (n_17546));
NAND2X1 g116653(.A (n_16267), .B (n_17051), .Y (n_17052));
INVX1 g116662(.A (n_17617), .Y (n_17048));
NAND2X1 g116670(.A (n_17056), .B (n_16390), .Y (n_17047));
NAND2X1 g116673(.A (n_34064), .B (n_17051), .Y (n_17539));
NAND2X1 g116674(.A (n_17045), .B (n_16609), .Y (n_17046));
NAND2X1 g116677(.A (n_35350), .B (n_17606), .Y (n_17536));
NAND2X1 g116684(.A (n_16602), .B (n_34065), .Y (n_17040));
NAND3X1 g116687(.A (n_16276), .B (n_11785), .C (n_16560), .Y(n_19397));
NAND2X1 g116693(.A (n_17057), .B (n_16591), .Y (n_17039));
NAND2X1 g116700(.A (n_34107), .B (n_35913), .Y (n_17532));
OR2X1 g116732(.A (n_17552), .B (n_16368), .Y (n_17038));
AND2X1 g116733(.A (n_34171), .B (n_17036), .Y (n_17037));
INVX1 g116754(.A (n_17035), .Y (n_17524));
NAND2X1 g116758(.A (n_35914), .B (n_17033), .Y (n_17034));
NAND2X1 g116760(.A (n_34065), .B (n_17057), .Y (n_17032));
NOR2X1 g116789(.A (n_17028), .B (n_16570), .Y (n_17029));
AND2X1 g116790(.A (n_17026), .B (n_17025), .Y (n_17027));
NOR2X1 g116810(.A (n_17024), .B (n_35882), .Y (n_17520));
NAND2X1 g116827(.A (n_17023), .B (n_17504), .Y (n_17515));
NAND2X1 g116832(.A (n_17022), .B (n_17021), .Y (n_17512));
NAND2X1 g116896(.A (n_18157), .B (n_19974), .Y (n_17020));
NAND3X1 g116897(.A (n_16073), .B (n_17018), .C (n_17017), .Y(n_32578));
NAND2X1 g116904(.A (n_16666), .B (n_16612), .Y (n_17507));
NAND2X1 g116907(.A (n_17015), .B (n_16690), .Y (n_17016));
NAND2X1 g116937(.A (n_16350), .B (n_22758), .Y (n_18190));
NAND2X1 g117033(.A (n_16344), .B (n_19410), .Y (n_18198));
NAND2X1 g117035(.A (n_16348), .B (n_19389), .Y (n_17501));
NAND2X1 g117036(.A (n_16342), .B (n_21874), .Y (n_18208));
NAND2X1 g117038(.A (n_16347), .B (n_22779), .Y (n_18205));
NAND2X1 g117040(.A (n_16346), .B (n_21545), .Y (n_18196));
CLKBUFX1 g117087(.A (n_17625), .Y (n_20012));
NAND2X1 g117097(.A (n_16377), .B (n_21875), .Y (n_18201));
NAND2X1 g117098(.A (n_16378), .B (n_13510), .Y (n_18203));
AOI21X1 g117113(.A0 (n_33769), .A1 (n_34581), .B0 (n_16946), .Y(n_17499));
OAI21X1 g117117(.A0 (n_17014), .A1 (n_17013), .B0 (n_15907), .Y(n_17497));
INVX1 g117127(.A (n_17610), .Y (n_17495));
OAI21X1 g117141(.A0 (n_16241), .A1 (n_32412), .B0 (n_16934), .Y(n_18194));
AOI21X1 g117154(.A0 (n_16337), .A1 (n_16260), .B0 (n_16944), .Y(n_17493));
NAND2X1 g117159(.A (n_16380), .B (n_21900), .Y (n_17491));
NOR2X1 g117162(.A (n_16383), .B (n_17012), .Y (n_18213));
NAND2X1 g117164(.A (n_16382), .B (n_19422), .Y (n_18219));
AOI22X1 g117226(.A0 (n_17007), .A1 (n_9624), .B0 (n_16349), .B1(n_17004), .Y (n_17010));
AOI22X1 g117227(.A0 (n_16577), .A1 (n_16644), .B0 (n_16643), .B1(n_16576), .Y (n_17009));
OAI21X1 g117254(.A0 (n_16569), .A1 (n_16664), .B0 (n_16530), .Y(n_17483));
AOI22X1 g117303(.A0 (n_17007), .A1 (n_16349), .B0 (n_9624), .B1(n_17004), .Y (n_17008));
INVX1 g117310(.A (n_16660), .Y (n_17003));
INVX1 g117314(.A (n_16659), .Y (n_17002));
AND2X1 g117323(.A (n_16360), .B (n_15938), .Y (n_17001));
NAND2X1 g117355(.A (n_10752), .B (n_16469), .Y (n_18695));
NAND2X1 g117361(.A (n_17000), .B (n_16468), .Y (n_18062));
INVX1 g117364(.A (n_34112), .Y (n_18097));
INVX1 g117374(.A (n_16999), .Y (n_18099));
NOR2X1 g117384(.A (n_18001), .B (n_18000), .Y (n_16998));
NAND2X1 g117391(.A (n_9761), .B (n_15798), .Y (n_16997));
INVX1 g117419(.A (n_17534), .Y (n_21047));
NAND2X1 g117426(.A (n_16593), .B (n_32982), .Y (n_16994));
NAND2X1 g117435(.A (n_9775), .B (n_16929), .Y (n_16993));
INVX1 g117464(.A (n_18096), .Y (n_16991));
INVX1 g117480(.A (n_16988), .Y (n_16989));
INVX1 g117489(.A (n_16987), .Y (n_17448));
NAND2X2 g117498(.A (n_8830), .B (n_16219), .Y (n_17446));
INVX1 g117502(.A (n_16986), .Y (n_17444));
NAND2X1 g117507(.A (n_16984), .B (n_33973), .Y (n_16985));
NAND2X1 g117510(.A (n_16983), .B (n_33968), .Y (n_17443));
INVX1 g117514(.A (n_16982), .Y (n_17442));
NAND2X1 g117521(.A (n_16585), .B (n_35686), .Y (n_17441));
NOR2X1 g117529(.A (n_10482), .B (n_17399), .Y (n_16980));
INVX1 g117540(.A (n_16099), .Y (n_17439));
NOR2X1 g117553(.A (n_9264), .B (n_16481), .Y (n_18583));
INVX1 g117560(.A (n_16973), .Y (n_16974));
NAND2X1 g117583(.A (n_10756), .B (n_17203), .Y (n_16970));
NAND2X1 g117591(.A (n_16968), .B (n_16488), .Y (n_19229));
NAND2X1 g117596(.A (n_17968), .B (n_17479), .Y (n_16967));
NOR2X1 g117613(.A (n_35600), .B (n_16320), .Y (n_16966));
NOR2X1 g117637(.A (n_35529), .B (n_16322), .Y (n_16965));
NAND2X1 g117638(.A (n_35736), .B (n_17479), .Y (n_16963));
NAND2X1 g117652(.A (n_16249), .B (n_16958), .Y (n_16960));
NAND2X1 g117653(.A (n_16250), .B (n_16958), .Y (n_16959));
AND2X1 g117678(.A (n_16242), .B (n_16955), .Y (n_17416));
NAND2X2 g117687(.A (n_32867), .B (n_35174), .Y (n_18774));
NOR2X1 g117701(.A (n_16197), .B (n_16294), .Y (n_18897));
NAND2X1 g117709(.A (n_17075), .B (n_16950), .Y (n_16951));
AND2X1 g117712(.A (n_33770), .B (n_35850), .Y (n_16949));
NOR2X1 g117714(.A (n_16946), .B (n_16046), .Y (n_16947));
NAND2X1 g117715(.A (n_16944), .B (n_16336), .Y (n_16945));
INVX1 g117723(.A (n_34843), .Y (n_16943));
NAND2X1 g117727(.A (n_20235), .B (n_16299), .Y (n_17406));
AND2X1 g117733(.A (n_15921), .B (n_16574), .Y (n_18599));
INVX1 g117750(.A (n_16618), .Y (n_19213));
NOR2X1 g117754(.A (n_16936), .B (n_16465), .Y (n_18146));
INVX1 g117755(.A (n_17578), .Y (n_16939));
NAND2X1 g117774(.A (n_35863), .B (n_18532), .Y (n_16938));
NAND2X1 g117795(.A (n_16229), .B (n_19957), .Y (n_18135));
NAND2X1 g117811(.A (n_32490), .B (n_16473), .Y (n_16937));
NOR2X1 g117822(.A (n_16936), .B (n_16197), .Y (n_18832));
NAND2X1 g117824(.A (n_16934), .B (n_16955), .Y (n_22978));
OR2X1 g117847(.A (n_32864), .B (n_16932), .Y (n_17395));
NAND2X1 g117868(.A (n_16929), .B (n_16646), .Y (n_18652));
OR2X1 g117894(.A (n_34383), .B (n_34385), .Y (n_17390));
AND2X1 g117899(.A (n_11787), .B (n_17922), .Y (n_16927));
NAND2X1 g117925(.A (n_16926), .B (n_16524), .Y (n_18069));
NAND2X1 g117966(.A (n_16922), .B (n_17045), .Y (n_21501));
NAND2X2 g117990(.A (n_10318), .B (n_33007), .Y (n_18691));
INVX1 g117996(.A (n_16598), .Y (n_17370));
NAND2X2 g117998(.A (n_16656), .B (n_16469), .Y (n_18717));
INVX1 g118008(.A (n_16594), .Y (n_17369));
INVX1 g118010(.A (n_16921), .Y (n_18151));
INVX1 g118012(.A (n_16920), .Y (n_18102));
INVX1 g118016(.A (n_16918), .Y (n_16917));
INVX1 g118026(.A (n_16915), .Y (n_17366));
INVX1 g118030(.A (n_16914), .Y (n_17365));
INVX1 g118033(.A (n_16589), .Y (n_17364));
NOR2X1 g118037(.A (n_10319), .B (n_33007), .Y (n_17363));
INVX1 g118039(.A (n_16912), .Y (n_17361));
INVX1 g118048(.A (n_18684), .Y (n_17360));
NAND2X1 g118050(.A (n_8384), .B (n_16219), .Y (n_19733));
NAND2X1 g118058(.A (n_16624), .B (n_33968), .Y (n_18711));
NAND2X2 g118060(.A (n_9623), .B (n_33973), .Y (n_18683));
INVX1 g118062(.A (n_16907), .Y (n_17357));
NAND2X1 g118069(.A (n_10271), .B (n_16542), .Y (n_17356));
NAND2X1 g118079(.A (n_9701), .B (n_17203), .Y (n_18106));
NAND2X1 g118082(.A (n_16904), .B (n_34357), .Y (n_16905));
NAND2X1 g118083(.A (n_9331), .B (n_16212), .Y (n_19242));
NAND2X1 g118087(.A (n_9627), .B (n_16488), .Y (n_18676));
NAND2X1 g118091(.A (n_16903), .B (n_16477), .Y (n_19245));
INVX1 g118095(.A (n_17549), .Y (n_16902));
INVX1 g118113(.A (n_16586), .Y (n_18127));
NAND2X1 g118137(.A (n_33770), .B (n_16060), .Y (n_16899));
NAND2X1 g118139(.A (n_17075), .B (n_16054), .Y (n_16898));
NAND2X1 g118167(.A (n_16506), .B (n_16249), .Y (n_16897));
NAND2X1 g118170(.A (n_16895), .B (n_35173), .Y (n_18855));
NAND2X1 g118171(.A (n_35175), .B (n_16932), .Y (n_16894));
NAND2X1 g118173(.A (n_16946), .B (n_16619), .Y (n_16893));
INVX1 g118175(.A (n_16892), .Y (n_17346));
INVX1 g118178(.A (n_33768), .Y (n_17344));
NOR2X1 g118199(.A (n_16256), .B (n_35218), .Y (n_16891));
NAND2X1 g118223(.A (n_10322), .B (n_17928), .Y (n_16890));
INVX1 g118232(.A (n_16886), .Y (n_16887));
INVX1 g118235(.A (n_35942), .Y (n_16885));
NOR2X1 g118281(.A (n_35555), .B (n_16318), .Y (n_16881));
NAND2X1 g118282(.A (n_18533), .B (n_17479), .Y (n_16880));
AND2X1 g118285(.A (n_16878), .B (n_32533), .Y (n_16879));
NOR2X1 g118288(.A (n_16944), .B (n_16071), .Y (n_18614));
NAND2X1 g118342(.A (n_16265), .B (n_17312), .Y (n_17326));
INVX2 g118344(.A (n_16559), .Y (n_18632));
INVX1 g118348(.A (n_16558), .Y (n_18046));
NAND2X1 g118361(.A (n_17317), .B (n_17312), .Y (n_17315));
INVX2 g118362(.A (n_16557), .Y (n_18060));
NAND2X1 g118365(.A (n_17330), .B (n_16540), .Y (n_17314));
NAND2X1 g118387(.A (n_35059), .B (n_35061), .Y (n_22706));
INVX1 g118562(.A (n_16876), .Y (n_18142));
OAI22X1 g118569(.A0 (n_34913), .A1 (n_349), .B0 (n_15985), .B1(n_7243), .Y (n_16875));
NAND2X1 g118578(.A (n_16258), .B (n_16065), .Y (n_16874));
AOI22X1 g118599(.A0 (n_8829), .A1 (n_32428), .B0 (n_10451), .B1(n_16546), .Y (n_16873));
INVX1 g118607(.A (n_16872), .Y (n_18149));
INVX1 g118608(.A (n_16871), .Y (n_18108));
INVX1 g118611(.A (n_18163), .Y (n_16870));
NAND2X1 g118722(.A (n_17767), .B (n_34720), .Y (n_16869));
INVX2 g118739(.A (n_16867), .Y (n_19523));
NAND2X1 g118749(.A (n_17273), .B (n_18399), .Y (n_16866));
NAND2X1 g118764(.A (n_11278), .B (n_35622), .Y (n_17256));
OR2X1 g118778(.A (n_18561), .B (n_19766), .Y (n_18517));
NAND2X1 g118779(.A (n_17273), .B (n_15089), .Y (n_16862));
OR2X1 g118799(.A (n_16518), .B (n_32745), .Y (n_16861));
NAND2X1 g118820(.A (n_18145), .B (n_16181), .Y (n_17884));
INVX2 g118843(.A (n_17372), .Y (n_17908));
INVX1 g118859(.A (n_17384), .Y (n_17251));
AND2X1 g118866(.A (n_35949), .B (n_17233), .Y (n_17250));
NAND2X1 g118867(.A (n_16857), .B (n_18262), .Y (n_16858));
NAND2X1 g118878(.A (n_16444), .B (n_33051), .Y (n_16855));
NAND2X1 g118897(.A (n_16854), .B (n_16169), .Y (n_19652));
INVX1 g118904(.A (n_16853), .Y (n_17246));
INVX1 g118919(.A (n_16851), .Y (n_17894));
INVX2 g118924(.A (n_16522), .Y (n_18580));
INVX1 g118927(.A (n_16958), .Y (n_17243));
AND2X1 g118930(.A (n_18091), .B (n_16845), .Y (n_19891));
INVX1 g118935(.A (n_16849), .Y (n_17242));
INVX1 g118938(.A (n_16847), .Y (n_16848));
AND2X1 g118948(.A (n_16845), .B (n_16170), .Y (n_17892));
INVX1 g118952(.A (n_35063), .Y (n_16844));
NAND2X1 g118962(.A (n_16450), .B (n_16843), .Y (n_20916));
NOR2X1 g118981(.A (n_16842), .B (n_16841), .Y (n_19238));
NOR2X1 g118991(.A (n_10309), .B (n_16181), .Y (n_16840));
NOR2X1 g118994(.A (n_16837), .B (n_16836), .Y (n_16838));
NOR2X1 g118995(.A (n_16842), .B (n_16835), .Y (n_19236));
NOR2X1 g118996(.A (n_11790), .B (n_16837), .Y (n_16834));
NOR2X1 g118997(.A (n_11483), .B (n_16836), .Y (n_16833));
OR2X1 g118998(.A (n_16854), .B (n_16835), .Y (n_16832));
INVX1 g119000(.A (n_16517), .Y (n_17236));
AND2X1 g119004(.A (n_16164), .B (n_16448), .Y (n_19724));
INVX1 g119015(.A (n_17343), .Y (n_17231));
NAND2X1 g119020(.A (n_17273), .B (n_20154), .Y (n_16831));
INVX1 g119025(.A (n_21395), .Y (n_16830));
NAND2X1 g119044(.A (n_16829), .B (n_16117), .Y (n_17230));
NAND2X1 g119085(.A (n_16417), .B (n_16505), .Y (n_17923));
NAND2X1 g119101(.A (n_18667), .B (n_16820), .Y (n_17228));
NAND2X1 g119109(.A (n_17253), .B (n_17221), .Y (n_16825));
NAND2X1 g119141(.A (n_35244), .B (n_16392), .Y (n_16823));
INVX1 g119153(.A (n_17885), .Y (n_16821));
NAND2X1 g119172(.A (n_17221), .B (n_16820), .Y (n_17224));
INVX1 g119179(.A (n_16497), .Y (n_17223));
NAND2X1 g119182(.A (n_16857), .B (n_25596), .Y (n_16819));
NAND2X1 g119184(.A (n_16857), .B (n_35528), .Y (n_16818));
INVX1 g119266(.A (n_16817), .Y (n_17219));
INVX1 g119329(.A (n_17398), .Y (n_19631));
INVX2 g119408(.A (n_16213), .Y (n_17203));
INVX1 g119418(.A (n_16808), .Y (n_20830));
INVX1 g119517(.A (n_19071), .Y (n_17970));
CLKBUFX1 g119532(.A (n_16801), .Y (n_17975));
INVX1 g119578(.A (n_16799), .Y (n_18511));
AOI22X1 g119688(.A0 (n_16796), .A1 (n_17150), .B0 (n_16460), .B1(n_16420), .Y (n_16797));
XOR2X1 g119711(.A (n_16734), .B (n_18164), .Y (n_16795));
OAI21X1 g119712(.A0 (n_16176), .A1 (n_16777), .B0 (n_16177), .Y(n_16794));
NAND2X1 g119719(.A (n_12349), .B (n_17172), .Y (n_16793));
INVX1 g119720(.A (n_18437), .Y (n_16792));
INVX1 g119728(.A (n_17860), .Y (n_16791));
INVX1 g119788(.A (n_35399), .Y (n_17763));
NAND2X1 g119801(.A (n_16419), .B (n_16403), .Y (n_18705));
NAND2X1 g119806(.A (n_15966), .B (n_10666), .Y (n_17820));
NAND2X1 g119813(.A (n_16778), .B (n_16777), .Y (n_16782));
NAND2X1 g119816(.A (n_16182), .B (n_16173), .Y (n_17165));
OR2X1 g119817(.A (n_16778), .B (n_16777), .Y (n_16779));
NOR2X1 g119821(.A (n_16176), .B (n_16400), .Y (n_16776));
NAND2X1 g119829(.A (n_16435), .B (n_17186), .Y (n_17161));
NAND2X1 g119838(.A (n_16446), .B (n_15955), .Y (n_18426));
INVX1 g119840(.A (n_17226), .Y (n_17866));
INVX1 g119846(.A (n_16773), .Y (n_17158));
NOR2X1 g119853(.A (n_16435), .B (n_16135), .Y (n_32382));
INVX1 g119858(.A (n_16771), .Y (n_17803));
NAND2X1 g119861(.A (n_16768), .B (n_16740), .Y (n_16770));
OR2X1 g119862(.A (n_16768), .B (n_16740), .Y (n_16769));
INVX1 g119865(.A (n_17249), .Y (n_16767));
NOR2X1 g119881(.A (n_16750), .B (n_15854), .Y (n_17777));
INVX1 g119884(.A (n_19186), .Y (n_19505));
NAND2X2 g119889(.A (n_16748), .B (n_16140), .Y (n_17735));
INVX1 g119893(.A (n_16764), .Y (n_17155));
INVX1 g119905(.A (n_16761), .Y (n_18320));
INVX1 g119906(.A (n_16761), .Y (n_16760));
INVX2 g119914(.A (n_16759), .Y (n_17740));
INVX1 g119931(.A (n_16757), .Y (n_18434));
INVX1 g119935(.A (n_16755), .Y (n_21748));
NAND2X1 g119939(.A (n_16754), .B (n_15852), .Y (n_18773));
NAND2X1 g119944(.A (n_17172), .B (n_16731), .Y (n_19187));
NAND2X1 g119947(.A (n_16747), .B (n_16745), .Y (n_20301));
NAND2X1 g119955(.A (n_16407), .B (n_16406), .Y (n_17822));
NAND2X1 g119961(.A (n_16750), .B (n_15854), .Y (n_19183));
NAND2X1 g119968(.A (n_16748), .B (n_16747), .Y (n_16749));
INVX1 g119969(.A (n_16746), .Y (n_17766));
NAND2X1 g119985(.A (n_11503), .B (n_16745), .Y (n_17136));
INVX1 g119993(.A (n_17222), .Y (n_16742));
NOR2X1 g119996(.A (n_16174), .B (n_16740), .Y (n_16741));
NAND2X1 g120001(.A (n_16738), .B (n_16402), .Y (n_16739));
NOR2X1 g120021(.A (n_17712), .B (n_16171), .Y (n_17125));
NOR2X1 g120022(.A (n_16740), .B (n_17639), .Y (n_16737));
NAND2X1 g120026(.A (n_15950), .B (n_16162), .Y (n_20102));
NAND2X1 g120031(.A (n_16735), .B (n_16777), .Y (n_32888));
NAND2X1 g120032(.A (n_16734), .B (n_16777), .Y (n_19162));
NAND2X1 g120035(.A (n_16732), .B (n_16731), .Y (n_16733));
CLKBUFX1 gbuf_d_390(.A(n_16152), .Y(d_out_390));
CLKBUFX1 gbuf_q_390(.A(q_in_390), .Y(P2_IR[22]));
CLKBUFX1 gbuf_d_391(.A(n_16151), .Y(d_out_391));
CLKBUFX1 gbuf_q_391(.A(q_in_391), .Y(P2_IR[30]));
CLKBUFX1 gbuf_d_392(.A(n_16145), .Y(d_out_392));
CLKBUFX1 gbuf_q_392(.A(q_in_392), .Y(P2_IR[31]));
INVX1 g120211(.A (n_18997), .Y (n_17117));
CLKBUFX1 gbuf_d_393(.A(n_16147), .Y(d_out_393));
CLKBUFX1 gbuf_q_393(.A(q_in_393), .Y(P3_IR[28]));
INVX1 g120221(.A (n_17647), .Y (n_17116));
CLKBUFX1 gbuf_d_394(.A(n_16146), .Y(d_out_394));
CLKBUFX1 gbuf_q_394(.A(q_in_394), .Y(P1_IR[29]));
INVX1 g120241(.A (n_16837), .Y (n_17800));
INVX1 g120250(.A (n_16836), .Y (n_17798));
INVX1 g120409(.A (n_16420), .Y (n_20741));
CLKBUFX1 g120430(.A (n_17174), .Y (n_18948));
CLKBUFX1 g120512(.A (n_16134), .Y (n_17680));
INVX1 g120528(.A (n_17130), .Y (n_17682));
INVX1 g120154(.A (n_17830), .Y (n_17092));
INVX1 g114913(.A (n_16701), .Y (n_16702));
OAI21X1 g116099(.A0 (n_34362), .A1 (n_16699), .B0 (n_35915), .Y(n_17082));
NAND2X1 g116316(.A (n_18824), .B (n_16359), .Y (n_32915));
INVX1 g116346(.A (n_16696), .Y (n_16697));
NAND3X1 g116394(.A (n_16694), .B (n_15804), .C (n_16693), .Y(n_16695));
NAND2X1 g116418(.A (n_35221), .B (n_18088), .Y (n_16692));
NAND2X1 g116420(.A (n_16371), .B (n_16690), .Y (n_16691));
NAND2X1 g116426(.A (n_16351), .B (n_16354), .Y (n_16689));
OR2X1 g116500(.A (n_11079), .B (n_16269), .Y (n_16688));
NAND2X1 g116512(.A (n_16374), .B (n_17036), .Y (n_16687));
NAND2X1 g116517(.A (n_16324), .B (n_16109), .Y (n_17059));
NAND2X1 g116519(.A (n_16107), .B (n_16685), .Y (n_16686));
INVX1 g116523(.A (n_16683), .Y (n_16684));
NAND2X1 g116527(.A (n_16066), .B (n_16367), .Y (n_16682));
NAND2X2 g116646(.A (n_16690), .B (n_18088), .Y (n_17053));
INVX1 g116657(.A (n_16388), .Y (n_17049));
NAND2X1 g116659(.A (n_16312), .B (n_17615), .Y (n_16680));
NAND2X1 g116660(.A (n_16311), .B (n_16678), .Y (n_16679));
NAND2X1 g116663(.A (n_17025), .B (n_16677), .Y (n_17617));
NAND2X1 g116664(.A (n_17552), .B (n_17025), .Y (n_16676));
INVX1 g116735(.A (n_17086), .Y (n_16675));
INVX1 g116750(.A (n_16673), .Y (n_16674));
NAND2X1 g116755(.A (n_17045), .B (n_16678), .Y (n_17035));
INVX1 g116772(.A (n_16672), .Y (n_18235));
INVX1 g116777(.A (n_16671), .Y (n_17030));
INVX1 g116782(.A (n_17085), .Y (n_16670));
NAND2X1 g116799(.A (n_35352), .B (n_16376), .Y (n_16669));
NAND2X1 g116899(.A (n_16666), .B (n_33977), .Y (n_16667));
AOI21X1 g116981(.A0 (n_16878), .A1 (n_15813), .B0 (n_32535), .Y(n_16665));
NAND2X2 g117088(.A (n_16074), .B (n_16664), .Y (n_17625));
NAND2X2 g117128(.A (n_16080), .B (n_16663), .Y (n_17610));
CLKBUFX1 gbuf_d_395(.A(n_15971), .Y(d_out_395));
CLKBUFX1 gbuf_q_395(.A(q_in_395), .Y(P1_IR[28]));
INVX1 g117184(.A (n_34545), .Y (n_16662));
AOI22X1 g117311(.A0 (n_16381), .A1 (n_7988), .B0 (n_11138), .B1(P3_reg3[0] ), .Y (n_16660));
AOI22X1 g117315(.A0 (n_16379), .A1 (n_7988), .B0 (n_11138), .B1(n_13675), .Y (n_16659));
NOR2X1 g117342(.A (n_35840), .B (n_15937), .Y (n_16658));
NAND2X2 g117347(.A (n_16656), .B (n_33905), .Y (n_19235));
INVX1 g117366(.A (n_17058), .Y (n_16655));
NAND2X2 g117370(.A (n_9274), .B (n_17997), .Y (n_17533));
INVX1 g117375(.A (n_16653), .Y (n_16999));
NOR2X1 g117383(.A (n_10699), .B (n_17997), .Y (n_16652));
INVX1 g117399(.A (n_16650), .Y (n_18071));
INVX2 g117415(.A (n_16647), .Y (n_17569));
INVX1 g117416(.A (n_16647), .Y (n_35632));
INVX1 g117420(.A (n_16366), .Y (n_17534));
NAND2X2 g117428(.A (n_16646), .B (n_16199), .Y (n_19304));
NAND2X1 g117437(.A (n_16644), .B (n_16643), .Y (n_16645));
INVX1 g117445(.A (n_16641), .Y (n_17543));
INVX1 g117455(.A (n_34107), .Y (n_16640));
NAND2X1 g117465(.A (n_9223), .B (n_32995), .Y (n_18096));
INVX2 g117470(.A (n_17024), .Y (n_21068));
NOR2X1 g117474(.A (n_9780), .B (n_16936), .Y (n_16637));
INVX1 g117479(.A (n_16635), .Y (n_16636));
INVX1 g117481(.A (n_16635), .Y (n_16988));
INVX1 g117490(.A (n_17022), .Y (n_16987));
INVX1 g117492(.A (n_18644), .Y (n_16633));
NAND2X1 g117499(.A (n_8384), .B (n_16218), .Y (n_19210));
NAND2X1 g117503(.A (n_9181), .B (n_33972), .Y (n_16986));
INVX1 g117515(.A (n_16631), .Y (n_16982));
INVX1 g117516(.A (n_16631), .Y (n_16632));
NAND2X1 g117522(.A (n_15824), .B (n_16590), .Y (n_16630));
INVX1 g117524(.A (n_16629), .Y (n_18735));
INVX1 g117527(.A (n_17603), .Y (n_18792));
INVX1 g117534(.A (n_21528), .Y (n_16978));
INVX1 g117549(.A (n_16626), .Y (n_16975));
NAND2X2 g117552(.A (n_16293), .B (n_35674), .Y (n_17570));
INVX2 g117557(.A (n_17023), .Y (n_19206));
NAND2X2 g117564(.A (n_16624), .B (n_33967), .Y (n_16973));
NAND2X2 g117572(.A (n_9627), .B (n_16222), .Y (n_16972));
NAND2X2 g117576(.A (n_9227), .B (n_16213), .Y (n_19208));
NAND2X2 g117590(.A (n_9331), .B (n_34357), .Y (n_19827));
INVX1 g117741(.A (n_16338), .Y (n_18192));
NAND2X1 g117751(.A (n_17334), .B (n_35175), .Y (n_16618));
INVX1 g117752(.A (n_17021), .Y (n_18620));
NAND2X1 g117756(.A (n_15912), .B (n_16042), .Y (n_17578));
INVX1 g117791(.A (n_16334), .Y (n_18144));
NAND2X1 g117829(.A (n_16616), .B (n_16214), .Y (n_19279));
INVX1 g117848(.A (n_17504), .Y (n_16615));
NAND2X1 g117852(.A (n_16263), .B (n_16613), .Y (n_16614));
INVX1 g117857(.A (n_16611), .Y (n_18166));
INVX1 g117863(.A (n_16610), .Y (n_16930));
INVX1 g117872(.A (n_16328), .Y (n_17584));
NOR2X1 g117931(.A (n_16209), .B (n_17993), .Y (n_16606));
OR2X1 g117934(.A (n_15739), .B (n_16202), .Y (n_16605));
NAND2X1 g117949(.A (n_35077), .B (n_16297), .Y (n_17510));
NAND2X1 g117963(.A (n_10758), .B (n_16025), .Y (n_35310));
INVX2 g117975(.A (n_16599), .Y (n_20033));
NAND2X1 g117997(.A (n_9792), .B (n_33905), .Y (n_16598));
NAND2X1 g118009(.A (n_16593), .B (n_32995), .Y (n_16594));
NOR2X1 g118011(.A (n_32995), .B (n_35253), .Y (n_16921));
INVX2 g118013(.A (n_16309), .Y (n_16920));
NAND2X1 g118017(.A (n_16375), .B (n_15800), .Y (n_16918));
INVX1 g118020(.A (n_16591), .Y (n_16916));
NAND2X1 g118027(.A (n_32857), .B (n_16590), .Y (n_16915));
NOR2X1 g118031(.A (n_34934), .B (n_16015), .Y (n_16914));
NAND2X1 g118034(.A (n_16357), .B (n_15896), .Y (n_16589));
NAND2X1 g118040(.A (n_34935), .B (n_16465), .Y (n_16912));
INVX1 g118042(.A (n_17067), .Y (n_16910));
NAND2X1 g118049(.A (n_8381), .B (n_19085), .Y (n_18684));
NAND2X1 g118063(.A (n_16331), .B (n_16197), .Y (n_16907));
NAND2X2 g118096(.A (n_9742), .B (n_16194), .Y (n_17549));
INVX1 g118098(.A (n_16301), .Y (n_16901));
NAND2X1 g118110(.A (n_9628), .B (n_15881), .Y (n_17576));
NAND2X1 g118114(.A (n_16585), .B (n_15801), .Y (n_16586));
INVX1 g118124(.A (n_16292), .Y (n_16900));
AND2X1 g118149(.A (n_16046), .B (n_32411), .Y (n_16584));
NAND2X2 g118164(.A (n_35864), .B (n_16800), .Y (n_18074));
NOR2X1 g118176(.A (n_16934), .B (n_16243), .Y (n_16892));
AND2X1 g118180(.A (n_16582), .B (n_11047), .Y (n_16583));
OR2X1 g118206(.A (n_10317), .B (n_32535), .Y (n_16580));
NAND2X1 g118212(.A (n_16577), .B (n_16576), .Y (n_16578));
NAND2X1 g118217(.A (n_16239), .B (n_16574), .Y (n_16575));
INVX1 g118219(.A (n_16572), .Y (n_16573));
INVX1 g118230(.A (n_16571), .Y (n_16888));
INVX1 g118233(.A (n_16570), .Y (n_16886));
INVX1 g118244(.A (n_16568), .Y (n_17585));
INVX1 g118246(.A (n_34546), .Y (n_16567));
INVX1 g118250(.A (n_16278), .Y (n_17568));
INVX1 g118254(.A (n_16566), .Y (n_18101));
NAND2X1 g118257(.A (n_9333), .B (n_16210), .Y (n_18161));
INVX1 g118269(.A (n_34064), .Y (n_18104));
NOR2X1 g118278(.A (n_35555), .B (n_15878), .Y (n_16565));
NOR2X1 g118283(.A (n_16286), .B (n_16054), .Y (n_16564));
NOR2X1 g118286(.A (n_16562), .B (n_16060), .Y (n_16563));
OR2X1 g118308(.A (n_16582), .B (n_16560), .Y (n_16561));
NAND2X2 g118345(.A (n_34741), .B (n_17317), .Y (n_16559));
NAND2X1 g118349(.A (n_34740), .B (n_35059), .Y (n_16558));
NAND2X1 g118363(.A (n_16613), .B (n_17482), .Y (n_16557));
OAI22X1 g118535(.A0 (n_33586), .A1 (n_16150), .B0 (n_16114), .B1(n_15864), .Y (n_16556));
OAI22X1 g118544(.A0 (n_3973), .A1 (n_16415), .B0 (n_16002), .B1(n_15864), .Y (n_16555));
OAI21X1 g118561(.A0 (n_16004), .A1 (n_31647), .B0 (n_3905), .Y(n_16553));
OAI21X1 g118563(.A0 (n_15810), .A1 (n_16552), .B0 (n_16234), .Y(n_16876));
OAI22X1 g118567(.A0 (n_15859), .A1 (n_34188), .B0 (n_4170), .B1(n_7062), .Y (n_16551));
MX2X1 g118568(.A (n_6375), .B (n_16254), .S0 (n_31490), .Y (n_16550));
MX2X1 g118570(.A (n_6292), .B (n_16266), .S0 (n_30702), .Y (n_16549));
XOR2X1 g118606(.A (n_20572), .B (n_17284), .Y (n_17623));
INVX1 g118614(.A (n_17591), .Y (n_16548));
NAND2X1 g118713(.A (n_16546), .B (n_32428), .Y (n_16547));
INVX1 g118714(.A (n_16543), .Y (n_16544));
NOR2X1 g118716(.A (n_17273), .B (n_32428), .Y (n_18041));
INVX1 g118740(.A (n_16542), .Y (n_16867));
INVX1 g118741(.A (n_16542), .Y (n_16541));
CLKBUFX1 g118754(.A (n_16540), .Y (n_17320));
NAND2X2 g118765(.A (n_17262), .B (n_16158), .Y (n_18012));
INVX1 g118768(.A (n_16539), .Y (n_16864));
AND2X1 g118771(.A (n_16181), .B (n_16275), .Y (n_18057));
NOR2X1 g118789(.A (n_17474), .B (n_35824), .Y (n_16537));
NAND2X1 g118790(.A (n_10669), .B (n_16518), .Y (n_16535));
NAND2X1 g118800(.A (n_15875), .B (n_32794), .Y (n_16532));
INVX1 g118804(.A (n_16530), .Y (n_16531));
NAND2X1 g118808(.A (n_16552), .B (n_17797), .Y (n_16529));
NAND2X1 g118825(.A (n_15825), .B (n_18909), .Y (n_16528));
NAND2X1 g118834(.A (n_16829), .B (n_16120), .Y (n_18038));
INVX2 g118844(.A (n_16526), .Y (n_17372));
INVX2 g118860(.A (n_16524), .Y (n_17384));
INVX1 g118872(.A (n_21149), .Y (n_16856));
NAND2X1 g118905(.A (n_16005), .B (n_15850), .Y (n_16853));
NAND2X1 g118920(.A (n_16115), .B (n_15850), .Y (n_16851));
NAND2X1 g118925(.A (n_9738), .B (n_16511), .Y (n_16522));
INVX1 g118936(.A (n_16521), .Y (n_16849));
INVX1 g118939(.A (n_16249), .Y (n_16847));
NOR2X1 g118973(.A (n_10669), .B (n_16518), .Y (n_16519));
CLKBUFX1 gbuf_d_396(.A(n_15976), .Y(d_out_396));
CLKBUFX1 gbuf_q_396(.A(q_in_396), .Y(P3_IR[24]));
NAND2X2 g119016(.A (n_9714), .B (n_15995), .Y (n_17343));
CLKBUFX1 g119026(.A (n_16514), .Y (n_21395));
NAND2X1 g119045(.A (n_16251), .B (n_16120), .Y (n_17878));
NAND2X1 g119048(.A (n_35245), .B (n_16511), .Y (n_32839));
INVX1 g119056(.A (n_16510), .Y (n_16826));
NAND2X1 g119058(.A (n_9700), .B (n_15868), .Y (n_18018));
NAND2X1 g119084(.A (n_12002), .B (n_16505), .Y (n_17918));
INVX1 g119128(.A (n_16231), .Y (n_16824));
NAND2X1 g119154(.A (n_16501), .B (n_16154), .Y (n_17885));
NAND2X1 g119163(.A (n_9785), .B (n_16501), .Y (n_16502));
INVX1 g119168(.A (n_17311), .Y (n_16500));
NAND2X1 g119180(.A (n_32356), .B (n_16061), .Y (n_16497));
AND2X1 g119194(.A (n_16339), .B (n_18909), .Y (n_16496));
NOR2X1 g119226(.A (n_15819), .B (n_16518), .Y (n_16495));
AND2X1 g119231(.A (n_15875), .B (n_18909), .Y (n_16494));
INVX1 g119267(.A (n_16488), .Y (n_16817));
INVX1 g119330(.A (n_16219), .Y (n_17398));
INVX1 g119364(.A (n_16481), .Y (n_19179));
INVX1 g119398(.A (n_16477), .Y (n_16810));
INVX1 g119419(.A (n_34357), .Y (n_16808));
INVX1 g119420(.A (n_34357), .Y (n_16475));
INVX1 g119450(.A (n_17473), .Y (n_18005));
CLKBUFX1 g119500(.A (n_18000), .Y (n_17451));
INVX1 g119507(.A (n_16202), .Y (n_16804));
CLKBUFX1 g119518(.A (n_16469), .Y (n_19071));
INVX2 g119526(.A (n_16468), .Y (n_17732));
INVX1 g119527(.A (n_16468), .Y (n_32602));
INVX1 g119533(.A (n_16929), .Y (n_16801));
INVX2 g119541(.A (n_18532), .Y (n_16800));
INVX1 g119579(.A (n_16197), .Y (n_16799));
INVX1 g119601(.A (n_20235), .Y (n_16798));
INVX1 g119609(.A (n_16465), .Y (n_18833));
AND2X1 g119721(.A (n_16460), .B (n_17150), .Y (n_18437));
OR2X1 g119722(.A (n_16460), .B (n_17150), .Y (n_17818));
OR2X1 g119723(.A (n_16184), .B (n_16457), .Y (n_16459));
NAND2X1 g119725(.A (n_16184), .B (n_16457), .Y (n_16458));
NAND2X1 g119726(.A (n_11333), .B (n_17178), .Y (n_16456));
NAND2X1 g119727(.A (n_16778), .B (n_16734), .Y (n_16455));
NOR2X1 g119729(.A (n_16768), .B (n_16454), .Y (n_17860));
NAND2X1 g119730(.A (n_16768), .B (n_16454), .Y (n_18421));
NAND2X1 g119731(.A (n_16176), .B (n_15838), .Y (n_18163));
NOR2X1 g119732(.A (n_16452), .B (n_16451), .Y (n_16871));
NAND2X1 g119733(.A (n_16452), .B (n_16451), .Y (n_16872));
INVX1 g119738(.A (n_16450), .Y (n_17786));
INVX1 g119750(.A (n_16448), .Y (n_19790));
NAND2X1 g119758(.A (n_16131), .B (n_16446), .Y (n_35896));
INVX1 g119762(.A (n_16820), .Y (n_16786));
NAND2X2 g119782(.A (n_9722), .B (n_15949), .Y (n_16785));
INVX1 g119793(.A (n_16444), .Y (n_16783));
NAND2X1 g119796(.A (n_16748), .B (n_16428), .Y (n_18395));
NOR2X1 g119800(.A (n_9198), .B (n_16434), .Y (n_17745));
AND2X1 g119802(.A (n_16167), .B (n_16427), .Y (n_19031));
OR2X1 g119823(.A (n_16442), .B (n_16172), .Y (n_16443));
INVX1 g119825(.A (n_17863), .Y (n_16440));
NOR2X1 g119831(.A (n_9745), .B (n_17139), .Y (n_16439));
INVX1 g119832(.A (n_17861), .Y (n_16438));
NAND2X1 g119841(.A (n_16188), .B (n_16130), .Y (n_17226));
INVX1 g119843(.A (n_18667), .Y (n_16774));
NAND2X1 g119847(.A (n_11246), .B (n_16130), .Y (n_16773));
INVX1 g119848(.A (n_17841), .Y (n_16436));
NAND2X1 g119851(.A (n_16137), .B (n_9746), .Y (n_16772));
NOR2X1 g119856(.A (n_16435), .B (n_16434), .Y (n_19225));
NAND2X2 g119859(.A (n_32582), .B (n_16186), .Y (n_16771));
NOR2X1 g119866(.A (n_16182), .B (n_15948), .Y (n_17249));
INVX1 g119867(.A (n_16835), .Y (n_16433));
NAND2X1 g119869(.A (n_10270), .B (n_16172), .Y (n_17843));
OR2X1 g119870(.A (n_9722), .B (n_15950), .Y (n_17847));
INVX1 g119873(.A (n_16845), .Y (n_16765));
NAND2X1 g119875(.A (n_16163), .B (n_19471), .Y (n_17846));
NAND2X2 g119885(.A (n_16754), .B (n_19474), .Y (n_19186));
INVX1 g119895(.A (n_16168), .Y (n_16764));
INVX1 g119898(.A (n_16166), .Y (n_17207));
INVX1 g119903(.A (n_16430), .Y (n_17206));
NAND2X1 g119907(.A (n_16428), .B (n_16429), .Y (n_16761));
NAND2X1 g119910(.A (n_16161), .B (n_15767), .Y (n_32362));
NAND2X1 g119915(.A (n_10666), .B (n_16427), .Y (n_16759));
NAND2X2 g119927(.A (n_11555), .B (n_15950), .Y (n_18969));
INVX1 g119933(.A (n_16425), .Y (n_16757));
INVX1 g119937(.A (n_17233), .Y (n_16755));
NOR2X1 g119943(.A (n_16452), .B (n_16423), .Y (n_16424));
AND2X1 g119970(.A (n_16165), .B (n_16138), .Y (n_16746));
NAND2X1 g119971(.A (n_10497), .B (n_16421), .Y (n_18428));
OR2X1 g119973(.A (n_8737), .B (n_16136), .Y (n_17526));
NAND2X1 g119986(.A (n_16750), .B (n_16420), .Y (n_18981));
INVX1 g119990(.A (n_34720), .Y (n_16743));
NAND2X1 g119994(.A (n_16419), .B (n_16134), .Y (n_17222));
CLKBUFX1 gbuf_d_397(.A(n_15969), .Y(d_out_397));
CLKBUFX1 gbuf_q_397(.A(q_in_397), .Y(P1_IR[30]));
CLKBUFX1 gbuf_d_398(.A(n_15974), .Y(d_out_398));
CLKBUFX1 gbuf_q_398(.A(q_in_398), .Y(P3_IR[30]));
CLKBUFX1 gbuf_d_399(.A(n_15972), .Y(d_out_399));
CLKBUFX1 gbuf_q_399(.A(q_in_399), .Y(P1_IR[23]));
CLKBUFX1 gbuf_d_400(.A(n_15982), .Y(d_out_400));
CLKBUFX1 gbuf_q_400(.A(q_in_400), .Y(P1_IR[31]));
CLKBUFX1 gbuf_d_401(.A(n_15988), .Y(d_out_401));
CLKBUFX1 gbuf_q_401(.A(q_in_401), .Y(P2_IR[28]));
INVX1 g120202(.A (n_18145), .Y (n_16728));
CLKBUFX1 gbuf_d_402(.A(n_15980), .Y(d_out_402));
CLKBUFX1 gbuf_q_402(.A(q_in_402), .Y(P3_IR[20]));
INVX1 g120212(.A (n_16181), .Y (n_18997));
CLKBUFX1 gbuf_d_403(.A(n_15983), .Y(d_out_403));
CLKBUFX1 gbuf_q_403(.A(q_in_403), .Y(n_1964));
INVX1 g120222(.A (n_17260), .Y (n_17647));
CLKBUFX1 gbuf_d_404(.A(n_15973), .Y(d_out_404));
CLKBUFX1 gbuf_q_404(.A(q_in_404), .Y(P1_IR[20]));
INVX1 g120260(.A (n_16417), .Y (n_18379));
INVX1 g120268(.A (n_16505), .Y (n_17814));
OAI22X1 g120292(.A0 (n_6256), .A1 (n_16415), .B0 (n_15830), .B1(n_15484), .Y (n_16416));
OAI22X1 g120355(.A0 (n_15828), .A1 (n_34188), .B0 (n_5874), .B1(n_7062), .Y (n_16414));
CLKBUFX1 gbuf_d_405(.A(n_15979), .Y(d_out_405));
CLKBUFX1 gbuf_q_405(.A(q_in_405), .Y(P3_IR[21]));
INVX1 g120431(.A (n_16745), .Y (n_17174));
INVX2 g120437(.A (n_16747), .Y (n_17715));
INVX1 g120447(.A (n_16407), .Y (n_18917));
INVX1 g120455(.A (n_16406), .Y (n_18288));
INVX1 g120491(.A (n_17592), .Y (n_17133));
INVX1 g120509(.A (n_17186), .Y (n_17678));
CLKBUFX1 g120529(.A (n_15955), .Y (n_17130));
INVX1 g120584(.A (n_16731), .Y (n_23778));
INVX1 g120589(.A (n_18275), .Y (n_16707));
CLKBUFX1 gbuf_d_406(.A(n_15977), .Y(d_out_406));
CLKBUFX1 gbuf_q_406(.A(q_in_406), .Y(P3_IR[22]));
INVX1 g120155(.A (n_16117), .Y (n_17830));
INVX1 g120144(.A (n_16392), .Y (n_17831));
NOR2X1 g115824(.A (n_16546), .B (n_16113), .Y (n_16701));
NOR2X1 g116347(.A (n_16098), .B (n_16391), .Y (n_16696));
NOR2X1 g116524(.A (n_16091), .B (n_16391), .Y (n_16683));
NAND2X1 g116558(.A (n_16699), .B (n_16390), .Y (n_20605));
INVX1 g116649(.A (n_17612), .Y (n_16389));
NAND2X1 g116658(.A (n_16387), .B (n_17614), .Y (n_16388));
NAND2X1 g116736(.A (n_16386), .B (n_16390), .Y (n_17086));
INVX1 g116751(.A (n_16385), .Y (n_16673));
NAND2X1 g116773(.A (n_16390), .B (n_16387), .Y (n_16672));
NAND2X1 g116778(.A (n_17033), .B (n_16386), .Y (n_16671));
NAND2X1 g116783(.A (n_17033), .B (n_16678), .Y (n_17085));
OAI21X1 g117195(.A0 (n_16878), .A1 (n_16060), .B0 (n_15902), .Y(n_17608));
AND2X1 g117334(.A (n_17968), .B (n_16349), .Y (n_16383));
NAND2X1 g117337(.A (n_17968), .B (n_16381), .Y (n_16382));
NAND2X1 g117338(.A (n_17968), .B (n_16379), .Y (n_16380));
NAND2X1 g117339(.A (n_35744), .B (n_16381), .Y (n_16378));
NAND2X1 g117343(.A (n_35816), .B (n_16379), .Y (n_16377));
INVX2 g117368(.A (n_16376), .Y (n_17058));
NOR2X1 g117371(.A (n_16375), .B (n_16365), .Y (n_17607));
NAND2X2 g117372(.A (n_16026), .B (n_9755), .Y (n_17545));
NAND2X1 g117376(.A (n_33999), .B (n_15798), .Y (n_16653));
INVX1 g117377(.A (n_16374), .Y (n_17026));
NOR2X1 g117382(.A (n_10314), .B (n_32496), .Y (n_16373));
INVX1 g117400(.A (n_16685), .Y (n_16650));
NAND2X1 g117407(.A (n_9962), .B (n_16320), .Y (n_16369));
INVX1 g117411(.A (n_16677), .Y (n_16368));
NAND2X1 g117414(.A (n_35713), .B (n_16027), .Y (n_32503));
INVX2 g117417(.A (n_16367), .Y (n_16647));
NAND2X1 g117421(.A (n_9336), .B (n_16317), .Y (n_16366));
NAND2X1 g117422(.A (n_16375), .B (n_16365), .Y (n_17605));
NAND2X2 g117423(.A (n_9706), .B (n_32489), .Y (n_17606));
INVX1 g117438(.A (n_16363), .Y (n_16364));
INVX1 g117446(.A (n_16361), .Y (n_16641));
NAND2X1 g117467(.A (n_12289), .B (n_16322), .Y (n_16360));
INVX2 g117472(.A (n_16101), .Y (n_17024));
INVX1 g117482(.A (n_16359), .Y (n_16635));
NAND2X2 g117491(.A (n_16357), .B (n_16034), .Y (n_17022));
NAND2X1 g117493(.A (n_8381), .B (n_16031), .Y (n_18644));
INVX1 g117517(.A (n_16355), .Y (n_16631));
INVX2 g117525(.A (n_16354), .Y (n_16629));
NAND2X1 g117528(.A (n_8788), .B (n_16353), .Y (n_17603));
NAND2X1 g117535(.A (n_16291), .B (n_16289), .Y (n_21528));
NAND2X1 g117536(.A (n_16079), .B (n_15889), .Y (n_32862));
INVX1 g117543(.A (n_16099), .Y (n_16628));
NAND2X2 g117550(.A (n_8851), .B (n_16290), .Y (n_16626));
NAND2X2 g117559(.A (n_9322), .B (n_16299), .Y (n_17023));
INVX2 g117567(.A (n_16351), .Y (n_17604));
NAND2X1 g117599(.A (n_35479), .B (n_16349), .Y (n_16350));
NAND2X1 g117601(.A (n_25599), .B (n_16381), .Y (n_16348));
NAND2X1 g117614(.A (n_18533), .B (n_16349), .Y (n_16347));
NAND2X1 g117618(.A (n_35540), .B (n_16379), .Y (n_16346));
NAND2X1 g117628(.A (n_35578), .B (n_16381), .Y (n_16344));
NAND2X1 g117633(.A (n_18533), .B (n_16379), .Y (n_16342));
AND2X1 g117657(.A (n_16694), .B (n_16663), .Y (n_16341));
INVX1 g117698(.A (n_17081), .Y (n_16621));
NAND2X2 g117742(.A (n_16337), .B (n_16336), .Y (n_16338));
NAND2X1 g117753(.A (n_34934), .B (n_16016), .Y (n_17021));
NAND2X1 g117792(.A (n_16048), .B (n_32868), .Y (n_16334));
NAND2X1 g117849(.A (n_8517), .B (n_16296), .Y (n_17504));
NAND2X2 g117854(.A (n_16331), .B (n_33985), .Y (n_16612));
INVX1 g117858(.A (n_33977), .Y (n_16611));
INVX1 g117864(.A (n_16666), .Y (n_16610));
NAND2X1 g117873(.A (n_34580), .B (n_35849), .Y (n_16328));
INVX1 g120179(.A (n_16339), .Y (n_16327));
INVX1 g117902(.A (n_16095), .Y (n_16609));
INVX1 g117908(.A (n_17614), .Y (n_16326));
INVX1 g117920(.A (n_16325), .Y (n_16607));
NOR2X1 g117940(.A (n_34934), .B (n_35110), .Y (n_32976));
INVX1 g117942(.A (n_16324), .Y (n_17015));
NAND2X1 g117945(.A (n_15937), .B (n_16322), .Y (n_16323));
NAND2X1 g117947(.A (n_16320), .B (n_16318), .Y (n_16321));
NAND2X1 g117950(.A (n_16084), .B (n_16318), .Y (n_16319));
INVX1 g117959(.A (n_16090), .Y (n_16602));
INVX2 g117968(.A (n_16315), .Y (n_17051));
NAND2X2 g117970(.A (n_16103), .B (n_32489), .Y (n_17057));
NAND2X2 g117971(.A (n_32500), .B (n_9706), .Y (n_18170));
INVX1 g117977(.A (n_16312), .Y (n_16599));
INVX2 g117981(.A (n_16086), .Y (n_17595));
INVX2 g117983(.A (n_16085), .Y (n_17056));
NAND2X2 g118014(.A (n_35214), .B (n_34163), .Y (n_16309));
NAND2X2 g118021(.A (n_9274), .B (n_16365), .Y (n_16591));
NAND2X1 g118022(.A (n_32858), .B (n_15894), .Y (n_18687));
NAND2X1 g118043(.A (n_8697), .B (n_16034), .Y (n_17067));
INVX1 g118044(.A (n_16305), .Y (n_16306));
NAND2X1 g118064(.A (n_33980), .B (n_33985), .Y (n_18682));
NAND2X1 g118099(.A (n_9322), .B (n_15897), .Y (n_16301));
NAND2X1 g118103(.A (n_8850), .B (n_16299), .Y (n_18093));
NAND2X1 g118109(.A (n_16297), .B (n_16296), .Y (n_16587));
NOR2X1 g118111(.A (n_16096), .B (n_16294), .Y (n_16295));
NAND2X1 g118115(.A (n_35675), .B (n_16293), .Y (n_35951));
NAND2X1 g118116(.A (n_16353), .B (n_35423), .Y (n_17073));
NAND2X1 g118125(.A (n_16291), .B (n_16290), .Y (n_16292));
NAND2X1 g118126(.A (n_8551), .B (n_16289), .Y (n_17064));
NAND2X1 g118141(.A (n_15911), .B (n_16694), .Y (n_16288));
AND2X1 g118162(.A (n_17013), .B (n_16336), .Y (n_18602));
NAND2X2 g118183(.A (n_16286), .B (n_16076), .Y (n_17076));
NAND2X1 g118198(.A (n_8356), .B (n_15889), .Y (n_17063));
NAND2X1 g118218(.A (n_16100), .B (n_16031), .Y (n_18685));
NOR2X1 g118220(.A (n_16052), .B (n_16285), .Y (n_16572));
NAND2X1 g118231(.A (n_16279), .B (n_16284), .Y (n_16571));
NAND2X1 g118234(.A (n_16574), .B (n_16613), .Y (n_16570));
INVX1 g118237(.A (n_17028), .Y (n_16283));
INVX1 g118241(.A (n_16281), .Y (n_32878));
NAND2X1 g118245(.A (n_34981), .B (n_16279), .Y (n_16568));
NAND2X1 g118251(.A (n_16047), .B (n_16044), .Y (n_16278));
NOR2X1 g118255(.A (n_35215), .B (n_34163), .Y (n_16566));
OAI22X1 g118559(.A0 (n_6069), .A1 (n_31105), .B0 (n_15860), .B1(n_15981), .Y (n_16277));
AOI22X1 g118576(.A0 (n_11249), .A1 (n_16275), .B0 (n_9640), .B1(n_16273), .Y (n_16276));
OAI22X1 g118596(.A0 (n_10303), .A1 (n_9640), .B0 (n_16275), .B1(n_16273), .Y (n_16274));
OAI22X1 g118597(.A0 (n_10303), .A1 (n_16275), .B0 (n_12827), .B1(n_16273), .Y (n_16272));
INVX1 g118610(.A (n_16269), .Y (n_16268));
INVX4 g120173(.A (n_16191), .Y (n_18561));
INVX1 g118703(.A (n_16267), .Y (n_16922));
INVX2 g118707(.A (n_16072), .Y (n_16944));
NAND2X1 g118715(.A (n_17630), .B (n_32426), .Y (n_16543));
NAND2X1 g118742(.A (n_16266), .B (n_16230), .Y (n_16542));
NAND2X1 g118755(.A (n_9714), .B (n_16257), .Y (n_16540));
NAND2X1 g118769(.A (n_16068), .B (n_15787), .Y (n_16539));
INVX1 g118773(.A (n_16265), .Y (n_16538));
INVX1 g118791(.A (n_16069), .Y (n_16946));
INVX1 g118794(.A (n_16261), .Y (n_16533));
NAND2X1 g118803(.A (n_16257), .B (n_15733), .Y (n_17922));
INVX1 g118805(.A (n_16260), .Y (n_16530));
NAND2X1 g118828(.A (n_16068), .B (n_16257), .Y (n_16258));
INVX1 g118829(.A (n_16255), .Y (n_16256));
NAND2X2 g118846(.A (n_15984), .B (n_16253), .Y (n_16526));
NAND2X2 g118855(.A (n_16253), .B (n_16254), .Y (n_33007));
INVX1 g118861(.A (n_16063), .Y (n_16524));
INVX1 g118873(.A (n_16252), .Y (n_21149));
NAND2X1 g118929(.A (n_16251), .B (n_16117), .Y (n_16958));
INVX1 g118931(.A (n_16250), .Y (n_18560));
NAND2X1 g118937(.A (n_16040), .B (n_35623), .Y (n_16521));
INVX2 g118974(.A (n_16245), .Y (n_17075));
NAND2X2 g119002(.A (n_9700), .B (n_16417), .Y (n_16517));
NAND2X1 g119007(.A (n_16064), .B (n_16257), .Y (n_18709));
INVX1 g119021(.A (n_16243), .Y (n_17928));
INVX1 g119022(.A (n_16243), .Y (n_16242));
NOR2X1 g119027(.A (n_10275), .B (n_15784), .Y (n_16514));
INVX1 g119028(.A (n_16241), .Y (n_16955));
INVX1 g119036(.A (n_16619), .Y (n_16512));
NAND2X1 g119057(.A (n_9036), .B (n_15989), .Y (n_16510));
NAND2X1 g119059(.A (n_11010), .B (n_16417), .Y (n_17312));
INVX1 g119074(.A (n_16238), .Y (n_16506));
NAND2X1 g119077(.A (n_11401), .B (n_32426), .Y (n_16237));
INVX1 g119086(.A (n_16043), .Y (n_16932));
INVX1 g119119(.A (n_16041), .Y (n_16504));
INVX1 g119124(.A (n_17330), .Y (n_32901));
NAND2X1 g119126(.A (n_10326), .B (n_15819), .Y (n_17298));
NAND2X1 g119129(.A (n_10274), .B (n_15784), .Y (n_16231));
INVX1 g119148(.A (n_16228), .Y (n_16229));
NAND2X2 g119169(.A (n_10322), .B (n_15992), .Y (n_17311));
NAND2X1 g119174(.A (n_32344), .B (n_15998), .Y (n_16499));
INVX1 g119227(.A (n_16582), .Y (n_16225));
NOR2X1 g119229(.A (n_15797), .B (n_15875), .Y (n_17335));
INVX1 g119268(.A (n_16222), .Y (n_16488));
INVX1 g119294(.A (n_16299), .Y (n_17411));
CLKBUFX1 g119299(.A (n_16936), .Y (n_17418));
INVX1 g119310(.A (n_16590), .Y (n_16486));
INVX1 g119324(.A (n_16218), .Y (n_16219));
INVX1 g119366(.A (n_16353), .Y (n_16481));
INVX1 g119372(.A (n_16616), .Y (n_17409));
INVX2 g119380(.A (n_16214), .Y (n_17399));
INVX1 g119399(.A (n_16028), .Y (n_16477));
INVX1 g119412(.A (n_34357), .Y (n_16212));
INVX1 g119451(.A (n_16210), .Y (n_17473));
INVX1 g119468(.A (n_17993), .Y (n_16474));
INVX1 g119484(.A (n_17997), .Y (n_16473));
INVX1 g119502(.A (n_16203), .Y (n_18000));
INVX1 g119519(.A (n_33905), .Y (n_16469));
NAND2X1 g119528(.A (n_33011), .B (n_33012), .Y (n_16468));
INVX1 g119534(.A (n_16199), .Y (n_16929));
INVX2 g119587(.A (n_16196), .Y (n_17413));
INVX2 g119602(.A (n_16194), .Y (n_20235));
NAND2X1 g119735(.A (n_9302), .B (n_16187), .Y (n_18353));
NAND2X1 g119740(.A (n_16011), .B (n_16171), .Y (n_16450));
NAND2X1 g119752(.A (n_9793), .B (n_15836), .Y (n_16448));
NAND2X1 g119759(.A (n_15701), .B (n_9745), .Y (n_17253));
NAND2X1 g119763(.A (n_16188), .B (n_16187), .Y (n_16820));
NAND2X1 g119764(.A (n_35311), .B (n_33964), .Y (n_17221));
NAND2X1 g119786(.A (n_16186), .B (n_15958), .Y (n_16445));
NAND2X1 g119794(.A (n_35321), .B (n_33964), .Y (n_16444));
OR2X1 g119818(.A (n_11057), .B (n_16172), .Y (n_18638));
NAND2X1 g119824(.A (n_11333), .B (n_15962), .Y (n_17591));
NOR2X1 g119826(.A (n_16184), .B (n_16183), .Y (n_17863));
NAND2X1 g119830(.A (n_9474), .B (n_16183), .Y (n_17864));
NOR2X1 g119833(.A (n_16182), .B (n_16173), .Y (n_17861));
INVX1 g119835(.A (n_16180), .Y (n_18435));
NAND2X2 g119844(.A (n_16012), .B (n_15955), .Y (n_18667));
NOR2X1 g119849(.A (n_35311), .B (n_33964), .Y (n_17841));
INVX1 g119854(.A (n_18061), .Y (n_16178));
NAND2X1 g119863(.A (n_16176), .B (n_16777), .Y (n_16177));
NOR2X1 g119864(.A (n_16174), .B (n_16173), .Y (n_17248));
NOR2X1 g119868(.A (n_10270), .B (n_16172), .Y (n_16835));
NAND2X1 g119871(.A (n_9722), .B (n_15950), .Y (n_18091));
NAND2X2 g119874(.A (n_9281), .B (n_16162), .Y (n_16845));
NAND2X1 g119876(.A (n_10718), .B (n_16171), .Y (n_17300));
INVX1 g119878(.A (n_16170), .Y (n_16841));
INVX1 g119882(.A (n_16842), .Y (n_16169));
NAND2X1 g119896(.A (n_16167), .B (n_15966), .Y (n_16168));
NAND2X1 g119899(.A (n_16165), .B (n_15965), .Y (n_16166));
NAND2X1 g119904(.A (n_10497), .B (n_16160), .Y (n_16430));
CLKBUFX1 g119908(.A (n_35000), .Y (n_17743));
INVX2 g119925(.A (n_16164), .Y (n_17240));
INVX1 g119929(.A (n_16843), .Y (n_18433));
NAND2X1 g119934(.A (n_16163), .B (n_16162), .Y (n_16425));
NAND2X2 g119938(.A (n_10717), .B (n_15952), .Y (n_17233));
NAND2X1 g119942(.A (n_15705), .B (n_16008), .Y (n_17767));
NAND2X1 g119953(.A (n_15701), .B (n_9746), .Y (n_33051));
INVX1 g120223(.A (n_16158), .Y (n_17260));
CLKBUFX1 gbuf_d_407(.A(n_15856), .Y(d_out_407));
CLKBUFX1 gbuf_q_407(.A(q_in_407), .Y(P1_IR[22]));
INVX1 g120164(.A (n_19766), .Y (n_19005));
CLKBUFX1 gbuf_d_408(.A(n_15863), .Y(d_out_408));
CLKBUFX1 gbuf_q_408(.A(q_in_408), .Y(P2_IR[23]));
CLKBUFX1 gbuf_d_409(.A(n_15862), .Y(d_out_409));
CLKBUFX1 gbuf_q_409(.A(q_in_409), .Y(P2_IR[21]));
CLKBUFX1 gbuf_d_410(.A(n_15855), .Y(d_out_410));
CLKBUFX1 gbuf_q_410(.A(q_in_410), .Y(P1_IR[24]));
INVX1 g120233(.A (n_17259), .Y (n_17794));
CLKBUFX1 g120243(.A (n_16501), .Y (n_16837));
CLKBUFX1 g120252(.A (n_16154), .Y (n_16836));
INVX2 g120261(.A (n_15868), .Y (n_16417));
OAI22X1 g120290(.A0 (n_4006), .A1 (n_16150), .B0 (n_15762), .B1(n_15864), .Y (n_16152));
OAI22X1 g120301(.A0 (n_6342), .A1 (n_16150), .B0 (n_15967), .B1(n_15864), .Y (n_16151));
INVX1 g120311(.A (n_16148), .Y (n_16149));
MX2X1 g120352(.A (n_4990), .B (n_15960), .S0 (n_15643), .Y (n_16147));
MX2X1 g120378(.A (n_6180), .B (n_15947), .S0 (n_15968), .Y (n_16146));
OAI22X1 g120385(.A0 (n_15951), .A1 (n_15484), .B0 (n_34947), .B1(n_31328), .Y (n_16145));
INVX2 g120393(.A (n_16423), .Y (n_17172));
INVX1 g120401(.A (n_17150), .Y (n_16411));
INVX1 g120432(.A (n_16428), .Y (n_16745));
INVX2 g120433(.A (n_16428), .Y (n_16140));
INVX1 g120438(.A (n_16427), .Y (n_16747));
INVX1 g120448(.A (n_16138), .Y (n_16407));
INVX1 g120456(.A (n_16421), .Y (n_16406));
INVX1 g120483(.A (n_16137), .Y (n_16738));
CLKBUFX1 g120492(.A (n_16136), .Y (n_17592));
INVX1 g120503(.A (n_16457), .Y (n_16404));
INVX1 g120506(.A (n_16434), .Y (n_16135));
CLKBUFX1 g120510(.A (n_16434), .Y (n_17186));
INVX1 g120514(.A (n_16134), .Y (n_16403));
INVX1 g120525(.A (n_17139), .Y (n_16402));
INVX1 g120537(.A (n_16130), .Y (n_17131));
INVX1 g120552(.A (n_16734), .Y (n_16400));
INVX1 g120574(.A (n_16126), .Y (n_16396));
INVX1 g120585(.A (n_16451), .Y (n_16731));
INVX1 g120590(.A (n_15950), .Y (n_18275));
INVX2 g120621(.A (n_16454), .Y (n_16740));
CLKBUFX1 gbuf_d_411(.A(n_15865), .Y(d_out_411));
CLKBUFX1 gbuf_q_411(.A(q_in_411), .Y(P2_IR[24]));
INVX1 g120145(.A (n_16511), .Y (n_16392));
INVX1 g120157(.A (n_16117), .Y (n_16120));
CLKBUFX1 gbuf_d_412(.A(n_15778), .Y(d_out_412));
CLKBUFX1 gbuf_q_412(.A(q_in_412), .Y(P3_IR[23]));
INVX1 g120135(.A (n_15943), .Y (n_17289));
NAND2X1 g116650(.A (n_17036), .B (n_17025), .Y (n_17612));
NAND2X1 g116752(.A (n_16690), .B (n_17036), .Y (n_16385));
INVX1 g120066(.A (n_16114), .Y (n_16115));
INVX1 g117331(.A (n_16113), .Y (n_17628));
NAND2X1 g117369(.A (n_16112), .B (n_15884), .Y (n_16376));
INVX1 g117378(.A (n_15940), .Y (n_16374));
INVX1 g117388(.A (n_34171), .Y (n_16371));
INVX1 g117392(.A (n_34004), .Y (n_16109));
INVX2 g117393(.A (n_34004), .Y (n_18088));
CLKBUFX3 g117397(.A (n_16107), .Y (n_17089));
NAND2X2 g117401(.A (n_8479), .B (n_16379), .Y (n_16685));
INVX1 g117405(.A (n_15936), .Y (n_16370));
INVX1 g117409(.A (n_16105), .Y (n_17552));
INVX1 g117412(.A (n_16391), .Y (n_16677));
NAND2X1 g117418(.A (n_8859), .B (n_16087), .Y (n_16367));
NOR2X1 g117439(.A (n_9269), .B (n_16381), .Y (n_16363));
NAND2X2 g117442(.A (n_32501), .B (n_16103), .Y (n_35352));
NAND2X1 g117447(.A (n_16102), .B (n_16089), .Y (n_16361));
NAND2X1 g117473(.A (n_8697), .B (n_15896), .Y (n_16101));
NAND2X1 g117483(.A (n_32859), .B (n_15894), .Y (n_16359));
INVX1 g117486(.A (n_15935), .Y (n_16358));
NAND2X1 g117518(.A (n_16100), .B (n_15893), .Y (n_16355));
NAND2X1 g117526(.A (n_8711), .B (n_34298), .Y (n_16354));
NAND2X1 g117544(.A (n_8850), .B (n_15897), .Y (n_16099));
NAND2X2 g117568(.A (n_8513), .B (n_16083), .Y (n_16351));
INVX1 g117699(.A (n_16098), .Y (n_17081));
INVX1 g117816(.A (n_16387), .Y (n_16097));
INVX1 g120183(.A (n_16275), .Y (n_16339));
NAND2X1 g117865(.A (n_16096), .B (n_15881), .Y (n_16666));
NAND2X1 g117903(.A (n_33999), .B (n_34002), .Y (n_16095));
NAND2X1 g117921(.A (n_8799), .B (n_16379), .Y (n_16325));
NAND2X1 g117941(.A (n_33999), .B (n_15878), .Y (n_16092));
INVX1 g117943(.A (n_15932), .Y (n_16324));
INVX1 g117951(.A (n_16091), .Y (n_17080));
NAND2X1 g117960(.A (n_9755), .B (n_16089), .Y (n_16090));
NOR2X1 g117969(.A (n_35713), .B (n_16087), .Y (n_16315));
INVX1 g117978(.A (n_15930), .Y (n_16312));
NAND2X1 g117982(.A (n_11404), .B (n_15877), .Y (n_16086));
NAND2X1 g117984(.A (n_16084), .B (n_15898), .Y (n_16085));
INVX1 g118002(.A (n_15926), .Y (n_16311));
NAND2X1 g118006(.A (n_34172), .B (n_15899), .Y (n_35915));
NAND2X1 g118046(.A (n_16079), .B (n_16083), .Y (n_16305));
INVX1 g118106(.A (n_15924), .Y (n_16298));
INVX4 g120116(.A (n_15819), .Y (n_17273));
NAND2X1 g118117(.A (n_8788), .B (n_34298), .Y (n_17084));
NAND2X1 g118169(.A (n_15804), .B (n_15910), .Y (n_16080));
NOR2X1 g118197(.A (n_16079), .B (n_16083), .Y (n_17055));
NAND2X1 g118238(.A (n_16078), .B (n_16336), .Y (n_17028));
NAND2X1 g118243(.A (n_16574), .B (n_16078), .Y (n_16281));
NAND2X1 g118284(.A (n_34548), .B (n_16284), .Y (n_16075));
NAND2X1 g118287(.A (n_17018), .B (n_16664), .Y (n_18157));
NAND2X1 g118289(.A (n_16073), .B (n_17018), .Y (n_16074));
NAND2X2 g118702(.A (n_15918), .B (n_35448), .Y (n_17045));
INVX1 g118704(.A (n_15922), .Y (n_16267));
NAND2X2 g118708(.A (n_10706), .B (n_32429), .Y (n_16072));
INVX2 g118710(.A (n_16337), .Y (n_16071));
NAND2X1 g118774(.A (n_15909), .B (n_15733), .Y (n_16265));
INVX1 g118785(.A (n_15921), .Y (n_16263));
NAND2X1 g118792(.A (n_34575), .B (n_16067), .Y (n_16069));
NAND2X1 g118795(.A (n_16068), .B (n_15733), .Y (n_16261));
INVX1 g118806(.A (n_15920), .Y (n_16260));
NAND2X2 g118812(.A (n_9720), .B (n_16067), .Y (n_17482));
INVX1 g118814(.A (n_16569), .Y (n_17017));
INVX1 g118830(.A (n_16066), .Y (n_16255));
NAND2X1 g118832(.A (n_16064), .B (n_17259), .Y (n_16065));
NAND2X1 g118862(.A (n_15841), .B (n_15858), .Y (n_16063));
NAND2X1 g118874(.A (n_9749), .B (n_15663), .Y (n_16252));
NOR2X1 g118880(.A (n_17474), .B (n_17472), .Y (n_16062));
NOR2X1 g118932(.A (n_32344), .B (n_16061), .Y (n_16250));
NAND2X1 g118941(.A (n_32344), .B (n_16061), .Y (n_16249));
INVX1 g118956(.A (n_34981), .Y (n_16060));
INVX1 g118975(.A (n_15913), .Y (n_16245));
INVX1 g118977(.A (n_16693), .Y (n_16054));
INVX1 g118988(.A (n_16052), .Y (n_16950));
INVX1 g119008(.A (n_17334), .Y (n_16051));
NAND2X1 g119019(.A (n_11010), .B (n_15868), .Y (n_35175));
INVX1 g119023(.A (n_16048), .Y (n_16243));
INVX1 g119029(.A (n_16047), .Y (n_16241));
NAND2X1 g119031(.A (n_15873), .B (n_8802), .Y (n_32412));
INVX1 g119032(.A (n_34581), .Y (n_16046));
CLKBUFX1 g119037(.A (n_16044), .Y (n_16619));
NAND2X2 g119054(.A (n_35270), .B (n_11280), .Y (n_17317));
INVX1 g119064(.A (n_15907), .Y (n_16239));
NAND2X1 g119075(.A (n_33227), .B (n_16039), .Y (n_16238));
INVX1 g119080(.A (n_19974), .Y (n_16234));
NAND2X1 g119087(.A (n_9036), .B (n_35270), .Y (n_16043));
NAND2X1 g119088(.A (n_16036), .B (n_10322), .Y (n_16934));
NAND2X1 g119120(.A (n_9640), .B (n_15753), .Y (n_16041));
NAND2X1 g119125(.A (n_16040), .B (n_16039), .Y (n_17330));
NOR2X1 g119149(.A (n_10312), .B (n_15943), .Y (n_16228));
INVX1 g120175(.A (n_35622), .Y (n_16191));
NAND2X1 g119208(.A (n_16275), .B (n_16273), .Y (n_16560));
NAND2X1 g119228(.A (n_15819), .B (n_15806), .Y (n_16582));
INVX1 g119242(.A (n_16322), .Y (n_17004));
INVX1 g119256(.A (n_16320), .Y (n_16643));
NAND3X1 g119270(.A (n_15688), .B (n_15681), .C (n_6822), .Y(n_16222));
INVX1 g119300(.A (n_16034), .Y (n_16936));
INVX1 g119311(.A (n_15894), .Y (n_16590));
INVX2 g119320(.A (n_16031), .Y (n_19085));
INVX1 g119333(.A (n_15891), .Y (n_16218));
INVX1 g119381(.A (n_16290), .Y (n_16214));
NAND3X1 g119400(.A (n_15690), .B (n_15680), .C (n_6803), .Y(n_16028));
NAND3X1 g119411(.A (n_15699), .B (n_15686), .C (n_6793), .Y(n_16213));
INVX1 g119452(.A (n_16027), .Y (n_16210));
INVX1 g119460(.A (n_16026), .Y (n_16209));
INVX1 g119469(.A (n_16317), .Y (n_17993));
INVX1 g119470(.A (n_16317), .Y (n_16025));
INVX4 g119485(.A (n_16365), .Y (n_17997));
INVX1 g119503(.A (n_34163), .Y (n_16203));
INVX1 g119510(.A (n_15798), .Y (n_16202));
NAND2X2 g119535(.A (n_15541), .B (n_15779), .Y (n_16199));
INVX1 g119581(.A (n_33985), .Y (n_16197));
INVX1 g119589(.A (n_16294), .Y (n_16196));
INVX1 g119603(.A (n_16296), .Y (n_16194));
INVX1 g119604(.A (n_16296), .Y (n_35077));
INVX2 g119613(.A (n_16016), .Y (n_16465));
INVX1 g119614(.A (n_16016), .Y (n_16015));
INVX1 g119639(.A (n_16318), .Y (n_16576));
NOR2X1 g119734(.A (n_9637), .B (n_15838), .Y (n_16269));
INVX1 g120107(.A (n_15797), .Y (n_16518));
NAND2X2 g119837(.A (n_9745), .B (n_16137), .Y (n_16180));
NAND2X2 g119855(.A (n_16012), .B (n_15840), .Y (n_18061));
NAND2X1 g119879(.A (n_16011), .B (n_16007), .Y (n_16170));
NAND2X1 g119880(.A (n_16010), .B (n_16009), .Y (n_16854));
NOR2X1 g119883(.A (n_16010), .B (n_16009), .Y (n_16842));
NAND2X1 g119921(.A (n_10718), .B (n_16007), .Y (n_35949));
NAND2X1 g119926(.A (n_9327), .B (n_16009), .Y (n_16164));
NAND2X1 g119930(.A (n_9280), .B (n_15832), .Y (n_16843));
INVX1 g120062(.A (n_16004), .Y (n_16005));
INVX1 g120064(.A (n_16002), .Y (n_16003));
INVX1 g120224(.A (n_16257), .Y (n_16158));
CLKBUFX1 gbuf_d_413(.A(n_15768), .Y(d_out_413));
CLKBUFX1 gbuf_q_413(.A(q_in_413), .Y(P1_IR[21]));
CLKBUFX1 gbuf_d_414(.A(n_15772), .Y(d_out_414));
CLKBUFX1 gbuf_q_414(.A(q_in_414), .Y(P1_IR[17]));
INVX1 g120165(.A (n_15998), .Y (n_19766));
CLKBUFX1 gbuf_d_415(.A(n_15771), .Y(d_out_415));
CLKBUFX1 gbuf_q_415(.A(q_in_415), .Y(P1_IR[18]));
CLKBUFX1 gbuf_d_416(.A(n_15773), .Y(d_out_416));
CLKBUFX1 gbuf_q_416(.A(q_in_416), .Y(P1_IR[16]));
INVX1 g120204(.A (n_15997), .Y (n_18145));
INVX1 g120214(.A (n_15996), .Y (n_16181));
CLKBUFX1 gbuf_d_417(.A(n_15776), .Y(d_out_417));
CLKBUFX1 gbuf_q_417(.A(q_in_417), .Y(P1_IR[14]));
CLKBUFX1 gbuf_d_418(.A(n_15775), .Y(d_out_418));
CLKBUFX1 gbuf_q_418(.A(q_in_418), .Y(P1_IR[15]));
CLKBUFX1 gbuf_d_419(.A(n_15769), .Y(d_out_419));
CLKBUFX1 gbuf_q_419(.A(q_in_419), .Y(P1_IR[19]));
INVX1 g120226(.A (n_16257), .Y (n_15995));
INVX2 g120234(.A (n_15787), .Y (n_17259));
INVX1 g120244(.A (n_15992), .Y (n_16501));
INVX1 g120253(.A (n_15784), .Y (n_16154));
INVX1 g120270(.A (n_15989), .Y (n_16505));
OAI22X1 g120291(.A0 (n_33583), .A1 (n_16150), .B0 (n_15853), .B1(n_15484), .Y (n_15988));
NAND3X1 g120312(.A (n_15601), .B (n_15677), .C (n_15596), .Y(n_16148));
INVX1 g120314(.A (n_15984), .Y (n_15985));
MX2X1 g120330(.A (n_34396), .B (n_15844), .S0 (n_15975), .Y(n_15983));
OAI22X1 g120336(.A0 (n_4901), .A1 (n_31105), .B0 (n_15671), .B1(n_15981), .Y (n_15982));
MX2X1 g120347(.A (n_32637), .B (n_15666), .S0 (n_15975), .Y(n_15980));
MX2X1 g120348(.A (n_6527), .B (n_15839), .S0 (n_15975), .Y (n_15979));
MX2X1 g120349(.A (n_6802), .B (n_15842), .S0 (n_15975), .Y (n_15977));
MX2X1 g120351(.A (n_34119), .B (n_15843), .S0 (n_15975), .Y(n_15976));
MX2X1 g120354(.A (n_5015), .B (n_15845), .S0 (n_15975), .Y (n_15974));
MX2X1 g120372(.A (n_6348), .B (n_15833), .S0 (n_31105), .Y (n_15973));
MX2X1 g120375(.A (n_6246), .B (n_15668), .S0 (n_15968), .Y (n_15972));
MX2X1 g120377(.A (n_6231), .B (n_15831), .S0 (n_31105), .Y (n_15971));
MX2X1 g120384(.A (n_35400), .B (n_15837), .S0 (n_15968), .Y(n_15969));
NOR2X1 g120395(.A (n_15967), .B (n_8424), .Y (n_16423));
NAND2X1 g120402(.A (n_15829), .B (n_15708), .Y (n_17150));
INVX1 g120413(.A (n_15854), .Y (n_16420));
INVX2 g120421(.A (n_15852), .Y (n_19474));
INVX2 g120434(.A (n_15851), .Y (n_16428));
INVX1 g120440(.A (n_15966), .Y (n_16427));
INVX1 g120449(.A (n_15965), .Y (n_16138));
INVX1 g120457(.A (n_16160), .Y (n_16421));
NAND2X1 g120493(.A (n_15827), .B (n_15959), .Y (n_16136));
INVX2 g120498(.A (n_15962), .Y (n_17178));
INVX2 g120504(.A (n_16183), .Y (n_16457));
NAND2X1 g120511(.A (n_15960), .B (n_15959), .Y (n_16434));
INVX1 g120516(.A (n_15958), .Y (n_16134));
INVX1 g120517(.A (n_15958), .Y (n_32582));
INVX1 g120526(.A (n_33964), .Y (n_17139));
INVX1 g120531(.A (n_15955), .Y (n_16131));
INVX2 g120538(.A (n_16187), .Y (n_16130));
INVX1 g120553(.A (n_15953), .Y (n_16734));
INVX1 g120558(.A (n_15952), .Y (n_17712));
INVX1 g120576(.A (n_16171), .Y (n_16126));
OR2X1 g120586(.A (n_15951), .B (n_8424), .Y (n_16451));
INVX1 g120592(.A (n_15950), .Y (n_15949));
INVX2 g120601(.A (n_16162), .Y (n_19471));
INVX2 g120615(.A (n_16173), .Y (n_17639));
INVX1 g120616(.A (n_16173), .Y (n_15948));
NAND2X1 g120623(.A (n_15947), .B (n_15946), .Y (n_16454));
INVX2 g120146(.A (n_15945), .Y (n_16511));
CLKBUFX1 gbuf_d_420(.A(n_15729), .Y(d_out_420));
CLKBUFX1 gbuf_q_420(.A(q_in_420), .Y(P2_IR[18]));
AOI21X1 g120067(.A0 (n_15676), .A1 (datao_1[27] ), .B0 (n_15678), .Y(n_16114));
NAND2X1 g117379(.A (n_15817), .B (n_15745), .Y (n_15940));
NAND2X1 g117395(.A (n_9953), .B (n_15937), .Y (n_15938));
NAND2X1 g117398(.A (n_9269), .B (n_15929), .Y (n_16107));
NAND2X1 g117406(.A (n_8231), .B (n_15928), .Y (n_15936));
NAND2X1 g117410(.A (n_8233), .B (n_15934), .Y (n_16105));
NOR2X1 g117413(.A (n_8233), .B (n_15934), .Y (n_16391));
NAND2X1 g117487(.A (n_32334), .B (n_15802), .Y (n_15935));
NOR2X1 g117700(.A (n_8086), .B (n_15931), .Y (n_16098));
NAND2X1 g117817(.A (n_8418), .B (n_15934), .Y (n_16387));
INVX1 g117831(.A (n_34362), .Y (n_16386));
NAND2X2 g117885(.A (n_8803), .B (n_15798), .Y (n_16678));
NAND2X2 g117910(.A (n_8518), .B (n_15931), .Y (n_17614));
NAND2X1 g117944(.A (n_8526), .B (n_15878), .Y (n_15932));
NAND2X1 g117952(.A (n_8086), .B (n_15931), .Y (n_16091));
NAND2X1 g117979(.A (n_7810), .B (n_15929), .Y (n_15930));
NAND2X2 g117980(.A (n_8479), .B (n_15928), .Y (n_17615));
NAND2X2 g117985(.A (n_15820), .B (n_15937), .Y (n_16390));
NAND2X2 g118000(.A (n_15815), .B (n_15878), .Y (n_17033));
NAND2X1 g118003(.A (n_8526), .B (n_15739), .Y (n_15926));
NAND2X1 g118107(.A (n_16096), .B (n_15795), .Y (n_15924));
INVX1 g118202(.A (n_16690), .Y (n_15923));
NAND2X1 g118705(.A (n_15919), .B (n_35343), .Y (n_15922));
NAND2X2 g118712(.A (n_32430), .B (n_15807), .Y (n_16337));
NAND2X1 g118743(.A (n_15809), .B (n_15757), .Y (n_16113));
CLKBUFX1 g118775(.A (n_18824), .Y (n_19957));
NAND2X1 g118786(.A (n_10303), .B (n_34978), .Y (n_15921));
NAND2X1 g118807(.A (n_35705), .B (n_15812), .Y (n_15920));
INVX2 g118815(.A (n_15814), .Y (n_16569));
NOR2X1 g118831(.A (n_15919), .B (n_15918), .Y (n_16066));
NAND2X1 g118968(.A (n_8729), .B (n_15592), .Y (n_16279));
NAND2X1 g118976(.A (n_8625), .B (n_32431), .Y (n_15913));
INVX2 g118979(.A (n_16285), .Y (n_16693));
INVX1 g118982(.A (n_15911), .Y (n_15912));
CLKBUFX1 g118984(.A (n_15910), .Y (n_16694));
INVX1 g118989(.A (n_16076), .Y (n_16052));
NAND2X2 g119010(.A (n_15909), .B (n_15787), .Y (n_17334));
NAND2X1 g119013(.A (n_11280), .B (n_15783), .Y (n_32868));
NAND2X1 g119024(.A (n_10275), .B (n_15784), .Y (n_16048));
NAND2X1 g119030(.A (n_9652), .B (n_15785), .Y (n_16047));
NAND2X1 g119038(.A (n_15908), .B (n_15791), .Y (n_16044));
NAND2X1 g119060(.A (n_8756), .B (n_15661), .Y (n_17013));
NAND2X1 g119065(.A (n_15906), .B (n_15592), .Y (n_15907));
NOR2X1 g119066(.A (n_15906), .B (n_15797), .Y (n_17014));
INVX2 g119071(.A (n_15905), .Y (n_16286));
NAND2X1 g119076(.A (n_10706), .B (n_17630), .Y (n_15904));
CLKBUFX1 g119081(.A (n_16073), .Y (n_19974));
INVX1 g119090(.A (n_15902), .Y (n_16562));
INVX1 g119094(.A (n_15900), .Y (n_16042));
NAND2X2 g119152(.A (n_10484), .B (n_15919), .Y (n_35221));
NAND2X1 g119166(.A (n_9730), .B (n_15821), .Y (n_16613));
INVX1 g119243(.A (n_15899), .Y (n_16322));
INVX1 g119257(.A (n_15898), .Y (n_16320));
INVX2 g119292(.A (n_15897), .Y (n_16299));
INVX2 g119302(.A (n_15896), .Y (n_16034));
INVX2 g119321(.A (n_15893), .Y (n_16031));
NAND3X1 g119334(.A (n_15626), .B (n_15623), .C (n_6528), .Y(n_15891));
INVX4 g119368(.A (n_34298), .Y (n_16353));
INVX1 g119370(.A (n_16083), .Y (n_15889));
INVX1 g119374(.A (n_16083), .Y (n_16616));
INVX1 g119377(.A (n_15887), .Y (n_16289));
CLKBUFX1 g119382(.A (n_15887), .Y (n_16290));
INVX1 g119453(.A (n_16087), .Y (n_16027));
INVX2 g119461(.A (n_16089), .Y (n_16026));
INVX2 g119471(.A (n_15884), .Y (n_16317));
INVX2 g119486(.A (n_15800), .Y (n_16365));
INVX1 g119590(.A (n_15881), .Y (n_16294));
INVX2 g119605(.A (n_15793), .Y (n_16296));
INVX1 g119615(.A (n_15879), .Y (n_16016));
INVX1 g119616(.A (n_15879), .Y (n_35110));
INVX1 g119631(.A (n_15878), .Y (n_17479));
INVX1 g119640(.A (n_15877), .Y (n_16318));
INVX1 g120049(.A (n_17474), .Y (n_16857));
AOI21X1 g120063(.A0 (n_15676), .A1 (n_641), .B0 (n_15703), .Y(n_16004));
AOI21X1 g120065(.A0 (n_15676), .A1 (n_12319), .B0 (n_15702), .Y(n_16002));
INVX1 g120167(.A (n_16061), .Y (n_15998));
NAND2X2 g120159(.A (n_15709), .B (n_8150), .Y (n_16117));
CLKBUFX1 gbuf_d_421(.A(n_15714), .Y(d_out_421));
CLKBUFX1 gbuf_q_421(.A(q_in_421), .Y(P1_IR[13]));
CLKBUFX1 gbuf_d_422(.A(n_15731), .Y(d_out_422));
CLKBUFX1 gbuf_q_422(.A(q_in_422), .Y(P2_IR[16]));
CLKBUFX1 gbuf_d_423(.A(n_15732), .Y(d_out_423));
CLKBUFX1 gbuf_q_423(.A(q_in_423), .Y(P2_IR[19]));
INVX1 g120205(.A (n_15873), .Y (n_15997));
CLKBUFX1 gbuf_d_424(.A(n_15718), .Y(d_out_424));
CLKBUFX1 gbuf_q_424(.A(q_in_424), .Y(P3_IR[15]));
CLKBUFX1 gbuf_d_425(.A(n_15715), .Y(d_out_425));
CLKBUFX1 gbuf_q_425(.A(q_in_425), .Y(P3_IR[19]));
INVX1 g120215(.A (n_16067), .Y (n_15996));
INVX2 g120225(.A (n_15872), .Y (n_16257));
INVX1 g120245(.A (n_16036), .Y (n_15992));
INVX1 g120271(.A (n_35270), .Y (n_15989));
OAI22X1 g120279(.A0 (n_34485), .A1 (n_16150), .B0 (n_15674), .B1(n_15864), .Y (n_15865));
OAI22X1 g120280(.A0 (n_32641), .A1 (n_16150), .B0 (n_15672), .B1(n_15864), .Y (n_15863));
OAI22X1 g120289(.A0 (n_6467), .A1 (n_16415), .B0 (n_15766), .B1(n_3185), .Y (n_15862));
INVX1 g120308(.A (n_15860), .Y (n_15861));
NAND3X1 g120313(.A (n_15506), .B (n_15612), .C (n_15501), .Y(n_16266));
NAND3X1 g120315(.A (n_15599), .B (n_15610), .C (n_15504), .Y(n_15984));
NAND3X1 g120316(.A (n_15598), .B (n_15609), .C (n_15502), .Y(n_16254));
INVX1 g120317(.A (n_15858), .Y (n_15859));
AOI21X1 g120323(.A0 (n_6281), .A1 (n_7793), .B0 (n_15679), .Y(n_33011));
MX2X1 g120374(.A (n_35390), .B (n_15764), .S0 (n_15968), .Y(n_15856));
MX2X1 g120376(.A (n_6214), .B (n_15765), .S0 (n_31105), .Y (n_15855));
NOR2X1 g120414(.A (n_15853), .B (n_7865), .Y (n_15854));
NAND2X1 g120422(.A (n_15675), .B (n_15708), .Y (n_15852));
NAND2X2 g120435(.A (n_15850), .B (n_15761), .Y (n_15851));
NAND2X2 g120441(.A (n_15673), .B (n_15850), .Y (n_15966));
INVX1 g120450(.A (n_15849), .Y (n_15965));
INVX1 g120459(.A (n_15767), .Y (n_16160));
NAND2X1 g120500(.A (n_15845), .B (n_15959), .Y (n_15962));
NAND2X1 g120505(.A (n_15844), .B (n_15959), .Y (n_16183));
NAND2X1 g120518(.A (n_15843), .B (n_15841), .Y (n_15958));
INVX1 g120532(.A (n_15840), .Y (n_15955));
NAND2X2 g120540(.A (n_15839), .B (n_15841), .Y (n_16187));
INVX1 g120545(.A (n_15838), .Y (n_16777));
AND2X1 g120554(.A (n_15837), .B (n_15946), .Y (n_15953));
INVX1 g120559(.A (n_16009), .Y (n_15952));
INVX4 g120566(.A (n_15835), .Y (n_16172));
INVX1 g120567(.A (n_15835), .Y (n_15836));
INVX2 g120577(.A (n_16007), .Y (n_16171));
NAND2X2 g120593(.A (n_15833), .B (n_16230), .Y (n_15950));
INVX1 g120602(.A (n_15832), .Y (n_16162));
NAND2X2 g120617(.A (n_15946), .B (n_15831), .Y (n_16173));
CLKBUFX1 gbuf_d_426(.A(n_15711), .Y(d_out_426));
CLKBUFX1 gbuf_q_426(.A(q_in_426), .Y(P1_IR[6]));
INVX1 g120882(.A (n_15829), .Y (n_15830));
INVX1 g120957(.A (n_15827), .Y (n_15828));
CLKBUFX1 gbuf_d_427(.A(n_15721), .Y(d_out_427));
CLKBUFX1 gbuf_q_427(.A(q_in_427), .Y(P3_IR[16]));
CLKBUFX1 gbuf_d_428(.A(n_15712), .Y(d_out_428));
CLKBUFX1 gbuf_q_428(.A(q_in_428), .Y(P1_IR[2]));
CLKBUFX1 gbuf_d_429(.A(n_15724), .Y(d_out_429));
CLKBUFX1 gbuf_q_429(.A(q_in_429), .Y(P1_IR[4]));
NAND2X2 g120147(.A (n_15710), .B (n_8153), .Y (n_15945));
INVX2 g120083(.A (n_15825), .Y (n_17284));
CLKBUFX1 gbuf_d_430(.A(n_15728), .Y(d_out_430));
CLKBUFX1 gbuf_q_430(.A(q_in_430), .Y(P2_IR[20]));
CLKBUFX1 gbuf_d_431(.A(n_15651), .Y(d_out_431));
CLKBUFX1 gbuf_q_431(.A(q_in_431), .Y(P3_IR[9]));
INVX1 g120137(.A (n_15824), .Y (n_15943));
INVX1 g120193(.A (n_16552), .Y (n_20572));
INVX2 g120128(.A (n_17630), .Y (n_16546));
CLKBUFX3 g120185(.A (n_15821), .Y (n_16275));
NAND2X2 g117386(.A (n_8465), .B (n_34358), .Y (n_17036));
NAND2X2 g117436(.A (n_15820), .B (n_34471), .Y (n_17025));
NAND2X1 g117986(.A (n_15817), .B (n_34471), .Y (n_16699));
NAND2X2 g118203(.A (n_15815), .B (n_15739), .Y (n_16690));
NOR2X1 g120177(.A (n_15706), .B (n_7609), .Y (n_16039));
NAND2X2 g118706(.A (n_33268), .B (n_15736), .Y (n_16664));
NAND2X1 g118718(.A (n_15805), .B (n_10006), .Y (n_16574));
NAND2X1 g118776(.A (n_8801), .B (n_15663), .Y (n_18824));
NAND2X1 g118816(.A (n_8829), .B (n_15811), .Y (n_15814));
NAND2X1 g118961(.A (n_15906), .B (n_15806), .Y (n_16878));
INVX1 g118963(.A (n_16284), .Y (n_15813));
NOR2X1 g118980(.A (n_15812), .B (n_15811), .Y (n_16285));
AND2X1 g118983(.A (n_15810), .B (n_15809), .Y (n_15911));
NAND2X1 g118985(.A (n_15492), .B (n_15749), .Y (n_15910));
CLKBUFX3 g118986(.A (n_15808), .Y (n_16663));
NAND2X2 g118990(.A (n_15807), .B (n_32432), .Y (n_16076));
NAND2X2 g119061(.A (n_9278), .B (n_15752), .Y (n_16336));
NAND2X1 g119067(.A (n_9292), .B (n_15806), .Y (n_16078));
NAND2X1 g119072(.A (n_15811), .B (n_15812), .Y (n_15905));
INVX1 g119082(.A (n_15747), .Y (n_16073));
NAND2X1 g119091(.A (n_9729), .B (n_15805), .Y (n_15902));
INVX1 g119096(.A (n_15804), .Y (n_15900));
INVX1 g119236(.A (n_15937), .Y (n_16349));
INVX1 g119244(.A (n_34167), .Y (n_15899));
CLKBUFX1 g119248(.A (n_15929), .Y (n_16381));
NAND2X2 g119252(.A (n_15381), .B (n_15654), .Y (n_16379));
INVX1 g119258(.A (n_15934), .Y (n_15898));
NAND3X1 g119297(.A (n_15569), .B (n_15567), .C (n_6715), .Y(n_15897));
NAND3X1 g119304(.A (n_15563), .B (n_15545), .C (n_6721), .Y(n_15896));
INVX1 g119313(.A (n_15802), .Y (n_15894));
NAND3X1 g119323(.A (n_15561), .B (n_15559), .C (n_6712), .Y(n_15893));
NAND3X1 g119360(.A (n_15557), .B (n_15544), .C (n_6714), .Y(n_15801));
NAND3X1 g119376(.A (n_15552), .B (n_15549), .C (n_6716), .Y(n_16083));
NAND3X1 g119383(.A (n_15548), .B (n_15546), .C (n_6545), .Y(n_15887));
NAND3X1 g119454(.A (n_15537), .B (n_15534), .C (n_7438), .Y(n_16087));
NAND3X1 g119463(.A (n_15533), .B (n_15531), .C (n_7436), .Y(n_16089));
NAND3X1 g119472(.A (n_15539), .B (n_15521), .C (n_7363), .Y(n_15884));
NAND2X2 g119478(.A (n_15529), .B (n_15652), .Y (n_32501));
NAND3X1 g119487(.A (n_15528), .B (n_15526), .C (n_7440), .Y(n_15800));
NAND3X1 g119499(.A (n_15524), .B (n_15522), .C (n_7441), .Y(n_32995));
INVX1 g119591(.A (n_15795), .Y (n_15881));
NAND3X1 g119606(.A (n_15573), .B (n_6725), .C (n_15572), .Y(n_15793));
NAND3X1 g119617(.A (n_15566), .B (n_6702), .C (n_15565), .Y(n_15879));
INVX2 g119632(.A (n_15739), .Y (n_15878));
INVX1 g119641(.A (n_15931), .Y (n_15877));
INVX1 g120050(.A (n_15919), .Y (n_17474));
INVX1 g120051(.A (n_15919), .Y (n_35448));
INVX1 g120098(.A (n_16273), .Y (n_15875));
CLKBUFX1 gbuf_d_432(.A(n_15633), .Y(d_out_432));
CLKBUFX1 gbuf_q_432(.A(q_in_432), .Y(P1_IR[9]));
CLKBUFX1 gbuf_d_433(.A(n_15634), .Y(d_out_433));
CLKBUFX1 gbuf_q_433(.A(q_in_433), .Y(P1_IR[8]));
CLKBUFX1 gbuf_d_434(.A(n_15636), .Y(d_out_434));
CLKBUFX1 gbuf_q_434(.A(q_in_434), .Y(P1_IR[12]));
CLKBUFX1 gbuf_d_435(.A(n_15655), .Y(d_out_435));
CLKBUFX1 gbuf_q_435(.A(q_in_435), .Y(P2_IR[13]));
CLKBUFX1 gbuf_d_436(.A(n_15657), .Y(d_out_436));
CLKBUFX1 gbuf_q_436(.A(q_in_436), .Y(P2_IR[14]));
CLKBUFX1 gbuf_d_437(.A(n_15659), .Y(d_out_437));
CLKBUFX1 gbuf_q_437(.A(q_in_437), .Y(P2_IR[17]));
INVX2 g120206(.A (n_15791), .Y (n_15873));
CLKBUFX1 gbuf_d_438(.A(n_15642), .Y(d_out_438));
CLKBUFX1 gbuf_q_438(.A(q_in_438), .Y(P3_IR[13]));
CLKBUFX1 gbuf_d_439(.A(n_15650), .Y(d_out_439));
CLKBUFX1 gbuf_q_439(.A(q_in_439), .Y(P3_IR[17]));
INVX1 g120216(.A (n_34579), .Y (n_16067));
CLKBUFX1 gbuf_d_440(.A(n_15639), .Y(d_out_440));
CLKBUFX1 gbuf_q_440(.A(q_in_440), .Y(P3_IR[8]));
CLKBUFX1 gbuf_d_441(.A(n_15638), .Y(d_out_441));
CLKBUFX1 gbuf_q_441(.A(q_in_441), .Y(P1_IR[10]));
CLKBUFX1 gbuf_d_442(.A(n_15637), .Y(d_out_442));
CLKBUFX1 gbuf_q_442(.A(q_in_442), .Y(P1_IR[11]));
CLKBUFX1 gbuf_d_443(.A(n_15649), .Y(d_out_443));
CLKBUFX1 gbuf_q_443(.A(q_in_443), .Y(P1_IR[7]));
NAND2X1 g120228(.A (n_15629), .B (n_7904), .Y (n_15872));
INVX2 g120246(.A (n_15785), .Y (n_16036));
INVX1 g120256(.A (n_15784), .Y (n_15870));
NAND2X2 g120265(.A (n_15627), .B (n_8344), .Y (n_15868));
INVX2 g120273(.A (n_15783), .Y (n_35270));
AOI21X1 g120309(.A0 (n_15236), .A1 (datao_2[27] ), .B0 (n_15613), .Y(n_15860));
OAI21X1 g120318(.A0 (n_15676), .A1 (n_45), .B0 (n_15614), .Y(n_15858));
AOI21X1 g120324(.A0 (n_4288), .A1 (n_7793), .B0 (n_15615), .Y(n_15779));
MX2X1 g120350(.A (n_6170), .B (n_15700), .S0 (n_15643), .Y (n_15778));
MX2X1 g120365(.A (n_33034), .B (n_15692), .S0 (n_15968), .Y(n_15776));
MX2X1 g120366(.A (n_4825), .B (n_15696), .S0 (n_30702), .Y (n_15775));
MX2X1 g120367(.A (n_4731), .B (n_15698), .S0 (n_15968), .Y (n_15773));
MX2X1 g120368(.A (n_4478), .B (n_34349), .S0 (n_31105), .Y (n_15772));
MX2X1 g120369(.A (n_8105), .B (n_15687), .S0 (n_15968), .Y (n_15771));
MX2X1 g120370(.A (n_6204), .B (n_15689), .S0 (n_15968), .Y (n_15769));
MX2X1 g120373(.A (n_6810), .B (n_15602), .S0 (n_15968), .Y (n_15768));
INVX1 g120452(.A (n_15705), .Y (n_15849));
NOR2X1 g120460(.A (n_15766), .B (n_8293), .Y (n_15767));
INVX2 g120487(.A (n_15701), .Y (n_16137));
NOR2X1 g120533(.A (n_15665), .B (n_8746), .Y (n_15840));
NAND2X1 g120546(.A (n_15670), .B (n_16230), .Y (n_15838));
NOR2X1 g120560(.A (n_15667), .B (n_15763), .Y (n_16009));
NAND2X1 g120568(.A (n_15765), .B (n_16230), .Y (n_15835));
NAND2X1 g120578(.A (n_15764), .B (n_16230), .Y (n_16007));
NOR2X1 g120603(.A (n_15603), .B (n_15763), .Y (n_15832));
AOI22X1 g120881(.A0 (n_15608), .A1 (n_4944), .B0 (n_15676), .B1(datao_1[30] ), .Y (n_15967));
MX2X1 g120883(.A (datao_1[29] ), .B (n_5928), .S0 (n_15427), .Y(n_15829));
INVX1 g120894(.A (n_15761), .Y (n_15762));
AOI22X1 g120926(.A0 (n_15427), .A1 (n_5112), .B0 (n_15676), .B1(datao_1[31] ), .Y (n_15951));
MX2X1 g120958(.A (si[31]), .B (n_4865), .S0 (n_15676), .Y (n_15827));
MX2X1 g120961(.A (si[28]), .B (n_5684), .S0 (n_15676), .Y (n_15960));
MX2X1 g120996(.A (n_5790), .B (datao_2[29] ), .S0 (n_15427), .Y(n_15947));
NAND2X1 g120168(.A (n_15631), .B (n_8365), .Y (n_16061));
CLKBUFX1 gbuf_d_444(.A(n_15640), .Y(d_out_444));
CLKBUFX1 gbuf_q_444(.A(q_in_444), .Y(P3_IR[18]));
CLKBUFX1 gbuf_d_445(.A(n_15645), .Y(d_out_445));
CLKBUFX1 gbuf_q_445(.A(q_in_445), .Y(P3_IR[12]));
CLKBUFX1 gbuf_d_446(.A(n_15646), .Y(d_out_446));
CLKBUFX1 gbuf_q_446(.A(q_in_446), .Y(P3_IR[11]));
CLKBUFX1 gbuf_d_447(.A(n_15632), .Y(d_out_447));
CLKBUFX1 gbuf_q_447(.A(q_in_447), .Y(P1_IR[5]));
CLKBUFX1 gbuf_d_448(.A(n_15641), .Y(d_out_448));
CLKBUFX1 gbuf_q_448(.A(q_in_448), .Y(P3_IR[14]));
CLKBUFX1 gbuf_d_449(.A(n_15647), .Y(d_out_449));
CLKBUFX1 gbuf_q_449(.A(q_in_449), .Y(P3_IR[10]));
CLKBUFX1 gbuf_d_450(.A(n_15658), .Y(d_out_450));
CLKBUFX1 gbuf_q_450(.A(q_in_450), .Y(P2_IR[15]));
INVX1 g120085(.A (n_15757), .Y (n_15825));
CLKBUFX1 gbuf_d_451(.A(n_15635), .Y(d_out_451));
CLKBUFX1 gbuf_q_451(.A(q_in_451), .Y(P1_IR[3]));
CLKBUFX1 gbuf_d_452(.A(n_15589), .Y(d_out_452));
CLKBUFX1 gbuf_q_452(.A(q_in_452), .Y(P2_IR[12]));
CLKBUFX3 g120099(.A (n_15805), .Y (n_16273));
CLKBUFX1 gbuf_d_453(.A(n_15591), .Y(d_out_453));
CLKBUFX1 gbuf_q_453(.A(q_in_453), .Y(P2_IR[10]));
CLKBUFX1 gbuf_d_454(.A(n_15584), .Y(d_out_454));
CLKBUFX1 gbuf_q_454(.A(q_in_454), .Y(P1_IR[0]));
INVX1 g120130(.A (n_15811), .Y (n_35705));
CLKBUFX1 gbuf_d_455(.A(n_15587), .Y(d_out_455));
CLKBUFX1 gbuf_q_455(.A(q_in_455), .Y(P2_IR[9]));
CLKBUFX1 g120129(.A (n_15811), .Y (n_17630));
INVX1 g120187(.A (n_15753), .Y (n_15821));
CLKBUFX3 g120120(.A (n_15752), .Y (n_15819));
NAND2X2 g118709(.A (n_15749), .B (n_15493), .Y (n_17018));
NAND2X2 g118964(.A (n_9278), .B (n_15661), .Y (n_16284));
NAND2X1 g118987(.A (n_33268), .B (n_15493), .Y (n_15808));
NAND2X1 g119083(.A (n_8784), .B (n_15746), .Y (n_15747));
NAND2X1 g119097(.A (n_9243), .B (n_15746), .Y (n_15804));
INVX1 g119232(.A (n_34471), .Y (n_15745));
INVX2 g119237(.A (n_34471), .Y (n_15937));
NAND2X1 g119249(.A (n_15339), .B (n_15586), .Y (n_15929));
AOI21X1 g119251(.A0 (n_15387), .A1 (n_15461), .B0 (n_15653), .Y(n_15928));
INVX2 g119259(.A (n_15743), .Y (n_15934));
AOI21X1 g119314(.A0 (n_15451), .A1 (n_15576), .B0 (n_15585), .Y(n_15802));
INVX1 g120110(.A (n_15806), .Y (n_15797));
INVX1 g119513(.A (n_34002), .Y (n_15798));
NAND3X1 g119593(.A (n_15445), .B (n_6538), .C (n_15444), .Y(n_15795));
INVX2 g119642(.A (n_15737), .Y (n_15931));
NAND2X2 g120052(.A (n_7437), .B (n_15520), .Y (n_15919));
INVX1 g120086(.A (n_15736), .Y (n_15757));
CLKBUFX1 gbuf_d_456(.A(n_15590), .Y(d_out_456));
CLKBUFX1 gbuf_q_456(.A(q_in_456), .Y(P2_IR[11]));
INVX2 g120238(.A (n_15733), .Y (n_15787));
NAND2X2 g120247(.A (n_15580), .B (n_7894), .Y (n_15785));
NAND2X2 g120257(.A (n_15579), .B (n_7879), .Y (n_15784));
NAND2X1 g120274(.A (n_15578), .B (n_7813), .Y (n_15783));
OAI22X1 g120275(.A0 (n_35180), .A1 (n_15477), .B0 (n_15513), .B1(n_15484), .Y (n_15732));
OAI22X1 g120285(.A0 (n_4724), .A1 (n_15477), .B0 (n_15630), .B1(n_15864), .Y (n_15731));
OAI22X1 g120286(.A0 (n_4086), .A1 (n_16150), .B0 (n_15511), .B1(n_15864), .Y (n_15729));
OAI22X1 g120288(.A0 (n_6313), .A1 (n_16150), .B0 (n_15509), .B1(n_15484), .Y (n_15728));
AOI21X1 g120320(.A0 (n_15717), .A1 (n_15725), .B0 (n_7598), .Y(n_15727));
AOI21X1 g120325(.A0 (n_15720), .A1 (n_15725), .B0 (n_7635), .Y(n_15726));
OAI22X1 g120331(.A0 (n_15433), .A1 (n_15723), .B0 (n_3170), .B1(n_15722), .Y (n_15724));
MX2X1 g120333(.A (n_32386), .B (n_15720), .S0 (n_15975), .Y(n_15721));
MX2X1 g120343(.A (n_4735), .B (n_15717), .S0 (n_15975), .Y (n_15718));
MX2X1 g120345(.A (n_4844), .B (n_15616), .S0 (n_15975), .Y (n_15715));
MX2X1 g120364(.A (n_3845), .B (n_15625), .S0 (n_15968), .Y (n_15714));
OAI22X1 g120379(.A0 (n_15431), .A1 (n_15723), .B0 (n_2878), .B1(n_15722), .Y (n_15712));
OAI22X1 g120381(.A0 (n_15432), .A1 (n_15723), .B0 (n_2962), .B1(n_15722), .Y (n_15711));
NAND2X1 g120423(.A (n_15514), .B (n_15704), .Y (n_15710));
NAND2X1 g120424(.A (n_15512), .B (n_15708), .Y (n_15709));
INVX1 g120426(.A (n_15706), .Y (n_15707));
NAND2X1 g120453(.A (n_15510), .B (n_15704), .Y (n_15705));
OAI21X1 g120478(.A0 (n_5270), .A1 (n_15240), .B0 (n_15517), .Y(n_15703));
OAI21X1 g120479(.A0 (n_5263), .A1 (n_15676), .B0 (n_15516), .Y(n_15702));
NAND2X1 g120488(.A (n_15700), .B (n_8039), .Y (n_15701));
NAND2X1 g120640(.A (n_15698), .B (n_34355), .Y (n_15699));
NAND2X1 g120643(.A (n_15692), .B (n_34296), .Y (n_15693));
NAND2X1 g120644(.A (n_15692), .B (n_15622), .Y (n_15691));
NAND2X1 g120653(.A (n_15689), .B (n_34355), .Y (n_15690));
NAND2X1 g120655(.A (n_15687), .B (n_34355), .Y (n_15688));
NAND2X1 g120656(.A (n_15698), .B (n_15685), .Y (n_15686));
NAND2X1 g120659(.A (n_15687), .B (n_15685), .Y (n_15681));
NAND2X1 g120660(.A (n_15689), .B (n_15685), .Y (n_15680));
NOR2X1 g120685(.A (n_15508), .B (n_7821), .Y (n_15679));
OAI21X1 g120707(.A0 (n_5192), .A1 (n_15676), .B0 (n_15518), .Y(n_15678));
NAND4X1 g120880(.A (n_4069), .B (n_15198), .C (n_4634), .D (n_4635),.Y (n_15677));
AOI22X1 g120884(.A0 (n_15608), .A1 (n_5831), .B0 (n_15676), .B1(datao_1[28] ), .Y (n_15853));
INVX1 g120885(.A (n_15674), .Y (n_15675));
MX2X1 g120895(.A (n_12188), .B (n_4310), .S0 (n_15427), .Y (n_15761));
INVX1 g120896(.A (n_15672), .Y (n_15673));
INVX1 g120927(.A (n_15670), .Y (n_15671));
MX2X1 g120929(.A (n_4993), .B (n_479), .S0 (n_15608), .Y (n_15837));
INVX1 g120931(.A (n_15667), .Y (n_15668));
MX2X1 g120959(.A (n_5269), .B (si[30]), .S0 (n_15608), .Y (n_15845));
MX2X1 g120960(.A (n_5893), .B (si[29]), .S0 (n_15608), .Y (n_15844));
NAND2X1 g120962(.A (n_15498), .B (n_15505), .Y (n_15843));
NAND2X1 g120979(.A (n_15499), .B (n_15422), .Y (n_15842));
NAND2X1 g120987(.A (n_15500), .B (n_15426), .Y (n_15839));
INVX1 g120988(.A (n_15665), .Y (n_15666));
NAND2X1 g120990(.A (n_15497), .B (n_15421), .Y (n_15833));
MX2X1 g120997(.A (n_491), .B (n_5492), .S0 (n_15198), .Y (n_15831));
NAND2X2 g120208(.A (n_15583), .B (n_7849), .Y (n_15791));
CLKBUFX1 gbuf_d_457(.A(n_15588), .Y(d_out_457));
CLKBUFX1 gbuf_q_457(.A(q_in_457), .Y(P2_IR[8]));
INVX1 g120194(.A (n_15809), .Y (n_16552));
INVX1 g120139(.A (n_15663), .Y (n_15824));
INVX2 g120131(.A (n_15593), .Y (n_15811));
CLKBUFX1 gbuf_d_458(.A(n_15476), .Y(d_out_458));
CLKBUFX1 gbuf_q_458(.A(q_in_458), .Y(P2_IR[3]));
CLKBUFX1 gbuf_d_459(.A(n_15485), .Y(d_out_459));
CLKBUFX1 gbuf_q_459(.A(q_in_459), .Y(P2_IR[1]));
NAND2X1 g120188(.A (n_15449), .B (n_7884), .Y (n_15753));
INVX2 g120121(.A (n_15661), .Y (n_15752));
INVX2 g120112(.A (n_15592), .Y (n_15806));
NAND2X1 g119261(.A (n_15380), .B (n_15473), .Y (n_15743));
NAND2X2 g119634(.A (n_15384), .B (n_15471), .Y (n_15739));
NAND2X1 g119643(.A (n_32042), .B (n_32043), .Y (n_15737));
NAND2X2 g120079(.A (n_15448), .B (n_8147), .Y (n_32432));
CLKBUFX1 gbuf_d_460(.A(n_15450), .Y(d_out_460));
CLKBUFX1 gbuf_q_460(.A(q_in_460), .Y(P2_IR[0]));
INVX2 g120101(.A (n_34978), .Y (n_15805));
AOI21X1 g120239(.A0 (n_15656), .A1 (n_15399), .B0 (n_7428), .Y(n_15733));
OAI22X1 g120276(.A0 (n_4340), .A1 (n_16150), .B0 (n_15440), .B1(n_15864), .Y (n_15659));
OAI22X1 g120278(.A0 (n_34078), .A1 (n_16150), .B0 (n_15436), .B1(n_15864), .Y (n_15658));
MX2X1 g120284(.A (n_6988), .B (n_15656), .S0 (n_15480), .Y (n_15657));
CLKBUFX1 gbuf_d_461(.A(n_15465), .Y(d_out_461));
CLKBUFX1 gbuf_q_461(.A(q_in_461), .Y(P3_IR[7]));
OAI22X1 g120300(.A0 (n_4210), .A1 (n_16415), .B0 (n_15434), .B1(n_15864), .Y (n_15655));
INVX1 g120305(.A (n_15653), .Y (n_15654));
AOI21X1 g120319(.A0 (n_15644), .A1 (n_15725), .B0 (n_7636), .Y(n_15652));
MX2X1 g120328(.A (n_3854), .B (n_15535), .S0 (n_15975), .Y (n_15651));
MX2X1 g120334(.A (n_4288), .B (n_15540), .S0 (n_15975), .Y (n_15650));
CLKBUFX1 gbuf_d_462(.A(n_15456), .Y(d_out_462));
CLKBUFX1 gbuf_q_462(.A(q_in_462), .Y(P3_IR[4]));
MX2X1 g120335(.A (n_35368), .B (n_15568), .S0 (n_15968), .Y(n_15649));
MX2X1 g120338(.A (n_3862), .B (n_15532), .S0 (n_15643), .Y (n_15647));
MX2X1 g120339(.A (n_4040), .B (n_15538), .S0 (n_15975), .Y (n_15646));
MX2X1 g120340(.A (n_10656), .B (n_15644), .S0 (n_15643), .Y(n_15645));
MX2X1 g120341(.A (n_32445), .B (n_15527), .S0 (n_13010), .Y(n_15642));
MX2X1 g120342(.A (n_4320), .B (n_15523), .S0 (n_15643), .Y (n_15641));
MX2X1 g120344(.A (n_33901), .B (n_15542), .S0 (n_15643), .Y(n_15640));
CLKBUFX1 gbuf_d_463(.A(n_15458), .Y(d_out_463));
CLKBUFX1 gbuf_q_463(.A(q_in_463), .Y(P3_IR[3]));
CLKBUFX1 gbuf_d_464(.A(n_15467), .Y(d_out_464));
CLKBUFX1 gbuf_q_464(.A(q_in_464), .Y(P3_IR[5]));
MX2X1 g120359(.A (n_4133), .B (n_15519), .S0 (n_15975), .Y (n_15639));
MX2X1 g120361(.A (n_3959), .B (n_15551), .S0 (n_15968), .Y (n_15638));
MX2X1 g120362(.A (n_4535), .B (n_15547), .S0 (n_15968), .Y (n_15637));
MX2X1 g120363(.A (n_4010), .B (n_15560), .S0 (n_15968), .Y (n_15636));
MX2X1 g120380(.A (n_3472), .B (n_15562), .S0 (n_30702), .Y (n_15635));
MX2X1 g120382(.A (n_8115), .B (n_15556), .S0 (n_15968), .Y (n_15634));
MX2X1 g120386(.A (n_3870), .B (n_34291), .S0 (n_31105), .Y (n_15633));
OAI22X1 g120387(.A0 (n_15366), .A1 (n_15723), .B0 (n_3483), .B1(n_15722), .Y (n_15632));
NAND2X1 g120425(.A (n_15441), .B (n_15628), .Y (n_15631));
NOR2X1 g120427(.A (n_15630), .B (n_7581), .Y (n_15706));
NAND2X1 g120470(.A (n_15437), .B (n_15628), .Y (n_15629));
NAND2X1 g120473(.A (n_15435), .B (n_15628), .Y (n_15627));
NAND2X1 g120638(.A (n_15625), .B (n_34296), .Y (n_15626));
NAND2X1 g120639(.A (n_15625), .B (n_15622), .Y (n_15623));
NAND2X1 g120665(.A (n_15619), .B (n_15720), .Y (n_15621));
NAND2X1 g120675(.A (n_15619), .B (n_15717), .Y (n_15620));
NAND2X1 g120684(.A (n_7641), .B (n_15616), .Y (n_33012));
NOR2X1 g120686(.A (n_15429), .B (n_7403), .Y (n_15615));
AOI22X1 g120705(.A0 (n_5435), .A1 (n_15198), .B0 (n_15360), .B1(n_4779), .Y (n_15614));
OAI21X1 g120717(.A0 (n_5583), .A1 (n_15608), .B0 (n_15442), .Y(n_15613));
INVX1 g120195(.A (n_15746), .Y (n_15809));
CLKBUFX1 gbuf_d_465(.A(n_15462), .Y(d_out_465));
CLKBUFX1 gbuf_q_465(.A(q_in_465), .Y(P3_IR[1]));
NAND4X1 g120876(.A (n_5182), .B (n_15676), .C (n_4321), .D (n_4322),.Y (n_15612));
NAND4X1 g120877(.A (n_5188), .B (n_15676), .C (n_5189), .D (n_5190),.Y (n_15610));
NAND4X1 g120878(.A (n_4637), .B (n_15676), .C (n_4638), .D (n_4639),.Y (n_15609));
AOI22X1 g120886(.A0 (n_15608), .A1 (n_5294), .B0 (n_15198), .B1(datao_1[24] ), .Y (n_15674));
AOI22X1 g120897(.A0 (n_15608), .A1 (n_4444), .B0 (n_15676), .B1(datao_1[23] ), .Y (n_15672));
AOI22X1 g120900(.A0 (n_15236), .A1 (n_5029), .B0 (n_15676), .B1(n_12026), .Y (n_15766));
MX2X1 g120928(.A (datao_2[31] ), .B (n_4782), .S0 (n_15676), .Y(n_15670));
MX2X1 g120930(.A (n_667), .B (n_5008), .S0 (n_15676), .Y (n_15765));
AOI21X1 g120932(.A0 (n_15676), .A1 (n_4296), .B0 (n_15424), .Y(n_15667));
MX2X1 g120956(.A (datao_2[22] ), .B (n_4181), .S0 (n_15676), .Y(n_15764));
AOI21X1 g120989(.A0 (n_15240), .A1 (n_5117), .B0 (n_15428), .Y(n_15665));
INVX1 g120992(.A (n_15602), .Y (n_15603));
NAND2X1 g121009(.A (n_15427), .B (datao_2[26] ), .Y (n_15601));
NAND2X1 g121023(.A (n_15427), .B (si[27]), .Y (n_15599));
NAND2X1 g121024(.A (n_15608), .B (si[26]), .Y (n_15598));
OR2X1 g121055(.A (n_4842), .B (n_15427), .Y (n_15596));
CLKBUFX1 gbuf_d_466(.A(n_15454), .Y(d_out_466));
CLKBUFX1 gbuf_q_466(.A(q_in_466), .Y(P3_IR[6]));
CLKBUFX1 gbuf_d_467(.A(n_15452), .Y(d_out_467));
CLKBUFX1 gbuf_q_467(.A(q_in_467), .Y(P1_IR[1]));
CLKBUFX1 gbuf_d_468(.A(n_15460), .Y(d_out_468));
CLKBUFX1 gbuf_q_468(.A(q_in_468), .Y(P3_IR[2]));
CLKBUFX1 gbuf_d_469(.A(n_15486), .Y(d_out_469));
CLKBUFX1 gbuf_q_469(.A(q_in_469), .Y(P2_IR[2]));
CLKBUFX1 gbuf_d_470(.A(n_15482), .Y(d_out_470));
CLKBUFX1 gbuf_q_470(.A(q_in_470), .Y(P2_IR[5]));
CLKBUFX1 gbuf_d_471(.A(n_15479), .Y(d_out_471));
CLKBUFX1 gbuf_q_471(.A(q_in_471), .Y(P2_IR[7]));
CLKBUFX1 gbuf_d_472(.A(n_15478), .Y(d_out_472));
CLKBUFX1 gbuf_q_472(.A(q_in_472), .Y(P2_IR[4]));
CLKBUFX1 gbuf_d_473(.A(n_15481), .Y(d_out_473));
CLKBUFX1 gbuf_q_473(.A(q_in_473), .Y(P2_IR[6]));
INVX1 g120087(.A (n_15493), .Y (n_15736));
NAND2X1 g120140(.A (n_15447), .B (n_8741), .Y (n_15663));
NAND2X2 g120123(.A (n_15395), .B (n_8139), .Y (n_15661));
NAND2X1 g120132(.A (n_15393), .B (n_8135), .Y (n_15593));
NAND2X2 g120113(.A (n_15398), .B (n_8048), .Y (n_15592));
OAI22X1 g120281(.A0 (n_3917), .A1 (n_16150), .B0 (n_15371), .B1(n_15864), .Y (n_15591));
OAI22X1 g120282(.A0 (n_4395), .A1 (n_16150), .B0 (n_15369), .B1(n_15484), .Y (n_15590));
OAI22X1 g120283(.A0 (n_4389), .A1 (n_16150), .B0 (n_15367), .B1(n_15864), .Y (n_15589));
OAI22X1 g120296(.A0 (n_4055), .A1 (n_16150), .B0 (n_15374), .B1(n_15864), .Y (n_15588));
OAI22X1 g120297(.A0 (n_3883), .A1 (n_16150), .B0 (n_15376), .B1(n_15864), .Y (n_15587));
AOI21X1 g120304(.A0 (n_33895), .A1 (n_32505), .B0 (n_15382), .Y(n_15586));
NAND2X1 g120306(.A (n_15379), .B (n_7179), .Y (n_15653));
NAND2X1 g120310(.A (n_15389), .B (n_6722), .Y (n_15585));
MX2X1 g120360(.A (n_7747), .B (n_15446), .S0 (n_35017), .Y (n_15584));
NAND2X1 g120468(.A (n_15377), .B (n_15581), .Y (n_15583));
NAND2X1 g120471(.A (n_15372), .B (n_15581), .Y (n_15580));
NAND2X1 g120472(.A (n_15370), .B (n_15581), .Y (n_15579));
NAND2X1 g120474(.A (n_15368), .B (n_15581), .Y (n_15578));
NAND2X1 g120624(.A (n_15574), .B (n_15576), .Y (n_15577));
NAND2X1 g120625(.A (n_15574), .B (n_15570), .Y (n_15575));
NAND2X1 g120628(.A (n_15571), .B (n_15576), .Y (n_15573));
NAND2X1 g120629(.A (n_15571), .B (n_15570), .Y (n_15572));
NAND2X1 g120630(.A (n_15568), .B (n_34354), .Y (n_15569));
NAND2X1 g120631(.A (n_15568), .B (n_15558), .Y (n_15567));
NAND2X1 g120632(.A (n_15564), .B (n_15576), .Y (n_15566));
NAND2X1 g120633(.A (n_15564), .B (n_15570), .Y (n_15565));
NAND2X1 g120634(.A (n_15562), .B (n_15576), .Y (n_15563));
NAND2X1 g120636(.A (n_15560), .B (n_34354), .Y (n_15561));
NAND2X1 g120637(.A (n_15560), .B (n_15558), .Y (n_15559));
NAND2X1 g120645(.A (n_15556), .B (n_34296), .Y (n_15557));
NAND2X1 g120648(.A (n_15551), .B (n_34354), .Y (n_15552));
NAND2X1 g120649(.A (n_15551), .B (n_15558), .Y (n_15549));
NAND2X1 g120650(.A (n_15547), .B (n_34296), .Y (n_15548));
NAND2X1 g120651(.A (n_15547), .B (n_15558), .Y (n_15546));
NAND2X1 g120652(.A (n_15562), .B (n_15570), .Y (n_15545));
NAND2X1 g120654(.A (n_15556), .B (n_15558), .Y (n_15544));
NAND2X1 g120662(.A (n_15619), .B (n_15540), .Y (n_15541));
NAND2X1 g120664(.A (n_15536), .B (n_15538), .Y (n_15539));
NAND2X1 g120666(.A (n_15536), .B (n_15535), .Y (n_15537));
NAND2X1 g120667(.A (n_15535), .B (n_15530), .Y (n_15534));
NAND2X1 g120668(.A (n_15536), .B (n_15532), .Y (n_15533));
NAND2X1 g120669(.A (n_15532), .B (n_15530), .Y (n_15531));
NAND2X1 g120670(.A (n_15619), .B (n_15644), .Y (n_15529));
NAND2X1 g120671(.A (n_15536), .B (n_15527), .Y (n_15528));
NAND2X1 g120672(.A (n_15527), .B (n_15725), .Y (n_15526));
NAND2X1 g120673(.A (n_15536), .B (n_15523), .Y (n_15524));
NAND2X1 g120674(.A (n_15523), .B (n_15725), .Y (n_15522));
NAND2X1 g120688(.A (n_15538), .B (n_15530), .Y (n_15521));
OAI21X1 g120749(.A0 (n_7640), .A1 (n_7457), .B0 (n_15519), .Y(n_15520));
NAND4X1 g120777(.A (n_15427), .B (n_4442), .C (n_4937), .D (n_4938),.Y (n_15518));
NAND4X1 g120799(.A (n_4851), .B (n_15427), .C (n_4852), .D (n_4853),.Y (n_15517));
NAND4X1 g120800(.A (n_15427), .B (n_4417), .C (n_4855), .D (n_4856),.Y (n_15516));
INVX1 g120887(.A (n_15513), .Y (n_15514));
INVX1 g120889(.A (n_15511), .Y (n_15512));
INVX1 g120898(.A (n_15509), .Y (n_15510));
NAND2X1 g120940(.A (n_15365), .B (n_15329), .Y (n_15687));
NAND2X1 g120949(.A (n_15363), .B (n_15324), .Y (n_15696));
NAND2X1 g120950(.A (n_15362), .B (n_15322), .Y (n_15692));
OAI22X1 g120978(.A0 (n_15198), .A1 (n_28), .B0 (n_15608), .B1(n_4454), .Y (n_15700));
INVX1 g120982(.A (n_15616), .Y (n_15508));
MX2X1 g120993(.A (datao_2[21] ), .B (n_4633), .S0 (n_15198), .Y(n_15602));
NAND2X1 g120994(.A (n_15356), .B (n_15316), .Y (n_15698));
NAND2X1 g120998(.A (n_15357), .B (n_15315), .Y (n_15689));
NAND2X1 g121001(.A (n_15236), .B (datao_2[25] ), .Y (n_15506));
NAND2X1 g121025(.A (n_15236), .B (si[24]), .Y (n_15505));
OAI21X1 g121056(.A0 (n_5115), .A1 (n_5191), .B0 (n_15676), .Y(n_15504));
OAI21X1 g121057(.A0 (n_4456), .A1 (n_4640), .B0 (n_15676), .Y(n_15502));
NAND2X1 g121073(.A (n_5183), .B (n_15676), .Y (n_15501));
NAND2X1 g121077(.A (n_15676), .B (n_5007), .Y (n_15500));
NAND2X1 g121093(.A (n_15676), .B (n_4503), .Y (n_15499));
NAND2X1 g121101(.A (n_15676), .B (n_5164), .Y (n_15498));
NAND2X1 g121142(.A (n_15676), .B (n_4666), .Y (n_15497));
CLKBUFX1 gbuf_d_474(.A(n_15403), .Y(d_out_474));
CLKBUFX1 gbuf_q_474(.A(q_in_474), .Y(P3_IR[0]));
NAND2X1 g120196(.A (n_15391), .B (n_8129), .Y (n_15746));
INVX2 g120080(.A (n_15492), .Y (n_15493));
NAND2X1 g118428(.A (n_15348), .B (n_33629), .Y (n_15491));
AOI21X1 g120038(.A0 (n_15262), .A1 (n_29133), .B0 (n_8614), .Y(n_15490));
AOI21X1 g120044(.A0 (n_15259), .A1 (n_26570), .B0 (n_8614), .Y(n_15487));
MX2X1 g120277(.A (n_6887), .B (n_15392), .S0 (n_15477), .Y (n_15486));
OAI22X1 g120287(.A0 (n_15239), .A1 (n_15484), .B0 (n_2824), .B1(n_31328), .Y (n_15485));
MX2X1 g120293(.A (n_6962), .B (n_15397), .S0 (n_15480), .Y (n_15482));
MX2X1 g120294(.A (n_6964), .B (n_15400), .S0 (n_15480), .Y (n_15481));
OAI22X1 g120295(.A0 (n_3863), .A1 (n_16150), .B0 (n_15334), .B1(n_15864), .Y (n_15479));
MX2X1 g120298(.A (n_6963), .B (n_15394), .S0 (n_15477), .Y (n_15478));
OAI22X1 g120299(.A0 (n_15332), .A1 (n_15484), .B0 (n_3665), .B1(n_31328), .Y (n_15476));
AOI21X1 g120303(.A0 (n_15470), .A1 (n_15466), .B0 (n_7341), .Y(n_15474));
AOI21X1 g120307(.A0 (n_15457), .A1 (n_34469), .B0 (n_7299), .Y(n_15473));
AOI21X1 g120326(.A0 (n_15453), .A1 (n_15470), .B0 (n_7339), .Y(n_15471));
AOI21X1 g120327(.A0 (n_15459), .A1 (n_34469), .B0 (n_7286), .Y(n_32042));
MX2X1 g120329(.A (n_10740), .B (n_15466), .S0 (n_7417), .Y (n_15467));
MX2X1 g120332(.A (n_3583), .B (n_15464), .S0 (n_7417), .Y (n_15465));
MX2X1 g120346(.A (n_3063), .B (n_15461), .S0 (n_15975), .Y (n_15462));
MX2X1 g120353(.A (n_2872), .B (n_15459), .S0 (n_15975), .Y (n_15460));
MX2X1 g120356(.A (n_3165), .B (n_15457), .S0 (n_15975), .Y (n_15458));
MX2X1 g120357(.A (n_3176), .B (n_34466), .S0 (n_15643), .Y (n_15456));
MX2X1 g120358(.A (n_3429), .B (n_15453), .S0 (n_15643), .Y (n_15454));
MX2X1 g120371(.A (n_2807), .B (n_15451), .S0 (n_15968), .Y (n_15452));
MX2X1 g120383(.A (n_1803), .B (n_15390), .S0 (n_15477), .Y (n_15450));
NAND2X1 g120461(.A (n_15335), .B (n_15396), .Y (n_15449));
NAND2X1 g120465(.A (n_15333), .B (n_7297), .Y (n_15448));
NAND2X1 g120569(.A (n_15446), .B (n_7139), .Y (n_15447));
NAND2X1 g120626(.A (n_15443), .B (n_15576), .Y (n_15445));
NAND2X1 g120627(.A (n_15443), .B (n_15570), .Y (n_15444));
NAND4X1 g120879(.A (n_4781), .B (n_15676), .C (n_5194), .D (n_5195),.Y (n_15442));
AOI22X1 g120888(.A0 (n_15236), .A1 (n_4455), .B0 (n_15676), .B1(datao_1[19] ), .Y (n_15513));
AOI22X1 g120890(.A0 (n_15608), .A1 (n_4290), .B0 (n_15198), .B1(n_693), .Y (n_15511));
INVX1 g120891(.A (n_15440), .Y (n_15441));
AOI22X1 g120893(.A0 (n_15427), .A1 (n_4303), .B0 (n_15198), .B1(n_12454), .Y (n_15630));
AOI22X1 g120899(.A0 (n_15427), .A1 (n_5116), .B0 (n_15198), .B1(n_12322), .Y (n_15509));
INVX1 g120915(.A (n_15436), .Y (n_15437));
INVX1 g120922(.A (n_15434), .Y (n_15435));
INVX1 g120933(.A (n_15574), .Y (n_15433));
INVX1 g120937(.A (n_15571), .Y (n_15432));
INVX1 g120941(.A (n_15564), .Y (n_15431));
NAND2X1 g120947(.A (n_15314), .B (n_15325), .Y (n_15625));
NAND2X1 g120969(.A (n_15201), .B (n_15320), .Y (n_15717));
INVX1 g120980(.A (n_15542), .Y (n_15430));
NAND2X1 g120983(.A (n_15222), .B (n_15318), .Y (n_15616));
INVX1 g120984(.A (n_15540), .Y (n_15429));
NAND2X1 g120986(.A (n_15313), .B (n_15317), .Y (n_15720));
AND2X1 g121011(.A (n_15427), .B (si[20]), .Y (n_15428));
NAND2X1 g121021(.A (n_15608), .B (si[21]), .Y (n_15426));
AND2X1 g121022(.A (n_15608), .B (datao_2[23] ), .Y (n_15424));
NAND2X1 g121037(.A (n_15608), .B (si[22]), .Y (n_15422));
NAND2X1 g121042(.A (n_15608), .B (datao_2[20] ), .Y (n_15421));
AND2X1 g121485(.A (n_15305), .B (n_34423), .Y (n_15419));
NAND2X2 g120090(.A (n_15340), .B (n_8143), .Y (n_15492));
NAND2X1 g118425(.A (n_15303), .B (n_33661), .Y (n_35704));
AOI21X1 g118426(.A0 (n_15117), .A1 (n_15415), .B0 (n_14641), .Y(n_15416));
NAND2X1 g118427(.A (n_15301), .B (n_15413), .Y (n_15414));
AOI21X1 g118430(.A0 (n_15114), .A1 (n_15409), .B0 (n_33713), .Y(n_15410));
AOI21X1 g118439(.A0 (n_15113), .A1 (n_15407), .B0 (n_33713), .Y(n_15408));
NAND4X1 g119423(.A (n_14844), .B (n_14638), .C (n_15405), .D(n_14764), .Y (n_15406));
NAND2X1 g120056(.A (n_15272), .B (n_15288), .Y (n_15404));
MX2X1 g120337(.A (n_32509), .B (n_15338), .S0 (n_349), .Y (n_15403));
NAND2X1 g120463(.A (n_15397), .B (n_15396), .Y (n_15398));
NAND2X1 g120464(.A (n_15394), .B (n_15396), .Y (n_15395));
NAND2X1 g120466(.A (n_15392), .B (n_15396), .Y (n_15393));
NAND2X1 g120594(.A (n_15390), .B (n_15396), .Y (n_15391));
NAND2X1 g120635(.A (n_15451), .B (n_6464), .Y (n_15389));
NAND2X1 g120663(.A (n_15387), .B (n_15459), .Y (n_32043));
NAND2X1 g120677(.A (n_7291), .B (n_15466), .Y (n_15385));
NAND2X1 g120678(.A (n_7291), .B (n_15453), .Y (n_15384));
NOR2X1 g120681(.A (n_15237), .B (n_34472), .Y (n_15382));
NAND2X1 g120682(.A (n_15387), .B (n_15461), .Y (n_15381));
NAND2X1 g120687(.A (n_15387), .B (n_15457), .Y (n_15380));
NAND2X1 g120689(.A (n_15461), .B (n_34469), .Y (n_15379));
NAND2X1 g120697(.A (n_15244), .B (n_8313), .Y (n_15378));
AOI22X1 g120892(.A0 (n_15608), .A1 (n_4956), .B0 (n_15240), .B1(n_475), .Y (n_15440));
INVX1 g120911(.A (n_15376), .Y (n_15377));
INVX1 g120913(.A (n_15374), .Y (n_15375));
AOI22X1 g120916(.A0 (n_15608), .A1 (n_3880), .B0 (n_15240), .B1(n_12028), .Y (n_15436));
OAI22X1 g120917(.A0 (n_15240), .A1 (n_3981), .B0 (n_15608), .B1(n_540), .Y (n_15656));
INVX1 g120918(.A (n_15371), .Y (n_15372));
INVX1 g120920(.A (n_15369), .Y (n_15370));
AOI22X1 g120923(.A0 (n_15608), .A1 (n_4291), .B0 (n_15240), .B1(n_12030), .Y (n_15434));
INVX1 g120924(.A (n_15367), .Y (n_15368));
NAND2X1 g120934(.A (n_15224), .B (n_15054), .Y (n_15574));
INVX1 g120935(.A (n_15443), .Y (n_15366));
NAND2X1 g120938(.A (n_15220), .B (n_15053), .Y (n_15571));
NAND2X1 g120939(.A (n_15218), .B (n_15052), .Y (n_15568));
NAND2X1 g120942(.A (n_15216), .B (n_15051), .Y (n_15564));
NAND2X1 g120943(.A (n_15213), .B (n_15049), .Y (n_15562));
NAND2X1 g120946(.A (n_15211), .B (n_15047), .Y (n_15560));
NAND2X1 g120951(.A (n_15210), .B (n_15234), .Y (n_15556));
NAND2X1 g120953(.A (n_15195), .B (n_15046), .Y (n_15551));
NAND2X1 g120954(.A (n_15208), .B (n_15231), .Y (n_15547));
NAND2X1 g120955(.A (n_15202), .B (n_15235), .Y (n_15523));
NAND2X1 g120963(.A (n_15206), .B (n_15230), .Y (n_15519));
NAND2X1 g120964(.A (n_15205), .B (n_15045), .Y (n_15535));
NAND2X1 g120965(.A (n_15212), .B (n_15043), .Y (n_15532));
NAND2X1 g120966(.A (n_15203), .B (n_15044), .Y (n_15538));
NAND2X1 g120967(.A (n_15214), .B (n_15229), .Y (n_15644));
NAND2X1 g120968(.A (n_15196), .B (n_15228), .Y (n_15527));
NAND2X1 g120981(.A (n_15199), .B (n_15227), .Y (n_15542));
NAND2X1 g120985(.A (n_15197), .B (n_15226), .Y (n_15540));
NAND2X1 g121085(.A (n_15676), .B (n_4033), .Y (n_15365));
NAND2X1 g121094(.A (n_15676), .B (n_3814), .Y (n_15363));
NAND2X1 g121095(.A (n_15198), .B (n_3617), .Y (n_15362));
NOR2X1 g121102(.A (n_5113), .B (n_15236), .Y (n_15360));
NAND2X1 g121103(.A (n_15198), .B (n_4538), .Y (n_15358));
NAND2X1 g121122(.A (n_15198), .B (n_4453), .Y (n_15357));
NAND2X1 g121126(.A (n_15676), .B (n_3976), .Y (n_15356));
OAI21X1 g121526(.A0 (n_14987), .A1 (n_15352), .B0 (n_14490), .Y(n_15353));
NAND2X1 g118413(.A (n_15128), .B (n_8313), .Y (n_15350));
NAND2X1 g119146(.A (n_15116), .B (n_15347), .Y (n_15348));
NAND2X1 g119645(.A (n_15118), .B (n_13662), .Y (n_15346));
AOI21X1 g120036(.A0 (n_14961), .A1 (n_33792), .B0 (n_14916), .Y(n_15345));
NAND2X1 g120039(.A (n_15095), .B (n_8313), .Y (n_15344));
AOI21X1 g120041(.A0 (n_14960), .A1 (n_29667), .B0 (n_9971), .Y(n_15342));
AOI21X1 g120043(.A0 (n_14958), .A1 (n_26558), .B0 (n_8614), .Y(n_15341));
NAND2X1 g120467(.A (n_15238), .B (n_15396), .Y (n_15340));
NAND2X1 g120680(.A (n_15387), .B (n_15338), .Y (n_15339));
NAND2X1 g120691(.A (n_15057), .B (n_8313), .Y (n_15337));
NAND2X1 g120715(.A (n_15088), .B (n_15110), .Y (n_15336));
INVX1 g120901(.A (n_15334), .Y (n_15335));
INVX1 g120906(.A (n_15332), .Y (n_15333));
AOI22X1 g120912(.A0 (n_15236), .A1 (n_4197), .B0 (n_15676), .B1(datao_1[9] ), .Y (n_15376));
AOI22X1 g120914(.A0 (n_15236), .A1 (n_3426), .B0 (n_15198), .B1(n_12184), .Y (n_15374));
AOI22X1 g120919(.A0 (n_15236), .A1 (n_3821), .B0 (n_15198), .B1(datao_1[10] ), .Y (n_15371));
AOI22X1 g120921(.A0 (n_15236), .A1 (n_3791), .B0 (n_15240), .B1(datao_1[11] ), .Y (n_15369));
AOI22X1 g120925(.A0 (n_15236), .A1 (n_4122), .B0 (n_15240), .B1(n_11802), .Y (n_15367));
NAND2X1 g120936(.A (n_15041), .B (n_14915), .Y (n_15443));
OAI22X1 g120944(.A0 (n_15198), .A1 (n_144), .B0 (n_15236), .B1(n_1131), .Y (n_15446));
NAND2X1 g121000(.A (n_15608), .B (datao_2[18] ), .Y (n_15329));
NAND2X1 g121007(.A (n_15608), .B (datao_2[17] ), .Y (n_15327));
NAND2X1 g121010(.A (n_15236), .B (datao_2[13] ), .Y (n_15325));
NAND2X1 g121014(.A (n_15608), .B (datao_2[15] ), .Y (n_15324));
NAND2X1 g121015(.A (n_15608), .B (datao_2[14] ), .Y (n_15322));
NAND2X1 g121030(.A (n_15236), .B (si[15]), .Y (n_15320));
NAND2X1 g121039(.A (n_15236), .B (si[19]), .Y (n_15318));
NAND2X1 g121041(.A (n_15236), .B (si[16]), .Y (n_15317));
NAND2X1 g121045(.A (n_15608), .B (datao_2[16] ), .Y (n_15316));
NAND2X1 g121047(.A (n_15608), .B (datao_2[19] ), .Y (n_15315));
NAND2X1 g121092(.A (n_15198), .B (n_4036), .Y (n_15314));
NAND2X1 g121118(.A (n_15198), .B (n_4191), .Y (n_15313));
AOI21X1 g121285(.A0 (n_8284), .A1 (n_13967), .B0 (n_14999), .Y(n_15311));
NAND2X1 g121520(.A (n_14994), .B (n_24028), .Y (n_32871));
AOI21X1 g121528(.A0 (n_10925), .A1 (n_19494), .B0 (n_14991), .Y(n_15306));
AOI22X1 g121846(.A0 (n_14534), .A1 (n_14496), .B0 (n_18289), .B1(n_14096), .Y (n_15305));
AOI21X1 g118414(.A0 (n_14752), .A1 (n_25151), .B0 (n_8614), .Y(n_15304));
OAI21X1 g119113(.A0 (n_15300), .A1 (n_35572), .B0 (n_15302), .Y(n_15303));
OAI21X1 g119144(.A0 (n_15300), .A1 (n_35829), .B0 (n_15299), .Y(n_15301));
OAI21X1 g119165(.A0 (n_15300), .A1 (n_14749), .B0 (n_15297), .Y(n_15298));
OAI21X1 g119424(.A0 (n_15300), .A1 (n_13163), .B0 (n_15295), .Y(n_15296));
AOI21X1 g119618(.A0 (n_15292), .A1 (n_23001), .B0 (n_14053), .Y(n_15294));
AOI21X1 g119646(.A0 (n_15292), .A1 (n_18384), .B0 (n_14304), .Y(n_15293));
AOI21X1 g119647(.A0 (n_15292), .A1 (n_32764), .B0 (n_14292), .Y(n_15291));
NAND2X1 g120042(.A (n_14970), .B (n_8313), .Y (n_15290));
NAND2X1 g120046(.A (n_14962), .B (n_15288), .Y (n_15289));
NAND2X1 g120054(.A (n_14977), .B (n_15110), .Y (n_15287));
NAND2X1 g120055(.A (n_14975), .B (n_15110), .Y (n_15285));
NAND2X1 g120061(.A (n_14964), .B (n_8313), .Y (n_15284));
AOI21X1 g120068(.A0 (n_15280), .A1 (n_23192), .B0 (n_13461), .Y(n_15282));
AOI21X1 g120093(.A0 (n_15280), .A1 (n_13274), .B0 (n_13863), .Y(n_15281));
AOI21X1 g120690(.A0 (n_14691), .A1 (n_26208), .B0 (n_8614), .Y(n_15279));
NAND2X1 g120694(.A (n_14932), .B (n_22821), .Y (n_15278));
AOI21X1 g120699(.A0 (n_14688), .A1 (n_26199), .B0 (n_8614), .Y(n_15277));
NAND2X1 g120708(.A (n_14951), .B (n_33629), .Y (n_15275));
NAND2X1 g120709(.A (n_14949), .B (n_15413), .Y (n_15273));
NAND2X1 g120710(.A (n_14957), .B (n_29666), .Y (n_15272));
NAND2X1 g120711(.A (n_14947), .B (n_15110), .Y (n_15271));
NAND2X1 g120712(.A (n_14945), .B (n_33661), .Y (n_15269));
NAND2X1 g120713(.A (n_14943), .B (n_15252), .Y (n_15267));
NAND2X1 g120719(.A (n_14940), .B (n_15413), .Y (n_15266));
NAND2X1 g120727(.A (n_14922), .B (n_22821), .Y (n_15264));
NAND2X1 g120740(.A (n_14931), .B (n_15110), .Y (n_15263));
NAND2X1 g120756(.A (n_15260), .B (n_17719), .Y (n_15262));
NAND2X1 g120758(.A (n_15260), .B (n_18384), .Y (n_15261));
NAND2X1 g120761(.A (n_15260), .B (n_32697), .Y (n_15259));
INVX1 g120772(.A (n_15257), .Y (n_15258));
OAI21X1 g120807(.A0 (n_14217), .A1 (n_23178), .B0 (n_25675), .Y(n_15256));
NAND2X1 g120811(.A (n_14873), .B (n_8313), .Y (n_15255));
OAI21X1 g120812(.A0 (n_14217), .A1 (n_17304), .B0 (n_25702), .Y(n_15254));
NAND2X1 g120826(.A (n_14903), .B (n_15252), .Y (n_15253));
NAND2X1 g120833(.A (n_14907), .B (n_33629), .Y (n_15251));
NAND2X1 g120835(.A (n_14891), .B (n_15110), .Y (n_15250));
NAND2X1 g120836(.A (n_14888), .B (n_15110), .Y (n_15249));
NAND2X1 g120838(.A (n_14886), .B (n_15413), .Y (n_15247));
NAND2X1 g120839(.A (n_14884), .B (n_15252), .Y (n_15245));
NAND2X1 g120857(.A (n_14908), .B (n_27384), .Y (n_15244));
AOI22X1 g120902(.A0 (n_15608), .A1 (n_3389), .B0 (n_15240), .B1(datao_1[7] ), .Y (n_15334));
OAI22X1 g120903(.A0 (n_15240), .A1 (n_3225), .B0 (n_15608), .B1(n_492), .Y (n_15400));
OAI22X1 g120904(.A0 (n_15240), .A1 (n_3788), .B0 (n_15427), .B1(n_602), .Y (n_15397));
OAI22X1 g120905(.A0 (n_15240), .A1 (n_2855), .B0 (n_15236), .B1(n_585), .Y (n_15394));
AOI22X1 g120907(.A0 (n_15427), .A1 (n_2813), .B0 (n_15240), .B1(n_12022), .Y (n_15332));
OAI22X1 g120908(.A0 (n_15676), .A1 (n_2543), .B0 (n_15236), .B1(n_294), .Y (n_15392));
INVX1 g120909(.A (n_15238), .Y (n_15239));
NAND2X1 g120945(.A (n_14904), .B (n_14913), .Y (n_15451));
NAND2X1 g120948(.A (n_14899), .B (n_14909), .Y (n_15453));
NAND2X1 g120971(.A (n_14900), .B (n_14910), .Y (n_15466));
NAND2X1 g120972(.A (n_14897), .B (n_14912), .Y (n_15464));
INVX1 g120973(.A (n_15338), .Y (n_15237));
NAND2X1 g120975(.A (n_14896), .B (n_14696), .Y (n_15461));
NAND2X1 g120976(.A (n_14895), .B (n_14693), .Y (n_15457));
NAND2X1 g120977(.A (n_14893), .B (n_14694), .Y (n_15459));
OAI22X1 g120991(.A0 (n_15240), .A1 (n_1686), .B0 (n_15236), .B1(n_275), .Y (n_15390));
NAND2X1 g120999(.A (n_15236), .B (si[14]), .Y (n_15235));
NAND2X1 g121016(.A (n_15236), .B (datao_2[8] ), .Y (n_15234));
NAND2X1 g121018(.A (n_15236), .B (datao_2[9] ), .Y (n_15232));
NAND2X1 g121019(.A (n_15236), .B (n_12458), .Y (n_15231));
NAND2X1 g121026(.A (n_15236), .B (si[8]), .Y (n_15230));
NAND2X1 g121028(.A (n_15236), .B (si[12]), .Y (n_15229));
NAND2X1 g121029(.A (n_15236), .B (si[13]), .Y (n_15228));
NAND2X1 g121038(.A (n_15427), .B (si[18]), .Y (n_15227));
NAND2X1 g121040(.A (n_15427), .B (si[17]), .Y (n_15226));
NAND2X1 g121075(.A (n_15240), .B (n_2638), .Y (n_15224));
NAND2X1 g121080(.A (n_15240), .B (n_4630), .Y (n_15222));
NAND2X1 g121081(.A (n_15198), .B (n_2887), .Y (n_15220));
NAND2X1 g121082(.A (n_15676), .B (n_3092), .Y (n_15218));
NAND2X1 g121084(.A (n_15240), .B (n_2167), .Y (n_15216));
NAND2X1 g121086(.A (n_15676), .B (n_4121), .Y (n_15214));
NAND2X1 g121088(.A (n_15240), .B (n_2456), .Y (n_15213));
NAND2X1 g121090(.A (n_15240), .B (n_3754), .Y (n_15212));
NAND2X1 g121091(.A (n_15676), .B (n_3809), .Y (n_15211));
NAND2X1 g121096(.A (n_15240), .B (n_3200), .Y (n_15210));
NAND2X1 g121097(.A (n_15676), .B (n_3967), .Y (n_15209));
NAND2X1 g121098(.A (n_15676), .B (n_3464), .Y (n_15208));
NAND2X1 g121104(.A (n_15240), .B (n_3469), .Y (n_15206));
NAND2X1 g121105(.A (n_15676), .B (n_4187), .Y (n_15205));
NAND2X1 g121106(.A (n_15198), .B (n_3790), .Y (n_15203));
NAND2X1 g121107(.A (n_15676), .B (n_4021), .Y (n_15202));
NAND2X1 g121108(.A (n_15676), .B (n_3948), .Y (n_15201));
NAND2X1 g121116(.A (n_15198), .B (n_4447), .Y (n_15199));
NAND2X1 g121117(.A (n_15198), .B (n_4813), .Y (n_15197));
NAND2X1 g121119(.A (n_15676), .B (n_4446), .Y (n_15196));
NAND2X1 g121121(.A (n_15676), .B (n_3525), .Y (n_15195));
AOI21X1 g121156(.A0 (n_14618), .A1 (n_22441), .B0 (n_8614), .Y(n_15194));
AOI21X1 g121158(.A0 (n_14616), .A1 (n_24121), .B0 (n_8614), .Y(n_15193));
AOI21X1 g121160(.A0 (n_14617), .A1 (n_24305), .B0 (n_8614), .Y(n_15192));
AOI21X1 g121165(.A0 (n_14615), .A1 (n_26200), .B0 (n_8614), .Y(n_15190));
NAND2X1 g121168(.A (n_14847), .B (n_14490), .Y (n_35636));
NAND2X1 g121171(.A (n_14861), .B (n_15252), .Y (n_15187));
NAND2X1 g121176(.A (n_14859), .B (n_15252), .Y (n_15186));
NAND2X1 g121178(.A (n_14855), .B (n_33629), .Y (n_15185));
NAND2X1 g121188(.A (n_14857), .B (n_15110), .Y (n_15184));
NAND2X1 g121207(.A (n_14843), .B (n_14490), .Y (n_15183));
OAI21X1 g121295(.A0 (n_23178), .A1 (n_15179), .B0 (n_23382), .Y(n_15182));
NOR2X1 g121301(.A (n_14191), .B (n_14834), .Y (n_15181));
OAI21X1 g121302(.A0 (n_15179), .A1 (n_14282), .B0 (n_23381), .Y(n_15180));
NAND2X1 g121309(.A (n_14813), .B (n_14490), .Y (n_15178));
NAND2X1 g121312(.A (n_14815), .B (n_14490), .Y (n_15177));
NAND2X1 g121314(.A (n_14827), .B (n_14743), .Y (n_15176));
NAND2X1 g121315(.A (n_14839), .B (n_15110), .Y (n_15175));
AOI21X1 g121316(.A0 (n_14569), .A1 (n_15173), .B0 (n_14641), .Y(n_15174));
NAND2X1 g121317(.A (n_14837), .B (n_15110), .Y (n_15172));
NAND3X1 g121321(.A (n_14585), .B (n_14576), .C (n_13734), .Y(n_15170));
NOR2X1 g121325(.A (n_14192), .B (n_14821), .Y (n_15169));
OAI21X1 g121337(.A0 (n_14589), .A1 (n_22477), .B0 (n_14956), .Y(n_15168));
AND2X1 g121483(.A (n_14774), .B (n_35046), .Y (n_15165));
NAND2X1 g121509(.A (n_14794), .B (n_8313), .Y (n_15164));
NAND2X1 g121511(.A (n_14802), .B (n_15110), .Y (n_15163));
NAND2X1 g121512(.A (n_14784), .B (n_24028), .Y (n_15162));
AOI21X1 g121514(.A0 (n_14547), .A1 (n_23542), .B0 (n_8614), .Y(n_15161));
AOI21X1 g121515(.A0 (n_14545), .A1 (n_26207), .B0 (n_8614), .Y(n_15160));
NAND2X1 g121516(.A (n_14804), .B (n_15110), .Y (n_15158));
NAND2X1 g121518(.A (n_14786), .B (n_8313), .Y (n_15157));
AOI21X1 g121524(.A0 (n_14540), .A1 (n_24896), .B0 (n_8614), .Y(n_15155));
AOI21X1 g121529(.A0 (n_14538), .A1 (n_24888), .B0 (n_8614), .Y(n_15154));
NAND2X1 g121538(.A (n_14798), .B (n_15110), .Y (n_15153));
NAND2X1 g121541(.A (n_14800), .B (n_15110), .Y (n_15152));
NAND2X1 g121543(.A (n_14796), .B (n_15252), .Y (n_15151));
NAND2X1 g121544(.A (n_14806), .B (n_15252), .Y (n_15150));
NAND2X1 g121545(.A (n_14808), .B (n_15252), .Y (n_15149));
NAND2X1 g121553(.A (n_14782), .B (n_15147), .Y (n_15148));
AOI21X1 g121566(.A0 (n_14536), .A1 (n_26193), .B0 (n_8614), .Y(n_15146));
INVX1 g121629(.A (n_14997), .Y (n_15145));
INVX1 g121637(.A (n_14996), .Y (n_15144));
NAND2X1 g121702(.A (n_14757), .B (n_20688), .Y (n_15143));
AOI21X1 g121709(.A0 (n_14492), .A1 (n_18815), .B0 (n_8614), .Y(n_15142));
AOI21X1 g120092(.A0 (n_15280), .A1 (n_14339), .B0 (n_14118), .Y(n_15141));
NAND2X1 g121769(.A (n_14756), .B (n_20688), .Y (n_15140));
NAND2X1 g121780(.A (n_14761), .B (n_24028), .Y (n_15139));
AOI21X1 g121787(.A0 (n_14509), .A1 (n_23043), .B0 (n_8614), .Y(n_15138));
AOI21X1 g121788(.A0 (n_14505), .A1 (n_24007), .B0 (n_8614), .Y(n_15136));
AOI21X1 g121792(.A0 (n_14504), .A1 (n_20021), .B0 (n_8614), .Y(n_15134));
AOI21X1 g121793(.A0 (n_14499), .A1 (n_23041), .B0 (n_8614), .Y(n_15133));
AOI21X1 g121795(.A0 (n_14498), .A1 (n_23242), .B0 (n_8614), .Y(n_15132));
NAND2X1 g122035(.A (n_26160), .B (n_14496), .Y (n_15131));
AOI21X1 g120091(.A0 (n_15280), .A1 (n_27091), .B0 (n_13494), .Y(n_15130));
AOI21X1 g119545(.A0 (n_15126), .A1 (n_25207), .B0 (n_13323), .Y(n_15129));
NAND2X1 g119546(.A (n_14753), .B (n_28556), .Y (n_15128));
AOI21X1 g119547(.A0 (n_15126), .A1 (n_17727), .B0 (n_13877), .Y(n_15127));
AOI21X1 g119548(.A0 (n_15121), .A1 (n_32764), .B0 (n_14291), .Y(n_15125));
AOI21X1 g119549(.A0 (n_15126), .A1 (n_13274), .B0 (n_13868), .Y(n_15123));
AOI21X1 g119621(.A0 (n_15121), .A1 (n_25290), .B0 (n_14054), .Y(n_15122));
AOI21X1 g119622(.A0 (n_15126), .A1 (n_14731), .B0 (n_15119), .Y(n_15120));
NAND2X1 g119717(.A (n_15292), .B (n_17719), .Y (n_15118));
NAND2X1 g119964(.A (n_15115), .B (n_35540), .Y (n_15117));
NAND2X1 g119972(.A (n_15115), .B (n_35736), .Y (n_15116));
NAND2X1 g119980(.A (n_15115), .B (n_18533), .Y (n_15114));
NAND2X1 g119997(.A (n_15115), .B (n_18546), .Y (n_15113));
NAND2X1 g120058(.A (n_14747), .B (n_15413), .Y (n_15112));
NAND2X1 g120059(.A (n_14750), .B (n_15110), .Y (n_15111));
NAND2X1 g120692(.A (n_14709), .B (n_14743), .Y (n_15109));
NAND2X1 g120693(.A (n_14712), .B (n_14956), .Y (n_15107));
AOI21X1 g120696(.A0 (n_14456), .A1 (n_26203), .B0 (n_8614), .Y(n_15106));
AOI21X1 g120701(.A0 (n_14455), .A1 (n_24895), .B0 (n_25067), .Y(n_15105));
AOI21X1 g120703(.A0 (n_14449), .A1 (n_34690), .B0 (n_8614), .Y(n_15104));
NAND2X1 g120704(.A (n_14705), .B (n_14956), .Y (n_15103));
NAND2X1 g120714(.A (n_14724), .B (n_15073), .Y (n_15101));
NAND2X1 g120716(.A (n_14722), .B (n_30530), .Y (n_32615));
NAND2X1 g120718(.A (n_14720), .B (n_15147), .Y (n_32908));
NAND2X1 g120721(.A (n_14728), .B (n_15110), .Y (n_15098));
NAND2X1 g120722(.A (n_14718), .B (n_11107), .Y (n_15097));
NAND2X1 g120724(.A (n_14726), .B (n_33722), .Y (n_15096));
NAND2X1 g120733(.A (n_14481), .B (n_14128), .Y (n_15095));
NAND2X1 g120741(.A (n_14703), .B (n_14956), .Y (n_15094));
AOI21X1 g120742(.A0 (n_14971), .A1 (n_25290), .B0 (n_14059), .Y(n_15092));
NAND3X1 g120767(.A (n_15090), .B (n_25309), .C (n_22821), .Y(n_27134));
NAND3X1 g120768(.A (n_15090), .B (n_15089), .C (n_22821), .Y(n_27118));
NAND2X1 g120770(.A (n_14684), .B (n_15087), .Y (n_15088));
NOR2X1 g120773(.A (n_14491), .B (n_14459), .Y (n_15257));
AOI21X1 g120803(.A0 (n_14424), .A1 (n_24190), .B0 (n_9458), .Y(n_15086));
AOI21X1 g120804(.A0 (n_15059), .A1 (n_25309), .B0 (n_14139), .Y(n_15085));
NAND2X1 g120808(.A (n_14648), .B (n_8313), .Y (n_15083));
AOI21X1 g120813(.A0 (n_14422), .A1 (n_27222), .B0 (n_8614), .Y(n_15082));
NAND2X1 g120817(.A (n_14668), .B (n_15110), .Y (n_15081));
AOI21X1 g120818(.A0 (n_14700), .A1 (n_32764), .B0 (n_14299), .Y(n_15079));
NAND2X1 g120825(.A (n_14664), .B (n_15076), .Y (n_15078));
NAND2X1 g120828(.A (n_14657), .B (n_15076), .Y (n_15077));
NAND2X1 g120831(.A (n_14645), .B (n_14743), .Y (n_15075));
NAND2X1 g120840(.A (n_14686), .B (n_15073), .Y (n_15074));
NAND2X1 g120841(.A (n_14666), .B (n_15147), .Y (n_15072));
NAND2X1 g120843(.A (n_14683), .B (n_15110), .Y (n_15071));
NAND2X1 g120845(.A (n_14675), .B (n_11107), .Y (n_15069));
NAND2X1 g120848(.A (n_14673), .B (n_15110), .Y (n_15067));
NAND2X1 g120849(.A (n_14653), .B (n_15076), .Y (n_15066));
NAND2X1 g120851(.A (n_14669), .B (n_33661), .Y (n_32231));
NAND2X1 g120852(.A (n_14652), .B (n_15076), .Y (n_15061));
AOI21X1 g120853(.A0 (n_15059), .A1 (n_15089), .B0 (n_14305), .Y(n_15060));
NAND2X1 g120854(.A (n_14677), .B (n_33629), .Y (n_15058));
NAND2X1 g120855(.A (n_14689), .B (n_27389), .Y (n_15057));
AOI21X1 g120870(.A0 (n_25290), .A1 (n_15059), .B0 (n_14055), .Y(n_15056));
AOI21X1 g120873(.A0 (n_14918), .A1 (n_25290), .B0 (n_14056), .Y(n_15055));
OAI22X1 g120910(.A0 (n_15240), .A1 (n_2051), .B0 (n_14695), .B1(n_451), .Y (n_15238));
NAND2X1 g120974(.A (n_14697), .B (n_14692), .Y (n_15338));
NAND2X1 g121002(.A (n_15236), .B (datao_2[4] ), .Y (n_15054));
NAND2X1 g121004(.A (n_15427), .B (datao_2[6] ), .Y (n_15053));
NAND2X1 g121005(.A (n_15608), .B (datao_2[7] ), .Y (n_15052));
NAND2X1 g121006(.A (n_15236), .B (datao_2[2] ), .Y (n_15051));
NAND2X1 g121008(.A (n_15427), .B (datao_2[3] ), .Y (n_15049));
NAND2X1 g121013(.A (n_15236), .B (n_12330), .Y (n_15047));
NAND2X1 g121020(.A (n_15236), .B (datao_2[10] ), .Y (n_15046));
NAND2X1 g121027(.A (n_15236), .B (si[9]), .Y (n_15045));
NAND2X1 g121044(.A (n_15608), .B (si[11]), .Y (n_15044));
NAND2X1 g121046(.A (n_15236), .B (si[10]), .Y (n_15043));
NAND2X1 g121076(.A (n_15198), .B (n_3479), .Y (n_15041));
NAND2X1 g121083(.A (n_14629), .B (n_15038), .Y (n_15039));
AOI21X1 g121149(.A0 (n_14391), .A1 (n_26209), .B0 (n_8614), .Y(n_15037));
NAND2X1 g121152(.A (n_14623), .B (n_8313), .Y (n_15036));
NAND2X1 g121155(.A (n_14637), .B (n_15110), .Y (n_15034));
NAND2X1 g121179(.A (n_14633), .B (n_30530), .Y (n_35441));
AOI21X1 g121181(.A0 (n_14386), .A1 (n_15031), .B0 (n_14641), .Y(n_15032));
NAND2X1 g121183(.A (n_14631), .B (n_15029), .Y (n_15030));
NAND2X1 g121186(.A (n_14628), .B (n_15110), .Y (n_15028));
AOI21X1 g121290(.A0 (n_14371), .A1 (n_27388), .B0 (n_15026), .Y(n_15027));
NAND2X1 g121294(.A (n_14596), .B (n_8313), .Y (n_15025));
AOI21X1 g121298(.A0 (n_14370), .A1 (n_24673), .B0 (n_15026), .Y(n_15024));
NAND3X1 g121299(.A (n_14355), .B (n_14365), .C (n_13728), .Y(n_15023));
AOI21X1 g121327(.A0 (n_14345), .A1 (n_15020), .B0 (n_14641), .Y(n_15021));
NAND2X1 g121328(.A (n_14613), .B (n_15029), .Y (n_15018));
NAND2X1 g121330(.A (n_14609), .B (n_33722), .Y (n_15017));
AOI21X1 g121332(.A0 (n_14367), .A1 (n_28542), .B0 (n_14916), .Y(n_15016));
INVX2 g121410(.A (n_15198), .Y (n_15427));
OAI21X1 g121523(.A0 (n_9563), .A1 (n_14172), .B0 (n_14554), .Y(n_15013));
AOI21X1 g121527(.A0 (n_33297), .A1 (n_32644), .B0 (n_14295), .Y(n_15011));
NAND2X1 g121531(.A (n_14559), .B (n_8313), .Y (n_15010));
NAND2X1 g121533(.A (n_14562), .B (n_15029), .Y (n_15009));
NAND2X1 g121546(.A (n_14556), .B (n_15110), .Y (n_15008));
NAND2X1 g121550(.A (n_14573), .B (n_15073), .Y (n_15007));
NAND2X1 g121554(.A (n_14571), .B (n_15029), .Y (n_15006));
NAND2X1 g121555(.A (n_14584), .B (n_15110), .Y (n_15005));
NAND2X1 g121556(.A (n_14568), .B (n_15110), .Y (n_15004));
NAND2X1 g121558(.A (n_14578), .B (n_30530), .Y (n_15003));
NAND2X1 g121559(.A (n_14566), .B (n_15110), .Y (n_15002));
NAND2X1 g121561(.A (n_14564), .B (n_15110), .Y (n_15001));
NAND2X1 g121579(.A (n_14558), .B (n_8313), .Y (n_15000));
NAND2X1 g121593(.A (n_13773), .B (n_14516), .Y (n_14999));
INVX1 g121627(.A (n_14811), .Y (n_14998));
AOI21X1 g121630(.A0 (n_14810), .A1 (n_13732), .B0 (n_14575), .Y(n_14997));
NAND2X1 g121638(.A (n_13776), .B (n_14580), .Y (n_14996));
NAND2X1 g121716(.A (n_14510), .B (n_8313), .Y (n_14995));
NAND2X1 g121814(.A (n_14543), .B (n_21550), .Y (n_14994));
OAI21X1 g121815(.A0 (n_14783), .A1 (n_32720), .B0 (n_21549), .Y(n_14993));
INVX1 g121829(.A (n_14777), .Y (n_14991));
AOI21X1 g121839(.A0 (n_9603), .A1 (n_14135), .B0 (n_14535), .Y(n_14990));
AOI21X1 g121840(.A0 (n_9603), .A1 (n_14133), .B0 (n_14529), .Y(n_14989));
NOR2X1 g121915(.A (n_14793), .B (n_32677), .Y (n_14987));
NAND2X1 g122285(.A (n_14494), .B (n_20019), .Y (n_14986));
NAND2X1 g122326(.A (n_14495), .B (n_23046), .Y (n_14985));
AOI21X1 g120037(.A0 (n_14271), .A1 (n_14983), .B0 (n_14641), .Y(n_14984));
NAND2X1 g120045(.A (n_14484), .B (n_15288), .Y (n_14982));
NAND2X1 g120053(.A (n_14483), .B (n_15076), .Y (n_14980));
AOI21X1 g120057(.A0 (n_14272), .A1 (n_14978), .B0 (n_33713), .Y(n_14979));
OAI21X1 g120388(.A0 (n_14016), .A1 (n_35485), .B0 (n_14976), .Y(n_14977));
OAI21X1 g120475(.A0 (n_33099), .A1 (n_35570), .B0 (n_14973), .Y(n_14975));
AOI21X1 g120695(.A0 (n_14971), .A1 (n_18384), .B0 (n_14306), .Y(n_14972));
OAI21X1 g120698(.A0 (n_14014), .A1 (n_32698), .B0 (n_23181), .Y(n_14970));
NAND2X1 g120702(.A (n_14476), .B (n_15076), .Y (n_14968));
NAND2X1 g120706(.A (n_14465), .B (n_15076), .Y (n_14967));
NAND2X1 g120720(.A (n_14464), .B (n_15288), .Y (n_14966));
NAND2X1 g120729(.A (n_14479), .B (n_11107), .Y (n_14965));
OAI21X1 g120730(.A0 (n_14014), .A1 (n_22042), .B0 (n_24890), .Y(n_14964));
NAND2X1 g120731(.A (n_14482), .B (n_26564), .Y (n_14963));
NAND2X1 g120736(.A (n_14480), .B (n_25683), .Y (n_14962));
NAND2X1 g120754(.A (n_14959), .B (n_23356), .Y (n_14961));
NAND2X1 g120759(.A (n_14959), .B (n_17713), .Y (n_14960));
NAND2X1 g120760(.A (n_14733), .B (n_32697), .Y (n_14958));
NAND2X1 g120763(.A (n_14959), .B (n_27950), .Y (n_14957));
NAND3X1 g120764(.A (n_14955), .B (n_24101), .C (n_14956), .Y(n_28993));
NAND3X1 g120769(.A (n_14955), .B (n_20178), .C (n_14956), .Y(n_28974));
NOR2X1 g120775(.A (n_14448), .B (n_14952), .Y (n_14953));
OAI21X1 g120778(.A0 (n_14717), .A1 (n_35494), .B0 (n_14950), .Y(n_14951));
OAI21X1 g120779(.A0 (n_14268), .A1 (n_35555), .B0 (n_14948), .Y(n_14949));
OAI21X1 g120780(.A0 (n_13796), .A1 (n_35538), .B0 (n_14946), .Y(n_14947));
NAND2X1 g120781(.A (n_14446), .B (n_14944), .Y (n_14945));
NAND3X1 g120783(.A (n_14955), .B (n_17340), .C (n_14956), .Y(n_28954));
OAI21X1 g120787(.A0 (n_13549), .A1 (n_35505), .B0 (n_14941), .Y(n_14943));
NAND2X1 g120790(.A (n_14445), .B (n_14939), .Y (n_14940));
NAND3X1 g120791(.A (n_14935), .B (n_35736), .C (n_15029), .Y(n_23201));
NAND3X1 g120797(.A (n_14935), .B (n_35540), .C (n_15110), .Y(n_22482));
NAND3X1 g120798(.A (n_14935), .B (n_18533), .C (n_11107), .Y(n_15405));
AND2X1 g120802(.A (n_14458), .B (n_28064), .Y (n_14933));
OAI21X1 g120810(.A0 (n_13551), .A1 (n_14042), .B0 (n_22839), .Y(n_14932));
NAND2X1 g120814(.A (n_14440), .B (n_14930), .Y (n_14931));
AND2X1 g120815(.A (n_14454), .B (n_28063), .Y (n_14929));
AND2X1 g120816(.A (n_14453), .B (n_24897), .Y (n_14928));
AOI21X1 g120820(.A0 (n_15059), .A1 (n_32697), .B0 (n_14100), .Y(n_14927));
AND2X1 g120821(.A (n_14450), .B (n_28061), .Y (n_14925));
AOI21X1 g120823(.A0 (n_14237), .A1 (n_25350), .B0 (n_14916), .Y(n_14924));
NAND2X1 g120832(.A (n_14431), .B (n_15076), .Y (n_14923));
OAI21X1 g120834(.A0 (n_13551), .A1 (n_22042), .B0 (n_22836), .Y(n_14922));
AOI21X1 g120846(.A0 (n_14225), .A1 (n_14920), .B0 (n_33713), .Y(n_14921));
AOI21X1 g120859(.A0 (n_14918), .A1 (n_32697), .B0 (n_14104), .Y(n_14919));
AOI21X1 g120865(.A0 (n_14234), .A1 (n_25713), .B0 (n_14916), .Y(n_14917));
NAND2X1 g121003(.A (n_14695), .B (datao_2[5] ), .Y (n_14915));
NAND2X1 g121012(.A (n_14695), .B (datao_2[1] ), .Y (n_14913));
NAND2X1 g121017(.A (n_14695), .B (si[7]), .Y (n_14912));
NAND2X1 g121031(.A (n_14695), .B (si[4]), .Y (n_14911));
NAND2X1 g121032(.A (n_14695), .B (si[5]), .Y (n_14910));
NAND2X1 g121033(.A (n_14695), .B (si[6]), .Y (n_14909));
NAND2X1 g121064(.A (n_14918), .B (n_15089), .Y (n_14908));
OAI21X1 g121079(.A0 (n_13399), .A1 (n_35546), .B0 (n_14905), .Y(n_14907));
NAND2X1 g121089(.A (n_15198), .B (n_2198), .Y (n_14904));
OAI21X1 g121099(.A0 (n_13784), .A1 (n_35505), .B0 (n_14902), .Y(n_14903));
NAND2X1 g121109(.A (n_15240), .B (n_2908), .Y (n_14901));
NAND2X1 g121110(.A (n_15240), .B (n_3966), .Y (n_14900));
NAND2X1 g121111(.A (n_15676), .B (n_3278), .Y (n_14899));
NAND2X1 g121112(.A (n_15676), .B (n_3359), .Y (n_14897));
NAND2X1 g121113(.A (n_13998), .B (n_2217), .Y (n_14896));
NAND2X1 g121114(.A (n_15240), .B (n_2768), .Y (n_14895));
NAND2X1 g121115(.A (n_15240), .B (n_2678), .Y (n_14893));
OAI21X1 g121124(.A0 (n_13531), .A1 (n_35459), .B0 (n_14889), .Y(n_14891));
OAI21X1 g121125(.A0 (n_14682), .A1 (n_35459), .B0 (n_14887), .Y(n_14888));
NAND2X1 g121128(.A (n_14417), .B (n_14885), .Y (n_14886));
OAI21X1 g121146(.A0 (n_13240), .A1 (n_35505), .B0 (n_14883), .Y(n_14884));
NAND2X1 g121157(.A (n_14423), .B (n_25351), .Y (n_14882));
NAND2X1 g121159(.A (n_14415), .B (n_15073), .Y (n_14881));
AOI21X1 g121162(.A0 (n_14655), .A1 (n_32777), .B0 (n_14112), .Y(n_14880));
NAND2X1 g121166(.A (n_14405), .B (n_14850), .Y (n_14879));
NAND2X1 g121167(.A (n_14411), .B (n_15110), .Y (n_14878));
NAND2X1 g121173(.A (n_14407), .B (n_15076), .Y (n_14877));
NAND2X1 g121174(.A (n_14403), .B (n_14956), .Y (n_14876));
NAND2X1 g121182(.A (n_14413), .B (n_33629), .Y (n_14875));
OAI21X1 g121192(.A0 (n_13536), .A1 (n_14282), .B0 (n_23136), .Y(n_14873));
NAND2X1 g121196(.A (n_14420), .B (n_23040), .Y (n_14872));
OAI21X1 g121197(.A0 (n_13536), .A1 (n_32803), .B0 (n_25264), .Y(n_14871));
AOI21X1 g121199(.A0 (n_14649), .A1 (n_32728), .B0 (n_14107), .Y(n_14870));
AOI21X1 g121200(.A0 (n_14865), .A1 (n_32794), .B0 (n_14297), .Y(n_14869));
OAI21X1 g121201(.A0 (n_13242), .A1 (n_32765), .B0 (n_23038), .Y(n_14868));
AOI21X1 g121205(.A0 (n_14862), .A1 (n_23725), .B0 (n_14303), .Y(n_14867));
AOI21X1 g121213(.A0 (n_14865), .A1 (n_18375), .B0 (n_14286), .Y(n_14866));
NAND2X1 g121214(.A (n_14421), .B (n_23045), .Y (n_14864));
AOI21X1 g121215(.A0 (n_14862), .A1 (n_18378), .B0 (n_14287), .Y(n_14863));
NAND2X1 g121228(.A (n_12297), .B (n_14418), .Y (n_15260));
OAI21X1 g121260(.A0 (n_13111), .A1 (n_35572), .B0 (n_14860), .Y(n_14861));
OAI21X1 g121264(.A0 (n_14636), .A1 (n_35459), .B0 (n_14858), .Y(n_14859));
OAI21X1 g121268(.A0 (n_13035), .A1 (n_35505), .B0 (n_14856), .Y(n_14857));
OAI21X1 g121269(.A0 (n_14385), .A1 (n_35468), .B0 (n_14854), .Y(n_14855));
NAND2X1 g121300(.A (n_14390), .B (n_21603), .Y (n_14853));
AND2X1 g121303(.A (n_14389), .B (n_24309), .Y (n_14852));
NAND2X1 g121304(.A (n_14374), .B (n_14850), .Y (n_14851));
AOI21X1 g121305(.A0 (n_14201), .A1 (n_23640), .B0 (n_14658), .Y(n_14849));
OAI21X1 g121307(.A0 (n_12975), .A1 (n_32765), .B0 (n_21602), .Y(n_14848));
OAI21X1 g121310(.A0 (n_15179), .A1 (n_32774), .B0 (n_23380), .Y(n_14847));
NAND2X1 g121322(.A (n_14383), .B (n_33661), .Y (n_14846));
NAND2X1 g121323(.A (n_14388), .B (n_33629), .Y (n_14845));
NOR2X1 g121326(.A (n_14197), .B (n_14372), .Y (n_14844));
OAI21X1 g121339(.A0 (n_15179), .A1 (n_19037), .B0 (n_14049), .Y(n_14843));
OAI21X1 g121492(.A0 (n_13497), .A1 (n_35459), .B0 (n_14838), .Y(n_14839));
OAI21X1 g121494(.A0 (n_13325), .A1 (n_35494), .B0 (n_14835), .Y(n_14837));
NAND2X1 g121513(.A (n_13964), .B (n_14318), .Y (n_14834));
NAND2X1 g121517(.A (n_14337), .B (n_14956), .Y (n_14833));
AND2X1 g121519(.A (n_14369), .B (n_28555), .Y (n_14832));
AOI21X1 g121522(.A0 (n_14179), .A1 (n_21941), .B0 (n_25563), .Y(n_14831));
NAND2X1 g121535(.A (n_14334), .B (n_15076), .Y (n_14829));
NAND2X1 g121536(.A (n_14332), .B (n_14743), .Y (n_14828));
OAI21X1 g121537(.A0 (n_13669), .A1 (n_13588), .B0 (n_28548), .Y(n_14827));
NAND2X1 g121542(.A (n_14330), .B (n_9436), .Y (n_14826));
NAND2X1 g121547(.A (n_14361), .B (n_15073), .Y (n_14825));
NAND2X1 g121548(.A (n_14359), .B (n_15073), .Y (n_14824));
NAND2X1 g121551(.A (n_14357), .B (n_15073), .Y (n_14823));
NAND2X1 g121552(.A (n_14348), .B (n_15073), .Y (n_14822));
NAND2X1 g121560(.A (n_13951), .B (n_14316), .Y (n_14821));
NAND2X1 g121562(.A (n_14363), .B (n_33629), .Y (n_14820));
OAI21X1 g121568(.A0 (n_14817), .A1 (n_23178), .B0 (n_22016), .Y(n_14819));
OAI21X1 g121570(.A0 (n_14817), .A1 (n_14042), .B0 (n_22015), .Y(n_14818));
NAND2X1 g121571(.A (n_14368), .B (n_23534), .Y (n_14816));
OAI21X1 g121573(.A0 (n_14817), .A1 (n_19037), .B0 (n_14089), .Y(n_14815));
OAI21X1 g121575(.A0 (n_13186), .A1 (n_32662), .B0 (n_23533), .Y(n_14814));
OAI21X1 g121576(.A0 (n_14817), .A1 (n_32774), .B0 (n_22013), .Y(n_14813));
NAND2X1 g121578(.A (n_14343), .B (n_15110), .Y (n_14812));
AOI21X1 g121628(.A0 (n_14810), .A1 (n_13727), .B0 (n_14350), .Y(n_14811));
NAND2X1 g121714(.A (n_14313), .B (n_15288), .Y (n_14809));
OAI21X1 g121715(.A0 (n_12830), .A1 (n_35505), .B0 (n_14807), .Y(n_14808));
OAI21X1 g121719(.A0 (n_12700), .A1 (n_35468), .B0 (n_14805), .Y(n_14806));
OAI21X1 g121730(.A0 (n_13072), .A1 (n_35505), .B0 (n_14803), .Y(n_14804));
OAI21X1 g121731(.A0 (n_12515), .A1 (n_35505), .B0 (n_14801), .Y(n_14802));
OAI21X1 g121732(.A0 (n_35394), .A1 (n_35538), .B0 (n_14799), .Y(n_14800));
OAI21X1 g121756(.A0 (n_12936), .A1 (n_35468), .B0 (n_14797), .Y(n_14798));
OAI21X1 g121775(.A0 (n_12774), .A1 (n_35505), .B0 (n_14795), .Y(n_14796));
OAI21X1 g121782(.A0 (n_14793), .A1 (n_17856), .B0 (n_27064), .Y(n_14794));
AOI21X1 g121790(.A0 (n_14131), .A1 (n_21890), .B0 (n_9971), .Y(n_14792));
AND2X1 g121797(.A (n_14326), .B (n_26202), .Y (n_14791));
AOI21X1 g121799(.A0 (n_14108), .A1 (n_20020), .B0 (n_8614), .Y(n_14790));
AOI21X1 g121800(.A0 (n_14102), .A1 (n_25051), .B0 (n_25563), .Y(n_14789));
AOI21X1 g121804(.A0 (n_14087), .A1 (n_21885), .B0 (n_9971), .Y(n_14788));
AOI21X1 g121807(.A0 (n_14076), .A1 (n_23638), .B0 (n_9971), .Y(n_14787));
NAND2X1 g121808(.A (n_14323), .B (n_24675), .Y (n_14786));
AOI21X1 g121810(.A0 (n_14079), .A1 (n_25047), .B0 (n_9971), .Y(n_14785));
OAI21X1 g121813(.A0 (n_14783), .A1 (n_23178), .B0 (n_21551), .Y(n_14784));
OAI21X1 g121826(.A0 (n_14779), .A1 (n_14635), .B0 (n_14781), .Y(n_14782));
OAI21X1 g121827(.A0 (n_14779), .A1 (n_35468), .B0 (n_14778), .Y(n_14780));
AOI22X1 g121830(.A0 (n_18289), .A1 (n_13893), .B0 (n_19494), .B1(n_10063), .Y (n_14777));
AOI21X1 g121842(.A0 (n_9603), .A1 (n_13645), .B0 (n_14322), .Y(n_14776));
AOI21X1 g121843(.A0 (n_9603), .A1 (P2_reg1[31] ), .B0 (n_14321), .Y(n_14775));
AOI22X1 g121844(.A0 (n_11610), .A1 (n_21240), .B0 (n_20218), .B1(P1_reg2[30] ), .Y (n_14774));
NAND2X1 g121909(.A (n_21677), .B (n_14121), .Y (n_14773));
NAND2X1 g121910(.A (n_21677), .B (n_14074), .Y (n_14772));
NAND2X1 g122007(.A (n_26160), .B (n_14121), .Y (n_14771));
NAND2X1 g122009(.A (n_26528), .B (n_14121), .Y (n_14769));
NAND2X1 g122011(.A (n_26160), .B (n_14074), .Y (n_14768));
NAND2X1 g122013(.A (n_26528), .B (n_14074), .Y (n_14765));
NAND3X1 g122270(.A (n_14635), .B (n_33629), .C (n_14317), .Y(n_14764));
NAND3X1 g122272(.A (n_14635), .B (P3_reg2[30] ), .C (n_33629), .Y(n_14763));
OAI21X1 g122277(.A0 (n_14503), .A1 (n_23178), .B0 (n_20022), .Y(n_14761));
OAI21X1 g122318(.A0 (n_14508), .A1 (n_32720), .B0 (n_23039), .Y(n_14759));
OAI21X1 g122319(.A0 (n_14511), .A1 (n_32698), .B0 (n_24005), .Y(n_14758));
OAI21X1 g122332(.A0 (n_14755), .A1 (n_14042), .B0 (n_17292), .Y(n_14757));
OAI21X1 g122333(.A0 (n_14755), .A1 (n_22042), .B0 (n_18809), .Y(n_14756));
NAND2X1 g119716(.A (n_15121), .B (n_18340), .Y (n_14753));
NAND2X1 g119718(.A (n_15121), .B (n_18384), .Y (n_14752));
NAND2X1 g120060(.A (n_14276), .B (n_15110), .Y (n_32297));
OAI21X1 g120389(.A0 (n_14016), .A1 (n_14749), .B0 (n_14748), .Y(n_14750));
OAI21X1 g120476(.A0 (n_33099), .A1 (n_35775), .B0 (n_14745), .Y(n_14747));
NAND2X1 g120700(.A (n_14263), .B (n_14743), .Y (n_14744));
NAND2X1 g120723(.A (n_14269), .B (n_33661), .Y (n_14742));
AOI21X1 g120726(.A0 (n_14022), .A1 (n_14740), .B0 (n_33713), .Y(n_14741));
AOI21X1 g120732(.A0 (n_14736), .A1 (n_21919), .B0 (n_13891), .Y(n_14738));
AOI21X1 g120738(.A0 (n_14736), .A1 (n_17674), .B0 (n_13484), .Y(n_14737));
NAND2X1 g120739(.A (n_14264), .B (n_15147), .Y (n_14735));
AOI21X1 g120743(.A0 (n_14733), .A1 (n_21185), .B0 (n_14072), .Y(n_14734));
AOI21X1 g120745(.A0 (n_14736), .A1 (n_14731), .B0 (n_13458), .Y(n_14732));
NAND2X2 g120747(.A (n_32899), .B (n_32900), .Y (n_15292));
INVX2 g120750(.A (n_14729), .Y (n_15300));
NAND2X2 g120753(.A (n_32051), .B (n_32052), .Y (n_15115));
OAI21X1 g120774(.A0 (n_13549), .A1 (n_14627), .B0 (n_14727), .Y(n_14728));
NAND2X1 g120776(.A (n_14252), .B (n_14725), .Y (n_14726));
NAND2X1 g120784(.A (n_14257), .B (n_14723), .Y (n_14724));
NAND2X1 g120786(.A (n_14256), .B (n_14721), .Y (n_14722));
NAND2X1 g120788(.A (n_14254), .B (n_14719), .Y (n_14720));
OAI21X1 g120792(.A0 (n_14717), .A1 (n_14749), .B0 (n_14716), .Y(n_14718));
AOI21X1 g120805(.A0 (n_14009), .A1 (n_14714), .B0 (n_33713), .Y(n_14715));
OAI21X1 g120809(.A0 (n_14708), .A1 (n_19330), .B0 (n_25852), .Y(n_14712));
AOI21X1 g120819(.A0 (n_14011), .A1 (n_24839), .B0 (n_28659), .Y(n_14711));
OAI21X1 g120822(.A0 (n_14708), .A1 (n_13781), .B0 (n_25849), .Y(n_14709));
AOI21X1 g120827(.A0 (n_14006), .A1 (n_14706), .B0 (n_14641), .Y(n_14707));
OAI21X1 g120829(.A0 (n_14708), .A1 (n_13588), .B0 (n_25850), .Y(n_14705));
NAND2X1 g120864(.A (n_14248), .B (n_15110), .Y (n_14704));
OAI21X1 g120868(.A0 (n_14708), .A1 (n_14702), .B0 (n_25856), .Y(n_14703));
AOI21X1 g120869(.A0 (n_14700), .A1 (n_18375), .B0 (n_14058), .Y(n_14701));
AOI21X1 g120871(.A0 (n_14457), .A1 (n_27770), .B0 (n_13464), .Y(n_14698));
NAND2X2 g120875(.A (n_32300), .B (n_32301), .Y (n_15280));
NAND2X1 g121034(.A (n_14695), .B (si[0]), .Y (n_14697));
NAND2X1 g121035(.A (n_14695), .B (si[1]), .Y (n_14696));
NAND2X1 g121036(.A (n_14695), .B (si[2]), .Y (n_14694));
NAND2X1 g121043(.A (n_14695), .B (si[3]), .Y (n_14693));
OR2X1 g121048(.A (n_1642), .B (n_14695), .Y (n_14692));
NAND2X1 g121059(.A (n_14687), .B (n_14690), .Y (n_14691));
NAND2X1 g121060(.A (n_14918), .B (n_18399), .Y (n_14689));
NAND2X1 g121067(.A (n_14687), .B (n_32777), .Y (n_14688));
NAND2X1 g121129(.A (n_14229), .B (n_14685), .Y (n_14686));
NAND2X1 g121130(.A (n_13996), .B (n_35790), .Y (n_14684));
OAI21X1 g121131(.A0 (n_14682), .A1 (n_35775), .B0 (n_14680), .Y(n_14683));
NAND2X1 g121134(.A (n_14224), .B (n_14678), .Y (n_14679));
NAND2X1 g121135(.A (n_14223), .B (n_14676), .Y (n_14677));
OAI21X1 g121136(.A0 (n_13399), .A1 (n_14749), .B0 (n_14674), .Y(n_14675));
OAI21X1 g121137(.A0 (n_13973), .A1 (n_14627), .B0 (n_14672), .Y(n_14673));
OAI21X1 g121139(.A0 (n_14682), .A1 (n_14384), .B0 (n_13902), .Y(n_14669));
OAI21X1 g121143(.A0 (n_13240), .A1 (n_14627), .B0 (n_14667), .Y(n_14668));
NAND2X1 g121147(.A (n_14227), .B (n_14665), .Y (n_14666));
OAI21X1 g121150(.A0 (n_13529), .A1 (n_14430), .B0 (n_25342), .Y(n_14664));
AND2X1 g121153(.A (n_14241), .B (n_25353), .Y (n_14663));
AND2X1 g121154(.A (n_14240), .B (n_25705), .Y (n_14662));
AOI21X1 g121161(.A0 (n_13986), .A1 (n_14660), .B0 (n_33713), .Y(n_14661));
AOI21X1 g121163(.A0 (n_13989), .A1 (n_22953), .B0 (n_14658), .Y(n_14659));
OAI21X1 g121172(.A0 (n_13970), .A1 (n_13432), .B0 (n_25684), .Y(n_14657));
AOI21X1 g121175(.A0 (n_14655), .A1 (n_18340), .B0 (n_13890), .Y(n_14656));
NAND2X1 g121180(.A (n_14220), .B (n_14956), .Y (n_14654));
OAI21X1 g121184(.A0 (n_13529), .A1 (n_13316), .B0 (n_25336), .Y(n_14653));
OAI21X1 g121185(.A0 (n_13970), .A1 (n_13316), .B0 (n_25679), .Y(n_14652));
AOI21X1 g121189(.A0 (n_14649), .A1 (n_25309), .B0 (n_14143), .Y(n_14650));
NAND2X1 g121191(.A (n_14239), .B (n_23042), .Y (n_14648));
AND2X1 g121193(.A (n_14238), .B (n_28213), .Y (n_14647));
AOI21X1 g121194(.A0 (n_14649), .A1 (n_23007), .B0 (n_14129), .Y(n_14646));
NAND2X1 g121203(.A (n_14232), .B (n_19492), .Y (n_14645));
AOI21X1 g121206(.A0 (n_14655), .A1 (n_18378), .B0 (n_14071), .Y(n_14644));
AOI21X1 g121211(.A0 (n_13985), .A1 (n_14642), .B0 (n_14641), .Y(n_14643));
AOI21X1 g121217(.A0 (n_14649), .A1 (n_18378), .B0 (n_14057), .Y(n_14640));
AND2X1 g121253(.A (n_14206), .B (n_14638), .Y (n_14639));
OAI21X1 g121256(.A0 (n_14636), .A1 (n_14635), .B0 (n_14634), .Y(n_14637));
NAND2X1 g121262(.A (n_14211), .B (n_14632), .Y (n_14633));
OAI21X1 g121278(.A0 (n_13111), .A1 (n_14627), .B0 (n_14630), .Y(n_14631));
NAND2X1 g121280(.A (n_14416), .B (n_18533), .Y (n_14629));
OAI21X1 g121281(.A0 (n_13035), .A1 (n_14627), .B0 (n_14626), .Y(n_14628));
AOI21X1 g121287(.A0 (n_13958), .A1 (n_14624), .B0 (n_14641), .Y(n_14625));
NAND2X1 g121293(.A (n_14214), .B (n_21604), .Y (n_14623));
NAND2X1 g121333(.A (n_14208), .B (n_11107), .Y (n_14622));
NAND2X1 g121338(.A (n_14212), .B (n_21609), .Y (n_14621));
INVX4 g121363(.A (n_15240), .Y (n_15236));
INVX4 g121388(.A (n_15676), .Y (n_15608));
OR2X1 g121464(.A (n_13227), .B (n_14282), .Y (n_14618));
OR2X1 g121466(.A (n_13227), .B (n_14537), .Y (n_14617));
OR2X1 g121467(.A (n_14614), .B (n_14544), .Y (n_14616));
OR2X1 g121475(.A (n_14614), .B (n_32646), .Y (n_14615));
OAI21X1 g121487(.A0 (n_13325), .A1 (n_14627), .B0 (n_14612), .Y(n_14613));
NAND2X1 g121497(.A (n_14199), .B (n_14610), .Y (n_14611));
NAND2X1 g121499(.A (n_14193), .B (n_14608), .Y (n_14609));
NAND2X1 g121507(.A (n_14196), .B (n_33722), .Y (n_32274));
AOI21X1 g121521(.A0 (n_13907), .A1 (n_14605), .B0 (n_33713), .Y(n_14606));
AOI21X1 g121525(.A0 (n_13927), .A1 (n_14603), .B0 (n_14641), .Y(n_14604));
NAND2X1 g121530(.A (n_14187), .B (n_14743), .Y (n_14602));
AOI21X1 g121557(.A0 (n_13909), .A1 (n_14600), .B0 (n_33713), .Y(n_14601));
NAND2X1 g121563(.A (n_14186), .B (n_15029), .Y (n_14599));
AOI21X1 g121565(.A0 (n_13930), .A1 (n_14597), .B0 (n_14641), .Y(n_14598));
NAND2X1 g121569(.A (n_14203), .B (n_23535), .Y (n_14596));
OAI21X1 g121577(.A0 (n_14373), .A1 (n_21243), .B0 (n_22842), .Y(n_14595));
OAI21X1 g121580(.A0 (n_13943), .A1 (n_14593), .B0 (n_14956), .Y(n_14594));
AOI21X1 g121581(.A0 (n_33297), .A1 (n_18375), .B0 (n_14051), .Y(n_14592));
NAND2X1 g121582(.A (n_14200), .B (n_23545), .Y (n_14590));
NOR2X1 g121692(.A (n_13669), .B (n_13147), .Y (n_14589));
NAND2X1 g121700(.A (n_14148), .B (n_14956), .Y (n_14587));
NAND2X1 g121705(.A (n_14579), .B (n_15110), .Y (n_14586));
NAND2X1 g121707(.A (n_8284), .B (n_14581), .Y (n_14585));
OAI21X1 g121721(.A0 (n_13072), .A1 (n_14635), .B0 (n_14583), .Y(n_14584));
NAND2X1 g121729(.A (n_29341), .B (n_14581), .Y (n_14582));
NAND2X1 g121736(.A (n_29505), .B (n_14579), .Y (n_14580));
NAND2X1 g121741(.A (n_14153), .B (n_14577), .Y (n_14578));
NAND2X1 g121748(.A (n_29505), .B (n_14581), .Y (n_14576));
AND2X1 g121749(.A (n_14349), .B (n_14581), .Y (n_14575));
NAND2X1 g121750(.A (n_14351), .B (n_14581), .Y (n_14574));
NAND2X1 g121755(.A (n_14152), .B (n_14572), .Y (n_14573));
OAI21X1 g121757(.A0 (n_12936), .A1 (n_14627), .B0 (n_14570), .Y(n_14571));
OR2X1 g121758(.A (n_14344), .B (n_35485), .Y (n_14569));
OAI21X1 g121759(.A0 (n_12515), .A1 (n_14635), .B0 (n_14567), .Y(n_14568));
OAI21X1 g121762(.A0 (n_12774), .A1 (n_14627), .B0 (n_14565), .Y(n_14566));
OAI21X1 g121771(.A0 (n_12700), .A1 (n_14635), .B0 (n_14563), .Y(n_14564));
OAI21X1 g121772(.A0 (n_12830), .A1 (n_14627), .B0 (n_14561), .Y(n_14562));
AOI21X1 g121796(.A0 (n_13871), .A1 (n_23641), .B0 (n_26372), .Y(n_14560));
NAND2X1 g121816(.A (n_14177), .B (n_21548), .Y (n_14559));
NAND2X1 g121823(.A (n_14176), .B (n_26216), .Y (n_14558));
OAI21X1 g121824(.A0 (n_14793), .A1 (n_21169), .B0 (n_27068), .Y(n_14557));
OAI21X1 g121825(.A0 (n_14779), .A1 (n_35775), .B0 (n_14555), .Y(n_14556));
AOI22X1 g121828(.A0 (n_10573), .A1 (n_13640), .B0 (n_14319), .B1(n_29199), .Y (n_14554));
AOI21X1 g121857(.A0 (n_14550), .A1 (P1_reg_180), .B0 (n_14164), .Y(n_14552));
AOI21X1 g121858(.A0 (n_14550), .A1 (n_13635), .B0 (n_14169), .Y(n_14551));
NAND2X1 g121903(.A (n_21677), .B (n_14533), .Y (n_14549));
NAND2X1 g121904(.A (n_21677), .B (n_14528), .Y (n_14548));
OR2X1 g121906(.A (n_14539), .B (n_14282), .Y (n_14547));
OR2X1 g121907(.A (n_13452), .B (n_14544), .Y (n_14545));
OR2X1 g121908(.A (n_14783), .B (n_14282), .Y (n_14543));
NAND2X1 g121912(.A (n_11356), .B (n_21240), .Y (n_14542));
OR2X1 g121913(.A (n_14539), .B (n_32770), .Y (n_14540));
OR2X1 g121916(.A (n_14539), .B (n_14537), .Y (n_14538));
NAND2X1 g121926(.A (n_14325), .B (n_14690), .Y (n_14536));
AND2X1 g121965(.A (n_14534), .B (n_14533), .Y (n_14535));
NAND2X1 g121966(.A (n_26160), .B (n_14533), .Y (n_14532));
NOR2X1 g121967(.A (n_18310), .B (n_8614), .Y (n_14531));
AND2X1 g121970(.A (n_14534), .B (n_14528), .Y (n_14529));
NAND2X1 g121972(.A (n_26160), .B (n_14528), .Y (n_14527));
NOR2X1 g121973(.A (n_20072), .B (n_8614), .Y (n_14526));
NAND2X1 g121974(.A (n_26528), .B (n_14528), .Y (n_14525));
NOR2X1 g122008(.A (n_13646), .B (n_8614), .Y (n_14524));
NOR2X1 g122012(.A (n_13622), .B (n_8614), .Y (n_14523));
NAND2X1 g122019(.A (n_9503), .B (n_21240), .Y (n_14522));
NAND2X1 g122037(.A (n_19494), .B (n_34802), .Y (n_14521));
NAND2X1 g122038(.A (n_19494), .B (n_14490), .Y (n_14520));
NAND2X1 g122039(.A (n_28785), .B (n_19494), .Y (n_14518));
NAND2X1 g122042(.A (n_26528), .B (n_14533), .Y (n_14517));
NAND2X1 g122242(.A (n_35485), .B (n_13341), .Y (n_15173));
NAND3X1 g122268(.A (n_35485), .B (n_29505), .C (n_14513), .Y(n_14516));
NAND3X1 g122269(.A (n_35555), .B (n_14513), .C (n_33629), .Y(n_14514));
OAI21X1 g122324(.A0 (n_14511), .A1 (n_21169), .B0 (n_24012), .Y(n_14512));
OAI21X1 g122335(.A0 (n_14755), .A1 (n_14036), .B0 (n_18814), .Y(n_14510));
OR2X1 g122435(.A (n_14508), .B (n_14537), .Y (n_14509));
OR2X1 g122450(.A (n_14511), .B (n_14537), .Y (n_14505));
OR2X1 g122489(.A (n_14503), .B (n_14544), .Y (n_14504));
OR2X1 g122540(.A (n_14508), .B (n_14544), .Y (n_14499));
OR2X1 g122548(.A (n_14511), .B (n_14282), .Y (n_14498));
OR2X1 g122649(.A (n_14508), .B (n_13823), .Y (n_14495));
OR2X1 g122672(.A (n_14503), .B (n_13823), .Y (n_14494));
OR2X1 g122813(.A (n_14755), .B (n_32677), .Y (n_14492));
NAND2X1 g122892(.A (n_32728), .B (n_14490), .Y (n_14491));
INVX1 g123273(.A (n_15089), .Y (n_17304));
NAND2X1 g120728(.A (n_14027), .B (n_13765), .Y (n_14486));
AOI21X1 g120734(.A0 (n_14274), .A1 (n_25198), .B0 (n_13880), .Y(n_14485));
OAI21X1 g120735(.A0 (n_13809), .A1 (n_17287), .B0 (n_27227), .Y(n_14484));
OAI21X1 g120737(.A0 (n_13809), .A1 (n_13434), .B0 (n_27217), .Y(n_14483));
NAND2X2 g120748(.A (n_32109), .B (n_32110), .Y (n_15126));
NAND2X1 g120752(.A (n_35434), .B (n_35435), .Y (n_14729));
NAND2X1 g120755(.A (n_14733), .B (n_17719), .Y (n_14482));
NAND2X1 g120757(.A (n_14733), .B (n_20050), .Y (n_14481));
NAND2X1 g120762(.A (n_14736), .B (n_13274), .Y (n_14480));
NAND2X1 g120796(.A (n_14019), .B (n_14478), .Y (n_14479));
AND2X1 g120806(.A (n_14026), .B (n_25706), .Y (n_14477));
OAI21X1 g120824(.A0 (n_32936), .A1 (n_13432), .B0 (n_25689), .Y(n_14476));
AOI21X1 g120837(.A0 (n_13803), .A1 (n_14473), .B0 (n_14641), .Y(n_14474));
AOI21X1 g120842(.A0 (n_13805), .A1 (n_24837), .B0 (n_14658), .Y(n_14471));
AND2X1 g120847(.A (n_14023), .B (n_25680), .Y (n_14470));
AND2X1 g120856(.A (n_14025), .B (n_28215), .Y (n_14469));
AOI21X1 g120858(.A0 (n_14466), .A1 (n_25198), .B0 (n_14080), .Y(n_14468));
AOI21X1 g120860(.A0 (n_14466), .A1 (n_23578), .B0 (n_13866), .Y(n_14467));
OAI21X1 g120861(.A0 (n_13799), .A1 (n_13432), .B0 (n_28202), .Y(n_14465));
OAI21X1 g120862(.A0 (n_13799), .A1 (n_17287), .B0 (n_28196), .Y(n_14464));
AOI21X1 g120863(.A0 (n_14466), .A1 (n_25098), .B0 (n_13485), .Y(n_14463));
AOI21X1 g120866(.A0 (n_13806), .A1 (n_24843), .B0 (n_29968), .Y(n_14462));
AND2X1 g120872(.A (n_14024), .B (n_28205), .Y (n_14461));
AOI21X1 g120874(.A0 (n_23192), .A1 (n_14466), .B0 (n_13466), .Y(n_14460));
INVX1 g121049(.A (n_14459), .Y (n_15090));
INVX1 g121051(.A (n_14259), .Y (n_14955));
INVX1 g121053(.A (n_14258), .Y (n_14935));
NAND2X1 g121058(.A (n_14457), .B (n_19577), .Y (n_14458));
NAND2X1 g121063(.A (n_14687), .B (n_20050), .Y (n_14456));
NAND2X1 g121065(.A (n_14452), .B (n_23001), .Y (n_14455));
NAND2X1 g121066(.A (n_14457), .B (n_18498), .Y (n_14454));
NAND2X1 g121068(.A (n_14452), .B (n_32652), .Y (n_14453));
NAND2X1 g121071(.A (n_14457), .B (n_17340), .Y (n_14450));
NAND2X1 g121072(.A (n_14687), .B (n_23001), .Y (n_14449));
NOR2X1 g121100(.A (n_14717), .B (n_13163), .Y (n_14448));
NAND2X1 g121127(.A (n_14444), .B (n_35500), .Y (n_14446));
NAND2X1 g121133(.A (n_14444), .B (n_35736), .Y (n_14445));
NAND2X1 g121141(.A (n_14444), .B (n_18533), .Y (n_14442));
NAND2X1 g121145(.A (n_14444), .B (n_14439), .Y (n_14440));
AOI21X1 g121170(.A0 (n_13789), .A1 (n_27710), .B0 (n_14916), .Y(n_14436));
AOI21X1 g121177(.A0 (n_13787), .A1 (n_22952), .B0 (n_14658), .Y(n_14435));
NAND2X1 g121187(.A (n_14002), .B (n_14956), .Y (n_14434));
AND2X1 g121195(.A (n_14012), .B (n_27716), .Y (n_14433));
AOI21X1 g121202(.A0 (n_14425), .A1 (n_27091), .B0 (n_13490), .Y(n_14432));
OAI21X1 g121204(.A0 (n_13785), .A1 (n_14430), .B0 (n_24299), .Y(n_14431));
AOI21X1 g121208(.A0 (n_13790), .A1 (n_25355), .B0 (n_14916), .Y(n_14429));
NAND2X1 g121210(.A (n_13999), .B (n_9436), .Y (n_14428));
AOI21X1 g121216(.A0 (n_14425), .A1 (n_14731), .B0 (n_13457), .Y(n_14426));
NAND2X1 g121229(.A (n_12151), .B (n_14008), .Y (n_14959));
NAND2X1 g121237(.A (n_14865), .B (n_18340), .Y (n_14424));
NAND2X1 g121241(.A (n_14655), .B (n_18384), .Y (n_14423));
NAND2X1 g121244(.A (n_14865), .B (n_18384), .Y (n_14422));
NAND2X1 g121248(.A (n_14419), .B (n_22786), .Y (n_14421));
NAND2X1 g121250(.A (n_14419), .B (n_20050), .Y (n_14420));
NAND2X1 g121255(.A (n_14260), .B (n_13966), .Y (n_14418));
NAND2X1 g121267(.A (n_14416), .B (n_35540), .Y (n_14417));
NAND2X1 g121270(.A (n_13984), .B (n_14414), .Y (n_14415));
NAND2X1 g121275(.A (n_13987), .B (n_14412), .Y (n_14413));
NAND2X1 g121277(.A (n_13981), .B (n_14410), .Y (n_14411));
AOI21X1 g121289(.A0 (n_13783), .A1 (n_23642), .B0 (n_14916), .Y(n_14409));
AND2X1 g121292(.A (n_13993), .B (n_25055), .Y (n_14408));
OAI21X1 g121296(.A0 (n_14001), .A1 (n_14430), .B0 (n_27709), .Y(n_14407));
AND2X1 g121297(.A (n_13991), .B (n_27718), .Y (n_14406));
OAI21X1 g121306(.A0 (n_14219), .A1 (n_14404), .B0 (n_24006), .Y(n_14405));
OAI21X1 g121308(.A0 (n_13992), .A1 (n_13434), .B0 (n_25345), .Y(n_14403));
NAND2X1 g121313(.A (n_13977), .B (n_9436), .Y (n_14401));
AOI21X1 g121318(.A0 (n_13779), .A1 (n_23637), .B0 (n_14658), .Y(n_14400));
NAND2X1 g121331(.A (n_13979), .B (n_14398), .Y (n_14399));
AOI21X1 g121334(.A0 (n_13780), .A1 (n_23647), .B0 (n_29968), .Y(n_14397));
OAI21X1 g121335(.A0 (n_13227), .A1 (n_24013), .B0 (n_24324), .Y(n_14395));
OAI21X1 g121336(.A0 (n_14614), .A1 (n_24013), .B0 (n_26197), .Y(n_14394));
INVX8 g121397(.A (n_14695), .Y (n_15676));
INVX4 g121401(.A (n_14695), .Y (n_15240));
INVX4 g121415(.A (n_14695), .Y (n_15198));
OR2X1 g121461(.A (n_14614), .B (n_13571), .Y (n_14391));
NAND2X1 g121468(.A (n_14213), .B (n_18918), .Y (n_14390));
NAND2X1 g121469(.A (n_13228), .B (n_32794), .Y (n_14389));
NAND2X1 g121481(.A (n_13955), .B (n_14387), .Y (n_14388));
OR2X1 g121486(.A (n_14385), .B (n_14384), .Y (n_14386));
NAND2X1 g121490(.A (n_13956), .B (n_14382), .Y (n_14383));
NAND2X1 g121508(.A (n_13945), .B (n_9436), .Y (n_14381));
NAND2X1 g121532(.A (n_13946), .B (n_14956), .Y (n_14380));
AOI21X1 g121534(.A0 (n_13755), .A1 (n_21939), .B0 (n_29968), .Y(n_14379));
NAND2X1 g121539(.A (n_13948), .B (n_15288), .Y (n_14377));
AOI21X1 g121564(.A0 (n_13717), .A1 (n_14375), .B0 (n_33713), .Y(n_14376));
OAI21X1 g121572(.A0 (n_14373), .A1 (n_14404), .B0 (n_22844), .Y(n_14374));
NAND2X1 g121610(.A (n_13959), .B (n_9034), .Y (n_14372));
NAND2X1 g121686(.A (n_33297), .B (n_17719), .Y (n_14371));
NAND2X1 g121688(.A (n_33297), .B (n_18384), .Y (n_14370));
NAND2X1 g121689(.A (n_14366), .B (n_28441), .Y (n_14369));
NAND2X1 g121690(.A (n_14202), .B (n_18918), .Y (n_14368));
NAND2X1 g121696(.A (n_14366), .B (n_23356), .Y (n_14367));
NAND2X1 g121698(.A (n_29505), .B (n_14353), .Y (n_14365));
NAND2X1 g121738(.A (n_13908), .B (n_14362), .Y (n_14363));
NAND2X1 g121739(.A (n_13935), .B (n_14360), .Y (n_14361));
NAND2X1 g121740(.A (n_13924), .B (n_14358), .Y (n_14359));
NAND2X1 g121743(.A (n_13919), .B (n_14356), .Y (n_14357));
NAND2X1 g121744(.A (n_13952), .B (n_14353), .Y (n_14355));
NAND2X1 g121745(.A (n_29341), .B (n_14353), .Y (n_14354));
NAND2X1 g121746(.A (n_14351), .B (n_14353), .Y (n_14352));
AND2X1 g121747(.A (n_14349), .B (n_14353), .Y (n_14350));
NAND2X1 g121752(.A (n_13914), .B (n_14347), .Y (n_14348));
NAND2X1 g121754(.A (n_13894), .B (n_15288), .Y (n_14346));
OR2X1 g121770(.A (n_14344), .B (n_14384), .Y (n_14345));
NAND2X1 g121781(.A (n_13939), .B (n_13518), .Y (n_14343));
AOI21X1 g121783(.A0 (n_13664), .A1 (n_23643), .B0 (n_14916), .Y(n_14342));
AOI21X1 g121784(.A0 (n_13660), .A1 (n_25056), .B0 (n_14916), .Y(n_14341));
AOI21X1 g121789(.A0 (n_13454), .A1 (n_14339), .B0 (n_13655), .Y(n_14340));
OAI21X1 g121791(.A0 (n_14331), .A1 (n_14404), .B0 (n_27717), .Y(n_14337));
NAND2X1 g121798(.A (n_13932), .B (n_14335), .Y (n_14336));
OAI21X1 g121802(.A0 (n_35944), .A1 (n_13434), .B0 (n_26787), .Y(n_14334));
AOI21X1 g121803(.A0 (n_13620), .A1 (n_21892), .B0 (n_14916), .Y(n_14333));
OAI21X1 g121805(.A0 (n_14331), .A1 (n_19165), .B0 (n_27708), .Y(n_14332));
OAI21X1 g121812(.A0 (n_14178), .A1 (n_14430), .B0 (n_21940), .Y(n_14330));
NAND2X1 g121818(.A (n_13896), .B (n_14743), .Y (n_14329));
AOI21X1 g121819(.A0 (n_13632), .A1 (n_25058), .B0 (n_29968), .Y(n_14328));
OAI21X1 g121822(.A0 (n_14539), .A1 (n_24013), .B0 (n_24894), .Y(n_14327));
NAND2X1 g121914(.A (n_14325), .B (n_32723), .Y (n_14326));
NAND2X1 g121923(.A (n_13455), .B (n_23270), .Y (n_14323));
AND2X1 g122006(.A (n_14534), .B (n_14121), .Y (n_14322));
AND2X1 g122010(.A (n_14534), .B (n_14074), .Y (n_14321));
NAND2X1 g122022(.A (n_14319), .B (n_26870), .Y (n_14320));
NAND2X1 g122202(.A (n_14384), .B (n_565), .Y (n_14781));
NAND2X1 g122233(.A (n_14635), .B (P3_reg2[29] ), .Y (n_15038));
NAND3X1 g122261(.A (n_14635), .B (n_14317), .C (n_8966), .Y(n_14318));
NAND3X1 g122271(.A (n_14635), .B (P3_reg2[30] ), .C (n_8966), .Y(n_14316));
OAI21X1 g122334(.A0 (n_14147), .A1 (n_14430), .B0 (n_19328), .Y(n_14313));
INVX1 g122437(.A (n_23535), .Y (n_14506));
INVX1 g122451(.A (n_14307), .Y (n_17292));
INVX1 g122478(.A (n_25590), .Y (n_14306));
INVX1 g122511(.A (n_26924), .Y (n_14305));
INVX1 g122517(.A (n_28554), .Y (n_14304));
INVX1 g122522(.A (n_25260), .Y (n_14303));
INVX1 g122575(.A (n_25696), .Y (n_14299));
INVX1 g122586(.A (n_20020), .Y (n_14298));
INVX1 g122592(.A (n_27219), .Y (n_14297));
INVX1 g122600(.A (n_27379), .Y (n_14295));
INVX1 g122611(.A (n_21549), .Y (n_14497));
INVX1 g122616(.A (n_14097), .Y (n_14496));
INVX1 g122653(.A (n_28549), .Y (n_14292));
INVX1 g122662(.A (n_28551), .Y (n_14291));
INVX1 g122721(.A (n_27059), .Y (n_15352));
INVX1 g122900(.A (n_25271), .Y (n_14287));
INVX1 g122916(.A (n_27230), .Y (n_14286));
INVX4 g123274(.A (n_14282), .Y (n_15089));
INVX2 g123662(.A (n_14690), .Y (n_14279));
INVX2 g123666(.A (n_22052), .Y (n_19024));
OAI21X1 g120477(.A0 (n_33099), .A1 (n_14267), .B0 (n_13911), .Y(n_14276));
AOI21X1 g120744(.A0 (n_14274), .A1 (n_23192), .B0 (n_13467), .Y(n_14275));
NAND2X1 g120746(.A (n_35698), .B (n_35699), .Y (n_15121));
NAND2X1 g120766(.A (n_13413), .B (n_13810), .Y (n_32899));
NAND2X1 g120785(.A (n_14270), .B (n_35816), .Y (n_14272));
NAND2X1 g120789(.A (n_14270), .B (n_14439), .Y (n_14271));
OAI21X1 g120793(.A0 (n_14268), .A1 (n_14267), .B0 (n_14266), .Y(n_14269));
NAND2X1 g120801(.A (n_13075), .B (n_13807), .Y (n_32051));
NAND2X1 g120830(.A (n_13811), .B (n_13520), .Y (n_14264));
OAI21X1 g120867(.A0 (n_32936), .A1 (n_14261), .B0 (n_25693), .Y(n_14263));
NAND3X1 g121050(.A (n_14260), .B (n_13407), .C (n_13548), .Y(n_14459));
NAND3X1 g121052(.A (n_14007), .B (n_13546), .C (n_13545), .Y(n_14259));
NAND2X1 g121054(.A (n_13791), .B (n_8744), .Y (n_14258));
OR2X1 g121074(.A (n_13549), .B (n_35775), .Y (n_14257));
OR2X1 g121078(.A (n_14268), .B (n_35840), .Y (n_14256));
NAND2X1 g121123(.A (n_13555), .B (n_13800), .Y (n_32300));
OR2X1 g121132(.A (n_13796), .B (n_35768), .Y (n_14254));
NAND2X1 g121140(.A (n_14018), .B (n_18533), .Y (n_14252));
NAND2X1 g121151(.A (n_13802), .B (n_14956), .Y (n_14249));
NAND2X1 g121169(.A (n_13804), .B (n_14247), .Y (n_14248));
AOI21X1 g121198(.A0 (n_14242), .A1 (n_25098), .B0 (n_13482), .Y(n_14246));
AOI21X1 g121209(.A0 (n_13542), .A1 (n_22960), .B0 (n_29968), .Y(n_14244));
AOI21X1 g121212(.A0 (n_14242), .A1 (n_23192), .B0 (n_13469), .Y(n_14243));
NAND2X1 g121238(.A (n_14236), .B (n_25554), .Y (n_14241));
NAND2X1 g121239(.A (n_14233), .B (n_28441), .Y (n_14240));
NAND2X1 g121240(.A (n_14419), .B (n_18399), .Y (n_14239));
NAND2X1 g121242(.A (n_14425), .B (n_24105), .Y (n_14238));
NAND2X1 g121246(.A (n_14236), .B (n_14235), .Y (n_14237));
NAND2X1 g121247(.A (n_14233), .B (n_14235), .Y (n_14234));
NAND2X1 g121251(.A (n_14425), .B (n_23578), .Y (n_14232));
NAND2X1 g121259(.A (n_14226), .B (n_18533), .Y (n_14230));
OR2X1 g121271(.A (n_13784), .B (n_35775), .Y (n_14229));
NAND2X1 g121272(.A (n_14226), .B (n_35822), .Y (n_14227));
NAND2X1 g121273(.A (n_13974), .B (n_13957), .Y (n_14225));
NAND2X1 g121274(.A (n_14416), .B (n_35794), .Y (n_14224));
OR2X1 g121276(.A (n_13240), .B (n_35719), .Y (n_14223));
NOR2X1 g121286(.A (n_13786), .B (n_14221), .Y (n_14222));
OAI21X1 g121320(.A0 (n_14219), .A1 (n_14218), .B0 (n_24003), .Y(n_14220));
INVX4 g121416(.A (n_13998), .Y (n_14695));
INVX1 g121432(.A (n_14700), .Y (n_14217));
NAND2X1 g121463(.A (n_14213), .B (n_18399), .Y (n_14214));
NAND2X1 g121473(.A (n_14213), .B (n_23791), .Y (n_14212));
OR2X1 g121496(.A (n_14636), .B (n_35775), .Y (n_14211));
NOR2X1 g121510(.A (n_13778), .B (n_14209), .Y (n_14210));
NAND2X1 g121549(.A (n_13767), .B (n_14207), .Y (n_14208));
AOI22X1 g121619(.A0 (n_14349), .A1 (n_13960), .B0 (n_11138), .B1(P3_reg2[30] ), .Y (n_14206));
AOI21X1 g121626(.A0 (n_14810), .A1 (n_14168), .B0 (n_13768), .Y(n_14204));
NAND2X1 g121687(.A (n_14202), .B (n_18399), .Y (n_14203));
OR2X1 g121691(.A (n_13782), .B (n_13845), .Y (n_14201));
NAND2X1 g121693(.A (n_14202), .B (n_23791), .Y (n_14200));
OR2X1 g121704(.A (n_13496), .B (n_35830), .Y (n_14199));
AOI21X1 g121713(.A0 (n_13470), .A1 (n_19327), .B0 (n_26372), .Y(n_14198));
INVX1 g121717(.A (n_13962), .Y (n_14197));
OAI21X1 g121760(.A0 (n_35394), .A1 (n_14267), .B0 (n_14194), .Y(n_14196));
NAND2X1 g121761(.A (n_13766), .B (n_18533), .Y (n_14193));
INVX1 g121763(.A (n_13953), .Y (n_14192));
INVX1 g121767(.A (n_13949), .Y (n_14191));
NOR2X1 g121773(.A (n_13372), .B (n_25881), .Y (n_14190));
AND2X1 g121786(.A (n_13760), .B (n_25053), .Y (n_14189));
AND2X1 g121801(.A (n_13757), .B (n_25048), .Y (n_14188));
OAI21X1 g121809(.A0 (n_14331), .A1 (n_13318), .B0 (n_27702), .Y(n_14187));
NAND2X1 g121817(.A (n_13712), .B (n_14185), .Y (n_14186));
AOI21X1 g121821(.A0 (n_13454), .A1 (n_24361), .B0 (n_14182), .Y(n_14184));
AOI21X1 g121835(.A0 (n_14550), .A1 (P1_reg1[30] ), .B0 (n_13749), .Y(n_14181));
AOI21X1 g121836(.A0 (n_14550), .A1 (n_13322), .B0 (n_13744), .Y(n_14180));
OR2X1 g121911(.A (n_14178), .B (n_17293), .Y (n_14179));
NAND2X1 g121919(.A (n_12775), .B (n_24984), .Y (n_14177));
NAND2X1 g121922(.A (n_14325), .B (n_23791), .Y (n_14176));
NAND2X1 g121936(.A (n_35600), .B (n_13388), .Y (n_28125));
NAND2X1 g121979(.A (n_13901), .B (n_13498), .Y (n_14563));
NAND2X1 g121985(.A (n_13901), .B (P3_reg2[10] ), .Y (n_14630));
NAND2X1 g121987(.A (n_35583), .B (n_13211), .Y (n_14801));
NAND2X1 g121991(.A (n_35602), .B (n_13351), .Y (n_14944));
NOR2X1 g122023(.A (n_14172), .B (n_9435), .Y (n_14173));
NAND2X1 g122024(.A (n_35590), .B (n_13365), .Y (n_14976));
NAND2X1 g122032(.A (n_35555), .B (n_13204), .Y (n_14860));
NAND2X1 g122048(.A (n_35529), .B (n_13213), .Y (n_14902));
NAND2X1 g122055(.A (n_35555), .B (n_13212), .Y (n_14858));
NAND2X1 g122060(.A (n_35590), .B (n_13359), .Y (n_14889));
NAND2X1 g122066(.A (n_35529), .B (n_13199), .Y (n_14941));
NOR2X1 g122067(.A (n_13748), .B (n_21293), .Y (n_14169));
AND2X1 g122074(.A (n_35514), .B (n_14168), .Y (n_14579));
NAND2X1 g122079(.A (n_35590), .B (n_13215), .Y (n_14778));
NAND2X1 g122081(.A (n_35485), .B (n_13373), .Y (n_14905));
NAND2X1 g122082(.A (n_35583), .B (n_13200), .Y (n_14797));
NAND2X1 g122084(.A (n_35463), .B (n_13203), .Y (n_14948));
NAND2X1 g122085(.A (n_35463), .B (n_13377), .Y (n_14950));
NAND2X1 g122086(.A (n_35602), .B (n_13216), .Y (n_14803));
NAND2X1 g122092(.A (n_35464), .B (n_13367), .Y (n_14799));
NAND2X1 g122094(.A (n_35464), .B (n_13357), .Y (n_14887));
NAND2X1 g122097(.A (n_35464), .B (n_13355), .Y (n_14973));
NAND2X1 g122100(.A (n_35580), .B (n_13354), .Y (n_14946));
NAND2X1 g122103(.A (n_35464), .B (n_13353), .Y (n_14838));
NAND2X1 g122105(.A (n_35583), .B (n_13348), .Y (n_15302));
NOR2X1 g122106(.A (n_13748), .B (n_22097), .Y (n_14164));
OR2X1 g122109(.A (n_14162), .B (n_22097), .Y (n_14163));
NOR2X1 g122110(.A (n_22097), .B (n_29968), .Y (n_14161));
NOR2X1 g122112(.A (n_14159), .B (n_22097), .Y (n_14160));
NAND2X1 g122114(.A (n_35463), .B (n_13330), .Y (n_14885));
NAND2X1 g122117(.A (n_35555), .B (n_13209), .Y (n_14795));
OR2X1 g122118(.A (n_14162), .B (n_21293), .Y (n_14158));
NOR2X1 g122119(.A (n_21293), .B (n_8945), .Y (n_14157));
NOR2X1 g122124(.A (n_14159), .B (n_21293), .Y (n_14155));
NAND2X1 g122127(.A (n_35580), .B (n_13208), .Y (n_14805));
NAND2X1 g122128(.A (n_35580), .B (n_13205), .Y (n_14835));
NAND2X1 g122130(.A (n_35580), .B (n_13207), .Y (n_14883));
NAND2X1 g122133(.A (n_35485), .B (n_13340), .Y (n_14854));
NAND2X1 g122135(.A (n_35583), .B (n_13206), .Y (n_14807));
INVX1 g122146(.A (n_26371), .Y (n_14154));
NAND2X1 g122151(.A (n_35555), .B (n_13202), .Y (n_14856));
NAND2X1 g122158(.A (n_13154), .B (n_35790), .Y (n_14153));
OR2X1 g122174(.A (n_12830), .B (n_35834), .Y (n_14152));
INVX1 g122178(.A (n_29694), .Y (n_14151));
INVX1 g122190(.A (n_14150), .Y (n_14581));
NAND2X1 g122195(.A (n_35463), .B (n_524), .Y (n_15415));
NAND2X1 g122207(.A (n_13901), .B (P3_reg2[13] ), .Y (n_14570));
NAND2X1 g122214(.A (n_13901), .B (n_13337), .Y (n_14567));
OAI21X1 g122328(.A0 (n_14147), .A1 (n_19330), .B0 (n_19329), .Y(n_14148));
INVX1 g122386(.A (n_34500), .Y (n_24190));
NAND2X1 g122392(.A (n_13820), .B (P2_reg_107), .Y (n_26564));
INVX1 g122399(.A (n_14141), .Y (n_19494));
INVX1 g122405(.A (n_26925), .Y (n_14139));
NAND2X1 g122410(.A (n_14123), .B (n_9132), .Y (n_28556));
AND2X1 g122422(.A (n_14134), .B (n_14135), .Y (n_14533));
NAND2X1 g122423(.A (n_26210), .B (n_14135), .Y (n_18310));
AND2X1 g122425(.A (n_14134), .B (n_14133), .Y (n_14528));
NAND2X1 g122426(.A (n_13817), .B (n_14133), .Y (n_20072));
INVX1 g122429(.A (n_21604), .Y (n_14311));
NAND2X1 g122438(.A (n_24889), .B (n_9597), .Y (n_23535));
INVX1 g122441(.A (n_23042), .Y (n_14309));
NAND2X2 g122445(.A (n_14134), .B (n_9592), .Y (n_23382));
AND2X1 g122453(.A (n_26204), .B (n_9590), .Y (n_14307));
NAND2X1 g122466(.A (n_13840), .B (P2_reg1[12] ), .Y (n_25351));
NAND2X1 g122479(.A (n_13838), .B (P2_reg1[15] ), .Y (n_25590));
NAND2X1 g122481(.A (n_13839), .B (P2_reg1[16] ), .Y (n_25702));
OR2X1 g122482(.A (n_14086), .B (n_14101), .Y (n_14131));
NAND2X1 g122503(.A (n_26204), .B (P2_reg1[23] ), .Y (n_14128));
NAND2X1 g122506(.A (n_14124), .B (n_9231), .Y (n_27384));
INVX1 g122507(.A (n_14125), .Y (n_14126));
INVX1 g122508(.A (n_14125), .Y (n_24673));
NAND2X1 g122512(.A (n_14124), .B (n_9142), .Y (n_26924));
NAND2X1 g122518(.A (n_14116), .B (n_9081), .Y (n_28554));
NAND2X1 g122523(.A (n_14123), .B (n_9773), .Y (n_25260));
INVX1 g122536(.A (n_14118), .Y (n_14117));
NAND2X1 g122541(.A (n_26204), .B (P2_reg1[6] ), .Y (n_23534));
NAND2X1 g122543(.A (n_14116), .B (n_4237), .Y (n_23040));
NAND2X1 g122544(.A (n_13842), .B (P2_reg1[8] ), .Y (n_23381));
INVX2 g122550(.A (n_20173), .Y (n_21240));
NAND2X2 g122553(.A (n_32675), .B (P2_reg2[10] ), .Y (n_24309));
NAND2X2 g122567(.A (n_32654), .B (n_4160), .Y (n_24896));
NAND2X1 g122568(.A (n_32709), .B (n_4367), .Y (n_25264));
INVX1 g122572(.A (n_14109), .Y (n_23181));
NAND2X1 g122576(.A (n_32767), .B (P2_reg2[16] ), .Y (n_25696));
NAND2X2 g122582(.A (n_14134), .B (n_9549), .Y (n_18809));
NAND2X2 g122583(.A (n_32654), .B (P2_reg2[19] ), .Y (n_26199));
NAND2X2 g122584(.A (n_32718), .B (P2_reg2[11] ), .Y (n_24897));
OR2X1 g122585(.A (n_14503), .B (n_32646), .Y (n_14108));
NAND2X1 g122587(.A (n_32649), .B (P2_reg2[1] ), .Y (n_20020));
INVX1 g122589(.A (n_27220), .Y (n_14107));
NAND2X1 g122594(.A (n_32720), .B (n_10610), .Y (n_27219));
NAND2X1 g122595(.A (n_32767), .B (n_10043), .Y (n_26558));
INVX1 g122596(.A (n_27380), .Y (n_14104));
OR2X1 g122599(.A (n_14078), .B (n_14101), .Y (n_14102));
NAND2X1 g122601(.A (n_32646), .B (n_10607), .Y (n_27379));
INVX1 g122603(.A (n_26923), .Y (n_14100));
NAND2X2 g122612(.A (n_32649), .B (P2_reg2[2] ), .Y (n_21549));
NAND2X1 g122617(.A (n_14096), .B (n_32711), .Y (n_14097));
NAND2X1 g122618(.A (n_32719), .B (P2_reg2[3] ), .Y (n_21602));
INVX1 g122619(.A (n_22013), .Y (n_14094));
NAND2X1 g122624(.A (n_32707), .B (n_3724), .Y (n_23533));
NAND2X1 g122625(.A (n_32719), .B (n_4344), .Y (n_23038));
NAND2X2 g122627(.A (n_32802), .B (P2_reg2[9] ), .Y (n_24005));
INVX1 g122641(.A (n_14090), .Y (n_22836));
NAND2X2 g122654(.A (n_32654), .B (n_10653), .Y (n_28549));
NAND2X1 g122663(.A (n_32720), .B (n_10602), .Y (n_28551));
OR2X1 g122665(.A (n_14086), .B (n_13437), .Y (n_14087));
NAND2X2 g122681(.A (n_14134), .B (n_9565), .Y (n_25675));
OR2X1 g122702(.A (n_14078), .B (n_13437), .Y (n_14079));
NAND2X1 g122706(.A (n_14116), .B (P2_reg1[3] ), .Y (n_21603));
NAND2X1 g122723(.A (n_32745), .B (n_10613), .Y (n_27059));
OR2X1 g122724(.A (n_13895), .B (n_13437), .Y (n_14076));
INVX1 g122739(.A (n_26569), .Y (n_14072));
INVX1 g122746(.A (n_25344), .Y (n_14071));
NAND2X1 g122896(.A (n_7664), .B (n_13826), .Y (n_24895));
NAND2X1 g122901(.A (n_3100), .B (n_13823), .Y (n_25271));
INVX1 g122902(.A (n_24892), .Y (n_14059));
INVX1 g122905(.A (n_34800), .Y (n_14058));
NAND2X1 g122918(.A (n_9209), .B (n_13823), .Y (n_27230));
INVX1 g122924(.A (n_26376), .Y (n_14057));
INVX1 g122926(.A (n_27377), .Y (n_14056));
INVX1 g122933(.A (n_26929), .Y (n_14055));
INVX1 g122937(.A (n_28572), .Y (n_14054));
INVX1 g122939(.A (n_28570), .Y (n_14053));
NAND2X1 g122954(.A (n_13826), .B (n_8193), .Y (n_23045));
NAND2X1 g122962(.A (n_13826), .B (n_8205), .Y (n_23545));
INVX1 g122967(.A (n_27399), .Y (n_14051));
INVX4 g123276(.A (n_14045), .Y (n_14282));
INVX2 g123283(.A (n_23270), .Y (n_14042));
INVX1 g123290(.A (n_18918), .Y (n_18429));
INVX2 g123293(.A (n_18918), .Y (n_14544));
INVX1 g123551(.A (n_14036), .Y (n_20154));
INVX2 g123552(.A (n_14036), .Y (n_18907));
INVX1 g123580(.A (n_22786), .Y (n_19037));
INVX1 g123589(.A (n_23001), .Y (n_17848));
INVX1 g123596(.A (n_18378), .Y (n_18441));
INVX1 g123631(.A (n_21627), .Y (n_14537));
INVX2 g123636(.A (n_22412), .Y (n_22042));
INVX1 g123649(.A (n_18340), .Y (n_17856));
INVX1 g123665(.A (n_14032), .Y (n_14690));
INVX1 g123667(.A (n_14032), .Y (n_22052));
INVX4 g123671(.A (n_25309), .Y (n_23178));
NAND2X1 g121311(.A (n_13526), .B (rd_3), .Y (rd));
NAND2X1 g120771(.A (n_13540), .B (n_13558), .Y (n_32109));
NAND2X1 g120782(.A (n_13416), .B (n_13557), .Y (n_35434));
OR2X1 g120795(.A (n_33099), .B (n_13214), .Y (n_14027));
OR2X1 g121061(.A (n_32936), .B (n_13990), .Y (n_14026));
OR2X1 g121062(.A (n_13553), .B (n_13283), .Y (n_14025));
NAND2X1 g121069(.A (n_13798), .B (n_27770), .Y (n_14024));
OR2X1 g121070(.A (n_32936), .B (n_13184), .Y (n_14023));
NAND2X1 g121087(.A (n_13793), .B (n_13957), .Y (n_14022));
NAND2X1 g121144(.A (n_14018), .B (n_14439), .Y (n_14019));
AOI21X1 g121190(.A0 (n_14010), .A1 (n_18065), .B0 (n_13491), .Y(n_14017));
NAND2X1 g121220(.A (n_35883), .B (n_35884), .Y (n_14736));
INVX1 g121224(.A (n_14270), .Y (n_14016));
INVX1 g121230(.A (n_14971), .Y (n_14014));
NAND2X1 g121243(.A (n_14242), .B (n_28441), .Y (n_14012));
NAND2X1 g121245(.A (n_14010), .B (n_17727), .Y (n_14011));
OR2X1 g121263(.A (n_13399), .B (n_35719), .Y (n_14009));
NAND2X1 g121266(.A (n_14007), .B (n_13525), .Y (n_14008));
NAND2X1 g121279(.A (n_13396), .B (n_13957), .Y (n_14006));
NAND2X1 g121283(.A (n_13530), .B (n_14439), .Y (n_14005));
AOI21X1 g121288(.A0 (n_13988), .A1 (n_18065), .B0 (n_13492), .Y(n_14003));
OAI21X1 g121329(.A0 (n_14001), .A1 (n_13317), .B0 (n_27705), .Y(n_14002));
OAI21X1 g121340(.A0 (n_14219), .A1 (n_13976), .B0 (n_24011), .Y(n_13999));
NAND2X2 g121417(.A (n_13524), .B (n_13537), .Y (n_13998));
NAND2X1 g121434(.A (n_11512), .B (n_13538), .Y (n_14700));
INVX1 g121436(.A (n_13996), .Y (n_14717));
NAND2X1 g121443(.A (n_11958), .B (n_13541), .Y (n_14457));
INVX1 g121444(.A (n_13994), .Y (n_14708));
NAND2X1 g121447(.A (n_32250), .B (n_32251), .Y (n_14444));
INVX1 g121454(.A (n_33746), .Y (n_17655));
OR2X1 g121462(.A (n_13992), .B (n_13283), .Y (n_13993));
OR2X1 g121465(.A (n_14001), .B (n_13990), .Y (n_13991));
NAND2X1 g121470(.A (n_13988), .B (n_17727), .Y (n_13989));
OR2X1 g121480(.A (n_13035), .B (n_35824), .Y (n_13987));
NAND2X1 g121484(.A (n_13983), .B (n_13957), .Y (n_13986));
NAND2X1 g121489(.A (n_13108), .B (n_13957), .Y (n_13985));
NAND2X1 g121495(.A (n_13983), .B (n_35744), .Y (n_13984));
OR2X1 g121498(.A (n_14385), .B (n_35766), .Y (n_13981));
NAND2X1 g121503(.A (n_13523), .B (n_14439), .Y (n_13979));
OAI21X1 g121567(.A0 (n_14373), .A1 (n_13317), .B0 (n_22760), .Y(n_13978));
OAI21X1 g121574(.A0 (n_14373), .A1 (n_13976), .B0 (n_22759), .Y(n_13977));
INVX1 g121603(.A (n_13974), .Y (n_13973));
INVX2 g121620(.A (n_14233), .Y (n_13970));
AOI21X1 g121625(.A0 (n_14349), .A1 (n_13967), .B0 (n_9548), .Y(n_13968));
XOR2X1 g121641(.A (n_18159), .B (n_13376), .Y (n_13966));
NAND2X1 g121699(.A (n_29695), .B (n_13963), .Y (n_13965));
NAND2X1 g121703(.A (n_29505), .B (n_13963), .Y (n_13964));
NAND2X1 g121718(.A (n_10917), .B (n_13963), .Y (n_13962));
NAND2X1 g121723(.A (n_14351), .B (n_13960), .Y (n_13961));
NAND2X1 g121724(.A (n_13963), .B (n_29523), .Y (n_13959));
NAND2X1 g121742(.A (n_13954), .B (n_13957), .Y (n_13958));
OR2X1 g121751(.A (n_14344), .B (n_35766), .Y (n_13956));
NAND2X1 g121753(.A (n_13954), .B (n_35744), .Y (n_13955));
NAND2X1 g121764(.A (n_13952), .B (n_13960), .Y (n_13953));
NAND2X1 g121765(.A (n_29505), .B (n_13960), .Y (n_13951));
NAND2X1 g121766(.A (n_29695), .B (n_13960), .Y (n_13950));
NAND2X1 g121768(.A (n_8284), .B (n_13963), .Y (n_13949));
OAI21X1 g121785(.A0 (n_35944), .A1 (n_13316), .B0 (n_24505), .Y(n_13948));
OAI21X1 g121794(.A0 (n_13759), .A1 (n_13317), .B0 (n_25682), .Y(n_13946));
OAI21X1 g121811(.A0 (n_14178), .A1 (n_13317), .B0 (n_21942), .Y(n_13945));
AND2X1 g121820(.A (n_13516), .B (n_25049), .Y (n_13944));
NOR2X1 g121918(.A (n_14331), .B (n_13147), .Y (n_13943));
INVX1 g121937(.A (n_21168), .Y (n_13942));
INVX1 g121941(.A (n_27225), .Y (n_13941));
INVX1 g121943(.A (n_26785), .Y (n_13940));
NAND2X1 g121946(.A (n_13154), .B (n_18262), .Y (n_13939));
NAND2X1 g121959(.A (n_17665), .B (P3_reg1[11] ), .Y (n_24760));
NAND2X1 g121960(.A (n_14267), .B (n_13366), .Y (n_14727));
INVX1 g121961(.A (n_33287), .Y (n_13938));
NAND2X1 g121968(.A (n_23034), .B (n_13515), .Y (n_15031));
INVX1 g121980(.A (n_25035), .Y (n_13937));
INVX1 g121999(.A (n_22813), .Y (n_13936));
OR2X1 g122002(.A (n_13072), .B (n_35719), .Y (n_13935));
NAND2X1 g122005(.A (n_14267), .B (n_13511), .Y (n_15020));
INVX1 g122014(.A (n_24090), .Y (n_13933));
NAND2X1 g122031(.A (n_13156), .B (n_13957), .Y (n_13932));
INVX1 g122040(.A (n_13720), .Y (n_13931));
NAND2X1 g122047(.A (n_13918), .B (n_13957), .Y (n_13930));
INVX1 g122058(.A (n_21666), .Y (n_13929));
INVX1 g122068(.A (n_21617), .Y (n_13928));
NAND2X1 g122076(.A (n_13913), .B (n_13957), .Y (n_13927));
NAND2X1 g122136(.A (n_13925), .B (n_2718), .Y (n_19389));
NAND2X1 g122138(.A (n_13901), .B (n_13721), .Y (n_24711));
NAND2X1 g122141(.A (n_17665), .B (n_13680), .Y (n_25387));
NAND2X1 g122147(.A (n_13925), .B (P3_reg1[18] ), .Y (n_26371));
NAND2X1 g122150(.A (n_13925), .B (n_13724), .Y (n_26776));
OR2X1 g122152(.A (n_12515), .B (n_35834), .Y (n_13924));
INVX1 g122153(.A (n_18939), .Y (n_13923));
INVX1 g122156(.A (n_27762), .Y (n_13922));
INVX1 g122164(.A (n_18936), .Y (n_13921));
INVX1 g122167(.A (n_20755), .Y (n_13920));
NAND2X1 g122175(.A (n_23034), .B (P3_reg2[15] ), .Y (n_14748));
NAND2X1 g122179(.A (n_13616), .B (n_13689), .Y (n_29694));
NAND2X1 g122184(.A (n_13918), .B (n_35744), .Y (n_13919));
INVX1 g122185(.A (n_13917), .Y (n_14353));
INVX1 g122188(.A (n_13686), .Y (n_13915));
NAND2X1 g122192(.A (n_17665), .B (n_13732), .Y (n_14150));
NAND2X1 g122201(.A (n_17665), .B (P3_reg1[9] ), .Y (n_24751));
NAND2X1 g122205(.A (n_13913), .B (n_35744), .Y (n_13914));
NAND2X1 g122211(.A (n_17665), .B (P3_reg1[17] ), .Y (n_26777));
INVX1 g122221(.A (n_13911), .Y (n_13912));
NAND2X1 g122231(.A (n_14267), .B (n_13338), .Y (n_14672));
NAND2X1 g122232(.A (n_12923), .B (n_13957), .Y (n_13909));
NAND2X1 g122236(.A (n_14267), .B (n_13332), .Y (n_14565));
NAND2X1 g122237(.A (n_14267), .B (n_13358), .Y (n_14626));
NAND2X1 g122243(.A (n_13716), .B (n_35816), .Y (n_13908));
NAND2X1 g122248(.A (n_12572), .B (n_13957), .Y (n_13907));
INVX1 g122251(.A (n_13905), .Y (n_13904));
INVX1 g122256(.A (n_13902), .Y (n_13903));
NAND2X1 g122259(.A (n_13901), .B (P3_reg1[1] ), .Y (n_21874));
INVX1 g122262(.A (n_24086), .Y (n_13900));
INVX1 g122264(.A (n_24709), .Y (n_13899));
INVX1 g122266(.A (n_24088), .Y (n_13898));
INVX1 g122273(.A (n_23130), .Y (n_13897));
OAI21X1 g122325(.A0 (n_13895), .A1 (n_14261), .B0 (n_23648), .Y(n_13896));
OAI21X1 g122338(.A0 (n_14147), .A1 (n_13316), .B0 (n_19325), .Y(n_13894));
INVX1 g122350(.A (n_13669), .Y (n_14366));
INVX1 g122382(.A (n_13667), .Y (n_14143));
NAND2X1 g122385(.A (n_13892), .B (n_9135), .Y (n_27064));
NAND2X1 g122395(.A (n_13813), .B (P2_reg_108), .Y (n_27389));
NAND2X1 g122402(.A (n_32711), .B (n_13893), .Y (n_14141));
NAND2X1 g122406(.A (n_13892), .B (n_9178), .Y (n_26925));
NAND2X1 g122430(.A (n_13892), .B (n_9599), .Y (n_21604));
NAND2X1 g122431(.A (n_13571), .B (n_10363), .Y (n_22016));
NAND2X1 g122433(.A (n_13850), .B (n_9634), .Y (n_21548));
NAND2X1 g122442(.A (n_13892), .B (n_9595), .Y (n_23042));
INVX1 g122443(.A (n_25704), .Y (n_13891));
INVX1 g122454(.A (n_25335), .Y (n_13890));
INVX1 g122460(.A (n_13888), .Y (n_22441));
INVX1 g122471(.A (n_13885), .Y (n_23542));
INVX1 g122486(.A (n_27717), .Y (n_13883));
INVX1 g122492(.A (n_13650), .Y (n_14129));
INVX1 g122494(.A (n_13881), .Y (n_24675));
INVX1 g122504(.A (n_27221), .Y (n_13880));
INVX1 g122509(.A (n_13648), .Y (n_14125));
INVX1 g122514(.A (n_13878), .Y (n_25151));
NAND2X1 g122524(.A (n_13873), .B (n_10886), .Y (n_28063));
INVX1 g122530(.A (n_13646), .Y (n_14121));
INVX1 g122532(.A (n_28325), .Y (n_13877));
INVX1 g122537(.A (n_26985), .Y (n_14118));
INVX1 g122545(.A (n_13875), .Y (n_23242));
NAND2X1 g122549(.A (n_32770), .B (n_10563), .Y (n_18815));
NAND2X1 g122552(.A (n_13873), .B (P1_reg2[30] ), .Y (n_20173));
INVX1 g122557(.A (n_14172), .Y (n_14319));
INVX1 g122563(.A (n_13639), .Y (n_14112));
INVX1 g122573(.A (n_13638), .Y (n_14109));
OR2X1 g122578(.A (n_13895), .B (n_19330), .Y (n_13871));
NAND2X1 g122579(.A (n_32648), .B (n_4475), .Y (n_26202));
NAND2X1 g122580(.A (n_32709), .B (P2_reg2[18] ), .Y (n_26200));
NAND2X1 g122590(.A (n_32720), .B (n_10047), .Y (n_27220));
NAND2X1 g122598(.A (n_32711), .B (n_10082), .Y (n_27380));
NAND2X1 g122604(.A (n_32767), .B (n_10604), .Y (n_26923));
NAND2X1 g122620(.A (n_32767), .B (n_3565), .Y (n_22013));
NAND2X1 g122622(.A (n_32719), .B (n_3709), .Y (n_23039));
NAND2X1 g122626(.A (n_32767), .B (P2_reg2[8] ), .Y (n_23380));
NAND2X1 g122628(.A (n_13850), .B (n_10562), .Y (n_18814));
NAND2X1 g122636(.A (n_13581), .B (P2_reg3[1] ), .Y (n_20019));
INVX1 g122637(.A (n_28324), .Y (n_13868));
AND2X1 g122643(.A (n_13862), .B (P2_reg_95), .Y (n_14090));
NAND2X1 g122647(.A (n_1183), .B (n_13854), .Y (n_14089));
INVX1 g122667(.A (n_19492), .Y (n_14084));
INVX1 g122687(.A (n_13628), .Y (n_14080));
INVX1 g122692(.A (n_13864), .Y (n_24121));
INVX1 g122708(.A (n_29014), .Y (n_13863));
NAND2X1 g122715(.A (n_13862), .B (n_9101), .Y (n_24890));
INVX1 g122729(.A (n_13622), .Y (n_14074));
NAND2X1 g122740(.A (n_10032), .B (n_13852), .Y (n_26569));
NAND2X1 g122747(.A (n_8185), .B (n_13581), .Y (n_25344));
INVX2 g122759(.A (n_18533), .Y (n_14635));
INVX2 g122791(.A (n_26234), .Y (n_14749));
INVX2 g122799(.A (n_22021), .Y (n_14627));
INVX2 g122806(.A (n_25072), .Y (n_14384));
NAND2X1 g122903(.A (n_8467), .B (n_13854), .Y (n_24892));
NAND2X1 g122910(.A (n_8164), .B (n_13854), .Y (n_26197));
NAND2X1 g122915(.A (n_10612), .B (n_13854), .Y (n_27068));
NAND2X1 g122925(.A (n_10041), .B (n_13852), .Y (n_26376));
NAND2X1 g122927(.A (n_10081), .B (n_13850), .Y (n_27377));
NAND2X1 g122934(.A (n_9345), .B (n_13852), .Y (n_26929));
NAND2X2 g122938(.A (n_10601), .B (n_13852), .Y (n_28572));
NAND2X2 g122940(.A (n_8447), .B (n_13852), .Y (n_28570));
NAND2X1 g122941(.A (n_13850), .B (n_7475), .Y (n_21609));
NAND2X1 g122949(.A (n_13581), .B (n_1911), .Y (n_23046));
NAND2X1 g122968(.A (n_9512), .B (n_13850), .Y (n_27399));
NAND2X1 g123096(.A (n_13581), .B (n_2784), .Y (n_24012));
NAND2X1 g123100(.A (n_8190), .B (n_13852), .Y (n_14049));
INVX2 g123251(.A (n_13843), .Y (n_20050));
INVX1 g123254(.A (n_13842), .Y (n_23007));
INVX1 g123259(.A (n_14116), .Y (n_22064));
INVX1 g123263(.A (n_13840), .Y (n_26412));
INVX1 g123265(.A (n_13839), .Y (n_22792));
INVX1 g123266(.A (n_13839), .Y (n_25297));
INVX1 g123267(.A (n_13839), .Y (n_25003));
INVX2 g123278(.A (n_13838), .Y (n_14045));
INVX2 g123285(.A (n_14124), .Y (n_23270));
INVX4 g123289(.A (n_26204), .Y (n_18918));
INVX1 g123412(.A (n_26631), .Y (n_21243));
CLKBUFX1 g123555(.A (n_13823), .Y (n_14036));
INVX2 g123560(.A (n_13826), .Y (n_25402));
INVX1 g123571(.A (n_24984), .Y (n_21169));
INVX2 g123581(.A (n_24893), .Y (n_22786));
INVX4 g123583(.A (n_13823), .Y (n_25290));
CLKBUFX1 g123588(.A (n_13822), .Y (n_17797));
CLKBUFX3 g123590(.A (n_13822), .Y (n_23001));
INVX2 g123597(.A (n_13821), .Y (n_18378));
INVX1 g123598(.A (n_13821), .Y (n_21185));
INVX1 g123599(.A (n_13821), .Y (n_23696));
INVX1 g123632(.A (n_13820), .Y (n_21627));
INVX2 g123637(.A (n_26210), .Y (n_22412));
CLKBUFX1 g123651(.A (n_34499), .Y (n_18340));
INVX1 g123655(.A (n_18399), .Y (n_17288));
INVX1 g123668(.A (n_25374), .Y (n_14032));
INVX4 g123672(.A (n_13817), .Y (n_25309));
NAND2X1 g122505(.A (n_13644), .B (n_11148), .Y (n_27221));
NAND2X1 g122497(.A (n_13637), .B (n_10893), .Y (n_27716));
NAND2X1 g122455(.A (n_13668), .B (n_9071), .Y (n_25335));
INVX1 g123264(.A (n_13602), .Y (n_13840));
INVX1 g123669(.A (n_13862), .Y (n_25374));
NAND2X1 g120765(.A (n_13413), .B (n_13418), .Y (n_35698));
INVX2 g123561(.A (n_13582), .Y (n_13826));
NAND2X1 g121120(.A (n_13552), .B (n_17968), .Y (n_13811));
MX2X1 g121219(.A (n_11500), .B (n_13114), .S0 (n_34615), .Y(n_13810));
INVX1 g121221(.A (n_14274), .Y (n_13809));
NAND2X1 g121226(.A (n_11277), .B (n_13417), .Y (n_14270));
NAND2X1 g121232(.A (n_35442), .B (n_35443), .Y (n_14971));
XOR2X1 g121236(.A (n_9883), .B (n_13245), .Y (n_13807));
NAND2X1 g121249(.A (n_14010), .B (n_14235), .Y (n_13806));
NAND2X1 g121252(.A (n_14010), .B (n_13274), .Y (n_13805));
NAND2X1 g121258(.A (n_14226), .B (n_14439), .Y (n_13804));
NAND2X1 g121282(.A (n_13533), .B (n_14439), .Y (n_13803));
OAI21X1 g121291(.A0 (n_14219), .A1 (n_24312), .B0 (n_24009), .Y(n_13802));
AND2X1 g121324(.A (n_13406), .B (n_24721), .Y (n_13801));
XOR2X1 g121418(.A (n_10771), .B (n_13231), .Y (n_13800));
NAND2X1 g121419(.A (n_11751), .B (n_13404), .Y (n_14918));
INVX1 g121420(.A (n_13798), .Y (n_13799));
NAND2X1 g121424(.A (n_11053), .B (n_13402), .Y (n_14466));
INVX1 g121427(.A (n_14018), .Y (n_13796));
NAND2X1 g121438(.A (n_11515), .B (n_13401), .Y (n_13996));
NAND2X1 g121439(.A (n_12299), .B (n_13403), .Y (n_15059));
OAI21X1 g121446(.A0 (n_7832), .A1 (n_13223), .B0 (n_11265), .Y(n_13994));
XOR2X1 g121456(.A (n_9482), .B (n_13233), .Y (n_13791));
OR2X1 g121471(.A (n_13992), .B (n_13788), .Y (n_13790));
OR2X1 g121472(.A (n_14001), .B (n_13788), .Y (n_13789));
NAND2X1 g121476(.A (n_13988), .B (n_13274), .Y (n_13787));
NOR2X1 g121500(.A (n_14385), .B (n_13163), .Y (n_13786));
NAND2X1 g121590(.A (n_11261), .B (n_13394), .Y (n_14425));
INVX1 g121591(.A (n_14242), .Y (n_13785));
INVX1 g121604(.A (n_13784), .Y (n_13974));
INVX1 g121617(.A (n_13529), .Y (n_14236));
INVX2 g121622(.A (n_13528), .Y (n_14233));
OR2X1 g121685(.A (n_13782), .B (n_13781), .Y (n_13783));
OR2X1 g121694(.A (n_13782), .B (n_13788), .Y (n_13780));
OR2X1 g121695(.A (n_13782), .B (n_14218), .Y (n_13779));
NOR2X1 g121711(.A (n_14344), .B (n_13163), .Y (n_13778));
NAND2X1 g121712(.A (n_14351), .B (n_13775), .Y (n_13777));
NAND2X1 g121720(.A (n_13775), .B (n_26548), .Y (n_13776));
NAND2X1 g121722(.A (n_29341), .B (n_13775), .Y (n_13774));
NAND2X1 g121726(.A (n_13967), .B (n_26548), .Y (n_13773));
NAND2X1 g121727(.A (n_8284), .B (n_13775), .Y (n_13771));
NAND2X1 g121734(.A (n_29695), .B (n_13967), .Y (n_13770));
NAND2X1 g121735(.A (n_14351), .B (n_13967), .Y (n_13769));
AND2X1 g121737(.A (n_14349), .B (n_13775), .Y (n_13768));
NAND2X1 g121774(.A (n_13766), .B (n_14439), .Y (n_13767));
NAND2X1 g122661(.A (n_13653), .B (n_10175), .Y (n_27709));
NAND2X1 g121885(.A (n_13736), .B (n_2721), .Y (n_14642));
INVX1 g121892(.A (n_13764), .Y (n_13765));
OR2X1 g121901(.A (n_13761), .B (n_34417), .Y (n_13763));
OR2X1 g121902(.A (n_13761), .B (n_18303), .Y (n_13762));
OR2X1 g121905(.A (n_13759), .B (n_13758), .Y (n_13760));
NAND2X1 g122648(.A (n_13437), .B (n_10150), .Y (n_24003));
OR2X1 g121920(.A (n_13759), .B (n_13434), .Y (n_13757));
OR2X1 g121921(.A (n_14178), .B (n_13788), .Y (n_13755));
NAND2X1 g121929(.A (n_35600), .B (n_13381), .Y (n_26398));
NAND2X1 g121930(.A (n_35485), .B (n_13389), .Y (n_26869));
NAND2X1 g121931(.A (n_35466), .B (n_7734), .Y (n_22758));
NAND2X1 g121932(.A (n_35600), .B (n_13383), .Y (n_28543));
NAND2X1 g121933(.A (n_35600), .B (n_13387), .Y (n_29545));
NAND2X1 g121934(.A (n_35485), .B (n_13380), .Y (n_27525));
NAND2X1 g121935(.A (n_35583), .B (n_3187), .Y (n_27711));
NAND2X1 g121938(.A (n_35600), .B (n_2721), .Y (n_21168));
NAND2X1 g121939(.A (n_35485), .B (n_13386), .Y (n_28322));
NAND2X1 g121940(.A (n_35583), .B (n_13385), .Y (n_27707));
NAND2X1 g121942(.A (n_35583), .B (n_3887), .Y (n_27225));
NAND2X1 g121944(.A (n_35485), .B (n_3072), .Y (n_26785));
NOR2X1 g121949(.A (n_13748), .B (n_34417), .Y (n_13749));
OR2X1 g121950(.A (n_14162), .B (n_34417), .Y (n_13747));
NOR2X1 g121951(.A (n_34417), .B (n_8945), .Y (n_13746));
NOR2X1 g121953(.A (n_14159), .B (n_34417), .Y (n_13745));
NOR2X1 g121954(.A (n_13748), .B (n_18303), .Y (n_13744));
OR2X1 g121955(.A (n_9172), .B (n_18303), .Y (n_13743));
NOR2X1 g121956(.A (n_18303), .B (n_8945), .Y (n_13742));
NOR2X1 g121957(.A (n_33505), .B (n_18303), .Y (n_13741));
NAND2X1 g121958(.A (n_35719), .B (P3_reg1[11] ), .Y (n_14723));
NAND2X1 g121963(.A (n_13739), .B (P3_reg2[18] ), .Y (n_14634));
NAND2X1 g121971(.A (n_13737), .B (n_13507), .Y (n_14716));
INVX1 g121975(.A (n_24060), .Y (n_13738));
NAND2X1 g121977(.A (n_35766), .B (n_13695), .Y (n_14610));
NAND2X1 g121981(.A (n_35600), .B (n_13327), .Y (n_25035));
NAND2X1 g121983(.A (n_13737), .B (P3_reg2[6] ), .Y (n_14612));
NAND2X1 g121986(.A (n_13696), .B (P3_reg1[3] ), .Y (n_22027));
NAND2X1 g121988(.A (n_13739), .B (P3_reg2[9] ), .Y (n_14561));
NAND2X1 g121992(.A (n_13737), .B (n_13329), .Y (n_14266));
NAND2X1 g121993(.A (n_13736), .B (n_13735), .Y (n_14624));
NAND3X1 g121994(.A (n_35719), .B (n_13732), .C (n_8316), .Y(n_13734));
NAND2X1 g122000(.A (n_35485), .B (n_13711), .Y (n_22813));
NAND3X1 g122001(.A (n_35813), .B (n_13727), .C (n_8316), .Y(n_13728));
NAND2X1 g122015(.A (n_35600), .B (n_13370), .Y (n_24090));
NAND2X1 g122016(.A (n_35600), .B (n_7755), .Y (n_24002));
NAND2X1 g122020(.A (n_35830), .B (n_13724), .Y (n_14721));
INVX1 g122026(.A (n_22776), .Y (n_13723));
NAND2X1 g122029(.A (n_35719), .B (n_13721), .Y (n_14414));
NAND2X1 g122033(.A (n_13737), .B (P3_reg1[6] ), .Y (n_23935));
NAND2X1 g122036(.A (n_35600), .B (n_13375), .Y (n_25793));
NAND3X1 g122041(.A (n_35768), .B (n_15147), .C (n_13732), .Y(n_13720));
NAND2X1 g122043(.A (n_35834), .B (P3_reg1[1] ), .Y (n_14358));
NAND2X1 g122044(.A (n_13737), .B (n_13361), .Y (n_14667));
NAND2X1 g122045(.A (n_35840), .B (n_13698), .Y (n_14719));
NAND2X1 g122046(.A (n_35600), .B (n_13379), .Y (n_28058));
NAND2X1 g122050(.A (n_13716), .B (n_14439), .Y (n_13717));
NAND2X1 g122051(.A (n_35830), .B (n_13681), .Y (n_14410));
NAND2X1 g122056(.A (n_13736), .B (n_10578), .Y (n_14603));
NAND2X1 g122059(.A (n_13696), .B (n_13692), .Y (n_21666));
INVX1 g122064(.A (n_25837), .Y (n_13714));
NAND2X1 g122069(.A (n_35485), .B (P3_reg3[2] ), .Y (n_21617));
NAND2X1 g122070(.A (n_13696), .B (P3_reg1[16] ), .Y (n_25839));
NAND2X1 g122071(.A (n_13737), .B (n_13343), .Y (n_14936));
NAND2X1 g122077(.A (n_13739), .B (n_13502), .Y (n_14583));
NAND2X1 g122078(.A (n_13696), .B (P3_reg1[4] ), .Y (n_22779));
NAND2X1 g122080(.A (n_13696), .B (n_13344), .Y (n_14608));
NAND2X1 g122091(.A (n_13701), .B (n_13699), .Y (n_27685));
NAND2X1 g122111(.A (n_12049), .B (n_14439), .Y (n_13712));
NAND2X1 g122115(.A (n_35583), .B (n_13378), .Y (n_25148));
NAND2X1 g122131(.A (n_13736), .B (n_13711), .Y (n_14706));
NAND2X1 g122139(.A (n_13739), .B (n_13709), .Y (n_25925));
NAND2X1 g122140(.A (n_35824), .B (n_13709), .Y (n_14714));
NAND2X1 g122142(.A (n_13737), .B (n_13679), .Y (n_25327));
NAND2X1 g122144(.A (n_35766), .B (P3_reg1[16] ), .Y (n_15087));
NAND2X1 g122145(.A (n_35834), .B (P3_reg1[17] ), .Y (n_14360));
NAND2X1 g122148(.A (n_35775), .B (P3_reg1[18] ), .Y (n_14632));
NAND2X1 g122154(.A (n_13696), .B (n_13687), .Y (n_18939));
NAND2X1 g122155(.A (n_35834), .B (n_13678), .Y (n_14978));
NAND2X1 g122157(.A (n_13701), .B (n_13673), .Y (n_27762));
NAND2X1 g122161(.A (n_35766), .B (n_13697), .Y (n_14680));
NAND2X1 g122163(.A (n_35766), .B (n_13699), .Y (n_14745));
NAND2X1 g122165(.A (n_13696), .B (n_13698), .Y (n_18936));
NAND2X1 g122166(.A (n_13701), .B (n_13697), .Y (n_27205));
NAND2X1 g122168(.A (n_13696), .B (n_13695), .Y (n_20755));
NAND2X1 g122169(.A (n_35583), .B (P3_reg3[0] ), .Y (n_19410));
NAND2X1 g122171(.A (n_35775), .B (P3_reg1[26] ), .Y (n_14939));
NAND2X1 g122172(.A (n_13696), .B (P3_reg2[28] ), .Y (n_15409));
NAND2X1 g122173(.A (n_35768), .B (n_13692), .Y (n_15299));
NAND2X1 g122176(.A (n_13737), .B (n_13690), .Y (n_29480));
NAND2X1 g122177(.A (n_35719), .B (n_13690), .Y (n_15347));
NAND2X1 g122180(.A (n_35766), .B (n_13689), .Y (n_14678));
NAND2X1 g122181(.A (n_35834), .B (P3_reg1[9] ), .Y (n_14572));
NAND2X1 g122182(.A (n_35775), .B (n_13687), .Y (n_14665));
NAND2X1 g122183(.A (n_13737), .B (n_13677), .Y (n_21601));
NAND2X1 g122187(.A (n_13701), .B (n_13727), .Y (n_13917));
NAND3X1 g122189(.A (n_35768), .B (n_13727), .C (n_15110), .Y(n_13686));
NAND2X1 g122193(.A (n_35824), .B (P3_reg1[3] ), .Y (n_14412));
NAND2X1 g122194(.A (n_35766), .B (P3_reg1[4] ), .Y (n_14382));
NAND2X1 g122196(.A (n_13696), .B (n_13683), .Y (n_23666));
NAND2X1 g122197(.A (n_35834), .B (n_13683), .Y (n_14347));
NAND2X1 g122198(.A (n_35766), .B (P3_reg1[6] ), .Y (n_14387));
NAND2X1 g122199(.A (n_13737), .B (P3_reg1[7] ), .Y (n_23401));
NAND2X1 g122200(.A (n_13696), .B (n_13681), .Y (n_24042));
NAND2X1 g122204(.A (n_35766), .B (n_13680), .Y (n_14362));
NAND2X1 g122210(.A (n_13739), .B (n_13342), .Y (n_14674));
NAND2X1 g122215(.A (n_35719), .B (n_13679), .Y (n_14685));
NAND2X1 g122217(.A (n_13739), .B (n_13678), .Y (n_26493));
NAND2X1 g122218(.A (n_13696), .B (n_13336), .Y (n_14670));
NAND2X1 g122219(.A (n_13696), .B (n_13368), .Y (n_14194));
NAND2X1 g122222(.A (n_13737), .B (n_13335), .Y (n_13911));
NAND2X1 g122225(.A (n_13696), .B (n_13334), .Y (n_14725));
NAND2X1 g122228(.A (n_35834), .B (n_13677), .Y (n_14356));
NAND2X1 g122229(.A (n_35485), .B (n_13675), .Y (n_21545));
NAND2X1 g122230(.A (n_13701), .B (n_13201), .Y (n_15297));
NAND2X1 g122249(.A (n_35824), .B (P3_reg1[7] ), .Y (n_14676));
NOR2X1 g122252(.A (n_13554), .B (n_290), .Y (n_13905));
NAND2X1 g122253(.A (n_35830), .B (n_13673), .Y (n_14577));
NAND2X1 g122257(.A (n_13737), .B (n_13352), .Y (n_13902));
NAND2X1 g122258(.A (n_13736), .B (P3_reg3[2] ), .Y (n_14597));
NAND2X1 g122263(.A (n_35600), .B (n_10097), .Y (n_24086));
NAND2X1 g122265(.A (n_35600), .B (n_10582), .Y (n_24709));
NAND2X1 g122267(.A (n_35583), .B (n_10100), .Y (n_24088));
NAND2X1 g122274(.A (n_35600), .B (n_34587), .Y (n_23130));
NAND2X1 g122275(.A (n_35600), .B (n_8055), .Y (n_25842));
OAI21X1 g122284(.A0 (n_14086), .A1 (n_14702), .B0 (n_21889), .Y(n_13670));
NOR2X1 g122351(.A (n_11727), .B (n_13297), .Y (n_13669));
NAND2X1 g122370(.A (n_13665), .B (n_9165), .Y (n_26209));
NAND2X1 g122373(.A (n_13665), .B (n_9139), .Y (n_26208));
NAND2X1 g122378(.A (n_13668), .B (n_10452), .Y (n_20022));
NAND2X1 g122383(.A (n_13661), .B (P2_reg_104), .Y (n_13667));
OR2X1 g122398(.A (n_13895), .B (n_13663), .Y (n_13664));
NAND2X1 g122403(.A (n_13665), .B (n_9794), .Y (n_27388));
NAND2X1 g122416(.A (n_13661), .B (n_9602), .Y (n_13662));
OR2X1 g122417(.A (n_14078), .B (n_13663), .Y (n_13660));
NAND2X1 g122418(.A (n_25054), .B (n_11136), .Y (n_19329));
NAND2X1 g122419(.A (n_13661), .B (n_9088), .Y (n_29133));
NAND2X1 g122420(.A (n_13657), .B (n_4151), .Y (n_25055));
NAND2X1 g122421(.A (n_13668), .B (n_10435), .Y (n_21551));
NAND2X1 g122424(.A (n_13657), .B (n_4590), .Y (n_25706));
NAND2X1 g122427(.A (n_13659), .B (n_4445), .Y (n_25353));
NAND2X1 g122432(.A (n_13651), .B (n_4213), .Y (n_25053));
NAND2X1 g122434(.A (n_13661), .B (n_10443), .Y (n_23043));
NAND2X1 g122439(.A (n_13659), .B (P1_reg2[14] ), .Y (n_25705));
NAND2X1 g122444(.A (n_13448), .B (n_4824), .Y (n_25704));
NAND2X1 g122448(.A (n_13665), .B (n_9121), .Y (n_24007));
NAND2X1 g122449(.A (n_13657), .B (P1_reg2[16] ), .Y (n_25852));
INVX1 g122457(.A (n_13655), .Y (n_24508));
AND2X1 g122462(.A (n_13654), .B (P2_reg1[10] ), .Y (n_13888));
NAND2X1 g122464(.A (n_13652), .B (P2_reg1[11] ), .Y (n_22839));
NAND2X1 g122467(.A (n_13659), .B (n_4277), .Y (n_27718));
AND2X1 g122473(.A (n_13654), .B (P2_reg1[13] ), .Y (n_13885));
NAND2X1 g122474(.A (n_13653), .B (n_10128), .Y (n_28202));
NAND2X1 g122476(.A (n_13652), .B (n_9586), .Y (n_23136));
NAND2X1 g122477(.A (n_13657), .B (P1_reg2[19] ), .Y (n_28215));
NAND2X1 g122480(.A (n_13627), .B (P1_reg2[1] ), .Y (n_21890));
NAND2X1 g122483(.A (n_13652), .B (P2_reg1[17] ), .Y (n_26207));
NAND2X1 g122484(.A (n_13651), .B (n_11120), .Y (n_28213));
NAND2X1 g122485(.A (n_13652), .B (P2_reg1[19] ), .Y (n_26203));
NAND2X1 g122487(.A (n_13657), .B (n_10897), .Y (n_27717));
NAND2X1 g122488(.A (n_13647), .B (P2_reg1[1] ), .Y (n_20021));
NAND2X1 g122493(.A (n_13652), .B (P2_reg1[20] ), .Y (n_13650));
AND2X1 g122496(.A (n_13652), .B (P2_reg1[21] ), .Y (n_13881));
NAND2X1 g122498(.A (n_13652), .B (P2_reg1[22] ), .Y (n_27222));
NAND2X1 g122510(.A (n_13564), .B (n_9097), .Y (n_13648));
AND2X1 g122515(.A (n_13641), .B (P2_reg1[27] ), .Y (n_13878));
NAND2X1 g122516(.A (n_13444), .B (n_10890), .Y (n_28555));
NAND2X1 g122521(.A (n_13647), .B (n_9092), .Y (n_29132));
NAND2X1 g122525(.A (n_13647), .B (P2_reg1[2] ), .Y (n_21550));
NAND2X1 g122531(.A (n_13647), .B (n_13645), .Y (n_13646));
NAND2X2 g122533(.A (n_13644), .B (n_11327), .Y (n_28325));
NAND2X1 g122534(.A (n_13647), .B (P2_reg1[4] ), .Y (n_22015));
NAND2X1 g122538(.A (n_13651), .B (n_11144), .Y (n_26985));
NAND2X1 g122539(.A (n_13652), .B (P2_reg1[5] ), .Y (n_23041));
AND2X1 g122547(.A (n_13641), .B (P2_reg1[9] ), .Y (n_13875));
NAND2X2 g122558(.A (n_13659), .B (n_13640), .Y (n_14172));
NAND2X1 g122564(.A (n_32711), .B (P2_reg2[12] ), .Y (n_13639));
NAND2X1 g122565(.A (n_13633), .B (n_10134), .Y (n_28061));
NAND2X1 g122566(.A (n_13637), .B (n_3470), .Y (n_22953));
NAND2X1 g122569(.A (n_13644), .B (n_3668), .Y (n_22844));
NAND2X1 g122574(.A (n_32648), .B (P2_reg2[15] ), .Y (n_13638));
NAND2X1 g122577(.A (n_13657), .B (n_3693), .Y (n_23641));
NAND2X1 g122581(.A (n_13651), .B (n_3416), .Y (n_23640));
NAND2X1 g122588(.A (n_13637), .B (n_4561), .Y (n_24839));
NAND2X1 g122591(.A (n_13657), .B (n_4230), .Y (n_24006));
NAND2X1 g122605(.A (n_13634), .B (n_10187), .Y (n_19328));
NAND2X1 g122609(.A (n_32707), .B (P2_reg2[29] ), .Y (n_26570));
NAND2X1 g122621(.A (n_13653), .B (n_10205), .Y (n_25345));
NAND2X1 g122629(.A (n_13665), .B (n_9067), .Y (n_24305));
NAND2X1 g122630(.A (n_13629), .B (n_13635), .Y (n_21293));
NAND2X1 g122631(.A (n_13653), .B (n_10201), .Y (n_25689));
NAND2X1 g122638(.A (n_13624), .B (n_10219), .Y (n_28324));
NAND2X1 g122639(.A (n_13634), .B (n_10156), .Y (n_25342));
NAND2X1 g122650(.A (n_13633), .B (n_10191), .Y (n_25048));
NAND2X1 g122656(.A (n_13634), .B (n_10189), .Y (n_25684));
OR2X1 g122657(.A (n_14078), .B (n_14261), .Y (n_13632));
NAND2X1 g122658(.A (n_13653), .B (n_10182), .Y (n_25683));
NAND2X1 g122659(.A (n_13637), .B (n_3259), .Y (n_21941));
NAND2X1 g122660(.A (n_13653), .B (n_10180), .Y (n_25850));
NAND2X1 g122668(.A (n_13434), .B (n_10171), .Y (n_19492));
NAND2X1 g122669(.A (n_13633), .B (n_10165), .Y (n_27708));
NAND2X1 g122673(.A (n_13634), .B (P1_reg_173), .Y (n_27217));
INVX1 g122677(.A (n_13487), .Y (n_13866));
NAND2X1 g122679(.A (n_13432), .B (n_10225), .Y (n_28548));
NAND2X1 g122680(.A (n_13624), .B (n_10211), .Y (n_29666));
NAND2X1 g122683(.A (n_13629), .B (P1_reg_180), .Y (n_22097));
NAND2X1 g122684(.A (n_13665), .B (n_9103), .Y (n_24888));
NAND2X1 g122688(.A (n_13627), .B (n_10858), .Y (n_13628));
NAND2X1 g122689(.A (n_13629), .B (n_10197), .Y (n_22952));
NAND2X1 g122690(.A (n_13653), .B (n_10178), .Y (n_26787));
AND2X1 g122693(.A (n_13654), .B (P2_reg1[18] ), .Y (n_13864));
NAND2X1 g122694(.A (n_13653), .B (n_10144), .Y (n_22842));
NAND2X1 g122695(.A (n_13624), .B (n_10221), .Y (n_23638));
NAND2X1 g122696(.A (n_13627), .B (P1_reg2[9] ), .Y (n_25051));
NAND2X1 g122697(.A (n_13629), .B (n_10140), .Y (n_23637));
NAND2X1 g122699(.A (n_13629), .B (n_10138), .Y (n_24837));
NAND2X1 g122701(.A (n_13435), .B (n_10154), .Y (n_25047));
NAND2X1 g122709(.A (n_13624), .B (n_10152), .Y (n_29014));
NAND2X1 g122730(.A (n_13647), .B (P2_reg1[31] ), .Y (n_13622));
NAND2X1 g122736(.A (n_13665), .B (n_9475), .Y (n_26193));
OR2X1 g122738(.A (n_14086), .B (n_13663), .Y (n_13620));
INVX8 g122765(.A (n_17665), .Y (n_18533));
INVX1 g122792(.A (n_13616), .Y (n_26234));
INVX4 g122800(.A (n_13901), .Y (n_22021));
INVX1 g122803(.A (n_13925), .Y (n_20133));
INVX1 g122805(.A (n_13616), .Y (n_25599));
INVX1 g122807(.A (n_13616), .Y (n_25072));
NAND2X1 g122895(.A (n_10617), .B (n_13613), .Y (n_24324));
NAND2X1 g122899(.A (n_2909), .B (n_13613), .Y (n_24894));
NAND2X1 g122907(.A (n_8458), .B (n_13613), .Y (n_26216));
INVX1 g123197(.A (n_18498), .Y (n_14101));
INVX1 g123201(.A (n_22032), .Y (n_17293));
INVX1 g123206(.A (n_14339), .Y (n_14404));
INVX1 g123217(.A (n_19330), .Y (n_20178));
INVX1 g123223(.A (n_17713), .Y (n_13845));
INVX2 g123252(.A (n_24249), .Y (n_13843));
INVX1 g123255(.A (n_13604), .Y (n_13842));
BUFX3 g123256(.A (n_13604), .Y (n_24446));
INVX2 g123258(.A (n_13602), .Y (n_14116));
INVX1 g123268(.A (n_13602), .Y (n_13839));
INVX2 g123279(.A (n_13601), .Y (n_13838));
INVX2 g123286(.A (n_13601), .Y (n_14124));
INVX4 g123292(.A (n_13600), .Y (n_26204));
INVX2 g123416(.A (n_18137), .Y (n_14430));
INVX1 g123436(.A (n_19597), .Y (n_19165));
INVX1 g123455(.A (n_23578), .Y (n_13588));
INVX2 g123548(.A (n_13584), .Y (n_26866));
INVX2 g123549(.A (n_13584), .Y (n_27470));
INVX1 g123567(.A (n_24013), .Y (n_18375));
INVX2 g123574(.A (n_13850), .Y (n_24984));
INVX1 g123582(.A (n_13582), .Y (n_24893));
INVX4 g123584(.A (n_13582), .Y (n_13823));
INVX1 g123591(.A (n_13854), .Y (n_13822));
CLKBUFX3 g123600(.A (n_13581), .Y (n_13821));
INVX2 g123603(.A (n_34688), .Y (n_13579));
CLKBUFX3 g123606(.A (n_34688), .Y (n_23791));
INVX1 g123609(.A (n_13581), .Y (n_25404));
INVX1 g123621(.A (n_23725), .Y (n_20054));
INVX2 g123625(.A (n_13574), .Y (n_14134));
INVX2 g123629(.A (n_13573), .Y (n_24889));
CLKBUFX3 g123630(.A (n_13573), .Y (n_27999));
INVX1 g123633(.A (n_13573), .Y (n_13820));
INVX1 g123635(.A (n_13572), .Y (n_14123));
INVX2 g123640(.A (n_13572), .Y (n_26210));
INVX1 g123645(.A (n_13571), .Y (n_24652));
INVX1 g123647(.A (n_34498), .Y (n_22414));
INVX4 g123659(.A (n_13813), .Y (n_18399));
CLKBUFX1 g123674(.A (n_13569), .Y (n_26530));
INVX2 g123682(.A (n_13569), .Y (n_13817));
CLKBUFX1 gbuf_d_475(.A(n_13195), .Y(d_out_475));
CLKBUFX1 gbuf_qn_475(.A(qn_in_475), .Y(addr_484));
CLKBUFX1 gbuf_d_476(.A(n_13193), .Y(d_out_476));
CLKBUFX1 gbuf_qn_476(.A(qn_in_476), .Y(addr_485));
CLKBUFX1 gbuf_d_477(.A(n_13188), .Y(d_out_477));
CLKBUFX1 gbuf_q_477(.A(q_in_477), .Y(n_3314));
CLKBUFX1 gbuf_d_478(.A(n_13198), .Y(d_out_478));
CLKBUFX1 gbuf_qn_478(.A(qn_in_478), .Y(addr_483));
INVX2 g123287(.A (n_13564), .Y (n_13601));
CLKBUFX3 g123683(.A (n_13426), .Y (n_13569));
INVX2 g123269(.A (n_13641), .Y (n_13602));
INVX1 g123257(.A (n_13641), .Y (n_13604));
INVX1 g123646(.A (n_34499), .Y (n_13571));
INVX1 g123644(.A (n_34499), .Y (n_13892));
CLKBUFX1 gbuf_d_479(.A(n_13191), .Y(d_out_479));
CLKBUFX1 gbuf_qn_479(.A(qn_in_479), .Y(addr_3));
INVX1 g123634(.A (n_13427), .Y (n_13573));
CLKBUFX1 g123233(.A (n_26315), .Y (n_22831));
INVX1 g123205(.A (n_13758), .Y (n_17727));
INVX1 g122908(.A (n_28569), .Y (n_22477));
INVX4 g123601(.A (n_34687), .Y (n_13581));
INVX4 g123585(.A (n_13429), .Y (n_13582));
INVX4 g123569(.A (n_13559), .Y (n_13850));
INVX4 g123568(.A (n_13559), .Y (n_24013));
CLKBUFX1 g123550(.A (n_13429), .Y (n_13584));
NAND2X1 g121218(.A (n_11966), .B (n_13251), .Y (n_14733));
OAI21X1 g121223(.A0 (n_13400), .A1 (n_13124), .B0 (n_11490), .Y(n_14274));
XOR2X1 g121234(.A (n_11720), .B (n_13126), .Y (n_13558));
XOR2X1 g121235(.A (n_9198), .B (n_13125), .Y (n_13557));
NAND2X1 g121261(.A (n_13555), .B (n_13238), .Y (n_35883));
INVX1 g121422(.A (n_13553), .Y (n_13798));
INVX1 g121425(.A (n_13552), .Y (n_14268));
NAND2X1 g121429(.A (n_11482), .B (n_13248), .Y (n_14018));
INVX2 g121430(.A (n_13411), .Y (n_14687));
INVX1 g121440(.A (n_14452), .Y (n_13551));
INVX1 g121452(.A (n_13549), .Y (n_13793));
NAND2X1 g121458(.A (n_13235), .B (n_16452), .Y (n_13548));
NAND2X1 g121459(.A (n_13544), .B (n_10799), .Y (n_13546));
OR2X1 g121460(.A (n_13544), .B (n_10799), .Y (n_13545));
NAND2X1 g121474(.A (n_13988), .B (n_14235), .Y (n_13542));
NAND2X1 g121482(.A (n_13540), .B (n_13225), .Y (n_13541));
NAND2X1 g121493(.A (n_8124), .B (n_13220), .Y (n_32250));
NAND2X1 g121502(.A (n_33290), .B (n_13221), .Y (n_13538));
NAND4X1 g121505(.A (n_13236), .B (n_3904), .C (n_3802), .D (n_3390),.Y (n_13537));
INVX8 g123454(.A (n_13434), .Y (n_23578));
NAND2X1 g121586(.A (n_11281), .B (n_13237), .Y (n_14649));
OAI21X1 g121592(.A0 (n_13296), .A1 (n_13087), .B0 (n_11260), .Y(n_14242));
INVX1 g121595(.A (n_14862), .Y (n_13536));
AOI22X1 g121605(.A0 (n_13409), .A1 (n_13086), .B0 (n_9754), .B1(n_13408), .Y (n_13784));
INVX1 g121606(.A (n_14226), .Y (n_13531));
INVX1 g121608(.A (n_14682), .Y (n_13530));
AOI22X1 g121618(.A0 (n_13393), .A1 (n_13084), .B0 (n_11092), .B1(n_13527), .Y (n_13529));
AOI22X1 g121623(.A0 (n_12954), .A1 (n_13082), .B0 (n_17955), .B1(n_13527), .Y (n_13528));
OAI21X1 g121624(.A0 (n_8745), .A1 (n_13090), .B0 (n_11750), .Y(n_14416));
XOR2X1 g121639(.A (n_13098), .B (n_13081), .Y (n_13526));
XOR2X1 g121642(.A (n_10745), .B (n_13096), .Y (n_13525));
NAND4X1 g121701(.A (n_13217), .B (n_3427), .C (n_3803), .D (n_3302),.Y (n_13524));
INVX1 g121837(.A (n_14636), .Y (n_13523));
INVX1 g121887(.A (n_13520), .Y (n_13521));
NOR2X1 g121893(.A (n_24965), .B (n_10114), .Y (n_13764));
INVX1 g121894(.A (n_13518), .Y (n_13519));
NOR2X1 g121898(.A (n_13957), .B (n_2096), .Y (n_14209));
NAND2X1 g121899(.A (n_13214), .B (n_3072), .Y (n_14335));
OR2X1 g121917(.A (n_13759), .B (n_13056), .Y (n_13516));
NOR2X1 g121928(.A (n_18262), .B (n_2975), .Y (n_14221));
NAND2X1 g121976(.A (n_35771), .B (n_13515), .Y (n_24060));
NAND2X1 g122640(.A (n_13179), .B (n_10223), .Y (n_27705));
NAND2X1 g121989(.A (n_13214), .B (n_13675), .Y (n_14605));
INVX1 g121997(.A (n_13372), .Y (n_13963));
NAND2X1 g122018(.A (n_35824), .B (P3_reg2[18] ), .Y (n_27204));
NAND2X1 g122027(.A (n_35771), .B (n_13511), .Y (n_22776));
INVX1 g122052(.A (n_13509), .Y (n_13510));
NAND2X1 g122065(.A (n_35824), .B (n_13507), .Y (n_25837));
NOR2X1 g122095(.A (n_13957), .B (n_3297), .Y (n_14952));
NAND2X1 g122137(.A (n_35824), .B (n_2718), .Y (n_14555));
INVX1 g122159(.A (n_13504), .Y (n_17012));
NAND2X1 g122162(.A (n_35766), .B (n_13502), .Y (n_26775));
NAND2X1 g122203(.A (n_35766), .B (P3_reg2[10] ), .Y (n_24713));
NAND2X1 g122239(.A (n_13214), .B (P3_reg3[0] ), .Y (n_14185));
INVX1 g122254(.A (n_13499), .Y (n_13960));
NAND2X1 g122260(.A (n_35844), .B (n_13498), .Y (n_23718));
INVX1 g122342(.A (n_13766), .Y (n_13497));
INVX1 g122343(.A (n_13766), .Y (n_13496));
INVX1 g122375(.A (n_13494), .Y (n_13493));
INVX1 g122390(.A (n_22954), .Y (n_13492));
INVX1 g122407(.A (n_24840), .Y (n_13491));
INVX1 g122446(.A (n_28195), .Y (n_13490));
AND2X1 g122459(.A (n_13489), .B (n_11141), .Y (n_13655));
NAND2X1 g122542(.A (n_13489), .B (n_10546), .Y (n_29667));
NAND2X1 g122664(.A (n_13488), .B (n_10173), .Y (n_21885));
NAND2X1 g122671(.A (n_13488), .B (P1_reg_172), .Y (n_24299));
NAND2X1 g122678(.A (n_13488), .B (P1_reg_174), .Y (n_13487));
NAND2X1 g122682(.A (n_13488), .B (n_10148), .Y (n_21940));
INVX1 g122718(.A (n_25681), .Y (n_13484));
INVX2 g122748(.A (n_25877), .Y (n_14267));
INVX4 g122763(.A (n_13554), .Y (n_17665));
INVX1 g122771(.A (n_26584), .Y (n_23034));
INVX4 g122783(.A (n_13701), .Y (n_28053));
CLKBUFX2 g122786(.A (n_13478), .Y (n_25596));
INVX2 g122793(.A (n_13478), .Y (n_13616));
INVX4 g122801(.A (n_13478), .Y (n_13901));
INVX1 g122804(.A (n_13478), .Y (n_13925));
OR2X1 g122889(.A (n_14147), .B (n_13183), .Y (n_13470));
INVX1 g122935(.A (n_35057), .Y (n_13466));
INVX1 g122950(.A (n_15119), .Y (n_21262));
INVX1 g122955(.A (n_29034), .Y (n_13461));
INVX1 g123028(.A (n_25690), .Y (n_13458));
INVX1 g123032(.A (n_28204), .Y (n_13457));
INVX2 g123117(.A (n_35945), .Y (n_13454));
INVX1 g123133(.A (n_14325), .Y (n_13452));
INVX1 g123179(.A (n_28734), .Y (n_13873));
INVX8 g123187(.A (n_13657), .Y (n_25554));
INVX2 g123198(.A (n_13644), .Y (n_18498));
INVX1 g123202(.A (n_13448), .Y (n_22032));
INVX1 g123204(.A (n_13758), .Y (n_24105));
INVX1 g123207(.A (n_13758), .Y (n_14339));
INVX2 g123209(.A (n_25054), .Y (n_25198));
INVX4 g123218(.A (n_25302), .Y (n_19330));
INVX4 g123224(.A (n_13444), .Y (n_17713));
INVX4 g123230(.A (n_26315), .Y (n_13990));
INVX1 g123253(.A (n_13641), .Y (n_24249));
INVX2 g123296(.A (n_13654), .Y (n_13600));
INVX8 g123306(.A (n_13647), .Y (n_18384));
INVX2 g123309(.A (n_13652), .Y (n_22406));
INVX4 g123401(.A (n_13653), .Y (n_18137));
INVX1 g123414(.A (n_13437), .Y (n_26631));
INVX1 g123421(.A (n_13633), .Y (n_27950));
INVX1 g123434(.A (n_14218), .Y (n_22080));
INVX1 g123437(.A (n_14218), .Y (n_19597));
INVX1 g123438(.A (n_14218), .Y (n_19595));
INVX1 g123442(.A (n_13435), .Y (n_23329));
INVX1 g123451(.A (n_13629), .Y (n_25193));
INVX1 g123466(.A (n_13432), .Y (n_17340));
CLKBUFX3 g123577(.A (n_13429), .Y (n_13852));
INVX2 g123592(.A (n_13428), .Y (n_13854));
INVX1 g123622(.A (n_13668), .Y (n_23725));
INVX1 g123627(.A (n_13665), .Y (n_13574));
INVX1 g123641(.A (n_13427), .Y (n_13572));
INVX1 g123660(.A (n_34499), .Y (n_13813));
INVX1 g123670(.A (n_13426), .Y (n_13862));
INVX2 g123688(.A (n_13661), .Y (n_17719));
INVX1 g123717(.A (n_24101), .Y (n_13425));
INVX2 g123297(.A (n_13280), .Y (n_13654));
CLKBUFX3 g123689(.A (n_34498), .Y (n_13661));
CLKBUFX1 gbuf_d_480(.A(n_13094), .Y(d_out_480));
CLKBUFX1 gbuf_q_480(.A(q_in_480), .Y(addr_425));
INVX2 g123628(.A (n_13264), .Y (n_13665));
INVX1 g123225(.A (n_13284), .Y (n_13444));
INVX2 g123211(.A (n_13285), .Y (n_13637));
CLKBUFX1 g123595(.A (n_34686), .Y (n_13613));
CLKBUFX3 g123576(.A (n_13421), .Y (n_13559));
INVX4 g122802(.A (n_13419), .Y (n_13478));
INVX4 g122778(.A (n_13311), .Y (n_13696));
XOR2X1 g121233(.A (n_11961), .B (n_13039), .Y (n_13418));
CLKBUFX3 g122774(.A (n_13312), .Y (n_13737));
NAND2X1 g121257(.A (n_13416), .B (n_13123), .Y (n_13417));
INVX4 g122752(.A (n_13415), .Y (n_25877));
CLKBUFX1 g122750(.A (n_13415), .Y (n_13739));
NAND2X1 g121284(.A (n_13413), .B (n_13121), .Y (n_35442));
INVX2 g123404(.A (n_13277), .Y (n_13624));
INVX2 g123460(.A (n_13412), .Y (n_13629));
AOI22X1 g121423(.A0 (n_13230), .A1 (n_13034), .B0 (n_11559), .B1(n_13112), .Y (n_13553));
OAI21X1 g121426(.A0 (n_33094), .A1 (n_13032), .B0 (n_11046), .Y(n_13552));
AOI22X1 g121431(.A0 (n_33290), .A1 (n_13031), .B0 (n_11987), .B1(n_32827), .Y (n_13411));
NAND2X1 g121442(.A (n_11965), .B (n_13128), .Y (n_14452));
OAI21X1 g121449(.A0 (n_35873), .A1 (n_7769), .B0 (n_11272), .Y(n_13410));
AOI22X1 g121453(.A0 (n_13409), .A1 (n_13028), .B0 (n_17468), .B1(n_13408), .Y (n_13549));
NAND2X1 g121457(.A (n_13234), .B (n_10472), .Y (n_13407));
OR2X1 g121477(.A (n_13992), .B (n_13318), .Y (n_13406));
NAND2X1 g121478(.A (n_13413), .B (n_13104), .Y (n_13404));
NAND2X1 g121479(.A (n_13413), .B (n_13100), .Y (n_13403));
NAND2X1 g121488(.A (n_12954), .B (n_13105), .Y (n_13402));
INVX1 g123443(.A (n_13412), .Y (n_13435));
NAND2X1 g121540(.A (n_8124), .B (n_13103), .Y (n_13401));
INVX2 g123415(.A (n_13277), .Y (n_13437));
OAI21X1 g121587(.A0 (n_7613), .A1 (n_12994), .B0 (n_12154), .Y(n_14865));
OAI21X1 g121594(.A0 (n_13400), .A1 (n_12991), .B0 (n_11480), .Y(n_14010));
NAND2X1 g121597(.A (n_12156), .B (n_13119), .Y (n_14862));
INVX1 g121600(.A (n_13399), .Y (n_13533));
OAI21X1 g121607(.A0 (n_33094), .A1 (n_12993), .B0 (n_11044), .Y(n_14226));
NOR2X1 g121609(.A (n_11245), .B (n_13117), .Y (n_14682));
NAND2X1 g121631(.A (n_11955), .B (n_13120), .Y (n_14655));
NAND2X1 g121725(.A (n_13393), .B (n_13088), .Y (n_13394));
NOR2X1 g121834(.A (n_11479), .B (n_13097), .Y (n_14614));
AOI22X1 g121838(.A0 (n_8124), .A1 (n_12987), .B0 (n_13102), .B1(n_13106), .Y (n_14636));
NAND2X1 g121886(.A (n_13736), .B (n_3887), .Y (n_14437));
NAND2X1 g121888(.A (n_13736), .B (n_13389), .Y (n_13520));
NAND2X1 g121889(.A (n_13166), .B (n_13388), .Y (n_15295));
NAND2X1 g121890(.A (n_13736), .B (n_13387), .Y (n_15407));
NAND2X1 g121891(.A (n_13736), .B (n_13386), .Y (n_14247));
NAND2X1 g121895(.A (n_13166), .B (n_13385), .Y (n_13518));
NAND2X1 g121896(.A (n_13736), .B (n_13383), .Y (n_14207));
NAND2X1 g121897(.A (n_13736), .B (n_13381), .Y (n_14398));
NAND2X1 g121900(.A (n_13736), .B (n_13380), .Y (n_14930));
NAND2X1 g121927(.A (n_13736), .B (n_13379), .Y (n_14478));
NAND2X1 g121947(.A (n_13736), .B (n_13378), .Y (n_14473));
NAND2X1 g121948(.A (n_35834), .B (P3_reg2[29] ), .Y (n_29690));
NAND2X1 g121952(.A (n_13374), .B (n_13377), .Y (n_25846));
NOR2X1 g121964(.A (n_12451), .B (n_13078), .Y (n_13376));
NAND2X1 g121969(.A (n_13736), .B (n_13375), .Y (n_14983));
NAND2X1 g121978(.A (n_13214), .B (n_10097), .Y (n_14740));
NAND2X1 g121982(.A (n_13214), .B (n_10582), .Y (n_14375));
NAND2X1 g121984(.A (n_13374), .B (n_13373), .Y (n_25847));
NAND2X1 g121998(.A (n_35719), .B (n_14317), .Y (n_13372));
NAND2X1 g122003(.A (n_35768), .B (P3_reg2[15] ), .Y (n_26074));
NAND2X1 g122004(.A (n_13214), .B (n_13370), .Y (n_14600));
NAND2X1 g122017(.A (n_35829), .B (n_13368), .Y (n_27756));
NAND2X1 g122021(.A (n_13736), .B (n_13367), .Y (n_27687));
NAND2X1 g122025(.A (n_35844), .B (n_13366), .Y (n_24785));
NAND2X1 g122030(.A (n_13374), .B (n_13365), .Y (n_26514));
NAND2X1 g122034(.A (n_35824), .B (P3_reg2[9] ), .Y (n_24764));
NOR2X1 g122054(.A (n_35816), .B (n_286), .Y (n_13509));
NAND2X1 g122072(.A (n_35766), .B (n_13361), .Y (n_23418));
NAND2X1 g122075(.A (n_13214), .B (n_10100), .Y (n_14660));
NAND2X1 g122089(.A (n_13736), .B (n_13359), .Y (n_28310));
NAND2X1 g122090(.A (n_35766), .B (n_13358), .Y (n_22024));
NAND2X1 g122093(.A (n_13736), .B (n_13357), .Y (n_27207));
NAND2X1 g122096(.A (n_13736), .B (n_13355), .Y (n_27686));
NAND2X1 g122098(.A (n_13736), .B (n_13354), .Y (n_28054));
NAND2X1 g122101(.A (n_13736), .B (n_13353), .Y (n_28538));
NAND2X1 g122104(.A (n_13736), .B (n_13351), .Y (n_27521));
INVX1 g122107(.A (n_13350), .Y (n_29576));
NAND2X1 g122113(.A (n_13736), .B (n_13348), .Y (n_28124));
INVX1 g122120(.A (n_13347), .Y (n_13967));
INVX1 g122122(.A (n_13346), .Y (n_13775));
NAND2X1 g122125(.A (n_35771), .B (n_13344), .Y (n_28532));
NAND2X1 g122132(.A (n_35840), .B (n_13343), .Y (n_27519));
NAND2X1 g122149(.A (n_35771), .B (n_13342), .Y (n_25838));
NAND2X1 g122160(.A (n_13736), .B (n_13341), .Y (n_13504));
NAND2X1 g122170(.A (n_13374), .B (n_13340), .Y (n_23996));
NAND2X1 g122206(.A (n_35844), .B (P3_reg2[13] ), .Y (n_25400));
NAND2X1 g122208(.A (n_35834), .B (n_13338), .Y (n_25329));
NAND2X1 g122213(.A (n_35719), .B (n_13337), .Y (n_21875));
NAND2X1 g122216(.A (n_35775), .B (n_13336), .Y (n_28302));
NAND2X1 g122220(.A (n_35775), .B (n_13335), .Y (n_27681));
NAND2X1 g122224(.A (n_35840), .B (n_13334), .Y (n_28083));
INVX1 g122226(.A (n_28153), .Y (n_13333));
NAND2X1 g122235(.A (n_35844), .B (n_13332), .Y (n_21600));
NAND2X1 g122238(.A (n_13736), .B (n_13330), .Y (n_29662));
NAND2X1 g122240(.A (n_35829), .B (P3_reg2[28] ), .Y (n_29478));
NAND2X1 g122241(.A (n_35840), .B (n_13329), .Y (n_26774));
NAND2X1 g122244(.A (n_35834), .B (P3_reg2[6] ), .Y (n_23932));
NAND2X1 g122246(.A (n_13214), .B (n_13327), .Y (n_14920));
NAND2X1 g122255(.A (n_35766), .B (P3_reg2[30] ), .Y (n_13499));
INVX1 g122339(.A (n_13954), .Y (n_13325));
OAI21X1 g122344(.A0 (n_16186), .A1 (n_12690), .B0 (n_13076), .Y(n_13766));
INVX1 g122371(.A (n_28327), .Y (n_13323));
INVX1 g122376(.A (n_34773), .Y (n_13494));
NAND2X1 g122389(.A (n_13321), .B (n_13322), .Y (n_18303));
NAND2X1 g122391(.A (n_13663), .B (n_3235), .Y (n_22954));
NAND2X1 g122393(.A (n_13321), .B (P1_reg1[14] ), .Y (n_25679));
NAND2X1 g122404(.A (n_13317), .B (n_3402), .Y (n_23642));
NAND2X1 g122408(.A (n_13316), .B (n_4554), .Y (n_24840));
NAND2X1 g122409(.A (n_13134), .B (n_4231), .Y (n_24009));
NAND2X1 g122447(.A (n_13137), .B (n_10167), .Y (n_28195));
INVX1 g122468(.A (n_13320), .Y (n_24505));
NAND2X1 g122623(.A (n_13318), .B (n_10158), .Y (n_27702));
NAND2X1 g122632(.A (n_13321), .B (P1_reg1[12] ), .Y (n_25336));
NAND2X1 g122635(.A (n_13299), .B (n_10566), .Y (n_21889));
NAND2X1 g122698(.A (n_13318), .B (n_10136), .Y (n_27227));
NAND2X1 g122703(.A (n_13318), .B (P1_reg1[0] ), .Y (n_19325));
NAND2X1 g122704(.A (n_13318), .B (P1_reg1[19] ), .Y (n_28196));
NAND2X1 g122707(.A (n_13318), .B (n_4534), .Y (n_25680));
INVX1 g122713(.A (n_13181), .Y (n_13485));
NAND2X1 g122716(.A (n_13321), .B (n_4215), .Y (n_25682));
NAND2X1 g122719(.A (n_13317), .B (n_4920), .Y (n_25681));
NAND2X1 g122720(.A (n_13134), .B (P1_reg1[16] ), .Y (n_25849));
INVX1 g122734(.A (n_13180), .Y (n_13482));
NAND2X1 g122737(.A (n_13316), .B (n_10161), .Y (n_28064));
INVX2 g122764(.A (n_13313), .Y (n_13554));
INVX2 g122770(.A (n_13312), .Y (n_26584));
CLKBUFX3 g122782(.A (n_13419), .Y (n_13701));
INVX1 g122890(.A (n_25693), .Y (n_13304));
NAND2X1 g122893(.A (n_7730), .B (n_13145), .Y (n_25350));
NAND2X1 g122894(.A (n_2911), .B (n_13299), .Y (n_25856));
INVX1 g122897(.A (n_26791), .Y (n_14182));
NAND2X1 g122909(.A (n_10889), .B (n_13056), .Y (n_28569));
INVX1 g122912(.A (n_27727), .Y (n_14593));
INVX1 g122922(.A (n_13175), .Y (n_13469));
INVX1 g122931(.A (n_13174), .Y (n_13467));
INVX1 g122947(.A (n_13171), .Y (n_13464));
INVX1 g122952(.A (n_13170), .Y (n_15119));
NAND2X2 g122956(.A (n_13301), .B (n_13147), .Y (n_29034));
NAND2X1 g122957(.A (n_13145), .B (n_7515), .Y (n_22960));
NAND2X1 g122960(.A (n_7737), .B (n_13147), .Y (n_25355));
NAND2X1 g122961(.A (n_7546), .B (n_13788), .Y (n_24843));
NAND2X1 g122963(.A (n_2138), .B (n_13299), .Y (n_24011));
NAND2X1 g122966(.A (n_7819), .B (n_13147), .Y (n_27710));
NAND2X1 g122969(.A (n_7575), .B (n_13145), .Y (n_25713));
AOI21X1 g122974(.A0 (n_12981), .A1 (n_12913), .B0 (n_13296), .Y(n_13297));
NAND2X1 g123029(.A (n_3105), .B (n_13143), .Y (n_25690));
NAND2X1 g123033(.A (n_7957), .B (n_13145), .Y (n_28204));
INVX1 g123113(.A (n_14793), .Y (n_13455));
NOR2X1 g123115(.A (n_11742), .B (n_13064), .Y (n_14539));
NAND2X1 g123134(.A (n_12147), .B (n_13049), .Y (n_14325));
INVX1 g123180(.A (n_13489), .Y (n_28734));
BUFX3 g123182(.A (n_13287), .Y (n_28441));
INVX4 g123192(.A (n_13287), .Y (n_13657));
INVX2 g123199(.A (n_13285), .Y (n_13644));
INVX1 g123203(.A (n_13285), .Y (n_13448));
INVX1 g123208(.A (n_13285), .Y (n_13758));
INVX1 g123210(.A (n_13285), .Y (n_25054));
BUFX1 g123219(.A (n_13284), .Y (n_25302));
INVX1 g123220(.A (n_13284), .Y (n_13659));
INVX4 g123234(.A (n_13283), .Y (n_26315));
INVX2 g123239(.A (n_13283), .Y (n_21919));
INVX1 g123241(.A (n_13284), .Y (n_13651));
INVX1 g123242(.A (n_13284), .Y (n_13627));
INVX2 g123270(.A (n_13281), .Y (n_13641));
INVX1 g123288(.A (n_13280), .Y (n_13564));
INVX4 g123307(.A (n_13279), .Y (n_13647));
INVX2 g123310(.A (n_13281), .Y (n_13652));
INVX1 g123405(.A (n_13277), .Y (n_13634));
INVX4 g123406(.A (n_13277), .Y (n_13653));
BUFX3 g123408(.A (n_13277), .Y (n_26637));
INVX1 g123422(.A (n_13277), .Y (n_13633));
INVX1 g123428(.A (n_13274), .Y (n_13273));
INVX2 g123435(.A (n_24348), .Y (n_14218));
INVX4 g123449(.A (n_13412), .Y (n_13434));
INVX2 g123467(.A (n_13412), .Y (n_13432));
INVX4 g123503(.A (n_13268), .Y (n_14261));
INVX1 g123531(.A (n_24361), .Y (n_13976));
INVX4 g123586(.A (n_13421), .Y (n_13429));
INVX1 g123594(.A (n_34686), .Y (n_13428));
INVX1 g123623(.A (n_13264), .Y (n_13668));
INVX1 g123642(.A (n_13264), .Y (n_13427));
INVX1 g123684(.A (n_34498), .Y (n_13426));
INVX1 g123696(.A (n_24312), .Y (n_25605));
INVX1 g123700(.A (n_24312), .Y (n_18294));
INVX1 g123701(.A (n_24312), .Y (n_17674));
INVX1 g123707(.A (n_13179), .Y (n_25734));
INVX1 g123708(.A (n_13179), .Y (n_25207));
INVX2 g123710(.A (n_13179), .Y (n_27091));
INVX2 g123727(.A (n_27422), .Y (n_13781));
INVX1 g123741(.A (n_13318), .Y (n_19577));
INVX2 g123759(.A (n_26676), .Y (n_17287));
CLKBUFX1 gbuf_d_481(.A(n_13092), .Y(d_out_481));
CLKBUFX1 gbuf_q_481(.A(q_in_481), .Y(n_482));
INVX1 g123737(.A (n_13317), .Y (n_25098));
CLKBUFX1 gbuf_d_482(.A(n_13017), .Y(d_out_482));
CLKBUFX1 gbuf_q_482(.A(q_in_482), .Y(n_9655));
CLKBUFX1 gbuf_d_483(.A(n_13027), .Y(d_out_483));
CLKBUFX1 gbuf_q_483(.A(q_in_483), .Y(addr_491));
CLKBUFX1 gbuf_d_484(.A(n_12996), .Y(d_out_484));
CLKBUFX1 gbuf_q_484(.A(q_in_484), .Y(addr_488));
CLKBUFX1 gbuf_d_485(.A(n_13000), .Y(d_out_485));
CLKBUFX1 gbuf_q_485(.A(q_in_485), .Y(addr_489));
CLKBUFX1 gbuf_d_486(.A(n_13004), .Y(d_out_486));
CLKBUFX1 gbuf_q_486(.A(q_in_486), .Y(n_1170));
CLKBUFX1 gbuf_d_487(.A(n_13025), .Y(d_out_487));
CLKBUFX1 gbuf_q_487(.A(q_in_487), .Y(addr_494));
CLKBUFX1 gbuf_d_488(.A(n_13015), .Y(d_out_488));
CLKBUFX1 gbuf_q_488(.A(q_in_488), .Y(addr_495));
CLKBUFX1 gbuf_d_489(.A(n_13022), .Y(d_out_489));
CLKBUFX1 gbuf_q_489(.A(q_in_489), .Y(n_9663));
CLKBUFX1 gbuf_d_490(.A(n_13006), .Y(d_out_490));
CLKBUFX1 gbuf_q_490(.A(q_in_490), .Y(n_9675));
CLKBUFX1 gbuf_d_491(.A(n_13011), .Y(d_out_491));
CLKBUFX1 gbuf_q_491(.A(q_in_491), .Y(addr_497));
CLKBUFX1 gbuf_d_492(.A(n_13020), .Y(d_out_492));
CLKBUFX1 gbuf_q_492(.A(q_in_492), .Y(addr_492));
CLKBUFX1 gbuf_d_493(.A(n_13013), .Y(d_out_493));
CLKBUFX1 gbuf_q_493(.A(q_in_493), .Y(addr_496));
INVX1 g123643(.A (n_34497), .Y (n_13264));
CLKBUFX1 gbuf_d_494(.A(n_12998), .Y(d_out_494));
CLKBUFX1 gbuf_q_494(.A(q_in_494), .Y(addr_490));
CLKBUFX1 gbuf_d_495(.A(n_13008), .Y(d_out_495));
CLKBUFX1 gbuf_q_495(.A(q_in_495), .Y(n_9658));
CLKBUFX1 gbuf_d_496(.A(n_13002), .Y(d_out_496));
CLKBUFX1 gbuf_q_496(.A(q_in_496), .Y(addr_487));
NAND2X1 g122914(.A (n_8207), .B (n_13183), .Y (n_27727));
NAND2X1 g122384(.A (n_13184), .B (n_3337), .Y (n_21942));
INVX2 g122810(.A (n_13252), .Y (n_13419));
CLKBUFX3 g122781(.A (n_13252), .Y (n_13311));
NAND2X1 g121254(.A (n_13413), .B (n_13038), .Y (n_13251));
INVX1 g122769(.A (n_13252), .Y (n_13313));
NAND2X1 g121491(.A (n_8124), .B (n_13033), .Y (n_13248));
NAND4X1 g121506(.A (n_13101), .B (n_16435), .C (n_32041), .D(n_17906), .Y (n_13245));
CLKBUFX1 g123440(.A (n_13243), .Y (n_24348));
INVX1 g121588(.A (n_14419), .Y (n_13242));
AOI22X1 g121601(.A0 (n_8124), .A1 (n_12952), .B0 (n_17467), .B1(n_13408), .Y (n_13399));
INVX1 g121613(.A (n_13240), .Y (n_13396));
INVX2 g123407(.A (n_13239), .Y (n_13277));
XOR2X1 g121633(.A (n_10658), .B (n_12973), .Y (n_13238));
NAND2X1 g121697(.A (n_33290), .B (n_13040), .Y (n_13237));
NOR2X1 g121710(.A (rd_2), .B (n_1170), .Y (n_13236));
INVX1 g121776(.A (n_13234), .Y (n_13235));
NAND4X1 g121778(.A (n_12563), .B (n_18164), .C (n_12840), .D(n_11548), .Y (n_13544));
NAND4X1 g121779(.A (n_12696), .B (n_11333), .C (n_13085), .D(n_13232), .Y (n_13233));
NAND3X1 g121806(.A (n_12203), .B (n_12449), .C (n_13222), .Y(n_13231));
AOI22X1 g121845(.A0 (n_13230), .A1 (n_12933), .B0 (n_10330), .B1(n_13527), .Y (n_14219));
INVX1 g121851(.A (n_13111), .Y (n_13983));
INVX1 g121854(.A (n_13228), .Y (n_13227));
XOR2X1 g121872(.A (n_34384), .B (n_12948), .Y (n_13225));
MX2X1 g121875(.A (n_18536), .B (n_11034), .S0 (n_13222), .Y(n_13223));
XOR2X1 g121877(.A (n_32349), .B (n_12947), .Y (n_13221));
XOR2X1 g121878(.A (n_17909), .B (n_12941), .Y (n_13220));
MX2X1 g121879(.A (n_9482), .B (n_8737), .S0 (n_12945), .Y (n_13219));
NOR2X1 g121990(.A (rd_1), .B (addr_442), .Y (n_13217));
NAND2X1 g122028(.A (n_13214), .B (n_13216), .Y (n_26780));
NAND2X1 g122049(.A (n_13214), .B (n_13215), .Y (n_19422));
NAND2X1 g122063(.A (n_13214), .B (n_13213), .Y (n_25396));
NAND2X1 g122087(.A (n_13214), .B (n_13212), .Y (n_26401));
NAND2X1 g122088(.A (n_13214), .B (n_13211), .Y (n_21900));
NOR2X1 g122108(.A (n_13131), .B (n_7043), .Y (n_13350));
NAND2X1 g122116(.A (n_13214), .B (n_13209), .Y (n_21622));
NAND2X1 g122121(.A (n_13214), .B (n_14513), .Y (n_13347));
NAND2X1 g122123(.A (n_13214), .B (n_14168), .Y (n_13346));
NAND2X1 g122126(.A (n_13214), .B (n_13208), .Y (n_23635));
NAND2X1 g122129(.A (n_13214), .B (n_13207), .Y (n_23379));
NAND2X1 g122134(.A (n_13214), .B (n_13206), .Y (n_24717));
NAND2X1 g122143(.A (n_13214), .B (n_13205), .Y (n_23904));
NAND2X1 g122209(.A (n_13214), .B (n_13204), .Y (n_24719));
NAND2X1 g122212(.A (n_13214), .B (n_13203), .Y (n_26854));
NAND2X1 g122223(.A (n_13214), .B (n_13202), .Y (n_22012));
NAND2X1 g122227(.A (n_35844), .B (n_13201), .Y (n_28153));
NAND2X1 g122245(.A (n_13214), .B (n_13200), .Y (n_25331));
NAND2X1 g122247(.A (n_13214), .B (n_13199), .Y (n_24718));
OAI21X1 g122296(.A0 (n_12921), .A1 (n_13197), .B0 (n_13196), .Y(n_13198));
OAI21X1 g122297(.A0 (n_12925), .A1 (n_13024), .B0 (n_13194), .Y(n_13195));
OAI21X1 g122298(.A0 (n_12920), .A1 (n_13024), .B0 (n_13192), .Y(n_13193));
OAI21X1 g122304(.A0 (n_12927), .A1 (n_13024), .B0 (n_13189), .Y(n_13191));
OAI21X1 g122315(.A0 (n_12918), .A1 (n_13197), .B0 (n_13187), .Y(n_13188));
INVX1 g122330(.A (n_14202), .Y (n_13186));
OAI21X1 g122341(.A0 (n_33094), .A1 (n_12915), .B0 (n_10747), .Y(n_13954));
NAND2X1 g122372(.A (n_24312), .B (n_10247), .Y (n_28327));
NAND2X1 g122394(.A (n_13185), .B (n_3333), .Y (n_22760));
NAND2X1 g122397(.A (n_13185), .B (n_3716), .Y (n_23643));
NAND2X1 g122411(.A (n_13184), .B (n_4011), .Y (n_25056));
NOR2X1 g122470(.A (n_13080), .B (n_182), .Y (n_13320));
NAND2X1 g122602(.A (n_13183), .B (n_11135), .Y (n_19327));
NAND2X1 g122651(.A (n_13056), .B (n_10854), .Y (n_21939));
NAND2X1 g122652(.A (n_24312), .B (P1_reg1[1] ), .Y (n_21892));
NAND2X1 g122655(.A (n_1003), .B (n_13183), .Y (n_22759));
NAND2X1 g122705(.A (n_24312), .B (n_3958), .Y (n_24721));
NAND2X1 g122714(.A (n_13179), .B (P1_reg1[24] ), .Y (n_13181));
NAND2X1 g122717(.A (n_13184), .B (n_10215), .Y (n_28542));
NAND2X1 g122735(.A (n_13179), .B (n_10217), .Y (n_13180));
INVX1 g122753(.A (n_13252), .Y (n_13415));
INVX1 g122775(.A (n_13252), .Y (n_13312));
NAND2X1 g122891(.A (n_7724), .B (n_13056), .Y (n_25693));
NAND2X1 g122898(.A (n_10822), .B (n_13183), .Y (n_26791));
NAND2X1 g122904(.A (n_8001), .B (n_13183), .Y (n_28205));
NAND2X1 g122923(.A (n_3372), .B (n_13056), .Y (n_13175));
NAND2X1 g122932(.A (n_13173), .B (n_13056), .Y (n_13174));
NAND2X1 g122948(.A (n_10885), .B (n_13056), .Y (n_13171));
NAND2X1 g122953(.A (n_13169), .B (n_13183), .Y (n_13170));
NAND2X1 g122958(.A (n_13167), .B (n_13183), .Y (n_23648));
NAND2X1 g122959(.A (n_10880), .B (n_13183), .Y (n_23647));
NAND2X1 g122964(.A (n_2601), .B (n_13056), .Y (n_25058));
INVX4 g122975(.A (n_13166), .Y (n_18546));
INVX2 g122987(.A (n_13163), .Y (n_13957));
INVX4 g122995(.A (n_13736), .Y (n_18262));
INVX4 g123017(.A (n_13736), .Y (n_17968));
INVX2 g123019(.A (n_13736), .Y (n_24965));
NAND2X1 g123035(.A (n_7706), .B (n_13183), .Y (n_25049));
AOI22X1 g123114(.A0 (n_33290), .A1 (n_12907), .B0 (n_11464), .B1(n_32827), .Y (n_14793));
AOI22X1 g123120(.A0 (n_13540), .A1 (n_12908), .B0 (n_11555), .B1(n_12953), .Y (n_14331));
INVX1 g123125(.A (n_35395), .Y (n_13154));
CLKBUFX1 g123181(.A (n_13152), .Y (n_13489));
INVX2 g123193(.A (n_13152), .Y (n_13287));
INVX2 g123212(.A (n_13151), .Y (n_13285));
INVX2 g123226(.A (n_13151), .Y (n_13284));
CLKBUFX3 g123240(.A (n_13151), .Y (n_13283));
INVX2 g123271(.A (n_13150), .Y (n_13281));
INVX1 g123298(.A (n_13150), .Y (n_13280));
INVX1 g123308(.A (n_13150), .Y (n_13279));
INVX1 g123425(.A (n_13243), .Y (n_13488));
BUFX3 g123433(.A (n_13243), .Y (n_13274));
INVX2 g123468(.A (n_13239), .Y (n_13412));
INVX1 g123484(.A (n_13299), .Y (n_25956));
INVX4 g123493(.A (n_13147), .Y (n_23192));
INVX1 g123495(.A (n_35054), .Y (n_14702));
INVX2 g123505(.A (n_13145), .Y (n_13268));
INVX1 g123509(.A (n_13788), .Y (n_26965));
INVX2 g123511(.A (n_13143), .Y (n_22994));
INVX1 g123519(.A (n_25694), .Y (n_14731));
INVX1 g123520(.A (n_25694), .Y (n_23149));
INVX1 g123521(.A (n_25694), .Y (n_23457));
CLKBUFX1 g123528(.A (n_24361), .Y (n_14235));
INVX2 g123587(.A (n_34685), .Y (n_13421));
INVX4 g123719(.A (n_13316), .Y (n_24101));
INVX1 g123728(.A (n_13137), .Y (n_27422));
INVX1 g123731(.A (n_13318), .Y (n_27089));
INVX1 g123744(.A (n_13318), .Y (n_18065));
INVX2 g123753(.A (n_13134), .Y (n_26676));
INVX1 g123757(.A (n_13663), .Y (n_22036));
INVX1 g123745(.A (n_13318), .Y (n_27747));
INVX4 g123738(.A (n_34418), .Y (n_13317));
INVX1 g123729(.A (n_13051), .Y (n_13137));
CLKBUFX1 gbuf_d_497(.A(n_12961), .Y(d_out_497));
CLKBUFX1 gbuf_qn_497(.A(qn_in_497), .Y(addr_444));
CLKBUFX1 gbuf_d_498(.A(n_12967), .Y(d_out_498));
CLKBUFX1 gbuf_q_498(.A(q_in_498), .Y(addr_446));
INVX2 g122990(.A (n_13130), .Y (n_13163));
INVX1 g122982(.A (n_13130), .Y (n_13374));
INVX1 g122978(.A (n_13130), .Y (n_13166));
CLKBUFX1 gbuf_d_499(.A(n_12963), .Y(d_out_499));
CLKBUFX1 gbuf_qn_499(.A(qn_in_499), .Y(addr_445));
INVX2 g123522(.A (n_13042), .Y (n_25694));
INVX2 g123510(.A (n_13058), .Y (n_13788));
INVX2 g123506(.A (n_13059), .Y (n_13145));
INVX4 g123494(.A (n_35053), .Y (n_13147));
INVX4 g123474(.A (n_13183), .Y (n_27770));
NAND2X1 g121501(.A (n_33290), .B (n_12974), .Y (n_13128));
INVX2 g123424(.A (n_13062), .Y (n_13239));
NAND3X1 g121584(.A (n_12972), .B (n_32221), .C (n_12790), .Y(n_13126));
NAND3X1 g121585(.A (n_13122), .B (n_35433), .C (n_12787), .Y(n_13125));
OAI21X1 g121589(.A0 (n_7613), .A1 (n_12869), .B0 (n_11738), .Y(n_14419));
AOI22X1 g121614(.A0 (n_13409), .A1 (n_12867), .B0 (n_9761), .B1(n_13408), .Y (n_13240));
AOI21X1 g121634(.A0 (n_12977), .A1 (n_12976), .B0 (n_12978), .Y(n_13124));
XOR2X1 g121635(.A (n_35860), .B (n_13122), .Y (n_13123));
XOR2X1 g121640(.A (n_11498), .B (n_12900), .Y (n_13121));
NAND2X1 g121706(.A (n_33290), .B (n_12949), .Y (n_13120));
NAND2X1 g121708(.A (n_33290), .B (n_12950), .Y (n_13119));
NOR2X1 g121733(.A (n_33094), .B (n_12951), .Y (n_13117));
NAND4X1 g121777(.A (n_12796), .B (n_18159), .C (n_12759), .D(n_13114), .Y (n_13234));
AOI22X1 g121841(.A0 (n_33290), .A1 (n_12852), .B0 (n_12827), .B1(n_32827), .Y (n_15179));
AOI22X1 g121847(.A0 (n_13230), .A1 (n_12850), .B0 (n_18584), .B1(n_12953), .Y (n_13992));
AOI22X1 g121848(.A0 (n_13230), .A1 (n_12846), .B0 (n_11034), .B1(n_13112), .Y (n_14001));
AOI22X1 g121852(.A0 (n_13409), .A1 (n_12848), .B0 (n_17472), .B1(n_13408), .Y (n_13111));
NAND2X1 g121856(.A (n_11504), .B (n_12971), .Y (n_13228));
AOI22X1 g121863(.A0 (n_8124), .A1 (n_12845), .B0 (n_10287), .B1(n_13106), .Y (n_14385));
XOR2X1 g121866(.A (n_16442), .B (n_34872), .Y (n_13105));
XOR2X1 g121867(.A (n_34610), .B (n_12862), .Y (n_13104));
XOR2X1 g121869(.A (n_13102), .B (n_13101), .Y (n_13103));
XOR2X1 g121871(.A (n_11716), .B (n_12861), .Y (n_13100));
INVX1 g121881(.A (rd_2), .Y (n_13098));
NOR2X1 g121945(.A (n_7613), .B (n_12934), .Y (n_13097));
OR4X1 g122099(.A (n_12702), .B (n_11571), .C (n_13095), .D (n_12720),.Y (n_13096));
OAI21X1 g122320(.A0 (n_12832), .A1 (n_31726), .B0 (n_13093), .Y(n_13094));
OAI21X1 g122321(.A0 (n_12831), .A1 (n_30783), .B0 (n_13091), .Y(n_13092));
OAI21X1 g122331(.A0 (n_7613), .A1 (n_12829), .B0 (n_11253), .Y(n_14202));
AOI21X1 g122346(.A0 (n_12939), .A1 (n_11333), .B0 (n_12940), .Y(n_13090));
XOR2X1 g122356(.A (n_9744), .B (n_12838), .Y (n_13088));
AOI21X1 g122357(.A0 (n_12943), .A1 (n_12942), .B0 (n_12944), .Y(n_13087));
XOR2X1 g122359(.A (n_35212), .B (n_13085), .Y (n_13086));
XOR2X1 g122364(.A (n_17955), .B (n_12844), .Y (n_13084));
XOR2X1 g122365(.A (n_10755), .B (n_12840), .Y (n_13082));
INVX1 g122367(.A (rd_1), .Y (n_13081));
INVX1 g123755(.A (n_13080), .Y (n_13321));
INVX2 g122811(.A (n_12989), .Y (n_13252));
NAND4X1 g122888(.A (n_12013), .B (n_11962), .C (n_11716), .D(n_12701), .Y (n_13078));
INVX8 g122996(.A (n_13131), .Y (n_13736));
INVX4 g123009(.A (n_13214), .Y (n_14439));
NAND2X1 g123030(.A (n_13075), .B (n_12916), .Y (n_13076));
INVX1 g123123(.A (n_13072), .Y (n_13156));
INVX1 g123194(.A (n_13068), .Y (n_13152));
INVX2 g123244(.A (n_13068), .Y (n_13151));
NAND2X1 g123316(.A (n_13054), .B (n_13067), .Y (n_13150));
NAND2X2 g123397(.A (n_13065), .B (n_13053), .Y (n_13066));
NOR2X1 g123398(.A (n_7613), .B (n_12912), .Y (n_13064));
CLKBUFX1 g123441(.A (n_13062), .Y (n_13243));
INVX1 g123485(.A (n_13060), .Y (n_13299));
INVX1 g123513(.A (n_13058), .Y (n_13143));
INVX4 g123533(.A (n_13056), .Y (n_24361));
NOR2X1 g123544(.A (n_7555), .B (n_12911), .Y (n_13055));
INVX1 g123703(.A (n_24312), .Y (n_21092));
INVX1 g123704(.A (n_24312), .Y (n_24386));
INVX2 g123722(.A (n_13051), .Y (n_13316));
INVX4 g123743(.A (n_34418), .Y (n_13318));
INVX2 g123751(.A (n_13184), .Y (n_23356));
INVX1 g123754(.A (n_13080), .Y (n_13134));
INVX1 g123758(.A (n_13080), .Y (n_13663));
NAND2X1 g123767(.A (n_33290), .B (n_12910), .Y (n_13049));
CLKBUFX1 gbuf_d_500(.A(n_12956), .Y(d_out_500));
CLKBUFX1 gbuf_q_500(.A(q_in_500), .Y(addr_461));
CLKBUFX1 gbuf_d_501(.A(n_12959), .Y(d_out_501));
CLKBUFX1 gbuf_q_501(.A(q_in_501), .Y(n_628));
CLKBUFX1 gbuf_d_502(.A(n_12970), .Y(d_out_502));
CLKBUFX1 gbuf_qn_502(.A(qn_in_502), .Y(addr_443));
CLKBUFX1 gbuf_d_503(.A(n_12965), .Y(d_out_503));
CLKBUFX1 gbuf_q_503(.A(q_in_503), .Y(addr_2));
CLKBUFX1 gbuf_d_504(.A(n_12893), .Y(d_out_504));
CLKBUFX1 gbuf_q_504(.A(q_in_504), .Y(addr_453));
INVX1 g123713(.A (n_13046), .Y (n_13179));
CLKBUFX1 gbuf_d_505(.A(n_12880), .Y(d_out_505));
CLKBUFX1 gbuf_q_505(.A(q_in_505), .Y(addr_457));
CLKBUFX1 gbuf_d_506(.A(n_12895), .Y(d_out_506));
CLKBUFX1 gbuf_q_506(.A(q_in_506), .Y(addr_450));
CLKBUFX1 gbuf_d_507(.A(n_12874), .Y(d_out_507));
CLKBUFX1 gbuf_q_507(.A(q_in_507), .Y(addr_454));
INVX4 g123699(.A (n_13046), .Y (n_24312));
CLKBUFX1 gbuf_d_508(.A(n_12823), .Y(d_out_508));
CLKBUFX1 gbuf_q_508(.A(q_in_508), .Y(addr_429));
INVX2 g123021(.A (n_13045), .Y (n_13131));
CLKBUFX1 gbuf_d_509(.A(n_12885), .Y(d_out_509));
CLKBUFX1 gbuf_q_509(.A(q_in_509), .Y(n_7839));
INVX1 g123245(.A (n_12931), .Y (n_13068));
CLKBUFX1 gbuf_d_510(.A(n_12891), .Y(d_out_510));
CLKBUFX1 gbuf_q_510(.A(q_in_510), .Y(n_7843));
CLKBUFX1 gbuf_d_511(.A(n_12887), .Y(d_out_511));
CLKBUFX1 gbuf_q_511(.A(q_in_511), .Y(n_481));
CLKBUFX1 g123752(.A (n_34416), .Y (n_13184));
CLKBUFX1 gbuf_d_512(.A(n_12897), .Y(d_out_512));
CLKBUFX1 gbuf_q_512(.A(q_in_512), .Y(addr_452));
CLKBUFX1 gbuf_d_513(.A(n_12876), .Y(d_out_513));
CLKBUFX1 gbuf_q_513(.A(q_in_513), .Y(n_8074));
CLKBUFX1 gbuf_d_514(.A(n_12882), .Y(d_out_514));
CLKBUFX1 gbuf_q_514(.A(q_in_514), .Y(addr_455));
CLKBUFX1 gbuf_d_515(.A(n_12815), .Y(d_out_515));
CLKBUFX1 gbuf_q_515(.A(q_in_515), .Y(addr_442));
CLKBUFX1 gbuf_d_516(.A(n_12809), .Y(d_out_516));
CLKBUFX1 gbuf_q_516(.A(q_in_516), .Y(addr_435));
CLKBUFX1 gbuf_d_517(.A(n_12817), .Y(d_out_517));
CLKBUFX1 gbuf_q_517(.A(q_in_517), .Y(addr_1));
CLKBUFX1 gbuf_d_518(.A(n_12825), .Y(d_out_518));
CLKBUFX1 gbuf_q_518(.A(q_in_518), .Y(n_8361));
CLKBUFX1 gbuf_d_519(.A(n_12872), .Y(d_out_519));
CLKBUFX1 gbuf_q_519(.A(q_in_519), .Y(addr_451));
CLKBUFX1 gbuf_d_520(.A(n_12878), .Y(d_out_520));
CLKBUFX1 gbuf_q_520(.A(q_in_520), .Y(addr_447));
AOI22X1 g123124(.A0 (n_8124), .A1 (n_12704), .B0 (n_35860), .B1(n_13408), .Y (n_13072));
CLKBUFX1 gbuf_d_521(.A(n_12807), .Y(d_out_521));
CLKBUFX1 gbuf_q_521(.A(q_in_521), .Y(addr_441));
INVX4 g123534(.A (n_13042), .Y (n_13056));
INVX1 g123514(.A (n_35052), .Y (n_13058));
CLKBUFX1 gbuf_d_522(.A(n_12821), .Y(d_out_522));
CLKBUFX1 gbuf_q_522(.A(q_in_522), .Y(addr_430));
XOR2X1 g122352(.A (n_11712), .B (n_12767), .Y (n_13040));
INVX1 g123486(.A (n_35052), .Y (n_13060));
NAND3X1 g121583(.A (n_12312), .B (n_12791), .C (n_12899), .Y(n_13039));
XOR2X1 g121632(.A (n_16754), .B (n_12793), .Y (n_13038));
CLKBUFX1 gbuf_d_523(.A(n_12811), .Y(d_out_523));
CLKBUFX1 gbuf_q_523(.A(q_in_523), .Y(addr_424));
INVX1 g121861(.A (n_13035), .Y (n_13108));
XOR2X1 g121864(.A (n_9722), .B (n_12780), .Y (n_13034));
XOR2X1 g121865(.A (n_10540), .B (n_12772), .Y (n_13033));
XOR2X1 g121868(.A (n_13071), .B (n_12777), .Y (n_13032));
XOR2X1 g121870(.A (n_11464), .B (n_12784), .Y (n_13031));
MX2X1 g121874(.A (n_10329), .B (n_11089), .S0 (n_12786), .Y(n_35873));
XOR2X1 g121876(.A (n_10757), .B (n_12782), .Y (n_13028));
CLKBUFX1 gbuf_d_524(.A(n_12819), .Y(d_out_524));
CLKBUFX1 gbuf_q_524(.A(q_in_524), .Y(addr_438));
CLKBUFX1 gbuf_d_525(.A(n_12856), .Y(d_out_525));
CLKBUFX1 gbuf_q_525(.A(q_in_525), .Y(rd_2));
CLKBUFX1 gbuf_d_526(.A(n_12813), .Y(d_out_526));
CLKBUFX1 gbuf_q_526(.A(q_in_526), .Y(addr_439));
OAI21X1 g122278(.A0 (n_12736), .A1 (n_13019), .B0 (n_13026), .Y(n_13027));
OAI21X1 g122282(.A0 (n_12749), .A1 (n_13024), .B0 (n_13023), .Y(n_13025));
OAI21X1 g122286(.A0 (n_12754), .A1 (n_13024), .B0 (n_34196), .Y(n_13022));
OAI21X1 g122287(.A0 (n_12746), .A1 (n_13019), .B0 (n_13018), .Y(n_13020));
OAI21X1 g122288(.A0 (n_12752), .A1 (n_13019), .B0 (n_13016), .Y(n_13017));
OAI21X1 g122289(.A0 (n_12744), .A1 (n_13010), .B0 (n_13014), .Y(n_13015));
OAI21X1 g122290(.A0 (n_12742), .A1 (n_31979), .B0 (n_13012), .Y(n_13013));
OAI21X1 g122291(.A0 (n_12750), .A1 (n_13010), .B0 (n_13009), .Y(n_13011));
OAI21X1 g122292(.A0 (n_12741), .A1 (n_13010), .B0 (n_13007), .Y(n_13008));
OAI21X1 g122293(.A0 (n_12751), .A1 (n_13010), .B0 (n_13005), .Y(n_13006));
OAI21X1 g122295(.A0 (n_12756), .A1 (n_13197), .B0 (n_13003), .Y(n_13004));
OAI21X1 g122299(.A0 (n_12740), .A1 (n_13024), .B0 (n_13001), .Y(n_13002));
OAI21X1 g122300(.A0 (n_12738), .A1 (n_13019), .B0 (n_12999), .Y(n_13000));
OAI21X1 g122301(.A0 (n_12737), .A1 (n_13024), .B0 (n_12997), .Y(n_12998));
OAI21X1 g122305(.A0 (n_12735), .A1 (n_13024), .B0 (n_12995), .Y(n_12996));
AOI21X1 g122353(.A0 (n_11503), .A1 (n_12863), .B0 (n_12865), .Y(n_12994));
XOR2X1 g122355(.A (n_12992), .B (n_12763), .Y (n_12993));
AOI22X1 g122362(.A0 (n_9264), .A1 (n_12765), .B0 (n_9741), .B1(n_12764), .Y (n_12991));
CLKBUFX1 gbuf_d_527(.A(n_12901), .Y(d_out_527));
CLKBUFX1 gbuf_q_527(.A(q_in_527), .Y(rd_1));
NAND2X1 g122812(.A (n_12836), .B (n_12938), .Y (n_12989));
INVX1 g122991(.A (n_13045), .Y (n_13130));
BUFX3 g123023(.A (n_13045), .Y (n_13214));
AOI22X1 g123116(.A0 (n_13230), .A1 (n_12706), .B0 (n_11089), .B1(n_12953), .Y (n_13759));
INVX1 g123131(.A (n_12936), .Y (n_13716));
XOR2X1 g123142(.A (n_12986), .B (n_12722), .Y (n_12987));
INVX1 g123470(.A (n_12930), .Y (n_13062));
INVX8 g123476(.A (n_12985), .Y (n_13183));
INVX1 g123507(.A (n_35052), .Y (n_13059));
INVX1 g123706(.A (n_13046), .Y (n_13185));
INVX1 g123730(.A (n_34416), .Y (n_13051));
INVX1 g123762(.A (n_34416), .Y (n_13080));
AOI22X1 g123778(.A0 (n_33290), .A1 (n_12697), .B0 (n_11797), .B1(n_32827), .Y (n_14511));
AOI22X1 g123789(.A0 (n_13230), .A1 (n_12698), .B0 (n_9741), .B1(n_13527), .Y (n_14078));
NAND2X1 g123958(.A (n_18496), .B (n_12802), .Y (n_12981));
NAND2X1 g124003(.A (n_12798), .B (n_9375), .Y (n_12979));
CLKBUFX1 gbuf_d_528(.A(n_12853), .Y(d_out_528));
CLKBUFX1 gbuf_q_528(.A(q_in_528), .Y(P3_d));
CLKBUFX1 gbuf_d_529(.A(n_12889), .Y(d_out_529));
CLKBUFX1 gbuf_q_529(.A(q_in_529), .Y(addr_456));
CLKBUFX1 gbuf_d_530(.A(n_12729), .Y(d_out_530));
CLKBUFX1 gbuf_q_530(.A(q_in_530), .Y(addr_432));
CLKBUFX1 gbuf_d_531(.A(n_12694), .Y(d_out_531));
CLKBUFX1 gbuf_q_531(.A(q_in_531), .Y(datao_2[26]));
CLKBUFX1 gbuf_d_532(.A(n_12717), .Y(d_out_532));
CLKBUFX1 gbuf_q_532(.A(q_in_532), .Y(addr_437));
CLKBUFX1 gbuf_d_533(.A(n_12770), .Y(d_out_533));
CLKBUFX1 gbuf_q_533(.A(q_in_533), .Y(P2_d));
CLKBUFX1 gbuf_d_534(.A(n_12713), .Y(d_out_534));
CLKBUFX1 gbuf_q_534(.A(q_in_534), .Y(addr_433));
CLKBUFX3 g123482(.A (n_35051), .Y (n_12985));
CLKBUFX1 gbuf_d_535(.A(n_12715), .Y(d_out_535));
CLKBUFX1 gbuf_q_535(.A(q_in_535), .Y(n_8117));
CLKBUFX1 gbuf_d_536(.A(n_12724), .Y(d_out_536));
CLKBUFX1 gbuf_q_536(.A(q_in_536), .Y(addr_434));
CLKBUFX1 gbuf_d_537(.A(n_12719), .Y(d_out_537));
CLKBUFX1 gbuf_q_537(.A(q_in_537), .Y(addr_436));
NOR2X1 g121728(.A (n_12977), .B (n_12976), .Y (n_12978));
CLKBUFX1 gbuf_d_538(.A(n_12731), .Y(d_out_538));
CLKBUFX1 gbuf_q_538(.A(q_in_538), .Y(addr_431));
INVX1 g121831(.A (n_14213), .Y (n_12975));
OAI21X1 g121833(.A0 (n_13400), .A1 (n_12688), .B0 (n_10761), .Y(n_13988));
AOI22X1 g121862(.A0 (n_13409), .A1 (n_12689), .B0 (n_9962), .B1(n_13408), .Y (n_13035));
XOR2X1 g121873(.A (n_16895), .B (n_12693), .Y (n_12974));
INVX1 g122061(.A (n_12972), .Y (n_12973));
NAND2X1 g122234(.A (n_33290), .B (n_12769), .Y (n_12971));
OAI21X1 g122279(.A0 (n_12681), .A1 (n_12969), .B0 (n_12968), .Y(n_12970));
OAI21X1 g122280(.A0 (n_12676), .A1 (n_12969), .B0 (n_12966), .Y(n_12967));
OAI21X1 g122302(.A0 (n_12680), .A1 (n_12969), .B0 (n_12964), .Y(n_12965));
OAI21X1 g122311(.A0 (n_12677), .A1 (n_12969), .B0 (n_12962), .Y(n_12963));
OAI21X1 g122317(.A0 (n_12675), .A1 (n_12969), .B0 (n_12960), .Y(n_12961));
OAI21X1 g122322(.A0 (n_12684), .A1 (n_34375), .B0 (n_34973), .Y(n_12959));
OAI21X1 g122323(.A0 (n_12683), .A1 (n_34375), .B0 (n_12955), .Y(n_12956));
AOI22X1 g122336(.A0 (n_12954), .A1 (n_12673), .B0 (n_12232), .B1(n_12953), .Y (n_14373));
CLKBUFX1 gbuf_d_539(.A(n_12733), .Y(d_out_539));
CLKBUFX1 gbuf_q_539(.A(q_in_539), .Y(addr_426));
AOI22X1 g122337(.A0 (n_13230), .A1 (n_12672), .B0 (n_10333), .B1(n_13112), .Y (n_13782));
XOR2X1 g122358(.A (n_10314), .B (n_12857), .Y (n_12952));
XOR2X1 g122360(.A (n_11481), .B (n_12686), .Y (n_12951));
MX2X1 g122363(.A (n_11012), .B (n_12003), .S0 (n_12860), .Y(n_12950));
MX2X1 g122366(.A (n_11010), .B (n_12002), .S0 (n_12866), .Y(n_12949));
NOR2X1 g122396(.A (n_12037), .B (n_12843), .Y (n_13222));
NOR2X1 g122465(.A (n_12562), .B (n_12841), .Y (n_12948));
INVX1 g122519(.A (n_34616), .Y (n_12947));
OAI21X1 g122970(.A0 (n_12658), .A1 (n_12537), .B0 (n_9375), .Y(n_12945));
NOR2X1 g122972(.A (n_12943), .B (n_12942), .Y (n_12944));
NAND3X1 g123024(.A (n_12757), .B (n_12937), .C (n_12834), .Y(n_13045));
NOR2X1 g123031(.A (n_12695), .B (n_12839), .Y (n_12941));
NOR2X1 g123034(.A (n_12939), .B (n_11333), .Y (n_12940));
AOI22X1 g123132(.A0 (n_13409), .A1 (n_12656), .B0 (n_10757), .B1(n_13408), .Y (n_12936));
MX2X1 g123141(.A (n_35245), .B (n_35244), .S0 (n_12669), .Y(n_12934));
XOR2X1 g123149(.A (n_18584), .B (n_34874), .Y (n_12933));
NAND2X1 g123246(.A (n_12726), .B (n_12711), .Y (n_12931));
NAND2X1 g123471(.A (n_12726), .B (n_12709), .Y (n_12930));
CLKBUFX3 g123535(.A (n_35051), .Y (n_13042));
CLKBUFX3 g123714(.A (n_34415), .Y (n_13046));
AOI21X1 g123777(.A0 (n_11573), .A1 (n_12926), .B0 (n_12734), .Y(n_12927));
AOI22X1 g123797(.A0 (n_12641), .A1 (n_12739), .B0 (n_11811), .B1(n_12755), .Y (n_12925));
AOI22X1 g123808(.A0 (n_12639), .A1 (n_12753), .B0 (n_11814), .B1(n_12917), .Y (n_12921));
AOI22X1 g123809(.A0 (n_12638), .A1 (n_12739), .B0 (n_11809), .B1(n_12755), .Y (n_12920));
AOI22X1 g123810(.A0 (n_12635), .A1 (n_12739), .B0 (n_11807), .B1(n_12917), .Y (n_12918));
XOR2X1 g123821(.A (n_11470), .B (n_12654), .Y (n_12916));
AOI22X1 g123825(.A0 (n_17480), .A1 (n_12582), .B0 (n_10287), .B1(n_12721), .Y (n_12915));
INVX2 g123943(.A (n_12826), .Y (n_13065));
NAND2X1 g123950(.A (n_11218), .B (n_12801), .Y (n_12913));
INVX2 g123971(.A (n_12805), .Y (n_13054));
MX2X1 g123991(.A (n_10826), .B (n_17261), .S0 (n_12631), .Y(n_12912));
XOR2X1 g123993(.A (n_11215), .B (n_12633), .Y (n_12911));
XOR2X1 g123994(.A (n_11987), .B (n_12799), .Y (n_12910));
XOR2X1 g123995(.A (n_17182), .B (n_12627), .Y (n_12908));
XOR2X1 g123998(.A (n_16748), .B (n_12629), .Y (n_12907));
NAND2X1 g124004(.A (n_12905), .B (n_11333), .Y (n_12906));
CLKBUFX1 gbuf_d_540(.A(n_12623), .Y(d_out_540));
CLKBUFX1 gbuf_q_540(.A(q_in_540), .Y(datao_2[25]));
CLKBUFX1 gbuf_d_541(.A(n_12621), .Y(d_out_541));
CLKBUFX1 gbuf_q_541(.A(q_in_541), .Y(n_491));
CLKBUFX1 gbuf_d_542(.A(n_12624), .Y(d_out_542));
CLKBUFX1 gbuf_q_542(.A(q_in_542), .Y(datao_2[8]));
CLKBUFX1 gbuf_d_543(.A(n_12687), .Y(d_out_543));
CLKBUFX1 gbuf_qn_543(.A(qn_in_543), .Y(rd_3));
NAND2X1 g123399(.A (n_12657), .B (n_15981), .Y (n_12901));
OAI21X1 g121832(.A0 (n_7613), .A1 (n_12618), .B0 (n_10770), .Y(n_14213));
INVX1 g121924(.A (n_12899), .Y (n_12900));
NOR2X1 g122062(.A (n_11792), .B (n_12785), .Y (n_12972));
OR2X1 g122073(.A (n_12691), .B (n_6621), .Y (n_32189));
NOR2X1 g122083(.A (n_12038), .B (n_12781), .Y (n_13122));
OAI21X1 g122281(.A0 (n_12595), .A1 (n_27698), .B0 (n_12896), .Y(n_12897));
OAI21X1 g122283(.A0 (n_12599), .A1 (n_27698), .B0 (n_12894), .Y(n_12895));
OAI21X1 g122294(.A0 (n_12609), .A1 (n_29285), .B0 (n_12892), .Y(n_12893));
OAI21X1 g122303(.A0 (n_12613), .A1 (n_29285), .B0 (n_12890), .Y(n_12891));
OAI21X1 g122306(.A0 (n_12602), .A1 (n_34375), .B0 (n_12888), .Y(n_12889));
OAI21X1 g122307(.A0 (n_12603), .A1 (n_27698), .B0 (n_12886), .Y(n_12887));
OAI21X1 g122308(.A0 (n_12607), .A1 (n_27698), .B0 (n_12883), .Y(n_12885));
OAI21X1 g122309(.A0 (n_12614), .A1 (n_33201), .B0 (n_12881), .Y(n_12882));
OAI21X1 g122310(.A0 (n_12598), .A1 (n_33201), .B0 (n_12879), .Y(n_12880));
OAI21X1 g122312(.A0 (n_12600), .A1 (n_27698), .B0 (n_12877), .Y(n_12878));
OAI21X1 g122313(.A0 (n_12612), .A1 (n_27698), .B0 (n_12875), .Y(n_12876));
OAI21X1 g122314(.A0 (n_12596), .A1 (n_33201), .B0 (n_12873), .Y(n_12874));
OAI21X1 g122316(.A0 (n_12605), .A1 (n_33201), .B0 (n_12871), .Y(n_12872));
AOI22X1 g122329(.A0 (n_33290), .A1 (n_12594), .B0 (n_10706), .B1(n_32827), .Y (n_14817));
AOI22X1 g122345(.A0 (n_13075), .A1 (n_12593), .B0 (n_9284), .B1(n_13408), .Y (n_14344));
AOI22X1 g122354(.A0 (n_9720), .A1 (n_12792), .B0 (n_11797), .B1(n_12617), .Y (n_12869));
XOR2X1 g122361(.A (n_17471), .B (n_12788), .Y (n_12867));
NOR2X1 g122741(.A (n_11503), .B (n_12863), .Y (n_12865));
NAND3X1 g122742(.A (n_12766), .B (n_12851), .C (n_12314), .Y(n_12862));
NOR2X1 g122887(.A (n_12795), .B (n_12860), .Y (n_12861));
NAND2X1 g122973(.A (n_12671), .B (n_6950), .Y (n_12858));
NOR2X1 g123025(.A (n_12857), .B (n_12450), .Y (n_13101));
NAND2X1 g123101(.A (n_12682), .B (n_31528), .Y (n_12856));
MX2X1 g123137(.A (n_12586), .B (P3_d), .S0 (n_12389), .Y (n_12853));
XOR2X1 g123144(.A (n_11791), .B (n_12851), .Y (n_12852));
XOR2X1 g123145(.A (n_11092), .B (n_12768), .Y (n_12850));
XOR2X1 g123146(.A (n_17467), .B (n_12760), .Y (n_12848));
XOR2X1 g123147(.A (n_11556), .B (n_12591), .Y (n_12846));
XOR2X1 g123148(.A (n_17472), .B (n_12771), .Y (n_12845));
INVX1 g123168(.A (n_12843), .Y (n_12844));
INVX2 g123172(.A (n_12841), .Y (n_12840));
INVX1 g123542(.A (n_12839), .Y (n_13085));
NAND3X1 g123545(.A (n_34874), .B (n_34863), .C (n_34866), .Y(n_12838));
AND2X1 g123692(.A (n_12835), .B (n_12834), .Y (n_12836));
AOI21X1 g123774(.A0 (n_11360), .A1 (n_8916), .B0 (n_12665), .Y(n_12832));
AOI21X1 g123775(.A0 (n_11357), .A1 (n_12664), .B0 (n_12663), .Y(n_12831));
INVX1 g123800(.A (n_12830), .Y (n_12923));
AOI22X1 g123823(.A0 (n_9730), .A1 (n_12667), .B0 (n_12827), .B1(n_12428), .Y (n_12829));
NAND3X1 g123944(.A (n_12804), .B (n_12566), .C (n_12121), .Y(n_12826));
NAND2X1 g123945(.A (n_12651), .B (n_12824), .Y (n_12825));
NAND2X1 g123946(.A (n_12650), .B (n_12822), .Y (n_12823));
NAND2X1 g123947(.A (n_12647), .B (n_12820), .Y (n_12821));
NAND2X1 g123951(.A (n_12645), .B (n_12818), .Y (n_12819));
NAND2X1 g123952(.A (n_12636), .B (n_12816), .Y (n_12817));
NAND2X1 g123962(.A (n_12642), .B (n_12814), .Y (n_12815));
NAND2X1 g123965(.A (n_12643), .B (n_12812), .Y (n_12813));
NAND2X1 g123966(.A (n_12640), .B (n_12810), .Y (n_12811));
NAND2X1 g123969(.A (n_12644), .B (n_12808), .Y (n_12809));
NAND2X1 g123970(.A (n_12646), .B (n_12806), .Y (n_12807));
NAND3X1 g123972(.A (n_12804), .B (n_12566), .C (n_12122), .Y(n_12805));
XOR2X1 g123997(.A (n_35318), .B (n_12568), .Y (n_12803));
INVX1 g124000(.A (n_12801), .Y (n_12802));
NAND2X1 g124002(.A (n_12452), .B (n_12799), .Y (n_12800));
INVX1 g124243(.A (n_12905), .Y (n_12798));
CLKBUFX1 gbuf_d_544(.A(n_12622), .Y(d_out_544));
CLKBUFX1 gbuf_q_544(.A(q_in_544), .Y(datao_2[27]));
NOR2X1 g124448(.A (n_12294), .B (n_12795), .Y (n_12796));
CLKBUFX1 gbuf_d_545(.A(n_12549), .Y(d_out_545));
CLKBUFX1 gbuf_q_545(.A(q_in_545), .Y(n_641));
CLKBUFX1 gbuf_d_546(.A(n_12556), .Y(d_out_546));
CLKBUFX1 gbuf_q_546(.A(q_in_546), .Y(datao_2[4]));
CLKBUFX1 gbuf_d_547(.A(n_12547), .Y(d_out_547));
CLKBUFX1 gbuf_q_547(.A(q_in_547), .Y(datao_1[28]));
CLKBUFX1 gbuf_d_548(.A(n_12570), .Y(d_out_548));
CLKBUFX1 gbuf_q_548(.A(q_in_548), .Y(P2_d_394));
CLKBUFX1 gbuf_d_549(.A(n_12557), .Y(d_out_549));
CLKBUFX1 gbuf_q_549(.A(q_in_549), .Y(datao_2[13]));
CLKBUFX1 gbuf_d_550(.A(n_12553), .Y(d_out_550));
CLKBUFX1 gbuf_q_550(.A(q_in_550), .Y(datao_2[21]));
AOI22X1 g123801(.A0 (n_8124), .A1 (n_12514), .B0 (n_17471), .B1(n_13408), .Y (n_12830));
NOR2X1 g121925(.A (n_12335), .B (n_12692), .Y (n_12899));
NAND3X1 g122057(.A (n_12783), .B (n_12792), .C (n_12791), .Y(n_12793));
NAND4X1 g122276(.A (n_12779), .B (n_12778), .C (n_12009), .D(n_12790), .Y (n_12976));
NAND4X1 g122327(.A (n_12788), .B (n_12776), .C (n_11530), .D(n_12787), .Y (n_12789));
INVX1 g122633(.A (n_12785), .Y (n_12786));
AND2X1 g122971(.A (n_12783), .B (n_12792), .Y (n_12784));
INVX1 g123026(.A (n_12781), .Y (n_12782));
NAND3X1 g123103(.A (n_12779), .B (n_12778), .C (n_12790), .Y(n_12780));
NAND3X1 g123104(.A (n_12788), .B (n_12776), .C (n_12787), .Y(n_12777));
INVX1 g123106(.A (n_14783), .Y (n_12775));
INVX1 g123109(.A (n_13918), .Y (n_12774));
NAND4X1 g123128(.A (n_12762), .B (n_12771), .C (n_12338), .D(n_12761), .Y (n_12772));
MX2X1 g123136(.A (P2_d), .B (n_12539), .S0 (n_12488), .Y (n_12770));
XOR2X1 g123143(.A (n_11790), .B (n_12685), .Y (n_12769));
NAND2X1 g123169(.A (n_34875), .B (n_11310), .Y (n_12843));
NAND2X2 g123173(.A (n_11308), .B (n_12768), .Y (n_12841));
NAND2X1 g123175(.A (n_12766), .B (n_12851), .Y (n_12767));
INVX1 g123537(.A (n_12764), .Y (n_12765));
NAND3X1 g123541(.A (n_12771), .B (n_12762), .C (n_12761), .Y(n_12763));
NAND2X1 g123543(.A (n_12760), .B (n_11539), .Y (n_12839));
NAND2X1 g123546(.A (n_12587), .B (n_12204), .Y (n_12942));
INVX1 g123765(.A (n_12860), .Y (n_12759));
INVX1 g123768(.A (n_33410), .Y (n_12938));
INVX1 g123769(.A (n_33410), .Y (n_12757));
NAND4X1 g123771(.A (n_12194), .B (n_13232), .C (n_11992), .D(n_12655), .Y (n_12939));
CLKBUFX1 gbuf_d_551(.A(n_12619), .Y(d_out_551));
CLKBUFX1 gbuf_q_551(.A(q_in_551), .Y(P1_d));
AOI22X1 g123793(.A0 (n_12535), .A1 (n_12739), .B0 (n_11391), .B1(n_12755), .Y (n_12756));
AOI22X1 g123794(.A0 (n_12528), .A1 (n_12753), .B0 (n_11372), .B1(n_12917), .Y (n_12754));
AOI22X1 g123795(.A0 (n_12531), .A1 (n_6354), .B0 (n_11386), .B1(n_10342), .Y (n_12752));
AOI22X1 g123796(.A0 (n_12530), .A1 (n_12739), .B0 (n_11374), .B1(n_12917), .Y (n_12751));
AOI22X1 g123802(.A0 (n_12520), .A1 (n_12739), .B0 (n_11378), .B1(n_6421), .Y (n_12750));
AOI22X1 g123803(.A0 (n_12523), .A1 (n_6354), .B0 (n_11384), .B1(n_10342), .Y (n_12749));
AOI22X1 g123804(.A0 (n_12527), .A1 (n_6354), .B0 (n_11388), .B1(n_12755), .Y (n_12746));
AOI22X1 g123805(.A0 (n_12522), .A1 (n_12753), .B0 (n_11382), .B1(n_6421), .Y (n_12744));
AOI22X1 g123806(.A0 (n_12521), .A1 (n_12753), .B0 (n_11380), .B1(n_12755), .Y (n_12742));
AOI22X1 g123807(.A0 (n_12519), .A1 (n_6354), .B0 (n_11376), .B1(n_10342), .Y (n_12741));
AOI22X1 g123811(.A0 (n_12518), .A1 (n_12739), .B0 (n_11370), .B1(n_12755), .Y (n_12740));
AOI22X1 g123812(.A0 (n_12525), .A1 (n_12739), .B0 (n_11366), .B1(n_12755), .Y (n_12738));
AOI22X1 g123813(.A0 (n_12526), .A1 (n_12739), .B0 (n_11364), .B1(n_12755), .Y (n_12737));
AOI22X1 g123814(.A0 (n_12516), .A1 (n_12739), .B0 (n_11362), .B1(n_10342), .Y (n_12736));
AOI22X1 g123815(.A0 (n_12517), .A1 (n_12739), .B0 (n_11368), .B1(n_6421), .Y (n_12735));
NOR2X1 g123941(.A (n_12585), .B (n_12926), .Y (n_12734));
NAND2X1 g123942(.A (n_12574), .B (n_12732), .Y (n_12733));
NAND2X1 g123948(.A (n_12580), .B (n_12730), .Y (n_12731));
NAND2X1 g123949(.A (n_12579), .B (n_12728), .Y (n_12729));
INVX1 g123954(.A (n_12725), .Y (n_12726));
NAND2X1 g123956(.A (n_12577), .B (n_12723), .Y (n_12724));
NOR2X1 g123959(.A (n_12334), .B (n_12721), .Y (n_12722));
NAND3X1 g123960(.A (n_16182), .B (n_16768), .C (n_12705), .Y(n_12720));
NAND2X1 g123963(.A (n_12576), .B (n_12718), .Y (n_12719));
NAND2X1 g123964(.A (n_12581), .B (n_12716), .Y (n_12717));
NAND2X1 g123967(.A (n_12575), .B (n_12714), .Y (n_12715));
NAND2X1 g123968(.A (n_12578), .B (n_12712), .Y (n_12713));
INVX1 g123975(.A (n_34982), .Y (n_12711));
NOR2X1 g123977(.A (n_32011), .B (n_12707), .Y (n_13053));
INVX1 g123978(.A (n_34413), .Y (n_12709));
NOR2X1 g123981(.A (n_12707), .B (n_12376), .Y (n_13067));
XOR2X1 g123992(.A (n_11285), .B (n_12705), .Y (n_12706));
XOR2X1 g123999(.A (n_12703), .B (n_12653), .Y (n_12704));
NOR2X1 g124001(.A (n_12702), .B (n_12632), .Y (n_12801));
NOR2X1 g124007(.A (n_11500), .B (n_12630), .Y (n_12701));
INVX1 g124058(.A (n_13913), .Y (n_12700));
XOR2X1 g124094(.A (n_10482), .B (n_12626), .Y (n_12698));
XOR2X1 g124097(.A (n_11275), .B (n_12628), .Y (n_12697));
NAND2X1 g124245(.A (n_12564), .B (n_11333), .Y (n_12905));
CLKBUFX1 gbuf_d_552(.A(n_12555), .Y(d_out_552));
CLKBUFX1 gbuf_q_552(.A(q_in_552), .Y(n_667));
NOR2X1 g124498(.A (n_12695), .B (n_10320), .Y (n_12696));
CLKBUFX1 gbuf_d_553(.A(n_12551), .Y(d_out_553));
CLKBUFX1 gbuf_q_553(.A(q_in_553), .Y(datao_2[16]));
MX2X1 g125265(.A (datao_2[26] ), .B (n_12546), .S0 (n_12464), .Y(n_12694));
CLKBUFX1 gbuf_d_554(.A(n_12466), .Y(d_out_554));
CLKBUFX1 gbuf_q_554(.A(q_in_554), .Y(datao_2[29]));
CLKBUFX1 gbuf_d_555(.A(n_12484), .Y(d_out_555));
CLKBUFX1 gbuf_q_555(.A(q_in_555), .Y(P2_d_393));
CLKBUFX1 gbuf_d_556(.A(n_12494), .Y(d_out_556));
CLKBUFX1 gbuf_q_556(.A(q_in_556), .Y(P2_d_390));
CLKBUFX1 gbuf_d_557(.A(n_12461), .Y(d_out_557));
CLKBUFX1 gbuf_q_557(.A(q_in_557), .Y(datao_2[10]));
CLKBUFX1 gbuf_d_558(.A(n_12487), .Y(d_out_558));
CLKBUFX1 gbuf_q_558(.A(q_in_558), .Y(P2_d_384));
CLKBUFX1 gbuf_d_559(.A(n_12479), .Y(d_out_559));
CLKBUFX1 gbuf_q_559(.A(q_in_559), .Y(P2_d_382));
CLKBUFX1 gbuf_d_560(.A(n_12500), .Y(d_out_560));
CLKBUFX1 gbuf_q_560(.A(q_in_560), .Y(P3_d_393));
CLKBUFX1 gbuf_d_561(.A(n_12493), .Y(d_out_561));
CLKBUFX1 gbuf_q_561(.A(q_in_561), .Y(P3_d_377));
CLKBUFX1 gbuf_d_562(.A(n_12511), .Y(d_out_562));
CLKBUFX1 gbuf_q_562(.A(q_in_562), .Y(P1_d_98));
CLKBUFX1 gbuf_d_563(.A(n_12462), .Y(d_out_563));
CLKBUFX1 gbuf_q_563(.A(q_in_563), .Y(datao_2[17]));
CLKBUFX1 gbuf_d_564(.A(n_12470), .Y(d_out_564));
CLKBUFX1 gbuf_q_564(.A(q_in_564), .Y(P2_d_388));
CLKBUFX1 gbuf_d_565(.A(n_12495), .Y(d_out_565));
CLKBUFX1 gbuf_q_565(.A(q_in_565), .Y(P2_d_391));
CLKBUFX1 gbuf_d_566(.A(n_12492), .Y(d_out_566));
CLKBUFX1 gbuf_q_566(.A(q_in_566), .Y(P3_d_398));
CLKBUFX1 gbuf_d_567(.A(n_12475), .Y(d_out_567));
CLKBUFX1 gbuf_q_567(.A(q_in_567), .Y(P2_d_397));
CLKBUFX1 gbuf_d_568(.A(n_12503), .Y(d_out_568));
CLKBUFX1 gbuf_q_568(.A(q_in_568), .Y(P3_d_407));
CLKBUFX1 gbuf_d_569(.A(n_12510), .Y(d_out_569));
CLKBUFX1 gbuf_q_569(.A(q_in_569), .Y(P2_d_387));
CLKBUFX1 gbuf_d_570(.A(n_12502), .Y(d_out_570));
CLKBUFX1 gbuf_q_570(.A(q_in_570), .Y(P2_d_392));
CLKBUFX1 gbuf_d_571(.A(n_12486), .Y(d_out_571));
CLKBUFX1 gbuf_q_571(.A(q_in_571), .Y(P2_d_389));
CLKBUFX1 gbuf_d_572(.A(n_12508), .Y(d_out_572));
CLKBUFX1 gbuf_q_572(.A(q_in_572), .Y(P2_d_381));
CLKBUFX1 gbuf_d_573(.A(n_12504), .Y(d_out_573));
CLKBUFX1 gbuf_q_573(.A(q_in_573), .Y(P2_d_402));
CLKBUFX1 gbuf_d_574(.A(n_12482), .Y(d_out_574));
CLKBUFX1 gbuf_q_574(.A(q_in_574), .Y(P2_d_398));
CLKBUFX1 gbuf_d_575(.A(n_12483), .Y(d_out_575));
CLKBUFX1 gbuf_q_575(.A(q_in_575), .Y(P2_d_396));
CLKBUFX1 gbuf_d_576(.A(n_12459), .Y(d_out_576));
CLKBUFX1 gbuf_q_576(.A(q_in_576), .Y(n_12458));
CLKBUFX1 gbuf_d_577(.A(n_12456), .Y(d_out_577));
CLKBUFX1 gbuf_q_577(.A(q_in_577), .Y(datao_2[20]));
CLKBUFX1 gbuf_d_578(.A(n_12455), .Y(d_out_578));
CLKBUFX1 gbuf_q_578(.A(q_in_578), .Y(n_12454));
CLKBUFX1 gbuf_d_579(.A(n_12473), .Y(d_out_579));
CLKBUFX1 gbuf_q_579(.A(q_in_579), .Y(P2_d_404));
NAND3X1 g123955(.A (n_35288), .B (n_35289), .C (n_11705), .Y(n_12725));
CLKBUFX1 gbuf_d_580(.A(n_12505), .Y(d_out_580));
CLKBUFX1 gbuf_q_580(.A(q_in_580), .Y(P2_d_399));
CLKBUFX1 gbuf_d_581(.A(n_12457), .Y(d_out_581));
CLKBUFX1 gbuf_q_581(.A(q_in_581), .Y(datao_2[22]));
CLKBUFX1 gbuf_d_582(.A(n_12496), .Y(d_out_582));
CLKBUFX1 gbuf_q_582(.A(q_in_582), .Y(P2_d_408));
NAND2X1 g122634(.A (n_12616), .B (n_11541), .Y (n_12785));
CLKBUFX1 gbuf_d_583(.A(n_12489), .Y(d_out_583));
CLKBUFX1 gbuf_q_583(.A(q_in_583), .Y(P2_d_407));
CLKBUFX1 gbuf_d_584(.A(n_12507), .Y(d_out_584));
CLKBUFX1 gbuf_q_584(.A(q_in_584), .Y(P2_d_401));
CLKBUFX1 gbuf_d_585(.A(n_12471), .Y(d_out_585));
CLKBUFX1 gbuf_q_585(.A(q_in_585), .Y(P2_d_403));
CLKBUFX1 gbuf_d_586(.A(n_12476), .Y(d_out_586));
CLKBUFX1 gbuf_q_586(.A(q_in_586), .Y(P2_d_378));
CLKBUFX1 gbuf_d_587(.A(n_12481), .Y(d_out_587));
CLKBUFX1 gbuf_q_587(.A(q_in_587), .Y(P2_d_405));
INVX1 g122744(.A (n_12692), .Y (n_12693));
NAND2X1 g123027(.A (n_12615), .B (n_11553), .Y (n_12781));
AOI22X1 g123105(.A0 (n_13230), .A1 (n_12422), .B0 (n_32856), .B1(n_13112), .Y (n_14178));
AOI22X1 g123107(.A0 (n_33290), .A1 (n_12425), .B0 (n_33268), .B1(n_32827), .Y (n_14783));
MX2X1 g123108(.A (n_1054), .B (n_12435), .S0 (n_11916), .Y (n_12691));
OAI22X1 g123111(.A0 (n_33094), .A1 (n_12419), .B0 (n_9219), .B1(n_12690), .Y (n_13918));
XOR2X1 g123139(.A (n_12289), .B (n_12432), .Y (n_12689));
XOR2X1 g123140(.A (n_10331), .B (n_12434), .Y (n_12688));
NAND2X1 g123170(.A (n_12592), .B (n_12001), .Y (n_12866));
NAND3X1 g123174(.A (n_12668), .B (n_12667), .C (n_12625), .Y(n_12863));
INVX1 g123538(.A (n_12779), .Y (n_12764));
NAND2X1 g123547(.A (n_12540), .B (n_31774), .Y (n_12687));
NAND2X1 g123616(.A (n_12589), .B (n_11779), .Y (n_12857));
NAND4X1 g123619(.A (n_12559), .B (n_12333), .C (n_12004), .D(n_12582), .Y (n_12686));
NAND2X1 g123766(.A (n_12685), .B (n_12180), .Y (n_12860));
AOI21X1 g123772(.A0 (n_10943), .A1 (n_35012), .B0 (n_12542), .Y(n_12684));
AOI21X1 g123773(.A0 (n_10973), .A1 (n_35012), .B0 (n_12543), .Y(n_12683));
AOI22X1 g123784(.A0 (n_12429), .A1 (n_8400), .B0 (n_31420), .B1(n_8413), .Y (n_12682));
AOI22X1 g123816(.A0 (n_12414), .A1 (n_12611), .B0 (n_11155), .B1(n_12678), .Y (n_12681));
AOI22X1 g123817(.A0 (n_12417), .A1 (n_12611), .B0 (n_11157), .B1(n_12678), .Y (n_12680));
AOI22X1 g123818(.A0 (n_12423), .A1 (n_12611), .B0 (n_11151), .B1(n_12678), .Y (n_12677));
AOI22X1 g123819(.A0 (n_12424), .A1 (n_12611), .B0 (n_11160), .B1(n_12678), .Y (n_12676));
AOI22X1 g123820(.A0 (n_12415), .A1 (n_12611), .B0 (n_11153), .B1(n_9937), .Y (n_12675));
MX2X1 g123824(.A (n_8687), .B (n_12381), .S0 (n_9813), .Y (n_12674));
XOR2X1 g123826(.A (n_9628), .B (n_12588), .Y (n_12673));
XOR2X1 g123828(.A (n_9788), .B (n_34940), .Y (n_12672));
MX2X1 g123829(.A (n_12670), .B (n_12427), .S0 (n_7860), .Y (n_12671));
AND2X1 g123924(.A (n_12668), .B (n_12667), .Y (n_12669));
NOR2X1 g123927(.A (n_12661), .B (n_12124), .Y (n_12835));
AOI21X1 g123937(.A0 (n_12379), .A1 (n_12662), .B0 (n_12664), .Y(n_12665));
AOI21X1 g123938(.A0 (n_12378), .A1 (n_12662), .B0 (n_12664), .Y(n_12663));
NOR2X1 g123961(.A (n_12661), .B (n_12228), .Y (n_12937));
NOR2X1 g123980(.A (n_11299), .B (n_12538), .Y (n_12658));
AOI22X1 g123986(.A0 (n_12369), .A1 (n_7860), .B0 (n_9382), .B1(n_7209), .Y (n_12657));
XOR2X1 g123996(.A (n_11276), .B (n_12655), .Y (n_12656));
NAND3X1 g124013(.A (n_12653), .B (n_12343), .C (n_12035), .Y(n_12654));
AOI22X1 g124033(.A0 (n_12360), .A1 (n_12649), .B0 (n_11834), .B1(n_12648), .Y (n_12651));
AOI22X1 g124034(.A0 (n_12359), .A1 (n_12649), .B0 (n_11831), .B1(n_12648), .Y (n_12650));
AOI22X1 g124035(.A0 (n_12358), .A1 (n_12649), .B0 (n_11829), .B1(n_12648), .Y (n_12647));
AOI22X1 g124038(.A0 (n_12356), .A1 (n_12649), .B0 (n_11821), .B1(n_12648), .Y (n_12646));
AOI22X1 g124041(.A0 (n_12353), .A1 (n_12649), .B0 (n_11823), .B1(n_12648), .Y (n_12645));
AOI22X1 g124042(.A0 (n_12354), .A1 (n_12649), .B0 (n_11826), .B1(n_12648), .Y (n_12644));
AOI22X1 g124043(.A0 (n_12355), .A1 (n_12649), .B0 (n_11819), .B1(n_12648), .Y (n_12643));
AOI22X1 g124046(.A0 (n_12357), .A1 (n_12649), .B0 (n_11817), .B1(n_12648), .Y (n_12642));
OAI22X1 g124060(.A0 (n_33094), .A1 (n_12351), .B0 (n_9624), .B1(n_12690), .Y (n_13913));
MX2X1 g124071(.A (n_11734), .B (n_12364), .S0 (n_7970), .Y (n_12641));
AOI22X1 g124074(.A0 (n_12361), .A1 (n_12649), .B0 (n_11805), .B1(n_12648), .Y (n_12640));
MX2X1 g124082(.A (n_11513), .B (n_12365), .S0 (n_7970), .Y (n_12639));
MX2X1 g124083(.A (n_11489), .B (n_12363), .S0 (n_11916), .Y(n_12638));
AOI22X1 g124087(.A0 (n_12366), .A1 (n_12649), .B0 (n_11596), .B1(n_12648), .Y (n_12636));
MX2X1 g124092(.A (n_11488), .B (n_12362), .S0 (n_7970), .Y (n_12635));
INVX1 g124198(.A (n_12632), .Y (n_12633));
INVX1 g124201(.A (n_12630), .Y (n_12631));
NOR2X1 g124204(.A (n_12341), .B (n_12628), .Y (n_12629));
NOR2X1 g124206(.A (n_12628), .B (n_12340), .Y (n_12799));
NOR2X1 g124226(.A (n_12045), .B (n_12626), .Y (n_12627));
CLKBUFX1 gbuf_d_588(.A(n_12477), .Y(d_out_588));
CLKBUFX1 gbuf_q_588(.A(q_in_588), .Y(P2_d_386));
CLKBUFX1 gbuf_d_589(.A(n_12460), .Y(d_out_589));
CLKBUFX1 gbuf_q_589(.A(q_in_589), .Y(datao_2[3]));
CLKBUFX1 gbuf_d_590(.A(n_12480), .Y(d_out_590));
CLKBUFX1 gbuf_q_590(.A(q_in_590), .Y(P3_d_384));
NAND4X1 g124633(.A (n_12173), .B (n_11747), .C (n_12169), .D(n_12625), .Y (n_12795));
CLKBUFX1 gbuf_d_591(.A(n_12491), .Y(d_out_591));
CLKBUFX1 gbuf_q_591(.A(q_in_591), .Y(P3_d_406));
MX2X1 g125269(.A (datao_2[8] ), .B (n_12442), .S0 (n_12464), .Y(n_12624));
MX2X1 g125281(.A (datao_2[25] ), .B (n_12445), .S0 (n_12488), .Y(n_12623));
MX2X1 g125284(.A (datao_2[27] ), .B (n_12446), .S0 (n_12464), .Y(n_12622));
MX2X1 g125285(.A (n_491), .B (n_12443), .S0 (n_12488), .Y (n_12621));
CLKBUFX1 gbuf_d_592(.A(n_12498), .Y(d_out_592));
CLKBUFX1 gbuf_q_592(.A(q_in_592), .Y(P2_d_383));
CLKBUFX1 gbuf_d_593(.A(n_12329), .Y(d_out_593));
CLKBUFX1 gbuf_q_593(.A(q_in_593), .Y(datao_2[14]));
CLKBUFX1 gbuf_d_594(.A(n_12331), .Y(d_out_594));
CLKBUFX1 gbuf_q_594(.A(q_in_594), .Y(n_12330));
CLKBUFX1 gbuf_d_595(.A(n_12386), .Y(d_out_595));
CLKBUFX1 gbuf_q_595(.A(q_in_595), .Y(P2_d_395));
CLKBUFX1 gbuf_d_596(.A(n_12320), .Y(d_out_596));
CLKBUFX1 gbuf_q_596(.A(q_in_596), .Y(n_12319));
CLKBUFX1 gbuf_d_597(.A(n_12321), .Y(d_out_597));
CLKBUFX1 gbuf_q_597(.A(q_in_597), .Y(datao_1[24]));
CLKBUFX1 gbuf_d_598(.A(n_12402), .Y(d_out_598));
CLKBUFX1 gbuf_q_598(.A(q_in_598), .Y(P3_d_392));
CLKBUFX1 gbuf_d_599(.A(n_12393), .Y(d_out_599));
CLKBUFX1 gbuf_q_599(.A(q_in_599), .Y(P3_d_402));
CLKBUFX1 gbuf_d_600(.A(n_12394), .Y(d_out_600));
CLKBUFX1 gbuf_q_600(.A(q_in_600), .Y(P3_d_401));
CLKBUFX1 gbuf_d_601(.A(n_12332), .Y(d_out_601));
CLKBUFX1 gbuf_q_601(.A(q_in_601), .Y(datao_2[6]));
CLKBUFX1 gbuf_d_602(.A(n_12398), .Y(d_out_602));
CLKBUFX1 gbuf_q_602(.A(q_in_602), .Y(P3_d_394));
CLKBUFX1 gbuf_d_603(.A(n_12395), .Y(d_out_603));
CLKBUFX1 gbuf_q_603(.A(q_in_603), .Y(P3_d_397));
CLKBUFX1 gbuf_d_604(.A(n_12396), .Y(d_out_604));
CLKBUFX1 gbuf_q_604(.A(q_in_604), .Y(P3_d_396));
CLKBUFX1 gbuf_d_605(.A(n_12397), .Y(d_out_605));
CLKBUFX1 gbuf_q_605(.A(q_in_605), .Y(P3_d_395));
CLKBUFX1 gbuf_d_606(.A(n_12318), .Y(d_out_606));
CLKBUFX1 gbuf_q_606(.A(q_in_606), .Y(n_475));
CLKBUFX1 gbuf_d_607(.A(n_12410), .Y(d_out_607));
CLKBUFX1 gbuf_q_607(.A(q_in_607), .Y(P3_d_389));
CLKBUFX1 gbuf_d_608(.A(n_12385), .Y(d_out_608));
CLKBUFX1 gbuf_q_608(.A(q_in_608), .Y(P2_d_379));
CLKBUFX1 gbuf_d_609(.A(n_12328), .Y(d_out_609));
CLKBUFX1 gbuf_q_609(.A(q_in_609), .Y(datao_2[23]));
CLKBUFX1 gbuf_d_610(.A(n_12408), .Y(d_out_610));
CLKBUFX1 gbuf_q_610(.A(q_in_610), .Y(P3_d_387));
CLKBUFX1 gbuf_d_611(.A(n_12400), .Y(d_out_611));
CLKBUFX1 gbuf_q_611(.A(q_in_611), .Y(P3_d_388));
CLKBUFX1 gbuf_d_612(.A(n_12391), .Y(d_out_612));
CLKBUFX1 gbuf_q_612(.A(q_in_612), .Y(P3_d_404));
CLKBUFX1 gbuf_d_613(.A(n_12403), .Y(d_out_613));
CLKBUFX1 gbuf_q_613(.A(q_in_613), .Y(P3_d_379));
CLKBUFX1 gbuf_d_614(.A(n_12388), .Y(d_out_614));
CLKBUFX1 gbuf_q_614(.A(q_in_614), .Y(P2_d_385));
CLKBUFX1 gbuf_d_615(.A(n_12342), .Y(d_out_615));
CLKBUFX1 gbuf_q_615(.A(q_in_615), .Y(datao_1[30]));
CLKBUFX1 gbuf_d_616(.A(n_12325), .Y(d_out_616));
CLKBUFX1 gbuf_q_616(.A(q_in_616), .Y(n_693));
CLKBUFX1 gbuf_d_617(.A(n_12326), .Y(d_out_617));
CLKBUFX1 gbuf_q_617(.A(q_in_617), .Y(datao_1[7]));
CLKBUFX1 gbuf_d_618(.A(n_12323), .Y(d_out_618));
CLKBUFX1 gbuf_q_618(.A(q_in_618), .Y(n_12322));
CLKBUFX1 gbuf_d_619(.A(n_12405), .Y(d_out_619));
CLKBUFX1 gbuf_q_619(.A(q_in_619), .Y(P2_d_380));
CLKBUFX1 gbuf_d_620(.A(n_12407), .Y(d_out_620));
CLKBUFX1 gbuf_q_620(.A(q_in_620), .Y(P1_d_111));
CLKBUFX1 gbuf_d_621(.A(n_12383), .Y(d_out_621));
CLKBUFX1 gbuf_q_621(.A(q_in_621), .Y(P2_d_406));
CLKBUFX1 gbuf_d_622(.A(n_12412), .Y(d_out_622));
CLKBUFX1 gbuf_q_622(.A(q_in_622), .Y(P2_d_400));
NAND2X1 g122745(.A (n_12545), .B (n_12008), .Y (n_12692));
MX2X1 g123135(.A (P1_d), .B (n_12292), .S0 (n_6435), .Y (n_12619));
XOR2X1 g123138(.A (n_10317), .B (n_12291), .Y (n_12618));
INVX1 g123176(.A (n_12792), .Y (n_12617));
CLKBUFX1 g123539(.A (n_12616), .Y (n_12779));
CLKBUFX1 g123617(.A (n_12615), .Y (n_12788));
AOI22X1 g123776(.A0 (n_12284), .A1 (n_12597), .B0 (n_10953), .B1(n_12601), .Y (n_12614));
AOI22X1 g123779(.A0 (n_12278), .A1 (n_12611), .B0 (n_10948), .B1(n_12678), .Y (n_12613));
AOI22X1 g123780(.A0 (n_12279), .A1 (n_12611), .B0 (n_10986), .B1(n_12678), .Y (n_12612));
AOI22X1 g123781(.A0 (n_12276), .A1 (n_12606), .B0 (n_10977), .B1(n_9937), .Y (n_12609));
AOI22X1 g123782(.A0 (n_12272), .A1 (n_12606), .B0 (n_10946), .B1(n_12601), .Y (n_12607));
AOI22X1 g123783(.A0 (n_12270), .A1 (n_12611), .B0 (n_10983), .B1(n_12601), .Y (n_12605));
AOI22X1 g123785(.A0 (n_12273), .A1 (n_12611), .B0 (n_10960), .B1(n_12678), .Y (n_12603));
AOI22X1 g123786(.A0 (n_12274), .A1 (n_12611), .B0 (n_10951), .B1(n_12601), .Y (n_12602));
AOI22X1 g123787(.A0 (n_12271), .A1 (n_12611), .B0 (n_10969), .B1(n_12601), .Y (n_12600));
AOI22X1 g123788(.A0 (n_12285), .A1 (n_12611), .B0 (n_10967), .B1(n_12678), .Y (n_12599));
AOI22X1 g123790(.A0 (n_12283), .A1 (n_12597), .B0 (n_10962), .B1(n_12601), .Y (n_12598));
AOI22X1 g123791(.A0 (n_12281), .A1 (n_12606), .B0 (n_10979), .B1(n_12601), .Y (n_12596));
AOI22X1 g123792(.A0 (n_12280), .A1 (n_12611), .B0 (n_10981), .B1(n_12601), .Y (n_12595));
XOR2X1 g123822(.A (n_9292), .B (n_12288), .Y (n_12594));
XOR2X1 g123827(.A (n_17007), .B (n_12544), .Y (n_12593));
NOR2X1 g123926(.A (n_11793), .B (n_12536), .Y (n_12760));
CLKBUFX1 g123928(.A (n_12592), .Y (n_12851));
NOR2X1 g123931(.A (n_34940), .B (n_35113), .Y (n_12591));
CLKBUFX1 g123932(.A (n_12589), .Y (n_12771));
NOR2X1 g123936(.A (n_34940), .B (n_11569), .Y (n_12768));
NOR2X1 g123957(.A (n_34940), .B (n_12347), .Y (n_12587));
AOI21X1 g123985(.A0 (n_12124), .A1 (n_8484), .B0 (n_9309), .Y(n_12586));
NAND3X1 g124006(.A (n_12210), .B (n_12212), .C (n_12213), .Y(n_12707));
NOR2X1 g124012(.A (n_11710), .B (n_12368), .Y (n_12834));
AOI21X1 g124020(.A0 (n_12227), .A1 (n_7970), .B0 (n_11952), .Y(n_12585));
INVX1 g124028(.A (n_12582), .Y (n_12721));
AOI22X1 g124032(.A0 (n_12220), .A1 (n_12649), .B0 (n_11592), .B1(n_12648), .Y (n_12581));
AOI22X1 g124036(.A0 (n_12224), .A1 (n_12649), .B0 (n_11607), .B1(n_12648), .Y (n_12580));
AOI22X1 g124037(.A0 (n_12223), .A1 (n_12649), .B0 (n_11605), .B1(n_12648), .Y (n_12579));
AOI22X1 g124039(.A0 (n_12222), .A1 (n_12649), .B0 (n_11594), .B1(n_12648), .Y (n_12578));
AOI22X1 g124040(.A0 (n_12221), .A1 (n_12649), .B0 (n_11599), .B1(n_12648), .Y (n_12577));
AOI22X1 g124044(.A0 (n_12218), .A1 (n_12649), .B0 (n_11588), .B1(n_12648), .Y (n_12576));
AOI22X1 g124045(.A0 (n_12225), .A1 (n_12649), .B0 (n_11601), .B1(n_12648), .Y (n_12575));
AOI22X1 g124047(.A0 (n_33290), .A1 (n_12209), .B0 (n_10669), .B1(n_32827), .Y (n_14508));
AOI22X1 g124048(.A0 (n_13393), .A1 (n_12207), .B0 (n_11759), .B1(n_13527), .Y (n_13895));
AOI22X1 g124072(.A0 (n_12226), .A1 (n_12649), .B0 (n_11584), .B1(n_12648), .Y (n_12574));
MX2X1 g124118(.A (P2_d_394), .B (n_12215), .S0 (n_12488), .Y(n_12570));
NAND2X1 g124199(.A (n_12468), .B (n_12044), .Y (n_12632));
NAND2X1 g124202(.A (n_12467), .B (n_12014), .Y (n_12630));
NOR2X1 g124222(.A (n_12344), .B (n_12512), .Y (n_12568));
INVX2 g124224(.A (n_12565), .Y (n_12566));
INVX2 g124228(.A (n_12469), .Y (n_12804));
NAND2X1 g124260(.A (n_12348), .B (n_12048), .Y (n_12564));
CLKBUFX1 gbuf_d_623(.A(n_12390), .Y(d_out_623));
CLKBUFX1 gbuf_q_623(.A(q_in_623), .Y(P3_d_382));
CLKBUFX1 gbuf_d_624(.A(n_12384), .Y(d_out_624));
CLKBUFX1 gbuf_q_624(.A(q_in_624), .Y(P3_d_383));
NOR2X1 g124478(.A (n_11731), .B (n_12562), .Y (n_12563));
AND2X1 g124802(.A (n_12336), .B (n_12311), .Y (n_12783));
NAND4X1 g124883(.A (n_12559), .B (n_17906), .C (n_12561), .D(n_12005), .Y (n_12695));
MX2X1 g125262(.A (datao_2[13] ), .B (n_12304), .S0 (n_12488), .Y(n_12557));
MX2X1 g125274(.A (datao_2[4] ), .B (n_12308), .S0 (n_12488), .Y(n_12556));
MX2X1 g125276(.A (n_667), .B (n_12309), .S0 (n_12464), .Y (n_12555));
MX2X1 g125277(.A (datao_2[21] ), .B (n_12305), .S0 (n_12488), .Y(n_12553));
MX2X1 g125287(.A (datao_2[16] ), .B (n_12310), .S0 (n_12488), .Y(n_12551));
CLKBUFX1 gbuf_d_625(.A(n_12404), .Y(d_out_625));
CLKBUFX1 gbuf_q_625(.A(q_in_625), .Y(P3_d_378));
MX2X1 g125411(.A (n_641), .B (n_12301), .S0 (n_6435), .Y (n_12549));
MX2X1 g125414(.A (datao_1[28] ), .B (n_12302), .S0 (n_12257), .Y(n_12547));
MX2X1 g126722(.A (n_11747), .B (datao_2[26] ), .S0 (n_8534), .Y(n_12546));
CLKBUFX1 gbuf_d_626(.A(n_12263), .Y(d_out_626));
CLKBUFX1 gbuf_q_626(.A(q_in_626), .Y(P1_d_115));
CLKBUFX1 gbuf_d_627(.A(n_12235), .Y(d_out_627));
CLKBUFX1 gbuf_q_627(.A(q_in_627), .Y(P3_d_380));
CLKBUFX1 gbuf_d_628(.A(n_12234), .Y(d_out_628));
CLKBUFX1 gbuf_q_628(.A(q_in_628), .Y(P3_d_381));
CLKBUFX1 gbuf_d_629(.A(n_12200), .Y(d_out_629));
CLKBUFX1 gbuf_q_629(.A(q_in_629), .Y(n_479));
CLKBUFX1 gbuf_d_630(.A(n_12261), .Y(d_out_630));
CLKBUFX1 gbuf_q_630(.A(q_in_630), .Y(P1_d_118));
CLKBUFX1 gbuf_d_631(.A(n_12185), .Y(d_out_631));
CLKBUFX1 gbuf_q_631(.A(q_in_631), .Y(n_12184));
CLKBUFX1 gbuf_d_632(.A(n_12262), .Y(d_out_632));
CLKBUFX1 gbuf_q_632(.A(q_in_632), .Y(P1_d_116));
CLKBUFX1 gbuf_d_633(.A(n_12187), .Y(d_out_633));
CLKBUFX1 gbuf_q_633(.A(q_in_633), .Y(datao_1[4]));
CLKBUFX1 gbuf_d_634(.A(n_12250), .Y(d_out_634));
CLKBUFX1 gbuf_q_634(.A(q_in_634), .Y(P1_d_125));
CLKBUFX1 gbuf_d_635(.A(n_12239), .Y(d_out_635));
CLKBUFX1 gbuf_q_635(.A(q_in_635), .Y(P3_d_400));
CLKBUFX1 gbuf_d_636(.A(n_12243), .Y(d_out_636));
CLKBUFX1 gbuf_q_636(.A(q_in_636), .Y(P3_d_399));
CLKBUFX1 gbuf_d_637(.A(n_12189), .Y(d_out_637));
CLKBUFX1 gbuf_q_637(.A(q_in_637), .Y(n_12188));
CLKBUFX1 gbuf_d_638(.A(n_12233), .Y(d_out_638));
CLKBUFX1 gbuf_q_638(.A(q_in_638), .Y(P3_d_391));
CLKBUFX1 gbuf_d_639(.A(n_12260), .Y(d_out_639));
CLKBUFX1 gbuf_q_639(.A(q_in_639), .Y(P1_d_117));
CLKBUFX1 gbuf_d_640(.A(n_12251), .Y(d_out_640));
CLKBUFX1 gbuf_q_640(.A(q_in_640), .Y(P1_d_124));
CLKBUFX1 gbuf_d_641(.A(n_12241), .Y(d_out_641));
CLKBUFX1 gbuf_q_641(.A(q_in_641), .Y(P3_d_386));
CLKBUFX1 gbuf_d_642(.A(n_12240), .Y(d_out_642));
CLKBUFX1 gbuf_q_642(.A(q_in_642), .Y(P3_d_390));
CLKBUFX1 gbuf_d_643(.A(n_12248), .Y(d_out_643));
CLKBUFX1 gbuf_q_643(.A(q_in_643), .Y(P1_d_101));
CLKBUFX1 gbuf_d_644(.A(n_12246), .Y(d_out_644));
CLKBUFX1 gbuf_q_644(.A(q_in_644), .Y(P1_d_126));
CLKBUFX1 gbuf_d_645(.A(n_12253), .Y(d_out_645));
CLKBUFX1 gbuf_q_645(.A(q_in_645), .Y(P1_d_123));
CLKBUFX1 gbuf_d_646(.A(n_12255), .Y(d_out_646));
CLKBUFX1 gbuf_q_646(.A(q_in_646), .Y(P1_d_122));
CLKBUFX1 gbuf_d_647(.A(n_12191), .Y(d_out_647));
CLKBUFX1 gbuf_q_647(.A(q_in_647), .Y(datao_2[15]));
CLKBUFX1 gbuf_d_648(.A(n_12186), .Y(d_out_648));
CLKBUFX1 gbuf_q_648(.A(q_in_648), .Y(n_804));
CLKBUFX1 gbuf_d_649(.A(n_12258), .Y(d_out_649));
CLKBUFX1 gbuf_q_649(.A(q_in_649), .Y(P1_d_119));
CLKBUFX1 gbuf_d_650(.A(n_12256), .Y(d_out_650));
CLKBUFX1 gbuf_q_650(.A(q_in_650), .Y(P1_d_120));
CLKBUFX1 gbuf_d_651(.A(n_12237), .Y(d_out_651));
CLKBUFX1 gbuf_q_651(.A(q_in_651), .Y(P3_d_403));
CLKBUFX1 gbuf_d_652(.A(n_12264), .Y(d_out_652));
CLKBUFX1 gbuf_q_652(.A(q_in_652), .Y(P1_d_112));
CLKBUFX1 gbuf_d_653(.A(n_12193), .Y(d_out_653));
CLKBUFX1 gbuf_q_653(.A(q_in_653), .Y(datao_2[7]));
NOR2X1 g123540(.A (n_11535), .B (n_12433), .Y (n_12616));
CLKBUFX1 gbuf_d_654(.A(n_12267), .Y(d_out_654));
CLKBUFX1 gbuf_q_654(.A(q_in_654), .Y(P1_d_109));
CLKBUFX1 gbuf_d_655(.A(n_12266), .Y(d_out_655));
CLKBUFX1 gbuf_q_655(.A(q_in_655), .Y(P1_d_110));
CLKBUFX1 gbuf_d_656(.A(n_12269), .Y(d_out_656));
CLKBUFX1 gbuf_q_656(.A(q_in_656), .Y(P1_d_107));
CLKBUFX1 gbuf_d_657(.A(n_12249), .Y(d_out_657));
CLKBUFX1 gbuf_q_657(.A(q_in_657), .Y(P1_d_100));
CLKBUFX1 g123177(.A (n_12545), .Y (n_12792));
NOR2X1 g123618(.A (n_11297), .B (n_12431), .Y (n_12615));
NOR2X1 g123925(.A (n_12428), .B (n_11996), .Y (n_12685));
INVX1 g123929(.A (n_12436), .Y (n_12592));
NOR2X1 g123933(.A (n_11077), .B (n_12544), .Y (n_12589));
AOI21X1 g123939(.A0 (n_9416), .A1 (n_12144), .B0 (n_9928), .Y(n_12543));
AOI21X1 g123940(.A0 (n_9415), .A1 (n_12126), .B0 (n_9928), .Y(n_12542));
AOI21X1 g123973(.A0 (n_6763), .A1 (n_8696), .B0 (n_12286), .Y(n_12540));
AOI21X1 g123984(.A0 (n_12121), .A1 (n_8400), .B0 (n_9828), .Y(n_12539));
INVX1 g124008(.A (n_12430), .Y (n_12659));
NAND3X1 g124014(.A (n_12078), .B (n_12103), .C (n_12101), .Y(n_12661));
AND2X1 g124017(.A (n_11633), .B (n_12367), .Y (n_12902));
NAND3X1 g124019(.A (n_35861), .B (n_12537), .C (n_11075), .Y(n_12538));
INVX1 g124029(.A (n_12536), .Y (n_12582));
MX2X1 g124065(.A (n_11725), .B (n_12108), .S0 (n_7970), .Y (n_12535));
AOI22X1 g124066(.A0 (n_33290), .A1 (n_12051), .B0 (n_15810), .B1(n_32827), .Y (n_14503));
AOI22X1 g124067(.A0 (n_13393), .A1 (n_12050), .B0 (n_12532), .B1(n_13527), .Y (n_14086));
MX2X1 g124068(.A (n_11740), .B (n_12112), .S0 (n_11916), .Y(n_12531));
MX2X1 g124069(.A (n_11737), .B (n_12104), .S0 (n_11916), .Y(n_12530));
MX2X1 g124070(.A (n_11736), .B (n_12115), .S0 (n_7970), .Y (n_12528));
MX2X1 g124073(.A (n_11478), .B (n_12113), .S0 (n_7970), .Y (n_12527));
MX2X1 g124075(.A (n_11506), .B (n_12106), .S0 (n_11916), .Y(n_12526));
MX2X1 g124076(.A (n_11491), .B (n_12114), .S0 (n_7970), .Y (n_12525));
MX2X1 g124077(.A (n_11497), .B (n_12111), .S0 (n_7970), .Y (n_12523));
MX2X1 g124078(.A (n_11496), .B (n_12110), .S0 (n_11916), .Y(n_12522));
MX2X1 g124079(.A (n_11495), .B (n_12117), .S0 (n_7970), .Y (n_12521));
MX2X1 g124080(.A (n_11493), .B (n_12118), .S0 (n_11916), .Y(n_12520));
MX2X1 g124081(.A (n_11492), .B (n_12109), .S0 (n_7970), .Y (n_12519));
MX2X1 g124084(.A (n_11487), .B (n_12107), .S0 (n_7970), .Y (n_12518));
MX2X1 g124085(.A (n_11957), .B (n_12105), .S0 (n_11916), .Y(n_12517));
MX2X1 g124086(.A (n_11486), .B (n_12116), .S0 (n_7970), .Y (n_12516));
INVX1 g124090(.A (n_12515), .Y (n_12572));
XOR2X1 g124100(.A (n_10315), .B (n_12512), .Y (n_12514));
MX2X1 g124117(.A (P1_d_98), .B (n_12100), .S0 (n_6435), .Y (n_12511));
MX2X1 g124122(.A (P2_d_387), .B (n_12075), .S0 (n_12464), .Y(n_12510));
MX2X1 g124129(.A (P2_d_381), .B (n_12093), .S0 (n_12488), .Y(n_12508));
MX2X1 g124134(.A (P2_d_401), .B (n_12071), .S0 (n_12464), .Y(n_12507));
CLKBUFX1 gbuf_d_658(.A(n_12242), .Y(d_out_658));
CLKBUFX1 gbuf_q_658(.A(q_in_658), .Y(P3_d_385));
MX2X1 g124138(.A (P2_d_399), .B (n_12086), .S0 (n_12488), .Y(n_12505));
MX2X1 g124142(.A (P2_d_402), .B (n_12063), .S0 (n_12464), .Y(n_12504));
MX2X1 g124144(.A (n_12077), .B (P3_d_407), .S0 (n_12389), .Y(n_12503));
MX2X1 g124146(.A (P2_d_392), .B (n_12066), .S0 (n_12464), .Y(n_12502));
MX2X1 g124147(.A (n_12079), .B (P3_d_393), .S0 (n_12389), .Y(n_12500));
MX2X1 g124149(.A (P2_d_383), .B (n_12094), .S0 (n_12488), .Y(n_12498));
MX2X1 g124150(.A (P2_d_408), .B (n_12062), .S0 (n_12464), .Y(n_12496));
MX2X1 g124152(.A (P2_d_391), .B (n_12087), .S0 (n_12488), .Y(n_12495));
MX2X1 g124154(.A (P2_d_390), .B (n_12070), .S0 (n_12464), .Y(n_12494));
MX2X1 g124161(.A (n_12097), .B (P3_d_377), .S0 (n_12389), .Y(n_12493));
MX2X1 g124164(.A (n_12060), .B (P3_d_398), .S0 (n_12389), .Y(n_12492));
MX2X1 g124171(.A (n_12068), .B (P3_d_406), .S0 (n_12389), .Y(n_12491));
MX2X1 g124175(.A (P2_d_407), .B (n_12069), .S0 (n_12488), .Y(n_12489));
MX2X1 g124177(.A (P2_d_384), .B (n_12084), .S0 (n_12488), .Y(n_12487));
MX2X1 g124181(.A (P2_d_389), .B (n_12057), .S0 (n_12464), .Y(n_12486));
MX2X1 g124182(.A (P2_d_393), .B (n_12089), .S0 (n_12464), .Y(n_12484));
MX2X1 g124183(.A (P2_d_396), .B (n_12091), .S0 (n_12464), .Y(n_12483));
MX2X1 g124184(.A (P2_d_398), .B (n_12064), .S0 (n_12464), .Y(n_12482));
MX2X1 g124185(.A (P2_d_405), .B (n_12090), .S0 (n_12464), .Y(n_12481));
MX2X1 g124187(.A (n_12073), .B (P3_d_384), .S0 (n_12389), .Y(n_12480));
MX2X1 g124188(.A (P2_d_382), .B (n_12096), .S0 (n_12464), .Y(n_12479));
MX2X1 g124189(.A (P2_d_386), .B (n_12061), .S0 (n_12464), .Y(n_12477));
MX2X1 g124190(.A (P2_d_378), .B (n_12099), .S0 (n_12488), .Y(n_12476));
MX2X1 g124191(.A (P2_d_397), .B (n_12082), .S0 (n_12464), .Y(n_12475));
MX2X1 g124193(.A (P2_d_404), .B (n_12083), .S0 (n_12488), .Y(n_12473));
MX2X1 g124194(.A (P2_d_403), .B (n_12081), .S0 (n_12488), .Y(n_12471));
MX2X1 g124196(.A (P2_d_388), .B (n_12056), .S0 (n_12488), .Y(n_12470));
NOR2X1 g124200(.A (n_12512), .B (n_12198), .Y (n_12653));
NOR2X1 g124219(.A (n_12352), .B (n_11572), .Y (n_12705));
NAND3X1 g124225(.A (n_12211), .B (n_11845), .C (n_12052), .Y(n_12565));
NAND3X1 g124229(.A (n_12217), .B (n_12053), .C (n_11874), .Y(n_12469));
INVX1 g124322(.A (n_12468), .Y (n_12626));
INVX1 g124325(.A (n_12467), .Y (n_12628));
CLKBUFX1 gbuf_d_659(.A(n_12190), .Y(d_out_659));
CLKBUFX1 gbuf_q_659(.A(q_in_659), .Y(datao_2[9]));
CLKBUFX1 gbuf_d_660(.A(n_12236), .Y(d_out_660));
CLKBUFX1 gbuf_q_660(.A(q_in_660), .Y(P3_d_405));
CLKBUFX1 gbuf_d_661(.A(n_12192), .Y(d_out_661));
CLKBUFX1 gbuf_q_661(.A(q_in_661), .Y(datao_2[18]));
NOR2X1 g124795(.A (n_34613), .B (n_12196), .Y (n_12766));
MX2X1 g124912(.A (datao_2[29] ), .B (n_12178), .S0 (n_12464), .Y(n_12466));
INVX1 g124982(.A (n_12339), .Y (n_32041));
NOR2X1 g125198(.A (n_12168), .B (n_12181), .Y (n_12668));
MX2X1 g125268(.A (datao_2[17] ), .B (n_12167), .S0 (n_12464), .Y(n_12462));
MX2X1 g125271(.A (datao_2[10] ), .B (n_12161), .S0 (n_12464), .Y(n_12461));
MX2X1 g125280(.A (datao_2[3] ), .B (n_12166), .S0 (n_12464), .Y(n_12460));
MX2X1 g125282(.A (n_12458), .B (n_12163), .S0 (n_12488), .Y(n_12459));
MX2X1 g125283(.A (datao_2[22] ), .B (n_12159), .S0 (n_12464), .Y(n_12457));
MX2X1 g125290(.A (datao_2[20] ), .B (n_12160), .S0 (n_12488), .Y(n_12456));
CLKBUFX1 gbuf_d_662(.A(n_12245), .Y(d_out_662));
CLKBUFX1 gbuf_q_662(.A(q_in_662), .Y(P1_d_105));
MX2X1 g125403(.A (n_12454), .B (n_12157), .S0 (n_6435), .Y (n_12455));
INVX1 g125473(.A (n_12451), .Y (n_12452));
NOR2X1 g125527(.A (n_11780), .B (n_12450), .Y (n_12762));
NOR2X1 g125553(.A (n_34873), .B (n_13095), .Y (n_12449));
CLKBUFX1 gbuf_d_663(.A(n_12247), .Y(d_out_663));
CLKBUFX1 gbuf_q_663(.A(q_in_663), .Y(P1_d_103));
CLKBUFX1 gbuf_d_664(.A(n_12137), .Y(d_out_664));
CLKBUFX1 gbuf_q_664(.A(q_in_664), .Y(P1_d_121));
MX2X1 g126716(.A (n_11716), .B (datao_2[27] ), .S0 (n_8534), .Y(n_12446));
MX2X1 g126724(.A (n_34609), .B (datao_2[25] ), .S0 (n_8534), .Y(n_12445));
MX2X1 g126730(.A (n_16796), .B (n_491), .S0 (n_8534), .Y (n_12443));
MX2X1 g126731(.A (n_11797), .B (datao_2[8] ), .S0 (n_8534), .Y(n_12442));
NAND2X1 g126793(.A (n_11747), .B (n_32827), .Y (n_35699));
CLKBUFX1 gbuf_d_665(.A(n_12042), .Y(d_out_665));
CLKBUFX1 gbuf_q_665(.A(q_in_665), .Y(datao_1[29]));
CLKBUFX1 gbuf_d_666(.A(n_12041), .Y(d_out_666));
CLKBUFX1 gbuf_q_666(.A(q_in_666), .Y(datao_1[31]));
CLKBUFX1 gbuf_d_667(.A(n_12021), .Y(d_out_667));
CLKBUFX1 gbuf_q_667(.A(q_in_667), .Y(datao_1[5]));
CLKBUFX1 gbuf_d_668(.A(n_12135), .Y(d_out_668));
CLKBUFX1 gbuf_q_668(.A(q_in_668), .Y(P1_d_128));
CLKBUFX1 gbuf_d_669(.A(n_12133), .Y(d_out_669));
CLKBUFX1 gbuf_q_669(.A(q_in_669), .Y(P1_d_102));
CLKBUFX1 gbuf_d_670(.A(n_12130), .Y(d_out_670));
CLKBUFX1 gbuf_q_670(.A(q_in_670), .Y(P1_d_99));
CLKBUFX1 gbuf_d_671(.A(n_12025), .Y(d_out_671));
CLKBUFX1 gbuf_q_671(.A(q_in_671), .Y(datao_1[27]));
CLKBUFX1 gbuf_d_672(.A(n_12033), .Y(d_out_672));
CLKBUFX1 gbuf_q_672(.A(q_in_672), .Y(datao_2[19]));
NAND2X1 g124882(.A (n_12015), .B (wr_3), .Y (wr));
CLKBUFX1 gbuf_d_673(.A(n_12043), .Y(d_out_673));
CLKBUFX1 gbuf_q_673(.A(q_in_673), .Y(datao_2[31]));
CLKBUFX1 gbuf_d_674(.A(n_12034), .Y(d_out_674));
CLKBUFX1 gbuf_q_674(.A(q_in_674), .Y(datao_2[5]));
CLKBUFX1 gbuf_d_675(.A(n_12018), .Y(d_out_675));
CLKBUFX1 gbuf_q_675(.A(q_in_675), .Y(datao_1[10]));
CLKBUFX1 gbuf_d_676(.A(n_12031), .Y(d_out_676));
CLKBUFX1 gbuf_q_676(.A(q_in_676), .Y(n_12030));
CLKBUFX1 gbuf_d_677(.A(n_12023), .Y(d_out_677));
CLKBUFX1 gbuf_q_677(.A(q_in_677), .Y(n_12022));
CLKBUFX1 gbuf_d_678(.A(n_12020), .Y(d_out_678));
CLKBUFX1 gbuf_q_678(.A(q_in_678), .Y(datao_1[9]));
AOI22X1 g124091(.A0 (n_13409), .A1 (n_11839), .B0 (n_12437), .B1(n_13408), .Y (n_12515));
CLKBUFX1 gbuf_d_679(.A(n_12138), .Y(d_out_679));
CLKBUFX1 gbuf_q_679(.A(q_in_679), .Y(P1_d_114));
CLKBUFX1 gbuf_d_680(.A(n_12139), .Y(d_out_680));
CLKBUFX1 gbuf_q_680(.A(q_in_680), .Y(P1_d_113));
CLKBUFX1 gbuf_d_681(.A(n_12128), .Y(d_out_681));
CLKBUFX1 gbuf_q_681(.A(q_in_681), .Y(P1_d_104));
CLKBUFX1 gbuf_d_682(.A(n_12027), .Y(d_out_682));
CLKBUFX1 gbuf_q_682(.A(q_in_682), .Y(n_12026));
CLKBUFX1 gbuf_d_683(.A(n_12141), .Y(d_out_683));
CLKBUFX1 gbuf_q_683(.A(q_in_683), .Y(P1_d_108));
NAND3X1 g124030(.A (n_10487), .B (n_12418), .C (n_11076), .Y(n_12536));
CLKBUFX1 gbuf_d_684(.A(n_12016), .Y(d_out_684));
CLKBUFX1 gbuf_q_684(.A(q_in_684), .Y(datao_1[19]));
CLKBUFX1 gbuf_d_685(.A(n_12029), .Y(d_out_685));
CLKBUFX1 gbuf_q_685(.A(q_in_685), .Y(n_12028));
NOR2X1 g123178(.A (n_11786), .B (n_12290), .Y (n_12545));
NAND2X1 g123930(.A (n_11529), .B (n_12287), .Y (n_12436));
AOI21X1 g123982(.A0 (n_11615), .A1 (n_27042), .B0 (n_12143), .Y(n_12435));
INVX1 g123988(.A (n_12433), .Y (n_12434));
INVX1 g123990(.A (n_12431), .Y (n_12432));
NAND3X1 g124009(.A (n_11882), .B (n_11884), .C (n_11883), .Y(n_12430));
NAND3X1 g124010(.A (n_35420), .B (n_11759), .C (n_12232), .Y(n_12588));
AOI21X1 g124018(.A0 (n_11925), .A1 (n_10635), .B0 (n_9937), .Y(n_12429));
INVX1 g124024(.A (n_12428), .Y (n_12667));
NAND4X1 g124031(.A (n_10800), .B (n_11926), .C (n_12426), .D(n_11393), .Y (n_12427));
XOR2X1 g124093(.A (n_11256), .B (n_11708), .Y (n_12425));
MX2X1 g124095(.A (n_8141), .B (n_11936), .S0 (n_9310), .Y (n_12424));
MX2X1 g124096(.A (n_8149), .B (n_11935), .S0 (n_9310), .Y (n_12423));
XOR2X1 g124098(.A (n_12232), .B (n_34938), .Y (n_12422));
XOR2X1 g124099(.A (n_16577), .B (n_12418), .Y (n_12419));
MX2X1 g124101(.A (n_8132), .B (n_11937), .S0 (n_9310), .Y (n_12417));
MX2X1 g124102(.A (n_8137), .B (n_11933), .S0 (n_9310), .Y (n_12415));
MX2X1 g124103(.A (n_8145), .B (n_11934), .S0 (n_9310), .Y (n_12414));
MX2X1 g124104(.A (P2_d_400), .B (n_11890), .S0 (n_12464), .Y(n_12412));
MX2X1 g124105(.A (n_11912), .B (P3_d_389), .S0 (n_12389), .Y(n_12410));
MX2X1 g124106(.A (n_11918), .B (P3_d_387), .S0 (n_12389), .Y(n_12408));
MX2X1 g124111(.A (P1_d_111), .B (n_11915), .S0 (n_12257), .Y(n_12407));
MX2X1 g124141(.A (P2_d_380), .B (n_11893), .S0 (n_12464), .Y(n_12405));
MX2X1 g124143(.A (n_11919), .B (P3_d_378), .S0 (n_12389), .Y(n_12404));
MX2X1 g124145(.A (n_11898), .B (P3_d_379), .S0 (n_12389), .Y(n_12403));
MX2X1 g124151(.A (n_11913), .B (P3_d_392), .S0 (n_12389), .Y(n_12402));
MX2X1 g124157(.A (n_11922), .B (P3_d_388), .S0 (n_12389), .Y(n_12400));
MX2X1 g124159(.A (n_11909), .B (P3_d_394), .S0 (n_12389), .Y(n_12398));
MX2X1 g124160(.A (n_11906), .B (P3_d_395), .S0 (n_12389), .Y(n_12397));
MX2X1 g124162(.A (n_11904), .B (P3_d_396), .S0 (n_12389), .Y(n_12396));
MX2X1 g124163(.A (n_11920), .B (P3_d_397), .S0 (n_12389), .Y(n_12395));
MX2X1 g124166(.A (n_11896), .B (P3_d_401), .S0 (n_12389), .Y(n_12394));
MX2X1 g124167(.A (n_11901), .B (P3_d_402), .S0 (n_12389), .Y(n_12393));
MX2X1 g124169(.A (n_11899), .B (P3_d_404), .S0 (n_12389), .Y(n_12391));
MX2X1 g124173(.A (n_11889), .B (P3_d_382), .S0 (n_12389), .Y(n_12390));
MX2X1 g124178(.A (P2_d_385), .B (n_11891), .S0 (n_12488), .Y(n_12388));
MX2X1 g124179(.A (P2_d_395), .B (n_11894), .S0 (n_12488), .Y(n_12386));
MX2X1 g124186(.A (P2_d_379), .B (n_11892), .S0 (n_12488), .Y(n_12385));
MX2X1 g124192(.A (n_11888), .B (P3_d_383), .S0 (n_12389), .Y(n_12384));
MX2X1 g124195(.A (P2_d_406), .B (n_11914), .S0 (n_12488), .Y(n_12383));
NAND4X1 g124197(.A (n_10625), .B (n_11928), .C (n_12380), .D(n_10123), .Y (n_12381));
NAND2X1 g124203(.A (n_12120), .B (n_7415), .Y (n_12379));
NAND2X1 g124205(.A (n_12119), .B (n_7415), .Y (n_12378));
NAND3X1 g124211(.A (n_12374), .B (n_12098), .C (n_12373), .Y(n_12376));
NAND3X1 g124213(.A (n_12374), .B (n_11396), .C (n_12373), .Y(n_32011));
INVX1 g124214(.A (n_34989), .Y (n_35288));
NOR2X1 g124220(.A (n_12512), .B (n_12039), .Y (n_12655));
AOI21X1 g124227(.A0 (n_11629), .A1 (n_11873), .B0 (n_12664), .Y(n_12369));
INVX1 g124231(.A (n_12367), .Y (n_12368));
NAND4X1 g124250(.A (n_11597), .B (n_11836), .C (n_11317), .D(n_10626), .Y (n_12366));
NAND4X1 g124256(.A (n_11188), .B (n_11815), .C (n_11099), .D(n_10918), .Y (n_12365));
NAND4X1 g124257(.A (n_11187), .B (n_11813), .C (n_11110), .D(n_10916), .Y (n_12364));
NAND4X1 g124258(.A (n_11186), .B (n_11810), .C (n_11109), .D(n_10915), .Y (n_12363));
NAND4X1 g124259(.A (n_11185), .B (n_11808), .C (n_11105), .D(n_10914), .Y (n_12362));
NAND4X1 g124261(.A (n_11587), .B (n_11806), .C (n_11318), .D(n_10637), .Y (n_12361));
NAND3X1 g124278(.A (n_11613), .B (n_11835), .C (n_10907), .Y(n_12360));
NAND3X1 g124280(.A (n_11611), .B (n_11833), .C (n_10934), .Y(n_12359));
NAND3X1 g124281(.A (n_11609), .B (n_11830), .C (n_10933), .Y(n_12358));
NAND3X1 g124286(.A (n_11590), .B (n_11818), .C (n_10923), .Y(n_12357));
NAND3X1 g124293(.A (n_11598), .B (n_11822), .C (n_10929), .Y(n_12356));
NAND3X1 g124297(.A (n_11614), .B (n_11820), .C (n_10908), .Y(n_12355));
NAND3X1 g124313(.A (n_11604), .B (n_11827), .C (n_10921), .Y(n_12354));
NAND3X1 g124320(.A (n_11591), .B (n_11824), .C (n_10912), .Y(n_12353));
INVX1 g124323(.A (n_12352), .Y (n_12468));
INVX1 g124326(.A (n_12216), .Y (n_12467));
AOI22X1 g124436(.A0 (n_9286), .A1 (n_11617), .B0 (n_9761), .B1(n_11837), .Y (n_12351));
NAND2X1 g124447(.A (n_12349), .B (n_16732), .Y (n_12350));
NAND3X1 g124487(.A (n_11568), .B (n_12047), .C (n_11269), .Y(n_12348));
OR4X1 g124610(.A (n_11250), .B (n_12347), .C (n_34869), .D (n_12046),.Y (n_12562));
CLKBUFX1 gbuf_d_686(.A(n_12136), .Y(d_out_686));
CLKBUFX1 gbuf_q_686(.A(q_in_686), .Y(P1_d_127));
NAND2X1 g124838(.A (n_12197), .B (n_12343), .Y (n_12344));
MX2X1 g124917(.A (datao_1[30] ), .B (n_11999), .S0 (n_6435), .Y(n_12342));
OR2X1 g124958(.A (n_12340), .B (n_12313), .Y (n_12341));
NAND3X1 g124983(.A (n_12761), .B (n_12338), .C (n_12337), .Y(n_12339));
CLKBUFX1 gbuf_d_687(.A(n_12131), .Y(d_out_687));
CLKBUFX1 gbuf_q_687(.A(q_in_687), .Y(P1_d_106));
NOR2X1 g125126(.A (n_12007), .B (n_12335), .Y (n_12336));
NAND2X1 g125142(.A (n_12333), .B (n_12559), .Y (n_12334));
MX2X1 g125263(.A (datao_2[6] ), .B (n_11981), .S0 (n_12488), .Y(n_12332));
MX2X1 g125267(.A (n_12330), .B (n_11985), .S0 (n_12464), .Y(n_12331));
MX2X1 g125275(.A (datao_2[14] ), .B (n_11978), .S0 (n_12464), .Y(n_12329));
MX2X1 g125288(.A (datao_2[23] ), .B (n_11982), .S0 (n_12488), .Y(n_12328));
MX2X1 g125397(.A (datao_1[7] ), .B (n_11968), .S0 (n_6435), .Y(n_12326));
MX2X1 g125404(.A (n_693), .B (n_11976), .S0 (n_6435), .Y (n_12325));
MX2X1 g125406(.A (n_12322), .B (n_11973), .S0 (n_6435), .Y (n_12323));
MX2X1 g125410(.A (datao_1[24] ), .B (n_11971), .S0 (n_6435), .Y(n_12321));
MX2X1 g125412(.A (n_12319), .B (n_11970), .S0 (n_6435), .Y (n_12320));
MX2X1 g125424(.A (n_475), .B (n_11977), .S0 (n_6435), .Y (n_12318));
OR2X1 g125474(.A (n_12313), .B (n_12176), .Y (n_12451));
AND2X1 g125511(.A (n_12171), .B (n_12311), .Y (n_12312));
NAND2X1 g126087(.A (n_11066), .B (n_11954), .Y (n_12450));
MX2X1 g126706(.A (n_11713), .B (datao_2[16] ), .S0 (n_8534), .Y(n_12310));
MX2X1 g126712(.A (n_11732), .B (n_667), .S0 (n_8534), .Y (n_12309));
MX2X1 g126713(.A (n_10669), .B (datao_2[4] ), .S0 (n_8534), .Y(n_12308));
MX2X1 g126717(.A (n_11988), .B (datao_2[21] ), .S0 (n_8534), .Y(n_12305));
MX2X1 g126720(.A (n_12002), .B (datao_2[13] ), .S0 (n_8534), .Y(n_12304));
MX2X1 g126749(.A (n_11730), .B (datao_1[28] ), .S0 (n_7871), .Y(n_12302));
OAI21X1 g126756(.A0 (n_16442), .A1 (n_7860), .B0 (n_8537), .Y(n_12301));
NAND2X1 g126808(.A (n_34609), .B (n_32827), .Y (n_12299));
NAND2X1 g126825(.A (n_16796), .B (n_32827), .Y (n_12297));
NAND2X1 g126880(.A (n_16796), .B (n_11716), .Y (n_12294));
NAND2X1 g126968(.A (n_12561), .B (n_13106), .Y (n_35435));
CLKBUFX1 gbuf_d_688(.A(n_11799), .Y(d_out_688));
CLKBUFX1 gbuf_q_688(.A(q_in_688), .Y(datao_1[23]));
CLKBUFX1 gbuf_d_689(.A(n_11801), .Y(d_out_689));
CLKBUFX1 gbuf_q_689(.A(q_in_689), .Y(datao_1[0]));
NAND3X1 g124324(.A (n_11062), .B (n_12206), .C (n_11536), .Y(n_12352));
CLKBUFX1 gbuf_d_690(.A(n_11804), .Y(d_out_690));
CLKBUFX1 gbuf_q_690(.A(q_in_690), .Y(datao_2[1]));
CLKBUFX1 gbuf_d_691(.A(n_11800), .Y(d_out_691));
CLKBUFX1 gbuf_q_691(.A(q_in_691), .Y(n_928));
CLKBUFX1 gbuf_d_692(.A(n_11803), .Y(d_out_692));
CLKBUFX1 gbuf_q_692(.A(q_in_692), .Y(n_11802));
AOI21X1 g123983(.A0 (n_11705), .A1 (n_8557), .B0 (n_8560), .Y(n_12292));
INVX1 g123989(.A (n_12290), .Y (n_12291));
NAND3X1 g124005(.A (n_9284), .B (n_12289), .C (n_11880), .Y(n_12544));
INVX1 g124015(.A (n_12287), .Y (n_12288));
AOI21X1 g124021(.A0 (n_11616), .A1 (n_11685), .B0 (n_8505), .Y(n_12286));
NAND3X1 g124025(.A (n_11507), .B (n_12127), .C (n_11528), .Y(n_12428));
MX2X1 g124049(.A (n_7892), .B (n_11686), .S0 (n_9310), .Y (n_12285));
MX2X1 g124050(.A (n_8347), .B (n_11687), .S0 (n_9310), .Y (n_12284));
MX2X1 g124051(.A (n_7907), .B (n_11689), .S0 (n_9310), .Y (n_12283));
MX2X1 g124052(.A (n_7816), .B (n_11700), .S0 (n_9310), .Y (n_12281));
MX2X1 g124053(.A (n_7897), .B (n_11690), .S0 (n_9310), .Y (n_12280));
MX2X1 g124054(.A (n_7902), .B (n_11704), .S0 (n_9310), .Y (n_12279));
MX2X1 g124055(.A (n_7887), .B (n_11694), .S0 (n_9310), .Y (n_12278));
MX2X1 g124056(.A (n_7882), .B (n_11696), .S0 (n_9310), .Y (n_12276));
MX2X1 g124057(.A (n_8430), .B (n_11703), .S0 (n_9310), .Y (n_12274));
MX2X1 g124061(.A (n_8435), .B (n_11695), .S0 (n_9310), .Y (n_12273));
MX2X1 g124062(.A (n_8367), .B (n_11699), .S0 (n_9310), .Y (n_12272));
MX2X1 g124063(.A (n_8051), .B (n_11698), .S0 (n_9310), .Y (n_12271));
MX2X1 g124064(.A (n_7852), .B (n_11697), .S0 (n_9310), .Y (n_12270));
MX2X1 g124107(.A (P1_d_107), .B (n_11654), .S0 (n_6435), .Y(n_12269));
MX2X1 g124109(.A (P1_d_109), .B (n_11683), .S0 (n_12257), .Y(n_12267));
MX2X1 g124110(.A (P1_d_110), .B (n_11682), .S0 (n_6435), .Y(n_12266));
MX2X1 g124112(.A (P1_d_112), .B (n_11680), .S0 (n_12257), .Y(n_12264));
MX2X1 g124115(.A (P1_d_115), .B (n_11679), .S0 (n_6435), .Y(n_12263));
MX2X1 g124116(.A (P1_d_116), .B (n_11677), .S0 (n_6435), .Y(n_12262));
MX2X1 g124119(.A (P1_d_118), .B (n_11657), .S0 (n_12257), .Y(n_12261));
MX2X1 g124120(.A (P1_d_117), .B (n_11676), .S0 (n_6435), .Y(n_12260));
MX2X1 g124121(.A (P1_d_119), .B (n_11675), .S0 (n_12257), .Y(n_12258));
MX2X1 g124123(.A (P1_d_120), .B (n_11674), .S0 (n_12257), .Y(n_12256));
MX2X1 g124125(.A (P1_d_122), .B (n_11672), .S0 (n_12257), .Y(n_12255));
MX2X1 g124126(.A (P1_d_123), .B (n_11670), .S0 (n_6435), .Y(n_12253));
MX2X1 g124127(.A (P1_d_124), .B (n_11668), .S0 (n_6435), .Y(n_12251));
MX2X1 g124128(.A (P1_d_125), .B (n_11667), .S0 (n_6435), .Y(n_12250));
MX2X1 g124132(.A (P1_d_100), .B (n_11665), .S0 (n_6435), .Y(n_12249));
MX2X1 g124133(.A (P1_d_101), .B (n_11664), .S0 (n_6435), .Y(n_12248));
MX2X1 g124136(.A (P1_d_103), .B (n_11655), .S0 (n_12257), .Y(n_12247));
MX2X1 g124137(.A (P1_d_126), .B (n_11666), .S0 (n_12257), .Y(n_12246));
MX2X1 g124139(.A (P1_d_105), .B (n_11662), .S0 (n_12257), .Y(n_12245));
MX2X1 g124148(.A (n_11652), .B (P3_d_399), .S0 (n_12389), .Y(n_12243));
MX2X1 g124153(.A (n_11661), .B (P3_d_385), .S0 (n_12389), .Y(n_12242));
MX2X1 g124156(.A (n_11646), .B (P3_d_386), .S0 (n_12389), .Y(n_12241));
MX2X1 g124158(.A (n_11644), .B (P3_d_390), .S0 (n_12389), .Y(n_12240));
MX2X1 g124165(.A (n_11640), .B (P3_d_400), .S0 (n_12389), .Y(n_12239));
MX2X1 g124168(.A (n_11638), .B (P3_d_403), .S0 (n_12389), .Y(n_12237));
MX2X1 g124170(.A (n_11659), .B (P3_d_405), .S0 (n_12389), .Y(n_12236));
MX2X1 g124172(.A (n_11648), .B (P3_d_380), .S0 (n_12389), .Y(n_12235));
MX2X1 g124176(.A (n_11650), .B (P3_d_381), .S0 (n_12389), .Y(n_12234));
MX2X1 g124180(.A (n_11642), .B (P3_d_391), .S0 (n_12389), .Y(n_12233));
NAND2X1 g124218(.A (n_12232), .B (n_34938), .Y (n_12433));
NAND2X2 g124221(.A (n_12418), .B (n_9284), .Y (n_12431));
NOR2X1 g124232(.A (n_11932), .B (n_11693), .Y (n_12367));
NAND4X1 g124249(.A (n_10959), .B (n_11574), .C (n_10840), .D(n_10642), .Y (n_12227));
NAND4X1 g124254(.A (n_11585), .B (n_11576), .C (n_11321), .D(n_10647), .Y (n_12226));
NAND3X1 g124279(.A (n_11602), .B (n_11577), .C (n_10910), .Y(n_12225));
NAND3X1 g124282(.A (n_11608), .B (n_11582), .C (n_10931), .Y(n_12224));
NAND3X1 g124283(.A (n_11606), .B (n_11581), .C (n_10930), .Y(n_12223));
NAND3X1 g124285(.A (n_11595), .B (n_11583), .C (n_10919), .Y(n_12222));
NAND3X1 g124289(.A (n_11600), .B (n_11578), .C (n_10920), .Y(n_12221));
NAND3X1 g124298(.A (n_11593), .B (n_11579), .C (n_10909), .Y(n_12220));
NAND3X1 g124315(.A (n_11589), .B (n_11580), .C (n_10924), .Y(n_12218));
NOR2X1 g124321(.A (n_12214), .B (n_11877), .Y (n_12217));
NAND3X1 g124327(.A (n_11508), .B (n_12208), .C (n_11783), .Y(n_12216));
MX2X1 g124340(.A (P2_d_394), .B (n_12214), .S0 (n_8534), .Y(n_12215));
NOR2X1 g124425(.A (n_11625), .B (n_11842), .Y (n_12213));
NOR2X1 g124432(.A (n_11857), .B (n_11854), .Y (n_12212));
NOR2X1 g124433(.A (n_11860), .B (n_11851), .Y (n_12211));
NOR2X1 g124434(.A (n_11863), .B (n_11871), .Y (n_12210));
XOR2X1 g124435(.A (n_11249), .B (n_12208), .Y (n_12209));
XOR2X1 g124437(.A (n_11022), .B (n_12206), .Y (n_12207));
INVX1 g124624(.A (n_12349), .Y (n_12345));
INVX1 g124796(.A (n_12204), .Y (n_35113));
NOR3X1 g124831(.A (n_16442), .B (n_16174), .C (n_34862), .Y(n_12203));
MX2X1 g124911(.A (n_479), .B (n_11789), .S0 (n_12488), .Y (n_12200));
INVX1 g124930(.A (n_12197), .Y (n_12198));
OR2X1 g124954(.A (n_12000), .B (n_12195), .Y (n_12196));
INVX1 g125158(.A (n_12036), .Y (n_12194));
MX2X1 g125264(.A (datao_2[7] ), .B (n_11766), .S0 (n_12488), .Y(n_12193));
MX2X1 g125273(.A (datao_2[18] ), .B (n_11764), .S0 (n_12464), .Y(n_12192));
MX2X1 g125279(.A (datao_2[15] ), .B (n_11763), .S0 (n_12464), .Y(n_12191));
MX2X1 g125286(.A (datao_2[9] ), .B (n_11769), .S0 (n_12488), .Y(n_12190));
MX2X1 g125408(.A (n_12188), .B (n_11762), .S0 (n_6435), .Y (n_12189));
MX2X1 g125417(.A (datao_1[4] ), .B (n_11760), .S0 (n_12257), .Y(n_12187));
MX2X1 g125419(.A (n_804), .B (n_11756), .S0 (n_12257), .Y (n_12186));
MX2X1 g125420(.A (n_12184), .B (n_11752), .S0 (n_6435), .Y (n_12185));
NOR2X1 g125431(.A (n_12183), .B (n_10666), .Y (n_12791));
NOR2X1 g125448(.A (n_12183), .B (n_35245), .Y (n_12625));
NAND2X1 g125465(.A (n_11995), .B (n_12180), .Y (n_12181));
NOR2X1 g125538(.A (n_11997), .B (n_11294), .Y (n_35433));
MX2X1 g125938(.A (n_13114), .B (datao_2[29] ), .S0 (n_8534), .Y(n_12178));
OR2X1 g126030(.A (n_12175), .B (n_12174), .Y (n_12176));
NOR2X1 g126031(.A (n_10666), .B (n_12174), .Y (n_12173));
NOR2X1 g126032(.A (n_12174), .B (n_34612), .Y (n_12171));
NOR2X1 g126033(.A (n_11771), .B (n_11953), .Y (n_12559));
NOR2X1 g126700(.A (n_11733), .B (n_12175), .Y (n_12314));
INVX1 g126702(.A (n_12168), .Y (n_12169));
MX2X1 g126705(.A (n_32350), .B (datao_2[17] ), .S0 (n_8400), .Y(n_12167));
MX2X1 g126707(.A (n_10706), .B (datao_2[3] ), .S0 (n_8534), .Y(n_12166));
MX2X1 g126709(.A (n_11790), .B (n_12458), .S0 (n_8534), .Y (n_12163));
MX2X1 g126715(.A (n_11483), .B (datao_2[10] ), .S0 (n_8400), .Y(n_12161));
MX2X1 g126725(.A (n_11464), .B (datao_2[20] ), .S0 (n_8534), .Y(n_12160));
MX2X1 g126729(.A (n_16748), .B (datao_2[22] ), .S0 (n_8534), .Y(n_12159));
MX2X1 g126738(.A (n_19666), .B (n_12454), .S0 (n_7871), .Y (n_12157));
NAND2X1 g126764(.A (n_12002), .B (n_32827), .Y (n_12156));
NAND2X1 g126780(.A (n_11988), .B (n_32827), .Y (n_12154));
NAND2X1 g126801(.A (n_11730), .B (n_12953), .Y (n_12151));
NAND2X1 g126929(.A (n_11713), .B (n_32827), .Y (n_12147));
CLKBUFX1 gbuf_d_693(.A(n_11564), .Y(d_out_693));
CLKBUFX1 gbuf_q_693(.A(q_in_693), .Y(datao_2[2]));
CLKBUFX1 gbuf_d_694(.A(n_11561), .Y(d_out_694));
CLKBUFX1 gbuf_q_694(.A(q_in_694), .Y(n_732));
NOR3X1 g124016(.A (n_10451), .B (n_10317), .C (n_11708), .Y(n_12287));
NAND2X1 g124234(.A (n_11701), .B (n_9310), .Y (n_12144));
NAND4X1 g124011(.A (n_11190), .B (n_12142), .C (n_11198), .D(n_9997), .Y (n_12143));
MX2X1 g124108(.A (P1_d_108), .B (n_11453), .S0 (n_6435), .Y(n_12141));
MX2X1 g124113(.A (P1_d_113), .B (n_11452), .S0 (n_6435), .Y(n_12139));
MX2X1 g124114(.A (P1_d_114), .B (n_11451), .S0 (n_6435), .Y(n_12138));
MX2X1 g124124(.A (P1_d_121), .B (n_11449), .S0 (n_12257), .Y(n_12137));
MX2X1 g124130(.A (P1_d_127), .B (n_11446), .S0 (n_12257), .Y(n_12136));
MX2X1 g124131(.A (P1_d_128), .B (n_11441), .S0 (n_6435), .Y(n_12135));
MX2X1 g124135(.A (P1_d_102), .B (n_11445), .S0 (n_6435), .Y(n_12133));
MX2X1 g124140(.A (P1_d_106), .B (n_11442), .S0 (n_6435), .Y(n_12131));
MX2X1 g124155(.A (P1_d_99), .B (n_11448), .S0 (n_6435), .Y (n_12130));
MX2X1 g124174(.A (P1_d_104), .B (n_11443), .S0 (n_6435), .Y(n_12128));
CLKBUFX1 gbuf_d_695(.A(n_11563), .Y(d_out_695));
CLKBUFX1 gbuf_q_695(.A(q_in_695), .Y(datao_1[11]));
NAND2X1 g124212(.A (n_10706), .B (n_12127), .Y (n_12290));
NAND2X1 g124235(.A (n_11688), .B (n_9310), .Y (n_12126));
INVX1 g124238(.A (n_12124), .Y (n_12228));
INVX1 g124241(.A (n_12122), .Y (n_12121));
NAND4X1 g124253(.A (n_11361), .B (n_11395), .C (n_10575), .D(n_10628), .Y (n_12120));
NAND4X1 g124255(.A (n_11358), .B (n_11394), .C (n_10574), .D(n_10627), .Y (n_12119));
NAND3X1 g124262(.A (n_11379), .B (n_11359), .C (n_11179), .Y(n_12118));
NAND3X1 g124263(.A (n_11381), .B (n_11355), .C (n_11176), .Y(n_12117));
NAND3X1 g124264(.A (n_11363), .B (n_11352), .C (n_11173), .Y(n_12116));
NAND3X1 g124265(.A (n_11373), .B (n_11351), .C (n_11171), .Y(n_12115));
NAND3X1 g124266(.A (n_11367), .B (n_11348), .C (n_11170), .Y(n_12114));
NAND3X1 g124267(.A (n_11390), .B (n_11347), .C (n_11163), .Y(n_12113));
NAND3X1 g124268(.A (n_11387), .B (n_11349), .C (n_11178), .Y(n_12112));
NAND3X1 g124269(.A (n_11385), .B (n_11346), .C (n_11168), .Y(n_12111));
NAND3X1 g124270(.A (n_11383), .B (n_11345), .C (n_11167), .Y(n_12110));
NAND3X1 g124271(.A (n_11377), .B (n_11344), .C (n_11174), .Y(n_12109));
NAND3X1 g124272(.A (n_11392), .B (n_11342), .C (n_11166), .Y(n_12108));
NAND3X1 g124273(.A (n_11371), .B (n_11340), .C (n_11164), .Y(n_12107));
NAND3X1 g124274(.A (n_11365), .B (n_11350), .C (n_11169), .Y(n_12106));
NAND3X1 g124275(.A (n_11369), .B (n_11343), .C (n_11165), .Y(n_12105));
NAND3X1 g124276(.A (n_11375), .B (n_11341), .C (n_11162), .Y(n_12104));
NAND2X1 g124277(.A (n_11184), .B (n_11619), .Y (n_12537));
NOR2X1 g124292(.A (n_11636), .B (n_11658), .Y (n_12103));
NOR2X1 g124308(.A (n_11622), .B (n_11645), .Y (n_12101));
NAND3X1 g124328(.A (n_11045), .B (n_11617), .C (n_11305), .Y(n_12512));
AOI21X1 g124331(.A0 (n_11196), .A1 (n_7860), .B0 (n_8550), .Y(n_12100));
AOI21X1 g124332(.A0 (n_12098), .A1 (n_9310), .B0 (n_9816), .Y(n_12099));
MX2X1 g124333(.A (P3_d_377), .B (n_11192), .S0 (n_7970), .Y(n_12097));
AOI21X1 g124335(.A0 (n_11870), .A1 (n_8400), .B0 (n_9618), .Y(n_12096));
AOI21X1 g124336(.A0 (n_11859), .A1 (n_8400), .B0 (n_9815), .Y(n_12094));
AOI21X1 g124337(.A0 (n_11846), .A1 (n_8400), .B0 (n_9800), .Y(n_12093));
AOI21X1 g124339(.A0 (n_11844), .A1 (n_8400), .B0 (n_9811), .Y(n_12091));
AOI21X1 g124343(.A0 (n_11869), .A1 (n_8400), .B0 (n_9825), .Y(n_12090));
AOI21X1 g124371(.A0 (n_11868), .A1 (n_8400), .B0 (n_9833), .Y(n_12089));
AOI21X1 g124378(.A0 (n_12374), .A1 (n_8400), .B0 (n_9820), .Y(n_12087));
AOI21X1 g124380(.A0 (n_11856), .A1 (n_8400), .B0 (n_9819), .Y(n_12086));
AOI21X1 g124381(.A0 (n_11855), .A1 (n_8400), .B0 (n_9807), .Y(n_12084));
AOI21X1 g124382(.A0 (n_11843), .A1 (n_8400), .B0 (n_9806), .Y(n_12083));
AOI21X1 g124383(.A0 (n_11862), .A1 (n_8400), .B0 (n_9826), .Y(n_12082));
AOI21X1 g124384(.A0 (n_11841), .A1 (n_8400), .B0 (n_9804), .Y(n_12081));
AOI21X1 g124392(.A0 (n_12078), .A1 (n_8484), .B0 (n_9299), .Y(n_12079));
AOI21X1 g124400(.A0 (n_33330), .A1 (n_8484), .B0 (n_9719), .Y(n_12077));
AOI21X1 g124402(.A0 (n_11849), .A1 (n_8400), .B0 (n_9834), .Y(n_12075));
AOI21X1 g124403(.A0 (n_33333), .A1 (n_11916), .B0 (n_9718), .Y(n_12073));
AOI21X1 g124404(.A0 (n_11867), .A1 (n_8400), .B0 (n_9809), .Y(n_12071));
AOI21X1 g124405(.A0 (n_11840), .A1 (n_8400), .B0 (n_9617), .Y(n_12070));
AOI21X1 g124406(.A0 (n_11852), .A1 (n_8400), .B0 (n_9830), .Y(n_12069));
AOI21X1 g124408(.A0 (n_33331), .A1 (n_8484), .B0 (n_9758), .Y(n_12068));
AOI21X1 g124409(.A0 (n_11847), .A1 (n_8400), .B0 (n_9827), .Y(n_12066));
AOI21X1 g124411(.A0 (n_11850), .A1 (n_8400), .B0 (n_9835), .Y(n_12064));
AOI21X1 g124412(.A0 (n_11876), .A1 (n_8400), .B0 (n_9837), .Y(n_12063));
AOI21X1 g124413(.A0 (n_11864), .A1 (n_8400), .B0 (n_9832), .Y(n_12062));
AOI21X1 g124415(.A0 (n_11861), .A1 (n_8400), .B0 (n_9836), .Y(n_12061));
AOI21X1 g124416(.A0 (n_33332), .A1 (n_8484), .B0 (n_9230), .Y(n_12060));
AOI21X1 g124418(.A0 (n_11865), .A1 (n_8400), .B0 (n_9812), .Y(n_12057));
AOI21X1 g124423(.A0 (n_11853), .A1 (n_9310), .B0 (n_9801), .Y(n_12056));
NAND2X1 g124428(.A (n_11627), .B (n_11626), .Y (n_12055));
NAND2X1 g124445(.A (n_16778), .B (n_16735), .Y (n_12054));
INVX1 g124471(.A (n_11866), .Y (n_12053));
INVX1 g124482(.A (n_11848), .Y (n_12052));
XOR2X1 g124489(.A (n_11401), .B (n_32371), .Y (n_12051));
XOR2X1 g124491(.A (n_9780), .B (n_32944), .Y (n_12050));
NAND2X1 g124499(.A (n_11566), .B (n_13230), .Y (n_14147));
INVX1 g124598(.A (n_12049), .Y (n_14779));
AOI22X1 g124625(.A0 (n_10836), .A1 (n_11551), .B0 (n_11181), .B1(n_16452), .Y (n_12349));
CLKBUFX1 gbuf_d_696(.A(n_11565), .Y(d_out_696));
CLKBUFX1 gbuf_q_696(.A(q_in_696), .Y(datao_2[0]));
INVX1 g124793(.A (n_12047), .Y (n_12048));
NOR2X1 g124797(.A (n_12046), .B (n_11570), .Y (n_12204));
NAND2X1 g124864(.A (n_12044), .B (n_12006), .Y (n_12045));
MX2X1 g124913(.A (datao_2[31] ), .B (n_11550), .S0 (n_12488), .Y(n_12043));
MX2X1 g124916(.A (datao_1[29] ), .B (n_11549), .S0 (n_6435), .Y(n_12042));
MX2X1 g124918(.A (datao_1[31] ), .B (n_11546), .S0 (n_6435), .Y(n_12041));
NOR2X1 g124931(.A (n_12039), .B (n_11991), .Y (n_12197));
NOR2X1 g124936(.A (n_11552), .B (n_12038), .Y (n_12776));
NAND3X1 g125159(.A (n_12343), .B (n_12035), .C (n_12337), .Y(n_12036));
MX2X1 g125266(.A (datao_2[5] ), .B (n_11527), .S0 (n_12464), .Y(n_12034));
MX2X1 g125270(.A (datao_2[19] ), .B (n_11456), .S0 (n_12464), .Y(n_12033));
MX2X1 g125400(.A (n_12030), .B (n_11525), .S0 (n_6435), .Y (n_12031));
MX2X1 g125402(.A (n_12028), .B (n_11523), .S0 (n_6435), .Y (n_12029));
MX2X1 g125407(.A (n_12026), .B (n_11520), .S0 (n_6435), .Y (n_12027));
MX2X1 g125413(.A (datao_1[27] ), .B (n_11457), .S0 (n_6435), .Y(n_12025));
MX2X1 g125416(.A (n_12022), .B (n_11519), .S0 (n_6435), .Y (n_12023));
MX2X1 g125418(.A (datao_1[5] ), .B (n_11518), .S0 (n_6435), .Y(n_12021));
MX2X1 g125421(.A (datao_1[9] ), .B (n_11458), .S0 (n_6435), .Y(n_12020));
MX2X1 g125422(.A (datao_1[10] ), .B (n_11526), .S0 (n_6435), .Y(n_12018));
MX2X1 g125423(.A (datao_1[19] ), .B (n_11521), .S0 (n_12257), .Y(n_12016));
XOR2X1 g125425(.A (wr_1), .B (wr_2), .Y (n_12015));
NAND2X1 g125464(.A (n_12014), .B (n_12013), .Y (n_12340));
AND2X1 g125471(.A (n_11543), .B (n_12009), .Y (n_32221));
INVX1 g125490(.A (n_12007), .Y (n_12008));
NAND2X1 g125534(.A (n_12006), .B (n_11545), .Y (n_12702));
AND2X1 g125556(.A (n_12004), .B (n_11993), .Y (n_12005));
NAND3X1 g125573(.A (n_12003), .B (n_12002), .C (n_11994), .Y(n_12335));
INVX1 g125577(.A (n_12000), .Y (n_12001));
MX2X1 g125942(.A (n_18164), .B (datao_1[30] ), .S0 (n_7860), .Y(n_11999));
NAND2X1 g126029(.A (n_10470), .B (n_12337), .Y (n_11997));
INVX1 g126039(.A (n_11995), .Y (n_11996));
AND2X1 g126041(.A (n_11777), .B (n_11994), .Y (n_12180));
AND2X1 g126043(.A (n_11477), .B (n_11993), .Y (n_12338));
INVX1 g126055(.A (n_11991), .Y (n_11992));
OR2X1 g126082(.A (n_11990), .B (n_11989), .Y (n_12313));
NAND3X1 g126092(.A (n_16165), .B (n_16748), .C (n_11988), .Y(n_12183));
NAND4X1 g126703(.A (n_11987), .B (n_32350), .C (n_12003), .D(n_11278), .Y (n_12168));
MX2X1 g126704(.A (n_16895), .B (n_12330), .S0 (n_8400), .Y (n_11985));
MX2X1 g126710(.A (n_11503), .B (datao_2[23] ), .S0 (n_8534), .Y(n_11982));
MX2X1 g126728(.A (n_11249), .B (datao_2[6] ), .S0 (n_8534), .Y(n_11981));
MX2X1 g126732(.A (n_17261), .B (datao_2[14] ), .S0 (n_8534), .Y(n_11978));
MX2X1 g126739(.A (n_11034), .B (n_475), .S0 (n_7871), .Y (n_11977));
MX2X1 g126740(.A (n_11559), .B (n_693), .S0 (n_7871), .Y (n_11976));
MX2X1 g126742(.A (n_11555), .B (n_12322), .S0 (n_7871), .Y (n_11973));
MX2X1 g126746(.A (n_12977), .B (datao_1[24] ), .S0 (n_7871), .Y(n_11971));
MX2X1 g126747(.A (n_18496), .B (n_12319), .S0 (n_7871), .Y (n_11970));
MX2X1 g126754(.A (n_10330), .B (datao_1[7] ), .S0 (n_7871), .Y(n_11968));
NAND2X1 g126774(.A (n_16748), .B (n_32827), .Y (n_11966));
NAND2X1 g126799(.A (n_11483), .B (n_32827), .Y (n_11965));
NOR2X1 g126806(.A (n_34992), .B (n_11961), .Y (n_11962));
NAND2X1 g126948(.A (n_11033), .B (n_12953), .Y (n_11958));
AOI21X1 g126959(.A0 (n_9644), .A1 (n_11213), .B0 (n_11916), .Y(n_11957));
NAND2X1 g126969(.A (n_17909), .B (n_13106), .Y (n_32052));
NAND2X1 g126980(.A (n_11790), .B (n_32827), .Y (n_11955));
INVX1 g126982(.A (n_11953), .Y (n_11954));
AOI21X1 g127404(.A0 (n_11211), .A1 (n_10289), .B0 (n_7970), .Y(n_11952));
CLKBUFX1 gbuf_d_697(.A(n_11311), .Y(d_out_697));
CLKBUFX1 gbuf_q_697(.A(q_in_697), .Y(datao_1[1]));
NAND4X1 g124242(.A (n_7977), .B (n_11191), .C (n_10988), .D (n_7806),.Y (n_12122));
NOR3X1 g124207(.A (n_11939), .B (n_11196), .C (n_11938), .Y(n_11941));
NOR3X1 g124217(.A (n_11939), .B (n_10648), .C (n_11938), .Y(n_11940));
NOR2X1 g124239(.A (n_7973), .B (n_11454), .Y (n_12124));
NAND4X1 g124246(.A (n_10956), .B (n_11159), .C (n_10064), .D(n_10913), .Y (n_11937));
NAND4X1 g124247(.A (n_10972), .B (n_11161), .C (n_10052), .D(n_10906), .Y (n_11936));
NAND4X1 g124248(.A (n_10941), .B (n_11152), .C (n_10071), .D(n_10922), .Y (n_11935));
NAND4X1 g124251(.A (n_10976), .B (n_11156), .C (n_10061), .D(n_10926), .Y (n_11934));
NAND4X1 g124252(.A (n_10942), .B (n_11154), .C (n_10056), .D(n_10911), .Y (n_11933));
NAND3X1 g124303(.A (n_11649), .B (n_11660), .C (n_11903), .Y(n_11932));
NAND3X1 g124311(.A (n_11911), .B (n_11887), .C (n_11917), .Y(n_11931));
NAND3X1 g124317(.A (n_11897), .B (n_11908), .C (n_11900), .Y(n_11930));
NAND3X1 g124318(.A (n_11905), .B (n_11921), .C (n_11651), .Y(n_11929));
AOI21X1 g124329(.A0 (n_11923), .A1 (n_8687), .B0 (n_10631), .Y(n_11928));
AOI21X1 g124330(.A0 (n_11628), .A1 (n_12670), .B0 (n_10903), .Y(n_11926));
AOI22X1 g124334(.A0 (n_10623), .A1 (n_8413), .B0 (n_11923), .B1(n_8413), .Y (n_11925));
AOI21X1 g124338(.A0 (n_11921), .A1 (n_11916), .B0 (n_9791), .Y(n_11922));
AOI21X1 g124341(.A0 (n_11634), .A1 (n_11916), .B0 (n_9320), .Y(n_11920));
AOI21X1 g124342(.A0 (n_11620), .A1 (n_11916), .B0 (n_9321), .Y(n_11919));
AOI21X1 g124344(.A0 (n_11917), .A1 (n_11916), .B0 (n_9329), .Y(n_11918));
MX2X1 g124348(.A (P1_d_111), .B (n_11939), .S0 (n_7860), .Y(n_11915));
AOI21X1 g124376(.A0 (n_11858), .A1 (n_8400), .B0 (n_9818), .Y(n_11914));
AOI21X1 g124379(.A0 (n_11709), .A1 (n_11916), .B0 (n_9797), .Y(n_11913));
AOI21X1 g124386(.A0 (n_11911), .A1 (n_7970), .B0 (n_9704), .Y(n_11912));
AOI21X1 g124393(.A0 (n_11908), .A1 (n_8484), .B0 (n_9789), .Y(n_11909));
AOI21X1 g124394(.A0 (n_11905), .A1 (n_8484), .B0 (n_9699), .Y(n_11906));
AOI21X1 g124395(.A0 (n_11903), .A1 (n_8484), .B0 (n_9300), .Y(n_11904));
AOI21X1 g124397(.A0 (n_11900), .A1 (n_11916), .B0 (n_9703), .Y(n_11901));
AOI21X1 g124399(.A0 (n_11692), .A1 (n_8484), .B0 (n_9713), .Y(n_11899));
AOI21X1 g124401(.A0 (n_11897), .A1 (n_11916), .B0 (n_9239), .Y(n_11898));
AOI21X1 g124407(.A0 (n_11621), .A1 (n_8484), .B0 (n_9709), .Y(n_11896));
AOI21X1 g124410(.A0 (n_11623), .A1 (n_8400), .B0 (n_9810), .Y(n_11894));
AOI21X1 g124414(.A0 (n_11624), .A1 (n_8400), .B0 (n_9822), .Y(n_11893));
AOI21X1 g124417(.A0 (n_11875), .A1 (n_8400), .B0 (n_9803), .Y(n_11892));
AOI21X1 g124419(.A0 (n_11631), .A1 (n_9310), .B0 (n_9823), .Y(n_11891));
AOI21X1 g124420(.A0 (n_11630), .A1 (n_9310), .B0 (n_9802), .Y(n_11890));
AOI21X1 g124421(.A0 (n_11635), .A1 (n_8484), .B0 (n_9182), .Y(n_11889));
AOI21X1 g124422(.A0 (n_11887), .A1 (n_8484), .B0 (n_9710), .Y(n_11888));
NOR2X1 g124426(.A (n_11440), .B (n_11437), .Y (n_11886));
NOR2X1 g124427(.A (n_11434), .B (n_11431), .Y (n_11885));
NOR2X1 g124429(.A (n_11207), .B (n_11422), .Y (n_11884));
NOR2X1 g124430(.A (n_11203), .B (n_11419), .Y (n_11883));
NOR2X1 g124431(.A (n_11413), .B (n_11416), .Y (n_11882));
CLKBUFX3 g124440(.A (n_11880), .Y (n_12418));
INVX1 g124443(.A (n_34937), .Y (n_35420));
NAND2X1 g124446(.A (n_11876), .B (n_11875), .Y (n_11877));
INVX1 g124451(.A (n_11632), .Y (n_11874));
AOI21X1 g124454(.A0 (n_11172), .A1 (n_7209), .B0 (n_11330), .Y(n_11873));
NAND2X1 g124467(.A (n_11870), .B (n_11869), .Y (n_11871));
AND2X1 g124470(.A (n_11868), .B (n_11867), .Y (n_12373));
NAND2X1 g124472(.A (n_11865), .B (n_11864), .Y (n_11866));
NAND2X1 g124473(.A (n_11862), .B (n_11861), .Y (n_11863));
NAND2X1 g124474(.A (n_11859), .B (n_11858), .Y (n_11860));
NAND2X1 g124475(.A (n_11856), .B (n_11855), .Y (n_11857));
NAND2X1 g124476(.A (n_11853), .B (n_11852), .Y (n_11854));
NAND2X1 g124479(.A (n_11850), .B (n_11849), .Y (n_11851));
NAND2X1 g124483(.A (n_11847), .B (n_11846), .Y (n_11848));
AND2X1 g124484(.A (n_11844), .B (n_11843), .Y (n_11845));
NAND2X1 g124485(.A (n_11841), .B (n_11840), .Y (n_11842));
XOR2X1 g124490(.A (n_16644), .B (n_11150), .Y (n_11839));
NAND2X1 g124500(.A (n_11324), .B (n_33290), .Y (n_14755));
AND2X1 g124599(.A (n_11329), .B (n_13416), .Y (n_12049));
AND2X1 g124618(.A (n_9612), .B (n_11315), .Y (n_11836));
AOI22X1 g124700(.A0 (n_11832), .A1 (n_11834), .B0 (n_11825), .B1(n_11834), .Y (n_11835));
AOI22X1 g124702(.A0 (n_11832), .A1 (n_11831), .B0 (n_11356), .B1(n_11831), .Y (n_11833));
AOI22X1 g124703(.A0 (n_11832), .A1 (n_11829), .B0 (n_11356), .B1(n_11829), .Y (n_11830));
AOI22X1 g124706(.A0 (n_11832), .A1 (n_11826), .B0 (n_11825), .B1(n_11826), .Y (n_11827));
AOI22X1 g124708(.A0 (n_11832), .A1 (n_11823), .B0 (n_11825), .B1(n_11823), .Y (n_11824));
AOI22X1 g124727(.A0 (n_11832), .A1 (n_11821), .B0 (n_11356), .B1(n_11821), .Y (n_11822));
AOI22X1 g124731(.A0 (n_11832), .A1 (n_11819), .B0 (n_11356), .B1(n_11819), .Y (n_11820));
AOI22X1 g124732(.A0 (n_11832), .A1 (n_11817), .B0 (n_11825), .B1(n_11817), .Y (n_11818));
NAND2X1 g124733(.A (n_11182), .B (n_11338), .Y (n_16732));
AOI21X1 g124794(.A0 (n_10542), .A1 (n_11816), .B0 (n_11334), .Y(n_12047));
AOI21X1 g124886(.A0 (n_11812), .A1 (n_11814), .B0 (n_11312), .Y(n_11815));
AOI21X1 g124887(.A0 (n_11812), .A1 (n_11811), .B0 (n_11313), .Y(n_11813));
AOI21X1 g124888(.A0 (n_11812), .A1 (n_11809), .B0 (n_11320), .Y(n_11810));
AOI21X1 g124889(.A0 (n_11812), .A1 (n_11807), .B0 (n_11314), .Y(n_11808));
AOI21X1 g124900(.A0 (n_11575), .A1 (n_11805), .B0 (n_11322), .Y(n_11806));
MX2X1 g125278(.A (datao_2[1] ), .B (n_11290), .S0 (n_12488), .Y(n_11804));
MX2X1 g125396(.A (n_11802), .B (n_11283), .S0 (n_6435), .Y (n_11803));
MX2X1 g125398(.A (datao_1[0] ), .B (n_11288), .S0 (n_6435), .Y(n_11801));
MX2X1 g125401(.A (n_928), .B (n_11286), .S0 (n_6435), .Y (n_11800));
MX2X1 g125409(.A (datao_1[23] ), .B (n_11209), .S0 (n_6435), .Y(n_11799));
NAND3X1 g125489(.A (n_11278), .B (n_12002), .C (n_11268), .Y(n_12195));
NAND3X1 g125491(.A (n_11790), .B (n_11797), .C (n_11784), .Y(n_12007));
NOR2X1 g125542(.A (n_11793), .B (n_11540), .Y (n_12333));
NOR2X1 g125550(.A (n_11542), .B (n_11792), .Y (n_12778));
NAND3X1 g125578(.A (n_11791), .B (n_11790), .C (n_11776), .Y(n_12000));
MX2X1 g125940(.A (n_18159), .B (n_479), .S0 (n_8534), .Y (n_11789));
NOR2X1 g126028(.A (n_11788), .B (n_11989), .Y (n_12311));
NOR2X1 g126035(.A (n_11788), .B (n_11787), .Y (n_12013));
OR2X1 g126038(.A (n_11785), .B (n_11047), .Y (n_11786));
AND2X1 g126040(.A (n_11784), .B (n_11783), .Y (n_11995));
OR2X1 g126045(.A (n_11782), .B (n_11781), .Y (n_12038));
INVX1 g126047(.A (n_11779), .Y (n_11780));
OR2X1 g126056(.A (n_11782), .B (n_11778), .Y (n_11991));
AND2X1 g126066(.A (n_11777), .B (n_11776), .Y (n_12014));
NOR2X1 g126073(.A (n_11775), .B (n_11266), .Y (n_12006));
NOR2X1 g126074(.A (n_11775), .B (n_11052), .Y (n_12009));
NOR2X1 g126075(.A (n_11774), .B (n_11773), .Y (n_12790));
NOR2X1 g126079(.A (n_11772), .B (n_11778), .Y (n_12787));
NOR2X1 g126080(.A (n_11771), .B (n_11770), .Y (n_12761));
NOR2X1 g126081(.A (n_11770), .B (n_11476), .Y (n_12004));
MX2X1 g126714(.A (n_11791), .B (datao_2[9] ), .S0 (n_8400), .Y(n_11769));
MX2X1 g126718(.A (n_12827), .B (datao_2[7] ), .S0 (n_8534), .Y(n_11766));
MX2X1 g126719(.A (n_11987), .B (datao_2[18] ), .S0 (n_8400), .Y(n_11764));
MX2X1 g126726(.A (n_12003), .B (datao_2[15] ), .S0 (n_8534), .Y(n_11763));
MX2X1 g126744(.A (n_17182), .B (n_12188), .S0 (n_7871), .Y (n_11762));
MX2X1 g126752(.A (n_11759), .B (datao_1[4] ), .S0 (n_7860), .Y(n_11760));
MX2X1 g126757(.A (n_11022), .B (n_804), .S0 (n_7871), .Y (n_11756));
MX2X1 g126758(.A (n_9741), .B (n_12184), .S0 (n_7860), .Y (n_11752));
NAND2X1 g126775(.A (n_11503), .B (n_32827), .Y (n_11751));
NAND2X1 g126791(.A (n_16435), .B (n_13106), .Y (n_11750));
NAND2X1 g126796(.A (n_11791), .B (n_11797), .Y (n_11748));
NAND2X1 g126812(.A (n_18496), .B (n_12953), .Y (n_32110));
NAND2X1 g126829(.A (n_17261), .B (n_32827), .Y (n_35443));
AND2X1 g126868(.A (n_16895), .B (n_32827), .Y (n_11742));
AOI21X1 g126919(.A0 (n_11007), .A1 (n_9204), .B0 (n_11916), .Y(n_11740));
NAND2X1 g126920(.A (n_11249), .B (n_32827), .Y (n_11738));
AOI21X1 g126928(.A0 (n_11042), .A1 (n_9169), .B0 (n_7970), .Y(n_11737));
AOI21X1 g126931(.A0 (n_11008), .A1 (n_9201), .B0 (n_7970), .Y(n_11736));
AOI21X1 g126933(.A0 (n_11006), .A1 (n_10286), .B0 (n_8484), .Y(n_11734));
NAND2X1 g126934(.A (n_11988), .B (n_11732), .Y (n_11733));
NAND2X1 g126960(.A (n_34384), .B (n_11730), .Y (n_11731));
NAND2X1 g126983(.A (n_35212), .B (n_35860), .Y (n_11953));
AND2X1 g126987(.A (n_12977), .B (n_13527), .Y (n_11727));
NAND2X1 g126998(.A (n_11732), .B (n_34608), .Y (n_12174));
AOI21X1 g127005(.A0 (n_11009), .A1 (n_9203), .B0 (n_7970), .Y(n_11725));
INVX1 g128296(.A (n_11498), .Y (n_11713));
NAND2X1 g124444(.A (n_11709), .B (n_11397), .Y (n_11710));
INVX1 g124439(.A (n_11708), .Y (n_12127));
INVX1 g124209(.A (n_34983), .Y (n_11705));
NAND3X1 g124284(.A (n_10987), .B (n_10938), .C (n_10643), .Y(n_11704));
NAND3X1 g124287(.A (n_10935), .B (n_10952), .C (n_10638), .Y(n_11703));
NAND3X1 g124288(.A (n_11447), .B (n_11450), .C (n_11671), .Y(n_11702));
NAND3X1 g124290(.A (n_10974), .B (n_10971), .C (n_10646), .Y(n_11701));
NAND3X1 g124291(.A (n_10980), .B (n_10966), .C (n_10257), .Y(n_11700));
NAND3X1 g124294(.A (n_10945), .B (n_10947), .C (n_10263), .Y(n_11699));
NAND3X1 g124295(.A (n_10955), .B (n_10970), .C (n_10641), .Y(n_11698));
NAND3X1 g124296(.A (n_10985), .B (n_10939), .C (n_10261), .Y(n_11697));
NAND3X1 g124299(.A (n_10978), .B (n_10964), .C (n_10260), .Y(n_11696));
NAND3X1 g124300(.A (n_10950), .B (n_10961), .C (n_10645), .Y(n_11695));
NAND3X1 g124302(.A (n_10940), .B (n_10949), .C (n_10256), .Y(n_11694));
NAND3X1 g124304(.A (n_11692), .B (n_11639), .C (n_11643), .Y(n_11693));
NAND3X1 g124305(.A (n_11647), .B (n_11637), .C (n_11641), .Y(n_11691));
NAND3X1 g124309(.A (n_10958), .B (n_10982), .C (n_10258), .Y(n_11690));
NAND3X1 g124310(.A (n_10963), .B (n_10957), .C (n_10259), .Y(n_11689));
NAND3X1 g124312(.A (n_10937), .B (n_10944), .C (n_10640), .Y(n_11688));
NAND3X1 g124314(.A (n_10954), .B (n_10936), .C (n_10639), .Y(n_11687));
NAND3X1 g124316(.A (n_10968), .B (n_10965), .C (n_10264), .Y(n_11686));
AOI21X1 g124319(.A0 (n_10990), .A1 (n_8696), .B0 (n_10899), .Y(n_11685));
AOI21X1 g124346(.A0 (n_11429), .A1 (n_8557), .B0 (n_8556), .Y(n_11683));
AOI21X1 g124347(.A0 (n_11414), .A1 (n_8557), .B0 (n_8369), .Y(n_11682));
AOI21X1 g124349(.A0 (n_11436), .A1 (n_8552), .B0 (n_8555), .Y(n_11680));
AOI21X1 g124352(.A0 (n_11415), .A1 (n_8552), .B0 (n_8370), .Y(n_11679));
AOI21X1 g124353(.A0 (n_11438), .A1 (n_8557), .B0 (n_8553), .Y(n_11677));
AOI21X1 g124354(.A0 (n_11421), .A1 (n_8557), .B0 (n_8395), .Y(n_11676));
AOI21X1 g124355(.A0 (n_11418), .A1 (n_8552), .B0 (n_8380), .Y(n_11675));
AOI21X1 g124356(.A0 (n_11430), .A1 (n_8552), .B0 (n_8379), .Y(n_11674));
AOI21X1 g124358(.A0 (n_11671), .A1 (n_8557), .B0 (n_8354), .Y(n_11672));
AOI21X1 g124359(.A0 (n_11411), .A1 (n_8557), .B0 (n_8493), .Y(n_11670));
AOI21X1 g124360(.A0 (n_11435), .A1 (n_8557), .B0 (n_8549), .Y(n_11668));
AOI21X1 g124361(.A0 (n_11420), .A1 (n_8552), .B0 (n_8376), .Y(n_11667));
AOI21X1 g124362(.A0 (n_11426), .A1 (n_8552), .B0 (n_8547), .Y(n_11666));
AOI21X1 g124365(.A0 (n_11412), .A1 (n_8557), .B0 (n_8542), .Y(n_11665));
AOI21X1 g124366(.A0 (n_11439), .A1 (n_8557), .B0 (n_8541), .Y(n_11664));
AOI21X1 g124369(.A0 (n_11433), .A1 (n_8552), .B0 (n_8838), .Y(n_11662));
AOI21X1 g124372(.A0 (n_11660), .A1 (n_11916), .B0 (n_9298), .Y(n_11661));
MX2X1 g124373(.A (P3_d_405), .B (n_11658), .S0 (n_7970), .Y(n_11659));
AOI21X1 g124374(.A0 (n_11423), .A1 (n_8552), .B0 (n_8849), .Y(n_11657));
AOI21X1 g124375(.A0 (n_11424), .A1 (n_8552), .B0 (n_8839), .Y(n_11655));
AOI21X1 g124377(.A0 (n_11427), .A1 (n_8557), .B0 (n_8559), .Y(n_11654));
AOI21X1 g124385(.A0 (n_11651), .A1 (n_11916), .B0 (n_9177), .Y(n_11652));
AOI21X1 g124387(.A0 (n_11649), .A1 (n_7970), .B0 (n_9726), .Y(n_11650));
AOI21X1 g124388(.A0 (n_11647), .A1 (n_8484), .B0 (n_9240), .Y(n_11648));
MX2X1 g124389(.A (P3_d_386), .B (n_11645), .S0 (n_7970), .Y(n_11646));
AOI21X1 g124390(.A0 (n_11643), .A1 (n_8484), .B0 (n_9711), .Y(n_11644));
AOI21X1 g124391(.A0 (n_11641), .A1 (n_8484), .B0 (n_9276), .Y(n_11642));
AOI21X1 g124396(.A0 (n_11639), .A1 (n_8484), .B0 (n_9763), .Y(n_11640));
AOI21X1 g124398(.A0 (n_11637), .A1 (n_11916), .B0 (n_9698), .Y(n_11638));
INVX1 g124441(.A (n_11405), .Y (n_11880));
NAND2X1 g124449(.A (n_11635), .B (n_11634), .Y (n_11636));
AND2X1 g124450(.A (n_11709), .B (n_11192), .Y (n_11633));
NAND2X1 g124452(.A (n_11631), .B (n_11630), .Y (n_11632));
NAND2X1 g124453(.A (n_11628), .B (n_7209), .Y (n_11629));
INVX1 g124459(.A (n_11428), .Y (n_11627));
INVX1 g124461(.A (n_11425), .Y (n_11626));
NAND2X1 g124480(.A (n_11624), .B (n_11623), .Y (n_11625));
NAND2X1 g124481(.A (n_11621), .B (n_11620), .Y (n_11622));
NAND4X1 g124486(.A (n_11183), .B (n_16186), .C (n_32885), .D(n_9268), .Y (n_11619));
NOR2X1 g124506(.A (n_11175), .B (n_33), .Y (n_12214));
AND2X1 g124561(.A (n_11078), .B (n_34933), .Y (n_12206));
INVX1 g124575(.A (n_11617), .Y (n_11837));
NOR2X1 g124603(.A (n_11293), .B (n_32373), .Y (n_12208));
OAI21X1 g124622(.A0 (n_11615), .A1 (n_10203), .B0 (n_8696), .Y(n_11616));
AOI22X1 g124626(.A0 (n_10834), .A1 (n_11080), .B0 (n_11339), .B1(n_16176), .Y (n_16778));
AOI22X1 g124627(.A0 (n_11612), .A1 (addr_439), .B0 (n_11610), .B1(n_11819), .Y (n_11614));
AOI22X1 g124630(.A0 (n_11612), .A1 (n_8361), .B0 (n_11610), .B1(n_11834), .Y (n_11613));
AOI22X1 g124631(.A0 (n_11612), .A1 (addr_429), .B0 (n_11610), .B1(n_11831), .Y (n_11611));
AOI22X1 g124632(.A0 (n_11612), .A1 (addr_430), .B0 (n_11610), .B1(n_11829), .Y (n_11609));
AOI22X1 g124634(.A0 (n_11612), .A1 (addr_431), .B0 (n_11610), .B1(n_11607), .Y (n_11608));
AOI22X1 g124635(.A0 (n_11612), .A1 (addr_432), .B0 (n_11610), .B1(n_11605), .Y (n_11606));
AOI22X1 g124640(.A0 (n_11612), .A1 (addr_435), .B0 (n_11610), .B1(n_11826), .Y (n_11604));
AOI22X1 g124642(.A0 (n_11612), .A1 (n_8117), .B0 (n_11610), .B1(n_11601), .Y (n_11602));
AOI22X1 g124645(.A0 (n_11612), .A1 (addr_434), .B0 (n_11610), .B1(n_11599), .Y (n_11600));
AOI22X1 g124650(.A0 (n_11612), .A1 (addr_441), .B0 (n_11610), .B1(n_11821), .Y (n_11598));
AOI22X1 g124671(.A0 (n_11832), .A1 (n_11596), .B0 (n_11586), .B1(n_11596), .Y (n_11597));
AOI22X1 g124675(.A0 (n_11612), .A1 (addr_433), .B0 (n_11610), .B1(n_11594), .Y (n_11595));
AOI22X1 g124688(.A0 (n_11612), .A1 (addr_437), .B0 (n_11610), .B1(n_11592), .Y (n_11593));
AOI22X1 g124690(.A0 (n_11612), .A1 (addr_438), .B0 (n_11610), .B1(n_11823), .Y (n_11591));
AOI22X1 g124691(.A0 (n_11612), .A1 (addr_442), .B0 (n_11610), .B1(n_11817), .Y (n_11590));
AOI22X1 g124694(.A0 (n_11612), .A1 (addr_436), .B0 (n_11610), .B1(n_11588), .Y (n_11589));
AOI22X1 g124695(.A0 (n_11832), .A1 (n_11805), .B0 (n_11586), .B1(n_11805), .Y (n_11587));
AOI22X1 g124698(.A0 (n_11832), .A1 (n_11584), .B0 (n_11586), .B1(n_11584), .Y (n_11585));
AOI22X1 g124701(.A0 (n_11832), .A1 (n_11594), .B0 (n_11586), .B1(n_11594), .Y (n_11583));
AOI22X1 g124704(.A0 (n_11832), .A1 (n_11607), .B0 (n_11586), .B1(n_11607), .Y (n_11582));
AOI22X1 g124705(.A0 (n_11832), .A1 (n_11605), .B0 (n_11586), .B1(n_11605), .Y (n_11581));
AOI22X1 g124711(.A0 (n_11832), .A1 (n_11588), .B0 (n_11586), .B1(n_11588), .Y (n_11580));
AOI22X1 g124728(.A0 (n_11832), .A1 (n_11592), .B0 (n_11586), .B1(n_11592), .Y (n_11579));
AOI22X1 g124729(.A0 (n_11832), .A1 (n_11599), .B0 (n_11586), .B1(n_11599), .Y (n_11578));
AOI22X1 g124730(.A0 (n_11832), .A1 (n_11601), .B0 (n_11586), .B1(n_11601), .Y (n_11577));
AOI21X1 g124881(.A0 (n_11575), .A1 (n_11584), .B0 (n_11112), .Y(n_11576));
AOI21X1 g124885(.A0 (n_11812), .A1 (n_11573), .B0 (n_11111), .Y(n_11574));
NOR2X1 g124932(.A (n_11572), .B (n_11571), .Y (n_12044));
OR2X1 g124933(.A (n_11307), .B (n_11569), .Y (n_11570));
NOR3X1 g125118(.A (n_35861), .B (n_11772), .C (n_11294), .Y(n_11568));
NAND2X1 g125228(.A (n_10038), .B (n_11096), .Y (n_11567));
AOI21X1 g125238(.A0 (n_32857), .A1 (n_10797), .B0 (n_32945), .Y(n_11566));
MX2X1 g125272(.A (datao_2[0] ), .B (n_11072), .S0 (n_12464), .Y(n_11565));
MX2X1 g125289(.A (datao_2[2] ), .B (n_11074), .S0 (n_12488), .Y(n_11564));
MX2X1 g125399(.A (datao_1[11] ), .B (n_11070), .S0 (n_6435), .Y(n_11563));
MX2X1 g125415(.A (n_732), .B (n_11069), .S0 (n_6435), .Y (n_11561));
NAND3X1 g125470(.A (n_17955), .B (n_10754), .C (n_11558), .Y(n_12037));
NAND3X1 g125520(.A (n_11558), .B (n_16904), .C (n_11559), .Y(n_12046));
NAND3X1 g125532(.A (n_11556), .B (n_11555), .C (n_34867), .Y(n_12347));
INVX1 g125540(.A (n_11552), .Y (n_11553));
NAND3X1 g125552(.A (n_17468), .B (n_9754), .C (n_11060), .Y(n_12039));
OAI21X1 g125937(.A0 (n_16452), .A1 (n_34651), .B0 (n_11003), .Y(n_11551));
MX2X1 g125939(.A (n_16452), .B (datao_2[31] ), .S0 (n_8534), .Y(n_11550));
MX2X1 g125941(.A (n_11548), .B (datao_1[29] ), .S0 (n_7871), .Y(n_11549));
MX2X1 g125943(.A (n_16176), .B (datao_1[31] ), .S0 (n_7871), .Y(n_11546));
CLKBUFX1 gbuf_d_698(.A(n_11040), .Y(d_out_698));
CLKBUFX1 gbuf_qn_698(.A(qn_in_698), .Y(wr_2));
NOR2X1 g126034(.A (n_11052), .B (n_11544), .Y (n_11545));
NOR2X1 g126036(.A (n_11544), .B (n_13095), .Y (n_11543));
NOR2X1 g126048(.A (n_11061), .B (n_11302), .Y (n_11779));
INVX1 g126049(.A (n_11541), .Y (n_11542));
INVX1 g126051(.A (n_11539), .Y (n_11540));
NAND2X1 g126053(.A (n_34931), .B (n_11536), .Y (n_11538));
NAND2X1 g126054(.A (n_11064), .B (n_11534), .Y (n_11535));
NAND2X1 g126059(.A (n_16796), .B (n_16460), .Y (n_11533));
AND2X1 g126096(.A (n_11528), .B (n_11783), .Y (n_11529));
MX2X1 g126708(.A (n_10326), .B (datao_2[5] ), .S0 (n_8534), .Y(n_11527));
MX2X1 g126735(.A (n_9725), .B (datao_1[10] ), .S0 (n_7871), .Y(n_11526));
MX2X1 g126736(.A (n_17955), .B (n_12030), .S0 (n_7871), .Y (n_11525));
MX2X1 g126737(.A (n_10755), .B (n_12028), .S0 (n_7871), .Y (n_11523));
MX2X1 g126741(.A (n_11556), .B (datao_1[19] ), .S0 (n_7871), .Y(n_11521));
MX2X1 g126743(.A (n_17162), .B (n_12026), .S0 (n_7871), .Y (n_11520));
MX2X1 g126751(.A (n_12232), .B (n_12022), .S0 (n_7860), .Y (n_11519));
MX2X1 g126753(.A (n_10333), .B (datao_1[5] ), .S0 (n_7871), .Y(n_11518));
NAND2X1 g126770(.A (n_35212), .B (n_13106), .Y (n_11515));
AOI21X1 g126776(.A0 (n_9542), .A1 (n_10697), .B0 (n_8484), .Y(n_11513));
NAND2X1 g126778(.A (n_12003), .B (n_32827), .Y (n_11512));
NAND2X1 g126781(.A (n_16165), .B (n_10497), .Y (n_11990));
NOR2X1 g126794(.A (n_10792), .B (n_10716), .Y (n_11508));
NOR2X1 g126800(.A (n_11256), .B (n_10317), .Y (n_11507));
NOR2X1 g126813(.A (n_10826), .B (n_11280), .Y (n_11994));
AOI21X1 g126832(.A0 (n_9645), .A1 (n_10675), .B0 (n_8484), .Y(n_11506));
NAND2X1 g126837(.A (n_11791), .B (n_32827), .Y (n_11504));
NAND2X1 g126867(.A (n_16748), .B (n_11503), .Y (n_12175));
NOR2X1 g126874(.A (n_10320), .B (n_10689), .Y (n_12337));
AND2X1 g126877(.A (n_19666), .B (n_12953), .Y (n_11501));
INVX1 g126913(.A (n_11500), .Y (n_13114));
AOI21X1 g126921(.A0 (n_9643), .A1 (n_10657), .B0 (n_8484), .Y(n_11497));
AOI21X1 g126922(.A0 (n_9544), .A1 (n_10684), .B0 (n_8484), .Y(n_11496));
AOI21X1 g126923(.A0 (n_9651), .A1 (n_10688), .B0 (n_8484), .Y(n_11495));
AOI21X1 g126925(.A0 (n_9650), .A1 (n_10682), .B0 (n_7970), .Y(n_11493));
AOI21X1 g126927(.A0 (n_9552), .A1 (n_10680), .B0 (n_11916), .Y(n_11492));
AOI21X1 g126930(.A0 (n_9648), .A1 (n_10678), .B0 (n_11916), .Y(n_11491));
NAND2X1 g126932(.A (n_17182), .B (n_12953), .Y (n_11490));
AOI21X1 g126935(.A0 (n_9641), .A1 (n_10693), .B0 (n_8484), .Y(n_11489));
AOI21X1 g126936(.A0 (n_9642), .A1 (n_10691), .B0 (n_8484), .Y(n_11488));
AOI21X1 g126938(.A0 (n_9578), .A1 (n_10741), .B0 (n_8484), .Y(n_11487));
AOI21X1 g126942(.A0 (n_9647), .A1 (n_10672), .B0 (n_8484), .Y(n_11486));
NOR2X1 g126943(.A (n_11790), .B (n_11483), .Y (n_11485));
NAND2X1 g126965(.A (n_11481), .B (n_13106), .Y (n_11482));
NAND2X1 g126970(.A (n_11022), .B (n_12953), .Y (n_11480));
AND2X1 g126984(.A (n_32350), .B (n_32827), .Y (n_11479));
AOI21X1 g126985(.A0 (n_9646), .A1 (n_10686), .B0 (n_8484), .Y(n_11478));
INVX1 g126992(.A (n_11476), .Y (n_11477));
INVX1 g128032(.A (n_11470), .Y (n_12561));
INVX1 g128142(.A (n_11730), .Y (n_11720));
INVX1 g128258(.A (n_11468), .Y (n_11716));
INVX1 g128319(.A (n_11988), .Y (n_11712));
MX2X1 g126755(.A (n_18584), .B (datao_1[9] ), .S0 (n_7871), .Y(n_11458));
MX2X1 g126748(.A (n_34384), .B (datao_1[27] ), .S0 (n_7871), .Y(n_11457));
MX2X1 g126711(.A (n_35244), .B (datao_2[19] ), .S0 (n_8534), .Y(n_11456));
NAND4X1 g124301(.A (n_10989), .B (n_7972), .C (n_8059), .D (n_10254),.Y (n_11454));
AOI21X1 g124345(.A0 (n_11417), .A1 (n_8557), .B0 (n_8558), .Y(n_11453));
AOI21X1 g124350(.A0 (n_11200), .A1 (n_8552), .B0 (n_8554), .Y(n_11452));
AOI21X1 g124351(.A0 (n_11450), .A1 (n_8552), .B0 (n_8596), .Y(n_11451));
AOI21X1 g124357(.A0 (n_11199), .A1 (n_8557), .B0 (n_8857), .Y(n_11449));
AOI21X1 g124363(.A0 (n_11447), .A1 (n_8557), .B0 (n_8473), .Y(n_11448));
AOI21X1 g124364(.A0 (n_11202), .A1 (n_8557), .B0 (n_8545), .Y(n_11446));
AOI21X1 g124367(.A0 (n_11205), .A1 (n_7860), .B0 (n_8357), .Y(n_11445));
AOI21X1 g124368(.A0 (n_11201), .A1 (n_7860), .B0 (n_8378), .Y(n_11443));
AOI21X1 g124370(.A0 (n_11206), .A1 (n_8552), .B0 (n_8540), .Y(n_11442));
AOI21X1 g124424(.A0 (n_11432), .A1 (n_8557), .B0 (n_8544), .Y(n_11441));
NAND2X1 g124455(.A (n_11439), .B (n_11438), .Y (n_11440));
NAND2X1 g124456(.A (n_11436), .B (n_11435), .Y (n_11437));
NAND2X1 g124457(.A (n_11433), .B (n_11432), .Y (n_11434));
NAND2X1 g124458(.A (n_11430), .B (n_11429), .Y (n_11431));
NAND2X1 g124460(.A (n_11427), .B (n_11426), .Y (n_11428));
NAND2X1 g124462(.A (n_11424), .B (n_11423), .Y (n_11425));
NAND2X1 g124463(.A (n_11421), .B (n_11420), .Y (n_11422));
NAND2X1 g124466(.A (n_11418), .B (n_11417), .Y (n_11419));
NAND2X1 g124468(.A (n_11415), .B (n_11414), .Y (n_11416));
NAND2X1 g124477(.A (n_11412), .B (n_11411), .Y (n_11413));
NAND2X1 g124503(.A (n_11410), .B (P2_d_389), .Y (n_11865));
NAND2X1 g124518(.A (n_11410), .B (P2_d_405), .Y (n_11869));
NAND2X1 g124533(.A (n_11410), .B (P2_d_393), .Y (n_11868));
NAND2X1 g124546(.A (n_11407), .B (P2_d_384), .Y (n_11855));
NAND2X1 g124547(.A (n_11407), .B (P2_d_408), .Y (n_11864));
NAND2X1 g124549(.A (n_33405), .B (P3_d_393), .Y (n_12078));
NAND2X1 g124550(.A (n_11399), .B (P2_d_392), .Y (n_11847));
NAND2X1 g124552(.A (n_11407), .B (P2_d_396), .Y (n_11844));
NAND2X1 g124553(.A (n_11404), .B (n_11402), .Y (n_11405));
NAND2X1 g124557(.A (n_11407), .B (P2_d_402), .Y (n_11876));
NAND2X1 g124558(.A (n_11403), .B (P2_d_391), .Y (n_12374));
NAND2X1 g124559(.A (n_11403), .B (P2_d_407), .Y (n_11852));
NAND2X1 g124562(.A (n_11410), .B (P2_d_386), .Y (n_11861));
NAND2X1 g124567(.A (n_11410), .B (P2_d_403), .Y (n_11841));
AND2X1 g124576(.A (n_10793), .B (n_11402), .Y (n_11617));
NAND2X1 g124578(.A (n_11399), .B (P2_d_398), .Y (n_11850));
NAND2X1 g124580(.A (n_11401), .B (n_32374), .Y (n_11708));
NAND2X2 g124581(.A (n_11407), .B (P2_d_383), .Y (n_11859));
NAND2X1 g124583(.A (n_11403), .B (P2_d_401), .Y (n_11867));
NAND2X1 g124585(.A (n_11399), .B (P2_d_404), .Y (n_11843));
NAND2X1 g124587(.A (n_11399), .B (P2_d_387), .Y (n_11849));
NAND2X1 g124588(.A (n_11403), .B (P2_d_388), .Y (n_11853));
NAND2X1 g124591(.A (n_11403), .B (P2_d_390), .Y (n_11840));
NAND2X1 g124594(.A (n_11410), .B (P2_d_397), .Y (n_11862));
NAND2X1 g124597(.A (n_11399), .B (P2_d_381), .Y (n_11846));
NAND2X1 g124602(.A (n_11410), .B (P2_d_382), .Y (n_11870));
NAND2X1 g124605(.A (n_11410), .B (P2_d_399), .Y (n_11856));
INVX1 g124612(.A (n_11396), .Y (n_12098));
AND2X1 g124614(.A (n_9615), .B (n_10872), .Y (n_11395));
AND2X1 g124615(.A (n_9614), .B (n_10871), .Y (n_11394));
AOI21X1 g124620(.A0 (n_10630), .A1 (n_12670), .B0 (n_11086), .Y(n_11393));
AOI22X1 g124653(.A0 (n_11389), .A1 (n_1170), .B0 (n_14349), .B1(n_11391), .Y (n_11392));
AOI22X1 g124656(.A0 (n_11389), .A1 (addr_492), .B0 (n_14349), .B1(n_11388), .Y (n_11390));
AOI22X1 g124657(.A0 (n_11389), .A1 (n_9655), .B0 (n_14349), .B1(n_11386), .Y (n_11387));
AOI22X1 g124658(.A0 (n_11389), .A1 (n_9670), .B0 (n_14349), .B1(n_11384), .Y (n_11385));
AOI22X1 g124659(.A0 (n_11389), .A1 (n_9653), .B0 (n_14349), .B1(n_11382), .Y (n_11383));
AOI22X1 g124660(.A0 (n_11389), .A1 (n_9672), .B0 (n_14349), .B1(n_11380), .Y (n_11381));
AOI22X1 g124661(.A0 (n_11389), .A1 (n_9667), .B0 (n_14349), .B1(n_11378), .Y (n_11379));
AOI22X1 g124663(.A0 (n_11389), .A1 (n_9658), .B0 (n_14349), .B1(n_11376), .Y (n_11377));
AOI22X1 g124664(.A0 (n_11389), .A1 (n_9675), .B0 (n_14349), .B1(n_11374), .Y (n_11375));
AOI22X1 g124665(.A0 (n_11389), .A1 (n_9663), .B0 (n_14349), .B1(n_11372), .Y (n_11373));
AOI22X1 g124666(.A0 (n_11389), .A1 (addr_487), .B0 (n_14349), .B1(n_11370), .Y (n_11371));
AOI22X1 g124667(.A0 (n_11389), .A1 (addr_488), .B0 (n_14349), .B1(n_11368), .Y (n_11369));
AOI22X1 g124668(.A0 (n_11389), .A1 (addr_489), .B0 (n_14349), .B1(n_11366), .Y (n_11367));
AOI22X1 g124669(.A0 (n_11389), .A1 (addr_490), .B0 (n_14349), .B1(n_11364), .Y (n_11365));
AOI22X1 g124670(.A0 (n_11389), .A1 (addr_491), .B0 (n_14349), .B1(n_11362), .Y (n_11363));
AOI22X1 g124696(.A0 (n_11832), .A1 (n_11360), .B0 (n_11356), .B1(n_11360), .Y (n_11361));
AOI22X1 g124697(.A0 (n_11354), .A1 (n_11378), .B0 (n_11353), .B1(n_11378), .Y (n_11359));
AOI22X1 g124699(.A0 (n_11832), .A1 (n_11357), .B0 (n_11356), .B1(n_11357), .Y (n_11358));
AOI22X1 g124707(.A0 (n_11354), .A1 (n_11380), .B0 (n_11353), .B1(n_11380), .Y (n_11355));
AOI22X1 g124709(.A0 (n_11354), .A1 (n_11362), .B0 (n_11353), .B1(n_11362), .Y (n_11352));
AOI22X1 g124710(.A0 (n_11354), .A1 (n_11372), .B0 (n_11353), .B1(n_11372), .Y (n_11351));
AOI22X1 g124712(.A0 (n_11354), .A1 (n_11364), .B0 (n_11353), .B1(n_11364), .Y (n_11350));
AOI22X1 g124713(.A0 (n_11354), .A1 (n_11386), .B0 (n_11353), .B1(n_11386), .Y (n_11349));
AOI22X1 g124714(.A0 (n_11354), .A1 (n_11366), .B0 (n_11353), .B1(n_11366), .Y (n_11348));
AOI22X1 g124715(.A0 (n_11354), .A1 (n_11388), .B0 (n_11353), .B1(n_11388), .Y (n_11347));
AOI22X1 g124716(.A0 (n_11354), .A1 (n_11384), .B0 (n_11353), .B1(n_11384), .Y (n_11346));
AOI22X1 g124717(.A0 (n_11354), .A1 (n_11382), .B0 (n_11353), .B1(n_11382), .Y (n_11345));
AOI22X1 g124718(.A0 (n_11354), .A1 (n_11376), .B0 (n_11353), .B1(n_11376), .Y (n_11344));
AOI22X1 g124723(.A0 (n_11354), .A1 (n_11368), .B0 (n_11353), .B1(n_11368), .Y (n_11343));
AOI22X1 g124724(.A0 (n_11354), .A1 (n_11391), .B0 (n_11353), .B1(n_11391), .Y (n_11342));
AOI22X1 g124725(.A0 (n_11354), .A1 (n_11374), .B0 (n_11353), .B1(n_11374), .Y (n_11341));
AOI22X1 g124726(.A0 (n_11354), .A1 (n_11370), .B0 (n_11353), .B1(n_11370), .Y (n_11340));
XOR2X1 g124734(.A (n_10745), .B (n_11339), .Y (n_16735));
NAND2X1 g124833(.A (n_10836), .B (n_10467), .Y (n_11338));
AOI21X1 g124928(.A0 (n_10795), .A1 (n_8436), .B0 (n_11333), .Y(n_11334));
AOI21X1 g125211(.A0 (n_29381), .A1 (n_34719), .B0 (n_8113), .Y(n_11330));
AOI21X1 g125217(.A0 (n_9219), .A1 (n_10505), .B0 (n_11402), .Y(n_11329));
AOI22X1 g125224(.A0 (n_20218), .A1 (n_11327), .B0 (n_13169), .B1(n_8946), .Y (n_11328));
NAND2X1 g125232(.A (n_10037), .B (n_10829), .Y (n_11326));
NAND2X1 g125246(.A (n_10031), .B (n_10831), .Y (n_11325));
AOI21X1 g125250(.A0 (n_15749), .A1 (n_10821), .B0 (n_32371), .Y(n_11324));
INVX1 g125302(.A (n_11140), .Y (n_11322));
AOI22X1 g125310(.A0 (n_11584), .A1 (n_25636), .B0 (n_14850), .B1(addr_426), .Y (n_11321));
INVX1 g125315(.A (n_11139), .Y (n_11320));
INVX1 g125317(.A (n_11137), .Y (n_11319));
AOI22X1 g125319(.A0 (n_11805), .A1 (n_25636), .B0 (n_14850), .B1(addr_424), .Y (n_11318));
AOI22X1 g125341(.A0 (n_11596), .A1 (n_25082), .B0 (n_20218), .B1(addr_1), .Y (n_11317));
AOI22X1 g125365(.A0 (n_11596), .A1 (n_28013), .B0 (n_15288), .B1(addr_1), .Y (n_11315));
INVX1 g125377(.A (n_11104), .Y (n_11314));
INVX1 g125383(.A (n_11101), .Y (n_11313));
INVX1 g125389(.A (n_11098), .Y (n_11312));
MX2X1 g125405(.A (datao_1[1] ), .B (n_10774), .S0 (n_6435), .Y(n_11311));
INVX1 g125508(.A (n_11309), .Y (n_11310));
INVX1 g125515(.A (n_11307), .Y (n_11308));
NAND3X1 g125541(.A (n_17471), .B (n_17467), .C (n_11306), .Y(n_11552));
CLKBUFX1 gbuf_d_699(.A(n_10744), .Y(d_out_699));
CLKBUFX1 gbuf_qn_699(.A(qn_in_699), .Y(wr_3));
NAND2X1 g126044(.A (n_11306), .B (n_11305), .Y (n_11793));
NOR2X1 g126050(.A (n_11304), .B (n_11303), .Y (n_11541));
NOR2X1 g126052(.A (n_11302), .B (n_11065), .Y (n_11539));
OR2X1 g126058(.A (n_11301), .B (n_11300), .Y (n_11792));
OR2X1 g126067(.A (n_11301), .B (n_11774), .Y (n_11571));
NAND3X1 g126070(.A (n_10335), .B (n_10712), .C (n_35203), .Y(n_11299));
OR2X1 g126076(.A (n_11296), .B (n_11295), .Y (n_11297));
INVX1 g126085(.A (n_11294), .Y (n_11530));
NOR2X1 g126093(.A (n_11772), .B (n_35404), .Y (n_12343));
NAND2X1 g126095(.A (n_11048), .B (n_11050), .Y (n_11293));
MX2X1 g126727(.A (n_33268), .B (datao_2[1] ), .S0 (n_8534), .Y(n_11290));
MX2X1 g126734(.A (n_12532), .B (datao_1[0] ), .S0 (n_7871), .Y(n_11288));
MX2X1 g126759(.A (n_11285), .B (n_928), .S0 (n_7871), .Y (n_11286));
MX2X1 g126761(.A (n_11089), .B (n_11802), .S0 (n_7860), .Y (n_11283));
NAND2X1 g126771(.A (n_35244), .B (n_32827), .Y (n_11281));
NOR2X1 g126782(.A (n_11275), .B (n_11280), .Y (n_11776));
NAND2X1 g126804(.A (n_32356), .B (n_11278), .Y (n_11788));
NAND2X1 g126807(.A (n_11276), .B (n_13106), .Y (n_11277));
NOR2X1 g126809(.A (n_15908), .B (n_11275), .Y (n_11784));
NOR2X1 g126820(.A (n_10309), .B (n_11797), .Y (n_11274));
NAND2X1 g126824(.A (n_9725), .B (n_13527), .Y (n_11272));
NAND2X1 g126831(.A (n_17906), .B (n_13106), .Y (n_32251));
NAND2X1 g126834(.A (n_12703), .B (n_11269), .Y (n_11771));
INVX1 g126854(.A (n_11787), .Y (n_11268));
INVX1 g126858(.A (n_11267), .Y (n_11773));
INVX1 g126859(.A (n_11267), .Y (n_11266));
NAND2X1 g126873(.A (n_10755), .B (n_12953), .Y (n_11265));
NAND2X1 g126879(.A (n_35202), .B (n_10768), .Y (n_11782));
NAND2X2 g126893(.A (n_10713), .B (n_35860), .Y (n_11778));
NOR2X1 g126903(.A (n_17468), .B (n_17467), .Y (n_11264));
INVX1 g126915(.A (n_16460), .Y (n_11500));
NAND2X1 g126918(.A (n_11556), .B (n_12953), .Y (n_11261));
NAND2X1 g126924(.A (n_17162), .B (n_12953), .Y (n_11260));
NAND2X1 g126937(.A (n_8829), .B (n_11256), .Y (n_11258));
NAND2X1 g126955(.A (n_10326), .B (n_32827), .Y (n_11253));
NOR2X1 g126964(.A (n_11030), .B (n_11010), .Y (n_11777));
NOR2X1 g126966(.A (n_16186), .B (n_9745), .Y (n_11993));
NAND2X1 g126967(.A (n_11033), .B (n_18496), .Y (n_11250));
NAND2X1 g126973(.A (n_11249), .B (n_12827), .Y (n_11785));
NAND2X1 g126975(.A (n_34384), .B (n_12953), .Y (n_32301));
INVX1 g126977(.A (n_11989), .Y (n_11247));
NAND2X1 g126993(.A (n_35318), .B (n_11246), .Y (n_11476));
NOR2X1 g126996(.A (n_10711), .B (n_12690), .Y (n_11245));
INVX1 g128259(.A (n_18475), .Y (n_11468));
INVX1 g127668(.A (n_11057), .Y (n_12977));
INVX1 g128026(.A (n_16796), .Y (n_11961));
CLKBUFX1 g128033(.A (n_10689), .Y (n_11470));
INVX1 g128143(.A (n_16174), .Y (n_11730));
INVX1 g128185(.A (n_11227), .Y (n_13102));
INVX1 g128231(.A (n_16754), .Y (n_11732));
INVX1 g128239(.A (n_34617), .Y (n_11226));
INVX1 g128249(.A (n_34992), .Y (n_11747));
INVX1 g128298(.A (n_11278), .Y (n_11498));
INVX1 g128312(.A (n_11222), .Y (n_11464));
CLKBUFX1 g128320(.A (n_10497), .Y (n_11988));
AOI22X1 g129127(.A0 (n_5356), .A1 (n_10676), .B0 (n_10671), .B1(n_3429), .Y (n_11213));
NAND3X1 g129326(.A (n_7550), .B (n_7549), .C (n_10676), .Y (n_11211));
NOR2X1 g126042(.A (n_11210), .B (n_10794), .Y (n_12035));
MX2X1 g126745(.A (n_12943), .B (datao_1[23] ), .S0 (n_7871), .Y(n_11209));
NAND2X1 g124584(.A (n_11208), .B (P2_d_379), .Y (n_11875));
INVX1 g124589(.A (n_10991), .Y (n_11939));
NAND2X1 g124565(.A (n_11208), .B (P2_d_385), .Y (n_11631));
NAND2X1 g124464(.A (n_11206), .B (n_11205), .Y (n_11207));
NAND2X1 g124465(.A (n_11202), .B (n_11201), .Y (n_11203));
NAND2X1 g124469(.A (n_11200), .B (n_11199), .Y (n_11938));
AOI21X1 g124488(.A0 (n_10050), .A1 (n_27042), .B0 (n_11197), .Y(n_11198));
NAND2X1 g124501(.A (n_11208), .B (P2_d_395), .Y (n_11623));
NAND2X1 g124504(.A (n_33405), .B (P3_d_396), .Y (n_11903));
NAND2X1 g124505(.A (n_11195), .B (P3_d_388), .Y (n_11921));
NAND2X1 g124512(.A (n_10655), .B (P3_d_401), .Y (n_11621));
NAND2X1 g124531(.A (n_11208), .B (P2_d_380), .Y (n_11624));
NAND2X1 g124548(.A (n_11194), .B (P3_d_392), .Y (n_11709));
NAND2X1 g124563(.A (n_11195), .B (P3_d_404), .Y (n_11692));
NAND2X1 g124568(.A (n_11194), .B (P3_d_387), .Y (n_11917));
NAND2X1 g124569(.A (n_11195), .B (P3_d_395), .Y (n_11905));
NAND2X1 g124570(.A (n_10655), .B (P3_d_397), .Y (n_11634));
NAND2X1 g124571(.A (n_11195), .B (P3_d_402), .Y (n_11900));
NAND2X1 g124572(.A (n_10655), .B (P3_d_378), .Y (n_11620));
NAND2X1 g124573(.A (n_11194), .B (P3_d_379), .Y (n_11897));
NAND2X1 g124577(.A (n_11195), .B (P3_d_394), .Y (n_11908));
NAND2X1 g124582(.A (n_11208), .B (P2_d_400), .Y (n_11630));
NAND2X1 g124593(.A (n_11194), .B (P3_d_383), .Y (n_11887));
NAND2X1 g124600(.A (n_10655), .B (P3_d_382), .Y (n_11635));
NAND2X2 g124604(.A (n_11208), .B (P2_d_406), .Y (n_11858));
NAND2X1 g124606(.A (n_11194), .B (P3_d_389), .Y (n_11911));
INVX1 g124608(.A (n_11192), .Y (n_11397));
NAND4X1 g124611(.A (n_10023), .B (n_34951), .C (n_34752), .D(n_8678), .Y (n_11923));
NAND3X1 g124613(.A (n_11191), .B (n_10249), .C (n_10035), .Y(n_11396));
NAND4X1 g124619(.A (n_9172), .B (n_21365), .C (n_35043), .D(n_25119), .Y (n_11628));
AOI22X1 g124621(.A0 (n_10514), .A1 (n_27042), .B0 (n_10204), .B1(n_27042), .Y (n_11190));
AOI22X1 g124719(.A0 (n_11354), .A1 (n_11814), .B0 (n_11353), .B1(n_11814), .Y (n_11188));
AOI22X1 g124720(.A0 (n_11354), .A1 (n_11811), .B0 (n_11353), .B1(n_11811), .Y (n_11187));
AOI22X1 g124721(.A0 (n_11354), .A1 (n_11809), .B0 (n_11353), .B1(n_11809), .Y (n_11186));
AOI22X1 g124722(.A0 (n_11354), .A1 (n_11807), .B0 (n_11353), .B1(n_11807), .Y (n_11185));
NAND2X1 g124799(.A (n_11183), .B (n_9375), .Y (n_11184));
NAND2X1 g124800(.A (n_11181), .B (n_34651), .Y (n_11182));
NAND2X1 g124804(.A (n_11177), .B (n_11378), .Y (n_11179));
NAND2X1 g124813(.A (n_11177), .B (n_11386), .Y (n_11178));
NAND2X1 g124814(.A (n_11177), .B (n_11380), .Y (n_11176));
INVX1 g124817(.A (n_11399), .Y (n_11175));
NAND2X1 g124823(.A (n_11177), .B (n_11376), .Y (n_11174));
NAND2X1 g124826(.A (n_11177), .B (n_11362), .Y (n_11173));
NAND3X1 g124827(.A (n_29388), .B (n_10629), .C (n_10776), .Y(n_11172));
NAND2X1 g124835(.A (n_11177), .B (n_11372), .Y (n_11171));
NAND2X1 g124840(.A (n_11177), .B (n_11366), .Y (n_11170));
NAND2X1 g124843(.A (n_11177), .B (n_11364), .Y (n_11169));
NAND2X1 g124846(.A (n_11177), .B (n_11384), .Y (n_11168));
NAND2X1 g124847(.A (n_11177), .B (n_11382), .Y (n_11167));
NAND2X1 g124848(.A (n_11177), .B (n_11391), .Y (n_11166));
NAND2X1 g124853(.A (n_11177), .B (n_11368), .Y (n_11165));
NAND2X1 g124854(.A (n_11177), .B (n_11370), .Y (n_11164));
NAND2X1 g124859(.A (n_11177), .B (n_11388), .Y (n_11163));
NAND2X1 g124860(.A (n_11177), .B (n_11374), .Y (n_11162));
AOI21X1 g124884(.A0 (n_11158), .A1 (n_11160), .B0 (n_10576), .Y(n_11161));
AOI21X1 g124891(.A0 (n_11158), .A1 (n_11157), .B0 (n_10553), .Y(n_11159));
AOI21X1 g124892(.A0 (n_11158), .A1 (n_11155), .B0 (n_10551), .Y(n_11156));
AOI21X1 g124893(.A0 (n_11158), .A1 (n_11153), .B0 (n_10552), .Y(n_11154));
AOI21X1 g124894(.A0 (n_11158), .A1 (n_11151), .B0 (n_10570), .Y(n_11152));
INVX1 g124921(.A (n_11402), .Y (n_11150));
INVX1 g125008(.A (n_13761), .Y (n_11825));
AOI22X1 g125221(.A0 (n_10573), .A1 (n_11148), .B0 (n_13173), .B1(n_8946), .Y (n_11149));
NAND2X1 g125234(.A (n_10036), .B (n_10545), .Y (n_11147));
AOI22X1 g125249(.A0 (n_10573), .A1 (n_11144), .B0 (n_13301), .B1(n_8946), .Y (n_11146));
AOI22X1 g125293(.A0 (n_10573), .A1 (n_11141), .B0 (n_10822), .B1(n_8946), .Y (n_11143));
AOI22X1 g125303(.A0 (n_11805), .A1 (n_25220), .B0 (n_10573), .B1(addr_424), .Y (n_11140));
AOI22X1 g125316(.A0 (n_11809), .A1 (n_21328), .B0 (n_11138), .B1(n_190), .Y (n_11139));
AOI22X1 g125318(.A0 (n_10573), .A1 (n_11136), .B0 (n_8946), .B1(n_11135), .Y (n_11137));
AOI22X1 g125320(.A0 (n_10573), .A1 (n_4445), .B0 (n_7730), .B1(n_8946), .Y (n_11134));
INVX1 g125324(.A (n_10862), .Y (n_11130));
AOI22X1 g125328(.A0 (n_10573), .A1 (n_4277), .B0 (n_7819), .B1(n_8946), .Y (n_11129));
AOI22X1 g125329(.A0 (n_10573), .A1 (P1_reg2[19] ), .B0 (n_11122),.B1 (n_8946), .Y (n_11124));
AOI22X1 g125332(.A0 (n_10573), .A1 (n_11120), .B0 (n_7957), .B1(n_8946), .Y (n_11121));
INVX1 g125336(.A (n_10856), .Y (n_11118));
INVX1 g125346(.A (n_10851), .Y (n_11117));
AOI22X1 g125348(.A0 (n_10573), .A1 (n_3668), .B0 (n_1003), .B1(n_8946), .Y (n_11116));
INVX1 g125354(.A (n_10843), .Y (n_11113));
INVX1 g125369(.A (n_10841), .Y (n_11112));
INVX1 g125372(.A (n_10839), .Y (n_11111));
AOI22X1 g125374(.A0 (n_11811), .A1 (n_33738), .B0 (n_11107), .B1(n_2772), .Y (n_11110));
AOI22X1 g125375(.A0 (n_11809), .A1 (n_33738), .B0 (n_11107), .B1(n_190), .Y (n_11109));
AOI22X1 g125376(.A0 (n_11807), .A1 (n_33738), .B0 (n_11107), .B1(n_3314), .Y (n_11105));
AOI22X1 g125378(.A0 (n_11807), .A1 (n_21328), .B0 (n_11138), .B1(n_3314), .Y (n_11104));
AOI22X1 g125384(.A0 (n_11811), .A1 (n_21328), .B0 (n_11138), .B1(n_2772), .Y (n_11101));
AOI22X1 g125385(.A0 (n_11814), .A1 (n_33738), .B0 (n_11107), .B1(n_11097), .Y (n_11099));
AOI22X1 g125390(.A0 (n_11814), .A1 (n_21328), .B0 (n_11138), .B1(n_11097), .Y (n_11098));
NAND2X1 g125438(.A (n_20218), .B (n_3693), .Y (n_11096));
NAND3X1 g125509(.A (n_11092), .B (n_11089), .C (n_11002), .Y(n_11309));
NAND3X1 g125512(.A (n_9725), .B (n_11089), .C (n_11088), .Y(n_11572));
NAND3X1 g125516(.A (n_10754), .B (n_11089), .C (n_11088), .Y(n_11307));
INVX1 g125530(.A (n_11086), .Y (n_11087));
XOR2X1 g125936(.A (n_10799), .B (n_11079), .Y (n_11080));
NOR2X1 g126057(.A (n_10769), .B (n_10764), .Y (n_11078));
NAND2X1 g126083(.A (n_11076), .B (n_11305), .Y (n_11077));
NAND2X2 g126086(.A (n_35407), .B (n_10753), .Y (n_11294));
NOR2X1 g126097(.A (n_10461), .B (n_10468), .Y (n_11075));
MX2X1 g126721(.A (n_11401), .B (datao_2[2] ), .S0 (n_8534), .Y(n_11074));
MX2X1 g126723(.A (n_15810), .B (datao_2[0] ), .S0 (n_8534), .Y(n_11072));
MX2X1 g126733(.A (n_11092), .B (datao_1[11] ), .S0 (n_7860), .Y(n_11070));
MX2X1 g126750(.A (n_10760), .B (n_732), .S0 (n_7871), .Y (n_11069));
OAI22X1 g126779(.A0 (n_8409), .A1 (n_8407), .B0 (n_10709), .B1(n_10708), .Y (n_32900));
INVX1 g126785(.A (n_11065), .Y (n_11066));
INVX1 g126787(.A (n_11063), .Y (n_11064));
NOR2X1 g126792(.A (n_10710), .B (n_9632), .Y (n_11062));
NOR2X1 g126811(.A (n_10792), .B (n_9292), .Y (n_11528));
INVX1 g126815(.A (n_11306), .Y (n_11061));
INVX1 g126851(.A (n_11302), .Y (n_11060));
NAND2X1 g126855(.A (n_16064), .B (n_16068), .Y (n_11787));
NOR2X1 g126860(.A (n_9627), .B (n_11058), .Y (n_11267));
OR2X1 g126864(.A (n_11057), .B (n_17392), .Y (n_11544));
NAND2X1 g126869(.A (n_11285), .B (n_12953), .Y (n_35884));
NOR2X1 g126875(.A (n_10658), .B (n_11055), .Y (n_11558));
NAND2X1 g126878(.A (n_10757), .B (n_9754), .Y (n_11781));
NAND2X1 g126939(.A (n_12943), .B (n_12953), .Y (n_11053));
INVX1 g126945(.A (n_11052), .Y (n_11254));
INVX1 g126951(.A (n_11050), .Y (n_11051));
INVX1 g126957(.A (n_11048), .Y (n_11047));
NAND2X1 g126972(.A (n_12703), .B (n_13106), .Y (n_11046));
NOR2X1 g126974(.A (n_9798), .B (n_9286), .Y (n_11045));
NAND2X1 g126978(.A (n_16829), .B (n_35244), .Y (n_11989));
NAND2X1 g126988(.A (n_12986), .B (n_13106), .Y (n_11044));
NOR2X1 g126990(.A (n_9730), .B (n_9720), .Y (n_11783));
NAND2X1 g126991(.A (n_34384), .B (n_18496), .Y (n_13095));
NOR2X1 g126995(.A (n_17472), .B (n_17471), .Y (n_11043));
NAND2X1 g129604(.A (n_6396), .B (n_10676), .Y (n_11042));
NOR2X1 g127283(.A (n_10324), .B (n_6446), .Y (n_11040));
INVX2 g128232(.A (n_11037), .Y (n_16754));
INVX1 g127703(.A (n_11033), .Y (n_16442));
INVX1 g127728(.A (n_10331), .Y (n_11759));
INVX1 g127770(.A (n_11030), .Y (n_11790));
INVX1 g127994(.A (n_11275), .Y (n_11483));
INVX1 g128027(.A (n_16750), .Y (n_16796));
INVX1 g128169(.A (n_9745), .Y (n_11481));
INVX1 g128186(.A (n_11269), .Y (n_11227));
INVX1 g128260(.A (n_17348), .Y (n_18475));
INVX1 g128313(.A (n_16165), .Y (n_11222));
INVX1 g128383(.A (n_11280), .Y (n_16895));
INVX1 g128552(.A (n_11559), .Y (n_11215));
INVX2 g128563(.A (n_16429), .Y (n_16748));
INVX1 g128585(.A (n_11010), .Y (n_12002));
NAND2X1 g129574(.A (n_6438), .B (n_10676), .Y (n_11009));
NAND2X1 g129603(.A (n_6818), .B (n_10676), .Y (n_11008));
NAND2X1 g129665(.A (n_6000), .B (n_10676), .Y (n_11007));
NAND2X1 g129676(.A (n_4167), .B (n_10676), .Y (n_11006));
NAND2X1 g126094(.A (n_16452), .B (n_34651), .Y (n_11003));
NAND2X1 g126046(.A (n_11002), .B (n_11536), .Y (n_11569));
NAND2X1 g124596(.A (n_10999), .B (P3_d_390), .Y (n_11643));
INVX1 g124922(.A (n_10819), .Y (n_11402));
NAND2X1 g124502(.A (n_10999), .B (P3_d_403), .Y (n_11637));
AOI22X1 g125247(.A0 (n_10573), .A1 (n_4151), .B0 (n_7737), .B1(n_8946), .Y (n_10998));
INVX1 g124816(.A (n_10927), .Y (n_11403));
NAND2X1 g124508(.A (n_10999), .B (P3_d_385), .Y (n_11660));
NAND2X1 g124509(.A (n_32550), .B (P1_d_103), .Y (n_11424));
NAND2X1 g124510(.A (n_32548), .B (P1_d_107), .Y (n_11427));
NAND2X1 g124513(.A (n_32548), .B (P1_d_109), .Y (n_11429));
NAND2X1 g124514(.A (n_32548), .B (P1_d_110), .Y (n_11414));
NAND2X1 g124515(.A (n_32550), .B (P1_d_112), .Y (n_11436));
NAND2X1 g124516(.A (n_10999), .B (P3_d_381), .Y (n_11649));
AND2X1 g124519(.A (n_10999), .B (P3_d_386), .Y (n_11645));
NAND2X1 g124521(.A (n_32548), .B (P1_d_115), .Y (n_11415));
NAND2X1 g124522(.A (n_32544), .B (P1_d_116), .Y (n_11438));
INVX1 g124525(.A (n_10648), .Y (n_11196));
NAND2X1 g124527(.A (n_32548), .B (P1_d_117), .Y (n_11421));
NAND2X1 g124528(.A (n_32548), .B (P1_d_118), .Y (n_11423));
NAND2X1 g124529(.A (n_32544), .B (P1_d_119), .Y (n_11418));
NAND2X1 g124530(.A (n_32550), .B (P1_d_120), .Y (n_11430));
NAND2X1 g124534(.A (n_32548), .B (P1_d_122), .Y (n_11671));
NAND2X1 g124535(.A (n_32544), .B (P1_d_123), .Y (n_11411));
NAND2X1 g124536(.A (n_32550), .B (P1_d_124), .Y (n_11435));
NAND2X1 g124537(.A (n_32544), .B (P1_d_125), .Y (n_11420));
NAND2X1 g124538(.A (n_32548), .B (P1_d_126), .Y (n_11426));
NAND2X1 g124541(.A (n_32544), .B (P1_d_100), .Y (n_11412));
NAND2X1 g124542(.A (n_32544), .B (P1_d_101), .Y (n_11439));
NAND2X1 g124545(.A (n_32544), .B (P1_d_105), .Y (n_11433));
NAND2X1 g124551(.A (n_10999), .B (P3_d_400), .Y (n_11639));
AND2X1 g124555(.A (n_10999), .B (P3_d_405), .Y (n_11658));
NAND2X1 g124556(.A (n_10999), .B (P3_d_399), .Y (n_11651));
NAND2X1 g124560(.A (n_10999), .B (P3_d_391), .Y (n_11641));
NAND2X1 g124579(.A (n_10999), .B (P3_d_380), .Y (n_11647));
NAND2X1 g124590(.A (n_32544), .B (P1_d_111), .Y (n_10991));
NAND3X1 g124592(.A (n_9404), .B (n_10049), .C (n_28528), .Y(n_10990));
NAND3X1 g124609(.A (n_10989), .B (n_9610), .C (n_9621), .Y (n_11192));
AOI21X1 g124617(.A0 (n_9609), .A1 (P2_d), .B0 (n_10034), .Y(n_10988));
AOI22X1 g124628(.A0 (n_10984), .A1 (n_8074), .B0 (n_14534), .B1(n_10986), .Y (n_10987));
AOI22X1 g124629(.A0 (n_10984), .A1 (addr_451), .B0 (n_14534), .B1(n_10983), .Y (n_10985));
AOI22X1 g124636(.A0 (n_10975), .A1 (n_10981), .B0 (n_21677), .B1(n_10981), .Y (n_10982));
AOI22X1 g124637(.A0 (n_10984), .A1 (n_7833), .B0 (n_14534), .B1(n_10979), .Y (n_10980));
AOI22X1 g124638(.A0 (n_10984), .A1 (addr_453), .B0 (n_14534), .B1(n_10977), .Y (n_10978));
AOI22X1 g124639(.A0 (n_10975), .A1 (n_11155), .B0 (n_21677), .B1(n_11155), .Y (n_10976));
AOI22X1 g124641(.A0 (n_10984), .A1 (addr_461), .B0 (n_14534), .B1(n_10973), .Y (n_10974));
AOI22X1 g124643(.A0 (n_10975), .A1 (n_11160), .B0 (n_21677), .B1(n_11160), .Y (n_10972));
AOI22X1 g124644(.A0 (n_10975), .A1 (n_10973), .B0 (n_21677), .B1(n_10973), .Y (n_10971));
AOI22X1 g124646(.A0 (n_10975), .A1 (n_10969), .B0 (n_21677), .B1(n_10969), .Y (n_10970));
AOI22X1 g124647(.A0 (n_10984), .A1 (addr_450), .B0 (n_14534), .B1(n_10967), .Y (n_10968));
AOI22X1 g124648(.A0 (n_10975), .A1 (n_10979), .B0 (n_21677), .B1(n_10979), .Y (n_10966));
AOI22X1 g124649(.A0 (n_10975), .A1 (n_10967), .B0 (n_21677), .B1(n_10967), .Y (n_10965));
AOI22X1 g124651(.A0 (n_10975), .A1 (n_10977), .B0 (n_21677), .B1(n_10977), .Y (n_10964));
AOI22X1 g124652(.A0 (n_10984), .A1 (n_7841), .B0 (n_14534), .B1(n_10962), .Y (n_10963));
AOI22X1 g124654(.A0 (n_10975), .A1 (n_10960), .B0 (n_21677), .B1(n_10960), .Y (n_10961));
AOI22X1 g124655(.A0 (n_11354), .A1 (n_11573), .B0 (n_11353), .B1(n_11573), .Y (n_10959));
AOI22X1 g124662(.A0 (n_10984), .A1 (addr_452), .B0 (n_14534), .B1(n_10981), .Y (n_10958));
AOI22X1 g124672(.A0 (n_10975), .A1 (n_10962), .B0 (n_21677), .B1(n_10962), .Y (n_10957));
AOI22X1 g124673(.A0 (n_10975), .A1 (n_11157), .B0 (n_21677), .B1(n_11157), .Y (n_10956));
AOI22X1 g124674(.A0 (n_10984), .A1 (addr_447), .B0 (n_14534), .B1(n_10969), .Y (n_10955));
AOI22X1 g124676(.A0 (n_10984), .A1 (n_8079), .B0 (n_14534), .B1(n_10953), .Y (n_10954));
AOI22X1 g124677(.A0 (n_10975), .A1 (n_10951), .B0 (n_21677), .B1(n_10951), .Y (n_10952));
AOI22X1 g124678(.A0 (n_10984), .A1 (n_481), .B0 (n_14534), .B1(n_10960), .Y (n_10950));
AOI22X1 g124679(.A0 (n_10975), .A1 (n_10948), .B0 (n_21677), .B1(n_10948), .Y (n_10949));
AOI22X1 g124680(.A0 (n_10975), .A1 (n_10946), .B0 (n_21677), .B1(n_10946), .Y (n_10947));
AOI22X1 g124681(.A0 (n_10984), .A1 (n_7839), .B0 (n_14534), .B1(n_10946), .Y (n_10945));
AOI22X1 g124682(.A0 (n_10975), .A1 (n_10943), .B0 (n_21677), .B1(n_10943), .Y (n_10944));
AOI22X1 g124683(.A0 (n_10975), .A1 (n_11153), .B0 (n_21677), .B1(n_11153), .Y (n_10942));
AOI22X1 g124684(.A0 (n_10975), .A1 (n_11151), .B0 (n_21677), .B1(n_11151), .Y (n_10941));
AOI22X1 g124685(.A0 (n_10984), .A1 (n_7843), .B0 (n_14534), .B1(n_10948), .Y (n_10940));
AOI22X1 g124686(.A0 (n_10975), .A1 (n_10983), .B0 (n_21677), .B1(n_10983), .Y (n_10939));
AOI22X1 g124687(.A0 (n_10975), .A1 (n_10986), .B0 (n_21677), .B1(n_10986), .Y (n_10938));
AOI22X1 g124689(.A0 (n_10984), .A1 (n_628), .B0 (n_14534), .B1(n_10943), .Y (n_10937));
AOI22X1 g124692(.A0 (n_10975), .A1 (n_10953), .B0 (n_21677), .B1(n_10953), .Y (n_10936));
AOI22X1 g124693(.A0 (n_10984), .A1 (n_8083), .B0 (n_14534), .B1(n_10951), .Y (n_10935));
NAND2X1 g124807(.A (n_10932), .B (n_11831), .Y (n_10934));
NAND2X1 g124808(.A (n_10932), .B (n_11829), .Y (n_10933));
NAND2X1 g124809(.A (n_10932), .B (n_11607), .Y (n_10931));
NAND2X1 g124810(.A (n_10932), .B (n_11605), .Y (n_10930));
NAND2X1 g124811(.A (n_10932), .B (n_11821), .Y (n_10929));
INVX2 g124819(.A (n_10927), .Y (n_11399));
NAND2X1 g124824(.A (n_10925), .B (n_11155), .Y (n_10926));
NAND2X1 g124829(.A (n_10932), .B (n_11588), .Y (n_10924));
NAND2X1 g124830(.A (n_10932), .B (n_11817), .Y (n_10923));
NAND2X1 g124836(.A (n_10925), .B (n_11151), .Y (n_10922));
NAND2X1 g124839(.A (n_10932), .B (n_11826), .Y (n_10921));
NAND2X1 g124841(.A (n_10932), .B (n_11599), .Y (n_10920));
NAND2X1 g124845(.A (n_10932), .B (n_11594), .Y (n_10919));
NAND2X1 g124849(.A (n_10917), .B (n_11814), .Y (n_10918));
NAND2X1 g124850(.A (n_10917), .B (n_11811), .Y (n_10916));
NAND2X1 g124851(.A (n_10917), .B (n_11809), .Y (n_10915));
NAND2X1 g124852(.A (n_10917), .B (n_11807), .Y (n_10914));
NAND2X1 g124855(.A (n_10925), .B (n_11157), .Y (n_10913));
NAND2X1 g124857(.A (n_10932), .B (n_11823), .Y (n_10912));
NAND2X1 g124861(.A (n_10925), .B (n_11153), .Y (n_10911));
NAND2X1 g124863(.A (n_10932), .B (n_11601), .Y (n_10910));
NAND2X1 g124866(.A (n_10932), .B (n_11592), .Y (n_10909));
NAND2X1 g124870(.A (n_10932), .B (n_11819), .Y (n_10908));
NAND2X1 g124871(.A (n_10932), .B (n_11834), .Y (n_10907));
NAND2X1 g124872(.A (n_10925), .B (n_11160), .Y (n_10906));
INVX2 g124896(.A (n_10905), .Y (n_11407));
INVX2 g124897(.A (n_10905), .Y (n_11410));
AOI21X1 g124914(.A0 (n_9998), .A1 (n_8981), .B0 (n_991), .Y(n_10903));
INVX1 g124942(.A (n_11610), .Y (n_13748));
INVX1 g125009(.A (n_11356), .Y (n_13761));
CLKBUFX1 g125010(.A (n_11356), .Y (n_11586));
NAND2X1 g125202(.A (n_9001), .B (n_10779), .Y (n_10901));
OR2X1 g125206(.A (n_14351), .B (n_20864), .Y (n_11615));
AOI21X1 g125213(.A0 (n_8927), .A1 (n_23138), .B0 (n_9676), .Y(n_10899));
AOI22X1 g125219(.A0 (n_10573), .A1 (n_10897), .B0 (n_8207), .B1(n_8946), .Y (n_10898));
AOI22X1 g125220(.A0 (n_10573), .A1 (n_10893), .B0 (n_3372), .B1(n_8946), .Y (n_32561));
AOI22X1 g125223(.A0 (n_10573), .A1 (n_10886), .B0 (n_10885), .B1(n_8946), .Y (n_10887));
AOI22X1 g125226(.A0 (n_10573), .A1 (n_3470), .B0 (n_8946), .B1(n_7515), .Y (n_10884));
AOI22X1 g125229(.A0 (n_10573), .A1 (n_3416), .B0 (n_10880), .B1(n_8946), .Y (n_10882));
AOI22X1 g125230(.A0 (n_10573), .A1 (n_4561), .B0 (n_7546), .B1(n_8946), .Y (n_10879));
NAND2X1 g125244(.A (n_9014), .B (n_10046), .Y (n_10875));
INVX1 g125295(.A (n_10583), .Y (n_10874));
INVX1 g125300(.A (n_10580), .Y (n_10873));
AOI22X1 g125308(.A0 (n_11360), .A1 (n_33784), .B0 (n_14743), .B1(addr_425), .Y (n_10872));
AOI22X1 g125311(.A0 (n_11357), .A1 (n_33784), .B0 (n_14743), .B1(n_482), .Y (n_10871));
AOI22X1 g125322(.A0 (n_10573), .A1 (n_4213), .B0 (n_7706), .B1(n_8946), .Y (n_10868));
AOI22X1 g125323(.A0 (n_10573), .A1 (P1_reg2[14] ), .B0 (n_7575), .B1(n_8946), .Y (n_10865));
AOI22X1 g125325(.A0 (n_10573), .A1 (n_4824), .B0 (n_3105), .B1(n_8946), .Y (n_10862));
INVX1 g125330(.A (n_10569), .Y (n_10860));
AOI22X1 g125335(.A0 (n_10573), .A1 (n_10858), .B0 (n_3184), .B1(n_8946), .Y (n_10859));
AOI22X1 g125337(.A0 (n_20218), .A1 (n_3259), .B0 (n_8946), .B1(n_10854), .Y (n_10856));
INVX1 g125339(.A (n_10561), .Y (n_10853));
INVX1 g125342(.A (n_10665), .Y (n_10852));
AOI22X1 g125347(.A0 (n_18289), .A1 (n_4367), .B0 (n_3100), .B1(n_10848), .Y (n_10851));
AOI22X1 g125349(.A0 (n_18289), .A1 (P2_reg2[15] ), .B0 (n_8467), .B1(n_10848), .Y (n_10847));
AOI22X1 g125355(.A0 (n_18289), .A1 (P2_reg2[1] ), .B0 (n_10848), .B1(P2_reg3[1] ), .Y (n_10843));
AOI22X1 g125370(.A0 (n_11584), .A1 (n_25220), .B0 (n_10573), .B1(addr_426), .Y (n_10841));
AOI22X1 g125371(.A0 (n_11573), .A1 (n_33738), .B0 (n_15110), .B1(n_10838), .Y (n_10840));
AOI22X1 g125373(.A0 (n_11573), .A1 (n_21328), .B0 (n_11138), .B1(n_10838), .Y (n_10839));
INVX1 g128377(.A (n_18496), .Y (n_11218));
INVX1 g125391(.A (n_10550), .Y (n_10837));
INVX1 g125426(.A (n_11181), .Y (n_10836));
INVX1 g125428(.A (n_11339), .Y (n_10834));
NAND2X1 g125432(.A (n_10573), .B (n_4590), .Y (n_10833));
NAND2X1 g125433(.A (n_10573), .B (P1_reg2[16] ), .Y (n_10831));
NAND2X1 g125453(.A (n_10573), .B (n_4230), .Y (n_10829));
INVX1 g128366(.A (n_17261), .Y (n_10826));
NAND2X1 g125499(.A (n_10573), .B (n_3105), .Y (n_10825));
NAND2X1 g125501(.A (n_10573), .B (n_10822), .Y (n_10823));
NOR2X1 g125503(.A (n_15749), .B (n_10821), .Y (n_32374));
NAND2X1 g125529(.A (n_34708), .B (n_12670), .Y (n_12426));
NOR2X1 g125531(.A (n_9983), .B (n_991), .Y (n_11086));
INVX1 g125825(.A (n_33494), .Y (n_25119));
CLKBUFX1 g125872(.A (n_10808), .Y (n_28275));
INVX1 g125879(.A (n_34752), .Y (n_26106));
INVX1 g125884(.A (n_24526), .Y (n_30138));
CLKBUFX1 gbuf_d_700(.A(n_9908), .Y(d_out_700));
CLKBUFX1 gbuf_qn_700(.A(qn_in_700), .Y(wr_1));
NAND2X1 g125948(.A (n_30399), .B (n_12670), .Y (n_10800));
NAND2X1 g125949(.A (n_10472), .B (n_34651), .Y (n_11181));
NAND2X1 g125950(.A (n_10799), .B (n_11079), .Y (n_11339));
INVX1 g126060(.A (n_10796), .Y (n_10797));
NOR2X1 g126072(.A (n_9684), .B (n_10794), .Y (n_10795));
NOR2X1 g126088(.A (n_11295), .B (n_10474), .Y (n_10793));
INVX4 g126210(.A (n_10790), .Y (n_29925));
INVX2 g126217(.A (n_10790), .Y (n_25988));
INVX1 g126220(.A (n_34708), .Y (n_27158));
INVX1 g126223(.A (n_34708), .Y (n_10785));
INVX4 g126230(.A (n_34709), .Y (n_27696));
INVX1 g126478(.A (n_10779), .Y (n_28915));
INVX1 g126484(.A (n_10776), .Y (n_25636));
INVX1 g126488(.A (n_9983), .Y (n_29908));
MX2X1 g126760(.A (n_32856), .B (datao_1[1] ), .S0 (n_7860), .Y(n_10774));
INVX1 g126765(.A (n_10771), .Y (n_11548));
NAND2X1 g126773(.A (n_11401), .B (n_32827), .Y (n_10770));
INVX1 g126783(.A (n_10769), .Y (n_11534));
NAND2X1 g126786(.A (n_9754), .B (n_10768), .Y (n_11065));
NAND2X1 g126788(.A (n_10767), .B (n_10330), .Y (n_11063));
INVX1 g126797(.A (n_10764), .Y (n_10765));
NOR2X1 g126816(.A (n_9798), .B (n_10315), .Y (n_11306));
NAND2X1 g126826(.A (n_9760), .B (n_10490), .Y (n_10763));
NAND2X1 g126833(.A (n_16446), .B (n_17916), .Y (n_11770));
NAND2X1 g126844(.A (n_10760), .B (n_12953), .Y (n_10761));
NAND2X1 g126849(.A (n_9814), .B (n_34706), .Y (n_10759));
NAND2X1 g126852(.A (n_10758), .B (n_10757), .Y (n_11302));
NAND2X1 g126862(.A (n_16163), .B (n_11555), .Y (n_11775));
NAND2X1 g126866(.A (n_16904), .B (n_10756), .Y (n_11774));
NAND2X2 g126870(.A (n_10755), .B (n_10754), .Y (n_11301));
NAND2X1 g126871(.A (n_11089), .B (n_17955), .Y (n_11300));
NAND2X1 g126872(.A (n_18584), .B (n_9741), .Y (n_11304));
NAND2X1 g126881(.A (n_10287), .B (n_9761), .Y (n_11296));
INVX1 g126889(.A (n_10753), .Y (n_11210));
NAND2X2 g126892(.A (n_17916), .B (n_10752), .Y (n_11772));
NAND3X1 g126917(.A (n_9693), .B (n_8910), .C (n_34650), .Y (n_16460));
NOR2X1 g126952(.A (n_8829), .B (n_10451), .Y (n_11050));
NOR2X1 g126958(.A (n_10317), .B (n_9292), .Y (n_11048));
NAND2X1 g126962(.A (n_9953), .B (n_13106), .Y (n_10747));
NAND2X1 g126994(.A (n_9771), .B (n_6806), .Y (n_10746));
INVX2 g127002(.A (n_10745), .Y (n_18164));
NOR2X1 g127251(.A (n_9871), .B (n_6763), .Y (n_10744));
NAND3X1 g127298(.A (n_10736), .B (n_13375), .C (n_8884), .Y(n_10743));
AOI22X1 g128994(.A0 (n_10696), .A1 (n_10740), .B0 (n_5301), .B1(n_10676), .Y (n_10741));
NAND3X1 g127351(.A (n_12739), .B (n_13724), .C (n_8884), .Y(n_10739));
NAND3X1 g127365(.A (n_10736), .B (n_13378), .C (n_8884), .Y(n_10737));
NAND3X1 g127370(.A (n_10736), .B (n_13327), .C (n_8884), .Y(n_10734));
INVX1 g127617(.A (n_17467), .Y (n_11036));
INVX1 g127686(.A (n_18536), .Y (n_11034));
INVX1 g127704(.A (n_17392), .Y (n_11033));
INVX1 g127771(.A (n_9785), .Y (n_11030));
CLKBUFX1 g127940(.A (n_16829), .Y (n_11987));
INVX1 g127995(.A (n_10322), .Y (n_11275));
NOR2X1 g128028(.A (n_9212), .B (n_9689), .Y (n_16750));
NAND2X1 g126946(.A (n_10718), .B (n_10717), .Y (n_11052));
INVX1 g128163(.A (n_10716), .Y (n_11791));
INVX1 g128184(.A (n_10712), .Y (n_10713));
INVX1 g128187(.A (n_10712), .Y (n_11269));
INVX1 g128195(.A (n_12992), .Y (n_10711));
INVX1 g128202(.A (n_10710), .Y (n_11022));
INVX1 g128224(.A (n_11058), .Y (n_11556));
NAND2X1 g128234(.A (n_9207), .B (n_9691), .Y (n_11037));
NOR2X1 g128261(.A (n_10709), .B (n_10708), .Y (n_17348));
INVX1 g128278(.A (n_10706), .Y (n_11256));
INVX2 g128300(.A (n_16040), .Y (n_11278));
INVX1 g128322(.A (n_10497), .Y (n_16161));
INVX1 g128337(.A (n_10792), .Y (n_11249));
INVX2 g128384(.A (n_9036), .Y (n_11280));
INVX2 g128490(.A (n_9720), .Y (n_11797));
INVX1 g128516(.A (n_12003), .Y (n_11012));
INVX1 g128565(.A (n_10292), .Y (n_16429));
INVX1 g128596(.A (n_18001), .Y (n_11276));
NAND2X1 g128690(.A (n_9679), .B (n_7876), .Y (n_11374));
NAND2X1 g128840(.A (n_9631), .B (n_7847), .Y (n_11388));
NAND2X1 g128841(.A (n_9657), .B (n_7877), .Y (n_11386));
NAND2X1 g128842(.A (n_9671), .B (n_7602), .Y (n_11384));
NAND2X1 g128843(.A (n_9673), .B (n_7655), .Y (n_11380));
NAND2X1 g128844(.A (n_9669), .B (n_7654), .Y (n_11378));
NAND2X1 g128845(.A (n_9659), .B (n_7870), .Y (n_11376));
NAND2X1 g128906(.A (n_9665), .B (n_7829), .Y (n_11372));
NAND2X1 g128907(.A (n_9662), .B (n_7964), .Y (n_11391));
NAND2X1 g128909(.A (n_9687), .B (n_7647), .Y (n_11370));
NAND2X1 g128910(.A (n_9682), .B (n_7612), .Y (n_11368));
NAND2X1 g128911(.A (n_10014), .B (n_7873), .Y (n_11366));
NAND2X1 g128912(.A (n_9666), .B (n_7651), .Y (n_11364));
NAND2X1 g128913(.A (n_9674), .B (n_7649), .Y (n_11362));
NAND2X1 g128916(.A (n_9654), .B (n_7648), .Y (n_11382));
AOI22X1 g128992(.A0 (n_10696), .A1 (n_3063), .B0 (n_4078), .B1(n_10676), .Y (n_10697));
AOI22X1 g128993(.A0 (n_10696), .A1 (n_3165), .B0 (n_4631), .B1(n_10676), .Y (n_10693));
AOI22X1 g128995(.A0 (n_10696), .A1 (n_3176), .B0 (n_4889), .B1(n_10676), .Y (n_10691));
INVX1 g128035(.A (n_10689), .Y (n_17337));
AOI22X1 g129118(.A0 (n_10696), .A1 (n_4320), .B0 (n_6074), .B1(n_10676), .Y (n_10688));
AOI22X1 g129119(.A0 (n_10696), .A1 (n_3862), .B0 (n_6064), .B1(n_10676), .Y (n_10686));
AOI22X1 g129122(.A0 (n_10696), .A1 (n_32445), .B0 (n_6135), .B1(n_10676), .Y (n_10684));
AOI22X1 g129123(.A0 (n_10696), .A1 (n_4735), .B0 (n_6186), .B1(n_10676), .Y (n_10682));
AOI22X1 g129124(.A0 (n_7641), .A1 (n_32386), .B0 (n_6327), .B1(n_10676), .Y (n_10680));
AOI22X1 g129128(.A0 (n_10671), .A1 (n_3583), .B0 (n_5284), .B1(n_10676), .Y (n_10678));
AOI22X1 g129129(.A0 (n_7641), .A1 (n_4133), .B0 (n_5610), .B1(n_10676), .Y (n_10675));
AOI22X1 g129130(.A0 (n_10671), .A1 (n_3854), .B0 (n_6035), .B1(n_10676), .Y (n_10672));
NOR2X1 g126876(.A (n_10755), .B (n_10754), .Y (n_10667));
INVX1 g128305(.A (n_10666), .Y (n_11503));
AOI22X1 g125343(.A0 (n_18289), .A1 (P2_reg2[12] ), .B0 (n_8185), .B1(n_10848), .Y (n_10665));
INVX2 g128586(.A (n_9700), .Y (n_11010));
INVX1 g127634(.A (n_16011), .Y (n_17182));
INVX1 g128572(.A (n_10658), .Y (n_19666));
AOI22X1 g129121(.A0 (n_10696), .A1 (n_10656), .B0 (n_6072), .B1(n_10676), .Y (n_10657));
INVX2 g124906(.A (n_33412), .Y (n_10655));
AOI22X1 g125239(.A0 (n_18289), .A1 (n_10653), .B0 (n_8447), .B1(n_18909), .Y (n_32223));
INVX2 g124820(.A (n_10262), .Y (n_10927));
CLKBUFX3 g128367(.A (n_16068), .Y (n_17261));
NAND2X1 g124511(.A (n_32543), .B (P1_d_108), .Y (n_11417));
NAND2X1 g124517(.A (n_32543), .B (P1_d_113), .Y (n_11200));
NAND2X1 g124520(.A (n_32543), .B (P1_d_114), .Y (n_11450));
NAND3X1 g124526(.A (n_7787), .B (n_9146), .C (n_9032), .Y (n_10648));
NAND2X1 g124532(.A (n_32543), .B (P1_d_121), .Y (n_11199));
NAND2X1 g124539(.A (n_32543), .B (P1_d_99), .Y (n_11447));
NAND2X1 g124540(.A (n_32543), .B (P1_d_127), .Y (n_11202));
NAND2X1 g124543(.A (n_32543), .B (P1_d_102), .Y (n_11205));
NAND2X1 g124544(.A (n_32543), .B (P1_d_104), .Y (n_11201));
NAND2X1 g124566(.A (n_32543), .B (P1_d_128), .Y (n_11432));
NAND2X1 g124601(.A (n_32543), .B (P1_d_106), .Y (n_11206));
NAND2X1 g124805(.A (n_9613), .B (n_11584), .Y (n_10647));
NAND2X1 g124825(.A (n_10644), .B (n_10973), .Y (n_10646));
NAND2X1 g124832(.A (n_10644), .B (n_10960), .Y (n_10645));
NAND2X1 g124837(.A (n_10644), .B (n_10986), .Y (n_10643));
NAND2X1 g124844(.A (n_10917), .B (n_11573), .Y (n_10642));
NAND2X1 g124862(.A (n_10644), .B (n_10969), .Y (n_10641));
NAND2X1 g124865(.A (n_10644), .B (n_10943), .Y (n_10640));
NAND2X1 g124868(.A (n_10644), .B (n_10953), .Y (n_10639));
NAND2X1 g124869(.A (n_10644), .B (n_10951), .Y (n_10638));
NAND2X1 g124873(.A (n_9613), .B (n_11805), .Y (n_10637));
NAND2X1 g125207(.A (n_10624), .B (n_8413), .Y (n_10635));
BUFX1 g124895(.A (n_10634), .Y (n_11208));
INVX2 g124898(.A (n_10634), .Y (n_10905));
INVX1 g124907(.A (n_33412), .Y (n_11194));
INVX1 g124908(.A (n_33412), .Y (n_11195));
AOI21X1 g124915(.A0 (n_9495), .A1 (n_8325), .B0 (n_7967), .Y(n_10631));
NAND2X1 g124938(.A (n_33807), .B (n_10629), .Y (n_10630));
NAND2X2 g124944(.A (n_35043), .B (n_9983), .Y (n_11610));
NAND2X1 g124949(.A (n_11575), .B (n_11360), .Y (n_10628));
NAND2X1 g124960(.A (n_11575), .B (n_11357), .Y (n_10627));
NAND3X1 g125011(.A (n_8718), .B (n_33807), .C (n_34719), .Y(n_11356));
NAND3X1 g125048(.A (n_33505), .B (n_29381), .C (n_33807), .Y(n_22244));
NAND2X1 g125083(.A (n_11575), .B (n_11596), .Y (n_10626));
NAND2X1 g125112(.A (n_10624), .B (n_8687), .Y (n_10625));
NAND3X1 g125205(.A (n_8671), .B (n_33340), .C (n_8668), .Y (n_10623));
NAND2X1 g125214(.A (n_9511), .B (n_9483), .Y (n_11183));
OAI21X1 g125215(.A0 (n_3493), .A1 (n_8309), .B0 (n_9528), .Y(n_10622));
OAI21X1 g125216(.A0 (n_8309), .A1 (P3_reg3[3] ), .B0 (n_9524), .Y(n_10621));
AOI22X1 g125225(.A0 (n_18289), .A1 (P2_reg2[10] ), .B0 (n_10617),.B1 (n_18909), .Y (n_10619));
NAND2X1 g125227(.A (n_9016), .B (n_9532), .Y (n_10616));
AOI22X1 g125231(.A0 (n_18289), .A1 (n_10613), .B0 (n_10612), .B1(n_10848), .Y (n_10615));
AOI22X1 g125233(.A0 (n_18289), .A1 (n_10610), .B0 (n_9209), .B1(n_10848), .Y (n_10611));
AOI22X1 g125235(.A0 (n_18289), .A1 (n_10607), .B0 (n_9512), .B1(n_10848), .Y (n_10608));
AOI22X1 g125236(.A0 (n_18289), .A1 (n_10604), .B0 (n_9345), .B1(n_18909), .Y (n_10606));
AOI22X1 g125237(.A0 (n_18289), .A1 (n_10602), .B0 (n_10601), .B1(n_10848), .Y (n_10603));
AOI22X1 g125240(.A0 (n_18289), .A1 (P2_reg2[3] ), .B0 (n_10848), .B1(n_7475), .Y (n_10600));
NAND2X1 g125241(.A (n_9517), .B (n_9531), .Y (n_10597));
AOI22X1 g125242(.A0 (n_18289), .A1 (n_3724), .B0 (n_10594), .B1(n_18909), .Y (n_10596));
AOI22X1 g125243(.A0 (n_18289), .A1 (n_4344), .B0 (n_8193), .B1(n_18909), .Y (n_10593));
NAND2X1 g125245(.A (n_9509), .B (n_9527), .Y (n_10590));
OAI21X1 g125248(.A0 (n_3573), .A1 (n_8309), .B0 (n_9525), .Y(n_10589));
OAI21X1 g125253(.A0 (n_3269), .A1 (n_8309), .B0 (n_9523), .Y(n_10588));
INVX1 g125291(.A (n_10102), .Y (n_10587));
AOI22X1 g125294(.A0 (n_18289), .A1 (n_4475), .B0 (n_8458), .B1(n_18909), .Y (n_10586));
AOI22X1 g125296(.A0 (n_11138), .A1 (P3_reg2[13] ), .B0 (n_10582),.B1 (n_19108), .Y (n_10583));
INVX1 g125297(.A (n_10098), .Y (n_10581));
AOI22X1 g125301(.A0 (n_11138), .A1 (n_13498), .B0 (n_10578), .B1(n_19108), .Y (n_10580));
INVX1 g125304(.A (n_10095), .Y (n_10577));
INVX1 g125306(.A (n_10094), .Y (n_10576));
AOI22X1 g125309(.A0 (n_11360), .A1 (n_25082), .B0 (n_10573), .B1(addr_425), .Y (n_10575));
AOI22X1 g125312(.A0 (n_11357), .A1 (n_25082), .B0 (n_10573), .B1(n_482), .Y (n_10574));
INVX1 g125313(.A (n_10093), .Y (n_10571));
INVX1 g125326(.A (n_10092), .Y (n_10570));
AOI22X1 g125331(.A0 (n_10573), .A1 (P1_reg2[1] ), .B0 (n_8946), .B1(n_10566), .Y (n_10569));
AOI22X1 g125338(.A0 (n_18289), .A1 (n_10563), .B0 (n_10848), .B1(n_10562), .Y (n_10565));
AOI22X1 g125340(.A0 (n_18289), .A1 (P2_reg2[11] ), .B0 (n_7664), .B1(n_10848), .Y (n_10561));
INVX1 g125350(.A (n_10088), .Y (n_10557));
INVX1 g125357(.A (n_10080), .Y (n_10556));
INVX1 g125359(.A (n_10079), .Y (n_10555));
INVX1 g125361(.A (n_10076), .Y (n_10554));
INVX1 g125366(.A (n_10069), .Y (n_10553));
INVX1 g125379(.A (n_10066), .Y (n_10552));
INVX1 g125386(.A (n_10059), .Y (n_10551));
AOI22X1 g125392(.A0 (n_11138), .A1 (P3_reg2[9] ), .B0 (n_13370), .B1(n_7988), .Y (n_10550));
INVX1 g125393(.A (n_10053), .Y (n_10548));
NAND2X1 g125441(.A (n_20218), .B (P1_reg2[9] ), .Y (n_10545));
NOR2X1 g125514(.A (n_8981), .B (P1_reg3[3] ), .Y (n_10543));
NAND2X1 g125536(.A (n_10504), .B (n_8799), .Y (n_10819));
NAND2X1 g125549(.A (n_9482), .B (n_9995), .Y (n_10542));
INVX4 g125697(.A (n_10023), .Y (n_20304));
INVX1 g125725(.A (n_21703), .Y (n_20727));
INVX4 g125742(.A (n_20399), .Y (n_20112));
INVX1 g125749(.A (n_21365), .Y (n_22139));
INVX1 g125752(.A (n_10525), .Y (n_21333));
INVX1 g125758(.A (n_21365), .Y (n_20473));
INVX1 g125764(.A (n_21365), .Y (n_20490));
INVX1 g125770(.A (n_21374), .Y (n_20478));
INVX1 g125776(.A (n_10525), .Y (n_21658));
INVX1 g125779(.A (n_10525), .Y (n_21694));
INVX1 g125821(.A (n_26662), .Y (n_30355));
INVX1 g125851(.A (n_26528), .Y (n_27564));
INVX1 g125877(.A (n_34752), .Y (n_28636));
INVX1 g125902(.A (n_30291), .Y (n_10517));
AOI21X1 g125935(.A0 (n_33094), .A1 (n_8399), .B0 (n_33713), .Y(n_10514));
NAND2X1 g126037(.A (n_8784), .B (n_9960), .Y (n_10821));
INVX1 g126061(.A (n_9638), .Y (n_10796));
INVX1 g126089(.A (n_10504), .Y (n_10505));
INVX1 g128327(.A (n_9730), .Y (n_12827));
INVX1 g126473(.A (n_28013), .Y (n_10779));
INVX1 g126486(.A (n_25980), .Y (n_10776));
NAND2X2 g128323(.A (n_8761), .B (n_9205), .Y (n_10497));
INVX1 g126766(.A (n_16768), .Y (n_10771));
NAND2X1 g126769(.A (n_9242), .B (n_10490), .Y (n_10491));
NAND2X1 g126772(.A (n_9235), .B (n_34706), .Y (n_10489));
NAND2X1 g126784(.A (n_16096), .B (n_16331), .Y (n_10769));
NOR2X1 g126795(.A (n_16577), .B (n_9624), .Y (n_10487));
NAND2X1 g126798(.A (n_34935), .B (n_10485), .Y (n_10764));
NOR2X1 g126805(.A (n_8803), .B (n_10484), .Y (n_11305));
NOR2X1 g126818(.A (n_9632), .B (n_10482), .Y (n_11002));
NOR2X1 g126819(.A (n_9788), .B (n_9264), .Y (n_11536));
NAND2X1 g126822(.A (n_9262), .B (n_10490), .Y (n_10481));
NAND2X1 g126823(.A (n_9338), .B (n_34706), .Y (n_10480));
NAND2X1 g126827(.A (n_9234), .B (n_34706), .Y (n_10478));
AND2X1 g126836(.A (n_9341), .B (n_10465), .Y (n_10477));
NAND2X1 g126845(.A (n_9152), .B (n_34706), .Y (n_10476));
INVX1 g126847(.A (n_10474), .Y (n_10475));
NOR2X1 g126850(.A (n_8851), .B (n_8830), .Y (n_11088));
INVX1 g128301(.A (n_33227), .Y (n_16040));
INVX2 g126885(.A (n_10472), .Y (n_16452));
INVX1 g126890(.A (n_9959), .Y (n_10753));
INVX1 g126898(.A (n_10794), .Y (n_10470));
NAND2X1 g126906(.A (n_16012), .B (n_17000), .Y (n_10468));
INVX1 g126909(.A (n_10467), .Y (n_18159));
NAND2X1 g126949(.A (n_11092), .B (n_9725), .Y (n_11303));
AND2X1 g126950(.A (n_9346), .B (n_10465), .Y (n_10466));
NAND2X1 g126953(.A (n_9340), .B (n_34706), .Y (n_10464));
NAND2X1 g126954(.A (n_9237), .B (n_6806), .Y (n_10463));
NAND2X1 g126963(.A (n_35314), .B (n_16188), .Y (n_10461));
NAND2X1 g126971(.A (n_9285), .B (n_6806), .Y (n_10460));
NAND2X1 g126976(.A (n_9161), .B (n_10490), .Y (n_10459));
NAND2X1 g126981(.A (n_9334), .B (n_10490), .Y (n_10458));
NAND2X1 g126986(.A (n_9294), .B (n_6806), .Y (n_10457));
NAND2X1 g126989(.A (n_9314), .B (n_10490), .Y (n_10456));
NAND2X1 g126997(.A (n_9249), .B (n_6806), .Y (n_10455));
INVX1 g127003(.A (n_11079), .Y (n_10745));
NAND3X1 g127185(.A (n_10449), .B (n_10452), .C (n_8393), .Y(n_10453));
NAND3X1 g127188(.A (n_10449), .B (P2_reg_106), .C (n_8393), .Y(n_10450));
NOR2X1 g127190(.A (n_9369), .B (n_12755), .Y (n_10448));
NOR2X1 g127193(.A (n_9332), .B (n_9946), .Y (n_10447));
NAND3X1 g127204(.A (n_10736), .B (n_13699), .C (n_8884), .Y(n_10445));
NAND3X1 g127205(.A (n_10449), .B (n_10443), .C (n_8393), .Y(n_10444));
NAND3X1 g127206(.A (n_6478), .B (n_13377), .C (n_8884), .Y (n_10441));
NAND3X1 g127211(.A (n_10736), .B (P3_reg2[29] ), .C (n_8884), .Y(n_10440));
NAND3X1 g127216(.A (n_12611), .B (n_10435), .C (n_8393), .Y(n_10436));
NOR2X1 g127217(.A (n_9263), .B (n_9946), .Y (n_10433));
NOR2X1 g127220(.A (n_9232), .B (n_10414), .Y (n_10432));
NAND3X1 g127221(.A (n_10736), .B (n_13203), .C (n_8884), .Y(n_10431));
NAND3X1 g127223(.A (n_10736), .B (n_13695), .C (n_8884), .Y(n_10429));
NOR2X1 g127224(.A (n_9366), .B (n_10399), .Y (n_10427));
NAND3X1 g127226(.A (n_12611), .B (P2_reg1[4] ), .C (n_8393), .Y(n_10426));
NAND3X1 g127233(.A (n_34706), .B (n_9634), .C (n_8393), .Y (n_10423));
NAND3X1 g127236(.A (n_12606), .B (P2_reg2[16] ), .C (n_8393), .Y(n_10420));
NAND3X1 g127238(.A (n_10449), .B (P2_reg1[1] ), .C (n_8393), .Y(n_10418));
NOR2X1 g127249(.A (n_9349), .B (n_12755), .Y (n_10416));
NOR2X1 g127252(.A (n_9297), .B (n_10414), .Y (n_10415));
NAND3X1 g127255(.A (n_12606), .B (P2_reg2[2] ), .C (n_8393), .Y(n_10413));
NAND3X1 g127261(.A (n_34706), .B (n_10562), .C (n_8393), .Y(n_10409));
NAND3X1 g127263(.A (n_10449), .B (n_8185), .C (n_8393), .Y (n_10407));
NAND3X1 g127264(.A (n_10449), .B (n_2909), .C (n_8393), .Y (n_10406));
NAND3X1 g127266(.A (n_10449), .B (n_8467), .C (n_8393), .Y (n_10405));
NAND3X1 g127268(.A (n_10449), .B (n_8458), .C (n_8393), .Y (n_10403));
NAND3X1 g127270(.A (n_10449), .B (n_8164), .C (n_8393), .Y (n_10402));
NAND3X1 g127271(.A (n_10449), .B (n_3191), .C (n_8393), .Y (n_10401));
NOR2X1 g127279(.A (n_9361), .B (n_10399), .Y (n_10400));
NAND3X1 g127280(.A (n_10449), .B (n_3100), .C (n_8393), .Y (n_10398));
NAND3X1 g127281(.A (n_10449), .B (n_1183), .C (n_8393), .Y (n_10397));
NOR2X1 g127282(.A (n_9357), .B (n_12926), .Y (n_10395));
NAND3X1 g127288(.A (n_10449), .B (n_7664), .C (n_8393), .Y (n_10394));
NOR2X1 g127290(.A (n_9348), .B (n_12917), .Y (n_10393));
NAND3X1 g127292(.A (n_6478), .B (P3_reg3[2] ), .C (n_8884), .Y(n_10392));
NOR2X1 g127295(.A (n_9363), .B (n_12755), .Y (n_10390));
NAND3X1 g127304(.A (n_6478), .B (n_13735), .C (n_8884), .Y (n_10389));
NOR2X1 g127305(.A (n_9355), .B (n_10342), .Y (n_10385));
NAND3X1 g127308(.A (n_12739), .B (n_13689), .C (n_8884), .Y(n_10384));
NAND3X1 g127310(.A (n_12606), .B (n_3709), .C (n_8393), .Y (n_10383));
NAND3X1 g127311(.A (n_12606), .B (P2_reg1[5] ), .C (n_8393), .Y(n_10381));
NAND3X1 g127312(.A (n_12739), .B (n_13687), .C (n_8884), .Y(n_10379));
NAND3X1 g127317(.A (n_12611), .B (P2_reg1[2] ), .C (n_8393), .Y(n_10378));
NAND3X1 g127324(.A (n_6478), .B (n_13675), .C (n_8884), .Y (n_10376));
NAND3X1 g127325(.A (n_34706), .B (P2_reg3[1] ), .C (n_8393), .Y(n_10375));
NOR2X1 g127328(.A (n_9372), .B (n_12755), .Y (n_10373));
NAND3X1 g127332(.A (n_6478), .B (n_13698), .C (n_8884), .Y (n_10372));
NOR2X1 g127334(.A (n_9419), .B (n_12755), .Y (n_10370));
NOR2X1 g127337(.A (n_9356), .B (n_12755), .Y (n_10369));
NAND3X1 g127340(.A (n_6478), .B (n_524), .C (n_8884), .Y (n_10368));
NAND3X1 g127341(.A (n_10736), .B (n_13692), .C (n_8884), .Y(n_10367));
NOR2X1 g127343(.A (n_9374), .B (n_12755), .Y (n_10366));
NAND3X1 g127345(.A (n_12611), .B (n_10363), .C (n_8393), .Y(n_10364));
NAND3X1 g127346(.A (n_10736), .B (n_13340), .C (n_8884), .Y(n_10362));
NOR2X1 g127347(.A (n_9035), .B (n_12755), .Y (n_10361));
NOR2X1 g127348(.A (n_9354), .B (n_12755), .Y (n_10360));
NOR2X1 g127352(.A (n_9352), .B (n_10399), .Y (n_10358));
NAND3X1 g127353(.A (n_12739), .B (n_13673), .C (n_8884), .Y(n_10357));
NAND3X1 g127354(.A (n_12739), .B (n_13690), .C (n_8884), .Y(n_10356));
NAND3X1 g127355(.A (n_10736), .B (n_13370), .C (n_8884), .Y(n_10355));
NOR2X1 g127360(.A (n_9368), .B (n_12755), .Y (n_10354));
NAND3X1 g127363(.A (n_6478), .B (n_13697), .C (n_8884), .Y (n_10352));
NOR2X1 g127366(.A (n_9350), .B (n_12755), .Y (n_10351));
NAND3X1 g127367(.A (n_31495), .B (P3_reg3[0] ), .C (n_9373), .Y(n_10349));
NOR2X1 g127368(.A (n_9358), .B (n_12755), .Y (n_10348));
NAND3X1 g127371(.A (n_6478), .B (P3_reg1[26] ), .C (n_8884), .Y(n_10346));
NAND3X1 g127373(.A (n_10736), .B (n_13711), .C (n_8884), .Y(n_10345));
NOR2X1 g127375(.A (n_9364), .B (n_10342), .Y (n_10343));
CLKBUFX1 g127660(.A (n_17916), .Y (n_12986));
INVX1 g127677(.A (n_10335), .Y (n_12703));
INVX1 g127706(.A (n_10272), .Y (n_10334));
CLKBUFX1 g128196(.A (n_11246), .Y (n_12992));
CLKBUFX1 g127822(.A (n_16446), .Y (n_13071));
CLKBUFX1 g127854(.A (n_10754), .Y (n_11285));
INVX1 g127941(.A (n_16251), .Y (n_16829));
INVX2 g128188(.A (n_10325), .Y (n_10712));
NAND2X1 g127971(.A (n_8393), .B (n_34700), .Y (n_10324));
INVX2 g128017(.A (n_10320), .Y (n_17909));
INVX1 g128037(.A (n_10319), .Y (n_10689));
INVX1 g128038(.A (n_10319), .Y (n_10318));
INVX1 g128050(.A (n_10317), .Y (n_10669));
INVX1 g128072(.A (n_10315), .Y (n_17468));
INVX1 g128114(.A (n_10312), .Y (n_12532));
INVX1 g128164(.A (n_10309), .Y (n_10716));
INVX1 g128203(.A (n_10767), .Y (n_10710));
INVX1 g128225(.A (n_17351), .Y (n_11058));
INVX1 g128306(.A (n_16167), .Y (n_10666));
INVX1 g128315(.A (n_16008), .Y (n_16165));
INVX1 g128338(.A (n_10303), .Y (n_10792));
INVX2 g128368(.A (n_15909), .Y (n_16068));
INVX1 g128380(.A (n_17380), .Y (n_10299));
INVX2 g128146(.A (n_16182), .Y (n_16174));
CLKBUFX1 g128517(.A (n_17262), .Y (n_12003));
INVX1 g128536(.A (n_10755), .Y (n_11055));
INVX1 g128545(.A (n_10757), .Y (n_10699));
CLKBUFX1 g128554(.A (n_16968), .Y (n_11559));
NAND3X1 g128566(.A (n_9210), .B (n_7830), .C (n_7912), .Y (n_10292));
INVX1 g128573(.A (n_10756), .Y (n_10658));
INVX2 g128597(.A (n_10768), .Y (n_18001));
NAND2X1 g128680(.A (n_9197), .B (n_7452), .Y (n_11814));
NAND2X1 g128681(.A (n_9190), .B (n_7454), .Y (n_11809));
NAND2X1 g128908(.A (n_9194), .B (n_7455), .Y (n_11807));
NAND2X1 g128915(.A (n_9173), .B (n_7458), .Y (n_11811));
INVX2 g126215(.A (n_28926), .Y (n_10790));
AOI22X1 g128950(.A0 (n_8739), .A1 (n_7217), .B0 (n_7641), .B1(n_32509), .Y (n_10289));
INVX1 g128106(.A (n_10287), .Y (n_17480));
AOI22X1 g129131(.A0 (n_4184), .A1 (n_9676), .B0 (n_10671), .B1(n_2872), .Y (n_10286));
NAND2X1 g126904(.A (n_9342), .B (n_34706), .Y (n_10283));
NOR2X1 g127358(.A (n_9362), .B (n_10342), .Y (n_10279));
NOR2X1 g126814(.A (n_17007), .B (n_9286), .Y (n_11076));
AOI21X1 g124616(.A0 (n_8695), .A1 (P1_d), .B0 (n_7788), .Y (n_10278));
NAND2X1 g126777(.A (n_9288), .B (n_34706), .Y (n_10277));
INVX2 g125868(.A (n_10276), .Y (n_10808));
INVX1 g125885(.A (n_34752), .Y (n_24526));
INVX1 g127773(.A (n_10275), .Y (n_10274));
INVX4 g125723(.A (n_10020), .Y (n_21703));
INVX1 g127723(.A (n_10273), .Y (n_12943));
INVX1 g127705(.A (n_10272), .Y (n_17392));
INVX1 g127707(.A (n_10272), .Y (n_10271));
INVX1 g127687(.A (n_16904), .Y (n_18536));
INVX1 g127672(.A (n_10270), .Y (n_11057));
OAI21X1 g125251(.A0 (n_9313), .A1 (n_8309), .B0 (n_9030), .Y(n_10268));
INVX1 g128412(.A (n_10267), .Y (n_12232));
NAND2X1 g124803(.A (n_10644), .B (n_10967), .Y (n_10264));
NAND2X1 g124812(.A (n_10644), .B (n_10946), .Y (n_10263));
NAND3X1 g124821(.A (n_35384), .B (n_10251), .C (n_10253), .Y(n_10262));
NAND2X1 g124822(.A (n_10644), .B (n_10983), .Y (n_10261));
NAND2X1 g124828(.A (n_10644), .B (n_10977), .Y (n_10260));
NAND2X1 g124834(.A (n_10644), .B (n_10962), .Y (n_10259));
NAND2X1 g124856(.A (n_10644), .B (n_10981), .Y (n_10258));
NAND2X1 g124858(.A (n_10644), .B (n_10979), .Y (n_10257));
NAND2X1 g124867(.A (n_10644), .B (n_10948), .Y (n_10256));
NAND2X1 g124890(.A (n_9145), .B (P3_d), .Y (n_10254));
NAND3X1 g124899(.A (n_35385), .B (n_10253), .C (n_10251), .Y(n_10634));
CLKBUFX3 g124901(.A (n_33404), .Y (n_10999));
NAND2X1 g124927(.A (n_32400), .B (P2_d_378), .Y (n_10249));
NAND2X1 g124946(.A (n_14550), .B (n_10247), .Y (n_10248));
AND2X1 g124953(.A (n_14550), .B (n_10245), .Y (n_10246));
AND2X1 g124955(.A (n_14550), .B (n_3337), .Y (n_10244));
NAND2X1 g124956(.A (n_14550), .B (n_4215), .Y (n_10242));
NAND2X1 g124963(.A (n_14550), .B (n_3235), .Y (n_10240));
NAND2X1 g124965(.A (n_14550), .B (n_3333), .Y (n_10238));
AND2X1 g124968(.A (n_14550), .B (n_3716), .Y (n_10236));
NAND2X1 g124970(.A (n_14550), .B (n_3402), .Y (n_10234));
NAND2X1 g124972(.A (n_14550), .B (n_4554), .Y (n_10232));
NAND2X1 g124974(.A (n_14550), .B (n_4231), .Y (n_10230));
AND2X1 g124976(.A (n_14550), .B (n_4011), .Y (n_10228));
NAND2X1 g124997(.A (n_14550), .B (n_10223), .Y (n_10224));
AND2X1 g124999(.A (n_14550), .B (n_10221), .Y (n_10222));
NAND2X1 g125019(.A (n_14550), .B (n_10219), .Y (n_10220));
NAND2X1 g125026(.A (n_14550), .B (n_10217), .Y (n_10218));
AND2X1 g125038(.A (n_14550), .B (n_4534), .Y (n_10214));
NAND2X1 g125046(.A (n_14550), .B (n_10211), .Y (n_10212));
NAND2X1 g125050(.A (n_14550), .B (P1_reg1[12] ), .Y (n_10210));
NAND2X1 g125051(.A (n_14550), .B (P1_reg1[19] ), .Y (n_10208));
NAND2X1 g125052(.A (n_14550), .B (n_10205), .Y (n_10206));
OR2X1 g125056(.A (n_10203), .B (n_11138), .Y (n_10204));
NAND2X1 g125057(.A (n_14550), .B (n_10201), .Y (n_10202));
NAND2X1 g125059(.A (n_14550), .B (P1_reg1[0] ), .Y (n_10200));
NAND2X1 g125064(.A (n_14550), .B (n_10197), .Y (n_10198));
OR2X1 g125066(.A (n_34753), .B (n_10196), .Y (n_10925));
INVX1 g125070(.A (n_34312), .Y (n_30445));
AND2X1 g125079(.A (n_14550), .B (n_10191), .Y (n_10192));
NAND2X1 g125081(.A (n_14550), .B (n_10189), .Y (n_10190));
NAND2X1 g125082(.A (n_14550), .B (n_10187), .Y (n_10188));
NAND2X1 g125110(.A (n_14550), .B (n_10182), .Y (n_10183));
AND2X1 g125111(.A (n_14550), .B (n_10180), .Y (n_10181));
NAND2X1 g125113(.A (n_14550), .B (n_10178), .Y (n_10179));
NAND2X1 g125115(.A (n_14550), .B (P1_reg1[24] ), .Y (n_10177));
NAND2X1 g125116(.A (n_14550), .B (n_10175), .Y (n_10176));
AND2X1 g125122(.A (n_14550), .B (n_10173), .Y (n_10174));
NAND2X1 g125127(.A (n_14550), .B (n_10171), .Y (n_10172));
NAND2X1 g125128(.A (n_14550), .B (n_10169), .Y (n_10170));
NAND2X1 g125129(.A (n_14550), .B (n_10167), .Y (n_10168));
NAND2X1 g125130(.A (n_14550), .B (n_10165), .Y (n_10166));
NAND2X1 g125132(.A (n_14550), .B (P1_reg_172), .Y (n_10164));
NAND2X1 g125133(.A (n_14550), .B (P1_reg_173), .Y (n_10163));
NAND2X1 g125136(.A (n_14550), .B (n_10161), .Y (n_10162));
NAND2X1 g125137(.A (n_14550), .B (P1_reg_174), .Y (n_10160));
NAND2X1 g125139(.A (n_14550), .B (n_10158), .Y (n_10159));
NAND2X1 g125140(.A (n_14550), .B (n_10156), .Y (n_10157));
AND2X1 g125141(.A (n_14550), .B (n_10154), .Y (n_10155));
NAND2X1 g125144(.A (n_14550), .B (n_10152), .Y (n_10153));
NAND2X1 g125146(.A (n_14550), .B (n_10150), .Y (n_10151));
AND2X1 g125153(.A (n_14550), .B (n_10148), .Y (n_10149));
NAND2X1 g125155(.A (n_14550), .B (n_3958), .Y (n_10147));
NAND2X1 g125163(.A (n_14550), .B (n_10144), .Y (n_10145));
AND2X1 g125165(.A (n_14550), .B (P1_reg1[16] ), .Y (n_10143));
NAND2X1 g125170(.A (n_14550), .B (n_10140), .Y (n_10141));
NAND2X1 g125173(.A (n_14550), .B (n_10138), .Y (n_10139));
NAND2X1 g125175(.A (n_14550), .B (n_10136), .Y (n_10137));
NAND2X1 g125181(.A (n_14550), .B (n_10134), .Y (n_10135));
NAND2X1 g125183(.A (n_14550), .B (P1_reg1[14] ), .Y (n_10133));
AND2X1 g125185(.A (n_14550), .B (n_4920), .Y (n_10131));
NAND2X1 g125187(.A (n_14550), .B (n_10128), .Y (n_10129));
NAND2X1 g125189(.A (n_14550), .B (n_4477), .Y (n_10127));
AND2X1 g125192(.A (n_14550), .B (P1_reg1[1] ), .Y (n_10126));
NAND2X1 g125201(.A (n_9625), .B (n_27045), .Y (n_10124));
OR2X1 g125203(.A (n_10203), .B (n_14351), .Y (n_11177));
AOI21X1 g125212(.A0 (n_9162), .A1 (n_8687), .B0 (n_9507), .Y(n_10123));
AOI22X1 g125218(.A0 (n_11138), .A1 (n_13511), .B0 (n_7734), .B1(n_7988), .Y (n_10122));
OAI21X1 g125254(.A0 (n_10119), .A1 (n_8309), .B0 (n_9031), .Y(n_10120));
OAI21X1 g125255(.A0 (n_10116), .A1 (n_8309), .B0 (n_9024), .Y(n_10117));
OAI21X1 g125256(.A0 (n_10114), .A1 (n_8309), .B0 (n_9023), .Y(n_10115));
OAI21X1 g125257(.A0 (n_10112), .A1 (n_8309), .B0 (n_9026), .Y(n_10113));
OAI21X1 g125258(.A0 (n_10110), .A1 (n_8309), .B0 (n_9025), .Y(n_10111));
AOI22X1 g125259(.A0 (n_11138), .A1 (n_13515), .B0 (n_7755), .B1(n_7988), .Y (n_10108));
OAI21X1 g125260(.A0 (n_4154), .A1 (n_8309), .B0 (n_9028), .Y(n_10105));
OAI21X1 g125261(.A0 (n_10103), .A1 (n_8309), .B0 (n_9027), .Y(n_10104));
AOI22X1 g125292(.A0 (n_11138), .A1 (P3_reg2[10] ), .B0 (n_10100),.B1 (n_7988), .Y (n_10102));
AOI22X1 g125298(.A0 (n_11138), .A1 (n_13366), .B0 (n_10097), .B1(n_7988), .Y (n_10098));
AOI22X1 g125299(.A0 (n_11138), .A1 (n_13507), .B0 (n_8055), .B1(n_7988), .Y (n_10096));
AOI22X1 g125305(.A0 (n_11138), .A1 (n_13361), .B0 (n_13711), .B1(n_7988), .Y (n_10095));
AOI22X1 g125307(.A0 (n_11160), .A1 (n_7587), .B0 (n_18289), .B1(addr_446), .Y (n_10094));
AOI22X1 g125314(.A0 (n_11138), .A1 (n_13338), .B0 (n_13327), .B1(n_7988), .Y (n_10093));
AOI22X1 g125327(.A0 (n_11151), .A1 (n_25111), .B0 (n_18289), .B1(n_233), .Y (n_10092));
INVX1 g125333(.A (n_9635), .Y (n_10090));
INVX1 g125344(.A (n_9541), .Y (n_10089));
AOI22X1 g125351(.A0 (n_18289), .A1 (P2_reg2[18] ), .B0 (n_8164), .B1(n_10848), .Y (n_10088));
INVX1 g125352(.A (n_9538), .Y (n_10084));
AOI22X1 g125356(.A0 (n_18289), .A1 (n_10082), .B0 (n_10081), .B1(n_18909), .Y (n_10083));
AOI22X1 g125358(.A0 (n_11138), .A1 (n_13332), .B0 (n_19108), .B1(P3_reg3[2] ), .Y (n_10080));
AOI22X1 g125360(.A0 (n_18289), .A1 (n_3565), .B0 (n_1183), .B1(n_18909), .Y (n_10079));
AOI22X1 g125362(.A0 (n_11138), .A1 (n_13337), .B0 (n_19108), .B1(n_13675), .Y (n_10076));
AOI22X1 g125363(.A0 (n_11138), .A1 (n_565), .B0 (n_7988), .B1(P3_reg3[0] ), .Y (n_10074));
AOI22X1 g125364(.A0 (n_11151), .A1 (n_10063), .B0 (n_22821), .B1(n_233), .Y (n_10071));
AOI22X1 g125367(.A0 (n_11157), .A1 (n_7587), .B0 (n_18289), .B1(addr_2), .Y (n_10069));
NAND4X1 g125368(.A (n_9441), .B (n_10067), .C (n_8942), .D (n_8305),.Y (n_10932));
CLKBUFX3 g128379(.A (n_17380), .Y (n_18496));
AOI22X1 g125380(.A0 (n_11153), .A1 (n_25111), .B0 (n_18289), .B1(n_130), .Y (n_10066));
AOI22X1 g125381(.A0 (n_11157), .A1 (n_10063), .B0 (n_8313), .B1(addr_2), .Y (n_10064));
AOI22X1 g125382(.A0 (n_11155), .A1 (n_10063), .B0 (n_22821), .B1(n_10057), .Y (n_10061));
AOI22X1 g125387(.A0 (n_11155), .A1 (n_7587), .B0 (n_18289), .B1(n_10057), .Y (n_10059));
AOI22X1 g125388(.A0 (n_11153), .A1 (n_29090), .B0 (n_8313), .B1(n_130), .Y (n_10056));
AOI22X1 g125394(.A0 (n_11138), .A1 (P3_reg2[6] ), .B0 (n_13735), .B1(n_7988), .Y (n_10053));
AOI22X1 g125395(.A0 (n_11160), .A1 (n_29090), .B0 (n_8313), .B1(addr_446), .Y (n_10052));
NAND2X1 g124798(.A (n_30230), .B (n_10049), .Y (n_10050));
NAND2X1 g125439(.A (n_18289), .B (n_10047), .Y (n_10048));
NAND2X1 g125444(.A (n_18289), .B (P2_reg2[8] ), .Y (n_10046));
NAND2X1 g125452(.A (n_18289), .B (n_10043), .Y (n_10044));
NAND2X1 g125467(.A (n_18289), .B (n_10041), .Y (n_10042));
NAND2X1 g125486(.A (n_7724), .B (n_8946), .Y (n_10040));
NAND2X1 g125492(.A (n_13167), .B (n_8946), .Y (n_10038));
NAND2X1 g125493(.A (n_2138), .B (n_8946), .Y (n_10037));
NAND2X1 g125494(.A (n_2601), .B (n_8946), .Y (n_10036));
NOR2X1 g125506(.A (n_9429), .B (n_10034), .Y (n_10035));
NAND2X1 g125507(.A (n_18289), .B (n_10032), .Y (n_10033));
NAND2X1 g125517(.A (n_2911), .B (n_8946), .Y (n_10031));
NOR2X1 g125548(.A (n_8325), .B (P2_reg3[3] ), .Y (n_10030));
INVX1 g128357(.A (n_17906), .Y (n_10540));
INVX1 g125743(.A (n_20864), .Y (n_20399));
INVX1 g125755(.A (n_33803), .Y (n_21201));
INVX1 g125762(.A (n_21365), .Y (n_22123));
INVX1 g125772(.A (n_33803), .Y (n_21374));
NOR2X1 g125786(.A (n_8946), .B (n_25942), .Y (n_10629));
AOI22X1 g129475(.A0 (n_3583), .A1 (n_10676), .B0 (n_9676), .B1(addr_489), .Y (n_10014));
INVX1 g125815(.A (n_33513), .Y (n_14159));
CLKBUFX1 g125852(.A (n_28785), .Y (n_26528));
INVX2 g128339(.A (n_10006), .Y (n_10303));
CLKBUFX1 g125900(.A (n_27462), .Y (n_29430));
INVX1 g125908(.A (n_8677), .Y (n_26132));
INVX1 g125909(.A (n_8677), .Y (n_28347));
INVX1 g125913(.A (n_10003), .Y (n_26255));
INVX1 g125916(.A (n_10002), .Y (n_27632));
INVX1 g125922(.A (n_8692), .Y (n_29427));
INVX1 g125925(.A (n_8692), .Y (n_29341));
INVX1 g125926(.A (n_8692), .Y (n_29695));
NAND2X1 g125934(.A (n_7862), .B (n_14956), .Y (n_9998));
NAND2X1 g125947(.A (n_27522), .B (n_27042), .Y (n_9997));
INVX1 g126063(.A (n_9994), .Y (n_13232));
INVX1 g126064(.A (n_9994), .Y (n_9995));
INVX4 g126219(.A (n_34719), .Y (n_28926));
INVX1 g126340(.A (n_27045), .Y (n_26535));
INVX1 g126481(.A (n_33784), .Y (n_9983));
CLKBUFX1 g126483(.A (n_33784), .Y (n_29455));
INVX1 g126539(.A (n_14956), .Y (n_29968));
INVX1 g126554(.A (n_9978), .Y (n_14916));
INVX1 g126557(.A (n_9978), .Y (n_26801));
INVX1 g126559(.A (n_9978), .Y (n_25368));
INVX1 g126570(.A (n_14743), .Y (n_9971));
INVX1 g126592(.A (n_25540), .Y (n_20887));
INVX1 g126609(.A (n_25540), .Y (n_30505));
AND2X1 g126830(.A (n_8868), .B (n_10465), .Y (n_9964));
AND2X1 g126835(.A (n_8867), .B (n_6389), .Y (n_9963));
NAND2X1 g126848(.A (n_16084), .B (n_9962), .Y (n_10474));
NAND2X1 g126863(.A (n_8809), .B (n_9909), .Y (n_9961));
INVX1 g126887(.A (n_9960), .Y (n_10472));
NAND2X1 g126891(.A (n_35663), .B (n_33963), .Y (n_9959));
NAND2X1 g126897(.A (n_9302), .B (n_9303), .Y (n_9958));
NAND2X2 g126900(.A (n_9956), .B (n_9277), .Y (n_10794));
NOR2X1 g126905(.A (n_9279), .B (n_9956), .Y (n_32885));
INVX1 g126910(.A (n_34651), .Y (n_10467));
NAND2X1 g126947(.A (n_8818), .B (n_9909), .Y (n_9955));
NAND2X1 g126979(.A (n_9953), .B (n_12289), .Y (n_11295));
INVX1 g127042(.A (n_8718), .Y (n_30399));
INVX1 g127044(.A (n_8718), .Y (n_26611));
INVX1 g127076(.A (n_29505), .Y (n_25376));
NOR2X1 g127186(.A (n_8858), .B (n_9946), .Y (n_9947));
NOR2X1 g127189(.A (n_8709), .B (n_10414), .Y (n_9945));
NOR2X1 g127195(.A (n_8837), .B (n_10414), .Y (n_9944));
NAND3X1 g127196(.A (n_9909), .B (n_4231), .C (n_8245), .Y (n_9943));
NOR2X1 g127199(.A (n_8791), .B (n_9946), .Y (n_9942));
NOR2X1 g127202(.A (n_8877), .B (n_10399), .Y (n_9940));
NOR2X1 g127207(.A (n_8853), .B (n_9937), .Y (n_9939));
NOR2X1 g127209(.A (n_8815), .B (n_9937), .Y (n_9938));
NOR2X1 g127210(.A (n_8847), .B (n_9934), .Y (n_9936));
NOR2X1 g127212(.A (n_8846), .B (n_9934), .Y (n_9935));
NOR2X1 g127213(.A (n_8843), .B (n_9937), .Y (n_9933));
NOR2X1 g127215(.A (n_8841), .B (n_9928), .Y (n_9932));
NOR2X1 g127218(.A (n_8840), .B (n_9934), .Y (n_9931));
NOR2X1 g127225(.A (n_8826), .B (n_9934), .Y (n_9930));
NOR2X1 g127227(.A (n_8794), .B (n_9928), .Y (n_9929));
NOR2X1 g127229(.A (n_8713), .B (n_10414), .Y (n_9927));
NOR2X1 g127230(.A (n_8833), .B (n_10414), .Y (n_9925));
NOR2X1 g127234(.A (n_8743), .B (n_9946), .Y (n_9924));
NOR2X1 g127235(.A (n_8878), .B (n_12755), .Y (n_9923));
NOR2X1 g127240(.A (n_8796), .B (n_9928), .Y (n_9922));
NOR2X1 g127241(.A (n_8886), .B (n_12755), .Y (n_9921));
NOR2X1 g127242(.A (n_8779), .B (n_9946), .Y (n_9920));
NAND3X1 g127244(.A (n_9909), .B (P1_reg1[1] ), .C (n_8245), .Y(n_9919));
NOR2X1 g127246(.A (n_8827), .B (n_10414), .Y (n_9917));
NAND3X1 g127247(.A (n_9909), .B (P1_reg2[9] ), .C (n_8245), .Y(n_9916));
NOR2X1 g127258(.A (n_8824), .B (n_9928), .Y (n_9912));
NOR2X1 g127265(.A (n_8817), .B (n_9934), .Y (n_9911));
NAND3X1 g127275(.A (n_9909), .B (n_10167), .C (n_8245), .Y (n_9910));
NAND3X1 g129319(.A (n_8734), .B (n_8433), .C (n_8431), .Y (n_10960));
NOR2X1 g127291(.A (n_8880), .B (n_7250), .Y (n_9908));
NOR2X1 g127297(.A (n_8835), .B (n_9934), .Y (n_9907));
NOR2X1 g127299(.A (n_8874), .B (n_12755), .Y (n_9906));
NOR2X1 g127300(.A (n_8750), .B (n_12917), .Y (n_9905));
NOR2X1 g127309(.A (n_8814), .B (n_9937), .Y (n_9903));
NOR2X1 g127313(.A (n_8869), .B (n_12755), .Y (n_9902));
NOR2X1 g127321(.A (n_8825), .B (n_9946), .Y (n_9900));
NOR2X1 g127322(.A (n_8875), .B (n_10342), .Y (n_9899));
NOR2X1 g127330(.A (n_8883), .B (n_12917), .Y (n_9898));
NOR2X1 g127331(.A (n_8873), .B (n_12755), .Y (n_9897));
NOR2X1 g127333(.A (n_8870), .B (n_12755), .Y (n_9896));
NOR2X1 g127339(.A (n_8785), .B (n_9946), .Y (n_9895));
NOR2X1 g127342(.A (n_8876), .B (n_12755), .Y (n_9894));
NOR2X1 g127349(.A (n_8872), .B (n_12755), .Y (n_9893));
NOR2X1 g127357(.A (n_8881), .B (n_12755), .Y (n_9891));
NOR2X1 g127359(.A (n_8885), .B (n_12755), .Y (n_9890));
NOR2X1 g127361(.A (n_8871), .B (n_12755), .Y (n_9889));
NOR2X1 g127372(.A (n_8816), .B (n_9937), .Y (n_9888));
NAND3X1 g127377(.A (n_9909), .B (n_10217), .C (n_8245), .Y (n_9887));
NAND2X1 g127409(.A (n_13727), .B (n_8884), .Y (n_9882));
NAND2X1 g127413(.A (n_8742), .B (n_8245), .Y (n_12662));
NAND2X1 g127416(.A (n_13515), .B (n_9859), .Y (n_9881));
NAND2X1 g127425(.A (n_13368), .B (n_9373), .Y (n_9880));
NAND2X1 g127429(.A (n_13205), .B (n_9859), .Y (n_9879));
NAND2X1 g127441(.A (n_13344), .B (n_9859), .Y (n_9878));
NAND2X1 g127450(.A (n_13507), .B (n_8884), .Y (n_9876));
NAND2X1 g127454(.A (n_565), .B (n_8884), .Y (n_9875));
NAND2X1 g127466(.A (n_13342), .B (n_8884), .Y (n_9873));
NAND2X1 g127468(.A (n_9373), .B (n_27232), .Y (n_9871));
NAND2X1 g127470(.A (n_14317), .B (n_8884), .Y (n_9869));
NAND2X1 g127471(.A (n_13212), .B (n_9859), .Y (n_9868));
NAND2X1 g127472(.A (n_13336), .B (n_9859), .Y (n_9867));
NAND2X1 g127474(.A (n_13511), .B (n_9373), .Y (n_9866));
NAND2X1 g127476(.A (n_13200), .B (n_9859), .Y (n_9864));
NAND2X1 g127479(.A (n_13330), .B (n_9859), .Y (n_9863));
NAND2X1 g127480(.A (n_2718), .B (n_9373), .Y (n_9862));
NAND2X1 g127481(.A (n_13206), .B (n_9859), .Y (n_9861));
NAND2X1 g127492(.A (n_13216), .B (n_9859), .Y (n_9860));
NAND2X1 g127500(.A (n_13352), .B (n_9859), .Y (n_9858));
NAND2X1 g127505(.A (n_13329), .B (n_8884), .Y (n_9857));
NAND2X1 g127506(.A (n_13211), .B (n_9859), .Y (n_9856));
NAND2X1 g127516(.A (n_13335), .B (n_9859), .Y (n_9855));
NAND2X1 g127517(.A (n_13334), .B (n_9859), .Y (n_9854));
NAND2X1 g127520(.A (n_13215), .B (n_8884), .Y (n_9853));
NAND2X1 g127522(.A (n_13213), .B (n_8884), .Y (n_9852));
NAND2X1 g127524(.A (P3_reg1[16] ), .B (n_8884), .Y (n_9851));
NAND2X1 g127526(.A (n_13681), .B (n_8884), .Y (n_9850));
NAND2X1 g127529(.A (n_13202), .B (n_9373), .Y (n_9849));
NAND2X1 g127530(.A (n_13208), .B (n_9859), .Y (n_9848));
NAND2X1 g127531(.A (n_13343), .B (n_9859), .Y (n_9847));
NAND2X1 g127533(.A (n_13207), .B (n_9373), .Y (n_9846));
NAND2X1 g127538(.A (n_13199), .B (n_9373), .Y (n_9845));
NAND2X1 g127542(.A (P3_reg1[18] ), .B (n_8884), .Y (n_9844));
NAND2X1 g127543(.A (P3_reg1[4] ), .B (n_9373), .Y (n_9843));
INVX1 g128226(.A (n_16903), .Y (n_17351));
NAND2X1 g127547(.A (n_13209), .B (n_9373), .Y (n_9842));
NAND2X1 g127548(.A (n_13204), .B (n_9373), .Y (n_9841));
NAND2X1 g127561(.A (P3_reg2[15] ), .B (n_9859), .Y (n_9840));
OR2X1 g127565(.A (n_9038), .B (n_8484), .Y (n_9839));
NAND2X1 g127566(.A (n_13732), .B (n_8884), .Y (n_9838));
NAND3X1 g127570(.A (n_8740), .B (n_7551), .C (n_7218), .Y (n_11573));
NOR2X1 g127575(.A (P2_d_402), .B (n_9310), .Y (n_9837));
NOR2X1 g127576(.A (P2_d_386), .B (n_9310), .Y (n_9836));
NOR2X1 g127577(.A (P2_d_398), .B (n_9310), .Y (n_9835));
NOR2X1 g127578(.A (P2_d_387), .B (n_9813), .Y (n_9834));
NOR2X1 g127579(.A (P2_d_393), .B (n_9813), .Y (n_9833));
NOR2X1 g127580(.A (P2_d_408), .B (n_9813), .Y (n_9832));
NOR2X1 g127581(.A (P2_d_407), .B (n_9813), .Y (n_9830));
NOR2X1 g127582(.A (P2_d), .B (n_8534), .Y (n_9828));
NOR2X1 g127583(.A (P2_d_392), .B (n_9813), .Y (n_9827));
NOR2X1 g127584(.A (P2_d_397), .B (n_9310), .Y (n_9826));
NOR2X1 g127585(.A (P2_d_405), .B (n_9310), .Y (n_9825));
NOR2X1 g127586(.A (P2_d_385), .B (n_9813), .Y (n_9823));
NOR2X1 g127587(.A (P2_d_380), .B (n_9310), .Y (n_9822));
NOR2X1 g127589(.A (P2_d_391), .B (n_9310), .Y (n_9820));
NOR2X1 g127591(.A (P2_d_399), .B (n_9310), .Y (n_9819));
NOR2X1 g127592(.A (P2_d_406), .B (n_9310), .Y (n_9818));
NOR2X1 g127593(.A (P2_d_378), .B (n_9310), .Y (n_9816));
NOR2X1 g127595(.A (P2_d_383), .B (n_9310), .Y (n_9815));
NOR2X1 g127596(.A (n_2979), .B (n_9813), .Y (n_9814));
NOR2X1 g127597(.A (P2_d_389), .B (n_9310), .Y (n_9812));
NOR2X1 g127602(.A (P2_d_396), .B (n_9813), .Y (n_9811));
NOR2X1 g127603(.A (P2_d_395), .B (n_9813), .Y (n_9810));
NOR2X1 g127605(.A (P2_d_401), .B (n_9310), .Y (n_9809));
NOR2X1 g127606(.A (P2_d_384), .B (n_9813), .Y (n_9807));
NOR2X1 g127607(.A (P2_d_404), .B (n_8534), .Y (n_9806));
NOR2X1 g127608(.A (P2_d_403), .B (n_8400), .Y (n_9804));
NOR2X1 g127609(.A (P2_d_379), .B (n_9310), .Y (n_9803));
NOR2X1 g127611(.A (P2_d_400), .B (n_8534), .Y (n_9802));
NOR2X1 g127613(.A (P2_d_388), .B (n_8534), .Y (n_9801));
NOR2X1 g127614(.A (P2_d_381), .B (n_9310), .Y (n_9800));
CLKBUFX1 g127619(.A (n_10758), .Y (n_17467));
INVX1 g127636(.A (n_16011), .Y (n_10718));
INVX1 g127643(.A (n_9798), .Y (n_17472));
NOR2X1 g127649(.A (P3_d_392), .B (n_8484), .Y (n_9797));
INVX4 g127661(.A (n_17000), .Y (n_17916));
NAND2X1 g127665(.A (n_9794), .B (n_8393), .Y (n_9795));
INVX2 g127673(.A (n_9793), .Y (n_10270));
INVX1 g127678(.A (n_9792), .Y (n_10335));
NOR2X1 g127692(.A (P3_d_388), .B (n_8484), .Y (n_9791));
NOR2X1 g127694(.A (P3_d_394), .B (n_8484), .Y (n_9789));
NAND2X1 g127708(.A (n_8178), .B (n_8762), .Y (n_10272));
INVX1 g127724(.A (n_10717), .Y (n_10273));
INVX1 g127756(.A (n_9788), .Y (n_10330));
INVX2 g127774(.A (n_9785), .Y (n_10275));
NAND2X1 g127788(.A (P2_reg1[19] ), .B (n_8393), .Y (n_9783));
INVX1 g127789(.A (n_9780), .Y (n_10760));
INVX2 g127823(.A (n_16012), .Y (n_16446));
INVX1 g127830(.A (n_11089), .Y (n_10329));
NAND2X1 g127836(.A (P2_reg2[15] ), .B (n_8393), .Y (n_9778));
INVX1 g127839(.A (n_8830), .Y (n_17955));
INVX1 g127853(.A (n_10754), .Y (n_9776));
INVX1 g128190(.A (n_16646), .Y (n_9775));
NAND2X1 g127860(.A (n_9773), .B (n_8393), .Y (n_9774));
NAND2X1 g127862(.A (n_10043), .B (n_8393), .Y (n_9772));
NOR2X1 g127863(.A (n_2096), .B (n_8484), .Y (n_9771));
NAND2X1 g127870(.A (n_14096), .B (n_8393), .Y (n_9770));
NAND2X1 g127872(.A (n_13893), .B (n_8393), .Y (n_9769));
NAND2X1 g127922(.A (P2_reg2[8] ), .B (n_8393), .Y (n_9767));
INVX1 g127931(.A (n_9292), .Y (n_10326));
NAND2X1 g127938(.A (n_13388), .B (n_8884), .Y (n_9766));
NAND2X1 g127947(.A (n_3887), .B (n_8884), .Y (n_9765));
NOR2X1 g127950(.A (P3_d_400), .B (n_8484), .Y (n_9763));
NOR2X1 g127989(.A (P3_reg3[3] ), .B (n_8484), .Y (n_9760));
NOR2X1 g127991(.A (P3_d_406), .B (n_8484), .Y (n_9758));
INVX1 g128018(.A (n_8436), .Y (n_10320));
INVX1 g128059(.A (n_16186), .Y (n_16419));
INVX1 g128063(.A (n_17471), .Y (n_10316));
INVX1 g128073(.A (n_9755), .Y (n_10315));
INVX1 g128082(.A (n_9754), .Y (n_10314));
NAND2X1 g128094(.A (P2_reg1[22] ), .B (n_8393), .Y (n_9752));
INVX1 g128107(.A (n_8803), .Y (n_10287));
INVX1 g128115(.A (n_9749), .Y (n_10312));
INVX2 g128147(.A (n_9238), .Y (n_16182));
NAND2X1 g128150(.A (n_3565), .B (n_8393), .Y (n_9748));
INVX1 g128166(.A (n_15908), .Y (n_10309));
INVX2 g128173(.A (n_9746), .Y (n_9745));
INVX1 g128181(.A (n_9744), .Y (n_17162));
INVX1 g128189(.A (n_16646), .Y (n_10325));
INVX1 g128197(.A (n_16188), .Y (n_11246));
CLKBUFX1 g128205(.A (n_9742), .Y (n_10767));
INVX2 g128280(.A (n_10706), .Y (n_10451));
NAND4X1 g128308(.A (n_7984), .B (n_8440), .C (n_7928), .D (n_8158),.Y (n_16167));
NOR2X1 g128316(.A (n_8757), .B (n_8457), .Y (n_16008));
INVX1 g128340(.A (n_10006), .Y (n_9729));
INVX2 g128369(.A (n_9253), .Y (n_15909));
NOR2X1 g128397(.A (P3_d_381), .B (n_8484), .Y (n_9726));
INVX1 g128413(.A (n_10485), .Y (n_10267));
NOR2X1 g128495(.A (P3_d_407), .B (n_8484), .Y (n_9719));
NOR2X1 g128496(.A (P3_d_384), .B (n_8484), .Y (n_9718));
CLKBUFX1 g128497(.A (n_8784), .Y (n_15810));
CLKBUFX1 g128518(.A (n_16064), .Y (n_17262));
INVX1 g128519(.A (n_16064), .Y (n_9714));
NOR2X1 g128524(.A (P3_d_404), .B (n_8484), .Y (n_9713));
NOR2X1 g128527(.A (P3_d_390), .B (n_8484), .Y (n_9711));
NOR2X1 g128530(.A (P3_d_383), .B (n_8484), .Y (n_9710));
NOR2X1 g128531(.A (P3_d_401), .B (n_8484), .Y (n_9709));
NAND2X1 g128533(.A (P2_reg1[18] ), .B (n_8393), .Y (n_9708));
CLKBUFX3 g128537(.A (n_16984), .Y (n_10755));
INVX2 g128542(.A (n_16103), .Y (n_9706));
NOR2X1 g128559(.A (P3_d_389), .B (n_8484), .Y (n_9704));
NOR2X1 g128560(.A (P3_d_402), .B (n_8484), .Y (n_9703));
NOR2X1 g128590(.A (P3_d_395), .B (n_8484), .Y (n_9699));
NOR2X1 g128592(.A (P3_d_403), .B (n_8484), .Y (n_9698));
NAND3X1 g128928(.A (n_8154), .B (n_6956), .C (n_8408), .Y (n_10973));
AOI21X1 g128978(.A0 (n_9097), .A1 (n_9692), .B0 (n_8754), .Y(n_32287));
AOI21X1 g128979(.A0 (n_9178), .A1 (n_8445), .B0 (n_8752), .Y(n_9695));
AOI21X1 g129070(.A0 (n_9092), .A1 (n_9692), .B0 (n_8755), .Y(n_9693));
AOI21X1 g129073(.A0 (P2_reg_108), .A1 (n_7983), .B0 (n_8925), .Y(n_9691));
NOR2X1 g129074(.A (n_8633), .B (n_8753), .Y (n_32286));
NAND2X1 g129096(.A (n_8749), .B (n_8446), .Y (n_9689));
NAND2X1 g129111(.A (n_8747), .B (n_7828), .Y (n_10708));
NAND3X1 g128927(.A (n_8151), .B (n_6954), .C (n_8410), .Y (n_10943));
INVX2 g128051(.A (n_9688), .Y (n_10317));
NAND3X1 g129261(.A (n_8735), .B (n_7900), .C (n_7898), .Y (n_10986));
AOI22X1 g129498(.A0 (n_10740), .A1 (n_10676), .B0 (n_9676), .B1(addr_487), .Y (n_9687));
INVX1 g128039(.A (n_9684), .Y (n_10319));
NAND3X1 g129402(.A (n_8738), .B (n_8049), .C (n_8047), .Y (n_10969));
INVX2 g129430(.A (n_9683), .Y (n_16253));
INVX1 g129431(.A (n_9683), .Y (n_15959));
AOI22X1 g129448(.A0 (n_3429), .A1 (n_9677), .B0 (n_9676), .B1(addr_488), .Y (n_9682));
AOI22X1 g129464(.A0 (n_4288), .A1 (n_9677), .B0 (n_9676), .B1(n_9675), .Y (n_9679));
AOI22X1 g129465(.A0 (n_3854), .A1 (n_10676), .B0 (n_9676), .B1(addr_491), .Y (n_9674));
AOI22X1 g129466(.A0 (n_4320), .A1 (n_10676), .B0 (n_9676), .B1(n_9672), .Y (n_9673));
AOI22X1 g129467(.A0 (n_10656), .A1 (n_9668), .B0 (n_9676), .B1(n_9670), .Y (n_9671));
AOI22X1 g129468(.A0 (n_4735), .A1 (n_9668), .B0 (n_9676), .B1(n_9667), .Y (n_9669));
AOI22X1 g129469(.A0 (n_4133), .A1 (n_9668), .B0 (n_9676), .B1(addr_490), .Y (n_9666));
AOI22X1 g129470(.A0 (n_33901), .A1 (n_9668), .B0 (n_9676), .B1(n_9663), .Y (n_9665));
AOI22X1 g129471(.A0 (n_4844), .A1 (n_9677), .B0 (n_9676), .B1(n_1170), .Y (n_9662));
AOI22X1 g129473(.A0 (n_32386), .A1 (n_10676), .B0 (n_9676), .B1(n_9658), .Y (n_9659));
AOI22X1 g129474(.A0 (n_4040), .A1 (n_10676), .B0 (n_9676), .B1(n_9655), .Y (n_9657));
AOI22X1 g129476(.A0 (n_32445), .A1 (n_10676), .B0 (n_9676), .B1(n_9653), .Y (n_9654));
INVX1 g127997(.A (n_9652), .Y (n_10322));
NAND2X1 g129804(.A (n_6058), .B (n_9676), .Y (n_9651));
NAND2X1 g129805(.A (n_6183), .B (n_9676), .Y (n_9650));
NAND2X1 g129807(.A (n_5561), .B (n_9676), .Y (n_9648));
NAND2X1 g129808(.A (n_6037), .B (n_9676), .Y (n_9647));
NAND2X1 g129809(.A (n_6024), .B (n_9676), .Y (n_9646));
NAND2X1 g129811(.A (n_5613), .B (n_9676), .Y (n_9645));
NAND2X1 g129812(.A (n_5531), .B (n_9676), .Y (n_9644));
NAND2X1 g129819(.A (n_5999), .B (n_9676), .Y (n_9643));
NAND2X1 g129822(.A (n_5003), .B (n_9676), .Y (n_9642));
NAND2X1 g129840(.A (n_4887), .B (n_9676), .Y (n_9641));
NOR2X1 g127942(.A (n_8759), .B (n_8758), .Y (n_16251));
INVX1 g126090(.A (n_9473), .Y (n_10504));
INVX2 g128331(.A (n_9730), .Y (n_9640));
NOR2X1 g127350(.A (n_8882), .B (n_12755), .Y (n_9639));
NAND2X1 g126062(.A (n_9211), .B (n_9637), .Y (n_9638));
CLKBUFX1 g125905(.A (n_27462), .Y (n_30291));
INVX2 g125874(.A (n_34753), .Y (n_10276));
CLKBUFX1 g125823(.A (n_33494), .Y (n_26662));
INVX1 g125781(.A (n_33803), .Y (n_10525));
AOI22X1 g125334(.A0 (n_18289), .A1 (P2_reg2[2] ), .B0 (n_10848), .B1(n_9634), .Y (n_9635));
INVX4 g125757(.A (n_33803), .Y (n_21365));
INVX1 g125727(.A (n_20864), .Y (n_10020));
INVX1 g125720(.A (n_20864), .Y (n_10021));
INVX1 g128351(.A (n_9632), .Y (n_18584));
AOI22X1 g129472(.A0 (n_3862), .A1 (n_9677), .B0 (n_9676), .B1(addr_492), .Y (n_9631));
INVX1 g127731(.A (n_16331), .Y (n_10331));
CLKBUFX1 g128599(.A (n_16593), .Y (n_10768));
INVX1 g127716(.A (n_9628), .Y (n_10333));
INVX1 g128574(.A (n_9701), .Y (n_10756));
INVX1 g128556(.A (n_9627), .Y (n_16968));
NAND2X1 g124939(.A (n_34752), .B (n_33340), .Y (n_14534));
INVX1 g128546(.A (n_16103), .Y (n_10757));
INVX1 g128538(.A (n_16984), .Y (n_9623));
NAND2X1 g125551(.A (n_10032), .B (n_18909), .Y (n_9622));
NOR2X1 g125533(.A (n_8936), .B (n_8058), .Y (n_9621));
NOR2X1 g127610(.A (P2_d_382), .B (n_9813), .Y (n_9618));
CLKBUFX1 g126492(.A (n_33784), .Y (n_29199));
NOR2X1 g127604(.A (P2_d_390), .B (n_9310), .Y (n_9617));
CLKBUFX1 g126487(.A (n_33784), .Y (n_25980));
BUFX3 g126480(.A (n_33784), .Y (n_28013));
INVX2 g128478(.A (n_9722), .Y (n_11555));
INVX1 g127074(.A (n_29505), .Y (n_9616));
NAND3X1 g127004(.A (n_8703), .B (n_7661), .C (n_8387), .Y (n_11079));
NAND2X1 g124801(.A (n_9613), .B (n_11360), .Y (n_9615));
NAND2X1 g124806(.A (n_9613), .B (n_11357), .Y (n_9614));
NAND2X1 g124842(.A (n_9613), .B (n_11596), .Y (n_9612));
NAND2X1 g124926(.A (n_32479), .B (P3_d_377), .Y (n_9610));
NAND2X1 g124934(.A (n_32401), .B (n_7692), .Y (n_9609));
NAND2X1 g124959(.A (n_9603), .B (P2_reg_104), .Y (n_9608));
NAND2X1 g124961(.A (n_9603), .B (P2_reg_106), .Y (n_9607));
NAND2X1 g124964(.A (n_9603), .B (P2_reg_107), .Y (n_9606));
NAND2X1 g124967(.A (n_21365), .B (n_33505), .Y (n_11832));
NAND2X1 g124969(.A (n_9603), .B (P2_reg_95), .Y (n_9605));
NAND2X1 g124977(.A (n_9603), .B (n_9602), .Y (n_9604));
NAND2X1 g124984(.A (n_9603), .B (n_9599), .Y (n_9601));
NAND2X1 g124989(.A (n_9603), .B (n_9597), .Y (n_9598));
NAND2X1 g124991(.A (n_9603), .B (n_9595), .Y (n_9596));
NAND2X1 g124992(.A (n_9603), .B (n_9592), .Y (n_9594));
NAND2X1 g124995(.A (n_9603), .B (n_9590), .Y (n_9591));
NAND2X1 g124998(.A (n_9603), .B (P2_reg1[12] ), .Y (n_9589));
NAND2X1 g125000(.A (n_9603), .B (n_9586), .Y (n_9587));
NAND2X1 g125002(.A (n_9603), .B (P2_reg1[16] ), .Y (n_9585));
NAND2X1 g125017(.A (n_9603), .B (P2_reg1[20] ), .Y (n_9583));
NAND2X1 g125018(.A (n_9603), .B (P2_reg1[23] ), .Y (n_35112));
NOR2X1 g125027(.A (n_9557), .B (n_290), .Y (n_9581));
NAND2X1 g125032(.A (n_9603), .B (P2_reg1[3] ), .Y (n_9580));
NAND2X1 g129815(.A (n_5330), .B (n_9676), .Y (n_9578));
NAND2X1 g125037(.A (n_9603), .B (P2_reg1[6] ), .Y (n_9577));
NAND2X1 g125039(.A (n_9603), .B (n_4237), .Y (n_9575));
NAND2X1 g125040(.A (n_9603), .B (P2_reg1[8] ), .Y (n_9573));
NAND2X1 g125044(.A (n_9603), .B (P2_reg1[11] ), .Y (n_9571));
NOR2X1 g125047(.A (n_9557), .B (P3_reg_146), .Y (n_9569));
NOR2X1 g125055(.A (n_9557), .B (P3_reg_150), .Y (n_9567));
NAND2X1 g125058(.A (n_9603), .B (n_9565), .Y (n_9566));
NAND2X1 g125061(.A (n_8998), .B (n_8678), .Y (n_10975));
INVX1 g125073(.A (n_30050), .Y (n_30171));
INVX4 g125102(.A (n_26382), .Y (n_24925));
NAND2X1 g125123(.A (n_8677), .B (n_7997), .Y (n_10917));
NOR2X1 g125124(.A (n_9557), .B (P3_reg_151), .Y (n_9562));
NAND2X1 g125138(.A (n_14810), .B (n_13215), .Y (n_9561));
NAND2X1 g125145(.A (n_9498), .B (n_8692), .Y (n_11354));
NOR2X1 g125152(.A (n_9557), .B (P3_reg_148), .Y (n_9559));
NOR2X1 g125157(.A (n_9557), .B (n_7043), .Y (n_9558));
NOR2X1 g125162(.A (n_9557), .B (P3_reg_145), .Y (n_9556));
NOR2X1 g125164(.A (n_9557), .B (P3_reg_149), .Y (n_9555));
NOR2X1 g125169(.A (n_9557), .B (P3_reg_153), .Y (n_9554));
NOR2X1 g125171(.A (n_9557), .B (P3_reg_152), .Y (n_9553));
NAND2X1 g129806(.A (n_6360), .B (n_9676), .Y (n_9552));
NAND2X1 g125184(.A (n_14810), .B (n_2718), .Y (n_9551));
NAND2X1 g125188(.A (n_9603), .B (n_9549), .Y (n_9550));
AND2X1 g125193(.A (n_14810), .B (n_14513), .Y (n_9548));
NOR2X1 g125195(.A (n_9557), .B (P3_reg_147), .Y (n_9547));
OR2X1 g125204(.A (n_14351), .B (n_8954), .Y (n_9546));
NAND2X2 g128381(.A (n_32562), .B (n_32563), .Y (n_17380));
NAND2X1 g129803(.A (n_6118), .B (n_9676), .Y (n_9544));
NAND3X1 g129407(.A (n_8705), .B (n_8345), .C (n_8343), .Y (n_10953));
NAND2X1 g129801(.A (n_3766), .B (n_9676), .Y (n_9542));
AOI22X1 g125345(.A0 (n_18289), .A1 (n_4160), .B0 (n_2909), .B1(n_18909), .Y (n_9541));
AOI22X1 g125353(.A0 (n_18289), .A1 (P2_reg2[19] ), .B0 (n_3191), .B1(n_18909), .Y (n_9538));
NAND3X1 g129406(.A (n_8736), .B (n_8428), .C (n_8427), .Y (n_10951));
NAND2X1 g125429(.A (n_11138), .B (P3_reg2[15] ), .Y (n_9534));
NAND2X1 g125437(.A (n_18289), .B (P2_reg2[16] ), .Y (n_9532));
NAND2X1 g125443(.A (n_18289), .B (n_3709), .Y (n_9531));
NAND2X1 g125445(.A (n_18289), .B (P2_reg3[1] ), .Y (n_9530));
NAND2X1 g125446(.A (n_11138), .B (n_13342), .Y (n_9529));
NAND2X1 g125447(.A (n_11138), .B (P3_reg2[18] ), .Y (n_9528));
NAND2X1 g125449(.A (n_18289), .B (P2_reg2[9] ), .Y (n_9527));
NAND2X1 g125450(.A (n_11138), .B (n_13201), .Y (n_9525));
NAND2X1 g125461(.A (n_11138), .B (n_13358), .Y (n_9524));
NAND2X1 g125462(.A (n_11138), .B (n_13502), .Y (n_9523));
NOR2X1 g125466(.A (n_9520), .B (n_2096), .Y (n_9522));
NOR2X1 g125472(.A (n_9520), .B (n_3269), .Y (n_9521));
NOR2X1 g125485(.A (n_9520), .B (n_3573), .Y (n_9519));
NAND2X1 g125498(.A (n_1911), .B (n_10848), .Y (n_9517));
NAND2X1 g125502(.A (n_18289), .B (n_2909), .Y (n_9516));
NAND2X1 g125504(.A (n_18289), .B (n_8164), .Y (n_9515));
NAND2X1 g125505(.A (n_18289), .B (n_3191), .Y (n_9514));
AND2X1 g125518(.A (n_18289), .B (n_9512), .Y (n_9513));
NAND2X1 g125522(.A (n_8980), .B (n_9199), .Y (n_9511));
NOR2X1 g125537(.A (n_9520), .B (n_3297), .Y (n_9510));
NAND2X1 g125539(.A (n_2784), .B (n_10848), .Y (n_9509));
INVX1 g125544(.A (n_9507), .Y (n_9508));
NOR2X1 g125572(.A (n_9520), .B (P3_reg3[3] ), .Y (n_9506));
NAND2X1 g125574(.A (n_10041), .B (n_18909), .Y (n_9505));
NAND2X1 g125575(.A (n_8981), .B (n_8945), .Y (n_11612));
INVX4 g125594(.A (n_9625), .Y (n_28864));
INVX1 g125600(.A (n_9625), .Y (n_26162));
INVX2 g125610(.A (n_9626), .Y (n_29061));
INVX1 g125639(.A (n_9503), .Y (n_9502));
NAND2X1 g125661(.A (n_9983), .B (n_10067), .Y (n_26978));
NAND2X1 g125662(.A (n_9441), .B (n_8305), .Y (n_11575));
OR2X1 g125666(.A (n_18909), .B (n_25228), .Y (n_10624));
INVX4 g125700(.A (n_9629), .Y (n_10023));
INVX4 g125744(.A (n_9498), .Y (n_20864));
NAND2X1 g125789(.A (n_8420), .B (n_14490), .Y (n_9495));
INVX1 g125792(.A (n_35043), .Y (n_24786));
CLKBUFX1 g125796(.A (n_35044), .Y (n_30668));
INVX1 g125802(.A (n_23487), .Y (n_29445));
INVX1 g125810(.A (n_9490), .Y (n_29191));
INVX1 g125895(.A (n_28874), .Y (n_29172));
INVX1 g125906(.A (n_8677), .Y (n_27462));
INVX1 g125915(.A (n_8989), .Y (n_10003));
INVX1 g125918(.A (n_8989), .Y (n_10002));
INVX1 g125930(.A (n_29427), .Y (n_25748));
NAND2X1 g125951(.A (n_9483), .B (n_9482), .Y (n_11816));
INVX1 g126024(.A (n_8981), .Y (n_20218));
AND2X1 g125200(.A (n_9122), .B (n_9475), .Y (n_9476));
NAND2X1 g126065(.A (n_8979), .B (n_9474), .Y (n_9994));
NAND2X1 g126091(.A (n_7810), .B (n_8277), .Y (n_9473));
INVX1 g126138(.A (n_26238), .Y (n_28747));
INVX1 g126165(.A (n_23138), .Y (n_28319));
INVX1 g126282(.A (n_8313), .Y (n_25862));
INVX1 g126283(.A (n_8313), .Y (n_15026));
INVX1 g126308(.A (n_8614), .Y (n_25229));
INVX1 g126309(.A (n_8614), .Y (n_20688));
INVX1 g126312(.A (n_9458), .Y (n_23176));
CLKBUFX1 g126330(.A (n_33378), .Y (n_28808));
CLKBUFX1 g126332(.A (n_10063), .Y (n_30197));
INVX1 g126334(.A (n_29604), .Y (n_9455));
INVX1 g126344(.A (n_28468), .Y (n_27045));
INVX1 g126367(.A (n_29523), .Y (n_27192));
INVX2 g126373(.A (n_33738), .Y (n_28528));
INVX1 g126465(.A (n_29405), .Y (n_22528));
INVX1 g126524(.A (n_14850), .Y (n_14658));
INVX1 g126542(.A (n_9435), .Y (n_15076));
INVX1 g126547(.A (n_9436), .Y (n_26372));
INVX1 g126549(.A (n_9435), .Y (n_15288));
NAND2X1 g126653(.A (n_8635), .B (n_8996), .Y (n_9429));
AND2X1 g127527(.A (n_13709), .B (n_9373), .Y (n_9428));
INVX1 g126304(.A (n_8614), .Y (n_24028));
NAND2X2 g126768(.A (n_8486), .B (n_8189), .Y (n_16768));
NAND2X1 g126821(.A (n_8527), .B (n_9909), .Y (n_9426));
INVX1 g126841(.A (n_10799), .Y (n_16176));
NAND2X1 g126853(.A (n_8525), .B (n_9909), .Y (n_9425));
NAND2X1 g126856(.A (n_8464), .B (n_9909), .Y (n_9424));
NAND2X1 g126857(.A (n_8524), .B (n_9909), .Y (n_9422));
NAND2X1 g126861(.A (n_8523), .B (n_9909), .Y (n_9421));
NAND2X1 g126865(.A (n_8425), .B (n_30881), .Y (n_9420));
NAND2X1 g127523(.A (n_13354), .B (n_9373), .Y (n_9419));
NAND2X1 g126901(.A (n_8535), .B (n_9909), .Y (n_9418));
NAND3X1 g127007(.A (n_8393), .B (n_8155), .C (n_9413), .Y (n_9416));
NAND3X1 g127008(.A (n_8393), .B (n_8152), .C (n_9413), .Y (n_9415));
INVX1 g127038(.A (n_29381), .Y (n_29040));
INVX1 g127039(.A (n_29381), .Y (n_27956));
CLKBUFX1 g127065(.A (n_29505), .Y (n_27109));
INVX1 g127118(.A (n_30836), .Y (n_9404));
INVX1 g127151(.A (n_33807), .Y (n_24629));
NOR2X1 g127197(.A (n_8564), .B (n_6436), .Y (n_35695));
NOR2X1 g127237(.A (n_8571), .B (n_6436), .Y (n_9392));
NAND3X1 g127253(.A (n_9909), .B (n_7724), .C (n_8245), .Y (n_9391));
NAND3X1 g127260(.A (n_9387), .B (n_3105), .C (n_8245), .Y (n_9390));
NAND3X1 g127267(.A (n_9387), .B (n_11122), .C (n_8245), .Y (n_9388));
NAND3X1 g127272(.A (n_9387), .B (n_7819), .C (n_8245), .Y (n_9386));
NOR2X1 g127273(.A (n_8350), .B (n_9382), .Y (n_9385));
NAND3X1 g127284(.A (n_9909), .B (n_1003), .C (n_8245), .Y (n_9384));
NOR2X1 g127285(.A (n_8576), .B (n_9382), .Y (n_9383));
NAND2X1 g128269(.A (n_8336), .B (n_8460), .Y (n_9738));
NOR2X1 g127306(.A (n_8573), .B (n_12664), .Y (n_9381));
NOR2X1 g127323(.A (n_8566), .B (n_9382), .Y (n_9380));
NAND3X1 g127327(.A (n_9387), .B (n_11135), .C (n_8245), .Y (n_9379));
NOR2X1 g127369(.A (n_8569), .B (n_29486), .Y (n_9378));
NOR2X1 g127376(.A (n_8579), .B (n_6436), .Y (n_9377));
INVX4 g127394(.A (n_9375), .Y (n_11333));
INVX1 g127400(.A (n_16184), .Y (n_9883));
NAND2X1 g127408(.A (n_14168), .B (n_9373), .Y (n_9374));
NAND2X1 g127411(.A (P3_reg1[7] ), .B (n_8884), .Y (n_9372));
NOR2X1 g127422(.A (P3_reg_152), .B (n_11916), .Y (n_9371));
NAND2X1 g127431(.A (P3_reg2[10] ), .B (n_9373), .Y (n_9369));
NAND2X1 g127433(.A (n_13338), .B (n_8884), .Y (n_9368));
NAND2X1 g127444(.A (P3_reg1[11] ), .B (n_9373), .Y (n_9366));
NAND2X1 g127456(.A (n_13337), .B (n_9373), .Y (n_9364));
NAND2X1 g127459(.A (P3_reg2[6] ), .B (n_9373), .Y (n_9363));
NAND2X1 g127484(.A (P3_reg1[6] ), .B (n_8884), .Y (n_9362));
NAND2X1 g127485(.A (P3_reg2[18] ), .B (n_9373), .Y (n_9361));
AND2X1 g127487(.A (n_13365), .B (n_9373), .Y (n_9360));
NAND2X1 g127501(.A (P3_reg2[9] ), .B (n_9373), .Y (n_9358));
NAND2X1 g127515(.A (n_13332), .B (n_9373), .Y (n_9357));
NAND2X1 g127525(.A (n_13351), .B (n_9373), .Y (n_9356));
NAND2X1 g127532(.A (n_13361), .B (n_9373), .Y (n_9355));
NAND2X1 g127535(.A (n_13680), .B (n_8884), .Y (n_9354));
AND2X1 g127541(.A (n_13341), .B (n_9373), .Y (n_9353));
NAND2X1 g127549(.A (P3_reg1[1] ), .B (n_9373), .Y (n_9352));
AND2X1 g127552(.A (n_13678), .B (n_9373), .Y (n_9351));
NAND2X1 g127555(.A (P3_reg1[9] ), .B (n_8884), .Y (n_9350));
NAND2X1 g127557(.A (P3_reg1[3] ), .B (n_9373), .Y (n_9349));
NAND2X1 g127563(.A (n_13348), .B (n_8884), .Y (n_9348));
AND2X1 g127571(.A (n_10612), .B (n_8393), .Y (n_9347));
AND2X1 g127588(.A (n_9345), .B (n_8393), .Y (n_9346));
NAND2X1 g127598(.A (n_10032), .B (n_8393), .Y (n_9343));
AND2X1 g127599(.A (n_10617), .B (n_8393), .Y (n_9342));
AND2X1 g127600(.A (n_10601), .B (n_8393), .Y (n_9341));
AND2X1 g127601(.A (n_8193), .B (n_8393), .Y (n_9340));
AND2X1 g127615(.A (n_9337), .B (n_8393), .Y (n_9338));
INVX1 g127621(.A (n_16112), .Y (n_9336));
NOR2X1 g127627(.A (n_10116), .B (n_11916), .Y (n_9335));
NOR2X1 g127632(.A (n_3297), .B (n_7970), .Y (n_9334));
INVX1 g127644(.A (n_9333), .Y (n_9798));
INVX1 g127654(.A (n_12289), .Y (n_9624));
INVX2 g127662(.A (n_8710), .Y (n_17000));
NAND2X1 g127664(.A (P2_reg_108), .B (n_8393), .Y (n_9332));
NOR2X1 g127674(.A (n_8471), .B (n_8470), .Y (n_9793));
INVX2 g127676(.A (n_10752), .Y (n_16656));
CLKBUFX1 g127679(.A (n_10752), .Y (n_9792));
INVX1 g127681(.A (n_9171), .Y (n_9331));
NOR2X1 g127699(.A (P3_d_387), .B (n_11916), .Y (n_9329));
INVX1 g127717(.A (n_16096), .Y (n_9628));
INVX1 g127726(.A (n_16010), .Y (n_9327));
INVX1 g127758(.A (n_9322), .Y (n_9788));
NOR2X1 g127762(.A (P3_d_378), .B (n_8484), .Y (n_9321));
NOR2X1 g127778(.A (P3_d_397), .B (n_8484), .Y (n_9320));
NOR2X1 g127786(.A (n_10119), .B (n_11916), .Y (n_9318));
INVX1 g127790(.A (n_34936), .Y (n_9780));
NOR2X1 g127802(.A (n_9313), .B (n_7970), .Y (n_9314));
OR2X1 g127805(.A (n_35), .B (n_9310), .Y (n_9311));
NOR2X1 g127806(.A (P3_d), .B (n_8484), .Y (n_9309));
OR2X1 g127808(.A (P2_reg1[29] ), .B (n_9310), .Y (n_9308));
NOR2X1 g127810(.A (n_10112), .B (n_11916), .Y (n_9307));
INVX2 g127824(.A (n_9303), .Y (n_16012));
INVX1 g128198(.A (n_9302), .Y (n_16188));
NOR2X1 g127851(.A (P3_d_396), .B (n_11916), .Y (n_9300));
NOR2X1 g127852(.A (P3_d_393), .B (n_8484), .Y (n_9299));
BUFX1 g127856(.A (n_16983), .Y (n_10754));
NOR2X1 g127867(.A (P3_d_385), .B (n_11916), .Y (n_9298));
NAND2X1 g127868(.A (n_10602), .B (n_8393), .Y (n_9297));
AND2X1 g127869(.A (P2_reg2[11] ), .B (n_8393), .Y (n_9295));
AND2X1 g127928(.A (n_10582), .B (n_8884), .Y (n_9294));
OR2X1 g127937(.A (n_8011), .B (n_9310), .Y (n_9291));
NAND2X1 g127945(.A (n_10041), .B (n_8393), .Y (n_9290));
AND2X1 g127956(.A (n_10594), .B (n_8393), .Y (n_9288));
INVX1 g128182(.A (n_16163), .Y (n_9744));
AND2X1 g127967(.A (n_10100), .B (n_8884), .Y (n_9285));
INVX1 g127977(.A (n_9284), .Y (n_16577));
INVX2 g127998(.A (n_9195), .Y (n_9652));
INVX1 g128177(.A (n_16163), .Y (n_9281));
INVX1 g128178(.A (n_16163), .Y (n_9280));
INVX1 g128040(.A (n_9279), .Y (n_9684));
INVX1 g128052(.A (n_9278), .Y (n_9688));
INVX2 g128060(.A (n_9277), .Y (n_16186));
INVX1 g128064(.A (n_10484), .Y (n_17471));
NOR2X1 g128068(.A (P3_d_391), .B (n_8484), .Y (n_9276));
INVX1 g128083(.A (n_9274), .Y (n_9754));
INVX1 g128097(.A (n_9953), .Y (n_17007));
NOR2X1 g128102(.A (n_10114), .B (n_11916), .Y (n_9272));
INVX1 g128120(.A (n_9269), .Y (n_12437));
INVX1 g128135(.A (n_9962), .Y (n_16644));
INVX2 g128167(.A (n_8802), .Y (n_15908));
INVX1 g128175(.A (n_35663), .Y (n_9268));
INVX2 g128191(.A (n_8797), .Y (n_16646));
INVX1 g128214(.A (n_9264), .Y (n_9741));
NAND2X1 g128221(.A (P2_reg1[21] ), .B (n_8393), .Y (n_9263));
NOR2X1 g128227(.A (n_7932), .B (n_8462), .Y (n_16903));
NOR2X1 g128228(.A (n_3493), .B (n_7970), .Y (n_9262));
NOR2X1 g128270(.A (n_10103), .B (n_11916), .Y (n_9260));
INVX4 g128281(.A (n_15807), .Y (n_10706));
INVX4 g128332(.A (n_9257), .Y (n_9730));
INVX1 g128341(.A (n_34979), .Y (n_10006));
INVX1 g128352(.A (n_8788), .Y (n_9632));
NAND2X1 g128370(.A (n_8181), .B (n_8672), .Y (n_9253));
NOR2X1 g128371(.A (P2_reg_112), .B (n_9310), .Y (n_9252));
NOR2X1 g128399(.A (n_2975), .B (n_7970), .Y (n_9249));
INVX1 g128404(.A (n_10482), .Y (n_9725));
INVX4 g128480(.A (n_9247), .Y (n_9722));
INVX4 g128493(.A (n_34575), .Y (n_9720));
NOR2X1 g128501(.A (n_3269), .B (n_7970), .Y (n_9242));
NOR2X1 g128504(.A (P3_d_380), .B (n_8484), .Y (n_9240));
NOR2X1 g128505(.A (P3_d_379), .B (n_8484), .Y (n_9239));
NOR2X1 g128148(.A (n_8351), .B (n_8474), .Y (n_9238));
AND2X1 g128507(.A (n_10097), .B (n_8884), .Y (n_9237));
NOR2X1 g128521(.A (n_10110), .B (n_11916), .Y (n_9236));
NOR2X1 g128522(.A (n_2693), .B (n_9310), .Y (n_9235));
NOR2X1 g128525(.A (n_2379), .B (n_9310), .Y (n_9234));
NAND2X1 g128526(.A (n_9231), .B (n_8393), .Y (n_9232));
NOR2X1 g128532(.A (P3_d_398), .B (n_11916), .Y (n_9230));
CLKBUFX1 g128539(.A (n_9180), .Y (n_16984));
INVX2 g128548(.A (n_8780), .Y (n_16103));
INVX2 g128557(.A (n_9228), .Y (n_9627));
INVX1 g128568(.A (n_9226), .Y (n_9227));
INVX1 g128576(.A (n_9226), .Y (n_9701));
AND2X1 g128578(.A (P2_reg2[12] ), .B (n_8393), .Y (n_9225));
NAND2X2 g128589(.A (n_8454), .B (n_8472), .Y (n_9700));
INVX1 g128595(.A (n_9223), .Y (n_35253));
INVX1 g128600(.A (n_9223), .Y (n_16593));
INVX1 g128127(.A (n_8799), .Y (n_9219));
OAI21X1 g128959(.A0 (P2_reg1[28] ), .A1 (n_8168), .B0 (n_8448), .Y(n_9212));
CLKBUFX1 g128116(.A (n_9211), .Y (n_9749));
NAND2X1 g128980(.A (n_8444), .B (n_8443), .Y (n_10709));
AOI21X1 g128981(.A0 (n_9209), .A1 (n_8442), .B0 (n_8441), .Y(n_9210));
NOR2X1 g129072(.A (n_8449), .B (n_8169), .Y (n_9207));
NOR2X1 g129075(.A (n_8451), .B (n_8066), .Y (n_9206));
NOR2X1 g129082(.A (n_8438), .B (n_8156), .Y (n_9205));
AOI22X1 g129120(.A0 (n_10696), .A1 (n_4040), .B0 (n_6051), .B1(n_9676), .Y (n_9204));
AOI22X1 g129126(.A0 (n_10671), .A1 (n_4844), .B0 (n_6382), .B1(n_9676), .Y (n_9203));
INVX2 g128074(.A (n_16102), .Y (n_9755));
AOI22X1 g129132(.A0 (n_10696), .A1 (n_33901), .B0 (n_6480), .B1(n_9676), .Y (n_9201));
NAND2X1 g129200(.A (n_8363), .B (n_7578), .Y (n_11834));
NAND2X1 g129203(.A (n_8412), .B (n_7630), .Y (n_11831));
NAND3X1 g129273(.A (n_8371), .B (n_7890), .C (n_7888), .Y (n_10967));
NAND3X1 g129313(.A (n_8331), .B (n_8366), .C (n_8364), .Y (n_10946));
NAND3X1 g129337(.A (n_8416), .B (n_7814), .C (n_7812), .Y (n_10979));
NAND3X1 g129363(.A (n_8421), .B (n_7880), .C (n_7878), .Y (n_10977));
NAND3X1 g129383(.A (n_8422), .B (n_7885), .C (n_7883), .Y (n_10948));
NAND3X1 g129398(.A (n_8417), .B (n_7850), .C (n_7848), .Y (n_10983));
NAND3X1 g129410(.A (n_8374), .B (n_7905), .C (n_7903), .Y (n_10962));
NAND3X1 g129411(.A (n_8332), .B (n_7895), .C (n_7893), .Y (n_10981));
AOI22X1 g129489(.A0 (n_3063), .A1 (n_10676), .B0 (n_9676), .B1(n_11097), .Y (n_9197));
AOI22X1 g129501(.A0 (n_3176), .A1 (n_10676), .B0 (n_9676), .B1(n_3314), .Y (n_9194));
NAND2X1 g128293(.A (n_32294), .B (n_32295), .Y (n_9733));
NAND4X1 g126888(.A (n_32254), .B (n_34650), .C (n_7674), .D(n_32255), .Y (n_9960));
INVX1 g127962(.A (n_9286), .Y (n_9761));
AOI22X1 g129492(.A0 (n_3165), .A1 (n_10676), .B0 (n_9676), .B1(n_190), .Y (n_9190));
AND2X1 g125160(.A (n_14810), .B (n_13330), .Y (n_9188));
NOR2X1 g127289(.A (n_8574), .B (n_8899), .Y (n_9186));
INVX2 g126018(.A (n_8981), .Y (n_10573));
NAND2X1 g125131(.A (n_14810), .B (n_13721), .Y (n_9185));
CLKBUFX1 g125928(.A (n_29427), .Y (n_29568));
INVX1 g125893(.A (n_8677), .Y (n_29684));
AND2X1 g125062(.A (n_14810), .B (n_13709), .Y (n_9184));
NAND2X2 g127777(.A (n_8182), .B (n_8455), .Y (n_9785));
INVX1 g125803(.A (n_23487), .Y (n_30184));
INVX1 g128206(.A (n_16297), .Y (n_9742));
INVX1 g127744(.A (n_8851), .Y (n_11092));
CLKBUFX3 g127725(.A (n_16010), .Y (n_10717));
NOR2X1 g128591(.A (P3_d_382), .B (n_11916), .Y (n_9182));
INVX1 g128534(.A (n_9180), .Y (n_9181));
NAND2X1 g124971(.A (n_9122), .B (n_9178), .Y (n_9179));
NOR2X1 g127695(.A (P3_d_399), .B (n_8484), .Y (n_9177));
NAND2X1 g124966(.A (n_9122), .B (P2_reg_108), .Y (n_9176));
AOI22X1 g129447(.A0 (n_2872), .A1 (n_10676), .B0 (n_9676), .B1(n_2772), .Y (n_9173));
INVX2 g125641(.A (n_9172), .Y (n_9503));
CLKBUFX1 g127689(.A (n_9171), .Y (n_16904));
AOI22X1 g129125(.A0 (n_10671), .A1 (n_4288), .B0 (n_6393), .B1(n_9676), .Y (n_9169));
AND2X1 g127666(.A (n_13387), .B (n_9373), .Y (n_9167));
AND2X1 g124945(.A (n_9122), .B (n_9165), .Y (n_9166));
INVX4 g125599(.A (n_29027), .Y (n_9625));
AND2X1 g125580(.A (n_18289), .B (n_9337), .Y (n_9163));
OR2X1 g124929(.A (n_9162), .B (n_28785), .Y (n_26756));
AND2X1 g128541(.A (n_10578), .B (n_8884), .Y (n_9161));
INVX2 g127638(.A (n_8860), .Y (n_16011));
AND2X1 g125543(.A (n_18289), .B (n_9345), .Y (n_9159));
INVX1 g126534(.A (n_14956), .Y (n_25563));
INVX1 g126528(.A (n_14956), .Y (n_28659));
INVX1 g127620(.A (n_16112), .Y (n_10758));
NAND2X2 g125513(.A (n_8981), .B (n_8644), .Y (n_14550));
INVX1 g127170(.A (n_33807), .Y (n_27234));
NAND2X2 g128520(.A (n_8173), .B (n_8468), .Y (n_16064));
OR2X1 g127594(.A (n_4130), .B (n_9310), .Y (n_9154));
NOR2X1 g127590(.A (P2_reg3[3] ), .B (n_9310), .Y (n_9152));
INVX1 g127058(.A (n_29505), .Y (n_22762));
AND2X1 g127567(.A (n_13201), .B (n_9373), .Y (n_9149));
CLKBUFX1 g128414(.A (n_16357), .Y (n_10485));
INVX2 g129432(.A (n_15841), .Y (n_9683));
NAND2X1 g124925(.A (n_32341), .B (P1_d_98), .Y (n_9146));
NAND2X1 g124935(.A (n_32480), .B (n_7975), .Y (n_9145));
NAND2X1 g124947(.A (n_9122), .B (n_9142), .Y (n_9143));
AND2X1 g124948(.A (n_9122), .B (n_9139), .Y (n_9141));
AND2X1 g124952(.A (n_9122), .B (n_10452), .Y (n_9137));
NAND2X1 g124957(.A (n_9122), .B (n_9135), .Y (n_9136));
NAND2X1 g124973(.A (n_9122), .B (n_9132), .Y (n_9133));
NOR2X1 g124975(.A (n_29427), .B (n_8989), .Y (n_10049));
AND2X1 g124978(.A (n_14810), .B (n_13213), .Y (n_9131));
AND2X1 g124979(.A (n_9122), .B (P2_reg1[13] ), .Y (n_9130));
AND2X1 g124980(.A (n_9122), .B (n_10435), .Y (n_9128));
NAND2X1 g124985(.A (n_9122), .B (n_10363), .Y (n_9127));
AND2X1 g124986(.A (n_9122), .B (n_10443), .Y (n_9126));
NAND2X1 g124987(.A (n_14810), .B (P3_reg1[7] ), .Y (n_9125));
NAND2X1 g124988(.A (n_14810), .B (n_13354), .Y (n_9124));
AND2X1 g124993(.A (n_9122), .B (n_9121), .Y (n_9123));
AND2X1 g124994(.A (n_14810), .B (n_13365), .Y (n_9120));
AND2X1 g124996(.A (n_9122), .B (P2_reg1[10] ), .Y (n_9119));
AND2X1 g125001(.A (n_9122), .B (P2_reg1[15] ), .Y (n_9117));
AND2X1 g125003(.A (n_9122), .B (P2_reg1[17] ), .Y (n_9114));
AND2X1 g125012(.A (n_14810), .B (n_13209), .Y (n_9111));
AND2X1 g125013(.A (n_14810), .B (n_13211), .Y (n_9110));
AND2X1 g125014(.A (n_9122), .B (P2_reg1[18] ), .Y (n_9109));
AND2X1 g125015(.A (n_9122), .B (P2_reg1[19] ), .Y (n_9108));
AND2X1 g125016(.A (n_9122), .B (P2_reg1[1] ), .Y (n_9106));
NAND2X1 g125020(.A (n_9122), .B (n_9231), .Y (n_9105));
AND2X1 g125021(.A (n_9122), .B (n_9103), .Y (n_9104));
AND2X1 g125022(.A (n_9122), .B (n_9101), .Y (n_9102));
NAND2X1 g125023(.A (n_14810), .B (P3_reg1[6] ), .Y (n_9100));
NAND2X1 g125024(.A (n_9122), .B (n_9097), .Y (n_9099));
AND2X1 g125025(.A (n_9122), .B (P2_reg1[27] ), .Y (n_9096));
AND2X1 g125028(.A (n_9122), .B (P2_reg1[22] ), .Y (n_9095));
AND2X1 g125029(.A (n_9122), .B (n_9773), .Y (n_9094));
AND2X1 g125030(.A (n_9122), .B (n_9092), .Y (n_9093));
AND2X1 g125031(.A (n_9122), .B (P2_reg1[2] ), .Y (n_9091));
NAND2X1 g125033(.A (n_9122), .B (P2_reg1[4] ), .Y (n_9090));
AND2X1 g125034(.A (n_9122), .B (n_9088), .Y (n_9089));
AND2X1 g125035(.A (n_9122), .B (P2_reg1[5] ), .Y (n_9087));
NAND2X1 g125041(.A (n_14810), .B (n_13683), .Y (n_9086));
AND2X1 g125042(.A (n_9122), .B (P2_reg1[9] ), .Y (n_9085));
AND2X1 g125043(.A (n_14810), .B (P3_reg1[16] ), .Y (n_9083));
AND2X1 g125045(.A (n_9122), .B (n_9081), .Y (n_9082));
AND2X1 g125049(.A (n_14810), .B (n_13216), .Y (n_9080));
AND2X1 g125053(.A (n_14810), .B (n_13678), .Y (n_9079));
AND2X1 g125060(.A (n_14810), .B (n_13203), .Y (n_9078));
NAND2X1 g125063(.A (n_14810), .B (n_13359), .Y (n_9077));
AND2X1 g125065(.A (n_14810), .B (n_13698), .Y (n_9076));
NOR2X1 g125077(.A (n_29427), .B (n_29505), .Y (n_30050));
AND2X1 g125078(.A (n_14810), .B (n_13681), .Y (n_9074));
NAND2X1 g125080(.A (n_14810), .B (n_13351), .Y (n_9073));
AND2X1 g125084(.A (n_9122), .B (n_9071), .Y (n_9072));
INVX4 g125094(.A (n_27100), .Y (n_26382));
AND2X1 g125114(.A (n_9122), .B (n_9067), .Y (n_9068));
NAND2X1 g125117(.A (n_14810), .B (P3_reg1[18] ), .Y (n_9066));
INVX1 g125120(.A (n_9613), .Y (n_9563));
NAND2X1 g125135(.A (n_9122), .B (n_9794), .Y (n_9065));
AND2X1 g125143(.A (n_14810), .B (n_13212), .Y (n_9064));
NAND2X1 g125147(.A (n_14810), .B (n_13367), .Y (n_9063));
NAND2X1 g125149(.A (n_14810), .B (n_13357), .Y (n_9062));
NAND2X1 g125150(.A (n_14810), .B (n_13355), .Y (n_9061));
NAND2X1 g125151(.A (n_14810), .B (n_13353), .Y (n_9060));
AND2X1 g125154(.A (n_14810), .B (P3_reg1[4] ), .Y (n_9059));
AND2X1 g125156(.A (n_14810), .B (n_13697), .Y (n_9058));
AND2X1 g125161(.A (n_14810), .B (n_13202), .Y (n_9057));
NAND2X1 g125166(.A (n_14810), .B (P3_reg1[11] ), .Y (n_9056));
NAND2X1 g125167(.A (n_14810), .B (n_13680), .Y (n_9055));
NAND2X1 g125168(.A (n_14810), .B (n_13679), .Y (n_9054));
AND2X1 g125172(.A (n_14810), .B (n_13724), .Y (n_9053));
AND2X1 g125174(.A (n_14810), .B (n_13692), .Y (n_9052));
AND2X1 g125176(.A (n_14810), .B (n_13690), .Y (n_9051));
NAND2X1 g125177(.A (n_14810), .B (P3_reg1[9] ), .Y (n_9050));
NAND2X1 g125178(.A (n_14810), .B (n_13677), .Y (n_9049));
NAND2X1 g125180(.A (n_14810), .B (P3_reg1[1] ), .Y (n_9048));
NAND2X1 g125182(.A (n_14810), .B (n_13673), .Y (n_9047));
AND2X1 g125186(.A (n_14810), .B (n_13341), .Y (n_9046));
NAND2X1 g125190(.A (n_14810), .B (P3_reg1[17] ), .Y (n_9045));
AND2X1 g125191(.A (n_14810), .B (n_13699), .Y (n_9044));
AND2X1 g125194(.A (n_14810), .B (n_13377), .Y (n_9043));
NAND2X1 g125196(.A (n_9122), .B (P2_reg1[21] ), .Y (n_9042));
NAND2X1 g125197(.A (n_14810), .B (P3_reg1[3] ), .Y (n_9041));
AND2X1 g125199(.A (n_14810), .B (n_13687), .Y (n_9040));
OAI22X1 g125252(.A0 (n_9520), .A1 (n_9038), .B0 (n_3601), .B1(n_8309), .Y (n_9039));
NAND2X1 g127546(.A (n_13721), .B (n_8884), .Y (n_9035));
NAND2X1 g125430(.A (n_11138), .B (n_14317), .Y (n_9034));
NOR2X1 g125434(.A (n_8642), .B (n_7745), .Y (n_9032));
NAND2X1 g125440(.A (n_11138), .B (n_13336), .Y (n_9031));
NAND2X1 g125454(.A (n_11138), .B (n_13329), .Y (n_9030));
NAND2X1 g125455(.A (n_11138), .B (n_13352), .Y (n_9028));
NAND2X1 g125456(.A (n_11138), .B (n_13334), .Y (n_9027));
NAND2X1 g125457(.A (n_11138), .B (n_13344), .Y (n_9026));
NAND2X1 g125458(.A (n_11138), .B (n_13343), .Y (n_9025));
NAND2X1 g125459(.A (n_11138), .B (n_13368), .Y (n_9024));
NAND2X1 g125460(.A (n_11138), .B (n_13335), .Y (n_9023));
INVX2 g128359(.A (n_16926), .Y (n_17906));
NAND2X1 g125487(.A (n_13378), .B (n_19108), .Y (n_9021));
AND2X1 g125488(.A (n_11138), .B (n_10578), .Y (n_9020));
NAND2X1 g125495(.A (n_13375), .B (n_19108), .Y (n_9019));
AND2X1 g125500(.A (n_18289), .B (n_10617), .Y (n_9018));
NAND2X1 g125510(.A (n_18289), .B (n_10601), .Y (n_9017));
NAND2X1 g125526(.A (n_9337), .B (n_10848), .Y (n_9016));
NAND2X1 g127006(.A (n_8390), .B (n_9909), .Y (n_9015));
NOR2X1 g125545(.A (n_8958), .B (n_7967), .Y (n_9507));
NAND2X1 g125547(.A (n_8190), .B (n_10848), .Y (n_9014));
AND2X1 g125571(.A (n_11138), .B (n_10100), .Y (n_9013));
AND2X1 g125576(.A (n_11138), .B (n_10582), .Y (n_9011));
AND2X1 g125579(.A (n_11138), .B (n_10097), .Y (n_9010));
INVX1 g125585(.A (n_26160), .Y (n_26748));
INVX1 g125586(.A (n_26160), .Y (n_9009));
INVX2 g125614(.A (n_34952), .Y (n_9626));
INVX1 g125624(.A (n_34771), .Y (n_9003));
INVX1 g125626(.A (n_9001), .Y (n_29065));
INVX1 g125629(.A (n_9001), .Y (n_30438));
INVX1 g125632(.A (n_9001), .Y (n_28948));
NAND2X1 g125663(.A (n_8309), .B (n_25881), .Y (n_11812));
NAND2X1 g125665(.A (n_25540), .B (n_8309), .Y (n_10203));
INVX8 g125708(.A (n_8998), .Y (n_9629));
CLKBUFX1 g125795(.A (n_35044), .Y (n_25968));
INVX1 g125801(.A (n_26660), .Y (n_9493));
INVX1 g125804(.A (n_26660), .Y (n_23487));
INVX1 g125812(.A (n_28431), .Y (n_9490));
CLKBUFX1 g125889(.A (n_8990), .Y (n_30454));
CLKBUFX1 g125896(.A (n_8990), .Y (n_28874));
CLKBUFX1 g125898(.A (n_8989), .Y (n_27614));
NOR2X1 g126071(.A (n_8979), .B (n_8426), .Y (n_8980));
INVX1 g126142(.A (n_29553), .Y (n_29955));
INVX1 g126166(.A (n_30200), .Y (n_23138));
CLKBUFX1 g126169(.A (n_26553), .Y (n_27842));
INVX1 g126172(.A (n_8966), .Y (n_26920));
INVX1 g126174(.A (n_8966), .Y (n_29000));
INVX1 g126321(.A (n_8958), .Y (n_26142));
INVX1 g126323(.A (n_8958), .Y (n_27326));
INVX1 g126324(.A (n_8958), .Y (n_25424));
INVX1 g126328(.A (n_33340), .Y (n_10063));
INVX1 g126345(.A (n_33340), .Y (n_28468));
CLKBUFX1 g126368(.A (n_33738), .Y (n_29523));
INVX1 g126385(.A (n_14641), .Y (n_15029));
INVX1 g126398(.A (n_33713), .Y (n_15073));
INVX1 g126409(.A (n_33713), .Y (n_15252));
INVX1 g126412(.A (n_8949), .Y (n_30530));
INVX1 g126459(.A (n_25881), .Y (n_30109));
NOR2X1 g126495(.A (n_6495), .B (n_8948), .Y (n_8947));
INVX1 g126513(.A (n_8946), .Y (n_9441));
INVX1 g126525(.A (n_8945), .Y (n_14850));
INVX1 g126561(.A (n_8945), .Y (n_9978));
INVX1 g126573(.A (n_8945), .Y (n_14743));
INVX8 g126618(.A (n_25540), .Y (n_21328));
INVX1 g126624(.A (n_26458), .Y (n_25867));
INVX2 g126636(.A (n_8942), .Y (n_9431));
INVX1 g126639(.A (n_25082), .Y (n_8940));
INVX1 g126647(.A (n_25942), .Y (n_9430));
BUFX3 g126649(.A (n_25942), .Y (n_25220));
NAND2X1 g126701(.A (n_8295), .B (n_8326), .Y (n_8936));
AND2X1 g126810(.A (n_8230), .B (n_8933), .Y (n_8935));
AND2X1 g126828(.A (n_8236), .B (n_8933), .Y (n_8934));
INVX1 g126292(.A (n_8313), .Y (n_25067));
INVX1 g127021(.A (n_8382), .Y (n_28798));
CLKBUFX1 g127036(.A (n_26665), .Y (n_30557));
INVX1 g127055(.A (n_8927), .Y (n_27522));
NOR2X1 g129328(.A (n_3343), .B (n_7998), .Y (n_8925));
CLKBUFX1 g127119(.A (n_13952), .Y (n_30836));
CLKBUFX1 g127147(.A (n_33802), .Y (n_27993));
INVX2 g127176(.A (n_30180), .Y (n_29388));
NOR2X1 g127183(.A (n_8258), .B (n_8916), .Y (n_8917));
NOR2X1 g127194(.A (n_8272), .B (n_8899), .Y (n_8915));
NOR2X1 g127201(.A (n_8267), .B (n_6436), .Y (n_8914));
NOR2X1 g127203(.A (n_8241), .B (n_8893), .Y (n_8912));
NOR2X1 g127208(.A (n_8254), .B (n_8893), .Y (n_8911));
NAND2X1 g129322(.A (P2_reg2[29] ), .B (n_7864), .Y (n_8910));
NOR2X1 g127219(.A (n_8255), .B (n_8893), .Y (n_8909));
NOR2X1 g127228(.A (n_8260), .B (n_8893), .Y (n_8906));
NOR2X1 g127232(.A (n_8262), .B (n_6436), .Y (n_8905));
NOR2X1 g127243(.A (n_8249), .B (n_12664), .Y (n_8903));
NOR2X1 g127274(.A (n_8280), .B (n_12664), .Y (n_8901));
NOR2X1 g127278(.A (n_8320), .B (n_8899), .Y (n_8900));
NOR2X1 g127293(.A (n_8240), .B (n_6436), .Y (n_8898));
NOR2X1 g127296(.A (n_8269), .B (n_6436), .Y (n_8897));
NOR2X1 g127302(.A (n_8252), .B (n_8916), .Y (n_8896));
NOR2X1 g127303(.A (n_8251), .B (n_6436), .Y (n_8895));
NOR2X1 g127320(.A (n_8281), .B (n_8893), .Y (n_8894));
NOR2X1 g127329(.A (n_8244), .B (n_8916), .Y (n_8892));
NOR2X1 g127335(.A (n_8029), .B (n_8916), .Y (n_8891));
NOR2X1 g127336(.A (n_8242), .B (n_6436), .Y (n_8890));
NOR2X1 g127338(.A (n_8248), .B (n_8893), .Y (n_8889));
NOR2X1 g127344(.A (n_8243), .B (n_8899), .Y (n_8888));
NOR2X1 g127362(.A (n_8247), .B (n_8899), .Y (n_8887));
INVX2 g127395(.A (n_9483), .Y (n_9375));
CLKBUFX1 g127401(.A (n_9474), .Y (n_16184));
NAND2X1 g127424(.A (n_13677), .B (n_8884), .Y (n_8886));
NAND2X1 g127438(.A (P3_reg2[13] ), .B (n_8884), .Y (n_8885));
NAND2X1 g127477(.A (n_13359), .B (n_8884), .Y (n_8883));
NAND2X1 g127478(.A (n_13357), .B (n_8884), .Y (n_8882));
NAND2X1 g127482(.A (n_13683), .B (n_8884), .Y (n_8881));
NAND2X1 g127489(.A (n_8245), .B (n_15723), .Y (n_8880));
NAND2X1 g127497(.A (n_13498), .B (n_8884), .Y (n_8878));
NAND2X1 g127509(.A (n_13358), .B (n_8884), .Y (n_8877));
NAND2X1 g127510(.A (n_14513), .B (n_8884), .Y (n_8876));
NAND2X1 g127518(.A (n_13353), .B (n_8884), .Y (n_8875));
NAND2X1 g127519(.A (n_13366), .B (n_8884), .Y (n_8874));
NAND2X1 g127521(.A (n_13367), .B (n_8884), .Y (n_8873));
NAND2X1 g127537(.A (n_13679), .B (n_8884), .Y (n_8872));
NAND2X1 g127556(.A (n_13502), .B (n_8884), .Y (n_8871));
NAND2X1 g127558(.A (n_13355), .B (n_8884), .Y (n_8870));
NAND2X1 g127560(.A (P3_reg1[17] ), .B (n_8884), .Y (n_8869));
AND2X1 g127572(.A (n_9209), .B (n_8393), .Y (n_8868));
AND2X1 g127612(.A (n_9512), .B (n_8393), .Y (n_8867));
INVX2 g127622(.A (n_8561), .Y (n_16112));
NAND2X1 g127624(.A (n_9139), .B (n_8393), .Y (n_8865));
NAND2X1 g127625(.A (P2_reg2[3] ), .B (n_8393), .Y (n_8864));
NAND2X1 g127629(.A (n_4160), .B (n_8393), .Y (n_8862));
NAND2X1 g127630(.A (P2_reg_104), .B (n_8393), .Y (n_8861));
NAND2X1 g127639(.A (n_8291), .B (n_8210), .Y (n_8860));
CLKBUFX1 g127645(.A (n_35714), .Y (n_9333));
INVX1 g127646(.A (n_35714), .Y (n_8859));
NAND2X1 g127648(.A (n_9135), .B (n_8393), .Y (n_8858));
INVX1 g127655(.A (n_15820), .Y (n_12289));
NOR2X1 g127675(.A (P1_d_121), .B (n_7871), .Y (n_8857));
NAND2X2 g127680(.A (n_7945), .B (n_8199), .Y (n_10752));
NAND2X1 g127690(.A (n_8172), .B (n_8176), .Y (n_9171));
NAND2X1 g127698(.A (n_14135), .B (n_8844), .Y (n_8856));
NAND2X1 g127739(.A (n_9592), .B (n_8393), .Y (n_8853));
NOR2X1 g127763(.A (P1_d_118), .B (n_7871), .Y (n_8849));
NAND2X1 g127764(.A (P2_reg1[11] ), .B (n_9413), .Y (n_8847));
NAND2X1 g127767(.A (P2_reg1[12] ), .B (n_9413), .Y (n_8846));
NAND2X1 g127779(.A (P2_reg1[13] ), .B (n_8844), .Y (n_8845));
NAND2X1 g127780(.A (n_9586), .B (n_8393), .Y (n_8843));
NAND2X1 g127781(.A (P2_reg1[15] ), .B (n_8844), .Y (n_8842));
NAND2X1 g127782(.A (P2_reg1[16] ), .B (n_8393), .Y (n_8841));
NAND2X1 g127799(.A (P2_reg1[23] ), .B (n_9413), .Y (n_8840));
NOR2X1 g127800(.A (P1_d_103), .B (n_7871), .Y (n_8839));
NOR2X1 g127803(.A (P1_d_105), .B (n_7871), .Y (n_8838));
NAND2X1 g127807(.A (n_9178), .B (n_8393), .Y (n_8837));
NAND2X1 g127819(.A (n_4237), .B (n_9413), .Y (n_8835));
NAND2X1 g127820(.A (P2_reg1[8] ), .B (n_8393), .Y (n_8833));
NAND2X1 g127821(.A (P2_reg1[9] ), .B (n_8844), .Y (n_8832));
NAND2X1 g127826(.A (n_10563), .B (n_8844), .Y (n_8831));
NAND2X1 g128199(.A (n_7942), .B (n_8195), .Y (n_9302));
CLKBUFX1 g127832(.A (n_8381), .Y (n_11089));
INVX1 g127848(.A (n_8829), .Y (n_11401));
CLKBUFX1 g127857(.A (n_8828), .Y (n_16983));
INVX1 g127858(.A (n_8828), .Y (n_16624));
NAND2X1 g127861(.A (n_10610), .B (n_8393), .Y (n_8827));
NAND2X1 g127864(.A (P2_reg1[3] ), .B (n_9413), .Y (n_8826));
NAND2X1 g127865(.A (n_10607), .B (n_8393), .Y (n_8825));
NAND2X1 g127871(.A (n_4475), .B (n_8393), .Y (n_8824));
NAND2X1 g127919(.A (n_9067), .B (n_8844), .Y (n_8823));
NAND2X1 g127921(.A (n_4344), .B (n_8393), .Y (n_8822));
NAND2X1 g127923(.A (P2_reg1[10] ), .B (n_8393), .Y (n_8821));
NAND2X1 g127924(.A (P2_reg2[9] ), .B (n_8393), .Y (n_8820));
NAND2X1 g127925(.A (n_9097), .B (n_8393), .Y (n_8819));
NOR2X1 g127926(.A (n_3157), .B (n_7871), .Y (n_8818));
INVX2 g127933(.A (n_15906), .Y (n_9292));
NAND2X1 g127936(.A (P2_reg2[10] ), .B (n_8393), .Y (n_8817));
NAND2X1 g127943(.A (n_9549), .B (n_9413), .Y (n_8816));
NAND2X1 g127949(.A (n_9590), .B (n_9413), .Y (n_8815));
NAND2X1 g127951(.A (n_9565), .B (n_9413), .Y (n_8814));
NAND2X1 g127952(.A (P2_reg2[19] ), .B (n_8844), .Y (n_8813));
NAND2X1 g127954(.A (P2_reg1[17] ), .B (n_8844), .Y (n_8812));
NAND2X1 g127969(.A (n_10047), .B (n_8393), .Y (n_8811));
NAND2X1 g127970(.A (n_9101), .B (n_8393), .Y (n_8810));
NOR2X1 g127988(.A (n_2553), .B (n_7871), .Y (n_8809));
NAND4X1 g128000(.A (n_32086), .B (n_7658), .C (n_32087), .D (n_7689),.Y (n_9195));
INVX1 g128008(.A (n_16435), .Y (n_9198));
INVX1 g128020(.A (n_8436), .Y (n_9199));
NAND2X2 g128333(.A (n_7940), .B (n_8194), .Y (n_9257));
NAND2X1 g128041(.A (n_7791), .B (n_8203), .Y (n_9279));
NAND2X1 g128061(.A (n_7721), .B (n_8202), .Y (n_9277));
INVX2 g128066(.A (n_35343), .Y (n_15918));
INVX2 g128076(.A (n_8522), .Y (n_16102));
NAND2X1 g128168(.A (n_7955), .B (n_8204), .Y (n_8802));
INVX1 g128117(.A (n_8801), .Y (n_9211));
INVX2 g128121(.A (n_7810), .Y (n_9269));
CLKBUFX1 g128136(.A (n_11404), .Y (n_9962));
NAND2X1 g128149(.A (n_9121), .B (n_8844), .Y (n_8798));
NAND2X2 g128183(.A (n_8208), .B (n_8170), .Y (n_16163));
NAND3X1 g128192(.A (n_8196), .B (n_7675), .C (n_7700), .Y (n_8797));
NAND2X1 g128200(.A (P2_reg2[1] ), .B (n_9413), .Y (n_8796));
INVX2 g128208(.A (n_8517), .Y (n_16297));
INVX1 g128215(.A (n_16585), .Y (n_9264));
NAND2X1 g128222(.A (P2_reg1[20] ), .B (n_8844), .Y (n_8795));
NAND2X1 g128253(.A (P2_reg1[6] ), .B (n_8393), .Y (n_8794));
NAND2X1 g128263(.A (n_9103), .B (n_8393), .Y (n_8793));
NAND2X1 g128271(.A (n_9165), .B (n_8393), .Y (n_8792));
INVX2 g128282(.A (n_8625), .Y (n_15807));
NAND2X1 g128344(.A (n_9132), .B (n_8393), .Y (n_8791));
NAND2X1 g128345(.A (n_10604), .B (n_8393), .Y (n_8790));
INVX1 g128346(.A (n_8788), .Y (n_35423));
NAND2X1 g128355(.A (n_9071), .B (n_8393), .Y (n_8787));
NAND2X2 g128389(.A (n_7936), .B (n_8186), .Y (n_9036));
INVX1 g128405(.A (n_16079), .Y (n_10482));
NAND2X1 g128472(.A (n_9142), .B (n_8393), .Y (n_8785));
INVX1 g128499(.A (n_8784), .Y (n_9243));
NAND2X1 g128502(.A (n_9597), .B (n_8844), .Y (n_8783));
NAND2X1 g128503(.A (n_10082), .B (n_9413), .Y (n_8782));
CLKBUFX1 g128099(.A (n_34172), .Y (n_9953));
NAND2X1 g128513(.A (n_9595), .B (n_8393), .Y (n_8781));
NAND2X1 g128540(.A (n_8054), .B (n_8187), .Y (n_9180));
NAND2X1 g128549(.A (n_32269), .B (n_32270), .Y (n_8780));
NAND2X1 g128567(.A (n_10613), .B (n_8393), .Y (n_8779));
NAND2X1 g128577(.A (n_8188), .B (n_7959), .Y (n_9226));
NAND2X1 g128579(.A (n_3724), .B (n_8393), .Y (n_8778));
NAND2X1 g128603(.A (P2_reg1[31] ), .B (n_8844), .Y (n_8777));
NAND2X1 g128604(.A (n_9475), .B (n_8844), .Y (n_8776));
INVX1 g128622(.A (n_35008), .Y (n_30537));
INVX1 g128637(.A (n_8719), .Y (n_31523));
INVX1 g128641(.A (n_8719), .Y (n_27557));
INVX1 g128645(.A (n_8719), .Y (n_31564));
INVX1 g128648(.A (n_31064), .Y (n_27008));
INVX1 g128651(.A (n_31064), .Y (n_29681));
INVX1 g128733(.A (n_11916), .Y (n_9859));
AOI21X1 g128960(.A0 (n_10890), .A1 (n_8485), .B0 (n_8166), .Y(n_8762));
AOI21X1 g128982(.A0 (P2_reg1[21] ), .A1 (n_9692), .B0 (n_8085), .Y(n_8761));
AOI21X1 g128991(.A0 (n_10886), .A1 (n_7694), .B0 (n_8016), .Y(n_32562));
NAND2X1 g129031(.A (n_7929), .B (n_8165), .Y (n_8759));
NAND2X1 g129077(.A (n_8162), .B (n_7668), .Y (n_8758));
NAND2X1 g129080(.A (n_8052), .B (n_8157), .Y (n_8757));
INVX2 g128084(.A (n_16375), .Y (n_9274));
INVX2 g128065(.A (n_35344), .Y (n_10484));
INVX2 g128053(.A (n_8756), .Y (n_9278));
NAND2X1 g129202(.A (n_8093), .B (n_7586), .Y (n_11823));
NAND2X1 g129210(.A (n_8116), .B (n_7626), .Y (n_11607));
NAND2X1 g129223(.A (n_8106), .B (n_7633), .Y (n_11821));
NOR2X1 g129247(.A (P2_reg_113), .B (n_8125), .Y (n_8755));
NAND2X1 g129251(.A (n_8102), .B (n_7629), .Y (n_11829));
NAND2X1 g129256(.A (n_8109), .B (n_7622), .Y (n_11594));
NAND3X1 g129264(.A (n_8033), .B (n_8148), .C (n_8146), .Y (n_11151));
NAND4X1 g129266(.A (n_8130), .B (n_8128), .C (n_8131), .D (n_7617),.Y (n_11157));
NAND2X1 g129323(.A (n_8099), .B (n_7628), .Y (n_11605));
NOR2X1 g129329(.A (n_3494), .B (n_7998), .Y (n_8754));
NOR2X1 g129331(.A (P2_reg_109), .B (n_8125), .Y (n_8753));
NOR2X1 g129333(.A (n_3449), .B (n_7998), .Y (n_8752));
NAND2X1 g127412(.A (P3_reg2[30] ), .B (n_8884), .Y (n_8750));
NAND3X1 g129367(.A (n_8015), .B (n_8140), .C (n_8138), .Y (n_11160));
NAND2X1 g129371(.A (n_8119), .B (n_7591), .Y (n_11601));
NAND2X1 g129377(.A (n_8112), .B (n_7634), .Y (n_11817));
NAND2X1 g129385(.A (n_8027), .B (n_7623), .Y (n_11599));
NAND2X1 g129391(.A (n_8020), .B (n_7625), .Y (n_11826));
NAND2X1 g129396(.A (n_10653), .B (n_7864), .Y (n_8749));
NAND2X1 g129401(.A (n_8096), .B (n_7624), .Y (n_11592));
NAND2X1 g129416(.A (n_10602), .B (n_7864), .Y (n_8747));
NAND2X1 g129419(.A (n_8090), .B (n_7631), .Y (n_11588));
NAND2X1 g129422(.A (n_8031), .B (n_7619), .Y (n_11819));
INVX1 g129442(.A (n_8744), .Y (n_8745));
NAND2X1 g128001(.A (n_4367), .B (n_9413), .Y (n_8743));
NAND4X1 g129479(.A (n_7041), .B (n_8453), .C (n_8741), .D (n_8452),.Y (n_8742));
AOI22X1 g129480(.A0 (n_10676), .A1 (n_32509), .B0 (n_9676), .B1(n_10838), .Y (n_8740));
AND2X1 g129538(.A (n_7216), .B (n_9676), .Y (n_8739));
AND2X1 g129797(.A (n_8078), .B (n_8050), .Y (n_8738));
CLKBUFX1 g127978(.A (n_16084), .Y (n_9284));
AND2X1 g129814(.A (n_8084), .B (n_8429), .Y (n_8736));
AND2X1 g129817(.A (n_8075), .B (n_7901), .Y (n_8735));
AND2X1 g129837(.A (n_8082), .B (n_8434), .Y (n_8734));
INVX1 g127964(.A (n_8526), .Y (n_9286));
NAND3X1 g129208(.A (n_8035), .B (n_8144), .C (n_8142), .Y (n_11155));
NAND2X1 g127948(.A (n_10081), .B (n_9413), .Y (n_8732));
INVX1 g127934(.A (n_15906), .Y (n_8729));
INVX1 g126842(.A (n_9637), .Y (n_10799));
NOR2X1 g127319(.A (n_8022), .B (n_8899), .Y (n_8726));
NAND2X1 g125121(.A (n_35043), .B (n_10067), .Y (n_9613));
NAND2X2 g127825(.A (n_35444), .B (n_35445), .Y (n_9303));
NOR2X1 g127262(.A (n_8259), .B (n_8893), .Y (n_8721));
CLKBUFX1 g125809(.A (n_28431), .Y (n_30559));
NAND2X1 g127709(.A (n_14133), .B (n_8844), .Y (n_8716));
NOR2X1 g127245(.A (n_8229), .B (n_12664), .Y (n_8715));
NOR2X1 g125745(.A (n_18218), .B (n_18227), .Y (n_9498));
INVX2 g127759(.A (n_8850), .Y (n_9322));
NOR2X1 g127239(.A (n_8214), .B (n_8893), .Y (n_8714));
NAND2X2 g127727(.A (n_8279), .B (n_8224), .Y (n_16010));
INVX1 g127040(.A (n_26665), .Y (n_29381));
INVX2 g128601(.A (n_8492), .Y (n_9223));
NAND2X1 g128593(.A (P2_reg_95), .B (n_9413), .Y (n_8713));
CLKBUFX1 g125643(.A (n_34770), .Y (n_28597));
INVX1 g125653(.A (n_34770), .Y (n_14162));
INVX1 g125633(.A (n_34770), .Y (n_9001));
INVX1 g128347(.A (n_8788), .Y (n_8711));
NAND2X1 g127663(.A (n_7943), .B (n_8198), .Y (n_8710));
NAND2X1 g127650(.A (P2_reg_107), .B (n_9413), .Y (n_8709));
NAND2X1 g128558(.A (n_8174), .B (n_7820), .Y (n_9228));
INVX2 g125605(.A (n_34951), .Y (n_29027));
INVX1 g125593(.A (n_34951), .Y (n_26160));
AND2X1 g129823(.A (n_8080), .B (n_8346), .Y (n_8705));
NAND2X1 g127631(.A (n_9599), .B (n_8393), .Y (n_8704));
CLKBUFX1 g126552(.A (n_8945), .Y (n_9435));
INVX4 g128395(.A (n_33268), .Y (n_15749));
INVX1 g126548(.A (n_8945), .Y (n_9436));
INVX4 g126541(.A (n_8945), .Y (n_14956));
INVX1 g128360(.A (n_9956), .Y (n_16926));
INVX1 g129003(.A (n_8469), .Y (n_8703));
INVX4 g126466(.A (n_25881), .Y (n_29405));
INVX1 g126457(.A (n_25881), .Y (n_27902));
INVX1 g126449(.A (n_25881), .Y (n_29155));
INVX1 g126316(.A (n_8313), .Y (n_9458));
NAND2X1 g128506(.A (n_13645), .B (n_8844), .Y (n_8699));
NAND2X2 g128482(.A (n_8179), .B (n_7958), .Y (n_9247));
CLKBUFX1 g125619(.A (n_34770), .Y (n_29068));
INVX1 g128415(.A (n_8697), .Y (n_16357));
INVX2 g129434(.A (n_8746), .Y (n_15841));
NAND2X1 g124937(.A (n_8677), .B (n_33734), .Y (n_14349));
NAND2X1 g124951(.A (n_8678), .B (n_8321), .Y (n_24563));
NAND2X1 g124981(.A (n_32342), .B (n_7333), .Y (n_8695));
NAND2X1 g128398(.A (P2_reg2[18] ), .B (n_8844), .Y (n_8693));
NAND3X1 g129423(.A (n_8122), .B (n_8136), .C (n_8134), .Y (n_11153));
NAND2X2 g125109(.A (n_8692), .B (n_8333), .Y (n_27100));
INVX1 g126337(.A (n_33340), .Y (n_29604));
NAND2X1 g125148(.A (n_8010), .B (n_8322), .Y (n_21677));
OR4X1 g125321(.A (n_8009), .B (n_10196), .C (n_7587), .D (n_34802),.Y (n_10644));
INVX4 g125480(.A (n_14810), .Y (n_9557));
NAND2X1 g125519(.A (n_28136), .B (n_27042), .Y (n_12142));
NOR2X1 g125521(.A (n_28528), .B (n_1054), .Y (n_11197));
NAND2X1 g125546(.A (n_28492), .B (n_8687), .Y (n_12380));
INVX1 g125554(.A (n_8686), .Y (n_14638));
INVX1 g125622(.A (n_34770), .Y (n_27169));
INVX4 g125642(.A (n_34770), .Y (n_9172));
INVX1 g125655(.A (n_27743), .Y (n_8682));
INVX1 g125657(.A (n_27256), .Y (n_24752));
OR2X1 g125664(.A (n_8009), .B (n_34802), .Y (n_11158));
NOR2X1 g125709(.A (n_8680), .B (n_7775), .Y (n_8998));
INVX1 g125813(.A (n_35043), .Y (n_28431));
INVX1 g128634(.A (n_34336), .Y (n_31544));
INVX2 g125856(.A (n_8678), .Y (n_28785));
INVX1 g125920(.A (n_8677), .Y (n_8989));
NOR2X1 g129088(.A (n_7915), .B (n_7697), .Y (n_8672));
INVX1 g126068(.A (n_9162), .Y (n_8671));
INVX1 g126108(.A (n_28492), .Y (n_8977));
INVX1 g126113(.A (n_8319), .Y (n_29619));
INVX1 g126117(.A (n_8668), .Y (n_29008));
INVX1 g126119(.A (n_8668), .Y (n_27340));
INVX1 g126132(.A (n_30563), .Y (n_8664));
CLKBUFX1 g126141(.A (n_26238), .Y (n_30636));
INVX1 g126145(.A (n_26238), .Y (n_29553));
INVX1 g126147(.A (n_8661), .Y (n_28374));
INVX1 g126148(.A (n_8661), .Y (n_29253));
INVX1 g126152(.A (n_33991), .Y (n_28523));
INVX1 g126154(.A (n_33991), .Y (n_27662));
INVX1 g126167(.A (n_29725), .Y (n_30200));
INVX1 g126171(.A (n_29725), .Y (n_26553));
INVX1 g126195(.A (n_28136), .Y (n_8965));
INVX1 g126254(.A (n_8314), .Y (n_18909));
INVX1 g126325(.A (n_33378), .Y (n_8958));
INVX4 g126404(.A (n_33713), .Y (n_15110));
INVX1 g126413(.A (n_15147), .Y (n_8949));
INVX1 g126429(.A (n_8309), .Y (n_19108));
BUFX3 g126516(.A (n_8643), .Y (n_8946));
INVX1 g126517(.A (n_8643), .Y (n_8644));
NAND2X1 g126574(.A (n_7994), .B (n_8283), .Y (n_8945));
INVX1 g126580(.A (n_8305), .Y (n_26870));
NAND2X1 g126584(.A (n_7822), .B (n_8008), .Y (n_8642));
INVX4 g126619(.A (n_8358), .Y (n_25540));
BUFX3 g126623(.A (n_8641), .Y (n_25942));
CLKBUFX1 g126625(.A (n_8641), .Y (n_26458));
INVX1 g126659(.A (n_26052), .Y (n_23771));
INVX1 g126683(.A (n_26052), .Y (n_24451));
INVX1 g126688(.A (n_26052), .Y (n_24247));
INVX4 g126303(.A (n_8614), .Y (n_22821));
NAND2X1 g126762(.A (n_7797), .B (P2_d_378), .Y (n_8635));
INVX2 g127032(.A (n_8382), .Y (n_25756));
NOR2X1 g129330(.A (P2_reg2[25] ), .B (n_7917), .Y (n_8633));
INVX1 g127134(.A (n_8284), .Y (n_30230));
NAND4X1 g128283(.A (n_7381), .B (n_7199), .C (n_7222), .D (n_7477),.Y (n_8625));
INVX4 g127177(.A (n_33807), .Y (n_30180));
NAND3X1 g127184(.A (n_9909), .B (n_10169), .C (n_8245), .Y (n_8623));
NAND3X1 g127187(.A (n_9909), .B (n_3337), .C (n_8245), .Y (n_8622));
NAND3X1 g127191(.A (n_9909), .B (n_10150), .C (n_8245), .Y (n_8619));
NAND3X1 g127192(.A (n_9909), .B (n_3716), .C (n_8245), .Y (n_8618));
NAND3X1 g127198(.A (n_9909), .B (n_4011), .C (n_8245), .Y (n_8616));
NAND3X1 g127214(.A (n_9909), .B (P1_reg2[1] ), .C (n_8245), .Y(n_8615));
NAND3X1 g127231(.A (n_9909), .B (n_3259), .C (n_8245), .Y (n_8613));
NAND3X1 g127250(.A (n_9909), .B (n_10221), .C (n_8245), .Y (n_8612));
NAND3X1 g127257(.A (n_9909), .B (n_10154), .C (n_8245), .Y (n_8611));
NAND3X1 g127259(.A (n_9909), .B (n_7706), .C (n_8245), .Y (n_8610));
INVX1 g126278(.A (n_8614), .Y (n_14490));
NAND3X1 g127269(.A (n_9909), .B (n_10566), .C (n_8245), .Y (n_8609));
NAND3X1 g127276(.A (n_9909), .B (n_3958), .C (n_8245), .Y (n_8606));
NAND3X1 g127277(.A (n_9909), .B (n_10148), .C (n_8245), .Y (n_8605));
NAND3X1 g127301(.A (n_9909), .B (n_10173), .C (n_8245), .Y (n_8604));
NAND3X1 g127307(.A (n_9909), .B (P1_reg_174), .C (n_8245), .Y(n_8603));
NAND3X1 g127326(.A (n_9909), .B (P1_reg1[24] ), .C (n_8245), .Y(n_8602));
NAND3X1 g127374(.A (n_9909), .B (n_4534), .C (n_8245), .Y (n_8601));
INVX1 g127383(.A (n_9482), .Y (n_8737));
NAND2X1 g127414(.A (n_10245), .B (n_8598), .Y (n_8600));
NAND2X1 g127423(.A (P1_reg2[19] ), .B (n_8598), .Y (n_8599));
NAND2X1 g127427(.A (n_4151), .B (n_8598), .Y (n_8597));
NOR2X1 g128254(.A (P1_d_114), .B (n_8557), .Y (n_8596));
NAND2X1 g127430(.A (n_4445), .B (n_8598), .Y (n_8595));
NAND2X1 g127436(.A (P1_reg2[14] ), .B (n_8598), .Y (n_8593));
NAND2X1 g127439(.A (n_11141), .B (n_8245), .Y (n_8592));
NAND2X1 g127442(.A (n_11120), .B (n_8245), .Y (n_8591));
NAND2X1 g127443(.A (n_3235), .B (n_8245), .Y (n_8589));
NAND2X1 g127446(.A (n_10893), .B (n_8245), .Y (n_8588));
NAND2X1 g127448(.A (n_11148), .B (n_8245), .Y (n_8587));
NAND2X1 g127449(.A (n_10858), .B (n_8598), .Y (n_8586));
NAND2X1 g127452(.A (n_11144), .B (n_8245), .Y (n_8585));
NAND2X1 g127453(.A (n_10546), .B (n_8245), .Y (n_8584));
NAND2X1 g127455(.A (P1_reg2[30] ), .B (n_8245), .Y (n_8582));
NAND2X1 g127458(.A (n_3470), .B (n_8598), .Y (n_8581));
NAND2X1 g127461(.A (n_3416), .B (n_8245), .Y (n_8580));
NAND2X1 g127462(.A (P1_reg1[12] ), .B (n_8575), .Y (n_8579));
NAND2X1 g127463(.A (n_4561), .B (n_8245), .Y (n_8578));
NAND2X1 g127467(.A (n_10215), .B (n_8598), .Y (n_8577));
NAND2X1 g127486(.A (n_10189), .B (n_8575), .Y (n_8576));
NAND2X1 g127488(.A (n_10182), .B (n_8245), .Y (n_8574));
NAND2X1 g127494(.A (P1_reg_173), .B (n_8575), .Y (n_8573));
NAND2X1 g127496(.A (P1_reg1[16] ), .B (n_8245), .Y (n_8572));
NAND2X1 g127499(.A (n_3693), .B (n_8245), .Y (n_8571));
NAND2X1 g127503(.A (P1_reg1[19] ), .B (n_8245), .Y (n_8569));
NAND2X1 g127504(.A (P1_reg2[16] ), .B (n_8245), .Y (n_8568));
NAND2X1 g127512(.A (n_13322), .B (n_8245), .Y (n_8567));
NAND2X1 g127513(.A (n_10175), .B (n_8575), .Y (n_8566));
NAND2X1 g127528(.A (n_13635), .B (n_8245), .Y (n_8565));
NAND2X1 g127540(.A (n_10136), .B (n_8245), .Y (n_8564));
NAND2X1 g127562(.A (n_10219), .B (n_8245), .Y (n_8562));
NAND2X1 g127623(.A (n_35925), .B (n_35926), .Y (n_8561));
INVX2 g127656(.A (n_8360), .Y (n_15820));
NOR2X1 g127696(.A (P1_d), .B (n_8552), .Y (n_8560));
NOR2X1 g127710(.A (P1_d_107), .B (n_8552), .Y (n_8559));
NOR2X1 g127713(.A (P1_d_108), .B (n_8557), .Y (n_8558));
NOR2X1 g127721(.A (P1_d_109), .B (n_8552), .Y (n_8556));
NOR2X1 g127737(.A (P1_d_112), .B (n_8552), .Y (n_8555));
NOR2X1 g127738(.A (P1_d_113), .B (n_8557), .Y (n_8554));
NOR2X1 g127741(.A (P1_d_116), .B (n_8552), .Y (n_8553));
INVX1 g127747(.A (n_16291), .Y (n_8551));
NOR2X1 g127749(.A (P1_d_98), .B (n_8552), .Y (n_8550));
INVX1 g127760(.A (n_8239), .Y (n_8850));
NOR2X1 g127783(.A (P1_d_124), .B (n_8552), .Y (n_8549));
NOR2X1 g127785(.A (P1_d_126), .B (n_8552), .Y (n_8547));
NOR2X1 g127795(.A (P1_d_127), .B (n_8552), .Y (n_8545));
NOR2X1 g127796(.A (P1_d_128), .B (n_8552), .Y (n_8544));
NOR2X1 g127797(.A (P1_d_100), .B (n_8557), .Y (n_8542));
NOR2X1 g127798(.A (P1_d_101), .B (n_8557), .Y (n_8541));
NOR2X1 g127804(.A (P1_d_106), .B (n_8552), .Y (n_8540));
NAND2X1 g127835(.A (n_8552), .B (n_641), .Y (n_8537));
INVX2 g127849(.A (n_15812), .Y (n_8829));
AND2X1 g127866(.A (n_7737), .B (n_8245), .Y (n_8535));
INVX1 g127883(.A (n_30569), .Y (n_31410));
INVX1 g127913(.A (n_8528), .Y (n_28588));
INVX1 g127914(.A (n_8528), .Y (n_30619));
AND2X1 g127927(.A (n_10822), .B (n_8245), .Y (n_8527));
NAND2X2 g127935(.A (n_7934), .B (n_7786), .Y (n_15906));
NOR2X1 g127972(.A (P1_reg3[3] ), .B (n_7415), .Y (n_8525));
AND2X1 g127985(.A (n_10880), .B (n_8245), .Y (n_8524));
AND2X1 g127986(.A (n_7546), .B (n_8245), .Y (n_8523));
NAND2X1 g128055(.A (n_7954), .B (n_7937), .Y (n_8756));
NAND2X1 g128077(.A (n_7783), .B (n_7717), .Y (n_8522));
NAND2X2 g128086(.A (n_7766), .B (n_7949), .Y (n_16375));
INVX1 g128118(.A (n_8232), .Y (n_8801));
INVX1 g128137(.A (n_8518), .Y (n_11404));
NAND2X2 g128209(.A (n_7723), .B (n_7960), .Y (n_8517));
INVX1 g128217(.A (n_8329), .Y (n_16293));
NOR2X1 g128223(.A (n_8515), .B (n_7415), .Y (n_8516));
NAND2X2 g128354(.A (n_7789), .B (n_7727), .Y (n_8788));
INVX1 g128407(.A (n_16079), .Y (n_8513));
NOR2X1 g128409(.A (n_8511), .B (n_7415), .Y (n_8512));
INVX1 g128437(.A (n_26002), .Y (n_8505));
INVX1 g128440(.A (n_26002), .Y (n_31620));
INVX1 g128447(.A (n_30099), .Y (n_29769));
INVX1 g128459(.A (n_31878), .Y (n_31936));
NOR2X1 g128523(.A (P1_d_123), .B (n_8557), .Y (n_8493));
NAND2X1 g128602(.A (n_35438), .B (n_35439), .Y (n_8492));
INVX1 g128615(.A (n_34336), .Y (n_27485));
INVX1 g128617(.A (n_34336), .Y (n_30956));
INVX1 g128633(.A (n_34336), .Y (n_30353));
INVX1 g128653(.A (n_31236), .Y (n_31064));
AOI21X1 g128657(.A0 (n_10546), .A1 (n_8485), .B0 (n_7963), .Y(n_8486));
INVX1 g128629(.A (n_34739), .Y (n_30914));
INVX2 g128130(.A (n_8479), .Y (n_8799));
INVX2 g128112(.A (n_33999), .Y (n_8803));
NAND2X1 g128990(.A (n_7693), .B (n_7914), .Y (n_8474));
NOR2X1 g128103(.A (P1_d_99), .B (n_8552), .Y (n_8473));
NOR2X1 g128996(.A (n_7911), .B (n_7596), .Y (n_8472));
NAND2X1 g129000(.A (n_7811), .B (n_7430), .Y (n_8471));
NAND2X1 g129001(.A (n_7695), .B (n_7919), .Y (n_8470));
NAND2X1 g129004(.A (n_7927), .B (n_7368), .Y (n_8469));
AOI21X1 g129010(.A0 (n_8467), .A1 (n_7476), .B0 (n_7909), .Y(n_8468));
INVX1 g128095(.A (n_35625), .Y (n_8465));
AND2X1 g127984(.A (n_13167), .B (n_8245), .Y (n_8464));
NAND2X1 g129035(.A (n_7316), .B (n_8002), .Y (n_8462));
NOR2X1 g129071(.A (n_7978), .B (n_7924), .Y (n_8460));
AOI21X1 g129079(.A0 (n_8458), .A1 (n_8163), .B0 (n_7918), .Y(n_32294));
NAND2X1 g129081(.A (n_7923), .B (n_7666), .Y (n_8457));
INVX1 g126190(.A (n_29725), .Y (n_8966));
INVX1 g129107(.A (n_8175), .Y (n_8455));
AOI21X1 g129114(.A0 (n_9103), .A1 (n_8335), .B0 (n_7799), .Y(n_8454));
INVX1 g126182(.A (n_29725), .Y (n_26548));
NAND2X1 g129194(.A (n_7856), .B (n_7284), .Y (n_11584));
NAND2X1 g129198(.A (n_7859), .B (n_6871), .Y (n_11357));
NAND3X1 g129214(.A (n_7285), .B (n_8453), .C (n_8452), .Y (n_11596));
NAND2X1 g129231(.A (n_7858), .B (n_7283), .Y (n_11805));
NOR2X1 g129240(.A (P2_reg2[26] ), .B (n_7917), .Y (n_8451));
NOR2X1 g129263(.A (P2_reg2[24] ), .B (n_7917), .Y (n_8449));
NAND2X1 g129316(.A (n_8447), .B (n_8442), .Y (n_8448));
NAND2X1 g129327(.A (n_9602), .B (n_8445), .Y (n_8446));
NAND2X1 g129334(.A (n_9132), .B (n_8445), .Y (n_8444));
NAND2X1 g129335(.A (n_10601), .B (n_8442), .Y (n_8443));
NOR2X1 g129345(.A (n_335), .B (n_7917), .Y (n_8441));
NAND2X1 g129347(.A (n_10032), .B (n_8442), .Y (n_8440));
NOR2X1 g129354(.A (n_242), .B (n_7917), .Y (n_8438));
NAND2X1 g128021(.A (n_7507), .B (n_7962), .Y (n_8436));
INVX1 g126162(.A (n_29725), .Y (n_28364));
INVX2 g129435(.A (n_8039), .Y (n_8746));
OR2X1 g129443(.A (n_7644), .B (n_9676), .Y (n_8744));
NAND4X1 g129457(.A (n_8434), .B (n_8433), .C (n_8432), .D (n_8431),.Y (n_8435));
NAND4X1 g129459(.A (n_8429), .B (n_8428), .C (n_7429), .D (n_8427),.Y (n_8430));
CLKBUFX1 g128009(.A (n_8979), .Y (n_16435));
CLKBUFX1 g127402(.A (n_8426), .Y (n_9474));
NAND4X1 g127396(.A (n_35453), .B (n_7545), .C (n_7504), .D (n_7204),.Y (n_9483));
NOR2X1 g127990(.A (n_2837), .B (n_7415), .Y (n_8425));
INVX1 g129551(.A (n_15850), .Y (n_8424));
AND2X1 g129796(.A (n_7844), .B (n_7886), .Y (n_8422));
AND2X1 g129798(.A (n_7836), .B (n_7881), .Y (n_8421));
NAND2X1 g129802(.A (n_6961), .B (n_8413), .Y (n_8420));
INVX1 g127979(.A (n_8418), .Y (n_16084));
AND2X1 g129818(.A (n_7869), .B (n_7851), .Y (n_8417));
AND2X1 g129820(.A (n_7834), .B (n_7815), .Y (n_8416));
NAND2X1 g129841(.A (n_6952), .B (n_8413), .Y (n_14260));
AOI21X1 g129846(.A0 (n_8113), .A1 (addr_429), .B0 (n_7845), .Y(n_8412));
AOI22X1 g129847(.A0 (n_6352), .A1 (n_8409), .B0 (n_7616), .B1(n_628), .Y (n_8410));
AOI22X1 g129850(.A0 (n_6332), .A1 (n_8407), .B0 (n_7616), .B1(addr_461), .Y (n_8408));
INVX2 g127957(.A (n_8526), .Y (n_15815));
INVX1 g126118(.A (n_8668), .Y (n_27335));
INVX1 g128465(.A (n_33123), .Y (n_8401));
INVX1 g130030(.A (n_8399), .Y (n_9668));
CLKBUFX1 g126326(.A (n_33378), .Y (n_29090));
INVX1 g128464(.A (n_33123), .Y (n_8397));
INVX1 g128446(.A (n_30099), .Y (n_31245));
NOR2X1 g127944(.A (P1_d_117), .B (n_8552), .Y (n_8395));
NAND3X1 g127364(.A (n_9909), .B (n_10854), .C (n_8245), .Y (n_8394));
NAND2X1 g129192(.A (n_7785), .B (n_6857), .Y (n_11360));
INVX1 g130031(.A (n_8399), .Y (n_9677));
NAND3X1 g127356(.A (n_9909), .B (n_10191), .C (n_8245), .Y (n_8392));
INVX1 g127905(.A (n_7827), .Y (n_31360));
AND2X1 g127920(.A (n_7575), .B (n_8245), .Y (n_8390));
INVX1 g127884(.A (n_30569), .Y (n_31178));
NAND3X1 g126843(.A (n_8387), .B (n_6973), .C (n_32892), .Y (n_9637));
NAND4X1 g127859(.A (n_32128), .B (n_32129), .C (n_7161), .D (n_7496),.Y (n_8828));
INVX2 g126026(.A (n_8324), .Y (n_8981));
INVX1 g127843(.A (n_8384), .Y (n_8830));
INVX1 g127827(.A (n_8381), .Y (n_16100));
NOR2X1 g127809(.A (P1_d_119), .B (n_8552), .Y (n_8380));
NOR2X1 g127811(.A (P1_d_120), .B (n_8552), .Y (n_8379));
NOR2X1 g127801(.A (P1_d_104), .B (n_8557), .Y (n_8378));
INVX1 g125897(.A (n_8677), .Y (n_8990));
INVX1 g128646(.A (n_8377), .Y (n_8719));
NOR2X1 g127784(.A (P1_d_125), .B (n_8552), .Y (n_8376));
INVX1 g128640(.A (n_8377), .Y (n_31402));
AND2X1 g129813(.A (n_7842), .B (n_7906), .Y (n_8374));
INVX1 g128618(.A (n_34336), .Y (n_30958));
NAND3X1 g127256(.A (n_9909), .B (n_7730), .C (n_8245), .Y (n_8372));
INVX1 g128619(.A (n_34336), .Y (n_30360));
INVX1 g125805(.A (n_35043), .Y (n_26660));
INVX1 g125794(.A (n_35043), .Y (n_28890));
AND2X1 g129810(.A (n_7966), .B (n_7891), .Y (n_8371));
INVX1 g127746(.A (n_16291), .Y (n_8851));
NOR2X1 g127740(.A (P1_d_115), .B (n_8552), .Y (n_8370));
NOR2X1 g128594(.A (P1_d_110), .B (n_8552), .Y (n_8369));
OR2X1 g125656(.A (n_33378), .B (n_10196), .Y (n_27743));
NAND4X1 g129450(.A (n_8330), .B (n_8366), .C (n_8365), .D (n_8364),.Y (n_8367));
AOI21X1 g129845(.A0 (n_8113), .A1 (n_8361), .B0 (n_7916), .Y(n_8363));
INVX1 g126692(.A (n_26052), .Y (n_25122));
INVX1 g127912(.A (n_8528), .Y (n_31482));
CLKBUFX1 g127657(.A (n_8360), .Y (n_15817));
CLKBUFX1 g126644(.A (n_8641), .Y (n_25082));
INVX1 g126637(.A (n_8641), .Y (n_8942));
NOR2X1 g127640(.A (P1_d_102), .B (n_8552), .Y (n_8357));
INVX1 g128400(.A (n_16079), .Y (n_8356));
INVX1 g125557(.A (n_8375), .Y (n_9122));
INVX1 g128466(.A (n_33123), .Y (n_8355));
NOR2X1 g127626(.A (P1_d_122), .B (n_8557), .Y (n_8354));
INVX1 g127136(.A (n_30230), .Y (n_29551));
INVX1 g127120(.A (n_8352), .Y (n_13952));
INVX4 g126460(.A (n_28158), .Y (n_25881));
INVX1 g127128(.A (n_8352), .Y (n_8922));
NAND2X1 g129116(.A (n_7921), .B (n_7566), .Y (n_8351));
NAND2X1 g127559(.A (P1_reg1[14] ), .B (n_8575), .Y (n_8350));
INVX2 g126418(.A (n_15110), .Y (n_14641));
NAND2X2 g128500(.A (n_8000), .B (n_7933), .Y (n_8784));
NAND4X1 g129454(.A (n_8346), .B (n_8345), .C (n_8344), .D (n_8343),.Y (n_8347));
INVX1 g128454(.A (n_31878), .Y (n_8340));
INVX1 g127048(.A (n_8718), .Y (n_26665));
INVX4 g126366(.A (n_28528), .Y (n_8954));
INVX1 g128416(.A (n_8337), .Y (n_8697));
AOI21X1 g129076(.A0 (n_9139), .A1 (n_8335), .B0 (n_7910), .Y(n_8336));
INVX1 g127026(.A (n_8382), .Y (n_26112));
INVX1 g130113(.A (n_9676), .Y (n_8696));
NAND2X1 g127554(.A (n_10152), .B (n_8245), .Y (n_8334));
NAND3X1 g125179(.A (n_8927), .B (n_8333), .C (n_29725), .Y (n_11353));
AND2X1 g129800(.A (n_7838), .B (n_7896), .Y (n_8332));
AND2X1 g129799(.A (n_7840), .B (n_8330), .Y (n_8331));
CLKBUFX1 g128216(.A (n_8329), .Y (n_16585));
NAND2X1 g125475(.A (n_8325), .B (n_7992), .Y (n_10984));
NAND2X2 g125484(.A (n_8004), .B (n_8309), .Y (n_14810));
NAND2X1 g128361(.A (n_7720), .B (n_7961), .Y (n_9956));
NAND2X1 g125528(.A (n_8004), .B (n_33713), .Y (n_11389));
NOR2X1 g125555(.A (n_3264), .B (n_8309), .Y (n_8686));
INVX1 g125563(.A (n_8375), .Y (n_9603));
NAND4X1 g125584(.A (n_7743), .B (n_7519), .C (n_8326), .D (n_7328),.Y (n_32481));
NAND2X1 g125618(.A (n_7997), .B (n_8306), .Y (n_14351));
NOR2X1 g125660(.A (n_33738), .B (n_33991), .Y (n_27256));
INVX4 g125998(.A (n_8325), .Y (n_18289));
AND2X1 g126027(.A (n_7752), .B (n_30897), .Y (n_8324));
NAND2X1 g126069(.A (n_8322), .B (n_8321), .Y (n_9162));
NAND2X1 g127539(.A (n_10140), .B (n_8245), .Y (n_8320));
INVX1 g126109(.A (n_8319), .Y (n_28492));
INVX1 g126124(.A (n_34693), .Y (n_8668));
BUFX3 g126146(.A (n_33991), .Y (n_26238));
INVX1 g126150(.A (n_33991), .Y (n_8661));
CLKBUFX1 g126197(.A (n_8316), .Y (n_28136));
NOR2X1 g126246(.A (n_7379), .B (n_7782), .Y (n_8680));
INVX1 g126261(.A (n_8314), .Y (n_10848));
INVX8 g126289(.A (n_8313), .Y (n_8614));
INVX1 g126381(.A (n_33713), .Y (n_11107));
NOR2X1 g126446(.A (n_7758), .B (n_7770), .Y (n_18227));
INVX4 g126469(.A (n_8306), .Y (n_28158));
NOR2X1 g126621(.A (n_7342), .B (n_7758), .Y (n_8358));
NOR2X1 g126652(.A (n_8304), .B (n_7759), .Y (n_8641));
INVX4 g126680(.A (n_8303), .Y (n_26052));
NAND2X1 g126763(.A (n_7744), .B (P3_d_377), .Y (n_8295));
INVX1 g127111(.A (n_8285), .Y (n_30369));
INVX1 g127099(.A (n_8286), .Y (n_28791));
AOI21X1 g128997(.A0 (P1_reg_172), .A1 (n_8177), .B0 (n_7699), .Y(n_8291));
INVX4 g127033(.A (n_26213), .Y (n_8382));
INVX4 g127049(.A (n_7981), .Y (n_8718));
INVX4 g127081(.A (n_8927), .Y (n_29505));
INVX2 g127093(.A (n_29150), .Y (n_26288));
NOR2X1 g128999(.A (n_7465), .B (n_7592), .Y (n_32269));
CLKBUFX1 g127101(.A (n_8286), .Y (n_30523));
INVX1 g127129(.A (n_8284), .Y (n_8352));
INVX1 g127141(.A (n_8283), .Y (n_8948));
NAND2X1 g127545(.A (n_10134), .B (n_8245), .Y (n_8281));
NAND2X1 g127511(.A (n_10156), .B (n_8245), .Y (n_8280));
AOI21X1 g129005(.A0 (P1_reg_173), .A1 (n_8177), .B0 (n_7703), .Y(n_8279));
INVX1 g127384(.A (n_8277), .Y (n_9482));
NAND4X1 g127403(.A (n_35453), .B (n_7203), .C (n_7196), .D (n_7158),.Y (n_8426));
NAND2X1 g127410(.A (n_10247), .B (n_8245), .Y (n_8275));
NAND2X1 g127417(.A (P1_reg1[30] ), .B (n_8245), .Y (n_8274));
AND2X1 g127418(.A (n_3333), .B (n_8245), .Y (n_8273));
NAND2X1 g127420(.A (n_3402), .B (n_8245), .Y (n_8272));
NAND2X1 g127421(.A (n_4554), .B (n_8245), .Y (n_8270));
NAND2X1 g127502(.A (n_10128), .B (n_8245), .Y (n_8269));
NAND2X1 g127426(.A (n_11136), .B (n_8245), .Y (n_8267));
NAND2X1 g127432(.A (n_4213), .B (n_8245), .Y (n_8266));
NAND2X1 g127434(.A (n_10171), .B (n_8245), .Y (n_8264));
NAND2X1 g127440(.A (n_4277), .B (n_8245), .Y (n_8263));
NAND2X1 g127457(.A (n_13640), .B (n_8245), .Y (n_8262));
NAND2X1 g127460(.A (n_3668), .B (n_8245), .Y (n_8261));
NAND2X1 g127469(.A (n_10205), .B (n_8245), .Y (n_8260));
NAND2X1 g127473(.A (n_10201), .B (n_8245), .Y (n_8259));
NAND2X1 g127475(.A (n_10161), .B (n_8245), .Y (n_8258));
NAND2X1 g127483(.A (P1_reg_180), .B (n_8245), .Y (n_8257));
NAND2X1 g127490(.A (n_10180), .B (n_8245), .Y (n_8256));
NAND2X1 g127491(.A (P1_reg1[0] ), .B (n_8245), .Y (n_8255));
NAND2X1 g127495(.A (n_10158), .B (n_8245), .Y (n_8254));
NAND2X1 g127507(.A (n_10165), .B (n_8245), .Y (n_8252));
NAND2X1 g127508(.A (P1_reg_172), .B (n_8245), .Y (n_8251));
NAND2X1 g127514(.A (n_10890), .B (n_8245), .Y (n_8250));
NAND2X1 g127534(.A (n_10144), .B (n_8245), .Y (n_8249));
NAND2X1 g127536(.A (n_10886), .B (n_8245), .Y (n_8248));
NAND2X1 g127544(.A (n_4215), .B (n_8245), .Y (n_8247));
AND2X1 g127550(.A (n_4920), .B (n_8245), .Y (n_8246));
NAND2X1 g127551(.A (n_10225), .B (n_8245), .Y (n_8244));
NAND2X1 g127553(.A (n_10197), .B (n_8245), .Y (n_8243));
NAND2X1 g127564(.A (n_10138), .B (n_8245), .Y (n_8242));
NAND2X1 g127568(.A (n_10223), .B (n_8245), .Y (n_8241));
NAND2X1 g127493(.A (n_10178), .B (n_8245), .Y (n_8240));
NAND2X2 g127658(.A (n_7514), .B (n_7735), .Y (n_8360));
NAND2X1 g128218(.A (n_7728), .B (n_7739), .Y (n_8329));
NAND2X2 g127748(.A (n_7725), .B (n_7569), .Y (n_16291));
NAND2X1 g127761(.A (n_7732), .B (n_7547), .Y (n_8239));
NAND3X1 g127834(.A (n_7731), .B (n_7502), .C (n_7145), .Y (n_8381));
NAND2X1 g127844(.A (n_35617), .B (n_35616), .Y (n_8384));
NAND2X1 g127850(.A (n_7513), .B (n_7713), .Y (n_15812));
NAND2X1 g127451(.A (n_11327), .B (n_8245), .Y (n_8238));
INVX1 g127877(.A (n_30403), .Y (n_30935));
INVX1 g127890(.A (n_31233), .Y (n_31160));
INVX1 g127903(.A (n_31360), .Y (n_31771));
AND2X1 g127946(.A (n_8207), .B (n_8245), .Y (n_8236));
AND2X1 g127953(.A (n_10885), .B (n_8245), .Y (n_8235));
NAND2X1 g127955(.A (n_13169), .B (n_8245), .Y (n_8234));
INVX1 g127981(.A (n_8233), .Y (n_8418));
NAND4X1 g128119(.A (n_7053), .B (n_7142), .C (n_7317), .D (n_7228),.Y (n_8232));
INVX8 g128719(.A (n_9373), .Y (n_11916));
INVX4 g128131(.A (n_8231), .Y (n_8479));
AND2X1 g128262(.A (n_10889), .B (n_8245), .Y (n_8230));
NAND2X1 g127465(.A (n_10187), .B (n_8245), .Y (n_8229));
NAND2X1 g127464(.A (n_4230), .B (n_8245), .Y (n_8228));
NAND2X2 g128408(.A (n_7712), .B (n_7738), .Y (n_16079));
NAND2X1 g128417(.A (n_7779), .B (n_7516), .Y (n_8337));
INVX1 g128430(.A (n_33125), .Y (n_30683));
INVX1 g128431(.A (n_33125), .Y (n_31099));
NAND2X1 g128528(.A (n_7957), .B (n_8245), .Y (n_8226));
NAND2X1 g128529(.A (n_13173), .B (n_8245), .Y (n_8225));
AOI21X1 g128953(.A0 (n_13173), .A1 (n_8209), .B0 (n_7435), .Y(n_8224));
INVX1 g128647(.A (n_35008), .Y (n_8377));
NAND2X1 g127445(.A (n_10897), .B (n_8245), .Y (n_8214));
AOI21X1 g128951(.A0 (n_3372), .A1 (n_8209), .B0 (n_7492), .Y(n_8210));
AOI21X1 g128952(.A0 (n_8207), .A1 (n_7638), .B0 (n_7606), .Y(n_8208));
AOI21X1 g128955(.A0 (n_8205), .A1 (n_8192), .B0 (n_7684), .Y(n_8206));
AOI21X1 g128962(.A0 (n_7444), .A1 (P2_reg2[9] ), .B0 (n_7590), .Y(n_8204));
NOR2X1 g128965(.A (n_7683), .B (n_7740), .Y (n_8203));
NOR2X1 g128966(.A (n_7463), .B (n_7682), .Y (n_8202));
NOR2X1 g128971(.A (n_7681), .B (n_7679), .Y (n_8200));
AOI21X1 g128972(.A0 (P3_reg2[18] ), .A1 (n_8183), .B0 (n_7678), .Y(n_8199));
AOI21X1 g128973(.A0 (n_13389), .A1 (n_8197), .B0 (n_7677), .Y(n_8198));
AOI21X1 g128974(.A0 (n_3072), .A1 (n_8197), .B0 (n_7574), .Y(n_8196));
NOR2X1 g128977(.A (n_7671), .B (n_7670), .Y (n_8195));
AOI21X1 g128983(.A0 (n_8193), .A1 (n_8192), .B0 (n_7687), .Y(n_8194));
AOI21X1 g128986(.A0 (n_8190), .A1 (n_7657), .B0 (n_7660), .Y(n_8191));
AOI22X1 g129012(.A0 (n_10211), .A1 (n_8177), .B0 (n_10245), .B1(n_7926), .Y (n_8189));
AOI21X1 g129018(.A0 (n_10180), .A1 (n_7722), .B0 (n_7594), .Y(n_8188));
NOR2X1 g129021(.A (n_7385), .B (n_7701), .Y (n_8187));
AOI21X1 g129023(.A0 (n_8185), .A1 (n_8192), .B0 (n_7663), .Y(n_8186));
AND2X1 g129026(.A (n_7258), .B (n_7665), .Y (n_8182));
AOI21X1 g129030(.A0 (n_9773), .A1 (n_8335), .B0 (n_7580), .Y(n_8181));
CLKBUFX1 g126198(.A (n_8316), .Y (n_29411));
AOI21X1 g129078(.A0 (P2_reg1[17] ), .A1 (n_7930), .B0 (n_7572), .Y(n_32295));
AOI21X1 g129091(.A0 (n_10171), .A1 (n_8177), .B0 (n_7698), .Y(n_8179));
AOI21X1 g129092(.A0 (n_10225), .A1 (n_8177), .B0 (n_7704), .Y(n_8178));
NOR2X1 g129103(.A (n_7360), .B (n_7696), .Y (n_8176));
NAND2X1 g129108(.A (n_7741), .B (n_7260), .Y (n_8175));
AOI21X1 g129109(.A0 (n_10175), .A1 (n_8177), .B0 (n_7608), .Y(n_8174));
AOI21X1 g129110(.A0 (P2_reg1[15] ), .A1 (n_7556), .B0 (n_7781), .Y(n_8173));
AOI21X1 g129115(.A0 (n_10178), .A1 (n_8177), .B0 (n_7656), .Y(n_8172));
NOR2X1 g129117(.A (n_7471), .B (n_7659), .Y (n_8170));
NOR2X1 g129168(.A (n_309), .B (n_8168), .Y (n_8169));
NAND2X1 g129197(.A (n_13893), .B (n_33225), .Y (n_32255));
NOR2X1 g129201(.A (n_3399), .B (n_7639), .Y (n_8166));
NAND2X1 g129239(.A (n_8164), .B (n_8163), .Y (n_8165));
NAND2X1 g128010(.A (n_7753), .B (n_7512), .Y (n_8979));
NAND2X1 g129338(.A (P2_reg2[18] ), .B (n_33225), .Y (n_8162));
NAND2X1 g129348(.A (n_10043), .B (n_7864), .Y (n_8158));
NAND2X1 g129351(.A (n_10041), .B (n_8163), .Y (n_8157));
NOR2X1 g129355(.A (n_341), .B (n_7807), .Y (n_8156));
NAND3X1 g129400(.A (n_7022), .B (n_8154), .C (n_8153), .Y (n_8155));
NAND3X1 g129415(.A (n_7133), .B (n_8151), .C (n_8150), .Y (n_8152));
NAND4X1 g129445(.A (n_8032), .B (n_8148), .C (n_8147), .D (n_8146),.Y (n_8149));
NAND4X1 g129446(.A (n_8034), .B (n_8144), .C (n_8143), .D (n_8142),.Y (n_8145));
NAND4X1 g129453(.A (n_8014), .B (n_8140), .C (n_8139), .D (n_8138),.Y (n_8141));
NAND4X1 g129462(.A (n_8121), .B (n_8136), .C (n_8135), .D (n_8134),.Y (n_8137));
NAND4X1 g129482(.A (n_8131), .B (n_8130), .C (n_8129), .D (n_8128),.Y (n_8132));
INVX4 g129554(.A (n_8293), .Y (n_15850));
INVX2 g129745(.A (n_8445), .Y (n_8125));
CLKBUFX1 g126134(.A (n_34693), .Y (n_30563));
INVX1 g129831(.A (n_33094), .Y (n_8124));
INVX1 g129833(.A (n_33094), .Y (n_13409));
AND2X1 g129839(.A (n_7614), .B (n_8121), .Y (n_8122));
AOI22X1 g129848(.A0 (n_4478), .A1 (n_8114), .B0 (n_8113), .B1(n_8117), .Y (n_8119));
AOI22X1 g129849(.A0 (n_8115), .A1 (n_8114), .B0 (n_8113), .B1(addr_431), .Y (n_8116));
AOI22X1 g129853(.A0 (n_6204), .A1 (n_8114), .B0 (n_8113), .B1(addr_442), .Y (n_8112));
AOI22X1 g129854(.A0 (n_3959), .A1 (n_8114), .B0 (n_8113), .B1(addr_433), .Y (n_8109));
AOI22X1 g129856(.A0 (n_8105), .A1 (n_8114), .B0 (n_8113), .B1(addr_441), .Y (n_8106));
NAND2X1 g127968(.A (n_13301), .B (n_8245), .Y (n_8103));
AOI22X1 g129857(.A0 (n_35368), .A1 (n_8114), .B0 (n_8113), .B1(addr_430), .Y (n_8102));
AOI22X1 g129859(.A0 (n_3870), .A1 (n_8114), .B0 (n_8113), .B1(addr_432), .Y (n_8099));
AOI22X1 g129860(.A0 (n_33034), .A1 (n_8114), .B0 (n_8113), .B1(addr_437), .Y (n_8096));
AOI22X1 g129861(.A0 (n_4825), .A1 (n_8114), .B0 (n_8113), .B1(addr_438), .Y (n_8093));
NAND2X2 g127966(.A (n_7361), .B (n_7715), .Y (n_8526));
AOI22X1 g129863(.A0 (n_3845), .A1 (n_8114), .B0 (n_8113), .B1(addr_436), .Y (n_8090));
INVX2 g128138(.A (n_8086), .Y (n_8518));
NOR2X1 g129353(.A (n_3198), .B (n_7998), .Y (n_8085));
NAND2X1 g129913(.A (n_7616), .B (n_8083), .Y (n_8084));
NAND2X1 g129918(.A (n_7616), .B (n_481), .Y (n_8082));
NAND2X1 g129931(.A (n_7616), .B (n_8079), .Y (n_8080));
NAND2X1 g129933(.A (n_7616), .B (addr_447), .Y (n_8078));
NAND2X1 g129936(.A (n_7616), .B (n_8074), .Y (n_8075));
INVX1 g128827(.A (n_8393), .Y (n_8400));
INVX2 g128460(.A (n_33125), .Y (n_31878));
INVX1 g130032(.A (n_10676), .Y (n_8399));
INVX1 g128812(.A (n_8393), .Y (n_8534));
INVX1 g128449(.A (n_33125), .Y (n_31689));
INVX1 g126103(.A (n_8319), .Y (n_28485));
CLKBUFX1 g128799(.A (n_8393), .Y (n_8844));
INVX1 g128433(.A (n_33125), .Y (n_24695));
INVX1 g128769(.A (n_8393), .Y (n_9813));
CLKBUFX1 g128770(.A (n_8393), .Y (n_9413));
INVX1 g127902(.A (n_31360), .Y (n_30380));
INVX1 g127897(.A (n_31041), .Y (n_31174));
INVX1 g127888(.A (n_31233), .Y (n_31240));
NOR2X1 g129170(.A (P2_reg1[26] ), .B (n_8168), .Y (n_8066));
INVX8 g128712(.A (n_8884), .Y (n_8484));
NOR2X1 g128976(.A (n_7673), .B (n_7570), .Y (n_35444));
INVX1 g125967(.A (n_11138), .Y (n_9520));
NAND3X1 g125933(.A (n_7165), .B (n_8060), .C (n_7794), .Y (n_8692));
NAND3X1 g125921(.A (n_7165), .B (n_8060), .C (n_7396), .Y (n_8677));
INVX4 g125857(.A (n_8007), .Y (n_8678));
INVX1 g128654(.A (n_35008), .Y (n_31236));
NOR2X1 g128508(.A (n_7967), .B (n_7692), .Y (n_10034));
INVX1 g127765(.A (n_8058), .Y (n_8059));
AOI21X1 g129065(.A0 (n_8055), .A1 (n_8197), .B0 (n_7676), .Y(n_8056));
AOI21X1 g129020(.A0 (n_10182), .A1 (n_7722), .B0 (n_7567), .Y(n_8054));
NAND2X1 g129350(.A (n_10047), .B (n_33225), .Y (n_8052));
NAND2X2 g127720(.A (n_7767), .B (n_7535), .Y (n_16096));
NAND4X1 g129449(.A (n_8050), .B (n_8049), .C (n_8048), .D (n_8047),.Y (n_8051));
INVX1 g127915(.A (n_8070), .Y (n_8528));
INVX1 g127887(.A (n_31233), .Y (n_30569));
NAND2X2 g129436(.A (n_7403), .B (n_7553), .Y (n_8039));
NOR2X1 g126518(.A (n_7762), .B (n_8304), .Y (n_8643));
INVX1 g126496(.A (n_8036), .Y (n_8037));
INVX1 g129829(.A (n_33094), .Y (n_13416));
AND2X1 g129816(.A (n_7615), .B (n_8034), .Y (n_8035));
INVX1 g129835(.A (n_33094), .Y (n_13075));
AND2X1 g129838(.A (n_7610), .B (n_8032), .Y (n_8033));
INVX1 g127100(.A (n_8286), .Y (n_27798));
AOI22X1 g129862(.A0 (n_4731), .A1 (n_8114), .B0 (n_8113), .B1(addr_439), .Y (n_8031));
INVX1 g126414(.A (n_33713), .Y (n_15147));
NAND2X1 g127498(.A (n_10211), .B (n_8245), .Y (n_8029));
INVX1 g126396(.A (n_33713), .Y (n_15413));
AOI21X1 g129098(.A0 (n_10134), .A1 (n_8177), .B0 (n_7593), .Y(n_32563));
INVX1 g128450(.A (n_33125), .Y (n_31555));
AOI22X1 g129858(.A0 (n_4535), .A1 (n_8114), .B0 (n_8113), .B1(addr_434), .Y (n_8027));
AND2X1 g127437(.A (n_4824), .B (n_8245), .Y (n_8024));
NAND2X1 g127428(.A (n_4590), .B (n_8245), .Y (n_8023));
NAND2X1 g127419(.A (n_4477), .B (n_8245), .Y (n_8022));
INVX1 g128438(.A (n_33125), .Y (n_26002));
AOI22X1 g129855(.A0 (n_4010), .A1 (n_8114), .B0 (n_8113), .B1(addr_435), .Y (n_8020));
INVX1 g128432(.A (n_33125), .Y (n_29633));
NOR2X1 g129417(.A (n_3453), .B (n_7637), .Y (n_8016));
AND2X1 g129795(.A (n_7618), .B (n_8014), .Y (n_8015));
NOR4X1 g125435(.A (n_113), .B (n_7024), .C (n_7527), .D (n_7346), .Y(n_8013));
NOR2X1 g125463(.A (n_7573), .B (n_34693), .Y (n_8010));
NOR2X1 g125570(.A (n_8003), .B (n_8009), .Y (n_8375));
NAND4X1 g125582(.A (n_7531), .B (n_7398), .C (n_8008), .D (n_7155),.Y (n_32343));
NOR2X1 g125858(.A (n_7386), .B (n_6833), .Y (n_8007));
BUFX3 g125975(.A (n_8005), .Y (n_11138));
INVX1 g125977(.A (n_8005), .Y (n_8004));
INVX1 g125999(.A (n_8003), .Y (n_8325));
NAND2X1 g129372(.A (n_8001), .B (n_7401), .Y (n_8002));
AOI21X1 g129029(.A0 (n_9590), .A1 (n_7953), .B0 (n_7375), .Y(n_8000));
INVX1 g126157(.A (n_33991), .Y (n_7997));
NAND2X1 g126202(.A (n_7994), .B (n_7993), .Y (n_10067));
AND2X1 g126203(.A (n_7166), .B (n_7763), .Y (n_10196));
INVX1 g126262(.A (n_8009), .Y (n_8314));
INVX4 g126319(.A (n_7992), .Y (n_8313));
NAND2X1 g126497(.A (n_7993), .B (n_7986), .Y (n_8036));
NAND2X1 g126519(.A (n_7987), .B (n_7986), .Y (n_8679));
INVX1 g126520(.A (n_18218), .Y (n_7985));
NAND2X1 g129346(.A (P2_reg_107), .B (n_7983), .Y (n_7984));
INVX1 g127098(.A (n_30063), .Y (n_29150));
INVX1 g127102(.A (n_30063), .Y (n_8286));
AND2X1 g127050(.A (n_7394), .B (n_7558), .Y (n_7981));
INVX1 g127139(.A (n_8333), .Y (n_8284));
AND2X1 g127142(.A (n_29944), .B (n_7393), .Y (n_8283));
NOR2X1 g129317(.A (n_352), .B (n_7917), .Y (n_7978));
NAND4X1 g127385(.A (n_35454), .B (n_7195), .C (n_7031), .D (n_6834),.Y (n_8277));
NAND2X1 g127415(.A (n_7967), .B (n_7691), .Y (n_10253));
AND2X1 g127691(.A (n_7526), .B (n_7976), .Y (n_7977));
NOR2X1 g127766(.A (n_1054), .B (n_7975), .Y (n_8058));
INVX1 g127873(.A (n_7603), .Y (n_31398));
NAND2X2 g128132(.A (n_35613), .B (n_35612), .Y (n_8231));
NAND2X2 g128139(.A (n_32049), .B (n_32050), .Y (n_8086));
INVX4 g128725(.A (n_7970), .Y (n_9373));
OR2X1 g128372(.A (n_7520), .B (n_7530), .Y (n_7973));
OR2X1 g128373(.A (n_65), .B (n_7521), .Y (n_7972));
INVX1 g129669(.A (n_12690), .Y (n_13408));
OR2X1 g128609(.A (n_7188), .B (n_7517), .Y (n_7971));
INVX8 g128715(.A (n_7970), .Y (n_8884));
INVX1 g128901(.A (n_8557), .Y (n_8575));
NAND2X1 g127447(.A (n_7805), .B (n_7967), .Y (n_11191));
NAND2X1 g129929(.A (n_7616), .B (addr_450), .Y (n_7966));
AOI22X1 g129503(.A0 (n_6335), .A1 (n_7653), .B0 (n_6299), .B1(n_33068), .Y (n_7964));
INVX1 g128944(.A (n_8387), .Y (n_7963));
NOR2X1 g128964(.A (n_7313), .B (n_7562), .Y (n_7962));
NOR2X1 g128967(.A (n_7485), .B (n_7483), .Y (n_7961));
NOR2X1 g128969(.A (n_7140), .B (n_7370), .Y (n_7960));
AOI21X1 g128987(.A0 (n_2911), .A1 (n_7956), .B0 (n_7462), .Y(n_7959));
AOI21X1 g129002(.A0 (n_7957), .A1 (n_7956), .B0 (n_7374), .Y(n_7958));
AOI21X1 g129017(.A0 (n_7939), .A1 (n_9121), .B0 (n_7501), .Y(n_7955));
AOI21X1 g129022(.A0 (P2_reg1[4] ), .A1 (n_7953), .B0 (n_7480), .Y(n_7954));
NOR2X1 g129041(.A (n_7206), .B (n_7499), .Y (n_7952));
NOR2X1 g129043(.A (n_7359), .B (n_7461), .Y (n_35925));
AOI21X1 g129047(.A0 (P3_reg2[13] ), .A1 (n_8183), .B0 (n_7460), .Y(n_7949));
AOI21X1 g129048(.A0 (n_13327), .A1 (n_7754), .B0 (n_7544), .Y(n_35439));
AOI21X1 g129049(.A0 (n_13213), .A1 (n_7716), .B0 (n_7498), .Y(n_35438));
AOI21X1 g129062(.A0 (P3_reg1[18] ), .A1 (n_7944), .B0 (n_7490), .Y(n_7945));
AOI21X1 g129063(.A0 (n_13724), .A1 (n_7944), .B0 (n_7372), .Y(n_7943));
AOI21X1 g129067(.A0 (n_13673), .A1 (n_7503), .B0 (n_7470), .Y(n_7942));
AOI21X1 g129083(.A0 (n_7939), .A1 (n_9595), .B0 (n_7408), .Y(n_7940));
AOI21X1 g129084(.A0 (P2_reg1[6] ), .A1 (n_7935), .B0 (n_7493), .Y(n_7938));
AOI21X1 g129085(.A0 (n_10363), .A1 (n_7307), .B0 (n_7479), .Y(n_7937));
AOI21X1 g129086(.A0 (P2_reg1[12] ), .A1 (n_7935), .B0 (n_7494), .Y(n_7936));
AOI21X1 g129095(.A0 (P2_reg1[5] ), .A1 (n_7935), .B0 (n_7478), .Y(n_7934));
AOI21X1 g129102(.A0 (n_10563), .A1 (n_7380), .B0 (n_7467), .Y(n_7933));
NAND2X1 g129113(.A (n_7500), .B (n_7236), .Y (n_7932));
NAND2X1 g129141(.A (P2_reg1[18] ), .B (n_7930), .Y (n_7929));
NAND2X1 g129152(.A (P2_reg1[23] ), .B (n_9692), .Y (n_7928));
NAND2X1 g129154(.A (P1_reg1[30] ), .B (n_7926), .Y (n_7927));
NAND2X1 g129157(.A (n_10247), .B (n_7926), .Y (n_7925));
NOR2X1 g129172(.A (n_358), .B (n_7823), .Y (n_7924));
NAND2X1 g129173(.A (P2_reg1[20] ), .B (n_7930), .Y (n_7923));
NAND2X1 g129180(.A (P2_reg1[31] ), .B (n_7255), .Y (n_32254));
NAND2X1 g129189(.A (n_10169), .B (n_7926), .Y (n_7921));
NAND2X1 g129193(.A (n_13169), .B (n_8209), .Y (n_7920));
NAND2X1 g129206(.A (n_3184), .B (n_8209), .Y (n_7919));
NOR2X1 g129221(.A (n_235), .B (n_7917), .Y (n_7918));
NOR2X1 g129907(.A (n_3483), .B (n_7432), .Y (n_7916));
NOR2X1 g129234(.A (n_382), .B (n_7445), .Y (n_7915));
NAND2X1 g129260(.A (n_13301), .B (n_8209), .Y (n_7914));
NAND2X1 g129289(.A (P2_reg_106), .B (n_7983), .Y (n_7912));
NOR2X1 g129311(.A (n_273), .B (n_33228), .Y (n_7911));
NOR2X1 g129336(.A (n_3160), .B (n_7798), .Y (n_7910));
NOR2X1 g129380(.A (n_70), .B (n_33228), .Y (n_7909));
NAND4X1 g129451(.A (n_7906), .B (n_7905), .C (n_7904), .D (n_7903),.Y (n_7907));
NAND4X1 g129452(.A (n_7901), .B (n_7900), .C (n_34977), .D (n_7898),.Y (n_7902));
NAND4X1 g129455(.A (n_7896), .B (n_7895), .C (n_7894), .D (n_7893),.Y (n_7897));
NAND4X1 g129456(.A (n_7891), .B (n_7890), .C (n_34578), .D (n_7888),.Y (n_7892));
NAND4X1 g129461(.A (n_7886), .B (n_7885), .C (n_7884), .D (n_7883),.Y (n_7887));
NAND4X1 g129463(.A (n_7881), .B (n_7880), .C (n_7879), .D (n_7878),.Y (n_7882));
AOI22X1 g129481(.A0 (n_5713), .A1 (n_33068), .B0 (n_5873), .B1(n_7653), .Y (n_7877));
AOI22X1 g129485(.A0 (n_6277), .A1 (n_33068), .B0 (n_6279), .B1(n_7653), .Y (n_7876));
AOI22X1 g129488(.A0 (n_5394), .A1 (n_33068), .B0 (n_5456), .B1(n_7653), .Y (n_7873));
AOI22X1 g129499(.A0 (n_6399), .A1 (n_33068), .B0 (n_6377), .B1(n_7653), .Y (n_7870));
NAND2X1 g129900(.A (n_7616), .B (addr_451), .Y (n_7869));
INVX2 g129556(.A (n_15704), .Y (n_8293));
NAND2X2 g127982(.A (n_7539), .B (n_7238), .Y (n_8233));
NAND3X1 g129821(.A (n_7432), .B (n_7209), .C (n_6959), .Y (n_7862));
AOI21X1 g129844(.A0 (n_8113), .A1 (n_482), .B0 (n_7431), .Y (n_7859));
INVX1 g128848(.A (n_7860), .Y (n_8598));
AOI22X1 g129851(.A0 (n_2807), .A1 (n_8114), .B0 (n_8113), .B1(addr_424), .Y (n_7858));
AOI22X1 g129852(.A0 (n_3472), .A1 (n_8114), .B0 (n_8113), .B1(addr_426), .Y (n_7856));
NAND4X1 g129460(.A (n_7851), .B (n_7850), .C (n_7849), .D (n_7848),.Y (n_7852));
AOI22X1 g129490(.A0 (n_6063), .A1 (n_7653), .B0 (n_6095), .B1(n_33068), .Y (n_7847));
NOR2X1 g129895(.A (n_2962), .B (n_7432), .Y (n_7845));
INVX1 g129711(.A (n_7998), .Y (n_8442));
NAND2X1 g129909(.A (n_7616), .B (n_7843), .Y (n_7844));
NAND2X1 g129912(.A (n_7616), .B (n_7841), .Y (n_7842));
NAND2X1 g129917(.A (n_7616), .B (n_7839), .Y (n_7840));
NAND2X1 g129924(.A (n_7616), .B (addr_452), .Y (n_7838));
NAND2X1 g129925(.A (n_7616), .B (addr_453), .Y (n_7836));
NAND2X1 g129930(.A (n_7616), .B (n_7833), .Y (n_7834));
INVX1 g129971(.A (n_13555), .Y (n_7832));
INVX1 g129981(.A (n_7613), .Y (n_13413));
INVX1 g126115(.A (n_34693), .Y (n_8319));
INVX8 g128797(.A (n_9310), .Y (n_8393));
NAND2X1 g129191(.A (P2_reg1[22] ), .B (n_9692), .Y (n_7830));
AOI22X1 g129486(.A0 (n_6455), .A1 (n_33068), .B0 (n_6395), .B1(n_7653), .Y (n_7829));
NAND2X1 g129187(.A (P2_reg1[27] ), .B (n_9692), .Y (n_7828));
INVX1 g127916(.A (n_7827), .Y (n_8070));
INVX1 g127898(.A (n_31628), .Y (n_31041));
INVX1 g126679(.A (n_8065), .Y (n_25228));
INVX1 g126665(.A (n_8065), .Y (n_25111));
NAND2X1 g126789(.A (n_7532), .B (P1_d_98), .Y (n_7822));
INVX1 g130033(.A (n_7821), .Y (n_10676));
AOI21X1 g129013(.A0 (n_7819), .A1 (n_7956), .B0 (n_7472), .Y(n_7820));
NAND4X1 g127818(.A (n_7491), .B (n_7202), .C (n_7148), .D (n_7005),.Y (n_32334));
AOI21X1 g129066(.A0 (n_13687), .A1 (n_7503), .B0 (n_7468), .Y(n_35445));
NAND4X1 g129458(.A (n_7815), .B (n_7814), .C (n_7813), .D (n_7812),.Y (n_7816));
NAND2X1 g129136(.A (P1_reg1[24] ), .B (n_7926), .Y (n_7811));
NAND2X2 g128125(.A (n_7193), .B (n_7509), .Y (n_7810));
AOI21X1 g129060(.A0 (n_13699), .A1 (n_7944), .B0 (n_7489), .Y(n_7809));
AOI21X1 g129039(.A0 (n_7348), .A1 (P3_reg2[9] ), .B0 (n_7482), .Y(n_35337));
INVX2 g129747(.A (n_7807), .Y (n_8445));
NAND2X1 g128580(.A (P2_d), .B (n_7805), .Y (n_7806));
AOI21X1 g129061(.A0 (n_10144), .A1 (n_7722), .B0 (n_7540), .Y(n_7804));
NAND2X2 g128581(.A (n_7805), .B (P2_B), .Y (n_10251));
INVX4 g127082(.A (n_7764), .Y (n_8927));
INVX4 g126662(.A (n_8065), .Y (n_8303));
INVX1 g127886(.A (n_31573), .Y (n_31233));
INVX1 g127875(.A (n_7603), .Y (n_30403));
INVX1 g129673(.A (n_12690), .Y (n_13106));
NOR2X1 g129361(.A (n_2910), .B (n_7798), .Y (n_7799));
INVX1 g128857(.A (n_8245), .Y (n_8552));
NAND2X1 g126582(.A (n_7994), .B (n_7987), .Y (n_8305));
INVX1 g128309(.A (n_7796), .Y (n_7797));
NAND2X1 g126470(.A (n_7773), .B (n_7794), .Y (n_8306));
INVX1 g127112(.A (n_30063), .Y (n_8285));
AOI21X1 g129036(.A0 (P3_reg1[26] ), .A1 (n_7503), .B0 (n_7404), .Y(n_7791));
AOI21X1 g128984(.A0 (n_7183), .A1 (P1_reg2[9] ), .B0 (n_7488), .Y(n_7789));
INVX1 g127573(.A (n_7787), .Y (n_7788));
AOI21X1 g128985(.A0 (n_1911), .A1 (n_7476), .B0 (n_7474), .Y(n_7786));
INVX4 g127034(.A (n_8322), .Y (n_26213));
AOI21X1 g129843(.A0 (n_8113), .A1 (addr_425), .B0 (n_7433), .Y(n_7785));
INVX1 g129624(.A (n_7863), .Y (n_10671));
AOI21X1 g129045(.A0 (P3_reg2[10] ), .A1 (n_7714), .B0 (n_7378), .Y(n_7783));
NOR2X1 g129374(.A (n_271), .B (n_7571), .Y (n_7781));
AOI21X1 g129032(.A0 (n_10197), .A1 (n_7722), .B0 (n_7257), .Y(n_7779));
INVX4 g126200(.A (n_8316), .Y (n_29725));
NOR2X1 g126243(.A (n_6387), .B (n_7777), .Y (n_7778));
INVX1 g126244(.A (n_7775), .Y (n_7776));
NOR2X1 g126263(.A (n_7379), .B (n_7774), .Y (n_8009));
AND2X1 g126424(.A (n_8060), .B (n_7771), .Y (n_7772));
NOR2X1 g126521(.A (n_7383), .B (n_7770), .Y (n_18218));
INVX2 g129653(.A (n_9692), .Y (n_8168));
INVX1 g129972(.A (n_7769), .Y (n_13555));
AOI21X1 g129006(.A0 (n_10221), .A1 (n_7722), .B0 (n_7323), .Y(n_7767));
AOI21X1 g128998(.A0 (n_13680), .A1 (n_7503), .B0 (n_7241), .Y(n_7766));
NOR2X1 g127083(.A (n_7335), .B (n_7173), .Y (n_7764));
INVX1 g127181(.A (n_7993), .Y (n_7762));
NAND3X1 g128945(.A (n_7736), .B (n_7760), .C (n_7761), .Y (n_8387));
INVX1 g127286(.A (n_7987), .Y (n_7759));
INVX1 g127314(.A (n_7794), .Y (n_7758));
AOI21X1 g128968(.A0 (n_7755), .A1 (n_7754), .B0 (n_7242), .Y(n_7756));
NOR2X1 g128963(.A (n_7338), .B (n_7314), .Y (n_7753));
AOI21X1 g127407(.A0 (n_6495), .A1 (n_7393), .B0 (n_7528), .Y(n_7752));
NOR2X1 g129298(.A (n_228), .B (n_7672), .Y (n_7750));
NAND2X1 g127569(.A (n_1054), .B (n_7748), .Y (n_10989));
OR2X1 g127574(.A (n_7541), .B (n_7333), .Y (n_7787));
NAND2X1 g127736(.A (P3_B), .B (n_7748), .Y (n_7749));
NAND2X1 g129932(.A (n_8114), .B (n_7747), .Y (n_8452));
INVX1 g127917(.A (n_7603), .Y (n_7827));
INVX1 g128219(.A (n_7745), .Y (n_7746));
AND2X1 g128310(.A (n_7405), .B (n_7522), .Y (n_7796));
INVX1 g128374(.A (n_7743), .Y (n_7744));
NOR2X1 g128658(.A (n_7331), .B (n_7525), .Y (n_8996));
NAND2X1 g129252(.A (P2_reg2[11] ), .B (n_33225), .Y (n_7741));
NOR2X1 g129281(.A (n_10110), .B (n_7685), .Y (n_7740));
AOI21X1 g128957(.A0 (n_2138), .A1 (n_7705), .B0 (n_7160), .Y(n_7739));
AOI21X1 g128958(.A0 (n_7737), .A1 (n_7736), .B0 (n_7050), .Y(n_7738));
AOI21X1 g128975(.A0 (n_7734), .A1 (n_7538), .B0 (n_7315), .Y(n_7735));
NOR2X1 g129008(.A (n_7057), .B (n_7322), .Y (n_7733));
AOI21X1 g129009(.A0 (n_10138), .A1 (n_7722), .B0 (n_7231), .Y(n_7732));
AOI21X1 g129014(.A0 (n_7730), .A1 (n_7736), .B0 (n_7186), .Y(n_7731));
AOI21X1 g129016(.A0 (n_10191), .A1 (n_7722), .B0 (n_7252), .Y(n_35616));
AOI21X1 g129024(.A0 (n_10150), .A1 (n_7722), .B0 (n_7194), .Y(n_7728));
AOI21X1 g129027(.A0 (n_7722), .A1 (n_10154), .B0 (n_7320), .Y(n_7727));
AOI21X1 g129028(.A0 (n_7736), .A1 (n_7724), .B0 (n_7182), .Y(n_7725));
AOI21X1 g129033(.A0 (n_10140), .A1 (n_7722), .B0 (n_7198), .Y(n_7723));
AOI21X1 g129037(.A0 (n_13698), .A1 (n_7503), .B0 (n_7302), .Y(n_7721));
AOI21X1 g129038(.A0 (n_13695), .A1 (n_7584), .B0 (n_7309), .Y(n_7720));
NAND2X1 g127435(.A (n_1054), .B (n_7422), .Y (n_7719));
AOI21X1 g129046(.A0 (n_13204), .A1 (n_7716), .B0 (n_7233), .Y(n_7717));
AOI21X1 g129051(.A0 (P3_reg2[6] ), .A1 (n_7714), .B0 (n_7311), .Y(n_7715));
AOI21X1 g129087(.A0 (P2_reg2[2] ), .A1 (n_33225), .B0 (n_7208), .Y(n_7713));
AOI21X1 g129089(.A0 (n_10205), .A1 (n_7722), .B0 (n_7240), .Y(n_7712));
AND2X1 g129090(.A (n_7318), .B (n_7308), .Y (n_7711));
INVX1 g129105(.A (n_7505), .Y (n_32892));
AOI21X1 g129112(.A0 (n_7706), .A1 (n_7705), .B0 (n_7149), .Y(n_35617));
NOR2X1 g129135(.A (P1_reg1[25] ), .B (n_7702), .Y (n_7704));
NOR2X1 g129139(.A (n_122), .B (n_7702), .Y (n_7703));
NOR2X1 g129149(.A (n_322), .B (n_7443), .Y (n_7701));
NAND2X1 g129165(.A (P3_reg1[17] ), .B (n_7503), .Y (n_7700));
NOR2X1 g129166(.A (n_201), .B (n_7702), .Y (n_7699));
NOR2X1 g129171(.A (n_361), .B (n_7607), .Y (n_7698));
NOR2X1 g129175(.A (n_41), .B (n_7595), .Y (n_7697));
NOR2X1 g129182(.A (n_182), .B (n_7607), .Y (n_7696));
NAND2X1 g129204(.A (n_10858), .B (n_7694), .Y (n_7695));
NAND2X1 g129207(.A (n_11144), .B (n_8485), .Y (n_7693));
INVX1 g128917(.A (n_7691), .Y (n_7692));
NAND2X1 g129216(.A (P2_reg2[10] ), .B (n_33225), .Y (n_7689));
NOR2X1 g129217(.A (n_103), .B (n_7662), .Y (n_7687));
NOR2X1 g129235(.A (n_3037), .B (n_7685), .Y (n_7686));
NOR2X1 g129238(.A (n_311), .B (n_7662), .Y (n_7684));
NOR2X1 g129280(.A (n_333), .B (n_7680), .Y (n_7683));
NOR2X1 g129282(.A (n_10103), .B (n_7685), .Y (n_7682));
NOR2X1 g129299(.A (n_338), .B (n_7680), .Y (n_7681));
NOR2X1 g129300(.A (n_10114), .B (n_7669), .Y (n_7679));
NOR2X1 g129301(.A (n_3493), .B (n_7214), .Y (n_7678));
NOR2X1 g129302(.A (n_5289), .B (n_7680), .Y (n_7677));
NOR2X1 g129303(.A (n_115), .B (n_7349), .Y (n_7676));
NAND2X1 g129305(.A (n_13216), .B (n_7034), .Y (n_7675));
NAND2X1 g129306(.A (n_14133), .B (n_8335), .Y (n_7674));
NOR2X1 g129307(.A (n_387), .B (n_7672), .Y (n_7673));
NOR2X1 g129309(.A (n_304), .B (n_7672), .Y (n_7671));
NOR2X1 g129310(.A (n_10116), .B (n_7669), .Y (n_7670));
NAND2X1 g129339(.A (n_9165), .B (n_8335), .Y (n_7668));
NAND2X1 g129352(.A (P2_reg_104), .B (n_8335), .Y (n_7666));
NAND2X1 g129364(.A (n_7664), .B (n_8192), .Y (n_7665));
NOR2X1 g129365(.A (n_49), .B (n_7662), .Y (n_7663));
NAND2X1 g129366(.A (P1_reg2[30] ), .B (n_8485), .Y (n_7661));
NOR2X1 g129370(.A (n_15), .B (n_7662), .Y (n_7660));
NOR2X1 g129413(.A (n_83), .B (n_7136), .Y (n_7659));
NAND2X1 g129428(.A (n_10617), .B (n_7657), .Y (n_7658));
NOR2X1 g129444(.A (n_3124), .B (n_7442), .Y (n_7656));
INVX1 g128902(.A (n_8245), .Y (n_8557));
AOI22X1 g129478(.A0 (n_6227), .A1 (n_33068), .B0 (n_6239), .B1(n_7653), .Y (n_7655));
AOI22X1 g129484(.A0 (n_6103), .A1 (n_33068), .B0 (n_6151), .B1(n_7653), .Y (n_7654));
AOI22X1 g129494(.A0 (n_5771), .A1 (n_33068), .B0 (n_5690), .B1(n_7653), .Y (n_7651));
INVX1 g128885(.A (n_8245), .Y (n_7871));
AOI22X1 g129495(.A0 (n_5868), .A1 (n_7653), .B0 (n_5871), .B1(n_33068), .Y (n_7649));
AOI22X1 g129496(.A0 (n_6185), .A1 (n_7653), .B0 (n_6165), .B1(n_33068), .Y (n_7648));
AOI22X1 g129497(.A0 (n_5666), .A1 (n_7653), .B0 (n_5648), .B1(n_33068), .Y (n_7647));
AOI21X1 g129011(.A0 (n_10148), .A1 (n_7722), .B0 (n_7321), .Y(n_7646));
AND2X1 g129548(.A (n_7653), .B (n_1054), .Y (n_7644));
INVX2 g129612(.A (n_7917), .Y (n_7864));
INVX1 g129626(.A (n_7641), .Y (n_7863));
INVX1 g129674(.A (n_7640), .Y (n_12690));
INVX2 g129718(.A (n_7798), .Y (n_8163));
INVX1 g129729(.A (n_7638), .Y (n_7639));
INVX1 g129730(.A (n_7638), .Y (n_7637));
INVX2 g129748(.A (n_7983), .Y (n_7807));
NOR2X1 g129775(.A (n_4345), .B (n_7597), .Y (n_7636));
NOR2X1 g129776(.A (n_32388), .B (n_33906), .Y (n_7635));
AOI21X1 g129865(.A0 (n_6452), .A1 (n_6856), .B0 (n_7272), .Y(n_7634));
AOI21X1 g129866(.A0 (n_6315), .A1 (n_6856), .B0 (n_7224), .Y(n_7633));
AOI21X1 g129867(.A0 (n_6234), .A1 (n_6856), .B0 (n_7219), .Y(n_7631));
AOI21X1 g129872(.A0 (n_5533), .A1 (n_6856), .B0 (n_7278), .Y(n_7630));
AOI21X1 g129874(.A0 (n_5534), .A1 (n_6856), .B0 (n_7276), .Y(n_7629));
AOI21X1 g129875(.A0 (n_6068), .A1 (n_6856), .B0 (n_7273), .Y(n_7628));
AOI21X1 g129876(.A0 (n_5920), .A1 (n_6856), .B0 (n_7351), .Y(n_7626));
AOI21X1 g129878(.A0 (n_6173), .A1 (n_6856), .B0 (n_7275), .Y(n_7625));
AOI21X1 g129879(.A0 (n_6238), .A1 (n_6856), .B0 (n_7269), .Y(n_7624));
AOI21X1 g129880(.A0 (n_5992), .A1 (n_6856), .B0 (n_7266), .Y(n_7623));
AOI21X1 g129881(.A0 (n_6120), .A1 (n_6856), .B0 (n_7268), .Y(n_7622));
INVX8 g128836(.A (n_7620), .Y (n_9310));
AOI21X1 g129884(.A0 (n_6519), .A1 (n_6856), .B0 (n_7352), .Y(n_7619));
NAND2X1 g129893(.A (n_7616), .B (addr_446), .Y (n_7618));
NAND2X1 g129904(.A (n_7616), .B (addr_2), .Y (n_7617));
NAND2X1 g129914(.A (n_7616), .B (n_10057), .Y (n_7615));
NAND2X1 g129935(.A (n_7616), .B (n_130), .Y (n_7614));
INVX1 g129968(.A (n_13296), .Y (n_13540));
INVX1 g129986(.A (n_33290), .Y (n_7613));
AOI22X1 g129491(.A0 (n_5400), .A1 (n_33068), .B0 (n_5297), .B1(n_7653), .Y (n_7612));
INVX1 g130034(.A (n_15725), .Y (n_7821));
NAND2X1 g129896(.A (n_7616), .B (n_233), .Y (n_7610));
INVX1 g130098(.A (n_8432), .Y (n_7609));
BUFX3 g130116(.A (n_7793), .Y (n_9676));
NOR2X1 g129185(.A (n_4045), .B (n_7607), .Y (n_7608));
NOR2X1 g129186(.A (n_279), .B (n_7607), .Y (n_7606));
INVX1 g129973(.A (n_7769), .Y (n_12954));
AND2X1 g130598(.A (n_1332), .B (n_7244), .Y (n_7604));
INVX1 g127899(.A (n_7603), .Y (n_31628));
INVX1 g127892(.A (n_7603), .Y (n_31573));
AOI22X1 g129483(.A0 (n_6094), .A1 (n_7653), .B0 (n_6067), .B1(n_33068), .Y (n_7602));
AND2X1 g126000(.A (n_7345), .B (n_6878), .Y (n_8003));
AND2X1 g125978(.A (n_7347), .B (n_7165), .Y (n_8005));
NOR2X1 g129774(.A (n_4772), .B (n_7597), .Y (n_7598));
CLKBUFX1 g129627(.A (n_7641), .Y (n_10696));
NOR2X1 g129158(.A (n_66), .B (n_7595), .Y (n_7596));
NOR2X1 g129155(.A (n_75), .B (n_7443), .Y (n_7594));
NOR2X1 g129143(.A (P1_reg1[26] ), .B (n_7702), .Y (n_7593));
NOR2X1 g129291(.A (n_2817), .B (n_7685), .Y (n_7592));
AOI21X1 g129882(.A0 (n_6280), .A1 (n_6856), .B0 (n_7225), .Y(n_7591));
NAND2X1 g127035(.A (n_7337), .B (n_7552), .Y (n_8322));
NOR2X1 g129362(.A (n_2693), .B (n_7998), .Y (n_7590));
AOI21X1 g129040(.A0 (n_7503), .A1 (P3_reg1[9] ), .B0 (n_7013), .Y(n_35338));
INVX4 g126698(.A (n_7587), .Y (n_8065));
AOI21X1 g129877(.A0 (n_6241), .A1 (n_6856), .B0 (n_7354), .Y(n_7586));
AOI21X1 g129042(.A0 (P3_reg1[11] ), .A1 (n_7584), .B0 (n_7212), .Y(n_35926));
INVX1 g128855(.A (n_8245), .Y (n_7860));
NAND2X1 g129392(.A (n_11327), .B (n_7694), .Y (n_7582));
INVX2 g129557(.A (n_7581), .Y (n_15704));
NAND3X1 g127140(.A (n_7232), .B (n_6347), .C (n_7395), .Y (n_8333));
NOR2X1 g129438(.A (n_3101), .B (n_7998), .Y (n_7580));
INVX4 g126444(.A (n_8309), .Y (n_7988));
INVX1 g127113(.A (n_8321), .Y (n_30063));
AOI21X1 g129871(.A0 (n_5397), .A1 (n_6856), .B0 (n_7279), .Y(n_7578));
AOI21X1 g129104(.A0 (P3_reg1[12] ), .A1 (n_7503), .B0 (n_7227), .Y(n_32270));
NAND2X1 g129437(.A (n_7575), .B (n_7956), .Y (n_32128));
NOR2X1 g129304(.A (n_4474), .B (n_7672), .Y (n_7574));
INVX1 g129569(.A (n_15708), .Y (n_7865));
INVX1 g127114(.A (n_8321), .Y (n_7573));
NOR2X1 g129340(.A (n_94), .B (n_7571), .Y (n_7572));
OAI21X1 g129842(.A0 (n_12670), .A1 (n_7432), .B0 (n_7209), .Y(n_14007));
NOR2X1 g129308(.A (n_10119), .B (n_7669), .Y (n_7570));
AOI21X1 g129068(.A0 (n_10201), .A1 (n_7722), .B0 (n_7319), .Y(n_7569));
AOI21X1 g129064(.A0 (P3_reg1[16] ), .A1 (n_7503), .B0 (n_7306), .Y(n_7568));
NOR2X1 g129212(.A (n_3024), .B (n_7290), .Y (n_7567));
NAND2X1 g129404(.A (n_10152), .B (n_8177), .Y (n_7566));
AOI21X1 g129053(.A0 (n_13711), .A1 (n_34590), .B0 (n_7207), .Y(n_7565));
NAND2X1 g129321(.A (n_10219), .B (n_8177), .Y (n_7563));
OR2X1 g126320(.A (n_6974), .B (n_7777), .Y (n_7992));
INVX1 g129970(.A (n_13230), .Y (n_13400));
NOR2X1 g129378(.A (n_3573), .B (n_7481), .Y (n_7562));
NOR2X1 g126245(.A (n_7782), .B (n_7561), .Y (n_7775));
AOI21X1 g129055(.A0 (n_13209), .A1 (n_6836), .B0 (n_7004), .Y(n_32050));
AND2X1 g128610(.A (n_6322), .B (n_7994), .Y (n_7559));
NOR2X1 g127182(.A (n_7558), .B (n_7393), .Y (n_7993));
NOR2X1 g126699(.A (n_7774), .B (n_7561), .Y (n_7587));
INVX1 g129652(.A (n_7556), .Y (n_7823));
INVX1 g129977(.A (n_13230), .Y (n_7555));
NAND3X1 g127115(.A (n_7552), .B (n_7353), .C (n_6975), .Y (n_8321));
NAND3X1 g129324(.A (n_7550), .B (n_7549), .C (n_7457), .Y (n_7551));
NOR2X1 g127316(.A (n_7232), .B (n_6347), .Y (n_7794));
AOI21X1 g128956(.A0 (n_7546), .A1 (n_7534), .B0 (n_7162), .Y(n_7547));
NAND2X1 g129312(.A (P3_reg2[30] ), .B (n_8183), .Y (n_7545));
NOR2X1 g129292(.A (n_205), .B (n_7484), .Y (n_7544));
INVX1 g129969(.A (n_13230), .Y (n_13296));
AND2X1 g127628(.A (n_6435), .B (n_7415), .Y (n_12649));
NAND2X1 g127711(.A (n_7397), .B (n_12670), .Y (n_7543));
NAND2X1 g127712(.A (n_7541), .B (n_7332), .Y (n_32245));
NOR2X1 g129332(.A (n_1004), .B (n_7049), .Y (n_7540));
INVX4 g129629(.A (n_7553), .Y (n_15619));
AOI21X1 g128961(.A0 (n_7538), .A1 (n_2721), .B0 (n_7150), .Y(n_7539));
AOI21X1 g128954(.A0 (n_13167), .A1 (n_7534), .B0 (n_7143), .Y(n_7535));
NOR2X1 g128608(.A (n_6283), .B (n_6974), .Y (n_7533));
INVX1 g128611(.A (n_7531), .Y (n_7532));
NOR2X1 g128659(.A (n_7008), .B (n_7530), .Y (n_8326));
INVX1 g128667(.A (n_7528), .Y (n_29944));
INVX1 g128671(.A (n_7527), .Y (n_27567));
INVX1 g128677(.A (n_7525), .Y (n_7526));
NAND2X1 g128679(.A (n_7523), .B (n_7329), .Y (n_7976));
NAND2X1 g128689(.A (n_7523), .B (n_7200), .Y (n_7524));
NOR2X1 g128837(.A (n_7523), .B (n_7334), .Y (n_7620));
INVX1 g128919(.A (n_7522), .Y (n_7691));
INVX1 g128921(.A (n_7748), .Y (n_7521));
INVX1 g128925(.A (n_7519), .Y (n_7520));
INVX2 g129628(.A (n_7553), .Y (n_7641));
INVX1 g128939(.A (n_7773), .Y (n_7517));
AOI21X1 g128988(.A0 (n_7534), .A1 (n_7515), .B0 (n_7127), .Y(n_7516));
AOI21X1 g129007(.A0 (P3_reg1[4] ), .A1 (n_34586), .B0 (n_7189), .Y(n_7514));
AOI21X1 g129015(.A0 (P2_reg1[2] ), .A1 (n_7255), .B0 (n_7011), .Y(n_7513));
AOI21X1 g129034(.A0 (n_13690), .A1 (n_34586), .B0 (n_7044), .Y(n_7512));
AOI21X1 g129052(.A0 (P3_reg1[7] ), .A1 (n_7584), .B0 (n_7046), .Y(n_7510));
NOR2X1 g129054(.A (n_7014), .B (n_7153), .Y (n_7509));
AOI21X1 g129056(.A0 (n_7376), .A1 (P3_reg3[2] ), .B0 (n_7009), .Y(n_32049));
AOI21X1 g129097(.A0 (n_13692), .A1 (n_7584), .B0 (n_7003), .Y(n_7507));
NAND2X1 g129106(.A (n_7054), .B (n_7163), .Y (n_7505));
NAND2X1 g129134(.A (n_13727), .B (n_7503), .Y (n_7504));
NAND2X1 g129148(.A (P1_reg1[12] ), .B (n_7495), .Y (n_7502));
NOR2X1 g129153(.A (n_7407), .B (n_36), .Y (n_7501));
NAND2X1 g129160(.A (P1_reg1[19] ), .B (n_7355), .Y (n_7500));
NOR2X1 g129161(.A (n_4132), .B (n_7497), .Y (n_7499));
NOR2X1 g129163(.A (n_274), .B (n_7497), .Y (n_7498));
NAND2X1 g129184(.A (P1_reg1[14] ), .B (n_7495), .Y (n_7496));
NOR2X1 g129195(.A (n_96), .B (n_7289), .Y (n_7494));
INVX1 g129975(.A (n_13230), .Y (n_7769));
NOR2X1 g129199(.A (n_101), .B (n_7289), .Y (n_7493));
NOR2X1 g129209(.A (n_372), .B (n_7434), .Y (n_7492));
OR2X1 g129228(.A (n_149), .B (n_7135), .Y (n_7491));
NOR2X1 g129232(.A (n_388), .B (n_7012), .Y (n_7490));
NOR2X1 g129242(.A (n_375), .B (n_7469), .Y (n_7489));
NOR2X1 g129246(.A (n_2563), .B (n_7369), .Y (n_7488));
NOR2X1 g129283(.A (n_318), .B (n_7484), .Y (n_7485));
NOR2X1 g129284(.A (n_10112), .B (n_7459), .Y (n_7483));
NOR2X1 g129286(.A (n_2914), .B (n_7481), .Y (n_7482));
NOR2X1 g129357(.A (n_277), .B (n_7473), .Y (n_7480));
NOR2X1 g129358(.A (n_1058), .B (n_7466), .Y (n_7479));
NOR2X1 g129360(.A (n_295), .B (n_7134), .Y (n_7478));
NAND2X1 g129368(.A (n_7476), .B (n_7475), .Y (n_7477));
NOR2X1 g129376(.A (n_143), .B (n_7473), .Y (n_7474));
NOR2X1 g129379(.A (n_323), .B (n_7295), .Y (n_7472));
NOR2X1 g129229(.A (n_225), .B (n_7295), .Y (n_7471));
NOR2X1 g129389(.A (n_156), .B (n_7469), .Y (n_7470));
NOR2X1 g129399(.A (n_261), .B (n_7469), .Y (n_7468));
NOR2X1 g129405(.A (n_5), .B (n_7466), .Y (n_7467));
NOR2X1 g129409(.A (n_79), .B (n_7484), .Y (n_7465));
NAND2X1 g129421(.A (n_9067), .B (n_7939), .Y (n_32086));
NOR2X1 g129425(.A (n_267), .B (n_7484), .Y (n_7463));
NOR2X1 g129427(.A (n_230), .B (n_7373), .Y (n_7462));
NOR2X1 g129439(.A (n_2832), .B (n_7481), .Y (n_7461));
NOR2X1 g129441(.A (n_3262), .B (n_7459), .Y (n_7460));
AOI22X1 g129477(.A0 (n_4190), .A1 (n_7457), .B0 (n_4176), .B1(n_33068), .Y (n_7458));
INVX8 g128891(.A (n_7415), .Y (n_8245));
AOI22X1 g129487(.A0 (n_4892), .A1 (n_33068), .B0 (n_4748), .B1(n_7457), .Y (n_7455));
AOI22X1 g129493(.A0 (n_4648), .A1 (n_33068), .B0 (n_4410), .B1(n_7457), .Y (n_7454));
AOI22X1 g129500(.A0 (n_3919), .A1 (n_33068), .B0 (n_3850), .B1(n_7457), .Y (n_7452));
INVX2 g129558(.A (n_15628), .Y (n_7581));
INVX1 g129563(.A (n_15763), .Y (n_15946));
CLKBUFX3 g129570(.A (n_15399), .Y (n_15708));
INVX1 g129614(.A (n_7444), .Y (n_7445));
CLKBUFX3 g129654(.A (n_7556), .Y (n_9692));
INVX2 g129656(.A (n_7595), .Y (n_7930));
INVX2 g129682(.A (n_7443), .Y (n_7926));
INVX2 g129720(.A (n_7657), .Y (n_7798));
INVX2 g129728(.A (n_7442), .Y (n_8209));
NAND2X1 g129754(.A (n_4320), .B (n_33897), .Y (n_7441));
NAND2X1 g129755(.A (n_32445), .B (n_33897), .Y (n_7440));
NAND2X1 g129772(.A (n_3854), .B (n_33897), .Y (n_7438));
NAND2X1 g129793(.A (n_3855), .B (n_33897), .Y (n_7437));
NAND2X1 g129794(.A (n_3862), .B (n_7362), .Y (n_7436));
NOR2X1 g129211(.A (n_381), .B (n_7434), .Y (n_7435));
NOR2X1 g129891(.A (n_2878), .B (n_7432), .Y (n_7433));
NOR2X1 g129894(.A (n_3170), .B (n_7432), .Y (n_7431));
NAND2X1 g129205(.A (P1_reg_174), .B (n_8177), .Y (n_7430));
CLKBUFX1 g129976(.A (n_13230), .Y (n_13393));
INVX1 g130067(.A (n_7428), .Y (n_7429));
NOR2X1 g130093(.A (n_6495), .B (n_7393), .Y (n_7427));
NAND2X1 g130096(.A (n_4205), .B (n_7426), .Y (n_8150));
NAND2X1 g130097(.A (n_34232), .B (n_7132), .Y (n_8365));
NAND2X1 g130100(.A (n_35188), .B (n_7426), .Y (n_8153));
INVX1 g128761(.A (n_7422), .Y (n_7975));
NAND2X2 g128759(.A (n_7156), .B (n_6971), .Y (n_7970));
NAND2X1 g130094(.A (n_4432), .B (n_7132), .Y (n_8344));
AOI22X1 g130601(.A0 (n_3517), .A1 (n_7418), .B0 (P3_reg3[24] ), .B1(n_7417), .Y (n_7420));
AOI22X1 g130602(.A0 (n_3519), .A1 (n_7418), .B0 (P3_reg3[20] ), .B1(n_7417), .Y (n_7419));
NAND2X1 g127918(.A (n_6336), .B (n_7415), .Y (n_7603));
AOI22X1 g130615(.A0 (n_4060), .A1 (n_6769), .B0 (P1_reg3[25] ), .B1(P1_n_449), .Y (n_7414));
AND2X1 g128375(.A (n_7259), .B (n_7326), .Y (n_7743));
AOI22X1 g130623(.A0 (n_4696), .A1 (n_6763), .B0 (P3_reg3[22] ), .B1(n_7390), .Y (n_7411));
NOR2X1 g129174(.A (n_207), .B (n_7407), .Y (n_7408));
NOR2X1 g129257(.A (n_192), .B (n_7469), .Y (n_7406));
INVX1 g128694(.A (n_7405), .Y (n_7805));
INVX4 g130036(.A (n_7403), .Y (n_15725));
NOR2X1 g129344(.A (n_229), .B (n_7469), .Y (n_7404));
AOI22X1 g130624(.A0 (n_4030), .A1 (n_7418), .B0 (P3_reg3[25] ), .B1(n_7417), .Y (n_7402));
NOR2X1 g127287(.A (n_7558), .B (n_6322), .Y (n_7987));
INVX1 g129731(.A (n_7442), .Y (n_7638));
NAND2X1 g130099(.A (n_4764), .B (n_7132), .Y (n_8432));
INVX1 g129732(.A (n_7442), .Y (n_7401));
NOR2X1 g128656(.A (n_7393), .B (n_8304), .Y (n_7400));
AND2X1 g127787(.A (n_7171), .B (n_7398), .Y (n_7399));
AND2X1 g128220(.A (n_7397), .B (n_7541), .Y (n_7745));
NAND2X2 g126445(.A (n_7396), .B (n_7395), .Y (n_8309));
NOR2X1 g128607(.A (n_7393), .B (n_7325), .Y (n_7394));
AOI22X1 g130603(.A0 (n_4368), .A1 (n_6763), .B0 (P3_reg3[27] ), .B1(n_7390), .Y (n_7391));
NAND2X1 g127697(.A (P1_d), .B (n_7397), .Y (n_7389));
INVX2 g130117(.A (n_33906), .Y (n_7793));
INVX2 g129749(.A (n_7571), .Y (n_7983));
NAND2X1 g129675(.A (n_7267), .B (n_33071), .Y (n_7640));
NOR2X1 g126201(.A (n_7387), .B (n_7770), .Y (n_8316));
OR2X1 g126583(.A (n_6387), .B (n_7561), .Y (n_7386));
NOR2X1 g129356(.A (n_114), .B (n_7373), .Y (n_7385));
NAND2X1 g129397(.A (P2_reg2[3] ), .B (n_7380), .Y (n_7381));
INVX1 g127086(.A (n_7379), .Y (n_7763));
INVX4 g129613(.A (n_7444), .Y (n_7917));
NOR2X1 g129440(.A (n_3295), .B (n_7007), .Y (n_7378));
AOI21X1 g129093(.A0 (n_7376), .A1 (n_13675), .B0 (n_7152), .Y(n_35612));
NOR2X1 g129414(.A (n_288), .B (n_7134), .Y (n_7375));
INVX1 g130214(.A (n_7616), .Y (n_8413));
NOR2X1 g129388(.A (n_142), .B (n_7373), .Y (n_7374));
NOR2X1 g129349(.A (n_173), .B (n_7012), .Y (n_7372));
NOR2X1 g129244(.A (n_2175), .B (n_7369), .Y (n_7370));
NAND2X1 g129426(.A (P1_reg_180), .B (n_8177), .Y (n_7368));
AOI21X1 g129058(.A0 (n_10854), .A1 (n_7534), .B0 (n_7146), .Y(n_7367));
AOI22X1 g130617(.A0 (n_3558), .A1 (n_6769), .B0 (P1_reg3[28] ), .B1(n_7245), .Y (n_32318));
NAND2X1 g129176(.A (P2_reg1[10] ), .B (n_7255), .Y (n_32087));
AOI22X1 g130613(.A0 (n_3651), .A1 (n_7418), .B0 (P3_reg3[23] ), .B1(n_7417), .Y (n_7364));
NAND2X1 g129773(.A (n_4040), .B (n_7362), .Y (n_7363));
AOI21X1 g129050(.A0 (P3_reg1[6] ), .A1 (n_34586), .B0 (n_7010), .Y(n_7361));
NOR2X1 g129386(.A (n_7), .B (n_7373), .Y (n_7360));
NOR2X1 g129375(.A (n_4039), .B (n_7205), .Y (n_7359));
NOR2X1 g129707(.A (n_3911), .B (n_7340), .Y (n_7358));
CLKBUFX1 g130002(.A (n_12953), .Y (n_13527));
INVX2 g129615(.A (n_7473), .Y (n_7444));
NAND2X1 g128926(.A (n_7327), .B (n_7025), .Y (n_7519));
NOR2X1 g129979(.A (n_6237), .B (n_6959), .Y (n_7354));
INVX1 g129565(.A (n_7298), .Y (n_16230));
NAND2X1 g127087(.A (n_7343), .B (n_7353), .Y (n_7379));
INVX1 g127088(.A (n_7387), .Y (n_7771));
OR2X1 g127146(.A (n_7343), .B (n_7353), .Y (n_7777));
NOR2X1 g129961(.A (n_6559), .B (n_6959), .Y (n_7352));
NOR2X1 g129959(.A (n_5937), .B (n_6959), .Y (n_7351));
INVX1 g129591(.A (n_7348), .Y (n_7349));
INVX1 g129580(.A (n_7434), .Y (n_8485));
NOR2X1 g127405(.A (n_7346), .B (n_7173), .Y (n_7347));
NOR2X1 g127406(.A (n_7344), .B (n_7343), .Y (n_7345));
NAND2X1 g129927(.A (n_3308), .B (n_7280), .Y (n_8048));
INVX1 g128948(.A (n_7395), .Y (n_7342));
NOR2X1 g129543(.A (n_3444), .B (n_7340), .Y (n_7341));
NOR2X1 g129544(.A (n_3471), .B (n_7340), .Y (n_7339));
CLKBUFX3 g129631(.A (n_7293), .Y (n_7553));
NOR2X1 g129276(.A (n_9038), .B (n_7312), .Y (n_7338));
INVX2 g129605(.A (n_7380), .Y (n_7662));
NOR2X1 g128605(.A (n_6283), .B (n_7782), .Y (n_7337));
OR2X1 g128606(.A (n_7188), .B (n_7770), .Y (n_7335));
NOR2X1 g128613(.A (n_6965), .B (n_7170), .Y (n_8008));
INVX1 g128668(.A (n_7558), .Y (n_7528));
NOR2X1 g128678(.A (n_7334), .B (n_35668), .Y (n_7525));
INVX1 g128683(.A (n_7332), .Y (n_7333));
NOR2X1 g128691(.A (n_6877), .B (n_35667), .Y (n_7331));
NAND2X1 g128695(.A (n_35667), .B (n_7329), .Y (n_7405));
NAND2X1 g128760(.A (n_7327), .B (n_7169), .Y (n_7328));
AND2X1 g128612(.A (n_7177), .B (n_7172), .Y (n_7531));
INVX1 g128922(.A (n_7326), .Y (n_7748));
INVX1 g128936(.A (n_7325), .Y (n_7986));
NOR2X1 g128940(.A (n_7024), .B (n_8060), .Y (n_7773));
NOR2X1 g129133(.A (n_137), .B (n_6868), .Y (n_7323));
NOR2X1 g129140(.A (n_210), .B (n_7190), .Y (n_7322));
NOR2X1 g129144(.A (n_154), .B (n_7230), .Y (n_7321));
NOR2X1 g129146(.A (n_7197), .B (n_172), .Y (n_7320));
NOR2X1 g129177(.A (n_198), .B (n_6868), .Y (n_7319));
NAND2X1 g129179(.A (P2_reg1[8] ), .B (n_7935), .Y (n_7318));
NAND2X1 g129225(.A (P1_reg2[0] ), .B (n_7201), .Y (n_7317));
NAND2X1 g129258(.A (P1_reg2[19] ), .B (n_7270), .Y (n_7316));
NOR2X1 g129265(.A (n_204), .B (n_7205), .Y (n_7315));
NOR2X1 g129277(.A (n_3601), .B (n_7310), .Y (n_7314));
NOR2X1 g129279(.A (n_127), .B (n_7312), .Y (n_7313));
NOR2X1 g129293(.A (n_2814), .B (n_7310), .Y (n_7311));
NOR2X1 g129318(.A (n_303), .B (n_7301), .Y (n_7309));
NAND2X1 g129373(.A (n_9592), .B (n_7307), .Y (n_7308));
NOR2X1 g129382(.A (n_373), .B (n_7301), .Y (n_7306));
NOR2X1 g129384(.A (n_300), .B (n_7205), .Y (n_7305));
NOR2X1 g129412(.A (n_268), .B (n_7301), .Y (n_7302));
NOR2X1 g129546(.A (n_3162), .B (n_6841), .Y (n_7299));
CLKBUFX3 g129560(.A (n_15396), .Y (n_15581));
CLKBUFX1 g129564(.A (n_7298), .Y (n_15763));
INVX2 g129571(.A (n_35154), .Y (n_15399));
INVX1 g129572(.A (n_35153), .Y (n_7297));
INVX1 g129582(.A (n_7295), .Y (n_7694));
INVX2 g129589(.A (n_7348), .Y (n_7672));
INVX2 g129590(.A (n_7348), .Y (n_7680));
INVX1 g129622(.A (n_7293), .Y (n_15536));
INVX2 g129634(.A (n_7293), .Y (n_7291));
INVX2 g129646(.A (n_7497), .Y (n_7944));
INVX2 g129678(.A (n_7355), .Y (n_7607));
INVX4 g129714(.A (n_7476), .Y (n_7998));
INVX1 g129724(.A (n_7369), .Y (n_7956));
INVX1 g129727(.A (n_7705), .Y (n_7290));
INVX2 g129739(.A (n_7289), .Y (n_8335));
INVX2 g129782(.A (n_7459), .Y (n_8197));
INVX4 g129787(.A (n_7287), .Y (n_7685));
NOR2X1 g129540(.A (n_3054), .B (n_6841), .Y (n_7286));
AOI21X1 g129824(.A0 (n_8113), .A1 (addr_1), .B0 (n_7040), .Y(n_7285));
AOI21X1 g129869(.A0 (n_4571), .A1 (n_6856), .B0 (n_6960), .Y(n_7284));
AOI21X1 g129873(.A0 (n_4009), .A1 (n_6856), .B0 (n_6993), .Y(n_7283));
NAND2X1 g129898(.A (n_3752), .B (n_7280), .Y (n_8147));
NAND2X1 g129921(.A (n_3240), .B (n_7280), .Y (n_8135));
NAND2X1 g129922(.A (n_6963), .B (n_7280), .Y (n_8139));
NAND2X1 g129926(.A (n_7280), .B (n_1803), .Y (n_8129));
NOR2X1 g129955(.A (n_4966), .B (n_6959), .Y (n_7279));
NOR2X1 g129956(.A (n_5508), .B (n_6959), .Y (n_7278));
NOR2X1 g129957(.A (n_5472), .B (n_6959), .Y (n_7276));
NOR2X1 g129958(.A (n_6194), .B (n_6959), .Y (n_7275));
NOR2X1 g129965(.A (n_6073), .B (n_6959), .Y (n_7273));
NOR2X1 g129967(.A (n_6453), .B (n_6959), .Y (n_7272));
NAND2X1 g129978(.A (n_7432), .B (n_7209), .Y (n_13230));
NAND2X1 g129236(.A (P1_reg2[14] ), .B (n_7270), .Y (n_32129));
NOR2X1 g130012(.A (n_6240), .B (n_6959), .Y (n_7269));
NOR2X1 g130020(.A (n_6122), .B (n_6959), .Y (n_7268));
INVX4 g130040(.A (n_15470), .Y (n_7403));
INVX1 g130044(.A (n_7267), .Y (n_15530));
NOR2X1 g130059(.A (n_6032), .B (n_6959), .Y (n_7266));
INVX1 g130191(.A (n_7432), .Y (n_8114));
INVX2 g129683(.A (n_7495), .Y (n_7443));
NOR2X1 g129248(.A (n_168), .B (n_7301), .Y (n_7262));
NAND2X1 g129285(.A (P2_reg_95), .B (n_7307), .Y (n_7260));
INVX1 g128762(.A (n_7259), .Y (n_7422));
NAND2X1 g129190(.A (P2_reg1[11] ), .B (n_7935), .Y (n_7258));
NOR2X1 g129188(.A (n_319), .B (n_6867), .Y (n_7257));
AOI22X1 g130599(.A0 (n_4147), .A1 (n_31536), .B0 (P3_reg3[26] ), .B1(n_31081), .Y (n_7254));
AOI22X1 g130600(.A0 (n_3965), .A1 (n_31536), .B0 (P3_reg3[21] ), .B1(n_31081), .Y (n_7253));
NOR2X1 g129181(.A (n_191), .B (n_7239), .Y (n_7252));
AOI22X1 g130605(.A0 (n_3455), .A1 (n_7250), .B0 (P1_reg3[27] ), .B1(P1_n_449), .Y (n_35265));
AOI22X1 g130607(.A0 (n_3645), .A1 (n_6436), .B0 (P1_reg3[24] ), .B1(n_7245), .Y (n_7249));
AOI22X1 g130611(.A0 (n_3268), .A1 (n_7250), .B0 (P1_reg3[23] ), .B1(P1_n_449), .Y (n_35924));
AOI22X1 g130626(.A0 (n_3808), .A1 (n_6436), .B0 (P1_reg3[22] ), .B1(n_7245), .Y (n_7246));
NAND3X1 g130832(.A (n_25823), .B (n_13387), .C (n_7243), .Y (n_7244));
NOR2X1 g129287(.A (P3_reg_148), .B (n_7301), .Y (n_7242));
NOR2X1 g129290(.A (P3_reg_153), .B (n_7301), .Y (n_7241));
NOR2X1 g129169(.A (n_362), .B (n_7239), .Y (n_7240));
AOI21X1 g129057(.A0 (P3_reg1[3] ), .A1 (n_7210), .B0 (n_6972), .Y(n_7238));
AOI22X1 g130608(.A0 (n_3602), .A1 (n_7250), .B0 (P1_reg3[21] ), .B1(P1_n_449), .Y (n_7237));
NAND2X1 g129274(.A (n_10128), .B (n_7722), .Y (n_7236));
INVX2 g129721(.A (n_7466), .Y (n_7657));
CLKBUFX3 g129655(.A (n_7255), .Y (n_7556));
NOR2X1 g129162(.A (n_376), .B (n_7137), .Y (n_7233));
CLKBUFX3 g129559(.A (n_15396), .Y (n_15628));
INVX1 g128672(.A (n_7232), .Y (n_7527));
INVX1 g128662(.A (n_7552), .Y (n_7536));
NOR2X1 g129142(.A (n_331), .B (n_7230), .Y (n_7231));
INVX2 g129733(.A (n_7705), .Y (n_7442));
NAND2X1 g129408(.A (n_11135), .B (n_7534), .Y (n_7228));
INVX1 g129777(.A (n_7754), .Y (n_7669));
NOR2X1 g129369(.A (P3_reg_152), .B (n_7301), .Y (n_7227));
INVX1 g130105(.A (n_7362), .Y (n_7597));
NOR2X1 g130054(.A (n_6265), .B (n_6959), .Y (n_7225));
NOR2X1 g130068(.A (n_4051), .B (n_7027), .Y (n_7428));
NOR2X1 g130021(.A (n_6333), .B (n_6959), .Y (n_7224));
CLKBUFX1 g130003(.A (n_12953), .Y (n_13112));
NAND2X1 g129928(.A (n_2950), .B (n_7280), .Y (n_8143));
INVX2 g129750(.A (n_7939), .Y (n_7571));
INVX1 g129677(.A (n_7355), .Y (n_7702));
NAND2X1 g129268(.A (n_9599), .B (n_7221), .Y (n_7222));
CLKBUFX1 g130215(.A (n_7426), .Y (n_7616));
NOR2X1 g129964(.A (n_6235), .B (n_6959), .Y (n_7219));
NAND3X1 g129325(.A (n_7217), .B (n_7216), .C (n_33068), .Y (n_7218));
INVX1 g127144(.A (n_7396), .Y (n_7383));
INVX1 g129778(.A (n_7754), .Y (n_7214));
CLKBUFX3 g129716(.A (n_7213), .Y (n_8192));
INVX1 g129658(.A (n_7255), .Y (n_7595));
NOR2X1 g129381(.A (P3_reg_151), .B (n_7301), .Y (n_7212));
AOI21X1 g129094(.A0 (n_7210), .A1 (P3_reg1[1] ), .B0 (n_6845), .Y(n_35613));
NOR2X1 g129420(.A (n_95), .B (n_7192), .Y (n_7208));
NOR2X1 g129294(.A (n_363), .B (n_7312), .Y (n_7207));
NOR2X1 g129288(.A (n_4265), .B (n_7205), .Y (n_7206));
NAND2X1 g129259(.A (n_14513), .B (n_7034), .Y (n_7204));
NAND2X1 g129275(.A (P3_reg2[29] ), .B (n_7714), .Y (n_7203));
NAND2X1 g129227(.A (P1_reg2[1] ), .B (n_7201), .Y (n_7202));
NAND2X1 g128920(.A (n_35667), .B (n_7200), .Y (n_7522));
NAND2X1 g129178(.A (P2_reg1[3] ), .B (n_7255), .Y (n_7199));
NOR2X1 g129164(.A (n_109), .B (n_7197), .Y (n_7198));
NAND2X1 g129159(.A (n_13689), .B (n_7584), .Y (n_7196));
NAND2X1 g129156(.A (n_13732), .B (n_7584), .Y (n_7195));
NOR2X1 g129151(.A (n_174), .B (n_7239), .Y (n_7194));
AOI21X1 g129101(.A0 (n_2718), .A1 (n_7210), .B0 (n_6838), .Y(n_7193));
INVX1 g129725(.A (n_7534), .Y (n_7369));
INVX1 g129717(.A (n_7192), .Y (n_7213));
NOR2X1 g130796(.A (n_3038), .B (n_7074), .Y (n_7191));
INVX2 g129685(.A (n_7190), .Y (n_7495));
NOR2X1 g129245(.A (n_346), .B (n_6762), .Y (n_7189));
NAND2X1 g127089(.A (n_7187), .B (n_7188), .Y (n_7387));
NOR2X1 g127145(.A (n_7187), .B (n_7188), .Y (n_7396));
NOR2X1 g129249(.A (n_324), .B (n_7181), .Y (n_7186));
OR2X1 g127294(.A (n_6977), .B (n_7353), .Y (n_7561));
INVX1 g129581(.A (n_7270), .Y (n_7434));
INVX2 g129583(.A (n_7270), .Y (n_7295));
NOR2X1 g129250(.A (n_85), .B (n_7181), .Y (n_7182));
OR2X1 g128941(.A (n_30897), .B (n_6441), .Y (n_8304));
NAND2X1 g130338(.A (n_6986), .B (n_4215), .Y (n_7180));
NAND2X1 g129542(.A (n_3063), .B (n_33895), .Y (n_7179));
INVX1 g128692(.A (n_7177), .Y (n_7397));
XOR2X1 g128669(.A (n_35390), .B (n_6724), .Y (n_7558));
NAND2X1 g130404(.A (n_6986), .B (n_10128), .Y (n_7175));
INVX1 g128673(.A (n_7173), .Y (n_7232));
INVX1 g128684(.A (n_7172), .Y (n_7332));
NAND2X1 g128686(.A (n_7154), .B (n_6985), .Y (n_7398));
INVX1 g128687(.A (n_7170), .Y (n_7171));
NAND2X1 g128763(.A (n_7168), .B (n_7169), .Y (n_7259));
NOR2X1 g128839(.A (n_6970), .B (n_7168), .Y (n_7530));
NOR2X1 g128949(.A (n_7165), .B (n_8060), .Y (n_7395));
OR2X1 g128937(.A (n_30897), .B (n_6495), .Y (n_7325));
AND2X1 g128933(.A (n_30897), .B (n_6495), .Y (n_7994));
NAND2X1 g129213(.A (n_13635), .B (n_7722), .Y (n_7163));
NOR2X1 g129220(.A (n_73), .B (n_7159), .Y (n_7162));
NAND2X1 g129237(.A (n_10189), .B (n_7722), .Y (n_7161));
NOR2X1 g129241(.A (n_151), .B (n_7159), .Y (n_7160));
NAND2X1 g129243(.A (n_13330), .B (n_7716), .Y (n_7158));
NAND2X1 g130317(.A (n_6979), .B (n_3333), .Y (n_7157));
INVX1 g129506(.A (n_7327), .Y (n_7156));
NAND2X1 g128914(.A (n_7154), .B (n_6983), .Y (n_7155));
NOR2X1 g129295(.A (n_286), .B (n_7151), .Y (n_7153));
NOR2X1 g129296(.A (n_289), .B (n_7151), .Y (n_7152));
NOR2X1 g129297(.A (n_389), .B (n_7151), .Y (n_7150));
NOR2X1 g129233(.A (n_164), .B (n_7159), .Y (n_7149));
NAND2X1 g129315(.A (n_10173), .B (n_7722), .Y (n_7148));
NOR2X1 g129222(.A (n_121), .B (n_7181), .Y (n_7146));
NAND2X1 g129230(.A (n_10156), .B (n_7722), .Y (n_7145));
NOR2X1 g129226(.A (P3_reg_145), .B (n_7042), .Y (n_7144));
NOR2X1 g129418(.A (n_365), .B (n_7159), .Y (n_7143));
NAND2X1 g129224(.A (n_10187), .B (n_7722), .Y (n_7142));
INVX2 g129636(.A (n_7092), .Y (n_15387));
INVX1 g129504(.A (n_35668), .Y (n_7523));
NOR2X1 g129218(.A (n_243), .B (n_7159), .Y (n_7140));
INVX1 g129566(.A (n_7139), .Y (n_7298));
INVX2 g129575(.A (n_7183), .Y (n_7373));
INVX2 g129598(.A (n_7714), .Y (n_7484));
INVX1 g129662(.A (n_7953), .Y (n_7407));
INVX4 g129698(.A (n_7136), .Y (n_8177));
INVX1 g129736(.A (n_7534), .Y (n_7135));
INVX4 g129740(.A (n_7307), .Y (n_7289));
INVX1 g129743(.A (n_7221), .Y (n_7134));
INVX1 g129783(.A (n_34590), .Y (n_7459));
CLKBUFX3 g129788(.A (n_7538), .Y (n_7287));
AOI22X1 g129883(.A0 (n_6398), .A1 (n_8409), .B0 (n_6302), .B1(n_8407), .Y (n_7133));
CLKBUFX1 g130005(.A (n_34355), .Y (n_12953));
NAND2X1 g130065(.A (n_4099), .B (n_7132), .Y (n_7894));
NAND2X1 g130102(.A (n_4632), .B (n_7132), .Y (n_7813));
NAND2X1 g130130(.A (n_4599), .B (n_7132), .Y (n_7879));
NOR2X1 g130131(.A (n_6387), .B (n_6283), .Y (n_7131));
NAND2X1 g130312(.A (P1_reg1[30] ), .B (n_7124), .Y (n_7128));
NOR2X1 g129196(.A (n_148), .B (n_7181), .Y (n_7127));
NAND2X1 g130333(.A (n_6986), .B (P1_reg_173), .Y (n_7126));
NAND2X1 g130336(.A (n_7124), .B (n_10886), .Y (n_7125));
NAND2X1 g130343(.A (n_6979), .B (n_4824), .Y (n_7123));
NAND2X1 g130398(.A (n_7120), .B (n_4561), .Y (n_7122));
NAND2X1 g130407(.A (n_7120), .B (P1_reg2[9] ), .Y (n_7121));
NAND2X1 g130409(.A (n_7120), .B (P1_reg1[24] ), .Y (n_7119));
NAND2X1 g130410(.A (n_7120), .B (n_10167), .Y (n_7118));
NAND2X1 g130419(.A (n_6979), .B (n_11120), .Y (n_35697));
NAND2X1 g130420(.A (n_6986), .B (n_10189), .Y (n_7116));
NAND2X1 g130422(.A (n_6979), .B (n_4534), .Y (n_7115));
NAND2X1 g130429(.A (n_6986), .B (n_10201), .Y (n_7113));
NAND2X1 g130442(.A (P1_reg2[30] ), .B (n_7124), .Y (n_7112));
NAND2X1 g130449(.A (n_6979), .B (n_11141), .Y (n_7111));
NAND2X1 g130451(.A (n_6979), .B (n_10191), .Y (n_7110));
NAND2X1 g130460(.A (n_6979), .B (n_10182), .Y (n_7109));
NAND2X1 g130481(.A (n_7120), .B (n_3958), .Y (n_7107));
INVX2 g129715(.A (n_7192), .Y (n_7476));
NAND2X1 g130538(.A (n_6986), .B (n_10144), .Y (n_7106));
NAND2X1 g130557(.A (n_6986), .B (n_10187), .Y (n_7105));
NAND2X1 g130567(.A (n_6986), .B (n_11136), .Y (n_7104));
NAND2X1 g130579(.A (n_6979), .B (n_4920), .Y (n_7103));
NAND2X1 g130592(.A (n_7124), .B (n_10161), .Y (n_7102));
AOI22X1 g130610(.A0 (n_3364), .A1 (n_6446), .B0 (P2_reg3[23] ), .B1(n_34375), .Y (n_35098));
AOI22X1 g130612(.A0 (n_3991), .A1 (n_6446), .B0 (P2_reg3[25] ), .B1(n_33350), .Y (n_7098));
AOI22X1 g130618(.A0 (n_3436), .A1 (n_6446), .B0 (P2_reg3[20] ), .B1(n_34375), .Y (n_7096));
AOI22X1 g130620(.A0 (n_3582), .A1 (n_6446), .B0 (P2_reg3[22] ), .B1(n_33350), .Y (n_7094));
CLKBUFX3 g129635(.A (n_7092), .Y (n_7293));
INVX4 g129641(.A (n_7137), .Y (n_7503));
NOR2X1 g130777(.A (n_3186), .B (n_7077), .Y (n_7091));
NOR2X1 g130782(.A (n_1985), .B (n_7077), .Y (n_7090));
NOR2X1 g130785(.A (n_879), .B (n_7074), .Y (n_7088));
NOR2X1 g130793(.A (n_3034), .B (n_7077), .Y (n_7086));
NOR2X1 g130795(.A (n_3387), .B (n_7077), .Y (n_7085));
NOR2X1 g130800(.A (n_3481), .B (n_7077), .Y (n_7084));
NOR2X1 g130801(.A (n_3161), .B (n_7074), .Y (n_7083));
NOR2X1 g130804(.A (n_3357), .B (n_7074), .Y (n_7082));
NOR3X1 g130805(.A (n_9909), .B (P1_reg3[3] ), .C (n_1587), .Y(n_7081));
NOR2X1 g130808(.A (n_2177), .B (n_8933), .Y (n_7079));
NOR2X1 g130810(.A (n_2608), .B (n_7077), .Y (n_7078));
NOR3X1 g130811(.A (n_12753), .B (n_9313), .C (n_7058), .Y (n_7076));
NOR2X1 g130812(.A (n_3691), .B (n_7074), .Y (n_7075));
NOR3X1 g130818(.A (n_10736), .B (n_2096), .C (n_7058), .Y (n_7073));
NOR3X1 g130819(.A (n_10736), .B (P3_reg3[3] ), .C (n_7062), .Y(n_7071));
NOR2X1 g130820(.A (n_3779), .B (n_7074), .Y (n_7069));
NOR2X1 g130821(.A (n_1722), .B (n_8933), .Y (n_7068));
NOR2X1 g130827(.A (n_3133), .B (n_7077), .Y (n_7065));
INVX2 g129647(.A (n_7584), .Y (n_7497));
CLKBUFX3 g129722(.A (n_7192), .Y (n_7466));
INVX4 g130041(.A (n_34472), .Y (n_15470));
CLKBUFX3 g129726(.A (n_7534), .Y (n_7736));
NOR3X1 g130783(.A (n_12753), .B (n_3269), .C (n_7058), .Y (n_7059));
INVX1 g128663(.A (n_7343), .Y (n_7552));
NOR2X1 g129215(.A (n_224), .B (n_7159), .Y (n_7057));
NAND2X1 g130395(.A (n_6979), .B (n_3693), .Y (n_7055));
NAND2X1 g129150(.A (n_13322), .B (n_7052), .Y (n_7054));
NAND2X1 g129145(.A (P1_reg1[0] ), .B (n_7052), .Y (n_7053));
AOI22X1 g130616(.A0 (n_4027), .A1 (n_6446), .B0 (P2_reg3[26] ), .B1(n_1336), .Y (n_7051));
NOR2X1 g129253(.A (n_384), .B (n_7159), .Y (n_7050));
NAND2X1 g130101(.A (n_4461), .B (n_7132), .Y (n_7884));
INVX1 g129735(.A (n_7534), .Y (n_7049));
NAND2X1 g130490(.A (P1_reg_180), .B (n_7124), .Y (n_7048));
NAND2X1 g130103(.A (n_4131), .B (n_7132), .Y (n_7849));
CLKBUFX2 g130045(.A (n_34472), .Y (n_7267));
INVX1 g130106(.A (n_33896), .Y (n_7362));
NOR2X1 g129424(.A (P3_reg_147), .B (n_7012), .Y (n_7046));
INVX1 g129595(.A (n_7205), .Y (n_8183));
NOR2X1 g129278(.A (n_7043), .B (n_7042), .Y (n_7044));
CLKBUFX3 g129751(.A (n_7221), .Y (n_7939));
INVX1 g130074(.A (n_7040), .Y (n_7041));
NAND2X1 g130127(.A (n_4911), .B (n_7132), .Y (n_7904));
AOI22X1 g130619(.A0 (n_4439), .A1 (n_6446), .B0 (P2_reg3[28] ), .B1(n_34375), .Y (n_35076));
INVX1 g129607(.A (n_33269), .Y (n_7380));
INVX2 g129680(.A (n_7197), .Y (n_7355));
CLKBUFX3 g129616(.A (n_33269), .Y (n_7473));
NOR2X1 g130826(.A (n_2929), .B (n_10736), .Y (n_7033));
NAND2X1 g130480(.A (n_7120), .B (n_11327), .Y (n_32272));
NAND2X1 g129270(.A (n_14168), .B (n_7716), .Y (n_7031));
NAND2X1 g130492(.A (n_7120), .B (P1_reg_174), .Y (n_7030));
NAND2X1 g130491(.A (n_7120), .B (n_10546), .Y (n_35641));
INVX1 g129784(.A (n_34590), .Y (n_7481));
INVX1 g130216(.A (n_7027), .Y (n_7426));
CLKBUFX3 g129734(.A (n_7534), .Y (n_7705));
NOR2X1 g130792(.A (n_3611), .B (n_10736), .Y (n_7026));
NAND2X1 g128923(.A (n_7168), .B (n_7025), .Y (n_7326));
INVX2 g129592(.A (n_7312), .Y (n_7348));
AOI22X1 g129864(.A0 (n_6321), .A1 (n_8409), .B0 (n_6271), .B1(n_8407), .Y (n_7022));
NOR2X1 g130823(.A (n_3550), .B (n_7074), .Y (n_7021));
NOR3X1 g130817(.A (n_9909), .B (n_2553), .C (n_31105), .Y (n_7020));
NOR2X1 g130822(.A (n_2823), .B (n_7077), .Y (n_7017));
NOR2X1 g130806(.A (n_3418), .B (n_8933), .Y (n_7016));
NOR2X1 g130784(.A (n_931), .B (n_7074), .Y (n_7015));
OR2X1 g128905(.A (n_7154), .B (n_6976), .Y (n_7415));
NOR2X1 g129403(.A (n_72), .B (n_34589), .Y (n_7014));
NOR2X1 g129393(.A (n_7012), .B (P3_reg_149), .Y (n_7013));
NOR2X1 g129359(.A (n_77), .B (n_6968), .Y (n_7011));
NOR2X1 g129314(.A (P3_reg_146), .B (n_7042), .Y (n_7010));
NOR2X1 g129272(.A (n_379), .B (n_7151), .Y (n_7009));
NOR2X1 g128924(.A (n_6832), .B (n_7168), .Y (n_7008));
INVX1 g129785(.A (n_34590), .Y (n_7007));
INVX2 g129779(.A (n_7310), .Y (n_7754));
NAND2X1 g129147(.A (P1_reg1[1] ), .B (n_7052), .Y (n_7005));
INVX2 g129561(.A (n_6861), .Y (n_15396));
NOR2X1 g129137(.A (n_209), .B (n_34585), .Y (n_7004));
INVX2 g129756(.A (n_7034), .Y (n_7469));
NOR2X1 g129390(.A (n_215), .B (n_7012), .Y (n_7003));
INVX4 g129737(.A (n_6785), .Y (n_7534));
NOR2X1 g130828(.A (n_3166), .B (n_6892), .Y (n_7001));
NAND2X1 g129567(.A (n_34353), .B (n_6547), .Y (n_7139));
NAND2X1 g129934(.A (n_6990), .B (n_1803), .Y (n_8128));
NOR2X1 g130815(.A (n_3281), .B (n_6901), .Y (n_6999));
NAND2X1 g129942(.A (n_4432), .B (n_6990), .Y (n_8343));
NOR2X1 g130809(.A (n_2730), .B (n_6996), .Y (n_6998));
NOR2X1 g130788(.A (n_3403), .B (n_6996), .Y (n_6997));
NOR2X1 g130787(.A (n_1735), .B (n_9909), .Y (n_6995));
NAND2X1 g130366(.A (n_6986), .B (n_4477), .Y (n_6994));
INVX2 g129686(.A (n_7052), .Y (n_7190));
NOR2X1 g129992(.A (n_4077), .B (n_6959), .Y (n_6993));
NAND2X1 g130319(.A (n_6979), .B (n_3716), .Y (n_6992));
INVX2 g129648(.A (n_34585), .Y (n_7584));
NAND2X1 g130060(.A (n_6149), .B (n_8409), .Y (n_8345));
INVX2 g129577(.A (n_7181), .Y (n_7183));
NAND2X1 g129949(.A (n_4764), .B (n_6990), .Y (n_8431));
NAND2X1 g129947(.A (n_4131), .B (n_6990), .Y (n_7848));
NAND2X1 g129938(.A (n_3752), .B (n_6990), .Y (n_8146));
NAND2X1 g129944(.A (n_6988), .B (n_6990), .Y (n_8427));
NAND2X1 g130322(.A (n_6986), .B (n_3402), .Y (n_6987));
NAND2X1 g128693(.A (n_6984), .B (n_6985), .Y (n_7177));
NAND2X1 g128685(.A (n_6984), .B (n_6983), .Y (n_7172));
NAND2X1 g130400(.A (n_6979), .B (P1_reg1[19] ), .Y (n_6982));
NAND2X1 g130394(.A (n_6979), .B (n_3668), .Y (n_6980));
INVX1 g128675(.A (n_7187), .Y (n_7173));
NOR2X1 g128688(.A (n_6976), .B (n_6984), .Y (n_7170));
INVX1 g129513(.A (n_7165), .Y (n_7024));
NAND2X1 g128938(.A (n_6797), .B (n_8060), .Y (n_7770));
INVX1 g128942(.A (n_6975), .Y (n_7774));
INVX1 g128931(.A (n_6974), .Y (n_7166));
NAND3X1 g129254(.A (n_13640), .B (n_6466), .C (n_6290), .Y (n_6973));
NOR2X1 g129262(.A (n_196), .B (n_6844), .Y (n_6972));
INVX1 g129535(.A (n_6970), .Y (n_6971));
NOR2X1 g129549(.A (n_6860), .B (n_6876), .Y (n_7200));
INVX2 g129596(.A (n_35940), .Y (n_7205));
INVX1 g129688(.A (n_7052), .Y (n_7230));
INVX2 g129752(.A (n_6968), .Y (n_7221));
INVX2 g129760(.A (n_7012), .Y (n_7034));
INVX4 g129767(.A (n_7716), .Y (n_7301));
NOR2X1 g128838(.A (n_6356), .B (n_6984), .Y (n_6965));
NAND2X1 g129902(.A (n_2950), .B (n_6990), .Y (n_8142));
NAND2X1 g129903(.A (n_6964), .B (n_6990), .Y (n_7898));
NAND2X1 g129906(.A (n_6963), .B (n_6990), .Y (n_8138));
NAND2X1 g129937(.A (n_6962), .B (n_6990), .Y (n_8047));
NAND2X1 g129939(.A (n_4599), .B (n_6990), .Y (n_7878));
NAND2X1 g129940(.A (n_4205), .B (n_6990), .Y (n_8151));
NAND2X1 g129943(.A (n_4301), .B (n_6990), .Y (n_7888));
NAND2X1 g129945(.A (n_4461), .B (n_6990), .Y (n_7883));
NAND2X1 g129946(.A (n_4911), .B (n_6990), .Y (n_7903));
NAND2X1 g129948(.A (n_35188), .B (n_6990), .Y (n_8154));
NAND2X1 g129950(.A (n_4099), .B (n_6990), .Y (n_7893));
NAND2X1 g129951(.A (n_4632), .B (n_6990), .Y (n_7812));
NOR2X1 g129952(.A (n_6990), .B (n_8409), .Y (n_6961));
NOR2X1 g129953(.A (n_4569), .B (n_6959), .Y (n_6960));
NAND2X1 g129954(.A (n_6093), .B (n_8409), .Y (n_7815));
NAND2X1 g129960(.A (n_6098), .B (n_8409), .Y (n_7881));
NAND2X1 g129962(.A (n_4894), .B (n_8409), .Y (n_8140));
NAND2X1 g129963(.A (n_5433), .B (n_8409), .Y (n_8049));
NAND2X1 g130019(.A (n_6127), .B (n_8409), .Y (n_7906));
NAND2X1 g130049(.A (n_6005), .B (n_8409), .Y (n_7896));
NAND2X1 g130050(.A (n_3636), .B (n_8409), .Y (n_8144));
NAND2X1 g130051(.A (n_5495), .B (n_8409), .Y (n_7885));
NAND2X1 g130053(.A (n_4743), .B (n_8409), .Y (n_8148));
NAND2X1 g130057(.A (n_6331), .B (n_8409), .Y (n_6956));
NAND2X1 g130062(.A (n_6031), .B (n_8409), .Y (n_7850));
NAND2X1 g130132(.A (n_5832), .B (n_8407), .Y (n_7891));
NAND2X1 g130134(.A (n_6137), .B (n_8407), .Y (n_7814));
NAND2X1 g130136(.A (n_6096), .B (n_8407), .Y (n_7895));
NAND2X1 g130137(.A (n_6033), .B (n_8407), .Y (n_7851));
NAND2X1 g130138(.A (n_6066), .B (n_8407), .Y (n_7880));
NAND2X1 g130139(.A (n_6338), .B (n_8407), .Y (n_6954));
NAND2X1 g130144(.A (n_6222), .B (n_8407), .Y (n_8330));
NAND2X1 g130145(.A (n_6182), .B (n_8407), .Y (n_7905));
NAND2X1 g130146(.A (n_6124), .B (n_8407), .Y (n_8346));
NAND2X1 g130147(.A (n_6200), .B (n_8407), .Y (n_8429));
NAND2X1 g130149(.A (n_5529), .B (n_8407), .Y (n_7901));
NAND2X1 g130150(.A (n_5546), .B (n_8407), .Y (n_8050));
NAND3X1 g130151(.A (n_6856), .B (n_2319), .C (n_2460), .Y (n_8453));
INVX1 g130220(.A (n_6463), .Y (n_7280));
NAND2X1 g129890(.A (n_7967), .B (n_6990), .Y (n_6952));
OR2X1 g130303(.A (n_6950), .B (P1_reg1[27] ), .Y (n_6951));
OR2X1 g130307(.A (n_6950), .B (P1_reg1[28] ), .Y (n_32884));
NAND2X1 g130313(.A (n_6986), .B (P1_reg1[12] ), .Y (n_6948));
NAND2X1 g130315(.A (n_6979), .B (n_3235), .Y (n_6947));
NAND2X1 g130324(.A (n_6979), .B (n_4554), .Y (n_6945));
NAND2X1 g130325(.A (n_6979), .B (n_4011), .Y (n_6944));
NAND2X1 g130328(.A (n_6986), .B (n_10197), .Y (n_6943));
NAND2X1 g130329(.A (n_6979), .B (n_4151), .Y (n_6942));
NAND2X1 g130332(.A (n_6979), .B (n_4445), .Y (n_35645));
NAND2X1 g130334(.A (n_6938), .B (n_3337), .Y (n_6940));
NAND2X1 g130345(.A (n_6938), .B (P1_reg2[16] ), .Y (n_6939));
NAND2X1 g130356(.A (n_6938), .B (n_10171), .Y (n_6937));
NAND2X1 g130357(.A (n_6979), .B (n_10893), .Y (n_6936));
NAND2X1 g130368(.A (n_6979), .B (n_11148), .Y (n_35132));
NAND2X1 g130370(.A (n_6938), .B (n_10858), .Y (n_35142));
NAND2X1 g130374(.A (n_6938), .B (n_10150), .Y (n_6933));
NAND2X1 g130381(.A (n_6938), .B (n_4231), .Y (n_6932));
NAND2X1 g130387(.A (n_6979), .B (n_3259), .Y (n_6931));
NAND2X1 g130388(.A (n_6979), .B (n_4277), .Y (n_35121));
NAND2X1 g130392(.A (n_6986), .B (n_13640), .Y (n_6929));
NAND2X1 g130393(.A (n_6979), .B (n_3470), .Y (n_6928));
NAND2X1 g130435(.A (n_6986), .B (n_10138), .Y (n_6927));
NAND2X1 g130439(.A (n_6979), .B (n_10897), .Y (n_6926));
NAND2X1 g130446(.A (n_6938), .B (n_10245), .Y (n_32894));
NAND2X1 g130448(.A (n_6986), .B (n_10156), .Y (n_6924));
NAND2X1 g130463(.A (n_6979), .B (n_10211), .Y (n_6923));
NAND2X1 g130063(.A (n_6123), .B (n_8409), .Y (n_8428));
NAND2X1 g130466(.A (n_6986), .B (n_10178), .Y (n_6922));
NAND2X1 g130469(.A (n_6979), .B (n_4213), .Y (n_6921));
NAND2X1 g130489(.A (n_6979), .B (n_10136), .Y (n_35330));
NAND2X1 g130494(.A (n_6979), .B (n_3416), .Y (n_6919));
NAND2X1 g130498(.A (n_6986), .B (P1_reg1[14] ), .Y (n_6918));
NAND2X1 g130512(.A (n_6979), .B (n_10217), .Y (n_6917));
NAND2X1 g130516(.A (n_6979), .B (n_10148), .Y (n_6916));
NAND2X1 g130523(.A (n_6986), .B (n_10223), .Y (n_6914));
NAND2X1 g130529(.A (n_6986), .B (P1_reg1[0] ), .Y (n_6913));
NAND2X1 g130531(.A (n_6979), .B (n_10154), .Y (n_6912));
NAND2X1 g130532(.A (n_6938), .B (n_13635), .Y (n_6911));
NAND2X1 g130547(.A (n_6938), .B (n_10173), .Y (n_6910));
NAND2X1 g130548(.A (n_6979), .B (n_13322), .Y (n_6909));
NAND2X1 g130552(.A (n_6938), .B (P1_reg1[1] ), .Y (n_6908));
NAND2X1 g130554(.A (n_6938), .B (P1_reg2[14] ), .Y (n_32284));
NAND2X1 g130556(.A (n_6979), .B (P1_reg1[16] ), .Y (n_6906));
NAND2X1 g130581(.A (n_6979), .B (n_10219), .Y (n_32926));
NAND2X1 g130582(.A (n_6979), .B (n_10225), .Y (n_6904));
INVX2 g129643(.A (n_7210), .Y (n_7137));
AOI22X1 g130609(.A0 (n_3782), .A1 (n_35007), .B0 (P2_reg3[21] ), .B1(P2_n_749), .Y (n_6903));
NOR2X1 g130780(.A (n_3549), .B (n_6901), .Y (n_6902));
NOR2X1 g130781(.A (n_3392), .B (n_6901), .Y (n_6900));
NOR2X1 g130791(.A (n_3516), .B (n_9909), .Y (n_6899));
NOR2X1 g130797(.A (n_3071), .B (n_9909), .Y (n_6897));
NOR2X1 g130803(.A (n_2843), .B (n_9909), .Y (n_6896));
NOR2X1 g130807(.A (n_1758), .B (n_9909), .Y (n_6895));
NOR2X1 g130813(.A (n_3434), .B (n_6901), .Y (n_6894));
INVX1 g129585(.A (n_7159), .Y (n_7270));
NOR2X1 g130830(.A (n_3180), .B (n_6892), .Y (n_6893));
INVX1 g130980(.A (n_6891), .Y (n_25823));
INVX1 g130983(.A (n_6806), .Y (n_7418));
NAND2X1 g130354(.A (n_6938), .B (P1_reg2[19] ), .Y (n_6888));
NAND2X1 g129908(.A (n_6887), .B (n_6990), .Y (n_8134));
NAND2X1 g130052(.A (n_6266), .B (n_8409), .Y (n_8366));
NAND2X2 g129723(.A (n_6848), .B (n_35348), .Y (n_7192));
AND2X1 g130614(.A (n_2050), .B (n_6493), .Y (n_6885));
INVX2 g129599(.A (n_7151), .Y (n_7714));
INVX1 g128664(.A (n_6977), .Y (n_7343));
INVX1 g129663(.A (n_6883), .Y (n_7953));
INVX1 g129661(.A (n_6883), .Y (n_7935));
INVX1 g130193(.A (n_15685), .Y (n_7432));
NAND3X1 g130069(.A (n_8409), .B (n_2248), .C (n_2076), .Y (n_8130));
NAND2X1 g130421(.A (n_6979), .B (n_10158), .Y (n_6882));
NAND2X1 g130443(.A (n_6938), .B (n_10221), .Y (n_6881));
INVX2 g129789(.A (n_34589), .Y (n_7538));
NAND2X1 g129966(.A (n_5496), .B (n_8409), .Y (n_7900));
NAND2X1 g129550(.A (n_6876), .B (n_6858), .Y (n_6877));
INVX1 g130124(.A (n_33895), .Y (n_7340));
NAND2X1 g129941(.A (n_4623), .B (n_6990), .Y (n_8364));
NAND2X1 g130569(.A (n_6979), .B (n_4230), .Y (n_6875));
INVX1 g129507(.A (n_7168), .Y (n_7327));
NAND2X1 g130055(.A (n_6400), .B (n_8409), .Y (n_8434));
INVX2 g129742(.A (n_6968), .Y (n_7307));
NAND2X1 g130331(.A (n_6979), .B (n_4590), .Y (n_6874));
AOI21X1 g129870(.A0 (n_4745), .A1 (n_6856), .B0 (n_6718), .Y(n_6871));
INVX2 g129681(.A (n_7052), .Y (n_7197));
NAND2X1 g130465(.A (n_6938), .B (n_10180), .Y (n_6870));
NAND2X1 g130133(.A (n_5562), .B (n_8407), .Y (n_7886));
NAND2X1 g130361(.A (n_6979), .B (n_10165), .Y (n_6869));
INVX1 g129687(.A (n_7052), .Y (n_6868));
INVX1 g129689(.A (n_7052), .Y (n_6867));
INVX1 g130088(.A (n_6865), .Y (n_7653));
INVX2 g129780(.A (n_7376), .Y (n_7310));
INVX2 g129699(.A (n_7722), .Y (n_7136));
INVX1 g129690(.A (n_7052), .Y (n_7239));
NAND2X1 g130382(.A (n_6938), .B (n_11144), .Y (n_32557));
INVX2 g129660(.A (n_6883), .Y (n_7255));
INVX1 g129579(.A (n_7159), .Y (n_7201));
NAND2X1 g130510(.A (n_6979), .B (P1_reg2[1] ), .Y (n_6863));
NOR2X1 g129562(.A (n_6445), .B (n_32835), .Y (n_6861));
NAND2X2 g129527(.A (n_6860), .B (n_6876), .Y (n_7334));
NOR2X1 g129526(.A (n_6858), .B (n_6876), .Y (n_7329));
AOI21X1 g129868(.A0 (n_4302), .A1 (n_6856), .B0 (n_6544), .Y(n_6857));
NOR2X1 g130789(.A (n_3778), .B (n_6892), .Y (n_6855));
NOR2X1 g130825(.A (n_3215), .B (n_6892), .Y (n_6854));
NAND2X1 g130541(.A (n_6979), .B (n_10134), .Y (n_6853));
NOR2X1 g130779(.A (n_2971), .B (n_6996), .Y (n_6852));
NOR2X1 g130778(.A (n_3218), .B (n_6996), .Y (n_6851));
NAND2X1 g130583(.A (n_6986), .B (n_10205), .Y (n_6850));
INVX1 g130218(.A (n_7132), .Y (n_7027));
NAND2X1 g130495(.A (n_6986), .B (P1_reg_172), .Y (n_6847));
NOR2X1 g129387(.A (n_146), .B (n_6844), .Y (n_6845));
NAND2X1 g130459(.A (n_6938), .B (n_10215), .Y (n_35277));
NAND2X1 g130433(.A (n_6986), .B (n_10140), .Y (n_6842));
INVX1 g130122(.A (n_33895), .Y (n_6841));
NAND2X1 g130135(.A (n_6459), .B (n_8407), .Y (n_8433));
NAND2X1 g130467(.A (n_6986), .B (n_10175), .Y (n_6840));
NOR2X1 g129219(.A (n_336), .B (n_6844), .Y (n_6838));
INVX2 g129593(.A (n_35941), .Y (n_7312));
NOR2X1 g130075(.A (n_2498), .B (n_6959), .Y (n_7040));
NAND2X1 g130061(.A (n_5769), .B (n_8409), .Y (n_7890));
NAND2X1 g128934(.A (n_6833), .B (n_6837), .Y (n_7782));
INVX2 g129637(.A (n_6767), .Y (n_7092));
INVX1 g130906(.A (n_6436), .Y (n_9387));
INVX2 g129586(.A (n_6796), .Y (n_7159));
NOR2X1 g128943(.A (n_6835), .B (n_6837), .Y (n_6975));
NOR2X1 g129539(.A (n_6831), .B (n_6798), .Y (n_7169));
INVX4 g129761(.A (n_6836), .Y (n_7012));
NAND2X1 g128932(.A (n_6835), .B (n_6387), .Y (n_6974));
NAND3X1 g129269(.A (n_14317), .B (n_34393), .C (n_6402), .Y (n_6834));
NAND2X2 g129508(.A (n_6376), .B (n_6469), .Y (n_7168));
INVX1 g129520(.A (n_6833), .Y (n_6878));
NAND2X1 g129531(.A (n_6831), .B (n_6316), .Y (n_6832));
NOR2X1 g129537(.A (n_6831), .B (n_6316), .Y (n_7025));
NAND2X2 g129664(.A (n_35340), .B (n_35347), .Y (n_6883));
INVX4 g129692(.A (n_34535), .Y (n_7052));
INVX4 g129702(.A (n_6829), .Y (n_7722));
OR2X1 g130073(.A (n_33042), .B (n_6823), .Y (n_6825));
INVX1 g130090(.A (n_7457), .Y (n_6865));
OR2X1 g130128(.A (n_4046), .B (n_6823), .Y (n_6822));
NAND2X1 g130140(.A (n_4697), .B (n_8407), .Y (n_8032));
NAND3X1 g130148(.A (n_8407), .B (n_2239), .C (n_2428), .Y (n_8131));
INVX1 g130702(.A (n_6950), .Y (n_7120));
XOR2X1 g130639(.A (n_6394), .B (n_6392), .Y (n_6818));
CLKBUFX2 g129644(.A (n_34584), .Y (n_7210));
NOR3X1 g130776(.A (n_12597), .B (P2_reg3[3] ), .C (n_16415), .Y(n_6814));
XOR2X1 g129885(.A (n_6810), .B (n_6723), .Y (n_30897));
INVX1 g130911(.A (n_9909), .Y (n_29486));
INVX1 g130913(.A (n_9387), .Y (n_31480));
INVX1 g130974(.A (n_6806), .Y (n_12926));
INVX1 g130977(.A (n_31495), .Y (n_31536));
INVX1 g131008(.A (n_10342), .Y (n_7074));
INVX1 g131067(.A (n_31740), .Y (n_7077));
OR2X1 g130066(.A (n_6208), .B (n_6823), .Y (n_6803));
XOR2X1 g128676(.A (n_6802), .B (n_6401), .Y (n_7187));
XOR2X1 g128666(.A (n_34092), .B (n_6407), .Y (n_6977));
CLKBUFX2 g129781(.A (n_34588), .Y (n_7376));
NAND2X1 g130142(.A (n_3715), .B (n_8407), .Y (n_8034));
INVX2 g129600(.A (n_6800), .Y (n_7151));
NAND2X1 g130141(.A (n_5042), .B (n_8407), .Y (n_8014));
CLKBUFX3 g130194(.A (n_15622), .Y (n_15685));
NAND2X1 g129536(.A (n_6831), .B (n_6798), .Y (n_6970));
INVX2 g129514(.A (n_6797), .Y (n_7165));
NAND2X1 g130058(.A (n_4183), .B (n_8409), .Y (n_8121));
INVX1 g129578(.A (n_6796), .Y (n_7181));
INVX1 g130973(.A (n_6806), .Y (n_10399));
OR2X1 g130081(.A (n_4385), .B (n_6823), .Y (n_6793));
NOR2X1 g130824(.A (n_3382), .B (n_6389), .Y (n_6792));
NAND2X2 g129753(.A (n_35339), .B (n_35655), .Y (n_6968));
INVX1 g130982(.A (n_6787), .Y (n_6891));
INVX2 g129762(.A (n_6836), .Y (n_7042));
NAND2X2 g129738(.A (n_6414), .B (n_34534), .Y (n_6785));
INVX1 g130706(.A (n_6950), .Y (n_7124));
NOR2X1 g130786(.A (n_3331), .B (n_12597), .Y (n_6783));
NOR2X1 g130794(.A (n_3046), .B (n_12597), .Y (n_6782));
INVX1 g129522(.A (n_6984), .Y (n_7154));
NOR3X1 g130816(.A (n_12606), .B (n_2979), .C (n_15477), .Y (n_6779));
NOR2X1 g130814(.A (n_1731), .B (n_6389), .Y (n_6774));
NOR2X1 g130790(.A (n_1775), .B (n_6389), .Y (n_6773));
INVX1 g130978(.A (n_31495), .Y (n_24484));
BUFX3 g130219(.A (n_6770), .Y (n_7132));
CLKBUFX1 g130944(.A (n_6436), .Y (n_7250));
INVX1 g130696(.A (n_6979), .Y (n_12257));
NAND2X1 g129638(.A (n_6522), .B (n_33072), .Y (n_6767));
NAND2X1 g130143(.A (n_4308), .B (n_8407), .Y (n_8136));
NOR2X1 g130798(.A (n_3540), .B (n_12597), .Y (n_6765));
INVX1 g131025(.A (n_6421), .Y (n_12753));
INVX1 g131017(.A (n_6763), .Y (n_10490));
INVX1 g130985(.A (n_6787), .Y (n_31819));
INVX1 g130986(.A (n_6787), .Y (n_31876));
INVX4 g129766(.A (n_6844), .Y (n_7716));
INVX1 g129763(.A (n_6836), .Y (n_6762));
NAND2X1 g130412(.A (n_6748), .B (n_524), .Y (n_6761));
NAND2X1 g130369(.A (n_6752), .B (P2_reg1[15] ), .Y (n_32875));
NAND2X1 g130371(.A (n_6738), .B (P3_reg2[28] ), .Y (n_32069));
NAND2X1 g130505(.A (n_6754), .B (n_13699), .Y (n_6757));
NAND2X1 g130575(.A (n_6666), .B (P3_reg2[9] ), .Y (n_6756));
NAND2X1 g130527(.A (n_6754), .B (n_13351), .Y (n_6755));
NAND2X1 g130555(.A (n_6752), .B (P2_reg1[9] ), .Y (n_6753));
NAND2X1 g130553(.A (n_13727), .B (n_6621), .Y (n_6751));
NAND2X1 g130535(.A (n_6658), .B (P2_reg1[3] ), .Y (n_6750));
NAND2X1 g130577(.A (n_6748), .B (n_13692), .Y (n_35417));
NAND2X1 g130513(.A (n_6754), .B (P3_reg1[11] ), .Y (n_6747));
NAND2X1 g130499(.A (n_6744), .B (n_9165), .Y (n_35140));
NAND2X1 g130497(.A (n_6744), .B (P2_reg1[31] ), .Y (n_6745));
NAND2X1 g130488(.A (n_6596), .B (P2_reg1[5] ), .Y (n_6743));
NAND2X1 g129541(.A (n_32311), .B (n_3973), .Y (n_35143));
NAND2X1 g130453(.A (n_6690), .B (n_14133), .Y (n_6741));
NAND2X1 g130447(.A (n_6621), .B (n_13709), .Y (n_6740));
NAND2X1 g130445(.A (n_6738), .B (n_13511), .Y (n_6739));
INVX2 g129705(.A (n_6468), .Y (n_6829));
NAND2X1 g130348(.A (n_6429), .B (n_9590), .Y (n_6737));
NAND2X1 g130408(.A (n_6666), .B (n_13681), .Y (n_6736));
NAND2X1 g130405(.A (n_6661), .B (n_10610), .Y (n_6735));
NAND2X1 g130397(.A (n_6658), .B (P2_reg2[1] ), .Y (n_6734));
NAND2X1 g130327(.A (n_6744), .B (n_9088), .Y (n_32249));
NAND2X1 g130377(.A (n_6676), .B (n_13690), .Y (n_6732));
NAND2X1 g130373(.A (n_6661), .B (n_9142), .Y (n_6731));
NAND2X1 g130359(.A (n_6661), .B (n_10607), .Y (n_6730));
NAND2X1 g130347(.A (n_6754), .B (n_13377), .Y (n_6728));
NAND2X1 g130344(.A (n_6631), .B (n_9592), .Y (n_6727));
NAND2X1 g130335(.A (n_6703), .B (n_4160), .Y (n_6726));
NAND2X1 g129901(.A (n_3045), .B (n_6524), .Y (n_6725));
AND2X1 g129910(.A (n_6810), .B (n_6723), .Y (n_6724));
NAND2X1 g129911(.A (n_2807), .B (n_6524), .Y (n_6722));
NAND2X1 g129915(.A (n_3472), .B (n_6524), .Y (n_6721));
NAND2X1 g129919(.A (n_3334), .B (n_6524), .Y (n_6720));
NOR2X1 g129980(.A (n_4607), .B (n_6959), .Y (n_6718));
NAND2X1 g130000(.A (n_6419), .B (n_6416), .Y (n_32835));
NAND2X1 g130070(.A (n_3959), .B (n_6524), .Y (n_6716));
NOR2X1 g130076(.A (n_6837), .B (n_7353), .Y (n_7344));
NAND2X1 g130078(.A (n_35368), .B (n_6524), .Y (n_6715));
NAND2X1 g130079(.A (n_3869), .B (n_6524), .Y (n_6714));
NAND2X1 g130080(.A (n_4010), .B (n_6524), .Y (n_6712));
NAND2X2 g130158(.A (n_6379), .B (n_6343), .Y (n_6848));
CLKBUFX1 g130172(.A (n_7066), .Y (n_6990));
NAND2X2 g130253(.A (n_6362), .B (n_6341), .Y (n_6876));
NAND2X1 g130304(.A (n_6698), .B (n_9067), .Y (n_6708));
NAND2X1 g130305(.A (n_12389), .B (P3_reg2[18] ), .Y (n_6707));
NAND2X1 g130308(.A (n_6738), .B (n_13199), .Y (n_6706));
NAND2X1 g130309(.A (n_6703), .B (n_10452), .Y (n_6704));
NAND2X1 g129892(.A (n_2943), .B (n_6524), .Y (n_6702));
NAND2X1 g130316(.A (n_6658), .B (P2_reg_107), .Y (n_6701));
NAND2X1 g130320(.A (n_6698), .B (n_9794), .Y (n_35102));
NAND2X1 g130321(.A (n_6666), .B (n_13365), .Y (n_6697));
NAND2X1 g130323(.A (n_6661), .B (n_9178), .Y (n_6696));
NAND2X1 g130326(.A (n_6748), .B (n_13205), .Y (n_6695));
NAND2X1 g130337(.A (n_6752), .B (n_10363), .Y (n_6693));
NAND2X1 g130340(.A (n_6631), .B (n_10443), .Y (n_6692));
NAND2X1 g130342(.A (n_6690), .B (n_9595), .Y (n_35432));
NAND2X1 g130346(.A (n_6703), .B (P2_reg1[13] ), .Y (n_6689));
NAND2X1 g130350(.A (n_12389), .B (n_13679), .Y (n_6688));
NAND2X1 g130358(.A (n_6631), .B (P2_reg1[16] ), .Y (n_6687));
NAND2X1 g130364(.A (n_6608), .B (n_13215), .Y (n_6685));
NAND2X1 g130365(.A (n_6754), .B (P3_reg1[4] ), .Y (n_6684));
NAND2X1 g130306(.A (n_6698), .B (n_9139), .Y (n_6683));
NAND2X1 g130372(.A (n_6698), .B (n_9103), .Y (n_35263));
NAND2X1 g130314(.A (n_6752), .B (P2_reg_106), .Y (n_6681));
NAND2X1 g130375(.A (n_12389), .B (n_13354), .Y (n_6680));
NAND2X1 g130376(.A (n_6698), .B (P2_reg1[27] ), .Y (n_35146));
NAND2X1 g130378(.A (n_6676), .B (n_13695), .Y (n_6677));
NAND2X1 g130379(.A (n_6661), .B (n_9132), .Y (n_6675));
NAND2X1 g130380(.A (n_6621), .B (n_2718), .Y (n_6674));
NAND2X1 g130384(.A (n_12389), .B (n_13367), .Y (n_6672));
NAND2X1 g130386(.A (n_6658), .B (P2_reg1[8] ), .Y (n_6671));
NAND2X1 g130389(.A (n_6668), .B (P3_reg2[29] ), .Y (n_32073));
NAND2X1 g130390(.A (n_6668), .B (n_13330), .Y (n_32253));
NAND2X1 g130391(.A (n_6666), .B (n_13336), .Y (n_6667));
NAND2X1 g130396(.A (n_12389), .B (n_14168), .Y (n_6665));
NAND2X1 g130399(.A (n_6754), .B (n_13355), .Y (n_6664));
NAND2X1 g130402(.A (n_6666), .B (n_13352), .Y (n_35693));
NAND2X1 g130403(.A (n_6661), .B (n_10613), .Y (n_6662));
NAND2X1 g130406(.A (n_6744), .B (n_10043), .Y (n_35104));
NAND2X1 g130413(.A (n_6658), .B (P2_reg1[11] ), .Y (n_6659));
NAND2X1 g130414(.A (n_14096), .B (n_6631), .Y (n_6657));
NAND2X1 g130415(.A (n_6703), .B (n_13893), .Y (n_6656));
NAND2X1 g130417(.A (n_6429), .B (P2_reg2[11] ), .Y (n_6655));
NAND2X1 g130418(.A (n_6661), .B (n_3565), .Y (n_6653));
NAND2X1 g130311(.A (n_6661), .B (n_9135), .Y (n_6652));
NAND2X1 g130423(.A (n_6703), .B (n_4344), .Y (n_6651));
NAND2X1 g130424(.A (n_6748), .B (P3_reg2[15] ), .Y (n_6650));
NAND2X1 g130426(.A (n_6748), .B (n_13335), .Y (n_32092));
NAND2X1 g130428(.A (P3_reg2[30] ), .B (n_6754), .Y (n_6648));
NAND2X1 g130430(.A (n_6738), .B (n_13724), .Y (n_6647));
NAND2X1 g130431(.A (n_6658), .B (n_4475), .Y (n_6646));
NAND2X1 g130432(.A (n_6658), .B (P2_reg2[10] ), .Y (n_6645));
NAND2X1 g130434(.A (n_6661), .B (P2_reg1[21] ), .Y (n_6644));
NAND2X1 g130437(.A (n_6744), .B (n_9101), .Y (n_6643));
NAND2X1 g130440(.A (n_6752), .B (P2_reg2[29] ), .Y (n_32282));
NAND2X1 g130441(.A (n_6596), .B (n_3709), .Y (n_6641));
NAND2X1 g130450(.A (n_6703), .B (n_10563), .Y (n_6639));
NAND2X1 g130452(.A (n_14135), .B (n_6631), .Y (n_6638));
NAND2X1 g130454(.A (n_12389), .B (n_13353), .Y (n_6637));
NAND2X1 g130455(.A (n_6668), .B (n_13689), .Y (n_32167));
NAND2X1 g130456(.A (n_6668), .B (n_13200), .Y (n_6634));
NAND2X1 g130461(.A (n_6661), .B (n_9231), .Y (n_6630));
NAND2X1 g130462(.A (n_6690), .B (n_10653), .Y (n_6629));
NAND2X1 g130468(.A (n_6631), .B (P2_reg2[12] ), .Y (n_6628));
NAND2X1 g130470(.A (n_6698), .B (P2_reg1[20] ), .Y (n_32160));
NAND2X1 g130472(.A (n_6668), .B (n_13698), .Y (n_6626));
NAND2X1 g130473(.A (n_13645), .B (n_6631), .Y (n_6625));
NAND2X1 g130477(.A (n_6661), .B (n_10602), .Y (n_6624));
NAND2X1 g130478(.A (n_6429), .B (n_9549), .Y (n_6623));
NAND2X1 g130479(.A (n_6621), .B (n_13373), .Y (n_6622));
NAND2X1 g130482(.A (n_6621), .B (n_13341), .Y (n_6620));
NAND2X1 g130483(.A (n_6754), .B (P3_reg1[6] ), .Y (n_6619));
NAND2X1 g130485(.A (n_6754), .B (n_13683), .Y (n_6618));
NAND2X1 g130486(.A (n_6690), .B (n_9071), .Y (n_35430));
NAND2X1 g130487(.A (n_6748), .B (n_13697), .Y (n_6616));
NAND2X1 g130496(.A (n_6621), .B (n_13678), .Y (n_6615));
NAND2X1 g130353(.A (n_6429), .B (P2_reg1[12] ), .Y (n_6614));
NAND2X1 g130501(.A (n_6596), .B (P2_reg2[15] ), .Y (n_6613));
NAND2X1 g130502(.A (n_6748), .B (n_13206), .Y (n_6612));
NAND2X1 g130504(.A (n_6596), .B (P2_reg1[17] ), .Y (n_35282));
NAND2X1 g130508(.A (n_6608), .B (n_13343), .Y (n_35907));
NAND2X1 g130509(.A (n_6608), .B (n_13329), .Y (n_6607));
NAND2X1 g130515(.A (n_6596), .B (P2_reg1[4] ), .Y (n_6606));
NAND2X1 g130517(.A (n_6754), .B (P3_reg2[6] ), .Y (n_6605));
NAND2X1 g130518(.A (n_6631), .B (P2_reg1[23] ), .Y (n_6604));
NAND2X1 g130521(.A (n_6676), .B (n_13673), .Y (n_6603));
NAND2X1 g130525(.A (n_6666), .B (n_13209), .Y (n_6602));
NAND2X1 g130526(.A (n_6668), .B (n_13687), .Y (n_6601));
NAND2X1 g130528(.A (n_6676), .B (n_13213), .Y (n_6600));
NAND2X1 g130530(.A (n_6676), .B (n_13203), .Y (n_6599));
NAND2X1 g130533(.A (n_12389), .B (P3_reg2[10] ), .Y (n_6598));
NAND2X1 g130534(.A (n_6596), .B (P2_reg1[2] ), .Y (n_6597));
NAND2X1 g130536(.A (n_6666), .B (n_13202), .Y (n_6595));
NAND2X1 g130537(.A (n_6690), .B (n_9475), .Y (n_35138));
NAND2X1 g130539(.A (n_6666), .B (P3_reg1[18] ), .Y (n_6593));
NAND2X1 g130540(.A (n_6631), .B (n_4367), .Y (n_6592));
NAND2X1 g130542(.A (n_6666), .B (n_13204), .Y (n_6591));
NAND2X1 g130544(.A (n_6668), .B (n_13732), .Y (n_6589));
NAND2X1 g130545(.A (n_12389), .B (P3_reg1[1] ), .Y (n_6588));
NAND2X1 g130549(.A (n_6676), .B (n_13208), .Y (n_6587));
NAND2X1 g130551(.A (n_6744), .B (n_9097), .Y (n_6585));
NAND2X1 g130558(.A (n_6676), .B (n_13212), .Y (n_6584));
NAND2X1 g130559(.A (n_12389), .B (n_13680), .Y (n_6583));
NAND2X1 g130560(.A (n_6608), .B (n_13507), .Y (n_6582));
NAND2X1 g130562(.A (n_12389), .B (n_13366), .Y (n_6581));
NAND2X1 g130563(.A (n_6666), .B (n_13340), .Y (n_6579));
NAND2X1 g130565(.A (n_6658), .B (n_9586), .Y (n_6577));
NAND2X1 g130566(.A (n_6596), .B (P2_reg2[2] ), .Y (n_6576));
NAND2X1 g130570(.A (n_6596), .B (P2_reg1[18] ), .Y (n_6575));
NAND2X1 g130571(.A (n_6666), .B (n_13358), .Y (n_6574));
NAND2X1 g130574(.A (n_6608), .B (n_13211), .Y (n_6572));
NAND2X1 g130578(.A (n_12389), .B (P3_reg1[9] ), .Y (n_6571));
NAND2X1 g130580(.A (n_6666), .B (n_13348), .Y (n_6570));
NAND2X1 g130584(.A (n_6666), .B (n_13498), .Y (n_6568));
NAND2X1 g130585(.A (n_12389), .B (n_13721), .Y (n_6566));
NAND2X1 g130587(.A (n_6666), .B (n_13502), .Y (n_6565));
NAND2X1 g130589(.A (n_6738), .B (n_13216), .Y (n_6564));
NAND2X1 g130591(.A (n_6631), .B (n_3724), .Y (n_6563));
NAND2X1 g130593(.A (n_6429), .B (n_9565), .Y (n_6562));
NAND2X1 g130352(.A (n_6698), .B (n_9092), .Y (n_32264));
NAND2X1 g130438(.A (n_6621), .B (n_13337), .Y (n_6560));
XOR2X1 g130643(.A (n_5205), .B (n_6329), .Y (n_6559));
INVX1 g129587(.A (n_6425), .Y (n_6796));
AND2X1 g130095(.A (n_8060), .B (n_6347), .Y (n_6556));
INVX1 g130927(.A (n_8899), .Y (n_6901));
INVX1 g131001(.A (n_12917), .Y (n_6892));
INVX1 g131010(.A (n_12739), .Y (n_10342));
INVX1 g131073(.A (n_10465), .Y (n_31131));
NAND2X1 g130310(.A (n_6744), .B (P2_reg_104), .Y (n_6551));
NAND2X1 g130355(.A (n_6596), .B (P2_reg1[1] ), .Y (n_6550));
NAND2X1 g130330(.A (n_6738), .B (n_13368), .Y (n_6549));
NAND2X1 g130484(.A (n_6666), .B (P3_reg1[7] ), .Y (n_6548));
INVX1 g130928(.A (n_8899), .Y (n_6996));
INVX1 g130195(.A (n_6547), .Y (n_15622));
NAND2X1 g130360(.A (n_6752), .B (n_10435), .Y (n_6546));
NAND2X1 g130072(.A (n_4535), .B (n_6524), .Y (n_6545));
NOR2X1 g130056(.A (n_4182), .B (n_6959), .Y (n_6544));
NAND2X1 g130475(.A (n_6658), .B (n_4237), .Y (n_6541));
INVX1 g129521(.A (n_6835), .Y (n_6833));
NAND2X1 g130362(.A (n_6690), .B (n_9773), .Y (n_6540));
NAND2X1 g130572(.A (n_12389), .B (n_13359), .Y (n_6539));
NAND2X1 g129897(.A (n_3367), .B (n_6524), .Y (n_6538));
NAND2X1 g130476(.A (n_6748), .B (n_13207), .Y (n_6537));
NAND2X1 g130474(.A (n_6668), .B (P3_reg1[26] ), .Y (n_6534));
NAND2X2 g129523(.A (n_6408), .B (n_6304), .Y (n_6984));
NAND2X1 g130401(.A (n_6690), .B (n_10047), .Y (n_6532));
NAND2X1 g130363(.A (n_6752), .B (P2_reg1[19] ), .Y (n_32206));
NAND2X1 g130493(.A (n_6744), .B (n_9121), .Y (n_35413));
NAND2X1 g130425(.A (n_6631), .B (P2_reg2[9] ), .Y (n_6529));
NAND2X1 g130129(.A (n_3845), .B (n_6524), .Y (n_6528));
AOI21X1 g129886(.A0 (n_6527), .A1 (n_6404), .B0 (n_6405), .Y(n_6797));
NAND2X1 g130427(.A (n_6429), .B (P2_reg_95), .Y (n_6526));
NAND2X1 g129905(.A (n_2779), .B (n_6524), .Y (n_8741));
INVX1 g130707(.A (n_6979), .Y (n_6950));
CLKBUFX3 g130010(.A (n_34352), .Y (n_15576));
INVX1 g130091(.A (n_6522), .Y (n_7457));
NAND2X1 g130576(.A (n_12389), .B (n_13338), .Y (n_6521));
NAND2X1 g130385(.A (n_6631), .B (P2_reg1[6] ), .Y (n_6520));
CLKBUFX1 g130698(.A (n_6979), .Y (n_6938));
XOR2X1 g130631(.A (n_5214), .B (n_6330), .Y (n_6519));
NAND2X1 g130506(.A (n_6754), .B (n_13361), .Y (n_6518));
NAND2X1 g130564(.A (n_6698), .B (n_9599), .Y (n_6517));
INVX2 g129770(.A (n_6473), .Y (n_6844));
NAND2X1 g130503(.A (n_6754), .B (n_13342), .Y (n_6515));
NAND2X1 g130471(.A (n_6621), .B (P3_reg1[17] ), .Y (n_6514));
INVX1 g130954(.A (n_9909), .Y (n_6769));
NAND2X1 g130500(.A (n_12389), .B (P3_reg1[3] ), .Y (n_6512));
CLKBUFX1 g130979(.A (n_6806), .Y (n_31495));
NAND2X1 g130457(.A (n_6631), .B (P2_reg2[19] ), .Y (n_6511));
NAND2X1 g130524(.A (n_6621), .B (n_13357), .Y (n_6510));
INVX1 g130240(.A (n_7209), .Y (n_8113));
NAND2X1 g130367(.A (n_6703), .B (P2_reg1[22] ), .Y (n_32057));
NAND2X1 g130514(.A (n_12389), .B (n_13677), .Y (n_6506));
NAND2X1 g130561(.A (n_6666), .B (P3_reg2[13] ), .Y (n_6504));
NAND2X1 g130520(.A (n_6676), .B (n_13515), .Y (n_6503));
NAND2X1 g130351(.A (n_14513), .B (n_6754), .Y (n_6502));
NAND2X1 g130568(.A (n_6608), .B (n_14317), .Y (n_6501));
NAND2X1 g130543(.A (n_6690), .B (n_9597), .Y (n_6500));
NAND2X1 g130550(.A (n_6596), .B (P2_reg2[16] ), .Y (n_6499));
NAND2X1 g130546(.A (n_6596), .B (P2_reg2[8] ), .Y (n_6496));
INVX1 g130224(.A (n_6463), .Y (n_6770));
NAND3X1 g130802(.A (n_35012), .B (n_10601), .C (n_3185), .Y (n_6493));
INVX2 g129601(.A (n_6443), .Y (n_6800));
NAND2X1 g130519(.A (n_6703), .B (P2_reg2[18] ), .Y (n_6491));
INVX1 g130987(.A (n_6806), .Y (n_6787));
NAND2X1 g130349(.A (n_6754), .B (n_13332), .Y (n_6488));
NAND2X1 g130511(.A (n_6608), .B (n_13334), .Y (n_32158));
NAND2X1 g130590(.A (n_6738), .B (P3_reg1[16] ), .Y (n_6484));
NAND2X1 g130444(.A (n_6752), .B (P2_reg1[10] ), .Y (n_6483));
NAND2X1 g130436(.A (n_6738), .B (n_565), .Y (n_6482));
NAND2X1 g130416(.A (n_6596), .B (P2_reg2[3] ), .Y (n_6481));
XOR2X1 g130633(.A (n_6454), .B (n_6328), .Y (n_6480));
INVX1 g131070(.A (n_6437), .Y (n_31129));
INVX1 g131018(.A (n_6478), .Y (n_6763));
NAND2X1 g130411(.A (n_6608), .B (n_13344), .Y (n_6477));
NAND2X1 g130588(.A (n_6661), .B (P2_reg_108), .Y (n_35881));
CLKBUFX3 g129764(.A (n_6473), .Y (n_6836));
OR2X1 g130586(.A (n_6409), .B (n_127), .Y (n_6471));
NAND2X1 g129532(.A (n_34179), .B (n_6372), .Y (n_35144));
NAND2X1 g129534(.A (n_4315), .B (n_6345), .Y (n_6469));
NOR2X1 g129706(.A (n_34531), .B (n_34534), .Y (n_6468));
XOR2X1 g129887(.A (n_6467), .B (n_6406), .Y (n_6835));
NOR2X1 g130064(.A (n_8060), .B (n_6347), .Y (n_7346));
NAND2X1 g130092(.A (n_35651), .B (n_6296), .Y (n_6522));
INVX1 g130153(.A (n_34532), .Y (n_6466));
CLKBUFX1 g130197(.A (n_6464), .Y (n_15558));
NAND2X1 g130225(.A (n_6339), .B (n_6383), .Y (n_6463));
NAND2X1 g130251(.A (n_6306), .B (n_6268), .Y (n_6831));
INVX1 g130196(.A (n_6464), .Y (n_6547));
XOR2X1 g130641(.A (n_5306), .B (n_6282), .Y (n_6459));
INVX1 g130747(.A (n_6429), .Y (n_12464));
XOR2X1 g130838(.A (n_6454), .B (n_6275), .Y (n_6455));
XOR2X1 g130849(.A (n_4998), .B (n_6274), .Y (n_6453));
XOR2X1 g130850(.A (n_5218), .B (n_6273), .Y (n_6452));
INVX1 g130921(.A (n_6448), .Y (n_9382));
INVX1 g130923(.A (n_6448), .Y (n_8893));
INVX1 g130936(.A (n_30881), .Y (n_31881));
INVX1 g130937(.A (n_30881), .Y (n_31199));
INVX1 g130941(.A (n_30881), .Y (n_31734));
INVX1 g130990(.A (n_6447), .Y (n_30447));
INVX1 g130992(.A (n_6447), .Y (n_31639));
INVX1 g130996(.A (n_6447), .Y (n_31680));
INVX1 g131028(.A (n_6421), .Y (n_10736));
INVX1 g131059(.A (n_6446), .Y (n_12597));
INVX1 g131086(.A (n_6437), .Y (n_9937));
INVX1 g131090(.A (n_6437), .Y (n_30731));
CLKBUFX1 g130174(.A (n_6445), .Y (n_7066));
INVX1 g130241(.A (n_6524), .Y (n_7209));
INVX1 g130930(.A (n_9909), .Y (n_8916));
NAND2X1 g129602(.A (n_34393), .B (n_34595), .Y (n_6443));
INVX1 g130263(.A (n_6441), .Y (n_6495));
NAND2X1 g130018(.A (n_35651), .B (n_6439), .Y (n_33072));
INVX1 g130917(.A (n_6448), .Y (n_12664));
XOR2X1 g130628(.A (n_6334), .B (n_6269), .Y (n_6438));
INVX1 g130918(.A (n_6448), .Y (n_31713));
INVX1 g130940(.A (n_30881), .Y (n_30691));
INVX1 g131091(.A (n_6437), .Y (n_31422));
INVX1 g131063(.A (n_6446), .Y (n_12606));
INVX1 g130948(.A (n_6436), .Y (n_8933));
INVX8 g130723(.A (n_6435), .Y (n_6979));
INVX1 g130744(.A (n_6429), .Y (n_12488));
INVX1 g130976(.A (n_12755), .Y (n_6806));
INVX1 g130995(.A (n_6447), .Y (n_31019));
INVX1 g130920(.A (n_6448), .Y (n_30811));
INVX1 g131089(.A (n_6437), .Y (n_30893));
INVX4 g130243(.A (n_6524), .Y (n_6823));
NAND2X1 g129588(.A (n_34531), .B (n_34533), .Y (n_6425));
INVX1 g130991(.A (n_6447), .Y (n_31834));
INVX1 g131019(.A (n_6421), .Y (n_6478));
INVX1 g131080(.A (n_6446), .Y (n_10449));
INVX1 g130170(.A (n_6419), .Y (n_8409));
INVX1 g131088(.A (n_6437), .Y (n_31740));
INVX1 g131077(.A (n_31420), .Y (n_10465));
INVX1 g131011(.A (n_6421), .Y (n_12739));
INVX1 g130228(.A (n_6416), .Y (n_8407));
INVX1 g130154(.A (n_34532), .Y (n_6414));
INVX1 g130993(.A (n_6447), .Y (n_28332));
INVX1 g130994(.A (n_6447), .Y (n_30886));
INVX1 g130997(.A (n_6447), .Y (n_31299));
INVX1 g130999(.A (n_6354), .Y (n_12917));
INVX1 g130939(.A (n_30881), .Y (n_30527));
INVX1 g130938(.A (n_30881), .Y (n_31414));
AND2X1 g129771(.A (n_34595), .B (n_34582), .Y (n_6473));
INVX8 g130731(.A (n_6986), .Y (n_6435));
INVX1 g130677(.A (n_6409), .Y (n_6608));
INVX1 g130766(.A (n_6460), .Y (n_6690));
NAND2X1 g129524(.A (n_4026), .B (n_6293), .Y (n_6408));
NOR2X1 g129899(.A (n_6467), .B (n_6406), .Y (n_6407));
NOR2X1 g129916(.A (n_6527), .B (n_6404), .Y (n_6405));
NAND2X1 g130171(.A (n_35161), .B (n_6233), .Y (n_6419));
INVX1 g130254(.A (n_35652), .Y (n_6403));
INVX1 g130299(.A (n_34583), .Y (n_6402));
NOR2X1 g129923(.A (n_4188), .B (n_6404), .Y (n_6401));
XOR2X1 g130636(.A (n_5499), .B (n_6252), .Y (n_6400));
XOR2X1 g130637(.A (n_6359), .B (n_6220), .Y (n_6399));
XOR2X1 g130638(.A (n_6351), .B (n_6251), .Y (n_6398));
INVX1 g130666(.A (n_6409), .Y (n_6676));
INVX1 g130667(.A (n_6409), .Y (n_6738));
INVX1 g130671(.A (n_6409), .Y (n_6754));
INVX1 g130684(.A (n_6409), .Y (n_6621));
INVX1 g130767(.A (n_6460), .Y (n_6703));
XOR2X1 g130839(.A (n_6278), .B (n_6244), .Y (n_6396));
XOR2X1 g130841(.A (n_6394), .B (n_6243), .Y (n_6395));
XOR2X1 g130845(.A (n_6276), .B (n_6221), .Y (n_6393));
NAND2X1 g130899(.A (n_6297), .B (n_6132), .Y (n_6392));
CLKBUFX1 g130925(.A (n_9909), .Y (n_6448));
INVX1 g131029(.A (n_6354), .Y (n_6421));
INVX1 g131040(.A (n_34738), .Y (n_31122));
INVX1 g131044(.A (n_6349), .Y (n_10414));
INVX1 g131054(.A (n_34738), .Y (n_12601));
INVX1 g130270(.A (n_6387), .Y (n_6837));
NOR2X1 g130175(.A (n_35161), .B (n_6383), .Y (n_6445));
INVX2 g130198(.A (n_6365), .Y (n_6464));
INVX1 g130956(.A (n_9909), .Y (n_6436));
INVX1 g130679(.A (n_6409), .Y (n_6748));
XOR2X1 g130627(.A (n_6298), .B (n_6253), .Y (n_6382));
NAND2X1 g130164(.A (n_6378), .B (n_6284), .Y (n_6379));
XOR2X1 g130642(.A (n_6326), .B (n_6247), .Y (n_6377));
INVX1 g131035(.A (n_6349), .Y (n_9934));
NAND2X1 g129547(.A (n_6375), .B (n_6344), .Y (n_6376));
INVX1 g130680(.A (n_6409), .Y (n_6668));
CLKBUFX1 g130185(.A (n_6374), .Y (n_6959));
INVX1 g130163(.A (n_6372), .Y (n_32311));
INVX1 g130659(.A (n_12648), .Y (n_6371));
INVX1 g130676(.A (n_6409), .Y (n_12389));
XOR2X1 g129502(.A (n_4994), .B (n_6259), .Y (so[19]));
CLKBUFX1 g130942(.A (n_9909), .Y (n_30881));
INVX1 g130206(.A (n_6368), .Y (n_6856));
INVX1 g130678(.A (n_6409), .Y (n_6666));
INVX1 g130742(.A (n_6460), .Y (n_6429));
INVX1 g130187(.A (n_6365), .Y (n_15570));
INVX1 g131051(.A (n_6389), .Y (n_9928));
INVX1 g131056(.A (n_34738), .Y (n_12678));
INVX4 g130244(.A (n_6385), .Y (n_6524));
INVX1 g130762(.A (n_6460), .Y (n_6661));
INVX1 g130765(.A (n_6460), .Y (n_6698));
INVX1 g130772(.A (n_6460), .Y (n_6631));
NAND2X1 g130281(.A (n_32224), .B (n_6346), .Y (n_6362));
NOR2X1 g129530(.A (n_6355), .B (n_6353), .Y (n_6983));
INVX1 g131078(.A (n_34706), .Y (n_31420));
INVX1 g131065(.A (n_34706), .Y (n_6446));
XOR2X1 g131110(.A (n_6359), .B (n_6236), .Y (n_6360));
INVX1 g131099(.A (n_35007), .Y (n_12611));
INVX1 g131092(.A (n_35007), .Y (n_6437));
INVX1 g130255(.A (n_35652), .Y (n_6357));
NAND2X1 g129533(.A (n_6355), .B (n_6262), .Y (n_6356));
INVX1 g130758(.A (n_6460), .Y (n_6596));
INVX1 g130769(.A (n_6460), .Y (n_6658));
CLKBUFX1 g130998(.A (n_6354), .Y (n_6447));
INVX1 g130770(.A (n_6460), .Y (n_6744));
INVX1 g130768(.A (n_6460), .Y (n_6752));
NAND2X1 g130229(.A (n_35162), .B (n_6232), .Y (n_6416));
NAND2X1 g129545(.A (n_6355), .B (n_6353), .Y (n_6976));
XOR2X1 g130632(.A (n_6351), .B (n_6250), .Y (n_6352));
NOR2X1 g129529(.A (n_6355), .B (n_6262), .Y (n_6985));
INVX1 g131038(.A (n_35013), .Y (n_31307));
INVX1 g131046(.A (n_6349), .Y (n_9946));
XOR2X1 g130265(.A (n_6348), .B (n_6209), .Y (n_6441));
AND2X1 g130265_and(.A (n_6348), .B (n_6209), .Y (n_6723));
INVX1 g130859(.A (n_6347), .Y (n_7188));
NAND2X1 g130271(.A (n_34483), .B (n_6346), .Y (n_6372));
INVX1 g130162(.A (n_6344), .Y (n_6345));
NAND2X1 g130165(.A (n_6342), .B (n_6285), .Y (n_6343));
NAND2X2 g130199(.A (n_6309), .B (n_6310), .Y (n_6365));
NAND2X1 g130280(.A (n_3739), .B (n_34483), .Y (n_6341));
INVX1 g130290(.A (n_35162), .Y (n_6339));
XOR2X1 g130635(.A (n_6301), .B (n_6213), .Y (n_6338));
INVX1 g130655(.A (n_6439), .Y (n_6337));
NOR2X1 g130689(.A (n_12755), .B (n_349), .Y (n_6409));
NAND2X1 g130733(.A (n_6336), .B (n_35024), .Y (n_6986));
XOR2X1 g130836(.A (n_6334), .B (n_6201), .Y (n_6335));
XOR2X1 g130842(.A (n_4768), .B (n_6202), .Y (n_6333));
XOR2X1 g130851(.A (n_6270), .B (n_6206), .Y (n_6332));
MX2X1 g130853(.A (n_34485), .B (n_6324), .S0 (n_6323), .Y (n_6858));
XOR2X1 g130854(.A (n_6320), .B (n_6203), .Y (n_6331));
NAND3X1 g130873(.A (n_5730), .B (n_5551), .C (n_6196), .Y (n_6330));
NAND3X1 g130875(.A (n_5732), .B (n_5553), .C (n_6169), .Y (n_6329));
NAND2X1 g130900(.A (n_6242), .B (n_6193), .Y (n_6328));
INVX4 g130957(.A (n_8899), .Y (n_9909));
XOR2X1 g131104(.A (n_6326), .B (n_6195), .Y (n_6327));
XOR2X1 g130292(.A (n_32637), .B (n_6289), .Y (n_8060));
MX2X1 g130852(.A (n_6324), .B (n_34485), .S0 (n_6323), .Y (n_6860));
INVX1 g130869(.A (n_7393), .Y (n_6322));
NOR2X1 g130660(.A (n_6336), .B (P1_n_449), .Y (n_12648));
XOR2X1 g130856(.A (n_6320), .B (n_6175), .Y (n_6321));
INVX1 g130650(.A (n_6316), .Y (n_6798));
XOR2X1 g130846(.A (n_4903), .B (n_6164), .Y (n_6315));
XOR2X1 g130287(.A (n_6313), .B (n_6272), .Y (n_6387));
NAND2X1 g130186(.A (n_35952), .B (n_6311), .Y (n_6374));
NAND2X1 g130207(.A (n_6311), .B (n_6310), .Y (n_6368));
NAND2X2 g130248(.A (n_6309), .B (n_35653), .Y (n_6385));
NOR2X1 g130773(.A (n_35007), .B (P2_n_749), .Y (n_6460));
INVX1 g131048(.A (n_35012), .Y (n_6349));
NAND2X1 g130278(.A (n_6291), .B (n_6230), .Y (n_6306));
INVX1 g131052(.A (n_35012), .Y (n_6389));
NAND2X1 g129525(.A (n_6303), .B (n_6224), .Y (n_6304));
XOR2X1 g130640(.A (n_6301), .B (n_6191), .Y (n_6302));
XOR2X1 g130837(.A (n_6298), .B (n_6128), .Y (n_6299));
AOI21X1 g131167(.A0 (n_5806), .A1 (n_6131), .B0 (n_6199), .Y(n_6297));
INVX1 g130656(.A (n_6296), .Y (n_6439));
NAND2X1 g130272(.A (n_6292), .B (n_6178), .Y (n_6293));
NAND2X1 g130275(.A (n_6291), .B (n_35392), .Y (n_6344));
INVX1 g130297(.A (n_34534), .Y (n_6290));
NAND2X1 g130341(.A (n_32637), .B (n_6289), .Y (n_6404));
INVX1 g130648(.A (n_34483), .Y (n_32224));
INVX1 g130294(.A (n_6285), .Y (n_6286));
INVX1 g130293(.A (n_6285), .Y (n_6284));
MX2X1 g130835(.A (n_6188), .B (n_34119), .S0 (n_6153), .Y (n_6316));
INVX1 g130864(.A (n_6283), .Y (n_7353));
NAND3X1 g130876(.A (n_5402), .B (n_5308), .C (n_6142), .Y (n_6282));
AOI21X1 g130962(.A0 (n_6204), .A1 (n_6207), .B0 (n_6205), .Y(n_7393));
OAI21X1 g130965(.A0 (n_6281), .A1 (n_6210), .B0 (n_6177), .Y(n_6347));
XOR2X1 g131103(.A (n_5092), .B (n_6138), .Y (n_6280));
XOR2X1 g131106(.A (n_6278), .B (n_6140), .Y (n_6279));
XOR2X1 g131107(.A (n_6276), .B (n_6121), .Y (n_6277));
NAND4X1 g131132(.A (n_6130), .B (n_6133), .C (n_5925), .D (n_5942),.Y (n_6275));
NAND3X1 g131152(.A (n_6167), .B (n_5856), .C (n_4767), .Y (n_6274));
NAND3X1 g131154(.A (n_6198), .B (n_5858), .C (n_4595), .Y (n_6273));
NAND2X1 g130339(.A (n_4285), .B (n_6272), .Y (n_6406));
XOR2X1 g130855(.A (n_6270), .B (n_6157), .Y (n_6271));
NAND3X1 g130874(.A (n_6212), .B (n_6126), .C (n_5940), .Y (n_6269));
INVX1 g130958(.A (n_6336), .Y (n_8899));
NAND2X1 g130279(.A (n_4170), .B (n_35392), .Y (n_6268));
XOR2X1 g131109(.A (n_5087), .B (n_6139), .Y (n_6266));
XOR2X1 g131105(.A (n_5133), .B (n_6116), .Y (n_6265));
MX2X1 g130252(.A (n_3687), .B (n_6292), .S0 (n_35709), .Y (n_6355));
INVX1 g130653(.A (n_6262), .Y (n_6353));
NAND4X1 g130152(.A (n_6106), .B (n_6109), .C (n_5144), .D (n_5829),.Y (n_6259));
NAND2X1 g130277(.A (n_32242), .B (n_5067), .Y (n_6258));
INVX1 g130295(.A (n_6215), .Y (n_6285));
NAND3X1 g130877(.A (n_6112), .B (n_6080), .C (n_5951), .Y (n_6253));
NAND3X1 g130878(.A (n_5498), .B (n_5557), .C (n_6076), .Y (n_6252));
NAND3X1 g130884(.A (n_6249), .B (n_6057), .C (n_6248), .Y (n_6251));
NAND3X1 g130896(.A (n_6249), .B (n_6046), .C (n_6248), .Y (n_6250));
NAND2X1 g130898(.A (n_6158), .B (n_5600), .Y (n_6247));
XOR2X1 g130959(.A (n_6246), .B (n_6101), .Y (n_6336));
XOR2X1 g130961(.A (n_35188), .B (n_6211), .Y (n_6283));
NAND2X1 g130964(.A (n_6155), .B (n_6070), .Y (n_6310));
INVX4 g131032(.A (n_6354), .Y (n_12755));
OAI21X1 g131124(.A0 (n_6034), .A1 (n_6008), .B0 (n_6119), .Y(n_6244));
NAND4X1 g131133(.A (n_6081), .B (n_6090), .C (n_4934), .D (n_5830),.Y (n_6243));
AOI21X1 g131168(.A0 (n_5623), .A1 (n_6192), .B0 (n_6115), .Y(n_6242));
XOR2X1 g131176(.A (n_5494), .B (n_6197), .Y (n_6241));
XOR2X1 g131179(.A (n_5509), .B (n_6091), .Y (n_6240));
OAI21X1 g131181(.A0 (n_6144), .A1 (n_6143), .B0 (n_6145), .Y(n_6239));
XOR2X1 g131188(.A (n_5634), .B (n_6092), .Y (n_6238));
XOR2X1 g131191(.A (n_5392), .B (n_6166), .Y (n_6237));
NAND2X1 g131209(.A (n_6086), .B (n_6114), .Y (n_6236));
XOR2X1 g131260(.A (n_4880), .B (n_6087), .Y (n_6235));
XOR2X1 g131273(.A (n_5050), .B (n_6088), .Y (n_6234));
INVX1 g130861(.A (n_6232), .Y (n_6233));
MX2X1 g130289(.A (n_6231), .B (n_33173), .S0 (n_35156), .Y (n_6309));
INVX1 g130651(.A (n_35393), .Y (n_6230));
MX2X1 g130288(.A (n_33173), .B (n_6231), .S0 (n_35155), .Y (n_6311));
XOR2X1 g129889(.A (n_5145), .B (n_6110), .Y (so[18]));
INVX1 g130860(.A (n_6232), .Y (n_6383));
OAI21X1 g131185(.A0 (n_6147), .A1 (n_6146), .B0 (n_6148), .Y(n_6227));
XOR2X1 g129888(.A (n_4981), .B (n_6111), .Y (so[17]));
NOR2X1 g130273(.A (n_3687), .B (n_35709), .Y (n_6224));
XOR2X1 g131108(.A (n_5084), .B (n_6100), .Y (n_6222));
OAI21X1 g131138(.A0 (n_6036), .A1 (n_5935), .B0 (n_6141), .Y(n_6221));
NAND2X1 g130894(.A (n_6154), .B (n_5753), .Y (n_6220));
NAND2X1 g130847(.A (n_6113), .B (n_6085), .Y (n_6296));
NAND2X1 g130276(.A (n_4990), .B (n_35658), .Y (n_6218));
NAND2X1 g130775(.A (n_35452), .B (n_4656), .Y (n_6215));
MX2X1 g130848(.A (n_33176), .B (n_6214), .S0 (n_35387), .Y (n_6262));
NAND3X1 g130883(.A (n_6190), .B (n_5974), .C (n_6189), .Y (n_6213));
AOI21X1 g131113(.A0 (n_6026), .A1 (n_5637), .B0 (n_6052), .Y(n_6212));
NOR2X1 g131118(.A (n_35180), .B (n_6211), .Y (n_6272));
NOR2X1 g131119(.A (n_4396), .B (n_6210), .Y (n_6289));
NOR2X1 g131120(.A (n_6208), .B (n_6207), .Y (n_6209));
NAND2X1 g131129(.A (n_6156), .B (n_6083), .Y (n_6206));
NOR2X1 g131131(.A (n_6204), .B (n_6207), .Y (n_6205));
NAND2X1 g131141(.A (n_6174), .B (n_6099), .Y (n_6203));
NAND4X1 g131150(.A (n_6040), .B (n_6016), .C (n_5132), .D (n_5950),.Y (n_6202));
NAND3X1 g131157(.A (n_6078), .B (n_5941), .C (n_6125), .Y (n_6201));
XOR2X1 g131174(.A (n_4916), .B (n_6050), .Y (n_6200));
NAND3X1 g131203(.A (n_6017), .B (n_5864), .C (n_6022), .Y (n_6199));
NAND3X1 g131208(.A (n_6197), .B (n_5938), .C (n_5857), .Y (n_6198));
NAND3X1 g131210(.A (n_5571), .B (n_6172), .C (n_5591), .Y (n_6196));
NAND2X1 g131214(.A (n_6027), .B (n_6089), .Y (n_6195));
XOR2X1 g131272(.A (n_5031), .B (n_6168), .Y (n_6194));
NAND4X1 g131346(.A (n_5624), .B (n_5566), .C (n_5228), .D (n_6192),.Y (n_6193));
NAND3X1 g130886(.A (n_6190), .B (n_5973), .C (n_6189), .Y (n_6191));
INVX1 g131164(.A (n_34484), .Y (n_6323));
XOR2X1 g131173(.A (n_6150), .B (n_6049), .Y (n_6186));
XOR2X1 g131183(.A (n_6134), .B (n_6019), .Y (n_6185));
XOR2X1 g131170(.A (n_6102), .B (n_6003), .Y (n_6183));
XOR2X1 g131187(.A (n_5380), .B (n_6004), .Y (n_6182));
NAND2X1 g130960(.A (n_6105), .B (n_5988), .Y (n_6232));
INVX1 g130654(.A (n_35710), .Y (n_6178));
NAND2X1 g131135(.A (n_4256), .B (n_6210), .Y (n_6177));
XOR2X1 g130161(.A (n_5304), .B (n_6009), .Y (so[16]));
NAND3X1 g131126(.A (n_6174), .B (n_6039), .C (n_5245), .Y (n_6175));
XOR2X1 g131259(.A (n_5186), .B (n_6172), .Y (n_6173));
XOR2X1 g131033(.A (n_6170), .B (n_5997), .Y (n_6354));
NAND3X1 g131221(.A (n_5489), .B (n_6168), .C (n_5552), .Y (n_6169));
NAND3X1 g131211(.A (n_6166), .B (n_5948), .C (n_5855), .Y (n_6167));
XOR2X1 g131180(.A (n_6117), .B (n_6020), .Y (n_6165));
NAND4X1 g131149(.A (n_6011), .B (n_6042), .C (n_5091), .D (n_5945),.Y (n_6164));
INVX1 g130657(.A (n_35657), .Y (n_32242));
NAND2X1 g130594(.A (n_6107), .B (n_35105), .Y (n_32289));
NAND2X1 g130664(.A (n_6180), .B (n_6179), .Y (n_6160));
AOI21X1 g131160(.A0 (n_5978), .A1 (n_5060), .B0 (n_5422), .Y(n_6158));
NAND3X1 g131134(.A (n_6156), .B (n_5898), .C (n_5247), .Y (n_6157));
NAND2X1 g131146(.A (n_5161), .B (n_6054), .Y (n_6155));
AOI21X1 g131161(.A0 (n_5980), .A1 (n_5048), .B0 (n_5658), .Y(n_6154));
INVX1 g131162(.A (n_34574), .Y (n_6153));
XOR2X1 g131171(.A (n_6150), .B (n_6077), .Y (n_6151));
XOR2X1 g131186(.A (n_4874), .B (n_5910), .Y (n_6149));
NAND2X1 g131206(.A (n_6147), .B (n_6146), .Y (n_6148));
NAND2X1 g131217(.A (n_6144), .B (n_6143), .Y (n_6145));
NAND3X1 g131226(.A (n_5479), .B (n_6136), .C (n_5420), .Y (n_6142));
AOI21X1 g131228(.A0 (n_5953), .A1 (n_5721), .B0 (n_5751), .Y(n_6141));
NAND3X1 g131233(.A (n_5909), .B (n_5930), .C (n_5706), .Y (n_6140));
NAND3X1 g131241(.A (n_5964), .B (n_5931), .C (n_5537), .Y (n_6139));
NAND3X1 g131244(.A (n_6030), .B (n_5939), .C (n_5646), .Y (n_6138));
XOR2X1 g131264(.A (n_4988), .B (n_6136), .Y (n_6137));
XOR2X1 g131271(.A (n_6134), .B (n_5965), .Y (n_6135));
NAND2X1 g131313(.A (n_6002), .B (n_5521), .Y (n_6133));
NAND4X1 g131345(.A (n_5807), .B (n_5564), .C (n_5439), .D (n_6131),.Y (n_6132));
AOI21X1 g131350(.A0 (n_6047), .A1 (n_5850), .B0 (n_6028), .Y(n_6130));
XOR2X1 g130257(.A (n_5177), .B (n_5991), .Y (so[15]));
NAND3X1 g131158(.A (n_5994), .B (n_5952), .C (n_6079), .Y (n_6128));
XOR2X1 g131177(.A (n_5336), .B (n_5896), .Y (n_6127));
NAND2X1 g131314(.A (n_6018), .B (n_6125), .Y (n_6126));
XOR2X1 g131184(.A (n_4908), .B (n_5981), .Y (n_6124));
XOR2X1 g131190(.A (n_4910), .B (n_5982), .Y (n_6123));
XOR2X1 g131261(.A (n_4712), .B (n_5916), .Y (n_6122));
NAND3X1 g131236(.A (n_5904), .B (n_5944), .C (n_5698), .Y (n_6121));
XOR2X1 g131276(.A (n_4730), .B (n_5958), .Y (n_6120));
AOI21X1 g131227(.A0 (n_5954), .A1 (n_5819), .B0 (n_5847), .Y(n_6119));
XOR2X1 g131269(.A (n_6117), .B (n_5901), .Y (n_6118));
NAND3X1 g131242(.A (n_6007), .B (n_5949), .C (n_5642), .Y (n_6116));
NAND3X1 g131220(.A (n_5946), .B (n_5959), .C (n_5927), .Y (n_6115));
AOI21X1 g131325(.A0 (n_5912), .A1 (n_5611), .B0 (n_5926), .Y(n_6114));
NAND2X1 g130879(.A (n_34915), .B (n_6056), .Y (n_6113));
AOI21X1 g131114(.A0 (n_5895), .A1 (n_5655), .B0 (n_6012), .Y(n_6112));
NAND3X1 g130249(.A (n_5891), .B (n_5890), .C (n_5682), .Y (n_6111));
NAND4X1 g130250(.A (n_5892), .B (n_4980), .C (n_5791), .D (n_5797),.Y (n_6110));
AOI21X1 g130283(.A0 (n_5990), .A1 (n_5793), .B0 (n_5989), .Y(n_6109));
INVX1 g130862(.A (n_6107), .Y (n_32889));
NAND3X1 g130274(.A (n_5586), .B (n_5888), .C (n_5585), .Y (n_6106));
NAND2X1 g131123(.A (n_6055), .B (n_5986), .Y (n_6105));
XOR2X1 g131169(.A (n_6102), .B (n_5993), .Y (n_6103));
NOR2X1 g131219(.A (n_5969), .B (n_6059), .Y (n_6101));
NOR2X1 g131231(.A (n_5921), .B (n_5996), .Y (n_6210));
NOR2X1 g131234(.A (n_5782), .B (n_5917), .Y (n_6248));
NAND3X1 g131243(.A (n_5924), .B (n_5886), .C (n_5506), .Y (n_6100));
AOI21X1 g131246(.A0 (n_6097), .A1 (n_6038), .B0 (n_5244), .Y(n_6099));
XOR2X1 g131254(.A (n_4962), .B (n_6097), .Y (n_6098));
XOR2X1 g131255(.A (n_4428), .B (n_5818), .Y (n_6096));
XOR2X1 g131262(.A (n_6023), .B (n_5826), .Y (n_6095));
OAI21X1 g131267(.A0 (n_5977), .A1 (n_6071), .B0 (n_5975), .Y(n_6094));
XOR2X1 g131275(.A (n_5047), .B (n_6075), .Y (n_6093));
OAI21X1 g131278(.A0 (n_5841), .A1 (n_5762), .B0 (n_5786), .Y(n_6092));
OAI21X1 g131284(.A0 (n_5842), .A1 (n_5759), .B0 (n_5779), .Y(n_6091));
NAND2X1 g131296(.A (n_5962), .B (n_5703), .Y (n_6166));
NAND2X1 g131319(.A (n_5960), .B (n_5459), .Y (n_6090));
AOI21X1 g131324(.A0 (n_5845), .A1 (n_5608), .B0 (n_6021), .Y(n_6089));
OAI21X1 g131381(.A0 (n_5837), .A1 (n_5747), .B0 (n_5719), .Y(n_6088));
OAI21X1 g131382(.A0 (n_5836), .A1 (n_5766), .B0 (n_5710), .Y(n_6087));
AOI21X1 g131478(.A0 (n_5332), .A1 (n_5738), .B0 (n_5936), .Y(n_6086));
NAND2X1 g130881(.A (n_34913), .B (n_34924), .Y (n_6085));
AOI21X1 g131245(.A0 (n_6065), .A1 (n_5897), .B0 (n_5246), .Y(n_6083));
AOI21X1 g131354(.A0 (n_6048), .A1 (n_5750), .B0 (n_5906), .Y(n_6081));
NAND2X1 g131316(.A (n_5947), .B (n_6079), .Y (n_6080));
OR2X1 g131196(.A (n_5652), .B (n_6077), .Y (n_6078));
NAND2X1 g131298(.A (n_5934), .B (n_5742), .Y (n_6197));
NAND3X1 g131205(.A (n_5563), .B (n_6075), .C (n_5555), .Y (n_6076));
XOR2X1 g131172(.A (n_6143), .B (n_5883), .Y (n_6074));
XOR2X1 g131362(.A (n_4540), .B (n_6006), .Y (n_6073));
XOR2X1 g131257(.A (n_6071), .B (n_5823), .Y (n_6072));
NAND2X1 g131147(.A (n_6069), .B (n_6053), .Y (n_6070));
XOR2X1 g131361(.A (n_4549), .B (n_6029), .Y (n_6068));
AOI21X1 g131230(.A0 (n_5821), .A1 (n_4688), .B0 (n_6060), .Y(n_6211));
OAI21X1 g131274(.A0 (n_5979), .A1 (n_5998), .B0 (n_5976), .Y(n_6067));
XOR2X1 g131270(.A (n_4960), .B (n_6065), .Y (n_6066));
OAI21X1 g131277(.A0 (n_5918), .A1 (n_6062), .B0 (n_5919), .Y(n_6064));
XOR2X1 g131263(.A (n_6062), .B (n_5828), .Y (n_6063));
NOR2X1 g131223(.A (n_5967), .B (n_6060), .Y (n_6061));
AOI21X1 g131215(.A0 (n_5862), .A1 (n_33250), .B0 (n_6059), .Y(n_6207));
XOR2X1 g131178(.A (n_6146), .B (n_5882), .Y (n_6058));
NAND3X1 g131326(.A (n_6044), .B (n_6045), .C (n_6043), .Y (n_6057));
INVX1 g131127(.A (n_34924), .Y (n_6056));
NAND2X2 g131137(.A (n_35158), .B (n_6055), .Y (n_6107));
INVX1 g131198(.A (n_6053), .Y (n_6054));
AOI21X1 g131237(.A0 (n_5717), .A1 (n_5839), .B0 (n_6025), .Y(n_6052));
NOR2X1 g131239(.A (n_5705), .B (n_5879), .Y (n_6189));
XOR2X1 g131266(.A (n_5712), .B (n_5700), .Y (n_6051));
OAI21X1 g131285(.A0 (n_5739), .A1 (n_5673), .B0 (n_5704), .Y(n_6050));
NOR2X1 g131289(.A (n_5774), .B (n_5840), .Y (n_6049));
AOI21X1 g131290(.A0 (n_5805), .A1 (n_5749), .B0 (n_6048), .Y(n_6144));
AOI21X1 g131291(.A0 (n_5761), .A1 (n_5849), .B0 (n_6047), .Y(n_6147));
NAND3X1 g131302(.A (n_6045), .B (n_6044), .C (n_6043), .Y (n_6046));
NAND3X1 g131305(.A (n_5957), .B (n_5956), .C (n_6010), .Y (n_6042));
XOR2X1 g130286(.A (n_5147), .B (n_5804), .Y (so[14]));
AOI21X1 g131352(.A0 (n_5913), .A1 (n_6015), .B0 (n_5780), .Y(n_6040));
AOI22X1 g131356(.A0 (n_5812), .A1 (n_6038), .B0 (n_5811), .B1(n_6038), .Y (n_6039));
OAI21X1 g131374(.A0 (n_6036), .A1 (n_5870), .B0 (n_5817), .Y(n_6037));
OAI21X1 g131375(.A0 (n_6034), .A1 (n_5867), .B0 (n_5865), .Y(n_6035));
XOR2X1 g131376(.A (n_4373), .B (n_5923), .Y (n_6033));
XOR2X1 g131377(.A (n_5062), .B (n_5961), .Y (n_6032));
XOR2X1 g131378(.A (n_4542), .B (n_5963), .Y (n_6031));
OR2X1 g131392(.A (n_5748), .B (n_6029), .Y (n_6030));
NAND2X1 g131406(.A (n_5854), .B (n_5408), .Y (n_6172));
NOR2X1 g131407(.A (n_5824), .B (n_6001), .Y (n_6028));
AOI21X1 g131484(.A0 (n_5569), .A1 (n_5663), .B0 (n_5834), .Y(n_6027));
NOR2X1 g131540(.A (n_4955), .B (n_6025), .Y (n_6026));
OAI21X1 g131265(.A0 (n_5877), .A1 (n_6023), .B0 (n_5878), .Y(n_6024));
AOI22X1 g131476(.A0 (n_6021), .A1 (n_5662), .B0 (n_4934), .B1(n_5514), .Y (n_6022));
AOI21X1 g131318(.A0 (n_5746), .A1 (n_5902), .B0 (n_5943), .Y(n_6020));
AOI21X1 g131312(.A0 (n_5745), .A1 (n_5907), .B0 (n_5929), .Y(n_6019));
NAND2X1 g131471(.A (n_5848), .B (n_6017), .Y (n_6018));
NAND3X1 g131306(.A (n_5915), .B (n_5914), .C (n_6015), .Y (n_6016));
XOR2X1 g130285(.A (n_4873), .B (n_5801), .Y (so[13]));
XOR2X1 g130284(.A (n_4793), .B (n_5809), .Y (so[11]));
AOI21X1 g131235(.A0 (n_5692), .A1 (n_5843), .B0 (n_5894), .Y(n_6012));
AOI21X1 g131351(.A0 (n_5955), .A1 (n_6010), .B0 (n_5787), .Y(n_6011));
NAND3X1 g130282(.A (n_5794), .B (n_5715), .C (n_5588), .Y (n_6009));
OR2X1 g131608(.A (n_5813), .B (n_5743), .Y (n_6008));
OR2X1 g131386(.A (n_5767), .B (n_6006), .Y (n_6007));
XOR2X1 g131249(.A (n_4588), .B (n_5776), .Y (n_6005));
OAI21X1 g131281(.A0 (n_5726), .A1 (n_5604), .B0 (n_5783), .Y(n_6004));
NOR2X1 g131283(.A (n_5723), .B (n_5844), .Y (n_6003));
NOR2X1 g131399(.A (n_5825), .B (n_6001), .Y (n_6002));
XOR2X1 g131256(.A (n_5872), .B (n_5785), .Y (n_6000));
NAND2X2 g131111(.A (n_35296), .B (n_35295), .Y (n_6179));
XOR2X1 g131253(.A (n_5998), .B (n_5773), .Y (n_5999));
NOR2X1 g131216(.A (n_5875), .B (n_5996), .Y (n_5997));
INVX1 g131199(.A (n_6053), .Y (n_5995));
OR2X1 g131197(.A (n_5661), .B (n_5993), .Y (n_5994));
XOR2X1 g131363(.A (n_5202), .B (n_5933), .Y (n_5992));
NAND2X1 g131435(.A (n_5852), .B (n_5288), .Y (n_6168));
AOI21X1 g130302(.A0 (n_5681), .A1 (n_5792), .B0 (n_5990), .Y(n_5991));
NOR2X1 g130464(.A (n_5808), .B (n_5887), .Y (n_5989));
NAND3X1 g131125(.A (n_33586), .B (n_35301), .C (n_4688), .Y (n_5988));
INVX1 g131193(.A (n_35157), .Y (n_5986));
INVX1 g131201(.A (n_5922), .Y (n_35082));
NAND2X1 g131229(.A (n_5789), .B (n_4688), .Y (n_35275));
OAI21X1 g131279(.A0 (n_5667), .A1 (n_5757), .B0 (n_5781), .Y(n_5982));
OAI21X1 g131288(.A0 (n_5616), .A1 (n_5632), .B0 (n_5626), .Y(n_5981));
NOR2X1 g131294(.A (n_5979), .B (n_5657), .Y (n_5980));
NOR2X1 g131303(.A (n_5977), .B (n_5469), .Y (n_5978));
NAND2X1 g131310(.A (n_5979), .B (n_5998), .Y (n_5976));
NAND2X1 g131311(.A (n_5977), .B (n_6071), .Y (n_5975));
NAND3X1 g131321(.A (n_5971), .B (n_5972), .C (n_5970), .Y (n_5974));
NAND3X1 g131327(.A (n_5972), .B (n_5971), .C (n_5970), .Y (n_5973));
AOI21X1 g131329(.A0 (n_5671), .A1 (n_5293), .B0 (n_5577), .Y(n_6077));
AOI21X1 g131353(.A0 (n_5536), .A1 (n_5548), .B0 (n_5778), .Y(n_6174));
AOI21X1 g131355(.A0 (n_5615), .A1 (n_5861), .B0 (n_4901), .Y(n_5969));
AOI21X1 g131359(.A0 (n_5677), .A1 (n_5820), .B0 (n_34947), .Y(n_5967));
NOR2X1 g131380(.A (n_5744), .B (n_5735), .Y (n_5965));
OR2X1 g131390(.A (n_5697), .B (n_5963), .Y (n_5964));
NAND3X1 g131403(.A (n_5961), .B (n_5541), .C (n_5702), .Y (n_5962));
NAND2X1 g131404(.A (n_5756), .B (n_5416), .Y (n_6136));
NAND2X1 g131411(.A (n_5775), .B (n_6043), .Y (n_6249));
NOR2X1 g131421(.A (n_3393), .B (n_5905), .Y (n_5960));
OR2X1 g131424(.A (n_5880), .B (n_5932), .Y (n_5959));
AOI21X1 g131453(.A0 (n_5957), .A1 (n_5956), .B0 (n_5955), .Y(n_5958));
OAI21X1 g131460(.A0 (n_5734), .A1 (n_5150), .B0 (n_5727), .Y(n_5954));
OAI21X1 g131461(.A0 (n_5736), .A1 (n_5210), .B0 (n_5693), .Y(n_5953));
AOI21X1 g131463(.A0 (n_5234), .A1 (n_5951), .B0 (n_5699), .Y(n_5952));
AOI22X1 g131464(.A0 (n_5731), .A1 (n_5547), .B0 (n_5204), .B1(n_5131), .Y (n_5950));
AOI21X1 g131468(.A0 (n_5701), .A1 (n_5948), .B0 (n_5711), .Y(n_5949));
NAND2X1 g131469(.A (n_5752), .B (n_5946), .Y (n_5947));
AOI22X1 g131472(.A0 (n_5729), .A1 (n_5590), .B0 (n_5213), .B1(n_5090), .Y (n_5945));
AOI21X1 g131473(.A0 (n_5943), .A1 (n_5903), .B0 (n_5649), .Y(n_5944));
AOI21X1 g131474(.A0 (n_5539), .A1 (n_5946), .B0 (n_5754), .Y(n_5942));
AOI21X1 g131475(.A0 (n_4923), .A1 (n_5940), .B0 (n_5707), .Y(n_5941));
AOI21X1 g131485(.A0 (n_5740), .A1 (n_5938), .B0 (n_5720), .Y(n_5939));
XOR2X1 g131492(.A (n_4790), .B (n_5851), .Y (n_5937));
NOR2X1 g131549(.A (n_5772), .B (n_5911), .Y (n_5936));
OR2X1 g131634(.A (n_5722), .B (n_5668), .Y (n_5935));
NAND3X1 g131422(.A (n_5933), .B (n_5543), .C (n_5741), .Y (n_5934));
NOR2X1 g131561(.A (n_5932), .B (n_5881), .Y (n_6192));
AOI21X1 g131470(.A0 (n_5457), .A1 (n_5549), .B0 (n_5688), .Y(n_5931));
AOI21X1 g131481(.A0 (n_5929), .A1 (n_5908), .B0 (n_5656), .Y(n_5930));
XOR2X1 g131189(.A (n_1078), .B (n_5680), .Y (n_5928));
AOI22X1 g131465(.A0 (n_5926), .A1 (n_5708), .B0 (n_5925), .B1(n_5341), .Y (n_5927));
OR2X1 g131389(.A (n_5633), .B (n_5923), .Y (n_5924));
INVX1 g131200(.A (n_5922), .Y (n_6053));
AND2X1 g131344(.A (n_5725), .B (n_5219), .Y (n_5921));
XOR2X1 g131491(.A (n_4721), .B (n_5853), .Y (n_5920));
NAND2X1 g131299(.A (n_5918), .B (n_6062), .Y (n_5919));
NAND2X1 g131295(.A (n_5685), .B (n_5085), .Y (n_5917));
AOI21X1 g131444(.A0 (n_5915), .A1 (n_5914), .B0 (n_5913), .Y(n_5916));
AOI21X1 g131349(.A0 (n_5505), .A1 (n_5417), .B0 (n_5784), .Y(n_6156));
NOR2X1 g131581(.A (n_5180), .B (n_5911), .Y (n_5912));
OAI21X1 g131282(.A0 (n_5621), .A1 (n_5696), .B0 (n_5687), .Y(n_5910));
NAND3X1 g131420(.A (n_5866), .B (n_5908), .C (n_5907), .Y (n_5909));
NOR2X1 g131412(.A (n_5827), .B (n_5905), .Y (n_5906));
NAND3X1 g131405(.A (n_5869), .B (n_5903), .C (n_5902), .Y (n_5904));
NOR2X1 g131379(.A (n_5669), .B (n_5737), .Y (n_5901));
AOI22X1 g131357(.A0 (n_5860), .A1 (n_5897), .B0 (n_5859), .B1(n_5897), .Y (n_5898));
OAI21X1 g131286(.A0 (n_5620), .A1 (n_5765), .B0 (n_5777), .Y(n_5896));
NOR2X1 g131579(.A (n_5101), .B (n_5894), .Y (n_5895));
XOR2X1 g131175(.A (n_1354), .B (n_5607), .Y (n_5893));
NAND3X1 g130597(.A (n_5803), .B (n_5795), .C (n_5802), .Y (n_5892));
NAND3X1 g130596(.A (n_5800), .B (n_5889), .C (n_5799), .Y (n_5891));
AOI21X1 g130622(.A0 (n_5798), .A1 (n_5889), .B0 (n_5454), .Y(n_5890));
INVX1 g130691(.A (n_5887), .Y (n_5888));
AOI21X1 g131480(.A0 (n_5568), .A1 (n_5418), .B0 (n_5627), .Y(n_5886));
OAI21X1 g131144(.A0 (n_33170), .A1 (n_5105), .B0 (n_4502), .Y(n_35296));
OAI21X1 g131280(.A0 (n_5565), .A1 (n_5815), .B0 (n_5863), .Y(n_5883));
OAI21X1 g131287(.A0 (n_5567), .A1 (n_5881), .B0 (n_5880), .Y(n_5882));
NAND2X1 g131297(.A (n_5678), .B (n_5129), .Y (n_5879));
NAND2X1 g131317(.A (n_5877), .B (n_6023), .Y (n_5878));
AOI21X1 g131330(.A0 (n_5481), .A1 (n_5389), .B0 (n_5581), .Y(n_5993));
AOI21X1 g131358(.A0 (n_5463), .A1 (n_5724), .B0 (n_5874), .Y(n_5875));
XOR2X1 g131366(.A (n_5872), .B (n_5670), .Y (n_5873));
XOR2X1 g131371(.A (n_5870), .B (n_5869), .Y (n_5871));
XOR2X1 g131372(.A (n_5867), .B (n_5866), .Y (n_5868));
NAND2X1 g131409(.A (n_6034), .B (n_5867), .Y (n_5865));
OR2X1 g131415(.A (n_5863), .B (n_5816), .Y (n_5864));
NAND2X1 g131419(.A (n_5675), .B (n_5861), .Y (n_5862));
NAND2X1 g131430(.A (n_5618), .B (n_5413), .Y (n_6075));
OR2X1 g131437(.A (n_5860), .B (n_5859), .Y (n_6065));
AOI21X1 g131477(.A0 (n_5645), .A1 (n_5857), .B0 (n_5001), .Y(n_5858));
AOI21X1 g131483(.A0 (n_5641), .A1 (n_5855), .B0 (n_5082), .Y(n_5856));
NAND3X1 g131534(.A (n_5853), .B (n_5406), .C (n_5491), .Y (n_5854));
NAND3X1 g131537(.A (n_5851), .B (n_5286), .C (n_5544), .Y (n_5852));
NAND2X1 g131551(.A (n_5850), .B (n_5849), .Y (n_6001));
NAND2X1 g131574(.A (n_5847), .B (n_4934), .Y (n_5848));
NOR2X1 g131578(.A (n_5385), .B (n_5833), .Y (n_5845));
INVX1 g131614(.A (n_5843), .Y (n_5844));
AND2X1 g131616(.A (n_5602), .B (n_5695), .Y (n_5842));
AND2X1 g131630(.A (n_5639), .B (n_5768), .Y (n_5841));
INVX1 g131638(.A (n_5839), .Y (n_5840));
AND2X1 g131799(.A (n_5640), .B (n_5664), .Y (n_5837));
AND2X1 g131817(.A (n_5638), .B (n_5630), .Y (n_5836));
XOR2X1 g130630(.A (n_5017), .B (n_5504), .Y (so[12]));
NOR2X1 g131541(.A (n_5822), .B (n_5833), .Y (n_5834));
AOI21X1 g131648(.A0 (n_2313), .A1 (n_5516), .B0 (n_5631), .Y(n_6006));
XOR2X1 g131493(.A (n_4707), .B (n_5755), .Y (n_5832));
AOI21X1 g131644(.A0 (n_2674), .A1 (n_5512), .B0 (n_5665), .Y(n_6029));
XOR2X1 g130843(.A (n_1329), .B (n_5452), .Y (n_5831));
AOI21X1 g131467(.A0 (n_5644), .A1 (n_6017), .B0 (n_5601), .Y(n_5830));
AOI21X1 g130621(.A0 (n_4818), .A1 (n_5149), .B0 (n_5683), .Y(n_5829));
OAI21X1 g131393(.A0 (n_5460), .A1 (n_3393), .B0 (n_5827), .Y(n_5828));
OAI21X1 g131387(.A0 (n_5522), .A1 (n_5825), .B0 (n_5824), .Y(n_5826));
NAND2X1 g131455(.A (n_5597), .B (n_5822), .Y (n_5823));
NAND2X1 g131446(.A (n_5599), .B (n_5820), .Y (n_5821));
NAND3X1 g131750(.A (n_5819), .B (n_6125), .C (n_4934), .Y (n_6025));
AOI21X1 g131443(.A0 (n_5971), .A1 (n_5972), .B0 (n_5814), .Y(n_5818));
NAND2X1 g131438(.A (n_6036), .B (n_5870), .Y (n_5817));
NOR2X1 g131587(.A (n_5816), .B (n_5815), .Y (n_6131));
NAND2X1 g131434(.A (n_5814), .B (n_5970), .Y (n_6190));
NAND2X1 g131726(.A (n_5819), .B (n_5327), .Y (n_5813));
OR2X1 g131431(.A (n_5812), .B (n_5811), .Y (n_6097));
OAI21X1 g131143(.A0 (n_33582), .A1 (n_5258), .B0 (n_4688), .Y(n_35274));
NAND2X1 g131202(.A (n_5629), .B (n_33250), .Y (n_5922));
NAND2X1 g130829(.A (n_5587), .B (n_5808), .Y (n_5809));
AOI21X1 g131395(.A0 (n_5440), .A1 (n_5807), .B0 (n_5806), .Y(n_5918));
OR2X1 g131559(.A (n_5474), .B (n_5487), .Y (n_5805));
AOI21X1 g130661(.A0 (n_5803), .A1 (n_5802), .B0 (n_5796), .Y(n_5804));
AOI21X1 g130662(.A0 (n_5800), .A1 (n_5799), .B0 (n_5798), .Y(n_5801));
NAND2X1 g130663(.A (n_5796), .B (n_5795), .Y (n_5797));
NAND3X1 g130665(.A (n_5503), .B (n_5714), .C (n_5502), .Y (n_5794));
NAND2X1 g130692(.A (n_5793), .B (n_5792), .Y (n_5887));
AOI21X1 g130833(.A0 (n_5437), .A1 (n_5272), .B0 (n_5589), .Y(n_5791));
XOR2X1 g131182(.A (n_1260), .B (n_5281), .Y (n_5790));
NAND2X1 g131339(.A (n_5582), .B (n_4591), .Y (n_5789));
NOR2X1 g131396(.A (n_5786), .B (n_5763), .Y (n_5787));
AOI21X1 g131418(.A0 (n_4127), .A1 (n_5636), .B0 (n_5716), .Y(n_5785));
NOR2X1 g131423(.A (n_5783), .B (n_5603), .Y (n_5784));
NOR2X1 g131429(.A (n_5781), .B (n_5758), .Y (n_5782));
NOR2X1 g131433(.A (n_5779), .B (n_5760), .Y (n_5780));
NOR2X1 g131436(.A (n_5777), .B (n_5764), .Y (n_5778));
AOI21X1 g131441(.A0 (n_5770), .A1 (n_4935), .B0 (n_5298), .Y(n_5979));
AOI21X1 g131450(.A0 (n_6045), .A1 (n_6044), .B0 (n_5775), .Y(n_5776));
AOI21X1 g131454(.A0 (n_5328), .A1 (n_5578), .B0 (n_5523), .Y(n_5774));
NAND2X1 g131457(.A (n_5478), .B (n_5772), .Y (n_5773));
XOR2X1 g131497(.A (n_5612), .B (n_5770), .Y (n_5771));
XOR2X1 g131498(.A (n_4799), .B (n_5617), .Y (n_5769));
OAI21X1 g131514(.A0 (n_4957), .A1 (n_5518), .B0 (n_5768), .Y(n_5955));
OR2X1 g131526(.A (n_5709), .B (n_5766), .Y (n_5767));
NOR2X1 g131529(.A (n_5765), .B (n_5764), .Y (n_6038));
NAND2X1 g131533(.A (n_5383), .B (n_5486), .Y (n_5933));
NOR2X1 g131536(.A (n_5763), .B (n_5762), .Y (n_6010));
OR2X1 g131543(.A (n_5526), .B (n_5466), .Y (n_5761));
NOR2X1 g131544(.A (n_5760), .B (n_5759), .Y (n_6015));
NOR2X1 g131555(.A (n_5758), .B (n_5757), .Y (n_6043));
NAND3X1 g131567(.A (n_5755), .B (n_5415), .C (n_5404), .Y (n_5756));
NOR2X1 g131569(.A (n_5753), .B (n_5596), .Y (n_5754));
NAND2X1 g131572(.A (n_5751), .B (n_5925), .Y (n_5752));
NAND2X1 g131576(.A (n_5750), .B (n_5749), .Y (n_5905));
OR2X1 g131585(.A (n_5718), .B (n_5747), .Y (n_5748));
NAND2X1 g131588(.A (n_5378), .B (n_5465), .Y (n_5961));
INVX1 g131591(.A (n_5672), .Y (n_5746));
INVX1 g131593(.A (n_5606), .Y (n_5745));
AOI21X1 g131601(.A0 (n_5395), .A1 (n_5429), .B0 (n_5743), .Y(n_5744));
AOI21X1 g131633(.A0 (n_5542), .A1 (n_5741), .B0 (n_5740), .Y(n_5742));
AND2X1 g131635(.A (n_5525), .B (n_5676), .Y (n_5739));
AOI21X1 g131640(.A0 (n_4258), .A1 (n_5239), .B0 (n_5560), .Y(n_5963));
NAND2X1 g131732(.A (n_5738), .B (n_5333), .Y (n_5911));
INVX1 g131802(.A (n_5736), .Y (n_5737));
INVX1 g131810(.A (n_5734), .Y (n_5735));
XOR2X1 g130840(.A (n_4469), .B (n_5800), .Y (so[9]));
INVX1 g131840(.A (n_5731), .Y (n_5732));
OAI21X1 g131837(.A0 (n_5410), .A1 (n_5089), .B0 (n_5643), .Y(n_6021));
AOI21X1 g131646(.A0 (n_4143), .A1 (n_5391), .B0 (n_5559), .Y(n_5923));
INVX1 g131822(.A (n_5729), .Y (n_5730));
XOR2X1 g130844(.A (n_4685), .B (n_5803), .Y (so[10]));
AND2X1 g131639(.A (n_5558), .B (n_5727), .Y (n_5839));
AND2X1 g131632(.A (n_5471), .B (n_5595), .Y (n_5726));
NAND2X1 g131458(.A (n_5573), .B (n_5724), .Y (n_5725));
AOI21X1 g131448(.A0 (n_5428), .A1 (n_5467), .B0 (n_5517), .Y(n_5723));
NAND2X1 g131757(.A (n_5721), .B (n_5346), .Y (n_5722));
AOI21X1 g131440(.A0 (n_5689), .A1 (n_4836), .B0 (n_5424), .Y(n_5977));
NOR2X1 g131586(.A (n_5719), .B (n_5718), .Y (n_5720));
NAND2X1 g131388(.A (n_5716), .B (n_5635), .Y (n_5717));
AOI21X1 g130834(.A0 (n_5501), .A1 (n_5714), .B0 (n_5352), .Y(n_5715));
XOR2X1 g131370(.A (n_5712), .B (n_5480), .Y (n_5713));
NOR2X1 g131562(.A (n_5710), .B (n_5709), .Y (n_5711));
NAND2X1 g131713(.A (n_5738), .B (n_5708), .Y (n_5932));
NOR2X1 g131545(.A (n_5706), .B (n_5650), .Y (n_5707));
NOR2X1 g131408(.A (n_5704), .B (n_5674), .Y (n_5705));
AOI21X1 g131609(.A0 (n_5540), .A1 (n_5702), .B0 (n_5701), .Y(n_5703));
AOI21X1 g131400(.A0 (n_4391), .A1 (n_5654), .B0 (n_5691), .Y(n_5700));
NOR2X1 g131532(.A (n_5698), .B (n_5659), .Y (n_5699));
OR2X1 g131527(.A (n_5686), .B (n_5696), .Y (n_5697));
OAI21X1 g131516(.A0 (n_5043), .A1 (n_5513), .B0 (n_5695), .Y(n_5913));
OAI21X1 g131240(.A0 (n_5347), .A1 (n_4467), .B0 (n_4502), .Y(n_35295));
AND2X1 g131615(.A (n_5554), .B (n_5693), .Y (n_5843));
NAND2X1 g131391(.A (n_5691), .B (n_5653), .Y (n_5692));
XOR2X1 g131495(.A (n_5609), .B (n_5689), .Y (n_5690));
NOR2X1 g131580(.A (n_5687), .B (n_5686), .Y (n_5688));
AOI22X1 g131482(.A0 (n_5497), .A1 (n_5475), .B0 (n_5055), .B1(n_5086), .Y (n_5685));
NAND3X1 g131716(.A (n_5721), .B (n_6079), .C (n_5925), .Y (n_5894));
XOR2X1 g130634(.A (n_2056), .B (n_5447), .Y (n_5684));
OAI21X1 g131823(.A0 (n_5493), .A1 (n_5592), .B0 (n_5538), .Y(n_5729));
NOR2X1 g130774(.A (n_5682), .B (n_5448), .Y (n_5683));
OR2X1 g130888(.A (n_5340), .B (n_5354), .Y (n_5681));
NAND4X1 g131348(.A (n_4101), .B (n_5262), .C (n_1328), .D (n_1164),.Y (n_5680));
AOI22X1 g131466(.A0 (n_5401), .A1 (n_5419), .B0 (n_5035), .B1(n_5083), .Y (n_5678));
NOR2X1 g131509(.A (n_5200), .B (n_5598), .Y (n_5677));
OAI21X1 g131517(.A0 (n_5093), .A1 (n_5278), .B0 (n_5619), .Y(n_5811));
OAI21X1 g131521(.A0 (n_5044), .A1 (n_5379), .B0 (n_5676), .Y(n_5814));
NOR2X1 g131552(.A (n_5614), .B (n_4584), .Y (n_5675));
NOR2X1 g131568(.A (n_5674), .B (n_5673), .Y (n_5970));
AOI21X1 g131592(.A0 (n_5647), .A1 (n_5254), .B0 (n_5253), .Y(n_5672));
INVX1 g131596(.A (n_5670), .Y (n_5671));
AOI21X1 g131605(.A0 (n_5242), .A1 (n_5425), .B0 (n_5668), .Y(n_5669));
AND2X1 g131628(.A (n_5321), .B (n_5483), .Y (n_5667));
AOI21X1 g131641(.A0 (n_4556), .A1 (n_5140), .B0 (n_5430), .Y(n_6034));
XOR2X1 g131666(.A (n_5300), .B (n_5605), .Y (n_5666));
OAI21X1 g131682(.A0 (n_4924), .A1 (n_5511), .B0 (n_5664), .Y(n_5665));
OAI21X1 g131699(.A0 (n_4744), .A1 (n_5172), .B0 (n_5446), .Y(n_5853));
OAI21X1 g131704(.A0 (n_4606), .A1 (n_5170), .B0 (n_5369), .Y(n_5851));
NOR2X1 g131707(.A (n_4986), .B (n_5349), .Y (n_5860));
NAND2X1 g131710(.A (n_5663), .B (n_5662), .Y (n_5816));
NOR2X1 g131718(.A (n_5660), .B (n_5580), .Y (n_5903));
NAND2X1 g131719(.A (n_5663), .B (n_5570), .Y (n_5833));
OR2X1 g131722(.A (n_5660), .B (n_5659), .Y (n_5661));
NOR2X1 g131738(.A (n_5290), .B (n_5657), .Y (n_5658));
NOR2X1 g131739(.A (n_5575), .B (n_5651), .Y (n_5656));
AND2X1 g131759(.A (n_5654), .B (n_5653), .Y (n_5655));
OR2X1 g131760(.A (n_5651), .B (n_5650), .Y (n_5652));
NOR2X1 g131761(.A (n_5579), .B (n_5660), .Y (n_5649));
AOI21X1 g131803(.A0 (n_5178), .A1 (n_5345), .B0 (n_5317), .Y(n_5736));
AOI21X1 g131811(.A0 (n_5168), .A1 (n_5326), .B0 (n_5319), .Y(n_5734));
XOR2X1 g131656(.A (n_5329), .B (n_5647), .Y (n_5648));
INVX1 g131824(.A (n_5645), .Y (n_5646));
OAI21X1 g131826(.A0 (n_5644), .A1 (n_5643), .B0 (n_5023), .Y(n_5847));
OAI21X1 g131841(.A0 (n_5225), .A1 (n_5510), .B0 (n_5535), .Y(n_5731));
INVX1 g131842(.A (n_5641), .Y (n_5642));
NAND2X1 g131919(.A (n_5396), .B (n_5358), .Y (n_5640));
NAND2X1 g131921(.A (n_5532), .B (n_5441), .Y (n_5639));
NAND2X1 g131923(.A (n_4965), .B (n_5357), .Y (n_5638));
AND2X1 g131737(.A (n_5636), .B (n_5635), .Y (n_5637));
NAND2X1 g132015(.A (n_5364), .B (n_5628), .Y (n_6102));
NOR2X1 g132020(.A (n_5644), .B (n_5410), .Y (n_5819));
AOI21X1 g131645(.A0 (n_4523), .A1 (n_4977), .B0 (n_5426), .Y(n_6036));
NOR2X1 g132416(.A (n_5342), .B (n_5593), .Y (n_5634));
OR2X1 g131528(.A (n_5625), .B (n_5632), .Y (n_5633));
OAI21X1 g131686(.A0 (n_4472), .A1 (n_5515), .B0 (n_5630), .Y(n_5631));
NAND3X1 g131335(.A (n_35871), .B (n_5266), .C (n_35872), .Y (n_5629));
OAI21X1 g131821(.A0 (n_5484), .A1 (n_5384), .B0 (n_5628), .Y(n_5926));
NOR2X1 g131535(.A (n_5626), .B (n_5625), .Y (n_5627));
AOI21X1 g131394(.A0 (n_5229), .A1 (n_5624), .B0 (n_5623), .Y(n_5877));
AOI21X1 g131621(.A0 (n_5432), .A1 (n_4963), .B0 (n_5375), .Y(n_5621));
AND2X1 g131612(.A (n_5303), .B (n_5619), .Y (n_5620));
NAND3X1 g131542(.A (n_5617), .B (n_5412), .C (n_5252), .Y (n_5618));
AOI21X1 g131610(.A0 (n_5545), .A1 (n_5187), .B0 (n_5373), .Y(n_5616));
NOR2X1 g131513(.A (n_34507), .B (n_5614), .Y (n_5615));
XOR2X1 g131499(.A (n_5612), .B (n_5611), .Y (n_5613));
XOR2X1 g131496(.A (n_5609), .B (n_5608), .Y (n_5610));
NAND3X1 g131292(.A (n_2211), .B (n_3510), .C (n_5261), .Y (n_5607));
AOI21X1 g131594(.A0 (n_5605), .A1 (n_5136), .B0 (n_5135), .Y(n_5606));
NOR2X1 g131583(.A (n_5604), .B (n_5603), .Y (n_5897));
NOR2X1 g131747(.A (n_5651), .B (n_5576), .Y (n_5908));
NAND2X1 g131914(.A (n_5507), .B (n_5359), .Y (n_5602));
NOR2X1 g131570(.A (n_5600), .B (n_5468), .Y (n_5601));
NOR2X1 g131571(.A (n_5598), .B (n_4582), .Y (n_5599));
NAND2X1 g131519(.A (n_5608), .B (n_5386), .Y (n_5597));
NOR2X1 g131731(.A (n_5657), .B (n_5596), .Y (n_5850));
OAI21X1 g131520(.A0 (n_4984), .A1 (n_5348), .B0 (n_5595), .Y(n_5859));
OAI21X1 g132114(.A0 (n_5221), .A1 (n_5593), .B0 (n_5592), .Y(n_5740));
NAND2X1 g131733(.A (n_5591), .B (n_5590), .Y (n_5763));
NOR2X1 g130890(.A (n_5588), .B (n_5500), .Y (n_5589));
NAND2X1 g131117(.A (n_5586), .B (n_5585), .Y (n_5587));
AOI21X1 g131334(.A0 (n_4780), .A1 (n_1357), .B0 (n_5196), .Y(n_5583));
NOR2X1 g131447(.A (n_3615), .B (n_33480), .Y (n_5582));
OAI21X1 g131504(.A0 (n_5431), .A1 (n_5580), .B0 (n_5579), .Y(n_5581));
OAI21X1 g131507(.A0 (n_4953), .A1 (n_5193), .B0 (n_5578), .Y(n_5716));
OAI21X1 g131512(.A0 (n_5443), .A1 (n_5576), .B0 (n_5575), .Y(n_5577));
NOR2X1 g131563(.A (n_5461), .B (n_4419), .Y (n_5573));
OAI21X1 g131590(.A0 (n_4917), .A1 (n_5126), .B0 (n_5255), .Y(n_5869));
AOI21X1 g131607(.A0 (n_5405), .A1 (n_5571), .B0 (n_5550), .Y(n_5786));
AOI21X1 g131620(.A0 (n_5343), .A1 (n_5570), .B0 (n_5569), .Y(n_5863));
AOI21X1 g131622(.A0 (n_5409), .A1 (n_5315), .B0 (n_5568), .Y(n_5783));
AOI21X1 g131623(.A0 (n_5530), .A1 (n_5566), .B0 (n_5174), .Y(n_5567));
AOI21X1 g131636(.A0 (n_5355), .A1 (n_5564), .B0 (n_5250), .Y(n_5565));
AOI21X1 g131637(.A0 (n_5411), .A1 (n_5563), .B0 (n_5556), .Y(n_5781));
XOR2X1 g131657(.A (n_4871), .B (n_5470), .Y (n_5562));
XOR2X1 g131663(.A (n_5393), .B (n_5427), .Y (n_5561));
OAI21X1 g131684(.A0 (n_4826), .A1 (n_5238), .B0 (n_5374), .Y(n_5560));
OAI21X1 g131685(.A0 (n_5041), .A1 (n_5054), .B0 (n_5224), .Y(n_5755));
OAI21X1 g131705(.A0 (n_5096), .A1 (n_5390), .B0 (n_5372), .Y(n_5559));
NOR2X1 g131706(.A (n_5095), .B (n_5279), .Y (n_5812));
OR2X1 g131711(.A (n_5318), .B (n_5150), .Y (n_5558));
NAND2X1 g131720(.A (n_5556), .B (n_5555), .Y (n_5557));
OR2X1 g131723(.A (n_5316), .B (n_5210), .Y (n_5554));
NAND2X1 g131724(.A (n_5488), .B (n_5552), .Y (n_5553));
NAND2X1 g131728(.A (n_5550), .B (n_5591), .Y (n_5551));
NAND2X1 g131730(.A (n_5549), .B (n_5548), .Y (n_5764));
NAND2X1 g131741(.A (n_5552), .B (n_5547), .Y (n_5760));
XOR2X1 g131660(.A (n_4235), .B (n_5545), .Y (n_5546));
NAND2X1 g131753(.A (n_5948), .B (n_5702), .Y (n_5709));
NOR2X1 g131755(.A (n_3289), .B (n_5163), .Y (n_5996));
NAND2X1 g131763(.A (n_5938), .B (n_5741), .Y (n_5718));
AOI21X1 g131774(.A0 (n_5368), .A1 (n_5544), .B0 (n_5287), .Y(n_5695));
AOI21X1 g131777(.A0 (n_5628), .A1 (n_5519), .B0 (n_5484), .Y(n_5753));
AOI21X1 g131778(.A0 (n_5485), .A1 (n_5543), .B0 (n_5542), .Y(n_5719));
AOI21X1 g131791(.A0 (n_5464), .A1 (n_5541), .B0 (n_5540), .Y(n_5710));
AOI21X1 g131797(.A0 (n_5410), .A1 (n_5023), .B0 (n_5644), .Y(n_5706));
OAI21X1 g131820(.A0 (n_5539), .A1 (n_5628), .B0 (n_5444), .Y(n_5751));
OAI21X1 g131825(.A0 (n_5538), .A1 (n_5240), .B0 (n_4997), .Y(n_5645));
INVX1 g131829(.A (n_5536), .Y (n_5537));
OAI21X1 g131843(.A0 (n_5535), .A1 (n_5226), .B0 (n_5038), .Y(n_5641));
XOR2X1 g131849(.A (n_5039), .B (n_5382), .Y (n_5534));
XOR2X1 g131873(.A (n_3838), .B (n_5532), .Y (n_5533));
OAI21X1 g131875(.A0 (n_5530), .A1 (n_5399), .B0 (n_5233), .Y(n_5531));
XOR2X1 g131879(.A (n_4186), .B (n_5524), .Y (n_5529));
NOR2X1 g131908(.A (n_5398), .B (n_5158), .Y (n_5526));
NAND2X1 g131910(.A (n_5524), .B (n_5208), .Y (n_5525));
INVX1 g131939(.A (n_5635), .Y (n_5523));
INVX1 g131942(.A (n_5521), .Y (n_5522));
NAND2X1 g131968(.A (n_5361), .B (n_5643), .Y (n_6150));
NOR2X1 g131969(.A (n_5484), .B (n_5519), .Y (n_5738));
NOR2X1 g131980(.A (n_5518), .B (n_4497), .Y (n_5957));
INVX1 g132010(.A (n_5653), .Y (n_5517));
NOR2X1 g132019(.A (n_4473), .B (n_5515), .Y (n_5516));
NOR2X1 g132030(.A (n_5644), .B (n_5514), .Y (n_6326));
NOR2X1 g132037(.A (n_5513), .B (n_4566), .Y (n_5915));
NOR2X1 g132049(.A (n_4925), .B (n_5511), .Y (n_5512));
OAI21X1 g132127(.A0 (n_5155), .A1 (n_5206), .B0 (n_5510), .Y(n_5701));
NAND2X1 g132375(.A (n_5510), .B (n_5027), .Y (n_5509));
XOR2X1 g131850(.A (n_3937), .B (n_5507), .Y (n_5508));
INVX1 g131838(.A (n_5505), .Y (n_5506));
AOI21X1 g130901(.A0 (n_5503), .A1 (n_5502), .B0 (n_5501), .Y(n_5504));
NOR2X1 g130891(.A (n_5350), .B (n_5500), .Y (n_5795));
NOR2X1 g132040(.A (n_5055), .B (n_5442), .Y (n_5499));
INVX1 g131831(.A (n_5497), .Y (n_5498));
XOR2X1 g131851(.A (n_4220), .B (n_5320), .Y (n_5496));
NOR2X1 g132056(.A (n_5539), .B (n_5484), .Y (n_5721));
XOR2X1 g131662(.A (n_4886), .B (n_5302), .Y (n_5495));
NOR2X1 g132021(.A (n_5148), .B (n_5493), .Y (n_5494));
XOR2X1 g130629(.A (n_1478), .B (n_5125), .Y (n_5492));
AOI21X1 g131807(.A0 (n_5445), .A1 (n_5491), .B0 (n_5407), .Y(n_5768));
OAI21X1 g130658(.A0 (n_5438), .A1 (n_5450), .B0 (n_5453), .Y(n_5990));
AOI21X1 g131631(.A0 (n_5285), .A1 (n_5489), .B0 (n_5488), .Y(n_5779));
AOI21X1 g131626(.A0 (n_4770), .A1 (n_5344), .B0 (n_5487), .Y(n_5827));
AOI21X1 g131787(.A0 (n_5370), .A1 (n_5381), .B0 (n_5485), .Y(n_5486));
AOI21X1 g131775(.A0 (n_5484), .A1 (n_5444), .B0 (n_5539), .Y(n_5698));
OAI21X1 g131515(.A0 (n_5021), .A1 (n_5227), .B0 (n_5483), .Y(n_5775));
OAI21X1 g131595(.A0 (n_4802), .A1 (n_5130), .B0 (n_5138), .Y(n_5866));
INVX1 g131598(.A (n_5480), .Y (n_5481));
AOI21X1 g131597(.A0 (n_5455), .A1 (n_4822), .B0 (n_5111), .Y(n_5670));
AOI21X1 g131617(.A0 (n_5414), .A1 (n_5479), .B0 (n_5307), .Y(n_5704));
NAND2X1 g131503(.A (n_5611), .B (n_5181), .Y (n_5478));
NAND2X1 g131746(.A (n_5555), .B (n_5475), .Y (n_5758));
NOR2X1 g131911(.A (n_5296), .B (n_5141), .Y (n_5474));
NOR2X1 g131725(.A (n_34234), .B (n_34947), .Y (n_6060));
XOR2X1 g131877(.A (n_5037), .B (n_5377), .Y (n_5472));
NAND2X1 g131708(.A (n_5549), .B (n_5458), .Y (n_5686));
NAND2X1 g131700(.A (n_5470), .B (n_5207), .Y (n_5471));
NOR2X1 g131749(.A (n_5469), .B (n_5468), .Y (n_5750));
OAI21X1 g131511(.A0 (n_5099), .A1 (n_5235), .B0 (n_5467), .Y(n_5691));
AOI21X1 g131625(.A0 (n_4804), .A1 (n_5325), .B0 (n_5466), .Y(n_5824));
AOI21X1 g131784(.A0 (n_5366), .A1 (n_5376), .B0 (n_5464), .Y(n_5465));
NOR2X1 g131508(.A (n_5462), .B (n_5461), .Y (n_5463));
INVX1 g131999(.A (n_5459), .Y (n_5460));
AOI21X1 g131627(.A0 (n_5337), .A1 (n_5458), .B0 (n_5457), .Y(n_5777));
XOR2X1 g131667(.A (n_5283), .B (n_5455), .Y (n_5456));
NOR2X1 g130895(.A (n_5453), .B (n_5451), .Y (n_5454));
NAND4X1 g131159(.A (n_696), .B (n_1783), .C (n_3251), .D (n_4848), .Y(n_5452));
NOR2X1 g130885(.A (n_5451), .B (n_5450), .Y (n_5889));
XOR2X1 g131251(.A (n_4526), .B (n_5503), .Y (so[8]));
NOR2X1 g130889(.A (n_5451), .B (n_5448), .Y (n_5793));
NAND3X1 g130870(.A (n_2442), .B (n_3786), .C (n_4949), .Y (n_5447));
AOI21X1 g132095(.A0 (n_4649), .A1 (n_5171), .B0 (n_5445), .Y(n_5446));
NAND2X1 g131941(.A (n_5444), .B (n_5628), .Y (n_5660));
OAI21X1 g131696(.A0 (n_5109), .A1 (n_5292), .B0 (n_5443), .Y(n_5929));
OAI21X1 g131830(.A0 (n_5442), .A1 (n_5353), .B0 (n_5211), .Y(n_5536));
INVX1 g132357(.A (n_5518), .Y (n_5441));
AND2X1 g132046(.A (n_5564), .B (n_5439), .Y (n_5440));
OAI21X1 g130871(.A0 (n_5122), .A1 (n_5312), .B0 (n_5351), .Y(n_5796));
OAI21X1 g130872(.A0 (n_5012), .A1 (n_5436), .B0 (n_5438), .Y(n_5798));
AOI21X1 g130904(.A0 (n_5271), .A1 (n_5273), .B0 (n_5437), .Y(n_5682));
NOR2X1 g131140(.A (n_5450), .B (n_5436), .Y (n_5792));
NAND3X1 g131155(.A (n_4968), .B (n_4682), .C (n_5124), .Y (n_5803));
NAND2X1 g131439(.A (n_4941), .B (n_5114), .Y (n_5435));
NAND4X1 g131449(.A (n_5259), .B (n_4936), .C (n_5260), .D (n_4315),.Y (n_32202));
OAI21X1 g131506(.A0 (n_5423), .A1 (n_5236), .B0 (n_5421), .Y(n_6048));
OAI21X1 g131518(.A0 (n_4845), .A1 (n_4863), .B0 (n_5173), .Y(n_5623));
XOR2X1 g131665(.A (n_4226), .B (n_5432), .Y (n_5433));
OAI21X1 g131678(.A0 (n_4893), .A1 (n_4914), .B0 (n_4970), .Y(n_5617));
OAI21X1 g131695(.A0 (n_5106), .A1 (n_5388), .B0 (n_5431), .Y(n_5943));
OAI21X1 g131697(.A0 (n_4900), .A1 (n_5139), .B0 (n_5429), .Y(n_5430));
NAND2X1 g131698(.A (n_5427), .B (n_5051), .Y (n_5428));
OAI21X1 g131702(.A0 (n_4899), .A1 (n_4976), .B0 (n_5425), .Y(n_5426));
OAI21X1 g131703(.A0 (n_5151), .A1 (n_5237), .B0 (n_5423), .Y(n_5424));
NAND2X1 g131735(.A (n_5080), .B (n_4942), .Y (n_5598));
NOR2X1 g131743(.A (n_5421), .B (n_5469), .Y (n_5422));
NAND2X1 g131745(.A (n_5420), .B (n_5419), .Y (n_5674));
NAND2X1 g131758(.A (n_5418), .B (n_5417), .Y (n_5603));
AOI21X1 g131781(.A0 (n_5222), .A1 (n_5275), .B0 (n_5338), .Y(n_5619));
AOI21X1 g131783(.A0 (n_5403), .A1 (n_5415), .B0 (n_5414), .Y(n_5416));
AOI21X1 g131790(.A0 (n_5251), .A1 (n_5412), .B0 (n_5411), .Y(n_5413));
AOI21X1 g131804(.A0 (n_5643), .A1 (n_5387), .B0 (n_5410), .Y(n_5600));
AOI21X1 g131809(.A0 (n_5334), .A1 (n_5230), .B0 (n_5409), .Y(n_5626));
AOI21X1 g131815(.A0 (n_5407), .A1 (n_5406), .B0 (n_5405), .Y(n_5408));
AOI21X1 g131816(.A0 (n_5223), .A1 (n_5404), .B0 (n_5403), .Y(n_5676));
INVX1 g131827(.A (n_5401), .Y (n_5402));
OAI21X1 g131839(.A0 (n_5305), .A1 (n_5197), .B0 (n_5056), .Y(n_5505));
XOR2X1 g131869(.A (n_5399), .B (n_5398), .Y (n_5400));
XOR2X1 g131876(.A (n_4146), .B (n_5396), .Y (n_5397));
NAND2X1 g131915(.A (n_5299), .B (n_5030), .Y (n_5395));
XOR2X1 g131655(.A (n_5393), .B (n_5322), .Y (n_5394));
NAND2X1 g131934(.A (n_5535), .B (n_5064), .Y (n_5392));
NOR2X1 g131945(.A (n_5098), .B (n_5390), .Y (n_5391));
NOR2X1 g131946(.A (n_5388), .B (n_5580), .Y (n_5389));
NOR2X1 g131958(.A (n_5410), .B (n_5387), .Y (n_5663));
INVX1 g132005(.A (n_5385), .Y (n_5386));
NAND2X1 g132013(.A (n_5628), .B (n_5384), .Y (n_5657));
NAND3X1 g132041(.A (n_5382), .B (n_5381), .C (n_5371), .Y (n_5383));
NOR2X1 g132045(.A (n_5198), .B (n_5045), .Y (n_5380));
NOR2X1 g132051(.A (n_5379), .B (n_4563), .Y (n_5971));
NAND3X1 g132058(.A (n_5377), .B (n_5376), .C (n_5367), .Y (n_5378));
INVX1 g132083(.A (n_5374), .Y (n_5375));
INVX1 g132092(.A (n_5372), .Y (n_5373));
AOI21X1 g132096(.A0 (n_4551), .A1 (n_5371), .B0 (n_5370), .Y(n_5664));
AOI21X1 g132102(.A0 (n_4573), .A1 (n_5199), .B0 (n_5368), .Y(n_5369));
AOI21X1 g132104(.A0 (n_4624), .A1 (n_5367), .B0 (n_5366), .Y(n_5630));
AND2X1 g132118(.A (n_5024), .B (n_5384), .Y (n_5693));
INVX1 g132216(.A (n_5484), .Y (n_5364));
INVX1 g132286(.A (n_5513), .Y (n_5359));
INVX1 g132297(.A (n_5511), .Y (n_5358));
INVX1 g132326(.A (n_5515), .Y (n_5357));
XOR2X1 g131857(.A (n_5295), .B (n_5355), .Y (n_5356));
AND2X1 g132128(.A (n_5065), .B (n_5089), .Y (n_5727));
AOI21X1 g130902(.A0 (n_4946), .A1 (n_5159), .B0 (n_5354), .Y(n_5808));
OAI21X1 g131832(.A0 (n_5335), .A1 (n_4800), .B0 (n_5353), .Y(n_5497));
NOR2X1 g130882(.A (n_5351), .B (n_5350), .Y (n_5352));
NAND3X1 g131818(.A (n_5081), .B (n_4710), .C (n_5152), .Y (n_5689));
OR2X1 g132033(.A (n_5348), .B (n_4985), .Y (n_5349));
NAND4X1 g131452(.A (n_33009), .B (n_4158), .C (n_3868), .D (n_33010),.Y (n_5347));
AND2X1 g132011(.A (n_5346), .B (n_5345), .Y (n_5653));
AND2X1 g132000(.A (n_5344), .B (n_4771), .Y (n_5459));
AOI21X1 g131801(.A0 (n_5009), .A1 (n_5331), .B0 (n_5343), .Y(n_5822));
INVX1 g132692(.A (n_5592), .Y (n_5342));
NOR2X1 g131982(.A (n_5539), .B (n_5341), .Y (n_6359));
NOR2X1 g131192(.A (n_5310), .B (n_4989), .Y (n_5340));
AOI21X1 g131785(.A0 (n_5338), .A1 (n_5274), .B0 (n_5337), .Y(n_5687));
NOR2X1 g131970(.A (n_5335), .B (n_4974), .Y (n_5336));
AOI21X1 g131782(.A0 (n_5280), .A1 (n_5231), .B0 (n_5334), .Y(n_5595));
AOI21X1 g131613(.A0 (n_5248), .A1 (n_5333), .B0 (n_5332), .Y(n_5880));
NAND2X1 g131949(.A (n_5331), .B (n_5570), .Y (n_5815));
XOR2X1 g131878(.A (n_5329), .B (n_5241), .Y (n_5330));
NAND2X1 g131679(.A (n_5282), .B (n_5004), .Y (n_5328));
AND2X1 g131940(.A (n_5327), .B (n_5326), .Y (n_5635));
AND2X1 g131943(.A (n_5325), .B (n_4805), .Y (n_5521));
NAND2X1 g131926(.A (n_5023), .B (n_5643), .Y (n_5651));
AOI21X1 g131599(.A0 (n_5322), .A1 (n_4807), .B0 (n_5108), .Y(n_5480));
NAND2X1 g131920(.A (n_5320), .B (n_5000), .Y (n_5321));
NAND3X1 g131145(.A (n_5119), .B (n_4786), .C (n_5014), .Y (n_5800));
INVX1 g132134(.A (n_5318), .Y (n_5319));
INVX1 g132125(.A (n_5316), .Y (n_5317));
NAND2X1 g131721(.A (n_5418), .B (n_5315), .Y (n_5625));
NOR2X1 g131136(.A (n_5350), .B (n_5312), .Y (n_5714));
XOR2X1 g131250(.A (n_4115), .B (n_5310), .Y (so[7]));
NAND2X1 g131709(.A (n_5307), .B (n_5420), .Y (n_5308));
NOR2X1 g131948(.A (n_5035), .B (n_5305), .Y (n_5306));
NAND2X1 g131729(.A (n_5078), .B (n_34434), .Y (n_5614));
NOR2X1 g131121(.A (n_5437), .B (n_5118), .Y (n_5304));
NAND2X1 g131689(.A (n_5302), .B (n_5059), .Y (n_5303));
XOR2X1 g131871(.A (n_5300), .B (n_5299), .Y (n_5301));
OAI21X1 g131694(.A0 (n_5142), .A1 (n_5277), .B0 (n_5291), .Y(n_5298));
OAI21X1 g131870(.A0 (n_5296), .A1 (n_5295), .B0 (n_5134), .Y(n_5297));
XOR2X1 g131373(.A (n_1339), .B (n_4815), .Y (n_5294));
NOR2X1 g131951(.A (n_5292), .B (n_5576), .Y (n_5293));
OAI21X1 g131505(.A0 (n_5291), .A1 (n_5276), .B0 (n_5290), .Y(n_6047));
OAI21X1 g131510(.A0 (n_4926), .A1 (n_5005), .B0 (n_5249), .Y(n_5806));
AOI22X1 g132176(.A0 (n_4720), .A1 (n_13329), .B0 (n_4844), .B1(n_5289), .Y (n_6334));
NAND3X1 g131819(.A (n_5088), .B (n_4671), .C (n_5143), .Y (n_5770));
AOI21X1 g131814(.A0 (n_5287), .A1 (n_5286), .B0 (n_5285), .Y(n_5288));
XOR2X1 g131658(.A (n_5283), .B (n_5282), .Y (n_5284));
NOR2X1 g131328(.A (n_4992), .B (n_2053), .Y (n_5281));
NAND2X1 g132012(.A (n_5444), .B (n_5946), .Y (n_5596));
AOI21X1 g132093(.A0 (n_4755), .A1 (n_5049), .B0 (n_5280), .Y(n_5372));
OR2X1 g132032(.A (n_5278), .B (n_5094), .Y (n_5279));
NOR2X1 g132009(.A (n_5277), .B (n_5276), .Y (n_5849));
NAND2X1 g132008(.A (n_5169), .B (n_5326), .Y (n_5743));
NAND2X1 g131927(.A (n_5275), .B (n_5274), .Y (n_5696));
AOI21X1 g132091(.A0 (n_4975), .A1 (n_5384), .B0 (n_5519), .Y(n_5579));
NAND2X1 g131139(.A (n_5273), .B (n_5272), .Y (n_5500));
AOI21X1 g131342(.A0 (n_5203), .A1 (n_5176), .B0 (n_5271), .Y(n_5588));
NOR2X1 g131347(.A (n_4788), .B (n_4854), .Y (n_5270));
XOR2X1 g131368(.A (n_1960), .B (n_4689), .Y (n_5269));
NOR2X1 g131524(.A (n_34507), .B (n_35167), .Y (n_35871));
NOR2X1 g131548(.A (n_4820), .B (n_5077), .Y (n_5266));
NOR2X1 g131582(.A (n_4943), .B (n_5079), .Y (n_32054));
AOI21X1 g131649(.A0 (n_4416), .A1 (n_1748), .B0 (n_4857), .Y(n_5263));
NAND4X1 g131650(.A (n_3506), .B (n_4334), .C (n_4100), .D (n_5028),.Y (n_5262));
NAND4X1 g131654(.A (n_4282), .B (n_2992), .C (n_3509), .D (n_5006),.Y (n_5261));
NAND2X1 g131756(.A (n_5260), .B (n_5259), .Y (n_5461));
NAND2X1 g131768(.A (n_4931), .B (n_4940), .Y (n_5258));
NAND4X1 g131769(.A (n_4723), .B (n_4355), .C (n_32241), .D (n_34120),.Y (n_5257));
AOI21X1 g131779(.A0 (n_5232), .A1 (n_5254), .B0 (n_5253), .Y(n_5255));
AOI21X1 g131780(.A0 (n_4969), .A1 (n_5252), .B0 (n_5251), .Y(n_5483));
INVX1 g131788(.A (n_5249), .Y (n_5250));
AOI21X1 g131812(.A0 (n_5104), .A1 (n_5167), .B0 (n_5248), .Y(n_5772));
INVX1 g131833(.A (n_5246), .Y (n_5247));
INVX1 g131835(.A (n_5244), .Y (n_5245));
NAND2X1 g131906(.A (n_5241), .B (n_4906), .Y (n_5242));
NOR2X1 g131930(.A (n_5240), .B (n_5493), .Y (n_5938));
NAND2X1 g131935(.A (n_5286), .B (n_5489), .Y (n_5759));
NOR2X1 g131938(.A (n_5493), .B (n_5593), .Y (n_5591));
NAND2X1 g131944(.A (n_5376), .B (n_5541), .Y (n_5766));
NOR2X1 g131963(.A (n_4828), .B (n_5238), .Y (n_5239));
NOR2X1 g131972(.A (n_5335), .B (n_5442), .Y (n_5549));
NOR2X1 g131975(.A (n_5237), .B (n_5236), .Y (n_5749));
NOR2X1 g131981(.A (n_5335), .B (n_4909), .Y (n_5555));
NAND2X1 g131988(.A (n_5274), .B (n_5458), .Y (n_5765));
NOR2X1 g131996(.A (n_5110), .B (n_5292), .Y (n_5907));
NOR2X1 g132001(.A (n_5235), .B (n_5100), .Y (n_5654));
NOR2X1 g132017(.A (n_5539), .B (n_5234), .Y (n_5708));
OR2X1 g132024(.A (n_4803), .B (n_5137), .Y (n_5605));
NAND2X1 g132026(.A (n_5530), .B (n_5399), .Y (n_5233));
OR2X1 g132028(.A (n_4918), .B (n_5232), .Y (n_5647));
NOR2X1 g132038(.A (n_5644), .B (n_4923), .Y (n_5662));
NAND2X1 g132039(.A (n_5231), .B (n_5230), .Y (n_5632));
AND2X1 g132043(.A (n_5566), .B (n_5228), .Y (n_5229));
NOR2X1 g132044(.A (n_5227), .B (n_4560), .Y (n_6045));
NAND2X1 g132048(.A (n_5412), .B (n_5563), .Y (n_5757));
NAND2X1 g132053(.A (n_5415), .B (n_5479), .Y (n_5673));
NOR2X1 g132055(.A (n_5226), .B (n_5225), .Y (n_5948));
NAND2X1 g132060(.A (n_5406), .B (n_5571), .Y (n_5762));
AOI21X1 g132081(.A0 (n_4725), .A1 (n_5053), .B0 (n_5223), .Y(n_5224));
AOI21X1 g132084(.A0 (n_4699), .A1 (n_4872), .B0 (n_5222), .Y(n_5374));
AOI21X1 g132101(.A0 (n_5073), .A1 (n_5089), .B0 (n_5387), .Y(n_5575));
OAI21X1 g132113(.A0 (n_5073), .A1 (n_5160), .B0 (n_5215), .Y(n_5569));
OAI21X1 g132117(.A0 (n_4861), .A1 (n_5061), .B0 (n_5156), .Y(n_5540));
OAI21X1 g132120(.A0 (n_5216), .A1 (n_5220), .B0 (n_5221), .Y(n_5550));
AND2X1 g132126(.A (n_4922), .B (n_5076), .Y (n_5316));
OAI21X1 g132133(.A0 (n_5185), .A1 (n_4982), .B0 (n_5220), .Y(n_5542));
INVX1 g132146(.A (n_5219), .Y (n_5874));
AOI22X1 g132161(.A0 (n_35180), .A1 (n_358), .B0 (n_35188), .B1(P2_reg1[19] ), .Y (n_6320));
XOR2X1 g132162(.A (P1_reg2[19] ), .B (n_6204), .Y (n_5218));
INVX1 g132235(.A (n_5023), .Y (n_5514));
INVX1 g132241(.A (n_5410), .Y (n_5361));
NOR2X1 g132254(.A (n_5216), .B (n_5593), .Y (n_5741));
NAND2X1 g132255(.A (n_4690), .B (n_5215), .Y (n_6134));
NOR2X1 g132275(.A (n_5387), .B (n_5127), .Y (n_6143));
NOR2X1 g132295(.A (n_5213), .B (n_5240), .Y (n_5214));
NAND2X1 g132298(.A (n_4552), .B (n_5371), .Y (n_5511));
NAND2X1 g132327(.A (n_4625), .B (n_5367), .Y (n_5515));
INVX1 g132368(.A (n_5346), .Y (n_5210));
INVX1 g132387(.A (n_5379), .Y (n_5208));
NOR2X1 g132396(.A (n_5519), .B (n_4834), .Y (n_6146));
INVX1 g132421(.A (n_5348), .Y (n_5207));
NAND2X1 g132735(.A (n_33034), .B (P1_reg1[14] ), .Y (n_5510));
NOR2X1 g132317(.A (n_5157), .B (n_5206), .Y (n_5702));
OR2X1 g132335(.A (n_5204), .B (n_5226), .Y (n_5205));
AOI21X1 g131338(.A0 (n_5120), .A1 (n_5146), .B0 (n_5203), .Y(n_5453));
NOR2X1 g132303(.A (n_4983), .B (n_4866), .Y (n_5202));
NAND2X1 g132287(.A (n_5544), .B (n_5199), .Y (n_5513));
OAI21X1 g131828(.A0 (n_5198), .A1 (n_4927), .B0 (n_5197), .Y(n_5401));
OAI22X1 g131487(.A0 (n_5195), .A1 (n_5194), .B0 (n_4781), .B1(n_1356), .Y (n_5196));
NOR2X1 g132052(.A (n_5193), .B (n_4954), .Y (n_5636));
AOI21X1 g131647(.A0 (n_4441), .A1 (n_1374), .B0 (n_4939), .Y(n_5192));
OAI22X1 g131459(.A0 (n_5190), .A1 (n_5189), .B0 (n_5188), .B1(n_1916), .Y (n_5191));
NOR2X1 g132036(.A (n_5107), .B (n_5388), .Y (n_5902));
INVX1 g132384(.A (n_5390), .Y (n_5187));
NOR2X1 g132755(.A (n_4839), .B (n_5185), .Y (n_5186));
NAND2X1 g132018(.A (n_5179), .B (n_5345), .Y (n_5668));
XOR2X1 g131364(.A (n_4013), .B (n_4967), .Y (so[6]));
OAI21X1 g131337(.A0 (n_5182), .A1 (n_428), .B0 (n_4881), .Y (n_5183));
NAND2X1 g132006(.A (n_5010), .B (n_5331), .Y (n_5385));
INVX1 g132003(.A (n_5180), .Y (n_5181));
NAND2X1 g132693(.A (n_33034), .B (P1_reg2[14] ), .Y (n_5592));
AOI21X1 g131800(.A0 (n_5011), .A1 (n_5179), .B0 (n_5178), .Y(n_5467));
NAND2X1 g131398(.A (n_4945), .B (n_5176), .Y (n_5177));
NAND3X1 g131796(.A (n_5175), .B (n_4418), .C (n_4508), .Y (n_5462));
INVX1 g131792(.A (n_5173), .Y (n_5174));
NOR2X1 g131974(.A (n_5225), .B (n_5206), .Y (n_5552));
NAND2X1 g132372(.A (n_4650), .B (n_5171), .Y (n_5172));
NAND2X1 g131965(.A (n_5381), .B (n_5543), .Y (n_5747));
NAND2X1 g132340(.A (n_4574), .B (n_5199), .Y (n_5170));
AOI21X1 g131776(.A0 (n_5074), .A1 (n_5169), .B0 (n_5168), .Y(n_5578));
NAND2X1 g131952(.A (n_5167), .B (n_5333), .Y (n_5881));
AOI22X1 g132164(.A0 (n_35180), .A1 (n_352), .B0 (n_35188), .B1(P2_reg2[19] ), .Y (n_6270));
XOR2X1 g131494(.A (n_1967), .B (n_4695), .Y (n_5164));
NAND2X1 g131932(.A (n_5023), .B (n_6017), .Y (n_5468));
NAND2X1 g131931(.A (n_5230), .B (n_5315), .Y (n_5604));
INVX1 g132147(.A (n_5219), .Y (n_5163));
NAND2X1 g132358(.A (n_5491), .B (n_5171), .Y (n_5518));
NOR2X1 g131600(.A (n_4346), .B (n_4812), .Y (n_32105));
AND2X1 g132135(.A (n_4904), .B (n_5160), .Y (n_5318));
AND2X1 g131204(.A (n_5159), .B (n_4947), .Y (n_5585));
OAI21X1 g131742(.A0 (n_4888), .A1 (n_4654), .B0 (n_4841), .Y(n_5608));
INVX1 g132419(.A (n_5325), .Y (n_5158));
NAND2X1 g131130(.A (n_5176), .B (n_5273), .Y (n_5451));
NOR2X1 g131142(.A (n_5436), .B (n_5013), .Y (n_5799));
OAI21X1 g132122(.A0 (n_5157), .A1 (n_5156), .B0 (n_5155), .Y(n_5488));
OAI21X1 g131717(.A0 (n_5002), .A1 (n_4652), .B0 (n_4811), .Y(n_5611));
NOR2X1 g131122(.A (n_5312), .B (n_5123), .Y (n_5802));
OAI21X1 g131691(.A0 (n_5152), .A1 (n_5052), .B0 (n_5151), .Y(n_5487));
INVX1 g132446(.A (n_5327), .Y (n_5150));
NAND2X1 g131414(.A (n_5272), .B (n_5149), .Y (n_5448));
INVX1 g132433(.A (n_5538), .Y (n_5148));
NAND2X1 g131416(.A (n_4823), .B (n_5146), .Y (n_5147));
AND2X1 g131417(.A (n_5144), .B (n_5149), .Y (n_5145));
OAI21X1 g131690(.A0 (n_5143), .A1 (n_5046), .B0 (n_5142), .Y(n_5466));
INVX1 g132354(.A (n_5344), .Y (n_5141));
NOR2X1 g131936(.A (n_4380), .B (n_5139), .Y (n_5140));
AOI21X1 g131805(.A0 (n_5137), .A1 (n_5136), .B0 (n_5135), .Y(n_5138));
OAI21X1 g132116(.A0 (n_4907), .A1 (n_5071), .B0 (n_4929), .Y(n_5307));
NAND2X1 g132031(.A (n_5296), .B (n_5295), .Y (n_5134));
NAND2X1 g132034(.A (n_5132), .B (n_5131), .Y (n_5133));
NOR2X1 g131971(.A (n_5198), .B (n_5305), .Y (n_5418));
NAND2X1 g131909(.A (n_4658), .B (n_5136), .Y (n_5130));
OAI21X1 g131834(.A0 (n_4932), .A1 (n_5129), .B0 (n_4361), .Y(n_5246));
NAND2X1 g131907(.A (n_4797), .B (n_5254), .Y (n_5126));
NAND3X1 g130903(.A (n_1550), .B (n_3527), .C (n_4646), .Y (n_5125));
OAI21X1 g131116(.A0 (n_5124), .A1 (n_5123), .B0 (n_5122), .Y(n_5501));
AOI21X1 g131151(.A0 (n_4792), .A1 (n_5016), .B0 (n_5121), .Y(n_5438));
AOI21X1 g131153(.A0 (n_5121), .A1 (n_4978), .B0 (n_5120), .Y(n_5351));
NAND3X1 g131195(.A (n_4868), .B (n_4642), .C (n_4307), .Y (n_5119));
INVX1 g131212(.A (n_5273), .Y (n_5118));
XOR2X1 g131258(.A (n_1684), .B (n_4948), .Y (n_5117));
XOR2X1 g131268(.A (n_1774), .B (n_4847), .Y (n_5116));
NOR2X1 g131564(.A (n_5188), .B (n_1250), .Y (n_5115));
AOI22X1 g131653(.A0 (n_4778), .A1 (n_4777), .B0 (n_5113), .B1(n_2178), .Y (n_5114));
XOR2X1 g131672(.A (n_714), .B (n_4628), .Y (n_5112));
OAI21X1 g131692(.A0 (n_4832), .A1 (n_5110), .B0 (n_5109), .Y(n_5111));
OAI21X1 g131693(.A0 (n_4829), .A1 (n_5107), .B0 (n_5106), .Y(n_5108));
NAND3X1 g131767(.A (n_34505), .B (n_4619), .C (n_34506), .Y (n_5105));
AOI21X1 g131793(.A0 (n_4810), .A1 (n_5022), .B0 (n_5104), .Y(n_5173));
INVX1 g131884(.A (n_33586), .Y (n_6055));
INVX1 g131897(.A (n_6069), .Y (n_5161));
OAI21X1 g131903(.A0 (n_5101), .A1 (n_5100), .B0 (n_5099), .Y(n_5427));
OAI21X1 g131904(.A0 (n_5098), .A1 (n_2428), .B0 (n_5096), .Y(n_5545));
OAI21X1 g131905(.A0 (n_5095), .A1 (n_5094), .B0 (n_5093), .Y(n_5302));
AND2X1 g131929(.A (n_5091), .B (n_5090), .Y (n_5092));
NOR2X1 g131957(.A (n_5240), .B (n_4867), .Y (n_5590));
NAND2X1 g131979(.A (n_5643), .B (n_5089), .Y (n_5469));
NOR2X1 g131987(.A (n_5305), .B (n_4933), .Y (n_5419));
NAND3X1 g132002(.A (n_4890), .B (n_4236), .C (n_4728), .Y (n_5088));
AND2X1 g132016(.A (n_5086), .B (n_5085), .Y (n_5087));
NOR2X1 g132027(.A (n_5226), .B (n_4791), .Y (n_5547));
AND2X1 g132047(.A (n_5083), .B (n_5129), .Y (n_5084));
NOR2X1 g132050(.A (n_5132), .B (n_4193), .Y (n_5082));
NAND3X1 g132054(.A (n_4746), .B (n_4083), .C (n_4794), .Y (n_5081));
INVX1 g132068(.A (n_5079), .Y (n_5080));
INVX1 g132071(.A (n_5077), .Y (n_5078));
AOI21X1 g132077(.A0 (n_5076), .A1 (n_4787), .B0 (n_5075), .Y(n_5431));
AOI21X1 g132087(.A0 (n_5063), .A1 (n_5075), .B0 (n_4975), .Y(n_5290));
AOI21X1 g132089(.A0 (n_4615), .A1 (n_4919), .B0 (n_5074), .Y(n_5429));
AOI21X1 g132099(.A0 (n_5215), .A1 (n_5072), .B0 (n_5073), .Y(n_5421));
AOI21X1 g132100(.A0 (n_5160), .A1 (n_4774), .B0 (n_5072), .Y(n_5443));
OAI21X1 g132111(.A0 (n_4609), .A1 (n_4961), .B0 (n_4972), .Y(n_5411));
OAI21X1 g132121(.A0 (n_4987), .A1 (n_5070), .B0 (n_5071), .Y(n_5409));
OAI21X1 g132130(.A0 (n_4544), .A1 (n_4959), .B0 (n_5070), .Y(n_5414));
XOR2X1 g132175(.A (n_13724), .B (n_4720), .Y (n_6298));
INVX1 g132197(.A (n_35400), .Y (n_32219));
OR2X1 g132253(.A (n_5387), .B (n_5215), .Y (n_5065));
INVX1 g132258(.A (n_5225), .Y (n_5064));
NAND2X1 g132266(.A (n_5063), .B (n_5384), .Y (n_5580));
NAND2X1 g132273(.A (n_4663), .B (n_5061), .Y (n_5062));
INVX1 g132280(.A (n_5236), .Y (n_5060));
INVX1 g132291(.A (n_5278), .Y (n_5059));
NOR2X1 g132293(.A (n_5073), .B (n_5072), .Y (n_5570));
INVX1 g132321(.A (n_5055), .Y (n_5211));
NAND2X1 g132353(.A (n_4726), .B (n_5053), .Y (n_5054));
NOR2X1 g132355(.A (n_5052), .B (n_4536), .Y (n_5344));
INVX1 g132362(.A (n_5235), .Y (n_5051));
NOR2X1 g132378(.A (n_4737), .B (n_5216), .Y (n_5050));
NAND2X1 g132385(.A (n_4756), .B (n_5049), .Y (n_5390));
INVX1 g132393(.A (n_5276), .Y (n_5048));
NOR2X1 g132404(.A (n_4741), .B (n_4973), .Y (n_5047));
NOR2X1 g132420(.A (n_5046), .B (n_4548), .Y (n_5325));
NAND2X1 g132422(.A (n_5231), .B (n_5049), .Y (n_5348));
INVX1 g132424(.A (n_5197), .Y (n_5045));
NAND2X1 g132434(.A (n_4825), .B (n_4824), .Y (n_5538));
NOR2X1 g132448(.A (n_5387), .B (n_5073), .Y (n_5327));
NAND2X1 g132492(.A (n_4733), .B (n_5044), .Y (n_5524));
NAND2X1 g132493(.A (n_4719), .B (n_5043), .Y (n_5507));
XOR2X1 g132589(.A (n_4028), .B (n_5041), .Y (n_5042));
NOR2X1 g132695(.A (n_4769), .B (n_5033), .Y (n_5039));
INVX1 g132742(.A (n_5204), .Y (n_5038));
NAND2X1 g132765(.A (n_5034), .B (n_4722), .Y (n_5037));
INVX1 g132306(.A (n_5056), .Y (n_5035));
OAI21X1 g132552(.A0 (n_4298), .A1 (n_4884), .B0 (n_5034), .Y(n_5368));
OAI21X1 g132549(.A0 (n_5032), .A1 (n_4885), .B0 (n_4714), .Y(n_5370));
OAI21X1 g131836(.A0 (n_4859), .A1 (n_5085), .B0 (n_4375), .Y(n_5244));
OAI21X1 g132543(.A0 (n_4242), .A1 (n_5033), .B0 (n_5032), .Y(n_5445));
OAI21X1 g132539(.A0 (n_5034), .A1 (n_4883), .B0 (n_4789), .Y(n_5366));
NAND2X1 g132811(.A (n_5156), .B (n_4572), .Y (n_5031));
INVX1 g132263(.A (n_5139), .Y (n_5030));
NOR2X1 g132262(.A (n_5072), .B (n_4742), .Y (n_6071));
XOR2X1 g131659(.A (n_1698), .B (n_5028), .Y (n_5029));
INVX1 g132780(.A (n_5206), .Y (n_5027));
NAND2X1 g131383(.A (n_4692), .B (n_4681), .Y (n_5503));
NAND2X1 g132251(.A (n_4825), .B (n_4920), .Y (n_5535));
OR2X1 g132250(.A (n_5519), .B (n_5063), .Y (n_5024));
INVX1 g132228(.A (n_5444), .Y (n_5341));
NOR2X1 g132218(.A (n_4772), .B (P3_reg1[15] ), .Y (n_5484));
NAND2X1 g131432(.A (n_5176), .B (n_5146), .Y (n_5350));
NAND2X1 g132004(.A (n_5022), .B (n_5167), .Y (n_5180));
NAND2X1 g132496(.A (n_4740), .B (n_5021), .Y (n_5320));
AND2X1 g131989(.A (n_5131), .B (n_4766), .Y (n_5855));
NAND2X1 g132223(.A (n_4772), .B (P3_reg1[15] ), .Y (n_5628));
NOR2X1 g131978(.A (n_4901), .B (n_4426), .Y (n_6059));
NAND2X1 g131207(.A (n_4698), .B (n_5016), .Y (n_5017));
INVX1 g132177(.A (n_34388), .Y (n_5015));
OAI21X1 g131115(.A0 (n_5014), .A1 (n_5013), .B0 (n_5012), .Y(n_5354));
AOI21X1 g132105(.A0 (n_4669), .A1 (n_4808), .B0 (n_5011), .Y(n_5425));
AOI21X1 g131789(.A0 (n_4840), .A1 (n_5010), .B0 (n_5009), .Y(n_5249));
XOR2X1 g131369(.A (n_1851), .B (n_4550), .Y (n_5008));
XOR2X1 g131664(.A (n_1655), .B (n_5006), .Y (n_5007));
INVX1 g132407(.A (n_5005), .Y (n_5564));
INVX1 g132405(.A (n_5193), .Y (n_5004));
OAI21X1 g132590(.A0 (n_5002), .A1 (n_4891), .B0 (n_4738), .Y(n_5003));
NOR2X1 g131960(.A (n_5091), .B (n_4902), .Y (n_5001));
NAND2X1 g132388(.A (n_5404), .B (n_5053), .Y (n_5379));
INVX1 g132443(.A (n_5227), .Y (n_5000));
OAI21X1 g132132(.A0 (n_4592), .A1 (n_4774), .B0 (n_4915), .Y(n_5343));
XOR2X1 g132163(.A (P1_reg1[19] ), .B (n_6208), .Y (n_4998));
INVX1 g132699(.A (n_5213), .Y (n_4997));
INVX1 g132148(.A (n_34920), .Y (n_5219));
XOR2X1 g131500(.A (n_1170), .B (n_4486), .Y (n_4994));
NOR2X1 g131322(.A (n_4491), .B (n_5123), .Y (n_5502));
NAND2X1 g132423(.A (n_5215), .B (n_5089), .Y (n_5576));
XOR2X1 g131360(.A (n_1480), .B (n_4533), .Y (n_4993));
OAI21X1 g131442(.A0 (n_2846), .A1 (n_4341), .B0 (n_4776), .Y(n_4992));
NOR2X1 g131740(.A (n_6375), .B (n_4990), .Y (n_4991));
INVX1 g131300(.A (n_5159), .Y (n_4989));
NOR2X1 g132429(.A (n_4739), .B (n_4987), .Y (n_4988));
OAI21X1 g131912(.A0 (n_4986), .A1 (n_4985), .B0 (n_4984), .Y(n_5470));
OAI21X1 g132129(.A0 (n_4750), .A1 (n_4983), .B0 (n_4982), .Y(n_5405));
AND2X1 g131428(.A (n_4980), .B (n_5272), .Y (n_4981));
NAND2X1 g131410(.A (n_5146), .B (n_4978), .Y (n_5450));
NOR2X1 g131947(.A (n_4262), .B (n_4976), .Y (n_4977));
OAI21X1 g132123(.A0 (n_4975), .A1 (n_5076), .B0 (n_5063), .Y(n_5332));
NOR2X1 g132376(.A (n_5075), .B (n_4706), .Y (n_5998));
OAI21X1 g132115(.A0 (n_4912), .A1 (n_4971), .B0 (n_4801), .Y(n_5556));
OAI21X1 g132124(.A0 (n_4612), .A1 (n_4862), .B0 (n_5061), .Y(n_5285));
INVX1 g132402(.A (n_5353), .Y (n_4974));
OAI21X1 g132112(.A0 (n_4973), .A1 (n_4972), .B0 (n_4971), .Y(n_5337));
NAND3X1 g132108(.A (n_4655), .B (n_4364), .C (n_4833), .Y (n_5455));
AOI21X1 g132086(.A0 (n_4643), .A1 (n_4913), .B0 (n_4969), .Y(n_4970));
NAND3X1 g131218(.A (n_4967), .B (n_4783), .C (n_4111), .Y (n_4968));
XOR2X1 g131848(.A (n_4150), .B (n_4965), .Y (n_4966));
NOR2X1 g132370(.A (n_5519), .B (n_4975), .Y (n_5346));
INVX1 g132359(.A (n_5238), .Y (n_4963));
NOR2X1 g132339(.A (n_4961), .B (n_4732), .Y (n_4962));
NOR2X1 g132256(.A (n_4959), .B (n_4693), .Y (n_4960));
NOR2X1 g132242(.A (n_4772), .B (P3_reg2[15] ), .Y (n_5410));
NOR2X1 g131937(.A (n_5198), .B (n_4928), .Y (n_5420));
NAND2X1 g132494(.A (n_4734), .B (n_4957), .Y (n_5532));
NOR2X1 g132057(.A (n_5442), .B (n_4860), .Y (n_5475));
NOR2X1 g132380(.A (n_4905), .B (n_4774), .Y (n_5331));
NAND2X1 g132261(.A (n_4921), .B (n_4481), .Y (n_5712));
XOR2X1 g131668(.A (n_2184), .B (n_4451), .Y (n_4956));
OAI21X1 g131918(.A0 (n_4955), .A1 (n_4954), .B0 (n_4953), .Y(n_5282));
NOR2X1 g132775(.A (n_4243), .B (n_5033), .Y (n_5171));
NAND2X1 g132069(.A (n_35090), .B (n_35621), .Y (n_5079));
NAND2X1 g131224(.A (n_5016), .B (n_4694), .Y (n_5436));
NAND4X1 g131248(.A (n_4948), .B (n_3785), .C (n_1796), .D (n_4280),.Y (n_4949));
AOI21X1 g131445(.A0 (n_5586), .A1 (n_4947), .B0 (n_4946), .Y(n_5310));
INVX1 g131553(.A (n_5271), .Y (n_4945));
NAND2X1 g131558(.A (n_4817), .B (n_9663), .Y (n_5149));
XOR2X1 g131670(.A (n_1362), .B (n_4449), .Y (n_4944));
NAND2X1 g131688(.A (n_4942), .B (n_4357), .Y (n_4943));
NAND2X1 g131748(.A (n_5113), .B (n_748), .Y (n_4941));
NAND3X1 g131813(.A (n_4581), .B (n_4940), .C (n_4617), .Y (n_5200));
OAI22X1 g131845(.A0 (n_4938), .A1 (n_4937), .B0 (n_4442), .B1(n_696), .Y (n_4939));
NOR2X1 g131983(.A (n_4007), .B (n_34118), .Y (n_4936));
NOR2X1 g131985(.A (n_5277), .B (n_5046), .Y (n_4935));
AND2X1 g132014(.A (n_4934), .B (n_6017), .Y (n_6278));
NOR2X1 g132022(.A (n_4933), .B (n_4932), .Y (n_5417));
NOR2X1 g132067(.A (n_34237), .B (n_4618), .Y (n_4931));
NAND2X1 g132074(.A (n_4212), .B (n_4580), .Y (n_4930));
NOR3X1 g132078(.A (n_4040), .B (n_4271), .C (n_4579), .Y (n_5259));
NAND3X1 g132109(.A (n_4532), .B (n_4422), .C (n_4830), .Y (n_5322));
OAI21X1 g132330(.A0 (n_4568), .A1 (n_4448), .B0 (n_4626), .Y(n_5377));
OAI21X1 g132131(.A0 (n_4929), .A1 (n_4928), .B0 (n_4927), .Y(n_5568));
NAND2X1 g132203(.A (n_4530), .B (n_4926), .Y (n_5355));
OAI21X1 g132208(.A0 (n_4925), .A1 (n_2460), .B0 (n_4924), .Y(n_5396));
NOR2X1 g132219(.A (n_32388), .B (P3_reg1[16] ), .Y (n_5539));
NAND2X1 g132229(.A (n_32388), .B (P3_reg1[16] ), .Y (n_5444));
OR2X1 g132246(.A (n_4921), .B (n_5075), .Y (n_4922));
NOR2X1 g132259(.A (n_4825), .B (n_4920), .Y (n_5225));
NAND2X1 g132264(.A (n_4616), .B (n_4919), .Y (n_5139));
NOR2X1 g132276(.A (n_4796), .B (n_4917), .Y (n_4918));
NAND2X1 g132281(.A (n_5215), .B (n_5160), .Y (n_5236));
NOR2X1 g132289(.A (n_4594), .B (n_4928), .Y (n_4916));
NAND2X1 g132312(.A (n_4915), .B (n_5160), .Y (n_5292));
NAND2X1 g132313(.A (n_4644), .B (n_4913), .Y (n_4914));
NOR2X1 g132323(.A (n_5072), .B (n_4774), .Y (n_5326));
NOR2X1 g132328(.A (n_4912), .B (n_4973), .Y (n_5563));
NOR2X1 g132333(.A (n_4911), .B (P2_reg1[15] ), .Y (n_5335));
NOR2X1 g132342(.A (n_4597), .B (n_4909), .Y (n_4910));
NOR2X1 g132374(.A (n_4598), .B (n_4907), .Y (n_4908));
INVX1 g132382(.A (n_4976), .Y (n_4906));
NAND2X1 g132390(.A (n_4921), .B (n_5076), .Y (n_5388));
NOR2X1 g132717(.A (n_4905), .B (n_4547), .Y (n_6062));
OR2X1 g132392(.A (n_4915), .B (n_5072), .Y (n_4904));
NAND2X1 g132403(.A (n_4911), .B (P2_reg1[15] ), .Y (n_5353));
NAND2X1 g132406(.A (n_5169), .B (n_4919), .Y (n_5193));
NOR2X1 g132412(.A (n_4961), .B (n_4973), .Y (n_5274));
NOR2X1 g132415(.A (n_4983), .B (n_5185), .Y (n_5543));
NOR2X1 g132426(.A (n_4611), .B (n_4961), .Y (n_5412));
NOR2X1 g132428(.A (n_4596), .B (n_4902), .Y (n_4903));
NAND2X1 g132451(.A (n_4557), .B (n_4900), .Y (n_5299));
NAND2X1 g132452(.A (n_4524), .B (n_4899), .Y (n_5241));
NAND2X1 g132072(.A (n_4521), .B (n_4515), .Y (n_5077));
AOI21X1 g132517(.A0 (n_4431), .A1 (n_4753), .B0 (n_4846), .Y(n_5142));
AOI21X1 g132518(.A0 (n_4424), .A1 (n_4718), .B0 (n_4864), .Y(n_5151));
OAI21X1 g132532(.A0 (n_4882), .A1 (n_4431), .B0 (n_4593), .Y(n_5178));
OAI21X1 g132540(.A0 (n_4905), .A1 (n_4424), .B0 (n_4592), .Y(n_5168));
OAI21X1 g132545(.A0 (n_4895), .A1 (n_4727), .B0 (n_4752), .Y(n_5280));
OAI21X1 g132548(.A0 (n_4674), .A1 (n_4798), .B0 (n_4754), .Y(n_5222));
OAI21X1 g132553(.A0 (n_4148), .A1 (n_4870), .B0 (n_4895), .Y(n_5223));
XOR2X1 g132575(.A (n_3997), .B (n_4893), .Y (n_4894));
XOR2X1 g132576(.A (n_4891), .B (n_4890), .Y (n_4892));
OAI21X1 g132581(.A0 (n_4888), .A1 (n_4747), .B0 (n_4586), .Y(n_4889));
NOR2X1 g132319(.A (n_4546), .B (n_4959), .Y (n_5415));
INVX1 g132681(.A (n_5089), .Y (n_5127));
XOR2X1 g132940(.A (n_4647), .B (n_4391), .Y (n_4887));
NOR2X1 g132743(.A (n_4385), .B (n_75), .Y (n_5204));
NOR2X1 g132760(.A (n_4629), .B (n_4675), .Y (n_4886));
NOR2X1 g132761(.A (n_5033), .B (n_4885), .Y (n_5371));
NOR2X1 g132840(.A (n_4884), .B (n_4883), .Y (n_5367));
NOR2X1 g132856(.A (n_4882), .B (n_4541), .Y (n_6023));
AOI21X1 g131486(.A0 (n_4463), .A1 (n_2146), .B0 (n_4323), .Y(n_4881));
OAI21X1 g132311(.A0 (n_4570), .A1 (n_4359), .B0 (n_4553), .Y(n_5382));
NAND2X1 g132290(.A (n_5155), .B (n_4388), .Y (n_4880));
NAND2X1 g132307(.A (n_4764), .B (P2_reg2[16] ), .Y (n_5056));
NOR2X1 g132066(.A (n_4509), .B (n_4749), .Y (n_4877));
NOR2X1 g132294(.A (n_4959), .B (n_4987), .Y (n_5230));
NOR2X1 g132347(.A (n_4585), .B (n_4912), .Y (n_4874));
NAND2X1 g131530(.A (n_4498), .B (n_4978), .Y (n_4873));
NAND2X1 g132292(.A (n_5275), .B (n_4872), .Y (n_5278));
NOR2X1 g132824(.A (n_4476), .B (n_4870), .Y (n_4871));
NOR2X1 g132284(.A (n_4751), .B (n_4983), .Y (n_5406));
XOR2X1 g131367(.A (n_3939), .B (n_4868), .Y (so[5]));
NOR2X1 g132042(.A (n_4867), .B (n_4902), .Y (n_5857));
INVX1 g132829(.A (n_4982), .Y (n_4866));
NOR2X1 g132790(.A (n_4299), .B (n_4884), .Y (n_5199));
XOR2X1 g131479(.A (n_496), .B (n_4360), .Y (n_4865));
NOR2X1 g132781(.A (n_33034), .B (P1_reg1[14] ), .Y (n_5206));
NOR2X1 g132800(.A (n_4382), .B (n_4864), .Y (n_5867));
INVX1 g132243(.A (n_4863), .Y (n_5566));
NOR2X1 g132252(.A (n_4862), .B (n_4861), .Y (n_5541));
NOR2X1 g132029(.A (n_4860), .B (n_4859), .Y (n_5548));
NOR2X1 g132764(.A (n_33034), .B (P1_reg2[14] ), .Y (n_5593));
OAI22X1 g131844(.A0 (n_4856), .A1 (n_4855), .B0 (n_4417), .B1(n_1373), .Y (n_4857));
NAND2X1 g132237(.A (n_32388), .B (n_13507), .Y (n_5023));
OAI22X1 g131488(.A0 (n_4853), .A1 (n_4852), .B0 (n_4851), .B1(n_611), .Y (n_4854));
NOR2X1 g132221(.A (n_32388), .B (n_13507), .Y (n_5644));
NAND3X1 g131307(.A (n_4847), .B (n_1903), .C (n_3250), .Y (n_4848));
NOR2X1 g132696(.A (n_4381), .B (n_4846), .Y (n_5870));
NAND2X1 g132205(.A (n_4429), .B (n_4845), .Y (n_5530));
INVX1 g132193(.A (n_4990), .Y (n_5067));
AOI21X1 g131456(.A0 (n_4073), .A1 (n_1223), .B0 (n_4636), .Y(n_4842));
NOR2X1 g131301(.A (n_5013), .B (n_4785), .Y (n_5159));
AND2X1 g131966(.A (n_5925), .B (n_5946), .Y (n_6276));
AOI21X1 g132103(.A0 (n_4576), .A1 (n_4835), .B0 (n_4840), .Y(n_4841));
INVX1 g133219(.A (n_5220), .Y (n_4839));
NAND2X1 g132444(.A (n_5252), .B (n_4913), .Y (n_5227));
AND2X1 g132322(.A (n_4764), .B (P2_reg1[16] ), .Y (n_5055));
NAND2X1 g132425(.A (n_4911), .B (P2_reg2[15] ), .Y (n_5197));
NOR2X1 g132700(.A (n_4385), .B (n_230), .Y (n_5213));
NOR2X1 g131928(.A (n_5237), .B (n_5052), .Y (n_4836));
NAND2X1 g132408(.A (n_5010), .B (n_4835), .Y (n_5005));
INVX1 g132683(.A (n_5384), .Y (n_4834));
OAI21X1 g131917(.A0 (n_4833), .A1 (n_4821), .B0 (n_4832), .Y(n_5135));
OAI21X1 g132136(.A0 (n_4593), .A1 (n_4787), .B0 (n_4921), .Y(n_5248));
OAI21X1 g131916(.A0 (n_4830), .A1 (n_4806), .B0 (n_4829), .Y(n_5253));
OAI21X1 g131913(.A0 (n_4828), .A1 (n_2076), .B0 (n_4826), .Y(n_5432));
NOR2X1 g132417(.A (n_4825), .B (n_4824), .Y (n_5493));
NAND2X1 g131213(.A (n_4814), .B (n_9658), .Y (n_5273));
INVX1 g131556(.A (n_5203), .Y (n_4823));
NOR2X1 g132350(.A (n_5110), .B (n_4821), .Y (n_4822));
NAND2X1 g131683(.A (n_34434), .B (n_4326), .Y (n_4820));
INVX1 g131538(.A (n_4980), .Y (n_4818));
OR2X1 g131531(.A (n_4817), .B (n_9663), .Y (n_5144));
NAND3X1 g131550(.A (n_2997), .B (n_4443), .C (n_3609), .Y (n_4815));
NOR2X1 g131222(.A (n_4814), .B (n_9658), .Y (n_5437));
NAND2X1 g131225(.A (n_4978), .B (n_5016), .Y (n_5312));
XOR2X1 g131671(.A (n_1482), .B (n_4470), .Y (n_4813));
NAND4X1 g131770(.A (n_35254), .B (n_4511), .C (n_32394), .D(n_32021), .Y (n_4812));
AOI21X1 g132107(.A0 (n_4494), .A1 (n_4703), .B0 (n_4810), .Y(n_4811));
NAND2X1 g132360(.A (n_4700), .B (n_4872), .Y (n_5238));
INVX1 g132189(.A (n_6256), .Y (n_6255));
NOR2X1 g132386(.A (n_5075), .B (n_4787), .Y (n_5345));
NOR2X1 g132367(.A (n_4975), .B (n_5075), .Y (n_5333));
NAND2X1 g132363(.A (n_5179), .B (n_4808), .Y (n_5235));
NOR2X1 g132351(.A (n_5107), .B (n_4806), .Y (n_4807));
NAND2X1 g132304(.A (n_4350), .B (n_5063), .Y (n_6117));
AOI21X1 g132288(.A0 (n_3463), .A1 (n_4805), .B0 (n_4804), .Y(n_5398));
NOR2X1 g132265(.A (n_4657), .B (n_4802), .Y (n_4803));
NOR2X1 g132379(.A (n_4711), .B (n_4862), .Y (n_5286));
NAND2X1 g132394(.A (n_5063), .B (n_5076), .Y (n_5276));
OAI21X1 g132119(.A0 (n_4801), .A1 (n_4909), .B0 (n_4800), .Y(n_5457));
NOR2X1 g132740(.A (n_4384), .B (n_4798), .Y (n_4799));
INVX1 g132885(.A (n_4796), .Y (n_4797));
NOR2X1 g131712(.A (n_4792), .B (n_4452), .Y (n_4793));
INVX1 g132364(.A (n_4791), .Y (n_5131));
NAND2X1 g133222(.A (n_4789), .B (n_4394), .Y (n_4790));
NOR2X1 g132356(.A (n_4907), .B (n_4928), .Y (n_5315));
NOR2X1 g131560(.A (n_4851), .B (n_2989), .Y (n_4788));
NOR2X1 g132377(.A (n_4362), .B (n_4932), .Y (n_6301));
AOI21X1 g132098(.A0 (n_4882), .A1 (n_4921), .B0 (n_4787), .Y(n_5291));
NAND2X1 g133220(.A (n_4010), .B (n_4445), .Y (n_5220));
OR2X1 g131320(.A (n_4641), .B (n_4785), .Y (n_4786));
XOR2X1 g131489(.A (n_698), .B (n_4297), .Y (n_4782));
OR2X1 g131539(.A (n_4665), .B (n_9675), .Y (n_4980));
INVX1 g131675(.A (n_4780), .Y (n_4781));
NAND2X1 g132830(.A (n_4535), .B (n_4590), .Y (n_4982));
NOR2X1 g131734(.A (n_4778), .B (n_4777), .Y (n_4779));
NAND3X1 g131651(.A (n_4343), .B (n_2844), .C (n_4024), .Y (n_4776));
NOR2X1 g132070(.A (n_4514), .B (n_4415), .Y (n_33009));
AOI21X1 g132082(.A0 (n_4905), .A1 (n_4915), .B0 (n_4774), .Y(n_5423));
NAND2X1 g133199(.A (n_4010), .B (P1_reg1[12] ), .Y (n_5156));
INVX1 g132183(.A (n_33583), .Y (n_35105));
NAND2X1 g132220(.A (n_4772), .B (P3_reg2[15] ), .Y (n_5643));
AOI21X1 g132245(.A0 (n_3467), .A1 (n_4771), .B0 (n_4770), .Y(n_5296));
NOR2X1 g132269(.A (n_4882), .B (n_4787), .Y (n_5167));
INVX1 g133191(.A (n_5032), .Y (n_4769));
NAND2X1 g132283(.A (n_4767), .B (n_4766), .Y (n_4768));
NOR2X1 g132308(.A (n_4911), .B (P2_reg2[15] ), .Y (n_5198));
NOR2X1 g132373(.A (n_4376), .B (n_4859), .Y (n_6351));
NAND2X1 g132383(.A (n_4670), .B (n_4808), .Y (n_4976));
NOR2X1 g132399(.A (n_4764), .B (P2_reg1[16] ), .Y (n_5442));
NOR2X1 g132401(.A (n_4402), .B (n_4821), .Y (n_5136));
NOR2X1 g132430(.A (n_4764), .B (P2_reg2[16] ), .Y (n_5305));
NOR2X1 g132791(.A (n_4731), .B (P1_reg1[16] ), .Y (n_5226));
NAND2X1 g132466(.A (n_32642), .B (n_4006), .Y (n_4762));
INVX1 g132479(.A (n_34118), .Y (n_4759));
NOR2X1 g132488(.A (n_33174), .B (n_35391), .Y (n_4757));
AOI21X1 g132506(.A0 (n_4578), .A1 (n_4756), .B0 (n_4755), .Y(n_4984));
OAI21X1 g132531(.A0 (n_4789), .A1 (n_4600), .B0 (n_4613), .Y(n_5287));
OAI21X1 g132537(.A0 (n_4754), .A1 (n_4555), .B0 (n_4610), .Y(n_5251));
OAI21X1 g132547(.A0 (n_4753), .A1 (n_4377), .B0 (n_4430), .Y(n_5011));
OAI21X1 g132551(.A0 (n_4752), .A1 (n_4378), .B0 (n_4545), .Y(n_5403));
OAI21X1 g132554(.A0 (n_4751), .A1 (n_4713), .B0 (n_4750), .Y(n_5485));
NOR2X1 g132073(.A (n_4749), .B (n_32023), .Y (n_5260));
XOR2X1 g132567(.A (n_4747), .B (n_4746), .Y (n_4748));
XOR2X1 g132568(.A (n_4058), .B (n_4744), .Y (n_4745));
XOR2X1 g132569(.A (n_4054), .B (n_5095), .Y (n_4743));
NOR2X1 g132672(.A (n_4701), .B (n_13338), .Y (n_5387));
INVX1 g132673(.A (n_5160), .Y (n_4742));
NOR2X1 g132689(.A (n_4753), .B (n_4405), .Y (n_5612));
INVX1 g132701(.A (n_4971), .Y (n_4741));
NAND2X1 g132705(.A (n_6044), .B (n_4559), .Y (n_4740));
INVX1 g132706(.A (n_5071), .Y (n_4739));
NAND2X1 g132714(.A (n_5002), .B (n_4891), .Y (n_4738));
INVX1 g132730(.A (n_5221), .Y (n_4737));
NAND2X1 g132796(.A (n_5956), .B (n_4496), .Y (n_4734));
NAND2X1 g132802(.A (n_5972), .B (n_4562), .Y (n_4733));
INVX1 g132805(.A (n_4972), .Y (n_4732));
NOR2X1 g132809(.A (n_4731), .B (P1_reg2[16] ), .Y (n_5240));
NAND2X1 g132812(.A (n_4750), .B (n_4339), .Y (n_4730));
NOR2X1 g132827(.A (n_4870), .B (n_4727), .Y (n_5049));
NOR2X1 g132834(.A (n_4185), .B (n_4870), .Y (n_5053));
AOI21X1 g132890(.A0 (n_4651), .A1 (n_4726), .B0 (n_4725), .Y(n_5044));
INVX1 g132974(.A (n_4764), .Y (n_4724));
INVX1 g133046(.A (n_4723), .Y (n_6802));
INVX1 g133139(.A (n_4884), .Y (n_4722));
NAND3X1 g131589(.A (n_4466), .B (n_4206), .C (n_4504), .Y (n_4967));
NOR2X1 g133205(.A (n_4436), .B (n_4885), .Y (n_4721));
INVX1 g132964(.A (n_4720), .Y (n_4844));
NAND2X1 g132835(.A (n_5914), .B (n_4565), .Y (n_4719));
OAI21X1 g132544(.A0 (n_4718), .A1 (n_4614), .B0 (n_4423), .Y(n_5074));
INVX1 g132606(.A (n_33173), .Y (n_6231));
NOR2X1 g132282(.A (n_4907), .B (n_4987), .Y (n_5479));
OAI21X1 g132538(.A0 (n_4864), .A1 (n_4423), .B0 (n_4424), .Y(n_5009));
INVX1 g132278(.A (n_4933), .Y (n_5083));
NAND2X1 g132848(.A (n_4535), .B (n_4534), .Y (n_5061));
OAI21X1 g132534(.A0 (n_4714), .A1 (n_4537), .B0 (n_4713), .Y(n_5407));
NOR2X1 g132808(.A (n_4708), .B (n_4404), .Y (n_5393));
NOR2X1 g132807(.A (n_4392), .B (n_4711), .Y (n_4712));
OR2X1 g132366(.A (n_4437), .B (n_4536), .Y (n_4710));
NOR2X1 g132267(.A (n_4912), .B (n_4909), .Y (n_5458));
AOI21X1 g132510(.A0 (n_4075), .A1 (n_4377), .B0 (n_4708), .Y(n_5143));
AOI21X1 g132519(.A0 (n_4592), .A1 (n_4864), .B0 (n_4905), .Y(n_5109));
NOR2X1 g132798(.A (n_4462), .B (n_4727), .Y (n_4707));
INVX1 g132658(.A (n_5076), .Y (n_4706));
OAI21X1 g132546(.A0 (n_4846), .A1 (n_4430), .B0 (n_4431), .Y(n_5104));
NAND2X1 g132244(.A (n_5022), .B (n_4703), .Y (n_4863));
INVX1 g132247(.A (n_4860), .Y (n_5086));
NAND2X1 g132684(.A (n_4701), .B (n_13679), .Y (n_5384));
AOI21X1 g132507(.A0 (n_4493), .A1 (n_4700), .B0 (n_4699), .Y(n_5093));
INVX1 g132232(.A (n_4934), .Y (n_4923));
INVX1 g131308(.A (n_5121), .Y (n_4698));
XOR2X1 g132585(.A (n_4223), .B (n_4986), .Y (n_4697));
NOR2X1 g132615(.A (n_4154), .B (n_4029), .Y (n_4696));
AOI21X1 g132497(.A0 (n_4593), .A1 (n_4846), .B0 (n_4882), .Y(n_5106));
NOR2X1 g132484(.A (n_4354), .B (n_4653), .Y (n_5175));
NOR2X1 g132686(.A (n_4718), .B (n_4386), .Y (n_5609));
NAND3X1 g131798(.A (n_3089), .B (n_4281), .C (n_3603), .Y (n_4695));
NAND2X1 g132194(.A (n_2203), .B (n_4372), .Y (n_4990));
AOI21X1 g131629(.A0 (n_4684), .A1 (n_4694), .B0 (n_4792), .Y(n_5122));
INVX1 g132711(.A (n_5070), .Y (n_4693));
INVX1 g131618(.A (n_4505), .Y (n_4692));
NOR2X1 g132445(.A (n_5216), .B (n_5185), .Y (n_5571));
NAND3X1 g131501(.A (n_2972), .B (n_4295), .C (n_4270), .Y (n_4689));
INVX1 g132158(.A (n_34947), .Y (n_4688));
NOR2X1 g131764(.A (n_4684), .B (n_4450), .Y (n_4685));
OR2X1 g131315(.A (n_4681), .B (n_4491), .Y (n_4682));
NOR2X1 g132675(.A (n_4701), .B (n_13679), .Y (n_5519));
INVX1 g132413(.A (n_4867), .Y (n_5090));
NAND2X1 g131573(.A (n_4677), .B (n_9672), .Y (n_5146));
NAND2X1 g132682(.A (n_4701), .B (n_13338), .Y (n_5089));
AOI21X1 g131687(.A0 (n_4165), .A1 (n_4179), .B0 (n_3792), .Y(n_5188));
NOR2X1 g132395(.A (n_4420), .B (n_4806), .Y (n_5254));
NOR2X1 g131557(.A (n_4677), .B (n_9672), .Y (n_5203));
NOR2X1 g131554(.A (n_4668), .B (n_9667), .Y (n_5271));
OAI21X1 g132541(.A0 (n_4251), .A1 (n_4675), .B0 (n_4674), .Y(n_4969));
AOI21X1 g131611(.A0 (n_4519), .A1 (n_4488), .B0 (n_4684), .Y(n_5012));
OR2X1 g132352(.A (n_4605), .B (n_4548), .Y (n_4671));
NAND2X1 g132397(.A (n_4478), .B (n_4477), .Y (n_5132));
AOI21X1 g132521(.A0 (n_4459), .A1 (n_4670), .B0 (n_4669), .Y(n_5099));
NAND2X1 g131575(.A (n_4668), .B (n_9667), .Y (n_5176));
INVX1 g133021(.A (n_33175), .Y (n_6246));
XOR2X1 g131252(.A (n_1184), .B (n_4645), .Y (n_4666));
NAND2X1 g131577(.A (n_4665), .B (n_9675), .Y (n_5272));
INVX1 g132757(.A (n_4862), .Y (n_4663));
INVX1 g132437(.A (n_33250), .Y (n_4901));
NOR2X1 g132418(.A (n_5157), .B (n_4861), .Y (n_5489));
NAND2X1 g132411(.A (n_4478), .B (n_11141), .Y (n_5091));
INVX1 g132887(.A (n_4657), .Y (n_4658));
INVX1 g132190(.A (n_4656), .Y (n_6256));
NAND2X1 g132751(.A (n_4409), .B (n_4403), .Y (n_4655));
NAND2X1 g132296(.A (n_4915), .B (n_4602), .Y (n_5872));
NAND2X1 g132336(.A (n_4577), .B (n_4835), .Y (n_4654));
NAND2X1 g131950(.A (n_5946), .B (n_5951), .Y (n_5659));
NAND2X1 g132110(.A (n_4283), .B (n_2811), .Y (n_5113));
INVX1 g133047(.A (n_4653), .Y (n_4723));
NOR2X1 g133228(.A (n_35368), .B (n_4561), .Y (n_5033));
NAND2X1 g132324(.A (n_4495), .B (n_4703), .Y (n_4652));
AOI21X1 g133275(.A0 (n_5972), .A1 (n_4347), .B0 (n_4651), .Y(n_5041));
AOI21X1 g132898(.A0 (n_4254), .A1 (n_4650), .B0 (n_4649), .Y(n_4957));
XOR2X1 g132933(.A (n_4531), .B (n_4647), .Y (n_4648));
NAND3X1 g132886(.A (n_3125), .B (n_4041), .C (n_3663), .Y (n_4796));
NAND4X1 g131247(.A (n_4645), .B (n_4037), .C (n_1494), .D (n_3526),.Y (n_4646));
AOI21X1 g132910(.A0 (n_4468), .A1 (n_4644), .B0 (n_4643), .Y(n_5021));
AOI21X1 g131336(.A0 (n_4117), .A1 (n_4356), .B0 (n_4525), .Y(n_5014));
OAI21X1 g131677(.A0 (n_4109), .A1 (n_1723), .B0 (n_3795), .Y(n_4780));
XOR2X1 g131365(.A (n_1804), .B (n_4070), .Y (n_4814));
INVX1 g131401(.A (n_4785), .Y (n_4642));
OAI21X1 g131413(.A0 (n_4134), .A1 (n_3943), .B0 (n_3942), .Y(n_4948));
OAI21X1 g131502(.A0 (n_4457), .A1 (n_4065), .B0 (n_4641), .Y(n_4946));
INVX1 g132180(.A (n_6378), .Y (n_6342));
OAI22X1 g131643(.A0 (n_4639), .A1 (n_4638), .B0 (n_4637), .B1(n_780), .Y (n_4640));
OAI22X1 g131652(.A0 (n_4635), .A1 (n_4634), .B0 (n_4069), .B1(n_1222), .Y (n_4636));
XOR2X1 g131661(.A (n_1226), .B (n_4342), .Y (n_4633));
INVX1 g132954(.A (n_4772), .Y (n_4735));
NOR2X1 g132703(.A (n_4632), .B (P2_reg1[12] ), .Y (n_4973));
XOR2X1 g132932(.A (n_4408), .B (n_4127), .Y (n_4631));
XOR2X1 g131866(.A (n_1847), .B (n_3989), .Y (n_4630));
INVX1 g133209(.A (n_4674), .Y (n_4629));
NAND2X1 g131925(.A (n_3673), .B (n_4152), .Y (n_4628));
NAND3X1 g132065(.A (n_4289), .B (n_2965), .C (n_4135), .Y (n_5028));
NOR3X1 g132106(.A (n_34014), .B (n_34073), .C (n_34081), .Y (n_4942));
INVX1 g132186(.A (n_34396), .Y (n_4627));
AOI21X1 g132896(.A0 (n_4259), .A1 (n_4625), .B0 (n_4624), .Y(n_4626));
NAND2X1 g132398(.A (n_4623), .B (n_4475), .Y (n_5129));
INVX1 g132468(.A (n_4520), .Y (n_4619));
INVX1 g132486(.A (n_4617), .Y (n_4618));
AOI21X1 g132499(.A0 (n_4708), .A1 (n_4430), .B0 (n_4753), .Y(n_4829));
AOI21X1 g132500(.A0 (n_4411), .A1 (n_4616), .B0 (n_4615), .Y(n_4953));
AOI21X1 g132524(.A0 (n_4433), .A1 (n_4614), .B0 (n_4589), .Y(n_5152));
OAI21X1 g132535(.A0 (n_4711), .A1 (n_4613), .B0 (n_4612), .Y(n_5464));
OAI21X1 g132542(.A0 (n_4708), .A1 (n_4398), .B0 (n_4377), .Y(n_4810));
INVX1 g132965(.A (n_6281), .Y (n_4720));
OAI21X1 g132550(.A0 (n_4611), .A1 (n_4610), .B0 (n_4609), .Y(n_5338));
NOR2X1 g132562(.A (n_3871), .B (n_4209), .Y (n_4608));
XOR2X1 g132584(.A (n_3994), .B (n_4606), .Y (n_4607));
OAI21X1 g132642(.A0 (n_4318), .A1 (n_4464), .B0 (n_4605), .Y(n_4804));
NAND2X1 g132659(.A (n_4601), .B (P3_reg1[12] ), .Y (n_5076));
NOR2X1 g132676(.A (n_4601), .B (n_13342), .Y (n_5072));
NOR2X1 g132704(.A (n_4883), .B (n_4600), .Y (n_5544));
NAND2X1 g132712(.A (n_4599), .B (P2_reg2[11] ), .Y (n_5070));
INVX1 g132718(.A (n_4929), .Y (n_4598));
NOR2X1 g132726(.A (n_4864), .B (n_4718), .Y (n_5010));
INVX1 g132732(.A (n_4800), .Y (n_4597));
INVX1 g132746(.A (n_4595), .Y (n_4596));
INVX1 g132768(.A (n_4927), .Y (n_4594));
NAND2X1 g132789(.A (n_4593), .B (n_4431), .Y (n_5107));
NAND2X1 g132801(.A (n_4592), .B (n_4424), .Y (n_5110));
NAND2X1 g132806(.A (n_4599), .B (P2_reg1[11] ), .Y (n_4972));
AND2X1 g132814(.A (n_4233), .B (n_4137), .Y (n_4591));
NOR2X1 g132817(.A (n_4535), .B (n_4590), .Y (n_4983));
NOR2X1 g132819(.A (n_4589), .B (n_4218), .Y (n_5283));
NAND2X1 g132820(.A (n_4609), .B (n_4264), .Y (n_4588));
NAND2X1 g132852(.A (n_4888), .B (n_4747), .Y (n_4586));
NOR2X1 g132853(.A (n_4718), .B (n_4589), .Y (n_4919));
INVX1 g132858(.A (n_4801), .Y (n_4585));
INVX1 g132863(.A (n_34504), .Y (n_4584));
INVX1 g132865(.A (n_4581), .Y (n_4582));
INVX1 g132876(.A (n_4579), .Y (n_4580));
AOI21X1 g132891(.A0 (n_4142), .A1 (n_4575), .B0 (n_4578), .Y(n_5096));
AOI21X1 g132899(.A0 (n_4247), .A1 (n_4577), .B0 (n_4576), .Y(n_4926));
NAND3X1 g132901(.A (n_3713), .B (n_4575), .C (n_3688), .Y (n_5098));
AOI21X1 g132908(.A0 (n_4019), .A1 (n_4574), .B0 (n_4573), .Y(n_5043));
INVX1 g133172(.A (n_4861), .Y (n_4572));
XOR2X1 g132928(.A (n_3866), .B (n_4570), .Y (n_4571));
XOR2X1 g132938(.A (n_3833), .B (n_4568), .Y (n_4569));
NOR2X1 g132414(.A (n_4478), .B (n_11141), .Y (n_4867));
NAND2X1 g133126(.A (n_35368), .B (n_4554), .Y (n_5034));
INVX1 g133154(.A (n_4565), .Y (n_4566));
INVX1 g133217(.A (n_4562), .Y (n_4563));
NAND2X1 g133192(.A (n_35368), .B (n_4561), .Y (n_5032));
INVX1 g133241(.A (n_4559), .Y (n_4560));
NAND2X1 g132843(.A (n_4379), .B (n_4556), .Y (n_4557));
NOR2X1 g132842(.A (n_4905), .B (n_4864), .Y (n_5169));
NOR2X1 g132836(.A (n_4798), .B (n_4555), .Y (n_5252));
NOR2X1 g133140(.A (n_35368), .B (n_4554), .Y (n_4884));
AOI21X1 g132892(.A0 (n_4399), .A1 (n_4552), .B0 (n_4551), .Y(n_4553));
NAND3X1 g131522(.A (n_3064), .B (n_4038), .C (n_3293), .Y (n_4550));
NAND2X1 g132825(.A (n_4211), .B (n_4713), .Y (n_4549));
INVX1 g132822(.A (n_4548), .Y (n_4728));
INVX1 g133095(.A (n_4592), .Y (n_4547));
OAI21X1 g132536(.A0 (n_4546), .A1 (n_4545), .B0 (n_4544), .Y(n_5334));
NAND2X1 g132845(.A (n_4180), .B (n_4610), .Y (n_4542));
OAI21X1 g132533(.A0 (n_4589), .A1 (n_4305), .B0 (n_4614), .Y(n_4840));
INVX1 g133101(.A (n_4593), .Y (n_4541));
NOR2X1 g132804(.A (n_4600), .B (n_4261), .Y (n_4540));
NOR2X1 g132841(.A (n_4882), .B (n_4846), .Y (n_5179));
XOR2X1 g131669(.A (n_1317), .B (n_4031), .Y (n_4538));
NOR2X1 g132833(.A (n_4252), .B (n_4675), .Y (n_4913));
NOR2X1 g132832(.A (n_4751), .B (n_4537), .Y (n_5381));
INVX1 g132794(.A (n_4536), .Y (n_4794));
NOR2X1 g132758(.A (n_4535), .B (n_4534), .Y (n_4862));
NAND4X1 g131624(.A (n_4202), .B (n_3487), .C (n_1928), .D (n_2418),.Y (n_4533));
NAND2X1 g132756(.A (n_4531), .B (n_4241), .Y (n_4532));
AOI21X1 g132508(.A0 (n_4589), .A1 (n_4423), .B0 (n_4718), .Y(n_4832));
NAND2X1 g132741(.A (n_5807), .B (n_5439), .Y (n_4530));
NOR2X1 g131309(.A (n_4499), .B (n_9670), .Y (n_5121));
NAND2X1 g132674(.A (n_4601), .B (n_13342), .Y (n_5160));
NOR2X1 g132478(.A (n_34440), .B (n_4336), .Y (n_4528));
NAND2X1 g132707(.A (n_4632), .B (P2_reg2[12] ), .Y (n_5071));
NOR2X1 g132694(.A (n_4885), .B (n_4537), .Y (n_5491));
NOR2X1 g132691(.A (n_4675), .B (n_4798), .Y (n_4872));
NOR2X1 g131397(.A (n_4525), .B (n_4306), .Y (n_4526));
NAND2X1 g132736(.A (n_4263), .B (n_4523), .Y (n_4524));
INVX1 g132669(.A (n_5073), .Y (n_4690));
OAI21X1 g132191(.A0 (n_4097), .A1 (n_2415), .B0 (n_2505), .Y(n_4656));
INVX1 g132470(.A (n_4520), .Y (n_4521));
AOI21X1 g131343(.A0 (n_4525), .A1 (n_4487), .B0 (n_4519), .Y(n_5124));
NAND2X1 g132467(.A (n_4396), .B (n_32388), .Y (n_4518));
INVX1 g132469(.A (n_4520), .Y (n_4516));
NAND2X1 g131984(.A (n_4287), .B (n_3355), .Y (n_5006));
INVX1 g132462(.A (n_4514), .Y (n_4515));
NAND2X1 g132455(.A (n_4155), .B (n_4511), .Y (n_4512));
XOR2X1 g131874(.A (n_1994), .B (n_4108), .Y (n_4817));
INVX1 g132460(.A (n_4508), .Y (n_4509));
NAND2X1 g131964(.A (n_6017), .B (n_5940), .Y (n_5650));
INVX1 g133016(.A (n_4507), .Y (n_4825));
AOI21X1 g131619(.A0 (n_3986), .A1 (n_4504), .B0 (n_4110), .Y(n_4505));
XOR2X1 g131865(.A (n_1533), .B (n_3996), .Y (n_4503));
INVX1 g132441(.A (n_33242), .Y (n_4502));
OAI21X1 g131384(.A0 (n_4050), .A1 (n_2397), .B0 (n_4293), .Y(n_4847));
NAND2X1 g132702(.A (n_4632), .B (P2_reg1[12] ), .Y (n_4971));
NAND2X1 g131293(.A (n_4499), .B (n_9670), .Y (n_5016));
NOR2X1 g132661(.A (n_4601), .B (P3_reg1[12] ), .Y (n_5075));
INVX1 g131751(.A (n_5120), .Y (n_4498));
NOR2X1 g132826(.A (n_4599), .B (P2_reg1[11] ), .Y (n_4961));
INVX1 g133200(.A (n_4496), .Y (n_4497));
AOI21X1 g132897(.A0 (n_4324), .A1 (n_4495), .B0 (n_4494), .Y(n_4845));
AOI21X1 g132903(.A0 (n_4257), .A1 (n_4414), .B0 (n_4493), .Y(n_4826));
INVX1 g131426(.A (n_4491), .Y (n_4783));
NOR2X1 g132687(.A (n_4599), .B (P2_reg2[11] ), .Y (n_4959));
NAND2X1 g132341(.A (n_4192), .B (n_609), .Y (n_35117));
NAND2X1 g131727(.A (n_4488), .B (n_4487), .Y (n_5013));
XOR2X1 g131882(.A (n_1802), .B (n_4061), .Y (n_4486));
INVX1 g132662(.A (n_4787), .Y (n_4481));
NAND2X1 g132731(.A (n_3845), .B (n_4213), .Y (n_5221));
NAND2X1 g133227(.A (n_4670), .B (n_4460), .Y (n_5100));
INVX1 g132224(.A (n_5234), .Y (n_5925));
NAND2X1 g132766(.A (n_3845), .B (n_4215), .Y (n_5155));
NAND2X1 g132389(.A (n_4592), .B (n_4915), .Y (n_5237));
NOR2X1 g132365(.A (n_4478), .B (n_4477), .Y (n_4791));
INVX1 g133150(.A (n_4895), .Y (n_4476));
NAND2X1 g131744(.A (n_4694), .B (n_4488), .Y (n_5123));
NAND2X1 g132337(.A (n_4623), .B (P2_reg1[17] ), .Y (n_5085));
NAND2X1 g132381(.A (n_4593), .B (n_4921), .Y (n_5277));
NOR2X1 g132279(.A (n_4623), .B (n_4475), .Y (n_4933));
NAND2X1 g132233(.A (n_4288), .B (n_4474), .Y (n_4934));
OAI21X1 g132202(.A0 (n_4473), .A1 (n_2497), .B0 (n_4472), .Y(n_4965));
INVX1 g132195(.A (n_6180), .Y (n_4471));
NAND3X1 g132888(.A (n_3678), .B (n_4082), .C (n_3745), .Y (n_4657));
NOR2X1 g132248(.A (n_4623), .B (P2_reg1[17] ), .Y (n_4860));
INVX1 g133448(.A (n_4601), .Y (n_10656));
NAND2X1 g132025(.A (n_4353), .B (n_3815), .Y (n_4470));
NOR2X1 g132007(.A (n_4519), .B (n_4114), .Y (n_4469));
AOI21X1 g133299(.A0 (n_6044), .A1 (n_4465), .B0 (n_4468), .Y(n_4893));
NAND3X1 g133284(.A (n_3627), .B (n_4400), .C (n_3822), .Y (n_4925));
OR2X1 g132850(.A (n_34503), .B (n_3545), .Y (n_4467));
OR2X1 g131701(.A (n_3738), .B (n_4042), .Y (n_4466));
AND2X1 g133242(.A (n_4465), .B (n_4644), .Y (n_4559));
OAI21X1 g132637(.A0 (n_3861), .A1 (n_4401), .B0 (n_4363), .Y(n_5137));
NOR2X1 g133221(.A (n_4319), .B (n_4464), .Y (n_4805));
INVX1 g131765(.A (n_5182), .Y (n_4463));
INVX1 g133128(.A (n_4752), .Y (n_4462));
NAND2X1 g133210(.A (n_4461), .B (n_4237), .Y (n_4674));
AOI21X1 g132916(.A0 (n_4304), .A1 (n_4460), .B0 (n_4459), .Y(n_4899));
NAND3X1 g131642(.A (n_3969), .B (n_3847), .C (n_4457), .Y (n_4868));
NOR2X1 g131714(.A (n_4637), .B (n_2173), .Y (n_4456));
NOR2X1 g131736(.A (n_4136), .B (n_3507), .Y (n_4851));
XOR2X1 g131847(.A (n_1900), .B (n_3864), .Y (n_4668));
XOR2X1 g131859(.A (n_1418), .B (n_3890), .Y (n_4665));
XOR2X1 g131863(.A (n_1287), .B (n_3974), .Y (n_4455));
XOR2X1 g131864(.A (n_1930), .B (n_3950), .Y (n_4454));
XOR2X1 g131880(.A (n_1951), .B (n_3903), .Y (n_4453));
INVX1 g131955(.A (n_4694), .Y (n_4452));
NOR2X1 g131990(.A (n_4335), .B (n_3577), .Y (n_4451));
INVX1 g131993(.A (n_4488), .Y (n_4450));
AOI21X1 g132080(.A0 (n_3940), .A1 (n_2851), .B0 (n_3949), .Y(n_4449));
NAND2X1 g133236(.A (n_4625), .B (n_4260), .Y (n_4448));
XOR2X1 g132167(.A (n_1558), .B (n_3888), .Y (n_4447));
XOR2X1 g132170(.A (n_1403), .B (n_4286), .Y (n_4446));
NOR2X1 g133193(.A (n_4010), .B (n_4445), .Y (n_5185));
NOR2X1 g132226(.A (n_4311), .B (P3_reg1[17] ), .Y (n_5234));
XOR2X1 g131846(.A (n_1185), .B (n_3952), .Y (n_4444));
AND2X1 g132361(.A (n_6125), .B (n_5940), .Y (n_6394));
INVX1 g132075(.A (n_4294), .Y (n_4443));
INVX1 g132512(.A (n_4441), .Y (n_4442));
NAND2X1 g133223(.A (n_4616), .B (n_4412), .Y (n_4954));
NOR2X1 g132614(.A (n_4130), .B (n_1633), .Y (n_4439));
NOR2X1 g132866(.A (n_4232), .B (n_35251), .Y (n_4581));
OAI21X1 g132625(.A0 (n_4300), .A1 (n_4195), .B0 (n_4437), .Y(n_4770));
OAI21X1 g132640(.A0 (n_3923), .A1 (n_4240), .B0 (n_4421), .Y(n_5232));
INVX1 g133591(.A (n_4714), .Y (n_4436));
INVX1 g132656(.A (n_4774), .Y (n_4602));
NOR2X1 g132685(.A (n_4632), .B (P2_reg2[12] ), .Y (n_4987));
NOR2X1 g133585(.A (n_4433), .B (n_4022), .Y (n_5295));
NAND2X1 g132719(.A (n_4432), .B (n_4160), .Y (n_4929));
NAND2X1 g132723(.A (n_4431), .B (n_4430), .Y (n_5046));
NOR2X1 g132737(.A (n_4433), .B (n_4589), .Y (n_4835));
NAND2X1 g132749(.A (n_5624), .B (n_5228), .Y (n_4429));
NAND2X1 g132759(.A (n_4544), .B (n_4094), .Y (n_4428));
AND2X1 g132762(.A (n_5861), .B (n_4426), .Y (n_35872));
NAND2X1 g132318(.A (n_3992), .B (n_4112), .Y (n_4425));
NAND2X1 g132795(.A (n_4305), .B (n_4614), .Y (n_4536));
NAND2X1 g132838(.A (n_4424), .B (n_4423), .Y (n_5052));
OR2X1 g132854(.A (n_4421), .B (n_4420), .Y (n_4422));
INVX1 g132861(.A (n_4418), .Y (n_4419));
INVX1 g132314(.A (n_4416), .Y (n_4417));
NAND2X1 g132877(.A (n_4345), .B (n_32435), .Y (n_4579));
NAND2X1 g132881(.A (n_3775), .B (n_33046), .Y (n_4415));
NAND2X1 g132859(.A (n_4432), .B (P2_reg1[13] ), .Y (n_4801));
NAND3X1 g132905(.A (n_3747), .B (n_4414), .C (n_3797), .Y (n_4828));
NAND2X1 g132857(.A (n_8105), .B (n_10223), .Y (n_4767));
NOR2X1 g133173(.A (n_4010), .B (P1_reg1[12] ), .Y (n_4861));
AOI21X1 g132917(.A0 (n_3920), .A1 (n_4412), .B0 (n_4411), .Y(n_4900));
XOR2X1 g132935(.A (n_4409), .B (n_4408), .Y (n_4410));
INVX1 g132982(.A (n_34078), .Y (n_4911));
INVX1 g133011(.A (n_34485), .Y (n_6324));
INVX1 g133098(.A (n_4430), .Y (n_4405));
INVX1 g133104(.A (n_4377), .Y (n_4404));
NOR2X1 g133142(.A (n_4402), .B (n_4401), .Y (n_4403));
NAND2X1 g133231(.A (n_4700), .B (n_4414), .Y (n_5094));
AOI21X1 g133280(.A0 (n_4081), .A1 (n_4400), .B0 (n_4399), .Y(n_4924));
OAI21X1 g133321(.A0 (n_4075), .A1 (n_4267), .B0 (n_4398), .Y(n_4669));
INVX1 g132966(.A (n_4396), .Y (n_6281));
INVX1 g133460(.A (n_4599), .Y (n_4395));
INVX1 g133588(.A (n_4883), .Y (n_4394));
NAND2X1 g133151(.A (n_4461), .B (n_4344), .Y (n_4895));
AND2X1 g133201(.A (n_4255), .B (n_4650), .Y (n_4496));
INVX1 g133147(.A (n_4612), .Y (n_4392));
INVX1 g133653(.A (n_5101), .Y (n_4391));
AND2X1 g132285(.A (n_6079), .B (n_5951), .Y (n_6454));
INVX1 g133465(.A (n_4632), .Y (n_4389));
NAND2X1 g132823(.A (n_4398), .B (n_4377), .Y (n_4548));
INVX1 g132815(.A (n_5157), .Y (n_4388));
INVX1 g133115(.A (n_4423), .Y (n_4386));
INVX1 g133455(.A (n_4385), .Y (n_4731));
INVX1 g133238(.A (n_4754), .Y (n_4384));
NOR2X1 g132813(.A (n_4611), .B (n_4555), .Y (n_5275));
NOR2X1 g132846(.A (n_4753), .B (n_4708), .Y (n_4808));
INVX1 g133214(.A (n_4379), .Y (n_4380));
NOR2X1 g132828(.A (n_4727), .B (n_4378), .Y (n_5404));
NAND2X1 g132785(.A (n_4377), .B (n_4430), .Y (n_4806));
INVX1 g132782(.A (n_4375), .Y (n_4376));
NAND2X1 g132777(.A (n_4096), .B (n_4545), .Y (n_4373));
NOR2X1 g132784(.A (n_4711), .B (n_4600), .Y (n_5376));
NAND2X1 g132249(.A (n_4032), .B (n_4371), .Y (n_4372));
NOR2X1 g132770(.A (n_6988), .B (n_4367), .Y (n_4928));
NOR2X1 g132611(.A (n_3573), .B (n_349), .Y (n_4368));
NAND2X1 g132752(.A (n_4614), .B (n_4423), .Y (n_4821));
NAND2X1 g132769(.A (n_6988), .B (n_4367), .Y (n_4927));
OR2X1 g132750(.A (n_4363), .B (n_4402), .Y (n_4364));
CLKBUFX1 g132955(.A (n_4511), .Y (n_4772));
INVX1 g132724(.A (n_4361), .Y (n_4362));
NOR2X1 g131806(.A (n_4052), .B (n_4125), .Y (n_4360));
NAND2X1 g133237(.A (n_4552), .B (n_4400), .Y (n_4359));
CLKBUFX1 g132976(.A (n_33485), .Y (n_4764));
NAND2X1 g131427(.A (n_4487), .B (n_4356), .Y (n_4491));
NOR2X1 g132748(.A (n_4846), .B (n_4753), .Y (n_5022));
NOR2X1 g132744(.A (n_4432), .B (P2_reg1[13] ), .Y (n_4912));
NAND2X1 g132747(.A (n_8105), .B (n_4277), .Y (n_4595));
NOR2X1 g132483(.A (n_4354), .B (n_32639), .Y (n_4355));
NAND2X1 g132733(.A (n_6988), .B (n_9586), .Y (n_4800));
NAND2X1 g132182(.A (n_2920), .B (n_4085), .Y (n_6378));
NAND2X1 g132196(.A (n_2322), .B (n_4002), .Y (n_6180));
NOR2X1 g131986(.A (n_2641), .B (n_4353), .Y (n_4777));
NAND2X1 g132471(.A (n_4351), .B (n_3776), .Y (n_4520));
INVX1 g132649(.A (n_4350), .Y (n_4975));
NOR2X1 g132459(.A (n_4328), .B (n_4219), .Y (n_4349));
NOR2X1 g132461(.A (n_32639), .B (n_4256), .Y (n_4508));
NOR2X1 g132720(.A (n_6988), .B (n_9586), .Y (n_4909));
AND2X1 g133218(.A (n_4347), .B (n_4726), .Y (n_4562));
NAND2X1 g132867(.A (n_3851), .B (n_4345), .Y (n_4346));
NOR2X1 g133204(.A (n_4461), .B (n_4344), .Y (n_4870));
NOR2X1 g131681(.A (n_4342), .B (n_4341), .Y (n_4343));
NAND2X1 g133526(.A (n_4139), .B (n_4398), .Y (n_5399));
INVX1 g133024(.A (n_4623), .Y (n_4340));
NAND2X1 g133048(.A (n_35335), .B (n_35336), .Y (n_4653));
INVX1 g133224(.A (n_4751), .Y (n_4339));
NOR2X1 g132670(.A (n_32442), .B (P3_reg2[13] ), .Y (n_5073));
NAND2X1 g131762(.A (n_4313), .B (n_9653), .Y (n_4978));
NAND2X1 g131402(.A (n_4118), .B (n_4356), .Y (n_4785));
INVX1 g133004(.A (n_6208), .Y (n_6204));
INVX1 g133017(.A (n_4336), .Y (n_4507));
NAND3X1 g131953(.A (n_4335), .B (n_4334), .C (n_2207), .Y (n_4852));
NAND2X1 g132465(.A (n_32394), .B (n_4266), .Y (n_32023));
NAND2X1 g132463(.A (n_4194), .B (n_4067), .Y (n_4514));
NOR2X1 g132487(.A (n_3881), .B (n_35195), .Y (n_4617));
INVX1 g132622(.A (n_4325), .Y (n_4326));
AOI21X1 g133314(.A0 (n_5624), .A1 (n_4095), .B0 (n_4324), .Y(n_5002));
NOR2X1 g131754(.A (n_4322), .B (n_4321), .Y (n_4323));
INVX1 g133428(.A (n_4320), .Y (n_4701));
OAI21X1 g133080(.A0 (n_5825), .A1 (n_4319), .B0 (n_4318), .Y(n_4890));
AND2X1 g133155(.A (n_4020), .B (n_4574), .Y (n_4565));
XOR2X1 g131858(.A (n_1912), .B (n_3980), .Y (n_4677));
INVX2 g133167(.A (n_4315), .Y (n_6375));
NOR2X1 g131752(.A (n_4313), .B (n_9653), .Y (n_5120));
NAND2X1 g132238(.A (n_4311), .B (P3_reg1[17] ), .Y (n_5946));
NAND2X1 g133162(.A (n_4756), .B (n_4575), .Y (n_4985));
XOR2X1 g131868(.A (n_1592), .B (n_3908), .Y (n_4310));
XOR2X1 g133397(.A (n_5972), .B (n_3689), .Y (n_4308));
AND2X1 g131973(.A (n_4307), .B (n_3968), .Y (n_4947));
NOR2X1 g131959(.A (n_4201), .B (addr_492), .Y (n_4684));
CLKBUFX1 g133025(.A (n_34232), .Y (n_4623));
OAI21X1 g133313(.A0 (n_4145), .A1 (n_4080), .B0 (n_4244), .Y(n_4649));
OAI21X1 g133312(.A0 (n_4225), .A1 (n_4162), .B0 (n_4253), .Y(n_4643));
INVX1 g131565(.A (n_4356), .Y (n_4306));
AOI21X1 g133282(.A0 (n_4278), .A1 (n_4305), .B0 (n_4433), .Y(n_4833));
AOI21X1 g133655(.A0 (n_3990), .A1 (n_4523), .B0 (n_4304), .Y(n_5101));
OAI21X1 g132943(.A0 (n_3695), .A1 (n_33579), .B0 (n_1473), .Y(n_4365));
NAND2X1 g133103(.A (n_4217), .B (n_13721), .Y (n_4593));
XOR2X1 g131852(.A (n_1772), .B (n_3741), .Y (n_4303));
XOR2X1 g133382(.A (n_3824), .B (n_5956), .Y (n_4302));
NAND2X1 g133129(.A (n_4301), .B (P2_reg2[8] ), .Y (n_4752));
OAI21X1 g133065(.A0 (n_3393), .A1 (n_4196), .B0 (n_4300), .Y(n_4746));
OAI21X1 g133324(.A0 (n_4250), .A1 (n_4299), .B0 (n_4298), .Y(n_4624));
NAND4X1 g131773(.A (n_3896), .B (n_3746), .C (n_2054), .D (n_2344),.Y (n_4297));
XOR2X1 g131855(.A (n_1120), .B (n_3727), .Y (n_4296));
OR2X1 g131902(.A (n_3895), .B (n_3945), .Y (n_4295));
NAND2X1 g133592(.A (n_8115), .B (n_4230), .Y (n_4714));
AOI21X1 g132076(.A0 (n_3789), .A1 (n_4293), .B0 (n_1902), .Y(n_4294));
XOR2X1 g132173(.A (n_1784), .B (n_3891), .Y (n_4291));
XOR2X1 g132174(.A (n_2287), .B (n_3767), .Y (n_4290));
NAND3X1 g132213(.A (n_3892), .B (n_2207), .C (n_2363), .Y (n_4289));
OR2X1 g132222(.A (n_4288), .B (n_4474), .Y (n_6017));
NAND3X1 g132277(.A (n_4286), .B (n_3353), .C (n_4014), .Y (n_4287));
INVX1 g132998(.A (n_4285), .Y (n_6313));
NAND2X1 g132477(.A (n_6467), .B (n_4003), .Y (n_4284));
OAI21X1 g132498(.A0 (n_3816), .A1 (n_3352), .B0 (n_4282), .Y(n_4283));
NAND2X1 g132523(.A (n_3944), .B (n_4280), .Y (n_4281));
MX2X1 g132603(.A (n_593), .B (P3_IR[27] ), .S0 (n_3777), .Y(n_4279));
OAI21X1 g133315(.A0 (n_4278), .A1 (n_3982), .B0 (n_4246), .Y(n_4576));
NOR2X1 g132722(.A (n_8105), .B (n_4277), .Y (n_4902));
NOR2X1 g132862(.A (n_4092), .B (n_4056), .Y (n_4418));
NAND2X1 g132875(.A (n_3599), .B (n_4068), .Y (n_4274));
NOR2X1 g132878(.A (n_33573), .B (n_4271), .Y (n_35254));
OR2X1 g132316(.A (n_3936), .B (n_3373), .Y (n_4416));
NAND2X1 g132555(.A (n_3946), .B (n_2900), .Y (n_4270));
OAI21X1 g133319(.A0 (n_4229), .A1 (n_4023), .B0 (n_4267), .Y(n_4494));
INVX2 g133168(.A (n_4043), .Y (n_4315));
CLKBUFX3 g132956(.A (n_4266), .Y (n_4511));
AND2X1 g133089(.A (n_4133), .B (n_4265), .Y (n_4718));
INVX1 g133131(.A (n_4611), .Y (n_4264));
AND2X1 g133146(.A (n_4248), .B (n_4577), .Y (n_5439));
INVX1 g133170(.A (n_4262), .Y (n_4263));
INVX1 g133181(.A (n_4613), .Y (n_4261));
NAND2X1 g133239(.A (n_4301), .B (P2_reg1[8] ), .Y (n_4754));
AOI21X1 g133274(.A0 (n_4059), .A1 (n_4260), .B0 (n_4259), .Y(n_4472));
AOI21X1 g133276(.A0 (n_3748), .A1 (n_4258), .B0 (n_4257), .Y(n_5095));
INVX1 g132967(.A (n_4256), .Y (n_4396));
AOI21X1 g133292(.A0 (n_5956), .A1 (n_4255), .B0 (n_4254), .Y(n_4744));
OAI21X1 g133311(.A0 (n_4253), .A1 (n_4252), .B0 (n_4251), .Y(n_4699));
OAI21X1 g133316(.A0 (n_4234), .A1 (n_4249), .B0 (n_4149), .Y(n_4725));
OAI21X1 g133317(.A0 (n_4119), .A1 (n_3832), .B0 (n_4250), .Y(n_4573));
OAI21X1 g133322(.A0 (n_4224), .A1 (n_4034), .B0 (n_4249), .Y(n_4578));
AOI21X1 g133326(.A0 (n_5807), .A1 (n_4248), .B0 (n_4247), .Y(n_4888));
OAI21X1 g133327(.A0 (n_4433), .A1 (n_4246), .B0 (n_4305), .Y(n_4615));
OAI21X1 g133328(.A0 (n_4244), .A1 (n_4243), .B0 (n_4242), .Y(n_4551));
NOR2X1 g133158(.A (n_4420), .B (n_4240), .Y (n_4241));
CLKBUFX1 g133449(.A (n_4345), .Y (n_4601));
NOR2X1 g133149(.A (n_4461), .B (n_4237), .Y (n_4675));
INVX1 g133519(.A (n_4464), .Y (n_4236));
NOR2X1 g133552(.A (n_4129), .B (n_3915), .Y (n_4747));
NAND2X1 g133555(.A (n_8115), .B (n_4231), .Y (n_4789));
NOR2X1 g133568(.A (n_3913), .B (n_4234), .Y (n_4235));
INVX1 g133251(.A (n_4232), .Y (n_4233));
NOR2X1 g133589(.A (n_8115), .B (n_4231), .Y (n_4883));
NOR2X1 g133600(.A (n_8115), .B (n_4230), .Y (n_4885));
NAND2X1 g132623(.A (n_3687), .B (n_6303), .Y (n_4325));
NOR2X1 g133607(.A (n_4229), .B (n_3953), .Y (n_5329));
NOR2X1 g133613(.A (n_4075), .B (n_4229), .Y (n_4670));
NOR2X1 g133621(.A (n_3922), .B (n_4225), .Y (n_4226));
NAND2X1 g133148(.A (n_3959), .B (n_3958), .Y (n_4612));
OAI21X1 g133661(.A0 (n_4072), .A1 (n_3701), .B0 (n_4224), .Y(n_4651));
AOI21X1 g133293(.A0 (n_4267), .A1 (n_4156), .B0 (n_4229), .Y(n_4605));
NOR2X1 g132831(.A (n_4075), .B (n_4708), .Y (n_4703));
NAND2X1 g133866(.A (n_4224), .B (n_3859), .Y (n_4223));
INVX1 g132987(.A (n_4351), .Y (n_4478));
NOR2X1 g133551(.A (n_3877), .B (n_4252), .Y (n_4220));
INVX1 g133456(.A (n_4219), .Y (n_4385));
INVX1 g133118(.A (n_4614), .Y (n_4218));
NOR2X1 g133120(.A (n_4217), .B (P3_reg2[10] ), .Y (n_4905));
AND2X1 g133215(.A (n_3921), .B (n_4412), .Y (n_4379));
NOR2X1 g132816(.A (n_3845), .B (n_4215), .Y (n_5157));
NOR2X1 g132818(.A (n_4546), .B (n_4378), .Y (n_5231));
NOR2X1 g132792(.A (n_3845), .B (n_4213), .Y (n_5216));
INVX1 g133111(.A (n_4424), .Y (n_4382));
NAND2X1 g133097(.A (n_4217), .B (P3_reg2[10] ), .Y (n_4592));
NOR2X1 g132563(.A (n_3856), .B (n_3853), .Y (n_4212));
INVX1 g133229(.A (n_4537), .Y (n_4211));
INVX1 g133470(.A (n_4432), .Y (n_4210));
NAND2X1 g132874(.A (n_3621), .B (n_4157), .Y (n_4209));
NAND2X1 g132652(.A (n_4200), .B (P3_reg1[11] ), .Y (n_4921));
OR2X1 g132035(.A (n_3737), .B (n_3926), .Y (n_4206));
NAND2X1 g132783(.A (n_4205), .B (P2_reg1[18] ), .Y (n_4375));
NOR2X1 g132767(.A (n_4205), .B (P2_reg1[18] ), .Y (n_4859));
NOR2X1 g133122(.A (n_4217), .B (n_13721), .Y (n_4882));
OR2X1 g131991(.A (n_3979), .B (n_3485), .Y (n_4202));
NAND2X1 g131994(.A (n_4201), .B (addr_492), .Y (n_4488));
NAND2X1 g132725(.A (n_4205), .B (P2_reg2[18] ), .Y (n_4361));
NOR2X1 g132657(.A (n_4200), .B (n_13366), .Y (n_4774));
OAI21X1 g131385(.A0 (n_3731), .A1 (n_2384), .B0 (n_3697), .Y(n_4645));
INVX1 g132475(.A (n_4749), .Y (n_32241));
NOR2X1 g132457(.A (n_6810), .B (n_6348), .Y (n_4198));
NOR2X1 g131967(.A (n_4164), .B (n_9655), .Y (n_4792));
XOR2X1 g132168(.A (n_1298), .B (n_4116), .Y (n_4197));
NOR2X1 g133211(.A (n_4196), .B (n_4195), .Y (n_4771));
INVX1 g133018(.A (n_4194), .Y (n_4336));
INVX1 g132697(.A (n_4766), .Y (n_4193));
OAI22X1 g133049(.A0 (n_3829), .A1 (n_241), .B0 (n_3830), .B1(P1_IR[30] ), .Y (n_4192));
XOR2X1 g131867(.A (n_1535), .B (n_3805), .Y (n_4191));
XOR2X1 g133393(.A (n_4166), .B (n_3467), .Y (n_4190));
MX2X1 g132602(.A (n_600), .B (P2_IR[27] ), .S0 (n_3828), .Y(n_4189));
NOR2X1 g131766(.A (n_3878), .B (n_2845), .Y (n_5182));
XOR2X1 g131490(.A (n_1873), .B (n_3708), .Y (n_4499));
INVX1 g133031(.A (n_4188), .Y (n_6527));
NOR2X1 g133225(.A (n_3959), .B (n_4151), .Y (n_4751));
XOR2X1 g132169(.A (n_1528), .B (n_4015), .Y (n_4187));
NOR2X1 g133548(.A (n_3886), .B (n_4185), .Y (n_4186));
XOR2X1 g133380(.A (n_4175), .B (n_5624), .Y (n_4184));
XOR2X1 g133388(.A (n_6044), .B (n_3799), .Y (n_4183));
XOR2X1 g133384(.A (n_3772), .B (n_5914), .Y (n_4182));
XOR2X1 g131860(.A (n_1193), .B (n_3813), .Y (n_4181));
INVX1 g133243(.A (n_4555), .Y (n_4180));
NAND3X1 g132331(.A (n_3842), .B (n_4179), .C (n_2792), .Y (n_5189));
INVX1 g133093(.A (n_4431), .Y (n_4381));
XOR2X1 g133386(.A (n_4175), .B (n_3463), .Y (n_4176));
INVX1 g132868(.A (n_34439), .Y (n_4174));
XOR2X1 g131854(.A (n_3669), .B (n_3985), .Y (so[4]));
INVX1 g133376(.A (n_4170), .Y (n_6291));
INVX1 g133013(.A (n_34482), .Y (n_4169));
XOR2X1 g133379(.A (n_5807), .B (n_4166), .Y (n_4167));
OR2X1 g132516(.A (n_3885), .B (n_3090), .Y (n_4165));
NAND2X1 g131956(.A (n_4164), .B (n_9655), .Y (n_4694));
NOR2X1 g133232(.A (n_4301), .B (P2_reg1[8] ), .Y (n_4798));
OAI21X1 g133325(.A0 (n_4053), .A1 (n_4005), .B0 (n_4162), .Y(n_4493));
OR2X1 g132514(.A (n_3910), .B (n_2891), .Y (n_4441));
NOR2X1 g132715(.A (n_4432), .B (n_4160), .Y (n_4907));
INVX1 g133005(.A (n_4328), .Y (n_6208));
MX2X1 g132579(.A (n_1890), .B (P1_IR[27] ), .S0 (n_33681), .Y(n_4159));
NOR2X1 g132664(.A (n_4200), .B (P3_reg1[11] ), .Y (n_4787));
AND2X1 g132870(.A (n_4157), .B (n_3957), .Y (n_4158));
NOR2X1 g133617(.A (n_4156), .B (n_3916), .Y (n_4891));
INVX1 g133429(.A (n_4155), .Y (n_4320));
NAND2X1 g132651(.A (n_32445), .B (n_3848), .Y (n_4350));
NAND3X1 g132338(.A (n_3897), .B (n_3951), .C (n_2188), .Y (n_4152));
NAND2X1 g133164(.A (n_3959), .B (n_4151), .Y (n_4750));
NAND2X1 g133612(.A (n_4250), .B (n_3873), .Y (n_4150));
OAI21X1 g133318(.A0 (n_4149), .A1 (n_4185), .B0 (n_4148), .Y(n_4755));
NOR2X1 g132199(.A (n_10110), .B (n_3964), .Y (n_4147));
NOR2X1 g133525(.A (n_3909), .B (n_4145), .Y (n_4146));
INVX1 g132946(.A (n_34119), .Y (n_6188));
AOI21X1 g133289(.A0 (n_3714), .A1 (n_4143), .B0 (n_4142), .Y(n_4986));
CLKBUFX1 g133467(.A (n_4141), .Y (n_4632));
OR2X1 g133117(.A (n_4133), .B (n_4265), .Y (n_4423));
NAND2X1 g132671(.A (n_32442), .B (P3_reg2[13] ), .Y (n_5215));
INVX1 g133934(.A (n_4075), .Y (n_4139));
AND2X1 g133161(.A (n_3863), .B (n_4137), .Y (n_4138));
NAND2X1 g133252(.A (n_3593), .B (n_3863), .Y (n_4232));
AOI21X1 g132097(.A0 (n_3578), .A1 (n_4135), .B0 (n_1917), .Y(n_4136));
AOI21X1 g131808(.A0 (n_4120), .A1 (n_3538), .B0 (n_3537), .Y(n_4134));
AND2X1 g133121(.A (n_4133), .B (n_4132), .Y (n_4753));
NOR2X1 g133244(.A (n_4131), .B (P2_reg1[9] ), .Y (n_4555));
INVX1 g133344(.A (n_8447), .Y (n_4130));
OAI21X1 g133323(.A0 (n_4129), .A1 (n_3983), .B0 (n_3982), .Y(n_4411));
NAND2X1 g133144(.A (n_4131), .B (P2_reg1[9] ), .Y (n_4610));
NAND2X1 g133544(.A (n_4246), .B (n_4305), .Y (n_4402));
INVX1 g133656(.A (n_4955), .Y (n_4127));
NOR2X1 g132325(.A (n_3794), .B (n_2535), .Y (n_4125));
NAND2X1 g133006(.A (n_1575), .B (n_3781), .Y (n_4328));
NOR2X1 g131673(.A (n_3453), .B (P1_n_449), .Y (n_4124));
XOR2X1 g131853(.A (n_1379), .B (n_4049), .Y (n_4122));
XOR2X1 g131862(.A (n_1568), .B (n_4120), .Y (n_4121));
NOR2X1 g133528(.A (n_4119), .B (n_4299), .Y (n_4625));
AOI21X1 g131961(.A0 (n_3675), .A1 (n_3894), .B0 (n_3893), .Y(n_4637));
AOI21X1 g132064(.A0 (n_4035), .A1 (n_2482), .B0 (n_3183), .Y(n_4342));
AOI21X1 g132079(.A0 (n_4012), .A1 (n_4118), .B0 (n_4117), .Y(n_4681));
NOR2X1 g132210(.A (n_4116), .B (n_2435), .Y (n_4335));
NAND2X1 g132260(.A (n_3750), .B (n_4118), .Y (n_4115));
INVX1 g132300(.A (n_4487), .Y (n_4114));
NAND2X1 g132302(.A (n_3817), .B (n_4112), .Y (n_4113));
INVX1 g132309(.A (n_4110), .Y (n_4111));
NOR2X1 g132456(.A (n_3876), .B (n_34092), .Y (n_4940));
NAND2X1 g132476(.A (n_3941), .B (n_33899), .Y (n_4749));
AOI21X1 g132526(.A0 (n_3902), .A1 (n_2642), .B0 (n_2880), .Y(n_4109));
NAND2X2 g132969(.A (n_35283), .B (n_35284), .Y (n_4256));
NAND4X1 g132565(.A (n_3753), .B (n_2148), .C (n_2580), .D (n_2728),.Y (n_4108));
NAND2X1 g133182(.A (n_3870), .B (n_4011), .Y (n_4613));
OR2X1 g132677(.A (n_3999), .B (P3_reg2[18] ), .Y (n_6125));
NOR2X1 g132721(.A (n_3564), .B (n_34178), .Y (n_4357));
NAND2X1 g132895(.A (n_3690), .B (n_4100), .Y (n_4101));
NOR2X1 g133132(.A (n_4099), .B (P2_reg1[10] ), .Y (n_4611));
AND2X1 g132979(.A (n_3783), .B (n_3634), .Y (n_4097));
INVX1 g133019(.A (n_3962), .Y (n_4194));
AOI21X1 g133646(.A0 (n_4091), .A1 (n_3899), .B0 (n_4079), .Y(n_4318));
NAND2X1 g133145(.A (n_4099), .B (P2_reg2[10] ), .Y (n_4544));
NOR2X1 g131584(.A (n_4017), .B (addr_490), .Y (n_4525));
INVX1 g133194(.A (n_4378), .Y (n_4096));
AND2X1 g133196(.A (n_4095), .B (n_4495), .Y (n_5228));
INVX1 g133247(.A (n_4546), .Y (n_4094));
INVX1 g133256(.A (n_4092), .Y (n_32021));
OAI21X1 g133320(.A0 (n_4156), .A1 (n_4091), .B0 (n_4023), .Y(n_4459));
INVX1 g133364(.A (n_3887), .Y (n_4154));
OAI21X1 g132844(.A0 (n_3614), .A1 (n_2627), .B0 (n_4371), .Y(n_4087));
INVX1 g133439(.A (n_4205), .Y (n_4086));
NAND2X1 g132299(.A (n_3784), .B (n_34946), .Y (n_4085));
NOR2X1 g133558(.A (n_4433), .B (n_4278), .Y (n_4616));
INVX1 g133609(.A (n_4195), .Y (n_4083));
NOR2X1 g133616(.A (n_4225), .B (n_4252), .Y (n_4700));
INVX1 g133625(.A (n_4401), .Y (n_4082));
INVX1 g133478(.A (n_4157), .Y (n_4535));
AOI21X1 g133644(.A0 (n_3639), .A1 (n_2674), .B0 (n_4081), .Y(n_4570));
OAI21X1 g133663(.A0 (n_3865), .A1 (n_4004), .B0 (n_4080), .Y(n_4399));
OAI21X1 g133667(.A0 (n_4079), .A1 (n_3663), .B0 (n_4091), .Y(n_4324));
OAI21X1 g133711(.A0 (n_3849), .A1 (n_4556), .B0 (n_3820), .Y(n_4078));
XOR2X1 g133712(.A (n_2313), .B (n_3562), .Y (n_4077));
NAND2X1 g133143(.A (n_3870), .B (P1_reg2[9] ), .Y (n_4713));
AOI21X1 g133277(.A0 (n_4229), .A1 (n_4398), .B0 (n_4075), .Y(n_4830));
AOI21X1 g133267(.A0 (n_3978), .A1 (n_3982), .B0 (n_4129), .Y(n_4363));
INVX1 g132988(.A (n_3930), .Y (n_4351));
NOR2X1 g133852(.A (n_4072), .B (n_3702), .Y (n_4347));
NOR2X1 g133137(.A (n_4301), .B (P2_reg2[8] ), .Y (n_4727));
NAND2X1 g133520(.A (n_4267), .B (n_4023), .Y (n_4464));
NAND3X1 g131523(.A (n_2904), .B (n_3676), .C (n_2112), .Y (n_4070));
NAND2X1 g133125(.A (n_4131), .B (P2_reg2[9] ), .Y (n_4545));
INVX1 g132061(.A (n_4073), .Y (n_4069));
INVX1 g133462(.A (n_4068), .Y (n_4599));
NAND2X1 g133119(.A (n_3911), .B (n_13361), .Y (n_4614));
INVX1 g133457(.A (n_4067), .Y (n_4219));
NOR2X1 g133604(.A (n_4145), .B (n_4243), .Y (n_4552));
NOR2X1 g133230(.A (n_3870), .B (P1_reg2[9] ), .Y (n_4537));
INVX2 g133450(.A (n_3987), .Y (n_4345));
NOR2X1 g133113(.A (n_4066), .B (P3_reg1[9] ), .Y (n_4846));
NOR2X1 g133107(.A (n_4066), .B (P3_reg2[9] ), .Y (n_4864));
NAND2X1 g133112(.A (n_4066), .B (P3_reg2[9] ), .Y (n_4424));
INVX1 g132271(.A (n_4307), .Y (n_4065));
NAND2X1 g133094(.A (n_4066), .B (P3_reg1[9] ), .Y (n_4431));
NOR2X1 g133088(.A (n_3911), .B (n_13361), .Y (n_4589));
OR2X1 g133100(.A (n_4133), .B (n_4132), .Y (n_4430));
AOI21X1 g132564(.A0 (n_2651), .A1 (n_3642), .B0 (n_3230), .Y(n_4061));
NOR2X1 g132613(.A (n_3399), .B (n_15968), .Y (n_4060));
AOI21X1 g133649(.A0 (n_3682), .A1 (n_2313), .B0 (n_4059), .Y(n_4568));
INVX1 g133430(.A (n_4271), .Y (n_4155));
NAND2X1 g133932(.A (n_4080), .B (n_3684), .Y (n_4058));
NOR2X1 g132763(.A (n_4056), .B (n_3743), .Y (n_32106));
INVX1 g133797(.A (n_4301), .Y (n_4055));
NAND2X1 g133917(.A (n_4053), .B (n_3703), .Y (n_4054));
NAND2X1 g132023(.A (n_3801), .B (n_2665), .Y (n_4052));
INVX1 g133421(.A (n_4051), .Y (n_6988));
AOI21X1 g131786(.A0 (n_4049), .A1 (n_2800), .B0 (n_2607), .Y(n_4050));
NOR2X1 g132713(.A (n_4205), .B (P2_reg2[18] ), .Y (n_4932));
NAND2X1 g133070(.A (n_3768), .B (n_1423), .Y (n_35335));
NAND2X1 g132698(.A (n_4046), .B (n_4045), .Y (n_4766));
NAND2X1 g133066(.A (n_3694), .B (n_609), .Y (n_33052));
NAND3X1 g133169(.A (n_3811), .B (n_1424), .C (n_3604), .Y (n_4043));
NAND2X1 g131998(.A (n_3984), .B (n_3433), .Y (n_4042));
INVX1 g133614(.A (n_4240), .Y (n_4041));
NOR2X1 g133573(.A (n_4234), .B (n_4185), .Y (n_4756));
OR2X1 g132647(.A (n_4040), .B (n_4039), .Y (n_4915));
NAND2X1 g131976(.A (n_3698), .B (n_4037), .Y (n_4038));
NAND2X1 g133233(.A (n_4099), .B (P2_reg1[10] ), .Y (n_4609));
NAND2X2 g132997(.A (n_1377), .B (n_3812), .Y (n_35195));
XOR2X1 g132172(.A (n_1073), .B (n_4035), .Y (n_4036));
NOR2X1 g133561(.A (n_4234), .B (n_4034), .Y (n_4726));
XOR2X1 g132166(.A (n_1137), .B (n_3606), .Y (n_4033));
MX2X1 g133052(.A (P3_IR[28] ), .B (n_1369), .S0 (n_3568), .Y(n_4032));
NOR2X1 g131954(.A (n_4025), .B (n_3456), .Y (n_4031));
NOR2X1 g132617(.A (n_10112), .B (n_4029), .Y (n_4030));
NAND2X1 g133521(.A (n_4249), .B (n_3758), .Y (n_4028));
AOI21X1 g133281(.A0 (n_4246), .A1 (n_4129), .B0 (n_4278), .Y(n_4437));
NOR2X1 g131674(.A (n_3449), .B (n_3834), .Y (n_4027));
NOR2X1 g132957(.A (n_886), .B (n_3819), .Y (n_4266));
INVX1 g133371(.A (n_6303), .Y (n_4026));
NAND3X1 g131933(.A (n_4025), .B (n_4024), .C (n_2292), .Y (n_4321));
INVX1 g133032(.A (n_4354), .Y (n_4188));
NAND2X1 g132665(.A (n_3999), .B (P3_reg1[18] ), .Y (n_5951));
AOI21X1 g133266(.A0 (n_4079), .A1 (n_4023), .B0 (n_4156), .Y(n_4421));
INVX1 g133868(.A (n_4305), .Y (n_4022));
XOR2X1 g132570(.A (n_1470), .B (n_3995), .Y (n_4021));
AOI21X1 g133265(.A0 (n_5914), .A1 (n_4020), .B0 (n_4019), .Y(n_4606));
INVX1 g132959(.A (n_34120), .Y (n_6170));
NAND2X1 g131566(.A (n_4017), .B (addr_490), .Y (n_4356));
NOR2X1 g133553(.A (n_4119), .B (n_3993), .Y (n_4574));
XOR2X1 g131881(.A (n_3524), .B (n_5586), .Y (so[3]));
NAND3X1 g132332(.A (n_4015), .B (n_3630), .C (n_4014), .Y (n_4353));
NOR2X1 g132427(.A (n_4012), .B (n_3787), .Y (n_4013));
NOR2X1 g133234(.A (n_3870), .B (n_4011), .Y (n_4600));
XOR2X1 g133708(.A (n_2460), .B (n_3628), .Y (n_4009));
INVX1 g133377(.A (n_4007), .Y (n_4170));
NOR2X1 g133208(.A (n_3836), .B (n_3472), .Y (n_5861));
NAND3X1 g133300(.A (n_3561), .B (n_4260), .C (n_3770), .Y (n_4473));
NOR2X1 g133916(.A (n_4079), .B (n_3760), .Y (n_4647));
NOR2X1 g133549(.A (n_4225), .B (n_4005), .Y (n_4644));
NOR2X1 g133576(.A (n_4145), .B (n_4004), .Y (n_4650));
INVX1 g132999(.A (n_4003), .Y (n_4285));
NAND2X1 g132400(.A (n_3704), .B (n_609), .Y (n_4002));
NAND2X1 g132678(.A (n_3999), .B (P3_reg2[18] ), .Y (n_5940));
NOR2X1 g133534(.A (n_4278), .B (n_3764), .Y (n_5300));
NAND2X1 g133572(.A (n_4162), .B (n_3685), .Y (n_3997));
XOR2X1 g132171(.A (n_1708), .B (n_3618), .Y (n_4313));
OAI21X1 g132501(.A0 (n_3995), .A1 (n_2899), .B0 (n_3532), .Y(n_3996));
NOR2X1 g133581(.A (n_4072), .B (n_4034), .Y (n_4575));
NOR2X1 g133892(.A (n_3751), .B (n_3993), .Y (n_3994));
MX2X1 g133051(.A (P3_IR[30] ), .B (n_594), .S0 (n_3646), .Y(n_3992));
OAI21X1 g133664(.A0 (n_3935), .A1 (n_3798), .B0 (n_4053), .Y(n_4468));
OR2X1 g132646(.A (n_3999), .B (P3_reg1[18] ), .Y (n_6079));
NOR2X1 g132609(.A (n_3494), .B (P2_n_749), .Y (n_3991));
NAND2X1 g133171(.A (n_3990), .B (n_4460), .Y (n_4262));
NAND2X1 g133106(.A (n_3911), .B (P3_reg1[7] ), .Y (n_4377));
NAND2X1 g132204(.A (n_3841), .B (n_3884), .Y (n_3989));
AOI21X1 g132088(.A0 (n_3938), .A1 (n_3954), .B0 (n_4012), .Y(n_4641));
NAND2X1 g131924(.A (n_3985), .B (n_3984), .Y (n_3986));
INVX1 g132971(.A (n_4288), .Y (n_4311));
NAND2X2 g133431(.A (n_32015), .B (n_32016), .Y (n_4271));
INVX1 g133458(.A (n_3774), .Y (n_4067));
NAND2X1 g133626(.A (n_3983), .B (n_3982), .Y (n_4401));
XOR2X1 g132591(.A (n_1811), .B (n_3907), .Y (n_3981));
OAI21X1 g132502(.A0 (n_3906), .A1 (n_2657), .B0 (n_2727), .Y(n_3980));
AND2X1 g132527(.A (n_3660), .B (n_3912), .Y (n_3979));
OAI21X1 g133660(.A0 (n_3978), .A1 (n_3745), .B0 (n_3983), .Y(n_4247));
MX2X1 g133494(.A (n_1107), .B (P1_IR[28] ), .S0 (n_3495), .Y(n_3977));
XOR2X1 g131872(.A (n_1144), .B (n_3395), .Y (n_3976));
NOR2X1 g132371(.A (n_3955), .B (n_3653), .Y (n_3974));
INVX1 g133187(.A (n_34179), .Y (n_3973));
AND2X1 g133179(.A (n_5820), .B (n_34234), .Y (n_32055));
CLKBUFX2 g133027(.A (n_3971), .Y (n_6810));
INVX1 g133036(.A (n_34092), .Y (n_4006));
NOR2X1 g133608(.A (n_4129), .B (n_3978), .Y (n_4412));
NOR2X1 g133872(.A (n_3831), .B (n_4004), .Y (n_4400));
NAND3X1 g131715(.A (n_3534), .B (n_3299), .C (n_3968), .Y (n_3969));
XOR2X1 g132165(.A (n_1248), .B (n_3806), .Y (n_3967));
XOR2X1 g132936(.A (n_1672), .B (n_3553), .Y (n_3966));
NOR2X1 g132619(.A (n_10116), .B (n_3964), .Y (n_3965));
NAND2X1 g133933(.A (n_4091), .B (n_3663), .Y (n_4319));
OAI21X1 g133020(.A0 (n_3501), .A1 (n_1645), .B0 (n_1172), .Y(n_3962));
NAND2X1 g133033(.A (n_1554), .B (n_3580), .Y (n_4354));
NOR2X1 g133579(.A (n_4278), .B (n_4129), .Y (n_4577));
OAI21X1 g133045(.A0 (n_3477), .A1 (n_33566), .B0 (n_718), .Y(n_3961));
INVX1 g133295(.A (n_3960), .Y (n_5724));
NOR2X1 g133174(.A (n_3959), .B (n_3958), .Y (n_4711));
INVX1 g133763(.A (n_3957), .Y (n_4010));
NAND2X1 g133523(.A (n_4267), .B (n_4398), .Y (n_4420));
NOR2X1 g133195(.A (n_4131), .B (P2_reg2[9] ), .Y (n_4378));
NAND3X1 g132268(.A (n_3955), .B (n_2188), .C (n_1961), .Y (n_4937));
AND2X1 g132272(.A (n_3954), .B (n_3928), .Y (n_4307));
NOR2X1 g132410(.A (n_3927), .B (addr_491), .Y (n_4519));
INVX1 g133808(.A (n_4267), .Y (n_3953));
AOI21X1 g132529(.A0 (n_3879), .A1 (n_3951), .B0 (n_3672), .Y(n_3952));
AOI21X1 g132530(.A0 (n_3947), .A1 (n_3800), .B0 (n_3793), .Y(n_3950));
NAND4X1 g132566(.A (n_3381), .B (n_1365), .C (n_3374), .D (n_2719),.Y (n_3949));
XOR2X1 g132592(.A (n_1446), .B (n_3947), .Y (n_3948));
NOR2X1 g132621(.A (n_3995), .B (n_3945), .Y (n_3946));
OAI21X1 g132633(.A0 (n_3804), .A1 (n_3943), .B0 (n_3942), .Y(n_3944));
INVX1 g132972(.A (n_3941), .Y (n_4288));
NOR2X1 g132738(.A (n_3671), .B (n_2569), .Y (n_3940));
NOR2X1 g132788(.A (n_3938), .B (n_3655), .Y (n_3939));
NAND2X1 g133518(.A (n_4298), .B (n_3643), .Y (n_3937));
AOI21X1 g132894(.A0 (n_3518), .A1 (n_2999), .B0 (n_2026), .Y(n_3936));
INVX1 g133444(.A (n_4040), .Y (n_4200));
NOR2X1 g133863(.A (n_3935), .B (n_3749), .Y (n_4465));
OR2X1 g133254(.A (n_3670), .B (n_3742), .Y (n_3933));
INVX1 g133290(.A (n_33681), .Y (n_3932));
OAI21X1 g132989(.A0 (n_3408), .A1 (n_3596), .B0 (n_985), .Y (n_3930));
AOI21X1 g132094(.A0 (n_3679), .A1 (n_3928), .B0 (n_3938), .Y(n_4504));
NAND2X1 g132301(.A (n_3927), .B (addr_491), .Y (n_4487));
INVX2 g133372(.A (n_3723), .Y (n_6303));
INVX1 g132348(.A (n_3984), .Y (n_3926));
CLKBUFX1 g133425(.A (n_3925), .Y (n_6348));
NAND2X1 g133537(.A (n_3664), .B (n_3923), .Y (n_4531));
INVX1 g133901(.A (n_4253), .Y (n_3922));
AOI21X1 g133658(.A0 (n_3921), .A1 (n_4556), .B0 (n_3920), .Y(n_4955));
OAI21X1 g133716(.A0 (n_3765), .A1 (n_4917), .B0 (n_3641), .Y(n_3919));
INVX1 g133785(.A (n_4099), .Y (n_3917));
INVX1 g133832(.A (n_4023), .Y (n_3916));
INVX1 g133842(.A (n_3982), .Y (n_3915));
INVX1 g133468(.A (n_3914), .Y (n_4141));
INVX1 g133875(.A (n_4149), .Y (n_3913));
OAI21X1 g132063(.A0 (n_3491), .A1 (n_1747), .B0 (n_3912), .Y(n_4073));
NOR2X1 g133923(.A (n_3978), .B (n_3635), .Y (n_4408));
NOR2X1 g133114(.A (n_3911), .B (P3_reg1[7] ), .Y (n_4708));
NAND2X1 g133452(.A (n_1267), .B (n_3650), .Y (n_3987));
INVX1 g134128(.A (n_3566), .Y (n_8115));
INVX1 g133463(.A (n_34014), .Y (n_4068));
NOR2X1 g132851(.A (n_3654), .B (n_1935), .Y (n_3910));
INVX1 g133819(.A (n_4244), .Y (n_3909));
AOI21X1 g132270(.A0 (n_3907), .A1 (n_2850), .B0 (n_3380), .Y(n_3908));
XOR2X1 g132586(.A (n_1602), .B (n_3906), .Y (n_4201));
NAND2X1 g132797(.A (n_6346), .B (n_31647), .Y (n_3905));
AOI21X1 g132525(.A0 (n_3556), .A1 (n_2707), .B0 (n_147), .Y (n_3904));
NOR2X1 g132257(.A (n_3666), .B (n_3902), .Y (n_3903));
NOR2X1 g133248(.A (n_4099), .B (P2_reg2[10] ), .Y (n_4546));
OAI21X1 g134047(.A0 (n_3125), .A1 (n_3899), .B0 (n_3663), .Y(n_4304));
NOR2X1 g132839(.A (n_3652), .B (n_2558), .Y (n_3897));
INVX1 g132882(.A (n_3796), .Y (n_3896));
AOI21X1 g132515(.A0 (n_3533), .A1 (n_3894), .B0 (n_3893), .Y(n_3895));
INVX1 g132913(.A (n_3891), .Y (n_3892));
NAND3X1 g132509(.A (n_2367), .B (n_3413), .C (n_2991), .Y (n_3890));
NAND3X1 g132727(.A (n_2913), .B (n_3512), .C (n_3674), .Y (n_3888));
NAND2X1 g132734(.A (n_3631), .B (n_3273), .Y (n_4286));
INVX1 g133887(.A (n_4148), .Y (n_3886));
NOR2X1 g132745(.A (n_3884), .B (n_2328), .Y (n_3885));
INVX1 g133409(.A (n_4046), .Y (n_8105));
INVX1 g133791(.A (n_4131), .Y (n_3883));
INVX1 g133406(.A (n_33176), .Y (n_6214));
INVX1 g133000(.A (n_3881), .Y (n_4003));
NAND2X1 g133615(.A (n_4091), .B (n_4023), .Y (n_4240));
NAND2X1 g133378(.A (n_3648), .B (n_3478), .Y (n_4007));
OAI21X1 g133030(.A0 (n_3500), .A1 (n_99), .B0 (n_1324), .Y (n_32639));
XOR2X1 g132571(.A (n_1740), .B (n_3879), .Y (n_3880));
AOI21X1 g131962(.A0 (n_3457), .A1 (n_3182), .B0 (n_1883), .Y(n_3878));
NAND2X1 g133257(.A (n_33140), .B (n_3852), .Y (n_4092));
INVX1 g133893(.A (n_4251), .Y (n_3877));
INVX1 g132949(.A (n_3876), .Y (n_6467));
INVX1 g133821(.A (n_4119), .Y (n_3873));
OR2X1 g133258(.A (n_3870), .B (n_3869), .Y (n_3871));
INVX1 g133259(.A (n_34502), .Y (n_3868));
NAND2X1 g133909(.A (n_3865), .B (n_3683), .Y (n_3866));
OAI21X1 g132522(.A0 (n_3860), .A1 (n_2649), .B0 (n_2864), .Y(n_3864));
INVX1 g133774(.A (n_3863), .Y (n_4461));
INVX1 g133768(.A (n_3862), .Y (n_4217));
NAND2X1 g133556(.A (n_3640), .B (n_3861), .Y (n_4409));
XOR2X1 g132583(.A (n_1378), .B (n_3860), .Y (n_4164));
INVX1 g134145(.A (n_4072), .Y (n_3859));
OR2X1 g133255(.A (n_3855), .B (n_3854), .Y (n_3856));
NAND2X1 g132872(.A (n_3852), .B (n_3851), .Y (n_3853));
XOR2X1 g133704(.A (n_4802), .B (n_3849), .Y (n_3850));
OR2X1 g132660(.A (n_32445), .B (n_3848), .Y (n_5063));
OR2X1 g131977(.A (n_3661), .B (n_3585), .Y (n_3847));
NOR2X1 g133522(.A (n_3935), .B (n_4005), .Y (n_4414));
INVX2 g133422(.A (n_34073), .Y (n_4051));
INVX1 g132773(.A (n_3841), .Y (n_3842));
INVX1 g133479(.A (n_34428), .Y (n_4157));
AOI21X1 g133643(.A0 (n_3983), .A1 (n_3759), .B0 (n_3978), .Y(n_4300));
NAND2X1 g133610(.A (n_4246), .B (n_3982), .Y (n_4195));
NAND2X1 g132310(.A (n_4118), .B (n_3954), .Y (n_4110));
NOR2X1 g133557(.A (n_3576), .B (n_4243), .Y (n_3838));
INVX1 g133559(.A (n_3836), .Y (n_3837));
NOR2X1 g133543(.A (n_3343), .B (n_3834), .Y (n_3835));
NOR2X1 g133862(.A (n_3629), .B (n_3826), .Y (n_3833));
OAI21X1 g133666(.A0 (n_3825), .A1 (n_3993), .B0 (n_3832), .Y(n_4259));
OAI21X1 g133668(.A0 (n_3831), .A1 (n_3823), .B0 (n_3865), .Y(n_4254));
AOI22X1 g133469(.A0 (n_3342), .A1 (n_852), .B0 (n_284), .B1(n_34093), .Y (n_3914));
INVX1 g133619(.A (n_3829), .Y (n_3830));
NAND3X1 g133286(.A (n_3590), .B (n_2387), .C (n_3591), .Y (n_3828));
NOR2X1 g133936(.A (n_3471), .B (P3_reg1[6] ), .Y (n_4075));
CLKBUFX1 g133441(.A (n_34231), .Y (n_4205));
OAI21X1 g133665(.A0 (n_3826), .A1 (n_3771), .B0 (n_3825), .Y(n_4019));
AND2X1 g134306(.A (n_3823), .B (n_3822), .Y (n_3824));
XOR2X1 g132939(.A (n_1272), .B (n_3530), .Y (n_3821));
NAND2X1 g133970(.A (n_3849), .B (n_4556), .Y (n_3820));
OAI21X1 g132950(.A0 (n_3347), .A1 (n_34093), .B0 (n_1237), .Y(n_3876));
AOI21X1 g133235(.A0 (n_3345), .A1 (n_3246), .B0 (n_3196), .Y(n_3819));
MX2X1 g132978(.A (n_1964), .B (n_212), .S0 (n_3338), .Y (n_3817));
OAI21X1 g134008(.A0 (n_3762), .A1 (n_3637), .B0 (n_3823), .Y(n_4081));
NOR2X1 g133160(.A (n_3815), .B (n_2278), .Y (n_3816));
XOR2X1 g132578(.A (n_1225), .B (n_3726), .Y (n_3814));
NOR2X1 g132453(.A (n_3423), .B (n_3659), .Y (n_3813));
NAND2X1 g133071(.A (n_3406), .B (n_3719), .Y (n_3812));
AOI21X1 g132915(.A0 (n_2798), .A1 (n_2595), .B0 (n_3551), .Y(n_4116));
NAND2X1 g133976(.A (n_1030), .B (n_3497), .Y (n_3811));
INVX1 g132921(.A (n_10110), .Y (n_13380));
XOR2X1 g131856(.A (n_1067), .B (n_3730), .Y (n_3809));
NOR2X1 g131900(.A (n_8511), .B (P1_n_449), .Y (n_3808));
NOR2X1 g132209(.A (n_3806), .B (n_2339), .Y (n_4025));
OAI21X1 g132212(.A0 (n_2645), .A1 (n_3468), .B0 (n_3804), .Y(n_3805));
AND2X1 g132349(.A (n_3928), .B (n_3680), .Y (n_3984));
NOR2X1 g133822(.A (n_3367), .B (n_3716), .Y (n_4119));
AOI21X1 g132503(.A0 (n_3315), .A1 (n_2588), .B0 (n_126), .Y (n_3803));
AOI21X1 g132520(.A0 (n_3388), .A1 (n_2610), .B0 (n_194), .Y (n_3802));
NAND4X1 g132528(.A (n_3947), .B (n_2536), .C (n_4179), .D (n_3800),.Y (n_3801));
AND2X1 g133859(.A (n_3798), .B (n_3797), .Y (n_3799));
AOI21X1 g132883(.A0 (n_3285), .A1 (n_3795), .B0 (n_3547), .Y(n_3796));
NOR2X1 g134223(.A (n_3899), .B (n_3589), .Y (n_4175));
AOI21X1 g132893(.A0 (n_3793), .A1 (n_4179), .B0 (n_3792), .Y(n_3794));
XOR2X1 g132580(.A (n_1475), .B (n_3594), .Y (n_3791));
XOR2X1 g132582(.A (n_1413), .B (n_3521), .Y (n_3790));
NAND2X1 g132643(.A (n_3740), .B (n_2789), .Y (n_3789));
XOR2X1 g132934(.A (n_1844), .B (n_3700), .Y (n_3788));
INVX1 g132728(.A (n_3954), .Y (n_3787));
NAND2X1 g132771(.A (n_3520), .B (n_3785), .Y (n_3786));
NAND3X1 g132774(.A (n_3522), .B (n_3188), .C (n_3001), .Y (n_3841));
MX2X1 g133050(.A (P2_IR[30] ), .B (n_100), .S0 (n_3304), .Y(n_3784));
OR2X1 g133054(.A (n_3505), .B (P2_IR[29] ), .Y (n_3783));
NOR2X1 g133057(.A (n_3198), .B (n_3834), .Y (n_3782));
NAND2X1 g133062(.A (n_3440), .B (n_609), .Y (n_3781));
NAND2X1 g133083(.A (n_3431), .B (n_1423), .Y (n_35283));
NAND2X1 g133127(.A (n_10582), .B (n_7243), .Y (n_3779));
NAND2X1 g133206(.A (n_13327), .B (n_7243), .Y (n_3778));
OAI21X1 g133347(.A0 (n_3404), .A1 (P2_reg3[28] ), .B0 (n_3405), .Y(n_8447));
NAND3X1 g133268(.A (n_3613), .B (n_2294), .C (n_3612), .Y (n_3777));
INVX1 g133411(.A (n_3736), .Y (n_3776));
INVX1 g133417(.A (n_3775), .Y (n_3845));
OAI21X1 g133459(.A0 (n_3303), .A1 (n_1277), .B0 (n_1117), .Y(n_3774));
INVX1 g133491(.A (n_33901), .Y (n_3999));
NAND2X1 g134308(.A (n_3771), .B (n_3770), .Y (n_3772));
NOR2X1 g133624(.A (n_4229), .B (n_4156), .Y (n_4495));
NAND2X1 g133681(.A (n_3391), .B (n_3528), .Y (n_3768));
NAND2X1 g132837(.A (n_3421), .B (n_3368), .Y (n_3767));
XOR2X1 g133715(.A (n_4523), .B (n_3765), .Y (n_3766));
CLKBUFX1 g133746(.A (n_3855), .Y (n_4133));
INVX1 g133756(.A (n_3854), .Y (n_4066));
INVX1 g133811(.A (n_4246), .Y (n_3764));
NAND2X1 g133876(.A (n_6962), .B (n_3709), .Y (n_4149));
NOR2X1 g133884(.A (n_3831), .B (n_3762), .Y (n_4255));
NOR2X1 g133889(.A (n_3307), .B (P2_reg1[6] ), .Y (n_4252));
NAND2X1 g133894(.A (n_6964), .B (P2_reg1[6] ), .Y (n_4251));
NOR2X1 g133928(.A (n_3308), .B (P2_reg1[5] ), .Y (n_4225));
NAND2X1 g133130(.A (n_3536), .B (n_3719), .Y (n_3761));
INVX1 g134154(.A (n_4091), .Y (n_3760));
NOR2X1 g134222(.A (n_3759), .B (n_3541), .Y (n_4166));
INVX1 g133940(.A (n_4034), .Y (n_3758));
XOR2X1 g132931(.A (n_1680), .B (n_3658), .Y (n_3754));
OR2X1 g132847(.A (n_2659), .B (n_3906), .Y (n_3753));
NAND2X1 g134162(.A (n_3752), .B (P2_reg1[3] ), .Y (n_4053));
OAI21X1 g133426(.A0 (n_3296), .A1 (n_3705), .B0 (n_1072), .Y(n_3925));
INVX1 g134160(.A (n_3832), .Y (n_3751));
INVX1 g132786(.A (n_4117), .Y (n_3750));
OAI21X1 g133669(.A0 (n_3749), .A1 (n_3231), .B0 (n_3798), .Y(n_4257));
OAI21X1 g134010(.A0 (n_3681), .A1 (n_3560), .B0 (n_3771), .Y(n_4059));
NAND2X1 g133902(.A (n_6962), .B (P2_reg1[5] ), .Y (n_4253));
AND2X1 g133890(.A (n_3747), .B (n_3797), .Y (n_3748));
NAND2X1 g134147(.A (n_3752), .B (P2_reg2[3] ), .Y (n_4224));
NAND3X1 g132345(.A (n_3548), .B (n_3725), .C (n_3283), .Y (n_3746));
NAND2X1 g133913(.A (n_3983), .B (n_3745), .Y (n_4196));
XOR2X1 g131861(.A (n_1504), .B (n_3707), .Y (n_4017));
OR2X1 g133246(.A (n_3583), .B (n_3743), .Y (n_3744));
CLKBUFX1 g133799(.A (n_3742), .Y (n_4301));
NOR2X1 g133926(.A (n_6964), .B (n_3724), .Y (n_4185));
AOI21X1 g132215(.A0 (n_2802), .A1 (n_3425), .B0 (n_3740), .Y(n_3741));
NOR2X1 g134146(.A (n_3752), .B (P2_reg2[3] ), .Y (n_4072));
NAND4X1 g132708(.A (n_3531), .B (n_3420), .C (n_2391), .D (n_2849),.Y (n_4855));
INVX1 g133067(.A (n_6346), .Y (n_3739));
OAI21X1 g132211(.A0 (n_3738), .A1 (n_3432), .B0 (n_3737), .Y(n_3985));
INVX1 g133410(.A (n_3736), .Y (n_4046));
NOR2X1 g133878(.A (n_3978), .B (n_3759), .Y (n_4248));
NAND2X1 g133185(.A (n_3452), .B (P2_IR[31] ), .Y (n_32579));
NAND2X1 g133820(.A (n_3367), .B (n_3693), .Y (n_4244));
AOI21X1 g131795(.A0 (n_3730), .A1 (n_2623), .B0 (n_2302), .Y(n_3731));
INVX2 g133775(.A (n_3728), .Y (n_3863));
AOI21X1 g132449(.A0 (n_3726), .A1 (n_3725), .B0 (n_3284), .Y(n_3727));
NAND2X1 g133560(.A (n_3170), .B (n_3546), .Y (n_3836));
NAND2X1 g133888(.A (n_6964), .B (n_3724), .Y (n_4148));
NAND2X1 g133870(.A (n_3471), .B (P3_reg2[6] ), .Y (n_4305));
MX2X1 g133373(.A (n_686), .B (P1_IR[26] ), .S0 (n_3288), .Y(n_3723));
INVX1 g133764(.A (n_34435), .Y (n_3957));
NAND2X1 g133085(.A (n_3502), .B (n_3719), .Y (n_3720));
NAND2X1 g133814(.A (n_3367), .B (n_3716), .Y (n_4250));
XOR2X1 g134097(.A (n_2428), .B (n_3270), .Y (n_3715));
INVX1 g133769(.A (n_3852), .Y (n_3862));
AND2X1 g133865(.A (n_3713), .B (n_3688), .Y (n_3714));
NOR2X1 g133927(.A (n_6962), .B (n_3709), .Y (n_4234));
MX2X1 g133366(.A (n_165), .B (P3_reg3[22] ), .S0 (n_3325), .Y(n_3887));
OAI21X1 g131680(.A0 (n_3707), .A1 (n_2457), .B0 (n_2690), .Y(n_3708));
NOR2X1 g133921(.A (n_3471), .B (P3_reg2[6] ), .Y (n_4433));
OAI21X1 g133028(.A0 (n_3348), .A1 (n_3705), .B0 (n_1207), .Y(n_3971));
OAI21X1 g132900(.A0 (n_2598), .A1 (n_2766), .B0 (n_3442), .Y(n_4015));
NAND2X1 g133261(.A (n_3586), .B (n_3447), .Y (n_4056));
MX2X1 g133007(.A (P1_IR[29] ), .B (n_252), .S0 (n_3351), .Y(n_3704));
INVX1 g134138(.A (n_3935), .Y (n_3703));
OAI21X1 g133662(.A0 (n_3702), .A1 (n_3350), .B0 (n_3701), .Y(n_4142));
AOI21X1 g132914(.A0 (n_3700), .A1 (n_2414), .B0 (n_3411), .Y(n_3891));
NAND2X1 g132511(.A (n_3529), .B (n_3697), .Y (n_3698));
MX2X1 g133687(.A (n_367), .B (P2_IR[23] ), .S0 (n_3341), .Y(n_3695));
MX2X1 g133683(.A (P1_IR[23] ), .B (n_211), .S0 (n_3326), .Y(n_3694));
NOR2X1 g133818(.A (n_3367), .B (n_3693), .Y (n_4145));
NAND3X1 g133296(.A (n_3201), .B (n_3162), .C (n_3490), .Y (n_3960));
NAND2X1 g133618(.A (n_10100), .B (n_7243), .Y (n_3691));
NOR2X1 g133611(.A (n_4156), .B (n_4079), .Y (n_4460));
NAND2X1 g133159(.A (n_3508), .B (n_1373), .Y (n_3690));
AND2X1 g133861(.A (n_3701), .B (n_3688), .Y (n_3689));
INVX1 g133074(.A (n_3687), .Y (n_6292));
AOI22X1 g132973(.A0 (n_3366), .A1 (n_3686), .B0 (P3_IR[17] ), .B1(n_1870), .Y (n_3941));
INVX1 g133911(.A (n_4005), .Y (n_3685));
OAI21X1 g133001(.A0 (n_3336), .A1 (n_1486), .B0 (n_1204), .Y(n_3881));
INVX1 g134170(.A (n_4004), .Y (n_3684));
INVX1 g134268(.A (n_3831), .Y (n_3683));
NAND2X1 g133412(.A (n_1275), .B (n_3311), .Y (n_3736));
NOR2X1 g134298(.A (n_3559), .B (n_3681), .Y (n_3682));
AOI21X1 g132090(.A0 (n_3523), .A1 (n_3680), .B0 (n_3679), .Y(n_4457));
NOR2X1 g134171(.A (n_3334), .B (n_3668), .Y (n_4004));
OAI21X1 g134033(.A0 (n_3678), .A1 (n_3759), .B0 (n_3745), .Y(n_3920));
OR2X1 g131922(.A (n_2459), .B (n_3707), .Y (n_3676));
OAI21X1 g132904(.A0 (n_3674), .A1 (n_2395), .B0 (n_2724), .Y(n_3675));
AOI22X1 g132919(.A0 (n_2560), .A1 (n_3209), .B0 (n_2447), .B1(n_3672), .Y (n_3673));
NOR2X1 g133912(.A (n_6963), .B (P2_reg1[4] ), .Y (n_4005));
INVX1 g133306(.A (n_3907), .Y (n_3671));
AOI21X1 g133971(.A0 (n_3663), .A1 (n_3362), .B0 (n_3899), .Y(n_3923));
CLKBUFX1 g133793(.A (n_3670), .Y (n_4131));
NOR2X1 g132343(.A (n_3679), .B (n_3361), .Y (n_3669));
NAND2X1 g133812(.A (n_3444), .B (n_13498), .Y (n_4246));
NAND2X1 g134163(.A (n_3334), .B (n_3668), .Y (n_4080));
NAND2X1 g133081(.A (n_3370), .B (n_3656), .Y (n_32215));
AOI21X1 g133294(.A0 (n_2932), .A1 (n_3252), .B0 (n_3335), .Y(n_3902));
NAND2X1 g132344(.A (n_2491), .B (n_3666), .Y (n_5194));
MX2X1 g132922(.A (P3_reg3[26] ), .B (n_3108), .S0 (n_3232), .Y(n_10110));
INVX1 g134686(.A (n_3752), .Y (n_3665));
NAND3X1 g133977(.A (n_3126), .B (n_3125), .C (n_3663), .Y (n_3664));
NAND2X1 g133844(.A (n_3450), .B (n_13511), .Y (n_3982));
NAND2X1 g132729(.A (n_3563), .B (addr_488), .Y (n_3954));
NAND2X1 g132391(.A (n_3300), .B (n_3661), .Y (n_5586));
NAND2X1 g132629(.A (n_3659), .B (n_3492), .Y (n_3660));
NAND4X1 g132927(.A (n_3658), .B (n_3511), .C (n_3386), .D (n_3894),.Y (n_4638));
NAND2X2 g133574(.A (n_3377), .B (n_3656), .Y (n_3657));
INVX1 g133212(.A (n_3928), .Y (n_3655));
AOI21X1 g133287(.A0 (n_3653), .A1 (n_1961), .B0 (n_3139), .Y(n_3654));
NOR2X1 g133910(.A (n_3826), .B (n_3681), .Y (n_4020));
INVX1 g133303(.A (n_3879), .Y (n_3652));
NOR2X1 g133496(.A (n_10114), .B (n_4029), .Y (n_3651));
NAND2X1 g133498(.A (n_3385), .B (n_33567), .Y (n_3650));
NAND2X1 g133540(.A (n_3306), .B (P3_IR[25] ), .Y (n_3648));
AND2X1 g133508(.A (n_9337), .B (n_34700), .Y (n_3647));
NAND4X1 g133571(.A (n_1965), .B (n_3310), .C (n_32450), .D (n_3309),.Y (n_3646));
NOR2X1 g133593(.A (n_8515), .B (P1_n_449), .Y (n_3645));
OR4X1 g133620(.A (n_3298), .B (n_2955), .C (P1_IR[29] ), .D(n_1108), .Y (n_3829));
OAI21X1 g133744(.A0 (n_3210), .A1 (n_3474), .B0 (n_861), .Y (n_3644));
INVX1 g133839(.A (n_4299), .Y (n_3643));
NAND2X1 g133919(.A (n_6963), .B (n_3565), .Y (n_4249));
INVX1 g133135(.A (n_3860), .Y (n_3642));
NAND2X1 g133990(.A (n_3765), .B (n_4917), .Y (n_3641));
AOI21X1 g133995(.A0 (n_3745), .A1 (n_3203), .B0 (n_3759), .Y(n_3861));
NAND3X1 g133999(.A (n_3204), .B (n_3678), .C (n_3745), .Y (n_3640));
NOR2X1 g134195(.A (n_3638), .B (n_3762), .Y (n_3639));
OAI21X1 g134011(.A0 (n_2460), .A1 (n_3638), .B0 (n_3637), .Y(n_5956));
XOR2X1 g134087(.A (n_2076), .B (n_3173), .Y (n_3636));
INVX1 g134136(.A (n_3983), .Y (n_3635));
OR2X1 g133055(.A (n_3504), .B (n_2504), .Y (n_3634));
NOR2X1 g133829(.A (n_3450), .B (n_13511), .Y (n_4129));
NAND3X1 g133270(.A (n_3552), .B (n_3630), .C (n_3441), .Y (n_3631));
INVX1 g134264(.A (n_3825), .Y (n_3629));
NAND2X1 g134315(.A (n_3627), .B (n_3637), .Y (n_3628));
INVX1 g133446(.A (n_4040), .Y (n_3851));
NAND3X1 g132912(.A (n_3328), .B (n_3094), .C (n_3159), .Y (n_4035));
NOR2X1 g133813(.A (n_3444), .B (n_13498), .Y (n_4278));
INVX1 g133781(.A (n_3621), .Y (n_3959));
NOR2X1 g132787(.A (n_3605), .B (addr_489), .Y (n_4117));
OAI21X1 g132620(.A0 (n_3145), .A1 (n_2405), .B0 (n_2590), .Y(n_3618));
AND2X1 g133184(.A (n_3356), .B (n_3087), .Y (n_3995));
XOR2X1 g132573(.A (n_1258), .B (n_3486), .Y (n_3617));
XOR2X1 g132572(.A (n_3738), .B (n_3243), .Y (so[2]));
OR2X1 g133652(.A (n_3241), .B (n_3340), .Y (n_3615));
NAND2X1 g133563(.A (n_3613), .B (n_3612), .Y (n_3614));
INVX1 g133770(.A (n_3445), .Y (n_3852));
NAND2X1 g133602(.A (n_8055), .B (n_7243), .Y (n_3611));
OR2X1 g132505(.A (n_2790), .B (n_3570), .Y (n_3609));
INVX1 g133418(.A (n_34437), .Y (n_3775));
NOR2X1 g133075(.A (n_3179), .B (n_3349), .Y (n_3687));
NAND2X1 g132709(.A (n_3277), .B (n_3023), .Y (n_3606));
NAND2X1 g132754(.A (n_3605), .B (addr_489), .Y (n_4118));
NAND2X1 g133929(.A (n_728), .B (n_3496), .Y (n_3604));
OR2X1 g132495(.A (n_2733), .B (n_3567), .Y (n_3603));
AND2X1 g133056(.A (n_8207), .B (n_35023), .Y (n_3602));
INVX1 g133332(.A (n_3601), .Y (n_13387));
NOR2X1 g134139(.A (n_3752), .B (P2_reg1[3] ), .Y (n_3935));
INVX1 g133787(.A (n_3599), .Y (n_4099));
NOR2X1 g133570(.A (n_3329), .B (n_3346), .Y (n_5820));
NAND2X1 g133834(.A (n_3450), .B (P3_reg1[4] ), .Y (n_4023));
INVX2 g133757(.A (n_33140), .Y (n_3854));
NOR2X1 g132641(.A (n_3594), .B (n_2567), .Y (n_3955));
INVX1 g133800(.A (n_3593), .Y (n_3742));
NOR2X1 g133896(.A (n_3826), .B (n_3993), .Y (n_4260));
OAI21X1 g133061(.A0 (n_3141), .A1 (n_2793), .B0 (n_3312), .Y(n_3884));
NAND2X1 g133536(.A (n_3591), .B (n_3590), .Y (n_3592));
INVX1 g133747(.A (n_3586), .Y (n_3855));
INVX1 g132431(.A (n_3968), .Y (n_3585));
INVX1 g133751(.A (n_3583), .Y (n_3911));
AND2X1 g131901(.A (n_9209), .B (n_34309), .Y (n_3582));
OAI21X1 g133777(.A0 (n_3258), .A1 (n_377), .B0 (n_858), .Y (n_3728));
NAND2X1 g133569(.A (n_3318), .B (n_1423), .Y (n_32015));
NAND2X1 g133078(.A (n_3282), .B (n_1423), .Y (n_3580));
NAND2X1 g132636(.A (n_3577), .B (n_2207), .Y (n_3578));
INVX1 g133815(.A (n_4242), .Y (n_3576));
NAND2X1 g133810(.A (n_3444), .B (P3_reg1[5] ), .Y (n_4267));
NAND2X1 g134161(.A (n_3334), .B (n_3333), .Y (n_3832));
XOR2X1 g132930(.A (n_1586), .B (n_3412), .Y (n_3927));
INVX1 g133352(.A (n_3573), .Y (n_13388));
NAND2X1 g132346(.A (n_3570), .B (n_3542), .Y (n_4049));
INVX1 g133335(.A (n_10112), .Y (n_13383));
NAND3X1 g133630(.A (n_2382), .B (n_1148), .C (n_3256), .Y (n_3568));
NAND2X1 g132329(.A (n_3567), .B (n_3207), .Y (n_4120));
INVX1 g134131(.A (n_3566), .Y (n_3869));
NOR2X1 g133941(.A (n_6963), .B (n_3565), .Y (n_4034));
NAND2X1 g133849(.A (n_6963), .B (P2_reg1[4] ), .Y (n_4162));
CLKBUFX1 g133068(.A (n_3564), .Y (n_6346));
NOR2X1 g132739(.A (n_3563), .B (addr_488), .Y (n_4012));
NAND2X1 g134194(.A (n_3561), .B (n_3560), .Y (n_3562));
OAI21X1 g134009(.A0 (n_2497), .A1 (n_3559), .B0 (n_3560), .Y(n_5914));
AND2X1 g132616(.A (n_13301), .B (n_35023), .Y (n_3558));
NOR2X1 g134278(.A (n_3759), .B (n_3203), .Y (n_3921));
NAND2X1 g134321(.A (n_3678), .B (n_3116), .Y (n_3849));
NAND3X1 g133368(.A (n_650), .B (n_3020), .C (addr_429), .Y (n_3556));
MX2X1 g133336(.A (P3_reg3[25] ), .B (n_158), .S0 (n_3059), .Y(n_10112));
INVX1 g133360(.A (n_10116), .Y (n_13385));
NAND2X1 g134300(.A (n_3472), .B (n_3470), .Y (n_3865));
INVX1 g134272(.A (n_3702), .Y (n_3688));
INVX1 g133633(.A (n_3552), .Y (n_3553));
INVX1 g134249(.A (n_3444), .Y (n_10740));
NAND3X1 g133304(.A (n_3169), .B (n_2959), .C (n_3193), .Y (n_3879));
OAI21X1 g133077(.A0 (n_3301), .A1 (n_2594), .B0 (n_3410), .Y(n_3551));
NAND2X1 g133582(.A (n_13375), .B (n_7243), .Y (n_3550));
NAND2X1 g132799(.A (n_11122), .B (n_15981), .Y (n_3549));
NOR2X1 g132849(.A (n_3360), .B (n_3547), .Y (n_3548));
INVX1 g133879(.A (n_3545), .Y (n_3546));
NOR2X1 g133904(.A (n_4079), .B (n_3899), .Y (n_4095));
AOI22X1 g133748(.A0 (n_3044), .A1 (n_33567), .B0 (n_434), .B1(n_33566), .Y (n_3586));
NOR2X1 g133836(.A (n_3045), .B (n_3416), .Y (n_4243));
OAI21X1 g133082(.A0 (n_3542), .A1 (n_2574), .B0 (n_2606), .Y(n_3740));
INVX1 g134528(.A (n_3745), .Y (n_3541));
NAND2X1 g133216(.A (n_8458), .B (n_1313), .Y (n_3540));
AOI21X1 g133648(.A0 (n_3206), .A1 (n_3538), .B0 (n_3537), .Y(n_3804));
MX2X1 g133803(.A (P2_IR[24] ), .B (n_561), .S0 (n_3026), .Y(n_3536));
XOR2X1 g133389(.A (n_3534), .B (n_3012), .Y (so[1]));
NAND2X1 g134156(.A (n_3162), .B (P3_reg1[3] ), .Y (n_4091));
AND2X1 g133198(.A (n_3223), .B (n_2421), .Y (n_3906));
INVX1 g133278(.A (n_3532), .Y (n_3533));
INVX1 g133514(.A (n_3530), .Y (n_3531));
NAND2X1 g132628(.A (n_3394), .B (n_2622), .Y (n_3529));
NAND2X1 g133937(.A (n_3245), .B (n_262), .Y (n_3528));
OAI21X1 g132860(.A0 (n_3065), .A1 (n_2483), .B0 (n_3526), .Y(n_3527));
XOR2X1 g132937(.A (n_1198), .B (n_3137), .Y (n_3525));
NAND2X1 g133183(.A (n_3190), .B (n_3143), .Y (n_3947));
NOR2X1 g133226(.A (n_3523), .B (n_3167), .Y (n_3524));
NOR2X1 g133245(.A (n_3451), .B (addr_487), .Y (n_3938));
INVX1 g133272(.A (n_3521), .Y (n_3522));
NAND2X1 g133298(.A (n_3220), .B (n_2775), .Y (n_3520));
NOR2X1 g133495(.A (n_10119), .B (n_4029), .Y (n_3519));
NAND2X1 g133500(.A (n_3419), .B (n_2391), .Y (n_3518));
AOI21X1 g132907(.A0 (n_3136), .A1 (n_3454), .B0 (n_3523), .Y(n_3737));
NOR2X1 g133511(.A (n_10103), .B (n_4029), .Y (n_3517));
NAND2X1 g133513(.A (n_2911), .B (n_15981), .Y (n_3516));
AND2X1 g133527(.A (n_3202), .B (n_3011), .Y (n_3514));
AND2X1 g133533(.A (n_7957), .B (n_35023), .Y (n_3513));
NAND2X1 g133587(.A (n_3153), .B (n_3511), .Y (n_3512));
NAND2X1 g133597(.A (n_3228), .B (n_3509), .Y (n_3510));
AOI21X1 g133631(.A0 (n_3507), .A1 (n_3506), .B0 (n_2282), .Y(n_3508));
INVX1 g133637(.A (n_3504), .Y (n_3505));
MX2X1 g133688(.A (n_516), .B (n_453), .S0 (n_3082), .Y (n_3502));
MX2X1 g133703(.A (n_1171), .B (P1_IR[15] ), .S0 (n_33674), .Y(n_3501));
MX2X1 g133720(.A (n_1323), .B (P3_IR[20] ), .S0 (n_3120), .Y(n_3500));
MX2X1 g133804(.A (P3_IR[24] ), .B (n_664), .S0 (n_3098), .Y(n_3498));
INVX1 g134240(.A (n_3397), .Y (n_6962));
INVX1 g134236(.A (n_3496), .Y (n_3497));
NAND3X1 g133962(.A (n_2001), .B (n_1360), .C (n_3056), .Y (n_3495));
INVX1 g133356(.A (n_3494), .Y (n_9512));
NAND2X1 g134028(.A (n_3177), .B (n_3678), .Y (n_5807));
NAND4X1 g132776(.A (n_3138), .B (n_3276), .C (n_2359), .D (n_3492),.Y (n_4634));
AOI21X1 g132918(.A0 (n_3275), .A1 (n_2359), .B0 (n_3375), .Y(n_3491));
INVX1 g133824(.A (n_3490), .Y (n_3743));
NAND2X1 g133817(.A (n_3045), .B (n_3402), .Y (n_4298));
MX2X1 g133333(.A (P3_reg3[28] ), .B (n_259), .S0 (n_3110), .Y(n_3601));
NAND2X2 g133447(.A (n_1212), .B (n_3224), .Y (n_4040));
INVX1 g134294(.A (n_3749), .Y (n_3797));
OR4X1 g132409(.A (n_3486), .B (n_3485), .C (n_1747), .D (n_3422), .Y(n_3487));
NAND2X1 g132855(.A (n_3191), .B (n_1313), .Y (n_3481));
XOR2X1 g132929(.A (n_1208), .B (n_3327), .Y (n_3479));
NAND2X1 g133541(.A (n_3305), .B (n_282), .Y (n_3478));
MX2X1 g133717(.A (n_439), .B (P3_IR[16] ), .S0 (n_3255), .Y(n_3477));
NAND2X1 g134265(.A (n_3472), .B (n_3235), .Y (n_3825));
INVX1 g134149(.A (n_3476), .Y (n_6964));
INVX1 g133801(.A (n_3280), .Y (n_3593));
INVX1 g133782(.A (n_3460), .Y (n_3621));
OAI21X1 g133069(.A0 (n_1487), .A1 (n_3226), .B0 (n_3227), .Y(n_3564));
NAND2X1 g133930(.A (n_3471), .B (P3_reg1[6] ), .Y (n_4398));
NOR2X1 g134269(.A (n_3472), .B (n_3470), .Y (n_3831));
XOR2X1 g132574(.A (n_1581), .B (n_3468), .Y (n_3469));
NAND2X1 g131997(.A (n_8164), .B (n_1313), .Y (n_3466));
INVX1 g133794(.A (n_34016), .Y (n_3670));
XOR2X1 g132577(.A (n_1262), .B (n_3320), .Y (n_3464));
INVX1 g134020(.A (n_3463), .Y (n_5825));
INVX4 g133736(.A (n_3462), .Y (n_3870));
NOR2X1 g134132(.A (n_715), .B (n_3249), .Y (n_3566));
NAND2X1 g132627(.A (n_3456), .B (n_2292), .Y (n_3457));
AND2X1 g132610(.A (n_13169), .B (n_35023), .Y (n_3455));
AND2X1 g132432(.A (n_3454), .B (n_3680), .Y (n_3968));
INVX1 g132143(.A (n_3453), .Y (n_10885));
MX2X1 g133710(.A (P2_IR[15] ), .B (n_632), .S0 (n_3379), .Y(n_3452));
NAND2X1 g133213(.A (n_3451), .B (addr_487), .Y (n_3928));
NOR2X1 g133827(.A (n_3450), .B (P3_reg1[4] ), .Y (n_4156));
AOI21X1 g132911(.A0 (n_835), .A1 (n_2496), .B0 (n_3194), .Y (n_3806));
INVX1 g132139(.A (n_3449), .Y (n_9345));
INVX1 g133752(.A (n_3447), .Y (n_3583));
OAI21X1 g133771(.A0 (n_3067), .A1 (n_33566), .B0 (n_1033), .Y(n_3445));
INVX1 g132558(.A (n_3372), .Y (n_8511));
NOR2X1 g133807(.A (n_3444), .B (P3_reg1[5] ), .Y (n_4229));
NAND3X1 g133629(.A (n_2032), .B (n_1091), .C (n_2998), .Y (n_3443));
AOI21X1 g133297(.A0 (n_3365), .A1 (n_3441), .B0 (n_3272), .Y(n_3442));
AND2X1 g133136(.A (n_3248), .B (n_2425), .Y (n_3860));
MX2X1 g133684(.A (P1_IR[19] ), .B (n_739), .S0 (n_3118), .Y(n_3440));
INVX1 g133788(.A (n_33540), .Y (n_3599));
INVX1 g134487(.A (n_3663), .Y (n_3589));
NAND2X1 g133505(.A (n_3181), .B (n_609), .Y (n_3438));
AND2X1 g133524(.A (n_10041), .B (n_3185), .Y (n_3436));
NAND2X1 g131992(.A (n_7819), .B (n_15981), .Y (n_3434));
INVX1 g133133(.A (n_3432), .Y (n_3433));
MX2X1 g133682(.A (P3_IR[19] ), .B (n_1666), .S0 (n_3074), .Y(n_3431));
AOI21X1 g133676(.A0 (n_3271), .A1 (n_4014), .B0 (n_3354), .Y(n_3815));
AOI21X1 g132334(.A0 (n_3096), .A1 (n_2552), .B0 (addr_461), .Y(n_3427));
XOR2X1 g132588(.A (n_1742), .B (n_3425), .Y (n_3426));
NOR2X1 g132632(.A (n_3486), .B (n_3422), .Y (n_3423));
NAND2X1 g134023(.A (n_3233), .B (n_3125), .Y (n_5624));
AOI21X1 g133271(.A0 (n_3323), .A1 (n_3420), .B0 (n_3419), .Y(n_3421));
NAND2X1 g133175(.A (n_10822), .B (n_3217), .Y (n_3418));
NAND2X1 g134137(.A (n_3162), .B (n_13358), .Y (n_3983));
NAND2X1 g133816(.A (n_3045), .B (n_3416), .Y (n_4242));
NOR2X1 g134167(.A (n_3162), .B (n_13358), .Y (n_3978));
OR2X1 g133177(.A (n_2407), .B (n_3412), .Y (n_3413));
INVX1 g134421(.A (n_3681), .Y (n_3770));
OAI21X1 g133084(.A0 (n_3410), .A1 (n_2434), .B0 (n_3316), .Y(n_3411));
MX2X1 g133686(.A (P3_IR[23] ), .B (n_545), .S0 (n_3062), .Y(n_3409));
MX2X1 g133695(.A (n_984), .B (P1_IR[17] ), .S0 (n_3115), .Y(n_3408));
MX2X1 g133353(.A (P3_reg3[27] ), .B (n_269), .S0 (n_3052), .Y(n_3573));
MX2X1 g133694(.A (P2_IR[19] ), .B (n_607), .S0 (n_3058), .Y(n_3406));
NAND2X1 g133601(.A (n_3404), .B (P2_reg3[28] ), .Y (n_3405));
NAND2X1 g132059(.A (n_7575), .B (n_3217), .Y (n_3403));
NAND3X1 g133307(.A (n_3008), .B (n_3114), .C (n_3146), .Y (n_3907));
NOR2X1 g133840(.A (n_3045), .B (n_3402), .Y (n_4299));
AND2X1 g133898(.A (n_3234), .B (n_3171), .Y (n_33010));
INVX1 g133339(.A (n_3399), .Y (n_10889));
INVX1 g134427(.A (n_3762), .Y (n_3822));
AOI21X1 g132214(.A0 (n_2466), .A1 (n_3199), .B0 (n_3394), .Y(n_3395));
XOR2X1 g133357(.A (P2_reg3[25] ), .B (n_2905), .Y (n_3494));
INVX1 g134017(.A (n_3393), .Y (n_3467));
NAND2X1 g133153(.A (n_3105), .B (n_15981), .Y (n_3392));
NAND2X1 g133848(.A (n_3244), .B (n_1878), .Y (n_3391));
NAND2X1 g132753(.A (n_3112), .B (n_2446), .Y (n_3390));
INVX1 g134361(.A (n_3471), .Y (n_3429));
XOR2X1 g133385(.A (n_1235), .B (n_3294), .Y (n_3389));
NOR2X1 g133825(.A (n_3192), .B (n_3257), .Y (n_3490));
NAND4X1 g133370(.A (n_3084), .B (addr_452), .C (addr_450), .D(addr_451), .Y (n_3388));
OAI21X1 g133358(.A0 (n_3003), .A1 (P1_reg3[28] ), .B0 (n_3004), .Y(n_13301));
MX2X1 g133361(.A (P3_reg3[21] ), .B (n_307), .S0 (n_2937), .Y(n_10116));
NOR2X1 g134422(.A (n_2943), .B (n_3337), .Y (n_3681));
NAND2X1 g131995(.A (n_3100), .B (n_3185), .Y (n_3387));
AOI21X1 g133279(.A0 (n_3254), .A1 (n_3386), .B0 (n_2725), .Y(n_3532));
NOR2X1 g134295(.A (n_6887), .B (P2_reg1[2] ), .Y (n_3749));
MX2X1 g134068(.A (P3_IR[12] ), .B (n_564), .S0 (n_2974), .Y(n_3385));
AOI22X1 g133753(.A0 (n_2934), .A1 (n_33567), .B0 (n_666), .B1(n_33566), .Y (n_3447));
INVX1 g134688(.A (n_34079), .Y (n_3752));
NAND2X1 g133180(.A (n_8467), .B (n_1313), .Y (n_3382));
NAND2X1 g133584(.A (n_2570), .B (n_3380), .Y (n_3381));
NAND4X1 g133638(.A (n_1391), .B (n_1623), .C (n_2830), .D (n_2876),.Y (n_3504));
NOR2X1 g133924(.A (n_1422), .B (n_3379), .Y (n_3590));
NOR2X1 g134273(.A (n_6887), .B (P2_reg2[2] ), .Y (n_3702));
MX2X1 g134093(.A (n_1646), .B (n_578), .S0 (n_3078), .Y (n_3377));
OR2X1 g133249(.A (n_3018), .B (n_3375), .Y (n_3659));
AOI21X1 g133659(.A0 (n_3373), .A1 (n_1989), .B0 (n_1914), .Y(n_3374));
MX2X1 g133697(.A (n_1401), .B (P1_IR[22] ), .S0 (n_2956), .Y(n_3370));
INVX1 g134150(.A (n_3307), .Y (n_3476));
NAND4X1 g134049(.A (n_3324), .B (n_3006), .C (n_2948), .D (n_3420),.Y (n_3368));
INVX1 g134353(.A (n_3367), .Y (n_3483));
MX2X1 g133685(.A (n_684), .B (P3_IR[17] ), .S0 (n_2915), .Y(n_3366));
OR2X1 g133634(.A (n_2599), .B (n_3365), .Y (n_3552));
AND2X1 g132612(.A (n_10032), .B (n_34309), .Y (n_3364));
NAND2X1 g132635(.A (n_3425), .B (n_2801), .Y (n_3570));
OR2X1 g134022(.A (n_3127), .B (n_3362), .Y (n_3463));
INVX1 g132778(.A (n_3680), .Y (n_3361));
INVX1 g133301(.A (n_3360), .Y (n_3726));
XOR2X1 g133340(.A (P1_reg3[25] ), .B (n_2896), .Y (n_3399));
XOR2X1 g133387(.A (n_1745), .B (n_3222), .Y (n_3563));
XOR2X1 g133398(.A (n_1611), .B (n_3313), .Y (n_3359));
NAND2X1 g133596(.A (n_13370), .B (n_7243), .Y (n_3357));
NAND3X1 g133635(.A (n_3107), .B (n_3050), .C (n_3086), .Y (n_3356));
AOI21X1 g133642(.A0 (n_3354), .A1 (n_3353), .B0 (n_3352), .Y(n_3355));
NAND4X1 g133647(.A (n_1657), .B (n_2135), .C (n_2806), .D (n_2834),.Y (n_3351));
OAI21X1 g134335(.A0 (n_2428), .A1 (n_3103), .B0 (n_3350), .Y(n_5972));
NAND2X1 g133677(.A (n_1309), .B (n_3027), .Y (n_3349));
MX2X1 g133692(.A (P1_IR[21] ), .B (n_1206), .S0 (n_2966), .Y(n_3348));
MX2X1 g133693(.A (P2_IR[21] ), .B (n_1236), .S0 (n_2967), .Y(n_3347));
NAND2X1 g133134(.A (n_3242), .B (n_3454), .Y (n_3432));
OR2X1 g133831(.A (n_3307), .B (n_34082), .Y (n_3346));
NAND2X1 g133858(.A (n_32951), .B (n_527), .Y (n_3345));
INVX1 g134105(.A (n_3343), .Y (n_10081));
NAND2X1 g134058(.A (n_3099), .B (n_2945), .Y (n_3342));
NAND2X1 g134142(.A (n_3075), .B (n_3057), .Y (n_3341));
OR2X1 g134183(.A (n_34082), .B (n_2663), .Y (n_3340));
NAND4X1 g133641(.A (n_1634), .B (n_1949), .C (n_2869), .D (n_2439),.Y (n_3338));
NOR2X1 g134279(.A (n_3899), .B (n_3362), .Y (n_3990));
NOR2X1 g134318(.A (n_3129), .B (n_3362), .Y (n_3765));
NAND2X1 g134434(.A (n_2943), .B (n_3337), .Y (n_3771));
INVX1 g134536(.A (n_3638), .Y (n_3627));
MX2X1 g133721(.A (n_287), .B (P2_IR[20] ), .S0 (n_2954), .Y(n_3336));
NAND2X1 g133497(.A (n_2794), .B (n_3091), .Y (n_3793));
OR2X1 g132772(.A (n_3468), .B (n_2280), .Y (n_3567));
INVX1 g133639(.A (n_3253), .Y (n_3335));
NOR2X1 g134158(.A (n_3334), .B (n_3333), .Y (n_3993));
NAND2X1 g133914(.A (n_8185), .B (n_1313), .Y (n_3331));
NAND2X1 g133725(.A (n_3048), .B (n_3010), .Y (n_13327));
OR2X1 g133905(.A (n_3308), .B (n_3239), .Y (n_3329));
NAND2X1 g133186(.A (n_3327), .B (n_2293), .Y (n_3328));
NAND2X1 g133880(.A (n_3147), .B (n_2962), .Y (n_3545));
NAND2X1 g134141(.A (n_3025), .B (n_3117), .Y (n_3326));
NAND3X1 g133853(.A (n_2361), .B (n_2360), .C (n_2767), .Y (n_3325));
NAND2X1 g134213(.A (n_6887), .B (P2_reg2[2] ), .Y (n_3701));
AOI21X1 g133515(.A0 (n_2949), .A1 (n_3324), .B0 (n_3323), .Y(n_3530));
MX2X1 g134133(.A (P1_IR[24] ), .B (n_658), .S0 (n_2884), .Y(n_3321));
OAI21X1 g133784(.A0 (n_2898), .A1 (n_998), .B0 (n_1020), .Y (n_3460));
NOR2X1 g132634(.A (n_3320), .B (n_2343), .Y (n_3666));
INVX1 g134115(.A (n_3184), .Y (n_8515));
NAND2X1 g132274(.A (n_3292), .B (n_3195), .Y (n_3730));
MX2X1 g134079(.A (P3_IR[14] ), .B (n_704), .S0 (n_32452), .Y(n_3318));
NAND2X1 g134429(.A (n_2943), .B (n_3259), .Y (n_3823));
OAI21X1 g133064(.A0 (n_3316), .A1 (n_2433), .B0 (n_2964), .Y(n_3577));
NAND4X1 g133369(.A (n_3070), .B (addr_488), .C (n_3314), .D(addr_487), .Y (n_3315));
XOR2X1 g133381(.A (n_1895), .B (n_3247), .Y (n_3605));
AOI21X1 g133273(.A0 (n_3313), .A1 (n_3189), .B0 (n_3142), .Y(n_3521));
XOR2X1 g132144(.A (P1_reg3[26] ), .B (n_2926), .Y (n_3453));
NOR2X1 g133567(.A (n_2644), .B (n_3002), .Y (n_3312));
NAND2X1 g133583(.A (n_3035), .B (n_3656), .Y (n_3311));
NAND3X1 g134237(.A (n_32450), .B (n_3310), .C (n_3309), .Y (n_3496));
NOR2X1 g133895(.A (n_3308), .B (n_3307), .Y (n_4137));
INVX1 g133873(.A (n_3305), .Y (n_3306));
NAND4X1 g133542(.A (n_1717), .B (n_2321), .C (n_2782), .D (n_1915),.Y (n_3304));
NOR2X1 g133860(.A (n_1583), .B (n_32951), .Y (n_3612));
NAND2X1 g134225(.A (n_6887), .B (P2_reg1[2] ), .Y (n_3798));
MX2X1 g134080(.A (n_488), .B (P1_IR[16] ), .S0 (n_3055), .Y(n_3303));
NAND2X1 g132710(.A (n_3047), .B (n_2413), .Y (n_3302));
NAND2X1 g133512(.A (n_2799), .B (n_3301), .Y (n_3700));
NAND2X1 g132688(.A (n_3534), .B (n_3299), .Y (n_3300));
NAND2X1 g134235(.A (n_1729), .B (n_3079), .Y (n_3298));
INVX2 g133737(.A (n_3151), .Y (n_3462));
MX2X1 g134112(.A (n_345), .B (P1_IR[20] ), .S0 (n_2885), .Y(n_3296));
INVX1 g134084(.A (n_3295), .Y (n_10100));
INVX1 g134440(.A (n_3559), .Y (n_3561));
AOI21X1 g133288(.A0 (n_3294), .A1 (n_3168), .B0 (n_2958), .Y(n_3594));
OR2X1 g132504(.A (n_2624), .B (n_3292), .Y (n_3293));
OAI21X1 g133538(.A0 (n_2444), .A1 (n_1841), .B0 (n_3152), .Y(n_3658));
NAND2X1 g133979(.A (n_3119), .B (n_609), .Y (n_3288));
NAND2X1 g133503(.A (n_3284), .B (n_3283), .Y (n_3285));
MX2X1 g133696(.A (n_657), .B (P3_IR[21] ), .S0 (n_2890), .Y(n_3282));
NAND2X1 g132201(.A (n_7737), .B (n_15981), .Y (n_3281));
OAI21X1 g133802(.A0 (n_2927), .A1 (n_3279), .B0 (n_752), .Y (n_3280));
XOR2X1 g133396(.A (n_1616), .B (n_3106), .Y (n_3278));
AOI21X1 g133269(.A0 (n_3043), .A1 (n_3276), .B0 (n_3275), .Y(n_3277));
AOI21X1 g132450(.A0 (n_2988), .A1 (n_3221), .B0 (n_2420), .Y(n_3707));
AOI21X1 g133283(.A0 (n_3272), .A1 (n_3630), .B0 (n_3271), .Y(n_3273));
NAND2X1 g134515(.A (n_3713), .B (n_3350), .Y (n_3270));
AND2X1 g132618(.A (n_13173), .B (n_35023), .Y (n_3268));
INVX1 g134241(.A (n_3308), .Y (n_3397));
NAND2X1 g133545(.A (n_3081), .B (n_33815), .Y (n_3266));
INVX1 g133622(.A (n_3263), .Y (n_3264));
INVX1 g133706(.A (n_3262), .Y (n_10582));
XOR2X1 g132140(.A (P2_reg3[26] ), .B (n_2977), .Y (n_3449));
NOR2X1 g134428(.A (n_2943), .B (n_3259), .Y (n_3762));
CLKBUFX1 g133403(.A (n_8001), .Y (n_11122));
MX2X1 g134397(.A (n_1800), .B (n_654), .S0 (n_2755), .Y (n_3258));
INVX1 g134362(.A (n_3257), .Y (n_3471));
INVX1 g134312(.A (n_3255), .Y (n_3256));
OAI21X1 g133367(.A0 (n_2917), .A1 (P1_reg3[27] ), .B0 (n_2918), .Y(n_13169));
AOI21X1 g133632(.A0 (n_3085), .A1 (n_2679), .B0 (n_3254), .Y(n_3674));
XOR2X1 g134106(.A (P2_reg3[24] ), .B (n_2758), .Y (n_3343));
AOI22X1 g133640(.A0 (n_2842), .A1 (n_2235), .B0 (n_3252), .B1(n_2841), .Y (n_3253));
AOI21X1 g133651(.A0 (n_2996), .A1 (n_3250), .B0 (n_1814), .Y(n_3251));
AOI21X1 g134282(.A0 (n_2836), .A1 (n_2743), .B0 (n_3596), .Y(n_3249));
NAND3X1 g133586(.A (n_3247), .B (n_2423), .C (n_2556), .Y (n_3248));
NAND2X1 g133899(.A (n_32950), .B (P3_IR[15] ), .Y (n_3246));
INVX1 g134275(.A (n_3244), .Y (n_3245));
NAND2X1 g133152(.A (n_2990), .B (n_3242), .Y (n_3243));
XOR2X1 g133699(.A (n_1840), .B (n_3144), .Y (n_3451));
OR2X1 g133854(.A (n_3240), .B (n_3239), .Y (n_3241));
INVX1 g134043(.A (n_3072), .Y (n_3269));
NOR2X1 g134289(.A (n_3472), .B (n_3235), .Y (n_3826));
AOI21X1 g133302(.A0 (n_3104), .A1 (n_2297), .B0 (n_2933), .Y(n_3360));
NAND4X1 g133965(.A (n_2984), .B (n_2976), .C (P2_reg3[27] ), .D(P2_reg3[26] ), .Y (n_3404));
AND2X1 g134303(.A (n_2654), .B (n_3148), .Y (n_3234));
NAND2X1 g134319(.A (n_4523), .B (n_3032), .Y (n_3233));
NAND4X1 g133636(.A (n_2362), .B (n_1461), .C (n_2767), .D (n_3109),.Y (n_3232));
OAI21X1 g134336(.A0 (n_2076), .A1 (n_2985), .B0 (n_3231), .Y(n_6044));
NAND3X1 g133598(.A (n_1993), .B (n_2865), .C (n_2759), .Y (n_3230));
NAND2X1 g132557(.A (n_2895), .B (n_2894), .Y (n_9209));
NAND2X1 g134006(.A (n_2993), .B (n_2776), .Y (n_3228));
XOR2X1 g132560(.A (P1_reg3[22] ), .B (n_2751), .Y (n_3372));
AOI22X1 g133678(.A0 (n_1367), .A1 (n_3226), .B0 (P2_IR[25] ), .B1(n_33579), .Y (n_3227));
XOR2X1 g133390(.A (n_1822), .B (n_3007), .Y (n_3225));
NAND2X1 g133506(.A (n_2903), .B (n_33567), .Y (n_3224));
NAND3X1 g133539(.A (n_3222), .B (n_2419), .C (n_3221), .Y (n_3223));
NAND2X1 g133590(.A (n_3088), .B (n_1796), .Y (n_3220));
NAND2X1 g133138(.A (n_7706), .B (n_3217), .Y (n_3218));
NAND2X1 g134165(.A (n_7755), .B (n_7243), .Y (n_3215));
INVX1 g134173(.A (n_4426), .Y (n_3212));
MX2X1 g134398(.A (n_1969), .B (n_603), .S0 (n_2861), .Y (n_3210));
NAND2X1 g134443(.A (n_2807), .B (P1_reg2[1] ), .Y (n_3637));
NAND2X1 g134489(.A (n_3054), .B (n_13677), .Y (n_3663));
NAND2X1 g133562(.A (n_2559), .B (n_2892), .Y (n_3209));
MX2X1 g134085(.A (P3_reg3[10] ), .B (n_301), .S0 (n_2687), .Y(n_3295));
NAND2X1 g132779(.A (n_3178), .B (n_3314), .Y (n_3680));
INVX1 g134323(.A (n_3206), .Y (n_3207));
NAND2X1 g133671(.A (n_2947), .B (n_2942), .Y (n_8207));
MX2X1 g133707(.A (P3_reg3[13] ), .B (n_272), .S0 (n_2778), .Y(n_3262));
NOR2X1 g133510(.A (n_2837), .B (n_7245), .Y (n_3205));
AOI21X1 g134018(.A0 (n_3204), .A1 (n_3678), .B0 (n_3203), .Y(n_3393));
AND2X1 g133900(.A (n_2771), .B (n_3201), .Y (n_3202));
XOR2X1 g132587(.A (n_1210), .B (n_3199), .Y (n_3200));
INVX1 g133674(.A (n_3198), .Y (n_10612));
INVX1 g134143(.A (n_3289), .Y (n_3197));
NOR2X1 g133874(.A (n_2987), .B (n_3196), .Y (n_3305));
OAI21X1 g133063(.A0 (n_3195), .A1 (n_2016), .B0 (n_2301), .Y(n_3394));
OAI21X1 g133060(.A0 (n_3039), .A1 (n_2495), .B0 (n_3093), .Y(n_3194));
OAI21X1 g133847(.A0 (n_3193), .A1 (n_2566), .B0 (n_2960), .Y(n_3653));
INVX1 g134251(.A (n_3192), .Y (n_3444));
NAND3X1 g133595(.A (n_3313), .B (n_3189), .C (n_3188), .Y (n_3190));
NAND2X1 g133197(.A (n_2909), .B (n_3185), .Y (n_3186));
OAI21X1 g133250(.A0 (n_3158), .A1 (n_2481), .B0 (n_3182), .Y(n_3183));
MX2X1 g134057(.A (n_668), .B (P1_IR[11] ), .S0 (n_33672), .Y(n_3181));
NAND2X1 g133886(.A (n_13378), .B (n_7243), .Y (n_3180));
AND2X1 g133922(.A (n_874), .B (n_2995), .Y (n_3179));
NOR2X1 g132690(.A (n_3178), .B (n_3314), .Y (n_3679));
NOR2X1 g134537(.A (n_2807), .B (P1_reg2[1] ), .Y (n_3638));
NAND2X1 g134320(.A (n_4556), .B (n_3116), .Y (n_3177));
INVX1 g134210(.A (n_3176), .Y (n_3450));
NAND2X1 g134530(.A (n_3054), .B (n_13332), .Y (n_3745));
INVX1 g134091(.A (n_8055), .Y (n_3297));
NOR2X1 g134441(.A (n_2807), .B (P1_reg1[1] ), .Y (n_3559));
INVX1 g134261(.A (n_3174), .Y (n_6963));
NAND2X1 g134503(.A (n_3747), .B (n_3231), .Y (n_3173));
NOR2X1 g134512(.A (n_3054), .B (n_13332), .Y (n_3759));
AND2X1 g134189(.A (n_3170), .B (n_2878), .Y (n_3171));
NAND3X1 g133550(.A (n_3294), .B (n_3168), .C (n_2957), .Y (n_3169));
INVX1 g133564(.A (n_3454), .Y (n_3167));
NAND2X1 g133903(.A (n_10097), .B (n_7243), .Y (n_3166));
NOR2X1 g134134(.A (n_3162), .B (P3_reg1[3] ), .Y (n_4079));
NAND2X1 g133881(.A (n_13735), .B (n_7243), .Y (n_3161));
INVX1 g133401(.A (n_3191), .Y (n_3160));
OAI21X1 g133076(.A0 (n_3159), .A1 (n_2480), .B0 (n_3158), .Y(n_3456));
MX2X1 g134366(.A (n_1018), .B (P1_IR[12] ), .S0 (n_2786), .Y(n_3156));
INVX1 g134036(.A (n_3493), .Y (n_13381));
INVX1 g133984(.A (n_3152), .Y (n_3153));
OAI21X1 g133738(.A0 (n_2826), .A1 (n_998), .B0 (n_763), .Y (n_3151));
AOI21X1 g133305(.A0 (n_2886), .A1 (n_2797), .B0 (n_2848), .Y(n_3486));
MX2X1 g134056(.A (n_551), .B (n_1175), .S0 (n_3121), .Y (n_3150));
INVX1 g134354(.A (n_3147), .Y (n_3367));
OAI21X1 g133846(.A0 (n_3146), .A1 (n_2781), .B0 (n_3000), .Y(n_3419));
AOI21X1 g133645(.A0 (n_3144), .A1 (n_3140), .B0 (n_2695), .Y(n_3145));
AOI21X1 g134002(.A0 (n_3142), .A1 (n_3188), .B0 (n_3141), .Y(n_3143));
AOI21X1 g133627(.A0 (n_2514), .A1 (n_3140), .B0 (n_2963), .Y(n_3412));
OR2X1 g133993(.A (n_2961), .B (n_3139), .Y (n_3672));
NAND2X1 g134445(.A (n_2807), .B (P1_reg1[1] ), .Y (n_3560));
NAND2X1 g134061(.A (n_2928), .B (n_2986), .Y (n_9337));
INVX1 g133516(.A (n_3137), .Y (n_3138));
AOI21X1 g132902(.A0 (n_3095), .A1 (n_3242), .B0 (n_3136), .Y(n_3661));
NOR2X1 g133623(.A (n_2087), .B (n_2939), .Y (n_3263));
NAND2X1 g133502(.A (n_2784), .B (n_1313), .Y (n_3133));
INVX1 g134405(.A (n_3125), .Y (n_3129));
NAND3X1 g134229(.A (n_1576), .B (n_2672), .C (n_1577), .Y (n_3507));
AND2X1 g134317(.A (n_3126), .B (n_3125), .Y (n_3127));
INVX1 g133701(.A (n_3124), .Y (n_10822));
NAND2X2 g134215(.A (n_2628), .B (n_3121), .Y (n_3379));
NAND3X1 g134270(.A (n_2130), .B (n_3097), .C (n_2380), .Y (n_3120));
INVX1 g134479(.A (n_3472), .Y (n_3148));
MX2X1 g133675(.A (P2_reg3[21] ), .B (n_19), .S0 (n_2653), .Y(n_3198));
INVX1 g134211(.A (n_3201), .Y (n_3176));
NAND2X1 g134207(.A (n_2550), .B (n_2921), .Y (n_3119));
NAND2X1 g134205(.A (n_3117), .B (n_2860), .Y (n_3118));
NAND2X1 g134188(.A (n_2839), .B (n_2475), .Y (n_3115));
NAND2X1 g134217(.A (n_2762), .B (n_3005), .Y (n_3114));
OAI21X1 g133947(.A0 (n_2528), .A1 (n_2131), .B0 (n_2871), .Y(n_3301));
XOR2X1 g134117(.A (P1_reg3[24] ), .B (n_2618), .Y (n_3184));
INVX1 g134679(.A (n_3170), .Y (n_3334));
NAND2X1 g132601(.A (n_2804), .B (n_2874), .Y (n_7819));
NAND2X1 g132626(.A (n_3199), .B (n_2465), .Y (n_3292));
AOI22X1 g133058(.A0 (n_2042), .A1 (n_2732), .B0 (n_2907), .B1(n_1882), .Y (n_3468));
OR4X1 g133202(.A (n_2835), .B (addr_492), .C (addr_490), .D(addr_491), .Y (n_3112));
NAND2X1 g134276(.A (n_3310), .B (n_32453), .Y (n_3244));
NAND2X1 g134252(.A (n_2859), .B (n_2795), .Y (n_3192));
INVX1 g134071(.A (n_2911), .Y (n_3157));
NAND4X1 g134003(.A (n_2857), .B (n_3109), .C (n_269), .D (n_3108), .Y(n_3110));
INVX1 g133973(.A (n_3106), .Y (n_3107));
NAND2X1 g133565(.A (n_3069), .B (n_190), .Y (n_3454));
AOI21X1 g133285(.A0 (n_3104), .A1 (n_2296), .B0 (n_2592), .Y(n_3320));
INVX1 g134704(.A (n_3103), .Y (n_3713));
OAI21X1 g133871(.A0 (n_2643), .A1 (n_3252), .B0 (n_2879), .Y(n_3284));
NAND2X1 g132594(.A (n_2746), .B (n_2808), .Y (n_7575));
INVX1 g132596(.A (n_3100), .Y (n_3101));
NAND2X1 g134187(.A (n_2852), .B (n_606), .Y (n_3099));
NAND3X1 g134285(.A (n_2300), .B (n_2381), .C (n_3097), .Y (n_3098));
OR4X1 g133163(.A (n_2763), .B (addr_452), .C (addr_450), .D(addr_451), .Y (n_3096));
NAND3X1 g134243(.A (n_2714), .B (n_827), .C (n_2640), .Y (n_3308));
OAI21X1 g133628(.A0 (n_2847), .A1 (n_2467), .B0 (n_3017), .Y(n_3275));
AOI21X1 g133650(.A0 (n_3534), .A1 (n_3068), .B0 (n_3095), .Y(n_3738));
OR2X1 g133566(.A (n_3093), .B (n_2338), .Y (n_3094));
XOR2X1 g133383(.A (n_1303), .B (n_3104), .Y (n_3092));
INVX1 g133981(.A (n_3090), .Y (n_3091));
INVX1 g133987(.A (n_3088), .Y (n_3089));
AOI21X1 g134001(.A0 (n_3049), .A1 (n_3086), .B0 (n_3085), .Y(n_3087));
AND2X1 g133975(.A (n_2875), .B (n_1083), .Y (n_3084));
NAND2X1 g134226(.A (n_2740), .B (n_2484), .Y (n_3082));
MX2X1 g134126(.A (n_1624), .B (n_549), .S0 (n_2632), .Y (n_3081));
NOR2X1 g134174(.A (n_2780), .B (n_2462), .Y (n_4426));
INVX1 g134463(.A (n_3078), .Y (n_3079));
NOR2X1 g134550(.A (n_1825), .B (n_32238), .Y (n_3075));
NAND2X1 g134287(.A (n_3061), .B (n_3060), .Y (n_3074));
AOI21X1 g134324(.A0 (n_2683), .A1 (n_1766), .B0 (n_2858), .Y(n_3206));
OAI21X1 g133952(.A0 (n_2673), .A1 (n_2252), .B0 (n_2822), .Y(n_3542));
NAND2X1 g133546(.A (n_7724), .B (n_3217), .Y (n_3071));
AOI21X1 g134326(.A0 (n_2828), .A1 (n_1789), .B0 (n_2753), .Y(n_3271));
AND2X1 g133992(.A (n_2754), .B (n_969), .Y (n_3070));
NOR2X1 g133554(.A (n_3069), .B (n_190), .Y (n_3523));
AND2X1 g133203(.A (n_3242), .B (n_3068), .Y (n_3299));
MX2X1 g134348(.A (P3_IR[10] ), .B (n_34849), .S0 (n_2682), .Y(n_3067));
OAI21X1 g133348(.A0 (n_2787), .A1 (P2_reg3[27] ), .B0 (n_2788), .Y(n_10601));
NOR2X1 g133504(.A (n_3064), .B (n_1627), .Y (n_3065));
NAND3X1 g134152(.A (n_2626), .B (n_1229), .C (n_2633), .Y (n_3307));
NOR3X1 g134144(.A (n_3063), .B (n_2872), .C (n_32505), .Y (n_3289));
NAND3X1 g134140(.A (n_3061), .B (n_3060), .C (n_3613), .Y (n_3062));
NAND4X1 g134050(.A (n_2936), .B (n_2938), .C (n_2474), .D (n_2084),.Y (n_3059));
MX2X1 g134108(.A (n_586), .B (P2_reg3[20] ), .S0 (n_2668), .Y(n_10041));
OAI33X1 g133310(.A0 (n_2208), .A1 (n_2099), .A2 (n_2490), .B0(n_2854), .B1 (n_2152), .B2 (n_1826), .Y (n_3425));
NAND2X1 g134227(.A (n_3057), .B (n_2764), .Y (n_3058));
INVX1 g134546(.A (n_3055), .Y (n_3056));
NOR2X1 g134545(.A (n_3054), .B (n_13677), .Y (n_3899));
NAND4X1 g133997(.A (n_2821), .B (n_2518), .C (n_2085), .D (n_809), .Y(n_3052));
CLKBUFX1 g134541(.A (n_3240), .Y (n_6887));
AOI21X1 g133985(.A0 (n_2969), .A1 (n_3050), .B0 (n_3049), .Y(n_3152));
NAND2X1 g133838(.A (n_3009), .B (P3_reg3[14] ), .Y (n_3048));
OR4X1 g133141(.A (n_2831), .B (addr_433), .C (addr_431), .D(addr_432), .Y (n_3047));
NAND2X1 g133606(.A (n_7664), .B (n_34309), .Y (n_3046));
OAI22X1 g134119(.A0 (n_2689), .A1 (P1_reg3[20] ), .B0 (n_2688), .B1(n_134), .Y (n_7957));
NAND2X1 g134313(.A (n_34412), .B (n_1955), .Y (n_3255));
AOI21X1 g133996(.A0 (n_2306), .A1 (n_1828), .B0 (n_2863), .Y(n_3365));
MX2X1 g134399(.A (n_34199), .B (n_434), .S0 (n_3097), .Y (n_3044));
AOI21X1 g133517(.A0 (n_2635), .A1 (n_3022), .B0 (n_3043), .Y(n_3137));
MX2X1 g134127(.A (P3_IR[18] ), .B (n_943), .S0 (n_2705), .Y(n_3042));
NAND2X1 g132599(.A (n_2748), .B (n_2752), .Y (n_8164));
INVX1 g134024(.A (n_13389), .Y (n_9313));
NAND2X1 g133499(.A (n_2631), .B (n_3039), .Y (n_3327));
NAND2X1 g133856(.A (n_10578), .B (n_7243), .Y (n_3038));
INVX1 g134110(.A (n_3037), .Y (n_13375));
MX2X1 g134094(.A (n_1012), .B (P1_IR[13] ), .S0 (n_2805), .Y(n_3036));
OAI22X1 g134092(.A0 (n_2856), .A1 (P3_reg3[16] ), .B0 (n_2652), .B1(n_17), .Y (n_8055));
MX2X1 g134125(.A (n_1274), .B (n_120), .S0 (n_2615), .Y (n_3035));
NAND2X1 g132200(.A (n_10617), .B (n_1313), .Y (n_3034));
INVX1 g134493(.A (n_3162), .Y (n_3165));
MX2X1 g134037(.A (P3_reg3[18] ), .B (n_320), .S0 (n_2722), .Y(n_3493));
INVX1 g134075(.A (n_10103), .Y (n_13379));
NAND2X1 g133938(.A (n_800), .B (n_2994), .Y (n_3027));
NAND4X1 g134238(.A (n_2953), .B (n_2952), .C (n_2951), .D (n_2031),.Y (n_3026));
NOR2X1 g134532(.A (n_2760), .B (n_33676), .Y (n_3025));
INVX1 g133730(.A (n_3105), .Y (n_3024));
NAND2X1 g133714(.A (n_2816), .B (n_2840), .Y (n_8458));
NAND4X1 g134048(.A (n_3022), .B (n_2542), .C (n_2634), .D (n_3276),.Y (n_3023));
XOR2X1 g133402(.A (P2_reg3[19] ), .B (n_2669), .Y (n_3191));
MX2X1 g134096(.A (n_764), .B (P2_IR[13] ), .S0 (n_2829), .Y(n_3021));
AND2X1 g133991(.A (n_2827), .B (n_812), .Y (n_3020));
NAND2X1 g133404(.A (n_2738), .B (n_2749), .Y (n_8001));
NOR2X1 g133580(.A (n_3017), .B (n_2468), .Y (n_3018));
INVX1 g134031(.A (n_10114), .Y (n_3187));
INVX1 g134039(.A (n_10119), .Y (n_13386));
MX2X1 g134363(.A (n_117), .B (n_1218), .S0 (n_2736), .Y (n_3257));
MX2X1 g134355(.A (n_32473), .B (n_32475), .S0 (n_2621), .Y (n_3147));
NOR2X1 g133883(.A (n_3095), .B (n_2774), .Y (n_3012));
INVX1 g134262(.A (n_3239), .Y (n_3174));
AND2X1 g134228(.A (n_3162), .B (n_2720), .Y (n_3011));
OR2X1 g133837(.A (n_3009), .B (P3_reg3[14] ), .Y (n_3010));
NAND3X1 g133594(.A (n_3007), .B (n_3006), .C (n_3005), .Y (n_3008));
NAND2X1 g133575(.A (n_3003), .B (P1_reg3[28] ), .Y (n_3004));
AOI21X1 g134000(.A0 (n_3141), .A1 (n_3001), .B0 (n_2791), .Y(n_3002));
OAI21X1 g133845(.A0 (n_3000), .A1 (n_2515), .B0 (n_2999), .Y(n_3380));
INVX2 g134245(.A (n_3029), .Y (n_2998));
OAI21X1 g133343(.A0 (n_2769), .A1 (P1_reg3[23] ), .B0 (n_2770), .Y(n_13173));
OAI21X1 g133949(.A0 (n_2660), .A1 (n_2263), .B0 (n_2862), .Y(n_3410));
INVX1 g134416(.A (n_3203), .Y (n_3116));
INVX1 g134232(.A (n_2996), .Y (n_2997));
INVX1 g134332(.A (n_2994), .Y (n_2995));
NAND2X1 g134314(.A (n_2810), .B (n_2992), .Y (n_2993));
AOI21X1 g134041(.A0 (n_2450), .A1 (n_2219), .B0 (n_2591), .Y(n_2991));
INVX1 g133577(.A (n_3136), .Y (n_2990));
NAND3X1 g134175(.A (n_1813), .B (n_2502), .C (n_2989), .Y (n_3373));
OAI21X1 g133308(.A0 (n_2916), .A1 (n_1941), .B0 (n_2508), .Y(n_2988));
NOR3X1 g134331(.A (n_1950), .B (n_2438), .C (n_32321), .Y (n_2987));
OR2X1 g134284(.A (n_2983), .B (P2_reg3[16] ), .Y (n_2986));
INVX1 g134718(.A (n_2985), .Y (n_3747));
NOR2X1 g134192(.A (n_2757), .B (n_2983), .Y (n_2984));
MX2X1 g134357(.A (n_1799), .B (P2_IR[10] ), .S0 (n_2417), .Y(n_2982));
AOI21X1 g133988(.A0 (n_2494), .A1 (n_2037), .B0 (n_2666), .Y(n_3088));
MX2X1 g134680(.A (n_32485), .B (n_32486), .S0 (n_2464), .Y (n_3170));
MX2X1 g134111(.A (P3_reg3[15] ), .B (n_231), .S0 (n_2820), .Y(n_3037));
NAND2X2 g134247(.A (n_2944), .B (n_1763), .Y (n_3029));
AOI21X1 g134212(.A0 (n_865), .A1 (n_33111), .B0 (n_2701), .Y(n_3201));
NAND4X1 g132889(.A (n_2726), .B (n_2255), .C (n_2976), .D (n_1499),.Y (n_2977));
NAND2X1 g132924(.A (n_2597), .B (n_2715), .Y (n_7737));
INVX1 g134468(.A (n_34412), .Y (n_2974));
AOI21X1 g134004(.A0 (n_2443), .A1 (n_2303), .B0 (n_790), .Y (n_2972));
AOI21X1 g133982(.A0 (n_2257), .A1 (n_1793), .B0 (n_2699), .Y(n_3090));
NAND2X1 g133851(.A (n_7730), .B (n_3217), .Y (n_2971));
OAI21X1 g133950(.A0 (n_2853), .A1 (n_2716), .B0 (n_2761), .Y(n_3323));
AOI21X1 g133974(.A0 (n_2100), .A1 (n_2912), .B0 (n_2969), .Y(n_3106));
MX2X1 g134076(.A (P3_reg3[24] ), .B (n_188), .S0 (n_2432), .Y(n_10103));
NOR2X1 g134164(.A (n_2485), .B (n_2739), .Y (n_2967));
NOR2X1 g134168(.A (n_2476), .B (n_2838), .Y (n_2966));
OR2X1 g134186(.A (n_2964), .B (n_2284), .Y (n_2965));
OAI21X1 g133826(.A0 (n_2877), .A1 (n_2383), .B0 (n_2694), .Y(n_2963));
INVX1 g134372(.A (n_2962), .Y (n_3045));
NOR2X1 g134286(.A (n_2960), .B (n_2516), .Y (n_2961));
NAND2X1 g134307(.A (n_2958), .B (n_2957), .Y (n_2959));
NOR2X1 g134256(.A (n_2955), .B (n_2783), .Y (n_2956));
MX2X1 g134032(.A (P3_reg3[23] ), .B (n_343), .S0 (n_2519), .Y(n_10114));
AOI21X1 g133980(.A0 (n_2931), .A1 (n_2044), .B0 (n_2698), .Y(n_3272));
NAND3X1 g134177(.A (n_2953), .B (n_2952), .C (n_2951), .Y (n_2954));
NAND2X1 g134717(.A (n_2950), .B (P2_reg2[1] ), .Y (n_3350));
AND2X1 g134800(.A (n_3006), .B (n_2948), .Y (n_2949));
NAND2X1 g133857(.A (n_2941), .B (P1_reg3[21] ), .Y (n_2947));
NAND2X1 g134179(.A (n_284), .B (n_2944), .Y (n_2945));
OR2X1 g133918(.A (n_2941), .B (P1_reg3[21] ), .Y (n_2942));
NAND2X1 g133939(.A (n_2777), .B (n_2938), .Y (n_2939));
MX2X1 g133702(.A (P1_reg3[17] ), .B (n_202), .S0 (n_2675), .Y(n_3124));
NAND3X1 g133920(.A (n_2936), .B (n_2938), .C (n_2474), .Y (n_2937));
AOI21X1 g133972(.A0 (n_2348), .A1 (n_1924), .B0 (n_2731), .Y(n_3254));
MX2X1 g134396(.A (n_666), .B (n_1753), .S0 (n_2477), .Y (n_2934));
NAND2X1 g134012(.A (n_2593), .B (n_2932), .Y (n_2933));
MX2X1 g134040(.A (P3_reg3[20] ), .B (n_354), .S0 (n_2437), .Y(n_10119));
NAND3X1 g134005(.A (n_2585), .B (n_2311), .C (n_2931), .Y (n_3313));
OAI21X1 g133956(.A0 (n_2241), .A1 (n_2329), .B0 (n_2686), .Y(n_3316));
NAND2X1 g133908(.A (n_2232), .B (n_2685), .Y (n_3222));
NAND2X1 g134200(.A (n_13711), .B (n_7243), .Y (n_2929));
NAND2X1 g134184(.A (n_2983), .B (P2_reg3[16] ), .Y (n_2928));
MX2X1 g134400(.A (n_562), .B (n_1720), .S0 (n_2952), .Y (n_2927));
NAND4X1 g132884(.A (n_2713), .B (n_2408), .C (n_2870), .D (n_1681),.Y (n_2926));
OAI21X1 g133877(.A0 (n_2873), .A1 (n_2017), .B0 (n_2734), .Y(n_3247));
INVX1 g134403(.A (n_3362), .Y (n_3032));
NAND3X1 g134542(.A (n_2403), .B (n_1455), .C (n_2471), .Y (n_3240));
INVX2 g134464(.A (n_2921), .Y (n_3078));
XOR2X1 g133731(.A (P1_reg3[15] ), .B (n_2561), .Y (n_3105));
NAND2X1 g135943(.A (P2_IR[30] ), .B (n_2415), .Y (n_2920));
NAND2X1 g133603(.A (n_2917), .B (P1_reg3[27] ), .Y (n_2918));
XOR2X1 g133391(.A (n_2271), .B (n_2916), .Y (n_3178));
NOR2X1 g134176(.A (n_2889), .B (n_2386), .Y (n_2915));
INVX1 g134123(.A (n_2914), .Y (n_13370));
NAND2X1 g134547(.A (n_2785), .B (n_1934), .Y (n_3055));
NAND4X1 g134102(.A (n_2100), .B (n_3050), .C (n_2912), .D (n_3511),.Y (n_2913));
INVX1 g133727(.A (n_2909), .Y (n_2910));
XOR2X1 g133394(.A (n_1530), .B (n_2907), .Y (n_2908));
OAI21X1 g133719(.A0 (n_2710), .A1 (P2_reg3[15] ), .B0 (n_2711), .Y(n_8467));
NAND3X1 g133994(.A (n_2586), .B (n_1491), .C (n_2352), .Y (n_2905));
NAND3X1 g134263(.A (n_2396), .B (n_1156), .C (n_2512), .Y (n_3239));
AOI21X1 g134046(.A0 (n_2215), .A1 (n_2333), .B0 (n_2691), .Y(n_2904));
NOR2X1 g134705(.A (n_2950), .B (P2_reg2[1] ), .Y (n_3103));
MX2X1 g134059(.A (n_34524), .B (n_1211), .S0 (n_34543), .Y (n_2903));
MX2X1 g134045(.A (n_330), .B (P3_reg3[17] ), .S0 (n_2517), .Y(n_3072));
NOR2X1 g134623(.A (n_2899), .B (n_2270), .Y (n_2900));
MX2X1 g134365(.A (n_1968), .B (P1_IR[10] ), .S0 (n_2473), .Y(n_2898));
XOR2X1 g132597(.A (P2_reg3[14] ), .B (n_2530), .Y (n_3100));
NAND2X1 g134389(.A (n_2616), .B (n_2636), .Y (n_8185));
NAND3X1 g133989(.A (n_2676), .B (n_1459), .C (n_2260), .Y (n_2896));
NAND2X1 g132803(.A (n_2893), .B (P2_reg3[22] ), .Y (n_2895));
OR2X1 g132810(.A (n_2893), .B (P2_reg3[22] ), .Y (n_2894));
NOR2X1 g133925(.A (n_2891), .B (n_1669), .Y (n_2892));
NOR2X1 g134166(.A (n_2889), .B (n_2546), .Y (n_2890));
MX2X1 g133342(.A (n_238), .B (P2_reg3[23] ), .S0 (n_2506), .Y(n_10032));
XOR2X1 g133399(.A (n_1081), .B (n_2886), .Y (n_2887));
NAND2X1 g134725(.A (n_2950), .B (P2_reg1[1] ), .Y (n_3231));
OAI21X1 g133943(.A0 (n_2812), .A1 (n_2120), .B0 (n_2661), .Y(n_3294));
NAND3X1 g134511(.A (n_2881), .B (n_2883), .C (n_2882), .Y (n_2885));
AOI21X1 g134328(.A0 (n_2612), .A1 (n_1931), .B0 (n_2735), .Y(n_3354));
NAND4X1 g134571(.A (n_2000), .B (n_2883), .C (n_2882), .D (n_2881),.Y (n_2884));
INVX1 g134301(.A (n_2879), .Y (n_2880));
OAI21X1 g133954(.A0 (n_2162), .A1 (n_1701), .B0 (n_2526), .Y(n_3039));
OAI21X1 g133944(.A0 (n_2221), .A1 (n_1692), .B0 (n_2493), .Y(n_3093));
NAND2X1 g134219(.A (n_2513), .B (n_2877), .Y (n_3144));
NAND3X1 g134334(.A (n_2202), .B (n_2876), .C (n_33376), .Y (n_3226));
AND2X1 g134327(.A (n_605), .B (n_2609), .Y (n_2875));
INVX1 g134683(.A (n_7755), .Y (n_2975));
OR2X1 g132638(.A (n_2803), .B (P1_reg3[18] ), .Y (n_2874));
XOR2X1 g134081(.A (n_2121), .B (n_2873), .Y (n_3069));
INVX1 g134904(.A (n_2872), .Y (n_3054));
NOR2X1 g134288(.A (n_2132), .B (n_2529), .Y (n_2871));
INVX1 g134652(.A (n_8190), .Y (n_2979));
NAND4X1 g133968(.A (n_2525), .B (n_2870), .C (P1_reg3[27] ), .D(P1_reg3[26] ), .Y (n_3003));
OR2X1 g134296(.A (n_1310), .B (n_2687), .Y (n_3009));
INVX1 g134446(.A (n_33564), .Y (n_2869));
INVX1 g134638(.A (n_2629), .Y (n_3057));
NAND2X2 g134293(.A (n_34543), .B (n_2670), .Y (n_32951));
OR2X1 g134231(.A (n_2864), .B (n_2650), .Y (n_2865));
OAI21X1 g134337(.A0 (n_2307), .A1 (n_2310), .B0 (n_1829), .Y(n_2863));
NOR2X1 g134181(.A (n_2049), .B (n_2503), .Y (n_2862));
INVX1 g134751(.A (n_2860), .Y (n_2861));
NAND2X1 g134847(.A (n_1228), .B (n_2532), .Y (n_2859));
INVX1 g134588(.A (n_2684), .Y (n_2858));
NOR2X1 g134206(.A (n_1868), .B (n_2856), .Y (n_2857));
XOR2X1 g133395(.A (n_1415), .B (n_2854), .Y (n_2855));
NAND2X1 g133960(.A (n_2479), .B (n_2853), .Y (n_3007));
INVX1 g134470(.A (n_2944), .Y (n_2852));
AND2X1 g134462(.A (n_2850), .B (n_2849), .Y (n_2851));
OAI21X1 g134013(.A0 (n_2729), .A1 (n_2796), .B0 (n_2847), .Y(n_2848));
INVX1 g134596(.A (n_2671), .Y (n_3061));
NOR2X1 g133578(.A (n_2773), .B (n_2772), .Y (n_3136));
AOI21X1 g134007(.A0 (n_2845), .A1 (n_2844), .B0 (n_2228), .Y(n_2846));
OAI33X1 g133309(.A0 (n_1927), .A1 (n_1400), .A2 (n_2083), .B0(n_2637), .B1 (n_1355), .B2 (n_1383), .Y (n_3199));
XOR2X1 g133728(.A (P2_reg3[13] ), .B (n_8212), .Y (n_2909));
NAND2X1 g133806(.A (n_7546), .B (n_3217), .Y (n_2843));
OR2X1 g134193(.A (n_2932), .B (n_2841), .Y (n_2842));
OAI21X1 g133953(.A0 (n_2004), .A1 (n_1823), .B0 (n_2436), .Y(n_3159));
OAI21X1 g133948(.A0 (n_2351), .A1 (n_1834), .B0 (n_2501), .Y(n_3195));
INVX1 g134600(.A (n_2648), .Y (n_3117));
OR2X1 g133931(.A (n_2815), .B (P2_reg3[17] ), .Y (n_2840));
INVX1 g134592(.A (n_2838), .Y (n_2839));
OR2X1 g134700(.A (n_2883), .B (n_2742), .Y (n_2836));
NAND4X1 g133966(.A (n_557), .B (n_2445), .C (n_50), .D (n_615), .Y(n_2835));
NAND3X1 g134333(.A (n_2136), .B (n_2834), .C (n_2825), .Y (n_2994));
NOR2X1 g133823(.A (n_2379), .B (n_33350), .Y (n_2833));
INVX1 g134375(.A (n_2832), .Y (n_10097));
NAND4X1 g133961(.A (n_588), .B (n_2412), .C (n_649), .D (n_638), .Y(n_2831));
INVX1 g134456(.A (n_2829), .Y (n_2830));
NAND2X1 g134519(.A (n_2581), .B (n_2828), .Y (n_3142));
NOR2X1 g134526(.A (n_2081), .B (n_2681), .Y (n_32453));
AND2X1 g134325(.A (n_472), .B (n_2706), .Y (n_2827));
MX2X1 g134373(.A (n_1858), .B (n_485), .S0 (n_2305), .Y (n_2962));
AOI21X1 g134566(.A0 (n_2330), .A1 (n_2133), .B0 (n_2712), .Y(n_3193));
OAI21X1 g133955(.A0 (n_2422), .A1 (n_2336), .B0 (n_2571), .Y(n_3158));
MX2X1 g134347(.A (n_618), .B (n_939), .S0 (n_2825), .Y (n_2826));
INVX1 g135261(.A (n_2950), .Y (n_2824));
OAI21X1 g133945(.A0 (n_1683), .A1 (n_1425), .B0 (n_2520), .Y(n_3064));
NAND2X1 g133805(.A (n_8193), .B (n_3185), .Y (n_2823));
NOR2X1 g134234(.A (n_2029), .B (n_2441), .Y (n_2822));
NOR2X1 g134190(.A (n_2820), .B (n_1320), .Y (n_2821));
MX2X1 g134356(.A (n_35865), .B (n_35867), .S0 (n_33376), .Y (n_2819));
INVX1 g134391(.A (n_2817), .Y (n_13378));
NAND2X1 g133906(.A (n_2815), .B (P2_reg3[17] ), .Y (n_2816));
INVX1 g134394(.A (n_2814), .Y (n_13735));
XOR2X1 g134099(.A (n_1922), .B (n_2812), .Y (n_2813));
INVX1 g134513(.A (n_2810), .Y (n_2811));
NOR2X1 g134719(.A (n_2950), .B (P2_reg1[1] ), .Y (n_2985));
OR2X1 g132645(.A (n_2745), .B (P1_reg3[14] ), .Y (n_2808));
INVX1 g134551(.A (n_2805), .Y (n_2806));
NAND2X1 g132630(.A (n_2803), .B (P1_reg3[18] ), .Y (n_2804));
NAND2X1 g134407(.A (n_2771), .B (P3_reg1[1] ), .Y (n_3125));
AND2X1 g134783(.A (n_2801), .B (n_2800), .Y (n_2802));
MX2X1 g134124(.A (P3_reg3[9] ), .B (n_1031), .S0 (n_2692), .Y(n_2914));
NAND2X1 g134450(.A (n_2540), .B (n_2798), .Y (n_2799));
NOR2X1 g134812(.A (n_2366), .B (n_2796), .Y (n_2797));
AOI22X1 g134667(.A0 (n_1011), .A1 (n_2531), .B0 (n_1227), .B1(n_33566), .Y (n_2795));
NAND3X1 g134255(.A (n_2793), .B (n_2792), .C (n_2791), .Y (n_2794));
NAND3X1 g134521(.A (n_2800), .B (n_2789), .C (n_1903), .Y (n_2790));
NAND2X1 g133599(.A (n_2787), .B (P2_reg3[27] ), .Y (n_2788));
INVX1 g134755(.A (n_2785), .Y (n_2786));
NAND2X1 g136256(.A (n_286), .B (n_32517), .Y (n_7549));
INVX2 g134465(.A (n_2783), .Y (n_2921));
INVX1 g134438(.A (n_2980), .Y (n_2782));
NOR2X1 g134823(.A (n_2541), .B (n_2781), .Y (n_3420));
OR2X1 g134424(.A (n_2943), .B (n_2779), .Y (n_2780));
INVX1 g134202(.A (n_2777), .Y (n_2778));
NAND2X1 g134619(.A (n_2533), .B (n_2776), .Y (n_3792));
NAND2X1 g134499(.A (n_2579), .B (n_2775), .Y (n_3893));
INVX1 g134304(.A (n_3068), .Y (n_2774));
NAND2X1 g133535(.A (n_2773), .B (n_2772), .Y (n_3242));
AND2X1 g134495(.A (n_2402), .B (n_2511), .Y (n_3162));
NOR2X1 g134417(.A (n_2771), .B (n_13337), .Y (n_3203));
NAND2X1 g133547(.A (n_2769), .B (P1_reg3[23] ), .Y (n_2770));
XOR2X1 g134098(.A (n_1570), .B (n_2584), .Y (n_2768));
NAND2X1 g134073(.A (n_2583), .B (n_2488), .Y (n_2911));
CLKBUFX1 g134377(.A (n_34587), .Y (n_10578));
NAND2X1 g134474(.A (n_2449), .B (n_3441), .Y (n_2766));
INVX1 g134741(.A (n_2764), .Y (n_32238));
NAND4X1 g133963(.A (n_466), .B (n_2551), .C (n_52), .D (n_563), .Y(n_2763));
INVX1 g134555(.A (n_2761), .Y (n_2762));
NAND2X1 g133723(.A (n_2545), .B (n_2575), .Y (n_7706));
INVX1 g134752(.A (n_2860), .Y (n_2760));
AOI21X1 g134657(.A0 (n_2368), .A1 (n_2218), .B0 (n_2149), .Y(n_2759));
OR2X1 g134420(.A (n_2548), .B (n_2757), .Y (n_2758));
NAND2X1 g134418(.A (n_2771), .B (n_13337), .Y (n_3678));
INVX1 g134742(.A (n_2764), .Y (n_2755));
AOI21X1 g134562(.A0 (n_2253), .A1 (n_2440), .B0 (n_2509), .Y(n_3146));
NOR2X1 g134404(.A (n_2771), .B (P3_reg1[1] ), .Y (n_3362));
AND2X1 g134329(.A (n_443), .B (n_2587), .Y (n_2754));
INVX1 g134603(.A (n_2704), .Y (n_2753));
OR2X1 g132639(.A (n_2747), .B (P2_reg3[18] ), .Y (n_2752));
NAND3X1 g134482(.A (n_2355), .B (n_1095), .C (n_2277), .Y (n_3472));
AND2X1 g133240(.A (n_2410), .B (n_2489), .Y (n_2751));
MX2X1 g134027(.A (n_56), .B (P3_reg3[19] ), .S0 (n_2378), .Y(n_13389));
AOI21X1 g134612(.A0 (n_2602), .A1 (n_2101), .B0 (n_2346), .Y(n_4135));
AOI21X1 g134602(.A0 (n_2662), .A1 (n_1996), .B0 (n_2564), .Y(n_2999));
NAND2X1 g134233(.A (n_2565), .B (n_2035), .Y (n_2996));
OAI21X1 g133946(.A0 (n_2126), .A1 (n_2204), .B0 (n_2534), .Y(n_3017));
OR2X1 g133509(.A (n_2737), .B (P1_reg3[19] ), .Y (n_2749));
NAND2X1 g132631(.A (n_2747), .B (P2_reg3[18] ), .Y (n_2748));
NAND2X1 g132644(.A (n_2745), .B (P1_reg3[14] ), .Y (n_2746));
NAND2X1 g134701(.A (n_2883), .B (n_2742), .Y (n_2743));
NOR2X1 g134432(.A (n_33924), .B (n_1801), .Y (n_3121));
INVX1 g134576(.A (n_2739), .Y (n_2740));
NAND2X1 g133507(.A (n_2737), .B (P1_reg3[19] ), .Y (n_2738));
NAND2X1 g134818(.A (n_32367), .B (n_1724), .Y (n_2736));
INVX1 g134669(.A (n_2573), .Y (n_2735));
AOI21X1 g134618(.A0 (n_2430), .A1 (n_2200), .B0 (n_2557), .Y(n_2734));
NAND3X1 g134625(.A (n_2537), .B (n_3538), .C (n_4280), .Y (n_2733));
AOI22X1 g134656(.A0 (n_1798), .A1 (n_1907), .B0 (n_2072), .B1(n_2071), .Y (n_3942));
AOI22X1 g134342(.A0 (n_2171), .A1 (n_1977), .B0 (n_2041), .B1(n_2169), .Y (n_2732));
NAND2X1 g134338(.A (n_1925), .B (n_2238), .Y (n_2731));
NAND2X1 g133079(.A (n_10880), .B (n_3217), .Y (n_2730));
OAI21X1 g133942(.A0 (n_2538), .A1 (n_2366), .B0 (n_2729), .Y(n_3043));
OR2X1 g134216(.A (n_2727), .B (n_2658), .Y (n_2728));
NAND2X1 g136209(.A (n_2718), .B (n_32509), .Y (n_7217));
INVX1 g133156(.A (n_2747), .Y (n_2726));
INVX1 g134497(.A (n_2724), .Y (n_2725));
INVX1 g134753(.A (n_2723), .Y (n_2860));
NAND4X1 g134659(.A (n_2374), .B (n_1311), .C (n_2721), .D (n_1691),.Y (n_2722));
INVX2 g134905(.A (n_2720), .Y (n_2872));
OR2X1 g134548(.A (n_2309), .B (n_733), .Y (n_2719));
OAI22X1 g134653(.A0 (n_1719), .A1 (n_1976), .B0 (n_2667), .B1(n_125), .Y (n_8190));
OR2X1 g136206(.A (n_2718), .B (n_32505), .Y (n_7216));
INVX1 g134996(.A (n_2716), .Y (n_3006));
OR2X1 g133165(.A (n_2596), .B (P1_reg3[10] ), .Y (n_2715));
OR2X1 g134883(.A (n_914), .B (n_2639), .Y (n_2714));
INVX1 g133123(.A (n_2803), .Y (n_2713));
NAND2X1 g134568(.A (n_2265), .B (n_1548), .Y (n_2958));
AOI21X1 g134622(.A0 (n_2712), .A1 (n_2115), .B0 (n_2603), .Y(n_2964));
NAND2X1 g133835(.A (n_2710), .B (P2_reg3[15] ), .Y (n_2711));
OAI21X1 g133951(.A0 (n_2455), .A1 (n_1885), .B0 (n_2222), .Y(n_3104));
OR2X1 g134792(.A (n_2388), .B (n_1076), .Y (n_2708));
INVX1 g134410(.A (n_2706), .Y (n_2707));
NAND3X1 g134442(.A (n_2082), .B (n_32368), .C (n_2194), .Y (n_2705));
AOI21X1 g134604(.A0 (n_2828), .A1 (n_2268), .B0 (n_2356), .Y(n_2704));
OAI22X1 g134668(.A0 (n_967), .A1 (n_33111), .B0 (n_34321), .B1(n_1724), .Y (n_2701));
NAND2X1 g134457(.A (n_2589), .B (n_33375), .Y (n_2829));
NAND2X1 g134346(.A (n_1769), .B (n_2258), .Y (n_2699));
OAI21X1 g134343(.A0 (n_2145), .A1 (n_1510), .B0 (n_1707), .Y(n_2698));
INVX1 g134634(.A (n_2694), .Y (n_2695));
AND2X1 g134471(.A (n_33237), .B (n_2033), .Y (n_2944));
INVX1 g134054(.A (n_2693), .Y (n_2784));
NOR2X1 g134203(.A (n_1173), .B (n_2692), .Y (n_2777));
NAND2X1 g134297(.A (n_2347), .B (n_2244), .Y (n_3139));
NOR2X1 g134299(.A (n_2690), .B (n_2458), .Y (n_2691));
INVX1 g134448(.A (n_2688), .Y (n_2689));
INVX1 g134453(.A (n_2687), .Y (n_2767));
NOR2X1 g134220(.A (n_2680), .B (n_11097), .Y (n_3095));
AOI22X1 g134640(.A0 (n_2205), .A1 (n_2124), .B0 (n_2079), .B1(n_2078), .Y (n_3697));
NOR2X1 g134248(.A (n_2156), .B (n_2242), .Y (n_2686));
NAND3X1 g134574(.A (n_35427), .B (n_34853), .C (n_2209), .Y (n_2889));
OAI21X1 g134583(.A0 (n_2500), .A1 (n_1881), .B0 (n_2170), .Y(n_2969));
AOI21X1 g134582(.A0 (n_2499), .A1 (n_2231), .B0 (n_2507), .Y(n_2685));
AOI21X1 g134589(.A0 (n_2683), .A1 (n_2364), .B0 (n_2220), .Y(n_2684));
INVX1 g134745(.A (n_2681), .Y (n_2682));
NAND2X1 g134305(.A (n_2680), .B (n_11097), .Y (n_3068));
NAND2X1 g134877(.A (n_3386), .B (n_2679), .Y (n_2899));
XOR2X1 g134078(.A (n_2067), .B (n_1841), .Y (n_2678));
INVX1 g134198(.A (n_2675), .Y (n_2676));
NAND2X1 g134214(.A (n_2283), .B (n_1373), .Y (n_2891));
AOI21X1 g134556(.A0 (n_2160), .A1 (n_2582), .B0 (n_2673), .Y(n_2761));
NAND2X1 g134888(.A (n_2245), .B (n_1609), .Y (n_2672));
NAND3X1 g134597(.A (n_1582), .B (n_2003), .C (n_2670), .Y (n_2671));
NOR2X1 g133915(.A (n_2394), .B (n_2196), .Y (n_2669));
NAND3X1 g134501(.A (n_2667), .B (n_2547), .C (n_1500), .Y (n_2668));
OAI21X1 g134339(.A0 (n_2095), .A1 (n_2578), .B0 (n_2038), .Y(n_2666));
AOI21X1 g134573(.A0 (n_1553), .A1 (n_1997), .B0 (n_2212), .Y(n_2665));
OR2X1 g134724(.A (n_2663), .B (n_1803), .Y (n_2664));
AOI21X1 g134611(.A0 (n_2426), .A1 (n_2182), .B0 (n_2662), .Y(n_4293));
NAND3X1 g134593(.A (n_1643), .B (n_2061), .C (n_2600), .Y (n_2838));
AOI21X1 g134567(.A0 (n_2075), .A1 (n_1502), .B0 (n_2611), .Y(n_3182));
AOI21X1 g134557(.A0 (n_1991), .A1 (n_2527), .B0 (n_2660), .Y(n_2661));
OR2X1 g134737(.A (n_2658), .B (n_2657), .Y (n_2659));
INVX1 g134730(.A (n_2654), .Y (n_2807));
NAND2X1 g134114(.A (n_2214), .B (n_2276), .Y (n_7664));
OR2X1 g134322(.A (n_2353), .B (n_2577), .Y (n_2653));
INVX1 g134543(.A (n_2856), .Y (n_2652));
NOR2X1 g134829(.A (n_2650), .B (n_2649), .Y (n_2651));
OR2X1 g134330(.A (n_2261), .B (n_2562), .Y (n_2941));
NAND2X2 g134466(.A (n_2233), .B (n_2472), .Y (n_2783));
NAND3X1 g134601(.A (n_33680), .B (n_2400), .C (n_33673), .Y (n_2648));
NAND2X1 g134854(.A (n_2281), .B (n_3538), .Y (n_2645));
NOR2X1 g134534(.A (n_2793), .B (n_3001), .Y (n_2644));
NAND2X1 g134533(.A (n_2642), .B (n_2236), .Y (n_2643));
NAND2X1 g134848(.A (n_4282), .B (n_3353), .Y (n_2641));
NAND2X1 g134760(.A (n_1016), .B (n_2639), .Y (n_2640));
NAND4X1 g133959(.A (n_1980), .B (n_1451), .C (n_2572), .D (n_954), .Y(n_2917));
XOR2X1 g133392(.A (n_1312), .B (n_2637), .Y (n_2638));
NAND2X1 g134514(.A (n_2372), .B (n_2109), .Y (n_2810));
OR2X1 g134435(.A (n_2620), .B (P2_reg3[12] ), .Y (n_2636));
AND2X1 g134774(.A (n_2542), .B (n_2634), .Y (n_2635));
NAND2X1 g134816(.A (n_1264), .B (n_2625), .Y (n_2633));
NAND3X1 g134506(.A (n_2331), .B (n_35278), .C (n_2064), .Y (n_2632));
NAND2X1 g134505(.A (n_2390), .B (n_835), .Y (n_2631));
NAND3X1 g134639(.A (n_1421), .B (n_2334), .C (n_2628), .Y (n_2629));
OR2X1 g134799(.A (n_2295), .B (n_1370), .Y (n_2627));
OR2X1 g134822(.A (n_1254), .B (n_2625), .Y (n_2626));
NAND3X1 g134496(.A (n_2623), .B (n_2622), .C (n_4037), .Y (n_2624));
OR2X1 g133176(.A (n_2256), .B (n_2605), .Y (n_2893));
NAND2X1 g134821(.A (n_2320), .B (P1_IR[31] ), .Y (n_2621));
OR2X1 g134467(.A (n_2620), .B (n_1215), .Y (n_2983));
INVX2 g134787(.A (n_33110), .Y (n_3097));
NOR2X1 g134423(.A (n_2227), .B (n_2524), .Y (n_2618));
NAND2X1 g134121(.A (n_2325), .B (n_2318), .Y (n_7724));
NAND2X1 g134444(.A (n_2365), .B (n_2349), .Y (n_3085));
NAND2X2 g134439(.A (n_1396), .B (n_33431), .Y (n_2980));
NOR2X1 g134756(.A (n_1987), .B (n_35160), .Y (n_2785));
NAND2X1 g134425(.A (n_2620), .B (P2_reg3[12] ), .Y (n_2616));
NAND2X1 g136303(.A (n_565), .B (n_32509), .Y (n_7550));
NAND3X1 g134485(.A (n_2234), .B (n_32482), .C (n_2048), .Y (n_2615));
INVX2 g134743(.A (n_33924), .Y (n_2764));
AND2X1 g134870(.A (n_2792), .B (n_3001), .Y (n_3800));
NAND2X1 g134553(.A (n_2269), .B (n_2612), .Y (n_3141));
OAI21X1 g134302(.A0 (n_2611), .A1 (n_1849), .B0 (n_2290), .Y(n_2879));
INVX1 g134408(.A (n_2609), .Y (n_2610));
NAND2X1 g133059(.A (n_10594), .B (n_3185), .Y (n_2608));
NAND2X1 g134500(.A (n_2254), .B (n_2683), .Y (n_3049));
MX2X1 g134376(.A (n_2), .B (P3_reg3[11] ), .S0 (n_2469), .Y(n_2832));
INVX1 g134598(.A (n_2606), .Y (n_2607));
NAND2X1 g134684(.A (n_2279), .B (n_2267), .Y (n_7755));
MX2X1 g132926(.A (n_334), .B (P2_reg3[10] ), .S0 (n_2605), .Y(n_10617));
MX2X1 g134392(.A (P3_reg3[12] ), .B (n_1032), .S0 (n_2554), .Y(n_2817));
INVX1 g134900(.A (n_2943), .Y (n_2878));
NOR2X1 g134569(.A (n_1492), .B (n_2340), .Y (n_8213));
AOI21X1 g134620(.A0 (n_2603), .A1 (n_2116), .B0 (n_2602), .Y(n_2960));
INVX1 g134065(.A (n_2601), .Y (n_2837));
NAND2X1 g134552(.A (n_2600), .B (n_2825), .Y (n_2805));
NOR2X1 g134507(.A (n_2448), .B (n_2598), .Y (n_2599));
NAND2X1 g133207(.A (n_2596), .B (P1_reg3[10] ), .Y (n_2597));
NOR2X1 g134475(.A (n_2539), .B (n_2594), .Y (n_2595));
NAND2X1 g134274(.A (n_2592), .B (n_2342), .Y (n_2593));
NOR2X1 g134309(.A (n_2590), .B (n_2406), .Y (n_2591));
MX2X1 g134395(.A (P3_reg3[6] ), .B (n_1027), .S0 (n_2549), .Y(n_2814));
NAND3X1 g134577(.A (n_35271), .B (n_1439), .C (n_2589), .Y (n_2739));
INVX1 g134412(.A (n_2587), .Y (n_2588));
INVX1 g134280(.A (n_2815), .Y (n_2586));
NAND3X1 g134218(.A (n_2584), .B (n_1561), .C (n_1526), .Y (n_2585));
NOR2X1 g134570(.A (n_1460), .B (n_2199), .Y (n_7761));
NAND2X1 g134387(.A (n_2062), .B (n_2176), .Y (n_7730));
NAND2X1 g134230(.A (n_2523), .B (P1_reg3[16] ), .Y (n_2583));
NAND2X1 g134997(.A (n_2582), .B (n_2098), .Y (n_2716));
NAND2X1 g134882(.A (n_2045), .B (n_1957), .Y (n_2581));
AOI22X1 g134665(.A0 (n_2111), .A1 (n_2332), .B0 (n_2011), .B1(n_1854), .Y (n_2580));
NAND2X1 g134866(.A (n_2010), .B (n_2578), .Y (n_2579));
AND2X1 g134795(.A (n_2642), .B (n_2341), .Y (n_3725));
OR2X1 g134281(.A (n_2165), .B (n_2577), .Y (n_2815));
OR2X1 g133841(.A (n_2544), .B (P1_reg3[13] ), .Y (n_2575));
INVX1 g135062(.A (n_2574), .Y (n_2800));
AOI22X1 g134670(.A0 (n_2404), .A1 (n_1942), .B0 (n_2612), .B1(n_1932), .Y (n_2573));
NAND3X1 g133897(.A (n_1451), .B (n_2486), .C (n_2572), .Y (n_2737));
NOR2X1 g134204(.A (n_1398), .B (n_2013), .Y (n_2571));
NOR2X1 g134483(.A (n_2569), .B (n_2026), .Y (n_2570));
OR2X1 g134820(.A (n_2399), .B (n_2566), .Y (n_2567));
AOI21X1 g134595(.A0 (n_2564), .A1 (n_1945), .B0 (n_1710), .Y(n_2565));
INVX1 g134066(.A (n_2563), .Y (n_2601));
OR2X1 g134199(.A (n_2021), .B (n_2562), .Y (n_2675));
NOR2X1 g134169(.A (n_1992), .B (n_1898), .Y (n_2561));
NAND3X1 g134180(.A (n_2559), .B (n_1670), .C (n_2558), .Y (n_2560));
AOI21X1 g134635(.A0 (n_2557), .A1 (n_2556), .B0 (n_2424), .Y(n_2694));
OR2X1 g134544(.A (n_2554), .B (n_1893), .Y (n_2856));
INVX1 g134508(.A (n_2551), .Y (n_2552));
NOR2X1 g134430(.A (n_2955), .B (n_1728), .Y (n_2550));
OR2X1 g134454(.A (n_2373), .B (n_2549), .Y (n_2687));
NAND2X1 g134838(.A (n_2667), .B (n_2547), .Y (n_2548));
NAND2X1 g134836(.A (n_2385), .B (n_2210), .Y (n_2546));
NAND2X1 g133830(.A (n_2544), .B (P1_reg3[13] ), .Y (n_2545));
XOR2X1 g134095(.A (n_1738), .B (n_3324), .Y (n_2543));
INVX1 g135033(.A (n_3005), .Y (n_2541));
INVX1 g134880(.A (n_2539), .Y (n_2540));
NAND2X1 g133967(.A (n_2134), .B (n_2538), .Y (n_2886));
INVX1 g135147(.A (n_2537), .Y (n_3943));
INVX1 g134878(.A (n_2535), .Y (n_2536));
NAND2X1 g134697(.A (n_2106), .B (n_2193), .Y (n_13711));
NOR2X1 g134221(.A (n_1910), .B (n_2127), .Y (n_2534));
NAND2X1 g134773(.A (n_2110), .B (n_2992), .Y (n_2533));
INVX1 g135028(.A (n_2531), .Y (n_2532));
NOR2X1 g133086(.A (n_2605), .B (n_1326), .Y (n_2530));
AOI21X1 g134626(.A0 (n_2528), .A1 (n_2229), .B0 (n_2527), .Y(n_2529));
OR2X1 g133157(.A (n_1874), .B (n_2605), .Y (n_2747));
NOR2X1 g134283(.A (n_1702), .B (n_2163), .Y (n_2526));
NOR2X1 g134254(.A (n_2524), .B (n_2523), .Y (n_2525));
NAND4X1 g133958(.A (n_2197), .B (n_2392), .C (n_1490), .D (n_711), .Y(n_2787));
NOR2X1 g134244(.A (n_1426), .B (n_2107), .Y (n_2520));
NAND4X1 g134671(.A (n_2377), .B (n_2376), .C (n_2375), .D (n_2518),.Y (n_2519));
NAND4X1 g134672(.A (n_2090), .B (n_1092), .C (n_2721), .D (n_2086),.Y (n_2517));
INVX1 g134721(.A (n_3063), .Y (n_2771));
NOR2X1 g134777(.A (n_2516), .B (n_2566), .Y (n_3951));
NOR2X1 g134793(.A (n_2515), .B (n_2781), .Y (n_2850));
INVX1 g134855(.A (n_2513), .Y (n_2514));
OR2X1 g134865(.A (n_893), .B (n_32375), .Y (n_2512));
AOI21X1 g134890(.A0 (n_34539), .A1 (n_33566), .B0 (n_2030), .Y(n_2511));
MX2X1 g134901(.A (n_1464), .B (n_371), .S0 (n_1727), .Y (n_2943));
NOR2X1 g134449(.A (n_2068), .B (n_2226), .Y (n_2688));
AOI21X1 g134599(.A0 (n_2509), .A1 (n_2312), .B0 (n_2427), .Y(n_2606));
INVX1 g135212(.A (n_2507), .Y (n_2508));
MX2X1 g134906(.A (n_32956), .B (n_32954), .S0 (n_1725), .Y (n_2720));
NAND2X1 g133124(.A (n_2409), .B (n_2489), .Y (n_2803));
NAND4X1 g133957(.A (n_1837), .B (n_2393), .C (n_1484), .D (n_1431),.Y (n_2506));
OR2X1 g135966(.A (n_2504), .B (n_34946), .Y (n_2505));
AOI21X1 g134575(.A0 (n_2660), .A1 (n_2190), .B0 (n_2264), .Y(n_2503));
NAND2X1 g134892(.A (n_2036), .B (n_1944), .Y (n_2502));
NOR2X1 g134277(.A (n_1809), .B (n_1999), .Y (n_2501));
OAI21X1 g133983(.A0 (n_1841), .A1 (n_1807), .B0 (n_2500), .Y(n_2907));
AOI21X1 g133978(.A0 (n_2478), .A1 (n_2230), .B0 (n_2499), .Y(n_2916));
OAI21X1 g135513(.A0 (P1_reg1[0] ), .A1 (n_7747), .B0 (n_2497), .Y(n_2498));
NOR2X1 g134484(.A (n_2389), .B (n_2495), .Y (n_2496));
AND2X1 g134498(.A (n_2073), .B (n_2494), .Y (n_2724));
NOR2X1 g134253(.A (n_1664), .B (n_1990), .Y (n_2493));
NAND2X2 g134746(.A (n_32369), .B (n_1449), .Y (n_2681));
AND2X1 g134759(.A (n_3283), .B (n_2642), .Y (n_2491));
AOI21X1 g134609(.A0 (n_2461), .A1 (n_2098), .B0 (n_2159), .Y(n_2490));
NAND2X1 g133087(.A (n_2489), .B (n_2192), .Y (n_2745));
CLKBUFX1 gbuf_d_701(.A(n_2189), .Y(d_out_701));
CLKBUFX1 gbuf_qn_701(.A(qn_in_701), .Y(P1_n_449));
OR2X1 g134201(.A (n_2523), .B (P1_reg3[16] ), .Y (n_2488));
NAND4X1 g133964(.A (n_1892), .B (n_2486), .C (n_1522), .D (n_1979),.Y (n_2769));
NAND2X1 g134831(.A (n_2484), .B (n_1411), .Y (n_2485));
OAI21X1 g134413(.A0 (n_1712), .A1 (n_567), .B0 (n_126), .Y (n_2587));
AOI21X1 g134560(.A0 (n_1417), .A1 (n_1494), .B0 (n_2483), .Y(n_3912));
NOR2X1 g134761(.A (n_2481), .B (n_2480), .Y (n_2482));
NAND2X1 g134185(.A (n_3324), .B (n_2948), .Y (n_2479));
NAND2X1 g134411(.A (n_2123), .B (n_147), .Y (n_2706));
XOR2X1 g134077(.A (n_1852), .B (n_2478), .Y (n_2773));
INVX1 g134833(.A (n_3060), .Y (n_2477));
NAND3X1 g134754(.A (n_32449), .B (n_32156), .C (n_647), .Y (n_2723));
NAND2X1 g134765(.A (n_2475), .B (n_1857), .Y (n_2476));
INVX1 g134517(.A (n_2692), .Y (n_2474));
INVX1 g134804(.A (n_2472), .Y (n_2473));
OR2X1 g135076(.A (n_1986), .B (n_33261), .Y (n_2471));
NAND2X1 g134436(.A (n_1617), .B (n_2469), .Y (n_2820));
OAI21X1 g134409(.A0 (n_1791), .A1 (n_417), .B0 (n_194), .Y (n_2609));
OR2X1 g134806(.A (n_2468), .B (n_2467), .Y (n_3422));
AND2X1 g134796(.A (n_2465), .B (n_2623), .Y (n_2466));
NAND2X1 g134980(.A (n_33358), .B (n_609), .Y (n_2464));
INVX1 g134731(.A (n_2462), .Y (n_2654));
AOI21X1 g134630(.A0 (n_2323), .A1 (n_2114), .B0 (n_2461), .Y(n_2853));
INVX1 g135273(.A (n_2460), .Y (n_2674));
OR2X1 g134775(.A (n_2458), .B (n_2457), .Y (n_2459));
XOR2X1 g134082(.A (n_1088), .B (n_2455), .Y (n_2456));
NAND2X1 g135928(.A (P3_IR[30] ), .B (n_1659), .Y (n_2454));
NOR2X1 g135004(.A (n_1762), .B (n_2034), .Y (n_2953));
NAND2X1 g134929(.A (n_2155), .B (n_852), .Y (n_2453));
CLKBUFX1 g134769(.A (n_33237), .Y (n_2952));
INVX2 g135150(.A (n_35159), .Y (n_2883));
AOI21X1 g134632(.A0 (n_2223), .A1 (n_2183), .B0 (n_2450), .Y(n_2864));
INVX1 g134863(.A (n_2448), .Y (n_2449));
NOR2X1 g134461(.A (n_2558), .B (n_1935), .Y (n_2447));
INVX1 g134539(.A (n_2445), .Y (n_2446));
NAND2X1 g134861(.A (n_3050), .B (n_2912), .Y (n_2444));
OAI21X1 g134645(.A0 (n_2442), .A1 (n_2055), .B0 (n_1936), .Y(n_2443));
AOI21X1 g134590(.A0 (n_2673), .A1 (n_2289), .B0 (n_2440), .Y(n_2441));
INVX1 g135019(.A (n_2438), .Y (n_2439));
NAND3X1 g134614(.A (n_2206), .B (n_2431), .C (n_1462), .Y (n_2437));
NAND2X1 g134559(.A (n_2080), .B (n_1705), .Y (n_3375));
NOR2X1 g134259(.A (n_1824), .B (n_2005), .Y (n_2436));
OR2X1 g134750(.A (n_2434), .B (n_2433), .Y (n_2435));
NAND3X1 g134629(.A (n_1869), .B (n_2206), .C (n_2431), .Y (n_2432));
AOI21X1 g134615(.A0 (n_2249), .A1 (n_2298), .B0 (n_2430), .Y(n_2877));
NAND2X1 g135879(.A (n_1964), .B (n_1659), .Y (n_2429));
INVX1 g135279(.A (n_2428), .Y (n_4143));
MX2X1 g134055(.A (n_1319), .B (n_316), .S0 (n_2577), .Y (n_2693));
AOI21X1 g134591(.A0 (n_2427), .A1 (n_2181), .B0 (n_2426), .Y(n_3000));
AOI21X1 g134584(.A0 (n_2424), .A1 (n_2423), .B0 (n_2224), .Y(n_2425));
OR2X1 g135897(.A (n_2718), .B (n_32517), .Y (n_4523));
CLKBUFX1 g135263(.A (n_2663), .Y (n_2950));
AOI21X1 g134564(.A0 (n_1700), .A1 (n_1963), .B0 (n_2422), .Y(n_2932));
AOI21X1 g134561(.A0 (n_1835), .A1 (n_1998), .B0 (n_2063), .Y(n_2847));
AOI21X1 g134628(.A0 (n_2420), .A1 (n_2419), .B0 (n_2324), .Y(n_2421));
OR2X1 g134257(.A (n_2015), .B (n_701), .Y (n_2418));
INVX1 g134813(.A (n_33431), .Y (n_2417));
NOR2X1 g134789(.A (n_2434), .B (n_2594), .Y (n_2414));
INVX1 g134459(.A (n_2412), .Y (n_2413));
AND2X1 g134714(.A (n_2409), .B (n_2408), .Y (n_2410));
OR2X1 g134808(.A (n_2406), .B (n_2405), .Y (n_2407));
NAND2X1 g134341(.A (n_1765), .B (n_1923), .Y (n_7546));
INVX1 g134771(.A (n_2195), .Y (n_3310));
INVX1 g135782(.A (n_3126), .Y (n_4917));
NAND2X1 g134794(.A (n_2404), .B (n_2243), .Y (n_2793));
OR2X1 g135017(.A (n_1906), .B (n_622), .Y (n_2403));
NAND2X1 g135104(.A (n_1064), .B (n_1861), .Y (n_2402));
INVX1 g136017(.A (n_3204), .Y (n_4802));
INVX1 g135088(.A (n_2399), .Y (n_2957));
NOR2X1 g135148(.A (n_2024), .B (n_2237), .Y (n_2537));
INVX1 g137874(.A (n_34946), .Y (n_2415));
INVX1 g135022(.A (n_2397), .Y (n_2789));
OR2X1 g134738(.A (n_1239), .B (n_33239), .Y (n_2396));
INVX1 g135142(.A (n_2395), .Y (n_3386));
NAND2X1 g134224(.A (n_2393), .B (n_2392), .Y (n_2394));
OR2X1 g134157(.A (n_1696), .B (n_1836), .Y (n_2710));
INVX1 g134966(.A (n_2515), .Y (n_2391));
INVX1 g134841(.A (n_2389), .Y (n_2390));
NAND2X1 g135026(.A (n_2387), .B (n_2504), .Y (n_2388));
INVX1 g135027(.A (n_2385), .Y (n_2386));
INVX1 g135014(.A (n_2622), .Y (n_2384));
INVX1 g135006(.A (n_2383), .Y (n_3140));
AND2X1 g135087(.A (n_2381), .B (n_2380), .Y (n_2382));
NAND3X1 g134504(.A (n_2377), .B (n_2376), .C (n_2375), .Y (n_2378));
NOR2X1 g134828(.A (n_1880), .B (n_2373), .Y (n_2374));
NAND2X1 g134875(.A (n_1795), .B (n_1785), .Y (n_2372));
OR2X1 g134531(.A (n_2275), .B (P3_reg3[5] ), .Y (n_2369));
INVX1 g135232(.A (n_2367), .Y (n_2368));
INVX1 g135046(.A (n_2366), .Y (n_2542));
OR2X1 g134862(.A (n_1768), .B (n_2364), .Y (n_2365));
NAND3X1 g134864(.A (n_2066), .B (n_1654), .C (n_1526), .Y (n_2448));
INVX1 g134956(.A (n_2433), .Y (n_2363));
NOR2X1 g134805(.A (n_32484), .B (n_1845), .Y (n_2472));
AND2X1 g134762(.A (n_2361), .B (n_2360), .Y (n_2362));
INVX1 g134998(.A (n_2468), .Y (n_2359));
OAI21X1 g135213(.A0 (n_2140), .A1 (n_1639), .B0 (n_1887), .Y(n_2507));
INVX1 g134310(.A (n_2544), .Y (n_7760));
OAI21X1 g135194(.A0 (n_2327), .A1 (n_1375), .B0 (n_1590), .Y(n_2662));
NAND2X1 g135805(.A (P3_reg3[3] ), .B (n_1017), .Y (n_13192));
AOI21X1 g134621(.A0 (n_1466), .A1 (n_2798), .B0 (n_2528), .Y(n_2812));
NAND2X1 g136351(.A (n_10563), .B (n_1803), .Y (n_2428));
INVX1 g134959(.A (n_2484), .Y (n_2639));
NOR2X1 g134889(.A (n_1790), .B (n_1956), .Y (n_2356));
CLKBUFX1 g133679(.A (n_8205), .Y (n_10594));
INVX1 g135029(.A (n_2385), .Y (n_2531));
NAND2X1 g134985(.A (n_1340), .B (n_32448), .Y (n_2355));
NAND2X1 g134785(.A (n_2164), .B (n_2352), .Y (n_2353));
AOI21X1 g134554(.A0 (n_1429), .A1 (n_2168), .B0 (n_2351), .Y(n_2729));
OAI21X1 g134581(.A0 (n_2349), .A1 (n_1973), .B0 (n_2348), .Y(n_3537));
AOI21X1 g134636(.A0 (n_2346), .A1 (n_1471), .B0 (n_1703), .Y(n_2347));
INVX1 g134662(.A (n_2138), .Y (n_2553));
NAND2X1 g134715(.A (n_2667), .B (n_2185), .Y (n_2620));
OAI21X1 g134734(.A0 (n_1838), .A1 (n_479), .B0 (n_1929), .Y (n_2344));
NAND2X1 g134740(.A (n_2342), .B (n_2341), .Y (n_2343));
NAND3X1 g134757(.A (P2_reg3[28] ), .B (n_2352), .C (n_1436), .Y(n_2340));
OR2X1 g134802(.A (n_2338), .B (n_2480), .Y (n_2339));
INVX1 g134834(.A (n_34542), .Y (n_3060));
OR2X1 g134860(.A (n_1839), .B (n_701), .Y (n_3547));
AOI21X1 g134885(.A0 (n_2012), .A1 (n_2336), .B0 (n_2065), .Y(n_3252));
NAND2X1 g134979(.A (n_2333), .B (n_2332), .Y (n_2658));
INVX1 g135056(.A (n_2331), .Y (n_2625));
AND2X1 g135055(.A (n_2240), .B (n_2329), .Y (n_2330));
INVX1 g135164(.A (n_2328), .Y (n_2792));
OAI21X1 g135221(.A0 (n_2186), .A1 (n_2286), .B0 (n_2327), .Y(n_2602));
NOR2X1 g134809(.A (n_2796), .B (n_2467), .Y (n_3276));
OR2X1 g134159(.A (n_2572), .B (n_2317), .Y (n_2325));
AOI21X1 g134627(.A0 (n_2324), .A1 (n_2069), .B0 (n_2216), .Y(n_2690));
AOI21X1 g133969(.A0 (n_3324), .A1 (n_2113), .B0 (n_2323), .Y(n_2854));
NAND2X1 g135823(.A (P1_IR[29] ), .B (n_998), .Y (n_2322));
INVX1 g134779(.A (n_2370), .Y (n_2321));
INVX1 g135082(.A (n_2475), .Y (n_2320));
OR2X1 g136066(.A (P1_reg2[0] ), .B (n_7747), .Y (n_2319));
NAND2X1 g134153(.A (n_2572), .B (n_2317), .Y (n_2318));
NAND2X1 g135063(.A (n_2288), .B (n_2312), .Y (n_2574));
NAND2X1 g134857(.A (n_1761), .B (n_2310), .Y (n_2311));
AOI21X1 g134886(.A0 (n_1782), .A1 (n_1952), .B0 (n_1913), .Y(n_2309));
NOR2X1 g134798(.A (n_2306), .B (n_1827), .Y (n_2307));
NAND2X1 g134748(.A (n_32483), .B (P1_IR[31] ), .Y (n_2305));
NAND3X1 g134879(.A (n_2303), .B (n_1958), .C (n_3509), .Y (n_2535));
INVX1 g134605(.A (n_2301), .Y (n_2302));
NOR2X1 g134768(.A (n_2129), .B (n_1757), .Y (n_2300));
NAND2X1 g134540(.A (n_1779), .B (n_1170), .Y (n_2445));
NAND3X1 g134856(.A (n_2291), .B (n_2250), .C (n_2298), .Y (n_2513));
AND2X1 g134786(.A (n_2296), .B (n_2342), .Y (n_2297));
NAND2X1 g134995(.A (n_2294), .B (n_212), .Y (n_2295));
NOR2X1 g134758(.A (n_2338), .B (n_2495), .Y (n_2293));
INVX1 g135121(.A (n_2481), .Y (n_2292));
XOR2X1 g134692(.A (n_2291), .B (n_1668), .Y (n_2680));
NOR2X1 g134522(.A (n_1884), .B (n_1818), .Y (n_2290));
INVX1 g133530(.A (n_2489), .Y (n_2596));
AND2X1 g135034(.A (n_2289), .B (n_2288), .Y (n_3005));
NOR2X1 g135465(.A (n_1947), .B (n_2286), .Y (n_2287));
NAND2X2 g134723(.A (n_1810), .B (n_1871), .Y (n_3063));
NAND2X1 g136401(.A (P1_reg2[0] ), .B (n_2779), .Y (n_2460));
AOI21X1 g134455(.A0 (n_1578), .A1 (n_3506), .B0 (n_2282), .Y(n_2283));
INVX1 g135172(.A (n_2280), .Y (n_2281));
NOR2X1 g134716(.A (n_2180), .B (n_2060), .Y (n_2825));
NAND2X1 g134819(.A (n_2266), .B (P3_reg3[8] ), .Y (n_2279));
INVX1 g135167(.A (n_2278), .Y (n_3353));
OR2X1 g135152(.A (n_999), .B (n_32448), .Y (n_2277));
NAND2X1 g134135(.A (n_2392), .B (n_2213), .Y (n_2276));
OR2X1 g134518(.A (n_2089), .B (n_2275), .Y (n_2692));
NAND2X1 g135789(.A (P1_IR[30] ), .B (n_998), .Y (n_35118));
NOR2X1 g135631(.A (n_1690), .B (n_2141), .Y (n_2271));
NAND2X1 g134520(.A (n_1454), .B (n_2306), .Y (n_2584));
INVX1 g135138(.A (n_3894), .Y (n_2270));
OR2X1 g134858(.A (n_1770), .B (n_2268), .Y (n_2269));
NAND3X1 g134732(.A (n_1974), .B (n_1351), .C (n_1445), .Y (n_2462));
OR2X1 g134766(.A (n_2266), .B (P3_reg3[8] ), .Y (n_2267));
NAND3X1 g134736(.A (n_2191), .B (n_2264), .C (n_2263), .Y (n_2265));
MX2X1 g134067(.A (P1_reg3[9] ), .B (n_169), .S0 (n_2562), .Y(n_2563));
NAND2X1 g134784(.A (n_2020), .B (n_2260), .Y (n_2261));
NAND2X1 g134510(.A (n_2275), .B (P3_reg3[5] ), .Y (n_2259));
AND2X1 g134859(.A (n_3086), .B (n_2679), .Y (n_3511));
OAI21X1 g134655(.A0 (n_2257), .A1 (n_2151), .B0 (n_1794), .Y(n_2258));
NAND2X1 g134733(.A (n_1875), .B (n_2255), .Y (n_2256));
NAND2X1 g134868(.A (n_1978), .B (n_2058), .Y (n_2254));
NAND2X1 g134509(.A (n_1788), .B (addr_461), .Y (n_2551));
AND2X1 g135103(.A (n_2252), .B (n_2288), .Y (n_2253));
AOI21X1 g134643(.A0 (n_2291), .A1 (n_2250), .B0 (n_2249), .Y(n_2873));
OR2X1 g136450(.A (n_9590), .B (n_1803), .Y (n_2248));
OR2X1 g135933(.A (n_1054), .B (n_7243), .Y (n_2247));
NAND2X1 g135032(.A (n_1704), .B (n_2244), .Y (n_2245));
OAI21X1 g134580(.A0 (n_2150), .A1 (n_2243), .B0 (n_2257), .Y(n_3352));
NAND2X1 g134565(.A (n_1695), .B (n_1687), .Y (n_2592));
AOI21X1 g134637(.A0 (n_2241), .A1 (n_2179), .B0 (n_2240), .Y(n_2242));
OR2X1 g136526(.A (n_10563), .B (n_1803), .Y (n_2239));
OAI21X1 g134666(.A0 (n_2348), .A1 (n_2237), .B0 (n_1797), .Y(n_2238));
NAND2X1 g134884(.A (n_1732), .B (n_2303), .Y (n_3945));
INVX1 g134790(.A (n_2235), .Y (n_2236));
AND2X1 g134977(.A (n_2233), .B (n_1846), .Y (n_2234));
NAND3X1 g134316(.A (n_2478), .B (n_2231), .C (n_2230), .Y (n_2232));
NAND3X1 g134881(.A (n_1737), .B (n_1110), .C (n_2229), .Y (n_2539));
NAND2X1 g135890(.A (n_286), .B (n_32509), .Y (n_4556));
AOI21X1 g134613(.A0 (n_1918), .A1 (n_2844), .B0 (n_2228), .Y(n_3795));
OR2X1 g134839(.A (n_2226), .B (n_1972), .Y (n_2227));
NOR2X1 g134178(.A (n_2577), .B (n_1771), .Y (n_8212));
NAND2X1 g135264(.A (n_1521), .B (n_1920), .Y (n_2663));
AOI21X1 g134572(.A0 (n_2224), .A1 (n_2187), .B0 (n_2223), .Y(n_2590));
AOI21X1 g134563(.A0 (n_1467), .A1 (n_2161), .B0 (n_2221), .Y(n_2222));
NAND2X1 g134558(.A (n_1850), .B (n_1919), .Y (n_2845));
NOR2X1 g134891(.A (n_1756), .B (n_2057), .Y (n_2220));
NAND2X1 g135016(.A (n_2219), .B (n_2218), .Y (n_2650));
XOR2X1 g134693(.A (n_2598), .B (n_1648), .Y (n_2217));
AOI21X1 g134578(.A0 (n_2216), .A1 (n_2122), .B0 (n_2215), .Y(n_2727));
OR2X1 g134172(.A (n_2392), .B (n_2213), .Y (n_2214));
NOR2X1 g134874(.A (n_1213), .B (n_2211), .Y (n_2212));
NAND2X1 g135020(.A (n_2210), .B (n_2209), .Y (n_2438));
NAND2X1 g134345(.A (n_1777), .B (n_1780), .Y (n_8193));
NOR2X1 g134825(.A (n_2461), .B (n_2158), .Y (n_2208));
NAND2X1 g134460(.A (n_1786), .B (addr_442), .Y (n_2412));
INVX1 g134990(.A (n_2284), .Y (n_2207));
NAND2X1 g134767(.A (n_2206), .B (n_1240), .Y (n_2554));
AND2X1 g135071(.A (n_2204), .B (n_2172), .Y (n_2205));
NAND2X1 g135778(.A (P3_IR[28] ), .B (n_1659), .Y (n_2203));
NOR2X1 g135174(.A (n_1610), .B (n_1937), .Y (n_3188));
NOR2X1 g135013(.A (n_1503), .B (n_1622), .Y (n_2202));
INVX1 g135057(.A (n_33434), .Y (n_2331));
NAND2X1 g135007(.A (n_2556), .B (n_2200), .Y (n_2383));
NAND3X1 g134735(.A (P1_reg3[28] ), .B (n_2260), .C (n_1308), .Y(n_2199));
XOR2X1 g134695(.A (n_707), .B (n_1140), .Y (n_2198));
NOR2X1 g134778(.A (n_1432), .B (n_2196), .Y (n_2197));
NAND3X1 g134772(.A (n_944), .B (n_2194), .C (n_721), .Y (n_2195));
NAND2X1 g134706(.A (n_2375), .B (n_2105), .Y (n_2193));
AND2X1 g135128(.A (n_2192), .B (n_965), .Y (n_2409));
AND2X1 g135117(.A (n_2191), .B (n_2190), .Y (n_3168));
NOR2X1 g135090(.A (n_1856), .B (n_1644), .Y (n_2834));
INVX1 g136970(.A (n_34668), .Y (n_2189));
NAND2X1 g135091(.A (n_2423), .B (n_2187), .Y (n_2405));
OAI21X1 g135181(.A0 (n_1865), .A1 (n_1536), .B0 (n_2186), .Y(n_2426));
NAND2X1 g135993(.A (P1_reg3[11] ), .B (n_2174), .Y (n_12723));
AND2X1 g135118(.A (n_2185), .B (n_1214), .Y (n_2547));
NAND2X1 g135630(.A (n_2186), .B (n_1302), .Y (n_2184));
NAND2X1 g135059(.A (n_2183), .B (n_2187), .Y (n_2649));
NAND2X1 g135023(.A (n_2182), .B (n_2181), .Y (n_2397));
INVX1 g135083(.A (n_2180), .Y (n_2475));
NAND2X1 g135037(.A (n_2191), .B (n_2179), .Y (n_2434));
AOI21X1 g135248(.A0 (n_1966), .A1 (n_1630), .B0 (n_2178), .Y(n_2775));
NAND2X1 g133828(.A (n_13167), .B (n_3217), .Y (n_2177));
OR2X1 g134419(.A (n_2137), .B (P1_reg3[12] ), .Y (n_2176));
INVX1 g133690(.A (n_2175), .Y (n_10880));
NAND2X1 g135889(.A (P1_reg3[7] ), .B (n_2174), .Y (n_12820));
AOI21X1 g135246(.A0 (n_2178), .A1 (n_2173), .B0 (n_1249), .Y(n_2776));
NAND2X1 g135000(.A (n_2172), .B (n_2077), .Y (n_2468));
OR2X1 g134827(.A (n_2170), .B (n_2169), .Y (n_2171));
NAND2X1 g135047(.A (n_2168), .B (n_1399), .Y (n_2366));
XOR2X1 g134101(.A (n_1257), .B (n_3022), .Y (n_2167));
INVX1 g134927(.A (n_2164), .Y (n_2165));
AOI21X1 g134617(.A0 (n_2162), .A1 (n_2147), .B0 (n_2161), .Y(n_2163));
AND2X1 g135111(.A (n_2159), .B (n_2158), .Y (n_2160));
NOR2X1 g135116(.A (n_2179), .B (n_2329), .Y (n_2156));
INVX1 g135289(.A (n_33921), .Y (n_2155));
OR2X1 g135165(.A (n_2151), .B (n_2150), .Y (n_2328));
NOR2X1 g135388(.A (n_2148), .B (n_1579), .Y (n_2149));
NAND3X1 g134842(.A (n_1255), .B (n_1139), .C (n_2147), .Y (n_2389));
OR2X1 g135185(.A (n_1434), .B (n_2146), .Y (n_2483));
NAND3X1 g133605(.A (n_1238), .B (n_1169), .C (n_1517), .Y (n_2605));
NOR2X1 g135133(.A (n_2094), .B (n_1518), .Y (n_4280));
NAND2X1 g135039(.A (n_2181), .B (n_2312), .Y (n_2781));
NOR2X1 g134749(.A (n_2931), .B (n_2052), .Y (n_2145));
NAND2X1 g134953(.A (n_2190), .B (n_2119), .Y (n_2594));
INVX1 g134960(.A (n_33373), .Y (n_2484));
INVX1 g134383(.A (n_1911), .Y (n_2379));
OAI21X1 g135224(.A0 (n_2117), .A1 (n_2141), .B0 (n_2140), .Y(n_2430));
OR2X1 g135168(.A (n_2150), .B (n_2097), .Y (n_2278));
OR2X1 g134549(.A (n_2137), .B (n_1437), .Y (n_2523));
AND2X1 g135051(.A (n_1817), .B (n_2074), .Y (n_2642));
AND2X1 g135049(.A (n_2600), .B (n_2135), .Y (n_2136));
AND2X1 g135015(.A (n_2172), .B (n_2125), .Y (n_2622));
AOI21X1 g133986(.A0 (n_3022), .A1 (n_1565), .B0 (n_2047), .Y(n_2637));
NAND2X1 g135888(.A (P1_reg3[18] ), .B (n_2091), .Y (n_12806));
NAND2X1 g134182(.A (n_3022), .B (n_2634), .Y (n_2134));
NAND2X1 g135089(.A (n_2133), .B (n_2179), .Y (n_2399));
NOR2X1 g135042(.A (n_2131), .B (n_2229), .Y (n_2132));
INVX1 g135093(.A (n_2129), .Y (n_2130));
INVX1 g135030(.A (n_34324), .Y (n_2385));
AOI21X1 g134607(.A0 (n_2126), .A1 (n_2125), .B0 (n_2124), .Y(n_2127));
NAND2X1 g133680(.A (n_1614), .B (n_1457), .Y (n_8205));
NAND3X1 g134867(.A (n_681), .B (n_1070), .C (addr_439), .Y (n_2123));
NAND2X1 g134983(.A (n_2333), .B (n_2122), .Y (n_2458));
NOR2X1 g135555(.A (n_1559), .B (n_2118), .Y (n_2121));
NAND2X1 g135085(.A (n_2119), .B (n_2229), .Y (n_2120));
NOR2X1 g135132(.A (n_1386), .B (n_2151), .Y (n_4282));
OAI21X1 g135200(.A0 (n_1608), .A1 (n_1901), .B0 (n_1867), .Y(n_2712));
OAI21X1 g135205(.A0 (n_1864), .A1 (n_2118), .B0 (n_2117), .Y(n_2499));
NAND2X1 g134958(.A (n_2116), .B (n_2115), .Y (n_2566));
AND2X1 g135068(.A (n_2114), .B (n_2113), .Y (n_2948));
INVX1 g135225(.A (n_2111), .Y (n_2112));
INVX1 g135237(.A (n_2109), .Y (n_2110));
INVX1 g134925(.A (n_1801), .Y (n_2334));
AOI21X1 g134608(.A0 (n_1683), .A1 (n_1632), .B0 (n_1416), .Y(n_2107));
OR2X1 g134712(.A (n_2375), .B (n_2105), .Y (n_2106));
NAND2X1 g136018(.A (n_565), .B (n_32517), .Y (n_3204));
OAI21X1 g134654(.A0 (n_1626), .A1 (n_10838), .B0 (n_3534), .Y(so[0]));
NAND2X1 g134993(.A (n_2101), .B (n_2116), .Y (n_2284));
NOR2X1 g135092(.A (n_2158), .B (n_2098), .Y (n_2099));
NAND2X1 g134824(.A (n_2097), .B (n_2243), .Y (n_2791));
INVX1 g134914(.A (n_1970), .Y (n_2400));
NOR2X1 g134763(.A (n_2494), .B (n_2094), .Y (n_2095));
NAND2X1 g135857(.A (P1_reg3[9] ), .B (n_2091), .Y (n_12728));
NOR2X1 g134707(.A (n_1689), .B (n_2089), .Y (n_2090));
NAND2X1 g135924(.A (P1_reg3[6] ), .B (n_2174), .Y (n_12822));
CLKBUFX1 gbuf_d_702(.A(n_1621), .Y(d_out_702));
CLKBUFX1 gbuf_qn_702(.A(qn_in_702), .Y(P2_n_749));
NAND2X1 g135964(.A (P1_reg3[15] ), .B (n_2174), .Y (n_12818));
OR2X1 g134311(.A (n_2562), .B (n_1805), .Y (n_2544));
NAND2X1 g135797(.A (n_10854), .B (n_2070), .Y (n_13093));
NAND4X1 g134586(.A (n_2086), .B (n_74), .C (n_2085), .D (n_2084), .Y(n_2087));
AOI21X1 g134633(.A0 (n_2046), .A1 (n_1399), .B0 (n_1428), .Y(n_2083));
NOR2X1 g135069(.A (n_2081), .B (n_1450), .Y (n_2082));
INVX1 g135277(.A (n_2497), .Y (n_2313));
NAND3X1 g134801(.A (n_2079), .B (n_2078), .C (n_2077), .Y (n_2080));
INVX1 g135281(.A (n_2076), .Y (n_4258));
AND2X1 g135048(.A (n_1501), .B (n_2074), .Y (n_2075));
NAND3X1 g134849(.A (n_2072), .B (n_2071), .C (n_2043), .Y (n_2073));
NAND2X1 g135816(.A (P1_reg3[3] ), .B (n_2070), .Y (n_12732));
NAND2X1 g134964(.A (n_2122), .B (n_2069), .Y (n_2657));
NOR2X1 g133531(.A (n_1525), .B (n_536), .Y (n_2489));
NAND2X1 g135796(.A (n_10566), .B (n_2070), .Y (n_12810));
NAND2X1 g135110(.A (n_2219), .B (n_2183), .Y (n_2406));
NAND2X1 g134747(.A (n_1971), .B (n_1682), .Y (n_2068));
NAND2X1 g135751(.A (n_1458), .B (n_2066), .Y (n_2067));
NOR2X1 g134791(.A (n_2065), .B (n_2059), .Y (n_2235));
NAND3X1 g134781(.A (n_608), .B (n_2064), .C (n_1541), .Y (n_2370));
AOI21X1 g134606(.A0 (n_2063), .A1 (n_1830), .B0 (n_2126), .Y(n_2301));
NAND2X1 g134433(.A (n_2137), .B (P1_reg3[12] ), .Y (n_2062));
INVX1 g134917(.A (n_2060), .Y (n_2061));
NAND2X1 g135123(.A (n_2074), .B (n_2059), .Y (n_2481));
NAND2X1 g135173(.A (n_2058), .B (n_2057), .Y (n_2280));
NOR2X1 g135722(.A (n_2055), .B (n_1448), .Y (n_2056));
NAND2X1 g134817(.A (n_1178), .B (n_2053), .Y (n_2054));
NOR2X1 g135064(.A (n_1412), .B (n_1440), .Y (n_2876));
NOR2X1 g135170(.A (n_1509), .B (n_2052), .Y (n_3189));
XOR2X1 g134694(.A (n_2798), .B (n_1111), .Y (n_2051));
NAND2X1 g135907(.A (P2_reg3[27] ), .B (n_1336), .Y (n_2050));
NOR2X1 g135070(.A (n_2263), .B (n_2190), .Y (n_2049));
NAND3X1 g134837(.A (n_741), .B (n_2048), .C (n_1289), .Y (n_2955));
AOI21X1 g134616(.A0 (n_2047), .A1 (n_1566), .B0 (n_2046), .Y(n_2538));
NOR2X1 g135158(.A (n_1511), .B (n_2044), .Y (n_2045));
NAND2X1 g135783(.A (n_2718), .B (n_32517), .Y (n_3126));
NAND2X1 g135143(.A (n_2043), .B (n_1907), .Y (n_2395));
NAND2X1 g134807(.A (n_2170), .B (n_2041), .Y (n_2042));
NAND2X1 g134957(.A (n_2133), .B (n_2115), .Y (n_2433));
INVX1 g134922(.A (n_33374), .Y (n_35271));
NAND2X1 g135155(.A (n_2037), .B (n_2094), .Y (n_2038));
NAND2X1 g135038(.A (n_1709), .B (n_2035), .Y (n_2036));
NAND2X1 g134826(.A (n_1879), .B (n_2721), .Y (n_2549));
INVX1 g135579(.A (n_2033), .Y (n_2034));
NOR2X1 g135134(.A (n_1564), .B (n_2169), .Y (n_3050));
AND2X1 g135114(.A (n_2031), .B (n_2951), .Y (n_2032));
AND2X1 g134810(.A (n_1618), .B (n_2375), .Y (n_2469));
AND2X1 g135177(.A (n_743), .B (n_1860), .Y (n_2030));
NAND2X1 g135878(.A (P1_reg3[5] ), .B (n_2091), .Y (n_12824));
NOR2X1 g134974(.A (n_2252), .B (n_2289), .Y (n_2029));
OR2X1 g135937(.A (n_600), .B (P2_IR[31] ), .Y (n_2028));
INVX1 g135078(.A (n_2849), .Y (n_2026));
NAND2X1 g136026(.A (P1_reg3[12] ), .B (n_2091), .Y (n_12808));
NOR2X1 g134948(.A (n_1397), .B (n_33432), .Y (n_35278));
INVX1 g134941(.A (n_2020), .Y (n_2021));
CLKBUFX1 gbuf_d_703(.A(n_349), .Y(d_out_703));
CLKBUFX1 gbuf_qn_703(.A(qn_in_703), .Y(n_349));
NAND2X1 g134986(.A (n_2200), .B (n_2298), .Y (n_2017));
INVX1 g135040(.A (n_2016), .Y (n_2623));
AOI21X1 g134658(.A0 (n_1549), .A1 (n_1754), .B0 (n_1477), .Y(n_2015));
NAND2X1 g135988(.A (P1_reg3[17] ), .B (n_2091), .Y (n_12714));
AOI21X1 g134631(.A0 (n_2422), .A1 (n_1438), .B0 (n_2012), .Y(n_2013));
NOR2X1 g135233(.A (n_1641), .B (n_2011), .Y (n_2367));
NOR2X1 g135139(.A (n_2009), .B (n_2094), .Y (n_3894));
NAND2X1 g135843(.A (P1_reg3[16] ), .B (n_2174), .Y (n_12812));
NOR2X1 g135180(.A (n_2037), .B (n_2009), .Y (n_2010));
INVX1 g134937(.A (n_34203), .Y (n_35427));
AOI21X1 g134610(.A0 (n_2004), .A1 (n_1962), .B0 (n_1699), .Y(n_2005));
NAND2X1 g135865(.A (P1_reg3[4] ), .B (n_2070), .Y (n_13091));
AND2X1 g135072(.A (n_2289), .B (n_2582), .Y (n_2801));
INVX1 g134935(.A (n_34536), .Y (n_2003));
AND2X1 g134954(.A (n_2000), .B (n_2882), .Y (n_2001));
NAND2X1 g135845(.A (P1_reg3[19] ), .B (n_2091), .Y (n_12814));
AOI21X1 g134587(.A0 (n_2351), .A1 (n_1808), .B0 (n_1998), .Y(n_1999));
AOI21X1 g135260(.A0 (n_1353), .A1 (n_1959), .B0 (n_1200), .Y(n_1997));
NAND2X1 g135822(.A (n_11135), .B (n_2070), .Y (n_12816));
AOI21X1 g135251(.A0 (n_1863), .A1 (n_1232), .B0 (n_1569), .Y(n_2500));
NAND2X1 g134968(.A (n_2182), .B (n_1996), .Y (n_2515));
NAND2X1 g135363(.A (n_1993), .B (n_1853), .Y (n_1994));
NAND2X1 g134527(.A (n_1451), .B (n_1522), .Y (n_1992));
AND2X1 g134976(.A (n_2131), .B (n_2119), .Y (n_1991));
NAND2X1 g135965(.A (P1_reg3[8] ), .B (n_2174), .Y (n_12730));
AOI21X1 g134579(.A0 (n_2221), .A1 (n_1663), .B0 (n_1693), .Y(n_1990));
INVX1 g134871(.A (n_2569), .Y (n_1989));
NAND2X1 g135779(.A (P1_reg3[13] ), .B (n_2174), .Y (n_12718));
NAND2X1 g135780(.A (P1_reg3[10] ), .B (n_2091), .Y (n_12712));
NOR2X1 g135036(.A (n_1933), .B (n_1987), .Y (n_2881));
NAND2X1 g135806(.A (P1_reg3[14] ), .B (n_2174), .Y (n_12716));
OR2X1 g135306(.A (n_35224), .B (n_33587), .Y (n_1986));
NAND2X1 g136107(.A (n_9634), .B (n_1313), .Y (n_1985));
NAND3X1 g134918(.A (n_32475), .B (n_33351), .C (n_629), .Y (n_2060));
AND2X1 g134984(.A (n_2486), .B (n_1979), .Y (n_1980));
NOR2X1 g135156(.A (n_1977), .B (n_2041), .Y (n_1978));
NAND3X1 g134585(.A (n_1484), .B (P2_reg3[7] ), .C (n_1976), .Y(n_2577));
OR2X1 g135544(.A (n_1133), .B (n_2779), .Y (n_1974));
NOR2X1 g135136(.A (n_1973), .B (n_1767), .Y (n_3538));
INVX1 g135112(.A (n_1971), .Y (n_1972));
NAND3X1 g134915(.A (n_1969), .B (n_1562), .C (n_1968), .Y (n_1970));
NOR2X1 g135699(.A (n_1966), .B (n_1044), .Y (n_1967));
NOR2X1 g134933(.A (n_1113), .B (n_1964), .Y (n_1965));
INVX1 g137452(.A (n_1444), .Y (n_7747));
AND2X1 g135120(.A (n_1963), .B (n_1962), .Y (n_2342));
INVX1 g135066(.A (n_2206), .Y (n_2266));
INVX1 g134950(.A (n_2516), .Y (n_1961));
AND2X1 g135686(.A (n_1959), .B (n_1958), .Y (n_1960));
AND2X1 g135137(.A (n_1957), .B (n_1956), .Y (n_3630));
NAND2X1 g135094(.A (n_1955), .B (n_34526), .Y (n_2129));
OAI21X1 g135195(.A0 (n_1886), .A1 (n_1572), .B0 (n_1894), .Y(n_2420));
AOI21X1 g134594(.A0 (n_856), .A1 (n_835), .B0 (n_2162), .Y (n_2455));
NAND3X1 g134872(.A (n_1749), .B (n_1778), .C (n_1952), .Y (n_2569));
NAND2X1 g135421(.A (n_1508), .B (n_1154), .Y (n_1951));
NAND2X1 g135050(.A (n_34853), .B (n_1949), .Y (n_1950));
INVX1 g136997(.A (n_35024), .Y (n_31470));
INVX1 g136101(.A (n_2327), .Y (n_1947));
AND2X1 g135079(.A (n_1945), .B (n_1944), .Y (n_2849));
NOR2X1 g135836(.A (n_991), .B (n_1677), .Y (n_1943));
NOR2X1 g135149(.A (n_1942), .B (n_2097), .Y (n_3001));
INVX1 g135610(.A (n_2231), .Y (n_1941));
NAND3X1 g135003(.A (n_34318), .B (n_1939), .C (n_33113), .Y (n_1940));
NAND2X1 g135991(.A (n_9634), .B (n_1336), .Y (n_12960));
NOR2X1 g135157(.A (n_1942), .B (n_1937), .Y (n_4014));
AND2X1 g135244(.A (n_1334), .B (n_1936), .Y (n_2211));
INVX1 g135010(.A (n_1935), .Y (n_2188));
INVX1 g135613(.A (n_1933), .Y (n_1934));
OR2X1 g135144(.A (n_1932), .B (n_1931), .Y (n_2404));
NOR2X1 g135754(.A (n_1263), .B (n_1495), .Y (n_1930));
NOR2X1 g135163(.A (n_1973), .B (n_2237), .Y (n_2679));
AOI21X1 g135249(.A0 (n_1928), .A1 (n_1479), .B0 (n_1000), .Y(n_1929));
NOR2X1 g134840(.A (n_2046), .B (n_1427), .Y (n_1927));
NAND2X1 g135986(.A (P2_reg3[19] ), .B (n_3834), .Y (n_12955));
NAND2X1 g135166(.A (n_1924), .B (n_2237), .Y (n_1925));
OR2X1 g134535(.A (n_1897), .B (P1_reg3[7] ), .Y (n_1923));
NAND2X1 g135491(.A (n_1759), .B (n_1168), .Y (n_1922));
OR2X1 g135828(.A (n_593), .B (n_4371), .Y (n_1921));
NOR2X1 g135646(.A (n_597), .B (n_915), .Y (n_2210));
NAND2X1 g135502(.A (n_1126), .B (n_32928), .Y (n_1920));
INVX1 g135187(.A (n_1918), .Y (n_1919));
INVX1 g135129(.A (n_4334), .Y (n_1917));
AND2X1 g135241(.A (n_1251), .B (n_1916), .Y (n_2442));
INVX1 g134920(.A (n_1733), .Y (n_1915));
NAND2X1 g134978(.A (n_1694), .B (n_1962), .Y (n_2338));
INVX1 g137030(.A (n_15968), .Y (n_31601));
AOI22X1 g134887(.A0 (n_1914), .A1 (n_1750), .B0 (n_735), .B1(n_1913), .Y (n_2559));
NAND2X1 g135508(.A (n_1908), .B (n_1371), .Y (n_1912));
NOR2X1 g135005(.A (n_2204), .B (n_2125), .Y (n_1910));
OAI21X1 g135226(.A0 (n_1908), .A1 (n_1468), .B0 (n_1899), .Y(n_2111));
OAI21X1 g135216(.A0 (n_1904), .A1 (n_1419), .B0 (n_1821), .Y(n_2660));
INVX1 g135709(.A (n_1907), .Y (n_2024));
INVX1 g134962(.A (n_2841), .Y (n_2341));
AND2X1 g135506(.A (n_1552), .B (n_1157), .Y (n_2288));
OAI21X1 g135204(.A0 (n_1697), .A1 (n_1588), .B0 (n_1593), .Y(n_2564));
OR2X1 g135523(.A (n_35223), .B (n_33814), .Y (n_1906));
OAI21X1 g135207(.A0 (n_1605), .A1 (n_1516), .B0 (n_1904), .Y(n_2461));
INVX1 g135125(.A (n_1902), .Y (n_1903));
OAI21X1 g135197(.A0 (n_1607), .A1 (n_1855), .B0 (n_1901), .Y(n_2509));
NAND2X1 g135641(.A (n_1899), .B (n_1115), .Y (n_1900));
NOR2X1 g134472(.A (n_1898), .B (n_1897), .Y (n_2572));
NAND2X1 g134699(.A (n_1688), .B (n_2721), .Y (n_2275));
NAND2X1 g135391(.A (n_1894), .B (n_1093), .Y (n_1895));
NOR2X1 g135086(.A (n_1241), .B (n_1893), .Y (n_2431));
NOR2X1 g134830(.A (n_1898), .B (n_1673), .Y (n_1892));
AND2X1 g135012(.A (n_1092), .B (n_2086), .Y (n_2936));
OR2X1 g136021(.A (n_1890), .B (n_1124), .Y (n_1891));
OAI21X1 g135214(.A0 (n_1675), .A1 (n_1651), .B0 (n_1872), .Y(n_2223));
NAND2X1 g136027(.A (P2_reg3[4] ), .B (n_1336), .Y (n_12966));
OAI21X1 g135215(.A0 (n_1887), .A1 (n_1595), .B0 (n_1886), .Y(n_2557));
NAND2X1 g135052(.A (n_1560), .B (n_2147), .Y (n_1885));
NOR2X1 g134739(.A (n_2611), .B (n_1848), .Y (n_1884));
INVX1 g136979(.A (n_15722), .Y (n_31092));
INVX1 g135080(.A (n_4024), .Y (n_1883));
NOR2X1 g135135(.A (n_1881), .B (n_2169), .Y (n_1882));
INVX1 g134909(.A (n_1879), .Y (n_1880));
AND2X1 g134916(.A (n_1123), .B (n_1878), .Y (n_3309));
NAND2X1 g135916(.A (n_33579), .B (P2_IR[24] ), .Y (n_1877));
INVX1 g134946(.A (n_1874), .Y (n_1875));
NAND2X1 g135334(.A (n_1872), .B (n_1321), .Y (n_1873));
AOI22X1 g135247(.A0 (n_724), .A1 (n_32505), .B0 (n_32938), .B1(n_1870), .Y (n_1871));
INVX1 g135145(.A (n_1868), .Y (n_1869));
OAI21X1 g135186(.A0 (n_1867), .A1 (n_1739), .B0 (n_1866), .Y(n_2427));
OAI21X1 g135196(.A0 (n_1715), .A1 (n_1488), .B0 (n_1908), .Y(n_2450));
OAI21X1 g135206(.A0 (n_1671), .A1 (n_1866), .B0 (n_1865), .Y(n_2603));
OAI21X1 g135220(.A0 (n_1667), .A1 (n_1327), .B0 (n_1864), .Y(n_2249));
OAI21X1 g135230(.A0 (n_1134), .A1 (n_1498), .B0 (n_1760), .Y(n_2528));
AOI21X1 g135245(.A0 (n_1653), .A1 (n_2066), .B0 (n_1863), .Y(n_2306));
INVX1 g135298(.A (n_1860), .Y (n_1861));
NOR2X1 g135301(.A (n_33362), .B (n_1858), .Y (n_32156));
INVX1 g135352(.A (n_1856), .Y (n_1857));
NAND2X1 g135606(.A (n_1284), .B (n_1855), .Y (n_2240));
AND2X1 g135546(.A (n_1854), .B (n_1853), .Y (n_2218));
NAND2X1 g135563(.A (n_1864), .B (n_1035), .Y (n_1852));
NOR2X1 g135404(.A (n_1350), .B (n_1496), .Y (n_1851));
NAND3X1 g134782(.A (n_1849), .B (n_1658), .C (n_1848), .Y (n_1850));
NOR2X1 g135692(.A (n_1341), .B (n_1551), .Y (n_1847));
INVX1 g135317(.A (n_1845), .Y (n_1846));
NAND2X1 g135556(.A (n_1904), .B (n_1100), .Y (n_1844));
INVX1 g134648(.A (n_1841), .Y (n_2100));
NAND2X1 g135532(.A (n_1887), .B (n_1160), .Y (n_1840));
NAND2X1 g134975(.A (n_1838), .B (n_1158), .Y (n_1839));
NOR2X1 g134797(.A (n_1836), .B (n_2196), .Y (n_1837));
NAND2X1 g135990(.A (n_1319), .B (n_1812), .Y (n_12871));
AND2X1 g135106(.A (n_1834), .B (n_1831), .Y (n_1835));
INVX1 g136999(.A (n_35024), .Y (n_31541));
NAND2X1 g135041(.A (n_1831), .B (n_1830), .Y (n_2016));
INVX1 g137000(.A (n_35024), .Y (n_31472));
NAND2X1 g135141(.A (n_1828), .B (n_1827), .Y (n_1829));
INVX1 g135398(.A (n_2114), .Y (n_1826));
INVX1 g135384(.A (n_1825), .Y (n_3591));
NOR2X1 g134988(.A (n_1962), .B (n_1823), .Y (n_1824));
NAND2X1 g135514(.A (n_1821), .B (n_1194), .Y (n_1822));
AOI21X1 g134869(.A0 (n_1849), .A1 (n_1848), .B0 (n_1817), .Y(n_1818));
NAND3X1 g135084(.A (n_474), .B (n_33355), .C (n_1444), .Y (n_2180));
AOI21X1 g134893(.A0 (n_2989), .A1 (n_1813), .B0 (n_1145), .Y(n_1814));
NAND2X1 g135861(.A (n_1976), .B (n_1812), .Y (n_12894));
OAI21X1 g135193(.A0 (n_1894), .A1 (n_1573), .B0 (n_1545), .Y(n_2424));
NAND2X1 g135323(.A (n_1867), .B (n_1061), .Y (n_1811));
NAND2X1 g135654(.A (n_1338), .B (n_32517), .Y (n_1810));
NOR2X1 g134987(.A (n_1834), .B (n_1808), .Y (n_1809));
NAND2X1 g134949(.A (n_1808), .B (n_1831), .Y (n_2796));
NOR2X1 g135131(.A (n_1881), .B (n_1807), .Y (n_2912));
NAND2X1 g136536(.A (P1_reg1[0] ), .B (n_2779), .Y (n_2497));
NOR2X1 g134942(.A (n_1805), .B (n_1307), .Y (n_2020));
OR2X1 g135534(.A (n_2011), .B (n_1640), .Y (n_1804));
NAND2X1 g136119(.A (n_9590), .B (n_1803), .Y (n_2076));
AOI22X1 g135757(.A0 (n_147), .A1 (n_194), .B0 (addr_442), .B1(addr_461), .Y (n_1802));
NOR2X1 g135345(.A (n_1166), .B (n_1346), .Y (n_2294));
NAND3X1 g134926(.A (n_33436), .B (n_1800), .C (n_1799), .Y (n_1801));
OAI21X1 g135209(.A0 (n_1604), .A1 (n_1580), .B0 (n_1297), .Y(n_2673));
NOR2X1 g135171(.A (n_1797), .B (n_1924), .Y (n_1798));
INVX1 g135740(.A (n_2009), .Y (n_1796));
NOR2X1 g135179(.A (n_1794), .B (n_1793), .Y (n_1795));
NAND2X1 g135901(.A (P2_reg3[17] ), .B (n_1812), .Y (n_12883));
OR2X1 g134907(.A (n_1347), .B (n_1787), .Y (n_1791));
NOR2X1 g135169(.A (n_2268), .B (n_1789), .Y (n_1790));
NAND4X1 g134764(.A (n_587), .B (n_1787), .C (n_555), .D (n_500), .Y(n_1788));
NAND2X1 g135119(.A (n_2069), .B (n_2419), .Y (n_2457));
NOR2X1 g135580(.A (n_1261), .B (n_35637), .Y (n_2033));
OR2X1 g135693(.A (n_2178), .B (n_748), .Y (n_4778));
NAND4X1 g134803(.A (n_494), .B (n_21), .C (n_558), .D (n_525), .Y(n_1786));
AND2X1 g135153(.A (n_2992), .B (n_1785), .Y (n_4179));
NAND2X1 g135390(.A (n_1901), .B (n_1157), .Y (n_1784));
INVX1 g135576(.A (n_1782), .Y (n_1783));
AND2X1 g135387(.A (n_1231), .B (n_1854), .Y (n_2332));
INVX1 g137166(.A (n_1659), .Y (n_4112));
OR2X1 g134538(.A (n_1300), .B (P2_reg3[7] ), .Y (n_1780));
NAND4X1 g134815(.A (n_412), .B (n_1711), .C (n_433), .D (n_596), .Y(n_1779));
AND2X1 g135098(.A (n_1944), .B (n_1778), .Y (n_3250));
NAND2X1 g134473(.A (n_1300), .B (P2_reg3[7] ), .Y (n_1777));
NAND2X1 g136509(.A (n_10562), .B (n_1313), .Y (n_1775));
NOR2X1 g135447(.A (n_1589), .B (n_1132), .Y (n_1774));
NAND2X1 g135493(.A (n_1865), .B (n_1068), .Y (n_1772));
NOR2X1 g134928(.A (n_1771), .B (n_1435), .Y (n_2164));
OR2X1 g135176(.A (n_1937), .B (n_1789), .Y (n_1770));
NAND2X1 g135161(.A (n_1793), .B (n_2151), .Y (n_1769));
OR2X1 g135178(.A (n_1767), .B (n_1766), .Y (n_1768));
NAND2X1 g134458(.A (n_1897), .B (P1_reg3[7] ), .Y (n_1765));
MX2X1 g134664(.A (n_321), .B (P1_reg3[8] ), .S0 (n_2226), .Y(n_2138));
INVX1 g135509(.A (n_1762), .Y (n_1763));
NOR2X1 g135154(.A (n_1828), .B (n_1746), .Y (n_1761));
OAI21X1 g135184(.A0 (n_1760), .A1 (n_1497), .B0 (n_1759), .Y(n_2323));
NAND2X1 g134832(.A (n_1003), .B (n_3217), .Y (n_1758));
INVX1 g135551(.A (n_1757), .Y (n_2380));
NOR2X1 g135159(.A (n_2364), .B (n_1766), .Y (n_1756));
NAND3X1 g134873(.A (n_1259), .B (n_3526), .C (n_1754), .Y (n_3485));
INVX1 g135463(.A (n_2098), .Y (n_2152));
NAND2X1 g135870(.A (P2_reg3[12] ), .B (n_1812), .Y (n_12873));
NOR2X1 g134502(.A (n_1836), .B (n_1300), .Y (n_2392));
MX2X1 g133691(.A (n_327), .B (P1_reg3[6] ), .S0 (n_1524), .Y(n_2175));
NAND2X1 g135109(.A (n_2125), .B (n_1830), .Y (n_2467));
NAND3X1 g134876(.A (n_1750), .B (n_1749), .C (n_4100), .Y (n_2558));
NOR2X1 g135522(.A (n_1748), .B (n_1612), .Y (n_4856));
INVX1 g135096(.A (n_1747), .Y (n_3492));
NOR2X1 g135160(.A (n_1746), .B (n_2052), .Y (n_3441));
NAND2X1 g135593(.A (n_1886), .B (n_1290), .Y (n_1745));
NOR2X1 g135629(.A (n_1333), .B (n_1537), .Y (n_1742));
NOR2X1 g135524(.A (n_1159), .B (n_1739), .Y (n_1740));
NAND2X1 g135527(.A (n_1760), .B (n_1737), .Y (n_1738));
NOR2X1 g135371(.A (n_1023), .B (n_1102), .Y (n_2387));
NAND2X1 g136535(.A (n_11135), .B (n_3217), .Y (n_1735));
NOR2X1 g135140(.A (n_1532), .B (n_2055), .Y (n_1732));
NAND2X1 g134811(.A (n_1183), .B (n_1313), .Y (n_1731));
NAND3X1 g134970(.A (n_33363), .B (n_33355), .C (n_33361), .Y(n_32484));
INVX1 g134939(.A (n_1728), .Y (n_1729));
NAND2X1 g135308(.A (n_33364), .B (P1_IR[31] ), .Y (n_1727));
NAND2X1 g135302(.A (n_1179), .B (n_1724), .Y (n_1725));
AND2X1 g135035(.A (n_1808), .B (n_2168), .Y (n_2465));
INVX1 g135024(.A (n_3283), .Y (n_1723));
INVX1 g135761(.A (n_7734), .Y (n_2096));
NOR2X1 g135175(.A (n_1447), .B (n_1767), .Y (n_3086));
NAND2X1 g136368(.A (n_10566), .B (n_1677), .Y (n_1722));
AND2X1 g136510(.A (n_10854), .B (n_15723), .Y (n_1721));
INVX1 g135256(.A (n_1719), .Y (n_2667));
OR2X1 g135795(.A (n_1107), .B (n_1124), .Y (n_1718));
NAND2X1 g135936(.A (P2_reg3[14] ), .B (n_1812), .Y (n_12888));
NOR2X1 g134934(.A (n_1220), .B (P2_IR[29] ), .Y (n_1717));
OAI21X1 g135222(.A0 (n_1872), .A1 (n_1652), .B0 (n_1715), .Y(n_2215));
AOI21X1 g135238(.A0 (n_1263), .A1 (n_1629), .B0 (n_1966), .Y(n_2109));
NAND2X1 g135892(.A (P2_reg3[16] ), .B (n_1812), .Y (n_12886));
OR2X1 g134908(.A (n_1056), .B (n_1711), .Y (n_1712));
INVX1 g135416(.A (n_1709), .Y (n_1710));
NAND2X1 g135320(.A (n_1715), .B (n_1114), .Y (n_1708));
NAND2X1 g135162(.A (n_2044), .B (n_2052), .Y (n_1707));
INVX1 g135520(.A (n_1703), .Y (n_1704));
NOR2X1 g135124(.A (n_1701), .B (n_2147), .Y (n_1702));
AND2X1 g135074(.A (n_1699), .B (n_1823), .Y (n_1700));
NOR2X1 g135456(.A (n_1202), .B (n_1697), .Y (n_1698));
OR2X1 g134476(.A (n_2196), .B (n_1300), .Y (n_1696));
NAND3X1 g134776(.A (n_1694), .B (n_1693), .C (n_1692), .Y (n_1695));
AND2X1 g134994(.A (n_1311), .B (n_1691), .Y (n_2361));
INVX1 g136421(.A (n_2140), .Y (n_1690));
INVX1 g134911(.A (n_1688), .Y (n_1689));
INVX1 g135182(.A (n_2004), .Y (n_1687));
XOR2X1 g135773(.A (si[0]), .B (n_275), .Y (n_1686));
NAND2X1 g135853(.A (P2_reg3[3] ), .B (P2_n_749), .Y (n_12962));
NOR2X1 g135731(.A (n_1620), .B (n_725), .Y (n_1684));
INVX1 g135218(.A (n_1683), .Y (n_1705));
NAND3X1 g135018(.A (n_1682), .B (n_457), .C (n_1681), .Y (n_2524));
NOR2X1 g135689(.A (n_844), .B (n_1523), .Y (n_1680));
NAND2X1 g135908(.A (n_10562), .B (P2_n_749), .Y (n_12964));
NOR2X1 g135067(.A (n_403), .B (n_1534), .Y (n_2206));
CLKBUFX1 g136974(.A (n_1677), .Y (n_31912));
OAI21X1 g135210(.A0 (n_1546), .A1 (n_1563), .B0 (n_1675), .Y(n_2216));
NAND2X1 g135849(.A (P2_reg3[1] ), .B (P2_n_749), .Y (n_12968));
NAND2X1 g135713(.A (n_922), .B (n_1393), .Y (n_1672));
NOR2X1 g135554(.A (n_1671), .B (n_1739), .Y (n_2115));
INVX1 g135286(.A (n_1669), .Y (n_1670));
NAND2X1 g135402(.A (n_1667), .B (n_927), .Y (n_1668));
NAND2X1 g136028(.A (P2_reg3[15] ), .B (n_1619), .Y (n_12879));
NAND3X1 g135552(.A (n_1104), .B (n_1666), .C (n_439), .Y (n_1757));
CLKBUFX1 g136975(.A (n_1677), .Y (n_31201));
NOR2X1 g135108(.A (n_1692), .B (n_1663), .Y (n_1664));
NAND2X1 g135984(.A (n_1661), .B (n_33579), .Y (n_1662));
OAI21X1 g134644(.A0 (n_706), .A1 (n_1190), .B0 (n_1667), .Y (n_2478));
INVX2 g137168(.A (n_4371), .Y (n_1659));
AND2X1 g135750(.A (n_780), .B (n_2173), .Y (n_4639));
AND2X1 g135025(.A (n_2844), .B (n_1658), .Y (n_3283));
AND2X1 g135531(.A (n_825), .B (n_1556), .Y (n_1657));
NAND2X1 g135638(.A (n_1615), .B (n_598), .Y (n_2440));
NOR2X1 g135719(.A (n_1385), .B (n_744), .Y (n_1655));
AOI21X1 g134649(.A0 (n_1453), .A1 (n_1654), .B0 (n_1653), .Y(n_1841));
NOR2X1 g135486(.A (n_1555), .B (n_1221), .Y (n_2074));
NOR2X1 g135350(.A (n_1652), .B (n_1651), .Y (n_2122));
NAND2X1 g135695(.A (n_794), .B (n_1654), .Y (n_1648));
NAND2X1 g135915(.A (n_1646), .B (n_1645), .Y (n_1647));
AOI21X1 g135254(.A0 (n_1234), .A1 (n_1230), .B0 (n_1527), .Y(n_2683));
INVX1 g135639(.A (n_1643), .Y (n_1644));
AOI21X1 g135763(.A0 (datao_1[0] ), .A1 (n_144), .B0 (n_2598), .Y(n_1642));
NOR2X1 g135401(.A (n_1899), .B (n_1640), .Y (n_1641));
NOR2X1 g135633(.A (n_806), .B (n_767), .Y (n_2031));
NOR2X1 g135611(.A (n_1639), .B (n_2141), .Y (n_2231));
INVX1 g137072(.A (n_34700), .Y (n_29285));
AND2X1 g135311(.A (n_934), .B (n_1345), .Y (n_1634));
INVX1 g137089(.A (n_1633), .Y (n_31534));
AND2X1 g135075(.A (n_2077), .B (n_1632), .Y (n_4037));
NAND2X1 g135742(.A (n_1630), .B (n_1629), .Y (n_2009));
NAND2X1 g134698(.A (n_1626), .B (n_10838), .Y (n_3534));
NAND2X1 g135842(.A (n_1624), .B (n_1407), .Y (n_1625));
INVX1 g135542(.A (n_1622), .Y (n_1623));
INVX1 g137095(.A (n_31493), .Y (n_1621));
NOR2X1 g135711(.A (n_2055), .B (n_795), .Y (n_3509));
NAND2X1 g136422(.A (addr_446), .B (n_482), .Y (n_2140));
AOI21X1 g135242(.A0 (n_1341), .A1 (n_1189), .B0 (n_1620), .Y(n_2257));
OR2X1 g135417(.A (n_2244), .B (n_962), .Y (n_1709));
NAND2X1 g136016(.A (P2_reg3[13] ), .B (n_1619), .Y (n_12881));
AND2X1 g135021(.A (n_1618), .B (n_1617), .Y (n_2377));
NAND2X1 g135700(.A (n_753), .B (n_1387), .Y (n_1616));
NAND2X1 g135425(.A (n_1615), .B (n_1855), .Y (n_2329));
NAND2X1 g133867(.A (n_1456), .B (P2_reg3[6] ), .Y (n_1614));
NOR2X1 g135734(.A (n_1247), .B (n_937), .Y (n_1611));
INVX1 g135680(.A (n_1956), .Y (n_1610));
NAND2X1 g135011(.A (n_3506), .B (n_1609), .Y (n_1935));
NAND2X1 g135441(.A (n_1821), .B (n_1603), .Y (n_2158));
INVX1 g137008(.A (n_1591), .Y (n_31726));
NOR2X1 g135326(.A (n_1608), .B (n_1607), .Y (n_2133));
NAND2X1 g135370(.A (n_1759), .B (n_1605), .Y (n_2527));
NAND2X1 g135468(.A (n_1604), .B (n_1603), .Y (n_2263));
NOR2X1 g135595(.A (n_1026), .B (n_1547), .Y (n_1602));
INVX1 g137120(.A (n_34309), .Y (n_31328));
INVX1 g137033(.A (n_31592), .Y (n_2070));
INVX1 g137119(.A (n_34309), .Y (n_27698));
NAND2X1 g135920(.A (P2_reg3[5] ), .B (n_1619), .Y (n_12877));
NAND2X1 g135982(.A (P2_reg3[10] ), .B (n_1619), .Y (n_12896));
NOR2X1 g135589(.A (n_2141), .B (n_2118), .Y (n_2298));
CLKBUFX1 g136993(.A (n_35024), .Y (n_31891));
NOR2X1 g135612(.A (n_1595), .B (n_1639), .Y (n_2200));
INVX1 g137019(.A (n_15981), .Y (n_31105));
NAND2X1 g135470(.A (n_761), .B (n_842), .Y (n_2081));
NOR2X1 g135521(.A (n_963), .B (n_1593), .Y (n_1703));
NAND2X1 g135408(.A (n_2244), .B (n_449), .Y (n_1592));
INVX1 g136980(.A (n_31845), .Y (n_15722));
NAND2X1 g135614(.A (n_1037), .B (n_1002), .Y (n_1933));
INVX1 g137009(.A (n_1591), .Y (n_31538));
OAI21X1 g135211(.A0 (n_1590), .A1 (n_1589), .B0 (n_1588), .Y(n_2346));
NAND2X1 g135359(.A (n_1615), .B (n_1271), .Y (n_2252));
INVX1 g137016(.A (n_1587), .Y (n_31894));
NOR2X1 g135592(.A (n_782), .B (n_1544), .Y (n_1586));
NAND2X1 g135987(.A (P2_reg3[6] ), .B (n_1619), .Y (n_12875));
INVX1 g135625(.A (n_1582), .Y (n_1583));
NAND2X1 g135730(.A (n_862), .B (n_1296), .Y (n_1581));
NOR2X1 g135377(.A (n_571), .B (n_1580), .Y (n_2191));
INVX1 g136435(.A (n_1853), .Y (n_1579));
NAND2X1 g135053(.A (n_1577), .B (n_1576), .Y (n_1578));
NAND2X1 g136012(.A (P1_IR[19] ), .B (n_1645), .Y (n_1575));
NOR2X1 g135644(.A (n_1573), .B (n_1572), .Y (n_2556));
CLKBUFX1 g136982(.A (n_31845), .Y (n_31205));
NOR2X1 g135718(.A (n_1569), .B (n_757), .Y (n_1570));
NOR2X1 g135755(.A (n_832), .B (n_1531), .Y (n_1568));
AND2X1 g134955(.A (n_1566), .B (n_1565), .Y (n_2634));
INVX1 g135736(.A (n_2058), .Y (n_1564));
NOR2X1 g135420(.A (n_1651), .B (n_1563), .Y (n_2187));
NAND2X1 g135637(.A (n_1562), .B (n_846), .Y (n_1987));
INVX1 g135732(.A (n_1746), .Y (n_1561));
NAND2X1 g134981(.A (n_1560), .B (n_1663), .Y (n_2495));
INVX1 g136288(.A (n_2117), .Y (n_1559));
NOR2X1 g135714(.A (n_1542), .B (n_833), .Y (n_1558));
NOR2X1 g135587(.A (n_824), .B (n_973), .Y (n_2185));
NOR2X1 g135564(.A (n_1082), .B (n_1009), .Y (n_2000));
NOR2X1 g135325(.A (n_1136), .B (n_1555), .Y (n_2172));
NOR2X1 g135570(.A (n_897), .B (n_399), .Y (n_2192));
NAND2X1 g135824(.A (P3_IR[21] ), .B (n_1512), .Y (n_1554));
NAND2X1 g135655(.A (n_817), .B (n_479), .Y (n_1553));
AND2X1 g135545(.A (n_1474), .B (n_1552), .Y (n_2179));
NAND2X1 g135726(.A (n_1244), .B (n_1551), .Y (n_2072));
INVX1 g135189(.A (n_1549), .Y (n_1550));
INVX1 g135202(.A (n_2241), .Y (n_1548));
OAI21X1 g135228(.A0 (n_1543), .A1 (n_1547), .B0 (n_1546), .Y(n_2224));
OAI21X1 g135229(.A0 (n_1545), .A1 (n_1544), .B0 (n_1543), .Y(n_2324));
AOI21X1 g135288(.A0 (n_1481), .A1 (n_1352), .B0 (n_1542), .Y(n_2243));
NAND2X1 g135364(.A (n_1316), .B (n_636), .Y (n_2124));
NAND3X1 g135385(.A (n_1541), .B (n_34090), .C (n_607), .Y (n_1825));
NAND2X1 g135430(.A (n_1604), .B (n_1537), .Y (n_2264));
NOR2X1 g135407(.A (n_2286), .B (n_1536), .Y (n_2116));
NOR2X1 g135729(.A (n_1182), .B (n_1040), .Y (n_1535));
NOR2X1 g134930(.A (n_1534), .B (P3_reg3[3] ), .Y (n_2375));
NOR2X1 g135656(.A (n_1368), .B (n_918), .Y (n_1533));
INVX1 g135683(.A (n_1532), .Y (n_3785));
AOI21X1 g135250(.A0 (n_1372), .A1 (n_1531), .B0 (n_1529), .Y(n_2349));
NOR2X1 g135745(.A (n_1394), .B (n_900), .Y (n_1530));
AOI21X1 g135239(.A0 (n_1469), .A1 (n_1529), .B0 (n_1381), .Y(n_2612));
NOR2X1 g135752(.A (n_912), .B (n_1527), .Y (n_1528));
INVX1 g135677(.A (n_1827), .Y (n_1526));
NAND2X1 g133907(.A (n_1524), .B (n_880), .Y (n_1525));
AOI21X1 g135253(.A0 (n_1344), .A1 (n_1527), .B0 (n_1523), .Y(n_2828));
NAND3X1 g134624(.A (n_1522), .B (P1_reg3[7] ), .C (P1_reg3[8] ), .Y(n_2562));
NAND2X1 g135422(.A (n_1125), .B (n_32927), .Y (n_1521));
NOR2X1 g135366(.A (n_1608), .B (n_1739), .Y (n_2312));
NAND2X1 g135931(.A (P1_IR[23] ), .B (n_998), .Y (n_33053));
INVX1 g136996(.A (n_35024), .Y (n_7245));
INVX1 g135663(.A (n_2043), .Y (n_1518));
NAND4X1 g135258(.A (n_1517), .B (P2_reg3[3] ), .C (P2_reg3[5] ), .D(P2_reg3[4] ), .Y (n_1719));
INVX1 g137127(.A (n_3185), .Y (n_31586));
NOR2X1 g135399(.A (n_1516), .B (n_1489), .Y (n_2114));
NAND2X1 g135999(.A (P3_IR[19] ), .B (n_1512), .Y (n_35284));
INVX1 g135661(.A (n_1510), .Y (n_1511));
NOR2X1 g135403(.A (n_940), .B (n_1099), .Y (n_2600));
INVX1 g135669(.A (n_1957), .Y (n_1509));
NAND2X1 g135518(.A (n_1508), .B (n_1555), .Y (n_2079));
INVX1 g137129(.A (n_3185), .Y (n_16415));
NOR2X1 g135410(.A (n_956), .B (n_1573), .Y (n_1504));
AND2X1 g135081(.A (n_1817), .B (n_1658), .Y (n_4024));
INVX1 g135347(.A (n_2589), .Y (n_1503));
AND2X1 g134989(.A (n_1502), .B (n_1501), .Y (n_2065));
NAND3X1 g135054(.A (n_1500), .B (n_1294), .C (n_1499), .Y (n_2757));
NOR2X1 g135607(.A (n_1498), .B (n_1497), .Y (n_2113));
NOR2X1 g135598(.A (n_959), .B (n_1096), .Y (n_2882));
OAI21X1 g135188(.A0 (n_1496), .A1 (n_1119), .B0 (n_1433), .Y(n_1918));
OR2X1 g135682(.A (n_1495), .B (n_918), .Y (n_2094));
NAND2X1 g135097(.A (n_1494), .B (n_1632), .Y (n_1747));
NAND3X1 g134971(.A (n_1491), .B (n_1490), .C (P2_reg3[27] ), .Y(n_1492));
NOR2X1 g135474(.A (n_1536), .B (n_1671), .Y (n_2181));
NOR2X1 g135710(.A (n_833), .B (n_1551), .Y (n_1907));
INVX1 g137133(.A (n_1812), .Y (n_31588));
NAND2X1 g135496(.A (n_1605), .B (n_1489), .Y (n_2131));
NOR2X1 g135519(.A (n_1488), .B (n_1652), .Y (n_2183));
NOR2X1 g135550(.A (n_1537), .B (n_1420), .Y (n_2190));
OR2X1 g136538(.A (n_150), .B (n_1486), .Y (n_1487));
AND2X1 g136210(.A (P2_reg3[1] ), .B (n_34309), .Y (n_1485));
INVX1 g134843(.A (n_1300), .Y (n_1484));
INVX1 g136991(.A (n_15723), .Y (n_2174));
NOR2X1 g135716(.A (n_1481), .B (n_758), .Y (n_1482));
NAND2X1 g135600(.A (n_1143), .B (n_497), .Y (n_2012));
AND2X1 g135485(.A (n_1479), .B (n_1838), .Y (n_1480));
NOR2X1 g135489(.A (n_925), .B (n_1477), .Y (n_1478));
NAND2X1 g135571(.A (n_1615), .B (n_1474), .Y (n_1475));
OR2X1 g135902(.A (n_367), .B (n_33815), .Y (n_1473));
INVX1 g137069(.A (n_34700), .Y (n_31149));
NAND2X1 g134952(.A (n_1471), .B (n_2101), .Y (n_2516));
OR2X1 g135739(.A (n_725), .B (n_1551), .Y (n_2150));
NAND2X1 g135688(.A (n_796), .B (n_1469), .Y (n_1470));
NAND2X1 g135787(.A (P2_reg3[7] ), .B (n_1619), .Y (n_12890));
NAND2X1 g135762(.A (n_787), .B (n_1006), .Y (n_7734));
NOR2X1 g135536(.A (n_1640), .B (n_1468), .Y (n_2219));
AND2X1 g134973(.A (n_1701), .B (n_1560), .Y (n_1467));
NOR2X1 g135537(.A (n_1498), .B (n_1135), .Y (n_1466));
XOR2X1 g134673(.A (n_339), .B (n_1007), .Y (n_1911));
NOR2X1 g135558(.A (n_1748), .B (n_2989), .Y (n_2282));
NAND2X1 g135304(.A (n_1464), .B (n_731), .Y (n_1465));
NOR2X1 g135619(.A (n_1468), .B (n_1488), .Y (n_2333));
NAND3X1 g135146(.A (n_1462), .B (n_972), .C (n_1461), .Y (n_1868));
AND2X1 g135043(.A (n_1694), .B (n_1663), .Y (n_2296));
NAND3X1 g135073(.A (n_1459), .B (n_544), .C (P1_reg3[27] ), .Y(n_1460));
INVX1 g135862(.A (n_1863), .Y (n_1458));
OR2X1 g133850(.A (n_1456), .B (P2_reg3[6] ), .Y (n_1457));
OR2X1 g135859(.A (n_622), .B (n_852), .Y (n_1455));
NAND3X1 g135353(.A (n_947), .B (n_739), .C (n_345), .Y (n_1856));
NAND3X1 g134853(.A (n_1453), .B (n_2066), .C (n_1654), .Y (n_1454));
INVX1 g135100(.A (n_1673), .Y (n_1451));
INVX1 g135321(.A (n_1449), .Y (n_1450));
NAND2X1 g136540(.A (si[17]), .B (n_475), .Y (n_2186));
INVX1 g135790(.A (n_1936), .Y (n_1448));
INVX1 g135671(.A (n_1447), .Y (n_2057));
NOR2X1 g135744(.A (n_1380), .B (n_1047), .Y (n_1446));
NAND3X1 g134947(.A (n_1325), .B (n_688), .C (n_982), .Y (n_1874));
NOR2X1 g135596(.A (n_1537), .B (n_1580), .Y (n_2582));
INVX1 g137138(.A (n_31328), .Y (n_31345));
INVX1 g137111(.A (n_1336), .Y (n_31647));
OR2X1 g135597(.A (n_986), .B (n_1444), .Y (n_1445));
INVX1 g135458(.A (n_1439), .Y (n_1440));
NAND2X1 g134963(.A (n_2059), .B (n_1438), .Y (n_2841));
NOR2X1 g135113(.A (n_1402), .B (n_1437), .Y (n_1971));
INVX1 g135561(.A (n_1435), .Y (n_1436));
NAND2X1 g135107(.A (n_1438), .B (n_1963), .Y (n_2480));
NOR2X1 g135479(.A (n_1433), .B (n_1177), .Y (n_1434));
NAND2X1 g135115(.A (n_2393), .B (n_1431), .Y (n_1432));
CLKBUFX1 g136976(.A (n_1677), .Y (n_31641));
AND2X1 g135105(.A (n_1428), .B (n_1427), .Y (n_1429));
NOR2X1 g134945(.A (n_1632), .B (n_1425), .Y (n_1426));
NAND3X1 g134921(.A (n_34090), .B (n_367), .C (n_1089), .Y (n_1733));
OR2X1 g135793(.A (n_727), .B (n_1423), .Y (n_1424));
CLKBUFX1 g137102(.A (n_1313), .Y (n_31528));
INVX1 g135515(.A (n_1421), .Y (n_1422));
NAND2X1 g135127(.A (n_1996), .B (n_1945), .Y (n_1902));
NOR2X1 g135464(.A (n_1420), .B (n_1419), .Y (n_2098));
NAND2X1 g135333(.A (n_2148), .B (n_1854), .Y (n_1418));
AND2X1 g134972(.A (n_1416), .B (n_1425), .Y (n_1417));
NOR2X1 g134910(.A (n_895), .B (P3_reg3[5] ), .Y (n_1879));
NOR2X1 g135492(.A (n_476), .B (n_1489), .Y (n_1415));
NAND2X1 g135833(.A (P3_IR[22] ), .B (n_1512), .Y (n_35336));
NAND2X1 g135668(.A (n_1343), .B (n_851), .Y (n_1413));
INVX1 g135525(.A (n_1411), .Y (n_1412));
CLKBUFX1 g137103(.A (n_1313), .Y (n_31965));
INVX1 g137124(.A (n_1409), .Y (n_30968));
NAND2X1 g135841(.A (P2_IR[15] ), .B (n_1407), .Y (n_32580));
NOR2X1 g135584(.A (n_1572), .B (n_1595), .Y (n_3221));
NAND2X1 g135860(.A (n_516), .B (n_1407), .Y (n_1405));
NOR2X1 g135675(.A (n_1529), .B (n_902), .Y (n_1403));
OR2X1 g134713(.A (n_2226), .B (n_1402), .Y (n_2137));
NAND2X1 g135707(.A (n_1268), .B (n_1495), .Y (n_2578));
NAND3X1 g134940(.A (n_1401), .B (n_211), .C (n_1359), .Y (n_1728));
NOR2X1 g135060(.A (n_1427), .B (n_1399), .Y (n_1400));
NOR2X1 g134965(.A (n_2336), .B (n_1438), .Y (n_1398));
INVX1 g135355(.A (n_1396), .Y (n_1397));
AOI21X1 g135240(.A0 (n_1394), .A1 (n_1393), .B0 (n_1388), .Y(n_2170));
INVX1 g135299(.A (n_34537), .Y (n_1860));
AND2X1 g135367(.A (n_908), .B (n_1101), .Y (n_1391));
NAND2X1 g135318(.A (n_33351), .B (n_1562), .Y (n_1845));
NAND2X1 g135944(.A (P2_reg3[11] ), .B (n_1619), .Y (n_12892));
AOI21X1 g135252(.A0 (n_1388), .A1 (n_1387), .B0 (n_1243), .Y(n_2931));
INVX1 g135724(.A (n_1785), .Y (n_1386));
AOI21X1 g135243(.A0 (n_1620), .A1 (n_1217), .B0 (n_1385), .Y(n_2494));
NOR2X1 g135061(.A (n_773), .B (P1_IR[29] ), .Y (n_1382));
AOI21X1 g135236(.A0 (n_1381), .A1 (n_1361), .B0 (n_1380), .Y(n_2348));
CLKBUFX1 g136977(.A (n_1677), .Y (n_31933));
INVX1 g136990(.A (n_15723), .Y (n_2091));
NAND2X1 g136083(.A (n_628), .B (addr_441), .Y (n_1993));
AND2X1 g135346(.A (n_1552), .B (n_1855), .Y (n_1379));
OR2X1 g135223(.A (n_926), .B (n_1477), .Y (n_2053));
NOR2X1 g135499(.A (n_1419), .B (n_1516), .Y (n_2119));
NOR2X1 g135586(.A (n_1489), .B (n_1497), .Y (n_2229));
NOR2X1 g135648(.A (n_840), .B (n_1563), .Y (n_1378));
NAND2X1 g135925(.A (P2_IR[19] ), .B (n_1486), .Y (n_1377));
NOR2X1 g135475(.A (n_1375), .B (n_2286), .Y (n_2182));
NOR2X1 g135577(.A (n_1374), .B (n_1373), .Y (n_1782));
AND2X1 g135622(.A (n_2989), .B (n_611), .Y (n_4853));
INVX1 g136984(.A (n_1677), .Y (n_30702));
NAND2X1 g136102(.A (si[18]), .B (n_693), .Y (n_2327));
NAND2X1 g135510(.A (n_951), .B (n_870), .Y (n_1762));
INVX1 g137132(.A (n_1812), .Y (n_31644));
AND2X1 g135130(.A (n_1471), .B (n_1609), .Y (n_4334));
CLKBUFX1 g137105(.A (n_1313), .Y (n_31677));
NAND2X1 g135746(.A (n_1469), .B (n_1372), .Y (n_1937));
XOR2X1 g134685(.A (n_830), .B (n_831), .Y (n_13167));
INVX1 g136186(.A (n_1488), .Y (n_1371));
NAND2X1 g136271(.A (n_130), .B (addr_425), .Y (n_1864));
NOR2X1 g135594(.A (n_1363), .B (n_1330), .Y (n_1962));
NAND2X1 g135293(.A (n_595), .B (n_1369), .Y (n_1370));
NOR2X1 g135665(.A (n_1368), .B (n_1385), .Y (n_1793));
AND2X1 g135898(.A (n_150), .B (n_1203), .Y (n_1367));
CLKBUFX1 g137094(.A (n_31097), .Y (n_31683));
AOI22X1 g135287(.A0 (n_1364), .A1 (n_734), .B0 (n_1365), .B1(n_1364), .Y (n_1669));
NAND2X1 g135624(.A (n_997), .B (n_1363), .Y (n_1998));
NAND2X1 g135324(.A (n_1364), .B (n_1750), .Y (n_1362));
NAND2X1 g135723(.A (n_1361), .B (n_1283), .Y (n_1942));
AND2X1 g135472(.A (n_1359), .B (n_1106), .Y (n_1360));
OAI21X1 g135190(.A0 (n_1357), .A1 (n_1222), .B0 (n_1356), .Y(n_1549));
INVX1 g136983(.A (n_34676), .Y (n_31845));
INVX1 g135603(.A (n_1566), .Y (n_1355));
OAI21X1 g135227(.A0 (n_1276), .A1 (n_855), .B0 (n_1256), .Y (n_2162));
AND2X1 g135702(.A (n_1353), .B (n_2303), .Y (n_1354));
AND2X1 g135439(.A (n_1142), .B (n_1315), .Y (n_2125));
INVX1 g137017(.A (n_15981), .Y (n_1587));
NAND2X1 g135720(.A (n_1352), .B (n_1282), .Y (n_2097));
OR2X1 g135918(.A (n_32397), .B (n_609), .Y (n_1351));
AND2X1 g135605(.A (n_1270), .B (n_1474), .Y (n_2289));
INVX1 g136304(.A (n_1433), .Y (n_1350));
NOR2X1 g135667(.A (n_1394), .B (n_1569), .Y (n_1828));
NOR2X1 g135749(.A (n_1314), .B (n_1523), .Y (n_1766));
OR2X1 g135766(.A (n_592), .B (n_554), .Y (n_1347));
INVX1 g137136(.A (n_34309), .Y (n_16150));
OAI21X1 g135198(.A0 (n_1331), .A1 (n_1224), .B0 (n_889), .Y (n_2126));
INVX1 g136354(.A (n_1345), .Y (n_1346));
NOR2X1 g135601(.A (n_760), .B (n_1069), .Y (n_1955));
NAND2X1 g135672(.A (n_1344), .B (n_1343), .Y (n_1447));
OR2X1 g135748(.A (n_1542), .B (n_1341), .Y (n_2071));
NOR2X1 g136402(.A (n_1094), .B (n_998), .Y (n_1340));
NAND2X1 g135543(.A (n_805), .B (n_1022), .Y (n_1622));
AND2X1 g135368(.A (n_708), .B (n_1576), .Y (n_1339));
INVX1 g135432(.A (n_1399), .Y (n_1383));
AND2X1 g136511(.A (n_32938), .B (n_1724), .Y (n_1338));
INVX1 g137108(.A (n_1313), .Y (n_1336));
OR2X1 g135691(.A (n_2055), .B (n_1916), .Y (n_1334));
INVX1 g136409(.A (n_1604), .Y (n_1333));
AND2X1 g135535(.A (n_584), .B (n_604), .Y (n_2147));
NAND2X1 g135979(.A (P3_reg3[28] ), .B (n_7390), .Y (n_1332));
OAI21X1 g135231(.A0 (n_1048), .A1 (n_1265), .B0 (n_1331), .Y(n_2422));
NOR2X1 g135378(.A (n_1330), .B (n_1266), .Y (n_1831));
NAND2X1 g135791(.A (n_116), .B (datao_1[28] ), .Y (n_1936));
INVX1 g136700(.A (n_1292), .Y (n_31958));
NOR2X1 g135427(.A (n_1363), .B (n_1299), .Y (n_1808));
AND2X1 g135628(.A (n_1952), .B (n_1328), .Y (n_1329));
NOR2X1 g135618(.A (n_1327), .B (n_2118), .Y (n_2230));
INVX1 g135329(.A (n_1325), .Y (n_1326));
OR2X1 g135858(.A (n_1323), .B (P3_IR[31] ), .Y (n_1324));
INVX1 g136411(.A (n_1651), .Y (n_1321));
INVX1 g135342(.A (n_1320), .Y (n_2376));
NAND3X1 g135685(.A (n_620), .B (P2_reg3[12] ), .C (n_1319), .Y(n_1771));
INVX1 g137079(.A (n_1409), .Y (n_31343));
INVX1 g137078(.A (n_1409), .Y (n_15477));
NAND2X1 g135328(.A (n_1316), .B (n_1315), .Y (n_1317));
NOR2X1 g135666(.A (n_1343), .B (n_1314), .Y (n_2364));
INVX1 g137090(.A (n_3185), .Y (n_1633));
AND2X1 g135681(.A (n_1343), .B (n_1195), .Y (n_1956));
NAND2X1 g135409(.A (n_1163), .B (n_584), .Y (n_1312));
NAND2X1 g135733(.A (n_1393), .B (n_1387), .Y (n_1746));
INVX1 g135567(.A (n_1310), .Y (n_1311));
OR2X1 g136022(.A (n_799), .B (n_609), .Y (n_1309));
INVX1 g135361(.A (n_1307), .Y (n_1308));
NOR2X1 g135348(.A (n_639), .B (n_1085), .Y (n_2589));
INVX1 g136978(.A (n_34676), .Y (n_1677));
NOR2X1 g135626(.A (n_1150), .B (n_915), .Y (n_1582));
AND2X1 g135820(.A (n_1304), .B (n_33815), .Y (n_1305));
NOR2X1 g135803(.A (n_138), .B (datao_2[25] ), .Y (n_2178));
NOR2X1 g135480(.A (n_395), .B (n_849), .Y (n_1303));
INVX1 g136506(.A (n_1536), .Y (n_1302));
OAI21X1 g135183(.A0 (n_1299), .A1 (n_1273), .B0 (n_1197), .Y(n_2004));
NAND2X1 g135436(.A (n_550), .B (n_1297), .Y (n_1298));
NAND2X1 g135694(.A (n_1246), .B (n_1296), .Y (n_2052));
NOR2X1 g135572(.A (n_409), .B (n_1199), .Y (n_2951));
INVX1 g135395(.A (n_1494), .Y (n_1627));
AND2X1 g135400(.A (n_981), .B (n_1294), .Y (n_2255));
INVX1 g136264(.A (n_1595), .Y (n_1290));
NAND2X1 g135557(.A (n_1590), .B (n_435), .Y (n_1287));
NOR2X1 g135476(.A (n_454), .B (n_869), .Y (n_2064));
NAND2X1 g135873(.A (P3_IR[14] ), .B (n_3196), .Y (n_32016));
INVX1 g136261(.A (n_1552), .Y (n_1284));
NAND2X1 g135706(.A (n_1283), .B (n_1282), .Y (n_2237));
NAND2X1 g135921(.A (P1_IR[11] ), .B (n_1277), .Y (n_1279));
NAND2X1 g135880(.A (datao_1[30] ), .B (n_380), .Y (n_1959));
OAI21X1 g134641(.A0 (n_707), .A1 (n_854), .B0 (n_1276), .Y (n_3022));
NAND2X1 g135922(.A (n_1274), .B (n_3705), .Y (n_1275));
OAI21X1 g135191(.A0 (n_1209), .A1 (n_1041), .B0 (n_1273), .Y(n_2351));
NAND2X1 g136193(.A (si[13]), .B (n_12030), .Y (n_1901));
NAND2X1 g135406(.A (n_1271), .B (n_1270), .Y (n_1272));
NOR2X1 g135698(.A (n_1314), .B (n_1531), .Y (n_1789));
NAND2X1 g135948(.A (P3_IR[12] ), .B (n_33566), .Y (n_1267));
OAI21X1 g135208(.A0 (n_1266), .A1 (n_1141), .B0 (n_1265), .Y(n_2063));
AND2X1 g135919(.A (n_1253), .B (n_852), .Y (n_1264));
NOR2X1 g135658(.A (n_1263), .B (n_1368), .Y (n_2037));
OR2X1 g135448(.A (n_679), .B (n_1363), .Y (n_1262));
NOR2X1 g135356(.A (n_950), .B (n_1261), .Y (n_1396));
NAND2X1 g135602(.A (n_1928), .B (n_1259), .Y (n_1260));
NAND2X1 g135617(.A (n_1331), .B (n_579), .Y (n_1258));
AND2X1 g135341(.A (n_1256), .B (n_1255), .Y (n_1257));
INVX1 g137010(.A (n_2091), .Y (n_1591));
OR2X1 g136249(.A (n_1253), .B (n_33587), .Y (n_1254));
NAND2X1 g135728(.A (n_1250), .B (n_1249), .Y (n_1251));
NOR2X1 g135676(.A (n_1481), .B (n_1282), .Y (n_1797));
NAND2X1 g135560(.A (n_414), .B (n_1273), .Y (n_1248));
NOR2X1 g135715(.A (n_1247), .B (n_1246), .Y (n_1977));
NOR2X1 g135657(.A (n_1243), .B (n_1247), .Y (n_2041));
INVX1 g136215(.A (n_1373), .Y (n_1612));
INVX1 g135565(.A (n_1240), .Y (n_1241));
OR2X1 g136495(.A (n_590), .B (n_33587), .Y (n_1239));
NAND3X1 g135747(.A (n_1238), .B (P2_reg3[10] ), .C (P2_reg3[7] ),.Y (n_1836));
OR2X1 g135705(.A (n_1394), .B (n_1233), .Y (n_2310));
INVX1 g137082(.A (n_33194), .Y (n_12969));
NAND2X1 g135701(.A (n_1469), .B (n_1361), .Y (n_1973));
OR2X1 g135911(.A (n_1236), .B (n_34946), .Y (n_1237));
NOR2X1 g135360(.A (n_599), .B (n_1420), .Y (n_1235));
NOR2X1 g135703(.A (n_1247), .B (n_1234), .Y (n_2044));
NAND2X1 g135932(.A (n_13675), .B (n_3964), .Y (n_13196));
NAND2X1 g135679(.A (n_1233), .B (n_1232), .Y (n_1827));
NOR2X1 g135322(.A (n_34409), .B (n_34528), .Y (n_1449));
INVX1 g136419(.A (n_1640), .Y (n_1231));
AND2X1 g135737(.A (n_1296), .B (n_1230), .Y (n_2058));
OR2X1 g135956(.A (n_1253), .B (n_33815), .Y (n_1229));
AND2X1 g136389(.A (n_1227), .B (n_1724), .Y (n_1228));
NAND3X1 g134982(.A (P2_reg3[11] ), .B (P2_reg3[12] ), .C (n_634),.Y (n_2196));
NAND2X1 g135653(.A (n_1079), .B (n_619), .Y (n_1226));
NOR2X1 g135379(.A (n_400), .B (n_1224), .Y (n_1225));
CLKBUFX1 g137109(.A (n_1313), .Y (n_31594));
NAND2X1 g135792(.A (P3_reg3[7] ), .B (n_3964), .Y (n_12999));
OAI21X1 g135199(.A0 (n_1223), .A1 (n_663), .B0 (n_1222), .Y (n_2228));
OAI21X1 g135235(.A0 (n_1508), .A1 (n_1221), .B0 (n_1080), .Y(n_2611));
NAND2X1 g135305(.A (n_366), .B (n_1090), .Y (n_1220));
NAND2X1 g135690(.A (n_1167), .B (n_1217), .Y (n_2151));
INVX1 g137023(.A (n_31105), .Y (n_3217));
INVX1 g135620(.A (n_1214), .Y (n_1215));
AND2X1 g136013(.A (datao_1[24] ), .B (n_171), .Y (n_1966));
NAND2X1 g135712(.A (n_1387), .B (n_1246), .Y (n_2169));
NAND2X1 g135673(.A (n_2303), .B (n_1958), .Y (n_1213));
NAND2X1 g135903(.A (n_1211), .B (n_3196), .Y (n_1212));
AND2X1 g135386(.A (n_1209), .B (n_397), .Y (n_1210));
NOR2X1 g135652(.A (n_640), .B (n_1162), .Y (n_1208));
OR2X1 g135971(.A (n_1206), .B (n_609), .Y (n_1207));
OR2X1 g135958(.A (n_287), .B (n_1203), .Y (n_1204));
INVX1 g136415(.A (n_1593), .Y (n_1202));
NOR2X1 g135457(.A (n_1958), .B (datao_1[30] ), .Y (n_1200));
NOR2X1 g135526(.A (n_683), .B (n_1199), .Y (n_1411));
NAND2X1 g135590(.A (n_1197), .B (n_513), .Y (n_1198));
NOR2X1 g135316(.A (n_489), .B (n_1001), .Y (n_2048));
INVX1 g137125(.A (P2_n_749), .Y (n_1409));
NOR2X1 g135863(.A (n_294), .B (datao_2[2] ), .Y (n_1863));
NAND2X1 g135674(.A (n_1195), .B (n_1372), .Y (n_1767));
INVX1 g136493(.A (n_1419), .Y (n_1194));
NAND2X1 g135438(.A (n_670), .B (n_955), .Y (n_1193));
NAND2X1 g135846(.A (P1_IR[22] ), .B (n_1277), .Y (n_32216));
CLKBUFX1 g137170(.A (n_1423), .Y (n_4371));
NAND3X1 g135753(.A (n_989), .B (P1_reg3[12] ), .C (P1_reg3[9] ), .Y(n_1805));
NOR2X1 g135642(.A (n_1327), .B (n_1190), .Y (n_2250));
NAND2X1 g135684(.A (n_1250), .B (n_2173), .Y (n_1532));
NAND2X1 g135985(.A (P3_reg3[2] ), .B (n_3964), .Y (n_13194));
AND2X1 g135664(.A (n_1217), .B (n_1189), .Y (n_2043));
AND2X1 g135670(.A (n_1344), .B (n_1230), .Y (n_1957));
NOR2X1 g135609(.A (n_34852), .B (n_1149), .Y (n_2670));
NOR2X1 g135516(.A (n_1075), .B (n_1199), .Y (n_1421));
NOR2X1 g135640(.A (n_1097), .B (n_1098), .Y (n_1643));
NAND2X1 g135635(.A (n_2035), .B (n_538), .Y (n_1185));
NOR2X1 g135380(.A (n_1223), .B (n_1052), .Y (n_4635));
NOR2X1 g135424(.A (n_1221), .B (n_665), .Y (n_1184));
NOR2X1 g135660(.A (n_1380), .B (n_1182), .Y (n_1931));
NOR2X1 g135687(.A (n_1481), .B (n_1182), .Y (n_1924));
NOR2X1 g135469(.A (n_1165), .B (n_546), .Y (n_2381));
NAND2X1 g135704(.A (n_2066), .B (n_1232), .Y (n_1807));
INVX1 g136290(.A (n_1939), .Y (n_1179));
AND2X1 g135484(.A (n_1259), .B (n_1838), .Y (n_1178));
NOR2X1 g135548(.A (n_2146), .B (n_1177), .Y (n_4322));
OAI21X1 g135192(.A0 (n_1256), .A1 (n_829), .B0 (n_1087), .Y (n_2047));
OR2X1 g135810(.A (n_1171), .B (n_609), .Y (n_1172));
INVX1 g134385(.A (n_1456), .Y (n_1169));
INVX1 g136173(.A (n_1497), .Y (n_1168));
NOR2X1 g135743(.A (n_1368), .B (n_1167), .Y (n_1794));
NOR2X1 g135497(.A (n_1166), .B (n_1165), .Y (n_1949));
NOR2X1 g135735(.A (n_1182), .B (n_1283), .Y (n_1932));
INVX1 g137034(.A (n_15968), .Y (n_31592));
INVX1 g135314(.A (n_1913), .Y (n_1164));
OR2X1 g135562(.A (n_992), .B (n_635), .Y (n_1435));
OAI21X1 g135201(.A0 (n_1163), .A1 (n_1162), .B0 (n_1066), .Y(n_2046));
INVX1 g137117(.A (P2_n_749), .Y (n_15864));
INVX1 g137134(.A (n_34309), .Y (n_1812));
INVX1 g136286(.A (n_1639), .Y (n_1160));
NAND2X1 g136289(.A (n_233), .B (addr_426), .Y (n_2117));
INVX1 g136333(.A (n_1866), .Y (n_1159));
INVX1 g137113(.A (n_1313), .Y (n_3834));
INVX1 g135615(.A (n_4341), .Y (n_1158));
INVX1 g136347(.A (n_1607), .Y (n_1157));
OR2X1 g135959(.A (n_590), .B (n_826), .Y (n_1156));
NOR2X1 g135504(.A (n_1036), .B (n_845), .Y (n_2233));
INVX1 g136273(.A (n_33436), .Y (n_35637));
INVX1 g136184(.A (n_1555), .Y (n_1154));
AND2X1 g135717(.A (n_1916), .B (n_1250), .Y (n_5190));
NOR2X1 g136360(.A (n_72), .B (n_7390), .Y (n_1153));
INVX1 g136702(.A (n_1292), .Y (n_13197));
NOR2X1 g135449(.A (n_1544), .B (n_1573), .Y (n_2419));
NOR2X1 g135500(.A (n_1150), .B (n_1149), .Y (n_2209));
AND2X1 g135443(.A (n_708), .B (n_611), .Y (n_1944));
AND2X1 g135426(.A (n_1112), .B (n_1121), .Y (n_1148));
INVX1 g137085(.A (n_15484), .Y (n_15480));
NAND2X1 g135721(.A (n_1393), .B (n_1233), .Y (n_1881));
INVX1 g135374(.A (n_1778), .Y (n_1145));
NAND2X1 g135393(.A (n_1143), .B (n_1142), .Y (n_1144));
NAND2X1 g135327(.A (n_1330), .B (n_1141), .Y (n_1699));
NAND2X1 g135503(.A (n_1276), .B (n_1139), .Y (n_1140));
NOR2X1 g135632(.A (n_1045), .B (n_1374), .Y (n_4938));
NOR2X1 g135419(.A (n_477), .B (n_1136), .Y (n_1137));
OAI21X1 g134642(.A0 (n_430), .A1 (n_1135), .B0 (n_1134), .Y (n_3324));
NAND3X1 g135102(.A (P1_reg3[11] ), .B (P1_reg3[12] ), .C (n_774),.Y (n_1673));
OR2X1 g136284(.A (n_32397), .B (n_998), .Y (n_1133));
INVX1 g136148(.A (n_1588), .Y (n_1132));
INVX1 g134851(.A (n_1522), .Y (n_1897));
XOR2X1 g135772(.A (si[0]), .B (n_144), .Y (n_1131));
INVX1 g136190(.A (n_1125), .Y (n_1126));
INVX1 g136812(.A (n_998), .Y (n_1124));
AND2X1 g135296(.A (n_545), .B (n_1121), .Y (n_1123));
NAND2X1 g135511(.A (n_685), .B (n_1119), .Y (n_1120));
NOR2X1 g135553(.A (n_801), .B (n_458), .Y (n_2408));
NOR2X1 g135738(.A (n_1195), .B (n_1531), .Y (n_2268));
OR2X1 g135983(.A (n_488), .B (n_609), .Y (n_1117));
INVX1 g136123(.A (n_1468), .Y (n_1115));
INVX1 g136381(.A (n_1652), .Y (n_1114));
NAND2X1 g135295(.A (n_1369), .B (n_1112), .Y (n_1113));
NOR2X1 g135434(.A (n_921), .B (n_406), .Y (n_2486));
INVX1 g136699(.A (n_1292), .Y (n_31569));
NAND2X1 g135415(.A (n_1134), .B (n_1110), .Y (n_1111));
NAND2X1 g135821(.A (P3_reg3[0] ), .B (n_3964), .Y (n_13189));
NAND2X1 g135291(.A (n_1107), .B (n_1106), .Y (n_1108));
CLKBUFX1 g137096(.A (n_31097), .Y (n_31493));
INVX1 g136458(.A (n_1101), .Y (n_1102));
INVX1 g136366(.A (n_1516), .Y (n_1100));
AOI21X1 g134912(.A0 (n_237), .A1 (P3_reg3[3] ), .B0 (P3_reg3[4] ),.Y (n_1688));
INVX1 g136454(.A (n_1498), .Y (n_1737));
OR2X1 g135808(.A (n_1094), .B (n_762), .Y (n_1095));
CLKBUFX1 g137093(.A (n_31097), .Y (n_31590));
NOR2X1 g135725(.A (n_1044), .B (n_1495), .Y (n_1785));
INVX1 g136327(.A (n_1572), .Y (n_1093));
INVX1 g135450(.A (n_1173), .Y (n_1092));
AND2X1 g135418(.A (n_1090), .B (n_1089), .Y (n_1091));
NAND2X1 g135397(.A (n_1087), .B (n_604), .Y (n_1088));
NOR2X1 g135528(.A (n_1085), .B (n_1074), .Y (n_2628));
INVX1 g135477(.A (n_1029), .Y (n_1083));
NOR2X1 g135373(.A (n_1082), .B (n_1042), .Y (n_2135));
NOR2X1 g136128(.A (n_1787), .B (n_21), .Y (n_2011));
OR2X1 g135662(.A (n_1234), .B (n_1296), .Y (n_1510));
NOR2X1 g135471(.A (n_390), .B (n_1357), .Y (n_5195));
NOR2X1 g135335(.A (n_572), .B (n_1065), .Y (n_1081));
OAI21X1 g135219(.A0 (n_979), .A1 (n_1080), .B0 (n_1079), .Y (n_1683));
AND2X1 g135530(.A (n_1365), .B (n_1749), .Y (n_1078));
NOR2X1 g135540(.A (n_1547), .B (n_1544), .Y (n_2423));
NAND2X1 g135307(.A (n_652), .B (n_366), .Y (n_1076));
NOR2X1 g135459(.A (n_1075), .B (n_1074), .Y (n_1439));
NOR2X1 g135382(.A (n_463), .B (n_1266), .Y (n_1073));
OR2X1 g135852(.A (n_345), .B (n_762), .Y (n_1072));
NAND2X1 g136436(.A (n_415), .B (n_680), .Y (n_1853));
INVX1 g135767(.A (n_828), .Y (n_1070));
INVX1 g137015(.A (n_15981), .Y (n_30783));
NOR2X1 g135354(.A (n_440), .B (n_1069), .Y (n_2194));
INVX1 g136395(.A (n_1671), .Y (n_1068));
NOR2X1 g135339(.A (n_1330), .B (n_394), .Y (n_1067));
OAI21X1 g135234(.A0 (n_1066), .A1 (n_1065), .B0 (n_949), .Y (n_2221));
NOR2X1 g136223(.A (n_34544), .B (n_33566), .Y (n_1064));
AND2X1 g135659(.A (n_1630), .B (n_2173), .Y (n_2992));
OR2X1 g135454(.A (n_679), .B (n_394), .Y (n_1823));
NOR2X1 g135461(.A (n_1547), .B (n_1563), .Y (n_2069));
INVX1 g136242(.A (n_1608), .Y (n_1061));
NAND3X1 g135727(.A (n_814), .B (P1_reg3[10] ), .C (P1_reg3[7] ), .Y(n_1898));
INVX1 g135283(.A (n_1183), .Y (n_1058));
NOR2X1 g135517(.A (n_539), .B (n_720), .Y (n_3613));
OAI21X1 g135203(.A0 (n_571), .A1 (n_1297), .B0 (n_1271), .Y (n_2241));
OR2X1 g135765(.A (n_523), .B (n_502), .Y (n_1056));
INVX1 g136717(.A (n_1049), .Y (n_13019));
NOR2X1 g136295(.A (si[18]), .B (n_693), .Y (n_2286));
INVX1 g137387(.A (n_1054), .Y (n_27042));
NAND2X1 g136318(.A (n_7841), .B (addr_438), .Y (n_1899));
INVX1 g136714(.A (n_983), .Y (n_31273));
NOR2X1 g135444(.A (n_978), .B (n_980), .Y (n_1632));
INVX1 g136718(.A (n_1049), .Y (n_13024));
OR2X1 g135310(.A (P3_reg3[4] ), .B (n_820), .Y (n_1534));
NOR2X1 g135529(.A (n_1048), .B (n_1266), .Y (n_1963));
INVX1 g135855(.A (n_1361), .Y (n_1047));
INVX1 g135882(.A (n_1044), .Y (n_1629));
INVX1 g136103(.A (n_1042), .Y (n_1043));
NOR2X1 g135585(.A (n_1299), .B (n_1041), .Y (n_1694));
NOR2X1 g136185(.A (si[19]), .B (datao_2[19] ), .Y (n_1555));
INVX1 g136014(.A (n_1283), .Y (n_1040));
INVX1 g136227(.A (n_1036), .Y (n_1037));
INVX1 g136032(.A (n_1327), .Y (n_1035));
INVX1 g137860(.A (n_1203), .Y (n_1486));
NAND2X1 g135483(.A (n_1508), .B (n_896), .Y (n_2078));
OR2X1 g135942(.A (n_34849), .B (n_33567), .Y (n_1033));
NAND3X1 g135452(.A (n_910), .B (n_1032), .C (n_1031), .Y (n_1173));
NOR2X1 g136507(.A (si[17]), .B (n_475), .Y (n_1536));
AND2X1 g136157(.A (P3_IR[26] ), .B (n_3686), .Y (n_1030));
NAND3X1 g135478(.A (addr_447), .B (addr_446), .C (addr_453), .Y(n_1029));
NOR2X1 g136243(.A (si[14]), .B (n_928), .Y (n_1608));
NAND3X1 g135507(.A (n_911), .B (n_1027), .C (n_2105), .Y (n_2373));
INVX1 g136519(.A (n_1546), .Y (n_1026));
NOR2X1 g136420(.A (n_481), .B (addr_439), .Y (n_1640));
INVX1 g136279(.A (n_1022), .Y (n_1023));
NAND2X1 g136293(.A (si[16]), .B (n_12454), .Y (n_1865));
NOR2X1 g136382(.A (n_8079), .B (addr_436), .Y (n_1652));
INVX1 g136733(.A (n_917), .Y (n_31388));
NAND2X1 g136416(.A (si[21]), .B (n_12026), .Y (n_1593));
NOR2X1 g135636(.A (n_1065), .B (n_1162), .Y (n_1560));
OR2X1 g135854(.A (n_1968), .B (n_609), .Y (n_1020));
AND2X1 g135446(.A (n_946), .B (n_994), .Y (n_2086));
OR2X1 g135832(.A (n_1018), .B (n_609), .Y (n_1019));
NAND2X1 g135809(.A (P3_reg3[19] ), .B (n_1017), .Y (n_13003));
NAND2X1 g136451(.A (si[30]), .B (n_479), .Y (n_1479));
AND2X1 g136007(.A (n_1015), .B (n_852), .Y (n_1016));
OR2X1 g135830(.A (n_1012), .B (n_873), .Y (n_1013));
NAND2X1 g136011(.A (P3_reg3[4] ), .B (n_1017), .Y (n_13187));
INVX1 g137851(.A (n_852), .Y (n_1407));
NOR2X1 g135645(.A (n_1374), .B (n_863), .Y (n_4100));
AND2X1 g135972(.A (n_34205), .B (n_33567), .Y (n_1011));
OR2X1 g136469(.A (P1_IR[23] ), .B (P1_IR[20] ), .Y (n_1009));
OR2X1 g134846(.A (n_1007), .B (n_110), .Y (n_1300));
OR2X1 g136136(.A (P3_reg3[4] ), .B (P3_reg3[3] ), .Y (n_1006));
INVX1 g135285(.A (n_1003), .Y (n_1004));
OR2X1 g135616(.A (n_1357), .B (n_925), .Y (n_4341));
INVX1 g136129(.A (n_1001), .Y (n_1002));
INVX1 g137076(.A (n_34700), .Y (n_1619));
NOR2X1 g135297(.A (n_1838), .B (si[30]), .Y (n_1000));
OR2X1 g135917(.A (n_653), .B (n_998), .Y (n_999));
NAND2X1 g135490(.A (n_997), .B (n_1197), .Y (n_1834));
OR2X1 g136262(.A (si[12]), .B (n_11802), .Y (n_1552));
NAND2X1 g135343(.A (n_994), .B (n_905), .Y (n_1320));
NOR2X1 g135312(.A (n_957), .B (n_992), .Y (n_2393));
NOR2X1 g136396(.A (si[16]), .B (n_12454), .Y (n_1671));
OR2X1 g136025(.A (n_32395), .B (n_998), .Y (n_986));
OR2X1 g135864(.A (n_984), .B (n_609), .Y (n_985));
INVX1 g136713(.A (n_983), .Y (n_31744));
AND2X1 g135488(.A (n_982), .B (n_981), .Y (n_1500));
NOR2X1 g135413(.A (n_878), .B (n_953), .Y (n_1459));
NOR2X1 g135414(.A (n_980), .B (n_979), .Y (n_1817));
NAND2X1 g136116(.A (n_7843), .B (addr_430), .Y (n_1894));
NAND2X1 g135582(.A (n_1603), .B (n_1420), .Y (n_2159));
NOR2X1 g135604(.A (n_1162), .B (n_716), .Y (n_1566));
NOR2X1 g135442(.A (n_1496), .B (n_978), .Y (n_1658));
NAND2X1 g136008(.A (P3_reg3[15] ), .B (n_1017), .Y (n_13009));
INVX1 g136679(.A (n_7058), .Y (n_31774));
NOR2X1 g135330(.A (n_736), .B (n_973), .Y (n_1325));
AND2X1 g135501(.A (n_746), .B (n_972), .Y (n_2360));
OR2X1 g134708(.A (n_1007), .B (n_339), .Y (n_1456));
NAND2X1 g135591(.A (n_1209), .B (n_847), .Y (n_1693));
INVX1 g135466(.A (n_614), .Y (n_969));
OR2X1 g135961(.A (n_864), .B (n_33566), .Y (n_967));
NOR2X1 g135392(.A (n_898), .B (n_802), .Y (n_965));
INVX1 g136723(.A (n_631), .Y (n_31081));
INVX2 g137171(.A (n_3196), .Y (n_1423));
NAND2X1 g135588(.A (n_929), .B (n_779), .Y (n_1893));
NOR2X1 g136494(.A (si[6]), .B (n_804), .Y (n_1419));
INVX1 g136689(.A (n_903), .Y (n_31783));
INVX1 g135905(.A (n_1263), .Y (n_1268));
NOR2X1 g135423(.A (n_963), .B (n_962), .Y (n_1945));
OR2X1 g135651(.A (n_781), .B (n_1576), .Y (n_1813));
NOR2X1 g136356(.A (si[8]), .B (n_12184), .Y (n_1537));
INVX1 g136719(.A (n_1049), .Y (n_31979));
NOR2X1 g135369(.A (n_963), .B (n_1697), .Y (n_1471));
NOR2X1 g135634(.A (n_1221), .B (n_979), .Y (n_2077));
INVX1 g136709(.A (n_983), .Y (n_30792));
NAND2X1 g135962(.A (P3_reg3[5] ), .B (n_1017), .Y (n_13001));
OR2X1 g136207(.A (P1_IR[19] ), .B (P1_IR[16] ), .Y (n_959));
NOR2X1 g135494(.A (n_497), .B (n_1224), .Y (n_1438));
NOR2X1 g136349(.A (si[13]), .B (n_12030), .Y (n_1607));
NAND2X1 g136216(.A (n_12319), .B (si[26]), .Y (n_1373));
NOR2X1 g135365(.A (n_957), .B (n_871), .Y (n_2352));
INVX1 g136429(.A (n_1545), .Y (n_956));
INVX1 g136825(.A (n_762), .Y (n_1645));
NAND2X1 g135405(.A (n_1079), .B (n_955), .Y (n_1848));
NOR2X1 g135599(.A (n_953), .B (n_543), .Y (n_954));
INVX1 g136238(.A (n_950), .Y (n_951));
NAND2X1 g135332(.A (n_949), .B (n_850), .Y (n_1427));
INVX1 g136431(.A (n_1096), .Y (n_947));
AND2X1 g135541(.A (n_266), .B (n_946), .Y (n_1617));
NOR2X1 g135375(.A (n_1748), .B (n_1374), .Y (n_1778));
AND2X1 g136281(.A (n_943), .B (n_1666), .Y (n_944));
NAND2X1 g135453(.A (n_980), .B (n_955), .Y (n_1849));
INVX1 g136331(.A (n_630), .Y (n_1562));
NAND2X1 g136467(.A (n_939), .B (n_1968), .Y (n_940));
NAND2X1 g136294(.A (n_8083), .B (addr_437), .Y (n_1908));
NOR2X1 g135650(.A (n_1589), .B (n_1697), .Y (n_1996));
INVX1 g135997(.A (n_1246), .Y (n_937));
NOR2X1 g135623(.A (n_1224), .B (n_1048), .Y (n_1830));
NOR2X1 g136443(.A (P3_IR[28] ), .B (P3_IR[27] ), .Y (n_934));
INVX1 g136126(.A (n_450), .Y (n_1541));
NAND2X1 g136440(.A (P3_reg3[2] ), .B (n_7243), .Y (n_931));
NAND2X1 g136149(.A (si[20]), .B (n_12322), .Y (n_1588));
AND2X1 g135608(.A (n_929), .B (n_747), .Y (n_1691));
NAND2X1 g136326(.A (si[14]), .B (n_928), .Y (n_1867));
INVX1 g136225(.A (n_1190), .Y (n_927));
NOR2X1 g136287(.A (addr_447), .B (n_8361), .Y (n_1639));
NAND2X1 g135930(.A (P3_reg3[14] ), .B (n_1017), .Y (n_13012));
NOR2X1 g135319(.A (n_1356), .B (n_925), .Y (n_926));
INVX1 g137880(.A (n_33579), .Y (n_3719));
NAND2X1 g136365(.A (n_8079), .B (addr_436), .Y (n_1715));
CLKBUFX1 g136750(.A (n_3964), .Y (n_31275));
OR2X1 g136191(.A (n_33371), .B (n_33587), .Y (n_1125));
NAND2X1 g136202(.A (si[11]), .B (datao_1[11] ), .Y (n_1615));
INVX1 g135934(.A (n_1388), .Y (n_922));
NOR2X1 g135429(.A (n_921), .B (n_877), .Y (n_2260));
INVX1 g136684(.A (n_811), .Y (n_31951));
INVX1 g135945(.A (n_1167), .Y (n_918));
INVX1 g136482(.A (n_915), .Y (n_1104));
OR2X1 g136522(.A (n_1015), .B (n_33587), .Y (n_914));
NOR2X1 g136355(.A (P3_IR[26] ), .B (P3_IR[25] ), .Y (n_1345));
INVX1 g135995(.A (n_1230), .Y (n_912));
AND2X1 g135566(.A (n_911), .B (n_910), .Y (n_1240));
INVX1 g136277(.A (n_34528), .Y (n_32566));
NOR2X1 g136044(.A (P2_IR[28] ), .B (P2_IR[27] ), .Y (n_908));
NOR2X1 g136459(.A (P2_IR[26] ), .B (P2_IR[25] ), .Y (n_1101));
AND2X1 g135455(.A (n_905), .B (n_892), .Y (n_2938));
OR2X1 g136194(.A (n_7839), .B (n_8117), .Y (n_1854));
INVX1 g135784(.A (n_1372), .Y (n_902));
INVX2 g136691(.A (n_903), .Y (n_31850));
INVX1 g135834(.A (n_1233), .Y (n_900));
INVX1 g136730(.A (n_392), .Y (n_15643));
OR2X1 g135336(.A (n_898), .B (n_897), .Y (n_1437));
NAND2X1 g135357(.A (n_1316), .B (n_896), .Y (n_1501));
INVX1 g135696(.A (n_441), .Y (n_895));
INVX1 g136712(.A (n_983), .Y (n_31278));
OR2X1 g135957(.A (n_589), .B (n_377), .Y (n_893));
AND2X1 g135583(.A (n_892), .B (n_808), .Y (n_2518));
INVX1 g135974(.A (n_1341), .Y (n_1244));
NAND2X1 g136410(.A (si[8]), .B (n_12184), .Y (n_1604));
NAND2X1 g135331(.A (n_1143), .B (n_889), .Y (n_2336));
OR2X1 g135896(.A (n_35867), .B (P2_IR[31] ), .Y (n_888));
AND2X1 g135847(.A (P3_IR[15] ), .B (n_33566), .Y (n_886));
NAND2X1 g135838(.A (P3_reg3[16] ), .B (n_1017), .Y (n_13007));
NAND4X1 g135259(.A (n_880), .B (P1_reg3[3] ), .C (P1_reg3[5] ), .D(P1_reg3[4] ), .Y (n_2226));
NAND2X1 g136172(.A (n_13675), .B (n_7243), .Y (n_879));
NOR2X1 g135643(.A (n_878), .B (n_877), .Y (n_1979));
AND2X1 g136406(.A (P1_IR[25] ), .B (n_873), .Y (n_874));
NAND2X1 g135910(.A (P3_reg3[6] ), .B (n_1017), .Y (n_12995));
NOR2X1 g135340(.A (n_810), .B (n_871), .Y (n_1431));
INVX1 g136087(.A (n_869), .Y (n_870));
INVX1 g137179(.A (P3_IR[31] ), .Y (n_1512));
AND2X1 g136321(.A (n_864), .B (n_1724), .Y (n_865));
NOR2X1 g135315(.A (n_696), .B (n_863), .Y (n_1913));
INVX1 g137035(.A (n_15981), .Y (n_15968));
INVX1 g135850(.A (n_1234), .Y (n_862));
OR2X1 g135798(.A (n_1969), .B (n_762), .Y (n_861));
NAND2X1 g136109(.A (si[22]), .B (n_12188), .Y (n_2244));
OR2X1 g135980(.A (n_1800), .B (P2_IR[31] ), .Y (n_858));
NOR2X1 g135473(.A (n_855), .B (n_854), .Y (n_856));
OR2X1 g135794(.A (n_1799), .B (n_852), .Y (n_853));
INVX1 g135268(.A (n_1453), .Y (n_2598));
INVX1 g135825(.A (n_1314), .Y (n_851));
NOR2X1 g135396(.A (n_1177), .B (n_1496), .Y (n_1494));
NOR2X1 g136093(.A (si[15]), .B (n_12028), .Y (n_1739));
NAND2X1 g135481(.A (n_850), .B (n_1209), .Y (n_1692));
NAND2X1 g136306(.A (si[12]), .B (n_11802), .Y (n_1855));
NAND2X1 g135435(.A (n_850), .B (n_849), .Y (n_1428));
NOR2X1 g135649(.A (n_847), .B (n_1041), .Y (n_2168));
INVX1 g136094(.A (n_845), .Y (n_846));
INVX1 g136000(.A (n_1344), .Y (n_844));
NOR2X1 g136151(.A (si[4]), .B (datao_1[4] ), .Y (n_1489));
NAND2X1 g135963(.A (P3_reg3[12] ), .B (n_1017), .Y (n_13023));
INVX1 g136445(.A (n_34527), .Y (n_842));
INVX1 g136706(.A (n_983), .Y (n_31605));
INVX1 g136341(.A (n_1675), .Y (n_840));
NAND2X1 g136465(.A (si[5]), .B (datao_1[5] ), .Y (n_1904));
NAND2X1 g135573(.A (n_1119), .B (n_955), .Y (n_1425));
NOR2X1 g135349(.A (n_733), .B (n_1328), .Y (n_1914));
NOR2X1 g136412(.A (n_7833), .B (addr_435), .Y (n_1651));
NAND2X1 g135989(.A (P3_reg3[13] ), .B (n_1017), .Y (n_13014));
NOR2X1 g135433(.A (n_1065), .B (n_849), .Y (n_1399));
NAND2X1 g136488(.A (n_7839), .B (n_8117), .Y (n_2148));
NAND2X1 g136305(.A (si[24]), .B (n_667), .Y (n_1433));
INVX1 g135812(.A (n_1352), .Y (n_833));
INVX1 g136019(.A (n_1195), .Y (n_832));
NOR2X1 g134702(.A (n_831), .B (n_830), .Y (n_1524));
NOR2X1 g135547(.A (n_855), .B (n_829), .Y (n_1565));
NAND4X1 g135768(.A (addr_438), .B (addr_437), .C (addr_435), .D(addr_436), .Y (n_828));
OR2X1 g135487(.A (n_536), .B (n_399), .Y (n_1402));
NOR2X1 g136455(.A (si[2]), .B (n_732), .Y (n_1498));
OR2X1 g135885(.A (n_1015), .B (n_826), .Y (n_827));
NOR2X1 g136470(.A (P1_IR[28] ), .B (P1_IR[27] ), .Y (n_825));
INVX1 g136339(.A (n_1238), .Y (n_824));
NAND2X1 g135929(.A (P3_reg3[10] ), .B (n_1017), .Y (n_13018));
OR2X1 g135428(.A (n_247), .B (n_820), .Y (n_2089));
INVX1 g135977(.A (n_1958), .Y (n_817));
INVX1 g135538(.A (n_651), .Y (n_812));
OR2X1 g135437(.A (n_2035), .B (n_788), .Y (n_1577));
INVX1 g136686(.A (n_811), .Y (n_31696));
NOR2X1 g135440(.A (n_810), .B (n_710), .Y (n_1491));
AND2X1 g135372(.A (n_809), .B (n_808), .Y (n_2084));
NAND2X1 g136023(.A (P3_reg3[11] ), .B (n_1017), .Y (n_13016));
NAND2X1 g135495(.A (n_1087), .B (n_1163), .Y (n_2161));
INVX1 g136528(.A (n_805), .Y (n_806));
NAND2X1 g136055(.A (si[25]), .B (n_641), .Y (n_2989));
NAND2X1 g136276(.A (si[6]), .B (n_804), .Y (n_1821));
AND2X1 g135505(.A (n_88), .B (n_911), .Y (n_1618));
NOR2X1 g135460(.A (n_802), .B (n_801), .Y (n_1682));
AND2X1 g135867(.A (n_799), .B (n_873), .Y (n_800));
NAND2X1 g136235(.A (n_8074), .B (addr_429), .Y (n_1886));
NOR2X1 g136265(.A (n_8074), .B (addr_429), .Y (n_1595));
INVX1 g135951(.A (n_1381), .Y (n_796));
NOR2X1 g136187(.A (n_8083), .B (addr_437), .Y (n_1488));
INVX1 g135801(.A (n_1250), .Y (n_795));
INVX1 g135817(.A (n_1653), .Y (n_794));
NOR2X1 g135389(.A (n_1136), .B (n_636), .Y (n_2059));
INVX1 g136738(.A (n_34188), .Y (n_15975));
NOR2X1 g134852(.A (n_831), .B (n_141), .Y (n_1522));
NAND2X1 g135376(.A (n_978), .B (n_1119), .Y (n_1416));
INVX1 g135839(.A (n_1353), .Y (n_790));
NAND2X1 g136024(.A (P3_reg3[17] ), .B (n_1017), .Y (n_13005));
NOR2X1 g135383(.A (n_1223), .B (n_1177), .Y (n_2844));
NOR2X1 g135445(.A (n_962), .B (n_788), .Y (n_1609));
INVX1 g136687(.A (n_811), .Y (n_31694));
NAND2X1 g136313(.A (P3_reg3[4] ), .B (P3_reg3[3] ), .Y (n_787));
NOR2X1 g136236(.A (addr_446), .B (n_482), .Y (n_2141));
NAND2X1 g135960(.A (P3_reg3[9] ), .B (n_1017), .Y (n_13026));
INVX1 g136703(.A (n_13010), .Y (n_1292));
INVX1 g136052(.A (n_1543), .Y (n_782));
NOR2X1 g136124(.A (n_7841), .B (addr_438), .Y (n_1468));
NOR2X1 g135647(.A (n_1748), .B (n_781), .Y (n_3506));
INVX1 g135969(.A (n_1249), .Y (n_780));
NAND2X1 g135569(.A (n_779), .B (n_910), .Y (n_1310));
NAND2X1 g136334(.A (si[15]), .B (n_12028), .Y (n_1866));
NAND2X1 g135362(.A (n_774), .B (n_405), .Y (n_1307));
NAND3X1 g135309(.A (n_1890), .B (n_1107), .C (n_241), .Y (n_773));
NOR2X1 g136174(.A (si[3]), .B (n_12022), .Y (n_1497));
XOR2X1 g135770(.A (n_263), .B (addr_1), .Y (n_1626));
INVX1 g136690(.A (n_903), .Y (n_31260));
OR2X1 g136120(.A (P2_IR[23] ), .B (P2_IR[20] ), .Y (n_767));
OR2X1 g135829(.A (n_764), .B (n_826), .Y (n_765));
OR2X1 g135894(.A (n_939), .B (n_762), .Y (n_763));
INVX1 g136533(.A (n_760), .Y (n_761));
INVX1 g136805(.A (n_3474), .Y (n_3656));
INVX1 g136749(.A (n_3964), .Y (n_27232));
INVX1 g135868(.A (n_1282), .Y (n_758));
AND2X1 g136357(.A (n_491), .B (si[28]), .Y (n_1477));
INVX1 g136003(.A (n_1232), .Y (n_757));
INVX1 g136685(.A (n_811), .Y (n_31922));
INVX1 g135954(.A (n_1243), .Y (n_753));
OR2X1 g135976(.A (n_1720), .B (n_826), .Y (n_752));
INVX1 g135876(.A (n_1630), .Y (n_748));
AND2X1 g135549(.A (n_747), .B (n_746), .Y (n_1462));
INVX1 g136681(.A (n_7062), .Y (n_30421));
NOR2X1 g135512(.A (n_849), .B (n_847), .Y (n_1663));
NAND2X1 g135578(.A (n_896), .B (n_1136), .Y (n_1502));
CLKBUFX1 g137098(.A (n_3185), .Y (n_31097));
INVX1 g136009(.A (n_1217), .Y (n_744));
AND2X1 g135866(.A (n_34544), .B (P3_IR[31] ), .Y (n_743));
NOR2X1 g135381(.A (n_1223), .B (n_1357), .Y (n_3526));
AND2X1 g136189(.A (n_120), .B (n_739), .Y (n_741));
NOR2X1 g135621(.A (n_687), .B (n_736), .Y (n_1214));
NAND2X1 g136397(.A (addr_447), .B (n_8361), .Y (n_1887));
NOR2X1 g135358(.A (n_734), .B (n_733), .Y (n_735));
NAND2X1 g136201(.A (si[2]), .B (n_732), .Y (n_1760));
NOR2X1 g136328(.A (n_7843), .B (addr_430), .Y (n_1572));
INVX1 g137086(.A (P2_n_749), .Y (n_15484));
INVX1 g136146(.A (n_33356), .Y (n_731));
NOR2X1 g135482(.A (n_1375), .B (n_1589), .Y (n_2101));
NAND2X1 g135351(.A (n_1316), .B (n_1143), .Y (n_2204));
NAND2X1 g136051(.A (si[3]), .B (n_12022), .Y (n_1759));
AND2X1 g135807(.A (n_727), .B (n_33567), .Y (n_728));
INVX1 g135939(.A (n_1189), .Y (n_725));
AND2X1 g135887(.A (n_32941), .B (P3_IR[31] ), .Y (n_724));
INVX2 g136291(.A (n_722), .Y (n_1939));
INVX1 g136489(.A (n_720), .Y (n_721));
NOR2X1 g136367(.A (si[5]), .B (datao_1[5] ), .Y (n_1516));
XOR2X1 g135769(.A (P2_reg3[4] ), .B (P2_reg3[3] ), .Y (n_1183));
OR2X1 g135994(.A (n_439), .B (n_33567), .Y (n_718));
NAND2X1 g135627(.A (n_1163), .B (n_716), .Y (n_1701));
AND2X1 g135848(.A (n_2742), .B (n_998), .Y (n_715));
NAND2X1 g136338(.A (n_7833), .B (addr_435), .Y (n_1872));
NAND2X1 g136002(.A (P3_reg3[8] ), .B (n_1017), .Y (n_12997));
XOR2X1 g135756(.A (si[31]), .B (datao_1[31] ), .Y (n_714));
NAND2X1 g135884(.A (n_12458), .B (n_13), .Y (n_1343));
NOR2X1 g135883(.A (datao_1[24] ), .B (n_171), .Y (n_1044));
INVX1 g136098(.A (n_710), .Y (n_711));
INVX1 g136831(.A (n_609), .Y (n_3705));
INVX1 g136282(.A (n_863), .Y (n_1952));
INVX1 g136372(.A (n_788), .Y (n_708));
INVX1 g135267(.A (n_707), .Y (n_835));
INVX1 g136806(.A (n_762), .Y (n_3474));
INVX1 g135274(.A (n_706), .Y (n_2291));
NAND2X1 g136337(.A (n_33568), .B (n_704), .Y (n_1149));
NOR2X1 g136047(.A (n_233), .B (addr_426), .Y (n_2118));
NOR2X1 g136096(.A (si[11]), .B (n_12458), .Y (n_1363));
INVX1 g136595(.A (P3_reg3[3] ), .Y (n_2721));
INVX1 g136695(.A (n_34188), .Y (n_7417));
INVX1 g136176(.A (n_701), .Y (n_1259));
XOR2X1 g135764(.A (si[31]), .B (datao_2[31] ), .Y (n_698));
NAND2X1 g136053(.A (addr_451), .B (addr_432), .Y (n_1543));
INVX1 g136133(.A (n_696), .Y (n_1045));
INVX1 g136688(.A (n_7243), .Y (n_811));
INVX1 g136057(.A (n_687), .Y (n_688));
AND2X1 g136408(.A (n_799), .B (n_686), .Y (n_1556));
AND2X1 g136059(.A (n_282), .B (n_664), .Y (n_1121));
INVX1 g136240(.A (n_978), .Y (n_685));
NAND2X1 g136483(.A (n_684), .B (n_943), .Y (n_915));
NAND2X1 g136140(.A (n_607), .B (n_287), .Y (n_683));
NAND2X1 g136088(.A (n_632), .B (n_682), .Y (n_869));
INVX1 g136822(.A (n_873), .Y (n_3596));
NOR2X1 g136418(.A (n_493), .B (n_680), .Y (n_681));
INVX1 g136437(.A (n_997), .Y (n_679));
NOR2X1 g136005(.A (n_535), .B (datao_2[16] ), .Y (n_1182));
INVX1 g136310(.A (n_854), .Y (n_1139));
NAND2X1 g135998(.A (n_68), .B (datao_2[7] ), .Y (n_1246));
NAND2X1 g135941(.A (n_547), .B (datao_2[20] ), .Y (n_1189));
NAND2X1 g135893(.A (n_625), .B (datao_2[26] ), .Y (n_2173));
INVX1 g136358(.A (n_980), .Y (n_670));
NAND2X1 g136444(.A (n_1018), .B (n_668), .Y (n_1099));
NOR2X1 g135837(.A (n_116), .B (datao_1[28] ), .Y (n_2055));
INVX1 g137960(.A (n_1753), .Y (n_666));
INVX1 g136121(.A (n_1080), .Y (n_665));
NOR2X1 g135926(.A (n_447), .B (datao_2[22] ), .Y (n_1368));
NAND2X1 g136061(.A (n_545), .B (n_664), .Y (n_1166));
INVX1 g136141(.A (n_663), .Y (n_2146));
NOR2X1 g135952(.A (n_540), .B (datao_2[14] ), .Y (n_1381));
XOR2X1 g135771(.A (P1_reg3[4] ), .B (P1_reg3[3] ), .Y (n_1003));
AND2X1 g136503(.A (n_799), .B (n_658), .Y (n_1359));
NOR2X1 g136508(.A (addr_451), .B (addr_432), .Y (n_1544));
NAND2X1 g136162(.A (n_1878), .B (n_657), .Y (n_1165));
NAND2X1 g136534(.A (n_564), .B (n_33568), .Y (n_760));
NAND2X1 g135802(.A (n_54), .B (datao_2[27] ), .Y (n_1250));
INVX1 g136860(.A (n_1800), .Y (n_654));
INVX1 g137190(.A (n_653), .Y (n_1094));
AND2X1 g136385(.A (n_100), .B (n_600), .Y (n_652));
INVX1 g138074(.A (n_120), .Y (n_1274));
NAND3X1 g135539(.A (addr_431), .B (addr_430), .C (addr_434), .Y(n_651));
NOR2X1 g135935(.A (n_602), .B (datao_2[5] ), .Y (n_1388));
NOR2X1 g136150(.A (n_649), .B (n_637), .Y (n_650));
NOR2X1 g135799(.A (datao_1[19] ), .B (n_612), .Y (n_1551));
NAND2X1 g136004(.A (n_455), .B (datao_2[3] ), .Y (n_1232));
NAND2X1 g135835(.A (n_585), .B (datao_2[4] ), .Y (n_1233));
NAND2X1 g136104(.A (n_211), .B (n_658), .Y (n_1042));
INVX1 g136170(.A (n_1066), .Y (n_640));
NAND2X1 g136164(.A (n_35868), .B (n_1799), .Y (n_639));
AND2X1 g136394(.A (n_637), .B (n_6), .Y (n_638));
INVX1 g136499(.A (n_636), .Y (n_1315));
NOR2X1 g136340(.A (n_125), .B (n_316), .Y (n_1238));
INVX1 g136197(.A (n_634), .Y (n_635));
NAND2X1 g136160(.A (n_632), .B (n_452), .Y (n_1075));
CLKBUFX1 g136721(.A (n_631), .Y (n_1049));
NAND2X2 g136332(.A (n_629), .B (n_218), .Y (n_630));
NOR2X1 g135970(.A (n_625), .B (datao_2[26] ), .Y (n_1249));
INVX1 g136800(.A (n_33261), .Y (n_622));
INVX1 g136244(.A (n_1135), .Y (n_1110));
INVX1 g136335(.A (n_973), .Y (n_620));
INVX1 g136250(.A (n_979), .Y (n_619));
INVX1 g137909(.A (n_939), .Y (n_618));
NAND2X1 g136084(.A (n_527), .B (n_704), .Y (n_1069));
AND2X1 g136453(.A (n_46), .B (n_69), .Y (n_615));
NAND3X1 g135467(.A (addr_491), .B (addr_489), .C (addr_490), .Y(n_614));
INVX1 g137861(.A (n_33814), .Y (n_1203));
AND2X1 g135975(.A (datao_1[19] ), .B (n_612), .Y (n_1341));
INVX1 g136039(.A (n_781), .Y (n_611));
AND2X1 g136320(.A (n_549), .B (n_607), .Y (n_608));
NAND2X1 g136239(.A (n_606), .B (n_764), .Y (n_950));
NOR2X1 g136541(.A (n_465), .B (n_464), .Y (n_605));
INVX1 g136246(.A (n_829), .Y (n_604));
INVX1 g136954(.A (n_1969), .Y (n_603));
NAND2X1 g135781(.A (n_602), .B (datao_2[5] ), .Y (n_1393));
AND2X1 g136487(.A (n_600), .B (n_1304), .Y (n_1090));
AND2X1 g136479(.A (n_1890), .B (n_686), .Y (n_1106));
INVX1 g136693(.A (n_7243), .Y (n_903));
INVX1 g136230(.A (n_1603), .Y (n_599));
INVX1 g136064(.A (n_1474), .Y (n_598));
NAND2X1 g136312(.A (n_1666), .B (n_1323), .Y (n_597));
AND2X1 g136531(.A (n_522), .B (n_521), .Y (n_596));
AND2X1 g136054(.A (n_594), .B (n_593), .Y (n_595));
OR2X1 g136067(.A (n_499), .B (n_498), .Y (n_592));
INVX1 g137605(.A (n_589), .Y (n_590));
AND2X1 g136518(.A (n_25), .B (n_60), .Y (n_588));
NAND2X1 g136115(.A (n_764), .B (n_682), .Y (n_1074));
NAND2X1 g135856(.A (n_515), .B (datao_2[15] ), .Y (n_1361));
AND2X1 g136468(.A (n_416), .B (n_415), .Y (n_587));
NOR2X1 g136434(.A (n_19), .B (n_586), .Y (n_1294));
NOR2X1 g135899(.A (n_585), .B (datao_2[4] ), .Y (n_1394));
NAND2X1 g135949(.A (n_492), .B (datao_2[6] ), .Y (n_1387));
INVX1 g136392(.A (n_716), .Y (n_584));
NOR2X1 g136063(.A (addr_450), .B (addr_431), .Y (n_1573));
CLKBUFX1 g136744(.A (n_392), .Y (n_31698));
NAND2X1 g136001(.A (datao_2[10] ), .B (n_1), .Y (n_1344));
INVX1 g136091(.A (n_1048), .Y (n_579));
NAND2X1 g136130(.A (n_1171), .B (n_578), .Y (n_1001));
NOR2X1 g135909(.A (n_528), .B (datao_2[18] ), .Y (n_1542));
AND2X1 g136370(.A (n_593), .B (n_727), .Y (n_1112));
INVX1 g136045(.A (n_949), .Y (n_572));
INVX1 g136204(.A (n_571), .Y (n_1270));
NAND2X1 g135950(.A (n_294), .B (datao_2[2] ), .Y (n_2066));
OR2X1 g136466(.A (n_411), .B (n_410), .Y (n_567));
NAND2X2 g136292(.A (n_34322), .B (n_34319), .Y (n_722));
AND2X1 g136255(.A (n_11), .B (n_34), .Y (n_563));
NAND2X1 g136020(.A (n_12330), .B (n_421), .Y (n_1195));
INVX1 g136957(.A (n_1720), .Y (n_562));
AND2X1 g136280(.A (n_367), .B (n_561), .Y (n_1022));
NOR2X1 g136226(.A (n_10057), .B (addr_424), .Y (n_1190));
AND2X1 g136502(.A (n_62), .B (n_40), .Y (n_558));
AND2X1 g136192(.A (n_442), .B (n_64), .Y (n_557));
NOR2X1 g136405(.A (addr_453), .B (addr_434), .Y (n_1563));
NAND2X1 g136520(.A (addr_452), .B (addr_433), .Y (n_1546));
AND2X1 g136460(.A (n_553), .B (n_552), .Y (n_555));
OR2X1 g136224(.A (n_553), .B (n_552), .Y (n_554));
INVX1 g136138(.A (n_855), .Y (n_1255));
NAND2X1 g136169(.A (n_606), .B (n_551), .Y (n_1085));
INVX1 g136071(.A (n_1580), .Y (n_550));
NAND2X1 g136523(.A (n_453), .B (n_549), .Y (n_1199));
NOR2X1 g136006(.A (n_547), .B (datao_2[20] ), .Y (n_1620));
NAND2X1 g136049(.A (n_545), .B (n_1323), .Y (n_546));
CLKBUFX1 g136745(.A (n_392), .Y (n_31781));
INVX4 g137172(.A (n_1724), .Y (n_3196));
INVX1 g136524(.A (n_543), .Y (n_544));
NAND2X1 g135953(.A (n_540), .B (datao_2[14] ), .Y (n_1469));
NAND2X1 g136188(.A (n_1878), .B (n_1666), .Y (n_539));
INVX1 g136751(.A (n_392), .Y (n_3964));
INVX1 g136112(.A (n_962), .Y (n_538));
NOR2X1 g135938(.A (n_529), .B (datao_2[13] ), .Y (n_1529));
INVX1 g136154(.A (n_536), .Y (n_814));
NAND2X1 g136015(.A (n_535), .B (datao_2[16] ), .Y (n_1283));
NAND2X1 g136260(.A (n_10057), .B (addr_424), .Y (n_1667));
NOR2X1 g135786(.A (n_424), .B (datao_2[17] ), .Y (n_1481));
INVX1 g137036(.A (P1_n_449), .Y (n_15981));
INVX1 g136678(.A (n_7243), .Y (n_7058));
NAND2X1 g136095(.A (n_1968), .B (n_668), .Y (n_845));
NAND2X1 g135785(.A (n_529), .B (datao_2[13] ), .Y (n_1372));
NAND2X1 g135814(.A (n_528), .B (datao_2[18] ), .Y (n_1352));
AND2X1 g135906(.A (datao_1[23] ), .B (n_32), .Y (n_1263));
NAND2X1 g136062(.A (n_527), .B (n_439), .Y (n_1150));
AND2X1 g136029(.A (n_10), .B (n_3), .Y (n_525));
NAND2X1 g135872(.A (n_275), .B (datao_2[0] ), .Y (n_1453));
OR2X1 g135978(.A (datao_1[30] ), .B (n_380), .Y (n_1958));
OR2X1 g136532(.A (n_522), .B (n_521), .Y (n_523));
NAND2X1 g136517(.A (n_1171), .B (n_488), .Y (n_1097));
INVX1 g136743(.A (n_392), .Y (n_7390));
INVX1 g137847(.A (n_852), .Y (n_3279));
NAND2X1 g135877(.A (n_138), .B (datao_2[25] ), .Y (n_1630));
NOR2X1 g135913(.A (n_515), .B (datao_2[15] ), .Y (n_1380));
NAND2X1 g136010(.A (n_393), .B (datao_2[21] ), .Y (n_1217));
INVX1 g136105(.A (n_1299), .Y (n_513));
NAND2X1 g136432(.A (n_984), .B (n_120), .Y (n_1096));
INVX1 g137564(.A (n_12670), .Y (n_991));
NOR2X1 g135900(.A (n_68), .B (datao_2[7] ), .Y (n_1247));
AND2X1 g136353(.A (n_150), .B (n_561), .Y (n_1089));
OR2X1 g136232(.A (n_432), .B (n_431), .Y (n_502));
AND2X1 g136060(.A (n_499), .B (n_498), .Y (n_500));
INVX1 g136463(.A (n_497), .Y (n_1142));
XOR2X1 g135774(.A (datao_1[31] ), .B (datao_2[31] ), .Y (n_496));
AND2X1 g136323(.A (n_493), .B (n_680), .Y (n_494));
NOR2X1 g135955(.A (n_492), .B (datao_2[6] ), .Y (n_1243));
INVX1 g136399(.A (n_1222), .Y (n_1052));
OR2X1 g135895(.A (n_54), .B (datao_2[27] ), .Y (n_1916));
NAND2X1 g136539(.A (n_1799), .B (n_551), .Y (n_1261));
NAND2X1 g136270(.A (n_984), .B (n_488), .Y (n_489));
INVX1 g137699(.A (n_1858), .Y (n_485));
INVX1 g136911(.A (n_34205), .Y (n_1227));
INVX1 g137115(.A (P2_n_749), .Y (n_1313));
NOR2X1 g135788(.A (datao_2[9] ), .B (n_153), .Y (n_1527));
NAND2X1 g136430(.A (addr_450), .B (addr_431), .Y (n_1545));
NOR2X1 g136033(.A (n_130), .B (addr_425), .Y (n_1327));
INVX1 g136195(.A (n_896), .Y (n_477));
INVX1 g136314(.A (n_1605), .Y (n_476));
NAND2X1 g136390(.A (n_1012), .B (n_578), .Y (n_1098));
OR2X1 g135912(.A (datao_1[29] ), .B (n_61), .Y (n_2303));
INVX1 g136504(.A (n_734), .Y (n_1750));
NOR2X1 g135851(.A (n_419), .B (datao_2[8] ), .Y (n_1234));
AND2X1 g136480(.A (n_32398), .B (n_32487), .Y (n_474));
NAND2X1 g135996(.A (datao_2[9] ), .B (n_153), .Y (n_1230));
NAND2X1 g136388(.A (n_1401), .B (n_1206), .Y (n_1082));
NOR2X1 g136516(.A (n_0), .B (n_22), .Y (n_472));
NOR2X1 g136253(.A (si[12]), .B (n_12330), .Y (n_1330));
AND2X1 g136529(.A (n_34090), .B (n_1236), .Y (n_805));
AND2X1 g136163(.A (n_465), .B (n_464), .Y (n_466));
INVX1 g136233(.A (n_1265), .Y (n_463));
INVX1 g136675(.A (n_7243), .Y (n_31490));
CLKBUFX1 g136716(.A (n_631), .Y (n_983));
INVX1 g136676(.A (n_7243), .Y (n_7062));
INVX1 g136300(.A (n_457), .Y (n_458));
NAND2X1 g136342(.A (addr_453), .B (addr_434), .Y (n_1675));
NOR2X1 g135811(.A (n_455), .B (datao_2[3] ), .Y (n_1569));
NAND2X1 g136497(.A (n_453), .B (n_452), .Y (n_454));
INVX1 g136477(.A (n_733), .Y (n_1749));
NOR2X1 g135818(.A (n_451), .B (datao_2[1] ), .Y (n_1653));
NAND2X1 g136127(.A (n_1236), .B (n_287), .Y (n_450));
INVX1 g136447(.A (n_963), .Y (n_449));
INVX1 g136704(.A (n_34188), .Y (n_13010));
NAND2X1 g135947(.A (n_447), .B (datao_2[22] ), .Y (n_1167));
NOR2X1 g136384(.A (n_442), .B (n_31), .Y (n_443));
AOI21X1 g135697(.A0 (P3_reg3[2] ), .A1 (P3_reg3[3] ), .B0(P3_reg3[4] ), .Y (n_441));
NAND2X1 g136428(.A (n_684), .B (n_439), .Y (n_440));
NOR2X1 g135826(.A (n_12458), .B (n_13), .Y (n_1314));
NOR2X1 g136097(.A (addr_452), .B (addr_433), .Y (n_1547));
INVX1 g136117(.A (n_1375), .Y (n_435));
INVX1 g136656(.A (n_34199), .Y (n_434));
AND2X1 g136501(.A (n_432), .B (n_431), .Y (n_433));
INVX1 g135269(.A (n_430), .Y (n_2798));
INVX1 g136343(.A (n_1177), .Y (n_428));
INVX1 g136267(.A (n_925), .Y (n_1754));
INVX1 g137440(.A (n_33371), .Y (n_1803));
NAND2X1 g135869(.A (n_424), .B (datao_2[17] ), .Y (n_1282));
INVX1 g137457(.A (n_1444), .Y (n_2779));
NOR2X1 g135981(.A (n_12330), .B (n_421), .Y (n_1531));
INVX1 g137099(.A (P2_n_749), .Y (n_3185));
NAND2X1 g135815(.A (n_419), .B (datao_2[8] ), .Y (n_1296));
OR2X1 g136110(.A (n_416), .B (n_415), .Y (n_417));
NAND2X1 g135840(.A (datao_1[29] ), .B (n_61), .Y (n_1353));
INVX1 g136030(.A (n_1041), .Y (n_414));
NAND2X1 g135927(.A (n_451), .B (datao_2[1] ), .Y (n_1654));
NAND2X1 g136490(.A (n_657), .B (n_1323), .Y (n_720));
AND2X1 g136070(.A (n_411), .B (n_410), .Y (n_412));
NAND2X1 g136515(.A (n_607), .B (n_452), .Y (n_409));
NOR2X1 g135914(.A (datao_2[10] ), .B (n_1), .Y (n_1523));
INVX1 g136423(.A (n_405), .Y (n_406));
NAND2X1 g136427(.A (n_2721), .B (n_2105), .Y (n_403));
INVX1 g136737(.A (n_349), .Y (n_917));
NOR2X1 g135844(.A (datao_1[23] ), .B (n_32), .Y (n_1495));
INVX1 g136219(.A (n_889), .Y (n_400));
INVX1 g136258(.A (n_399), .Y (n_989));
INVX1 g136375(.A (n_847), .Y (n_397));
AND2X1 g136361(.A (n_1206), .B (n_345), .Y (n_1289));
INVX1 g136829(.A (n_609), .Y (n_1277));
INVX1 g136898(.A (n_396), .Y (n_1253));
INVX1 g136456(.A (n_850), .Y (n_395));
INVX1 g136484(.A (n_1141), .Y (n_394));
NOR2X1 g135827(.A (n_393), .B (datao_2[21] ), .Y (n_1385));
NAND2X1 g136228(.A (n_1018), .B (n_1012), .Y (n_1036));
INVX1 g136752(.A (n_392), .Y (n_4029));
INVX1 g136179(.A (n_1356), .Y (n_390));
NAND2X1 g136111(.A (si[1]), .B (datao_1[1] ), .Y (n_1134));
NAND2X1 g136383(.A (si[1]), .B (datao_2[1] ), .Y (n_1276));
INVX1 g137292(.A (n_34524), .Y (n_1211));
NOR2X1 g136252(.A (P3_reg3[8] ), .B (P3_reg3[9] ), .Y (n_911));
NOR2X1 g136283(.A (datao_1[28] ), .B (si[28]), .Y (n_863));
CLKBUFX1 g136861(.A (n_33559), .Y (n_1800));
NOR2X1 g136461(.A (si[7]), .B (datao_2[7] ), .Y (n_849));
AND2X1 g136108(.A (P2_reg3[17] ), .B (P2_reg3[16] ), .Y (n_982));
NAND2X1 g136259(.A (P1_reg3[10] ), .B (P1_reg3[11] ), .Y (n_399));
NAND2X1 g136336(.A (P2_reg3[10] ), .B (P2_reg3[11] ), .Y (n_973));
AND2X1 g136079(.A (P1_reg3[24] ), .B (P1_reg3[25] ), .Y (n_2870));
NAND2X1 g136363(.A (si[19]), .B (datao_1[19] ), .Y (n_1590));
NOR2X1 g136359(.A (si[22]), .B (datao_2[22] ), .Y (n_980));
INVX1 g136849(.A (n_34321), .Y (n_864));
INVX1 g137461(.A (n_1464), .Y (n_371));
NAND2X1 g136090(.A (P1_reg3[17] ), .B (P1_reg3[16] ), .Y (n_802));
NAND2X1 g136155(.A (P1_reg3[8] ), .B (P1_reg3[9] ), .Y (n_536));
NOR2X1 g136248(.A (si[3]), .B (datao_2[3] ), .Y (n_829));
NOR2X1 g136221(.A (si[6]), .B (datao_2[6] ), .Y (n_1065));
NOR2X1 g136285(.A (si[13]), .B (datao_2[13] ), .Y (n_1266));
AND2X1 g136424(.A (P1_reg3[15] ), .B (P1_reg3[16] ), .Y (n_405));
NAND2X1 g136068(.A (P1_reg3[23] ), .B (P1_reg3[24] ), .Y (n_953));
NOR2X1 g136178(.A (P3_reg3[18] ), .B (P3_reg3[17] ), .Y (n_905));
NAND2X1 g136231(.A (si[7]), .B (datao_1[7] ), .Y (n_1603));
INVX1 g137595(.A (n_431), .Y (n_9670));
INVX1 g137510(.A (n_553), .Y (n_8079));
INVX1 g137042(.A (n_552), .Y (n_7833));
NOR2X1 g136125(.A (P3_reg3[14] ), .B (P3_reg3[13] ), .Y (n_946));
AND2X1 g136222(.A (P2_reg3[25] ), .B (P2_reg3[26] ), .Y (n_1490));
NAND2X1 g136143(.A (P2_reg3[3] ), .B (P2_reg3[4] ), .Y (n_1007));
NAND2X1 g136317(.A (P1_reg3[21] ), .B (P1_reg3[22] ), .Y (n_878));
OR2X1 g136065(.A (si[11]), .B (datao_1[11] ), .Y (n_1474));
NOR2X1 g136311(.A (si[1]), .B (datao_2[1] ), .Y (n_854));
NAND2X1 g136400(.A (datao_2[26] ), .B (si[26]), .Y (n_1222));
NOR2X1 g136442(.A (P3_reg3[24] ), .B (P3_reg3[23] ), .Y (n_809));
NOR2X1 g136441(.A (n_12319), .B (si[26]), .Y (n_1748));
NAND2X1 g136211(.A (P2_reg3[12] ), .B (P2_reg3[13] ), .Y (n_736));
OR2X1 g136082(.A (P3_reg3[6] ), .B (P3_reg3[5] ), .Y (n_820));
NAND2X1 g136156(.A (si[17]), .B (datao_2[17] ), .Y (n_1316));
NAND2X1 g136234(.A (si[13]), .B (datao_2[13] ), .Y (n_1265));
NOR2X1 g136475(.A (si[21]), .B (n_12026), .Y (n_1697));
NOR2X1 g136100(.A (P3_reg3[19] ), .B (P3_reg3[20] ), .Y (n_892));
NAND2X1 g136263(.A (P1_reg3[18] ), .B (P1_reg3[19] ), .Y (n_801));
NAND2X1 g136122(.A (si[20]), .B (datao_2[20] ), .Y (n_1080));
NAND2X1 g136171(.A (si[5]), .B (datao_2[5] ), .Y (n_1066));
NAND2X1 g136069(.A (P1_reg3[12] ), .B (P1_reg3[13] ), .Y (n_897));
NAND2X1 g136329(.A (P1_reg3[14] ), .B (P1_reg3[15] ), .Y (n_898));
NOR2X1 g136505(.A (si[30]), .B (datao_1[30] ), .Y (n_734));
INVX4 g136819(.A (n_998), .Y (n_609));
AND2X1 g136345(.A (P2_reg3[6] ), .B (P2_reg3[7] ), .Y (n_1517));
NOR2X1 g136042(.A (si[25]), .B (n_641), .Y (n_781));
AND2X1 g136208(.A (P1_reg3[6] ), .B (P1_reg3[7] ), .Y (n_880));
NAND2X1 g136080(.A (si[21]), .B (datao_2[21] ), .Y (n_1079));
AND2X1 g136449(.A (P1_reg3[13] ), .B (P1_reg3[14] ), .Y (n_774));
NAND2X1 g136525(.A (P1_reg3[25] ), .B (P1_reg3[26] ), .Y (n_543));
NOR2X1 g136177(.A (si[29]), .B (datao_2[29] ), .Y (n_701));
NOR2X1 g136205(.A (si[10]), .B (datao_1[10] ), .Y (n_571));
NAND2X1 g136492(.A (si[0]), .B (datao_1[0] ), .Y (n_430));
NOR2X1 g136106(.A (si[10]), .B (datao_2[10] ), .Y (n_1299));
NAND2X1 g136056(.A (si[23]), .B (datao_2[23] ), .Y (n_1119));
INVX1 g138004(.A (n_606), .Y (n_284));
INVX1 g137835(.A (n_578), .Y (n_1646));
NAND2X1 g136403(.A (addr_1), .B (addr_2), .Y (n_706));
NOR2X1 g136373(.A (si[24]), .B (datao_1[24] ), .Y (n_788));
NOR2X1 g136183(.A (P3_reg3[11] ), .B (P3_reg3[12] ), .Y (n_266));
INVX1 g137990(.A (n_33257), .Y (n_265));
NAND2X1 g136086(.A (si[24]), .B (datao_1[24] ), .Y (n_1576));
NAND2X1 g136324(.A (si[2]), .B (datao_2[2] ), .Y (n_1256));
NOR2X1 g136471(.A (P3_reg3[21] ), .B (P3_reg3[22] ), .Y (n_808));
INVX1 g136663(.A (n_1878), .Y (n_262));
NOR2X1 g136089(.A (P3_reg3[11] ), .B (P3_reg3[10] ), .Y (n_910));
NOR2X1 g136241(.A (si[23]), .B (datao_2[23] ), .Y (n_978));
INVX1 g137447(.A (n_629), .Y (n_2742));
AND2X1 g136404(.A (P2_reg3[22] ), .B (P2_reg3[23] ), .Y (n_1499));
NOR2X1 g136350(.A (datao_2[27] ), .B (si[27]), .Y (n_1357));
NOR2X1 g136139(.A (si[2]), .B (datao_2[2] ), .Y (n_855));
AND2X1 g136301(.A (P1_reg3[21] ), .B (P1_reg3[20] ), .Y (n_457));
NOR2X1 g136050(.A (si[24]), .B (n_667), .Y (n_1496));
OR2X1 g136272(.A (P3_reg3[7] ), .B (P3_reg3[8] ), .Y (n_247));
INVX1 g136726(.A (n_349), .Y (n_631));
NAND2X1 g136134(.A (datao_1[27] ), .B (si[27]), .Y (n_696));
OR2X1 g136322(.A (si[30]), .B (n_479), .Y (n_1838));
AND2X1 g136198(.A (P2_reg3[13] ), .B (P2_reg3[14] ), .Y (n_634));
NOR2X1 g136135(.A (P3_reg3[20] ), .B (P3_reg3[21] ), .Y (n_972));
NAND2X1 g136486(.A (si[12]), .B (n_12330), .Y (n_1141));
NOR2X1 g136268(.A (n_491), .B (si[28]), .Y (n_925));
OR2X1 g136199(.A (P3_reg3[2] ), .B (n_13675), .Y (n_237));
INVX1 g137157(.A (n_1870), .Y (n_3686));
NAND2X1 g136352(.A (si[19]), .B (datao_2[19] ), .Y (n_1508));
NAND2X1 g136158(.A (si[29]), .B (datao_2[29] ), .Y (n_1928));
NAND2X1 g136269(.A (si[23]), .B (datao_1[23] ), .Y (n_2035));
NAND2X1 g136220(.A (si[15]), .B (datao_2[15] ), .Y (n_889));
NOR2X1 g136500(.A (si[17]), .B (datao_2[17] ), .Y (n_636));
INVX1 g137868(.A (n_33587), .Y (n_826));
CLKBUFX3 g137910(.A (n_218), .Y (n_939));
NOR2X1 g136464(.A (si[16]), .B (datao_2[16] ), .Y (n_497));
NAND2X1 g136315(.A (si[4]), .B (datao_1[4] ), .Y (n_1605));
CLKBUFX1 g137962(.A (n_216), .Y (n_1753));
NAND2X1 g136046(.A (si[6]), .B (datao_2[6] ), .Y (n_949));
AND2X1 g136076(.A (P2_reg3[18] ), .B (P2_reg3[19] ), .Y (n_981));
CLKBUFX1 g137458(.A (n_203), .Y (n_1444));
CLKBUFX1 g136958(.A (n_200), .Y (n_1720));
CLKBUFX1 g137333(.A (n_33562), .Y (n_1015));
INVX1 g136753(.A (n_349), .Y (n_392));
INVX1 g136935(.A (n_453), .Y (n_516));
NOR2X1 g136374(.A (datao_2[26] ), .B (si[26]), .Y (n_1223));
NOR2X1 g136527(.A (P3_reg3[13] ), .B (P3_reg3[12] ), .Y (n_779));
NAND2X1 g136182(.A (si[0]), .B (datao_2[0] ), .Y (n_707));
NOR2X1 g136448(.A (si[22]), .B (n_12188), .Y (n_963));
NAND2X1 g136237(.A (si[10]), .B (datao_1[10] ), .Y (n_1271));
INVX1 g137639(.A (n_7967), .Y (n_8687));
INVX1 g136871(.A (n_551), .Y (n_1175));
NOR2X1 g136537(.A (P3_reg3[14] ), .B (P3_reg3[15] ), .Y (n_929));
NOR2X1 g136376(.A (si[8]), .B (datao_2[8] ), .Y (n_847));
AND2X1 g136514(.A (P1_reg3[22] ), .B (P1_reg3[23] ), .Y (n_1681));
NAND2X1 g136439(.A (si[11]), .B (n_12458), .Y (n_997));
NAND2X1 g136417(.A (P2_reg3[19] ), .B (P2_reg3[20] ), .Y (n_871));
NAND2X1 g136137(.A (P1_reg3[19] ), .B (P1_reg3[20] ), .Y (n_877));
INVX1 g137210(.A (n_499), .Y (n_7841));
NOR2X1 g136362(.A (P3_reg3[16] ), .B (P3_reg3[15] ), .Y (n_994));
NAND2X1 g136180(.A (datao_2[27] ), .B (si[27]), .Y (n_1356));
NAND2X1 g136058(.A (P2_reg3[15] ), .B (P2_reg3[14] ), .Y (n_687));
NAND2X1 g136217(.A (P2_reg3[15] ), .B (P2_reg3[16] ), .Y (n_992));
NAND2X1 g136407(.A (datao_1[28] ), .B (si[28]), .Y (n_1328));
INVX1 g138036(.A (n_452), .Y (n_1661));
NAND2X1 g136142(.A (si[25]), .B (datao_2[25] ), .Y (n_663));
INVX1 g137700(.A (n_167), .Y (n_1858));
NOR2X1 g136254(.A (si[5]), .B (datao_2[5] ), .Y (n_1162));
NOR2X1 g136218(.A (P3_reg3[24] ), .B (P3_reg3[25] ), .Y (n_3109));
NOR2X1 g136038(.A (datao_1[27] ), .B (si[27]), .Y (n_1374));
NOR2X1 g136346(.A (si[20]), .B (n_12322), .Y (n_1589));
NAND2X1 g136369(.A (si[3]), .B (datao_2[3] ), .Y (n_1087));
NOR2X1 g136113(.A (si[23]), .B (datao_1[23] ), .Y (n_962));
NAND2X1 g136325(.A (si[29]), .B (datao_1[29] ), .Y (n_1365));
INVX1 g136694(.A (n_349), .Y (n_7243));
INVX2 g137848(.A (n_377), .Y (n_852));
NAND2X1 g136114(.A (si[10]), .B (datao_2[10] ), .Y (n_1197));
NAND2X1 g136319(.A (P1_reg3[5] ), .B (P1_reg3[6] ), .Y (n_141));
NOR2X1 g136031(.A (si[9]), .B (datao_2[9] ), .Y (n_1041));
NAND2X1 g136316(.A (si[30]), .B (datao_1[30] ), .Y (n_1364));
INVX1 g136899(.A (n_33560), .Y (n_396));
NAND2X1 g136380(.A (si[8]), .B (datao_2[8] ), .Y (n_1209));
INVX1 g137588(.A (n_521), .Y (n_9672));
INVX1 g137606(.A (n_33561), .Y (n_589));
AND2X1 g136307(.A (P2_reg3[24] ), .B (P2_reg3[25] ), .Y (n_2976));
NOR2X1 g136393(.A (si[4]), .B (datao_2[4] ), .Y (n_716));
NAND2X1 g136048(.A (P2_reg3[17] ), .B (P2_reg3[18] ), .Y (n_957));
NOR2X1 g136478(.A (si[29]), .B (datao_1[29] ), .Y (n_733));
NOR2X1 g136496(.A (si[20]), .B (datao_2[20] ), .Y (n_1221));
NOR2X1 g136078(.A (P3_reg3[26] ), .B (P3_reg3[25] ), .Y (n_2085));
NAND2X1 g136196(.A (si[18]), .B (datao_2[18] ), .Y (n_896));
NAND2X1 g136099(.A (P2_reg3[23] ), .B (P2_reg3[24] ), .Y (n_710));
CLKBUFX1 g136955(.A (n_118), .Y (n_1969));
INVX1 g136633(.A (n_117), .Y (n_1218));
INVX2 g136807(.A (n_998), .Y (n_762));
NOR2X1 g136344(.A (si[25]), .B (datao_2[25] ), .Y (n_1177));
NAND2X1 g136491(.A (P2_reg3[5] ), .B (P2_reg3[6] ), .Y (n_110));
NAND2X1 g136200(.A (si[14]), .B (datao_2[14] ), .Y (n_1331));
NOR2X1 g136118(.A (si[19]), .B (datao_1[19] ), .Y (n_1375));
CLKBUFX1 g136742(.A (n_349), .Y (n_1017));
NOR2X1 g136302(.A (si[15]), .B (datao_2[15] ), .Y (n_1224));
INVX1 g137191(.A (n_647), .Y (n_653));
INVX1 g137765(.A (P2_reg3[3] ), .Y (n_7475));
INVX4 g137163(.A (n_99), .Y (n_1724));
NOR2X1 g136181(.A (P3_reg3[18] ), .B (P3_reg3[19] ), .Y (n_746));
INVX1 g136901(.A (n_432), .Y (n_9653));
NAND2X1 g136457(.A (si[7]), .B (datao_2[7] ), .Y (n_850));
NAND2X1 g136165(.A (P1_reg3[3] ), .B (P1_reg3[4] ), .Y (n_831));
NOR2X1 g136245(.A (si[1]), .B (datao_1[1] ), .Y (n_1135));
NAND2X1 g136512(.A (si[16]), .B (datao_2[16] ), .Y (n_1143));
INVX1 g136891(.A (n_498), .Y (n_8083));
NOR2X1 g136433(.A (P3_reg3[16] ), .B (P3_reg3[17] ), .Y (n_747));
NAND2X1 g136081(.A (si[9]), .B (datao_2[9] ), .Y (n_1273));
NAND2X1 g136521(.A (P1_reg3[17] ), .B (P1_reg3[18] ), .Y (n_921));
NOR2X1 g136152(.A (P3_reg3[10] ), .B (P3_reg3[7] ), .Y (n_88));
INVX1 g137995(.A (n_549), .Y (n_1624));
NOR2X1 g136072(.A (si[9]), .B (datao_1[9] ), .Y (n_1580));
NAND2X1 g136161(.A (si[4]), .B (datao_2[4] ), .Y (n_1163));
NOR2X1 g136077(.A (P3_reg3[23] ), .B (P3_reg3[22] ), .Y (n_1461));
NAND2X1 g136043(.A (P2_reg3[21] ), .B (P2_reg3[22] ), .Y (n_810));
NAND2X1 g136530(.A (si[22]), .B (datao_2[22] ), .Y (n_955));
NAND2X1 g136212(.A (si[9]), .B (datao_1[9] ), .Y (n_1297));
NOR2X1 g136229(.A (si[18]), .B (datao_2[18] ), .Y (n_1136));
NOR2X1 g136251(.A (si[21]), .B (datao_2[21] ), .Y (n_979));
INVX1 g136823(.A (n_998), .Y (n_873));
NOR2X1 g136092(.A (si[14]), .B (datao_2[14] ), .Y (n_1048));
NOR2X1 g136168(.A (si[7]), .B (datao_1[7] ), .Y (n_1420));
NOR2X1 g136159(.A (P3_reg3[27] ), .B (P3_reg3[28] ), .Y (n_74));
INVX1 g137975(.A (n_522), .Y (n_9667));
INVX1 g137911(.A (P1_IR[9] ), .Y (n_218));
INVX1 g137511(.A (addr_455), .Y (n_553));
INVX1 g136877(.A (P3_IR[21] ), .Y (n_657));
INVX1 g136904(.A (n_9663), .Y (n_410));
INVX1 g137225(.A (P1_reg3[11] ), .Y (n_2317));
INVX1 g137657(.A (P1_IR[23] ), .Y (n_211));
INVX1 g137525(.A (P3_reg3[0] ), .Y (n_72));
INVX1 g137041(.A (P3_reg3[23] ), .Y (n_343));
INVX1 g137566(.A (n_12670), .Y (n_7541));
INVX1 g137594(.A (n_7839), .Y (n_416));
INVX1 g137148(.A (P1_IR[29] ), .Y (n_252));
INVX1 g136884(.A (n_1319), .Y (n_316));
INVX1 g137898(.A (n_4344), .Y (n_103));
INVX1 g137844(.A (P3_reg3[22] ), .Y (n_165));
INVX1 g137208(.A (n_3337), .Y (n_154));
INVX1 g137244(.A (n_10435), .Y (n_77));
INVX1 g137651(.A (n_13358), .Y (n_389));
INVX1 g136792(.A (P2_reg2[15] ), .Y (n_70));
INVX1 g136836(.A (n_3314), .Y (n_69));
CLKBUFX1 g137825(.A (P3_reg1[15] ), .Y (n_13678));
INVX1 g136648(.A (n_13348), .Y (n_215));
INVX1 g137318(.A (datao_1[7] ), .Y (n_68));
INVX1 g137047(.A (addr_485), .Y (n_190));
INVX1 g137189(.A (P3_IR[14] ), .Y (n_704));
INVX1 g137228(.A (n_4231), .Y (n_174));
INVX1 g137708(.A (n_13352), .Y (n_228));
INVX1 g136623(.A (addr_442), .Y (n_147));
INVX1 g137216(.A (datao_2[0] ), .Y (n_144));
INVX1 g137557(.A (P1_reg_175), .Y (n_10225));
INVX1 g137477(.A (P2_reg_112), .Y (n_9602));
INVX1 g136887(.A (n_4230), .Y (n_151));
INVX1 g137052(.A (P2_reg3[20] ), .Y (n_586));
INVX1 g137950(.A (P3_IR[15] ), .Y (n_527));
INVX1 g137329(.A (P2_reg1[13] ), .Y (n_66));
INVX1 g137623(.A (P3_d), .Y (n_65));
INVX1 g136859(.A (P1_reg2[29] ), .Y (n_10546));
INVX1 g137661(.A (n_4215), .Y (n_191));
INVX1 g138066(.A (n_3259), .Y (n_121));
INVX1 g136640(.A (n_4475), .Y (n_235));
INVX1 g137622(.A (addr_489), .Y (n_64));
INVX1 g138033(.A (n_4237), .Y (n_207));
INVX1 g138017(.A (P3_reg3[26] ), .Y (n_3108));
INVX1 g136777(.A (P2_reg2[19] ), .Y (n_352));
INVX1 g137727(.A (P2_reg2[26] ), .Y (n_10604));
INVX1 g137486(.A (addr_436), .Y (n_62));
INVX4 g136833(.A (P1_IR[31] ), .Y (n_998));
INVX1 g136557(.A (n_9135), .Y (n_341));
INVX1 g137591(.A (n_10167), .Y (n_361));
INVX1 g137840(.A (P3_reg3[6] ), .Y (n_1027));
INVX1 g137514(.A (n_12030), .Y (n_529));
INVX1 g138071(.A (n_12322), .Y (n_547));
INVX1 g136644(.A (P2_reg3[5] ), .Y (n_339));
INVX1 g137830(.A (datao_1[1] ), .Y (n_451));
INVX1 g136959(.A (P2_IR[8] ), .Y (n_200));
INVX1 g137055(.A (datao_2[29] ), .Y (n_61));
INVX1 g137375(.A (addr_429), .Y (n_60));
INVX1 g137355(.A (P3_reg2[28] ), .Y (n_9038));
INVX1 g137747(.A (n_4920), .Y (n_322));
INVX1 g136548(.A (P3_reg_153), .Y (n_13200));
INVX1 g137668(.A (P3_reg2[29] ), .Y (n_113));
INVX1 g137484(.A (n_13342), .Y (n_79));
INVX1 g137154(.A (P3_reg3[13] ), .Y (n_272));
INVX1 g137666(.A (n_9071), .Y (n_96));
INVX1 g136610(.A (n_13515), .Y (n_4265));
INVX1 g137420(.A (P2_reg2[25] ), .Y (n_10607));
INVX1 g137736(.A (reset), .Y (n_32010));
INVX1 g137715(.A (n_693), .Y (n_528));
INVX1 g137342(.A (P3_reg_147), .Y (n_13207));
INVX1 g137698(.A (n_3709), .Y (n_143));
INVX1 g136552(.A (P2_reg1[25] ), .Y (n_9097));
INVX2 g137462(.A (P1_IR[2] ), .Y (n_1464));
INVX1 g137596(.A (addr_494), .Y (n_431));
INVX1 g137308(.A (P3_reg3[19] ), .Y (n_56));
INVX1 g136637(.A (n_12028), .Y (n_515));
INVX1 g137927(.A (P3_reg3[17] ), .Y (n_330));
INVX1 g137278(.A (n_10613), .Y (n_242));
INVX1 g138011(.A (P1_IR[30] ), .Y (n_241));
INVX1 g137459(.A (P1_IR[0] ), .Y (n_203));
INVX1 g137235(.A (n_13368), .Y (n_304));
INVX1 g137555(.A (P1_reg2[24] ), .Y (n_10858));
INVX1 g136952(.A (n_4151), .Y (n_384));
INVX1 g137266(.A (n_9675), .Y (n_411));
INVX1 g137509(.A (P1_reg3[3] ), .Y (n_7515));
INVX1 g137359(.A (P1_reg1[27] ), .Y (n_10247));
INVX1 g137059(.A (P3_reg3[18] ), .Y (n_320));
INVX1 g137615(.A (n_12319), .Y (n_625));
INVX1 g137264(.A (datao_2[19] ), .Y (n_612));
INVX1 g136786(.A (datao_1[27] ), .Y (n_54));
INVX1 g137586(.A (n_928), .Y (n_540));
INVX1 g137777(.A (n_4367), .Y (n_382));
INVX1 g137701(.A (P1_IR[6] ), .Y (n_167));
INVX1 g136902(.A (addr_495), .Y (n_432));
INVX1 g137787(.A (n_4445), .Y (n_324));
INVX1 g136892(.A (addr_456), .Y (n_498));
INVX1 g137204(.A (P2_IR[21] ), .Y (n_1236));
INVX1 g136929(.A (n_3402), .Y (n_109));
INVX1 g136896(.A (P2_IR[20] ), .Y (n_287));
INVX1 g137816(.A (P1_IR[25] ), .Y (n_799));
INVX1 g137057(.A (P2_IR[14] ), .Y (n_682));
INVX1 g136948(.A (addr_447), .Y (n_52));
INVX1 g136555(.A (P1_reg3[9] ), .Y (n_169));
INVX1 g137062(.A (P3_IR[27] ), .Y (n_593));
INVX1 g138056(.A (addr_488), .Y (n_50));
INVX1 g137986(.A (P3_reg3[27] ), .Y (n_269));
INVX1 g137710(.A (P1_IR[12] ), .Y (n_1018));
INVX1 g137761(.A (P2_reg2[12] ), .Y (n_49));
INVX1 g137681(.A (addr_444), .Y (n_130));
INVX1 g137321(.A (n_8117), .Y (n_493));
INVX1 g137632(.A (P1_reg2[27] ), .Y (n_11327));
INVX1 g138037(.A (P2_IR[16] ), .Y (n_452));
INVX1 g138005(.A (P2_IR[12] ), .Y (n_606));
INVX1 g137742(.A (n_475), .Y (n_424));
INVX1 g137239(.A (addr_487), .Y (n_46));
INVX1 g137066(.A (si[25]), .Y (n_45));
INVX1 g137694(.A (n_10610), .Y (n_335));
INVX1 g137332(.A (n_3693), .Y (n_365));
INVX1 g137419(.A (n_13361), .Y (n_363));
INVX1 g137426(.A (n_12188), .Y (n_447));
INVX1 g137577(.A (n_12022), .Y (n_455));
INVX1 g137956(.A (P3_IR[12] ), .Y (n_564));
INVX1 g137732(.A (P3_IR[19] ), .Y (n_1666));
INVX1 g137676(.A (P1_reg1[29] ), .Y (n_10245));
INVX1 g137976(.A (addr_497), .Y (n_522));
INVX1 g137280(.A (P1_IR[13] ), .Y (n_1012));
INVX1 g137809(.A (addr_443), .Y (n_10057));
INVX1 g137270(.A (n_1964), .Y (n_212));
INVX1 g137248(.A (n_3716), .Y (n_137));
INVX1 g137467(.A (n_13203), .Y (n_173));
INVX1 g137272(.A (n_12184), .Y (n_419));
INVX1 g137610(.A (P2_reg1[29] ), .Y (n_9092));
INVX1 g136874(.A (n_13215), .Y (n_336));
INVX1 g137195(.A (P3_reg_148), .Y (n_13340));
INVX1 g136774(.A (n_13366), .Y (n_4039));
INVX1 g137211(.A (addr_457), .Y (n_499));
INVX1 g137339(.A (n_9586), .Y (n_41));
INVX1 g137401(.A (n_13332), .Y (n_379));
INVX1 g137530(.A (n_4561), .Y (n_73));
INVX1 g136865(.A (P2_IR[30] ), .Y (n_100));
INVX1 g137412(.A (n_524), .Y (n_7043));
CLKBUFX1 g137728(.A (P1_reg2[0] ), .Y (n_11136));
INVX1 g136857(.A (n_4160), .Y (n_273));
INVX1 g137546(.A (P1_reg1[26] ), .Y (n_10161));
INVX1 g137967(.A (addr_435), .Y (n_40));
INVX1 g137549(.A (P3_IR[24] ), .Y (n_664));
INVX1 g137630(.A (n_3668), .Y (n_224));
INVX1 g136854(.A (n_14096), .Y (n_185));
INVX1 g136576(.A (P1_IR[21] ), .Y (n_1206));
INVX1 g137371(.A (n_13645), .Y (n_296));
INVX1 g136655(.A (n_13677), .Y (n_209));
INVX1 g137598(.A (n_9101), .Y (n_271));
INVX1 g137892(.A (n_7843), .Y (n_465));
INVX1 g138027(.A (n_13202), .Y (n_196));
INVX1 g137202(.A (P1_IR[24] ), .Y (n_658));
INVX1 g137618(.A (P3_IR[20] ), .Y (n_1323));
INVX1 g136588(.A (P2_IR[27] ), .Y (n_600));
INVX1 g137908(.A (n_3235), .Y (n_319));
INVX1 g137769(.A (P1_reg3[20] ), .Y (n_134));
INVX1 g137348(.A (n_4554), .Y (n_331));
INVX1 g136626(.A (n_13502), .Y (n_4474));
INVX1 g137674(.A (datao_1[4] ), .Y (n_585));
INVX1 g136788(.A (P1_reg_179), .Y (n_10211));
INVX1 g136762(.A (P2_reg1[9] ), .Y (n_36));
INVX1 g136568(.A (P2_reg2[28] ), .Y (n_10653));
INVX1 g137545(.A (P2_reg1[27] ), .Y (n_35));
INVX1 g137431(.A (addr_453), .Y (n_34));
INVX1 g137772(.A (n_4277), .Y (n_323));
INVX1 g136915(.A (n_10443), .Y (n_295));
INVX1 g138054(.A (P2_d_394), .Y (n_33));
INVX1 g136879(.A (n_12454), .Y (n_535));
INVX1 g137481(.A (datao_2[23] ), .Y (n_32));
INVX1 g137805(.A (n_13211), .Y (n_146));
INVX1 g137704(.A (n_3724), .Y (n_311));
INVX1 g136870(.A (P2_reg_111), .Y (n_9132));
INVX1 g137259(.A (datao_1[9] ), .Y (n_153));
INVX1 g137323(.A (n_10136), .Y (n_122));
INVX1 g137213(.A (addr_492), .Y (n_31));
INVX1 g136563(.A (addr_445), .Y (n_233));
INVX1 g137774(.A (n_10158), .Y (n_279));
INVX1 g137689(.A (n_11802), .Y (n_421));
INVX1 g137959(.A (n_13357), .Y (n_192));
INVX1 g137199(.A (P1_IR[17] ), .Y (n_984));
INVX1 g136758(.A (P3_reg3[21] ), .Y (n_307));
INVX1 g136631(.A (n_479), .Y (n_380));
INVX1 g137963(.A (P3_IR[7] ), .Y (n_216));
INVX2 g137174(.A (P3_IR[31] ), .Y (n_99));
INVX1 g137613(.A (n_4213), .Y (n_164));
INVX1 g136652(.A (n_9231), .Y (n_309));
INVX1 g137918(.A (n_13201), .Y (n_127));
INVX1 g137993(.A (addr_484), .Y (n_2772));
INVX1 g137490(.A (datao_1[0] ), .Y (n_275));
INVX1 g137261(.A (si[23]), .Y (n_28));
INVX1 g137218(.A (P1_reg3[5] ), .Y (n_830));
INVX1 g137795(.A (n_4534), .Y (n_198));
INVX1 g138030(.A (P3_IR[25] ), .Y (n_282));
INVX1 g137904(.A (P2_IR[29] ), .Y (n_2504));
INVX1 g137792(.A (P2_reg_110), .Y (n_9178));
INVX1 g136956(.A (P1_IR[7] ), .Y (n_118));
INVX1 g137049(.A (P3_reg3[25] ), .Y (n_158));
INVX1 g137790(.A (P1_IR[16] ), .Y (n_488));
INVX1 g137534(.A (n_4477), .Y (n_182));
INVX1 g136798(.A (P1_reg1[25] ), .Y (n_10215));
INVX1 g136764(.A (n_8074), .Y (n_464));
INVX1 g137834(.A (n_13359), .Y (n_261));
INVX2 g137448(.A (P1_IR[8] ), .Y (n_629));
INVX1 g137895(.A (n_13337), .Y (n_289));
INVX1 g136941(.A (P3_reg3[20] ), .Y (n_354));
INVX1 g137520(.A (n_13334), .Y (n_267));
INVX1 g137379(.A (n_804), .Y (n_492));
INVX2 g137220(.A (P2_IR[10] ), .Y (n_1799));
INVX1 g137692(.A (P3_reg_146), .Y (n_13205));
INVX1 g137932(.A (n_482), .Y (n_637));
INVX1 g137537(.A (addr_483), .Y (n_11097));
INVX1 g136866(.A (P2_reg_109), .Y (n_9794));
CLKBUFX1 g136614(.A (P3_reg1[5] ), .Y (n_13683));
INVX1 g136768(.A (P3_IR[23] ), .Y (n_545));
INVX1 g136868(.A (addr_430), .Y (n_25));
INVX1 g137313(.A (P3_reg_152), .Y (n_13373));
INVX1 g137823(.A (n_481), .Y (n_1787));
INVX1 g137460(.A (P2_reg1[26] ), .Y (n_9142));
INVX1 g137887(.A (n_13680), .Y (n_3848));
INVX1 g138024(.A (P3_IR[17] ), .Y (n_684));
INVX1 g137579(.A (n_12026), .Y (n_393));
INVX1 g137836(.A (P1_IR[14] ), .Y (n_578));
INVX1 g136839(.A (n_10566), .Y (n_149));
INVX1 g137937(.A (n_565), .Y (n_286));
INVX1 g137223(.A (n_13343), .Y (n_333));
INVX1 g137735(.A (P2_reg1[28] ), .Y (n_9081));
INVX1 g137784(.A (P1_IR[26] ), .Y (n_686));
INVX1 g137325(.A (P1_reg3[17] ), .Y (n_202));
INVX1 g137589(.A (addr_496), .Y (n_521));
INVX1 g136608(.A (n_13365), .Y (n_168));
INVX1 g138063(.A (n_9597), .Y (n_101));
INVX1 g137721(.A (P2_IR[13] ), .Y (n_764));
INVX1 g136872(.A (P2_IR[11] ), .Y (n_551));
INVX1 g137946(.A (P3_reg_149), .Y (n_13206));
INVX1 g138042(.A (P1_IR[11] ), .Y (n_668));
INVX1 g137978(.A (addr_432), .Y (n_22));
INVX1 g137832(.A (P1_reg2[26] ), .Y (n_10886));
INVX1 g137899(.A (addr_439), .Y (n_21));
INVX1 g136852(.A (P1_IR[10] ), .Y (n_1968));
INVX1 g137602(.A (n_491), .Y (n_116));
INVX1 g138021(.A (n_641), .Y (n_138));
INVX1 g137718(.A (n_3958), .Y (n_362));
INVX1 g137922(.A (addr_461), .Y (n_194));
INVX2 g137192(.A (P1_IR[3] ), .Y (n_647));
INVX1 g137470(.A (n_13344), .Y (n_318));
INVX1 g136917(.A (P3_reg3[15] ), .Y (n_231));
INVX1 g138001(.A (n_628), .Y (n_415));
INVX1 g136605(.A (P2_reg_113), .Y (n_9088));
INVX1 g137151(.A (P1_IR[28] ), .Y (n_1107));
INVX1 g136910(.A (addr_2), .Y (n_263));
INVX1 g138044(.A (P1_reg_176), .Y (n_10134));
INVX1 g137996(.A (P2_IR[18] ), .Y (n_549));
INVX1 g137838(.A (n_10893), .Y (n_372));
INVX1 g137303(.A (n_13507), .Y (n_115));
INVX1 g137518(.A (P2_reg3[21] ), .Y (n_19));
INVX1 g138076(.A (P1_IR[18] ), .Y (n_120));
INVX1 g137913(.A (n_11120), .Y (n_142));
INVX1 g137145(.A (P1_reg_177), .Y (n_10219));
INVX1 g137757(.A (P2_reg3[23] ), .Y (n_238));
INVX1 g136670(.A (P2_IR[24] ), .Y (n_561));
INVX1 g137947(.A (P3_reg3[16] ), .Y (n_17));
INVX1 g137446(.A (n_13679), .Y (n_274));
INVX1 g137527(.A (n_13336), .Y (n_387));
INVX1 g136943(.A (P3_reg3[10] ), .Y (n_301));
INVX1 g136551(.A (n_11148), .Y (n_381));
INVX1 g137797(.A (n_9549), .Y (n_288));
INVX1 g137393(.A (n_13335), .Y (n_338));
INVX1 g136573(.A (P2_IR[23] ), .Y (n_367));
INVX1 g137751(.A (n_10165), .Y (n_83));
INVX1 g137686(.A (datao_1[5] ), .Y (n_602));
INVX1 g137543(.A (P3_reg_150), .Y (n_13204));
INVX1 g138007(.A (n_13377), .Y (n_373));
INVX1 g137307(.A (P2_IR[19] ), .Y (n_607));
INVX1 g136619(.A (n_13498), .Y (n_300));
INVX1 g137827(.A (P1_reg2[16] ), .Y (n_230));
INVX1 g137814(.A (P3_reg1[26] ), .Y (n_290));
INVX1 g137779(.A (P2_IR[26] ), .Y (n_1304));
INVX1 g138069(.A (P2_reg2[8] ), .Y (n_15));
INVX1 g136946(.A (n_13511), .Y (n_204));
INVX1 g136968(.A (n_13351), .Y (n_229));
INVX1 g137643(.A (P2_reg1[19] ), .Y (n_358));
INVX1 g136600(.A (P3_IR[30] ), .Y (n_594));
INVX1 g137365(.A (P1_reg1[28] ), .Y (n_10169));
INVX1 g136613(.A (n_4590), .Y (n_85));
INVX1 g136771(.A (P3_reg_151), .Y (n_13199));
INVX1 g137065(.A (n_3333), .Y (n_210));
INVX1 g138040(.A (n_3565), .Y (n_277));
INVX1 g137251(.A (P1_reg3[6] ), .Y (n_327));
INVX1 g136919(.A (P1_IR[15] ), .Y (n_1171));
INVX1 g137344(.A (P3_reg3[7] ), .Y (n_2105));
INVX1 g137285(.A (n_732), .Y (n_294));
INVX1 g137989(.A (n_10897), .Y (n_225));
INVX1 g137646(.A (P2_reg2[29] ), .Y (n_8011));
INVX1 g137574(.A (datao_1[11] ), .Y (n_13));
INVX1 g138048(.A (P1_IR[20] ), .Y (n_345));
INVX1 g137551(.A (n_13681), .Y (n_4132));
INVX1 g137940(.A (n_9475), .Y (n_94));
INVX1 g137197(.A (P3_IR[26] ), .Y (n_727));
INVX1 g137568(.A (n_9658), .Y (n_1711));
INVX1 g137233(.A (addr_446), .Y (n_11));
INVX1 g136582(.A (n_667), .Y (n_171));
INVX1 g137300(.A (P1_IR[19] ), .Y (n_739));
INVX1 g137391(.A (P3_B), .Y (n_1054));
INVX1 g137744(.A (n_9655), .Y (n_442));
INVX1 g137257(.A (addr_3), .Y (n_10838));
INVX1 g136584(.A (n_10217), .Y (n_201));
INVX1 g138058(.A (P1_reg2[25] ), .Y (n_10890));
INVX1 g136794(.A (P3_reg3[24] ), .Y (n_188));
INVX1 g137414(.A (P2_reg3[10] ), .Y (n_334));
INVX1 g136665(.A (P3_IR[22] ), .Y (n_1878));
INVX1 g137807(.A (n_13341), .Y (n_346));
INVX1 g137653(.A (addr_438), .Y (n_10));
INVX1 g136662(.A (n_3470), .Y (n_148));
INVX1 g137570(.A (n_8361), .Y (n_649));
INVX1 g137627(.A (n_9634), .Y (n_95));
INVX1 g137664(.A (n_13355), .Y (n_375));
INVX1 g137242(.A (P3_IR[16] ), .Y (n_439));
INVX1 g137726(.A (P3_IR[28] ), .Y (n_1369));
INVX1 g137754(.A (n_3416), .Y (n_243));
INVX1 g137361(.A (P1_reg1[16] ), .Y (n_75));
INVX1 g137706(.A (n_13353), .Y (n_303));
INVX1 g137353(.A (P3_IR[18] ), .Y (n_943));
INVX1 g137434(.A (n_13721), .Y (n_376));
INVX1 g137315(.A (P2_reg3[11] ), .Y (n_2213));
INVX1 g137237(.A (n_13354), .Y (n_268));
INVX1 g138061(.A (P3_reg_145), .Y (n_13208));
INVX1 g137398(.A (P1_reg2[28] ), .Y (n_11144));
INVX1 g137291(.A (n_1170), .Y (n_126));
INVX1 g137407(.A (n_13367), .Y (n_156));
INVX1 g136907(.A (n_4824), .Y (n_114));
INVX1 g137802(.A (P2_IR[15] ), .Y (n_632));
INVX2 g137855(.A (P2_IR[31] ), .Y (n_377));
INVX1 g136926(.A (n_11141), .Y (n_7));
INVX1 g136965(.A (P2_IR[25] ), .Y (n_150));
INVX1 g137424(.A (n_4011), .Y (n_172));
INVX1 g136846(.A (P2_IR[28] ), .Y (n_366));
INVX1 g137296(.A (n_10223), .Y (n_4045));
INVX1 g136668(.A (n_13338), .Y (n_205));
INVX1 g136936(.A (P2_IR[17] ), .Y (n_453));
INVX1 g137953(.A (P3_reg3[28] ), .Y (n_259));
INVX1 g136544(.A (n_1976), .Y (n_125));
INVX1 g137156(.A (P1_reg_178), .Y (n_10152));
INVX1 g138014(.A (n_13212), .Y (n_388));
INVX1 g137943(.A (P1_IR[22] ), .Y (n_1401));
INVX1 g137337(.A (P3_reg3[12] ), .Y (n_1032));
CLKBUFX1 g137695(.A (P3_reg1[12] ), .Y (n_13709));
INVX1 g137317(.A (addr_434), .Y (n_6));
INVX1 g137620(.A (n_10562), .Y (n_5));
INVX1 g136672(.A (P1_IR[27] ), .Y (n_1890));
INVX1 g137421(.A (P2_reg2[24] ), .Y (n_10082));
INVX1 g137043(.A (addr_454), .Y (n_552));
INVX1 g136889(.A (addr_441), .Y (n_680));
INVX1 g137965(.A (addr_437), .Y (n_3));
INVX2 g136634(.A (P3_IR[6] ), .Y (n_117));
INVX1 g136923(.A (n_13329), .Y (n_5289));
INVX1 g136938(.A (P3_reg3[9] ), .Y (n_1031));
INVX1 g137416(.A (P1_reg3[8] ), .Y (n_321));
INVX1 g138067(.A (P3_reg3[11] ), .Y (n_2));
INVX1 g138079(.A (P2_reg2[27] ), .Y (n_10602));
INVX1 g136602(.A (datao_1[10] ), .Y (n_1));
INVX1 g137159(.A (P3_IR[31] ), .Y (n_1870));
INVX1 g137915(.A (addr_433), .Y (n_0));
INVX1 g137640(.A (P2_B), .Y (n_7967));
INVX1 g138783(.A (n_33141), .Y (n_32321));
INVX1 g138798(.A (n_32340), .Y (n_32339));
INVX1 g138799(.A (n_32342), .Y (n_32341));
CLKBUFX1 g138800(.A (n_32343), .Y (n_32342));
INVX1 g138805(.A (n_32350), .Y (n_32349));
CLKBUFX1 g138810(.A (n_32356), .Y (n_32350));
INVX1 g138812(.A (n_32344), .Y (n_32356));
INVX1 g138813(.A (n_9733), .Y (n_32344));
INVX1 g138814(.A (n_32359), .Y (n_32358));
CLKBUFX3 g138816(.A (n_32362), .Y (n_32361));
INVX1 g138817(.A (n_32364), .Y (n_32363));
CLKBUFX1 g138818(.A (n_32366), .Y (n_32364));
INVX1 g138819(.A (n_32366), .Y (n_32365));
INVX1 g138820(.A (n_32368), .Y (n_32367));
CLKBUFX1 g138821(.A (n_32369), .Y (n_32368));
INVX2 g138822(.A (n_1940), .Y (n_32369));
INVX1 g138824(.A (n_32373), .Y (n_32371));
INVX1 g138826(.A (n_32374), .Y (n_32373));
INVX1 g138827(.A (n_33239), .Y (n_32375));
CLKBUFX1 g138829(.A (n_32379), .Y (n_32378));
INVX1 g138831(.A (n_32382), .Y (n_32381));
INVX1 g138835(.A (n_32388), .Y (n_32386));
CLKBUFX3 g138842(.A (n_32394), .Y (n_32388));
INVX2 g138843(.A (n_3961), .Y (n_32394));
INVX1 g138844(.A (n_32397), .Y (n_32395));
CLKBUFX1 g138846(.A (n_32398), .Y (n_32397));
CLKBUFX2 g138847(.A (n_32399), .Y (n_32398));
INVX2 g138848(.A (P1_IR[1] ), .Y (n_32399));
INVX1 g138849(.A (n_32401), .Y (n_32400));
CLKBUFX1 g138850(.A (n_35384), .Y (n_32401));
INVX1 g138856(.A (n_29845), .Y (n_32409));
CLKBUFX1 g138858(.A (n_32412), .Y (n_32411));
INVX1 g138863(.A (n_32428), .Y (n_32417));
INVX1 g138871(.A (n_32428), .Y (n_32426));
CLKBUFX1 g138873(.A (n_32429), .Y (n_32428));
INVX1 g138874(.A (n_32430), .Y (n_32429));
INVX2 g138875(.A (n_32432), .Y (n_32430));
INVX1 g138876(.A (n_32432), .Y (n_32431));
CLKBUFX1 g138877(.A (n_34807), .Y (n_32433));
INVX1 g138878(.A (n_33573), .Y (n_32435));
INVX1 g138885(.A (n_32445), .Y (n_32442));
CLKBUFX1 g138889(.A (n_33573), .Y (n_32445));
CLKBUFX1 g138890(.A (n_32449), .Y (n_32448));
INVX1 g138891(.A (n_1465), .Y (n_32449));
INVX2 g138892(.A (n_32452), .Y (n_32450));
INVX2 g138894(.A (n_32453), .Y (n_32452));
INVX1 g138906(.A (n_32475), .Y (n_32473));
CLKBUFX1 g138908(.A (n_32476), .Y (n_32475));
INVX1 g138909(.A (P1_IR[5] ), .Y (n_32476));
INVX1 g138911(.A (n_32480), .Y (n_32479));
CLKBUFX1 g138912(.A (n_32481), .Y (n_32480));
INVX1 g138913(.A (n_32483), .Y (n_32482));
CLKBUFX1 g138914(.A (n_32484), .Y (n_32483));
INVX1 g138915(.A (n_32486), .Y (n_32485));
CLKBUFX1 g138916(.A (n_32487), .Y (n_32486));
CLKBUFX2 g138917(.A (n_32488), .Y (n_32487));
INVX2 g138918(.A (P1_IR[4] ), .Y (n_32488));
INVX2 g138919(.A (n_32501), .Y (n_32489));
INVX1 g138920(.A (n_32496), .Y (n_32490));
CLKBUFX1 g138929(.A (n_32500), .Y (n_32496));
CLKBUFX1 g138930(.A (n_32501), .Y (n_32500));
INVX2 g138933(.A (n_32517), .Y (n_32505));
INVX1 g138937(.A (n_32517), .Y (n_32509));
CLKBUFX1 g138956(.A (n_34320), .Y (n_32517));
INVX1 g138960(.A (n_32535), .Y (n_32533));
CLKBUFX1 g138962(.A (n_32537), .Y (n_32535));
INVX1 g138964(.A (n_16279), .Y (n_32537));
CLKBUFX3 g138966(.A (n_35166), .Y (n_32543));
CLKBUFX3 g138967(.A (n_35165), .Y (n_32544));
INVX4 g138968(.A (n_32552), .Y (n_32548));
INVX2 g138969(.A (n_32552), .Y (n_32550));
INVX2 g138971(.A (n_35165), .Y (n_32552));
CLKBUFX1 g138983(.A (n_32639), .Y (n_32637));
CLKBUFX1 g138986(.A (n_32642), .Y (n_32641));
INVX2 g138987(.A (n_4365), .Y (n_32642));
INVX1 g138988(.A (n_32646), .Y (n_32644));
CLKBUFX3 g138991(.A (n_32648), .Y (n_32646));
CLKBUFX2 g138992(.A (n_32648), .Y (n_32649));
CLKBUFX3 g138993(.A (n_32710), .Y (n_32648));
INVX1 g138995(.A (n_32654), .Y (n_32652));
INVX4 g138997(.A (n_32683), .Y (n_32654));
INVX2 g139004(.A (n_32664), .Y (n_32662));
INVX4 g139009(.A (n_32675), .Y (n_32664));
INVX1 g139010(.A (n_32664), .Y (n_32669));
INVX1 g139012(.A (n_32664), .Y (n_32673));
INVX1 g139016(.A (n_32664), .Y (n_32677));
INVX2 g139021(.A (n_32683), .Y (n_32675));
INVX2 g139022(.A (n_32710), .Y (n_32683));
INVX4 g139027(.A (n_32707), .Y (n_32685));
INVX1 g139028(.A (n_32685), .Y (n_32690));
INVX2 g139034(.A (n_32698), .Y (n_32697));
INVX4 g139035(.A (n_32685), .Y (n_32698));
CLKBUFX3 g139042(.A (n_32710), .Y (n_32707));
CLKBUFX1 g139043(.A (n_32710), .Y (n_32709));
CLKBUFX3 g139044(.A (n_32710), .Y (n_32711));
INVX4 g139045(.A (n_32818), .Y (n_32710));
INVX1 g139049(.A (n_32718), .Y (n_32715));
CLKBUFX1 g139050(.A (n_32719), .Y (n_32718));
INVX1 g139053(.A (n_32720), .Y (n_32723));
CLKBUFX3 g139055(.A (n_32719), .Y (n_32720));
INVX2 g139056(.A (n_32745), .Y (n_32728));
INVX4 g139064(.A (n_32745), .Y (n_32739));
INVX4 g139068(.A (n_32746), .Y (n_32745));
INVX2 g139069(.A (n_32719), .Y (n_32746));
INVX2 g139070(.A (n_32818), .Y (n_32719));
INVX2 g139072(.A (n_32764), .Y (n_32748));
INVX1 g139087(.A (n_32764), .Y (n_32765));
INVX4 g139088(.A (n_32767), .Y (n_32764));
INVX4 g139089(.A (n_32768), .Y (n_32767));
CLKBUFX1 g139090(.A (n_32767), .Y (n_32770));
INVX2 g139092(.A (n_32817), .Y (n_32768));
INVX1 g139095(.A (n_32777), .Y (n_32774));
INVX4 g139102(.A (n_32791), .Y (n_32777));
INVX1 g139104(.A (n_32786), .Y (n_32784));
CLKBUFX3 g139107(.A (n_32777), .Y (n_32786));
CLKBUFX3 g139110(.A (n_32817), .Y (n_32791));
INVX4 g139115(.A (n_32802), .Y (n_32794));
INVX2 g139118(.A (n_32802), .Y (n_32798));
INVX4 g139119(.A (n_32794), .Y (n_32803));
INVX1 g139127(.A (n_32815), .Y (n_32812));
INVX2 g139129(.A (n_32802), .Y (n_32815));
CLKBUFX3 g139130(.A (n_32817), .Y (n_32802));
INVX2 g139131(.A (n_32818), .Y (n_32817));
INVX4 g139132(.A (n_13066), .Y (n_32818));
BUFX3 g139138(.A (n_32834), .Y (n_32827));
CLKBUFX2 g139139(.A (n_32835), .Y (n_32834));
INVX1 g139140(.A (n_32837), .Y (n_32836));
CLKBUFX2 g139141(.A (n_32838), .Y (n_32837));
CLKBUFX2 g139142(.A (n_32839), .Y (n_32838));
INVX1 g139144(.A (n_33092), .Y (n_32841));
INVX1 g139145(.A (n_32844), .Y (n_32843));
CLKBUFX1 g139146(.A (n_33648), .Y (n_32844));
INVX1 g139147(.A (n_33648), .Y (n_32845));
INVX1 g139149(.A (n_20921), .Y (n_32847));
CLKBUFX1 g139150(.A (n_32851), .Y (n_32850));
INVX2 g139155(.A (n_32857), .Y (n_32856));
INVX2 g139156(.A (n_32858), .Y (n_32857));
INVX2 g139157(.A (n_32859), .Y (n_32858));
INVX2 g139158(.A (n_32334), .Y (n_32859));
INVX1 g139161(.A (n_32867), .Y (n_32864));
CLKBUFX2 g139164(.A (n_32868), .Y (n_32867));
CLKBUFX2 g139165(.A (n_32870), .Y (n_32869));
INVX1 g139166(.A (n_32928), .Y (n_32927));
CLKBUFX1 g139167(.A (n_32929), .Y (n_32928));
INVX2 g139168(.A (P2_IR[1] ), .Y (n_32929));
INVX1 g139169(.A (n_32932), .Y (n_32930));
CLKBUFX1 g139171(.A (n_32933), .Y (n_32932));
INVX1 g139172(.A (n_32935), .Y (n_32934));
INVX2 g139173(.A (n_13410), .Y (n_32936));
INVX1 g139174(.A (n_32941), .Y (n_32938));
CLKBUFX1 g139177(.A (n_34323), .Y (n_32941));
INVX1 g139180(.A (n_32945), .Y (n_32944));
CLKBUFX1 g139181(.A (n_34933), .Y (n_32945));
INVX1 g139183(.A (n_32949), .Y (n_32947));
INVX1 g139185(.A (n_32951), .Y (n_32950));
INVX1 g139187(.A (n_32956), .Y (n_32954));
INVX2 g139189(.A (n_32957), .Y (n_32956));
INVX2 g139190(.A (P3_IR[2] ), .Y (n_32957));
INVX1 g139192(.A (n_16772), .Y (n_32959));
INVX1 g139199(.A (n_19331), .Y (n_32967));
CLKBUFX1 g139200(.A (n_32969), .Y (n_32968));
CLKBUFX1 g139201(.A (n_32971), .Y (n_32970));
INVX1 g139206(.A (n_32978), .Y (n_32977));
CLKBUFX1 g139207(.A (n_32979), .Y (n_32978));
INVX1 g139209(.A (n_32995), .Y (n_32982));
INVX1 g139218(.A (n_32984), .Y (n_32992));
CLKBUFX1 g139219(.A (n_32995), .Y (n_32984));
INVX4 g139227(.A (n_33004), .Y (n_33000));
INVX2 g139228(.A (n_33006), .Y (n_33004));
INVX1 g139230(.A (n_33007), .Y (n_33006));
INVX1 g139236(.A (n_33025), .Y (n_33024));
CLKBUFX1 g139237(.A (n_33027), .Y (n_33025));
INVX1 g139238(.A (n_33027), .Y (n_33026));
INVX1 g139242(.A (n_33032), .Y (n_33031));
CLKBUFX3 g139243(.A (n_34999), .Y (n_33032));
INVX1 g139244(.A (n_33042), .Y (n_33034));
CLKBUFX1 g139255(.A (n_33046), .Y (n_33042));
INVX2 g139256(.A (n_34440), .Y (n_33046));
INVX2 g139264(.A (n_33071), .Y (n_33068));
CLKBUFX1 g139266(.A (n_33072), .Y (n_33071));
NAND4X1 g37(.A (n_33078), .B (n_33082), .C (n_32606), .D (n_33085),.Y (n_33086));
AOI21X1 g39(.A0 (n_14679), .A1 (n_15413), .B0 (n_33077), .Y(n_33078));
INVX1 g45(.A (n_32607), .Y (n_33077));
AND2X1 g38(.A (n_33079), .B (n_33081), .Y (n_33082));
NAND2X1 g43(.A (n_30079), .B (n_8954), .Y (n_33079));
NOR2X1 g40(.A (n_33080), .B (n_20123), .Y (n_33081));
AND2X1 g42(.A (n_14810), .B (n_13689), .Y (n_33080));
OR2X1 g41(.A (n_25881), .B (n_33084), .Y (n_33085));
INVX1 g44(.A (n_30079), .Y (n_33084));
NAND3X1 g48(.A (n_35286), .B (n_35287), .C (n_33091), .Y (n_33092));
NAND3X1 g52(.A (n_22870), .B (n_22887), .C (n_22888), .Y (n_35287));
NAND4X1 g49(.A (n_33088), .B (n_24915), .C (n_24170), .D (n_33089),.Y (n_35286));
OAI21X1 g50(.A0 (n_21087), .A1 (n_21085), .B0 (n_26641), .Y(n_33088));
AND2X1 g53(.A (n_22564), .B (n_22501), .Y (n_33089));
NAND3X1 g51(.A (n_23236), .B (n_22851), .C (n_24170), .Y (n_33091));
NOR2X1 g139267(.A (n_33093), .B (n_33098), .Y (n_33099));
NOR2X1 g34(.A (n_12690), .B (n_35315), .Y (n_33093));
OAI21X1 g139268(.A0 (n_12789), .A1 (n_33095), .B0 (n_33097), .Y(n_33098));
OR2X1 g139269(.A (n_33094), .B (n_16419), .Y (n_33095));
NOR2X1 g33(.A (n_7793), .B (n_7457), .Y (n_33094));
NAND3X1 g139270(.A (n_12789), .B (n_16419), .C (n_8124), .Y(n_33097));
NAND3X1 g139279(.A (n_33401), .B (n_34408), .C (n_34410), .Y(n_33110));
INVX1 g139280(.A (n_34405), .Y (n_33111));
INVX1 g139281(.A (n_33112), .Y (n_33113));
NAND2X1 g48_dup(.A (n_34321), .B (n_34201), .Y (n_33112));
OAI21X1 g139282(.A0 (n_33117), .A1 (n_33121), .B0 (n_33123), .Y(n_33124));
NAND3X1 g139283(.A (n_33114), .B (n_33115), .C (n_33116), .Y(n_33117));
INVX1 g139284(.A (n_28762), .Y (n_33114));
INVX1 g139285(.A (n_28748), .Y (n_33115));
AND2X1 g139286(.A (n_19849), .B (n_27611), .Y (n_33116));
NAND2X1 g139287(.A (n_33118), .B (n_33120), .Y (n_33121));
INVX1 g139288(.A (n_28186), .Y (n_33118));
NOR2X1 g139289(.A (n_33119), .B (n_29240), .Y (n_33120));
NAND2X1 g139290(.A (n_9534), .B (n_9019), .Y (n_33119));
BUFX3 g139291(.A (n_30099), .Y (n_33123));
AND2X1 g139292(.A (n_7970), .B (n_6354), .Y (n_30099));
INVX4 g139293(.A (n_30099), .Y (n_33125));
NAND4X1 g139294(.A (n_35249), .B (n_35250), .C (n_33131), .D(n_33132), .Y (n_33133));
AOI21X1 g139295(.A0 (n_20694), .A1 (n_21658), .B0 (n_28664), .Y(n_35250));
NOR2X1 g139296(.A (n_33127), .B (n_30208), .Y (n_35249));
NOR2X1 g139297(.A (n_34719), .B (n_30203), .Y (n_33127));
NAND2X1 g139298(.A (n_33129), .B (n_33546), .Y (n_33131));
NAND2X2 g139299(.A (n_29596), .B (n_14117), .Y (n_33129));
NAND2X1 g139301(.A (n_33129), .B (n_30180), .Y (n_33132));
AOI22X1 g139302(.A0 (n_33136), .A1 (n_33566), .B0 (P3_IR[31] ), .B1(n_33139), .Y (n_33140));
INVX1 g139303(.A (n_33135), .Y (n_33136));
CLKBUFX1 g139304(.A (n_34850), .Y (n_33135));
XOR2X1 g139307(.A (n_33135), .B (n_33138), .Y (n_33139));
NOR2X1 g33_dup(.A (n_34203), .B (n_34324), .Y (n_33138));
NOR2X1 g139309(.A (n_34203), .B (n_34324), .Y (n_33141));
NAND4X1 g60(.A (n_35255), .B (n_33161), .C (n_35256), .D (n_35168),.Y (n_33170));
NOR2X1 g70(.A (n_33156), .B (n_33157), .Y (n_35256));
NAND2X1 g73(.A (n_1891), .B (n_1718), .Y (n_33156));
NOR2X1 g72(.A (n_998), .B (n_3977), .Y (n_33157));
NAND2X1 g75(.A (n_33159), .B (n_1124), .Y (n_33161));
INVX1 g80(.A (n_4159), .Y (n_33159));
NOR2X1 g77(.A (n_2779), .B (n_4325), .Y (n_35255));
NAND2X1 g63(.A (n_33167), .B (n_33052), .Y (n_33168));
INVX1 g64(.A (n_33166), .Y (n_33167));
NAND2X1 g65(.A (n_33163), .B (n_33165), .Y (n_33166));
NAND2X1 g76(.A (n_3321), .B (n_1124), .Y (n_33163));
AND2X1 g69(.A (n_33053), .B (n_33164), .Y (n_33165));
NAND2X1 g74(.A (n_998), .B (P1_IR[24] ), .Y (n_33164));
AND2X1 g66(.A (n_33161), .B (n_1891), .Y (n_6069));
AND2X1 g67(.A (n_33172), .B (n_1718), .Y (n_33173));
INVX1 g71(.A (n_33157), .Y (n_33172));
INVX1 g78(.A (n_33174), .Y (n_33175));
NAND2X1 g79(.A (n_33052), .B (n_33053), .Y (n_33174));
AND2X1 g68(.A (n_33163), .B (n_33164), .Y (n_33176));
INVX1 g139315(.A (n_22530), .Y (n_33180));
INVX1 g139316(.A (n_21472), .Y (n_33181));
INVX1 g139317(.A (n_20494), .Y (n_33183));
INVX1 g36(.A (n_33184), .Y (n_33185));
OAI21X1 g139318(.A0 (n_20342), .A1 (n_20341), .B0 (n_20254), .Y(n_33184));
NAND2X1 g55(.A (n_33195), .B (n_33199), .Y (n_33200));
NAND4X1 g57(.A (n_33188), .B (n_9310), .C (n_34706), .D (n_33194), .Y(n_33195));
NAND3X1 g139319(.A (n_31049), .B (n_31023), .C (n_30533), .Y(n_33188));
INVX1 g139324(.A (P2_n_749), .Y (n_33194));
AOI21X1 g56(.A0 (n_6631), .A1 (n_9081), .B0 (n_33198), .Y (n_33199));
NOR2X1 g58(.A (n_33197), .B (n_9310), .Y (n_33198));
NAND2X1 g59(.A (n_33196), .B (n_33194), .Y (n_33197));
NOR2X1 g139325(.A (P2_reg1[28] ), .B (n_35007), .Y (n_33196));
INVX1 g139326(.A (n_33194), .Y (n_33201));
NAND2X1 g139329(.A (n_33213), .B (n_33217), .Y (n_33218));
NAND3X1 g139330(.A (n_33209), .B (n_8719), .C (n_34308), .Y(n_33213));
NAND2X1 g139331(.A (n_30772), .B (n_30007), .Y (n_33209));
NOR2X1 g139335(.A (n_33214), .B (n_33216), .Y (n_33217));
AND2X1 g139336(.A (n_6429), .B (n_10604), .Y (n_33214));
NOR2X1 g139337(.A (n_33215), .B (n_8790), .Y (n_33216));
OR2X1 g139338(.A (P2_n_749), .B (n_9934), .Y (n_33215));
NAND4X1 g139340(.A (n_33220), .B (n_33221), .C (n_33222), .D(n_33226), .Y (n_33227));
NAND2X1 g139341(.A (n_8163), .B (n_9337), .Y (n_33220));
NAND2X1 g139342(.A (n_7930), .B (P2_reg1[16] ), .Y (n_33221));
NAND2X1 g139343(.A (n_8335), .B (n_9565), .Y (n_33222));
NAND2X1 g139344(.A (n_33225), .B (P2_reg2[16] ), .Y (n_33226));
INVX2 g139345(.A (n_33265), .Y (n_33225));
INVX1 g139348(.A (n_33225), .Y (n_33228));
MX2X1 g17(.A (n_33231), .B (n_33230), .S0 (n_33232), .Y (n_33233));
INVX1 g19(.A (n_33230), .Y (n_33231));
OR2X1 g20(.A (n_19031), .B (n_18373), .Y (n_33230));
NAND2X1 g18(.A (n_22620), .B (n_23483), .Y (n_33232));
AND2X1 g139350(.A (n_35285), .B (n_35225), .Y (n_33237));
NOR2X1 g139351(.A (n_33234), .B (n_33563), .Y (n_35285));
NAND2X1 g139352(.A (n_33257), .B (n_33918), .Y (n_33234));
NAND2X1 g139354(.A (n_35224), .B (n_33238), .Y (n_33239));
INVX1 g139355(.A (n_33234), .Y (n_33238));
NAND3X1 g139359(.A (n_3932), .B (n_609), .C (n_1382), .Y (n_33242));
NAND4X1 g139361(.A (n_4757), .B (n_4198), .C (n_4528), .D (n_4516),.Y (n_33243));
NAND4X1 g139362(.A (n_4608), .B (n_4349), .C (n_33246), .D (n_4174),.Y (n_33247));
INVX1 g54(.A (n_33245), .Y (n_33246));
NAND3X1 g139363(.A (n_3837), .B (n_33244), .C (n_35380), .Y(n_33245));
NOR2X1 g139364(.A (n_3472), .B (n_3212), .Y (n_33244));
INVX1 g139365(.A (n_33242), .Y (n_33250));
INVX1 g139375(.A (P2_IR[3] ), .Y (n_33257));
INVX1 g139376(.A (n_33918), .Y (n_33261));
NAND2X2 g139378(.A (n_33264), .B (n_33267), .Y (n_33268));
AOI22X1 g139379(.A0 (n_7213), .A1 (P2_reg3[1] ), .B0 (n_7221), .B1(n_10452), .Y (n_33264));
AOI22X1 g139380(.A0 (P2_reg1[1] ), .A1 (n_7255), .B0 (n_33225), .B1(P2_reg2[1] ), .Y (n_33267));
NAND2X1 g33_dup139382(.A (n_35655), .B (n_6848), .Y (n_33265));
NAND2X1 g139383(.A (n_35656), .B (n_6848), .Y (n_33269));
NAND2X2 g21(.A (n_33270), .B (n_33273), .Y (n_33274));
NAND2X1 g139385(.A (n_16791), .B (n_18421), .Y (n_33270));
NAND2X1 g23(.A (n_33272), .B (n_32141), .Y (n_33273));
INVX1 g139386(.A (n_33271), .Y (n_33272));
NAND2X1 g139387(.A (n_32142), .B (n_22214), .Y (n_33271));
NAND3X1 g22(.A (n_33275), .B (n_32141), .C (n_33276), .Y (n_33277));
INVX1 g139388(.A (n_33271), .Y (n_33275));
INVX1 g139389(.A (n_33270), .Y (n_33276));
OAI21X1 g139390(.A0 (n_35532), .A1 (n_33286), .B0 (n_33287), .Y(n_33288));
NOR2X1 g139395(.A (n_33410), .B (n_33280), .Y (n_33281));
NAND2X1 g139397(.A (n_12835), .B (n_12902), .Y (n_33280));
XOR2X1 g139398(.A (n_17016), .B (n_22365), .Y (n_33286));
NAND2X1 g139399(.A (n_35600), .B (n_13735), .Y (n_33287));
NAND2X1 g139401(.A (n_33293), .B (n_33296), .Y (n_33297));
AOI21X1 g139402(.A0 (n_11732), .A1 (n_32827), .B0 (n_33292), .Y(n_33293));
NOR2X1 g139403(.A (n_33291), .B (n_12800), .Y (n_33292));
NAND2X1 g139404(.A (n_34992), .B (n_33290), .Y (n_33291));
OR2X1 g139405(.A (n_7066), .B (n_7426), .Y (n_33290));
NAND2X1 g139406(.A (n_12800), .B (n_33295), .Y (n_33296));
NOR2X1 g139407(.A (n_7613), .B (n_34992), .Y (n_33295));
INVX1 g139410(.A (n_33299), .Y (n_33300));
NAND3X1 g139411(.A (n_4991), .B (n_33298), .C (n_4759), .Y (n_33299));
AND2X1 g139412(.A (n_5175), .B (n_32106), .Y (n_33298));
NOR2X1 g139413(.A (n_33301), .B (n_33302), .Y (n_33303));
NAND4X1 g139414(.A (n_3514), .B (n_34913), .C (n_4170), .D (n_32517),.Y (n_33301));
NAND2X1 g139415(.A (n_32105), .B (n_4877), .Y (n_33302));
NAND2X1 g139418(.A (n_4087), .B (n_33304), .Y (n_33305));
INVX1 g61(.A (n_1659), .Y (n_33304));
NAND2X2 g139419(.A (n_33314), .B (n_33318), .Y (n_33319));
NAND4X1 g139420(.A (n_33310), .B (n_22880), .C (n_33312), .D(n_33313), .Y (n_33314));
NAND2X1 g139421(.A (n_24289), .B (n_33309), .Y (n_33310));
OR2X1 g139422(.A (n_19898), .B (n_24095), .Y (n_33309));
AOI21X1 g139423(.A0 (n_21289), .A1 (n_19608), .B0 (n_33311), .Y(n_33312));
INVX1 g139424(.A (n_19591), .Y (n_33311));
AOI21X1 g139425(.A0 (n_11559), .A1 (n_17219), .B0 (n_19703), .Y(n_33313));
AOI21X1 g139426(.A0 (n_33315), .A1 (n_22518), .B0 (n_33317), .Y(n_33318));
AND2X1 g139427(.A (n_22880), .B (n_22877), .Y (n_33315));
AOI21X1 g139428(.A0 (n_22956), .A1 (n_17390), .B0 (n_33316), .Y(n_33317));
AND2X1 g139429(.A (n_22293), .B (n_22228), .Y (n_33316));
NAND2X1 g139439(.A (n_33329), .B (P3_d_407), .Y (n_33330));
CLKBUFX1 g139440(.A (n_33405), .Y (n_33329));
NAND2X1 g139441(.A (n_33329), .B (P3_d_406), .Y (n_33331));
NAND2X1 g139442(.A (n_33329), .B (P3_d_398), .Y (n_33332));
NAND2X1 g139443(.A (n_33329), .B (P3_d_384), .Y (n_33333));
NAND3X1 g139444(.A (n_33336), .B (n_33337), .C (n_33338), .Y(n_33339));
OAI21X1 g139445(.A0 (n_34952), .A1 (n_33378), .B0 (n_33335), .Y(n_33336));
NAND2X2 g139447(.A (n_26404), .B (n_26929), .Y (n_33335));
NAND2X1 g139448(.A (n_34753), .B (n_35630), .Y (n_33337));
AOI21X1 g139449(.A0 (n_20195), .A1 (n_10848), .B0 (n_9159), .Y(n_33338));
INVX4 g139450(.A (n_33378), .Y (n_33340));
NAND2X1 g139451(.A (n_33345), .B (n_33348), .Y (n_33349));
NAND3X1 g139452(.A (n_33341), .B (n_8719), .C (n_34700), .Y(n_33345));
NAND2X1 g139453(.A (n_31218), .B (n_31266), .Y (n_33341));
AND2X1 g139457(.A (n_33346), .B (n_33347), .Y (n_33348));
NAND3X1 g139458(.A (n_9252), .B (n_10465), .C (n_34700), .Y(n_33346));
OR2X1 g139459(.A (P2_reg_112), .B (n_6460), .Y (n_33347));
INVX1 g139460(.A (n_34700), .Y (n_33350));
NAND2X1 g139462(.A (n_33351), .B (n_33352), .Y (n_33353));
AND2X1 g139463(.A (n_118), .B (n_167), .Y (n_33351));
AND2X1 g40_dup(.A (n_32476), .B (n_32488), .Y (n_33352));
NAND2X2 g139464(.A (n_33355), .B (n_33357), .Y (n_33358));
INVX2 g139465(.A (n_33354), .Y (n_33355));
NAND2X2 g139466(.A (n_647), .B (n_1464), .Y (n_33354));
INVX1 g139467(.A (n_33356), .Y (n_33357));
NAND2X2 g139468(.A (n_32399), .B (n_203), .Y (n_33356));
INVX1 g139470(.A (n_33361), .Y (n_33362));
AND2X1 g139471(.A (n_32476), .B (n_32488), .Y (n_33361));
INVX1 g139472(.A (n_33363), .Y (n_33364));
INVX1 g139473(.A (n_33356), .Y (n_33363));
OAI21X1 g139474(.A0 (n_33365), .A1 (n_33366), .B0 (n_33367), .Y(n_33368));
MX2X1 g139475(.A (n_17150), .B (n_16411), .S0 (n_16460), .Y(n_33365));
NAND3X1 g139476(.A (n_32210), .B (n_22519), .C (n_32211), .Y(n_33366));
NAND2X1 g139477(.A (n_33365), .B (n_33366), .Y (n_33367));
CLKBUFX1 g2(.A (n_33375), .Y (n_33376));
NOR2X1 g26(.A (n_33374), .B (n_33373), .Y (n_33375));
NAND4X1 g27(.A (n_33369), .B (n_33371), .C (n_32929), .D (n_33561),.Y (n_33373));
AND2X1 g139478(.A (n_33257), .B (n_33918), .Y (n_33369));
CLKBUFX3 g139479(.A (n_33370), .Y (n_33371));
INVX1 g139480(.A (P2_IR[0] ), .Y (n_33370));
NAND3X1 g139482(.A (n_1720), .B (n_1015), .C (n_35447), .Y (n_33374));
NAND4X1 g139483(.A (n_33380), .B (n_33381), .C (n_20151), .D(n_9017), .Y (n_33382));
NAND2X1 g139484(.A (n_33377), .B (n_33379), .Y (n_33380));
NAND2X1 g139485(.A (n_27471), .B (n_28572), .Y (n_33377));
OR2X1 g139486(.A (n_33378), .B (n_34952), .Y (n_33379));
NOR2X1 g139487(.A (n_7774), .B (n_7777), .Y (n_33378));
NAND2X1 g139488(.A (n_29378), .B (n_34753), .Y (n_33381));
INVX1 g139505(.A (n_34405), .Y (n_33401));
NAND3X1 g139506(.A (n_33402), .B (n_33403), .C (n_33409), .Y(n_33410));
NOR2X1 g139507(.A (n_11929), .B (n_11931), .Y (n_33402));
INVX1 g139508(.A (n_11930), .Y (n_33403));
NOR2X1 g139509(.A (n_33408), .B (n_11691), .Y (n_33409));
NAND2X1 g139510(.A (n_33406), .B (n_33407), .Y (n_33408));
AOI22X1 g139511(.A0 (P3_d_384), .A1 (n_33405), .B0 (n_33405), .B1(P3_d_407), .Y (n_33406));
CLKBUFX3 g139512(.A (n_33404), .Y (n_33405));
NAND3X1 g139513(.A (n_32481), .B (n_7749), .C (n_7719), .Y (n_33404));
OAI21X1 g139514(.A0 (P3_d_406), .A1 (P3_d_398), .B0 (n_33405), .Y(n_33407));
INVX2 g139515(.A (n_33411), .Y (n_33412));
NAND3X1 g139516(.A (n_32481), .B (n_7749), .C (n_7719), .Y (n_33411));
NAND2X1 g139521(.A (n_33415), .B (n_20153), .Y (n_33416));
NAND2X1 g139522(.A (n_29925), .B (n_35058), .Y (n_33415));
NAND2X1 g139526(.A (n_34770), .B (n_35058), .Y (n_33419));
INVX1 g139527(.A (n_18931), .Y (n_33420));
NOR2X1 g139530(.A (n_33426), .B (n_33430), .Y (n_33431));
NAND2X1 g139531(.A (n_33923), .B (n_33369), .Y (n_33426));
NAND2X1 g139532(.A (n_35225), .B (n_33429), .Y (n_33430));
NOR2X1 g25(.A (n_35712), .B (n_33427), .Y (n_33429));
NAND2X2 g139533(.A (n_35868), .B (n_200), .Y (n_33427));
INVX1 g24(.A (n_33429), .Y (n_33432));
NAND2X1 g139535(.A (n_33433), .B (n_35225), .Y (n_33434));
INVX1 g139536(.A (n_33426), .Y (n_33433));
INVX1 g139537(.A (n_35711), .Y (n_35447));
INVX1 g139538(.A (n_33427), .Y (n_33436));
NAND3X1 g139545(.A (n_33445), .B (n_33446), .C (n_33447), .Y(n_33448));
OAI21X1 g139546(.A0 (n_29199), .A1 (n_34770), .B0 (n_33444), .Y(n_33445));
NAND2X1 g139547(.A (n_27481), .B (n_28555), .Y (n_33444));
NAND2X1 g139548(.A (n_24786), .B (n_29357), .Y (n_33446));
AOI22X1 g139549(.A0 (n_10889), .A1 (n_8946), .B0 (n_20218), .B1(n_10890), .Y (n_33447));
NAND2X1 g139551(.A (n_33454), .B (n_33457), .Y (n_33458));
NAND3X1 g139552(.A (n_33450), .B (n_31573), .C (n_35024), .Y(n_33454));
NAND2X1 g139553(.A (n_30986), .B (n_30391), .Y (n_33450));
AND2X1 g139557(.A (n_33455), .B (n_33456), .Y (n_33457));
NAND3X1 g139558(.A (n_8235), .B (n_30881), .C (n_35024), .Y(n_33455));
AOI22X1 g139559(.A0 (P1_reg3[26] ), .A1 (n_2091), .B0 (n_6769), .B1(n_4124), .Y (n_33456));
NAND4X1 g139571(.A (n_33473), .B (n_33478), .C (n_33479), .D(n_33592), .Y (n_33480));
NOR2X1 g139572(.A (n_34073), .B (n_35259), .Y (n_33473));
INVX1 g139576(.A (n_33477), .Y (n_33478));
NAND2X1 g139577(.A (n_32579), .B (n_33476), .Y (n_33477));
NOR2X1 g139578(.A (n_33474), .B (n_33475), .Y (n_33476));
INVX1 g139579(.A (n_32580), .Y (n_33474));
INVX1 g139580(.A (n_1662), .Y (n_33475));
INVX1 g139581(.A (n_4141), .Y (n_33479));
NOR2X1 g139582(.A (n_33481), .B (n_33477), .Y (n_35090));
INVX1 g139583(.A (n_33592), .Y (n_33481));
NAND2X1 g139584(.A (n_34016), .B (n_34009), .Y (n_35251));
NAND2X1 g139586(.A (n_33592), .B (n_1662), .Y (n_33485));
NAND2X1 g139593(.A (n_33496), .B (n_33500), .Y (n_33501));
OAI21X1 g139594(.A0 (n_33492), .A1 (n_33494), .B0 (n_33495), .Y(n_33496));
OR2X1 g139595(.A (n_30557), .B (n_30180), .Y (n_33492));
INVX1 g139596(.A (n_33505), .Y (n_33494));
NAND2X1 g139598(.A (n_29075), .B (n_28324), .Y (n_33495));
AOI21X1 g139599(.A0 (n_21246), .A1 (n_22123), .B0 (n_33499), .Y(n_33500));
AND2X1 g139600(.A (n_34708), .B (n_33498), .Y (n_33499));
NAND2X1 g139602(.A (n_27767), .B (n_28324), .Y (n_33498));
NAND2X1 g139604(.A (n_33507), .B (n_33511), .Y (n_33512));
NAND2X1 g139605(.A (n_33503), .B (n_33506), .Y (n_33507));
NAND2X1 g139606(.A (n_29085), .B (n_28327), .Y (n_33503));
NAND2X1 g139607(.A (n_33504), .B (n_33505), .Y (n_33506));
NOR2X1 g139608(.A (n_30557), .B (n_30180), .Y (n_33504));
NAND3X1 g139609(.A (n_7987), .B (n_30897), .C (n_6441), .Y (n_33505));
AOI21X1 g139610(.A0 (n_21255), .A1 (n_21694), .B0 (n_33510), .Y(n_33511));
AND2X1 g139611(.A (n_34708), .B (n_33509), .Y (n_33510));
NAND2X1 g139613(.A (n_27804), .B (n_28327), .Y (n_33509));
INVX1 g139614(.A (n_33505), .Y (n_33513));
INVX1 g139637(.A (n_853), .Y (n_33535));
NOR2X1 g139638(.A (n_34093), .B (n_2982), .Y (n_33536));
INVX1 g139639(.A (n_34011), .Y (n_4432));
INVX1 g139640(.A (n_34009), .Y (n_33540));
NAND3X1 g139641(.A (n_33542), .B (n_33545), .C (n_33547), .Y(n_33548));
AOI21X1 g139642(.A0 (n_30180), .A1 (n_33541), .B0 (n_27517), .Y(n_33542));
NAND2X1 g139643(.A (n_29079), .B (n_21262), .Y (n_33541));
NOR2X1 g139644(.A (n_29105), .B (n_33544), .Y (n_33545));
OAI21X1 g139645(.A0 (n_29093), .A1 (n_27696), .B0 (n_33543), .Y(n_33544));
NAND2X1 g139646(.A (n_21263), .B (n_21694), .Y (n_33543));
NAND2X1 g139647(.A (n_33546), .B (n_33541), .Y (n_33547));
NAND2X2 g139648(.A (n_8718), .B (n_33505), .Y (n_33546));
MX2X1 g139649(.A (n_33551), .B (n_33550), .S0 (n_33554), .Y(n_33555));
INVX1 g139651(.A (n_33551), .Y (n_33550));
NAND2X2 g139652(.A (n_15946), .B (n_16148), .Y (n_33551));
NAND3X1 g139653(.A (n_33552), .B (n_33553), .C (n_21311), .Y(n_33554));
AND2X1 g139654(.A (n_17125), .B (n_21385), .Y (n_33552));
NOR2X1 g139655(.A (n_20545), .B (n_21161), .Y (n_33553));
INVX1 g139656(.A (n_33551), .Y (n_33556));
NAND2X1 g139657(.A (n_21311), .B (n_33552), .Y (n_33557));
INVX1 g139658(.A (n_33553), .Y (n_33558));
NAND4X1 g139659(.A (n_33559), .B (n_33560), .C (n_33561), .D(n_33562), .Y (n_33563));
INVX2 g139660(.A (P2_IR[7] ), .Y (n_33559));
INVX2 g139661(.A (P2_IR[6] ), .Y (n_33560));
INVX2 g139662(.A (P2_IR[4] ), .Y (n_33561));
INVX2 g139663(.A (P2_IR[5] ), .Y (n_33562));
NAND3X1 g139664(.A (n_33570), .B (n_33571), .C (n_33572), .Y(n_33573));
NAND3X1 g139665(.A (n_2869), .B (n_33567), .C (P3_IR[13] ), .Y(n_33570));
NAND2X1 g139667(.A (n_34853), .B (n_33141), .Y (n_33564));
INVX4 g139668(.A (n_33566), .Y (n_33567));
INVX4 g139669(.A (P3_IR[31] ), .Y (n_33566));
INVX1 g139671(.A (P3_IR[13] ), .Y (n_33568));
NAND3X1 g139672(.A (n_33564), .B (n_33567), .C (n_33568), .Y(n_33571));
OR2X1 g139673(.A (n_33568), .B (n_33567), .Y (n_33572));
NAND3X1 g139674(.A (n_33577), .B (n_33578), .C (n_33581), .Y(n_33582));
NOR2X1 g139675(.A (n_33576), .B (n_35116), .Y (n_33577));
NAND4X1 g139676(.A (n_32642), .B (n_2028), .C (n_33574), .D(n_33371), .Y (n_35116));
OR2X1 g139677(.A (n_366), .B (n_3719), .Y (n_33574));
NOR2X1 g139678(.A (n_2415), .B (n_4189), .Y (n_33576));
AND2X1 g139679(.A (n_4357), .B (n_4169), .Y (n_33578));
OR2X1 g139680(.A (n_33579), .B (n_33580), .Y (n_33581));
INVX1 g139681(.A (P2_IR[31] ), .Y (n_33579));
MX2X1 g139682(.A (n_366), .B (P2_IR[28] ), .S0 (n_3443), .Y(n_33580));
AND2X1 g139683(.A (n_33581), .B (n_33574), .Y (n_33583));
NAND2X1 g139684(.A (n_4169), .B (n_32642), .Y (n_33584));
NOR2X1 g139685(.A (n_33585), .B (n_33576), .Y (n_33586));
INVX1 g139686(.A (n_2028), .Y (n_33585));
INVX1 g139687(.A (P2_IR[31] ), .Y (n_33587));
NAND2X2 g13(.A (n_33590), .B (n_34946), .Y (n_33592));
NAND2X1 g14(.A (n_33588), .B (n_33589), .Y (n_33590));
NAND2X1 g16(.A (n_2998), .B (n_1661), .Y (n_33588));
NAND2X1 g15(.A (n_452), .B (n_3029), .Y (n_33589));
NAND3X1 g139704(.A (n_33608), .B (n_33612), .C (n_33614), .Y(n_33615));
NAND2X1 g139705(.A (n_21755), .B (n_22626), .Y (n_33608));
NAND2X1 g139706(.A (n_33609), .B (n_33611), .Y (n_33612));
NOR2X1 g139707(.A (n_21762), .B (n_21754), .Y (n_33609));
CLKBUFX1 g139708(.A (n_33610), .Y (n_33611));
NAND2X1 g139709(.A (n_20025), .B (n_20026), .Y (n_33610));
AOI21X1 g139710(.A0 (n_22552), .A1 (n_22352), .B0 (n_33613), .Y(n_33614));
NAND2X1 g139711(.A (n_20356), .B (n_32589), .Y (n_33613));
NAND2X2 g139712(.A (n_33623), .B (n_33625), .Y (n_33626));
NAND2X2 g139713(.A (n_33620), .B (n_33622), .Y (n_33623));
NAND2X2 g139714(.A (n_33616), .B (n_33619), .Y (n_33620));
NAND3X1 g139715(.A (n_23925), .B (n_20418), .C (n_20998), .Y(n_33616));
AOI21X1 g139716(.A0 (n_20414), .A1 (n_20825), .B0 (n_33618), .Y(n_33619));
NAND3X1 g139717(.A (n_20999), .B (n_18666), .C (n_33617), .Y(n_33618));
INVX1 g139718(.A (n_17248), .Y (n_33617));
CLKBUFX1 g139719(.A (n_33621), .Y (n_33622));
NAND2X1 g139720(.A (n_16770), .B (n_16769), .Y (n_33621));
NAND3X1 g139721(.A (n_33624), .B (n_33619), .C (n_33616), .Y(n_33625));
INVX1 g139722(.A (n_33622), .Y (n_33624));
NAND4X1 g139723(.A (n_33631), .B (n_33634), .C (n_33635), .D(n_33636), .Y (n_33637));
AOI21X1 g139724(.A0 (n_33627), .A1 (n_33629), .B0 (n_33630), .Y(n_33631));
NAND2X1 g139725(.A (n_14005), .B (n_14437), .Y (n_33627));
INVX1 g139726(.A (n_33713), .Y (n_33629));
NAND2X1 g139728(.A (n_27914), .B (n_27915), .Y (n_33630));
NOR2X1 g139729(.A (n_33633), .B (n_29003), .Y (n_33634));
NAND2X1 g139730(.A (n_27913), .B (n_33632), .Y (n_33633));
NAND2X1 g139731(.A (n_17139), .B (n_7988), .Y (n_33632));
AOI21X1 g139732(.A0 (n_8954), .A1 (n_28020), .B0 (n_20161), .Y(n_33635));
AOI22X1 g139733(.A0 (n_27522), .A1 (n_27261), .B0 (n_11138), .B1(n_3887), .Y (n_33636));
NAND2X2 g139734(.A (n_33641), .B (n_33643), .Y (n_33644));
NAND2X1 g139735(.A (n_33638), .B (n_33640), .Y (n_33641));
NAND2X1 g139737(.A (n_16445), .B (n_17222), .Y (n_33638));
NAND3X1 g139738(.A (n_32096), .B (n_23310), .C (n_32097), .Y(n_33640));
NAND4X1 g139739(.A (n_32096), .B (n_23310), .C (n_32097), .D(n_33642), .Y (n_33643));
INVX1 g139740(.A (n_33638), .Y (n_33642));
OAI21X1 g139741(.A0 (n_33645), .A1 (n_33646), .B0 (n_33647), .Y(n_33648));
NAND3X1 g139742(.A (n_32575), .B (n_32576), .C (n_23141), .Y(n_33645));
NAND2X1 g139743(.A (n_19331), .B (n_18069), .Y (n_33646));
NAND2X1 g139744(.A (n_33646), .B (n_33645), .Y (n_33647));
NAND3X1 g139745(.A (n_33649), .B (n_33651), .C (n_33654), .Y(n_33655));
OR2X1 g139746(.A (n_10779), .B (n_29012), .Y (n_33649));
AOI21X1 g139747(.A0 (n_29878), .A1 (n_33650), .B0 (n_15016), .Y(n_33651));
OR2X1 g139748(.A (n_35044), .B (n_30399), .Y (n_33650));
AOI21X1 g139749(.A0 (n_29615), .A1 (n_30438), .B0 (n_33653), .Y(n_33654));
INVX1 g139750(.A (n_33652), .Y (n_33653));
AOI22X1 g139751(.A0 (n_25942), .A1 (n_24904), .B0 (n_14550), .B1(n_10215), .Y (n_33652));
NAND2X1 g139752(.A (n_33658), .B (n_33662), .Y (n_33663));
AOI21X1 g139753(.A0 (n_28696), .A1 (n_33656), .B0 (n_33657), .Y(n_33658));
OR2X1 g139754(.A (n_33991), .B (n_29155), .Y (n_33656));
AND2X1 g139755(.A (n_28874), .B (n_28052), .Y (n_33657));
NAND2X1 g139756(.A (n_33659), .B (n_33661), .Y (n_33662));
NAND2X1 g139757(.A (n_14442), .B (n_14936), .Y (n_33659));
INVX1 g139758(.A (n_33713), .Y (n_33661));
NAND4X1 g139760(.A (n_35331), .B (n_35332), .C (n_33670), .D(n_29566), .Y (n_33671));
INVX1 g139761(.A (n_33666), .Y (n_35332));
NAND2X1 g139762(.A (n_33664), .B (n_33665), .Y (n_33666));
NAND2X1 g139763(.A (n_29955), .B (n_29565), .Y (n_33664));
NAND2X1 g139764(.A (n_29405), .B (n_29565), .Y (n_33665));
AND2X1 g139765(.A (n_33668), .B (n_21701), .Y (n_35331));
AOI21X1 g139766(.A0 (n_14810), .A1 (n_13695), .B0 (n_29169), .Y(n_33668));
NAND2X1 g139767(.A (n_14611), .B (n_15147), .Y (n_33670));
NAND4X1 g139768(.A (n_33675), .B (n_33679), .C (n_33680), .D(n_1556), .Y (n_33681));
INVX1 g139769(.A (n_33674), .Y (n_33675));
NAND2X1 g139770(.A (n_33673), .B (n_33672), .Y (n_33674));
NOR2X1 g139771(.A (n_1970), .B (n_2723), .Y (n_33672));
NOR2X1 g139772(.A (n_1098), .B (n_1099), .Y (n_33673));
INVX1 g139773(.A (n_33678), .Y (n_33679));
NAND2X1 g139774(.A (n_33677), .B (n_1043), .Y (n_33678));
INVX1 g139775(.A (n_33676), .Y (n_33677));
NAND3X1 g139776(.A (n_739), .B (n_1289), .C (n_1401), .Y (n_33676));
NOR2X1 g139777(.A (n_1096), .B (n_1097), .Y (n_33680));
NAND3X1 g139798(.A (n_33706), .B (n_33708), .C (n_33709), .Y(n_33710));
NAND4X1 g139799(.A (n_34281), .B (n_21008), .C (n_19437), .D(n_33705), .Y (n_33706));
NAND2X1 g139801(.A (n_20988), .B (n_21007), .Y (n_33703));
NOR2X1 g139802(.A (n_16697), .B (n_17612), .Y (n_33705));
INVX1 g139803(.A (n_33707), .Y (n_33708));
OAI21X1 g45_dup(.A0 (n_21944), .A1 (n_20394), .B0 (n_21860), .Y(n_33707));
NAND2X1 g139804(.A (n_34281), .B (n_21612), .Y (n_33709));
OAI21X1 g139805(.A0 (n_21944), .A1 (n_20394), .B0 (n_21860), .Y(n_33711));
NAND2X1 g139806(.A (n_33716), .B (n_33720), .Y (n_33721));
NAND2X1 g139807(.A (n_33712), .B (n_33722), .Y (n_33716));
NAND2X1 g139808(.A (n_14230), .B (n_14670), .Y (n_33712));
NAND2X2 g139811(.A (n_7771), .B (n_7773), .Y (n_33713));
AND2X1 g139812(.A (n_33718), .B (n_33719), .Y (n_33720));
NAND2X1 g139813(.A (n_29401), .B (n_33717), .Y (n_33718));
OR2X1 g139814(.A (n_33991), .B (n_28158), .Y (n_33717));
NAND2X1 g139815(.A (n_28840), .B (n_30454), .Y (n_33719));
INVX1 g139816(.A (n_33713), .Y (n_33722));
OR2X1 g139817(.A (n_33725), .B (n_33727), .Y (n_33728));
OAI21X1 g139818(.A0 (n_8250), .A1 (n_33723), .B0 (n_33724), .Y(n_33725));
OR2X1 g139819(.A (P1_n_449), .B (n_9382), .Y (n_33723));
NAND2X1 g139820(.A (n_6986), .B (n_10890), .Y (n_33724));
AOI21X1 g139821(.A0 (n_31319), .A1 (n_31138), .B0 (n_33726), .Y(n_33727));
OR2X1 g139822(.A (P1_n_449), .B (n_8070), .Y (n_33726));
INVX1 g139823(.A (P1_n_449), .Y (n_15723));
OAI21X1 g139824(.A0 (n_33733), .A1 (n_33734), .B0 (n_33736), .Y(n_33737));
INVX1 g139825(.A (n_33732), .Y (n_33733));
NAND2X1 g139826(.A (n_33730), .B (n_33731), .Y (n_33732));
NAND2X2 g139827(.A (n_35736), .B (n_26236), .Y (n_33730));
NAND2X1 g139828(.A (n_35829), .B (n_13352), .Y (n_33731));
OR2X1 g139830(.A (n_7387), .B (n_7342), .Y (n_33734));
NAND2X1 g139831(.A (n_19555), .B (n_21328), .Y (n_33736));
INVX8 g139832(.A (n_33734), .Y (n_33738));
NAND2X2 g139833(.A (n_35333), .B (n_35334), .Y (n_33748));
OAI21X1 g139834(.A0 (n_33739), .A1 (n_33741), .B0 (n_17133), .Y(n_35334));
INVX1 g139835(.A (n_12979), .Y (n_33739));
NAND2X1 g139836(.A (n_12906), .B (n_17178), .Y (n_33741));
OAI21X1 g139838(.A0 (n_33739), .A1 (n_33744), .B0 (n_33746), .Y(n_35333));
NAND2X1 g139839(.A (n_12906), .B (n_17178), .Y (n_33744));
AOI21X1 g139841(.A0 (n_13219), .A1 (n_12798), .B0 (n_33745), .Y(n_33746));
AND2X1 g139842(.A (n_8737), .B (n_12905), .Y (n_33745));
NAND2X1 g139843(.A (n_17133), .B (n_15962), .Y (n_33749));
NAND2X1 g139844(.A (n_12979), .B (n_12906), .Y (n_33750));
CLKBUFX1 g139845(.A (n_33754), .Y (n_33755));
OAI21X1 g139846(.A0 (n_33751), .A1 (n_33752), .B0 (n_33753), .Y(n_33754));
NAND3X1 g139847(.A (n_32173), .B (n_23409), .C (n_32174), .Y(n_33751));
NAND2X1 g139848(.A (n_17931), .B (n_18691), .Y (n_33752));
NAND2X1 g139849(.A (n_33751), .B (n_33752), .Y (n_33753));
AOI21X1 g139859(.A0 (n_34841), .A1 (n_33767), .B0 (n_33771), .Y(n_33772));
OAI21X1 g139862(.A0 (n_32537), .A1 (n_34548), .B0 (n_16878), .Y(n_33767));
NAND2X2 g139863(.A (n_33768), .B (n_33770), .Y (n_33771));
NAND2X2 g139864(.A (n_16562), .B (n_35849), .Y (n_33768));
INVX1 g139865(.A (n_33769), .Y (n_33770));
AND2X1 g139866(.A (n_15821), .B (n_9257), .Y (n_33769));
OAI21X1 g139867(.A0 (n_33775), .A1 (n_33776), .B0 (n_33780), .Y(n_33781));
NAND3X1 g139868(.A (n_35671), .B (n_35666), .C (n_33774), .Y(n_33775));
INVX2 g139870(.A (n_18843), .Y (n_33774));
AOI21X1 g139871(.A0 (n_20044), .A1 (n_17089), .B0 (n_21110), .Y(n_33776));
AOI21X1 g139872(.A0 (n_33777), .A1 (n_33778), .B0 (n_35938), .Y(n_33780));
NAND2X2 g139873(.A (n_18876), .B (n_19311), .Y (n_33777));
NOR2X1 g139874(.A (n_18843), .B (n_35670), .Y (n_33778));
CLKBUFX1 g139876(.A (n_33776), .Y (n_33782));
NAND3X1 g139877(.A (n_33786), .B (n_33788), .C (n_33789), .Y(n_33790));
NAND2X1 g139878(.A (n_33783), .B (n_33785), .Y (n_33786));
NAND2X1 g139879(.A (n_27465), .B (n_28548), .Y (n_33783));
BUFX3 g139880(.A (n_33784), .Y (n_33785));
NOR2X1 g139881(.A (n_8304), .B (n_8948), .Y (n_33784));
AOI21X1 g139882(.A0 (n_24903), .A1 (n_25942), .B0 (n_33787), .Y(n_33788));
AND2X1 g139883(.A (n_14550), .B (n_10225), .Y (n_33787));
NAND2X1 g139884(.A (n_29191), .B (n_29889), .Y (n_33789));
AOI21X1 g139886(.A0 (n_33801), .A1 (n_33802), .B0 (n_33805), .Y(n_33806));
INVX1 g139887(.A (n_33800), .Y (n_33801));
NOR2X1 g139888(.A (n_33793), .B (n_33799), .Y (n_33800));
INVX1 g139889(.A (n_33792), .Y (n_33793));
NAND2X1 g139890(.A (n_13185), .B (n_10245), .Y (n_33792));
AOI21X1 g139891(.A0 (n_33277), .A1 (n_33274), .B0 (n_13318), .Y(n_33799));
AND2X1 g139897(.A (n_7400), .B (n_29944), .Y (n_33802));
AOI21X1 g139898(.A0 (n_18281), .A1 (n_33792), .B0 (n_21365), .Y(n_33805));
NAND2X2 g139900(.A (n_8036), .B (n_8679), .Y (n_33803));
INVX4 g139901(.A (n_33802), .Y (n_33807));
NAND2X2 g139902(.A (n_33274), .B (n_33277), .Y (n_33808));
MX2X1 g139903(.A (n_33810), .B (n_33809), .S0 (n_33811), .Y(n_33812));
INVX1 g139904(.A (n_33809), .Y (n_33810));
NAND2X1 g139905(.A (n_33051), .B (n_16180), .Y (n_33809));
NAND2X1 g139906(.A (n_22669), .B (n_23522), .Y (n_33811));
MX2X1 g139909(.A (P2_IR[14] ), .B (n_682), .S0 (n_2980), .Y(n_33813));
INVX1 g139910(.A (n_33814), .Y (n_33815));
INVX1 g139911(.A (P2_IR[31] ), .Y (n_33814));
AND2X1 g139912(.A (n_34093), .B (P2_IR[14] ), .Y (n_33816));
AOI21X1 g139934(.A0 (n_33852), .A1 (n_33857), .B0 (n_33858), .Y(n_33859));
INVX1 g139935(.A (n_33851), .Y (n_33852));
AOI21X1 g139936(.A0 (n_18185), .A1 (n_18775), .B0 (n_21059), .Y(n_33851));
INVX1 g139937(.A (n_35396), .Y (n_33857));
AND2X1 g139939(.A (n_19235), .B (n_18062), .Y (n_33853));
NAND2X1 g139941(.A (n_19304), .B (n_34107), .Y (n_33854));
NAND2X1 g139942(.A (n_20535), .B (n_20424), .Y (n_33858));
INVX1 g139943(.A (n_33853), .Y (n_33860));
INVX1 g139968(.A (n_33904), .Y (n_33905));
AOI21X1 g139969(.A0 (n_15619), .A1 (n_15542), .B0 (n_33903), .Y(n_33904));
OAI21X1 g139970(.A0 (n_7403), .A1 (n_15430), .B0 (n_33902), .Y(n_33903));
NAND2X1 g139971(.A (n_33897), .B (n_33901), .Y (n_33902));
INVX2 g139972(.A (n_33896), .Y (n_33897));
INVX1 g139973(.A (n_33895), .Y (n_33896));
INVX2 g139974(.A (n_33894), .Y (n_33895));
NAND2X1 g139975(.A (n_6357), .B (n_6439), .Y (n_33894));
INVX1 g139976(.A (n_33899), .Y (n_33901));
AOI21X1 g139978(.A0 (n_3042), .A1 (n_33567), .B0 (n_33898), .Y(n_33899));
AND2X1 g139979(.A (n_33566), .B (P3_IR[18] ), .Y (n_33898));
INVX2 g139980(.A (n_33897), .Y (n_33906));
NAND2X2 g139981(.A (n_33910), .B (n_33916), .Y (n_33917));
AOI21X1 g139982(.A0 (n_20402), .A1 (n_34491), .B0 (n_33909), .Y(n_33910));
NAND2X1 g139983(.A (n_20992), .B (n_33908), .Y (n_33909));
NOR2X1 g139984(.A (n_17745), .B (n_33907), .Y (n_33908));
INVX1 g139985(.A (n_18738), .Y (n_33907));
NAND3X1 g139986(.A (n_33911), .B (n_34487), .C (n_33915), .Y(n_33916));
NAND2X2 g139987(.A (n_23612), .B (n_22628), .Y (n_33911));
INVX1 g139988(.A (n_33914), .Y (n_33915));
NAND2X1 g139989(.A (n_20401), .B (n_33912), .Y (n_33914));
AND2X1 g139991(.A (n_32381), .B (n_19255), .Y (n_33912));
NAND3X1 g139992(.A (n_33921), .B (n_33922), .C (n_33923), .Y(n_33924));
NOR2X1 g139993(.A (n_33261), .B (n_33920), .Y (n_33921));
INVX1 g139995(.A (P2_IR[2] ), .Y (n_33918));
NAND2X2 g139996(.A (n_32929), .B (n_33370), .Y (n_33920));
NOR2X1 g139997(.A (n_265), .B (n_396), .Y (n_33922));
AND2X1 g139998(.A (n_33562), .B (n_33561), .Y (n_33923));
NAND2X2 g140025(.A (n_33961), .B (n_33962), .Y (n_33963));
AOI21X1 g140026(.A0 (n_7503), .A1 (n_13697), .B0 (n_7750), .Y(n_33961));
AOI21X1 g140027(.A0 (n_3887), .A1 (n_8197), .B0 (n_7406), .Y(n_33962));
NAND2X2 g140028(.A (n_15841), .B (n_15842), .Y (n_33964));
NAND2X1 g140030(.A (n_33973), .B (n_33968), .Y (n_33976));
INVX1 g140031(.A (n_33967), .Y (n_33968));
NAND3X1 g140032(.A (n_15693), .B (n_15691), .C (n_6825), .Y(n_33967));
INVX2 g140035(.A (n_33972), .Y (n_33973));
NAND3X1 g140036(.A (n_33969), .B (n_33970), .C (n_33971), .Y(n_33972));
NAND2X1 g140037(.A (n_34355), .B (n_15696), .Y (n_33969));
NAND2X1 g140038(.A (n_15685), .B (n_15696), .Y (n_33970));
OR2X1 g140039(.A (n_4507), .B (n_6823), .Y (n_33971));
NAND2X1 g140040(.A (n_16611), .B (n_33982), .Y (n_33983));
NOR2X1 g140042(.A (n_16096), .B (n_15881), .Y (n_33977));
NAND2X1 g140043(.A (n_33980), .B (n_33981), .Y (n_33982));
INVX1 g140044(.A (n_33979), .Y (n_33980));
NAND2X1 g36_dup(.A (n_7733), .B (n_7804), .Y (n_33979));
NAND3X1 g140045(.A (n_15577), .B (n_6720), .C (n_15575), .Y(n_33981));
NAND2X1 g140046(.A (n_7804), .B (n_7733), .Y (n_16331));
INVX1 g140047(.A (n_33981), .Y (n_33985));
NAND4X1 g140048(.A (n_33986), .B (n_33989), .C (n_33996), .D(n_33997), .Y (n_33998));
NAND2X1 g140049(.A (n_15298), .B (n_33629), .Y (n_33986));
NAND2X1 g140050(.A (n_29125), .B (n_28347), .Y (n_33989));
INVX1 g140053(.A (n_33995), .Y (n_33996));
AOI21X1 g140054(.A0 (n_28528), .A1 (n_7997), .B0 (n_33994), .Y(n_33995));
AND2X1 g140057(.A (n_7773), .B (n_7396), .Y (n_33991));
INVX2 g140058(.A (n_33993), .Y (n_33994));
NAND2X2 g140059(.A (n_28154), .B (n_28153), .Y (n_33993));
AOI21X1 g140060(.A0 (n_30109), .A1 (n_33993), .B0 (n_22108), .Y(n_33997));
NOR2X1 g140061(.A (n_33999), .B (n_34003), .Y (n_34004));
NAND2X2 g140062(.A (n_7565), .B (n_7510), .Y (n_33999));
INVX1 g140063(.A (n_34002), .Y (n_34003));
NAND2X1 g140064(.A (n_34000), .B (n_34001), .Y (n_34002));
AOI21X1 g140065(.A0 (n_34469), .A1 (n_15464), .B0 (n_7358), .Y(n_34000));
NAND2X1 g140066(.A (n_7291), .B (n_15464), .Y (n_34001));
NAND4X1 g140067(.A (n_34008), .B (n_34009), .C (n_34011), .D(n_34012), .Y (n_35259));
NOR2X1 g140068(.A (n_34005), .B (n_34007), .Y (n_34008));
NOR2X1 g140069(.A (n_377), .B (n_2819), .Y (n_34005));
NAND2X1 g140070(.A (n_888), .B (n_34006), .Y (n_34007));
NAND2X1 g140071(.A (n_33814), .B (n_1175), .Y (n_34006));
NOR2X1 g140072(.A (n_33535), .B (n_33536), .Y (n_34009));
INVX2 g140073(.A (n_34010), .Y (n_34011));
OAI21X1 g140074(.A0 (n_3021), .A1 (n_3279), .B0 (n_765), .Y(n_34010));
NAND2X1 g140075(.A (n_3150), .B (n_852), .Y (n_34012));
NAND2X1 g140076(.A (n_34012), .B (n_34006), .Y (n_34014));
NOR2X1 g140077(.A (n_34015), .B (n_34005), .Y (n_34016));
INVX1 g140078(.A (n_888), .Y (n_34015));
INVX1 g140113(.A (n_34067), .Y (n_34068));
NAND2X1 g140114(.A (n_34063), .B (n_34066), .Y (n_34067));
INVX1 g140115(.A (n_34062), .Y (n_34063));
NAND2X2 g140116(.A (n_17045), .B (n_17051), .Y (n_34062));
AND2X1 g140117(.A (n_34064), .B (n_34065), .Y (n_34066));
NAND2X2 g140118(.A (n_16026), .B (n_16102), .Y (n_34064));
NAND2X1 g140119(.A (n_16317), .B (n_16112), .Y (n_34065));
NAND4X1 g140120(.A (n_34076), .B (n_34077), .C (n_34078), .D(n_34079), .Y (n_34080));
NOR2X1 g140121(.A (n_4274), .B (n_34075), .Y (n_34076));
NAND2X1 g140122(.A (n_34070), .B (n_4051), .Y (n_34075));
INVX1 g140123(.A (n_34069), .Y (n_34070));
NAND2X1 g64_dup(.A (n_34011), .B (n_3914), .Y (n_34069));
NAND2X2 g140125(.A (n_34071), .B (n_34072), .Y (n_34073));
NAND2X1 g140126(.A (n_33813), .B (n_33815), .Y (n_34071));
INVX1 g140127(.A (n_33816), .Y (n_34072));
INVX1 g140128(.A (n_3933), .Y (n_34077));
AND2X1 g140129(.A (n_32579), .B (n_32580), .Y (n_34078));
XOR2X1 g140130(.A (n_265), .B (n_2453), .Y (n_34079));
NAND2X1 g140131(.A (n_3914), .B (n_34011), .Y (n_34081));
INVX1 g140132(.A (n_34079), .Y (n_34082));
NAND2X2 g140133(.A (n_34088), .B (n_34091), .Y (n_34092));
AOI21X1 g140134(.A0 (n_377), .A1 (P2_IR[22] ), .B0 (n_34087), .Y(n_34088));
NOR2X1 g140136(.A (n_2980), .B (n_34086), .Y (n_34087));
NAND3X1 g140137(.A (n_2321), .B (n_34946), .C (P2_IR[22] ), .Y(n_34086));
NAND3X1 g140140(.A (n_34089), .B (n_34946), .C (n_34090), .Y(n_34091));
OR2X1 g140141(.A (n_2980), .B (n_2370), .Y (n_34089));
INVX1 g140142(.A (P2_IR[22] ), .Y (n_34090));
INVX1 g140143(.A (n_34946), .Y (n_34093));
INVX1 g140145(.A (n_34094), .Y (n_34095));
OAI22X1 g140146(.A0 (n_20744), .A1 (n_10320), .B0 (n_18371), .B1(n_17909), .Y (n_34094));
NAND3X1 g140147(.A (n_34096), .B (n_34099), .C (n_34100), .Y(n_34101));
NAND3X1 g140148(.A (n_23729), .B (n_22889), .C (n_23521), .Y(n_34096));
NOR2X1 g140149(.A (n_34098), .B (n_20898), .Y (n_34099));
INVX1 g140150(.A (n_34097), .Y (n_34098));
AOI21X1 g140151(.A0 (n_18626), .A1 (n_32967), .B0 (n_17887), .Y(n_34097));
NAND2X1 g140152(.A (n_22668), .B (n_22889), .Y (n_34100));
NAND2X1 g140153(.A (n_34108), .B (n_34110), .Y (n_34111));
NAND2X1 g140154(.A (n_35936), .B (n_34107), .Y (n_34108));
NAND2X2 g140156(.A (n_35864), .B (n_34106), .Y (n_34107));
NAND2X2 g140158(.A (n_8056), .B (n_7568), .Y (n_34104));
NAND2X1 g140159(.A (n_15621), .B (n_15726), .Y (n_34106));
INVX1 g140160(.A (n_34109), .Y (n_34110));
NOR2X1 g140161(.A (n_34106), .B (n_35864), .Y (n_34109));
INVX2 g140162(.A (n_35937), .Y (n_34112));
NAND2X2 g140163(.A (n_15621), .B (n_15726), .Y (n_18532));
NAND4X1 g140164(.A (n_34114), .B (n_34115), .C (n_34116), .D(n_34117), .Y (n_34118));
NAND2X1 g140165(.A (n_3498), .B (n_3686), .Y (n_34114));
NAND2X1 g140166(.A (n_3409), .B (n_3686), .Y (n_34115));
NAND2X1 g140167(.A (n_3196), .B (P3_IR[24] ), .Y (n_34116));
NAND2X1 g140168(.A (n_33566), .B (P3_IR[23] ), .Y (n_34117));
NAND2X1 g140169(.A (n_34114), .B (n_34116), .Y (n_34119));
AND2X1 g140170(.A (n_34115), .B (n_34117), .Y (n_34120));
NAND2X2 g140196(.A (n_34159), .B (n_34160), .Y (n_35215));
AOI21X1 g140197(.A0 (n_7944), .A1 (P3_reg1[15] ), .B0 (n_7686), .Y(n_34159));
AOI21X1 g140198(.A0 (P3_reg2[15] ), .A1 (n_8183), .B0 (n_7262), .Y(n_34160));
NAND2X2 g140199(.A (n_15620), .B (n_15727), .Y (n_34163));
NAND2X1 g140201(.A (n_34167), .B (n_35624), .Y (n_34171));
INVX1 g140202(.A (n_34358), .Y (n_34167));
CLKBUFX1 g140207(.A (n_35625), .Y (n_34172));
NAND3X1 g140208(.A (n_34173), .B (n_34175), .C (n_34177), .Y(n_34178));
OR2X1 g140209(.A (n_852), .B (n_1304), .Y (n_34173));
NAND4X1 g140210(.A (n_2782), .B (n_34946), .C (n_2321), .D (n_34174),.Y (n_34175));
AND2X1 g140211(.A (n_1915), .B (P2_IR[26] ), .Y (n_34174));
NAND2X1 g140212(.A (n_34176), .B (n_1305), .Y (n_34177));
NAND3X1 g140213(.A (n_2782), .B (n_2321), .C (n_1915), .Y (n_34176));
CLKBUFX1 g140214(.A (n_34178), .Y (n_34179));
MX2X1 g140215(.A (n_34181), .B (n_34180), .S0 (n_34289), .Y(n_34187));
INVX1 g140216(.A (n_34180), .Y (n_34181));
OAI22X1 g140217(.A0 (n_33004), .A1 (n_12561), .B0 (n_33000), .B1(n_11470), .Y (n_34180));
NAND2X1 g140223(.A (n_34190), .B (n_34194), .Y (n_34195));
NAND2X1 g29(.A (n_34188), .B (n_34189), .Y (n_34190));
INVX1 g140224(.A (n_349), .Y (n_34188));
NAND2X1 g140225(.A (n_31248), .B (n_10481), .Y (n_34189));
NOR2X1 g140226(.A (n_34191), .B (n_34193), .Y (n_34194));
AND2X1 g140227(.A (n_1017), .B (P3_reg3[18] ), .Y (n_34191));
NOR2X1 g28(.A (n_34192), .B (n_12753), .Y (n_34193));
OR2X1 g30(.A (n_7062), .B (n_3493), .Y (n_34192));
INVX1 g31(.A (n_34191), .Y (n_34196));
NAND3X1 g140228(.A (n_34410), .B (n_34199), .C (n_34201), .Y(n_34203));
INVX2 g140232(.A (P3_IR[8] ), .Y (n_34199));
INVX2 g140234(.A (P3_IR[5] ), .Y (n_34201));
CLKBUFX1 g140236(.A (n_34201), .Y (n_34205));
OAI21X1 g140237(.A0 (n_34207), .A1 (n_34206), .B0 (n_34208), .Y(n_34209));
NAND2X1 g140238(.A (n_16771), .B (n_18705), .Y (n_34206));
NAND3X1 g140239(.A (n_33058), .B (n_33055), .C (n_33059), .Y(n_34207));
NAND2X1 g140240(.A (n_34206), .B (n_34207), .Y (n_34208));
NAND2X1 g140241(.A (n_34215), .B (n_35736), .Y (n_34220));
NAND2X1 g140242(.A (n_34212), .B (n_34214), .Y (n_34215));
NAND2X1 g140243(.A (n_34210), .B (n_34211), .Y (n_34212));
NAND3X1 g140244(.A (n_32019), .B (n_22216), .C (n_32020), .Y(n_34210));
NAND2X1 g140245(.A (n_16440), .B (n_17864), .Y (n_34211));
NAND4X1 g140246(.A (n_32019), .B (n_22216), .C (n_32020), .D(n_34213), .Y (n_34214));
INVX1 g140247(.A (n_34211), .Y (n_34213));
NAND3X1 g140251(.A (n_12938), .B (n_12937), .C (n_12902), .Y(n_34216));
NAND4X1 g140252(.A (n_34221), .B (n_34223), .C (n_34225), .D(n_34227), .Y (n_34228));
OR2X1 g140253(.A (n_9172), .B (n_32339), .Y (n_34221));
AOI21X1 g140254(.A0 (n_28926), .A1 (n_32340), .B0 (n_34222), .Y(n_34223));
NOR2X1 g140255(.A (n_28659), .B (n_15282), .Y (n_34222));
NOR2X1 g140256(.A (n_21202), .B (n_34224), .Y (n_34225));
INVX1 g140257(.A (n_27511), .Y (n_34224));
OAI21X1 g140258(.A0 (n_30180), .A1 (n_34226), .B0 (n_30874), .Y(n_34227));
OR2X1 g140259(.A (n_30557), .B (n_33494), .Y (n_34226));
NAND3X1 g140260(.A (n_34229), .B (n_34230), .C (n_34235), .Y(n_34236));
NOR2X1 g140261(.A (n_4284), .B (n_4762), .Y (n_34229));
NOR2X1 g140262(.A (n_35195), .B (n_33485), .Y (n_34230));
AND2X1 g140263(.A (n_35620), .B (n_34234), .Y (n_34235));
NAND2X2 g140265(.A (n_3266), .B (n_1625), .Y (n_34231));
NAND2X2 g140266(.A (n_3720), .B (n_1405), .Y (n_34232));
NOR2X1 g140267(.A (n_2664), .B (n_3240), .Y (n_34234));
INVX1 g140268(.A (n_35620), .Y (n_34237));
INVX1 g140291(.A (n_29924), .Y (n_34258));
NOR2X1 g140292(.A (n_21657), .B (n_25561), .Y (n_34259));
INVX1 g140299(.A (n_30342), .Y (n_34264));
NAND4X1 g140311(.A (n_34285), .B (n_34286), .C (n_34287), .D(n_34288), .Y (n_34289));
NAND3X1 g140312(.A (n_34280), .B (n_34281), .C (n_34284), .Y(n_34285));
NAND2X1 g57_dup(.A (n_21611), .B (n_20624), .Y (n_34280));
INVX1 g140313(.A (n_33703), .Y (n_34281));
NOR2X1 g140314(.A (n_20995), .B (n_34283), .Y (n_34284));
INVX1 g140315(.A (n_34282), .Y (n_34283));
NOR2X1 g140316(.A (n_17760), .B (n_33860), .Y (n_34282));
NAND2X1 g140317(.A (n_20996), .B (n_33711), .Y (n_34286));
NAND2X1 g140318(.A (n_22678), .B (n_20375), .Y (n_34287));
AOI21X1 g140319(.A0 (n_20407), .A1 (n_19041), .B0 (n_20993), .Y(n_34288));
NAND2X1 g140320(.A (n_21611), .B (n_20624), .Y (n_34290));
NAND2X2 g140321(.A (n_34293), .B (n_34297), .Y (n_34298));
AOI21X1 g140322(.A0 (n_15622), .A1 (n_34291), .B0 (n_34292), .Y(n_34293));
NAND2X1 g140323(.A (n_15232), .B (n_15209), .Y (n_34291));
AND2X1 g140324(.A (n_6524), .B (n_3870), .Y (n_34292));
NAND2X1 g140325(.A (n_34291), .B (n_34296), .Y (n_34297));
INVX1 g140326(.A (n_34353), .Y (n_34296));
NAND2X1 g140329(.A (n_34302), .B (n_34306), .Y (n_34307));
NAND2X1 g140330(.A (n_34299), .B (n_34301), .Y (n_34302));
NAND2X1 g140331(.A (n_31377), .B (n_31258), .Y (n_34299));
NOR2X1 g140332(.A (n_34300), .B (n_31564), .Y (n_34301));
CLKBUFX1 g140333(.A (P2_n_749), .Y (n_34300));
AND2X1 g140334(.A (n_34304), .B (n_34305), .Y (n_34306));
OR2X1 g140335(.A (n_34303), .B (n_8732), .Y (n_34304));
OR2X1 g140336(.A (n_34300), .B (n_10414), .Y (n_34303));
AOI22X1 g140337(.A0 (P2_reg3[24] ), .A1 (n_1336), .B0 (n_6446), .B1(n_3835), .Y (n_34305));
INVX1 g140338(.A (n_34300), .Y (n_34308));
INVX1 g140339(.A (P2_n_749), .Y (n_34309));
NAND2X1 g140341(.A (n_28570), .B (n_27469), .Y (n_34310));
AOI21X1 g140343(.A0 (n_28618), .A1 (n_28570), .B0 (n_30445), .Y(n_34314));
NAND2X1 g140345(.A (n_8678), .B (n_8322), .Y (n_34312));
AND2X1 g140347(.A (n_27469), .B (n_28570), .Y (n_34317));
NAND4X1 g140348(.A (n_34318), .B (n_34320), .C (n_34321), .D(n_34323), .Y (n_34324));
AND2X1 g140349(.A (n_32957), .B (n_34538), .Y (n_34318));
CLKBUFX1 g140350(.A (n_34319), .Y (n_34320));
INVX1 g140351(.A (P3_IR[0] ), .Y (n_34319));
INVX2 g140352(.A (P3_IR[4] ), .Y (n_34321));
CLKBUFX1 g140353(.A (n_34322), .Y (n_34323));
INVX2 g140354(.A (P3_IR[1] ), .Y (n_34322));
INVX1 g140359(.A (n_32226), .Y (n_34326));
AND2X1 g140363(.A (n_34310), .B (n_34693), .Y (n_34330));
INVX1 g140366(.A (n_35008), .Y (n_34336));
NAND2X2 g140379(.A (n_34351), .B (n_34356), .Y (n_34357));
AOI21X1 g140380(.A0 (n_15685), .A1 (n_34349), .B0 (n_34350), .Y(n_34351));
NAND2X1 g140381(.A (n_15327), .B (n_15358), .Y (n_34349));
NOR2X1 g140382(.A (n_4351), .B (n_6823), .Y (n_34350));
NAND2X1 g140383(.A (n_34355), .B (n_34349), .Y (n_34356));
CLKBUFX2 g140384(.A (n_34354), .Y (n_34355));
INVX2 g140385(.A (n_34353), .Y (n_34354));
INVX2 g140386(.A (n_34352), .Y (n_34353));
NAND2X2 g140387(.A (n_6368), .B (n_6374), .Y (n_34352));
NOR2X1 g140388(.A (n_34358), .B (n_35624), .Y (n_34362));
NAND2X2 g140389(.A (n_15385), .B (n_15474), .Y (n_34358));
NOR2X1 g140391(.A (n_7144), .B (n_7305), .Y (n_34359));
NAND2X1 g140395(.A (n_34363), .B (n_29910), .Y (n_34364));
INVX1 g140396(.A (n_25539), .Y (n_34363));
NAND2X2 g140402(.A (n_34377), .B (n_34381), .Y (n_34382));
NAND3X1 g140403(.A (n_34372), .B (n_8719), .C (n_34700), .Y(n_34377));
NAND2X1 g140404(.A (n_31378), .B (n_30960), .Y (n_34372));
INVX1 g140407(.A (n_34700), .Y (n_34375));
NOR2X1 g140409(.A (n_34378), .B (n_34380), .Y (n_34381));
AND2X1 g140410(.A (n_6429), .B (n_10082), .Y (n_34378));
NOR2X1 g140411(.A (n_34379), .B (n_8782), .Y (n_34380));
OR2X1 g140412(.A (P2_n_749), .B (n_9934), .Y (n_34379));
NAND2X1 g140413(.A (n_34384), .B (n_34385), .Y (n_34386));
CLKBUFX1 g140414(.A (n_34383), .Y (n_34384));
NAND4X1 g140415(.A (n_7563), .B (n_7925), .C (n_7920), .D (n_7582),.Y (n_34383));
NAND2X1 g140416(.A (n_15861), .B (n_16230), .Y (n_34385));
INVX1 g140417(.A (n_34385), .Y (n_34387));
XOR2X1 g140418(.A (n_34388), .B (n_34392), .Y (n_34393));
AND2X1 g140419(.A (n_2454), .B (n_4425), .Y (n_34388));
NAND2X2 g140420(.A (n_34389), .B (n_34391), .Y (n_34392));
NAND2X1 g140421(.A (n_33300), .B (n_33303), .Y (n_34389));
NOR2X1 g140422(.A (n_34390), .B (n_34920), .Y (n_34391));
AND2X1 g140423(.A (n_2429), .B (n_4113), .Y (n_34390));
AOI21X1 g140425(.A0 (n_33300), .A1 (n_33303), .B0 (n_34920), .Y(n_34395));
INVX1 g140426(.A (n_34390), .Y (n_34396));
NAND4X1 g140427(.A (n_35897), .B (n_34399), .C (n_35898), .D(n_34403), .Y (n_35933));
INVX1 g140428(.A (n_34364), .Y (n_35898));
NOR2X1 g140429(.A (n_34398), .B (n_33416), .Y (n_34399));
NAND2X1 g140430(.A (n_30187), .B (n_33420), .Y (n_34398));
NOR2X1 g140431(.A (n_34400), .B (n_34401), .Y (n_35897));
AOI21X1 g140432(.A0 (n_8718), .A1 (n_30355), .B0 (n_30478), .Y(n_34400));
INVX1 g140433(.A (n_33419), .Y (n_34401));
NAND2X1 g140434(.A (n_29767), .B (n_33802), .Y (n_34403));
NOR2X1 g140435(.A (n_34405), .B (n_34411), .Y (n_34412));
NAND3X1 g140436(.A (n_1939), .B (n_32957), .C (n_34538), .Y(n_34405));
NAND3X1 g140437(.A (n_34526), .B (n_34408), .C (n_34410), .Y(n_34411));
INVX1 g140439(.A (n_34407), .Y (n_34408));
NAND2X1 g140440(.A (n_34321), .B (n_34201), .Y (n_34407));
INVX2 g140441(.A (n_34409), .Y (n_34410));
NAND2X2 g140442(.A (n_117), .B (n_216), .Y (n_34409));
NAND2X1 g140443(.A (n_34416), .B (P1_reg1[30] ), .Y (n_34417));
INVX2 g140444(.A (n_34415), .Y (n_34416));
NOR2X1 g140445(.A (n_34413), .B (n_34987), .Y (n_34415));
NAND2X1 g140446(.A (n_12659), .B (n_11940), .Y (n_34413));
INVX2 g140449(.A (n_34416), .Y (n_34418));
NAND4X1 g140450(.A (n_34421), .B (n_34422), .C (n_30026), .D(n_34426), .Y (n_34427));
AOI21X1 g140451(.A0 (n_30027), .A1 (n_34952), .B0 (n_34420), .Y(n_34421));
INVX1 g140452(.A (n_30004), .Y (n_34420));
AOI21X1 g140453(.A0 (n_26571), .A1 (n_8303), .B0 (n_15487), .Y(n_34422));
AOI21X1 g140454(.A0 (n_30005), .A1 (n_25756), .B0 (n_34425), .Y(n_34426));
NAND2X1 g140455(.A (n_34423), .B (n_34424), .Y (n_34425));
NAND3X1 g140456(.A (n_10848), .B (n_8212), .C (n_8213), .Y (n_34423));
OR4X1 g140457(.A (n_8011), .B (n_7344), .C (n_6833), .D (n_7536), .Y(n_34424));
NOR2X1 g140458(.A (n_34428), .B (n_34433), .Y (n_34434));
NAND2X1 g140459(.A (n_3438), .B (n_1279), .Y (n_34428));
NAND3X1 g140460(.A (n_34431), .B (n_34432), .C (n_3657), .Y(n_34433));
NOR2X1 g140461(.A (n_34429), .B (n_34430), .Y (n_34431));
NAND3X1 g140462(.A (n_1647), .B (n_1019), .C (n_1013), .Y (n_34429));
NOR2X1 g140463(.A (n_3474), .B (n_3036), .Y (n_34430));
OR2X1 g140464(.A (n_3596), .B (n_3156), .Y (n_34432));
NAND2X1 g140465(.A (n_3957), .B (n_34438), .Y (n_34439));
OAI21X1 g140467(.A0 (n_3156), .A1 (n_3596), .B0 (n_1019), .Y(n_34435));
INVX1 g140468(.A (n_34437), .Y (n_34438));
OAI21X1 g140469(.A0 (n_3036), .A1 (n_3474), .B0 (n_1013), .Y(n_34437));
NAND2X2 g140470(.A (n_3657), .B (n_1647), .Y (n_34440));
NOR2X1 g140473(.A (n_34722), .B (n_19091), .Y (n_34441));
INVX1 g140478(.A (n_34445), .Y (n_34446));
NAND2X1 g140479(.A (n_34724), .B (n_19302), .Y (n_34445));
AND2X1 g140480(.A (n_34807), .B (n_34808), .Y (n_34450));
NOR2X1 g140483(.A (n_34451), .B (n_34452), .Y (n_34453));
NOR2X1 g140484(.A (n_9009), .B (n_29923), .Y (n_34451));
AOI21X1 g140485(.A0 (n_30445), .A1 (n_8285), .B0 (n_34264), .Y(n_34452));
NAND2X1 g140487(.A (n_34753), .B (n_30342), .Y (n_34455));
NAND3X1 g140495(.A (n_34465), .B (n_34467), .C (n_34470), .Y(n_34471));
OR2X1 g140496(.A (n_3450), .B (n_7340), .Y (n_34465));
NAND2X1 g140497(.A (n_15387), .B (n_34466), .Y (n_34467));
NAND2X1 g140498(.A (n_14911), .B (n_14901), .Y (n_34466));
NAND2X1 g140499(.A (n_34469), .B (n_34466), .Y (n_34470));
INVX4 g140500(.A (n_34468), .Y (n_34469));
NAND2X2 g140501(.A (n_6403), .B (n_6337), .Y (n_34468));
INVX4 g140502(.A (n_34469), .Y (n_34472));
AND2X1 g140503(.A (n_34948), .B (n_34482), .Y (n_34483));
NAND2X1 g140513(.A (n_3761), .B (n_1877), .Y (n_34482));
INVX1 g140514(.A (n_34948), .Y (n_34484));
INVX1 g140515(.A (n_34482), .Y (n_34485));
NAND3X1 g140517(.A (n_34489), .B (n_34490), .C (n_34492), .Y(n_34493));
NAND2X1 g140518(.A (n_34487), .B (n_34488), .Y (n_34489));
NOR2X1 g140519(.A (n_19915), .B (n_17224), .Y (n_34487));
OAI21X1 g140520(.A0 (n_23047), .A1 (n_21425), .B0 (n_22212), .Y(n_34488));
NAND3X1 g140521(.A (n_23360), .B (n_34487), .C (n_20948), .Y(n_34490));
INVX1 g140522(.A (n_34491), .Y (n_34492));
OAI21X1 g140523(.A0 (n_20356), .A1 (n_19915), .B0 (n_20355), .Y(n_34491));
AOI21X1 g140524(.A0 (n_34496), .A1 (n_34499), .B0 (n_34500), .Y(n_34501));
NAND2X2 g140525(.A (n_34494), .B (n_34495), .Y (n_34496));
NAND2X1 g140526(.A (n_24257), .B (n_18345), .Y (n_34494));
NAND2X1 g140527(.A (n_23225), .B (n_34765), .Y (n_34495));
INVX2 g140528(.A (n_34498), .Y (n_34499));
CLKBUFX3 g140529(.A (n_34497), .Y (n_34498));
NAND2X2 g140530(.A (n_13065), .B (n_13067), .Y (n_34497));
AND2X1 g140531(.A (n_13665), .B (P2_reg_106), .Y (n_34500));
NAND3X1 g140532(.A (n_34504), .B (n_34505), .C (n_34506), .Y(n_34507));
NOR2X1 g140533(.A (n_34502), .B (n_34503), .Y (n_34504));
NAND2X1 g140534(.A (n_3621), .B (n_3462), .Y (n_34502));
NAND2X1 g140535(.A (n_35380), .B (n_3566), .Y (n_34503));
NOR2X1 g140536(.A (n_3971), .B (n_35391), .Y (n_34505));
NOR2X1 g140537(.A (n_3925), .B (n_4328), .Y (n_34506));
NOR2X1 g140538(.A (n_34508), .B (n_34513), .Y (n_34514));
NAND3X1 g140539(.A (n_21418), .B (n_21489), .C (n_19256), .Y(n_34508));
AOI21X1 g140540(.A0 (n_23676), .A1 (n_22351), .B0 (n_34512), .Y(n_34513));
NAND2X1 g140541(.A (n_19059), .B (n_34511), .Y (n_34512));
NAND2X1 g140543(.A (n_19230), .B (n_18466), .Y (n_34509));
AND2X1 g140544(.A (n_20411), .B (n_20408), .Y (n_34511));
NAND2X1 g140545(.A (n_23676), .B (n_22351), .Y (n_34515));
NAND3X1 g140546(.A (n_34518), .B (n_34519), .C (n_34520), .Y(n_34521));
NAND2X1 g140547(.A (n_34516), .B (n_34517), .Y (n_34518));
NAND2X1 g23_dup(.A (n_22713), .B (n_21930), .Y (n_34516));
AND2X1 g140548(.A (n_21472), .B (n_35179), .Y (n_34517));
OR2X1 g140549(.A (n_33180), .B (n_33181), .Y (n_34519));
AND2X1 g140550(.A (n_33185), .B (n_33183), .Y (n_34520));
NAND2X1 g140551(.A (n_21930), .B (n_22713), .Y (n_34522));
INVX1 g140552(.A (n_34525), .Y (n_34526));
NAND4X1 g140553(.A (n_34849), .B (n_34524), .C (n_34199), .D(n_34850), .Y (n_34525));
INVX1 g140555(.A (P3_IR[11] ), .Y (n_34524));
NAND2X1 g140556(.A (n_34849), .B (n_34524), .Y (n_34527));
NAND2X1 g140557(.A (n_34199), .B (n_34850), .Y (n_34528));
NAND2X1 g140558(.A (n_34532), .B (n_34534), .Y (n_34535));
INVX2 g140559(.A (n_34531), .Y (n_34532));
NAND2X2 g140560(.A (n_34529), .B (n_34530), .Y (n_34531));
NAND2X1 g140561(.A (n_35401), .B (n_6160), .Y (n_34529));
NAND3X1 g140562(.A (n_6180), .B (n_32219), .C (n_6179), .Y (n_34530));
INVX2 g140563(.A (n_34533), .Y (n_34534));
MX2X1 g140564(.A (n_4471), .B (n_6180), .S0 (n_6179), .Y (n_34533));
NOR2X1 g140565(.A (n_34536), .B (n_34542), .Y (n_34543));
NAND3X1 g35(.A (n_32566), .B (n_1753), .C (n_34849), .Y (n_34536));
NAND3X1 g140566(.A (n_34537), .B (n_34540), .C (n_34541), .Y(n_34542));
NOR2X1 g140567(.A (n_32956), .B (n_722), .Y (n_34537));
NOR2X1 g140568(.A (n_1218), .B (n_34539), .Y (n_34540));
INVX1 g140569(.A (n_34538), .Y (n_34539));
INVX1 g140570(.A (P3_IR[3] ), .Y (n_34538));
INVX1 g140571(.A (n_34407), .Y (n_34541));
INVX1 g140572(.A (n_34539), .Y (n_34544));
OAI21X1 g140574(.A0 (n_16285), .A1 (n_15808), .B0 (n_15905), .Y(n_34545));
AND2X1 g140575(.A (n_16076), .B (n_16284), .Y (n_34546));
NAND2X1 g140576(.A (n_34547), .B (n_34548), .Y (n_34549));
NAND2X1 g140577(.A (n_16245), .B (n_16284), .Y (n_34547));
NAND2X1 g140578(.A (n_15752), .B (n_9688), .Y (n_34548));
NAND3X1 g140579(.A (n_35266), .B (n_34555), .C (n_35267), .Y(n_34557));
OR2X1 g140580(.A (n_34551), .B (n_34552), .Y (n_35267));
AOI21X1 g140581(.A0 (n_34545), .A1 (n_34546), .B0 (n_34549), .Y(n_34551));
NAND2X1 g140582(.A (n_17585), .B (n_17584), .Y (n_34552));
INVX1 g140583(.A (n_34554), .Y (n_34555));
NAND2X1 g140584(.A (n_17609), .B (n_17499), .Y (n_34554));
NAND3X1 g140585(.A (n_18134), .B (n_19407), .C (n_16042), .Y(n_35266));
NAND2X2 g140594(.A (n_34919), .B (n_34573), .Y (n_34574));
NAND4X1 g140597(.A (n_34568), .B (n_34569), .C (n_34571), .D(n_34572), .Y (n_34573));
NOR2X1 g140598(.A (n_4512), .B (n_5257), .Y (n_34568));
INVX1 g140599(.A (n_4930), .Y (n_34569));
NOR2X1 g140600(.A (n_34570), .B (n_4518), .Y (n_34571));
NAND2X1 g140601(.A (n_3289), .B (n_3162), .Y (n_34570));
NOR2X1 g140602(.A (n_3176), .B (n_3744), .Y (n_34572));
CLKBUFX1 g140603(.A (n_34580), .Y (n_34581));
NAND2X1 g140604(.A (n_9720), .B (n_34579), .Y (n_34580));
NAND2X2 g140606(.A (n_8191), .B (n_7711), .Y (n_34575));
NAND2X1 g140607(.A (n_34577), .B (n_34578), .Y (n_34579));
NAND2X1 g140608(.A (n_15581), .B (n_15375), .Y (n_34577));
NAND2X1 g140609(.A (n_4301), .B (n_7132), .Y (n_34578));
AOI21X1 g140610(.A0 (n_34586), .A1 (P3_reg1[5] ), .B0 (n_34591), .Y(n_34592));
INVX1 g140611(.A (n_34585), .Y (n_34586));
INVX1 g140612(.A (n_34584), .Y (n_34585));
AND2X1 g140613(.A (n_34582), .B (n_34583), .Y (n_34584));
MX2X1 g140614(.A (n_5015), .B (n_34388), .S0 (n_34392), .Y (n_34582));
MX2X1 g140615(.A (n_34396), .B (n_4627), .S0 (n_34395), .Y (n_34583));
AND2X1 g140616(.A (n_34587), .B (n_34590), .Y (n_34591));
NAND2X1 g140617(.A (n_2369), .B (n_2259), .Y (n_34587));
INVX2 g140618(.A (n_34589), .Y (n_34590));
INVX2 g140619(.A (n_34588), .Y (n_34589));
AND2X1 g140620(.A (n_34393), .B (n_34583), .Y (n_34588));
MX2X1 g140621(.A (n_4627), .B (n_34396), .S0 (n_34395), .Y (n_34595));
NAND3X1 g140624(.A (n_34598), .B (n_34600), .C (n_34603), .Y(n_34604));
NAND2X1 g140625(.A (n_34597), .B (n_22374), .Y (n_34598));
INVX1 g140626(.A (n_34596), .Y (n_34597));
NAND2X1 g140627(.A (n_19046), .B (n_19047), .Y (n_34596));
INVX1 g140628(.A (n_34599), .Y (n_34600));
NAND2X1 g140629(.A (n_19757), .B (n_20493), .Y (n_34599));
NAND3X1 g140630(.A (n_34602), .B (n_21363), .C (n_34557), .Y(n_34603));
NOR2X1 g140631(.A (n_34601), .B (n_34596), .Y (n_34602));
NAND2X1 g140632(.A (n_35001), .B (n_19306), .Y (n_34601));
AND2X1 g140633(.A (n_21363), .B (n_34557), .Y (n_34605));
INVX1 g140634(.A (n_34601), .Y (n_34606));
NAND4X1 g140635(.A (n_34611), .B (n_12314), .C (n_34614), .D(n_16796), .Y (n_34615));
NOR3X1 g140636(.A (n_34610), .B (n_12195), .C (n_12866), .Y(n_34611));
INVX2 g140637(.A (n_34609), .Y (n_34610));
CLKBUFX1 g140638(.A (n_34608), .Y (n_34609));
CLKBUFX1 g140639(.A (n_34607), .Y (n_34608));
NAND2X2 g140640(.A (n_32286), .B (n_32287), .Y (n_34607));
NOR2X1 g140641(.A (n_34612), .B (n_34613), .Y (n_34614));
NAND2X1 g140642(.A (n_11747), .B (n_18475), .Y (n_34612));
NAND3X1 g140643(.A (n_11247), .B (n_32350), .C (n_11464), .Y(n_34613));
NOR2X1 g140644(.A (n_12195), .B (n_12866), .Y (n_34616));
INVX2 g140645(.A (n_34607), .Y (n_34617));
CLKBUFX1 g140669(.A (n_34645), .Y (n_34646));
NAND2X1 g140670(.A (n_35086), .B (n_35087), .Y (n_34645));
NAND2X1 g140671(.A (n_34641), .B (n_34642), .Y (n_35087));
NAND2X1 g140672(.A (n_16695), .B (n_16662), .Y (n_34641));
NOR2X1 g140673(.A (n_16568), .B (n_16567), .Y (n_34642));
AOI21X1 g140674(.A0 (n_17585), .A1 (n_34549), .B0 (n_17608), .Y(n_35086));
NAND3X1 g140676(.A (n_34648), .B (n_34649), .C (n_34650), .Y(n_34651));
AOI21X1 g140677(.A0 (n_14135), .A1 (n_7983), .B0 (n_34647), .Y(n_34648));
NOR2X1 g140678(.A (n_296), .B (n_7823), .Y (n_34647));
OR2X1 g140679(.A (n_185), .B (n_7917), .Y (n_34649));
NAND3X1 g140680(.A (n_8213), .B (n_8212), .C (n_7476), .Y (n_34650));
NAND2X2 g140693(.A (n_34673), .B (n_34674), .Y (n_34675));
NAND2X1 g140694(.A (n_34668), .B (n_34672), .Y (n_34673));
INVX1 g140695(.A (n_35017), .Y (n_34668));
NAND2X1 g140699(.A (n_31638), .B (n_34671), .Y (n_34672));
NAND2X1 g140700(.A (n_34669), .B (n_34670), .Y (n_34671));
INVX1 g140701(.A (n_8334), .Y (n_34669));
INVX1 g140702(.A (n_31881), .Y (n_34670));
NAND2X1 g140703(.A (n_6979), .B (n_10152), .Y (n_34674));
INVX1 g140704(.A (n_35023), .Y (n_34676));
AOI21X1 g140705(.A0 (n_34677), .A1 (n_34678), .B0 (n_34682), .Y(n_34683));
NOR2X1 g140706(.A (n_17314), .B (n_17326), .Y (n_34677));
NAND2X2 g140707(.A (n_19655), .B (n_18860), .Y (n_34678));
NAND2X2 g140708(.A (n_34679), .B (n_34681), .Y (n_34682));
NAND2X1 g140709(.A (n_18578), .B (n_19198), .Y (n_34679));
INVX1 g140710(.A (n_34680), .Y (n_34681));
OAI21X1 g140711(.A0 (n_32901), .A1 (n_18012), .B0 (n_17256), .Y(n_34680));
NAND2X1 g140712(.A (n_34692), .B (n_34694), .Y (n_34695));
INVX1 g140713(.A (n_34691), .Y (n_34692));
AND2X1 g140714(.A (n_34689), .B (n_34690), .Y (n_34691));
NAND2X1 g140715(.A (n_34684), .B (n_34688), .Y (n_34689));
MX2X1 g140716(.A (n_19051), .B (n_20241), .S0 (n_23890), .Y(n_34684));
CLKBUFX3 g140717(.A (n_34687), .Y (n_34688));
INVX2 g140718(.A (n_34686), .Y (n_34687));
CLKBUFX3 g140719(.A (n_34685), .Y (n_34686));
NAND2X2 g140720(.A (n_13054), .B (n_13053), .Y (n_34685));
NAND2X1 g140721(.A (n_13854), .B (n_3191), .Y (n_34690));
CLKBUFX1 g140722(.A (n_34693), .Y (n_34694));
NOR2X1 g140723(.A (n_7782), .B (n_7777), .Y (n_34693));
INVX2 g140724(.A (n_34684), .Y (n_34696));
NAND2X2 g140725(.A (n_34702), .B (n_34703), .Y (n_34704));
NAND4X1 g140726(.A (n_34697), .B (n_34698), .C (n_34699), .D(n_34701), .Y (n_34702));
NAND2X1 g140727(.A (n_31548), .B (n_31453), .Y (n_34697));
OR2X1 g140728(.A (n_32641), .B (n_6061), .Y (n_34698));
NAND2X1 g140729(.A (n_6061), .B (n_32641), .Y (n_34699));
CLKBUFX1 g140730(.A (n_34700), .Y (n_34701));
INVX1 g140731(.A (P2_n_749), .Y (n_34700));
AOI22X1 g140732(.A0 (n_6460), .A1 (n_12674), .B0 (n_1812), .B1(n_8687), .Y (n_34703));
INVX1 g140734(.A (n_35007), .Y (n_34706));
NOR2X1 g140735(.A (n_34711), .B (n_34716), .Y (n_34717));
AOI21X1 g140736(.A0 (n_27710), .A1 (n_27131), .B0 (n_27696), .Y(n_34711));
BUFX3 g140739(.A (n_34708), .Y (n_34709));
NOR2X1 g140740(.A (n_7325), .B (n_8948), .Y (n_34708));
NOR2X1 g140741(.A (n_34713), .B (n_34715), .Y (n_34716));
INVX1 g140742(.A (n_34712), .Y (n_34713));
NAND2X2 g140743(.A (n_33807), .B (n_33505), .Y (n_34712));
INVX1 g140744(.A (n_34714), .Y (n_34715));
NAND2X1 g140745(.A (n_26656), .B (n_27710), .Y (n_34714));
NAND2X1 g140746(.A (n_27131), .B (n_27710), .Y (n_34718));
INVX4 g140747(.A (n_34708), .Y (n_34719));
AND2X1 g140748(.A (n_34723), .B (n_34724), .Y (n_34725));
INVX1 g140749(.A (n_34722), .Y (n_34723));
NAND2X2 g140750(.A (n_34720), .B (n_34721), .Y (n_34722));
NAND2X1 g140751(.A (n_16161), .B (n_16160), .Y (n_34720));
NAND2X2 g140752(.A (n_16140), .B (n_16429), .Y (n_34721));
AND2X1 g140753(.A (n_17767), .B (n_32839), .Y (n_34724));
NAND2X1 g140754(.A (n_34732), .B (n_34736), .Y (n_34737));
OAI21X1 g140755(.A0 (n_35084), .A1 (n_35085), .B0 (n_34731), .Y(n_34732));
NAND4X1 g140756(.A (n_32571), .B (n_34726), .C (n_30064), .D(n_32112), .Y (n_35085));
AND2X1 g140757(.A (n_30017), .B (n_27794), .Y (n_34726));
NAND2X1 g140758(.A (n_32570), .B (n_30567), .Y (n_35084));
CLKBUFX1 g140759(.A (n_35008), .Y (n_34731));
NAND2X1 g140762(.A (n_34733), .B (n_6349), .Y (n_34736));
NOR2X1 g140763(.A (P2_reg_113), .B (n_9310), .Y (n_34733));
INVX1 g140766(.A (n_35012), .Y (n_34738));
INVX1 g140767(.A (n_34731), .Y (n_34739));
NOR2X1 g140768(.A (n_34743), .B (n_34744), .Y (n_34745));
INVX1 g140769(.A (n_34742), .Y (n_34743));
AND2X1 g140770(.A (n_34740), .B (n_34741), .Y (n_34742));
NAND2X2 g140771(.A (n_16036), .B (n_9652), .Y (n_34740));
NAND2X1 g140772(.A (n_15870), .B (n_10275), .Y (n_34741));
NAND2X1 g140773(.A (n_35059), .B (n_17482), .Y (n_34744));
INVX1 g140774(.A (n_34740), .Y (n_34746));
OR2X1 g140779(.A (n_34326), .B (n_21656), .Y (n_34749));
NAND2X1 g140781(.A (n_28618), .B (n_28570), .Y (n_34751));
INVX4 g140782(.A (n_34752), .Y (n_34753));
NAND3X1 g140783(.A (n_7763), .B (n_6878), .C (n_6837), .Y (n_34752));
NAND2X1 g140784(.A (n_34758), .B (n_34764), .Y (n_34765));
AOI21X1 g140785(.A0 (n_20307), .A1 (n_21406), .B0 (n_34757), .Y(n_34758));
NAND2X1 g53_dup(.A (n_34756), .B (n_19033), .Y (n_34757));
OR2X1 g140786(.A (n_16869), .B (n_20970), .Y (n_34756));
OAI21X1 g140787(.A0 (n_34762), .A1 (n_22540), .B0 (n_34763), .Y(n_34764));
NOR2X1 g140788(.A (n_20255), .B (n_34761), .Y (n_34762));
NAND2X1 g140789(.A (n_20011), .B (n_34760), .Y (n_34761));
NAND2X1 g140791(.A (n_20519), .B (n_19344), .Y (n_34760));
NOR2X1 g140792(.A (n_20960), .B (n_19201), .Y (n_34763));
NAND2X1 g140793(.A (n_19033), .B (n_34756), .Y (n_34766));
CLKBUFX1 g140794(.A (n_34760), .Y (n_34767));
NOR2X1 g140795(.A (n_34768), .B (n_20255), .Y (n_34769));
INVX1 g140796(.A (n_20011), .Y (n_34768));
NOR2X1 g140797(.A (n_34771), .B (n_34775), .Y (n_34776));
INVX1 g140798(.A (n_34770), .Y (n_34771));
NAND2X2 g140799(.A (n_10067), .B (n_8305), .Y (n_34770));
INVX1 g140800(.A (n_34774), .Y (n_34775));
NAND2X2 g140801(.A (n_34772), .B (n_34773), .Y (n_34774));
NAND2X2 g140802(.A (n_21092), .B (n_27983), .Y (n_34772));
NAND2X1 g140803(.A (n_13185), .B (n_10169), .Y (n_34773));
OAI21X1 g140804(.A0 (n_34930), .A1 (n_34781), .B0 (n_35009), .Y(n_34784));
OAI21X1 g140806(.A0 (n_34317), .A1 (n_34779), .B0 (n_34780), .Y(n_34781));
INVX1 g140808(.A (n_30197), .Y (n_34779));
AOI21X1 g140809(.A0 (n_34751), .A1 (n_30369), .B0 (n_34330), .Y(n_34780));
NAND2X1 g140825(.A (n_34801), .B (n_34802), .Y (n_34803));
NAND2X2 g140826(.A (n_34799), .B (n_34800), .Y (n_34801));
NAND2X2 g140827(.A (n_25290), .B (n_25298), .Y (n_34799));
NAND2X1 g140828(.A (n_13850), .B (n_9337), .Y (n_34800));
NOR2X1 g140829(.A (n_6974), .B (n_7561), .Y (n_34802));
NAND3X1 g140830(.A (n_34804), .B (n_34806), .C (n_34809), .Y(n_34810));
NAND2X1 g140831(.A (n_22733), .B (n_34441), .Y (n_34804));
INVX1 g140832(.A (n_34805), .Y (n_34806));
NAND2X1 g140833(.A (n_20303), .B (n_19542), .Y (n_34805));
NAND4X1 g140834(.A (n_34807), .B (n_34441), .C (n_34808), .D(n_34446), .Y (n_34809));
NAND3X1 g140835(.A (n_20616), .B (n_21071), .C (n_20522), .Y(n_34807));
NOR2X1 g140836(.A (n_18628), .B (n_18636), .Y (n_34808));
OAI21X1 g140837(.A0 (n_34814), .A1 (n_34817), .B0 (n_35008), .Y(n_34819));
NAND4X1 g140838(.A (n_35073), .B (n_32187), .C (n_34813), .D(n_35074), .Y (n_34814));
INVX1 g140839(.A (n_28339), .Y (n_35074));
NOR2X1 g140840(.A (n_34812), .B (n_28251), .Y (n_34813));
NAND2X1 g140841(.A (n_10033), .B (n_17698), .Y (n_34812));
NAND2X1 g140842(.A (n_34815), .B (n_34816), .Y (n_34817));
AOI21X1 g140843(.A0 (n_28864), .A1 (n_28850), .B0 (n_28253), .Y(n_34815));
AOI21X1 g140844(.A0 (n_29008), .A1 (n_28850), .B0 (n_26012), .Y(n_34816));
NAND3X1 g140846(.A (n_34820), .B (n_34821), .C (n_34833), .Y(n_34834));
NAND2X1 g140847(.A (n_22508), .B (n_23552), .Y (n_34820));
NAND2X1 g140848(.A (n_22939), .B (n_21766), .Y (n_34821));
AND2X1 g140849(.A (n_34827), .B (n_34832), .Y (n_34833));
NAND2X1 g140850(.A (n_34823), .B (n_34826), .Y (n_34827));
NAND2X1 g140851(.A (n_34822), .B (n_18425), .Y (n_34823));
OR2X1 g140852(.A (n_21813), .B (n_17241), .Y (n_34822));
INVX1 g140853(.A (n_34825), .Y (n_34826));
NAND2X1 g140854(.A (n_34824), .B (n_19236), .Y (n_34825));
AND2X1 g140855(.A (n_17356), .B (n_17901), .Y (n_34824));
NOR2X1 g140856(.A (n_34828), .B (n_34831), .Y (n_34832));
OAI21X1 g140857(.A0 (n_19799), .A1 (n_19294), .B0 (n_18479), .Y(n_34828));
NOR2X1 g140858(.A (n_34829), .B (n_34830), .Y (n_34831));
INVX1 g140859(.A (n_34824), .Y (n_34829));
AND2X1 g140860(.A (n_16832), .B (n_17843), .Y (n_34830));
MX2X1 g140861(.A (n_34836), .B (n_34835), .S0 (n_34837), .Y(n_34838));
INVX1 g140862(.A (n_34835), .Y (n_34836));
NAND2X1 g140863(.A (n_16450), .B (n_35949), .Y (n_34835));
NAND2X1 g140864(.A (n_23267), .B (n_23520), .Y (n_34837));
INVX2 g140865(.A (n_34844), .Y (n_34845));
OR2X1 g140866(.A (n_34842), .B (n_34843), .Y (n_34844));
INVX1 g140867(.A (n_34841), .Y (n_34842));
AND2X1 g140868(.A (n_35849), .B (n_34981), .Y (n_34841));
NAND2X2 g140869(.A (n_9730), .B (n_15753), .Y (n_35849));
NAND2X1 g140871(.A (n_16619), .B (n_34581), .Y (n_34843));
NOR2X1 g140875(.A (n_34851), .B (n_34852), .Y (n_34853));
NAND2X1 g140876(.A (n_34849), .B (n_34850), .Y (n_34851));
INVX2 g140877(.A (P3_IR[10] ), .Y (n_34849));
INVX1 g140878(.A (P3_IR[9] ), .Y (n_34850));
NAND2X1 g140879(.A (n_564), .B (n_34524), .Y (n_34852));
NAND3X1 g140880(.A (n_34856), .B (n_34857), .C (n_34858), .Y(n_34859));
NAND2X1 g140881(.A (n_34854), .B (n_34855), .Y (n_34856));
NAND2X1 g33_dup140882(.A (n_23656), .B (n_33859), .Y (n_34854));
AND2X1 g140883(.A (n_21415), .B (n_21416), .Y (n_34855));
AOI21X1 g140884(.A0 (n_20993), .A1 (n_20406), .B0 (n_20343), .Y(n_34857));
NAND2X1 g140885(.A (n_21297), .B (n_21415), .Y (n_34858));
NAND2X1 g140886(.A (n_33859), .B (n_23656), .Y (n_34860));
OR2X1 g140887(.A (n_34865), .B (n_34871), .Y (n_34872));
NAND3X1 g140888(.A (n_34861), .B (n_34863), .C (n_34864), .Y(n_34865));
INVX1 g140889(.A (n_12588), .Y (n_34861));
INVX1 g140890(.A (n_34862), .Y (n_34863));
NAND3X1 g140891(.A (n_11267), .B (n_11555), .C (n_16904), .Y(n_34862));
INVX1 g140892(.A (n_11538), .Y (n_34864));
NAND2X1 g140893(.A (n_34866), .B (n_34870), .Y (n_34871));
NOR2X1 g140894(.A (n_11309), .B (n_12037), .Y (n_34866));
NOR2X1 g140895(.A (n_34868), .B (n_34869), .Y (n_34870));
INVX1 g140896(.A (n_34867), .Y (n_34868));
NOR2X1 g140897(.A (n_9744), .B (n_16011), .Y (n_34867));
NAND2X1 g140898(.A (n_12977), .B (n_12943), .Y (n_34869));
INVX1 g140899(.A (n_34870), .Y (n_34873));
NOR2X1 g59_dup(.A (n_12588), .B (n_11538), .Y (n_34874));
NOR2X1 g140900(.A (n_12588), .B (n_11538), .Y (n_34875));
INVX1 g140922(.A (n_34913), .Y (n_34915));
INVX2 g47(.A (n_34912), .Y (n_34913));
OAI21X1 g140924(.A0 (n_4279), .A1 (n_1659), .B0 (n_1921), .Y(n_34912));
AOI21X1 g43_dup(.A0 (n_34916), .A1 (n_34918), .B0 (n_34920), .Y(n_34921));
INVX1 g140925(.A (n_32202), .Y (n_34916));
NOR2X1 g49_dup(.A (n_34917), .B (n_5462), .Y (n_34918));
OR2X1 g140926(.A (n_3960), .B (n_3197), .Y (n_34917));
INVX1 g140927(.A (n_34919), .Y (n_34920));
OAI21X1 g140928(.A0 (n_4371), .A1 (n_4087), .B0 (n_33305), .Y(n_34919));
AOI21X1 g140929(.A0 (n_34916), .A1 (n_34923), .B0 (n_34920), .Y(n_34924));
NOR2X1 g140930(.A (n_34917), .B (n_5462), .Y (n_34923));
NAND4X1 g140931(.A (n_34925), .B (n_34926), .C (n_34927), .D(n_34929), .Y (n_34930));
OR2X1 g140932(.A (n_9009), .B (n_34317), .Y (n_34925));
NOR2X1 g140933(.A (n_34749), .B (n_34314), .Y (n_34926));
NAND2X1 g140934(.A (n_34753), .B (n_34751), .Y (n_34927));
INVX1 g140935(.A (n_34928), .Y (n_34929));
OAI21X1 g140936(.A0 (n_15294), .A1 (n_8614), .B0 (n_25222), .Y(n_34928));
NAND3X1 g140937(.A (n_34938), .B (n_34931), .C (n_34939), .Y(n_34940));
NOR2X1 g140938(.A (n_9628), .B (n_10710), .Y (n_34931));
INVX2 g140939(.A (n_34937), .Y (n_34938));
NAND2X2 g140940(.A (n_34933), .B (n_34936), .Y (n_34937));
INVX2 g140941(.A (n_34932), .Y (n_34933));
NAND2X2 g140942(.A (n_32856), .B (n_10796), .Y (n_34932));
CLKBUFX1 g140943(.A (n_34935), .Y (n_34936));
CLKBUFX1 g140944(.A (n_34934), .Y (n_34935));
NAND2X2 g140945(.A (n_7367), .B (n_7646), .Y (n_34934));
NOR2X1 g140946(.A (n_10331), .B (n_10267), .Y (n_34939));
AOI21X1 g140947(.A0 (n_34941), .A1 (n_34943), .B0 (n_34947), .Y(n_34948));
INVX1 g140948(.A (n_34236), .Y (n_34941));
NOR2X1 g140949(.A (n_34942), .B (n_34080), .Y (n_34943));
NAND2X1 g140950(.A (n_4138), .B (n_3174), .Y (n_34942));
NAND3X1 g140951(.A (n_34944), .B (n_34945), .C (n_34946), .Y(n_34947));
INVX1 g140952(.A (n_3592), .Y (n_34944));
INVX1 g140953(.A (n_2708), .Y (n_34945));
CLKBUFX3 g140954(.A (P2_IR[31] ), .Y (n_34946));
NAND3X1 g140956(.A (n_34954), .B (n_34957), .C (n_34961), .Y(n_34962));
NOR2X1 g140957(.A (n_34953), .B (n_30604), .Y (n_34954));
AND2X1 g140958(.A (n_34950), .B (n_34952), .Y (n_34953));
NAND2X1 g140959(.A (n_28633), .B (n_29132), .Y (n_34950));
INVX4 g140960(.A (n_34951), .Y (n_34952));
NOR2X1 g140961(.A (n_34802), .B (n_10196), .Y (n_34951));
AND2X1 g140962(.A (n_34955), .B (n_34956), .Y (n_34957));
NAND2X1 g140963(.A (n_26572), .B (n_8303), .Y (n_34955));
NAND2X1 g140964(.A (n_25756), .B (n_30013), .Y (n_34956));
AND2X1 g140965(.A (n_34959), .B (n_34960), .Y (n_34961));
INVX1 g140966(.A (n_34958), .Y (n_34959));
AOI21X1 g140967(.A0 (n_15261), .A1 (n_29132), .B0 (n_8614), .Y(n_34958));
INVX1 g140968(.A (n_9093), .Y (n_34960));
AND2X1 g140969(.A (n_28633), .B (n_29132), .Y (n_34963));
OAI21X1 g140977(.A0 (n_34971), .A1 (n_31343), .B0 (n_34974), .Y(n_34975));
AND2X1 g140978(.A (n_31073), .B (n_10402), .Y (n_34971));
AND2X1 g140979(.A (n_34972), .B (n_34973), .Y (n_34974));
OR2X1 g140980(.A (n_3466), .B (n_6389), .Y (n_34972));
NAND2X1 g140981(.A (n_1619), .B (P2_reg3[18] ), .Y (n_34973));
NAND2X2 g140982(.A (n_35436), .B (n_34978), .Y (n_34981));
NAND2X2 g140983(.A (n_34976), .B (n_34977), .Y (n_34978));
NAND2X1 g140984(.A (n_15399), .B (n_15400), .Y (n_34976));
NAND2X1 g140985(.A (n_7132), .B (n_3307), .Y (n_34977));
INVX1 g140986(.A (n_34979), .Y (n_35436));
NAND2X1 g140987(.A (n_8206), .B (n_7938), .Y (n_34979));
NAND2X1 g140989(.A (n_11941), .B (n_12659), .Y (n_34982));
NAND4X1 g140990(.A (n_34984), .B (n_34985), .C (n_34986), .D(n_11885), .Y (n_34987));
AND2X1 g140991(.A (n_11886), .B (n_34983), .Y (n_34984));
NAND4X1 g140992(.A (n_10278), .B (n_7746), .C (n_7399), .D (n_7389),.Y (n_34983));
INVX1 g140993(.A (n_11702), .Y (n_34985));
INVX1 g140994(.A (n_12055), .Y (n_34986));
NAND2X1 g140995(.A (n_11885), .B (n_11886), .Y (n_34989));
NOR2X1 g140996(.A (n_11702), .B (n_12055), .Y (n_35289));
NAND2X1 g140997(.A (n_34995), .B (n_34996), .Y (n_34997));
NAND2X1 g140998(.A (n_34992), .B (n_34998), .Y (n_34995));
INVX2 g140999(.A (n_34991), .Y (n_34992));
NAND2X2 g141000(.A (n_9695), .B (n_9206), .Y (n_34991));
NAND2X1 g141002(.A (n_15850), .B (n_16003), .Y (n_34993));
NAND2X1 g141003(.A (n_34617), .B (n_17246), .Y (n_34996));
INVX2 g141004(.A (n_34993), .Y (n_34998));
NOR2X1 g141005(.A (n_35002), .B (n_35003), .Y (n_35179));
INVX1 g141006(.A (n_35001), .Y (n_35002));
AND2X1 g141007(.A (n_34999), .B (n_35000), .Y (n_35001));
NAND2X1 g141008(.A (n_35245), .B (n_15945), .Y (n_34999));
NAND2X1 g141009(.A (n_15849), .B (n_16008), .Y (n_35000));
NAND2X1 g141010(.A (n_16761), .B (n_32362), .Y (n_35003));
NAND2X1 g141011(.A (n_35010), .B (n_35014), .Y (n_35015));
OAI21X1 g141012(.A0 (n_35005), .A1 (n_35006), .B0 (n_35009), .Y(n_35010));
NAND3X1 g141013(.A (n_34453), .B (n_32222), .C (n_32223), .Y(n_35005));
NAND3X1 g141014(.A (n_34258), .B (n_34259), .C (n_34455), .Y(n_35006));
CLKBUFX1 g141015(.A (n_35008), .Y (n_35009));
NOR2X1 g141016(.A (n_35007), .B (n_7620), .Y (n_35008));
AND2X1 g141017(.A (n_34698), .B (n_34699), .Y (n_35007));
NAND2X1 g141018(.A (n_35011), .B (n_35013), .Y (n_35014));
NOR2X1 g141019(.A (P2_reg2[28] ), .B (n_9310), .Y (n_35011));
INVX1 g141020(.A (n_35012), .Y (n_35013));
CLKBUFX1 g141021(.A (n_35007), .Y (n_35012));
NAND2X1 g141022(.A (n_35019), .B (n_35021), .Y (n_35022));
INVX1 g141023(.A (n_35018), .Y (n_35019));
AOI21X1 g141024(.A0 (n_31325), .A1 (n_35016), .B0 (n_35017), .Y(n_35018));
OR2X1 g141025(.A (n_31713), .B (n_8226), .Y (n_35016));
CLKBUFX1 g141026(.A (P1_n_449), .Y (n_35017));
AOI21X1 g141027(.A0 (n_6769), .A1 (n_3513), .B0 (n_35020), .Y(n_35021));
AND2X1 g141028(.A (n_35017), .B (P1_reg3[20] ), .Y (n_35020));
INVX1 g141029(.A (n_35017), .Y (n_35023));
INVX1 g141030(.A (P1_n_449), .Y (n_35024));
NAND2X1 g141041(.A (n_35038), .B (n_35039), .Y (n_35040));
NAND2X1 g141042(.A (n_35036), .B (n_35037), .Y (n_35038));
INVX1 g141043(.A (n_35035), .Y (n_35036));
NAND2X1 g141044(.A (n_32902), .B (n_32903), .Y (n_35035));
AND2X1 g141045(.A (n_17847), .B (n_18091), .Y (n_35037));
NAND2X1 g141046(.A (n_24521), .B (n_35041), .Y (n_35039));
INVX1 g141047(.A (n_35037), .Y (n_35041));
NAND2X1 g141048(.A (n_35045), .B (n_35049), .Y (n_35050));
NAND2X1 g141049(.A (n_35042), .B (n_35044), .Y (n_35045));
NAND2X2 g141050(.A (n_29187), .B (n_29667), .Y (n_35042));
INVX1 g141051(.A (n_35043), .Y (n_35044));
NAND3X1 g141052(.A (n_7993), .B (n_6441), .C (n_30897), .Y (n_35043));
AOI21X1 g141053(.A0 (n_32851), .A1 (n_28013), .B0 (n_35048), .Y(n_35049));
NAND2X1 g141054(.A (n_35046), .B (n_35047), .Y (n_35048));
NAND3X1 g141055(.A (n_8946), .B (n_7760), .C (n_7761), .Y (n_35046));
NAND2X1 g141056(.A (n_20218), .B (n_10546), .Y (n_35047));
NAND2X1 g141057(.A (n_35056), .B (n_35057), .Y (n_35058));
NAND2X1 g141058(.A (n_35054), .B (n_35055), .Y (n_35056));
BUFX3 g141059(.A (n_35053), .Y (n_35054));
INVX2 g141060(.A (n_35052), .Y (n_35053));
INVX2 g141061(.A (n_35051), .Y (n_35052));
NOR2X1 g141062(.A (n_34982), .B (n_34987), .Y (n_35051));
MX2X1 g141063(.A (n_17781), .B (n_21390), .S0 (n_25827), .Y(n_35055));
NAND2X1 g141064(.A (n_13299), .B (n_3184), .Y (n_35057));
NAND2X1 g141065(.A (n_35060), .B (n_35061), .Y (n_35062));
NAND3X1 g141066(.A (n_35059), .B (n_15996), .C (n_11797), .Y(n_35060));
NAND2X2 g141067(.A (n_15873), .B (n_15908), .Y (n_35059));
NAND2X2 g141068(.A (n_15997), .B (n_10309), .Y (n_35061));
AND2X1 g141069(.A (n_11797), .B (n_15996), .Y (n_35063));
MX2X1 g141079(.A (n_20776), .B (n_20775), .S0 (n_24388), .Y(n_35151));
MX2X1 g111095_dup(.A (n_20776), .B (n_20775), .S0 (n_24388), .Y(n_35152));
NOR2X1 g141080(.A (n_7066), .B (n_32834), .Y (n_35153));
NOR2X1 g129573_dup(.A (n_7066), .B (n_32834), .Y (n_35154));
NAND2X1 g141081(.A (n_35082), .B (n_5161), .Y (n_35155));
NAND2X1 g131148_dup(.A (n_35082), .B (n_5161), .Y (n_35156));
AND2X1 g141082(.A (n_35301), .B (n_4688), .Y (n_35157));
AND2X1 g131194_dup(.A (n_35302), .B (n_4688), .Y (n_35158));
OR2X1 g141083(.A (n_33353), .B (n_33358), .Y (n_35159));
OR2X1 g139461_dup(.A (n_33353), .B (n_33358), .Y (n_35160));
NAND2X1 g141084(.A (n_35946), .B (n_32289), .Y (n_35161));
NAND2X1 g130291_dup(.A (n_35947), .B (n_32289), .Y (n_35162));
MX2X1 g141085(.A (n_20266), .B (n_22511), .S0 (n_24329), .Y(n_35163));
MX2X1 g111094_dup(.A (n_20266), .B (n_22511), .S0 (n_24329), .Y(n_35164));
NAND3X1 g141086(.A (n_32343), .B (n_7543), .C (n_32245), .Y(n_35165));
NAND3X1 g124880_dup(.A (n_32343), .B (n_7543), .C (n_32245), .Y(n_35166));
INVX1 g141087(.A (n_35168), .Y (n_35167));
INVX1 g141088(.A (n_33168), .Y (n_35168));
INVX1 g141090(.A (n_35173), .Y (n_35171));
CLKBUFX1 g141092(.A (n_35174), .Y (n_35173));
CLKBUFX1 g141093(.A (n_35175), .Y (n_35174));
INVX1 g141094(.A (n_35304), .Y (n_35176));
INVX1 g141096(.A (n_35188), .Y (n_35180));
CLKBUFX1 g141109(.A (n_35195), .Y (n_35188));
INVX1 g141111(.A (n_35198), .Y (n_35196));
CLKBUFX1 g141112(.A (n_35198), .Y (n_35197));
INVX1 g141113(.A (n_35201), .Y (n_35199));
INVX1 g141115(.A (n_35203), .Y (n_35202));
CLKBUFX1 g141116(.A (n_35205), .Y (n_35203));
INVX1 g141117(.A (n_35205), .Y (n_35446));
INVX2 g141118(.A (n_35215), .Y (n_35205));
INVX2 g141119(.A (n_35208), .Y (n_35206));
CLKBUFX1 g141124(.A (n_35208), .Y (n_35212));
CLKBUFX1 g141125(.A (n_35214), .Y (n_35208));
CLKBUFX2 g141126(.A (n_35215), .Y (n_35214));
INVX1 g141127(.A (n_35217), .Y (n_35216));
INVX1 g141128(.A (n_19712), .Y (n_35217));
INVX1 g141129(.A (n_35221), .Y (n_35218));
INVX1 g141132(.A (n_35224), .Y (n_35223));
CLKBUFX1 g141133(.A (n_35225), .Y (n_35224));
INVX2 g141134(.A (n_33920), .Y (n_35225));
CLKBUFX1 g141137(.A (n_35231), .Y (n_35230));
INVX2 g141149(.A (n_35245), .Y (n_35244));
INVX2 g141150(.A (n_9738), .Y (n_35245));
INVX1 g141151(.A (n_35248), .Y (n_35247));
NAND3X1 g141152(.A (n_32054), .B (n_32055), .C (n_35659), .Y(n_35301));
NAND3X1 g131323_dup(.A (n_32054), .B (n_32055), .C (n_35660), .Y(n_35302));
NOR2X1 g141153(.A (n_18038), .B (n_33031), .Y (n_35303));
NOR2X1 g118240_dup(.A (n_18038), .B (n_33031), .Y (n_35304));
NAND2X1 g141154(.A (n_21116), .B (n_19439), .Y (n_35305));
NAND2X1 g114156_dup(.A (n_21116), .B (n_19439), .Y (n_35306));
NAND2X1 g141155(.A (n_29557), .B (n_29690), .Y (n_35307));
NAND2X1 g107502_dup(.A (n_29557), .B (n_29690), .Y (n_35308));
INVX1 g141156(.A (n_35310), .Y (n_35309));
INVX2 g141157(.A (n_35313), .Y (n_35311));
CLKBUFX3 g141159(.A (n_33963), .Y (n_35313));
INVX1 g141160(.A (n_35321), .Y (n_35314));
INVX1 g141161(.A (n_35318), .Y (n_35315));
CLKBUFX1 g141165(.A (n_35321), .Y (n_35318));
CLKBUFX2 g141167(.A (n_33963), .Y (n_35321));
MX2X1 g141169(.A (n_6378), .B (n_6342), .S0 (n_6286), .Y (n_35339));
MX2X1 g130157_dup(.A (n_6378), .B (n_6342), .S0 (n_6286), .Y(n_35340));
MX2X1 g141170(.A (n_34095), .B (n_34094), .S0 (n_34101), .Y(n_35341));
MX2X1 g140144_dup(.A (n_34095), .B (n_34094), .S0 (n_34101), .Y(n_35342));
NAND2X1 g141171(.A (n_7756), .B (n_7952), .Y (n_35343));
NAND2X1 g128067_dup(.A (n_7756), .B (n_7952), .Y (n_35344));
NOR2X1 g141172(.A (n_17058), .B (n_17545), .Y (n_35345));
NOR2X1 g116529_dup(.A (n_17545), .B (n_17058), .Y (n_35346));
MX2X1 g141173(.A (n_6255), .B (n_6256), .S0 (n_32406), .Y (n_35347));
MX2X1 g130646_dup(.A (n_6255), .B (n_6256), .S0 (n_32406), .Y(n_35348));
INVX1 g141174(.A (n_35350), .Y (n_35349));
CLKBUFX1 g141175(.A (n_35351), .Y (n_35350));
CLKBUFX2 g141176(.A (n_35352), .Y (n_35351));
CLKBUFX1 g141177(.A (n_35355), .Y (n_35353));
INVX1 g141178(.A (n_35355), .Y (n_35354));
INVX1 g141179(.A (n_35357), .Y (n_35356));
INVX2 g141181(.A (n_35364), .Y (n_35360));
INVX1 g141182(.A (n_35364), .Y (n_35361));
CLKBUFX3 g141185(.A (n_35366), .Y (n_35364));
INVX1 g141186(.A (n_35366), .Y (n_35882));
INVX2 g141187(.A (n_32976), .Y (n_35366));
INVX1 g141189(.A (n_35380), .Y (n_35368));
INVX2 g141201(.A (n_3644), .Y (n_35380));
NAND4X1 g141202(.A (n_7796), .B (n_7976), .C (n_8996), .D (n_7524),.Y (n_35384));
NAND4X1 g125788_dup(.A (n_7796), .B (n_7976), .C (n_8996), .D(n_7524), .Y (n_35385));
NOR2X1 g141203(.A (n_33242), .B (n_35661), .Y (n_35386));
NOR2X1 g139358_dup(.A (n_33242), .B (n_35662), .Y (n_35387));
NAND2X1 g141204(.A (n_23072), .B (n_22297), .Y (n_35388));
NAND2X1 g112730_dup(.A (n_23072), .B (n_22297), .Y (n_35389));
NAND2X1 g141205(.A (n_32215), .B (n_32216), .Y (n_35390));
NAND2X1 g132958_dup(.A (n_32215), .B (n_32216), .Y (n_35391));
NOR2X1 g141206(.A (n_6188), .B (n_34574), .Y (n_35392));
NOR2X1 g130880_dup(.A (n_6188), .B (n_34574), .Y (n_35393));
AOI22X1 g141207(.A0 (n_8124), .A1 (n_12803), .B0 (n_13071), .B1(n_13106), .Y (n_35394));
AOI22X1 g123127_dup(.A0 (n_8124), .A1 (n_12803), .B0 (n_13071), .B1(n_13106), .Y (n_35395));
NAND2X1 g141208(.A (n_35903), .B (n_33853), .Y (n_35396));
NAND2X1 g139938_dup(.A (n_33853), .B (n_35902), .Y (n_35397));
OR2X1 g141209(.A (n_35313), .B (n_33964), .Y (n_35398));
OR2X1 g140024_dup(.A (n_35313), .B (n_33964), .Y (n_35399));
NAND2X1 g141210(.A (n_35117), .B (n_35118), .Y (n_35400));
NAND2X1 g132198_dup(.A (n_35117), .B (n_35118), .Y (n_35401));
NAND2X1 g141211(.A (n_20034), .B (n_21062), .Y (n_35402));
NAND2X1 g114269_dup(.A (n_20034), .B (n_21062), .Y (n_35403));
INVX1 g141212(.A (n_35407), .Y (n_35404));
INVX1 g141215(.A (n_9958), .Y (n_35407));
NAND2X1 g141216(.A (n_35274), .B (n_35275), .Y (n_32406));
NAND2X1 g131112_dup(.A (n_35275), .B (n_35274), .Y (n_35452));
NAND2X1 g141217(.A (n_7287), .B (n_3263), .Y (n_35453));
NAND2X1 g129271_dup(.A (n_7287), .B (n_3263), .Y (n_35454));
NAND2X1 g141218(.A (n_24082), .B (n_25214), .Y (n_35455));
NAND2X1 g109005_dup(.A (n_24082), .B (n_25214), .Y (n_35456));
CLKBUFX3 g141219(.A (n_35467), .Y (n_35457));
INVX1 g141220(.A (n_35462), .Y (n_35459));
INVX1 g141222(.A (n_35463), .Y (n_35462));
CLKBUFX3 g141223(.A (n_35463), .Y (n_35464));
CLKBUFX3 g141224(.A (n_35466), .Y (n_35463));
INVX2 g141225(.A (n_35467), .Y (n_35466));
INVX1 g141226(.A (n_35473), .Y (n_35468));
INVX2 g141234(.A (n_35478), .Y (n_35473));
INVX2 g141235(.A (n_35467), .Y (n_35478));
CLKBUFX3 g141237(.A (n_35467), .Y (n_35479));
CLKBUFX3 g141238(.A (n_35524), .Y (n_35467));
INVX2 g141244(.A (n_35524), .Y (n_35485));
INVX2 g141245(.A (n_35500), .Y (n_35494));
INVX2 g141252(.A (n_35523), .Y (n_35500));
INVX2 g141254(.A (n_35508), .Y (n_35505));
CLKBUFX1 g141256(.A (n_35519), .Y (n_35508));
INVX1 g141259(.A (n_35515), .Y (n_35514));
CLKBUFX1 g141260(.A (n_35519), .Y (n_35515));
INVX4 g141263(.A (n_35519), .Y (n_35520));
INVX4 g141265(.A (n_35523), .Y (n_35519));
INVX2 g141266(.A (n_35524), .Y (n_35523));
INVX2 g141267(.A (n_35606), .Y (n_35524));
INVX2 g141271(.A (n_35528), .Y (n_35529));
INVX4 g141272(.A (n_35532), .Y (n_35528));
INVX2 g141273(.A (n_35537), .Y (n_35532));
INVX2 g141277(.A (n_35540), .Y (n_35538));
INVX8 g141279(.A (n_35570), .Y (n_35540));
INVX1 g141283(.A (n_35540), .Y (n_35546));
INVX4 g141293(.A (n_35540), .Y (n_35555));
INVX4 g141305(.A (n_35537), .Y (n_35570));
INVX2 g141306(.A (n_35606), .Y (n_35537));
INVX1 g141308(.A (n_35576), .Y (n_35572));
INVX2 g141312(.A (n_35583), .Y (n_35576));
INVX1 g141314(.A (n_35578), .Y (n_35580));
INVX2 g141315(.A (n_35583), .Y (n_35578));
CLKBUFX1 g141320(.A (n_35583), .Y (n_35590));
BUFX3 g141321(.A (n_35606), .Y (n_35583));
CLKBUFX3 g141322(.A (n_35600), .Y (n_35596));
CLKBUFX1 g141325(.A (n_35600), .Y (n_35602));
BUFX3 g141326(.A (n_35606), .Y (n_35600));
INVX2 g141327(.A (n_33281), .Y (n_35606));
NOR2X1 g141328(.A (n_34231), .B (n_34232), .Y (n_35620));
NOR2X1 g140264_dup(.A (n_34231), .B (n_34232), .Y (n_35621));
NAND2X1 g141329(.A (n_15707), .B (n_8432), .Y (n_35622));
NAND2X1 g120176_dup(.A (n_15707), .B (n_8432), .Y (n_35623));
NAND2X1 g141330(.A (n_34359), .B (n_34592), .Y (n_35624));
NAND2X1 g140390_dup(.A (n_34359), .B (n_34592), .Y (n_35625));
INVX1 g141331(.A (n_35630), .Y (n_35626));
INVX1 g141332(.A (n_35630), .Y (n_35627));
INVX1 g141334(.A (n_35630), .Y (n_35629));
NAND2X1 g141335(.A (n_32196), .B (n_32197), .Y (n_35649));
NAND2X1 g110248_dup(.A (n_32196), .B (n_32197), .Y (n_35650));
NAND2X1 g141336(.A (n_6258), .B (n_6218), .Y (n_35651));
NAND2X1 g130256_dup(.A (n_6218), .B (n_6258), .Y (n_35652));
MX2X1 g141337(.A (n_5161), .B (n_6069), .S0 (n_5995), .Y (n_35653));
MX2X1 g130963_dup(.A (n_5161), .B (n_6069), .S0 (n_5995), .Y(n_35952));
MX2X1 g141338(.A (n_6256), .B (n_6255), .S0 (n_32406), .Y (n_35655));
MX2X1 g130647_dup(.A (n_6256), .B (n_6255), .S0 (n_32406), .Y(n_35656));
NAND2X1 g141339(.A (n_34915), .B (n_34921), .Y (n_35657));
NAND2X1 g140921_dup(.A (n_34915), .B (n_34921), .Y (n_35658));
NOR2X1 g141340(.A (n_33584), .B (n_5200), .Y (n_35659));
NOR2X1 g131525_dup(.A (n_33584), .B (n_5200), .Y (n_35660));
NOR2X1 g141341(.A (n_33243), .B (n_33247), .Y (n_35661));
NOR2X1 g139360_dup(.A (n_33243), .B (n_33247), .Y (n_35662));
NAND2X1 g141342(.A (n_7809), .B (n_8200), .Y (n_35663));
NAND2X2 g128176_dup(.A (n_7809), .B (n_8200), .Y (n_9746));
NOR2X1 g141343(.A (n_16674), .B (n_17573), .Y (n_35665));
NOR2X1 g115865_dup(.A (n_16674), .B (n_17573), .Y (n_35666));
NAND2X1 g141344(.A (n_35143), .B (n_35144), .Y (n_35667));
NAND2X1 g129505_dup(.A (n_35143), .B (n_35144), .Y (n_35668));
INVX1 g141345(.A (n_35672), .Y (n_35670));
CLKBUFX1 g141346(.A (n_35672), .Y (n_35671));
INVX2 g141347(.A (n_16669), .Y (n_35672));
INVX1 g141349(.A (n_35675), .Y (n_35674));
INVX2 g141353(.A (n_35686), .Y (n_35679));
CLKBUFX3 g141360(.A (n_35675), .Y (n_35686));
INVX2 g141361(.A (n_15801), .Y (n_35675));
CLKBUFX1 g141362(.A (n_35689), .Y (n_35688));
OR2X1 g141363(.A (n_17218), .B (n_18412), .Y (n_35707));
OR2X1 g118537_dup(.A (n_17218), .B (n_18412), .Y (n_35708));
NAND2X2 g141364(.A (n_6214), .B (n_35386), .Y (n_35709));
NAND2X1 g130887_dup(.A (n_6214), .B (n_35386), .Y (n_35710));
NAND2X1 g141365(.A (n_33559), .B (n_33560), .Y (n_35711));
NAND2X1 g139534_dup(.A (n_33559), .B (n_33560), .Y (n_35712));
NAND2X1 g141366(.A (n_35338), .B (n_35337), .Y (n_35713));
NAND2X1 g127647_dup(.A (n_35338), .B (n_35337), .Y (n_35714));
NAND2X1 g141367(.A (n_17542), .B (n_16255), .Y (n_35715));
NAND2X1 g116171_dup(.A (n_17542), .B (n_16255), .Y (n_35716));
OAI21X1 g141368(.A0 (n_18482), .A1 (n_18684), .B0 (n_19733), .Y(n_35717));
OAI21X1 g116078_dup(.A0 (n_18482), .A1 (n_18684), .B0 (n_19733), .Y(n_35718));
INVX8 g141379(.A (n_35719), .Y (n_35736));
BUFX3 g141383(.A (n_35818), .Y (n_35719));
INVX4 g141386(.A (n_35771), .Y (n_35744));
INVX1 g141397(.A (n_35766), .Y (n_35761));
INVX4 g141399(.A (n_35767), .Y (n_35766));
CLKBUFX3 g141401(.A (n_35771), .Y (n_35768));
INVX4 g141403(.A (n_35767), .Y (n_35771));
INVX4 g141404(.A (n_35818), .Y (n_35767));
INVX1 g141405(.A (n_35775), .Y (n_35776));
INVX4 g141414(.A (n_35775), .Y (n_35790));
INVX1 g141415(.A (n_35775), .Y (n_35794));
BUFX3 g141420(.A (n_35818), .Y (n_35775));
INVX4 g141432(.A (n_35813), .Y (n_35816));
CLKBUFX1 g141433(.A (n_35818), .Y (n_35813));
INVX4 g141439(.A (n_35822), .Y (n_35824));
INVX4 g141440(.A (n_35829), .Y (n_35822));
CLKBUFX1 g141442(.A (n_35829), .Y (n_35830));
CLKBUFX3 g141443(.A (n_35818), .Y (n_35829));
INVX2 g141447(.A (n_35767), .Y (n_35834));
INVX1 g141449(.A (n_35840), .Y (n_35842));
INVX2 g141450(.A (n_35767), .Y (n_35840));
INVX2 g141452(.A (n_35767), .Y (n_35844));
CLKBUFX3 g141454(.A (n_34216), .Y (n_35818));
CLKBUFX1 g141455(.A (n_35849), .Y (n_35850));
INVX2 g141464(.A (n_35861), .Y (n_35860));
CLKBUFX3 g141465(.A (n_35864), .Y (n_35861));
INVX1 g141466(.A (n_35864), .Y (n_35863));
INVX4 g141467(.A (n_34104), .Y (n_35864));
INVX1 g141468(.A (n_35867), .Y (n_35865));
CLKBUFX1 g141470(.A (n_35868), .Y (n_35867));
INVX1 g141471(.A (P2_IR[9] ), .Y (n_35868));
INVX1 g141475(.A (n_35896), .Y (n_35895));
INVX1 g141476(.A (n_35903), .Y (n_35901));
CLKBUFX1 g141477(.A (n_35903), .Y (n_35902));
INVX1 g141478(.A (n_33854), .Y (n_35903));
NAND2X1 g141479(.A (n_35205), .B (n_34163), .Y (n_35912));
NAND2X1 g140194_dup(.A (n_35205), .B (n_34163), .Y (n_35913));
INVX1 g141480(.A (n_35915), .Y (n_35914));
NAND2X1 g141482(.A (n_20036), .B (n_18865), .Y (n_35934));
NAND2X1 g114412_dup(.A (n_20036), .B (n_18865), .Y (n_35935));
AND2X1 g141483(.A (n_35446), .B (n_16203), .Y (n_35936));
AND2X1 g140155_dup(.A (n_35446), .B (n_16203), .Y (n_35937));
NAND2X1 g141484(.A (n_32293), .B (n_19816), .Y (n_35938));
NAND2X1 g139875_dup(.A (n_32293), .B (n_19816), .Y (n_35939));
CLKBUFX1 g141485(.A (n_6800), .Y (n_35940));
CLKBUFX1 g129597_dup(.A (n_6800), .Y (n_35941));
NOR2X1 g141486(.A (n_16569), .B (n_16071), .Y (n_35942));
NOR2X1 g118236_dup(.A (n_16569), .B (n_16071), .Y (n_35943));
NOR2X1 g141487(.A (n_11501), .B (n_13055), .Y (n_35944));
NOR2X1 g123119_dup(.A (n_11501), .B (n_13055), .Y (n_35945));
NAND2X1 g141488(.A (n_32889), .B (n_33583), .Y (n_35946));
NAND2X1 g130595_dup(.A (n_32889), .B (n_33583), .Y (n_35947));
CLKBUFX1 g141490(.A (n_35951), .Y (n_35950));
endmodule
