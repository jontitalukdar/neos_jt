module gcm_aes_v0 ( clk, rst, dii_data, dii_data_vld, dii_data_type,dii_data_not_ready, dii_last_word, dii_data_size, cii_ctl_vld,cii_IV_vld, cii_K, Out_data, Out_vld, Out_data_size, Out_last_word,Tag_vld );
input [127:0] dii_data;
input [3:0] dii_data_size;
input [127:0] cii_K;
output [127:0] Out_data;
output [3:0] Out_data_size;
input clk, rst, dii_data_vld, dii_data_type, dii_last_word, cii_ctl_vld,cii_IV_vld;
output dii_data_not_ready, Out_vld, Out_last_word, Tag_vld;
wire   aes_done, aes_kld, N2027, N2028, N2029, N2030, N2031, N2032, N2033,N2034, N2035, N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043,N2044, N2045, N2046, N2047, N2048, N2049, N2050, N2051, N2052, N2053,N2054, N2055, N2056, N2057, N2058, N2059, N2060, N2061, N2062, N2063,N2064, N2065, N2066, N2067, N2068, N2069, N2070, N2071, N2072, N2073,N2074, N2075, N2076, N2077, N2078, N2079, N2080, N2081, N2082, N2083,N2084, N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092, N2093,N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102, N2103,N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112, N2113,N2114, N2115, N2116, N2117, N2118, N2119, N2120, N2121, N2122, N2123,N2124, N2125, N2126, N2127, N2128, N2129, N2130, N2131, N2132, N2133,N2134, N2135, N2136, N2137, N2138, N2139, N2140, N2141, N2142, N2143,N2144, N2145, N2146, N2147, N2148, N2149, N2150, N2151, N2152, N2153,N2154, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357,N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367,N2368, N2369, N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377,N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387,N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397,N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407,N2408, N2409, N2410, N2411, N2412, N2479, N2480, N2481, N2482, N2483,N2484, N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493,N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503,N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513,N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523,N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533,N2534, N2535, N2536, N2537, N2538, N2539, N2540, N2541, N2542, N2815,N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825,N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835,N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845,N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855,N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863, N2864, N2865,N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875,N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, N2885,N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895,N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905,N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915,N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925,N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935,N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945,N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955,N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965,N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975,N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985,N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995,N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005,N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015,N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025,N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035,N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045,N3046, N3047, N3048, N3049, N3050, N3051, N3052, N3053, N3054, N3055,N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065,N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075,N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085,N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095,N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105,N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115,N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123, N3124, N3125,N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133, N3134, N3135,N3136, N3137, N3138, N3139, N3140, N3141, N3142, N3143, N3144, N3145,N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155,N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165,N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, N3175,N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, N3185,N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195,N3196, N3197, N3198, n5326, n5327, n5328, n5329, n5330, n5331, n5332,n5333, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5358,n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5374, n5375, n5376,n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,n5437, n5438, n5439, n5440, n5441, n5442, n5444, n5445, n5446, n5447,n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,n5568, n5569, n5570, n5571, n5574, n5575, n5576, n5577, n5578, n5579,n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,n6290, n6291, n6292, n6293, n6294, n6295, n6850, n6859, n11921,n11922, n11923, n11924, n11926, n11927, n11928, n11929, n11930,n11931, n11935, n11936, n11937, n11939, n11940, n11941, n11942,n11943, n11944, n11946, n11947, n11948, n11949, n11950, n11953,n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11970,n11971, n11973, n11976, n11979, n11980, n11981, n11982, n11983,n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,n12496, n12497, n12498, n12499, n12500, n12501, n12502, n13019,n13020, n13023, n13024, n13025, n13026, n13027, n13028, n13029,n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,n13278, n13279, n13280, n13281, n13284, n13285, n13286, n13287,n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,n13656, n13657, n13658, n13659, n13661, n13662, n13663, n13664,n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,n14025, n14026, n14155, n14157, n14158, n14159, n14160, n14161,n14162, n14163, n14164, n14166, n14167, n14168, n14169, n14170,n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,n14387, n14388, n14389, n14391, n14393, n14394, n14395, n14396,n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14773,n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,n14942, n14943, n14944, n14945, n14946, n14947, n14949, n14950,n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15504,n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,n15529, n15530, n15532, n15533, n15534, n15535, n15536, n15537,n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,n15546, n15547, n15548, n15549, n15550, n15551, n15553, n15554,n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,n15571, n15572, n15574, n15575, n15576, n15577, n15578, n15579,n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,n15588, n15589, n15590, n15591, n15592, n15593, n15595, n15596,n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,n16437, n16438, n16439, n16440, n16443, n16444, n16445, n16446,n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,n16455, n16458, n16459, n16460, n16461, n16462, n16463, n16464,n16465, n16466, n16467, n16468, n16471, n16472, n16473, n16474,n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16484,n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,n16493, n16494, n16497, n16498, n16499, n16500, n16501, n16502,n16503, n16504, n16505, n16506, n16507, n16510, n16511, n16512,n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,n16531, n16532, n16533, n16536, n16537, n16538, n16539, n16540,n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,n16549, n16550, n16551, n16553, n16554, n16555, n16556, n16558,n16559, n16560, n16561, n16563, n16564, n16565, n16566, n16568,n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,n16833, n16834, n16835, n16836, n16837, n16838, n16839, n17024,n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17041,n17043, n17045, n17047, n17049, n17051, n17053, n17055, n17057,n17059, n17061, n17063, n17065, n17067, n17069, n17071, n17073,n17075, n17077, n17079, n17081, n17083, n17085, n17087, n17089,n17091, n17093, n17095, n17097, n17099, n17101, n17103, n17105,n17107, n17109, n17111, n17113, n17115, n17117, n17119, n17121,n17123, n17125, n17127, n17129, n17131, n17133, n17135, n17137,n17139, n17141, n17143, n17145, n17147, n17149, n17151, n17153,n17155, n17157, n17159, n17161, n17163, n17165, n17167, n17169,n17171, n17173, n17175, n17177, n17179, n17181, n17183, n17185,n17187, n17189, n17191, n17193, n17195, n17197, n17199, n17201,n17203, n17205, n17207, n17209, n17211, n17213, n17215, n17217,n17219, n17221, n17223, n17225, n17227, n17229, n17231, n17233,n17235, n17237, n17239, n17241, n17243, n17245, n17247, n17249,n17251, n17253, n17255, n17257, n17259, n17261, n17263, n17264,n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,n19201, n19202, n19203, n19204, n19205, n19206, \GFM/n2699 ,\GFM/n26980 , \GFM/n2697 , \GFM/n2696 , \GFM/n2695 , \GFM/n26940 ,\GFM/n26930 , \GFM/n26921 , \GFM/n26910 , \GFM/n26900 , \GFM/n2689 ,\GFM/n2688 , \GFM/n26870 , \GFM/n26860 , \GFM/n2685 , \GFM/n26840 ,\GFM/n2683 , \GFM/n26820 , \GFM/n26810 , \GFM/n26801 , \GFM/n2679 ,\GFM/n2678 , \GFM/n26770 , \GFM/n26760 , \GFM/n2675 , \GFM/n26740 ,\GFM/n26730 , \GFM/n2672 , \GFM/n2671 , \GFM/n26700 , \GFM/n26690 ,\GFM/n2668 , \GFM/n26670 , \GFM/n2666 , \GFM/n2665 , \GFM/n2664 ,\GFM/n26630 , \GFM/n26620 , \GFM/n26611 , \GFM/n26600 , \GFM/n26590 ,\GFM/n2658 , \GFM/n2657 , \GFM/n26560 , \GFM/n26550 , \GFM/n2654 ,\GFM/n26530 , \GFM/n2652 , \GFM/n26510 , \GFM/n26500 , \GFM/n2649 ,\GFM/n2648 , \GFM/n2647 , \GFM/n26460 , \GFM/n26450 , \GFM/n2644 ,\GFM/n26430 , \GFM/n26420 , \GFM/n2641 , \GFM/n26401 , \GFM/n26390 ,\GFM/n26380 , \GFM/n2637 , \GFM/n26360 , \GFM/n2635 , \GFM/n2634 ,\GFM/n2633 , \GFM/n26320 , \GFM/n26310 , \GFM/n26301 , \GFM/n26290 ,\GFM/n26280 , \GFM/n2627 , \GFM/n2626 , \GFM/n26250 , \GFM/n26240 ,\GFM/n2623 , \GFM/n26220 , \GFM/n2621 , \GFM/n26200 , \GFM/n26190 ,\GFM/n2618 , \GFM/n2617 , \GFM/n2616 , \GFM/n26150 , \GFM/n26140 ,\GFM/n2613 , \GFM/n26120 , \GFM/n26110 , \GFM/n2610 , \GFM/n2609 ,\GFM/n26080 , \GFM/n26070 , \GFM/n2606 , \GFM/n26050 , \GFM/n2604 ,\GFM/n2603 , \GFM/n2602 , \GFM/n26010 , \GFM/n26000 , \GFM/n2599 ,\GFM/n25980 , \GFM/n25970 , \GFM/n2596 , \GFM/n2595 , \GFM/n25940 ,\GFM/n25930 , \GFM/n2592 , \GFM/n25910 , \GFM/n25901 , \GFM/n25890 ,\GFM/n25880 , \GFM/n2587 , \GFM/n2586 , \GFM/n2585 , \GFM/n25840 ,\GFM/n25830 , \GFM/n25821 , \GFM/n25810 , \GFM/n25800 , \GFM/n2579 ,\GFM/n2578 , \GFM/n25770 , \GFM/n25760 , \GFM/n2575 , \GFM/n25740 ,\GFM/n2573 , \GFM/n2572 , \GFM/n2571 , \GFM/n25700 , \GFM/n25690 ,\GFM/n2568 , \GFM/n25670 , \GFM/n25660 , \GFM/n2565 , \GFM/n2564 ,\GFM/n25630 , \GFM/n25620 , \GFM/n25611 , \GFM/n25600 , \GFM/n2559 ,\GFM/n25580 , \GFM/n25570 , \GFM/n2556 , \GFM/n2555 , \GFM/n2554 ,\GFM/n25530 , \GFM/n25520 , \GFM/n25511 , \GFM/n25500 , \GFM/n25490 ,\GFM/n2548 , \GFM/n2547 , \GFM/n25460 , \GFM/n25450 , \GFM/n2544 ,\GFM/n25430 , \GFM/n2542 , \GFM/n2541 , \GFM/n2540 , \GFM/n25390 ,\GFM/n25380 , \GFM/n2537 , \GFM/n25360 , \GFM/n25350 , \GFM/n2534 ,\GFM/n2533 , \GFM/n25320 , \GFM/n25310 , \GFM/n2530 , \GFM/n25290 ,\GFM/n2528 , \GFM/n25270 , \GFM/n25260 , \GFM/n2525 , \GFM/n2524 ,\GFM/n2523 , \GFM/n25220 , \GFM/n25210 , \GFM/n25201 , \GFM/n25190 ,\GFM/n25180 , \GFM/n2517 , \GFM/n2516 , \GFM/n25150 , \GFM/n25140 ,\GFM/n2513 , \GFM/n25120 , \GFM/n2511 , \GFM/n25101 , \GFM/n2509 ,\GFM/n25080 , \GFM/n25070 , \GFM/n2506 , \GFM/n25050 , \GFM/n25040 ,\GFM/n2503 , \GFM/n2502 , \GFM/n25010 , \GFM/n25000 , \GFM/n2499 ,\GFM/n24980 , \GFM/n2497 , \GFM/n24960 , \GFM/n24950 , \GFM/n2494 ,\GFM/n2493 , \GFM/n24921 , \GFM/n24910 , \GFM/n24900 , \GFM/n2489 ,\GFM/n24880 , \GFM/n24870 , \GFM/n2486 , \GFM/n2485 , \GFM/n24840 ,\GFM/n24830 , \GFM/n2482 , \GFM/n24810 , \GFM/n2480 , \GFM/n2479 ,\GFM/n2478 , \GFM/n24770 , \GFM/n24760 , \GFM/n2475 , \GFM/n24740 ,\GFM/n24730 , \GFM/n2472 , \GFM/n2471 , \GFM/n24700 , \GFM/n24690 ,\GFM/n2468 , \GFM/n24670 , \GFM/n2466 , \GFM/n24650 , \GFM/n24640 ,\GFM/n2463 , \GFM/n2462 , \GFM/n2461 , \GFM/n24600 , \GFM/n24590 ,\GFM/n2458 , \GFM/n24570 , \GFM/n24560 , \GFM/n2455 , \GFM/n2454 ,\GFM/n24530 , \GFM/n24520 , \GFM/n24511 , \GFM/n24500 , \GFM/n2449 ,\GFM/n2448 , \GFM/n2447 , \GFM/n24460 , \GFM/n24450 , \GFM/n2444 ,\GFM/n24430 , \GFM/n24420 , \GFM/n2441 , \GFM/n24401 , \GFM/n24390 ,\GFM/n24380 , \GFM/n2437 , \GFM/n24360 , \GFM/n2435 , \GFM/n24340 ,\GFM/n24330 , \GFM/n2432 , \GFM/n2431 , \GFM/n2430 , \GFM/n24290 ,\GFM/n24280 , \GFM/n2427 , \GFM/n24260 , \GFM/n24250 , \GFM/n2424 ,\GFM/n2423 , \GFM/n24220 , \GFM/n24210 , \GFM/n24201 , \GFM/n24190 ,\GFM/n2418 , \GFM/n2417 , \GFM/n2416 , \GFM/n24150 , \GFM/n24140 ,\GFM/n2413 , \GFM/n24120 , \GFM/n24110 , \GFM/n24101 , \GFM/n2409 ,\GFM/n24080 , \GFM/n24070 , \GFM/n2406 , \GFM/n24050 , \GFM/n2404 ,\GFM/n24030 , \GFM/n24020 , \GFM/n2401 , \GFM/n2400 , \GFM/n2399 ,\GFM/n23980 , \GFM/n23970 , \GFM/n2396 , \GFM/n23950 , \GFM/n23940 ,\GFM/n2393 , \GFM/n2392 , \GFM/n23910 , \GFM/n23900 , \GFM/n2389 ,\GFM/n23880 , \GFM/n2387 , \GFM/n21360 , \GFM/n21350 , \GFM/n2134 ,\GFM/n21330 , \GFM/n21320 , \GFM/n2131 , \GFM/n21301 , \GFM/n21290 ,\GFM/n21280 , \GFM/n2127 , \GFM/n21260 , \GFM/n2125 , \GFM/n21240 ,\GFM/n21230 , \GFM/n2122 , \GFM/n2121 , \GFM/n184 , \GFM/n18310 ,\GFM/n18210 , \GFM/n181 , \GFM/n18011 , \GFM/n17911 , \GFM/n178 ,\GFM/n177 , \GFM/n17611 , \GFM/n17511 , \GFM/n174 , \GFM/n17310 ,\GFM/n172 , \GFM/n17110 , \GFM/n17011 , \GFM/n2120 , \GFM/n21190 ,\GFM/n21180 , \GFM/n2117 , \GFM/n21160 , \GFM/n21150 , \GFM/n2114 ,\GFM/n2113 , \GFM/n21120 , \GFM/n21110 , \GFM/n21101 , \GFM/n21090 ,\GFM/n2108 , \GFM/n2107 , \GFM/n2106 , \GFM/n21050 , \GFM/n21040 ,\GFM/n2103 , \GFM/n21020 , \GFM/n21010 , \GFM/n21001 , \GFM/n2099 ,\GFM/n20980 , \GFM/n20970 , \GFM/n2096 , \GFM/n20950 , \GFM/n2094 ,\GFM/n20930 , \GFM/n20920 , \GFM/n2091 , \GFM/n2090 , \GFM/n2089 ,\GFM/n20880 , \GFM/n20870 , \GFM/n2086 , \GFM/n20850 , \GFM/n20840 ,\GFM/n2083 , \GFM/n2082 , \GFM/n20810 , \GFM/n20800 , \GFM/n2079 ,\GFM/n20780 , \GFM/n2077 , \GFM/n2076 , \GFM/n2075 , \GFM/n20740 ,\GFM/n20730 , \GFM/n20721 , \GFM/n20710 , \GFM/n20700 , \GFM/n2069 ,\GFM/n2068 , \GFM/n20670 , \GFM/n20660 , \GFM/n2065 , \GFM/n20640 ,\GFM/n2063 , \GFM/n20620 , \GFM/n20610 , \GFM/n20601 , \GFM/n2059 ,\GFM/n2058 , \GFM/n20570 , \GFM/n20560 , \GFM/n2055 , \GFM/n20540 ,\GFM/n20530 , \GFM/n2052 , \GFM/n2051 , \GFM/n20500 , \GFM/n20490 ,\GFM/n2048 , \GFM/n20470 , \GFM/n2046 , \GFM/n2045 , \GFM/n2044 ,\GFM/n20430 , \GFM/n20420 , \GFM/n20411 , \GFM/n20400 , \GFM/n20390 ,\GFM/n2038 , \GFM/n2037 , \GFM/n20360 , \GFM/n20350 , \GFM/n2034 ,\GFM/n20330 , \GFM/n2032 , \GFM/n20310 , \GFM/n20300 , \GFM/n2029 ,\GFM/n2028 , \GFM/n2027 , \GFM/n20260 , \GFM/n20250 , \GFM/n2024 ,\GFM/n20230 , \GFM/n20220 , \GFM/n2021 , \GFM/n20201 , \GFM/n20190 ,\GFM/n20180 , \GFM/n2017 , \GFM/n20160 , \GFM/n2015 , \GFM/n2014 ,\GFM/n2013 , \GFM/n20120 , \GFM/n20110 , \GFM/n20101 , \GFM/n20090 ,\GFM/n20080 , \GFM/n2007 , \GFM/n2006 , \GFM/n20050 , \GFM/n20040 ,\GFM/n2003 , \GFM/n20020 , \GFM/n2001 , \GFM/n20000 , \GFM/n19990 ,\GFM/n1998 , \GFM/n1997 , \GFM/n1996 , \GFM/n19950 , \GFM/n19940 ,\GFM/n1993 , \GFM/n19920 , \GFM/n19910 , \GFM/n1990 , \GFM/n1989 ,\GFM/n19880 , \GFM/n19870 , \GFM/n1986 , \GFM/n19850 , \GFM/n1984 ,\GFM/n1983 , \GFM/n1982 , \GFM/n19810 , \GFM/n19800 , \GFM/n1979 ,\GFM/n19780 , \GFM/n19770 , \GFM/n1976 , \GFM/n1975 , \GFM/n19740 ,\GFM/n19730 , \GFM/n1972 , \GFM/n19710 , \GFM/n19701 , \GFM/n19690 ,\GFM/n19680 , \GFM/n1967 , \GFM/n1966 , \GFM/n1965 , \GFM/n19640 ,\GFM/n19630 , \GFM/n19621 , \GFM/n19610 , \GFM/n19600 , \GFM/n1959 ,\GFM/n1958 , \GFM/n19570 , \GFM/n19560 , \GFM/n1955 , \GFM/n19540 ,\GFM/n1953 , \GFM/n1952 , \GFM/n1951 , \GFM/n19500 , \GFM/n19490 ,\GFM/n1948 , \GFM/n19470 , \GFM/n19460 , \GFM/n1945 , \GFM/n1944 ,\GFM/n19430 , \GFM/n19420 , \GFM/n19411 , \GFM/n19400 , \GFM/n1939 ,\GFM/n19380 , \GFM/n19370 , \GFM/n1936 , \GFM/n1935 , \GFM/n1934 ,\GFM/n19330 , \GFM/n19320 , \GFM/n19311 , \GFM/n19300 , \GFM/n19290 ,\GFM/n1928 , \GFM/n1927 , \GFM/n19260 , \GFM/n19250 , \GFM/n1924 ,\GFM/n19230 , \GFM/n1922 , \GFM/n1921 , \GFM/n1920 , \GFM/n19190 ,\GFM/n19180 , \GFM/n1917 , \GFM/n19160 , \GFM/n19150 , \GFM/n1914 ,\GFM/n1913 , \GFM/n19120 , \GFM/n19110 , \GFM/n1910 , \GFM/n19090 ,\GFM/n1908 , \GFM/n19070 , \GFM/n19060 , \GFM/n1905 , \GFM/n1904 ,\GFM/n1903 , \GFM/n19020 , \GFM/n19010 , \GFM/n19001 , \GFM/n18990 ,\GFM/n18980 , \GFM/n1897 , \GFM/n1896 , \GFM/n18950 , \GFM/n18940 ,\GFM/n1893 , \GFM/n18920 , \GFM/n1891 , \GFM/n18901 , \GFM/n1889 ,\GFM/n18880 , \GFM/n18870 , \GFM/n1886 , \GFM/n18850 , \GFM/n18840 ,\GFM/n1883 , \GFM/n1882 , \GFM/n18810 , \GFM/n18800 , \GFM/n1879 ,\GFM/n18780 , \GFM/n1877 , \GFM/n18760 , \GFM/n18750 , \GFM/n1874 ,\GFM/n1873 , \GFM/n18721 , \GFM/n18710 , \GFM/n18700 , \GFM/n1869 ,\GFM/n18680 , \GFM/n18670 , \GFM/n1866 , \GFM/n1865 , \GFM/n18640 ,\GFM/n18630 , \GFM/n1862 , \GFM/n18610 , \GFM/n1860 , \GFM/n1859 ,\GFM/n1858 , \GFM/n18570 , \GFM/n18560 , \GFM/n1855 , \GFM/n18540 ,\GFM/n18530 , \GFM/n1852 , \GFM/n1851 , \GFM/n18500 , \GFM/n18490 ,\GFM/n1848 , \GFM/n18470 , \GFM/n1846 , \GFM/n18450 , \GFM/n18440 ,\GFM/n1843 , \GFM/n1842 , \GFM/n1841 , \GFM/n18400 , \GFM/n18390 ,\GFM/n1838 , \GFM/n18370 , \GFM/n18360 , \GFM/n1835 , \GFM/n1834 ,\GFM/n18330 , \GFM/n18320 , \GFM/n1831 , \GFM/n18300 , \GFM/n1829 ,\GFM/n1828 , \GFM/n1827 , \GFM/n18260 , \GFM/n18250 , \GFM/n1824 ,\GFM/n18230 , \GFM/n18220 , \GFM/n1821 , \GFM/n1820 , \GFM/n18190 ,\GFM/n18180 , \GFM/n1817 , \GFM/n18160 , \GFM/n1815 , \GFM/n18140 ,\GFM/n18130 , \GFM/n1812 , \GFM/n1811 , \GFM/n1810 , \GFM/n18090 ,\GFM/n18080 , \GFM/n1807 , \GFM/n18060 , \GFM/n18050 , \GFM/n1804 ,\GFM/n1803 , \GFM/n18020 , \GFM/n18010 , \GFM/n1800 , \GFM/n17990 ,\GFM/n1798 , \GFM/n1797 , \GFM/n1796 , \GFM/n17950 , \GFM/n17940 ,\GFM/n1793 , \GFM/n17920 , \GFM/n17910 , \GFM/n1790 , \GFM/n1789 ,\GFM/n17880 , \GFM/n17870 , \GFM/n1786 , \GFM/n17850 , \GFM/n1784 ,\GFM/n17830 , \GFM/n17820 , \GFM/n1781 , \GFM/n1780 , \GFM/n1779 ,\GFM/n17780 , \GFM/n17770 , \GFM/n1776 , \GFM/n17750 , \GFM/n17740 ,\GFM/n1773 , \GFM/n1772 , \GFM/n17710 , \GFM/n17700 , \GFM/n1769 ,\GFM/n17680 , \GFM/n1767 , \GFM/n1766 , \GFM/n1765 , \GFM/n17640 ,\GFM/n17630 , \GFM/n1762 , \GFM/n17610 , \GFM/n17600 , \GFM/n1759 ,\GFM/n1758 , \GFM/n17570 , \GFM/n17560 , \GFM/n1755 , \GFM/n17540 ,\GFM/n1753 , \GFM/n17520 , \GFM/n17510 , \GFM/n1750 , \GFM/n1749 ,\GFM/n1748 , \GFM/n17470 , \GFM/n17460 , \GFM/n1745 , \GFM/n17440 ,\GFM/n17430 , \GFM/n1742 , \GFM/n1741 , \GFM/n17400 , \GFM/n17390 ,\GFM/n1738 , \GFM/n17370 , \GFM/n1736 , \GFM/n1735 , \GFM/n1734 ,\GFM/n17330 , \GFM/n17320 , \GFM/n1731 , \GFM/n17300 , \GFM/n17290 ,\GFM/n1728 , \GFM/n1727 , \GFM/n17260 , \GFM/n17250 , \GFM/n1724 ,\GFM/n17230 , \GFM/n1722 , \GFM/n17210 , \GFM/n17200 , \GFM/n1719 ,\GFM/n1718 , \GFM/n1717 , \GFM/n17160 , \GFM/n17150 , \GFM/n1714 ,\GFM/n17130 , \GFM/n17120 , \GFM/n1711 , \GFM/n1710 , \GFM/n17090 ,\GFM/n17080 , \GFM/n1707 , \GFM/n17060 , \GFM/n1705 , \GFM/n1704 ,\GFM/n1703 , \GFM/n17020 , \GFM/n17010 , \GFM/n1700 , \GFM/n16990 ,\GFM/n16980 , \GFM/n1697 , \GFM/n1696 , \GFM/n16950 , \GFM/n16940 ,\GFM/n1693 , \GFM/n16920 , \GFM/n1691 , \GFM/n16900 , \GFM/n16890 ,\GFM/n1688 , \GFM/n1687 , \GFM/n1686 , \GFM/n16850 , \GFM/n16840 ,\GFM/n1683 , \GFM/n16820 , \GFM/n16810 , \GFM/n1680 , \GFM/n1679 ,\GFM/n16780 , \GFM/n16770 , \GFM/n1676 , \GFM/n16750 , \GFM/n1674 ,\GFM/n1673 , \GFM/n1672 , \GFM/n16710 , \GFM/n16700 , \GFM/n1669 ,\GFM/n16680 , \GFM/n16670 , \GFM/n1666 , \GFM/n1665 , \GFM/n16640 ,\GFM/n16630 , \GFM/n1662 , \GFM/n16610 , \GFM/n1660 , \GFM/n16590 ,\GFM/n16580 , \GFM/n1657 , \GFM/n1656 , \GFM/n1655 , \GFM/n16540 ,\GFM/n16530 , \GFM/n1652 , \GFM/n16510 , \GFM/n16500 , \GFM/n1649 ,\GFM/n1648 , \GFM/n16470 , \GFM/n16460 , \GFM/n1645 , \GFM/n16440 ,\GFM/n1643 , \GFM/n1642 , \GFM/n1641 , \GFM/n16400 , \GFM/n16390 ,\GFM/n1638 , \GFM/n16370 , \GFM/n16360 , \GFM/n1635 , \GFM/n1634 ,\GFM/n16330 , \GFM/n16320 , \GFM/n1631 , \GFM/n16300 , \GFM/n1629 ,\GFM/n16280 , \GFM/n16270 , \GFM/n1626 , \GFM/n1625 , \GFM/n1624 ,\GFM/n16230 , \GFM/n16220 , \GFM/n1621 , \GFM/n16200 , \GFM/n16190 ,\GFM/n1618 , \GFM/n1617 , \GFM/n16160 , \GFM/n16150 , \GFM/n1614 ,\GFM/n16130 , \GFM/n1612 , \GFM/n1611 , \GFM/n1610 , \GFM/n16090 ,\GFM/n16080 , \GFM/n1607 , \GFM/n16060 , \GFM/n16050 , \GFM/n1604 ,\GFM/n1603 , \GFM/n16020 , \GFM/n16010 , \GFM/n1600 , \GFM/n15990 ,\GFM/n1598 , \GFM/n15970 , \GFM/n15960 , \GFM/n1595 , \GFM/n1594 ,\GFM/n1593 , \GFM/n15920 , \GFM/n15910 , \GFM/n1590 , \GFM/n15890 ,\GFM/n15880 , \GFM/n1587 , \GFM/n1586 , \GFM/n15850 , \GFM/n15840 ,\GFM/n1583 , \GFM/n15820 , \GFM/n1581 , \GFM/n1580 , \GFM/n1579 ,\GFM/n15780 , \GFM/n15770 , \GFM/n1576 , \GFM/n15750 , \GFM/n15740 ,\GFM/n1573 , \GFM/n1572 , \GFM/n15710 , \GFM/n15700 , \GFM/n1569 ,\GFM/n15680 , \GFM/n1567 , \GFM/n15660 , \GFM/n15650 , \GFM/n1564 ,\GFM/n1563 , \GFM/n1562 , \GFM/n15610 , \GFM/n15600 , \GFM/n1559 ,\GFM/n15580 , \GFM/n15570 , \GFM/n1556 , \GFM/n1555 , \GFM/n15540 ,\GFM/n15530 , \GFM/n1552 , \GFM/n15510 , \GFM/n1550 , \GFM/n1549 ,\GFM/n1548 , \GFM/n15470 , \GFM/n15460 , \GFM/n1545 , \GFM/n15440 ,\GFM/n15430 , \GFM/n1542 , \GFM/n1541 , \GFM/n15400 , \GFM/n15390 ,\GFM/n1538 , \GFM/n15370 , \GFM/n1536 , \GFM/n15350 , \GFM/n15340 ,\GFM/n1533 , \GFM/n1532 , \GFM/n1531 , \GFM/n15300 , \GFM/n15290 ,\GFM/n1528 , \GFM/n15270 , \GFM/n15260 , \GFM/n1525 , \GFM/n1524 ,\GFM/n15230 , \GFM/n15220 , \GFM/n1521 , \GFM/n15200 , \GFM/n1519 ,\GFM/n1518 , \GFM/n1517 , \GFM/n15160 , \GFM/n15150 , \GFM/n1514 ,\GFM/n15130 , \GFM/n15120 , \GFM/n1511 , \GFM/n1510 , \GFM/n15090 ,\GFM/n15080 , \GFM/n1507 , \GFM/n15060 , \GFM/n1505 , \GFM/n15040 ,\GFM/n15030 , \GFM/n1502 , \GFM/n1501 , \GFM/n1500 , \GFM/n14990 ,\GFM/n14980 , \GFM/n1497 , \GFM/n14960 , \GFM/n14950 , \GFM/n1494 ,\GFM/n1493 , \GFM/n14920 , \GFM/n14910 , \GFM/n1490 , \GFM/n14890 ,\GFM/n1488 , \GFM/n1487 , \GFM/n1486 , \GFM/n14850 , \GFM/n14840 ,\GFM/n1483 , \GFM/n14820 , \GFM/n14810 , \GFM/n1480 , \GFM/n1479 ,\GFM/n14780 , \GFM/n14770 , \GFM/n1476 , \GFM/n14750 , \GFM/n1474 ,\GFM/n14730 , \GFM/n14720 , \GFM/n1471 , \GFM/n1470 , \GFM/n1469 ,\GFM/n14680 , \GFM/n14670 , \GFM/n1466 , \GFM/n14650 , \GFM/n14640 ,\GFM/n1463 , \GFM/n1462 , \GFM/n14610 , \GFM/n14600 , \GFM/n1459 ,\GFM/n14580 , \GFM/n1457 , \GFM/n1456 , \GFM/n1455 , \GFM/n14540 ,\GFM/n14530 , \GFM/n1452 , \GFM/n14510 , \GFM/n14500 , \GFM/n1449 ,\GFM/n1448 , \GFM/n14470 , \GFM/n14460 , \GFM/n1445 , \GFM/n14440 ,\GFM/n1443 , \GFM/n14420 , \GFM/n14410 , \GFM/n1440 , \GFM/n1439 ,\GFM/n1438 , \GFM/n14370 , \GFM/n14360 , \GFM/n1435 , \GFM/n14340 ,\GFM/n14330 , \GFM/n1432 , \GFM/n1431 , \GFM/n14300 , \GFM/n14290 ,\GFM/n1428 , \GFM/n14270 , \GFM/n1426 , \GFM/n1425 , \GFM/n1424 ,\GFM/n14230 , \GFM/n14220 , \GFM/n1421 , \GFM/n14200 , \GFM/n14190 ,\GFM/n1418 , \GFM/n1417 , \GFM/n14160 , \GFM/n14150 , \GFM/n1414 ,\GFM/n14130 , \GFM/n1412 , \GFM/n14110 , \GFM/n14100 , \GFM/n1409 ,\GFM/n1408 , \GFM/n1407 , \GFM/n14060 , \GFM/n14050 , \GFM/n1404 ,\GFM/n14030 , \GFM/n14020 , \GFM/n1401 , \GFM/n1400 , \GFM/n13990 ,\GFM/n13980 , \GFM/n1397 , \GFM/n13960 , \GFM/n1395 , \GFM/n1394 ,\GFM/n1393 , \GFM/n13920 , \GFM/n13910 , \GFM/n1390 , \GFM/n13890 ,\GFM/n13880 , \GFM/n1387 , \GFM/n1386 , \GFM/n13850 , \GFM/n13840 ,\GFM/n1383 , \GFM/n13820 , \GFM/n1381 , \GFM/n13800 , \GFM/n13790 ,\GFM/n1378 , \GFM/n1377 , \GFM/n1376 , \GFM/n13750 , \GFM/n13740 ,\GFM/n1373 , \GFM/n13720 , \GFM/n13710 , \GFM/n1370 , \GFM/n1369 ,\GFM/n13680 , \GFM/n13670 , \GFM/n1366 , \GFM/n13650 , \GFM/n1364 ,\GFM/n1363 , \GFM/n1362 , \GFM/n13610 , \GFM/n13600 , \GFM/n1359 ,\GFM/n13580 , \GFM/n13570 , \GFM/n1356 , \GFM/n1355 , \GFM/n13540 ,\GFM/n13530 , \GFM/n1352 , \GFM/n13510 , \GFM/n1350 , \GFM/n13490 ,\GFM/n13480 , \GFM/n1347 , \GFM/n1346 , \GFM/n1345 , \GFM/n13440 ,\GFM/n13430 , \GFM/n1342 , \GFM/n13410 , \GFM/n13400 , \GFM/n1339 ,\GFM/n1338 , \GFM/n13370 , \GFM/n13360 , \GFM/n1335 , \GFM/n13340 ,\GFM/n1333 , \GFM/n1332 , \GFM/n1331 , \GFM/n13300 , \GFM/n13290 ,\GFM/n1328 , \GFM/n13270 , \GFM/n13260 , \GFM/n1325 , \GFM/n1324 ,\GFM/n13230 , \GFM/n13220 , \GFM/n1321 , \GFM/n13200 , \GFM/n1319 ,\GFM/n13180 , \GFM/n13170 , \GFM/n1316 , \GFM/n1315 , \GFM/n1314 ,\GFM/n13130 , \GFM/n13120 , \GFM/n1311 , \GFM/n13100 , \GFM/n13090 ,\GFM/n1308 , \GFM/n1307 , \GFM/n13060 , \GFM/n13050 , \GFM/n1304 ,\GFM/n13030 , \GFM/n1302 , \GFM/n1301 , \GFM/n1300 , \GFM/n12990 ,\GFM/n12980 , \GFM/n1297 , \GFM/n12960 , \GFM/n12950 , \GFM/n1294 ,\GFM/n1293 , \GFM/n12920 , \GFM/n12910 , \GFM/n1290 , \GFM/n12890 ,\GFM/n1288 , \GFM/n12870 , \GFM/n12860 , \GFM/n1285 , \GFM/n1284 ,\GFM/n1283 , \GFM/n12820 , \GFM/n12810 , \GFM/n1280 , \GFM/n12790 ,\GFM/n12780 , \GFM/n1277 , \GFM/n1276 , \GFM/n12750 , \GFM/n12740 ,\GFM/n1273 , \GFM/n12720 , \GFM/n1271 , \GFM/n1270 , \GFM/n1269 ,\GFM/n12680 , \GFM/n12670 , \GFM/n1266 , \GFM/n12650 , \GFM/n12640 ,\GFM/n1263 , \GFM/n1262 , \GFM/n12610 , \GFM/n12600 , \GFM/n1259 ,\GFM/n12580 , \GFM/n1257 , \GFM/n12560 , \GFM/n12550 , \GFM/n1254 ,\GFM/n1253 , \GFM/n1252 , \GFM/n12510 , \GFM/n12500 , \GFM/n1249 ,\GFM/n12480 , \GFM/n12470 , \GFM/n1246 , \GFM/n1245 , \GFM/n12440 ,\GFM/n12430 , \GFM/n1242 , \GFM/n12410 , \GFM/n1240 , \GFM/n1239 ,\GFM/n1238 , \GFM/n12370 , \GFM/n12360 , \GFM/n1235 , \GFM/n12340 ,\GFM/n12330 , \GFM/n1232 , \GFM/n1231 , \GFM/n12300 , \GFM/n12290 ,\GFM/n1228 , \GFM/n12270 , \GFM/n1226 , \GFM/n12250 , \GFM/n12240 ,\GFM/n1223 , \GFM/n1222 , \GFM/n1221 , \GFM/n12200 , \GFM/n12190 ,\GFM/n1218 , \GFM/n12170 , \GFM/n12160 , \GFM/n1215 , \GFM/n1214 ,\GFM/n12130 , \GFM/n12120 , \GFM/n1211 , \GFM/n12100 , \GFM/n1209 ,\GFM/n1208 , \GFM/n1207 , \GFM/n12060 , \GFM/n12050 , \GFM/n1204 ,\GFM/n12030 , \GFM/n12020 , \GFM/n1201 , \GFM/n1200 , \GFM/n11990 ,\GFM/n11980 , \GFM/n1197 , \GFM/n11960 , \GFM/n1195 , \GFM/n11940 ,\GFM/n11930 , \GFM/n1192 , \GFM/n1191 , \GFM/n1190 , \GFM/n11890 ,\GFM/n11880 , \GFM/n1187 , \GFM/n11860 , \GFM/n11850 , \GFM/n1184 ,\GFM/n1183 , \GFM/n11820 , \GFM/n11810 , \GFM/n1180 , \GFM/n11790 ,\GFM/n1178 , \GFM/n1177 , \GFM/n1176 , \GFM/n11750 , \GFM/n11740 ,\GFM/n1173 , \GFM/n11720 , \GFM/n11710 , \GFM/n1170 , \GFM/n1169 ,\GFM/n11680 , \GFM/n11670 , \GFM/n1166 , \GFM/n11650 , \GFM/n1164 ,\GFM/n11630 , \GFM/n11620 , \GFM/n1161 , \GFM/n1160 , \GFM/n1159 ,\GFM/n11580 , \GFM/n11570 , \GFM/n1156 , \GFM/n11550 , \GFM/n11540 ,\GFM/n1153 , \GFM/n1152 , \GFM/n11510 , \GFM/n11500 , \GFM/n1149 ,\GFM/n11480 , \GFM/n1147 , \GFM/n1146 , \GFM/n1145 , \GFM/n11440 ,\GFM/n11430 , \GFM/n1142 , \GFM/n11410 , \GFM/n11400 , \GFM/n1139 ,\GFM/n1138 , \GFM/n11370 , \GFM/n11360 , \GFM/n1135 , \GFM/n11340 ,\GFM/n1133 , \GFM/n11320 , \GFM/n11310 , \GFM/n1130 , \GFM/n1129 ,\GFM/n1128 , \GFM/n11270 , \GFM/n11260 , \GFM/n1125 , \GFM/n11240 ,\GFM/n11230 , \GFM/n1122 , \GFM/n1121 , \GFM/n11200 , \GFM/n11190 ,\GFM/n1118 , \GFM/n11170 , \GFM/n1116 , \GFM/n1115 , \GFM/n1114 ,\GFM/n11130 , \GFM/n11120 , \GFM/n1111 , \GFM/n11100 , \GFM/n11090 ,\GFM/n1108 , \GFM/n1107 , \GFM/n11060 , \GFM/n11050 , \GFM/n1104 ,\GFM/n11030 , \GFM/n1102 , \GFM/n11010 , \GFM/n11000 , \GFM/n1099 ,\GFM/n1098 , \GFM/n1097 , \GFM/n10960 , \GFM/n10950 , \GFM/n1094 ,\GFM/n10930 , \GFM/n10920 , \GFM/n1091 , \GFM/n1090 , \GFM/n10890 ,\GFM/n10880 , \GFM/n1087 , \GFM/n10860 , \GFM/n1085 , \GFM/n1084 ,\GFM/n1083 , \GFM/n10820 , \GFM/n10810 , \GFM/n1080 , \GFM/n10790 ,\GFM/n10780 , \GFM/n1077 , \GFM/n1076 , \GFM/n10750 , \GFM/n10740 ,\GFM/n1073 , \GFM/n10720 , \GFM/n1071 , \GFM/n10700 , \GFM/n10690 ,\GFM/n1068 , \GFM/n1067 , \GFM/n1066 , \GFM/n10650 , \GFM/n10640 ,\GFM/n1063 , \GFM/n10620 , \GFM/n10610 , \GFM/n1060 , \GFM/n1059 ,\GFM/n10580 , \GFM/n10570 , \GFM/n1056 , \GFM/n10550 , \GFM/n1054 ,\GFM/n1053 , \GFM/n1052 , \GFM/n10510 , \GFM/n10500 , \GFM/n1049 ,\GFM/n10480 , \GFM/n10470 , \GFM/n1046 , \GFM/n1045 , \GFM/n10440 ,\GFM/n10430 , \GFM/n1042 , \GFM/n10410 , \GFM/n1040 , \GFM/n10390 ,\GFM/n10380 , \GFM/n1037 , \GFM/n1036 , \GFM/n1035 , \GFM/n10340 ,\GFM/n10330 , \GFM/n1032 , \GFM/n10310 , \GFM/n10300 , \GFM/n1029 ,\GFM/n1028 , \GFM/n10270 , \GFM/n10260 , \GFM/n1025 , \GFM/n10240 ,\GFM/n1023 , \GFM/n1022 , \GFM/n1021 , \GFM/n10200 , \GFM/n10190 ,\GFM/n1018 , \GFM/n10170 , \GFM/n10160 , \GFM/n1015 , \GFM/n1014 ,\GFM/n10130 , \GFM/n10120 , \GFM/n1011 , \GFM/n10100 , \GFM/n1009 ,\GFM/n10080 , \GFM/n10070 , \GFM/n1006 , \GFM/n1005 , \GFM/n1004 ,\GFM/n10030 , \GFM/n10020 , \GFM/n1001 , \GFM/n10000 , \GFM/n9990 ,\GFM/n998 , \GFM/n997 , \GFM/n9960 , \GFM/n9950 , \GFM/n994 ,\GFM/n9930 , \GFM/n992 , \GFM/n991 , \GFM/n990 , \GFM/n9890 ,\GFM/n9880 , \GFM/n987 , \GFM/n9860 , \GFM/n9850 , \GFM/n984 ,\GFM/n983 , \GFM/n9820 , \GFM/n9810 , \GFM/n980 , \GFM/n9790 ,\GFM/n978 , \GFM/n9770 , \GFM/n9760 , \GFM/n975 , \GFM/n974 ,\GFM/n973 , \GFM/n9720 , \GFM/n9710 , \GFM/n970 , \GFM/n9690 ,\GFM/n9680 , \GFM/n967 , \GFM/n966 , \GFM/n9650 , \GFM/n9640 ,\GFM/n963 , \GFM/n9620 , \GFM/n961 , \GFM/n960 , \GFM/n959 ,\GFM/n9580 , \GFM/n9570 , \GFM/n956 , \GFM/n9550 , \GFM/n9540 ,\GFM/n953 , \GFM/n952 , \GFM/n9510 , \GFM/n9500 , \GFM/n949 ,\GFM/n9480 , \GFM/n947 , \GFM/n9460 , \GFM/n9450 , \GFM/n944 ,\GFM/n943 , \GFM/n942 , \GFM/n9410 , \GFM/n9400 , \GFM/n939 ,\GFM/n9380 , \GFM/n9370 , \GFM/n936 , \GFM/n935 , \GFM/n9340 ,\GFM/n9330 , \GFM/n932 , \GFM/n9310 , \GFM/n930 , \GFM/n929 ,\GFM/n928 , \GFM/n9270 , \GFM/n9260 , \GFM/n925 , \GFM/n9240 ,\GFM/n9230 , \GFM/n922 , \GFM/n921 , \GFM/n9200 , \GFM/n9190 ,\GFM/n918 , \GFM/n9170 , \GFM/n916 , \GFM/n9150 , \GFM/n9140 ,\GFM/n913 , \GFM/n912 , \GFM/n911 , \GFM/n9100 , \GFM/n9090 ,\GFM/n908 , \GFM/n9070 , \GFM/n9060 , \GFM/n905 , \GFM/n904 ,\GFM/n9030 , \GFM/n9020 , \GFM/n901 , \GFM/n9000 , \GFM/n899 ,\GFM/n898 , \GFM/n897 , \GFM/n8960 , \GFM/n8950 , \GFM/n894 ,\GFM/n8930 , \GFM/n8920 , \GFM/n891 , \GFM/n890 , \GFM/n8890 ,\GFM/n8880 , \GFM/n887 , \GFM/n8860 , \GFM/n885 , \GFM/n8840 ,\GFM/n8830 , \GFM/n882 , \GFM/n881 , \GFM/n880 , \GFM/n8790 ,\GFM/n8780 , \GFM/n877 , \GFM/n8760 , \GFM/n8750 , \GFM/n874 ,\GFM/n873 , \GFM/n8720 , \GFM/n8710 , \GFM/n870 , \GFM/n8690 ,\GFM/n868 , \GFM/n867 , \GFM/n866 , \GFM/n8650 , \GFM/n8640 ,\GFM/n863 , \GFM/n8620 , \GFM/n8610 , \GFM/n860 , \GFM/n859 ,\GFM/n8580 , \GFM/n8570 , \GFM/n856 , \GFM/n8550 , \GFM/n854 ,\GFM/n8530 , \GFM/n8520 , \GFM/n851 , \GFM/n850 , \GFM/n849 ,\GFM/n8480 , \GFM/n8470 , \GFM/n846 , \GFM/n8450 , \GFM/n8440 ,\GFM/n843 , \GFM/n842 , \GFM/n8410 , \GFM/n8400 , \GFM/n839 ,\GFM/n8380 , \GFM/n837 , \GFM/n836 , \GFM/n835 , \GFM/n8340 ,\GFM/n8330 , \GFM/n832 , \GFM/n8310 , \GFM/n8300 , \GFM/n829 ,\GFM/n828 , \GFM/n8270 , \GFM/n8260 , \GFM/n825 , \GFM/n8240 ,\GFM/n823 , \GFM/n8220 , \GFM/n8210 , \GFM/n820 , \GFM/n819 ,\GFM/n818 , \GFM/n8170 , \GFM/n8160 , \GFM/n815 , \GFM/n8140 ,\GFM/n8130 , \GFM/n812 , \GFM/n811 , \GFM/n8100 , \GFM/n8090 ,\GFM/n808 , \GFM/n8070 , \GFM/n806 , \GFM/n805 , \GFM/n804 ,\GFM/n8030 , \GFM/n8020 , \GFM/n801 , \GFM/n8000 , \GFM/n7990 ,\GFM/n798 , \GFM/n797 , \GFM/n7960 , \GFM/n7950 , \GFM/n794 ,\GFM/n7930 , \GFM/n792 , \GFM/n7910 , \GFM/n7900 , \GFM/n789 ,\GFM/n788 , \GFM/n787 , \GFM/n7860 , \GFM/n7850 , \GFM/n784 ,\GFM/n7830 , \GFM/n7820 , \GFM/n781 , \GFM/n780 , \GFM/n7790 ,\GFM/n7780 , \GFM/n777 , \GFM/n7760 , \GFM/n775 , \GFM/n774 ,\GFM/n773 , \GFM/n7720 , \GFM/n7710 , \GFM/n770 , \GFM/n7690 ,\GFM/n7680 , \GFM/n767 , \GFM/n766 , \GFM/n7650 , \GFM/n7640 ,\GFM/n763 , \GFM/n7620 , \GFM/n761 , \GFM/n7600 , \GFM/n7590 ,\GFM/n758 , \GFM/n757 , \GFM/n756 , \GFM/n7550 , \GFM/n7540 ,\GFM/n753 , \GFM/n7520 , \GFM/n7510 , \GFM/n750 , \GFM/n749 ,\GFM/n7480 , \GFM/n7470 , \GFM/n746 , \GFM/n7450 , \GFM/n744 ,\GFM/n743 , \GFM/n742 , \GFM/n7410 , \GFM/n7400 , \GFM/n739 ,\GFM/n7380 , \GFM/n7370 , \GFM/n736 , \GFM/n735 , \GFM/n7340 ,\GFM/n7330 , \GFM/n732 , \GFM/n7310 , \GFM/n730 , \GFM/n7290 ,\GFM/n7280 , \GFM/n727 , \GFM/n726 , \GFM/n725 , \GFM/n7240 ,\GFM/n7230 , \GFM/n722 , \GFM/n7210 , \GFM/n7200 , \GFM/n719 ,\GFM/n718 , \GFM/n7170 , \GFM/n7160 , \GFM/n715 , \GFM/n7140 ,\GFM/n713 , \GFM/n712 , \GFM/n711 , \GFM/n7100 , \GFM/n7090 ,\GFM/n708 , \GFM/n7070 , \GFM/n7060 , \GFM/n705 , \GFM/n704 ,\GFM/n7030 , \GFM/n7020 , \GFM/n701 , \GFM/n7000 , \GFM/n699 ,\GFM/n6980 , \GFM/n6970 , \GFM/n696 , \GFM/n695 , \GFM/n694 ,\GFM/n6930 , \GFM/n6920 , \GFM/n691 , \GFM/n6900 , \GFM/n6890 ,\GFM/n688 , \GFM/n687 , \GFM/n6860 , \GFM/n6850 , \GFM/n684 ,\GFM/n6830 , \GFM/n682 , \GFM/n681 , \GFM/n680 , \GFM/n6790 ,\GFM/n6780 , \GFM/n677 , \GFM/n6760 , \GFM/n6750 , \GFM/n674 ,\GFM/n673 , \GFM/n6720 , \GFM/n6710 , \GFM/n670 , \GFM/n6690 ,\GFM/n668 , \GFM/n6670 , \GFM/n6660 , \GFM/n665 , \GFM/n664 ,\GFM/n663 , \GFM/n6620 , \GFM/n6610 , \GFM/n660 , \GFM/n6590 ,\GFM/n6580 , \GFM/n657 , \GFM/n656 , \GFM/n6550 , \GFM/n6540 ,\GFM/n653 , \GFM/n6520 , \GFM/n651 , \GFM/n650 , \GFM/n649 ,\GFM/n6480 , \GFM/n6470 , \GFM/n646 , \GFM/n6450 , \GFM/n6440 ,\GFM/n643 , \GFM/n642 , \GFM/n6410 , \GFM/n6400 , \GFM/n639 ,\GFM/n6380 , \GFM/n637 , \GFM/n6360 , \GFM/n6350 , \GFM/n634 ,\GFM/n633 , \GFM/n632 , \GFM/n6310 , \GFM/n6300 , \GFM/n629 ,\GFM/n6280 , \GFM/n6270 , \GFM/n626 , \GFM/n625 , \GFM/n6240 ,\GFM/n6230 , \GFM/n622 , \GFM/n6210 , \GFM/n620 , \GFM/n619 ,\GFM/n618 , \GFM/n6170 , \GFM/n6160 , \GFM/n615 , \GFM/n6140 ,\GFM/n6130 , \GFM/n612 , \GFM/n611 , \GFM/n6100 , \GFM/n6090 ,\GFM/n608 , \GFM/n6070 , \GFM/n606 , \GFM/n6050 , \GFM/n6040 ,\GFM/n603 , \GFM/n602 , \GFM/n601 , \GFM/n6000 , \GFM/n5990 ,\GFM/n598 , \GFM/n5970 , \GFM/n5960 , \GFM/n595 , \GFM/n594 ,\GFM/n5930 , \GFM/n5920 , \GFM/n591 , \GFM/n5900 , \GFM/n589 ,\GFM/n588 , \GFM/n587 , \GFM/n5860 , \GFM/n5850 , \GFM/n584 ,\GFM/n5830 , \GFM/n5820 , \GFM/n581 , \GFM/n580 , \GFM/n5790 ,\GFM/n5780 , \GFM/n577 , \GFM/n5760 , \GFM/n575 , \GFM/n5740 ,\GFM/n5730 , \GFM/n572 , \GFM/n571 , \GFM/n570 , \GFM/n5690 ,\GFM/n5680 , \GFM/n567 , \GFM/n5660 , \GFM/n5650 , \GFM/n564 ,\GFM/n563 , \GFM/n5620 , \GFM/n5610 , \GFM/n560 , \GFM/n5590 ,\GFM/n558 , \GFM/n557 , \GFM/n556 , \GFM/n5550 , \GFM/n5540 ,\GFM/n553 , \GFM/n5520 , \GFM/n5510 , \GFM/n550 , \GFM/n549 ,\GFM/n5480 , \GFM/n5470 , \GFM/n546 , \GFM/n5450 , \GFM/n544 ,\GFM/n5430 , \GFM/n5420 , \GFM/n541 , \GFM/n540 , \GFM/n539 ,\GFM/n5380 , \GFM/n5370 , \GFM/n536 , \GFM/n5350 , \GFM/n5340 ,\GFM/n533 , \GFM/n532 , \GFM/n5310 , \GFM/n5300 , \GFM/n529 ,\GFM/n5280 , \GFM/n527 , \GFM/n526 , \GFM/n525 , \GFM/n5240 ,\GFM/n5230 , \GFM/n522 , \GFM/n5210 , \GFM/n5200 , \GFM/n519 ,\GFM/n518 , \GFM/n5170 , \GFM/n5160 , \GFM/n515 , \GFM/n5140 ,\GFM/n513 , \GFM/n5120 , \GFM/n5110 , \GFM/n510 , \GFM/n509 ,\GFM/n508 , \GFM/n5070 , \GFM/n5060 , \GFM/n505 , \GFM/n5040 ,\GFM/n5030 , \GFM/n502 , \GFM/n501 , \GFM/n5000 , \GFM/n4990 ,\GFM/n498 , \GFM/n4970 , \GFM/n496 , \GFM/n495 , \GFM/n494 ,\GFM/n4930 , \GFM/n4920 , \GFM/n491 , \GFM/n4900 , \GFM/n4890 ,\GFM/n488 , \GFM/n487 , \GFM/n4860 , \GFM/n4850 , \GFM/n484 ,\GFM/n4830 , \GFM/n482 , \GFM/n4810 , \GFM/n4800 , \GFM/n479 ,\GFM/n478 , \GFM/n477 , \GFM/n4760 , \GFM/n4750 , \GFM/n474 ,\GFM/n4730 , \GFM/n4720 , \GFM/n471 , \GFM/n470 , \GFM/n4690 ,\GFM/n4680 , \GFM/n467 , \GFM/n4660 , \GFM/n465 , \GFM/n464 ,\GFM/n463 , \GFM/n4620 , \GFM/n4610 , \GFM/n460 , \GFM/n4590 ,\GFM/n4580 , \GFM/n457 , \GFM/n456 , \GFM/n4550 , \GFM/n4540 ,\GFM/n453 , \GFM/n4520 , \GFM/n451 , \GFM/n4500 , \GFM/n4490 ,\GFM/n448 , \GFM/n447 , \GFM/n446 , \GFM/n4450 , \GFM/n4440 ,\GFM/n443 , \GFM/n4420 , \GFM/n4410 , \GFM/n440 , \GFM/n439 ,\GFM/n4380 , \GFM/n4370 , \GFM/n436 , \GFM/n4350 , \GFM/n434 ,\GFM/n433 , \GFM/n432 , \GFM/n4310 , \GFM/n4301 , \GFM/n429 ,\GFM/n4280 , \GFM/n4270 , \GFM/n426 , \GFM/n425 , \GFM/n4241 ,\GFM/n4230 , \GFM/n422 , \GFM/n4211 , \GFM/n420 , \GFM/n4190 ,\GFM/n4180 , \GFM/n417 , \GFM/n416 , \GFM/n415 , \GFM/n4140 ,\GFM/n4130 , \GFM/n412 , \GFM/n4110 , \GFM/n4100 , \GFM/n409 ,\GFM/n408 , \GFM/n4070 , \GFM/n4060 , \GFM/n405 , \GFM/n4040 ,\GFM/n403 , \GFM/n402 , \GFM/n401 , \GFM/n4000 , \GFM/n3991 ,\GFM/n398 , \GFM/n3970 , \GFM/n3960 , \GFM/n395 , \GFM/n394 ,\GFM/n3930 , \GFM/n3920 , \GFM/n391 , \GFM/n3900 , \GFM/n389 ,\GFM/n3880 , \GFM/n3870 , \GFM/n386 , \GFM/n385 , \GFM/n384 ,\GFM/n3830 , \GFM/n3820 , \GFM/n381 , \GFM/n3800 , \GFM/n3790 ,\GFM/n378 , \GFM/n377 , \GFM/n3760 , \GFM/n3751 , \GFM/n374 ,\GFM/n3730 , \GFM/n372 , \GFM/n371 , \GFM/n370 , \GFM/n3691 ,\GFM/n3680 , \GFM/n367 , \GFM/n3660 , \GFM/n3650 , \GFM/n364 ,\GFM/n363 , \GFM/n3621 , \GFM/n3610 , \GFM/n360 , \GFM/n3590 ,\GFM/n358 , \GFM/n3570 , \GFM/n3560 , \GFM/n355 , \GFM/n354 ,\GFM/n353 , \GFM/n3520 , \GFM/n3510 , \GFM/n350 , \GFM/n3490 ,\GFM/n3480 , \GFM/n347 , \GFM/n346 , \GFM/n3451 , \GFM/n3440 ,\GFM/n343 , \GFM/n3420 , \GFM/n341 , \GFM/n340 , \GFM/n339 ,\GFM/n3381 , \GFM/n3370 , \GFM/n336 , \GFM/n3350 , \GFM/n3342 ,\GFM/n333 , \GFM/n332 , \GFM/n3310 , \GFM/n3300 , \GFM/n329 ,\GFM/n3281 , \GFM/n327 , \GFM/n3260 , \GFM/n3250 , \GFM/n324 ,\GFM/n323 , \GFM/n322 , \GFM/n3210 , \GFM/n3202 , \GFM/n319 ,\GFM/n3181 , \GFM/n3171 , \GFM/n316 , \GFM/n315 , \GFM/n3140 ,\GFM/n3130 , \GFM/n312 , \GFM/n3112 , \GFM/n310 , \GFM/n309 ,\GFM/n308 , \GFM/n3071 , \GFM/n3060 , \GFM/n305 , \GFM/n3040 ,\GFM/n3030 , \GFM/n302 , \GFM/n301 , \GFM/n3002 , \GFM/n2990 ,\GFM/n298 , \GFM/n2971 , \GFM/n296 , \GFM/n2950 , \GFM/n2940 ,\GFM/n293 , \GFM/n292 , \GFM/n291 , \GFM/n2900 , \GFM/n2892 ,\GFM/n288 , \GFM/n2871 , \GFM/n2861 , \GFM/n285 , \GFM/n284 ,\GFM/n2830 , \GFM/n2820 , \GFM/n281 , \GFM/n2802 , \GFM/n279 ,\GFM/n278 , \GFM/n277 , \GFM/n2761 , \GFM/n2750 , \GFM/n274 ,\GFM/n2730 , \GFM/n2720 , \GFM/n271 , \GFM/n270 , \GFM/n26920 ,\GFM/n26800 , \GFM/n267 , \GFM/n26610 , \GFM/n265 , \GFM/n26400 ,\GFM/n26300 , \GFM/n262 , \GFM/n261 , \GFM/n260 , \GFM/n25900 ,\GFM/n25820 , \GFM/n257 , \GFM/n25610 , \GFM/n25510 , \GFM/n254 ,\GFM/n253 , \GFM/n25200 , \GFM/n25100 , \GFM/n250 , \GFM/n24920 ,\GFM/n248 , \GFM/n247 , \GFM/n246 , \GFM/n24510 , \GFM/n24400 ,\GFM/n243 , \GFM/n24200 , \GFM/n24100 , \GFM/n240 , \GFM/n239 ,\GFM/n2382 , \GFM/n2370 , \GFM/n236 , \GFM/n2351 , \GFM/n234 ,\GFM/n2330 , \GFM/n2320 , \GFM/n231 , \GFM/n230 , \GFM/n229 ,\GFM/n2280 , \GFM/n2272 , \GFM/n226 , \GFM/n2251 , \GFM/n2241 ,\GFM/n223 , \GFM/n222 , \GFM/n2210 , \GFM/n2200 , \GFM/n219 ,\GFM/n2182 , \GFM/n217 , \GFM/n216 , \GFM/n215 , \GFM/n2141 ,\GFM/n21300 , \GFM/n212 , \GFM/n21100 , \GFM/n21000 , \GFM/n209 ,\GFM/n208 , \GFM/n20720 , \GFM/n20600 , \GFM/n205 , \GFM/n20410 ,\GFM/n203 , \GFM/n20200 , \GFM/n20100 , \GFM/n200 , \GFM/n199 ,\GFM/n198 , \GFM/n19700 , \GFM/n19620 , \GFM/n195 , \GFM/n19410 ,\GFM/n19310 , \GFM/n192 , \GFM/n191 , \GFM/n19000 , \GFM/n18900 ,\GFM/n188 , \GFM/n18720 , \GFM/n186 , \GFM/n185 , \GFM/N4349 ,\GFM/N4348 , \GFM/N4346 , \GFM/N4345 , \GFM/N4342 , \GFM/N4341 ,\GFM/N4339 , \GFM/N4337 , \GFM/N4336 , \GFM/N4332 , \GFM/N4331 ,\GFM/N4329 , \GFM/N4328 , \GFM/N4325 , \GFM/N4324 , \GFM/N4322 ,\GFM/N4318 , \GFM/N4316 , \GFM/N4313 , \GFM/N4311 , \GFM/N4307 ,\GFM/N4305 , \GFM/N4302 , \GFM/N4300 , \GFM/N4295 , \GFM/N4293 ,\GFM/N4290 , \GFM/N4288 , \GFM/N4284 , \GFM/N4282 , \GFM/N4279 ,\GFM/N4276 , \GFM/N4272 , \GFM/N4269 , \GFM/N4265 , \GFM/N4263 ,\GFM/N4258 , \GFM/N4257 , \GFM/N4255 , \GFM/N4254 , \GFM/N4251 ,\GFM/N4250 , \GFM/N4249 , \GFM/N4248 , \GFM/N4243 , \GFM/N4242 ,\GFM/N4240 , \GFM/N4239 , \GFM/N4236 , \GFM/N4235 , \GFM/N4233 ,\GFM/N4232 , \GFM/N4228 , \GFM/N4227 , \GFM/N4225 , \GFM/N4224 ,\GFM/N4221 , \GFM/N4218 , \GFM/N4213 , \GFM/N4210 , \GFM/N4206 ,\GFM/N4203 , \GFM/N4198 , \GFM/N4195 , \GFM/N4191 , \GFM/N4188 ,\GFM/N4182 , \GFM/N4179 , \GFM/N4175 , \GFM/N4172 , \GFM/N4167 ,\GFM/N4164 , \GFM/N4160 , \GFM/N4159 , \GFM/N4154 , \GFM/N4151 ,\GFM/N4147 , \GFM/N4144 , \GFM/N4139 , \GFM/N4136 , \GFM/N4132 ,\GFM/N4129 , \GFM/N4123 , \GFM/N4120 , \GFM/N4116 , \GFM/N4113 ,\GFM/N4108 , \GFM/N4106 , \GFM/N4103 , \GFM/N4102 , \GFM/N4097 ,\GFM/N4094 , \GFM/N4090 , \GFM/N4087 , \GFM/N4082 , \GFM/N4079 ,\GFM/N4075 , \GFM/N4072 , \GFM/N4066 , \GFM/N4063 , \GFM/N4059 ,\GFM/N4057 , \GFM/N4052 , \GFM/N4050 , \GFM/N4049 , \GFM/N4047 ,\GFM/N4042 , \GFM/N4039 , \GFM/N4035 , \GFM/N4032 , \GFM/N4027 ,\GFM/N4024 , \GFM/N4020 , \GFM/N4017 , \GFM/N4012 , \GFM/N4007 ,\GFM/N4006 , \GFM/N4004 , \GFM/N3999 , \GFM/N3997 , \GFM/N3996 ,\GFM/N3994 , \GFM/N3990 , \GFM/N3985 , \GFM/N3981 , \GFM/N3975 ,\GFM/N3971 , \GFM/N3966 , \GFM/N3962 , \GFM/N3955 , \GFM/N3951 ,\GFM/N3946 , \GFM/N3944 , \GFM/N3939 , \GFM/N3936 , \GFM/N3934 ,\GFM/N3931 , \GFM/N3928 , \GFM/N3923 , \GFM/N3918 , \GFM/N3914 ,\GFM/N3908 , \GFM/N3904 , \GFM/N3899 , \GFM/N3895 , \GFM/N3889 ,\GFM/N3883 , \GFM/N3881 , \GFM/N3879 , \GFM/N3874 , \GFM/N3871 ,\GFM/N3869 , \GFM/N3865 , \GFM/N3864 , \GFM/N3859 , \GFM/N3854 ,\GFM/N3850 , \GFM/N3844 , \GFM/N3840 , \GFM/N3835 , \GFM/N3831 ,\GFM/N3825 , \GFM/N3821 , \GFM/N3818 , \GFM/N3816 , \GFM/N3812 ,\GFM/N3809 , \GFM/N3808 , \GFM/N3804 , \GFM/N3803 , \GFM/N3798 ,\GFM/N3793 , \GFM/N3789 , \GFM/N3783 , \GFM/N3780 , \GFM/N3775 ,\GFM/N3771 , \GFM/N3764 , \GFM/N3762 , \GFM/N3759 , \GFM/N3756 ,\GFM/N3754 , \GFM/N3750 , \GFM/N3748 , \GFM/N3747 , \GFM/N3745 ,\GFM/N3740 , \GFM/N3735 , \GFM/N3731 , \GFM/N3725 , \GFM/N3723 ,\GFM/N3719 , \GFM/N3715 , \GFM/N3708 , \GFM/N3706 , \GFM/N3703 ,\GFM/N3701 , \GFM/N3699 , \GFM/N3695 , \GFM/N3693 , \GFM/N3692 ,\GFM/N3690 , \GFM/N3685 , \GFM/N3681 , \GFM/N3674 , \GFM/N3672 ,\GFM/N3670 , \GFM/N3666 , \GFM/N3662 , \GFM/N3655 , \GFM/N3653 ,\GFM/N3649 , \GFM/N3648 , \GFM/N3647 , \GFM/N3643 , \GFM/N3641 ,\GFM/N3640 , \GFM/N3638 , \GFM/N3633 , \GFM/N3629 , \GFM/N3623 ,\GFM/N3620 , \GFM/N3618 , \GFM/N3615 , \GFM/N3611 , \GFM/N3605 ,\GFM/N3603 , \GFM/N3600 , \GFM/N3598 , \GFM/N3597 , \GFM/N3594 ,\GFM/N3592 , \GFM/N3591 , \GFM/N3589 , \GFM/N3584 , \GFM/N3580 ,\GFM/N3574 , \GFM/N3571 , \GFM/N3569 , \GFM/N3566 , \GFM/N3563 ,\GFM/N3558 , \GFM/N3556 , \GFM/N3554 , \GFM/N3552 , \GFM/N3551 ,\GFM/N3548 , \GFM/N3546 , \GFM/N3545 , \GFM/N3543 , \GFM/N3538 ,\GFM/N3534 , \GFM/N3529 , \GFM/N3527 , \GFM/N3524 , \GFM/N3521 ,\GFM/N3519 , \GFM/N3514 , \GFM/N3513 , \GFM/N3511 , \GFM/N3509 ,\GFM/N3508 , \GFM/N3505 , \GFM/N3503 , \GFM/N3502 , \GFM/N3500 ,\GFM/N3495 , \GFM/N3491 , \GFM/N3489 , \GFM/N3484 , \GFM/N3483 ,\GFM/N3482 , \GFM/N3479 , \GFM/N3477 , \GFM/N3472 , \GFM/N3471 ,\GFM/N3469 , \GFM/N3467 , \GFM/N3466 , \GFM/N3463 , \GFM/N3462 ,\GFM/N3460 , \GFM/N3455 , \GFM/N3452 , \GFM/N3450 , \GFM/N3446 ,\GFM/N3444 , \GFM/N3443 , \GFM/N3441 , \GFM/N3439 , \GFM/N3434 ,\GFM/N3433 , \GFM/N3431 , \GFM/N3429 , \GFM/N3428 , \GFM/N3425 ,\GFM/N3424 , \GFM/N3422 , \GFM/N3418 , \GFM/N3415 , \GFM/N3413 ,\GFM/N3409 , \GFM/N3407 , \GFM/N3406 , \GFM/N3404 , \GFM/N3402 ,\GFM/N3398 , \GFM/N3397 , \GFM/N3395 , \GFM/N3393 , \GFM/N3392 ,\GFM/N3389 , \GFM/N3388 , \GFM/N3386 , \GFM/N3383 , \GFM/N3380 ,\GFM/N3378 , \GFM/N3374 , \GFM/N3373 , \GFM/N3371 , \GFM/N3369 ,\GFM/N3368 , \GFM/N3364 , \GFM/N3363 , \GFM/N3361 , \GFM/N3359 ,\GFM/N3358 , \GFM/N3355 , \GFM/N3354 , \GFM/N3352 , \GFM/N3349 ,\GFM/N3346 , \GFM/N3345 , \GFM/N3341 , \GFM/N3340 , \GFM/N3338 ,\GFM/N3336 , \GFM/N3335 , \GFM/N3331 , \GFM/N3330 , \GFM/N3328 ,\GFM/N3326 , \GFM/N3325 , \GFM/N3322 , \GFM/N3321 , \GFM/N3319 ,\GFM/N3316 , \GFM/N3313 , \GFM/N3312 , \GFM/N3309 , \GFM/N3308 ,\GFM/N3306 , \GFM/N3304 , \GFM/N3303 , \GFM/N3299 , \GFM/N3298 ,\GFM/N3296 , \GFM/N3294 , \GFM/N3293 , \GFM/N3290 , \GFM/N3289 ,\GFM/N3287 , \GFM/N3283 , \GFM/N3282 , \GFM/N3280 , \GFM/N3279 ,\GFM/N3276 , \GFM/N3275 , \GFM/N3273 , \GFM/N3271 , \GFM/N3270 ,\GFM/N3266 , \GFM/N3265 , \GFM/N3263 , \GFM/N3262 , \GFM/N3259 ,\GFM/N3258 , \GFM/N3256 , \GFM/N3252 , \GFM/N3251 , \GFM/N3249 ,\GFM/N3248 , \GFM/N3245 , \GFM/N3244 , \GFM/N3242 , \GFM/N3240 ,\GFM/N3239 , \GFM/N3235 , \GFM/N3234 , \GFM/N3232 , \GFM/N3231 ,\GFM/N3228 , \GFM/N3227 , \GFM/N3225 , \GFM/N3221 , \GFM/N3220 ,\GFM/N3218 , \GFM/N3217 , \GFM/N3214 , \GFM/N3213 , \GFM/N3211 ,\GFM/N3209 , \GFM/N3208 , \GFM/N3204 , \GFM/N3203 , \GFM/N3201 ,\GFM/N3200 , \GFM/N3197 , \GFM/N3196 , \GFM/N3194 , \GFM/N3190 ,\GFM/N3189 , \GFM/N3187 , \GFM/N3186 , \GFM/N3183 , \GFM/N3182 ,\GFM/N3180 , \GFM/N3178 , \GFM/N3177 , \GFM/N3173 , \GFM/N3172 ,\GFM/N3170 , \GFM/N3169 , \GFM/N3166 , \GFM/N3165 , \GFM/N3163 ,\GFM/N3159 , \GFM/N3158 , \GFM/N3156 , \GFM/N3155 , \GFM/N3152 ,\GFM/N3151 , \GFM/N3149 , \GFM/N3147 , \GFM/N3146 , \GFM/N3142 ,\GFM/N3141 , \GFM/N3139 , \GFM/N3138 , \GFM/N3135 , \GFM/N3134 ,\GFM/N3132 , \GFM/N3128 , \GFM/N3127 , \GFM/N3125 , \GFM/N3124 ,\GFM/N3121 , \GFM/N3120 , \GFM/N3118 , \GFM/N3116 , \GFM/N3115 ,\GFM/N3111 , \GFM/N3110 , \GFM/N3108 , \GFM/N3107 , \GFM/N3104 ,\GFM/N3103 , \GFM/N3101 , \GFM/N3097 , \GFM/N3096 , \GFM/N3094 ,\GFM/N3093 , \GFM/N3090 , \GFM/N3089 , \GFM/N3087 , \GFM/N3085 ,\GFM/N3084 , \GFM/N3080 , \GFM/N3079 , \GFM/N3077 , \GFM/N3076 ,\GFM/N3073 , \GFM/N3072 , \GFM/N3070 , \GFM/N3066 , \GFM/N3065 ,\GFM/N3063 , \GFM/N3062 , \GFM/N3059 , \GFM/N3058 , \GFM/N3056 ,\GFM/N3054 , \GFM/N3053 , \GFM/N3049 , \GFM/N3048 , \GFM/N3046 ,\GFM/N3045 , \GFM/N3042 , \GFM/N3041 , \GFM/N3039 , \GFM/N3035 ,\GFM/N3034 , \GFM/N3032 , \GFM/N3031 , \GFM/N3028 , \GFM/N3027 ,\GFM/N3025 , \GFM/N3023 , \GFM/N3022 , \GFM/N3018 , \GFM/N3017 ,\GFM/N3015 , \GFM/N3014 , \GFM/N3011 , \GFM/N3010 , \GFM/N3008 ,\GFM/N3004 , \GFM/N3003 , \GFM/N3001 , \GFM/N3000 , \GFM/N2997 ,\GFM/N2996 , \GFM/N2994 , \GFM/N2992 , \GFM/N2991 , \GFM/N2987 ,\GFM/N2986 , \GFM/N2984 , \GFM/N2983 , \GFM/N2980 , \GFM/N2979 ,\GFM/N2977 , \GFM/N2973 , \GFM/N2972 , \GFM/N2970 , \GFM/N2969 ,\GFM/N2966 , \GFM/N2965 , \GFM/N2963 , \GFM/N2961 , \GFM/N2960 ,\GFM/N2956 , \GFM/N2955 , \GFM/N2953 , \GFM/N2952 , \GFM/N2949 ,\GFM/N2948 , \GFM/N2946 , \GFM/N2942 , \GFM/N2941 , \GFM/N2939 ,\GFM/N2938 , \GFM/N2935 , \GFM/N2934 , \GFM/N2932 , \GFM/N2930 ,\GFM/N2929 , \GFM/N2925 , \GFM/N2924 , \GFM/N2922 , \GFM/N2921 ,\GFM/N2918 , \GFM/N2917 , \GFM/N2915 , \GFM/N2911 , \GFM/N2910 ,\GFM/N2908 , \GFM/N2907 , \GFM/N2904 , \GFM/N2903 , \GFM/N2901 ,\GFM/N2899 , \GFM/N2898 , \GFM/N2894 , \GFM/N2893 , \GFM/N2891 ,\GFM/N2890 , \GFM/N2887 , \GFM/N2886 , \GFM/N2884 , \GFM/N2880 ,\GFM/N2879 , \GFM/N2877 , \GFM/N2876 , \GFM/N2873 , \GFM/N2872 ,\GFM/N2870 , \GFM/N2868 , \GFM/N2867 , \GFM/N2863 , \GFM/N2862 ,\GFM/N2860 , \GFM/N2859 , \GFM/N2856 , \GFM/N2855 , \GFM/N2853 ,\GFM/N2849 , \GFM/N2848 , \GFM/N2846 , \GFM/N2845 , \GFM/N2842 ,\GFM/N2841 , \GFM/N2839 , \GFM/N2837 , \GFM/N2836 , \GFM/N2832 ,\GFM/N2831 , \GFM/N2829 , \GFM/N2828 , \GFM/N2825 , \GFM/N2824 ,\GFM/N2822 , \GFM/N2818 , \GFM/N2817 , \GFM/N2815 , \GFM/N2814 ,\GFM/N2811 , \GFM/N2810 , \GFM/N2808 , \GFM/N2806 , \GFM/N2805 ,\GFM/N2801 , \GFM/N2800 , \GFM/N2798 , \GFM/N2797 , \GFM/N2794 ,\GFM/N2793 , \GFM/N2791 , \GFM/N2787 , \GFM/N2786 , \GFM/N2784 ,\GFM/N2783 , \GFM/N2780 , \GFM/N2779 , \GFM/N2777 , \GFM/N2775 ,\GFM/N2774 , \GFM/N2770 , \GFM/N2769 , \GFM/N2767 , \GFM/N2766 ,\GFM/N2763 , \GFM/N2762 , \GFM/N2760 , \GFM/N2756 , \GFM/N2755 ,\GFM/N2753 , \GFM/N2752 , \GFM/N2749 , \GFM/N2748 , \GFM/N2746 ,\GFM/N2744 , \GFM/N2743 , \GFM/N2739 , \GFM/N2738 , \GFM/N2736 ,\GFM/N2735 , \GFM/N2732 , \GFM/N2731 , \GFM/N2729 , \GFM/N2725 ,\GFM/N2724 , \GFM/N2722 , \GFM/N2721 , \GFM/N2718 , \GFM/N2717 ,\GFM/N2715 , \GFM/N2713 , \GFM/N2712 , \GFM/N2708 , \GFM/N2707 ,\GFM/N2705 , \GFM/N2704 , \GFM/N2701 , \GFM/N2700 , \GFM/N2698 ,\GFM/N2694 , \GFM/N2693 , \GFM/N2691 , \GFM/N2690 , \GFM/N2687 ,\GFM/N2686 , \GFM/N2684 , \GFM/N2682 , \GFM/N2681 , \GFM/N2677 ,\GFM/N2676 , \GFM/N2674 , \GFM/N2673 , \GFM/N2670 , \GFM/N2669 ,\GFM/N2667 , \GFM/N2663 , \GFM/N2662 , \GFM/N2660 , \GFM/N2659 ,\GFM/N2656 , \GFM/N2655 , \GFM/N2653 , \GFM/N2651 , \GFM/N2650 ,\GFM/N2646 , \GFM/N2645 , \GFM/N2643 , \GFM/N2642 , \GFM/N2639 ,\GFM/N2638 , \GFM/N2636 , \GFM/N2632 , \GFM/N2631 , \GFM/N2629 ,\GFM/N2628 , \GFM/N2625 , \GFM/N2624 , \GFM/N2622 , \GFM/N2620 ,\GFM/N2619 , \GFM/N2615 , \GFM/N2614 , \GFM/N2612 , \GFM/N2611 ,\GFM/N2608 , \GFM/N2607 , \GFM/N2605 , \GFM/N2601 , \GFM/N2600 ,\GFM/N2598 , \GFM/N2597 , \GFM/N2594 , \GFM/N2593 , \GFM/N2591 ,\GFM/N2589 , \GFM/N2588 , \GFM/N2584 , \GFM/N2583 , \GFM/N2581 ,\GFM/N2580 , \GFM/N2577 , \GFM/N2576 , \GFM/N2574 , \GFM/N2570 ,\GFM/N2569 , \GFM/N2567 , \GFM/N2566 , \GFM/N2563 , \GFM/N2562 ,\GFM/N2560 , \GFM/N2558 , \GFM/N2557 , \GFM/N2553 , \GFM/N2552 ,\GFM/N2550 , \GFM/N2549 , \GFM/N2546 , \GFM/N2545 , \GFM/N2543 ,\GFM/N2539 , \GFM/N2538 , \GFM/N2536 , \GFM/N2535 , \GFM/N2532 ,\GFM/N2531 , \GFM/N2529 , \GFM/N2527 , \GFM/N2526 , \GFM/N2522 ,\GFM/N2521 , \GFM/N2519 , \GFM/N2518 , \GFM/N2515 , \GFM/N2514 ,\GFM/N2512 , \GFM/N2508 , \GFM/N2507 , \GFM/N2505 , \GFM/N2504 ,\GFM/N2501 , \GFM/N2500 , \GFM/N2498 , \GFM/N2496 , \GFM/N2495 ,\GFM/N2491 , \GFM/N2490 , \GFM/N2488 , \GFM/N2487 , \GFM/N2484 ,\GFM/N2483 , \GFM/N2481 , \GFM/N2477 , \GFM/N2476 , \GFM/N2474 ,\GFM/N2473 , \GFM/N2470 , \GFM/N2469 , \GFM/N2467 , \GFM/N2465 ,\GFM/N2464 , \GFM/N2460 , \GFM/N2459 , \GFM/N2457 , \GFM/N2456 ,\GFM/N2453 , \GFM/N2452 , \GFM/N2450 , \GFM/N2446 , \GFM/N2445 ,\GFM/N2443 , \GFM/N2442 , \GFM/N2439 , \GFM/N2438 , \GFM/N2436 ,\GFM/N2434 , \GFM/N2433 , \GFM/N2429 , \GFM/N2428 , \GFM/N2426 ,\GFM/N2425 , \GFM/N2422 , \GFM/N2421 , \GFM/N2419 , \GFM/N2415 ,\GFM/N2414 , \GFM/N2412 , \GFM/N2411 , \GFM/N2408 , \GFM/N2407 ,\GFM/N2405 , \GFM/N2403 , \GFM/N2402 , \GFM/N2398 , \GFM/N2397 ,\GFM/N2395 , \GFM/N2394 , \GFM/N2391 , \GFM/N2390 , \GFM/N2388 ,\GFM/N2384 , \GFM/N2383 , \GFM/N2381 , \GFM/N2380 , \GFM/N2377 ,\GFM/N2376 , \GFM/N2374 , \GFM/N2372 , \GFM/N2371 , \GFM/N2367 ,\GFM/N2366 , \GFM/N2364 , \GFM/N2363 , \GFM/N2360 , \GFM/N2359 ,\GFM/N2357 , \GFM/N2353 , \GFM/N2352 , \GFM/N2350 , \GFM/N2349 ,\GFM/N2346 , \GFM/N2345 , \GFM/N2343 , \GFM/N2341 , \GFM/N2340 ,\GFM/N2336 , \GFM/N2335 , \GFM/N2333 , \GFM/N2332 , \GFM/N2329 ,\GFM/N2328 , \GFM/N2326 , \GFM/N2322 , \GFM/N2321 , \GFM/N2319 ,\GFM/N2318 , \GFM/N2315 , \GFM/N2314 , \GFM/N2312 , \GFM/N2310 ,\GFM/N2309 , \GFM/N2305 , \GFM/N2304 , \GFM/N2302 , \GFM/N2301 ,\GFM/N2298 , \GFM/N2297 , \GFM/N2295 , \GFM/N2291 , \GFM/N2290 ,\GFM/N2288 , \GFM/N2287 , \GFM/N2284 , \GFM/N2283 , \GFM/N2281 ,\GFM/N2279 , \GFM/N2278 , \GFM/N2274 , \GFM/N2273 , \GFM/N2271 ,\GFM/N2270 , \GFM/N2267 , \GFM/N2266 , \GFM/N2264 , \GFM/N2260 ,\GFM/N2259 , \GFM/N2257 , \GFM/N2256 , \GFM/N2253 , \GFM/N2252 ,\GFM/N2250 , \GFM/N2248 , \GFM/N2247 , \GFM/N2243 , \GFM/N2242 ,\GFM/N2240 , \GFM/N2239 , \GFM/N2236 , \GFM/N2235 , \GFM/N2233 ,\GFM/N2229 , \GFM/N2228 , \GFM/N2226 , \GFM/N2225 , \GFM/N2222 ,\GFM/N2221 , \GFM/N2219 , \GFM/N2217 , \GFM/N2216 , \GFM/N2212 ,\GFM/N2211 , \GFM/N2209 , \GFM/N2208 , \GFM/N2205 , \GFM/N2204 ,\GFM/N2202 , \GFM/N2198 , \GFM/N2197 , \GFM/N2195 , \GFM/N2194 ,\GFM/N2191 , \GFM/N2190 , \GFM/N2188 , \GFM/N2186 , \GFM/N2185 ,\GFM/N2181 , \GFM/N2180 , \GFM/N2178 , \GFM/N2177 , \GFM/N2174 ,\GFM/N2173 , \GFM/N2171 , \GFM/N2167 , \GFM/N2166 , \GFM/N2164 ,\GFM/N2163 , \GFM/N2160 , \GFM/N2159 , \GFM/N2157 , \GFM/N2155 ,\GFM/N2154 , \GFM/N2150 , \GFM/N2149 , \GFM/N2147 , \GFM/N2146 ,\GFM/N2143 , \GFM/N2142 , \GFM/N2140 , \GFM/N2136 , \GFM/N2135 ,\GFM/N2133 , \GFM/N2132 , \GFM/N2129 , \GFM/N2128 , \GFM/N2126 ,\GFM/N2124 , \GFM/N2123 , \GFM/N2119 , \GFM/N2118 , \GFM/N2116 ,\GFM/N2115 , \GFM/N2112 , \GFM/N2111 , \GFM/N2109 , \GFM/N2105 ,\GFM/N2104 , \GFM/N2102 , \GFM/N2101 , \GFM/N2098 , \GFM/N2097 ,\GFM/N2095 , \GFM/N2093 , \GFM/N2092 , \GFM/N2088 , \GFM/N2087 ,\GFM/N2085 , \GFM/N2084 , \GFM/N2081 , \GFM/N2080 , \GFM/N2078 ,\GFM/N2074 , \GFM/N2073 , \GFM/N2071 , \GFM/N2070 , \GFM/N2067 ,\GFM/N2066 , \GFM/N2064 , \GFM/N2062 , \GFM/N2061 , \GFM/N2057 ,\GFM/N2056 , \GFM/N2054 , \GFM/N2053 , \GFM/N2050 , \GFM/N2049 ,\GFM/N2047 , \GFM/N2043 , \GFM/N2042 , \GFM/N2040 , \GFM/N2039 ,\GFM/N2036 , \GFM/N2035 , \GFM/N2033 , \GFM/N2031 , \GFM/N2030 ,\GFM/N2026 , \GFM/N2025 , \GFM/N2023 , \GFM/N2022 , \GFM/N2019 ,\GFM/N2018 , \GFM/N2016 , \GFM/N2012 , \GFM/N2011 , \GFM/N2009 ,\GFM/N2008 , \GFM/N2005 , \GFM/N2004 , \GFM/N2002 , \GFM/N2000 ,\GFM/N1999 , \GFM/N1995 , \GFM/N1994 , \GFM/N1992 , \GFM/N1991 ,\GFM/N1988 , \GFM/N1987 , \GFM/N1985 , \GFM/N1981 , \GFM/N1980 ,\GFM/N1978 , \GFM/N1977 , \GFM/N1974 , \GFM/N1973 , \GFM/N1971 ,\GFM/N1969 , \GFM/N1968 , \GFM/N1964 , \GFM/N1963 , \GFM/N1961 ,\GFM/N1960 , \GFM/N1957 , \GFM/N1956 , \GFM/N1954 , \GFM/N1950 ,\GFM/N1949 , \GFM/N1947 , \GFM/N1946 , \GFM/N1943 , \GFM/N1942 ,\GFM/N1940 , \GFM/N1938 , \GFM/N1937 , \GFM/N1933 , \GFM/N1932 ,\GFM/N1930 , \GFM/N1929 , \GFM/N1926 , \GFM/N1925 , \GFM/N1923 ,\GFM/N1919 , \GFM/N1918 , \GFM/N1916 , \GFM/N1915 , \GFM/N1912 ,\GFM/N1911 , \GFM/N1909 , \GFM/N1907 , \GFM/N1906 , \GFM/N1902 ,\GFM/N1901 , \GFM/N1899 , \GFM/N1898 , \GFM/N1895 , \GFM/N1894 ,\GFM/N1892 , \GFM/N1888 , \GFM/N1887 , \GFM/N1885 , \GFM/N1884 ,\GFM/N1881 , \GFM/N1880 , \GFM/N1878 , \GFM/N1876 , \GFM/N1875 ,\GFM/N1871 , \GFM/N1870 , \GFM/N1868 , \GFM/N1867 , \GFM/N1864 ,\GFM/N1863 , \GFM/N1861 , \GFM/N1857 , \GFM/N1856 , \GFM/N1854 ,\GFM/N1853 , \GFM/N1850 , \GFM/N1849 , \GFM/N1847 , \GFM/N1845 ,\GFM/N1844 , \GFM/N1840 , \GFM/N1839 , \GFM/N1837 , \GFM/N1836 ,\GFM/N1833 , \GFM/N1832 , \GFM/N1830 , \GFM/N1826 , \GFM/N1825 ,\GFM/N1823 , \GFM/N1822 , \GFM/N1819 , \GFM/N1818 , \GFM/N1816 ,\GFM/N1814 , \GFM/N1813 , \GFM/N1809 , \GFM/N1808 , \GFM/N1806 ,\GFM/N1805 , \GFM/N1802 , \GFM/N1801 , \GFM/N1799 , \GFM/N1795 ,\GFM/N1794 , \GFM/N1792 , \GFM/N1791 , \GFM/N1788 , \GFM/N1787 ,\GFM/N1785 , \GFM/N1783 , \GFM/N1782 , \GFM/N1778 , \GFM/N1777 ,\GFM/N1775 , \GFM/N1774 , \GFM/N1771 , \GFM/N1770 , \GFM/N1768 ,\GFM/N1764 , \GFM/N1763 , \GFM/N1761 , \GFM/N1760 , \GFM/N1757 ,\GFM/N1756 , \GFM/N1754 , \GFM/N1752 , \GFM/N1751 , \GFM/N1747 ,\GFM/N1746 , \GFM/N1744 , \GFM/N1743 , \GFM/N1740 , \GFM/N1739 ,\GFM/N1737 , \GFM/N1733 , \GFM/N1732 , \GFM/N1730 , \GFM/N1729 ,\GFM/N1726 , \GFM/N1725 , \GFM/N1723 , \GFM/N1721 , \GFM/N1720 ,\GFM/N1716 , \GFM/N1715 , \GFM/N1713 , \GFM/N1712 , \GFM/N1709 ,\GFM/N1708 , \GFM/N1706 , \GFM/N1702 , \GFM/N1701 , \GFM/N1699 ,\GFM/N1698 , \GFM/N1695 , \GFM/N1694 , \GFM/N1692 , \GFM/N1690 ,\GFM/N1689 , \GFM/N1685 , \GFM/N1684 , \GFM/N1682 , \GFM/N1681 ,\GFM/N1678 , \GFM/N1677 , \GFM/N1675 , \GFM/N1671 , \GFM/N1670 ,\GFM/N1668 , \GFM/N1667 , \GFM/N1664 , \GFM/N1663 , \GFM/N1661 ,\GFM/N1659 , \GFM/N1658 , \GFM/N1654 , \GFM/N1653 , \GFM/N1651 ,\GFM/N1650 , \GFM/N1647 , \GFM/N1646 , \GFM/N1644 , \GFM/N1640 ,\GFM/N1639 , \GFM/N1637 , \GFM/N1636 , \GFM/N1633 , \GFM/N1632 ,\GFM/N1630 , \GFM/N1628 , \GFM/N1627 , \GFM/N1623 , \GFM/N1622 ,\GFM/N1620 , \GFM/N1619 , \GFM/N1616 , \GFM/N1615 , \GFM/N1613 ,\GFM/N1609 , \GFM/N1608 , \GFM/N1606 , \GFM/N1605 , \GFM/N1602 ,\GFM/N1601 , \GFM/N1599 , \GFM/N1597 , \GFM/N1596 , \GFM/N1592 ,\GFM/N1591 , \GFM/N1589 , \GFM/N1588 , \GFM/N1585 , \GFM/N1584 ,\GFM/N1582 , \GFM/N1578 , \GFM/N1577 , \GFM/N1575 , \GFM/N1574 ,\GFM/N1571 , \GFM/N1570 , \GFM/N1568 , \GFM/N1566 , \GFM/N1565 ,\GFM/N1561 , \GFM/N1560 , \GFM/N1558 , \GFM/N1557 , \GFM/N1554 ,\GFM/N1553 , \GFM/N1551 , \GFM/N1547 , \GFM/N1546 , \GFM/N1544 ,\GFM/N1543 , \GFM/N1540 , \GFM/N1539 , \GFM/N1537 , \GFM/N1535 ,\GFM/N1534 , \GFM/N1530 , \GFM/N1529 , \GFM/N1527 , \GFM/N1526 ,\GFM/N1523 , \GFM/N1522 , \GFM/N1520 , \GFM/N1516 , \GFM/N1515 ,\GFM/N1513 , \GFM/N1512 , \GFM/N1509 , \GFM/N1508 , \GFM/N1506 ,\GFM/N1504 , \GFM/N1503 , \GFM/N1499 , \GFM/N1498 , \GFM/N1496 ,\GFM/N1495 , \GFM/N1492 , \GFM/N1491 , \GFM/N1489 , \GFM/N1485 ,\GFM/N1484 , \GFM/N1482 , \GFM/N1481 , \GFM/N1478 , \GFM/N1477 ,\GFM/N1475 , \GFM/N1473 , \GFM/N1472 , \GFM/N1468 , \GFM/N1467 ,\GFM/N1465 , \GFM/N1464 , \GFM/N1461 , \GFM/N1460 , \GFM/N1458 ,\GFM/N1454 , \GFM/N1453 , \GFM/N1451 , \GFM/N1450 , \GFM/N1447 ,\GFM/N1446 , \GFM/N1444 , \GFM/N1442 , \GFM/N1441 , \GFM/N1437 ,\GFM/N1436 , \GFM/N1434 , \GFM/N1433 , \GFM/N1430 , \GFM/N1429 ,\GFM/N1427 , \GFM/N1423 , \GFM/N1422 , \GFM/N1420 , \GFM/N1419 ,\GFM/N1416 , \GFM/N1415 , \GFM/N1413 , \GFM/N1411 , \GFM/N1410 ,\GFM/N1406 , \GFM/N1405 , \GFM/N1403 , \GFM/N1402 , \GFM/N1399 ,\GFM/N1398 , \GFM/N1396 , \GFM/N1392 , \GFM/N1391 , \GFM/N1389 ,\GFM/N1388 , \GFM/N1385 , \GFM/N1384 , \GFM/N1382 , \GFM/N1380 ,\GFM/N1379 , \GFM/N1375 , \GFM/N1374 , \GFM/N1372 , \GFM/N1371 ,\GFM/N1368 , \GFM/N1367 , \GFM/N1365 , \GFM/N1361 , \GFM/N1360 ,\GFM/N1358 , \GFM/N1357 , \GFM/N1354 , \GFM/N1353 , \GFM/N1351 ,\GFM/N1349 , \GFM/N1348 , \GFM/N1344 , \GFM/N1343 , \GFM/N1341 ,\GFM/N1340 , \GFM/N1337 , \GFM/N1336 , \GFM/N1334 , \GFM/N1330 ,\GFM/N1329 , \GFM/N1327 , \GFM/N1326 , \GFM/N1323 , \GFM/N1322 ,\GFM/N1320 , \GFM/N1318 , \GFM/N1317 , \GFM/N1313 , \GFM/N1312 ,\GFM/N1310 , \GFM/N1309 , \GFM/N1306 , \GFM/N1305 , \GFM/N1303 ,\GFM/N1299 , \GFM/N1298 , \GFM/N1296 , \GFM/N1295 , \GFM/N1292 ,\GFM/N1291 , \GFM/N1289 , \GFM/N1287 , \GFM/N1286 , \GFM/N1282 ,\GFM/N1281 , \GFM/N1279 , \GFM/N1278 , \GFM/N1275 , \GFM/N1274 ,\GFM/N1272 , \GFM/N1268 , \GFM/N1267 , \GFM/N1265 , \GFM/N1264 ,\GFM/N1261 , \GFM/N1260 , \GFM/N1258 , \GFM/N1256 , \GFM/N1255 ,\GFM/N1251 , \GFM/N1250 , \GFM/N1248 , \GFM/N1247 , \GFM/N1244 ,\GFM/N1243 , \GFM/N1241 , \GFM/N1237 , \GFM/N1236 , \GFM/N1234 ,\GFM/N1233 , \GFM/N1230 , \GFM/N1229 , \GFM/N1227 , \GFM/N1225 ,\GFM/N1224 , \GFM/N1220 , \GFM/N1219 , \GFM/N1217 , \GFM/N1216 ,\GFM/N1213 , \GFM/N1212 , \GFM/N1210 , \GFM/N1206 , \GFM/N1205 ,\GFM/N1203 , \GFM/N1202 , \GFM/N1199 , \GFM/N1198 , \GFM/N1196 ,\GFM/N1194 , \GFM/N1193 , \GFM/N1189 , \GFM/N1188 , \GFM/N1186 ,\GFM/N1185 , \GFM/N1182 , \GFM/N1181 , \GFM/N1179 , \GFM/N1175 ,\GFM/N1174 , \GFM/N1172 , \GFM/N1171 , \GFM/N1168 , \GFM/N1167 ,\GFM/N1165 , \GFM/N1163 , \GFM/N1162 , \GFM/N1158 , \GFM/N1157 ,\GFM/N1155 , \GFM/N1154 , \GFM/N1151 , \GFM/N1150 , \GFM/N1148 ,\GFM/N1144 , \GFM/N1143 , \GFM/N1141 , \GFM/N1140 , \GFM/N1137 ,\GFM/N1136 , \GFM/N1134 , \GFM/N1132 , \GFM/N1131 , \GFM/N1127 ,\GFM/N1126 , \GFM/N1124 , \GFM/N1123 , \GFM/N1120 , \GFM/N1119 ,\GFM/N1117 , \GFM/N1113 , \GFM/N1112 , \GFM/N1110 , \GFM/N1109 ,\GFM/N1106 , \GFM/N1105 , \GFM/N1103 , \GFM/N1101 , \GFM/N1100 ,\GFM/N1096 , \GFM/N1095 , \GFM/N1093 , \GFM/N1092 , \GFM/N1089 ,\GFM/N1088 , \GFM/N1086 , \GFM/N1082 , \GFM/N1081 , \GFM/N1079 ,\GFM/N1078 , \GFM/N1075 , \GFM/N1074 , \GFM/N1072 , \GFM/N1070 ,\GFM/N1069 , \GFM/N1065 , \GFM/N1064 , \GFM/N1062 , \GFM/N1061 ,\GFM/N1058 , \GFM/N1057 , \GFM/N1055 , \GFM/N1051 , \GFM/N1050 ,\GFM/N1048 , \GFM/N1047 , \GFM/N1044 , \GFM/N1043 , \GFM/N1041 ,\GFM/N1039 , \GFM/N1038 , \GFM/N1034 , \GFM/N1033 , \GFM/N1031 ,\GFM/N1030 , \GFM/N1027 , \GFM/N1026 , \GFM/N1024 , \GFM/N1020 ,\GFM/N1019 , \GFM/N1017 , \GFM/N1016 , \GFM/N1013 , \GFM/N1012 ,\GFM/N1010 , \GFM/N1008 , \GFM/N1007 , \GFM/N1003 , \GFM/N1002 ,\GFM/N1000 , \GFM/N999 , \GFM/N996 , \GFM/N995 , \GFM/N993 ,\GFM/N989 , \GFM/N988 , \GFM/N986 , \GFM/N985 , \GFM/N982 ,\GFM/N981 , \GFM/N979 , \GFM/N977 , \GFM/N976 , \GFM/N972 ,\GFM/N971 , \GFM/N969 , \GFM/N968 , \GFM/N965 , \GFM/N964 ,\GFM/N962 , \GFM/N958 , \GFM/N957 , \GFM/N955 , \GFM/N954 ,\GFM/N951 , \GFM/N950 , \GFM/N948 , \GFM/N946 , \GFM/N945 ,\GFM/N941 , \GFM/N940 , \GFM/N938 , \GFM/N937 , \GFM/N934 ,\GFM/N933 , \GFM/N931 , \GFM/N927 , \GFM/N926 , \GFM/N924 ,\GFM/N923 , \GFM/N920 , \GFM/N919 , \GFM/N917 , \GFM/N915 ,\GFM/N914 , \GFM/N910 , \GFM/N909 , \GFM/N907 , \GFM/N906 ,\GFM/N903 , \GFM/N902 , \GFM/N900 , \GFM/N896 , \GFM/N895 ,\GFM/N893 , \GFM/N892 , \GFM/N889 , \GFM/N888 , \GFM/N886 ,\GFM/N884 , \GFM/N883 , \GFM/N879 , \GFM/N878 , \GFM/N876 ,\GFM/N875 , \GFM/N872 , \GFM/N871 , \GFM/N869 , \GFM/N865 ,\GFM/N864 , \GFM/N862 , \GFM/N861 , \GFM/N858 , \GFM/N857 ,\GFM/N855 , \GFM/N853 , \GFM/N852 , \GFM/N848 , \GFM/N847 ,\GFM/N845 , \GFM/N844 , \GFM/N841 , \GFM/N840 , \GFM/N838 ,\GFM/N834 , \GFM/N833 , \GFM/N831 , \GFM/N830 , \GFM/N827 ,\GFM/N826 , \GFM/N824 , \GFM/N822 , \GFM/N821 , \GFM/N817 ,\GFM/N816 , \GFM/N814 , \GFM/N813 , \GFM/N810 , \GFM/N809 ,\GFM/N807 , \GFM/N803 , \GFM/N802 , \GFM/N800 , \GFM/N799 ,\GFM/N796 , \GFM/N795 , \GFM/N793 , \GFM/N791 , \GFM/N790 ,\GFM/N786 , \GFM/N785 , \GFM/N783 , \GFM/N782 , \GFM/N779 ,\GFM/N778 , \GFM/N776 , \GFM/N772 , \GFM/N771 , \GFM/N769 ,\GFM/N768 , \GFM/N765 , \GFM/N764 , \GFM/N762 , \GFM/N760 ,\GFM/N759 , \GFM/N755 , \GFM/N754 , \GFM/N752 , \GFM/N751 ,\GFM/N748 , \GFM/N747 , \GFM/N745 , \GFM/N741 , \GFM/N740 ,\GFM/N738 , \GFM/N737 , \GFM/N734 , \GFM/N733 , \GFM/N731 ,\GFM/N729 , \GFM/N728 , \GFM/N724 , \GFM/N723 , \GFM/N721 ,\GFM/N720 , \GFM/N717 , \GFM/N716 , \GFM/N714 , \GFM/N710 ,\GFM/N709 , \GFM/N707 , \GFM/N706 , \GFM/N703 , \GFM/N702 ,\GFM/N700 , \GFM/N698 , \GFM/N697 , \GFM/N693 , \GFM/N692 ,\GFM/N690 , \GFM/N689 , \GFM/N686 , \GFM/N685 , \GFM/N683 ,\GFM/N679 , \GFM/N678 , \GFM/N676 , \GFM/N675 , \GFM/N672 ,\GFM/N671 , \GFM/N669 , \GFM/N667 , \GFM/N666 , \GFM/N662 ,\GFM/N661 , \GFM/N659 , \GFM/N658 , \GFM/N655 , \GFM/N654 ,\GFM/N652 , \GFM/N648 , \GFM/N647 , \GFM/N645 , \GFM/N644 ,\GFM/N641 , \GFM/N640 , \GFM/N638 , \GFM/N636 , \GFM/N635 ,\GFM/N631 , \GFM/N630 , \GFM/N628 , \GFM/N627 , \GFM/N624 ,\GFM/N623 , \GFM/N621 , \GFM/N617 , \GFM/N616 , \GFM/N614 ,\GFM/N613 , \GFM/N610 , \GFM/N609 , \GFM/N607 , \GFM/N605 ,\GFM/N604 , \GFM/N600 , \GFM/N599 , \GFM/N597 , \GFM/N596 ,\GFM/N593 , \GFM/N592 , \GFM/N590 , \GFM/N586 , \GFM/N585 ,\GFM/N583 , \GFM/N582 , \GFM/N579 , \GFM/N578 , \GFM/N576 ,\GFM/N574 , \GFM/N573 , \GFM/N569 , \GFM/N568 , \GFM/N566 ,\GFM/N565 , \GFM/N562 , \GFM/N561 , \GFM/N559 , \GFM/N555 ,\GFM/N554 , \GFM/N552 , \GFM/N551 , \GFM/N548 , \GFM/N547 ,\GFM/N545 , \GFM/N543 , \GFM/N542 , \GFM/N538 , \GFM/N537 ,\GFM/N535 , \GFM/N534 , \GFM/N531 , \GFM/N530 , \GFM/N528 ,\GFM/N524 , \GFM/N523 , \GFM/N521 , \GFM/N520 , \GFM/N517 ,\GFM/N516 , \GFM/N514 , \GFM/N512 , \GFM/N511 , \GFM/N507 ,\GFM/N506 , \GFM/N504 , \GFM/N503 , \GFM/N500 , \GFM/N499 ,\GFM/N497 , \GFM/N493 , \GFM/N492 , \GFM/N490 , \GFM/N489 ,\GFM/N486 , \GFM/N485 , \GFM/N483 , \GFM/N481 , \GFM/N480 ,\GFM/N476 , \GFM/N475 , \GFM/N473 , \GFM/N472 , \GFM/N469 ,\GFM/N468 , \GFM/N466 , \GFM/N462 , \GFM/N461 , \GFM/N459 ,\GFM/N458 , \GFM/N455 , \GFM/N454 , \GFM/N452 , \GFM/N450 ,\GFM/N449 , \GFM/N445 , \GFM/N444 , \GFM/N442 , \GFM/N441 ,\GFM/N438 , \GFM/N437 , \GFM/N435 , \GFM/N431 , \GFM/N430 ,\GFM/N428 , \GFM/N427 , \GFM/N424 , \GFM/N423 , \GFM/N421 ,\GFM/N419 , \GFM/N418 , \GFM/N414 , \GFM/N413 , \GFM/N411 ,\GFM/N410 , \GFM/N407 , \GFM/N406 , \GFM/N404 , \GFM/N400 ,\GFM/N399 , \GFM/N397 , \GFM/N396 , \GFM/N393 , \GFM/N392 ,\GFM/N390 , \GFM/N388 , \GFM/N387 , \GFM/N383 , \GFM/N382 ,\GFM/N380 , \GFM/N379 , \GFM/N376 , \GFM/N375 , \GFM/N373 ,\GFM/N369 , \GFM/N368 , \GFM/N366 , \GFM/N365 , \GFM/N362 ,\GFM/N361 , \GFM/N359 , \GFM/N357 , \GFM/N356 , \GFM/N352 ,\GFM/N351 , \GFM/N349 , \GFM/N348 , \GFM/N345 , \GFM/N344 ,\GFM/N342 , \GFM/N338 , \GFM/N337 , \GFM/N335 , \GFM/N334 ,\GFM/N331 , \GFM/N330 , \GFM/N328 , \GFM/N326 , \GFM/N325 ,\GFM/N321 , \GFM/N320 , \GFM/N318 , \GFM/N317 , \GFM/N314 ,\GFM/N313 , \GFM/N311 , \GFM/N307 , \GFM/N306 , \GFM/N304 ,\GFM/N303 , \GFM/N300 , \GFM/N299 , \GFM/N297 , \GFM/N295 ,\GFM/N294 , \GFM/N290 , \GFM/N289 , \GFM/N287 , \GFM/N286 ,\GFM/N283 , \GFM/N282 , \GFM/N280 , \GFM/N276 , \GFM/N275 ,\GFM/N273 , \GFM/N272 , \GFM/N269 , \GFM/N268 , \GFM/N266 ,\GFM/N264 , \GFM/N263 , \GFM/N259 , \GFM/N258 , \GFM/N256 ,\GFM/N255 , \GFM/N252 , \GFM/N251 , \GFM/N249 , \GFM/N245 ,\GFM/N244 , \GFM/N242 , \GFM/N241 , \GFM/N238 , \GFM/N237 ,\GFM/N235 , \GFM/N233 , \GFM/N232 , \GFM/N228 , \GFM/N227 ,\GFM/N225 , \GFM/N224 , \GFM/N221 , \GFM/N220 , \GFM/N218 ,\GFM/N214 , \GFM/N213 , \GFM/N211 , \GFM/N210 , \GFM/N207 ,\GFM/N206 , \GFM/N204 , \GFM/N202 , \GFM/N201 , \GFM/N197 ,\GFM/N196 , \GFM/N194 , \GFM/N193 , \GFM/N190 , \GFM/N189 ,\GFM/N187 , \GFM/N183 , \GFM/N182 , \GFM/N180 , \GFM/N179 ,\GFM/N176 , \GFM/N175 , \GFM/N173 , \GFM/N171 , \GFM/N170 ,\GFM/N166 , \GFM/N165 , \GFM/N163 , \GFM/N162 , \GFM/N159 ,\GFM/N158 , \GFM/N156 , \GFM/N152 , \GFM/N151 , \GFM/N149 ,\GFM/N148 , \GFM/N145 , \GFM/N144 , \GFM/N142 , \GFM/N140 ,\GFM/N139 , \GFM/N135 , \GFM/N134 , \GFM/N132 , \GFM/N131 ,\GFM/N128 , \GFM/N127 , \GFM/N125 , \GFM/N121 , \GFM/N120 ,\GFM/N118 , \GFM/N117 , \GFM/N114 , \GFM/N113 , \GFM/N111 ,\GFM/N109 , \GFM/N108 , \GFM/N104 , \GFM/N103 , \GFM/N101 ,\GFM/N100 , \GFM/N97 , \GFM/N96 , \GFM/N94 , \GFM/N90 , \GFM/N89 ,\GFM/N87 , \GFM/N86 , \GFM/N83 , \GFM/N82 , \GFM/N80 , \GFM/N78 ,\GFM/N77 , \GFM/N73 , \GFM/N72 , \GFM/N70 , \GFM/N69 , \GFM/N66 ,\GFM/N65 , \GFM/N63 , \GFM/N59 , \GFM/N58 , \GFM/N56 , \GFM/N55 ,\GFM/N52 , \GFM/N51 , \GFM/N49 , \GFM/N47 , \GFM/N46 , \GFM/N42 ,\GFM/N41 , \GFM/N39 , \GFM/N38 , \GFM/N35 , \GFM/N34 , \GFM/N32 ,\GFM/N28 , \GFM/N27 , \GFM/N25 , \GFM/N24 , \GFM/N21 , \GFM/N20 ,\GFM/N18 , \GFM/N16 , \GFM/N15 , \GFM/N11 , \GFM/N10 , \GFM/N8 ,\GFM/N7 , \GFM/N4 , \GFM/N3 , \GFM/N1 , \AES_ENC/n1267 ,\AES_ENC/n1266 , \AES_ENC/n1265 , \AES_ENC/n1264 , \AES_ENC/n1263 ,\AES_ENC/n1262 , \AES_ENC/n1261 , \AES_ENC/n12601 , \AES_ENC/n1259 ,\AES_ENC/n1258 , \AES_ENC/n1257 , \AES_ENC/n1256 , \AES_ENC/n1255 ,\AES_ENC/n1254 , \AES_ENC/n1253 , \AES_ENC/n1252 , \AES_ENC/n1251 ,\AES_ENC/n1250 , \AES_ENC/n1249 , \AES_ENC/n1248 , \AES_ENC/n1247 ,\AES_ENC/n1246 , \AES_ENC/n1245 , \AES_ENC/n1244 , \AES_ENC/n1243 ,\AES_ENC/n1242 , \AES_ENC/n1241 , \AES_ENC/n1240 , \AES_ENC/n1239 ,\AES_ENC/n1238 , \AES_ENC/n1237 , \AES_ENC/n1236 , \AES_ENC/n1235 ,\AES_ENC/n1234 , \AES_ENC/n1233 , \AES_ENC/n1232 , \AES_ENC/n1231 ,\AES_ENC/n793 , \AES_ENC/n794 , \AES_ENC/n792 , \AES_ENC/n791 ,\AES_ENC/n7901 , \AES_ENC/n7891 , \AES_ENC/n6601 , \AES_ENC/n659 ,\AES_ENC/n658 , \AES_ENC/n657 , \AES_ENC/n656 , \AES_ENC/n655 ,\AES_ENC/n654 , \AES_ENC/n653 , \AES_ENC/n652 , \AES_ENC/n651 ,\AES_ENC/n6501 , \AES_ENC/n649 , \AES_ENC/n648 , \AES_ENC/n647 ,\AES_ENC/n646 , \AES_ENC/n645 , \AES_ENC/n644 , \AES_ENC/n643 ,\AES_ENC/n642 , \AES_ENC/n641 , \AES_ENC/n6401 , \AES_ENC/n639 ,\AES_ENC/n638 , \AES_ENC/n637 , \AES_ENC/n636 , \AES_ENC/n635 ,\AES_ENC/n634 , \AES_ENC/n633 , \AES_ENC/n632 , \AES_ENC/n631 ,\AES_ENC/n6301 , \AES_ENC/n629 , \AES_ENC/n628 , \AES_ENC/n627 ,\AES_ENC/n626 , \AES_ENC/n625 , \AES_ENC/n624 , \AES_ENC/n623 ,\AES_ENC/n622 , \AES_ENC/n621 , \AES_ENC/n6201 , \AES_ENC/n619 ,\AES_ENC/n618 , \AES_ENC/n617 , \AES_ENC/n616 , \AES_ENC/n615 ,\AES_ENC/n614 , \AES_ENC/n613 , \AES_ENC/n612 , \AES_ENC/n611 ,\AES_ENC/n610 , \AES_ENC/n609 , \AES_ENC/n608 , \AES_ENC/n607 ,\AES_ENC/n606 , \AES_ENC/n605 , \AES_ENC/n604 , \AES_ENC/n603 ,\AES_ENC/n602 , \AES_ENC/n601 , \AES_ENC/n600 , \AES_ENC/n599 ,\AES_ENC/n598 , \AES_ENC/n597 , \AES_ENC/n596 , \AES_ENC/n595 ,\AES_ENC/n594 , \AES_ENC/n593 , \AES_ENC/n592 , \AES_ENC/n591 ,\AES_ENC/n590 , \AES_ENC/n589 , \AES_ENC/n588 , \AES_ENC/n587 ,\AES_ENC/n586 , \AES_ENC/n585 , \AES_ENC/n584 , \AES_ENC/n583 ,\AES_ENC/n582 , \AES_ENC/n581 , \AES_ENC/n580 , \AES_ENC/n579 ,\AES_ENC/n578 , \AES_ENC/n577 , \AES_ENC/n576 , \AES_ENC/n575 ,\AES_ENC/n574 , \AES_ENC/n573 , \AES_ENC/n572 , \AES_ENC/n571 ,\AES_ENC/n570 , \AES_ENC/n569 , \AES_ENC/n568 , \AES_ENC/n567 ,\AES_ENC/n566 , \AES_ENC/n565 , \AES_ENC/n564 , \AES_ENC/n563 ,\AES_ENC/n562 , \AES_ENC/n561 , \AES_ENC/n560 , \AES_ENC/n559 ,\AES_ENC/n558 , \AES_ENC/n557 , \AES_ENC/n556 , \AES_ENC/n555 ,\AES_ENC/n554 , \AES_ENC/n553 , \AES_ENC/n552 , \AES_ENC/n551 ,\AES_ENC/n550 , \AES_ENC/n549 , \AES_ENC/n548 , \AES_ENC/n547 ,\AES_ENC/n546 , \AES_ENC/n545 , \AES_ENC/n544 , \AES_ENC/n543 ,\AES_ENC/n542 , \AES_ENC/n541 , \AES_ENC/n540 , \AES_ENC/n539 ,\AES_ENC/n538 , \AES_ENC/n537 , \AES_ENC/n536 , \AES_ENC/n535 ,\AES_ENC/n534 , \AES_ENC/n533 , \AES_ENC/n532 , \AES_ENC/n531 ,\AES_ENC/n5301 , \AES_ENC/n529 , \AES_ENC/n528 , \AES_ENC/n527 ,\AES_ENC/n526 , \AES_ENC/n525 , \AES_ENC/n524 , \AES_ENC/n523 ,\AES_ENC/n522 , \AES_ENC/n521 , \AES_ENC/n5201 , \AES_ENC/n519 ,\AES_ENC/n518 , \AES_ENC/n517 , \AES_ENC/n516 , \AES_ENC/n515 ,\AES_ENC/n514 , \AES_ENC/n513 , \AES_ENC/n512 , \AES_ENC/n511 ,\AES_ENC/n5101 , \AES_ENC/n509 , \AES_ENC/n508 , \AES_ENC/n507 ,\AES_ENC/n506 , \AES_ENC/n505 , \AES_ENC/n504 , \AES_ENC/n503 ,\AES_ENC/n5021 , \AES_ENC/n5010 , \AES_ENC/n5000 , \AES_ENC/n4990 ,\AES_ENC/n4980 , \AES_ENC/n4970 , \AES_ENC/n4960 , \AES_ENC/n4950 ,\AES_ENC/n4940 , \AES_ENC/n4930 , \AES_ENC/n4920 , \AES_ENC/n4911 ,\AES_ENC/n4900 , \AES_ENC/n4890 , \AES_ENC/n4880 , \AES_ENC/n4870 ,\AES_ENC/n4860 , \AES_ENC/n4850 , \AES_ENC/n4840 , \AES_ENC/n4830 ,\AES_ENC/n4820 , \AES_ENC/n4811 , \AES_ENC/n4800 , \AES_ENC/n4790 ,\AES_ENC/n4780 , \AES_ENC/n4770 , \AES_ENC/n4760 , \AES_ENC/n4750 ,\AES_ENC/n4740 , \AES_ENC/n4730 , \AES_ENC/n4720 , \AES_ENC/n4711 ,\AES_ENC/n4700 , \AES_ENC/n4690 , \AES_ENC/n4680 , \AES_ENC/n4670 ,\AES_ENC/n4660 , \AES_ENC/n4650 , \AES_ENC/n4640 , \AES_ENC/n4630 ,\AES_ENC/n4620 , \AES_ENC/n4611 , \AES_ENC/n4600 , \AES_ENC/n4590 ,\AES_ENC/n4580 , \AES_ENC/n4570 , \AES_ENC/n4560 , \AES_ENC/n4550 ,\AES_ENC/n4540 , \AES_ENC/n4530 , \AES_ENC/n4520 , \AES_ENC/n4510 ,\AES_ENC/n4500 , \AES_ENC/n4490 , \AES_ENC/n4480 , \AES_ENC/n4470 ,\AES_ENC/n4460 , \AES_ENC/n4450 , \AES_ENC/n4440 , \AES_ENC/n4430 ,\AES_ENC/n4420 , \AES_ENC/n4410 , \AES_ENC/n4400 , \AES_ENC/n4390 ,\AES_ENC/n4380 , \AES_ENC/n4370 , \AES_ENC/n4360 , \AES_ENC/n4350 ,\AES_ENC/n4340 , \AES_ENC/n4330 , \AES_ENC/n4320 , \AES_ENC/n4310 ,\AES_ENC/n4300 , \AES_ENC/n4290 , \AES_ENC/n4280 , \AES_ENC/n4270 ,\AES_ENC/n4260 , \AES_ENC/n4250 , \AES_ENC/n4240 , \AES_ENC/n4230 ,\AES_ENC/n4220 , \AES_ENC/n4210 , \AES_ENC/n4200 , \AES_ENC/n4190 ,\AES_ENC/n4180 , \AES_ENC/n4170 , \AES_ENC/n4160 , \AES_ENC/n4150 ,\AES_ENC/n4140 , \AES_ENC/n4130 , \AES_ENC/n4120 , \AES_ENC/n4110 ,\AES_ENC/n4100 , \AES_ENC/n4090 , \AES_ENC/n4080 , \AES_ENC/n4070 ,\AES_ENC/n4060 , \AES_ENC/n4050 , \AES_ENC/n4040 , \AES_ENC/n4030 ,\AES_ENC/n4020 , \AES_ENC/n4010 , \AES_ENC/n4000 , \AES_ENC/n3990 ,\AES_ENC/n3980 , \AES_ENC/n3970 , \AES_ENC/n3960 , \AES_ENC/n3950 ,\AES_ENC/n3940 , \AES_ENC/n3930 , \AES_ENC/n3920 , \AES_ENC/n3910 ,\AES_ENC/n3900 , \AES_ENC/n3890 , \AES_ENC/n3880 , \AES_ENC/n3870 ,\AES_ENC/n3860 , \AES_ENC/n3850 , \AES_ENC/n3840 , \AES_ENC/n3830 ,\AES_ENC/n3820 , \AES_ENC/n3810 , \AES_ENC/n3800 , \AES_ENC/n3790 ,\AES_ENC/n3780 , \AES_ENC/n3770 , \AES_ENC/n3760 , \AES_ENC/n3750 ,\AES_ENC/n3740 , \AES_ENC/n373 , \AES_ENC/n372 , \AES_ENC/n371 ,\AES_ENC/n3701 , \AES_ENC/n369 , \AES_ENC/n368 , \AES_ENC/n367 ,\AES_ENC/n366 , \AES_ENC/n365 , \AES_ENC/n364 , \AES_ENC/n363 ,\AES_ENC/n362 , \AES_ENC/n361 , \AES_ENC/n3601 , \AES_ENC/n359 ,\AES_ENC/n358 , \AES_ENC/n357 , \AES_ENC/n356 , \AES_ENC/n355 ,\AES_ENC/n354 , \AES_ENC/n353 , \AES_ENC/n352 , \AES_ENC/n351 ,\AES_ENC/n3501 , \AES_ENC/n349 , \AES_ENC/n348 , \AES_ENC/n347 ,\AES_ENC/n346 , \AES_ENC/n345 , \AES_ENC/n344 , \AES_ENC/n343 ,\AES_ENC/n342 , \AES_ENC/n341 , \AES_ENC/n3401 , \AES_ENC/n339 ,\AES_ENC/n338 , \AES_ENC/n337 , \AES_ENC/n336 , \AES_ENC/n335 ,\AES_ENC/n334 , \AES_ENC/n333 , \AES_ENC/n332 , \AES_ENC/n331 ,\AES_ENC/n3301 , \AES_ENC/n329 , \AES_ENC/n328 , \AES_ENC/n327 ,\AES_ENC/n326 , \AES_ENC/n325 , \AES_ENC/n324 , \AES_ENC/n323 ,\AES_ENC/n322 , \AES_ENC/n321 , \AES_ENC/n3201 , \AES_ENC/n319 ,\AES_ENC/n318 , \AES_ENC/n317 , \AES_ENC/n316 , \AES_ENC/n315 ,\AES_ENC/n314 , \AES_ENC/n313 , \AES_ENC/n312 , \AES_ENC/n311 ,\AES_ENC/n3101 , \AES_ENC/n309 , \AES_ENC/n308 , \AES_ENC/n307 ,\AES_ENC/n306 , \AES_ENC/n305 , \AES_ENC/n304 , \AES_ENC/n303 ,\AES_ENC/n302 , \AES_ENC/n301 , \AES_ENC/n3001 , \AES_ENC/n299 ,\AES_ENC/n298 , \AES_ENC/n297 , \AES_ENC/n296 , \AES_ENC/n295 ,\AES_ENC/n294 , \AES_ENC/n293 , \AES_ENC/n292 , \AES_ENC/n291 ,\AES_ENC/n290 , \AES_ENC/n289 , \AES_ENC/n288 , \AES_ENC/n287 ,\AES_ENC/n286 , \AES_ENC/n285 , \AES_ENC/n284 , \AES_ENC/n283 ,\AES_ENC/n282 , \AES_ENC/n281 , \AES_ENC/n280 , \AES_ENC/n279 ,\AES_ENC/n278 , \AES_ENC/n2770 , \AES_ENC/n2760 , \AES_ENC/n2750 ,\AES_ENC/n2740 , \AES_ENC/n2730 , \AES_ENC/n2720 , \AES_ENC/n2710 ,\AES_ENC/n2700 , \AES_ENC/n269 , \AES_ENC/n268 , \AES_ENC/n267 ,\AES_ENC/n266 , \AES_ENC/n265 , \AES_ENC/n264 , \AES_ENC/n263 ,\AES_ENC/n262 , \AES_ENC/n2610 , \AES_ENC/n2600 , \AES_ENC/n2590 ,\AES_ENC/n2580 , \AES_ENC/n2570 , \AES_ENC/n2560 , \AES_ENC/n2550 ,\AES_ENC/n2540 , \AES_ENC/n253 , \AES_ENC/n252 , \AES_ENC/n251 ,\AES_ENC/n250 , \AES_ENC/n249 , \AES_ENC/n248 , \AES_ENC/n247 ,\AES_ENC/n246 , \AES_ENC/n2450 , \AES_ENC/n2440 , \AES_ENC/n2430 ,\AES_ENC/n2420 , \AES_ENC/n2410 , \AES_ENC/n2400 , \AES_ENC/n2390 ,\AES_ENC/n2380 , \AES_ENC/n237 , \AES_ENC/n236 , \AES_ENC/n235 ,\AES_ENC/n234 , \AES_ENC/n233 , \AES_ENC/n232 , \AES_ENC/n231 ,\AES_ENC/n230 , \AES_ENC/n2290 , \AES_ENC/n2280 , \AES_ENC/n2270 ,\AES_ENC/n2260 , \AES_ENC/n2250 , \AES_ENC/n2240 , \AES_ENC/n2230 ,\AES_ENC/n2220 , \AES_ENC/n221 , \AES_ENC/n220 , \AES_ENC/n219 ,\AES_ENC/n218 , \AES_ENC/n217 , \AES_ENC/n216 , \AES_ENC/n215 ,\AES_ENC/n214 , \AES_ENC/n2130 , \AES_ENC/n2120 , \AES_ENC/n2110 ,\AES_ENC/n2100 , \AES_ENC/n2090 , \AES_ENC/n2080 , \AES_ENC/n2070 ,\AES_ENC/n2060 , \AES_ENC/n205 , \AES_ENC/n204 , \AES_ENC/n203 ,\AES_ENC/n202 , \AES_ENC/n201 , \AES_ENC/n200 , \AES_ENC/n199 ,\AES_ENC/n1981 , \AES_ENC/n1970 , \AES_ENC/n1960 , \AES_ENC/n1950 ,\AES_ENC/n1940 , \AES_ENC/n1930 , \AES_ENC/n1920 , \AES_ENC/n1910 ,\AES_ENC/n1900 , \AES_ENC/n189 , \AES_ENC/n188 , \AES_ENC/n187 ,\AES_ENC/n186 , \AES_ENC/n185 , \AES_ENC/n184 , \AES_ENC/n183 ,\AES_ENC/n182 , \AES_ENC/n1810 , \AES_ENC/n1800 , \AES_ENC/n1790 ,\AES_ENC/n1780 , \AES_ENC/n1770 , \AES_ENC/n1760 , \AES_ENC/n1750 ,\AES_ENC/n1740 , \AES_ENC/n173 , \AES_ENC/n172 , \AES_ENC/n171 ,\AES_ENC/n170 , \AES_ENC/n169 , \AES_ENC/n168 , \AES_ENC/n167 ,\AES_ENC/n166 , \AES_ENC/n1650 , \AES_ENC/n1640 , \AES_ENC/n1630 ,\AES_ENC/n1620 , \AES_ENC/n1610 , \AES_ENC/n1600 , \AES_ENC/n1590 ,\AES_ENC/n1580 , \AES_ENC/n157 , \AES_ENC/n156 , \AES_ENC/n155 ,\AES_ENC/n154 , \AES_ENC/n153 , \AES_ENC/n152 , \AES_ENC/n151 ,\AES_ENC/n150 , \AES_ENC/n1490 , \AES_ENC/n1480 , \AES_ENC/n1470 ,\AES_ENC/n1460 , \AES_ENC/n1450 , \AES_ENC/n1440 , \AES_ENC/n1430 ,\AES_ENC/n1420 , \AES_ENC/n141 , \AES_ENC/n140 , \AES_ENC/n139 ,\AES_ENC/n138 , \AES_ENC/n137 , \AES_ENC/n136 , \AES_ENC/n135 ,\AES_ENC/n134 , \AES_ENC/n1330 , \AES_ENC/n1320 , \AES_ENC/n1310 ,\AES_ENC/n1300 , \AES_ENC/n1290 , \AES_ENC/n1280 , \AES_ENC/n1270 ,\AES_ENC/n12600 , \AES_ENC/n125 , \AES_ENC/n124 , \AES_ENC/n123 ,\AES_ENC/n122 , \AES_ENC/n121 , \AES_ENC/n120 , \AES_ENC/n119 ,\AES_ENC/n118 , \AES_ENC/n11710 , \AES_ENC/n11610 , \AES_ENC/n11510 ,\AES_ENC/n11410 , \AES_ENC/n11310 , \AES_ENC/n11210 ,\AES_ENC/n11110 , \AES_ENC/n11010 , \AES_ENC/n109 , \AES_ENC/n108 ,\AES_ENC/n107 , \AES_ENC/n106 , \AES_ENC/n105 , \AES_ENC/n104 ,\AES_ENC/n103 , \AES_ENC/n102 , \AES_ENC/n10110 , \AES_ENC/n10010 ,\AES_ENC/n9910 , \AES_ENC/n9810 , \AES_ENC/n9710 , \AES_ENC/n9610 ,\AES_ENC/n9510 , \AES_ENC/n9410 , \AES_ENC/n93 , \AES_ENC/n92 ,\AES_ENC/n91 , \AES_ENC/n90 , \AES_ENC/n89 , \AES_ENC/n88 ,\AES_ENC/n87 , \AES_ENC/n86 , \AES_ENC/n8510 , \AES_ENC/n8410 ,\AES_ENC/n8310 , \AES_ENC/n8210 , \AES_ENC/n8110 , \AES_ENC/n8010 ,\AES_ENC/n7900 , \AES_ENC/n7890 , \AES_ENC/n77 , \AES_ENC/n76 ,\AES_ENC/n75 , \AES_ENC/n74 , \AES_ENC/n73 , \AES_ENC/n72 ,\AES_ENC/n71 , \AES_ENC/n70 , \AES_ENC/n6910 , \AES_ENC/n6810 ,\AES_ENC/n6710 , \AES_ENC/n6600 , \AES_ENC/n6500 , \AES_ENC/n6400 ,\AES_ENC/n6300 , \AES_ENC/n6200 , \AES_ENC/n61 , \AES_ENC/n60 ,\AES_ENC/n59 , \AES_ENC/n58 , \AES_ENC/n57 , \AES_ENC/n56 ,\AES_ENC/n55 , \AES_ENC/n54 , \AES_ENC/n5300 , \AES_ENC/n5200 ,\AES_ENC/n5100 , \AES_ENC/n5020 , \AES_ENC/n4910 , \AES_ENC/n4810 ,\AES_ENC/n4710 , \AES_ENC/n4610 , \AES_ENC/n45 , \AES_ENC/n44 ,\AES_ENC/n43 , \AES_ENC/n42 , \AES_ENC/n41 , \AES_ENC/n40 ,\AES_ENC/n39 , \AES_ENC/n38 , \AES_ENC/n3700 , \AES_ENC/n3600 ,\AES_ENC/n3500 , \AES_ENC/n3400 , \AES_ENC/n3300 , \AES_ENC/n3200 ,\AES_ENC/n3100 , \AES_ENC/n3000 , \AES_ENC/n29 , \AES_ENC/n28 ,\AES_ENC/n27 , \AES_ENC/n26 , \AES_ENC/n25 , \AES_ENC/n24 ,\AES_ENC/n23 , \AES_ENC/n22 , \AES_ENC/n21 , \AES_ENC/n20 ,\AES_ENC/n1980 , \AES_ENC/n18 , \AES_ENC/n17 , \AES_ENC/n16 ,\AES_ENC/n15 , \AES_ENC/n14 , \AES_ENC/n13 , \AES_ENC/n12 ,\AES_ENC/n11 , \AES_ENC/n2 , \AES_ENC/n1230 , \AES_ENC/n1229 ,\AES_ENC/n1228 , \AES_ENC/n1227 , \AES_ENC/n1226 , \AES_ENC/n1225 ,\AES_ENC/n1224 , \AES_ENC/n1223 , \AES_ENC/n1222 , \AES_ENC/n1221 ,\AES_ENC/n1220 , \AES_ENC/n1219 , \AES_ENC/n1218 , \AES_ENC/n1217 ,\AES_ENC/n1216 , \AES_ENC/n1215 , \AES_ENC/n1214 , \AES_ENC/n1213 ,\AES_ENC/n1212 , \AES_ENC/n1211 , \AES_ENC/n1210 , \AES_ENC/n1209 ,\AES_ENC/n1208 , \AES_ENC/n1207 , \AES_ENC/n1206 , \AES_ENC/n1205 ,\AES_ENC/n1204 , \AES_ENC/n1203 , \AES_ENC/n1202 , \AES_ENC/n1201 ,\AES_ENC/n1200 , \AES_ENC/n1199 , \AES_ENC/n1198 , \AES_ENC/n1197 ,\AES_ENC/n1196 , \AES_ENC/n1195 , \AES_ENC/n1194 , \AES_ENC/n1193 ,\AES_ENC/n1192 , \AES_ENC/n1191 , \AES_ENC/n1190 , \AES_ENC/n1189 ,\AES_ENC/n1188 , \AES_ENC/n1187 , \AES_ENC/n1186 , \AES_ENC/n1185 ,\AES_ENC/n1184 , \AES_ENC/n1183 , \AES_ENC/n1182 , \AES_ENC/n1181 ,\AES_ENC/n1180 , \AES_ENC/n1179 , \AES_ENC/n1178 , \AES_ENC/n1177 ,\AES_ENC/n1176 , \AES_ENC/n1175 , \AES_ENC/n1174 , \AES_ENC/n1173 ,\AES_ENC/n1172 , \AES_ENC/n1171 , \AES_ENC/n1170 , \AES_ENC/n1169 ,\AES_ENC/n1168 , \AES_ENC/n1167 , \AES_ENC/n1166 , \AES_ENC/n1165 ,\AES_ENC/n1164 , \AES_ENC/n1163 , \AES_ENC/n1162 , \AES_ENC/n1161 ,\AES_ENC/n1160 , \AES_ENC/n1159 , \AES_ENC/n1158 , \AES_ENC/n1157 ,\AES_ENC/n1156 , \AES_ENC/n1155 , \AES_ENC/n1154 , \AES_ENC/n1153 ,\AES_ENC/n1152 , \AES_ENC/n1151 , \AES_ENC/n1150 , \AES_ENC/n1149 ,\AES_ENC/n1148 , \AES_ENC/n1147 , \AES_ENC/n1146 , \AES_ENC/n1145 ,\AES_ENC/n1144 , \AES_ENC/n1143 , \AES_ENC/n1142 , \AES_ENC/n1141 ,\AES_ENC/n1140 , \AES_ENC/n1139 , \AES_ENC/n1138 , \AES_ENC/n1137 ,\AES_ENC/n1136 , \AES_ENC/n1135 , \AES_ENC/n1134 , \AES_ENC/n1133 ,\AES_ENC/n1132 , \AES_ENC/n1131 , \AES_ENC/n1130 , \AES_ENC/n1129 ,\AES_ENC/n1128 , \AES_ENC/n1127 , \AES_ENC/n1126 , \AES_ENC/n1125 ,\AES_ENC/n1124 , \AES_ENC/n1123 , \AES_ENC/n1122 , \AES_ENC/n1121 ,\AES_ENC/n1120 , \AES_ENC/n1119 , \AES_ENC/n1118 , \AES_ENC/n1117 ,\AES_ENC/n1116 , \AES_ENC/n1115 , \AES_ENC/n1114 , \AES_ENC/n1113 ,\AES_ENC/n1112 , \AES_ENC/n1111 , \AES_ENC/n1110 , \AES_ENC/n1109 ,\AES_ENC/n1108 , \AES_ENC/n1107 , \AES_ENC/n1106 , \AES_ENC/n1105 ,\AES_ENC/n1104 , \AES_ENC/n1103 , \AES_ENC/n1102 , \AES_ENC/n1101 ,\AES_ENC/n1100 , \AES_ENC/n1099 , \AES_ENC/n1098 , \AES_ENC/n1097 ,\AES_ENC/n1096 , \AES_ENC/n1095 , \AES_ENC/n1094 , \AES_ENC/n1093 ,\AES_ENC/n1092 , \AES_ENC/n1091 , \AES_ENC/n1090 , \AES_ENC/n1089 ,\AES_ENC/n1088 , \AES_ENC/n1087 , \AES_ENC/n1086 , \AES_ENC/n1085 ,\AES_ENC/n1084 , \AES_ENC/n1083 , \AES_ENC/n1082 , \AES_ENC/n1081 ,\AES_ENC/n1080 , \AES_ENC/n1079 , \AES_ENC/n1078 , \AES_ENC/n1077 ,\AES_ENC/n1076 , \AES_ENC/n1075 , \AES_ENC/n1074 , \AES_ENC/n1073 ,\AES_ENC/n1072 , \AES_ENC/n1071 , \AES_ENC/n1070 , \AES_ENC/n1069 ,\AES_ENC/n1068 , \AES_ENC/n1067 , \AES_ENC/n1066 , \AES_ENC/n1065 ,\AES_ENC/n1064 , \AES_ENC/n1063 , \AES_ENC/n1062 , \AES_ENC/n1061 ,\AES_ENC/n1060 , \AES_ENC/n1059 , \AES_ENC/n1058 , \AES_ENC/n1057 ,\AES_ENC/n1056 , \AES_ENC/n1055 , \AES_ENC/n1054 , \AES_ENC/n1053 ,\AES_ENC/n1052 , \AES_ENC/n1051 , \AES_ENC/n1050 , \AES_ENC/n1049 ,\AES_ENC/n1048 , \AES_ENC/n1047 , \AES_ENC/n1046 , \AES_ENC/n1045 ,\AES_ENC/n1044 , \AES_ENC/n1043 , \AES_ENC/n1042 , \AES_ENC/n1041 ,\AES_ENC/n1040 , \AES_ENC/n1039 , \AES_ENC/n1038 , \AES_ENC/n1037 ,\AES_ENC/n1036 , \AES_ENC/n1035 , \AES_ENC/n1034 , \AES_ENC/n1033 ,\AES_ENC/n1032 , \AES_ENC/n1031 , \AES_ENC/n1030 , \AES_ENC/n1029 ,\AES_ENC/n1028 , \AES_ENC/n1027 , \AES_ENC/n1026 , \AES_ENC/n1025 ,\AES_ENC/n1024 , \AES_ENC/n1023 , \AES_ENC/n1022 , \AES_ENC/n1021 ,\AES_ENC/n1020 , \AES_ENC/n1019 , \AES_ENC/n1018 , \AES_ENC/n1017 ,\AES_ENC/n1016 , \AES_ENC/n1015 , \AES_ENC/n1014 , \AES_ENC/n1013 ,\AES_ENC/n1012 , \AES_ENC/n1011 , \AES_ENC/n1010 , \AES_ENC/n1009 ,\AES_ENC/n1008 , \AES_ENC/n1007 , \AES_ENC/n1006 , \AES_ENC/n1005 ,\AES_ENC/n1004 , \AES_ENC/n1003 , \AES_ENC/n1002 , \AES_ENC/n1001 ,\AES_ENC/n1000 , \AES_ENC/n999 , \AES_ENC/n998 , \AES_ENC/n997 ,\AES_ENC/n996 , \AES_ENC/n995 , \AES_ENC/n994 , \AES_ENC/n993 ,\AES_ENC/n992 , \AES_ENC/n991 , \AES_ENC/n990 , \AES_ENC/n989 ,\AES_ENC/n988 , \AES_ENC/n987 , \AES_ENC/n986 , \AES_ENC/n985 ,\AES_ENC/n984 , \AES_ENC/n983 , \AES_ENC/n982 , \AES_ENC/n981 ,\AES_ENC/n980 , \AES_ENC/n979 , \AES_ENC/n978 , \AES_ENC/n977 ,\AES_ENC/n976 , \AES_ENC/n975 , \AES_ENC/n974 , \AES_ENC/n973 ,\AES_ENC/n972 , \AES_ENC/n971 , \AES_ENC/n970 , \AES_ENC/n969 ,\AES_ENC/n968 , \AES_ENC/n967 , \AES_ENC/n966 , \AES_ENC/n965 ,\AES_ENC/n964 , \AES_ENC/n963 , \AES_ENC/n962 , \AES_ENC/n961 ,\AES_ENC/n960 , \AES_ENC/n959 , \AES_ENC/n958 , \AES_ENC/n957 ,\AES_ENC/n956 , \AES_ENC/n955 , \AES_ENC/n954 , \AES_ENC/n953 ,\AES_ENC/n952 , \AES_ENC/n951 , \AES_ENC/n950 , \AES_ENC/n949 ,\AES_ENC/n948 , \AES_ENC/n947 , \AES_ENC/n946 , \AES_ENC/n945 ,\AES_ENC/n944 , \AES_ENC/n943 , \AES_ENC/n942 , \AES_ENC/n941 ,\AES_ENC/n940 , \AES_ENC/n939 , \AES_ENC/n938 , \AES_ENC/n937 ,\AES_ENC/n936 , \AES_ENC/n935 , \AES_ENC/n934 , \AES_ENC/n933 ,\AES_ENC/n932 , \AES_ENC/n931 , \AES_ENC/n930 , \AES_ENC/n929 ,\AES_ENC/n928 , \AES_ENC/n927 , \AES_ENC/n926 , \AES_ENC/n925 ,\AES_ENC/n924 , \AES_ENC/n923 , \AES_ENC/n922 , \AES_ENC/n921 ,\AES_ENC/n920 , \AES_ENC/n919 , \AES_ENC/n918 , \AES_ENC/n917 ,\AES_ENC/n916 , \AES_ENC/n915 , \AES_ENC/n914 , \AES_ENC/n913 ,\AES_ENC/n912 , \AES_ENC/n911 , \AES_ENC/n910 , \AES_ENC/n909 ,\AES_ENC/n908 , \AES_ENC/n907 , \AES_ENC/n906 , \AES_ENC/n905 ,\AES_ENC/n904 , \AES_ENC/n903 , \AES_ENC/n902 , \AES_ENC/n901 ,\AES_ENC/n900 , \AES_ENC/n899 , \AES_ENC/n898 , \AES_ENC/n897 ,\AES_ENC/n896 , \AES_ENC/n895 , \AES_ENC/n894 , \AES_ENC/n893 ,\AES_ENC/n892 , \AES_ENC/n891 , \AES_ENC/n890 , \AES_ENC/n889 ,\AES_ENC/n888 , \AES_ENC/n887 , \AES_ENC/n886 , \AES_ENC/n885 ,\AES_ENC/n884 , \AES_ENC/n883 , \AES_ENC/n882 , \AES_ENC/n881 ,\AES_ENC/n880 , \AES_ENC/n879 , \AES_ENC/n878 , \AES_ENC/n877 ,\AES_ENC/n876 , \AES_ENC/n875 , \AES_ENC/n874 , \AES_ENC/n873 ,\AES_ENC/n872 , \AES_ENC/n871 , \AES_ENC/n870 , \AES_ENC/n869 ,\AES_ENC/n868 , \AES_ENC/n867 , \AES_ENC/n866 , \AES_ENC/n865 ,\AES_ENC/n864 , \AES_ENC/n863 , \AES_ENC/n862 , \AES_ENC/n861 ,\AES_ENC/n860 , \AES_ENC/n859 , \AES_ENC/n858 , \AES_ENC/n857 ,\AES_ENC/n856 , \AES_ENC/n855 , \AES_ENC/n854 , \AES_ENC/n853 ,\AES_ENC/n852 , \AES_ENC/n851 , \AES_ENC/n850 , \AES_ENC/n849 ,\AES_ENC/n848 , \AES_ENC/n847 , \AES_ENC/n846 , \AES_ENC/n845 ,\AES_ENC/n844 , \AES_ENC/n843 , \AES_ENC/n842 , \AES_ENC/n841 ,\AES_ENC/n840 , \AES_ENC/n839 , \AES_ENC/n838 , \AES_ENC/n837 ,\AES_ENC/n836 , \AES_ENC/n835 , \AES_ENC/n834 , \AES_ENC/n833 ,\AES_ENC/n832 , \AES_ENC/n831 , \AES_ENC/n830 , \AES_ENC/n829 ,\AES_ENC/n828 , \AES_ENC/n827 , \AES_ENC/n826 , \AES_ENC/n825 ,\AES_ENC/n824 , \AES_ENC/n823 , \AES_ENC/n822 , \AES_ENC/n821 ,\AES_ENC/n820 , \AES_ENC/n819 , \AES_ENC/n818 , \AES_ENC/n817 ,\AES_ENC/n816 , \AES_ENC/n815 , \AES_ENC/n814 , \AES_ENC/n813 ,\AES_ENC/n812 , \AES_ENC/n811 , \AES_ENC/n810 , \AES_ENC/n809 ,\AES_ENC/n808 , \AES_ENC/n807 , \AES_ENC/n806 , \AES_ENC/n805 ,\AES_ENC/n804 , \AES_ENC/n803 , \AES_ENC/n802 , \AES_ENC/n801 ,\AES_ENC/n800 , \AES_ENC/n799 , \AES_ENC/n798 , \AES_ENC/n797 ,\AES_ENC/n796 , \AES_ENC/n795 , \AES_ENC/n788 , \AES_ENC/n787 ,\AES_ENC/n786 , \AES_ENC/n785 , \AES_ENC/n784 , \AES_ENC/n783 ,\AES_ENC/n782 , \AES_ENC/n781 , \AES_ENC/n780 , \AES_ENC/n779 ,\AES_ENC/n778 , \AES_ENC/n777 , \AES_ENC/n776 , \AES_ENC/n775 ,\AES_ENC/n774 , \AES_ENC/n773 , \AES_ENC/n772 , \AES_ENC/n771 ,\AES_ENC/n770 , \AES_ENC/n769 , \AES_ENC/n768 , \AES_ENC/n767 ,\AES_ENC/n766 , \AES_ENC/n765 , \AES_ENC/n764 , \AES_ENC/n763 ,\AES_ENC/n762 , \AES_ENC/n761 , \AES_ENC/n760 , \AES_ENC/n759 ,\AES_ENC/n758 , \AES_ENC/n757 , \AES_ENC/n756 , \AES_ENC/n755 ,\AES_ENC/n754 , \AES_ENC/n753 , \AES_ENC/n752 , \AES_ENC/n751 ,\AES_ENC/n750 , \AES_ENC/n749 , \AES_ENC/n748 , \AES_ENC/n747 ,\AES_ENC/n746 , \AES_ENC/n745 , \AES_ENC/n744 , \AES_ENC/n743 ,\AES_ENC/n742 , \AES_ENC/n741 , \AES_ENC/n740 , \AES_ENC/n739 ,\AES_ENC/n738 , \AES_ENC/n737 , \AES_ENC/n736 , \AES_ENC/n735 ,\AES_ENC/n734 , \AES_ENC/n733 , \AES_ENC/n732 , \AES_ENC/n731 ,\AES_ENC/n730 , \AES_ENC/n729 , \AES_ENC/n728 , \AES_ENC/n727 ,\AES_ENC/n726 , \AES_ENC/n725 , \AES_ENC/n724 , \AES_ENC/n723 ,\AES_ENC/n722 , \AES_ENC/n721 , \AES_ENC/n720 , \AES_ENC/n719 ,\AES_ENC/n718 , \AES_ENC/n717 , \AES_ENC/n716 , \AES_ENC/n715 ,\AES_ENC/n714 , \AES_ENC/n713 , \AES_ENC/n712 , \AES_ENC/n711 ,\AES_ENC/n710 , \AES_ENC/n709 , \AES_ENC/n708 , \AES_ENC/n707 ,\AES_ENC/n706 , \AES_ENC/n705 , \AES_ENC/n704 , \AES_ENC/n703 ,\AES_ENC/n702 , \AES_ENC/n701 , \AES_ENC/n700 , \AES_ENC/n699 ,\AES_ENC/n698 , \AES_ENC/n697 , \AES_ENC/n696 , \AES_ENC/n695 ,\AES_ENC/n694 , \AES_ENC/n693 , \AES_ENC/n692 , \AES_ENC/n691 ,\AES_ENC/n690 , \AES_ENC/n689 , \AES_ENC/n688 , \AES_ENC/n687 ,\AES_ENC/n686 , \AES_ENC/n685 , \AES_ENC/n684 , \AES_ENC/n683 ,\AES_ENC/n682 , \AES_ENC/n681 , \AES_ENC/n680 , \AES_ENC/n679 ,\AES_ENC/n678 , \AES_ENC/n677 , \AES_ENC/n676 , \AES_ENC/n675 ,\AES_ENC/n674 , \AES_ENC/n673 , \AES_ENC/n672 , \AES_ENC/n671 ,\AES_ENC/n670 , \AES_ENC/n669 , \AES_ENC/n668 , \AES_ENC/n667 ,\AES_ENC/n666 , \AES_ENC/n665 , \AES_ENC/n664 , \AES_ENC/n663 ,\AES_ENC/n662 , \AES_ENC/n661 , \AES_ENC/N501 , \AES_ENC/N500 ,\AES_ENC/N499 , \AES_ENC/N498 , \AES_ENC/N497 , \AES_ENC/N496 ,\AES_ENC/N495 , \AES_ENC/N494 , \AES_ENC/N493 , \AES_ENC/N492 ,\AES_ENC/N491 , \AES_ENC/N490 , \AES_ENC/N489 , \AES_ENC/N488 ,\AES_ENC/N487 , \AES_ENC/N486 , \AES_ENC/N485 , \AES_ENC/N484 ,\AES_ENC/N483 , \AES_ENC/N482 , \AES_ENC/N481 , \AES_ENC/N480 ,\AES_ENC/N479 , \AES_ENC/N478 , \AES_ENC/N477 , \AES_ENC/N476 ,\AES_ENC/N475 , \AES_ENC/N474 , \AES_ENC/N473 , \AES_ENC/N472 ,\AES_ENC/N471 , \AES_ENC/N470 , \AES_ENC/N469 , \AES_ENC/N468 ,\AES_ENC/N467 , \AES_ENC/N466 , \AES_ENC/N465 , \AES_ENC/N464 ,\AES_ENC/N463 , \AES_ENC/N462 , \AES_ENC/N461 , \AES_ENC/N460 ,\AES_ENC/N459 , \AES_ENC/N458 , \AES_ENC/N457 , \AES_ENC/N456 ,\AES_ENC/N455 , \AES_ENC/N454 , \AES_ENC/N453 , \AES_ENC/N452 ,\AES_ENC/N451 , \AES_ENC/N450 , \AES_ENC/N449 , \AES_ENC/N448 ,\AES_ENC/N447 , \AES_ENC/N446 , \AES_ENC/N445 , \AES_ENC/N444 ,\AES_ENC/N443 , \AES_ENC/N442 , \AES_ENC/N441 , \AES_ENC/N440 ,\AES_ENC/N439 , \AES_ENC/N438 , \AES_ENC/N437 , \AES_ENC/N436 ,\AES_ENC/N435 , \AES_ENC/N434 , \AES_ENC/N433 , \AES_ENC/N432 ,\AES_ENC/N431 , \AES_ENC/N430 , \AES_ENC/N429 , \AES_ENC/N428 ,\AES_ENC/N427 , \AES_ENC/N426 , \AES_ENC/N425 , \AES_ENC/N424 ,\AES_ENC/N423 , \AES_ENC/N422 , \AES_ENC/N421 , \AES_ENC/N420 ,\AES_ENC/N419 , \AES_ENC/N418 , \AES_ENC/N417 , \AES_ENC/N416 ,\AES_ENC/N415 , \AES_ENC/N414 , \AES_ENC/N413 , \AES_ENC/N412 ,\AES_ENC/N411 , \AES_ENC/N410 , \AES_ENC/N409 , \AES_ENC/N408 ,\AES_ENC/N407 , \AES_ENC/N406 , \AES_ENC/N405 , \AES_ENC/N404 ,\AES_ENC/N403 , \AES_ENC/N402 , \AES_ENC/N401 , \AES_ENC/N400 ,\AES_ENC/N399 , \AES_ENC/N398 , \AES_ENC/N397 , \AES_ENC/N396 ,\AES_ENC/N395 , \AES_ENC/N394 , \AES_ENC/N393 , \AES_ENC/N392 ,\AES_ENC/N391 , \AES_ENC/N390 , \AES_ENC/N389 , \AES_ENC/N388 ,\AES_ENC/N387 , \AES_ENC/N386 , \AES_ENC/N385 , \AES_ENC/N384 ,\AES_ENC/N383 , \AES_ENC/N382 , \AES_ENC/N381 , \AES_ENC/N380 ,\AES_ENC/N379 , \AES_ENC/N378 , \AES_ENC/N377 , \AES_ENC/N376 ,\AES_ENC/N375 , \AES_ENC/N374 , \AES_ENC/sa33_sub[0] ,\AES_ENC/sa33_sub[1] , \AES_ENC/sa33_sub[2] , \AES_ENC/sa33_sub[3] ,\AES_ENC/sa33_sub[4] , \AES_ENC/sa33_sub[5] , \AES_ENC/sa33_sub[6] ,\AES_ENC/sa33_sub[7] , \AES_ENC/sa32_sub[0] , \AES_ENC/sa32_sub[1] ,\AES_ENC/sa32_sub[2] , \AES_ENC/sa32_sub[3] , \AES_ENC/sa32_sub[4] ,\AES_ENC/sa32_sub[5] , \AES_ENC/sa32_sub[6] , \AES_ENC/sa32_sub[7] ,\AES_ENC/sa31_sub[0] , \AES_ENC/sa31_sub[1] , \AES_ENC/sa31_sub[2] ,\AES_ENC/sa31_sub[3] , \AES_ENC/sa31_sub[4] , \AES_ENC/sa31_sub[5] ,\AES_ENC/sa31_sub[6] , \AES_ENC/sa31_sub[7] , \AES_ENC/sa30_sub[0] ,\AES_ENC/sa30_sub[1] , \AES_ENC/sa30_sub[2] , \AES_ENC/sa30_sub[3] ,\AES_ENC/sa30_sub[4] , \AES_ENC/sa30_sub[5] , \AES_ENC/sa30_sub[6] ,\AES_ENC/sa30_sub[7] , \AES_ENC/sa23_sub[0] , \AES_ENC/sa23_sub[1] ,\AES_ENC/sa23_sub[2] , \AES_ENC/sa23_sub[3] , \AES_ENC/sa23_sub[4] ,\AES_ENC/sa23_sub[5] , \AES_ENC/sa23_sub[6] , \AES_ENC/sa23_sub[7] ,\AES_ENC/sa22_sub[0] , \AES_ENC/sa22_sub[1] , \AES_ENC/sa22_sub[2] ,\AES_ENC/sa22_sub[3] , \AES_ENC/sa22_sub[4] , \AES_ENC/sa22_sub[5] ,\AES_ENC/sa22_sub[6] , \AES_ENC/sa22_sub[7] , \AES_ENC/sa21_sub[0] ,\AES_ENC/sa21_sub[1] , \AES_ENC/sa21_sub[2] , \AES_ENC/sa21_sub[3] ,\AES_ENC/sa21_sub[4] , \AES_ENC/sa21_sub[5] , \AES_ENC/sa21_sub[6] ,\AES_ENC/sa21_sub[7] , \AES_ENC/sa20_sub[0] , \AES_ENC/sa20_sub[1] ,\AES_ENC/sa20_sub[2] , \AES_ENC/sa20_sub[3] , \AES_ENC/sa20_sub[4] ,\AES_ENC/sa20_sub[5] , \AES_ENC/sa20_sub[6] , \AES_ENC/sa20_sub[7] ,\AES_ENC/sa13_sub[0] , \AES_ENC/sa13_sub[1] , \AES_ENC/sa13_sub[2] ,\AES_ENC/sa13_sub[3] , \AES_ENC/sa13_sub[4] , \AES_ENC/sa13_sub[5] ,\AES_ENC/sa13_sub[6] , \AES_ENC/sa13_sub[7] , \AES_ENC/sa12_sub[0] ,\AES_ENC/sa12_sub[1] , \AES_ENC/sa12_sub[2] , \AES_ENC/sa12_sub[3] ,\AES_ENC/sa12_sub[4] , \AES_ENC/sa12_sub[5] , \AES_ENC/sa12_sub[6] ,\AES_ENC/sa12_sub[7] , \AES_ENC/sa11_sub[0] , \AES_ENC/sa11_sub[1] ,\AES_ENC/sa11_sub[2] , \AES_ENC/sa11_sub[3] , \AES_ENC/sa11_sub[4] ,\AES_ENC/sa11_sub[5] , \AES_ENC/sa11_sub[6] , \AES_ENC/sa11_sub[7] ,\AES_ENC/sa10_sub[0] , \AES_ENC/sa10_sub[1] , \AES_ENC/sa10_sub[2] ,\AES_ENC/sa10_sub[3] , \AES_ENC/sa10_sub[4] , \AES_ENC/sa10_sub[5] ,\AES_ENC/sa10_sub[6] , \AES_ENC/sa10_sub[7] , \AES_ENC/sa03_sub[0] ,\AES_ENC/sa03_sub[1] , \AES_ENC/sa03_sub[2] , \AES_ENC/sa03_sub[3] ,\AES_ENC/sa03_sub[4] , \AES_ENC/sa03_sub[5] , \AES_ENC/sa03_sub[6] ,\AES_ENC/sa03_sub[7] , \AES_ENC/sa02_sub[0] , \AES_ENC/sa02_sub[1] ,\AES_ENC/sa02_sub[2] , \AES_ENC/sa02_sub[3] , \AES_ENC/sa02_sub[4] ,\AES_ENC/sa02_sub[5] , \AES_ENC/sa02_sub[6] , \AES_ENC/sa02_sub[7] ,\AES_ENC/sa01_sub[0] , \AES_ENC/sa01_sub[1] , \AES_ENC/sa01_sub[2] ,\AES_ENC/sa01_sub[3] , \AES_ENC/sa01_sub[4] , \AES_ENC/sa01_sub[5] ,\AES_ENC/sa01_sub[6] , \AES_ENC/sa01_sub[7] , \AES_ENC/sa00_sub[0] ,\AES_ENC/sa00_sub[1] , \AES_ENC/sa00_sub[2] , \AES_ENC/sa00_sub[3] ,\AES_ENC/sa00_sub[4] , \AES_ENC/sa00_sub[5] , \AES_ENC/sa00_sub[6] ,\AES_ENC/sa00_sub[7] , \AES_ENC/N277 , \AES_ENC/N276 , \AES_ENC/N275 ,\AES_ENC/N274 , \AES_ENC/N273 , \AES_ENC/N272 , \AES_ENC/N271 ,\AES_ENC/N270 , \AES_ENC/N261 , \AES_ENC/N260 , \AES_ENC/N259 ,\AES_ENC/N258 , \AES_ENC/N257 , \AES_ENC/N256 , \AES_ENC/N255 ,\AES_ENC/N254 , \AES_ENC/N245 , \AES_ENC/N244 , \AES_ENC/N243 ,\AES_ENC/N242 , \AES_ENC/N241 , \AES_ENC/N240 , \AES_ENC/N239 ,\AES_ENC/N238 , \AES_ENC/N229 , \AES_ENC/N228 , \AES_ENC/N227 ,\AES_ENC/N226 , \AES_ENC/N225 , \AES_ENC/N224 , \AES_ENC/N223 ,\AES_ENC/N222 , \AES_ENC/w0[0] , \AES_ENC/w0[1] , \AES_ENC/w0[2] ,\AES_ENC/w0[3] , \AES_ENC/w0[4] , \AES_ENC/w0[5] , \AES_ENC/w0[6] ,\AES_ENC/w0[7] , \AES_ENC/w0[8] , \AES_ENC/w0[9] , \AES_ENC/w0[10] ,\AES_ENC/w0[11] , \AES_ENC/w0[12] , \AES_ENC/w0[13] ,\AES_ENC/w0[14] , \AES_ENC/w0[15] , \AES_ENC/w0[16] ,\AES_ENC/w0[17] , \AES_ENC/w0[18] , \AES_ENC/w0[19] ,\AES_ENC/w0[20] , \AES_ENC/w0[21] , \AES_ENC/w0[22] ,\AES_ENC/w0[23] , \AES_ENC/w0[24] , \AES_ENC/w0[25] ,\AES_ENC/w0[26] , \AES_ENC/w0[27] , \AES_ENC/w0[28] ,\AES_ENC/w0[29] , \AES_ENC/w0[30] , \AES_ENC/w0[31] , \AES_ENC/N213 ,\AES_ENC/N212 , \AES_ENC/N211 , \AES_ENC/N210 , \AES_ENC/N209 ,\AES_ENC/N208 , \AES_ENC/N207 , \AES_ENC/N206 , \AES_ENC/N197 ,\AES_ENC/N196 , \AES_ENC/N195 , \AES_ENC/N194 , \AES_ENC/N193 ,\AES_ENC/N192 , \AES_ENC/N191 , \AES_ENC/N190 , \AES_ENC/N181 ,\AES_ENC/N180 , \AES_ENC/N179 , \AES_ENC/N178 , \AES_ENC/N177 ,\AES_ENC/N176 , \AES_ENC/N175 , \AES_ENC/N174 , \AES_ENC/N165 ,\AES_ENC/N164 , \AES_ENC/N163 , \AES_ENC/N162 , \AES_ENC/N161 ,\AES_ENC/N160 , \AES_ENC/N159 , \AES_ENC/N158 , \AES_ENC/w1[0] ,\AES_ENC/w1[1] , \AES_ENC/w1[2] , \AES_ENC/w1[3] , \AES_ENC/w1[4] ,\AES_ENC/w1[5] , \AES_ENC/w1[6] , \AES_ENC/w1[7] , \AES_ENC/w1[8] ,\AES_ENC/w1[9] , \AES_ENC/w1[10] , \AES_ENC/w1[11] , \AES_ENC/w1[12] ,\AES_ENC/w1[13] , \AES_ENC/w1[14] , \AES_ENC/w1[15] ,\AES_ENC/w1[16] , \AES_ENC/w1[17] , \AES_ENC/w1[18] ,\AES_ENC/w1[19] , \AES_ENC/w1[20] , \AES_ENC/w1[21] ,\AES_ENC/w1[22] , \AES_ENC/w1[23] , \AES_ENC/w1[24] ,\AES_ENC/w1[25] , \AES_ENC/w1[26] , \AES_ENC/w1[27] ,\AES_ENC/w1[28] , \AES_ENC/w1[29] , \AES_ENC/w1[30] ,\AES_ENC/w1[31] , \AES_ENC/N149 , \AES_ENC/N148 , \AES_ENC/N147 ,\AES_ENC/N146 , \AES_ENC/N145 , \AES_ENC/N144 , \AES_ENC/N143 ,\AES_ENC/N142 , \AES_ENC/N133 , \AES_ENC/N132 , \AES_ENC/N131 ,\AES_ENC/N130 , \AES_ENC/N129 , \AES_ENC/N128 , \AES_ENC/N127 ,\AES_ENC/N126 , \AES_ENC/N117 , \AES_ENC/N116 , \AES_ENC/N115 ,\AES_ENC/N114 , \AES_ENC/N113 , \AES_ENC/N112 , \AES_ENC/N111 ,\AES_ENC/N110 , \AES_ENC/N101 , \AES_ENC/N100 , \AES_ENC/N99 ,\AES_ENC/N98 , \AES_ENC/N97 , \AES_ENC/N96 , \AES_ENC/N95 ,\AES_ENC/N94 , \AES_ENC/w2[0] , \AES_ENC/w2[1] , \AES_ENC/w2[2] ,\AES_ENC/w2[3] , \AES_ENC/w2[4] , \AES_ENC/w2[5] , \AES_ENC/w2[6] ,\AES_ENC/w2[7] , \AES_ENC/w2[8] , \AES_ENC/w2[9] , \AES_ENC/w2[10] ,\AES_ENC/w2[11] , \AES_ENC/w2[12] , \AES_ENC/w2[13] ,\AES_ENC/w2[14] , \AES_ENC/w2[15] , \AES_ENC/w2[16] ,\AES_ENC/w2[17] , \AES_ENC/w2[18] , \AES_ENC/w2[19] ,\AES_ENC/w2[20] , \AES_ENC/w2[21] , \AES_ENC/w2[22] ,\AES_ENC/w2[23] , \AES_ENC/w2[24] , \AES_ENC/w2[25] ,\AES_ENC/w2[26] , \AES_ENC/w2[27] , \AES_ENC/w2[28] ,\AES_ENC/w2[29] , \AES_ENC/w2[30] , \AES_ENC/w2[31] , \AES_ENC/N85 ,\AES_ENC/N84 , \AES_ENC/N83 , \AES_ENC/N82 , \AES_ENC/N81 ,\AES_ENC/N80 , \AES_ENC/N79 , \AES_ENC/N78 , \AES_ENC/N69 ,\AES_ENC/N68 , \AES_ENC/N67 , \AES_ENC/N66 , \AES_ENC/N65 ,\AES_ENC/N64 , \AES_ENC/N63 , \AES_ENC/N62 , \AES_ENC/N53 ,\AES_ENC/N52 , \AES_ENC/N51 , \AES_ENC/N50 , \AES_ENC/N49 ,\AES_ENC/N48 , \AES_ENC/N47 , \AES_ENC/N46 , \AES_ENC/N37 ,\AES_ENC/N36 , \AES_ENC/N35 , \AES_ENC/N34 , \AES_ENC/N33 ,\AES_ENC/N32 , \AES_ENC/N31 , \AES_ENC/N30 , \AES_ENC/w3[0] ,\AES_ENC/w3[1] , \AES_ENC/w3[2] , \AES_ENC/w3[3] , \AES_ENC/w3[4] ,\AES_ENC/w3[5] , \AES_ENC/w3[6] , \AES_ENC/w3[7] , \AES_ENC/w3[8] ,\AES_ENC/w3[9] , \AES_ENC/w3[10] , \AES_ENC/w3[11] , \AES_ENC/w3[12] ,\AES_ENC/w3[13] , \AES_ENC/w3[14] , \AES_ENC/w3[15] ,\AES_ENC/w3[16] , \AES_ENC/w3[17] , \AES_ENC/w3[18] ,\AES_ENC/w3[19] , \AES_ENC/w3[20] , \AES_ENC/w3[21] ,\AES_ENC/w3[22] , \AES_ENC/w3[23] , \AES_ENC/w3[24] ,\AES_ENC/w3[25] , \AES_ENC/w3[26] , \AES_ENC/w3[27] ,\AES_ENC/w3[28] , \AES_ENC/w3[29] , \AES_ENC/w3[30] ,\AES_ENC/w3[31] , \AES_ENC/text_in_r[0] , \AES_ENC/text_in_r[1] ,\AES_ENC/text_in_r[2] , \AES_ENC/text_in_r[3] ,\AES_ENC/text_in_r[4] , \AES_ENC/text_in_r[5] ,\AES_ENC/text_in_r[6] , \AES_ENC/text_in_r[7] ,\AES_ENC/text_in_r[8] , \AES_ENC/text_in_r[9] ,\AES_ENC/text_in_r[10] , \AES_ENC/text_in_r[11] ,\AES_ENC/text_in_r[12] , \AES_ENC/text_in_r[13] ,\AES_ENC/text_in_r[14] , \AES_ENC/text_in_r[15] ,\AES_ENC/text_in_r[16] , \AES_ENC/text_in_r[17] ,\AES_ENC/text_in_r[18] , \AES_ENC/text_in_r[19] ,\AES_ENC/text_in_r[20] , \AES_ENC/text_in_r[21] ,\AES_ENC/text_in_r[22] , \AES_ENC/text_in_r[23] ,\AES_ENC/text_in_r[24] , \AES_ENC/text_in_r[25] ,\AES_ENC/text_in_r[26] , \AES_ENC/text_in_r[27] ,\AES_ENC/text_in_r[28] , \AES_ENC/text_in_r[29] ,\AES_ENC/text_in_r[30] , \AES_ENC/text_in_r[31] ,\AES_ENC/text_in_r[32] , \AES_ENC/text_in_r[33] ,\AES_ENC/text_in_r[34] , \AES_ENC/text_in_r[35] ,\AES_ENC/text_in_r[36] , \AES_ENC/text_in_r[37] ,\AES_ENC/text_in_r[38] , \AES_ENC/text_in_r[39] ,\AES_ENC/text_in_r[40] , \AES_ENC/text_in_r[41] ,\AES_ENC/text_in_r[42] , \AES_ENC/text_in_r[43] ,\AES_ENC/text_in_r[44] , \AES_ENC/text_in_r[45] ,\AES_ENC/text_in_r[46] , \AES_ENC/text_in_r[47] ,\AES_ENC/text_in_r[48] , \AES_ENC/text_in_r[49] ,\AES_ENC/text_in_r[50] , \AES_ENC/text_in_r[51] ,\AES_ENC/text_in_r[52] , \AES_ENC/text_in_r[53] ,\AES_ENC/text_in_r[54] , \AES_ENC/text_in_r[55] ,\AES_ENC/text_in_r[56] , \AES_ENC/text_in_r[57] ,\AES_ENC/text_in_r[58] , \AES_ENC/text_in_r[59] ,\AES_ENC/text_in_r[60] , \AES_ENC/text_in_r[61] ,\AES_ENC/text_in_r[62] , \AES_ENC/text_in_r[63] ,\AES_ENC/text_in_r[64] , \AES_ENC/text_in_r[65] ,\AES_ENC/text_in_r[66] , \AES_ENC/text_in_r[67] ,\AES_ENC/text_in_r[68] , \AES_ENC/text_in_r[69] ,\AES_ENC/text_in_r[70] , \AES_ENC/text_in_r[71] ,\AES_ENC/text_in_r[72] , \AES_ENC/text_in_r[73] ,\AES_ENC/text_in_r[74] , \AES_ENC/text_in_r[75] ,\AES_ENC/text_in_r[76] , \AES_ENC/text_in_r[77] ,\AES_ENC/text_in_r[78] , \AES_ENC/text_in_r[79] ,\AES_ENC/text_in_r[80] , \AES_ENC/text_in_r[81] ,\AES_ENC/text_in_r[82] , \AES_ENC/text_in_r[83] ,\AES_ENC/text_in_r[84] , \AES_ENC/text_in_r[85] ,\AES_ENC/text_in_r[86] , \AES_ENC/text_in_r[87] ,\AES_ENC/text_in_r[88] , \AES_ENC/text_in_r[89] ,\AES_ENC/text_in_r[90] , \AES_ENC/text_in_r[91] ,\AES_ENC/text_in_r[92] , \AES_ENC/text_in_r[93] ,\AES_ENC/text_in_r[94] , \AES_ENC/text_in_r[95] ,\AES_ENC/text_in_r[96] , \AES_ENC/text_in_r[97] ,\AES_ENC/text_in_r[98] , \AES_ENC/text_in_r[99] ,\AES_ENC/text_in_r[100] , \AES_ENC/text_in_r[101] ,\AES_ENC/text_in_r[102] , \AES_ENC/text_in_r[103] ,\AES_ENC/text_in_r[104] , \AES_ENC/text_in_r[105] ,\AES_ENC/text_in_r[106] , \AES_ENC/text_in_r[107] ,\AES_ENC/text_in_r[108] , \AES_ENC/text_in_r[109] ,\AES_ENC/text_in_r[110] , \AES_ENC/text_in_r[111] ,\AES_ENC/text_in_r[112] , \AES_ENC/text_in_r[113] ,\AES_ENC/text_in_r[114] , \AES_ENC/text_in_r[115] ,\AES_ENC/text_in_r[116] , \AES_ENC/text_in_r[117] ,\AES_ENC/text_in_r[118] , \AES_ENC/text_in_r[119] ,\AES_ENC/text_in_r[120] , \AES_ENC/text_in_r[121] ,\AES_ENC/text_in_r[122] , \AES_ENC/text_in_r[123] ,\AES_ENC/text_in_r[124] , \AES_ENC/text_in_r[125] ,\AES_ENC/text_in_r[126] , \AES_ENC/text_in_r[127] , \AES_ENC/N19 ,\AES_ENC/u0/n325 , \AES_ENC/u0/n324 , \AES_ENC/u0/n323 ,\AES_ENC/u0/n322 , \AES_ENC/u0/n321 , \AES_ENC/u0/n320 ,\AES_ENC/u0/n319 , \AES_ENC/u0/n318 , \AES_ENC/u0/n317 ,\AES_ENC/u0/n316 , \AES_ENC/u0/n315 , \AES_ENC/u0/n314 ,\AES_ENC/u0/n281 , \AES_ENC/u0/n280 , \AES_ENC/u0/n279 ,\AES_ENC/u0/n278 , \AES_ENC/u0/n277 , \AES_ENC/u0/n276 ,\AES_ENC/u0/n275 , \AES_ENC/u0/n274 , \AES_ENC/u0/n273 ,\AES_ENC/u0/n272 , \AES_ENC/u0/n2710 , \AES_ENC/u0/n2700 ,\AES_ENC/u0/n2690 , \AES_ENC/u0/n2680 , \AES_ENC/u0/n2670 ,\AES_ENC/u0/n2660 , \AES_ENC/u0/n2650 , \AES_ENC/u0/n2640 ,\AES_ENC/u0/n2630 , \AES_ENC/u0/n2620 , \AES_ENC/u0/n2610 ,\AES_ENC/u0/n2600 , \AES_ENC/u0/n2590 , \AES_ENC/u0/n2580 ,\AES_ENC/u0/n2570 , \AES_ENC/u0/n2560 , \AES_ENC/u0/n2550 ,\AES_ENC/u0/n2540 , \AES_ENC/u0/n2530 , \AES_ENC/u0/n2520 ,\AES_ENC/u0/n2510 , \AES_ENC/u0/n2500 , \AES_ENC/u0/n2490 ,\AES_ENC/u0/n2480 , \AES_ENC/u0/n2470 , \AES_ENC/u0/n2460 ,\AES_ENC/u0/n2450 , \AES_ENC/u0/n2440 , \AES_ENC/u0/n2430 ,\AES_ENC/u0/n2420 , \AES_ENC/u0/n2410 , \AES_ENC/u0/n2400 ,\AES_ENC/u0/n2390 , \AES_ENC/u0/n2380 , \AES_ENC/u0/n2370 ,\AES_ENC/u0/n2360 , \AES_ENC/u0/n2350 , \AES_ENC/u0/n2340 ,\AES_ENC/u0/n2330 , \AES_ENC/u0/n2320 , \AES_ENC/u0/n2310 ,\AES_ENC/u0/n2300 , \AES_ENC/u0/n2290 , \AES_ENC/u0/n2280 ,\AES_ENC/u0/n2270 , \AES_ENC/u0/n2260 , \AES_ENC/u0/n2250 ,\AES_ENC/u0/n2240 , \AES_ENC/u0/n2230 , \AES_ENC/u0/n2220 ,\AES_ENC/u0/n2210 , \AES_ENC/u0/n2200 , \AES_ENC/u0/n2190 ,\AES_ENC/u0/n2180 , \AES_ENC/u0/n2170 , \AES_ENC/u0/n2160 ,\AES_ENC/u0/n2150 , \AES_ENC/u0/n2140 , \AES_ENC/u0/n2130 ,\AES_ENC/u0/n2120 , \AES_ENC/u0/n2110 , \AES_ENC/u0/n2100 ,\AES_ENC/u0/n2090 , \AES_ENC/u0/n2080 , \AES_ENC/u0/n207 ,\AES_ENC/u0/n206 , \AES_ENC/u0/n2050 , \AES_ENC/u0/n2040 ,\AES_ENC/u0/n2030 , \AES_ENC/u0/n2020 , \AES_ENC/u0/n2010 ,\AES_ENC/u0/n2000 , \AES_ENC/u0/n1990 , \AES_ENC/u0/n1980 ,\AES_ENC/u0/n1970 , \AES_ENC/u0/n1960 , \AES_ENC/u0/n1950 ,\AES_ENC/u0/n1940 , \AES_ENC/u0/n1930 , \AES_ENC/u0/n1920 ,\AES_ENC/u0/n1910 , \AES_ENC/u0/n1900 , \AES_ENC/u0/n1890 ,\AES_ENC/u0/n1880 , \AES_ENC/u0/n1870 , \AES_ENC/u0/n1860 ,\AES_ENC/u0/n1850 , \AES_ENC/u0/n1840 , \AES_ENC/u0/n1830 ,\AES_ENC/u0/n1820 , \AES_ENC/u0/n1810 , \AES_ENC/u0/n1800 ,\AES_ENC/u0/n1790 , \AES_ENC/u0/n1780 , \AES_ENC/u0/n1770 ,\AES_ENC/u0/n1760 , \AES_ENC/u0/n1750 , \AES_ENC/u0/n1740 ,\AES_ENC/u0/n1730 , \AES_ENC/u0/n1720 , \AES_ENC/u0/n1711 ,\AES_ENC/u0/n1700 , \AES_ENC/u0/n1690 , \AES_ENC/u0/n1680 ,\AES_ENC/u0/n1670 , \AES_ENC/u0/n1660 , \AES_ENC/u0/n1650 ,\AES_ENC/u0/n1640 , \AES_ENC/u0/n1630 , \AES_ENC/u0/n1620 ,\AES_ENC/u0/n1611 , \AES_ENC/u0/n1600 , \AES_ENC/u0/n1590 ,\AES_ENC/u0/n1580 , \AES_ENC/u0/n1570 , \AES_ENC/u0/n1560 ,\AES_ENC/u0/n1550 , \AES_ENC/u0/n1540 , \AES_ENC/u0/n1530 ,\AES_ENC/u0/n1520 , \AES_ENC/u0/n1511 , \AES_ENC/u0/n1500 ,\AES_ENC/u0/n1490 , \AES_ENC/u0/n1480 , \AES_ENC/u0/n1470 ,\AES_ENC/u0/n1460 , \AES_ENC/u0/n1450 , \AES_ENC/u0/n1440 ,\AES_ENC/u0/n1430 , \AES_ENC/u0/n1420 , \AES_ENC/u0/n141 ,\AES_ENC/u0/n1401 , \AES_ENC/u0/n1390 , \AES_ENC/u0/n1380 ,\AES_ENC/u0/n1370 , \AES_ENC/u0/n1360 , \AES_ENC/u0/n1350 ,\AES_ENC/u0/n1340 , \AES_ENC/u0/n1330 , \AES_ENC/u0/n1320 ,\AES_ENC/u0/n1311 , \AES_ENC/u0/n1300 , \AES_ENC/u0/n1290 ,\AES_ENC/u0/n1280 , \AES_ENC/u0/n1270 , \AES_ENC/u0/n1260 ,\AES_ENC/u0/n1250 , \AES_ENC/u0/n1240 , \AES_ENC/u0/n1230 ,\AES_ENC/u0/n1220 , \AES_ENC/u0/n1211 , \AES_ENC/u0/n1200 ,\AES_ENC/u0/n1190 , \AES_ENC/u0/n1180 , \AES_ENC/u0/n1170 ,\AES_ENC/u0/n1160 , \AES_ENC/u0/n1150 , \AES_ENC/u0/n1140 ,\AES_ENC/u0/n1130 , \AES_ENC/u0/n1120 , \AES_ENC/u0/n1111 ,\AES_ENC/u0/n1100 , \AES_ENC/u0/n1090 , \AES_ENC/u0/n1080 ,\AES_ENC/u0/n1070 , \AES_ENC/u0/n1060 , \AES_ENC/u0/n1050 ,\AES_ENC/u0/n1040 , \AES_ENC/u0/n1030 , \AES_ENC/u0/n1020 ,\AES_ENC/u0/n1011 , \AES_ENC/u0/n1000 , \AES_ENC/u0/n990 ,\AES_ENC/u0/n980 , \AES_ENC/u0/n970 , \AES_ENC/u0/n960 ,\AES_ENC/u0/n950 , \AES_ENC/u0/n940 , \AES_ENC/u0/n930 ,\AES_ENC/u0/n920 , \AES_ENC/u0/n910 , \AES_ENC/u0/n900 ,\AES_ENC/u0/n890 , \AES_ENC/u0/n880 , \AES_ENC/u0/n870 ,\AES_ENC/u0/n860 , \AES_ENC/u0/n850 , \AES_ENC/u0/n840 ,\AES_ENC/u0/n830 , \AES_ENC/u0/n820 , \AES_ENC/u0/n810 ,\AES_ENC/u0/n800 , \AES_ENC/u0/n790 , \AES_ENC/u0/n780 ,\AES_ENC/u0/n770 , \AES_ENC/u0/n760 , \AES_ENC/u0/n75 ,\AES_ENC/u0/n74 , \AES_ENC/u0/n730 , \AES_ENC/u0/n720 ,\AES_ENC/u0/n710 , \AES_ENC/u0/n700 , \AES_ENC/u0/n690 ,\AES_ENC/u0/n680 , \AES_ENC/u0/n670 , \AES_ENC/u0/n660 ,\AES_ENC/u0/n650 , \AES_ENC/u0/n640 , \AES_ENC/u0/n630 ,\AES_ENC/u0/n620 , \AES_ENC/u0/n610 , \AES_ENC/u0/n600 ,\AES_ENC/u0/n590 , \AES_ENC/u0/n580 , \AES_ENC/u0/n570 ,\AES_ENC/u0/n560 , \AES_ENC/u0/n550 , \AES_ENC/u0/n540 ,\AES_ENC/u0/n530 , \AES_ENC/u0/n520 , \AES_ENC/u0/n510 ,\AES_ENC/u0/n500 , \AES_ENC/u0/n490 , \AES_ENC/u0/n480 ,\AES_ENC/u0/n470 , \AES_ENC/u0/n460 , \AES_ENC/u0/n450 ,\AES_ENC/u0/n440 , \AES_ENC/u0/n430 , \AES_ENC/u0/n420 ,\AES_ENC/u0/n41 , \AES_ENC/u0/n40 , \AES_ENC/u0/n39 ,\AES_ENC/u0/n38 , \AES_ENC/u0/n37 , \AES_ENC/u0/n36 ,\AES_ENC/u0/n35 , \AES_ENC/u0/n34 , \AES_ENC/u0/n33 ,\AES_ENC/u0/n32 , \AES_ENC/u0/n31 , \AES_ENC/u0/n30 ,\AES_ENC/u0/n29 , \AES_ENC/u0/n28 , \AES_ENC/u0/n27 ,\AES_ENC/u0/n26 , \AES_ENC/u0/n25 , \AES_ENC/u0/n24 ,\AES_ENC/u0/n23 , \AES_ENC/u0/n22 , \AES_ENC/u0/n21 ,\AES_ENC/u0/n20 , \AES_ENC/u0/n19 , \AES_ENC/u0/n18 ,\AES_ENC/u0/n1710 , \AES_ENC/u0/n1610 , \AES_ENC/u0/n1510 ,\AES_ENC/u0/n1400 , \AES_ENC/u0/n1310 , \AES_ENC/u0/n1210 ,\AES_ENC/u0/n1110 , \AES_ENC/u0/n1010 , \AES_ENC/u0/n9 ,\AES_ENC/u0/n8 , \AES_ENC/u0/n7 , \AES_ENC/u0/n6 , \AES_ENC/u0/n5 ,\AES_ENC/u0/n4 , \AES_ENC/u0/n3 , \AES_ENC/u0/n2 , \AES_ENC/u0/n313 ,\AES_ENC/u0/n312 , \AES_ENC/u0/n311 , \AES_ENC/u0/n310 ,\AES_ENC/u0/n309 , \AES_ENC/u0/n308 , \AES_ENC/u0/n307 ,\AES_ENC/u0/n306 , \AES_ENC/u0/n305 , \AES_ENC/u0/n304 ,\AES_ENC/u0/n303 , \AES_ENC/u0/n302 , \AES_ENC/u0/n301 ,\AES_ENC/u0/n300 , \AES_ENC/u0/n299 , \AES_ENC/u0/n298 ,\AES_ENC/u0/n297 , \AES_ENC/u0/n296 , \AES_ENC/u0/n295 ,\AES_ENC/u0/n294 , \AES_ENC/u0/n293 , \AES_ENC/u0/n292 ,\AES_ENC/u0/n291 , \AES_ENC/u0/n290 , \AES_ENC/u0/n289 ,\AES_ENC/u0/n288 , \AES_ENC/u0/n287 , \AES_ENC/u0/n286 ,\AES_ENC/u0/n285 , \AES_ENC/u0/n284 , \AES_ENC/u0/n283 ,\AES_ENC/u0/n282 , \AES_ENC/u0/N271 , \AES_ENC/u0/N270 ,\AES_ENC/u0/N269 , \AES_ENC/u0/N268 , \AES_ENC/u0/N267 ,\AES_ENC/u0/N266 , \AES_ENC/u0/N265 , \AES_ENC/u0/N264 ,\AES_ENC/u0/N263 , \AES_ENC/u0/N262 , \AES_ENC/u0/N261 ,\AES_ENC/u0/N260 , \AES_ENC/u0/N259 , \AES_ENC/u0/N258 ,\AES_ENC/u0/N257 , \AES_ENC/u0/N256 , \AES_ENC/u0/N255 ,\AES_ENC/u0/N254 , \AES_ENC/u0/N253 , \AES_ENC/u0/N252 ,\AES_ENC/u0/N251 , \AES_ENC/u0/N250 , \AES_ENC/u0/N249 ,\AES_ENC/u0/N248 , \AES_ENC/u0/N247 , \AES_ENC/u0/N246 ,\AES_ENC/u0/N245 , \AES_ENC/u0/N244 , \AES_ENC/u0/N243 ,\AES_ENC/u0/N242 , \AES_ENC/u0/N241 , \AES_ENC/u0/N240 ,\AES_ENC/u0/N239 , \AES_ENC/u0/N238 , \AES_ENC/u0/N237 ,\AES_ENC/u0/N236 , \AES_ENC/u0/N235 , \AES_ENC/u0/N234 ,\AES_ENC/u0/N233 , \AES_ENC/u0/N232 , \AES_ENC/u0/N231 ,\AES_ENC/u0/N230 , \AES_ENC/u0/N229 , \AES_ENC/u0/N228 ,\AES_ENC/u0/N227 , \AES_ENC/u0/N226 , \AES_ENC/u0/N225 ,\AES_ENC/u0/N224 , \AES_ENC/u0/N223 , \AES_ENC/u0/N222 ,\AES_ENC/u0/N221 , \AES_ENC/u0/N220 , \AES_ENC/u0/N219 ,\AES_ENC/u0/N218 , \AES_ENC/u0/N217 , \AES_ENC/u0/N216 ,\AES_ENC/u0/N215 , \AES_ENC/u0/N214 , \AES_ENC/u0/N213 ,\AES_ENC/u0/N212 , \AES_ENC/u0/N211 , \AES_ENC/u0/N210 ,\AES_ENC/u0/N209 , \AES_ENC/u0/N208 , \AES_ENC/u0/N205 ,\AES_ENC/u0/N204 , \AES_ENC/u0/N203 , \AES_ENC/u0/N202 ,\AES_ENC/u0/N201 , \AES_ENC/u0/N200 , \AES_ENC/u0/N199 ,\AES_ENC/u0/N198 , \AES_ENC/u0/N197 , \AES_ENC/u0/N196 ,\AES_ENC/u0/N195 , \AES_ENC/u0/N194 , \AES_ENC/u0/N193 ,\AES_ENC/u0/N192 , \AES_ENC/u0/N191 , \AES_ENC/u0/N190 ,\AES_ENC/u0/N189 , \AES_ENC/u0/N188 , \AES_ENC/u0/N187 ,\AES_ENC/u0/N186 , \AES_ENC/u0/N185 , \AES_ENC/u0/N184 ,\AES_ENC/u0/N183 , \AES_ENC/u0/N182 , \AES_ENC/u0/N181 ,\AES_ENC/u0/N180 , \AES_ENC/u0/N179 , \AES_ENC/u0/N178 ,\AES_ENC/u0/N177 , \AES_ENC/u0/N176 , \AES_ENC/u0/N175 ,\AES_ENC/u0/N174 , \AES_ENC/u0/N173 , \AES_ENC/u0/N172 ,\AES_ENC/u0/N171 , \AES_ENC/u0/N170 , \AES_ENC/u0/N169 ,\AES_ENC/u0/N168 , \AES_ENC/u0/N167 , \AES_ENC/u0/N166 ,\AES_ENC/u0/N165 , \AES_ENC/u0/N164 , \AES_ENC/u0/N163 ,\AES_ENC/u0/N162 , \AES_ENC/u0/N161 , \AES_ENC/u0/N160 ,\AES_ENC/u0/N159 , \AES_ENC/u0/N158 , \AES_ENC/u0/N157 ,\AES_ENC/u0/N156 , \AES_ENC/u0/N155 , \AES_ENC/u0/N154 ,\AES_ENC/u0/N153 , \AES_ENC/u0/N152 , \AES_ENC/u0/N151 ,\AES_ENC/u0/N150 , \AES_ENC/u0/N149 , \AES_ENC/u0/N148 ,\AES_ENC/u0/N147 , \AES_ENC/u0/N146 , \AES_ENC/u0/N145 ,\AES_ENC/u0/N144 , \AES_ENC/u0/N143 , \AES_ENC/u0/N142 ,\AES_ENC/u0/N139 , \AES_ENC/u0/N138 , \AES_ENC/u0/N137 ,\AES_ENC/u0/N136 , \AES_ENC/u0/N135 , \AES_ENC/u0/N134 ,\AES_ENC/u0/N133 , \AES_ENC/u0/N132 , \AES_ENC/u0/N131 ,\AES_ENC/u0/N130 , \AES_ENC/u0/N129 , \AES_ENC/u0/N128 ,\AES_ENC/u0/N127 , \AES_ENC/u0/N126 , \AES_ENC/u0/N125 ,\AES_ENC/u0/N124 , \AES_ENC/u0/N123 , \AES_ENC/u0/N122 ,\AES_ENC/u0/N121 , \AES_ENC/u0/N120 , \AES_ENC/u0/N119 ,\AES_ENC/u0/N118 , \AES_ENC/u0/N117 , \AES_ENC/u0/N116 ,\AES_ENC/u0/N115 , \AES_ENC/u0/N114 , \AES_ENC/u0/N113 ,\AES_ENC/u0/N112 , \AES_ENC/u0/N111 , \AES_ENC/u0/N110 ,\AES_ENC/u0/N109 , \AES_ENC/u0/N108 , \AES_ENC/u0/N107 ,\AES_ENC/u0/N106 , \AES_ENC/u0/N105 , \AES_ENC/u0/N104 ,\AES_ENC/u0/N103 , \AES_ENC/u0/N102 , \AES_ENC/u0/N101 ,\AES_ENC/u0/N100 , \AES_ENC/u0/N99 , \AES_ENC/u0/N98 ,\AES_ENC/u0/N97 , \AES_ENC/u0/N96 , \AES_ENC/u0/N95 ,\AES_ENC/u0/N94 , \AES_ENC/u0/N93 , \AES_ENC/u0/N92 ,\AES_ENC/u0/N91 , \AES_ENC/u0/N90 , \AES_ENC/u0/N89 ,\AES_ENC/u0/N88 , \AES_ENC/u0/N87 , \AES_ENC/u0/N86 ,\AES_ENC/u0/N85 , \AES_ENC/u0/N84 , \AES_ENC/u0/N83 ,\AES_ENC/u0/N82 , \AES_ENC/u0/N81 , \AES_ENC/u0/N80 ,\AES_ENC/u0/N79 , \AES_ENC/u0/N78 , \AES_ENC/u0/N77 ,\AES_ENC/u0/N76 , \AES_ENC/u0/N73 , \AES_ENC/u0/N72 ,\AES_ENC/u0/N71 , \AES_ENC/u0/N70 , \AES_ENC/u0/N69 ,\AES_ENC/u0/N68 , \AES_ENC/u0/N67 , \AES_ENC/u0/N66 ,\AES_ENC/u0/N65 , \AES_ENC/u0/N64 , \AES_ENC/u0/N63 ,\AES_ENC/u0/N62 , \AES_ENC/u0/N61 , \AES_ENC/u0/N60 ,\AES_ENC/u0/N59 , \AES_ENC/u0/N58 , \AES_ENC/u0/N57 ,\AES_ENC/u0/N56 , \AES_ENC/u0/N55 , \AES_ENC/u0/N54 ,\AES_ENC/u0/N53 , \AES_ENC/u0/N52 , \AES_ENC/u0/N51 ,\AES_ENC/u0/N50 , \AES_ENC/u0/N49 , \AES_ENC/u0/N48 ,\AES_ENC/u0/N47 , \AES_ENC/u0/N46 , \AES_ENC/u0/N45 ,\AES_ENC/u0/N44 , \AES_ENC/u0/N43 , \AES_ENC/u0/N42 ,\AES_ENC/u0/N17 , \AES_ENC/u0/N16 , \AES_ENC/u0/N15 ,\AES_ENC/u0/N14 , \AES_ENC/u0/N13 , \AES_ENC/u0/N12 ,\AES_ENC/u0/N11 , \AES_ENC/u0/N10 , \AES_ENC/u0/subword[0] ,\AES_ENC/u0/subword[1] , \AES_ENC/u0/subword[2] ,\AES_ENC/u0/subword[3] , \AES_ENC/u0/subword[4] ,\AES_ENC/u0/subword[5] , \AES_ENC/u0/subword[6] ,\AES_ENC/u0/subword[7] , \AES_ENC/u0/subword[8] ,\AES_ENC/u0/subword[9] , \AES_ENC/u0/subword[10] ,\AES_ENC/u0/subword[11] , \AES_ENC/u0/subword[12] ,\AES_ENC/u0/subword[13] , \AES_ENC/u0/subword[14] ,\AES_ENC/u0/subword[15] , \AES_ENC/u0/subword[16] ,\AES_ENC/u0/subword[17] , \AES_ENC/u0/subword[18] ,\AES_ENC/u0/subword[19] , \AES_ENC/u0/subword[20] ,\AES_ENC/u0/subword[21] , \AES_ENC/u0/subword[22] ,\AES_ENC/u0/subword[23] , \AES_ENC/u0/subword[24] ,\AES_ENC/u0/subword[25] , \AES_ENC/u0/subword[26] ,\AES_ENC/u0/subword[27] , \AES_ENC/u0/subword[28] ,\AES_ENC/u0/subword[29] , \AES_ENC/u0/subword[30] ,\AES_ENC/u0/subword[31] , \AES_ENC/u0/u0/n1135 ,\AES_ENC/u0/u0/n1134 , \AES_ENC/u0/u0/n1133 , \AES_ENC/u0/u0/n1132 ,\AES_ENC/u0/u0/n1131 , \AES_ENC/u0/u0/n1130 , \AES_ENC/u0/u0/n1129 ,\AES_ENC/u0/u0/n1128 , \AES_ENC/u0/u0/n1127 , \AES_ENC/u0/u0/n1126 ,\AES_ENC/u0/u0/n1125 , \AES_ENC/u0/u0/n1124 , \AES_ENC/u0/u0/n1123 ,\AES_ENC/u0/u0/n1122 , \AES_ENC/u0/u0/n1121 , \AES_ENC/u0/u0/n1120 ,\AES_ENC/u0/u0/n1119 , \AES_ENC/u0/u0/n1118 , \AES_ENC/u0/u0/n1117 ,\AES_ENC/u0/u0/n1116 , \AES_ENC/u0/u0/n1115 , \AES_ENC/u0/u0/n1114 ,\AES_ENC/u0/u0/n1113 , \AES_ENC/u0/u0/n1112 , \AES_ENC/u0/u0/n1111 ,\AES_ENC/u0/u0/n1110 , \AES_ENC/u0/u0/n1109 , \AES_ENC/u0/u0/n1108 ,\AES_ENC/u0/u0/n1107 , \AES_ENC/u0/u0/n1106 , \AES_ENC/u0/u0/n1105 ,\AES_ENC/u0/u0/n1104 , \AES_ENC/u0/u0/n1103 , \AES_ENC/u0/u0/n1102 ,\AES_ENC/u0/u0/n1101 , \AES_ENC/u0/u0/n1100 , \AES_ENC/u0/u0/n1099 ,\AES_ENC/u0/u0/n1098 , \AES_ENC/u0/u0/n1097 , \AES_ENC/u0/u0/n1096 ,\AES_ENC/u0/u0/n1095 , \AES_ENC/u0/u0/n1094 , \AES_ENC/u0/u0/n1093 ,\AES_ENC/u0/u0/n1092 , \AES_ENC/u0/u0/n1091 , \AES_ENC/u0/u0/n1090 ,\AES_ENC/u0/u0/n1089 , \AES_ENC/u0/u0/n1088 , \AES_ENC/u0/u0/n1087 ,\AES_ENC/u0/u0/n1086 , \AES_ENC/u0/u0/n1085 , \AES_ENC/u0/u0/n1084 ,\AES_ENC/u0/u0/n1083 , \AES_ENC/u0/u0/n1082 , \AES_ENC/u0/u0/n1081 ,\AES_ENC/u0/u0/n1080 , \AES_ENC/u0/u0/n1079 , \AES_ENC/u0/u0/n1078 ,\AES_ENC/u0/u0/n1077 , \AES_ENC/u0/u0/n1076 , \AES_ENC/u0/u0/n1075 ,\AES_ENC/u0/u0/n1074 , \AES_ENC/u0/u0/n1073 , \AES_ENC/u0/u0/n1072 ,\AES_ENC/u0/u0/n1071 , \AES_ENC/u0/u0/n1070 , \AES_ENC/u0/u0/n1069 ,\AES_ENC/u0/u0/n1068 , \AES_ENC/u0/u0/n1067 , \AES_ENC/u0/u0/n1066 ,\AES_ENC/u0/u0/n1065 , \AES_ENC/u0/u0/n1064 , \AES_ENC/u0/u0/n1063 ,\AES_ENC/u0/u0/n1062 , \AES_ENC/u0/u0/n1061 , \AES_ENC/u0/u0/n1060 ,\AES_ENC/u0/u0/n1059 , \AES_ENC/u0/u0/n1058 , \AES_ENC/u0/u0/n1057 ,\AES_ENC/u0/u0/n1056 , \AES_ENC/u0/u0/n1055 , \AES_ENC/u0/u0/n1054 ,\AES_ENC/u0/u0/n1053 , \AES_ENC/u0/u0/n1052 , \AES_ENC/u0/u0/n1051 ,\AES_ENC/u0/u0/n1050 , \AES_ENC/u0/u0/n1049 , \AES_ENC/u0/u0/n1048 ,\AES_ENC/u0/u0/n1047 , \AES_ENC/u0/u0/n1046 , \AES_ENC/u0/u0/n1045 ,\AES_ENC/u0/u0/n1044 , \AES_ENC/u0/u0/n1043 , \AES_ENC/u0/u0/n1042 ,\AES_ENC/u0/u0/n1041 , \AES_ENC/u0/u0/n1040 , \AES_ENC/u0/u0/n1039 ,\AES_ENC/u0/u0/n1038 , \AES_ENC/u0/u0/n1037 , \AES_ENC/u0/u0/n1036 ,\AES_ENC/u0/u0/n1035 , \AES_ENC/u0/u0/n1034 , \AES_ENC/u0/u0/n1033 ,\AES_ENC/u0/u0/n1032 , \AES_ENC/u0/u0/n1031 , \AES_ENC/u0/u0/n1030 ,\AES_ENC/u0/u0/n1029 , \AES_ENC/u0/u0/n1028 , \AES_ENC/u0/u0/n1027 ,\AES_ENC/u0/u0/n1026 , \AES_ENC/u0/u0/n1025 , \AES_ENC/u0/u0/n1024 ,\AES_ENC/u0/u0/n1023 , \AES_ENC/u0/u0/n1022 , \AES_ENC/u0/u0/n1021 ,\AES_ENC/u0/u0/n1020 , \AES_ENC/u0/u0/n1019 , \AES_ENC/u0/u0/n1018 ,\AES_ENC/u0/u0/n1017 , \AES_ENC/u0/u0/n1016 , \AES_ENC/u0/u0/n1015 ,\AES_ENC/u0/u0/n1014 , \AES_ENC/u0/u0/n1013 , \AES_ENC/u0/u0/n1012 ,\AES_ENC/u0/u0/n1011 , \AES_ENC/u0/u0/n1010 , \AES_ENC/u0/u0/n1009 ,\AES_ENC/u0/u0/n1008 , \AES_ENC/u0/u0/n1007 , \AES_ENC/u0/u0/n1006 ,\AES_ENC/u0/u0/n1005 , \AES_ENC/u0/u0/n1004 , \AES_ENC/u0/u0/n1003 ,\AES_ENC/u0/u0/n1002 , \AES_ENC/u0/u0/n1001 , \AES_ENC/u0/u0/n1000 ,\AES_ENC/u0/u0/n999 , \AES_ENC/u0/u0/n998 , \AES_ENC/u0/u0/n997 ,\AES_ENC/u0/u0/n996 , \AES_ENC/u0/u0/n995 , \AES_ENC/u0/u0/n994 ,\AES_ENC/u0/u0/n993 , \AES_ENC/u0/u0/n992 , \AES_ENC/u0/u0/n991 ,\AES_ENC/u0/u0/n990 , \AES_ENC/u0/u0/n989 , \AES_ENC/u0/u0/n988 ,\AES_ENC/u0/u0/n987 , \AES_ENC/u0/u0/n986 , \AES_ENC/u0/u0/n985 ,\AES_ENC/u0/u0/n984 , \AES_ENC/u0/u0/n983 , \AES_ENC/u0/u0/n982 ,\AES_ENC/u0/u0/n981 , \AES_ENC/u0/u0/n980 , \AES_ENC/u0/u0/n979 ,\AES_ENC/u0/u0/n978 , \AES_ENC/u0/u0/n977 , \AES_ENC/u0/u0/n976 ,\AES_ENC/u0/u0/n975 , \AES_ENC/u0/u0/n974 , \AES_ENC/u0/u0/n973 ,\AES_ENC/u0/u0/n972 , \AES_ENC/u0/u0/n971 , \AES_ENC/u0/u0/n970 ,\AES_ENC/u0/u0/n969 , \AES_ENC/u0/u0/n968 , \AES_ENC/u0/u0/n967 ,\AES_ENC/u0/u0/n966 , \AES_ENC/u0/u0/n965 , \AES_ENC/u0/u0/n964 ,\AES_ENC/u0/u0/n963 , \AES_ENC/u0/u0/n962 , \AES_ENC/u0/u0/n961 ,\AES_ENC/u0/u0/n960 , \AES_ENC/u0/u0/n959 , \AES_ENC/u0/u0/n958 ,\AES_ENC/u0/u0/n957 , \AES_ENC/u0/u0/n956 , \AES_ENC/u0/u0/n955 ,\AES_ENC/u0/u0/n954 , \AES_ENC/u0/u0/n953 , \AES_ENC/u0/u0/n952 ,\AES_ENC/u0/u0/n951 , \AES_ENC/u0/u0/n950 , \AES_ENC/u0/u0/n949 ,\AES_ENC/u0/u0/n948 , \AES_ENC/u0/u0/n947 , \AES_ENC/u0/u0/n946 ,\AES_ENC/u0/u0/n945 , \AES_ENC/u0/u0/n944 , \AES_ENC/u0/u0/n943 ,\AES_ENC/u0/u0/n942 , \AES_ENC/u0/u0/n941 , \AES_ENC/u0/u0/n940 ,\AES_ENC/u0/u0/n939 , \AES_ENC/u0/u0/n938 , \AES_ENC/u0/u0/n937 ,\AES_ENC/u0/u0/n936 , \AES_ENC/u0/u0/n935 , \AES_ENC/u0/u0/n934 ,\AES_ENC/u0/u0/n933 , \AES_ENC/u0/u0/n932 , \AES_ENC/u0/u0/n931 ,\AES_ENC/u0/u0/n930 , \AES_ENC/u0/u0/n929 , \AES_ENC/u0/u0/n928 ,\AES_ENC/u0/u0/n927 , \AES_ENC/u0/u0/n926 , \AES_ENC/u0/u0/n925 ,\AES_ENC/u0/u0/n924 , \AES_ENC/u0/u0/n923 , \AES_ENC/u0/u0/n922 ,\AES_ENC/u0/u0/n921 , \AES_ENC/u0/u0/n920 , \AES_ENC/u0/u0/n919 ,\AES_ENC/u0/u0/n918 , \AES_ENC/u0/u0/n917 , \AES_ENC/u0/u0/n916 ,\AES_ENC/u0/u0/n915 , \AES_ENC/u0/u0/n914 , \AES_ENC/u0/u0/n913 ,\AES_ENC/u0/u0/n912 , \AES_ENC/u0/u0/n911 , \AES_ENC/u0/u0/n910 ,\AES_ENC/u0/u0/n909 , \AES_ENC/u0/u0/n908 , \AES_ENC/u0/u0/n907 ,\AES_ENC/u0/u0/n906 , \AES_ENC/u0/u0/n905 , \AES_ENC/u0/u0/n904 ,\AES_ENC/u0/u0/n903 , \AES_ENC/u0/u0/n902 , \AES_ENC/u0/u0/n901 ,\AES_ENC/u0/u0/n900 , \AES_ENC/u0/u0/n899 , \AES_ENC/u0/u0/n898 ,\AES_ENC/u0/u0/n897 , \AES_ENC/u0/u0/n896 , \AES_ENC/u0/u0/n895 ,\AES_ENC/u0/u0/n894 , \AES_ENC/u0/u0/n893 , \AES_ENC/u0/u0/n892 ,\AES_ENC/u0/u0/n891 , \AES_ENC/u0/u0/n890 , \AES_ENC/u0/u0/n889 ,\AES_ENC/u0/u0/n888 , \AES_ENC/u0/u0/n887 , \AES_ENC/u0/u0/n886 ,\AES_ENC/u0/u0/n885 , \AES_ENC/u0/u0/n884 , \AES_ENC/u0/u0/n883 ,\AES_ENC/u0/u0/n882 , \AES_ENC/u0/u0/n881 , \AES_ENC/u0/u0/n880 ,\AES_ENC/u0/u0/n879 , \AES_ENC/u0/u0/n878 , \AES_ENC/u0/u0/n877 ,\AES_ENC/u0/u0/n876 , \AES_ENC/u0/u0/n875 , \AES_ENC/u0/u0/n874 ,\AES_ENC/u0/u0/n873 , \AES_ENC/u0/u0/n872 , \AES_ENC/u0/u0/n871 ,\AES_ENC/u0/u0/n870 , \AES_ENC/u0/u0/n869 , \AES_ENC/u0/u0/n868 ,\AES_ENC/u0/u0/n867 , \AES_ENC/u0/u0/n866 , \AES_ENC/u0/u0/n865 ,\AES_ENC/u0/u0/n864 , \AES_ENC/u0/u0/n863 , \AES_ENC/u0/u0/n862 ,\AES_ENC/u0/u0/n861 , \AES_ENC/u0/u0/n860 , \AES_ENC/u0/u0/n859 ,\AES_ENC/u0/u0/n858 , \AES_ENC/u0/u0/n857 , \AES_ENC/u0/u0/n856 ,\AES_ENC/u0/u0/n855 , \AES_ENC/u0/u0/n854 , \AES_ENC/u0/u0/n853 ,\AES_ENC/u0/u0/n852 , \AES_ENC/u0/u0/n851 , \AES_ENC/u0/u0/n850 ,\AES_ENC/u0/u0/n849 , \AES_ENC/u0/u0/n848 , \AES_ENC/u0/u0/n847 ,\AES_ENC/u0/u0/n846 , \AES_ENC/u0/u0/n845 , \AES_ENC/u0/u0/n844 ,\AES_ENC/u0/u0/n843 , \AES_ENC/u0/u0/n842 , \AES_ENC/u0/u0/n841 ,\AES_ENC/u0/u0/n840 , \AES_ENC/u0/u0/n839 , \AES_ENC/u0/u0/n838 ,\AES_ENC/u0/u0/n837 , \AES_ENC/u0/u0/n836 , \AES_ENC/u0/u0/n835 ,\AES_ENC/u0/u0/n834 , \AES_ENC/u0/u0/n833 , \AES_ENC/u0/u0/n832 ,\AES_ENC/u0/u0/n831 , \AES_ENC/u0/u0/n830 , \AES_ENC/u0/u0/n829 ,\AES_ENC/u0/u0/n828 , \AES_ENC/u0/u0/n827 , \AES_ENC/u0/u0/n826 ,\AES_ENC/u0/u0/n825 , \AES_ENC/u0/u0/n824 , \AES_ENC/u0/u0/n823 ,\AES_ENC/u0/u0/n822 , \AES_ENC/u0/u0/n821 , \AES_ENC/u0/u0/n820 ,\AES_ENC/u0/u0/n819 , \AES_ENC/u0/u0/n818 , \AES_ENC/u0/u0/n817 ,\AES_ENC/u0/u0/n816 , \AES_ENC/u0/u0/n815 , \AES_ENC/u0/u0/n814 ,\AES_ENC/u0/u0/n813 , \AES_ENC/u0/u0/n812 , \AES_ENC/u0/u0/n811 ,\AES_ENC/u0/u0/n810 , \AES_ENC/u0/u0/n809 , \AES_ENC/u0/u0/n808 ,\AES_ENC/u0/u0/n807 , \AES_ENC/u0/u0/n806 , \AES_ENC/u0/u0/n805 ,\AES_ENC/u0/u0/n804 , \AES_ENC/u0/u0/n803 , \AES_ENC/u0/u0/n802 ,\AES_ENC/u0/u0/n801 , \AES_ENC/u0/u0/n800 , \AES_ENC/u0/u0/n799 ,\AES_ENC/u0/u0/n798 , \AES_ENC/u0/u0/n797 , \AES_ENC/u0/u0/n796 ,\AES_ENC/u0/u0/n795 , \AES_ENC/u0/u0/n794 , \AES_ENC/u0/u0/n793 ,\AES_ENC/u0/u0/n792 , \AES_ENC/u0/u0/n791 , \AES_ENC/u0/u0/n790 ,\AES_ENC/u0/u0/n789 , \AES_ENC/u0/u0/n788 , \AES_ENC/u0/u0/n787 ,\AES_ENC/u0/u0/n786 , \AES_ENC/u0/u0/n785 , \AES_ENC/u0/u0/n784 ,\AES_ENC/u0/u0/n783 , \AES_ENC/u0/u0/n782 , \AES_ENC/u0/u0/n781 ,\AES_ENC/u0/u0/n780 , \AES_ENC/u0/u0/n779 , \AES_ENC/u0/u0/n778 ,\AES_ENC/u0/u0/n777 , \AES_ENC/u0/u0/n776 , \AES_ENC/u0/u0/n775 ,\AES_ENC/u0/u0/n774 , \AES_ENC/u0/u0/n773 , \AES_ENC/u0/u0/n772 ,\AES_ENC/u0/u0/n771 , \AES_ENC/u0/u0/n770 , \AES_ENC/u0/u0/n769 ,\AES_ENC/u0/u0/n768 , \AES_ENC/u0/u0/n767 , \AES_ENC/u0/u0/n766 ,\AES_ENC/u0/u0/n765 , \AES_ENC/u0/u0/n764 , \AES_ENC/u0/u0/n763 ,\AES_ENC/u0/u0/n762 , \AES_ENC/u0/u0/n761 , \AES_ENC/u0/u0/n760 ,\AES_ENC/u0/u0/n759 , \AES_ENC/u0/u0/n758 , \AES_ENC/u0/u0/n757 ,\AES_ENC/u0/u0/n756 , \AES_ENC/u0/u0/n755 , \AES_ENC/u0/u0/n754 ,\AES_ENC/u0/u0/n753 , \AES_ENC/u0/u0/n752 , \AES_ENC/u0/u0/n751 ,\AES_ENC/u0/u0/n750 , \AES_ENC/u0/u0/n749 , \AES_ENC/u0/u0/n748 ,\AES_ENC/u0/u0/n747 , \AES_ENC/u0/u0/n746 , \AES_ENC/u0/u0/n745 ,\AES_ENC/u0/u0/n744 , \AES_ENC/u0/u0/n743 , \AES_ENC/u0/u0/n742 ,\AES_ENC/u0/u0/n741 , \AES_ENC/u0/u0/n740 , \AES_ENC/u0/u0/n739 ,\AES_ENC/u0/u0/n738 , \AES_ENC/u0/u0/n737 , \AES_ENC/u0/u0/n736 ,\AES_ENC/u0/u0/n735 , \AES_ENC/u0/u0/n734 , \AES_ENC/u0/u0/n733 ,\AES_ENC/u0/u0/n732 , \AES_ENC/u0/u0/n731 , \AES_ENC/u0/u0/n730 ,\AES_ENC/u0/u0/n729 , \AES_ENC/u0/u0/n728 , \AES_ENC/u0/u0/n727 ,\AES_ENC/u0/u0/n726 , \AES_ENC/u0/u0/n725 , \AES_ENC/u0/u0/n724 ,\AES_ENC/u0/u0/n723 , \AES_ENC/u0/u0/n722 , \AES_ENC/u0/u0/n721 ,\AES_ENC/u0/u0/n720 , \AES_ENC/u0/u0/n719 , \AES_ENC/u0/u0/n718 ,\AES_ENC/u0/u0/n717 , \AES_ENC/u0/u0/n716 , \AES_ENC/u0/u0/n715 ,\AES_ENC/u0/u0/n714 , \AES_ENC/u0/u0/n713 , \AES_ENC/u0/u0/n712 ,\AES_ENC/u0/u0/n711 , \AES_ENC/u0/u0/n710 , \AES_ENC/u0/u0/n709 ,\AES_ENC/u0/u0/n708 , \AES_ENC/u0/u0/n707 , \AES_ENC/u0/u0/n706 ,\AES_ENC/u0/u0/n705 , \AES_ENC/u0/u0/n704 , \AES_ENC/u0/u0/n703 ,\AES_ENC/u0/u0/n702 , \AES_ENC/u0/u0/n701 , \AES_ENC/u0/u0/n700 ,\AES_ENC/u0/u0/n699 , \AES_ENC/u0/u0/n698 , \AES_ENC/u0/u0/n697 ,\AES_ENC/u0/u0/n696 , \AES_ENC/u0/u0/n695 , \AES_ENC/u0/u0/n694 ,\AES_ENC/u0/u0/n693 , \AES_ENC/u0/u0/n692 , \AES_ENC/u0/u0/n691 ,\AES_ENC/u0/u0/n690 , \AES_ENC/u0/u0/n689 , \AES_ENC/u0/u0/n688 ,\AES_ENC/u0/u0/n687 , \AES_ENC/u0/u0/n686 , \AES_ENC/u0/u0/n685 ,\AES_ENC/u0/u0/n684 , \AES_ENC/u0/u0/n683 , \AES_ENC/u0/u0/n682 ,\AES_ENC/u0/u0/n681 , \AES_ENC/u0/u0/n680 , \AES_ENC/u0/u0/n679 ,\AES_ENC/u0/u0/n678 , \AES_ENC/u0/u0/n677 , \AES_ENC/u0/u0/n676 ,\AES_ENC/u0/u0/n675 , \AES_ENC/u0/u0/n674 , \AES_ENC/u0/u0/n673 ,\AES_ENC/u0/u0/n672 , \AES_ENC/u0/u0/n671 , \AES_ENC/u0/u0/n670 ,\AES_ENC/u0/u0/n669 , \AES_ENC/u0/u0/n668 , \AES_ENC/u0/u0/n667 ,\AES_ENC/u0/u0/n666 , \AES_ENC/u0/u0/n665 , \AES_ENC/u0/u0/n664 ,\AES_ENC/u0/u0/n663 , \AES_ENC/u0/u0/n662 , \AES_ENC/u0/u0/n661 ,\AES_ENC/u0/u0/n660 , \AES_ENC/u0/u0/n659 , \AES_ENC/u0/u0/n658 ,\AES_ENC/u0/u0/n657 , \AES_ENC/u0/u0/n656 , \AES_ENC/u0/u0/n655 ,\AES_ENC/u0/u0/n654 , \AES_ENC/u0/u0/n653 , \AES_ENC/u0/u0/n652 ,\AES_ENC/u0/u0/n651 , \AES_ENC/u0/u0/n650 , \AES_ENC/u0/u0/n649 ,\AES_ENC/u0/u0/n648 , \AES_ENC/u0/u0/n647 , \AES_ENC/u0/u0/n646 ,\AES_ENC/u0/u0/n645 , \AES_ENC/u0/u0/n644 , \AES_ENC/u0/u0/n643 ,\AES_ENC/u0/u0/n642 , \AES_ENC/u0/u0/n641 , \AES_ENC/u0/u0/n640 ,\AES_ENC/u0/u0/n639 , \AES_ENC/u0/u0/n638 , \AES_ENC/u0/u0/n637 ,\AES_ENC/u0/u0/n636 , \AES_ENC/u0/u0/n635 , \AES_ENC/u0/u0/n634 ,\AES_ENC/u0/u0/n633 , \AES_ENC/u0/u0/n632 , \AES_ENC/u0/u0/n631 ,\AES_ENC/u0/u0/n630 , \AES_ENC/u0/u0/n629 , \AES_ENC/u0/u0/n628 ,\AES_ENC/u0/u0/n627 , \AES_ENC/u0/u0/n626 , \AES_ENC/u0/u0/n625 ,\AES_ENC/u0/u0/n624 , \AES_ENC/u0/u0/n623 , \AES_ENC/u0/u0/n622 ,\AES_ENC/u0/u0/n621 , \AES_ENC/u0/u0/n620 , \AES_ENC/u0/u0/n619 ,\AES_ENC/u0/u0/n618 , \AES_ENC/u0/u0/n617 , \AES_ENC/u0/u0/n616 ,\AES_ENC/u0/u0/n615 , \AES_ENC/u0/u0/n614 , \AES_ENC/u0/u0/n613 ,\AES_ENC/u0/u0/n612 , \AES_ENC/u0/u0/n611 , \AES_ENC/u0/u0/n610 ,\AES_ENC/u0/u0/n609 , \AES_ENC/u0/u0/n608 , \AES_ENC/u0/u0/n607 ,\AES_ENC/u0/u0/n606 , \AES_ENC/u0/u0/n605 , \AES_ENC/u0/u0/n604 ,\AES_ENC/u0/u0/n603 , \AES_ENC/u0/u0/n602 , \AES_ENC/u0/u0/n601 ,\AES_ENC/u0/u0/n600 , \AES_ENC/u0/u0/n599 , \AES_ENC/u0/u0/n598 ,\AES_ENC/u0/u0/n597 , \AES_ENC/u0/u0/n596 , \AES_ENC/u0/u0/n595 ,\AES_ENC/u0/u0/n594 , \AES_ENC/u0/u0/n593 , \AES_ENC/u0/u0/n592 ,\AES_ENC/u0/u0/n591 , \AES_ENC/u0/u0/n590 , \AES_ENC/u0/u0/n589 ,\AES_ENC/u0/u0/n588 , \AES_ENC/u0/u0/n587 , \AES_ENC/u0/u0/n586 ,\AES_ENC/u0/u0/n585 , \AES_ENC/u0/u0/n584 , \AES_ENC/u0/u0/n583 ,\AES_ENC/u0/u0/n582 , \AES_ENC/u0/u0/n581 , \AES_ENC/u0/u0/n580 ,\AES_ENC/u0/u0/n579 , \AES_ENC/u0/u0/n578 , \AES_ENC/u0/u0/n577 ,\AES_ENC/u0/u0/n576 , \AES_ENC/u0/u0/n575 , \AES_ENC/u0/u0/n574 ,\AES_ENC/u0/u0/n573 , \AES_ENC/u0/u0/n572 , \AES_ENC/u0/u0/n571 ,\AES_ENC/u0/u0/n570 , \AES_ENC/u0/u0/n569 , \AES_ENC/u0/u1/n1135 ,\AES_ENC/u0/u1/n1134 , \AES_ENC/u0/u1/n1133 , \AES_ENC/u0/u1/n1132 ,\AES_ENC/u0/u1/n1131 , \AES_ENC/u0/u1/n1130 , \AES_ENC/u0/u1/n1129 ,\AES_ENC/u0/u1/n1128 , \AES_ENC/u0/u1/n1127 , \AES_ENC/u0/u1/n1126 ,\AES_ENC/u0/u1/n1125 , \AES_ENC/u0/u1/n1124 , \AES_ENC/u0/u1/n1123 ,\AES_ENC/u0/u1/n1122 , \AES_ENC/u0/u1/n1121 , \AES_ENC/u0/u1/n1120 ,\AES_ENC/u0/u1/n1119 , \AES_ENC/u0/u1/n1118 , \AES_ENC/u0/u1/n1117 ,\AES_ENC/u0/u1/n1116 , \AES_ENC/u0/u1/n1115 , \AES_ENC/u0/u1/n1114 ,\AES_ENC/u0/u1/n1113 , \AES_ENC/u0/u1/n1112 , \AES_ENC/u0/u1/n1111 ,\AES_ENC/u0/u1/n1110 , \AES_ENC/u0/u1/n1109 , \AES_ENC/u0/u1/n1108 ,\AES_ENC/u0/u1/n1107 , \AES_ENC/u0/u1/n1106 , \AES_ENC/u0/u1/n1105 ,\AES_ENC/u0/u1/n1104 , \AES_ENC/u0/u1/n1103 , \AES_ENC/u0/u1/n1102 ,\AES_ENC/u0/u1/n1101 , \AES_ENC/u0/u1/n1100 , \AES_ENC/u0/u1/n1099 ,\AES_ENC/u0/u1/n1098 , \AES_ENC/u0/u1/n1097 , \AES_ENC/u0/u1/n1096 ,\AES_ENC/u0/u1/n1095 , \AES_ENC/u0/u1/n1094 , \AES_ENC/u0/u1/n1093 ,\AES_ENC/u0/u1/n1092 , \AES_ENC/u0/u1/n1091 , \AES_ENC/u0/u1/n1090 ,\AES_ENC/u0/u1/n1089 , \AES_ENC/u0/u1/n1088 , \AES_ENC/u0/u1/n1087 ,\AES_ENC/u0/u1/n1086 , \AES_ENC/u0/u1/n1085 , \AES_ENC/u0/u1/n1084 ,\AES_ENC/u0/u1/n1083 , \AES_ENC/u0/u1/n1082 , \AES_ENC/u0/u1/n1081 ,\AES_ENC/u0/u1/n1080 , \AES_ENC/u0/u1/n1079 , \AES_ENC/u0/u1/n1078 ,\AES_ENC/u0/u1/n1077 , \AES_ENC/u0/u1/n1076 , \AES_ENC/u0/u1/n1075 ,\AES_ENC/u0/u1/n1074 , \AES_ENC/u0/u1/n1073 , \AES_ENC/u0/u1/n1072 ,\AES_ENC/u0/u1/n1071 , \AES_ENC/u0/u1/n1070 , \AES_ENC/u0/u1/n1069 ,\AES_ENC/u0/u1/n1068 , \AES_ENC/u0/u1/n1067 , \AES_ENC/u0/u1/n1066 ,\AES_ENC/u0/u1/n1065 , \AES_ENC/u0/u1/n1064 , \AES_ENC/u0/u1/n1063 ,\AES_ENC/u0/u1/n1062 , \AES_ENC/u0/u1/n1061 , \AES_ENC/u0/u1/n1060 ,\AES_ENC/u0/u1/n1059 , \AES_ENC/u0/u1/n1058 , \AES_ENC/u0/u1/n1057 ,\AES_ENC/u0/u1/n1056 , \AES_ENC/u0/u1/n1055 , \AES_ENC/u0/u1/n1054 ,\AES_ENC/u0/u1/n1053 , \AES_ENC/u0/u1/n1052 , \AES_ENC/u0/u1/n1051 ,\AES_ENC/u0/u1/n1050 , \AES_ENC/u0/u1/n1049 , \AES_ENC/u0/u1/n1048 ,\AES_ENC/u0/u1/n1047 , \AES_ENC/u0/u1/n1046 , \AES_ENC/u0/u1/n1045 ,\AES_ENC/u0/u1/n1044 , \AES_ENC/u0/u1/n1043 , \AES_ENC/u0/u1/n1042 ,\AES_ENC/u0/u1/n1041 , \AES_ENC/u0/u1/n1040 , \AES_ENC/u0/u1/n1039 ,\AES_ENC/u0/u1/n1038 , \AES_ENC/u0/u1/n1037 , \AES_ENC/u0/u1/n1036 ,\AES_ENC/u0/u1/n1035 , \AES_ENC/u0/u1/n1034 , \AES_ENC/u0/u1/n1033 ,\AES_ENC/u0/u1/n1032 , \AES_ENC/u0/u1/n1031 , \AES_ENC/u0/u1/n1030 ,\AES_ENC/u0/u1/n1029 , \AES_ENC/u0/u1/n1028 , \AES_ENC/u0/u1/n1027 ,\AES_ENC/u0/u1/n1026 , \AES_ENC/u0/u1/n1025 , \AES_ENC/u0/u1/n1024 ,\AES_ENC/u0/u1/n1023 , \AES_ENC/u0/u1/n1022 , \AES_ENC/u0/u1/n1021 ,\AES_ENC/u0/u1/n1020 , \AES_ENC/u0/u1/n1019 , \AES_ENC/u0/u1/n1018 ,\AES_ENC/u0/u1/n1017 , \AES_ENC/u0/u1/n1016 , \AES_ENC/u0/u1/n1015 ,\AES_ENC/u0/u1/n1014 , \AES_ENC/u0/u1/n1013 , \AES_ENC/u0/u1/n1012 ,\AES_ENC/u0/u1/n1011 , \AES_ENC/u0/u1/n1010 , \AES_ENC/u0/u1/n1009 ,\AES_ENC/u0/u1/n1008 , \AES_ENC/u0/u1/n1007 , \AES_ENC/u0/u1/n1006 ,\AES_ENC/u0/u1/n1005 , \AES_ENC/u0/u1/n1004 , \AES_ENC/u0/u1/n1003 ,\AES_ENC/u0/u1/n1002 , \AES_ENC/u0/u1/n1001 , \AES_ENC/u0/u1/n1000 ,\AES_ENC/u0/u1/n999 , \AES_ENC/u0/u1/n998 , \AES_ENC/u0/u1/n997 ,\AES_ENC/u0/u1/n996 , \AES_ENC/u0/u1/n995 , \AES_ENC/u0/u1/n994 ,\AES_ENC/u0/u1/n993 , \AES_ENC/u0/u1/n992 , \AES_ENC/u0/u1/n991 ,\AES_ENC/u0/u1/n990 , \AES_ENC/u0/u1/n989 , \AES_ENC/u0/u1/n988 ,\AES_ENC/u0/u1/n987 , \AES_ENC/u0/u1/n986 , \AES_ENC/u0/u1/n985 ,\AES_ENC/u0/u1/n984 , \AES_ENC/u0/u1/n983 , \AES_ENC/u0/u1/n982 ,\AES_ENC/u0/u1/n981 , \AES_ENC/u0/u1/n980 , \AES_ENC/u0/u1/n979 ,\AES_ENC/u0/u1/n978 , \AES_ENC/u0/u1/n977 , \AES_ENC/u0/u1/n976 ,\AES_ENC/u0/u1/n975 , \AES_ENC/u0/u1/n974 , \AES_ENC/u0/u1/n973 ,\AES_ENC/u0/u1/n972 , \AES_ENC/u0/u1/n971 , \AES_ENC/u0/u1/n970 ,\AES_ENC/u0/u1/n969 , \AES_ENC/u0/u1/n968 , \AES_ENC/u0/u1/n967 ,\AES_ENC/u0/u1/n966 , \AES_ENC/u0/u1/n965 , \AES_ENC/u0/u1/n964 ,\AES_ENC/u0/u1/n963 , \AES_ENC/u0/u1/n962 , \AES_ENC/u0/u1/n961 ,\AES_ENC/u0/u1/n960 , \AES_ENC/u0/u1/n959 , \AES_ENC/u0/u1/n958 ,\AES_ENC/u0/u1/n957 , \AES_ENC/u0/u1/n956 , \AES_ENC/u0/u1/n955 ,\AES_ENC/u0/u1/n954 , \AES_ENC/u0/u1/n953 , \AES_ENC/u0/u1/n952 ,\AES_ENC/u0/u1/n951 , \AES_ENC/u0/u1/n950 , \AES_ENC/u0/u1/n949 ,\AES_ENC/u0/u1/n948 , \AES_ENC/u0/u1/n947 , \AES_ENC/u0/u1/n946 ,\AES_ENC/u0/u1/n945 , \AES_ENC/u0/u1/n944 , \AES_ENC/u0/u1/n943 ,\AES_ENC/u0/u1/n942 , \AES_ENC/u0/u1/n941 , \AES_ENC/u0/u1/n940 ,\AES_ENC/u0/u1/n939 , \AES_ENC/u0/u1/n938 , \AES_ENC/u0/u1/n937 ,\AES_ENC/u0/u1/n936 , \AES_ENC/u0/u1/n935 , \AES_ENC/u0/u1/n934 ,\AES_ENC/u0/u1/n933 , \AES_ENC/u0/u1/n932 , \AES_ENC/u0/u1/n931 ,\AES_ENC/u0/u1/n930 , \AES_ENC/u0/u1/n929 , \AES_ENC/u0/u1/n928 ,\AES_ENC/u0/u1/n927 , \AES_ENC/u0/u1/n926 , \AES_ENC/u0/u1/n925 ,\AES_ENC/u0/u1/n924 , \AES_ENC/u0/u1/n923 , \AES_ENC/u0/u1/n922 ,\AES_ENC/u0/u1/n921 , \AES_ENC/u0/u1/n920 , \AES_ENC/u0/u1/n919 ,\AES_ENC/u0/u1/n918 , \AES_ENC/u0/u1/n917 , \AES_ENC/u0/u1/n916 ,\AES_ENC/u0/u1/n915 , \AES_ENC/u0/u1/n914 , \AES_ENC/u0/u1/n913 ,\AES_ENC/u0/u1/n912 , \AES_ENC/u0/u1/n911 , \AES_ENC/u0/u1/n910 ,\AES_ENC/u0/u1/n909 , \AES_ENC/u0/u1/n908 , \AES_ENC/u0/u1/n907 ,\AES_ENC/u0/u1/n906 , \AES_ENC/u0/u1/n905 , \AES_ENC/u0/u1/n904 ,\AES_ENC/u0/u1/n903 , \AES_ENC/u0/u1/n902 , \AES_ENC/u0/u1/n901 ,\AES_ENC/u0/u1/n900 , \AES_ENC/u0/u1/n899 , \AES_ENC/u0/u1/n898 ,\AES_ENC/u0/u1/n897 , \AES_ENC/u0/u1/n896 , \AES_ENC/u0/u1/n895 ,\AES_ENC/u0/u1/n894 , \AES_ENC/u0/u1/n893 , \AES_ENC/u0/u1/n892 ,\AES_ENC/u0/u1/n891 , \AES_ENC/u0/u1/n890 , \AES_ENC/u0/u1/n889 ,\AES_ENC/u0/u1/n888 , \AES_ENC/u0/u1/n887 , \AES_ENC/u0/u1/n886 ,\AES_ENC/u0/u1/n885 , \AES_ENC/u0/u1/n884 , \AES_ENC/u0/u1/n883 ,\AES_ENC/u0/u1/n882 , \AES_ENC/u0/u1/n881 , \AES_ENC/u0/u1/n880 ,\AES_ENC/u0/u1/n879 , \AES_ENC/u0/u1/n878 , \AES_ENC/u0/u1/n877 ,\AES_ENC/u0/u1/n876 , \AES_ENC/u0/u1/n875 , \AES_ENC/u0/u1/n874 ,\AES_ENC/u0/u1/n873 , \AES_ENC/u0/u1/n872 , \AES_ENC/u0/u1/n871 ,\AES_ENC/u0/u1/n870 , \AES_ENC/u0/u1/n869 , \AES_ENC/u0/u1/n868 ,\AES_ENC/u0/u1/n867 , \AES_ENC/u0/u1/n866 , \AES_ENC/u0/u1/n865 ,\AES_ENC/u0/u1/n864 , \AES_ENC/u0/u1/n863 , \AES_ENC/u0/u1/n862 ,\AES_ENC/u0/u1/n861 , \AES_ENC/u0/u1/n860 , \AES_ENC/u0/u1/n859 ,\AES_ENC/u0/u1/n858 , \AES_ENC/u0/u1/n857 , \AES_ENC/u0/u1/n856 ,\AES_ENC/u0/u1/n855 , \AES_ENC/u0/u1/n854 , \AES_ENC/u0/u1/n853 ,\AES_ENC/u0/u1/n852 , \AES_ENC/u0/u1/n851 , \AES_ENC/u0/u1/n850 ,\AES_ENC/u0/u1/n849 , \AES_ENC/u0/u1/n848 , \AES_ENC/u0/u1/n847 ,\AES_ENC/u0/u1/n846 , \AES_ENC/u0/u1/n845 , \AES_ENC/u0/u1/n844 ,\AES_ENC/u0/u1/n843 , \AES_ENC/u0/u1/n842 , \AES_ENC/u0/u1/n841 ,\AES_ENC/u0/u1/n840 , \AES_ENC/u0/u1/n839 , \AES_ENC/u0/u1/n838 ,\AES_ENC/u0/u1/n837 , \AES_ENC/u0/u1/n836 , \AES_ENC/u0/u1/n835 ,\AES_ENC/u0/u1/n834 , \AES_ENC/u0/u1/n833 , \AES_ENC/u0/u1/n832 ,\AES_ENC/u0/u1/n831 , \AES_ENC/u0/u1/n830 , \AES_ENC/u0/u1/n829 ,\AES_ENC/u0/u1/n828 , \AES_ENC/u0/u1/n827 , \AES_ENC/u0/u1/n826 ,\AES_ENC/u0/u1/n825 , \AES_ENC/u0/u1/n824 , \AES_ENC/u0/u1/n823 ,\AES_ENC/u0/u1/n822 , \AES_ENC/u0/u1/n821 , \AES_ENC/u0/u1/n820 ,\AES_ENC/u0/u1/n819 , \AES_ENC/u0/u1/n818 , \AES_ENC/u0/u1/n817 ,\AES_ENC/u0/u1/n816 , \AES_ENC/u0/u1/n815 , \AES_ENC/u0/u1/n814 ,\AES_ENC/u0/u1/n813 , \AES_ENC/u0/u1/n812 , \AES_ENC/u0/u1/n811 ,\AES_ENC/u0/u1/n810 , \AES_ENC/u0/u1/n809 , \AES_ENC/u0/u1/n808 ,\AES_ENC/u0/u1/n807 , \AES_ENC/u0/u1/n806 , \AES_ENC/u0/u1/n805 ,\AES_ENC/u0/u1/n804 , \AES_ENC/u0/u1/n803 , \AES_ENC/u0/u1/n802 ,\AES_ENC/u0/u1/n801 , \AES_ENC/u0/u1/n800 , \AES_ENC/u0/u1/n799 ,\AES_ENC/u0/u1/n798 , \AES_ENC/u0/u1/n797 , \AES_ENC/u0/u1/n796 ,\AES_ENC/u0/u1/n795 , \AES_ENC/u0/u1/n794 , \AES_ENC/u0/u1/n793 ,\AES_ENC/u0/u1/n792 , \AES_ENC/u0/u1/n791 , \AES_ENC/u0/u1/n790 ,\AES_ENC/u0/u1/n789 , \AES_ENC/u0/u1/n788 , \AES_ENC/u0/u1/n787 ,\AES_ENC/u0/u1/n786 , \AES_ENC/u0/u1/n785 , \AES_ENC/u0/u1/n784 ,\AES_ENC/u0/u1/n783 , \AES_ENC/u0/u1/n782 , \AES_ENC/u0/u1/n781 ,\AES_ENC/u0/u1/n780 , \AES_ENC/u0/u1/n779 , \AES_ENC/u0/u1/n778 ,\AES_ENC/u0/u1/n777 , \AES_ENC/u0/u1/n776 , \AES_ENC/u0/u1/n775 ,\AES_ENC/u0/u1/n774 , \AES_ENC/u0/u1/n773 , \AES_ENC/u0/u1/n772 ,\AES_ENC/u0/u1/n771 , \AES_ENC/u0/u1/n770 , \AES_ENC/u0/u1/n769 ,\AES_ENC/u0/u1/n768 , \AES_ENC/u0/u1/n767 , \AES_ENC/u0/u1/n766 ,\AES_ENC/u0/u1/n765 , \AES_ENC/u0/u1/n764 , \AES_ENC/u0/u1/n763 ,\AES_ENC/u0/u1/n762 , \AES_ENC/u0/u1/n761 , \AES_ENC/u0/u1/n760 ,\AES_ENC/u0/u1/n759 , \AES_ENC/u0/u1/n758 , \AES_ENC/u0/u1/n757 ,\AES_ENC/u0/u1/n756 , \AES_ENC/u0/u1/n755 , \AES_ENC/u0/u1/n754 ,\AES_ENC/u0/u1/n753 , \AES_ENC/u0/u1/n752 , \AES_ENC/u0/u1/n751 ,\AES_ENC/u0/u1/n750 , \AES_ENC/u0/u1/n749 , \AES_ENC/u0/u1/n748 ,\AES_ENC/u0/u1/n747 , \AES_ENC/u0/u1/n746 , \AES_ENC/u0/u1/n745 ,\AES_ENC/u0/u1/n744 , \AES_ENC/u0/u1/n743 , \AES_ENC/u0/u1/n742 ,\AES_ENC/u0/u1/n741 , \AES_ENC/u0/u1/n740 , \AES_ENC/u0/u1/n739 ,\AES_ENC/u0/u1/n738 , \AES_ENC/u0/u1/n737 , \AES_ENC/u0/u1/n736 ,\AES_ENC/u0/u1/n735 , \AES_ENC/u0/u1/n734 , \AES_ENC/u0/u1/n733 ,\AES_ENC/u0/u1/n732 , \AES_ENC/u0/u1/n731 , \AES_ENC/u0/u1/n730 ,\AES_ENC/u0/u1/n729 , \AES_ENC/u0/u1/n728 , \AES_ENC/u0/u1/n727 ,\AES_ENC/u0/u1/n726 , \AES_ENC/u0/u1/n725 , \AES_ENC/u0/u1/n724 ,\AES_ENC/u0/u1/n723 , \AES_ENC/u0/u1/n722 , \AES_ENC/u0/u1/n721 ,\AES_ENC/u0/u1/n720 , \AES_ENC/u0/u1/n719 , \AES_ENC/u0/u1/n718 ,\AES_ENC/u0/u1/n717 , \AES_ENC/u0/u1/n716 , \AES_ENC/u0/u1/n715 ,\AES_ENC/u0/u1/n714 , \AES_ENC/u0/u1/n713 , \AES_ENC/u0/u1/n712 ,\AES_ENC/u0/u1/n711 , \AES_ENC/u0/u1/n710 , \AES_ENC/u0/u1/n709 ,\AES_ENC/u0/u1/n708 , \AES_ENC/u0/u1/n707 , \AES_ENC/u0/u1/n706 ,\AES_ENC/u0/u1/n705 , \AES_ENC/u0/u1/n704 , \AES_ENC/u0/u1/n703 ,\AES_ENC/u0/u1/n702 , \AES_ENC/u0/u1/n701 , \AES_ENC/u0/u1/n700 ,\AES_ENC/u0/u1/n699 , \AES_ENC/u0/u1/n698 , \AES_ENC/u0/u1/n697 ,\AES_ENC/u0/u1/n696 , \AES_ENC/u0/u1/n695 , \AES_ENC/u0/u1/n694 ,\AES_ENC/u0/u1/n693 , \AES_ENC/u0/u1/n692 , \AES_ENC/u0/u1/n691 ,\AES_ENC/u0/u1/n690 , \AES_ENC/u0/u1/n689 , \AES_ENC/u0/u1/n688 ,\AES_ENC/u0/u1/n687 , \AES_ENC/u0/u1/n686 , \AES_ENC/u0/u1/n685 ,\AES_ENC/u0/u1/n684 , \AES_ENC/u0/u1/n683 , \AES_ENC/u0/u1/n682 ,\AES_ENC/u0/u1/n681 , \AES_ENC/u0/u1/n680 , \AES_ENC/u0/u1/n679 ,\AES_ENC/u0/u1/n678 , \AES_ENC/u0/u1/n677 , \AES_ENC/u0/u1/n676 ,\AES_ENC/u0/u1/n675 , \AES_ENC/u0/u1/n674 , \AES_ENC/u0/u1/n673 ,\AES_ENC/u0/u1/n672 , \AES_ENC/u0/u1/n671 , \AES_ENC/u0/u1/n670 ,\AES_ENC/u0/u1/n669 , \AES_ENC/u0/u1/n668 , \AES_ENC/u0/u1/n667 ,\AES_ENC/u0/u1/n666 , \AES_ENC/u0/u1/n665 , \AES_ENC/u0/u1/n664 ,\AES_ENC/u0/u1/n663 , \AES_ENC/u0/u1/n662 , \AES_ENC/u0/u1/n661 ,\AES_ENC/u0/u1/n660 , \AES_ENC/u0/u1/n659 , \AES_ENC/u0/u1/n658 ,\AES_ENC/u0/u1/n657 , \AES_ENC/u0/u1/n656 , \AES_ENC/u0/u1/n655 ,\AES_ENC/u0/u1/n654 , \AES_ENC/u0/u1/n653 , \AES_ENC/u0/u1/n652 ,\AES_ENC/u0/u1/n651 , \AES_ENC/u0/u1/n650 , \AES_ENC/u0/u1/n649 ,\AES_ENC/u0/u1/n648 , \AES_ENC/u0/u1/n647 , \AES_ENC/u0/u1/n646 ,\AES_ENC/u0/u1/n645 , \AES_ENC/u0/u1/n644 , \AES_ENC/u0/u1/n643 ,\AES_ENC/u0/u1/n642 , \AES_ENC/u0/u1/n641 , \AES_ENC/u0/u1/n640 ,\AES_ENC/u0/u1/n639 , \AES_ENC/u0/u1/n638 , \AES_ENC/u0/u1/n637 ,\AES_ENC/u0/u1/n636 , \AES_ENC/u0/u1/n635 , \AES_ENC/u0/u1/n634 ,\AES_ENC/u0/u1/n633 , \AES_ENC/u0/u1/n632 , \AES_ENC/u0/u1/n631 ,\AES_ENC/u0/u1/n630 , \AES_ENC/u0/u1/n629 , \AES_ENC/u0/u1/n628 ,\AES_ENC/u0/u1/n627 , \AES_ENC/u0/u1/n626 , \AES_ENC/u0/u1/n625 ,\AES_ENC/u0/u1/n624 , \AES_ENC/u0/u1/n623 , \AES_ENC/u0/u1/n622 ,\AES_ENC/u0/u1/n621 , \AES_ENC/u0/u1/n620 , \AES_ENC/u0/u1/n619 ,\AES_ENC/u0/u1/n618 , \AES_ENC/u0/u1/n617 , \AES_ENC/u0/u1/n616 ,\AES_ENC/u0/u1/n615 , \AES_ENC/u0/u1/n614 , \AES_ENC/u0/u1/n613 ,\AES_ENC/u0/u1/n612 , \AES_ENC/u0/u1/n611 , \AES_ENC/u0/u1/n610 ,\AES_ENC/u0/u1/n609 , \AES_ENC/u0/u1/n608 , \AES_ENC/u0/u1/n607 ,\AES_ENC/u0/u1/n606 , \AES_ENC/u0/u1/n605 , \AES_ENC/u0/u1/n604 ,\AES_ENC/u0/u1/n603 , \AES_ENC/u0/u1/n602 , \AES_ENC/u0/u1/n601 ,\AES_ENC/u0/u1/n600 , \AES_ENC/u0/u1/n599 , \AES_ENC/u0/u1/n598 ,\AES_ENC/u0/u1/n597 , \AES_ENC/u0/u1/n596 , \AES_ENC/u0/u1/n595 ,\AES_ENC/u0/u1/n594 , \AES_ENC/u0/u1/n593 , \AES_ENC/u0/u1/n592 ,\AES_ENC/u0/u1/n591 , \AES_ENC/u0/u1/n590 , \AES_ENC/u0/u1/n589 ,\AES_ENC/u0/u1/n588 , \AES_ENC/u0/u1/n587 , \AES_ENC/u0/u1/n586 ,\AES_ENC/u0/u1/n585 , \AES_ENC/u0/u1/n584 , \AES_ENC/u0/u1/n583 ,\AES_ENC/u0/u1/n582 , \AES_ENC/u0/u1/n581 , \AES_ENC/u0/u1/n580 ,\AES_ENC/u0/u1/n579 , \AES_ENC/u0/u1/n578 , \AES_ENC/u0/u1/n577 ,\AES_ENC/u0/u1/n576 , \AES_ENC/u0/u1/n575 , \AES_ENC/u0/u1/n574 ,\AES_ENC/u0/u1/n573 , \AES_ENC/u0/u1/n572 , \AES_ENC/u0/u1/n571 ,\AES_ENC/u0/u1/n570 , \AES_ENC/u0/u1/n569 , \AES_ENC/u0/u2/n1135 ,\AES_ENC/u0/u2/n1134 , \AES_ENC/u0/u2/n1133 , \AES_ENC/u0/u2/n1132 ,\AES_ENC/u0/u2/n1131 , \AES_ENC/u0/u2/n1130 , \AES_ENC/u0/u2/n1129 ,\AES_ENC/u0/u2/n1128 , \AES_ENC/u0/u2/n1127 , \AES_ENC/u0/u2/n1126 ,\AES_ENC/u0/u2/n1125 , \AES_ENC/u0/u2/n1124 , \AES_ENC/u0/u2/n1123 ,\AES_ENC/u0/u2/n1122 , \AES_ENC/u0/u2/n1121 , \AES_ENC/u0/u2/n1120 ,\AES_ENC/u0/u2/n1119 , \AES_ENC/u0/u2/n1118 , \AES_ENC/u0/u2/n1117 ,\AES_ENC/u0/u2/n1116 , \AES_ENC/u0/u2/n1115 , \AES_ENC/u0/u2/n1114 ,\AES_ENC/u0/u2/n1113 , \AES_ENC/u0/u2/n1112 , \AES_ENC/u0/u2/n1111 ,\AES_ENC/u0/u2/n1110 , \AES_ENC/u0/u2/n1109 , \AES_ENC/u0/u2/n1108 ,\AES_ENC/u0/u2/n1107 , \AES_ENC/u0/u2/n1106 , \AES_ENC/u0/u2/n1105 ,\AES_ENC/u0/u2/n1104 , \AES_ENC/u0/u2/n1103 , \AES_ENC/u0/u2/n1102 ,\AES_ENC/u0/u2/n1101 , \AES_ENC/u0/u2/n1100 , \AES_ENC/u0/u2/n1099 ,\AES_ENC/u0/u2/n1098 , \AES_ENC/u0/u2/n1097 , \AES_ENC/u0/u2/n1096 ,\AES_ENC/u0/u2/n1095 , \AES_ENC/u0/u2/n1094 , \AES_ENC/u0/u2/n1093 ,\AES_ENC/u0/u2/n1092 , \AES_ENC/u0/u2/n1091 , \AES_ENC/u0/u2/n1090 ,\AES_ENC/u0/u2/n1089 , \AES_ENC/u0/u2/n1088 , \AES_ENC/u0/u2/n1087 ,\AES_ENC/u0/u2/n1086 , \AES_ENC/u0/u2/n1085 , \AES_ENC/u0/u2/n1084 ,\AES_ENC/u0/u2/n1083 , \AES_ENC/u0/u2/n1082 , \AES_ENC/u0/u2/n1081 ,\AES_ENC/u0/u2/n1080 , \AES_ENC/u0/u2/n1079 , \AES_ENC/u0/u2/n1078 ,\AES_ENC/u0/u2/n1077 , \AES_ENC/u0/u2/n1076 , \AES_ENC/u0/u2/n1075 ,\AES_ENC/u0/u2/n1074 , \AES_ENC/u0/u2/n1073 , \AES_ENC/u0/u2/n1072 ,\AES_ENC/u0/u2/n1071 , \AES_ENC/u0/u2/n1070 , \AES_ENC/u0/u2/n1069 ,\AES_ENC/u0/u2/n1068 , \AES_ENC/u0/u2/n1067 , \AES_ENC/u0/u2/n1066 ,\AES_ENC/u0/u2/n1065 , \AES_ENC/u0/u2/n1064 , \AES_ENC/u0/u2/n1063 ,\AES_ENC/u0/u2/n1062 , \AES_ENC/u0/u2/n1061 , \AES_ENC/u0/u2/n1060 ,\AES_ENC/u0/u2/n1059 , \AES_ENC/u0/u2/n1058 , \AES_ENC/u0/u2/n1057 ,\AES_ENC/u0/u2/n1056 , \AES_ENC/u0/u2/n1055 , \AES_ENC/u0/u2/n1054 ,\AES_ENC/u0/u2/n1053 , \AES_ENC/u0/u2/n1052 , \AES_ENC/u0/u2/n1051 ,\AES_ENC/u0/u2/n1050 , \AES_ENC/u0/u2/n1049 , \AES_ENC/u0/u2/n1048 ,\AES_ENC/u0/u2/n1047 , \AES_ENC/u0/u2/n1046 , \AES_ENC/u0/u2/n1045 ,\AES_ENC/u0/u2/n1044 , \AES_ENC/u0/u2/n1043 , \AES_ENC/u0/u2/n1042 ,\AES_ENC/u0/u2/n1041 , \AES_ENC/u0/u2/n1040 , \AES_ENC/u0/u2/n1039 ,\AES_ENC/u0/u2/n1038 , \AES_ENC/u0/u2/n1037 , \AES_ENC/u0/u2/n1036 ,\AES_ENC/u0/u2/n1035 , \AES_ENC/u0/u2/n1034 , \AES_ENC/u0/u2/n1033 ,\AES_ENC/u0/u2/n1032 , \AES_ENC/u0/u2/n1031 , \AES_ENC/u0/u2/n1030 ,\AES_ENC/u0/u2/n1029 , \AES_ENC/u0/u2/n1028 , \AES_ENC/u0/u2/n1027 ,\AES_ENC/u0/u2/n1026 , \AES_ENC/u0/u2/n1025 , \AES_ENC/u0/u2/n1024 ,\AES_ENC/u0/u2/n1023 , \AES_ENC/u0/u2/n1022 , \AES_ENC/u0/u2/n1021 ,\AES_ENC/u0/u2/n1020 , \AES_ENC/u0/u2/n1019 , \AES_ENC/u0/u2/n1018 ,\AES_ENC/u0/u2/n1017 , \AES_ENC/u0/u2/n1016 , \AES_ENC/u0/u2/n1015 ,\AES_ENC/u0/u2/n1014 , \AES_ENC/u0/u2/n1013 , \AES_ENC/u0/u2/n1012 ,\AES_ENC/u0/u2/n1011 , \AES_ENC/u0/u2/n1010 , \AES_ENC/u0/u2/n1009 ,\AES_ENC/u0/u2/n1008 , \AES_ENC/u0/u2/n1007 , \AES_ENC/u0/u2/n1006 ,\AES_ENC/u0/u2/n1005 , \AES_ENC/u0/u2/n1004 , \AES_ENC/u0/u2/n1003 ,\AES_ENC/u0/u2/n1002 , \AES_ENC/u0/u2/n1001 , \AES_ENC/u0/u2/n1000 ,\AES_ENC/u0/u2/n999 , \AES_ENC/u0/u2/n998 , \AES_ENC/u0/u2/n997 ,\AES_ENC/u0/u2/n996 , \AES_ENC/u0/u2/n995 , \AES_ENC/u0/u2/n994 ,\AES_ENC/u0/u2/n993 , \AES_ENC/u0/u2/n992 , \AES_ENC/u0/u2/n991 ,\AES_ENC/u0/u2/n990 , \AES_ENC/u0/u2/n989 , \AES_ENC/u0/u2/n988 ,\AES_ENC/u0/u2/n987 , \AES_ENC/u0/u2/n986 , \AES_ENC/u0/u2/n985 ,\AES_ENC/u0/u2/n984 , \AES_ENC/u0/u2/n983 , \AES_ENC/u0/u2/n982 ,\AES_ENC/u0/u2/n981 , \AES_ENC/u0/u2/n980 , \AES_ENC/u0/u2/n979 ,\AES_ENC/u0/u2/n978 , \AES_ENC/u0/u2/n977 , \AES_ENC/u0/u2/n976 ,\AES_ENC/u0/u2/n975 , \AES_ENC/u0/u2/n974 , \AES_ENC/u0/u2/n973 ,\AES_ENC/u0/u2/n972 , \AES_ENC/u0/u2/n971 , \AES_ENC/u0/u2/n970 ,\AES_ENC/u0/u2/n969 , \AES_ENC/u0/u2/n968 , \AES_ENC/u0/u2/n967 ,\AES_ENC/u0/u2/n966 , \AES_ENC/u0/u2/n965 , \AES_ENC/u0/u2/n964 ,\AES_ENC/u0/u2/n963 , \AES_ENC/u0/u2/n962 , \AES_ENC/u0/u2/n961 ,\AES_ENC/u0/u2/n960 , \AES_ENC/u0/u2/n959 , \AES_ENC/u0/u2/n958 ,\AES_ENC/u0/u2/n957 , \AES_ENC/u0/u2/n956 , \AES_ENC/u0/u2/n955 ,\AES_ENC/u0/u2/n954 , \AES_ENC/u0/u2/n953 , \AES_ENC/u0/u2/n952 ,\AES_ENC/u0/u2/n951 , \AES_ENC/u0/u2/n950 , \AES_ENC/u0/u2/n949 ,\AES_ENC/u0/u2/n948 , \AES_ENC/u0/u2/n947 , \AES_ENC/u0/u2/n946 ,\AES_ENC/u0/u2/n945 , \AES_ENC/u0/u2/n944 , \AES_ENC/u0/u2/n943 ,\AES_ENC/u0/u2/n942 , \AES_ENC/u0/u2/n941 , \AES_ENC/u0/u2/n940 ,\AES_ENC/u0/u2/n939 , \AES_ENC/u0/u2/n938 , \AES_ENC/u0/u2/n937 ,\AES_ENC/u0/u2/n936 , \AES_ENC/u0/u2/n935 , \AES_ENC/u0/u2/n934 ,\AES_ENC/u0/u2/n933 , \AES_ENC/u0/u2/n932 , \AES_ENC/u0/u2/n931 ,\AES_ENC/u0/u2/n930 , \AES_ENC/u0/u2/n929 , \AES_ENC/u0/u2/n928 ,\AES_ENC/u0/u2/n927 , \AES_ENC/u0/u2/n926 , \AES_ENC/u0/u2/n925 ,\AES_ENC/u0/u2/n924 , \AES_ENC/u0/u2/n923 , \AES_ENC/u0/u2/n922 ,\AES_ENC/u0/u2/n921 , \AES_ENC/u0/u2/n920 , \AES_ENC/u0/u2/n919 ,\AES_ENC/u0/u2/n918 , \AES_ENC/u0/u2/n917 , \AES_ENC/u0/u2/n916 ,\AES_ENC/u0/u2/n915 , \AES_ENC/u0/u2/n914 , \AES_ENC/u0/u2/n913 ,\AES_ENC/u0/u2/n912 , \AES_ENC/u0/u2/n911 , \AES_ENC/u0/u2/n910 ,\AES_ENC/u0/u2/n909 , \AES_ENC/u0/u2/n908 , \AES_ENC/u0/u2/n907 ,\AES_ENC/u0/u2/n906 , \AES_ENC/u0/u2/n905 , \AES_ENC/u0/u2/n904 ,\AES_ENC/u0/u2/n903 , \AES_ENC/u0/u2/n902 , \AES_ENC/u0/u2/n901 ,\AES_ENC/u0/u2/n900 , \AES_ENC/u0/u2/n899 , \AES_ENC/u0/u2/n898 ,\AES_ENC/u0/u2/n897 , \AES_ENC/u0/u2/n896 , \AES_ENC/u0/u2/n895 ,\AES_ENC/u0/u2/n894 , \AES_ENC/u0/u2/n893 , \AES_ENC/u0/u2/n892 ,\AES_ENC/u0/u2/n891 , \AES_ENC/u0/u2/n890 , \AES_ENC/u0/u2/n889 ,\AES_ENC/u0/u2/n888 , \AES_ENC/u0/u2/n887 , \AES_ENC/u0/u2/n886 ,\AES_ENC/u0/u2/n885 , \AES_ENC/u0/u2/n884 , \AES_ENC/u0/u2/n883 ,\AES_ENC/u0/u2/n882 , \AES_ENC/u0/u2/n881 , \AES_ENC/u0/u2/n880 ,\AES_ENC/u0/u2/n879 , \AES_ENC/u0/u2/n878 , \AES_ENC/u0/u2/n877 ,\AES_ENC/u0/u2/n876 , \AES_ENC/u0/u2/n875 , \AES_ENC/u0/u2/n874 ,\AES_ENC/u0/u2/n873 , \AES_ENC/u0/u2/n872 , \AES_ENC/u0/u2/n871 ,\AES_ENC/u0/u2/n870 , \AES_ENC/u0/u2/n869 , \AES_ENC/u0/u2/n868 ,\AES_ENC/u0/u2/n867 , \AES_ENC/u0/u2/n866 , \AES_ENC/u0/u2/n865 ,\AES_ENC/u0/u2/n864 , \AES_ENC/u0/u2/n863 , \AES_ENC/u0/u2/n862 ,\AES_ENC/u0/u2/n861 , \AES_ENC/u0/u2/n860 , \AES_ENC/u0/u2/n859 ,\AES_ENC/u0/u2/n858 , \AES_ENC/u0/u2/n857 , \AES_ENC/u0/u2/n856 ,\AES_ENC/u0/u2/n855 , \AES_ENC/u0/u2/n854 , \AES_ENC/u0/u2/n853 ,\AES_ENC/u0/u2/n852 , \AES_ENC/u0/u2/n851 , \AES_ENC/u0/u2/n850 ,\AES_ENC/u0/u2/n849 , \AES_ENC/u0/u2/n848 , \AES_ENC/u0/u2/n847 ,\AES_ENC/u0/u2/n846 , \AES_ENC/u0/u2/n845 , \AES_ENC/u0/u2/n844 ,\AES_ENC/u0/u2/n843 , \AES_ENC/u0/u2/n842 , \AES_ENC/u0/u2/n841 ,\AES_ENC/u0/u2/n840 , \AES_ENC/u0/u2/n839 , \AES_ENC/u0/u2/n838 ,\AES_ENC/u0/u2/n837 , \AES_ENC/u0/u2/n836 , \AES_ENC/u0/u2/n835 ,\AES_ENC/u0/u2/n834 , \AES_ENC/u0/u2/n833 , \AES_ENC/u0/u2/n832 ,\AES_ENC/u0/u2/n831 , \AES_ENC/u0/u2/n830 , \AES_ENC/u0/u2/n829 ,\AES_ENC/u0/u2/n828 , \AES_ENC/u0/u2/n827 , \AES_ENC/u0/u2/n826 ,\AES_ENC/u0/u2/n825 , \AES_ENC/u0/u2/n824 , \AES_ENC/u0/u2/n823 ,\AES_ENC/u0/u2/n822 , \AES_ENC/u0/u2/n821 , \AES_ENC/u0/u2/n820 ,\AES_ENC/u0/u2/n819 , \AES_ENC/u0/u2/n818 , \AES_ENC/u0/u2/n817 ,\AES_ENC/u0/u2/n816 , \AES_ENC/u0/u2/n815 , \AES_ENC/u0/u2/n814 ,\AES_ENC/u0/u2/n813 , \AES_ENC/u0/u2/n812 , \AES_ENC/u0/u2/n811 ,\AES_ENC/u0/u2/n810 , \AES_ENC/u0/u2/n809 , \AES_ENC/u0/u2/n808 ,\AES_ENC/u0/u2/n807 , \AES_ENC/u0/u2/n806 , \AES_ENC/u0/u2/n805 ,\AES_ENC/u0/u2/n804 , \AES_ENC/u0/u2/n803 , \AES_ENC/u0/u2/n802 ,\AES_ENC/u0/u2/n801 , \AES_ENC/u0/u2/n800 , \AES_ENC/u0/u2/n799 ,\AES_ENC/u0/u2/n798 , \AES_ENC/u0/u2/n797 , \AES_ENC/u0/u2/n796 ,\AES_ENC/u0/u2/n795 , \AES_ENC/u0/u2/n794 , \AES_ENC/u0/u2/n793 ,\AES_ENC/u0/u2/n792 , \AES_ENC/u0/u2/n791 , \AES_ENC/u0/u2/n790 ,\AES_ENC/u0/u2/n789 , \AES_ENC/u0/u2/n788 , \AES_ENC/u0/u2/n787 ,\AES_ENC/u0/u2/n786 , \AES_ENC/u0/u2/n785 , \AES_ENC/u0/u2/n784 ,\AES_ENC/u0/u2/n783 , \AES_ENC/u0/u2/n782 , \AES_ENC/u0/u2/n781 ,\AES_ENC/u0/u2/n780 , \AES_ENC/u0/u2/n779 , \AES_ENC/u0/u2/n778 ,\AES_ENC/u0/u2/n777 , \AES_ENC/u0/u2/n776 , \AES_ENC/u0/u2/n775 ,\AES_ENC/u0/u2/n774 , \AES_ENC/u0/u2/n773 , \AES_ENC/u0/u2/n772 ,\AES_ENC/u0/u2/n771 , \AES_ENC/u0/u2/n770 , \AES_ENC/u0/u2/n769 ,\AES_ENC/u0/u2/n768 , \AES_ENC/u0/u2/n767 , \AES_ENC/u0/u2/n766 ,\AES_ENC/u0/u2/n765 , \AES_ENC/u0/u2/n764 , \AES_ENC/u0/u2/n763 ,\AES_ENC/u0/u2/n762 , \AES_ENC/u0/u2/n761 , \AES_ENC/u0/u2/n760 ,\AES_ENC/u0/u2/n759 , \AES_ENC/u0/u2/n758 , \AES_ENC/u0/u2/n757 ,\AES_ENC/u0/u2/n756 , \AES_ENC/u0/u2/n755 , \AES_ENC/u0/u2/n754 ,\AES_ENC/u0/u2/n753 , \AES_ENC/u0/u2/n752 , \AES_ENC/u0/u2/n751 ,\AES_ENC/u0/u2/n750 , \AES_ENC/u0/u2/n749 , \AES_ENC/u0/u2/n748 ,\AES_ENC/u0/u2/n747 , \AES_ENC/u0/u2/n746 , \AES_ENC/u0/u2/n745 ,\AES_ENC/u0/u2/n744 , \AES_ENC/u0/u2/n743 , \AES_ENC/u0/u2/n742 ,\AES_ENC/u0/u2/n741 , \AES_ENC/u0/u2/n740 , \AES_ENC/u0/u2/n739 ,\AES_ENC/u0/u2/n738 , \AES_ENC/u0/u2/n737 , \AES_ENC/u0/u2/n736 ,\AES_ENC/u0/u2/n735 , \AES_ENC/u0/u2/n734 , \AES_ENC/u0/u2/n733 ,\AES_ENC/u0/u2/n732 , \AES_ENC/u0/u2/n731 , \AES_ENC/u0/u2/n730 ,\AES_ENC/u0/u2/n729 , \AES_ENC/u0/u2/n728 , \AES_ENC/u0/u2/n727 ,\AES_ENC/u0/u2/n726 , \AES_ENC/u0/u2/n725 , \AES_ENC/u0/u2/n724 ,\AES_ENC/u0/u2/n723 , \AES_ENC/u0/u2/n722 , \AES_ENC/u0/u2/n721 ,\AES_ENC/u0/u2/n720 , \AES_ENC/u0/u2/n719 , \AES_ENC/u0/u2/n718 ,\AES_ENC/u0/u2/n717 , \AES_ENC/u0/u2/n716 , \AES_ENC/u0/u2/n715 ,\AES_ENC/u0/u2/n714 , \AES_ENC/u0/u2/n713 , \AES_ENC/u0/u2/n712 ,\AES_ENC/u0/u2/n711 , \AES_ENC/u0/u2/n710 , \AES_ENC/u0/u2/n709 ,\AES_ENC/u0/u2/n708 , \AES_ENC/u0/u2/n707 , \AES_ENC/u0/u2/n706 ,\AES_ENC/u0/u2/n705 , \AES_ENC/u0/u2/n704 , \AES_ENC/u0/u2/n703 ,\AES_ENC/u0/u2/n702 , \AES_ENC/u0/u2/n701 , \AES_ENC/u0/u2/n700 ,\AES_ENC/u0/u2/n699 , \AES_ENC/u0/u2/n698 , \AES_ENC/u0/u2/n697 ,\AES_ENC/u0/u2/n696 , \AES_ENC/u0/u2/n695 , \AES_ENC/u0/u2/n694 ,\AES_ENC/u0/u2/n693 , \AES_ENC/u0/u2/n692 , \AES_ENC/u0/u2/n691 ,\AES_ENC/u0/u2/n690 , \AES_ENC/u0/u2/n689 , \AES_ENC/u0/u2/n688 ,\AES_ENC/u0/u2/n687 , \AES_ENC/u0/u2/n686 , \AES_ENC/u0/u2/n685 ,\AES_ENC/u0/u2/n684 , \AES_ENC/u0/u2/n683 , \AES_ENC/u0/u2/n682 ,\AES_ENC/u0/u2/n681 , \AES_ENC/u0/u2/n680 , \AES_ENC/u0/u2/n679 ,\AES_ENC/u0/u2/n678 , \AES_ENC/u0/u2/n677 , \AES_ENC/u0/u2/n676 ,\AES_ENC/u0/u2/n675 , \AES_ENC/u0/u2/n674 , \AES_ENC/u0/u2/n673 ,\AES_ENC/u0/u2/n672 , \AES_ENC/u0/u2/n671 , \AES_ENC/u0/u2/n670 ,\AES_ENC/u0/u2/n669 , \AES_ENC/u0/u2/n668 , \AES_ENC/u0/u2/n667 ,\AES_ENC/u0/u2/n666 , \AES_ENC/u0/u2/n665 , \AES_ENC/u0/u2/n664 ,\AES_ENC/u0/u2/n663 , \AES_ENC/u0/u2/n662 , \AES_ENC/u0/u2/n661 ,\AES_ENC/u0/u2/n660 , \AES_ENC/u0/u2/n659 , \AES_ENC/u0/u2/n658 ,\AES_ENC/u0/u2/n657 , \AES_ENC/u0/u2/n656 , \AES_ENC/u0/u2/n655 ,\AES_ENC/u0/u2/n654 , \AES_ENC/u0/u2/n653 , \AES_ENC/u0/u2/n652 ,\AES_ENC/u0/u2/n651 , \AES_ENC/u0/u2/n650 , \AES_ENC/u0/u2/n649 ,\AES_ENC/u0/u2/n648 , \AES_ENC/u0/u2/n647 , \AES_ENC/u0/u2/n646 ,\AES_ENC/u0/u2/n645 , \AES_ENC/u0/u2/n644 , \AES_ENC/u0/u2/n643 ,\AES_ENC/u0/u2/n642 , \AES_ENC/u0/u2/n641 , \AES_ENC/u0/u2/n640 ,\AES_ENC/u0/u2/n639 , \AES_ENC/u0/u2/n638 , \AES_ENC/u0/u2/n637 ,\AES_ENC/u0/u2/n636 , \AES_ENC/u0/u2/n635 , \AES_ENC/u0/u2/n634 ,\AES_ENC/u0/u2/n633 , \AES_ENC/u0/u2/n632 , \AES_ENC/u0/u2/n631 ,\AES_ENC/u0/u2/n630 , \AES_ENC/u0/u2/n629 , \AES_ENC/u0/u2/n628 ,\AES_ENC/u0/u2/n627 , \AES_ENC/u0/u2/n626 , \AES_ENC/u0/u2/n625 ,\AES_ENC/u0/u2/n624 , \AES_ENC/u0/u2/n623 , \AES_ENC/u0/u2/n622 ,\AES_ENC/u0/u2/n621 , \AES_ENC/u0/u2/n620 , \AES_ENC/u0/u2/n619 ,\AES_ENC/u0/u2/n618 , \AES_ENC/u0/u2/n617 , \AES_ENC/u0/u2/n616 ,\AES_ENC/u0/u2/n615 , \AES_ENC/u0/u2/n614 , \AES_ENC/u0/u2/n613 ,\AES_ENC/u0/u2/n612 , \AES_ENC/u0/u2/n611 , \AES_ENC/u0/u2/n610 ,\AES_ENC/u0/u2/n609 , \AES_ENC/u0/u2/n608 , \AES_ENC/u0/u2/n607 ,\AES_ENC/u0/u2/n606 , \AES_ENC/u0/u2/n605 , \AES_ENC/u0/u2/n604 ,\AES_ENC/u0/u2/n603 , \AES_ENC/u0/u2/n602 , \AES_ENC/u0/u2/n601 ,\AES_ENC/u0/u2/n600 , \AES_ENC/u0/u2/n599 , \AES_ENC/u0/u2/n598 ,\AES_ENC/u0/u2/n597 , \AES_ENC/u0/u2/n596 , \AES_ENC/u0/u2/n595 ,\AES_ENC/u0/u2/n594 , \AES_ENC/u0/u2/n593 , \AES_ENC/u0/u2/n592 ,\AES_ENC/u0/u2/n591 , \AES_ENC/u0/u2/n590 , \AES_ENC/u0/u2/n589 ,\AES_ENC/u0/u2/n588 , \AES_ENC/u0/u2/n587 , \AES_ENC/u0/u2/n586 ,\AES_ENC/u0/u2/n585 , \AES_ENC/u0/u2/n584 , \AES_ENC/u0/u2/n583 ,\AES_ENC/u0/u2/n582 , \AES_ENC/u0/u2/n581 , \AES_ENC/u0/u2/n580 ,\AES_ENC/u0/u2/n579 , \AES_ENC/u0/u2/n578 , \AES_ENC/u0/u2/n577 ,\AES_ENC/u0/u2/n576 , \AES_ENC/u0/u2/n575 , \AES_ENC/u0/u2/n574 ,\AES_ENC/u0/u2/n573 , \AES_ENC/u0/u2/n572 , \AES_ENC/u0/u2/n571 ,\AES_ENC/u0/u2/n570 , \AES_ENC/u0/u2/n569 , \AES_ENC/u0/u3/n1135 ,\AES_ENC/u0/u3/n1134 , \AES_ENC/u0/u3/n1133 , \AES_ENC/u0/u3/n1132 ,\AES_ENC/u0/u3/n1131 , \AES_ENC/u0/u3/n1130 , \AES_ENC/u0/u3/n1129 ,\AES_ENC/u0/u3/n1128 , \AES_ENC/u0/u3/n1127 , \AES_ENC/u0/u3/n1126 ,\AES_ENC/u0/u3/n1125 , \AES_ENC/u0/u3/n1124 , \AES_ENC/u0/u3/n1123 ,\AES_ENC/u0/u3/n1122 , \AES_ENC/u0/u3/n1121 , \AES_ENC/u0/u3/n1120 ,\AES_ENC/u0/u3/n1119 , \AES_ENC/u0/u3/n1118 , \AES_ENC/u0/u3/n1117 ,\AES_ENC/u0/u3/n1116 , \AES_ENC/u0/u3/n1115 , \AES_ENC/u0/u3/n1114 ,\AES_ENC/u0/u3/n1113 , \AES_ENC/u0/u3/n1112 , \AES_ENC/u0/u3/n1111 ,\AES_ENC/u0/u3/n1110 , \AES_ENC/u0/u3/n1109 , \AES_ENC/u0/u3/n1108 ,\AES_ENC/u0/u3/n1107 , \AES_ENC/u0/u3/n1106 , \AES_ENC/u0/u3/n1105 ,\AES_ENC/u0/u3/n1104 , \AES_ENC/u0/u3/n1103 , \AES_ENC/u0/u3/n1102 ,\AES_ENC/u0/u3/n1101 , \AES_ENC/u0/u3/n1100 , \AES_ENC/u0/u3/n1099 ,\AES_ENC/u0/u3/n1098 , \AES_ENC/u0/u3/n1097 , \AES_ENC/u0/u3/n1096 ,\AES_ENC/u0/u3/n1095 , \AES_ENC/u0/u3/n1094 , \AES_ENC/u0/u3/n1093 ,\AES_ENC/u0/u3/n1092 , \AES_ENC/u0/u3/n1091 , \AES_ENC/u0/u3/n1090 ,\AES_ENC/u0/u3/n1089 , \AES_ENC/u0/u3/n1088 , \AES_ENC/u0/u3/n1087 ,\AES_ENC/u0/u3/n1086 , \AES_ENC/u0/u3/n1085 , \AES_ENC/u0/u3/n1084 ,\AES_ENC/u0/u3/n1083 , \AES_ENC/u0/u3/n1082 , \AES_ENC/u0/u3/n1081 ,\AES_ENC/u0/u3/n1080 , \AES_ENC/u0/u3/n1079 , \AES_ENC/u0/u3/n1078 ,\AES_ENC/u0/u3/n1077 , \AES_ENC/u0/u3/n1076 , \AES_ENC/u0/u3/n1075 ,\AES_ENC/u0/u3/n1074 , \AES_ENC/u0/u3/n1073 , \AES_ENC/u0/u3/n1072 ,\AES_ENC/u0/u3/n1071 , \AES_ENC/u0/u3/n1070 , \AES_ENC/u0/u3/n1069 ,\AES_ENC/u0/u3/n1068 , \AES_ENC/u0/u3/n1067 , \AES_ENC/u0/u3/n1066 ,\AES_ENC/u0/u3/n1065 , \AES_ENC/u0/u3/n1064 , \AES_ENC/u0/u3/n1063 ,\AES_ENC/u0/u3/n1062 , \AES_ENC/u0/u3/n1061 , \AES_ENC/u0/u3/n1060 ,\AES_ENC/u0/u3/n1059 , \AES_ENC/u0/u3/n1058 , \AES_ENC/u0/u3/n1057 ,\AES_ENC/u0/u3/n1056 , \AES_ENC/u0/u3/n1055 , \AES_ENC/u0/u3/n1054 ,\AES_ENC/u0/u3/n1053 , \AES_ENC/u0/u3/n1052 , \AES_ENC/u0/u3/n1051 ,\AES_ENC/u0/u3/n1050 , \AES_ENC/u0/u3/n1049 , \AES_ENC/u0/u3/n1048 ,\AES_ENC/u0/u3/n1047 , \AES_ENC/u0/u3/n1046 , \AES_ENC/u0/u3/n1045 ,\AES_ENC/u0/u3/n1044 , \AES_ENC/u0/u3/n1043 , \AES_ENC/u0/u3/n1042 ,\AES_ENC/u0/u3/n1041 , \AES_ENC/u0/u3/n1040 , \AES_ENC/u0/u3/n1039 ,\AES_ENC/u0/u3/n1038 , \AES_ENC/u0/u3/n1037 , \AES_ENC/u0/u3/n1036 ,\AES_ENC/u0/u3/n1035 , \AES_ENC/u0/u3/n1034 , \AES_ENC/u0/u3/n1033 ,\AES_ENC/u0/u3/n1032 , \AES_ENC/u0/u3/n1031 , \AES_ENC/u0/u3/n1030 ,\AES_ENC/u0/u3/n1029 , \AES_ENC/u0/u3/n1028 , \AES_ENC/u0/u3/n1027 ,\AES_ENC/u0/u3/n1026 , \AES_ENC/u0/u3/n1025 , \AES_ENC/u0/u3/n1024 ,\AES_ENC/u0/u3/n1023 , \AES_ENC/u0/u3/n1022 , \AES_ENC/u0/u3/n1021 ,\AES_ENC/u0/u3/n1020 , \AES_ENC/u0/u3/n1019 , \AES_ENC/u0/u3/n1018 ,\AES_ENC/u0/u3/n1017 , \AES_ENC/u0/u3/n1016 , \AES_ENC/u0/u3/n1015 ,\AES_ENC/u0/u3/n1014 , \AES_ENC/u0/u3/n1013 , \AES_ENC/u0/u3/n1012 ,\AES_ENC/u0/u3/n1011 , \AES_ENC/u0/u3/n1010 , \AES_ENC/u0/u3/n1009 ,\AES_ENC/u0/u3/n1008 , \AES_ENC/u0/u3/n1007 , \AES_ENC/u0/u3/n1006 ,\AES_ENC/u0/u3/n1005 , \AES_ENC/u0/u3/n1004 , \AES_ENC/u0/u3/n1003 ,\AES_ENC/u0/u3/n1002 , \AES_ENC/u0/u3/n1001 , \AES_ENC/u0/u3/n1000 ,\AES_ENC/u0/u3/n999 , \AES_ENC/u0/u3/n998 , \AES_ENC/u0/u3/n997 ,\AES_ENC/u0/u3/n996 , \AES_ENC/u0/u3/n995 , \AES_ENC/u0/u3/n994 ,\AES_ENC/u0/u3/n993 , \AES_ENC/u0/u3/n992 , \AES_ENC/u0/u3/n991 ,\AES_ENC/u0/u3/n990 , \AES_ENC/u0/u3/n989 , \AES_ENC/u0/u3/n988 ,\AES_ENC/u0/u3/n987 , \AES_ENC/u0/u3/n986 , \AES_ENC/u0/u3/n985 ,\AES_ENC/u0/u3/n984 , \AES_ENC/u0/u3/n983 , \AES_ENC/u0/u3/n982 ,\AES_ENC/u0/u3/n981 , \AES_ENC/u0/u3/n980 , \AES_ENC/u0/u3/n979 ,\AES_ENC/u0/u3/n978 , \AES_ENC/u0/u3/n977 , \AES_ENC/u0/u3/n976 ,\AES_ENC/u0/u3/n975 , \AES_ENC/u0/u3/n974 , \AES_ENC/u0/u3/n973 ,\AES_ENC/u0/u3/n972 , \AES_ENC/u0/u3/n971 , \AES_ENC/u0/u3/n970 ,\AES_ENC/u0/u3/n969 , \AES_ENC/u0/u3/n968 , \AES_ENC/u0/u3/n967 ,\AES_ENC/u0/u3/n966 , \AES_ENC/u0/u3/n965 , \AES_ENC/u0/u3/n964 ,\AES_ENC/u0/u3/n963 , \AES_ENC/u0/u3/n962 , \AES_ENC/u0/u3/n961 ,\AES_ENC/u0/u3/n960 , \AES_ENC/u0/u3/n959 , \AES_ENC/u0/u3/n958 ,\AES_ENC/u0/u3/n957 , \AES_ENC/u0/u3/n956 , \AES_ENC/u0/u3/n955 ,\AES_ENC/u0/u3/n954 , \AES_ENC/u0/u3/n953 , \AES_ENC/u0/u3/n952 ,\AES_ENC/u0/u3/n951 , \AES_ENC/u0/u3/n950 , \AES_ENC/u0/u3/n949 ,\AES_ENC/u0/u3/n948 , \AES_ENC/u0/u3/n947 , \AES_ENC/u0/u3/n946 ,\AES_ENC/u0/u3/n945 , \AES_ENC/u0/u3/n944 , \AES_ENC/u0/u3/n943 ,\AES_ENC/u0/u3/n942 , \AES_ENC/u0/u3/n941 , \AES_ENC/u0/u3/n940 ,\AES_ENC/u0/u3/n939 , \AES_ENC/u0/u3/n938 , \AES_ENC/u0/u3/n937 ,\AES_ENC/u0/u3/n936 , \AES_ENC/u0/u3/n935 , \AES_ENC/u0/u3/n934 ,\AES_ENC/u0/u3/n933 , \AES_ENC/u0/u3/n932 , \AES_ENC/u0/u3/n931 ,\AES_ENC/u0/u3/n930 , \AES_ENC/u0/u3/n929 , \AES_ENC/u0/u3/n928 ,\AES_ENC/u0/u3/n927 , \AES_ENC/u0/u3/n926 , \AES_ENC/u0/u3/n925 ,\AES_ENC/u0/u3/n924 , \AES_ENC/u0/u3/n923 , \AES_ENC/u0/u3/n922 ,\AES_ENC/u0/u3/n921 , \AES_ENC/u0/u3/n920 , \AES_ENC/u0/u3/n919 ,\AES_ENC/u0/u3/n918 , \AES_ENC/u0/u3/n917 , \AES_ENC/u0/u3/n916 ,\AES_ENC/u0/u3/n915 , \AES_ENC/u0/u3/n914 , \AES_ENC/u0/u3/n913 ,\AES_ENC/u0/u3/n912 , \AES_ENC/u0/u3/n911 , \AES_ENC/u0/u3/n910 ,\AES_ENC/u0/u3/n909 , \AES_ENC/u0/u3/n908 , \AES_ENC/u0/u3/n907 ,\AES_ENC/u0/u3/n906 , \AES_ENC/u0/u3/n905 , \AES_ENC/u0/u3/n904 ,\AES_ENC/u0/u3/n903 , \AES_ENC/u0/u3/n902 , \AES_ENC/u0/u3/n901 ,\AES_ENC/u0/u3/n900 , \AES_ENC/u0/u3/n899 , \AES_ENC/u0/u3/n898 ,\AES_ENC/u0/u3/n897 , \AES_ENC/u0/u3/n896 , \AES_ENC/u0/u3/n895 ,\AES_ENC/u0/u3/n894 , \AES_ENC/u0/u3/n893 , \AES_ENC/u0/u3/n892 ,\AES_ENC/u0/u3/n891 , \AES_ENC/u0/u3/n890 , \AES_ENC/u0/u3/n889 ,\AES_ENC/u0/u3/n888 , \AES_ENC/u0/u3/n887 , \AES_ENC/u0/u3/n886 ,\AES_ENC/u0/u3/n885 , \AES_ENC/u0/u3/n884 , \AES_ENC/u0/u3/n883 ,\AES_ENC/u0/u3/n882 , \AES_ENC/u0/u3/n881 , \AES_ENC/u0/u3/n880 ,\AES_ENC/u0/u3/n879 , \AES_ENC/u0/u3/n878 , \AES_ENC/u0/u3/n877 ,\AES_ENC/u0/u3/n876 , \AES_ENC/u0/u3/n875 , \AES_ENC/u0/u3/n874 ,\AES_ENC/u0/u3/n873 , \AES_ENC/u0/u3/n872 , \AES_ENC/u0/u3/n871 ,\AES_ENC/u0/u3/n870 , \AES_ENC/u0/u3/n869 , \AES_ENC/u0/u3/n868 ,\AES_ENC/u0/u3/n867 , \AES_ENC/u0/u3/n866 , \AES_ENC/u0/u3/n865 ,\AES_ENC/u0/u3/n864 , \AES_ENC/u0/u3/n863 , \AES_ENC/u0/u3/n862 ,\AES_ENC/u0/u3/n861 , \AES_ENC/u0/u3/n860 , \AES_ENC/u0/u3/n859 ,\AES_ENC/u0/u3/n858 , \AES_ENC/u0/u3/n857 , \AES_ENC/u0/u3/n856 ,\AES_ENC/u0/u3/n855 , \AES_ENC/u0/u3/n854 , \AES_ENC/u0/u3/n853 ,\AES_ENC/u0/u3/n852 , \AES_ENC/u0/u3/n851 , \AES_ENC/u0/u3/n850 ,\AES_ENC/u0/u3/n849 , \AES_ENC/u0/u3/n848 , \AES_ENC/u0/u3/n847 ,\AES_ENC/u0/u3/n846 , \AES_ENC/u0/u3/n845 , \AES_ENC/u0/u3/n844 ,\AES_ENC/u0/u3/n843 , \AES_ENC/u0/u3/n842 , \AES_ENC/u0/u3/n841 ,\AES_ENC/u0/u3/n840 , \AES_ENC/u0/u3/n839 , \AES_ENC/u0/u3/n838 ,\AES_ENC/u0/u3/n837 , \AES_ENC/u0/u3/n836 , \AES_ENC/u0/u3/n835 ,\AES_ENC/u0/u3/n834 , \AES_ENC/u0/u3/n833 , \AES_ENC/u0/u3/n832 ,\AES_ENC/u0/u3/n831 , \AES_ENC/u0/u3/n830 , \AES_ENC/u0/u3/n829 ,\AES_ENC/u0/u3/n828 , \AES_ENC/u0/u3/n827 , \AES_ENC/u0/u3/n826 ,\AES_ENC/u0/u3/n825 , \AES_ENC/u0/u3/n824 , \AES_ENC/u0/u3/n823 ,\AES_ENC/u0/u3/n822 , \AES_ENC/u0/u3/n821 , \AES_ENC/u0/u3/n820 ,\AES_ENC/u0/u3/n819 , \AES_ENC/u0/u3/n818 , \AES_ENC/u0/u3/n817 ,\AES_ENC/u0/u3/n816 , \AES_ENC/u0/u3/n815 , \AES_ENC/u0/u3/n814 ,\AES_ENC/u0/u3/n813 , \AES_ENC/u0/u3/n812 , \AES_ENC/u0/u3/n811 ,\AES_ENC/u0/u3/n810 , \AES_ENC/u0/u3/n809 , \AES_ENC/u0/u3/n808 ,\AES_ENC/u0/u3/n807 , \AES_ENC/u0/u3/n806 , \AES_ENC/u0/u3/n805 ,\AES_ENC/u0/u3/n804 , \AES_ENC/u0/u3/n803 , \AES_ENC/u0/u3/n802 ,\AES_ENC/u0/u3/n801 , \AES_ENC/u0/u3/n800 , \AES_ENC/u0/u3/n799 ,\AES_ENC/u0/u3/n798 , \AES_ENC/u0/u3/n797 , \AES_ENC/u0/u3/n796 ,\AES_ENC/u0/u3/n795 , \AES_ENC/u0/u3/n794 , \AES_ENC/u0/u3/n793 ,\AES_ENC/u0/u3/n792 , \AES_ENC/u0/u3/n791 , \AES_ENC/u0/u3/n790 ,\AES_ENC/u0/u3/n789 , \AES_ENC/u0/u3/n788 , \AES_ENC/u0/u3/n787 ,\AES_ENC/u0/u3/n786 , \AES_ENC/u0/u3/n785 , \AES_ENC/u0/u3/n784 ,\AES_ENC/u0/u3/n783 , \AES_ENC/u0/u3/n782 , \AES_ENC/u0/u3/n781 ,\AES_ENC/u0/u3/n780 , \AES_ENC/u0/u3/n779 , \AES_ENC/u0/u3/n778 ,\AES_ENC/u0/u3/n777 , \AES_ENC/u0/u3/n776 , \AES_ENC/u0/u3/n775 ,\AES_ENC/u0/u3/n774 , \AES_ENC/u0/u3/n773 , \AES_ENC/u0/u3/n772 ,\AES_ENC/u0/u3/n771 , \AES_ENC/u0/u3/n770 , \AES_ENC/u0/u3/n769 ,\AES_ENC/u0/u3/n768 , \AES_ENC/u0/u3/n767 , \AES_ENC/u0/u3/n766 ,\AES_ENC/u0/u3/n765 , \AES_ENC/u0/u3/n764 , \AES_ENC/u0/u3/n763 ,\AES_ENC/u0/u3/n762 , \AES_ENC/u0/u3/n761 , \AES_ENC/u0/u3/n760 ,\AES_ENC/u0/u3/n759 , \AES_ENC/u0/u3/n758 , \AES_ENC/u0/u3/n757 ,\AES_ENC/u0/u3/n756 , \AES_ENC/u0/u3/n755 , \AES_ENC/u0/u3/n754 ,\AES_ENC/u0/u3/n753 , \AES_ENC/u0/u3/n752 , \AES_ENC/u0/u3/n751 ,\AES_ENC/u0/u3/n750 , \AES_ENC/u0/u3/n749 , \AES_ENC/u0/u3/n748 ,\AES_ENC/u0/u3/n747 , \AES_ENC/u0/u3/n746 , \AES_ENC/u0/u3/n745 ,\AES_ENC/u0/u3/n744 , \AES_ENC/u0/u3/n743 , \AES_ENC/u0/u3/n742 ,\AES_ENC/u0/u3/n741 , \AES_ENC/u0/u3/n740 , \AES_ENC/u0/u3/n739 ,\AES_ENC/u0/u3/n738 , \AES_ENC/u0/u3/n737 , \AES_ENC/u0/u3/n736 ,\AES_ENC/u0/u3/n735 , \AES_ENC/u0/u3/n734 , \AES_ENC/u0/u3/n733 ,\AES_ENC/u0/u3/n732 , \AES_ENC/u0/u3/n731 , \AES_ENC/u0/u3/n730 ,\AES_ENC/u0/u3/n729 , \AES_ENC/u0/u3/n728 , \AES_ENC/u0/u3/n727 ,\AES_ENC/u0/u3/n726 , \AES_ENC/u0/u3/n725 , \AES_ENC/u0/u3/n724 ,\AES_ENC/u0/u3/n723 , \AES_ENC/u0/u3/n722 , \AES_ENC/u0/u3/n721 ,\AES_ENC/u0/u3/n720 , \AES_ENC/u0/u3/n719 , \AES_ENC/u0/u3/n718 ,\AES_ENC/u0/u3/n717 , \AES_ENC/u0/u3/n716 , \AES_ENC/u0/u3/n715 ,\AES_ENC/u0/u3/n714 , \AES_ENC/u0/u3/n713 , \AES_ENC/u0/u3/n712 ,\AES_ENC/u0/u3/n711 , \AES_ENC/u0/u3/n710 , \AES_ENC/u0/u3/n709 ,\AES_ENC/u0/u3/n708 , \AES_ENC/u0/u3/n707 , \AES_ENC/u0/u3/n706 ,\AES_ENC/u0/u3/n705 , \AES_ENC/u0/u3/n704 , \AES_ENC/u0/u3/n703 ,\AES_ENC/u0/u3/n702 , \AES_ENC/u0/u3/n701 , \AES_ENC/u0/u3/n700 ,\AES_ENC/u0/u3/n699 , \AES_ENC/u0/u3/n698 , \AES_ENC/u0/u3/n697 ,\AES_ENC/u0/u3/n696 , \AES_ENC/u0/u3/n695 , \AES_ENC/u0/u3/n694 ,\AES_ENC/u0/u3/n693 , \AES_ENC/u0/u3/n692 , \AES_ENC/u0/u3/n691 ,\AES_ENC/u0/u3/n690 , \AES_ENC/u0/u3/n689 , \AES_ENC/u0/u3/n688 ,\AES_ENC/u0/u3/n687 , \AES_ENC/u0/u3/n686 , \AES_ENC/u0/u3/n685 ,\AES_ENC/u0/u3/n684 , \AES_ENC/u0/u3/n683 , \AES_ENC/u0/u3/n682 ,\AES_ENC/u0/u3/n681 , \AES_ENC/u0/u3/n680 , \AES_ENC/u0/u3/n679 ,\AES_ENC/u0/u3/n678 , \AES_ENC/u0/u3/n677 , \AES_ENC/u0/u3/n676 ,\AES_ENC/u0/u3/n675 , \AES_ENC/u0/u3/n674 , \AES_ENC/u0/u3/n673 ,\AES_ENC/u0/u3/n672 , \AES_ENC/u0/u3/n671 , \AES_ENC/u0/u3/n670 ,\AES_ENC/u0/u3/n669 , \AES_ENC/u0/u3/n668 , \AES_ENC/u0/u3/n667 ,\AES_ENC/u0/u3/n666 , \AES_ENC/u0/u3/n665 , \AES_ENC/u0/u3/n664 ,\AES_ENC/u0/u3/n663 , \AES_ENC/u0/u3/n662 , \AES_ENC/u0/u3/n661 ,\AES_ENC/u0/u3/n660 , \AES_ENC/u0/u3/n659 , \AES_ENC/u0/u3/n658 ,\AES_ENC/u0/u3/n657 , \AES_ENC/u0/u3/n656 , \AES_ENC/u0/u3/n655 ,\AES_ENC/u0/u3/n654 , \AES_ENC/u0/u3/n653 , \AES_ENC/u0/u3/n652 ,\AES_ENC/u0/u3/n651 , \AES_ENC/u0/u3/n650 , \AES_ENC/u0/u3/n649 ,\AES_ENC/u0/u3/n648 , \AES_ENC/u0/u3/n647 , \AES_ENC/u0/u3/n646 ,\AES_ENC/u0/u3/n645 , \AES_ENC/u0/u3/n644 , \AES_ENC/u0/u3/n643 ,\AES_ENC/u0/u3/n642 , \AES_ENC/u0/u3/n641 , \AES_ENC/u0/u3/n640 ,\AES_ENC/u0/u3/n639 , \AES_ENC/u0/u3/n638 , \AES_ENC/u0/u3/n637 ,\AES_ENC/u0/u3/n636 , \AES_ENC/u0/u3/n635 , \AES_ENC/u0/u3/n634 ,\AES_ENC/u0/u3/n633 , \AES_ENC/u0/u3/n632 , \AES_ENC/u0/u3/n631 ,\AES_ENC/u0/u3/n630 , \AES_ENC/u0/u3/n629 , \AES_ENC/u0/u3/n628 ,\AES_ENC/u0/u3/n627 , \AES_ENC/u0/u3/n626 , \AES_ENC/u0/u3/n625 ,\AES_ENC/u0/u3/n624 , \AES_ENC/u0/u3/n623 , \AES_ENC/u0/u3/n622 ,\AES_ENC/u0/u3/n621 , \AES_ENC/u0/u3/n620 , \AES_ENC/u0/u3/n619 ,\AES_ENC/u0/u3/n618 , \AES_ENC/u0/u3/n617 , \AES_ENC/u0/u3/n616 ,\AES_ENC/u0/u3/n615 , \AES_ENC/u0/u3/n614 , \AES_ENC/u0/u3/n613 ,\AES_ENC/u0/u3/n612 , \AES_ENC/u0/u3/n611 , \AES_ENC/u0/u3/n610 ,\AES_ENC/u0/u3/n609 , \AES_ENC/u0/u3/n608 , \AES_ENC/u0/u3/n607 ,\AES_ENC/u0/u3/n606 , \AES_ENC/u0/u3/n605 , \AES_ENC/u0/u3/n604 ,\AES_ENC/u0/u3/n603 , \AES_ENC/u0/u3/n602 , \AES_ENC/u0/u3/n601 ,\AES_ENC/u0/u3/n600 , \AES_ENC/u0/u3/n599 , \AES_ENC/u0/u3/n598 ,\AES_ENC/u0/u3/n597 , \AES_ENC/u0/u3/n596 , \AES_ENC/u0/u3/n595 ,\AES_ENC/u0/u3/n594 , \AES_ENC/u0/u3/n593 , \AES_ENC/u0/u3/n592 ,\AES_ENC/u0/u3/n591 , \AES_ENC/u0/u3/n590 , \AES_ENC/u0/u3/n589 ,\AES_ENC/u0/u3/n588 , \AES_ENC/u0/u3/n587 , \AES_ENC/u0/u3/n586 ,\AES_ENC/u0/u3/n585 , \AES_ENC/u0/u3/n584 , \AES_ENC/u0/u3/n583 ,\AES_ENC/u0/u3/n582 , \AES_ENC/u0/u3/n581 , \AES_ENC/u0/u3/n580 ,\AES_ENC/u0/u3/n579 , \AES_ENC/u0/u3/n578 , \AES_ENC/u0/u3/n577 ,\AES_ENC/u0/u3/n576 , \AES_ENC/u0/u3/n575 , \AES_ENC/u0/u3/n574 ,\AES_ENC/u0/u3/n573 , \AES_ENC/u0/u3/n572 , \AES_ENC/u0/u3/n571 ,\AES_ENC/u0/u3/n570 , \AES_ENC/u0/u3/n569 , \AES_ENC/u0/r0/n38 ,\AES_ENC/u0/r0/n37 , \AES_ENC/u0/r0/n36 , \AES_ENC/u0/r0/n35 ,\AES_ENC/u0/r0/n34 , \AES_ENC/u0/r0/n33 , \AES_ENC/u0/r0/n29 ,\AES_ENC/u0/r0/n28 , \AES_ENC/u0/r0/n27 , \AES_ENC/u0/r0/n26 ,\AES_ENC/u0/r0/n25 , \AES_ENC/u0/r0/n24 , \AES_ENC/u0/r0/n23 ,\AES_ENC/u0/r0/n22 , \AES_ENC/u0/r0/n21 , \AES_ENC/u0/r0/n20 ,\AES_ENC/u0/r0/n19 , \AES_ENC/u0/r0/n18 , \AES_ENC/u0/r0/n17 ,\AES_ENC/u0/r0/n16 , \AES_ENC/u0/r0/n15 , \AES_ENC/u0/r0/n14 ,\AES_ENC/u0/r0/n13 , \AES_ENC/u0/r0/n12 , \AES_ENC/u0/r0/n11 ,\AES_ENC/u0/r0/n10 , \AES_ENC/u0/r0/n9 , \AES_ENC/u0/r0/n8 ,\AES_ENC/u0/r0/n7 , \AES_ENC/u0/r0/n32 , \AES_ENC/u0/r0/N55 ,\AES_ENC/u0/r0/N54 , \AES_ENC/u0/r0/N53 , \AES_ENC/u0/r0/rcnt[0] ,\AES_ENC/u0/r0/rcnt[1] , \AES_ENC/u0/r0/rcnt[2] , \AES_ENC/u0/r0/N51 ,\AES_ENC/u0/r0/N50 , \AES_ENC/u0/r0/N49 , \AES_ENC/u0/r0/N48 ,\AES_ENC/u0/r0/N47 , \AES_ENC/u0/r0/N46 , \AES_ENC/u0/r0/N45 ,\AES_ENC/u0/r0/N44 , \AES_ENC/us00/n627 , \AES_ENC/us00/n626 ,\AES_ENC/us00/n625 , \AES_ENC/us00/n624 , \AES_ENC/us00/n623 ,\AES_ENC/us00/n622 , \AES_ENC/us00/n621 , \AES_ENC/us00/n620 ,\AES_ENC/us00/n619 , \AES_ENC/us00/n618 , \AES_ENC/us00/n617 ,\AES_ENC/us00/n616 , \AES_ENC/us00/n615 , \AES_ENC/us00/n614 ,\AES_ENC/us00/n613 , \AES_ENC/us00/n612 , \AES_ENC/us00/n611 ,\AES_ENC/us00/n610 , \AES_ENC/us00/n609 , \AES_ENC/us00/n608 ,\AES_ENC/us00/n607 , \AES_ENC/us00/n606 , \AES_ENC/us00/n605 ,\AES_ENC/us00/n604 , \AES_ENC/us00/n603 , \AES_ENC/us00/n602 ,\AES_ENC/us00/n601 , \AES_ENC/us00/n600 , \AES_ENC/us00/n599 ,\AES_ENC/us00/n598 , \AES_ENC/us00/n597 , \AES_ENC/us00/n596 ,\AES_ENC/us00/n595 , \AES_ENC/us00/n594 , \AES_ENC/us00/n593 ,\AES_ENC/us00/n592 , \AES_ENC/us00/n591 , \AES_ENC/us00/n590 ,\AES_ENC/us00/n589 , \AES_ENC/us00/n588 , \AES_ENC/us00/n587 ,\AES_ENC/us00/n586 , \AES_ENC/us00/n585 , \AES_ENC/us00/n584 ,\AES_ENC/us00/n583 , \AES_ENC/us00/n582 , \AES_ENC/us00/n581 ,\AES_ENC/us00/n580 , \AES_ENC/us00/n579 , \AES_ENC/us00/n578 ,\AES_ENC/us00/n577 , \AES_ENC/us00/n576 , \AES_ENC/us00/n575 ,\AES_ENC/us00/n574 , \AES_ENC/us00/n573 , \AES_ENC/us00/n572 ,\AES_ENC/us00/n571 , \AES_ENC/us00/n570 , \AES_ENC/us00/n569 ,\AES_ENC/us00/n568 , \AES_ENC/us00/n567 , \AES_ENC/us00/n566 ,\AES_ENC/us00/n565 , \AES_ENC/us00/n564 , \AES_ENC/us00/n563 ,\AES_ENC/us00/n562 , \AES_ENC/us00/n561 , \AES_ENC/us00/n560 ,\AES_ENC/us00/n559 , \AES_ENC/us00/n558 , \AES_ENC/us00/n557 ,\AES_ENC/us00/n556 , \AES_ENC/us00/n555 , \AES_ENC/us00/n554 ,\AES_ENC/us00/n553 , \AES_ENC/us00/n552 , \AES_ENC/us00/n551 ,\AES_ENC/us00/n550 , \AES_ENC/us00/n549 , \AES_ENC/us00/n548 ,\AES_ENC/us00/n547 , \AES_ENC/us00/n546 , \AES_ENC/us00/n545 ,\AES_ENC/us00/n544 , \AES_ENC/us00/n543 , \AES_ENC/us00/n542 ,\AES_ENC/us00/n541 , \AES_ENC/us00/n540 , \AES_ENC/us00/n539 ,\AES_ENC/us00/n538 , \AES_ENC/us00/n537 , \AES_ENC/us00/n536 ,\AES_ENC/us00/n535 , \AES_ENC/us00/n534 , \AES_ENC/us00/n533 ,\AES_ENC/us00/n532 , \AES_ENC/us00/n531 , \AES_ENC/us00/n530 ,\AES_ENC/us00/n529 , \AES_ENC/us00/n528 , \AES_ENC/us00/n527 ,\AES_ENC/us00/n526 , \AES_ENC/us00/n525 , \AES_ENC/us00/n524 ,\AES_ENC/us00/n523 , \AES_ENC/us00/n522 , \AES_ENC/us00/n521 ,\AES_ENC/us00/n520 , \AES_ENC/us00/n519 , \AES_ENC/us00/n518 ,\AES_ENC/us00/n517 , \AES_ENC/us00/n516 , \AES_ENC/us00/n515 ,\AES_ENC/us00/n514 , \AES_ENC/us00/n513 , \AES_ENC/us00/n512 ,\AES_ENC/us00/n511 , \AES_ENC/us00/n510 , \AES_ENC/us00/n509 ,\AES_ENC/us00/n508 , \AES_ENC/us00/n507 , \AES_ENC/us00/n506 ,\AES_ENC/us00/n505 , \AES_ENC/us00/n504 , \AES_ENC/us00/n503 ,\AES_ENC/us00/n502 , \AES_ENC/us00/n501 , \AES_ENC/us00/n500 ,\AES_ENC/us00/n499 , \AES_ENC/us00/n498 , \AES_ENC/us00/n497 ,\AES_ENC/us00/n496 , \AES_ENC/us00/n495 , \AES_ENC/us00/n494 ,\AES_ENC/us00/n493 , \AES_ENC/us00/n492 , \AES_ENC/us00/n491 ,\AES_ENC/us00/n490 , \AES_ENC/us00/n489 , \AES_ENC/us00/n488 ,\AES_ENC/us00/n487 , \AES_ENC/us00/n486 , \AES_ENC/us00/n485 ,\AES_ENC/us00/n484 , \AES_ENC/us00/n483 , \AES_ENC/us00/n482 ,\AES_ENC/us00/n481 , \AES_ENC/us00/n480 , \AES_ENC/us00/n479 ,\AES_ENC/us00/n478 , \AES_ENC/us00/n477 , \AES_ENC/us00/n476 ,\AES_ENC/us00/n475 , \AES_ENC/us00/n474 , \AES_ENC/us00/n473 ,\AES_ENC/us00/n472 , \AES_ENC/us00/n471 , \AES_ENC/us00/n470 ,\AES_ENC/us00/n469 , \AES_ENC/us00/n468 , \AES_ENC/us00/n467 ,\AES_ENC/us00/n466 , \AES_ENC/us00/n465 , \AES_ENC/us00/n464 ,\AES_ENC/us00/n463 , \AES_ENC/us00/n462 , \AES_ENC/us00/n461 ,\AES_ENC/us00/n460 , \AES_ENC/us00/n459 , \AES_ENC/us00/n458 ,\AES_ENC/us00/n457 , \AES_ENC/us00/n456 , \AES_ENC/us00/n455 ,\AES_ENC/us00/n454 , \AES_ENC/us00/n453 , \AES_ENC/us00/n452 ,\AES_ENC/us00/n451 , \AES_ENC/us00/n450 , \AES_ENC/us00/n449 ,\AES_ENC/us00/n448 , \AES_ENC/us00/n447 , \AES_ENC/us00/n446 ,\AES_ENC/us00/n445 , \AES_ENC/us00/n444 , \AES_ENC/us00/n443 ,\AES_ENC/us00/n442 , \AES_ENC/us00/n441 , \AES_ENC/us00/n440 ,\AES_ENC/us00/n439 , \AES_ENC/us00/n438 , \AES_ENC/us00/n437 ,\AES_ENC/us00/n436 , \AES_ENC/us00/n435 , \AES_ENC/us00/n434 ,\AES_ENC/us00/n433 , \AES_ENC/us00/n432 , \AES_ENC/us00/n431 ,\AES_ENC/us00/n430 , \AES_ENC/us00/n429 , \AES_ENC/us00/n428 ,\AES_ENC/us00/n427 , \AES_ENC/us00/n426 , \AES_ENC/us00/n425 ,\AES_ENC/us00/n424 , \AES_ENC/us00/n423 , \AES_ENC/us00/n422 ,\AES_ENC/us00/n421 , \AES_ENC/us00/n420 , \AES_ENC/us00/n419 ,\AES_ENC/us00/n418 , \AES_ENC/us00/n417 , \AES_ENC/us00/n416 ,\AES_ENC/us00/n415 , \AES_ENC/us00/n414 , \AES_ENC/us00/n413 ,\AES_ENC/us00/n412 , \AES_ENC/us00/n411 , \AES_ENC/us00/n410 ,\AES_ENC/us00/n409 , \AES_ENC/us00/n408 , \AES_ENC/us00/n407 ,\AES_ENC/us00/n406 , \AES_ENC/us00/n405 , \AES_ENC/us00/n404 ,\AES_ENC/us00/n403 , \AES_ENC/us00/n402 , \AES_ENC/us00/n401 ,\AES_ENC/us00/n400 , \AES_ENC/us00/n399 , \AES_ENC/us00/n398 ,\AES_ENC/us00/n397 , \AES_ENC/us00/n396 , \AES_ENC/us00/n395 ,\AES_ENC/us00/n394 , \AES_ENC/us00/n393 , \AES_ENC/us00/n392 ,\AES_ENC/us00/n391 , \AES_ENC/us00/n390 , \AES_ENC/us00/n389 ,\AES_ENC/us00/n388 , \AES_ENC/us00/n387 , \AES_ENC/us00/n386 ,\AES_ENC/us00/n385 , \AES_ENC/us00/n384 , \AES_ENC/us00/n383 ,\AES_ENC/us00/n382 , \AES_ENC/us00/n381 , \AES_ENC/us00/n380 ,\AES_ENC/us00/n379 , \AES_ENC/us00/n378 , \AES_ENC/us00/n377 ,\AES_ENC/us00/n376 , \AES_ENC/us00/n375 , \AES_ENC/us00/n374 ,\AES_ENC/us00/n373 , \AES_ENC/us00/n372 , \AES_ENC/us00/n371 ,\AES_ENC/us00/n370 , \AES_ENC/us00/n369 , \AES_ENC/us00/n368 ,\AES_ENC/us00/n367 , \AES_ENC/us00/n366 , \AES_ENC/us00/n365 ,\AES_ENC/us00/n364 , \AES_ENC/us00/n363 , \AES_ENC/us00/n362 ,\AES_ENC/us00/n361 , \AES_ENC/us00/n360 , \AES_ENC/us00/n359 ,\AES_ENC/us00/n358 , \AES_ENC/us00/n357 , \AES_ENC/us00/n356 ,\AES_ENC/us00/n355 , \AES_ENC/us00/n354 , \AES_ENC/us00/n353 ,\AES_ENC/us00/n352 , \AES_ENC/us00/n351 , \AES_ENC/us00/n350 ,\AES_ENC/us00/n349 , \AES_ENC/us00/n348 , \AES_ENC/us00/n347 ,\AES_ENC/us00/n346 , \AES_ENC/us00/n345 , \AES_ENC/us00/n344 ,\AES_ENC/us00/n343 , \AES_ENC/us00/n342 , \AES_ENC/us00/n341 ,\AES_ENC/us00/n340 , \AES_ENC/us00/n339 , \AES_ENC/us00/n338 ,\AES_ENC/us00/n337 , \AES_ENC/us00/n336 , \AES_ENC/us00/n335 ,\AES_ENC/us00/n334 , \AES_ENC/us00/n333 , \AES_ENC/us00/n332 ,\AES_ENC/us00/n331 , \AES_ENC/us00/n330 , \AES_ENC/us00/n329 ,\AES_ENC/us00/n328 , \AES_ENC/us00/n327 , \AES_ENC/us00/n326 ,\AES_ENC/us00/n325 , \AES_ENC/us00/n324 , \AES_ENC/us00/n323 ,\AES_ENC/us00/n322 , \AES_ENC/us00/n321 , \AES_ENC/us00/n320 ,\AES_ENC/us00/n319 , \AES_ENC/us00/n318 , \AES_ENC/us00/n317 ,\AES_ENC/us00/n316 , \AES_ENC/us00/n315 , \AES_ENC/us00/n314 ,\AES_ENC/us00/n313 , \AES_ENC/us00/n312 , \AES_ENC/us00/n311 ,\AES_ENC/us00/n310 , \AES_ENC/us00/n309 , \AES_ENC/us00/n308 ,\AES_ENC/us00/n307 , \AES_ENC/us00/n306 , \AES_ENC/us00/n305 ,\AES_ENC/us00/n304 , \AES_ENC/us00/n303 , \AES_ENC/us00/n302 ,\AES_ENC/us00/n301 , \AES_ENC/us00/n300 , \AES_ENC/us00/n299 ,\AES_ENC/us00/n298 , \AES_ENC/us00/n297 , \AES_ENC/us00/n296 ,\AES_ENC/us00/n295 , \AES_ENC/us00/n294 , \AES_ENC/us00/n293 ,\AES_ENC/us00/n292 , \AES_ENC/us00/n291 , \AES_ENC/us00/n290 ,\AES_ENC/us00/n289 , \AES_ENC/us00/n288 , \AES_ENC/us00/n287 ,\AES_ENC/us00/n286 , \AES_ENC/us00/n285 , \AES_ENC/us00/n284 ,\AES_ENC/us00/n283 , \AES_ENC/us00/n282 , \AES_ENC/us00/n281 ,\AES_ENC/us00/n280 , \AES_ENC/us00/n279 , \AES_ENC/us00/n278 ,\AES_ENC/us00/n277 , \AES_ENC/us00/n276 , \AES_ENC/us00/n275 ,\AES_ENC/us00/n274 , \AES_ENC/us00/n273 , \AES_ENC/us00/n272 ,\AES_ENC/us00/n271 , \AES_ENC/us00/n270 , \AES_ENC/us00/n269 ,\AES_ENC/us00/n268 , \AES_ENC/us00/n267 , \AES_ENC/us00/n266 ,\AES_ENC/us00/n265 , \AES_ENC/us00/n264 , \AES_ENC/us00/n263 ,\AES_ENC/us00/n262 , \AES_ENC/us00/n261 , \AES_ENC/us00/n260 ,\AES_ENC/us00/n259 , \AES_ENC/us00/n258 , \AES_ENC/us00/n257 ,\AES_ENC/us00/n256 , \AES_ENC/us00/n255 , \AES_ENC/us00/n254 ,\AES_ENC/us00/n253 , \AES_ENC/us00/n252 , \AES_ENC/us00/n251 ,\AES_ENC/us00/n250 , \AES_ENC/us00/n249 , \AES_ENC/us00/n248 ,\AES_ENC/us00/n247 , \AES_ENC/us00/n246 , \AES_ENC/us00/n245 ,\AES_ENC/us00/n244 , \AES_ENC/us00/n243 , \AES_ENC/us00/n242 ,\AES_ENC/us00/n241 , \AES_ENC/us00/n240 , \AES_ENC/us00/n239 ,\AES_ENC/us00/n238 , \AES_ENC/us00/n237 , \AES_ENC/us00/n235 ,\AES_ENC/us00/n234 , \AES_ENC/us00/n233 , \AES_ENC/us00/n232 ,\AES_ENC/us00/n231 , \AES_ENC/us00/n230 , \AES_ENC/us00/n229 ,\AES_ENC/us00/n228 , \AES_ENC/us00/n227 , \AES_ENC/us00/n226 ,\AES_ENC/us00/n225 , \AES_ENC/us00/n224 , \AES_ENC/us00/n223 ,\AES_ENC/us00/n222 , \AES_ENC/us00/n221 , \AES_ENC/us00/n220 ,\AES_ENC/us00/n219 , \AES_ENC/us00/n218 , \AES_ENC/us00/n217 ,\AES_ENC/us00/n216 , \AES_ENC/us00/n215 , \AES_ENC/us00/n214 ,\AES_ENC/us00/n213 , \AES_ENC/us00/n212 , \AES_ENC/us00/n211 ,\AES_ENC/us00/n210 , \AES_ENC/us00/n209 , \AES_ENC/us00/n208 ,\AES_ENC/us00/n207 , \AES_ENC/us00/n206 , \AES_ENC/us00/n205 ,\AES_ENC/us00/n204 , \AES_ENC/us00/n203 , \AES_ENC/us00/n202 ,\AES_ENC/us00/n201 , \AES_ENC/us00/n200 , \AES_ENC/us00/n199 ,\AES_ENC/us00/n198 , \AES_ENC/us00/n197 , \AES_ENC/us00/n196 ,\AES_ENC/us00/n195 , \AES_ENC/us00/n194 , \AES_ENC/us00/n193 ,\AES_ENC/us00/n192 , \AES_ENC/us00/n191 , \AES_ENC/us00/n190 ,\AES_ENC/us00/n189 , \AES_ENC/us00/n188 , \AES_ENC/us00/n187 ,\AES_ENC/us00/n186 , \AES_ENC/us00/n185 , \AES_ENC/us00/n184 ,\AES_ENC/us00/n183 , \AES_ENC/us00/n182 , \AES_ENC/us00/n181 ,\AES_ENC/us00/n180 , \AES_ENC/us00/n179 , \AES_ENC/us00/n178 ,\AES_ENC/us00/n177 , \AES_ENC/us00/n176 , \AES_ENC/us00/n175 ,\AES_ENC/us00/n174 , \AES_ENC/us00/n173 , \AES_ENC/us00/n172 ,\AES_ENC/us00/n171 , \AES_ENC/us00/n170 , \AES_ENC/us00/n168 ,\AES_ENC/us00/n167 , \AES_ENC/us00/n166 , \AES_ENC/us00/n165 ,\AES_ENC/us00/n164 , \AES_ENC/us00/n163 , \AES_ENC/us00/n162 ,\AES_ENC/us00/n161 , \AES_ENC/us00/n160 , \AES_ENC/us00/n159 ,\AES_ENC/us00/n158 , \AES_ENC/us00/n157 , \AES_ENC/us00/n156 ,\AES_ENC/us00/n155 , \AES_ENC/us00/n154 , \AES_ENC/us00/n153 ,\AES_ENC/us00/n152 , \AES_ENC/us00/n151 , \AES_ENC/us00/n150 ,\AES_ENC/us00/n149 , \AES_ENC/us00/n148 , \AES_ENC/us00/n147 ,\AES_ENC/us00/n146 , \AES_ENC/us00/n145 , \AES_ENC/us00/n144 ,\AES_ENC/us00/n143 , \AES_ENC/us00/n142 , \AES_ENC/us00/n141 ,\AES_ENC/us00/n140 , \AES_ENC/us00/n139 , \AES_ENC/us00/n138 ,\AES_ENC/us00/n137 , \AES_ENC/us00/n136 , \AES_ENC/us00/n135 ,\AES_ENC/us00/n134 , \AES_ENC/us00/n133 , \AES_ENC/us00/n132 ,\AES_ENC/us00/n131 , \AES_ENC/us00/n130 , \AES_ENC/us00/n129 ,\AES_ENC/us00/n128 , \AES_ENC/us00/n127 , \AES_ENC/us00/n126 ,\AES_ENC/us00/n125 , \AES_ENC/us00/n124 , \AES_ENC/us00/n123 ,\AES_ENC/us00/n122 , \AES_ENC/us00/n121 , \AES_ENC/us00/n120 ,\AES_ENC/us00/n119 , \AES_ENC/us00/n118 , \AES_ENC/us00/n117 ,\AES_ENC/us00/n116 , \AES_ENC/us00/n115 , \AES_ENC/us00/n114 ,\AES_ENC/us00/n113 , \AES_ENC/us00/n112 , \AES_ENC/us00/n111 ,\AES_ENC/us00/n110 , \AES_ENC/us00/n109 , \AES_ENC/us00/n108 ,\AES_ENC/us00/n107 , \AES_ENC/us00/n106 , \AES_ENC/us00/n105 ,\AES_ENC/us00/n104 , \AES_ENC/us00/n103 , \AES_ENC/us00/n102 ,\AES_ENC/us00/n101 , \AES_ENC/us00/n100 , \AES_ENC/us00/n99 ,\AES_ENC/us00/n97 , \AES_ENC/us00/n96 , \AES_ENC/us00/n95 ,\AES_ENC/us00/n94 , \AES_ENC/us00/n93 , \AES_ENC/us00/n92 ,\AES_ENC/us00/n91 , \AES_ENC/us00/n90 , \AES_ENC/us00/n89 ,\AES_ENC/us00/n88 , \AES_ENC/us00/n87 , \AES_ENC/us00/n86 ,\AES_ENC/us00/n85 , \AES_ENC/us00/n84 , \AES_ENC/us00/n83 ,\AES_ENC/us00/n82 , \AES_ENC/us00/n81 , \AES_ENC/us00/n80 ,\AES_ENC/us00/n79 , \AES_ENC/us00/n78 , \AES_ENC/us00/n77 ,\AES_ENC/us00/n76 , \AES_ENC/us00/n75 , \AES_ENC/us00/n74 ,\AES_ENC/us00/n73 , \AES_ENC/us00/n72 , \AES_ENC/us00/n71 ,\AES_ENC/us00/n70 , \AES_ENC/us00/n69 , \AES_ENC/us00/n68 ,\AES_ENC/us00/n67 , \AES_ENC/us00/n66 , \AES_ENC/us00/n65 ,\AES_ENC/us00/n64 , \AES_ENC/us00/n63 , \AES_ENC/us00/n62 ,\AES_ENC/us00/n61 , \AES_ENC/us00/n60 , \AES_ENC/us00/n59 ,\AES_ENC/us00/n58 , \AES_ENC/us01/n1135 , \AES_ENC/us01/n1134 ,\AES_ENC/us01/n1133 , \AES_ENC/us01/n1132 , \AES_ENC/us01/n1131 ,\AES_ENC/us01/n1130 , \AES_ENC/us01/n1129 , \AES_ENC/us01/n1128 ,\AES_ENC/us01/n1127 , \AES_ENC/us01/n1126 , \AES_ENC/us01/n1125 ,\AES_ENC/us01/n1124 , \AES_ENC/us01/n1123 , \AES_ENC/us01/n1122 ,\AES_ENC/us01/n1121 , \AES_ENC/us01/n1120 , \AES_ENC/us01/n1119 ,\AES_ENC/us01/n1118 , \AES_ENC/us01/n1117 , \AES_ENC/us01/n1116 ,\AES_ENC/us01/n1115 , \AES_ENC/us01/n1114 , \AES_ENC/us01/n1113 ,\AES_ENC/us01/n1112 , \AES_ENC/us01/n1111 , \AES_ENC/us01/n1110 ,\AES_ENC/us01/n1109 , \AES_ENC/us01/n1108 , \AES_ENC/us01/n1107 ,\AES_ENC/us01/n1106 , \AES_ENC/us01/n1105 , \AES_ENC/us01/n1104 ,\AES_ENC/us01/n1103 , \AES_ENC/us01/n1102 , \AES_ENC/us01/n1101 ,\AES_ENC/us01/n1100 , \AES_ENC/us01/n1099 , \AES_ENC/us01/n1098 ,\AES_ENC/us01/n1097 , \AES_ENC/us01/n1096 , \AES_ENC/us01/n1095 ,\AES_ENC/us01/n1094 , \AES_ENC/us01/n1093 , \AES_ENC/us01/n1092 ,\AES_ENC/us01/n1091 , \AES_ENC/us01/n1090 , \AES_ENC/us01/n1089 ,\AES_ENC/us01/n1088 , \AES_ENC/us01/n1087 , \AES_ENC/us01/n1086 ,\AES_ENC/us01/n1085 , \AES_ENC/us01/n1084 , \AES_ENC/us01/n1083 ,\AES_ENC/us01/n1082 , \AES_ENC/us01/n1081 , \AES_ENC/us01/n1080 ,\AES_ENC/us01/n1079 , \AES_ENC/us01/n1078 , \AES_ENC/us01/n1077 ,\AES_ENC/us01/n1076 , \AES_ENC/us01/n1075 , \AES_ENC/us01/n1074 ,\AES_ENC/us01/n1073 , \AES_ENC/us01/n1072 , \AES_ENC/us01/n1071 ,\AES_ENC/us01/n1070 , \AES_ENC/us01/n1069 , \AES_ENC/us01/n1068 ,\AES_ENC/us01/n1067 , \AES_ENC/us01/n1066 , \AES_ENC/us01/n1065 ,\AES_ENC/us01/n1064 , \AES_ENC/us01/n1063 , \AES_ENC/us01/n1062 ,\AES_ENC/us01/n1061 , \AES_ENC/us01/n1060 , \AES_ENC/us01/n1059 ,\AES_ENC/us01/n1058 , \AES_ENC/us01/n1057 , \AES_ENC/us01/n1056 ,\AES_ENC/us01/n1055 , \AES_ENC/us01/n1054 , \AES_ENC/us01/n1053 ,\AES_ENC/us01/n1052 , \AES_ENC/us01/n1051 , \AES_ENC/us01/n1050 ,\AES_ENC/us01/n1049 , \AES_ENC/us01/n1048 , \AES_ENC/us01/n1047 ,\AES_ENC/us01/n1046 , \AES_ENC/us01/n1045 , \AES_ENC/us01/n1044 ,\AES_ENC/us01/n1043 , \AES_ENC/us01/n1042 , \AES_ENC/us01/n1041 ,\AES_ENC/us01/n1040 , \AES_ENC/us01/n1039 , \AES_ENC/us01/n1038 ,\AES_ENC/us01/n1037 , \AES_ENC/us01/n1036 , \AES_ENC/us01/n1035 ,\AES_ENC/us01/n1034 , \AES_ENC/us01/n1033 , \AES_ENC/us01/n1032 ,\AES_ENC/us01/n1031 , \AES_ENC/us01/n1030 , \AES_ENC/us01/n1029 ,\AES_ENC/us01/n1028 , \AES_ENC/us01/n1027 , \AES_ENC/us01/n1026 ,\AES_ENC/us01/n1025 , \AES_ENC/us01/n1024 , \AES_ENC/us01/n1023 ,\AES_ENC/us01/n1022 , \AES_ENC/us01/n1021 , \AES_ENC/us01/n1020 ,\AES_ENC/us01/n1019 , \AES_ENC/us01/n1018 , \AES_ENC/us01/n1017 ,\AES_ENC/us01/n1016 , \AES_ENC/us01/n1015 , \AES_ENC/us01/n1014 ,\AES_ENC/us01/n1013 , \AES_ENC/us01/n1012 , \AES_ENC/us01/n1011 ,\AES_ENC/us01/n1010 , \AES_ENC/us01/n1009 , \AES_ENC/us01/n1008 ,\AES_ENC/us01/n1007 , \AES_ENC/us01/n1006 , \AES_ENC/us01/n1005 ,\AES_ENC/us01/n1004 , \AES_ENC/us01/n1003 , \AES_ENC/us01/n1002 ,\AES_ENC/us01/n1001 , \AES_ENC/us01/n1000 , \AES_ENC/us01/n999 ,\AES_ENC/us01/n998 , \AES_ENC/us01/n997 , \AES_ENC/us01/n996 ,\AES_ENC/us01/n995 , \AES_ENC/us01/n994 , \AES_ENC/us01/n993 ,\AES_ENC/us01/n992 , \AES_ENC/us01/n991 , \AES_ENC/us01/n990 ,\AES_ENC/us01/n989 , \AES_ENC/us01/n988 , \AES_ENC/us01/n987 ,\AES_ENC/us01/n986 , \AES_ENC/us01/n985 , \AES_ENC/us01/n984 ,\AES_ENC/us01/n983 , \AES_ENC/us01/n982 , \AES_ENC/us01/n981 ,\AES_ENC/us01/n980 , \AES_ENC/us01/n979 , \AES_ENC/us01/n978 ,\AES_ENC/us01/n977 , \AES_ENC/us01/n976 , \AES_ENC/us01/n975 ,\AES_ENC/us01/n974 , \AES_ENC/us01/n973 , \AES_ENC/us01/n972 ,\AES_ENC/us01/n971 , \AES_ENC/us01/n970 , \AES_ENC/us01/n969 ,\AES_ENC/us01/n968 , \AES_ENC/us01/n967 , \AES_ENC/us01/n966 ,\AES_ENC/us01/n965 , \AES_ENC/us01/n964 , \AES_ENC/us01/n963 ,\AES_ENC/us01/n962 , \AES_ENC/us01/n961 , \AES_ENC/us01/n960 ,\AES_ENC/us01/n959 , \AES_ENC/us01/n958 , \AES_ENC/us01/n957 ,\AES_ENC/us01/n956 , \AES_ENC/us01/n955 , \AES_ENC/us01/n954 ,\AES_ENC/us01/n953 , \AES_ENC/us01/n952 , \AES_ENC/us01/n951 ,\AES_ENC/us01/n950 , \AES_ENC/us01/n949 , \AES_ENC/us01/n948 ,\AES_ENC/us01/n947 , \AES_ENC/us01/n946 , \AES_ENC/us01/n945 ,\AES_ENC/us01/n944 , \AES_ENC/us01/n943 , \AES_ENC/us01/n942 ,\AES_ENC/us01/n941 , \AES_ENC/us01/n940 , \AES_ENC/us01/n939 ,\AES_ENC/us01/n938 , \AES_ENC/us01/n937 , \AES_ENC/us01/n936 ,\AES_ENC/us01/n935 , \AES_ENC/us01/n934 , \AES_ENC/us01/n933 ,\AES_ENC/us01/n932 , \AES_ENC/us01/n931 , \AES_ENC/us01/n930 ,\AES_ENC/us01/n929 , \AES_ENC/us01/n928 , \AES_ENC/us01/n927 ,\AES_ENC/us01/n926 , \AES_ENC/us01/n925 , \AES_ENC/us01/n924 ,\AES_ENC/us01/n923 , \AES_ENC/us01/n922 , \AES_ENC/us01/n921 ,\AES_ENC/us01/n920 , \AES_ENC/us01/n919 , \AES_ENC/us01/n918 ,\AES_ENC/us01/n917 , \AES_ENC/us01/n916 , \AES_ENC/us01/n915 ,\AES_ENC/us01/n914 , \AES_ENC/us01/n913 , \AES_ENC/us01/n912 ,\AES_ENC/us01/n911 , \AES_ENC/us01/n910 , \AES_ENC/us01/n909 ,\AES_ENC/us01/n908 , \AES_ENC/us01/n907 , \AES_ENC/us01/n906 ,\AES_ENC/us01/n905 , \AES_ENC/us01/n904 , \AES_ENC/us01/n903 ,\AES_ENC/us01/n902 , \AES_ENC/us01/n901 , \AES_ENC/us01/n900 ,\AES_ENC/us01/n899 , \AES_ENC/us01/n898 , \AES_ENC/us01/n897 ,\AES_ENC/us01/n896 , \AES_ENC/us01/n895 , \AES_ENC/us01/n894 ,\AES_ENC/us01/n893 , \AES_ENC/us01/n892 , \AES_ENC/us01/n891 ,\AES_ENC/us01/n890 , \AES_ENC/us01/n889 , \AES_ENC/us01/n888 ,\AES_ENC/us01/n887 , \AES_ENC/us01/n886 , \AES_ENC/us01/n885 ,\AES_ENC/us01/n884 , \AES_ENC/us01/n883 , \AES_ENC/us01/n882 ,\AES_ENC/us01/n881 , \AES_ENC/us01/n880 , \AES_ENC/us01/n879 ,\AES_ENC/us01/n878 , \AES_ENC/us01/n877 , \AES_ENC/us01/n876 ,\AES_ENC/us01/n875 , \AES_ENC/us01/n874 , \AES_ENC/us01/n873 ,\AES_ENC/us01/n872 , \AES_ENC/us01/n871 , \AES_ENC/us01/n870 ,\AES_ENC/us01/n869 , \AES_ENC/us01/n868 , \AES_ENC/us01/n867 ,\AES_ENC/us01/n866 , \AES_ENC/us01/n865 , \AES_ENC/us01/n864 ,\AES_ENC/us01/n863 , \AES_ENC/us01/n862 , \AES_ENC/us01/n861 ,\AES_ENC/us01/n860 , \AES_ENC/us01/n859 , \AES_ENC/us01/n858 ,\AES_ENC/us01/n857 , \AES_ENC/us01/n856 , \AES_ENC/us01/n855 ,\AES_ENC/us01/n854 , \AES_ENC/us01/n853 , \AES_ENC/us01/n852 ,\AES_ENC/us01/n851 , \AES_ENC/us01/n850 , \AES_ENC/us01/n849 ,\AES_ENC/us01/n848 , \AES_ENC/us01/n847 , \AES_ENC/us01/n846 ,\AES_ENC/us01/n845 , \AES_ENC/us01/n844 , \AES_ENC/us01/n843 ,\AES_ENC/us01/n842 , \AES_ENC/us01/n841 , \AES_ENC/us01/n840 ,\AES_ENC/us01/n839 , \AES_ENC/us01/n838 , \AES_ENC/us01/n837 ,\AES_ENC/us01/n836 , \AES_ENC/us01/n835 , \AES_ENC/us01/n834 ,\AES_ENC/us01/n833 , \AES_ENC/us01/n832 , \AES_ENC/us01/n831 ,\AES_ENC/us01/n830 , \AES_ENC/us01/n829 , \AES_ENC/us01/n828 ,\AES_ENC/us01/n827 , \AES_ENC/us01/n826 , \AES_ENC/us01/n825 ,\AES_ENC/us01/n824 , \AES_ENC/us01/n823 , \AES_ENC/us01/n822 ,\AES_ENC/us01/n821 , \AES_ENC/us01/n820 , \AES_ENC/us01/n819 ,\AES_ENC/us01/n818 , \AES_ENC/us01/n817 , \AES_ENC/us01/n816 ,\AES_ENC/us01/n815 , \AES_ENC/us01/n814 , \AES_ENC/us01/n813 ,\AES_ENC/us01/n812 , \AES_ENC/us01/n811 , \AES_ENC/us01/n810 ,\AES_ENC/us01/n809 , \AES_ENC/us01/n808 , \AES_ENC/us01/n807 ,\AES_ENC/us01/n806 , \AES_ENC/us01/n805 , \AES_ENC/us01/n804 ,\AES_ENC/us01/n803 , \AES_ENC/us01/n802 , \AES_ENC/us01/n801 ,\AES_ENC/us01/n800 , \AES_ENC/us01/n799 , \AES_ENC/us01/n798 ,\AES_ENC/us01/n797 , \AES_ENC/us01/n796 , \AES_ENC/us01/n795 ,\AES_ENC/us01/n794 , \AES_ENC/us01/n793 , \AES_ENC/us01/n792 ,\AES_ENC/us01/n791 , \AES_ENC/us01/n790 , \AES_ENC/us01/n789 ,\AES_ENC/us01/n788 , \AES_ENC/us01/n787 , \AES_ENC/us01/n786 ,\AES_ENC/us01/n785 , \AES_ENC/us01/n784 , \AES_ENC/us01/n783 ,\AES_ENC/us01/n782 , \AES_ENC/us01/n781 , \AES_ENC/us01/n780 ,\AES_ENC/us01/n779 , \AES_ENC/us01/n778 , \AES_ENC/us01/n777 ,\AES_ENC/us01/n776 , \AES_ENC/us01/n775 , \AES_ENC/us01/n774 ,\AES_ENC/us01/n773 , \AES_ENC/us01/n772 , \AES_ENC/us01/n771 ,\AES_ENC/us01/n770 , \AES_ENC/us01/n769 , \AES_ENC/us01/n768 ,\AES_ENC/us01/n767 , \AES_ENC/us01/n766 , \AES_ENC/us01/n765 ,\AES_ENC/us01/n764 , \AES_ENC/us01/n763 , \AES_ENC/us01/n762 ,\AES_ENC/us01/n761 , \AES_ENC/us01/n760 , \AES_ENC/us01/n759 ,\AES_ENC/us01/n758 , \AES_ENC/us01/n757 , \AES_ENC/us01/n756 ,\AES_ENC/us01/n755 , \AES_ENC/us01/n754 , \AES_ENC/us01/n753 ,\AES_ENC/us01/n752 , \AES_ENC/us01/n751 , \AES_ENC/us01/n750 ,\AES_ENC/us01/n749 , \AES_ENC/us01/n748 , \AES_ENC/us01/n747 ,\AES_ENC/us01/n746 , \AES_ENC/us01/n745 , \AES_ENC/us01/n744 ,\AES_ENC/us01/n743 , \AES_ENC/us01/n742 , \AES_ENC/us01/n741 ,\AES_ENC/us01/n740 , \AES_ENC/us01/n739 , \AES_ENC/us01/n738 ,\AES_ENC/us01/n737 , \AES_ENC/us01/n736 , \AES_ENC/us01/n735 ,\AES_ENC/us01/n734 , \AES_ENC/us01/n733 , \AES_ENC/us01/n732 ,\AES_ENC/us01/n731 , \AES_ENC/us01/n730 , \AES_ENC/us01/n729 ,\AES_ENC/us01/n728 , \AES_ENC/us01/n727 , \AES_ENC/us01/n726 ,\AES_ENC/us01/n725 , \AES_ENC/us01/n724 , \AES_ENC/us01/n723 ,\AES_ENC/us01/n722 , \AES_ENC/us01/n721 , \AES_ENC/us01/n720 ,\AES_ENC/us01/n719 , \AES_ENC/us01/n718 , \AES_ENC/us01/n717 ,\AES_ENC/us01/n716 , \AES_ENC/us01/n715 , \AES_ENC/us01/n714 ,\AES_ENC/us01/n713 , \AES_ENC/us01/n712 , \AES_ENC/us01/n711 ,\AES_ENC/us01/n710 , \AES_ENC/us01/n709 , \AES_ENC/us01/n708 ,\AES_ENC/us01/n707 , \AES_ENC/us01/n706 , \AES_ENC/us01/n705 ,\AES_ENC/us01/n704 , \AES_ENC/us01/n703 , \AES_ENC/us01/n702 ,\AES_ENC/us01/n701 , \AES_ENC/us01/n700 , \AES_ENC/us01/n699 ,\AES_ENC/us01/n698 , \AES_ENC/us01/n697 , \AES_ENC/us01/n696 ,\AES_ENC/us01/n695 , \AES_ENC/us01/n694 , \AES_ENC/us01/n693 ,\AES_ENC/us01/n692 , \AES_ENC/us01/n691 , \AES_ENC/us01/n690 ,\AES_ENC/us01/n689 , \AES_ENC/us01/n688 , \AES_ENC/us01/n687 ,\AES_ENC/us01/n686 , \AES_ENC/us01/n685 , \AES_ENC/us01/n684 ,\AES_ENC/us01/n683 , \AES_ENC/us01/n682 , \AES_ENC/us01/n681 ,\AES_ENC/us01/n680 , \AES_ENC/us01/n679 , \AES_ENC/us01/n678 ,\AES_ENC/us01/n677 , \AES_ENC/us01/n676 , \AES_ENC/us01/n675 ,\AES_ENC/us01/n674 , \AES_ENC/us01/n673 , \AES_ENC/us01/n672 ,\AES_ENC/us01/n671 , \AES_ENC/us01/n670 , \AES_ENC/us01/n669 ,\AES_ENC/us01/n668 , \AES_ENC/us01/n667 , \AES_ENC/us01/n666 ,\AES_ENC/us01/n665 , \AES_ENC/us01/n664 , \AES_ENC/us01/n663 ,\AES_ENC/us01/n662 , \AES_ENC/us01/n661 , \AES_ENC/us01/n660 ,\AES_ENC/us01/n659 , \AES_ENC/us01/n658 , \AES_ENC/us01/n657 ,\AES_ENC/us01/n656 , \AES_ENC/us01/n655 , \AES_ENC/us01/n654 ,\AES_ENC/us01/n653 , \AES_ENC/us01/n652 , \AES_ENC/us01/n651 ,\AES_ENC/us01/n650 , \AES_ENC/us01/n649 , \AES_ENC/us01/n648 ,\AES_ENC/us01/n647 , \AES_ENC/us01/n646 , \AES_ENC/us01/n645 ,\AES_ENC/us01/n644 , \AES_ENC/us01/n643 , \AES_ENC/us01/n642 ,\AES_ENC/us01/n641 , \AES_ENC/us01/n640 , \AES_ENC/us01/n639 ,\AES_ENC/us01/n638 , \AES_ENC/us01/n637 , \AES_ENC/us01/n636 ,\AES_ENC/us01/n635 , \AES_ENC/us01/n634 , \AES_ENC/us01/n633 ,\AES_ENC/us01/n632 , \AES_ENC/us01/n631 , \AES_ENC/us01/n630 ,\AES_ENC/us01/n629 , \AES_ENC/us01/n628 , \AES_ENC/us01/n627 ,\AES_ENC/us01/n626 , \AES_ENC/us01/n625 , \AES_ENC/us01/n624 ,\AES_ENC/us01/n623 , \AES_ENC/us01/n622 , \AES_ENC/us01/n621 ,\AES_ENC/us01/n620 , \AES_ENC/us01/n619 , \AES_ENC/us01/n618 ,\AES_ENC/us01/n617 , \AES_ENC/us01/n616 , \AES_ENC/us01/n615 ,\AES_ENC/us01/n614 , \AES_ENC/us01/n613 , \AES_ENC/us01/n612 ,\AES_ENC/us01/n611 , \AES_ENC/us01/n610 , \AES_ENC/us01/n609 ,\AES_ENC/us01/n608 , \AES_ENC/us01/n607 , \AES_ENC/us01/n606 ,\AES_ENC/us01/n605 , \AES_ENC/us01/n604 , \AES_ENC/us01/n603 ,\AES_ENC/us01/n602 , \AES_ENC/us01/n601 , \AES_ENC/us01/n600 ,\AES_ENC/us01/n599 , \AES_ENC/us01/n598 , \AES_ENC/us01/n597 ,\AES_ENC/us01/n596 , \AES_ENC/us01/n595 , \AES_ENC/us01/n594 ,\AES_ENC/us01/n593 , \AES_ENC/us01/n592 , \AES_ENC/us01/n591 ,\AES_ENC/us01/n590 , \AES_ENC/us01/n589 , \AES_ENC/us01/n588 ,\AES_ENC/us01/n587 , \AES_ENC/us01/n586 , \AES_ENC/us01/n585 ,\AES_ENC/us01/n584 , \AES_ENC/us01/n583 , \AES_ENC/us01/n582 ,\AES_ENC/us01/n581 , \AES_ENC/us01/n580 , \AES_ENC/us01/n579 ,\AES_ENC/us01/n578 , \AES_ENC/us01/n577 , \AES_ENC/us01/n576 ,\AES_ENC/us01/n575 , \AES_ENC/us01/n574 , \AES_ENC/us01/n573 ,\AES_ENC/us01/n572 , \AES_ENC/us01/n571 , \AES_ENC/us01/n570 ,\AES_ENC/us01/n569 , \AES_ENC/us02/n1135 , \AES_ENC/us02/n1134 ,\AES_ENC/us02/n1133 , \AES_ENC/us02/n1132 , \AES_ENC/us02/n1131 ,\AES_ENC/us02/n1130 , \AES_ENC/us02/n1129 , \AES_ENC/us02/n1128 ,\AES_ENC/us02/n1127 , \AES_ENC/us02/n1126 , \AES_ENC/us02/n1125 ,\AES_ENC/us02/n1124 , \AES_ENC/us02/n1123 , \AES_ENC/us02/n1122 ,\AES_ENC/us02/n1121 , \AES_ENC/us02/n1120 , \AES_ENC/us02/n1119 ,\AES_ENC/us02/n1118 , \AES_ENC/us02/n1117 , \AES_ENC/us02/n1116 ,\AES_ENC/us02/n1115 , \AES_ENC/us02/n1114 , \AES_ENC/us02/n1113 ,\AES_ENC/us02/n1112 , \AES_ENC/us02/n1111 , \AES_ENC/us02/n1110 ,\AES_ENC/us02/n1109 , \AES_ENC/us02/n1108 , \AES_ENC/us02/n1107 ,\AES_ENC/us02/n1106 , \AES_ENC/us02/n1105 , \AES_ENC/us02/n1104 ,\AES_ENC/us02/n1103 , \AES_ENC/us02/n1102 , \AES_ENC/us02/n1101 ,\AES_ENC/us02/n1100 , \AES_ENC/us02/n1099 , \AES_ENC/us02/n1098 ,\AES_ENC/us02/n1097 , \AES_ENC/us02/n1096 , \AES_ENC/us02/n1095 ,\AES_ENC/us02/n1094 , \AES_ENC/us02/n1093 , \AES_ENC/us02/n1092 ,\AES_ENC/us02/n1091 , \AES_ENC/us02/n1090 , \AES_ENC/us02/n1089 ,\AES_ENC/us02/n1088 , \AES_ENC/us02/n1087 , \AES_ENC/us02/n1086 ,\AES_ENC/us02/n1085 , \AES_ENC/us02/n1084 , \AES_ENC/us02/n1083 ,\AES_ENC/us02/n1082 , \AES_ENC/us02/n1081 , \AES_ENC/us02/n1080 ,\AES_ENC/us02/n1079 , \AES_ENC/us02/n1078 , \AES_ENC/us02/n1077 ,\AES_ENC/us02/n1076 , \AES_ENC/us02/n1075 , \AES_ENC/us02/n1074 ,\AES_ENC/us02/n1073 , \AES_ENC/us02/n1072 , \AES_ENC/us02/n1071 ,\AES_ENC/us02/n1070 , \AES_ENC/us02/n1069 , \AES_ENC/us02/n1068 ,\AES_ENC/us02/n1067 , \AES_ENC/us02/n1066 , \AES_ENC/us02/n1065 ,\AES_ENC/us02/n1064 , \AES_ENC/us02/n1063 , \AES_ENC/us02/n1062 ,\AES_ENC/us02/n1061 , \AES_ENC/us02/n1060 , \AES_ENC/us02/n1059 ,\AES_ENC/us02/n1058 , \AES_ENC/us02/n1057 , \AES_ENC/us02/n1056 ,\AES_ENC/us02/n1055 , \AES_ENC/us02/n1054 , \AES_ENC/us02/n1053 ,\AES_ENC/us02/n1052 , \AES_ENC/us02/n1051 , \AES_ENC/us02/n1050 ,\AES_ENC/us02/n1049 , \AES_ENC/us02/n1048 , \AES_ENC/us02/n1047 ,\AES_ENC/us02/n1046 , \AES_ENC/us02/n1045 , \AES_ENC/us02/n1044 ,\AES_ENC/us02/n1043 , \AES_ENC/us02/n1042 , \AES_ENC/us02/n1041 ,\AES_ENC/us02/n1040 , \AES_ENC/us02/n1039 , \AES_ENC/us02/n1038 ,\AES_ENC/us02/n1037 , \AES_ENC/us02/n1036 , \AES_ENC/us02/n1035 ,\AES_ENC/us02/n1034 , \AES_ENC/us02/n1033 , \AES_ENC/us02/n1032 ,\AES_ENC/us02/n1031 , \AES_ENC/us02/n1030 , \AES_ENC/us02/n1029 ,\AES_ENC/us02/n1028 , \AES_ENC/us02/n1027 , \AES_ENC/us02/n1026 ,\AES_ENC/us02/n1025 , \AES_ENC/us02/n1024 , \AES_ENC/us02/n1023 ,\AES_ENC/us02/n1022 , \AES_ENC/us02/n1021 , \AES_ENC/us02/n1020 ,\AES_ENC/us02/n1019 , \AES_ENC/us02/n1018 , \AES_ENC/us02/n1017 ,\AES_ENC/us02/n1016 , \AES_ENC/us02/n1015 , \AES_ENC/us02/n1014 ,\AES_ENC/us02/n1013 , \AES_ENC/us02/n1012 , \AES_ENC/us02/n1011 ,\AES_ENC/us02/n1010 , \AES_ENC/us02/n1009 , \AES_ENC/us02/n1008 ,\AES_ENC/us02/n1007 , \AES_ENC/us02/n1006 , \AES_ENC/us02/n1005 ,\AES_ENC/us02/n1004 , \AES_ENC/us02/n1003 , \AES_ENC/us02/n1002 ,\AES_ENC/us02/n1001 , \AES_ENC/us02/n1000 , \AES_ENC/us02/n999 ,\AES_ENC/us02/n998 , \AES_ENC/us02/n997 , \AES_ENC/us02/n996 ,\AES_ENC/us02/n995 , \AES_ENC/us02/n994 , \AES_ENC/us02/n993 ,\AES_ENC/us02/n992 , \AES_ENC/us02/n991 , \AES_ENC/us02/n990 ,\AES_ENC/us02/n989 , \AES_ENC/us02/n988 , \AES_ENC/us02/n987 ,\AES_ENC/us02/n986 , \AES_ENC/us02/n985 , \AES_ENC/us02/n984 ,\AES_ENC/us02/n983 , \AES_ENC/us02/n982 , \AES_ENC/us02/n981 ,\AES_ENC/us02/n980 , \AES_ENC/us02/n979 , \AES_ENC/us02/n978 ,\AES_ENC/us02/n977 , \AES_ENC/us02/n976 , \AES_ENC/us02/n975 ,\AES_ENC/us02/n974 , \AES_ENC/us02/n973 , \AES_ENC/us02/n972 ,\AES_ENC/us02/n971 , \AES_ENC/us02/n970 , \AES_ENC/us02/n969 ,\AES_ENC/us02/n968 , \AES_ENC/us02/n967 , \AES_ENC/us02/n966 ,\AES_ENC/us02/n965 , \AES_ENC/us02/n964 , \AES_ENC/us02/n963 ,\AES_ENC/us02/n962 , \AES_ENC/us02/n961 , \AES_ENC/us02/n960 ,\AES_ENC/us02/n959 , \AES_ENC/us02/n958 , \AES_ENC/us02/n957 ,\AES_ENC/us02/n956 , \AES_ENC/us02/n955 , \AES_ENC/us02/n954 ,\AES_ENC/us02/n953 , \AES_ENC/us02/n952 , \AES_ENC/us02/n951 ,\AES_ENC/us02/n950 , \AES_ENC/us02/n949 , \AES_ENC/us02/n948 ,\AES_ENC/us02/n947 , \AES_ENC/us02/n946 , \AES_ENC/us02/n945 ,\AES_ENC/us02/n944 , \AES_ENC/us02/n943 , \AES_ENC/us02/n942 ,\AES_ENC/us02/n941 , \AES_ENC/us02/n940 , \AES_ENC/us02/n939 ,\AES_ENC/us02/n938 , \AES_ENC/us02/n937 , \AES_ENC/us02/n936 ,\AES_ENC/us02/n935 , \AES_ENC/us02/n934 , \AES_ENC/us02/n933 ,\AES_ENC/us02/n932 , \AES_ENC/us02/n931 , \AES_ENC/us02/n930 ,\AES_ENC/us02/n929 , \AES_ENC/us02/n928 , \AES_ENC/us02/n927 ,\AES_ENC/us02/n926 , \AES_ENC/us02/n925 , \AES_ENC/us02/n924 ,\AES_ENC/us02/n923 , \AES_ENC/us02/n922 , \AES_ENC/us02/n921 ,\AES_ENC/us02/n920 , \AES_ENC/us02/n919 , \AES_ENC/us02/n918 ,\AES_ENC/us02/n917 , \AES_ENC/us02/n916 , \AES_ENC/us02/n915 ,\AES_ENC/us02/n914 , \AES_ENC/us02/n913 , \AES_ENC/us02/n912 ,\AES_ENC/us02/n911 , \AES_ENC/us02/n910 , \AES_ENC/us02/n909 ,\AES_ENC/us02/n908 , \AES_ENC/us02/n907 , \AES_ENC/us02/n906 ,\AES_ENC/us02/n905 , \AES_ENC/us02/n904 , \AES_ENC/us02/n903 ,\AES_ENC/us02/n902 , \AES_ENC/us02/n901 , \AES_ENC/us02/n900 ,\AES_ENC/us02/n899 , \AES_ENC/us02/n898 , \AES_ENC/us02/n897 ,\AES_ENC/us02/n896 , \AES_ENC/us02/n895 , \AES_ENC/us02/n894 ,\AES_ENC/us02/n893 , \AES_ENC/us02/n892 , \AES_ENC/us02/n891 ,\AES_ENC/us02/n890 , \AES_ENC/us02/n889 , \AES_ENC/us02/n888 ,\AES_ENC/us02/n887 , \AES_ENC/us02/n886 , \AES_ENC/us02/n885 ,\AES_ENC/us02/n884 , \AES_ENC/us02/n883 , \AES_ENC/us02/n882 ,\AES_ENC/us02/n881 , \AES_ENC/us02/n880 , \AES_ENC/us02/n879 ,\AES_ENC/us02/n878 , \AES_ENC/us02/n877 , \AES_ENC/us02/n876 ,\AES_ENC/us02/n875 , \AES_ENC/us02/n874 , \AES_ENC/us02/n873 ,\AES_ENC/us02/n872 , \AES_ENC/us02/n871 , \AES_ENC/us02/n870 ,\AES_ENC/us02/n869 , \AES_ENC/us02/n868 , \AES_ENC/us02/n867 ,\AES_ENC/us02/n866 , \AES_ENC/us02/n865 , \AES_ENC/us02/n864 ,\AES_ENC/us02/n863 , \AES_ENC/us02/n862 , \AES_ENC/us02/n861 ,\AES_ENC/us02/n860 , \AES_ENC/us02/n859 , \AES_ENC/us02/n858 ,\AES_ENC/us02/n857 , \AES_ENC/us02/n856 , \AES_ENC/us02/n855 ,\AES_ENC/us02/n854 , \AES_ENC/us02/n853 , \AES_ENC/us02/n852 ,\AES_ENC/us02/n851 , \AES_ENC/us02/n850 , \AES_ENC/us02/n849 ,\AES_ENC/us02/n848 , \AES_ENC/us02/n847 , \AES_ENC/us02/n846 ,\AES_ENC/us02/n845 , \AES_ENC/us02/n844 , \AES_ENC/us02/n843 ,\AES_ENC/us02/n842 , \AES_ENC/us02/n841 , \AES_ENC/us02/n840 ,\AES_ENC/us02/n839 , \AES_ENC/us02/n838 , \AES_ENC/us02/n837 ,\AES_ENC/us02/n836 , \AES_ENC/us02/n835 , \AES_ENC/us02/n834 ,\AES_ENC/us02/n833 , \AES_ENC/us02/n832 , \AES_ENC/us02/n831 ,\AES_ENC/us02/n830 , \AES_ENC/us02/n829 , \AES_ENC/us02/n828 ,\AES_ENC/us02/n827 , \AES_ENC/us02/n826 , \AES_ENC/us02/n825 ,\AES_ENC/us02/n824 , \AES_ENC/us02/n823 , \AES_ENC/us02/n822 ,\AES_ENC/us02/n821 , \AES_ENC/us02/n820 , \AES_ENC/us02/n819 ,\AES_ENC/us02/n818 , \AES_ENC/us02/n817 , \AES_ENC/us02/n816 ,\AES_ENC/us02/n815 , \AES_ENC/us02/n814 , \AES_ENC/us02/n813 ,\AES_ENC/us02/n812 , \AES_ENC/us02/n811 , \AES_ENC/us02/n810 ,\AES_ENC/us02/n809 , \AES_ENC/us02/n808 , \AES_ENC/us02/n807 ,\AES_ENC/us02/n806 , \AES_ENC/us02/n805 , \AES_ENC/us02/n804 ,\AES_ENC/us02/n803 , \AES_ENC/us02/n802 , \AES_ENC/us02/n801 ,\AES_ENC/us02/n800 , \AES_ENC/us02/n799 , \AES_ENC/us02/n798 ,\AES_ENC/us02/n797 , \AES_ENC/us02/n796 , \AES_ENC/us02/n795 ,\AES_ENC/us02/n794 , \AES_ENC/us02/n793 , \AES_ENC/us02/n792 ,\AES_ENC/us02/n791 , \AES_ENC/us02/n790 , \AES_ENC/us02/n789 ,\AES_ENC/us02/n788 , \AES_ENC/us02/n787 , \AES_ENC/us02/n786 ,\AES_ENC/us02/n785 , \AES_ENC/us02/n784 , \AES_ENC/us02/n783 ,\AES_ENC/us02/n782 , \AES_ENC/us02/n781 , \AES_ENC/us02/n780 ,\AES_ENC/us02/n779 , \AES_ENC/us02/n778 , \AES_ENC/us02/n777 ,\AES_ENC/us02/n776 , \AES_ENC/us02/n775 , \AES_ENC/us02/n774 ,\AES_ENC/us02/n773 , \AES_ENC/us02/n772 , \AES_ENC/us02/n771 ,\AES_ENC/us02/n770 , \AES_ENC/us02/n769 , \AES_ENC/us02/n768 ,\AES_ENC/us02/n767 , \AES_ENC/us02/n766 , \AES_ENC/us02/n765 ,\AES_ENC/us02/n764 , \AES_ENC/us02/n763 , \AES_ENC/us02/n762 ,\AES_ENC/us02/n761 , \AES_ENC/us02/n760 , \AES_ENC/us02/n759 ,\AES_ENC/us02/n758 , \AES_ENC/us02/n757 , \AES_ENC/us02/n756 ,\AES_ENC/us02/n755 , \AES_ENC/us02/n754 , \AES_ENC/us02/n753 ,\AES_ENC/us02/n752 , \AES_ENC/us02/n751 , \AES_ENC/us02/n750 ,\AES_ENC/us02/n749 , \AES_ENC/us02/n748 , \AES_ENC/us02/n747 ,\AES_ENC/us02/n746 , \AES_ENC/us02/n745 , \AES_ENC/us02/n744 ,\AES_ENC/us02/n743 , \AES_ENC/us02/n742 , \AES_ENC/us02/n741 ,\AES_ENC/us02/n740 , \AES_ENC/us02/n739 , \AES_ENC/us02/n738 ,\AES_ENC/us02/n737 , \AES_ENC/us02/n736 , \AES_ENC/us02/n735 ,\AES_ENC/us02/n734 , \AES_ENC/us02/n733 , \AES_ENC/us02/n732 ,\AES_ENC/us02/n731 , \AES_ENC/us02/n730 , \AES_ENC/us02/n729 ,\AES_ENC/us02/n728 , \AES_ENC/us02/n727 , \AES_ENC/us02/n726 ,\AES_ENC/us02/n725 , \AES_ENC/us02/n724 , \AES_ENC/us02/n723 ,\AES_ENC/us02/n722 , \AES_ENC/us02/n721 , \AES_ENC/us02/n720 ,\AES_ENC/us02/n719 , \AES_ENC/us02/n718 , \AES_ENC/us02/n717 ,\AES_ENC/us02/n716 , \AES_ENC/us02/n715 , \AES_ENC/us02/n714 ,\AES_ENC/us02/n713 , \AES_ENC/us02/n712 , \AES_ENC/us02/n711 ,\AES_ENC/us02/n710 , \AES_ENC/us02/n709 , \AES_ENC/us02/n708 ,\AES_ENC/us02/n707 , \AES_ENC/us02/n706 , \AES_ENC/us02/n705 ,\AES_ENC/us02/n704 , \AES_ENC/us02/n703 , \AES_ENC/us02/n702 ,\AES_ENC/us02/n701 , \AES_ENC/us02/n700 , \AES_ENC/us02/n699 ,\AES_ENC/us02/n698 , \AES_ENC/us02/n697 , \AES_ENC/us02/n696 ,\AES_ENC/us02/n695 , \AES_ENC/us02/n694 , \AES_ENC/us02/n693 ,\AES_ENC/us02/n692 , \AES_ENC/us02/n691 , \AES_ENC/us02/n690 ,\AES_ENC/us02/n689 , \AES_ENC/us02/n688 , \AES_ENC/us02/n687 ,\AES_ENC/us02/n686 , \AES_ENC/us02/n685 , \AES_ENC/us02/n684 ,\AES_ENC/us02/n683 , \AES_ENC/us02/n682 , \AES_ENC/us02/n681 ,\AES_ENC/us02/n680 , \AES_ENC/us02/n679 , \AES_ENC/us02/n678 ,\AES_ENC/us02/n677 , \AES_ENC/us02/n676 , \AES_ENC/us02/n675 ,\AES_ENC/us02/n674 , \AES_ENC/us02/n673 , \AES_ENC/us02/n672 ,\AES_ENC/us02/n671 , \AES_ENC/us02/n670 , \AES_ENC/us02/n669 ,\AES_ENC/us02/n668 , \AES_ENC/us02/n667 , \AES_ENC/us02/n666 ,\AES_ENC/us02/n665 , \AES_ENC/us02/n664 , \AES_ENC/us02/n663 ,\AES_ENC/us02/n662 , \AES_ENC/us02/n661 , \AES_ENC/us02/n660 ,\AES_ENC/us02/n659 , \AES_ENC/us02/n658 , \AES_ENC/us02/n657 ,\AES_ENC/us02/n656 , \AES_ENC/us02/n655 , \AES_ENC/us02/n654 ,\AES_ENC/us02/n653 , \AES_ENC/us02/n652 , \AES_ENC/us02/n651 ,\AES_ENC/us02/n650 , \AES_ENC/us02/n649 , \AES_ENC/us02/n648 ,\AES_ENC/us02/n647 , \AES_ENC/us02/n646 , \AES_ENC/us02/n645 ,\AES_ENC/us02/n644 , \AES_ENC/us02/n643 , \AES_ENC/us02/n642 ,\AES_ENC/us02/n641 , \AES_ENC/us02/n640 , \AES_ENC/us02/n639 ,\AES_ENC/us02/n638 , \AES_ENC/us02/n637 , \AES_ENC/us02/n636 ,\AES_ENC/us02/n635 , \AES_ENC/us02/n634 , \AES_ENC/us02/n633 ,\AES_ENC/us02/n632 , \AES_ENC/us02/n631 , \AES_ENC/us02/n630 ,\AES_ENC/us02/n629 , \AES_ENC/us02/n628 , \AES_ENC/us02/n627 ,\AES_ENC/us02/n626 , \AES_ENC/us02/n625 , \AES_ENC/us02/n624 ,\AES_ENC/us02/n623 , \AES_ENC/us02/n622 , \AES_ENC/us02/n621 ,\AES_ENC/us02/n620 , \AES_ENC/us02/n619 , \AES_ENC/us02/n618 ,\AES_ENC/us02/n617 , \AES_ENC/us02/n616 , \AES_ENC/us02/n615 ,\AES_ENC/us02/n614 , \AES_ENC/us02/n613 , \AES_ENC/us02/n612 ,\AES_ENC/us02/n611 , \AES_ENC/us02/n610 , \AES_ENC/us02/n609 ,\AES_ENC/us02/n608 , \AES_ENC/us02/n607 , \AES_ENC/us02/n606 ,\AES_ENC/us02/n605 , \AES_ENC/us02/n604 , \AES_ENC/us02/n603 ,\AES_ENC/us02/n602 , \AES_ENC/us02/n601 , \AES_ENC/us02/n600 ,\AES_ENC/us02/n599 , \AES_ENC/us02/n598 , \AES_ENC/us02/n597 ,\AES_ENC/us02/n596 , \AES_ENC/us02/n595 , \AES_ENC/us02/n594 ,\AES_ENC/us02/n593 , \AES_ENC/us02/n592 , \AES_ENC/us02/n591 ,\AES_ENC/us02/n590 , \AES_ENC/us02/n589 , \AES_ENC/us02/n588 ,\AES_ENC/us02/n587 , \AES_ENC/us02/n586 , \AES_ENC/us02/n585 ,\AES_ENC/us02/n584 , \AES_ENC/us02/n583 , \AES_ENC/us02/n582 ,\AES_ENC/us02/n581 , \AES_ENC/us02/n580 , \AES_ENC/us02/n579 ,\AES_ENC/us02/n578 , \AES_ENC/us02/n577 , \AES_ENC/us02/n576 ,\AES_ENC/us02/n575 , \AES_ENC/us02/n574 , \AES_ENC/us02/n573 ,\AES_ENC/us02/n572 , \AES_ENC/us02/n571 , \AES_ENC/us02/n570 ,\AES_ENC/us02/n569 , \AES_ENC/us03/n1135 , \AES_ENC/us03/n1134 ,\AES_ENC/us03/n1133 , \AES_ENC/us03/n1132 , \AES_ENC/us03/n1131 ,\AES_ENC/us03/n1130 , \AES_ENC/us03/n1129 , \AES_ENC/us03/n1128 ,\AES_ENC/us03/n1127 , \AES_ENC/us03/n1126 , \AES_ENC/us03/n1125 ,\AES_ENC/us03/n1124 , \AES_ENC/us03/n1123 , \AES_ENC/us03/n1122 ,\AES_ENC/us03/n1121 , \AES_ENC/us03/n1120 , \AES_ENC/us03/n1119 ,\AES_ENC/us03/n1118 , \AES_ENC/us03/n1117 , \AES_ENC/us03/n1116 ,\AES_ENC/us03/n1115 , \AES_ENC/us03/n1114 , \AES_ENC/us03/n1113 ,\AES_ENC/us03/n1112 , \AES_ENC/us03/n1111 , \AES_ENC/us03/n1110 ,\AES_ENC/us03/n1109 , \AES_ENC/us03/n1108 , \AES_ENC/us03/n1107 ,\AES_ENC/us03/n1106 , \AES_ENC/us03/n1105 , \AES_ENC/us03/n1104 ,\AES_ENC/us03/n1103 , \AES_ENC/us03/n1102 , \AES_ENC/us03/n1101 ,\AES_ENC/us03/n1100 , \AES_ENC/us03/n1099 , \AES_ENC/us03/n1098 ,\AES_ENC/us03/n1097 , \AES_ENC/us03/n1096 , \AES_ENC/us03/n1095 ,\AES_ENC/us03/n1094 , \AES_ENC/us03/n1093 , \AES_ENC/us03/n1092 ,\AES_ENC/us03/n1091 , \AES_ENC/us03/n1090 , \AES_ENC/us03/n1089 ,\AES_ENC/us03/n1088 , \AES_ENC/us03/n1087 , \AES_ENC/us03/n1086 ,\AES_ENC/us03/n1085 , \AES_ENC/us03/n1084 , \AES_ENC/us03/n1083 ,\AES_ENC/us03/n1082 , \AES_ENC/us03/n1081 , \AES_ENC/us03/n1080 ,\AES_ENC/us03/n1079 , \AES_ENC/us03/n1078 , \AES_ENC/us03/n1077 ,\AES_ENC/us03/n1076 , \AES_ENC/us03/n1075 , \AES_ENC/us03/n1074 ,\AES_ENC/us03/n1073 , \AES_ENC/us03/n1072 , \AES_ENC/us03/n1071 ,\AES_ENC/us03/n1070 , \AES_ENC/us03/n1069 , \AES_ENC/us03/n1068 ,\AES_ENC/us03/n1067 , \AES_ENC/us03/n1066 , \AES_ENC/us03/n1065 ,\AES_ENC/us03/n1064 , \AES_ENC/us03/n1063 , \AES_ENC/us03/n1062 ,\AES_ENC/us03/n1061 , \AES_ENC/us03/n1060 , \AES_ENC/us03/n1059 ,\AES_ENC/us03/n1058 , \AES_ENC/us03/n1057 , \AES_ENC/us03/n1056 ,\AES_ENC/us03/n1055 , \AES_ENC/us03/n1054 , \AES_ENC/us03/n1053 ,\AES_ENC/us03/n1052 , \AES_ENC/us03/n1051 , \AES_ENC/us03/n1050 ,\AES_ENC/us03/n1049 , \AES_ENC/us03/n1048 , \AES_ENC/us03/n1047 ,\AES_ENC/us03/n1046 , \AES_ENC/us03/n1045 , \AES_ENC/us03/n1044 ,\AES_ENC/us03/n1043 , \AES_ENC/us03/n1042 , \AES_ENC/us03/n1041 ,\AES_ENC/us03/n1040 , \AES_ENC/us03/n1039 , \AES_ENC/us03/n1038 ,\AES_ENC/us03/n1037 , \AES_ENC/us03/n1036 , \AES_ENC/us03/n1035 ,\AES_ENC/us03/n1034 , \AES_ENC/us03/n1033 , \AES_ENC/us03/n1032 ,\AES_ENC/us03/n1031 , \AES_ENC/us03/n1030 , \AES_ENC/us03/n1029 ,\AES_ENC/us03/n1028 , \AES_ENC/us03/n1027 , \AES_ENC/us03/n1026 ,\AES_ENC/us03/n1025 , \AES_ENC/us03/n1024 , \AES_ENC/us03/n1023 ,\AES_ENC/us03/n1022 , \AES_ENC/us03/n1021 , \AES_ENC/us03/n1020 ,\AES_ENC/us03/n1019 , \AES_ENC/us03/n1018 , \AES_ENC/us03/n1017 ,\AES_ENC/us03/n1016 , \AES_ENC/us03/n1015 , \AES_ENC/us03/n1014 ,\AES_ENC/us03/n1013 , \AES_ENC/us03/n1012 , \AES_ENC/us03/n1011 ,\AES_ENC/us03/n1010 , \AES_ENC/us03/n1009 , \AES_ENC/us03/n1008 ,\AES_ENC/us03/n1007 , \AES_ENC/us03/n1006 , \AES_ENC/us03/n1005 ,\AES_ENC/us03/n1004 , \AES_ENC/us03/n1003 , \AES_ENC/us03/n1002 ,\AES_ENC/us03/n1001 , \AES_ENC/us03/n1000 , \AES_ENC/us03/n999 ,\AES_ENC/us03/n998 , \AES_ENC/us03/n997 , \AES_ENC/us03/n996 ,\AES_ENC/us03/n995 , \AES_ENC/us03/n994 , \AES_ENC/us03/n993 ,\AES_ENC/us03/n992 , \AES_ENC/us03/n991 , \AES_ENC/us03/n990 ,\AES_ENC/us03/n989 , \AES_ENC/us03/n988 , \AES_ENC/us03/n987 ,\AES_ENC/us03/n986 , \AES_ENC/us03/n985 , \AES_ENC/us03/n984 ,\AES_ENC/us03/n983 , \AES_ENC/us03/n982 , \AES_ENC/us03/n981 ,\AES_ENC/us03/n980 , \AES_ENC/us03/n979 , \AES_ENC/us03/n978 ,\AES_ENC/us03/n977 , \AES_ENC/us03/n976 , \AES_ENC/us03/n975 ,\AES_ENC/us03/n974 , \AES_ENC/us03/n973 , \AES_ENC/us03/n972 ,\AES_ENC/us03/n971 , \AES_ENC/us03/n970 , \AES_ENC/us03/n969 ,\AES_ENC/us03/n968 , \AES_ENC/us03/n967 , \AES_ENC/us03/n966 ,\AES_ENC/us03/n965 , \AES_ENC/us03/n964 , \AES_ENC/us03/n963 ,\AES_ENC/us03/n962 , \AES_ENC/us03/n961 , \AES_ENC/us03/n960 ,\AES_ENC/us03/n959 , \AES_ENC/us03/n958 , \AES_ENC/us03/n957 ,\AES_ENC/us03/n956 , \AES_ENC/us03/n955 , \AES_ENC/us03/n954 ,\AES_ENC/us03/n953 , \AES_ENC/us03/n952 , \AES_ENC/us03/n951 ,\AES_ENC/us03/n950 , \AES_ENC/us03/n949 , \AES_ENC/us03/n948 ,\AES_ENC/us03/n947 , \AES_ENC/us03/n946 , \AES_ENC/us03/n945 ,\AES_ENC/us03/n944 , \AES_ENC/us03/n943 , \AES_ENC/us03/n942 ,\AES_ENC/us03/n941 , \AES_ENC/us03/n940 , \AES_ENC/us03/n939 ,\AES_ENC/us03/n938 , \AES_ENC/us03/n937 , \AES_ENC/us03/n936 ,\AES_ENC/us03/n935 , \AES_ENC/us03/n934 , \AES_ENC/us03/n933 ,\AES_ENC/us03/n932 , \AES_ENC/us03/n931 , \AES_ENC/us03/n930 ,\AES_ENC/us03/n929 , \AES_ENC/us03/n928 , \AES_ENC/us03/n927 ,\AES_ENC/us03/n926 , \AES_ENC/us03/n925 , \AES_ENC/us03/n924 ,\AES_ENC/us03/n923 , \AES_ENC/us03/n922 , \AES_ENC/us03/n921 ,\AES_ENC/us03/n920 , \AES_ENC/us03/n919 , \AES_ENC/us03/n918 ,\AES_ENC/us03/n917 , \AES_ENC/us03/n916 , \AES_ENC/us03/n915 ,\AES_ENC/us03/n914 , \AES_ENC/us03/n913 , \AES_ENC/us03/n912 ,\AES_ENC/us03/n911 , \AES_ENC/us03/n910 , \AES_ENC/us03/n909 ,\AES_ENC/us03/n908 , \AES_ENC/us03/n907 , \AES_ENC/us03/n906 ,\AES_ENC/us03/n905 , \AES_ENC/us03/n904 , \AES_ENC/us03/n903 ,\AES_ENC/us03/n902 , \AES_ENC/us03/n901 , \AES_ENC/us03/n900 ,\AES_ENC/us03/n899 , \AES_ENC/us03/n898 , \AES_ENC/us03/n897 ,\AES_ENC/us03/n896 , \AES_ENC/us03/n895 , \AES_ENC/us03/n894 ,\AES_ENC/us03/n893 , \AES_ENC/us03/n892 , \AES_ENC/us03/n891 ,\AES_ENC/us03/n890 , \AES_ENC/us03/n889 , \AES_ENC/us03/n888 ,\AES_ENC/us03/n887 , \AES_ENC/us03/n886 , \AES_ENC/us03/n885 ,\AES_ENC/us03/n884 , \AES_ENC/us03/n883 , \AES_ENC/us03/n882 ,\AES_ENC/us03/n881 , \AES_ENC/us03/n880 , \AES_ENC/us03/n879 ,\AES_ENC/us03/n878 , \AES_ENC/us03/n877 , \AES_ENC/us03/n876 ,\AES_ENC/us03/n875 , \AES_ENC/us03/n874 , \AES_ENC/us03/n873 ,\AES_ENC/us03/n872 , \AES_ENC/us03/n871 , \AES_ENC/us03/n870 ,\AES_ENC/us03/n869 , \AES_ENC/us03/n868 , \AES_ENC/us03/n867 ,\AES_ENC/us03/n866 , \AES_ENC/us03/n865 , \AES_ENC/us03/n864 ,\AES_ENC/us03/n863 , \AES_ENC/us03/n862 , \AES_ENC/us03/n861 ,\AES_ENC/us03/n860 , \AES_ENC/us03/n859 , \AES_ENC/us03/n858 ,\AES_ENC/us03/n857 , \AES_ENC/us03/n856 , \AES_ENC/us03/n855 ,\AES_ENC/us03/n854 , \AES_ENC/us03/n853 , \AES_ENC/us03/n852 ,\AES_ENC/us03/n851 , \AES_ENC/us03/n850 , \AES_ENC/us03/n849 ,\AES_ENC/us03/n848 , \AES_ENC/us03/n847 , \AES_ENC/us03/n846 ,\AES_ENC/us03/n845 , \AES_ENC/us03/n844 , \AES_ENC/us03/n843 ,\AES_ENC/us03/n842 , \AES_ENC/us03/n841 , \AES_ENC/us03/n840 ,\AES_ENC/us03/n839 , \AES_ENC/us03/n838 , \AES_ENC/us03/n837 ,\AES_ENC/us03/n836 , \AES_ENC/us03/n835 , \AES_ENC/us03/n834 ,\AES_ENC/us03/n833 , \AES_ENC/us03/n832 , \AES_ENC/us03/n831 ,\AES_ENC/us03/n830 , \AES_ENC/us03/n829 , \AES_ENC/us03/n828 ,\AES_ENC/us03/n827 , \AES_ENC/us03/n826 , \AES_ENC/us03/n825 ,\AES_ENC/us03/n824 , \AES_ENC/us03/n823 , \AES_ENC/us03/n822 ,\AES_ENC/us03/n821 , \AES_ENC/us03/n820 , \AES_ENC/us03/n819 ,\AES_ENC/us03/n818 , \AES_ENC/us03/n817 , \AES_ENC/us03/n816 ,\AES_ENC/us03/n815 , \AES_ENC/us03/n814 , \AES_ENC/us03/n813 ,\AES_ENC/us03/n812 , \AES_ENC/us03/n811 , \AES_ENC/us03/n810 ,\AES_ENC/us03/n809 , \AES_ENC/us03/n808 , \AES_ENC/us03/n807 ,\AES_ENC/us03/n806 , \AES_ENC/us03/n805 , \AES_ENC/us03/n804 ,\AES_ENC/us03/n803 , \AES_ENC/us03/n802 , \AES_ENC/us03/n801 ,\AES_ENC/us03/n800 , \AES_ENC/us03/n799 , \AES_ENC/us03/n798 ,\AES_ENC/us03/n797 , \AES_ENC/us03/n796 , \AES_ENC/us03/n795 ,\AES_ENC/us03/n794 , \AES_ENC/us03/n793 , \AES_ENC/us03/n792 ,\AES_ENC/us03/n791 , \AES_ENC/us03/n790 , \AES_ENC/us03/n789 ,\AES_ENC/us03/n788 , \AES_ENC/us03/n787 , \AES_ENC/us03/n786 ,\AES_ENC/us03/n785 , \AES_ENC/us03/n784 , \AES_ENC/us03/n783 ,\AES_ENC/us03/n782 , \AES_ENC/us03/n781 , \AES_ENC/us03/n780 ,\AES_ENC/us03/n779 , \AES_ENC/us03/n778 , \AES_ENC/us03/n777 ,\AES_ENC/us03/n776 , \AES_ENC/us03/n775 , \AES_ENC/us03/n774 ,\AES_ENC/us03/n773 , \AES_ENC/us03/n772 , \AES_ENC/us03/n771 ,\AES_ENC/us03/n770 , \AES_ENC/us03/n769 , \AES_ENC/us03/n768 ,\AES_ENC/us03/n767 , \AES_ENC/us03/n766 , \AES_ENC/us03/n765 ,\AES_ENC/us03/n764 , \AES_ENC/us03/n763 , \AES_ENC/us03/n762 ,\AES_ENC/us03/n761 , \AES_ENC/us03/n760 , \AES_ENC/us03/n759 ,\AES_ENC/us03/n758 , \AES_ENC/us03/n757 , \AES_ENC/us03/n756 ,\AES_ENC/us03/n755 , \AES_ENC/us03/n754 , \AES_ENC/us03/n753 ,\AES_ENC/us03/n752 , \AES_ENC/us03/n751 , \AES_ENC/us03/n750 ,\AES_ENC/us03/n749 , \AES_ENC/us03/n748 , \AES_ENC/us03/n747 ,\AES_ENC/us03/n746 , \AES_ENC/us03/n745 , \AES_ENC/us03/n744 ,\AES_ENC/us03/n743 , \AES_ENC/us03/n742 , \AES_ENC/us03/n741 ,\AES_ENC/us03/n740 , \AES_ENC/us03/n739 , \AES_ENC/us03/n738 ,\AES_ENC/us03/n737 , \AES_ENC/us03/n736 , \AES_ENC/us03/n735 ,\AES_ENC/us03/n734 , \AES_ENC/us03/n733 , \AES_ENC/us03/n732 ,\AES_ENC/us03/n731 , \AES_ENC/us03/n730 , \AES_ENC/us03/n729 ,\AES_ENC/us03/n728 , \AES_ENC/us03/n727 , \AES_ENC/us03/n726 ,\AES_ENC/us03/n725 , \AES_ENC/us03/n724 , \AES_ENC/us03/n723 ,\AES_ENC/us03/n722 , \AES_ENC/us03/n721 , \AES_ENC/us03/n720 ,\AES_ENC/us03/n719 , \AES_ENC/us03/n718 , \AES_ENC/us03/n717 ,\AES_ENC/us03/n716 , \AES_ENC/us03/n715 , \AES_ENC/us03/n714 ,\AES_ENC/us03/n713 , \AES_ENC/us03/n712 , \AES_ENC/us03/n711 ,\AES_ENC/us03/n710 , \AES_ENC/us03/n709 , \AES_ENC/us03/n708 ,\AES_ENC/us03/n707 , \AES_ENC/us03/n706 , \AES_ENC/us03/n705 ,\AES_ENC/us03/n704 , \AES_ENC/us03/n703 , \AES_ENC/us03/n702 ,\AES_ENC/us03/n701 , \AES_ENC/us03/n700 , \AES_ENC/us03/n699 ,\AES_ENC/us03/n698 , \AES_ENC/us03/n697 , \AES_ENC/us03/n696 ,\AES_ENC/us03/n695 , \AES_ENC/us03/n694 , \AES_ENC/us03/n693 ,\AES_ENC/us03/n692 , \AES_ENC/us03/n691 , \AES_ENC/us03/n690 ,\AES_ENC/us03/n689 , \AES_ENC/us03/n688 , \AES_ENC/us03/n687 ,\AES_ENC/us03/n686 , \AES_ENC/us03/n685 , \AES_ENC/us03/n684 ,\AES_ENC/us03/n683 , \AES_ENC/us03/n682 , \AES_ENC/us03/n681 ,\AES_ENC/us03/n680 , \AES_ENC/us03/n679 , \AES_ENC/us03/n678 ,\AES_ENC/us03/n677 , \AES_ENC/us03/n676 , \AES_ENC/us03/n675 ,\AES_ENC/us03/n674 , \AES_ENC/us03/n673 , \AES_ENC/us03/n672 ,\AES_ENC/us03/n671 , \AES_ENC/us03/n670 , \AES_ENC/us03/n669 ,\AES_ENC/us03/n668 , \AES_ENC/us03/n667 , \AES_ENC/us03/n666 ,\AES_ENC/us03/n665 , \AES_ENC/us03/n664 , \AES_ENC/us03/n663 ,\AES_ENC/us03/n662 , \AES_ENC/us03/n661 , \AES_ENC/us03/n660 ,\AES_ENC/us03/n659 , \AES_ENC/us03/n658 , \AES_ENC/us03/n657 ,\AES_ENC/us03/n656 , \AES_ENC/us03/n655 , \AES_ENC/us03/n654 ,\AES_ENC/us03/n653 , \AES_ENC/us03/n652 , \AES_ENC/us03/n651 ,\AES_ENC/us03/n650 , \AES_ENC/us03/n649 , \AES_ENC/us03/n648 ,\AES_ENC/us03/n647 , \AES_ENC/us03/n646 , \AES_ENC/us03/n645 ,\AES_ENC/us03/n644 , \AES_ENC/us03/n643 , \AES_ENC/us03/n642 ,\AES_ENC/us03/n641 , \AES_ENC/us03/n640 , \AES_ENC/us03/n639 ,\AES_ENC/us03/n638 , \AES_ENC/us03/n637 , \AES_ENC/us03/n636 ,\AES_ENC/us03/n635 , \AES_ENC/us03/n634 , \AES_ENC/us03/n633 ,\AES_ENC/us03/n632 , \AES_ENC/us03/n631 , \AES_ENC/us03/n630 ,\AES_ENC/us03/n629 , \AES_ENC/us03/n628 , \AES_ENC/us03/n627 ,\AES_ENC/us03/n626 , \AES_ENC/us03/n625 , \AES_ENC/us03/n624 ,\AES_ENC/us03/n623 , \AES_ENC/us03/n622 , \AES_ENC/us03/n621 ,\AES_ENC/us03/n620 , \AES_ENC/us03/n619 , \AES_ENC/us03/n618 ,\AES_ENC/us03/n617 , \AES_ENC/us03/n616 , \AES_ENC/us03/n615 ,\AES_ENC/us03/n614 , \AES_ENC/us03/n613 , \AES_ENC/us03/n612 ,\AES_ENC/us03/n611 , \AES_ENC/us03/n610 , \AES_ENC/us03/n609 ,\AES_ENC/us03/n608 , \AES_ENC/us03/n607 , \AES_ENC/us03/n606 ,\AES_ENC/us03/n605 , \AES_ENC/us03/n604 , \AES_ENC/us03/n603 ,\AES_ENC/us03/n602 , \AES_ENC/us03/n601 , \AES_ENC/us03/n600 ,\AES_ENC/us03/n599 , \AES_ENC/us03/n598 , \AES_ENC/us03/n597 ,\AES_ENC/us03/n596 , \AES_ENC/us03/n595 , \AES_ENC/us03/n594 ,\AES_ENC/us03/n593 , \AES_ENC/us03/n592 , \AES_ENC/us03/n591 ,\AES_ENC/us03/n590 , \AES_ENC/us03/n589 , \AES_ENC/us03/n588 ,\AES_ENC/us03/n587 , \AES_ENC/us03/n586 , \AES_ENC/us03/n585 ,\AES_ENC/us03/n584 , \AES_ENC/us03/n583 , \AES_ENC/us03/n582 ,\AES_ENC/us03/n581 , \AES_ENC/us03/n580 , \AES_ENC/us03/n579 ,\AES_ENC/us03/n578 , \AES_ENC/us03/n577 , \AES_ENC/us03/n576 ,\AES_ENC/us03/n575 , \AES_ENC/us03/n574 , \AES_ENC/us03/n573 ,\AES_ENC/us03/n572 , \AES_ENC/us03/n571 , \AES_ENC/us03/n570 ,\AES_ENC/us03/n569 , \AES_ENC/us10/n1135 , \AES_ENC/us10/n1134 ,\AES_ENC/us10/n1133 , \AES_ENC/us10/n1132 , \AES_ENC/us10/n1131 ,\AES_ENC/us10/n1130 , \AES_ENC/us10/n1129 , \AES_ENC/us10/n1128 ,\AES_ENC/us10/n1127 , \AES_ENC/us10/n1126 , \AES_ENC/us10/n1125 ,\AES_ENC/us10/n1124 , \AES_ENC/us10/n1123 , \AES_ENC/us10/n1122 ,\AES_ENC/us10/n1121 , \AES_ENC/us10/n1120 , \AES_ENC/us10/n1119 ,\AES_ENC/us10/n1118 , \AES_ENC/us10/n1117 , \AES_ENC/us10/n1116 ,\AES_ENC/us10/n1115 , \AES_ENC/us10/n1114 , \AES_ENC/us10/n1113 ,\AES_ENC/us10/n1112 , \AES_ENC/us10/n1111 , \AES_ENC/us10/n1110 ,\AES_ENC/us10/n1109 , \AES_ENC/us10/n1108 , \AES_ENC/us10/n1107 ,\AES_ENC/us10/n1106 , \AES_ENC/us10/n1105 , \AES_ENC/us10/n1104 ,\AES_ENC/us10/n1103 , \AES_ENC/us10/n1102 , \AES_ENC/us10/n1101 ,\AES_ENC/us10/n1100 , \AES_ENC/us10/n1099 , \AES_ENC/us10/n1098 ,\AES_ENC/us10/n1097 , \AES_ENC/us10/n1096 , \AES_ENC/us10/n1095 ,\AES_ENC/us10/n1094 , \AES_ENC/us10/n1093 , \AES_ENC/us10/n1092 ,\AES_ENC/us10/n1091 , \AES_ENC/us10/n1090 , \AES_ENC/us10/n1089 ,\AES_ENC/us10/n1088 , \AES_ENC/us10/n1087 , \AES_ENC/us10/n1086 ,\AES_ENC/us10/n1085 , \AES_ENC/us10/n1084 , \AES_ENC/us10/n1083 ,\AES_ENC/us10/n1082 , \AES_ENC/us10/n1081 , \AES_ENC/us10/n1080 ,\AES_ENC/us10/n1079 , \AES_ENC/us10/n1078 , \AES_ENC/us10/n1077 ,\AES_ENC/us10/n1076 , \AES_ENC/us10/n1075 , \AES_ENC/us10/n1074 ,\AES_ENC/us10/n1073 , \AES_ENC/us10/n1072 , \AES_ENC/us10/n1071 ,\AES_ENC/us10/n1070 , \AES_ENC/us10/n1069 , \AES_ENC/us10/n1068 ,\AES_ENC/us10/n1067 , \AES_ENC/us10/n1066 , \AES_ENC/us10/n1065 ,\AES_ENC/us10/n1064 , \AES_ENC/us10/n1063 , \AES_ENC/us10/n1062 ,\AES_ENC/us10/n1061 , \AES_ENC/us10/n1060 , \AES_ENC/us10/n1059 ,\AES_ENC/us10/n1058 , \AES_ENC/us10/n1057 , \AES_ENC/us10/n1056 ,\AES_ENC/us10/n1055 , \AES_ENC/us10/n1054 , \AES_ENC/us10/n1053 ,\AES_ENC/us10/n1052 , \AES_ENC/us10/n1051 , \AES_ENC/us10/n1050 ,\AES_ENC/us10/n1049 , \AES_ENC/us10/n1048 , \AES_ENC/us10/n1047 ,\AES_ENC/us10/n1046 , \AES_ENC/us10/n1045 , \AES_ENC/us10/n1044 ,\AES_ENC/us10/n1043 , \AES_ENC/us10/n1042 , \AES_ENC/us10/n1041 ,\AES_ENC/us10/n1040 , \AES_ENC/us10/n1039 , \AES_ENC/us10/n1038 ,\AES_ENC/us10/n1037 , \AES_ENC/us10/n1036 , \AES_ENC/us10/n1035 ,\AES_ENC/us10/n1034 , \AES_ENC/us10/n1033 , \AES_ENC/us10/n1032 ,\AES_ENC/us10/n1031 , \AES_ENC/us10/n1030 , \AES_ENC/us10/n1029 ,\AES_ENC/us10/n1028 , \AES_ENC/us10/n1027 , \AES_ENC/us10/n1026 ,\AES_ENC/us10/n1025 , \AES_ENC/us10/n1024 , \AES_ENC/us10/n1023 ,\AES_ENC/us10/n1022 , \AES_ENC/us10/n1021 , \AES_ENC/us10/n1020 ,\AES_ENC/us10/n1019 , \AES_ENC/us10/n1018 , \AES_ENC/us10/n1017 ,\AES_ENC/us10/n1016 , \AES_ENC/us10/n1015 , \AES_ENC/us10/n1014 ,\AES_ENC/us10/n1013 , \AES_ENC/us10/n1012 , \AES_ENC/us10/n1011 ,\AES_ENC/us10/n1010 , \AES_ENC/us10/n1009 , \AES_ENC/us10/n1008 ,\AES_ENC/us10/n1007 , \AES_ENC/us10/n1006 , \AES_ENC/us10/n1005 ,\AES_ENC/us10/n1004 , \AES_ENC/us10/n1003 , \AES_ENC/us10/n1002 ,\AES_ENC/us10/n1001 , \AES_ENC/us10/n1000 , \AES_ENC/us10/n999 ,\AES_ENC/us10/n998 , \AES_ENC/us10/n997 , \AES_ENC/us10/n996 ,\AES_ENC/us10/n995 , \AES_ENC/us10/n994 , \AES_ENC/us10/n993 ,\AES_ENC/us10/n992 , \AES_ENC/us10/n991 , \AES_ENC/us10/n990 ,\AES_ENC/us10/n989 , \AES_ENC/us10/n988 , \AES_ENC/us10/n987 ,\AES_ENC/us10/n986 , \AES_ENC/us10/n985 , \AES_ENC/us10/n984 ,\AES_ENC/us10/n983 , \AES_ENC/us10/n982 , \AES_ENC/us10/n981 ,\AES_ENC/us10/n980 , \AES_ENC/us10/n979 , \AES_ENC/us10/n978 ,\AES_ENC/us10/n977 , \AES_ENC/us10/n976 , \AES_ENC/us10/n975 ,\AES_ENC/us10/n974 , \AES_ENC/us10/n973 , \AES_ENC/us10/n972 ,\AES_ENC/us10/n971 , \AES_ENC/us10/n970 , \AES_ENC/us10/n969 ,\AES_ENC/us10/n968 , \AES_ENC/us10/n967 , \AES_ENC/us10/n966 ,\AES_ENC/us10/n965 , \AES_ENC/us10/n964 , \AES_ENC/us10/n963 ,\AES_ENC/us10/n962 , \AES_ENC/us10/n961 , \AES_ENC/us10/n960 ,\AES_ENC/us10/n959 , \AES_ENC/us10/n958 , \AES_ENC/us10/n957 ,\AES_ENC/us10/n956 , \AES_ENC/us10/n955 , \AES_ENC/us10/n954 ,\AES_ENC/us10/n953 , \AES_ENC/us10/n952 , \AES_ENC/us10/n951 ,\AES_ENC/us10/n950 , \AES_ENC/us10/n949 , \AES_ENC/us10/n948 ,\AES_ENC/us10/n947 , \AES_ENC/us10/n946 , \AES_ENC/us10/n945 ,\AES_ENC/us10/n944 , \AES_ENC/us10/n943 , \AES_ENC/us10/n942 ,\AES_ENC/us10/n941 , \AES_ENC/us10/n940 , \AES_ENC/us10/n939 ,\AES_ENC/us10/n938 , \AES_ENC/us10/n937 , \AES_ENC/us10/n936 ,\AES_ENC/us10/n935 , \AES_ENC/us10/n934 , \AES_ENC/us10/n933 ,\AES_ENC/us10/n932 , \AES_ENC/us10/n931 , \AES_ENC/us10/n930 ,\AES_ENC/us10/n929 , \AES_ENC/us10/n928 , \AES_ENC/us10/n927 ,\AES_ENC/us10/n926 , \AES_ENC/us10/n925 , \AES_ENC/us10/n924 ,\AES_ENC/us10/n923 , \AES_ENC/us10/n922 , \AES_ENC/us10/n921 ,\AES_ENC/us10/n920 , \AES_ENC/us10/n919 , \AES_ENC/us10/n918 ,\AES_ENC/us10/n917 , \AES_ENC/us10/n916 , \AES_ENC/us10/n915 ,\AES_ENC/us10/n914 , \AES_ENC/us10/n913 , \AES_ENC/us10/n912 ,\AES_ENC/us10/n911 , \AES_ENC/us10/n910 , \AES_ENC/us10/n909 ,\AES_ENC/us10/n908 , \AES_ENC/us10/n907 , \AES_ENC/us10/n906 ,\AES_ENC/us10/n905 , \AES_ENC/us10/n904 , \AES_ENC/us10/n903 ,\AES_ENC/us10/n902 , \AES_ENC/us10/n901 , \AES_ENC/us10/n900 ,\AES_ENC/us10/n899 , \AES_ENC/us10/n898 , \AES_ENC/us10/n897 ,\AES_ENC/us10/n896 , \AES_ENC/us10/n895 , \AES_ENC/us10/n894 ,\AES_ENC/us10/n893 , \AES_ENC/us10/n892 , \AES_ENC/us10/n891 ,\AES_ENC/us10/n890 , \AES_ENC/us10/n889 , \AES_ENC/us10/n888 ,\AES_ENC/us10/n887 , \AES_ENC/us10/n886 , \AES_ENC/us10/n885 ,\AES_ENC/us10/n884 , \AES_ENC/us10/n883 , \AES_ENC/us10/n882 ,\AES_ENC/us10/n881 , \AES_ENC/us10/n880 , \AES_ENC/us10/n879 ,\AES_ENC/us10/n878 , \AES_ENC/us10/n877 , \AES_ENC/us10/n876 ,\AES_ENC/us10/n875 , \AES_ENC/us10/n874 , \AES_ENC/us10/n873 ,\AES_ENC/us10/n872 , \AES_ENC/us10/n871 , \AES_ENC/us10/n870 ,\AES_ENC/us10/n869 , \AES_ENC/us10/n868 , \AES_ENC/us10/n867 ,\AES_ENC/us10/n866 , \AES_ENC/us10/n865 , \AES_ENC/us10/n864 ,\AES_ENC/us10/n863 , \AES_ENC/us10/n862 , \AES_ENC/us10/n861 ,\AES_ENC/us10/n860 , \AES_ENC/us10/n859 , \AES_ENC/us10/n858 ,\AES_ENC/us10/n857 , \AES_ENC/us10/n856 , \AES_ENC/us10/n855 ,\AES_ENC/us10/n854 , \AES_ENC/us10/n853 , \AES_ENC/us10/n852 ,\AES_ENC/us10/n851 , \AES_ENC/us10/n850 , \AES_ENC/us10/n849 ,\AES_ENC/us10/n848 , \AES_ENC/us10/n847 , \AES_ENC/us10/n846 ,\AES_ENC/us10/n845 , \AES_ENC/us10/n844 , \AES_ENC/us10/n843 ,\AES_ENC/us10/n842 , \AES_ENC/us10/n841 , \AES_ENC/us10/n840 ,\AES_ENC/us10/n839 , \AES_ENC/us10/n838 , \AES_ENC/us10/n837 ,\AES_ENC/us10/n836 , \AES_ENC/us10/n835 , \AES_ENC/us10/n834 ,\AES_ENC/us10/n833 , \AES_ENC/us10/n832 , \AES_ENC/us10/n831 ,\AES_ENC/us10/n830 , \AES_ENC/us10/n829 , \AES_ENC/us10/n828 ,\AES_ENC/us10/n827 , \AES_ENC/us10/n826 , \AES_ENC/us10/n825 ,\AES_ENC/us10/n824 , \AES_ENC/us10/n823 , \AES_ENC/us10/n822 ,\AES_ENC/us10/n821 , \AES_ENC/us10/n820 , \AES_ENC/us10/n819 ,\AES_ENC/us10/n818 , \AES_ENC/us10/n817 , \AES_ENC/us10/n816 ,\AES_ENC/us10/n815 , \AES_ENC/us10/n814 , \AES_ENC/us10/n813 ,\AES_ENC/us10/n812 , \AES_ENC/us10/n811 , \AES_ENC/us10/n810 ,\AES_ENC/us10/n809 , \AES_ENC/us10/n808 , \AES_ENC/us10/n807 ,\AES_ENC/us10/n806 , \AES_ENC/us10/n805 , \AES_ENC/us10/n804 ,\AES_ENC/us10/n803 , \AES_ENC/us10/n802 , \AES_ENC/us10/n801 ,\AES_ENC/us10/n800 , \AES_ENC/us10/n799 , \AES_ENC/us10/n798 ,\AES_ENC/us10/n797 , \AES_ENC/us10/n796 , \AES_ENC/us10/n795 ,\AES_ENC/us10/n794 , \AES_ENC/us10/n793 , \AES_ENC/us10/n792 ,\AES_ENC/us10/n791 , \AES_ENC/us10/n790 , \AES_ENC/us10/n789 ,\AES_ENC/us10/n788 , \AES_ENC/us10/n787 , \AES_ENC/us10/n786 ,\AES_ENC/us10/n785 , \AES_ENC/us10/n784 , \AES_ENC/us10/n783 ,\AES_ENC/us10/n782 , \AES_ENC/us10/n781 , \AES_ENC/us10/n780 ,\AES_ENC/us10/n779 , \AES_ENC/us10/n778 , \AES_ENC/us10/n777 ,\AES_ENC/us10/n776 , \AES_ENC/us10/n775 , \AES_ENC/us10/n774 ,\AES_ENC/us10/n773 , \AES_ENC/us10/n772 , \AES_ENC/us10/n771 ,\AES_ENC/us10/n770 , \AES_ENC/us10/n769 , \AES_ENC/us10/n768 ,\AES_ENC/us10/n767 , \AES_ENC/us10/n766 , \AES_ENC/us10/n765 ,\AES_ENC/us10/n764 , \AES_ENC/us10/n763 , \AES_ENC/us10/n762 ,\AES_ENC/us10/n761 , \AES_ENC/us10/n760 , \AES_ENC/us10/n759 ,\AES_ENC/us10/n758 , \AES_ENC/us10/n757 , \AES_ENC/us10/n756 ,\AES_ENC/us10/n755 , \AES_ENC/us10/n754 , \AES_ENC/us10/n753 ,\AES_ENC/us10/n752 , \AES_ENC/us10/n751 , \AES_ENC/us10/n750 ,\AES_ENC/us10/n749 , \AES_ENC/us10/n748 , \AES_ENC/us10/n747 ,\AES_ENC/us10/n746 , \AES_ENC/us10/n745 , \AES_ENC/us10/n744 ,\AES_ENC/us10/n743 , \AES_ENC/us10/n742 , \AES_ENC/us10/n741 ,\AES_ENC/us10/n740 , \AES_ENC/us10/n739 , \AES_ENC/us10/n738 ,\AES_ENC/us10/n737 , \AES_ENC/us10/n736 , \AES_ENC/us10/n735 ,\AES_ENC/us10/n734 , \AES_ENC/us10/n733 , \AES_ENC/us10/n732 ,\AES_ENC/us10/n731 , \AES_ENC/us10/n730 , \AES_ENC/us10/n729 ,\AES_ENC/us10/n728 , \AES_ENC/us10/n727 , \AES_ENC/us10/n726 ,\AES_ENC/us10/n725 , \AES_ENC/us10/n724 , \AES_ENC/us10/n723 ,\AES_ENC/us10/n722 , \AES_ENC/us10/n721 , \AES_ENC/us10/n720 ,\AES_ENC/us10/n719 , \AES_ENC/us10/n718 , \AES_ENC/us10/n717 ,\AES_ENC/us10/n716 , \AES_ENC/us10/n715 , \AES_ENC/us10/n714 ,\AES_ENC/us10/n713 , \AES_ENC/us10/n712 , \AES_ENC/us10/n711 ,\AES_ENC/us10/n710 , \AES_ENC/us10/n709 , \AES_ENC/us10/n708 ,\AES_ENC/us10/n707 , \AES_ENC/us10/n706 , \AES_ENC/us10/n705 ,\AES_ENC/us10/n704 , \AES_ENC/us10/n703 , \AES_ENC/us10/n702 ,\AES_ENC/us10/n701 , \AES_ENC/us10/n700 , \AES_ENC/us10/n699 ,\AES_ENC/us10/n698 , \AES_ENC/us10/n697 , \AES_ENC/us10/n696 ,\AES_ENC/us10/n695 , \AES_ENC/us10/n694 , \AES_ENC/us10/n693 ,\AES_ENC/us10/n692 , \AES_ENC/us10/n691 , \AES_ENC/us10/n690 ,\AES_ENC/us10/n689 , \AES_ENC/us10/n688 , \AES_ENC/us10/n687 ,\AES_ENC/us10/n686 , \AES_ENC/us10/n685 , \AES_ENC/us10/n684 ,\AES_ENC/us10/n683 , \AES_ENC/us10/n682 , \AES_ENC/us10/n681 ,\AES_ENC/us10/n680 , \AES_ENC/us10/n679 , \AES_ENC/us10/n678 ,\AES_ENC/us10/n677 , \AES_ENC/us10/n676 , \AES_ENC/us10/n675 ,\AES_ENC/us10/n674 , \AES_ENC/us10/n673 , \AES_ENC/us10/n672 ,\AES_ENC/us10/n671 , \AES_ENC/us10/n670 , \AES_ENC/us10/n669 ,\AES_ENC/us10/n668 , \AES_ENC/us10/n667 , \AES_ENC/us10/n666 ,\AES_ENC/us10/n665 , \AES_ENC/us10/n664 , \AES_ENC/us10/n663 ,\AES_ENC/us10/n662 , \AES_ENC/us10/n661 , \AES_ENC/us10/n660 ,\AES_ENC/us10/n659 , \AES_ENC/us10/n658 , \AES_ENC/us10/n657 ,\AES_ENC/us10/n656 , \AES_ENC/us10/n655 , \AES_ENC/us10/n654 ,\AES_ENC/us10/n653 , \AES_ENC/us10/n652 , \AES_ENC/us10/n651 ,\AES_ENC/us10/n650 , \AES_ENC/us10/n649 , \AES_ENC/us10/n648 ,\AES_ENC/us10/n647 , \AES_ENC/us10/n646 , \AES_ENC/us10/n645 ,\AES_ENC/us10/n644 , \AES_ENC/us10/n643 , \AES_ENC/us10/n642 ,\AES_ENC/us10/n641 , \AES_ENC/us10/n640 , \AES_ENC/us10/n639 ,\AES_ENC/us10/n638 , \AES_ENC/us10/n637 , \AES_ENC/us10/n636 ,\AES_ENC/us10/n635 , \AES_ENC/us10/n634 , \AES_ENC/us10/n633 ,\AES_ENC/us10/n632 , \AES_ENC/us10/n631 , \AES_ENC/us10/n630 ,\AES_ENC/us10/n629 , \AES_ENC/us10/n628 , \AES_ENC/us10/n627 ,\AES_ENC/us10/n626 , \AES_ENC/us10/n625 , \AES_ENC/us10/n624 ,\AES_ENC/us10/n623 , \AES_ENC/us10/n622 , \AES_ENC/us10/n621 ,\AES_ENC/us10/n620 , \AES_ENC/us10/n619 , \AES_ENC/us10/n618 ,\AES_ENC/us10/n617 , \AES_ENC/us10/n616 , \AES_ENC/us10/n615 ,\AES_ENC/us10/n614 , \AES_ENC/us10/n613 , \AES_ENC/us10/n612 ,\AES_ENC/us10/n611 , \AES_ENC/us10/n610 , \AES_ENC/us10/n609 ,\AES_ENC/us10/n608 , \AES_ENC/us10/n607 , \AES_ENC/us10/n606 ,\AES_ENC/us10/n605 , \AES_ENC/us10/n604 , \AES_ENC/us10/n603 ,\AES_ENC/us10/n602 , \AES_ENC/us10/n601 , \AES_ENC/us10/n600 ,\AES_ENC/us10/n599 , \AES_ENC/us10/n598 , \AES_ENC/us10/n597 ,\AES_ENC/us10/n596 , \AES_ENC/us10/n595 , \AES_ENC/us10/n594 ,\AES_ENC/us10/n593 , \AES_ENC/us10/n592 , \AES_ENC/us10/n591 ,\AES_ENC/us10/n590 , \AES_ENC/us10/n589 , \AES_ENC/us10/n588 ,\AES_ENC/us10/n587 , \AES_ENC/us10/n586 , \AES_ENC/us10/n585 ,\AES_ENC/us10/n584 , \AES_ENC/us10/n583 , \AES_ENC/us10/n582 ,\AES_ENC/us10/n581 , \AES_ENC/us10/n580 , \AES_ENC/us10/n579 ,\AES_ENC/us10/n578 , \AES_ENC/us10/n577 , \AES_ENC/us10/n576 ,\AES_ENC/us10/n575 , \AES_ENC/us10/n574 , \AES_ENC/us10/n573 ,\AES_ENC/us10/n572 , \AES_ENC/us10/n571 , \AES_ENC/us10/n570 ,\AES_ENC/us10/n569 , \AES_ENC/us11/n1135 , \AES_ENC/us11/n1134 ,\AES_ENC/us11/n1133 , \AES_ENC/us11/n1132 , \AES_ENC/us11/n1131 ,\AES_ENC/us11/n1130 , \AES_ENC/us11/n1129 , \AES_ENC/us11/n1128 ,\AES_ENC/us11/n1127 , \AES_ENC/us11/n1126 , \AES_ENC/us11/n1125 ,\AES_ENC/us11/n1124 , \AES_ENC/us11/n1123 , \AES_ENC/us11/n1122 ,\AES_ENC/us11/n1121 , \AES_ENC/us11/n1120 , \AES_ENC/us11/n1119 ,\AES_ENC/us11/n1118 , \AES_ENC/us11/n1117 , \AES_ENC/us11/n1116 ,\AES_ENC/us11/n1115 , \AES_ENC/us11/n1114 , \AES_ENC/us11/n1113 ,\AES_ENC/us11/n1112 , \AES_ENC/us11/n1111 , \AES_ENC/us11/n1110 ,\AES_ENC/us11/n1109 , \AES_ENC/us11/n1108 , \AES_ENC/us11/n1107 ,\AES_ENC/us11/n1106 , \AES_ENC/us11/n1105 , \AES_ENC/us11/n1104 ,\AES_ENC/us11/n1103 , \AES_ENC/us11/n1102 , \AES_ENC/us11/n1101 ,\AES_ENC/us11/n1100 , \AES_ENC/us11/n1099 , \AES_ENC/us11/n1098 ,\AES_ENC/us11/n1097 , \AES_ENC/us11/n1096 , \AES_ENC/us11/n1095 ,\AES_ENC/us11/n1094 , \AES_ENC/us11/n1093 , \AES_ENC/us11/n1092 ,\AES_ENC/us11/n1091 , \AES_ENC/us11/n1090 , \AES_ENC/us11/n1089 ,\AES_ENC/us11/n1088 , \AES_ENC/us11/n1087 , \AES_ENC/us11/n1086 ,\AES_ENC/us11/n1085 , \AES_ENC/us11/n1084 , \AES_ENC/us11/n1083 ,\AES_ENC/us11/n1082 , \AES_ENC/us11/n1081 , \AES_ENC/us11/n1080 ,\AES_ENC/us11/n1079 , \AES_ENC/us11/n1078 , \AES_ENC/us11/n1077 ,\AES_ENC/us11/n1076 , \AES_ENC/us11/n1075 , \AES_ENC/us11/n1074 ,\AES_ENC/us11/n1073 , \AES_ENC/us11/n1072 , \AES_ENC/us11/n1071 ,\AES_ENC/us11/n1070 , \AES_ENC/us11/n1069 , \AES_ENC/us11/n1068 ,\AES_ENC/us11/n1067 , \AES_ENC/us11/n1066 , \AES_ENC/us11/n1065 ,\AES_ENC/us11/n1064 , \AES_ENC/us11/n1063 , \AES_ENC/us11/n1062 ,\AES_ENC/us11/n1061 , \AES_ENC/us11/n1060 , \AES_ENC/us11/n1059 ,\AES_ENC/us11/n1058 , \AES_ENC/us11/n1057 , \AES_ENC/us11/n1056 ,\AES_ENC/us11/n1055 , \AES_ENC/us11/n1054 , \AES_ENC/us11/n1053 ,\AES_ENC/us11/n1052 , \AES_ENC/us11/n1051 , \AES_ENC/us11/n1050 ,\AES_ENC/us11/n1049 , \AES_ENC/us11/n1048 , \AES_ENC/us11/n1047 ,\AES_ENC/us11/n1046 , \AES_ENC/us11/n1045 , \AES_ENC/us11/n1044 ,\AES_ENC/us11/n1043 , \AES_ENC/us11/n1042 , \AES_ENC/us11/n1041 ,\AES_ENC/us11/n1040 , \AES_ENC/us11/n1039 , \AES_ENC/us11/n1038 ,\AES_ENC/us11/n1037 , \AES_ENC/us11/n1036 , \AES_ENC/us11/n1035 ,\AES_ENC/us11/n1034 , \AES_ENC/us11/n1033 , \AES_ENC/us11/n1032 ,\AES_ENC/us11/n1031 , \AES_ENC/us11/n1030 , \AES_ENC/us11/n1029 ,\AES_ENC/us11/n1028 , \AES_ENC/us11/n1027 , \AES_ENC/us11/n1026 ,\AES_ENC/us11/n1025 , \AES_ENC/us11/n1024 , \AES_ENC/us11/n1023 ,\AES_ENC/us11/n1022 , \AES_ENC/us11/n1021 , \AES_ENC/us11/n1020 ,\AES_ENC/us11/n1019 , \AES_ENC/us11/n1018 , \AES_ENC/us11/n1017 ,\AES_ENC/us11/n1016 , \AES_ENC/us11/n1015 , \AES_ENC/us11/n1014 ,\AES_ENC/us11/n1013 , \AES_ENC/us11/n1012 , \AES_ENC/us11/n1011 ,\AES_ENC/us11/n1010 , \AES_ENC/us11/n1009 , \AES_ENC/us11/n1008 ,\AES_ENC/us11/n1007 , \AES_ENC/us11/n1006 , \AES_ENC/us11/n1005 ,\AES_ENC/us11/n1004 , \AES_ENC/us11/n1003 , \AES_ENC/us11/n1002 ,\AES_ENC/us11/n1001 , \AES_ENC/us11/n1000 , \AES_ENC/us11/n999 ,\AES_ENC/us11/n998 , \AES_ENC/us11/n997 , \AES_ENC/us11/n996 ,\AES_ENC/us11/n995 , \AES_ENC/us11/n994 , \AES_ENC/us11/n993 ,\AES_ENC/us11/n992 , \AES_ENC/us11/n991 , \AES_ENC/us11/n990 ,\AES_ENC/us11/n989 , \AES_ENC/us11/n988 , \AES_ENC/us11/n987 ,\AES_ENC/us11/n986 , \AES_ENC/us11/n985 , \AES_ENC/us11/n984 ,\AES_ENC/us11/n983 , \AES_ENC/us11/n982 , \AES_ENC/us11/n981 ,\AES_ENC/us11/n980 , \AES_ENC/us11/n979 , \AES_ENC/us11/n978 ,\AES_ENC/us11/n977 , \AES_ENC/us11/n976 , \AES_ENC/us11/n975 ,\AES_ENC/us11/n974 , \AES_ENC/us11/n973 , \AES_ENC/us11/n972 ,\AES_ENC/us11/n971 , \AES_ENC/us11/n970 , \AES_ENC/us11/n969 ,\AES_ENC/us11/n968 , \AES_ENC/us11/n967 , \AES_ENC/us11/n966 ,\AES_ENC/us11/n965 , \AES_ENC/us11/n964 , \AES_ENC/us11/n963 ,\AES_ENC/us11/n962 , \AES_ENC/us11/n961 , \AES_ENC/us11/n960 ,\AES_ENC/us11/n959 , \AES_ENC/us11/n958 , \AES_ENC/us11/n957 ,\AES_ENC/us11/n956 , \AES_ENC/us11/n955 , \AES_ENC/us11/n954 ,\AES_ENC/us11/n953 , \AES_ENC/us11/n952 , \AES_ENC/us11/n951 ,\AES_ENC/us11/n950 , \AES_ENC/us11/n949 , \AES_ENC/us11/n948 ,\AES_ENC/us11/n947 , \AES_ENC/us11/n946 , \AES_ENC/us11/n945 ,\AES_ENC/us11/n944 , \AES_ENC/us11/n943 , \AES_ENC/us11/n942 ,\AES_ENC/us11/n941 , \AES_ENC/us11/n940 , \AES_ENC/us11/n939 ,\AES_ENC/us11/n938 , \AES_ENC/us11/n937 , \AES_ENC/us11/n936 ,\AES_ENC/us11/n935 , \AES_ENC/us11/n934 , \AES_ENC/us11/n933 ,\AES_ENC/us11/n932 , \AES_ENC/us11/n931 , \AES_ENC/us11/n930 ,\AES_ENC/us11/n929 , \AES_ENC/us11/n928 , \AES_ENC/us11/n927 ,\AES_ENC/us11/n926 , \AES_ENC/us11/n925 , \AES_ENC/us11/n924 ,\AES_ENC/us11/n923 , \AES_ENC/us11/n922 , \AES_ENC/us11/n921 ,\AES_ENC/us11/n920 , \AES_ENC/us11/n919 , \AES_ENC/us11/n918 ,\AES_ENC/us11/n917 , \AES_ENC/us11/n916 , \AES_ENC/us11/n915 ,\AES_ENC/us11/n914 , \AES_ENC/us11/n913 , \AES_ENC/us11/n912 ,\AES_ENC/us11/n911 , \AES_ENC/us11/n910 , \AES_ENC/us11/n909 ,\AES_ENC/us11/n908 , \AES_ENC/us11/n907 , \AES_ENC/us11/n906 ,\AES_ENC/us11/n905 , \AES_ENC/us11/n904 , \AES_ENC/us11/n903 ,\AES_ENC/us11/n902 , \AES_ENC/us11/n901 , \AES_ENC/us11/n900 ,\AES_ENC/us11/n899 , \AES_ENC/us11/n898 , \AES_ENC/us11/n897 ,\AES_ENC/us11/n896 , \AES_ENC/us11/n895 , \AES_ENC/us11/n894 ,\AES_ENC/us11/n893 , \AES_ENC/us11/n892 , \AES_ENC/us11/n891 ,\AES_ENC/us11/n890 , \AES_ENC/us11/n889 , \AES_ENC/us11/n888 ,\AES_ENC/us11/n887 , \AES_ENC/us11/n886 , \AES_ENC/us11/n885 ,\AES_ENC/us11/n884 , \AES_ENC/us11/n883 , \AES_ENC/us11/n882 ,\AES_ENC/us11/n881 , \AES_ENC/us11/n880 , \AES_ENC/us11/n879 ,\AES_ENC/us11/n878 , \AES_ENC/us11/n877 , \AES_ENC/us11/n876 ,\AES_ENC/us11/n875 , \AES_ENC/us11/n874 , \AES_ENC/us11/n873 ,\AES_ENC/us11/n872 , \AES_ENC/us11/n871 , \AES_ENC/us11/n870 ,\AES_ENC/us11/n869 , \AES_ENC/us11/n868 , \AES_ENC/us11/n867 ,\AES_ENC/us11/n866 , \AES_ENC/us11/n865 , \AES_ENC/us11/n864 ,\AES_ENC/us11/n863 , \AES_ENC/us11/n862 , \AES_ENC/us11/n861 ,\AES_ENC/us11/n860 , \AES_ENC/us11/n859 , \AES_ENC/us11/n858 ,\AES_ENC/us11/n857 , \AES_ENC/us11/n856 , \AES_ENC/us11/n855 ,\AES_ENC/us11/n854 , \AES_ENC/us11/n853 , \AES_ENC/us11/n852 ,\AES_ENC/us11/n851 , \AES_ENC/us11/n850 , \AES_ENC/us11/n849 ,\AES_ENC/us11/n848 , \AES_ENC/us11/n847 , \AES_ENC/us11/n846 ,\AES_ENC/us11/n845 , \AES_ENC/us11/n844 , \AES_ENC/us11/n843 ,\AES_ENC/us11/n842 , \AES_ENC/us11/n841 , \AES_ENC/us11/n840 ,\AES_ENC/us11/n839 , \AES_ENC/us11/n838 , \AES_ENC/us11/n837 ,\AES_ENC/us11/n836 , \AES_ENC/us11/n835 , \AES_ENC/us11/n834 ,\AES_ENC/us11/n833 , \AES_ENC/us11/n832 , \AES_ENC/us11/n831 ,\AES_ENC/us11/n830 , \AES_ENC/us11/n829 , \AES_ENC/us11/n828 ,\AES_ENC/us11/n827 , \AES_ENC/us11/n826 , \AES_ENC/us11/n825 ,\AES_ENC/us11/n824 , \AES_ENC/us11/n823 , \AES_ENC/us11/n822 ,\AES_ENC/us11/n821 , \AES_ENC/us11/n820 , \AES_ENC/us11/n819 ,\AES_ENC/us11/n818 , \AES_ENC/us11/n817 , \AES_ENC/us11/n816 ,\AES_ENC/us11/n815 , \AES_ENC/us11/n814 , \AES_ENC/us11/n813 ,\AES_ENC/us11/n812 , \AES_ENC/us11/n811 , \AES_ENC/us11/n810 ,\AES_ENC/us11/n809 , \AES_ENC/us11/n808 , \AES_ENC/us11/n807 ,\AES_ENC/us11/n806 , \AES_ENC/us11/n805 , \AES_ENC/us11/n804 ,\AES_ENC/us11/n803 , \AES_ENC/us11/n802 , \AES_ENC/us11/n801 ,\AES_ENC/us11/n800 , \AES_ENC/us11/n799 , \AES_ENC/us11/n798 ,\AES_ENC/us11/n797 , \AES_ENC/us11/n796 , \AES_ENC/us11/n795 ,\AES_ENC/us11/n794 , \AES_ENC/us11/n793 , \AES_ENC/us11/n792 ,\AES_ENC/us11/n791 , \AES_ENC/us11/n790 , \AES_ENC/us11/n789 ,\AES_ENC/us11/n788 , \AES_ENC/us11/n787 , \AES_ENC/us11/n786 ,\AES_ENC/us11/n785 , \AES_ENC/us11/n784 , \AES_ENC/us11/n783 ,\AES_ENC/us11/n782 , \AES_ENC/us11/n781 , \AES_ENC/us11/n780 ,\AES_ENC/us11/n779 , \AES_ENC/us11/n778 , \AES_ENC/us11/n777 ,\AES_ENC/us11/n776 , \AES_ENC/us11/n775 , \AES_ENC/us11/n774 ,\AES_ENC/us11/n773 , \AES_ENC/us11/n772 , \AES_ENC/us11/n771 ,\AES_ENC/us11/n770 , \AES_ENC/us11/n769 , \AES_ENC/us11/n768 ,\AES_ENC/us11/n767 , \AES_ENC/us11/n766 , \AES_ENC/us11/n765 ,\AES_ENC/us11/n764 , \AES_ENC/us11/n763 , \AES_ENC/us11/n762 ,\AES_ENC/us11/n761 , \AES_ENC/us11/n760 , \AES_ENC/us11/n759 ,\AES_ENC/us11/n758 , \AES_ENC/us11/n757 , \AES_ENC/us11/n756 ,\AES_ENC/us11/n755 , \AES_ENC/us11/n754 , \AES_ENC/us11/n753 ,\AES_ENC/us11/n752 , \AES_ENC/us11/n751 , \AES_ENC/us11/n750 ,\AES_ENC/us11/n749 , \AES_ENC/us11/n748 , \AES_ENC/us11/n747 ,\AES_ENC/us11/n746 , \AES_ENC/us11/n745 , \AES_ENC/us11/n744 ,\AES_ENC/us11/n743 , \AES_ENC/us11/n742 , \AES_ENC/us11/n741 ,\AES_ENC/us11/n740 , \AES_ENC/us11/n739 , \AES_ENC/us11/n738 ,\AES_ENC/us11/n737 , \AES_ENC/us11/n736 , \AES_ENC/us11/n735 ,\AES_ENC/us11/n734 , \AES_ENC/us11/n733 , \AES_ENC/us11/n732 ,\AES_ENC/us11/n731 , \AES_ENC/us11/n730 , \AES_ENC/us11/n729 ,\AES_ENC/us11/n728 , \AES_ENC/us11/n727 , \AES_ENC/us11/n726 ,\AES_ENC/us11/n725 , \AES_ENC/us11/n724 , \AES_ENC/us11/n723 ,\AES_ENC/us11/n722 , \AES_ENC/us11/n721 , \AES_ENC/us11/n720 ,\AES_ENC/us11/n719 , \AES_ENC/us11/n718 , \AES_ENC/us11/n717 ,\AES_ENC/us11/n716 , \AES_ENC/us11/n715 , \AES_ENC/us11/n714 ,\AES_ENC/us11/n713 , \AES_ENC/us11/n712 , \AES_ENC/us11/n711 ,\AES_ENC/us11/n710 , \AES_ENC/us11/n709 , \AES_ENC/us11/n708 ,\AES_ENC/us11/n707 , \AES_ENC/us11/n706 , \AES_ENC/us11/n705 ,\AES_ENC/us11/n704 , \AES_ENC/us11/n703 , \AES_ENC/us11/n702 ,\AES_ENC/us11/n701 , \AES_ENC/us11/n700 , \AES_ENC/us11/n699 ,\AES_ENC/us11/n698 , \AES_ENC/us11/n697 , \AES_ENC/us11/n696 ,\AES_ENC/us11/n695 , \AES_ENC/us11/n694 , \AES_ENC/us11/n693 ,\AES_ENC/us11/n692 , \AES_ENC/us11/n691 , \AES_ENC/us11/n690 ,\AES_ENC/us11/n689 , \AES_ENC/us11/n688 , \AES_ENC/us11/n687 ,\AES_ENC/us11/n686 , \AES_ENC/us11/n685 , \AES_ENC/us11/n684 ,\AES_ENC/us11/n683 , \AES_ENC/us11/n682 , \AES_ENC/us11/n681 ,\AES_ENC/us11/n680 , \AES_ENC/us11/n679 , \AES_ENC/us11/n678 ,\AES_ENC/us11/n677 , \AES_ENC/us11/n676 , \AES_ENC/us11/n675 ,\AES_ENC/us11/n674 , \AES_ENC/us11/n673 , \AES_ENC/us11/n672 ,\AES_ENC/us11/n671 , \AES_ENC/us11/n670 , \AES_ENC/us11/n669 ,\AES_ENC/us11/n668 , \AES_ENC/us11/n667 , \AES_ENC/us11/n666 ,\AES_ENC/us11/n665 , \AES_ENC/us11/n664 , \AES_ENC/us11/n663 ,\AES_ENC/us11/n662 , \AES_ENC/us11/n661 , \AES_ENC/us11/n660 ,\AES_ENC/us11/n659 , \AES_ENC/us11/n658 , \AES_ENC/us11/n657 ,\AES_ENC/us11/n656 , \AES_ENC/us11/n655 , \AES_ENC/us11/n654 ,\AES_ENC/us11/n653 , \AES_ENC/us11/n652 , \AES_ENC/us11/n651 ,\AES_ENC/us11/n650 , \AES_ENC/us11/n649 , \AES_ENC/us11/n648 ,\AES_ENC/us11/n647 , \AES_ENC/us11/n646 , \AES_ENC/us11/n645 ,\AES_ENC/us11/n644 , \AES_ENC/us11/n643 , \AES_ENC/us11/n642 ,\AES_ENC/us11/n641 , \AES_ENC/us11/n640 , \AES_ENC/us11/n639 ,\AES_ENC/us11/n638 , \AES_ENC/us11/n637 , \AES_ENC/us11/n636 ,\AES_ENC/us11/n635 , \AES_ENC/us11/n634 , \AES_ENC/us11/n633 ,\AES_ENC/us11/n632 , \AES_ENC/us11/n631 , \AES_ENC/us11/n630 ,\AES_ENC/us11/n629 , \AES_ENC/us11/n628 , \AES_ENC/us11/n627 ,\AES_ENC/us11/n626 , \AES_ENC/us11/n625 , \AES_ENC/us11/n624 ,\AES_ENC/us11/n623 , \AES_ENC/us11/n622 , \AES_ENC/us11/n621 ,\AES_ENC/us11/n620 , \AES_ENC/us11/n619 , \AES_ENC/us11/n618 ,\AES_ENC/us11/n617 , \AES_ENC/us11/n616 , \AES_ENC/us11/n615 ,\AES_ENC/us11/n614 , \AES_ENC/us11/n613 , \AES_ENC/us11/n612 ,\AES_ENC/us11/n611 , \AES_ENC/us11/n610 , \AES_ENC/us11/n609 ,\AES_ENC/us11/n608 , \AES_ENC/us11/n607 , \AES_ENC/us11/n606 ,\AES_ENC/us11/n605 , \AES_ENC/us11/n604 , \AES_ENC/us11/n603 ,\AES_ENC/us11/n602 , \AES_ENC/us11/n601 , \AES_ENC/us11/n600 ,\AES_ENC/us11/n599 , \AES_ENC/us11/n598 , \AES_ENC/us11/n597 ,\AES_ENC/us11/n596 , \AES_ENC/us11/n595 , \AES_ENC/us11/n594 ,\AES_ENC/us11/n593 , \AES_ENC/us11/n592 , \AES_ENC/us11/n591 ,\AES_ENC/us11/n590 , \AES_ENC/us11/n589 , \AES_ENC/us11/n588 ,\AES_ENC/us11/n587 , \AES_ENC/us11/n586 , \AES_ENC/us11/n585 ,\AES_ENC/us11/n584 , \AES_ENC/us11/n583 , \AES_ENC/us11/n582 ,\AES_ENC/us11/n581 , \AES_ENC/us11/n580 , \AES_ENC/us11/n579 ,\AES_ENC/us11/n578 , \AES_ENC/us11/n577 , \AES_ENC/us11/n576 ,\AES_ENC/us11/n575 , \AES_ENC/us11/n574 , \AES_ENC/us11/n573 ,\AES_ENC/us11/n572 , \AES_ENC/us11/n571 , \AES_ENC/us11/n570 ,\AES_ENC/us11/n569 , \AES_ENC/us12/n1135 , \AES_ENC/us12/n1134 ,\AES_ENC/us12/n1133 , \AES_ENC/us12/n1132 , \AES_ENC/us12/n1131 ,\AES_ENC/us12/n1130 , \AES_ENC/us12/n1129 , \AES_ENC/us12/n1128 ,\AES_ENC/us12/n1127 , \AES_ENC/us12/n1126 , \AES_ENC/us12/n1125 ,\AES_ENC/us12/n1124 , \AES_ENC/us12/n1123 , \AES_ENC/us12/n1122 ,\AES_ENC/us12/n1121 , \AES_ENC/us12/n1120 , \AES_ENC/us12/n1119 ,\AES_ENC/us12/n1118 , \AES_ENC/us12/n1117 , \AES_ENC/us12/n1116 ,\AES_ENC/us12/n1115 , \AES_ENC/us12/n1114 , \AES_ENC/us12/n1113 ,\AES_ENC/us12/n1112 , \AES_ENC/us12/n1111 , \AES_ENC/us12/n1110 ,\AES_ENC/us12/n1109 , \AES_ENC/us12/n1108 , \AES_ENC/us12/n1107 ,\AES_ENC/us12/n1106 , \AES_ENC/us12/n1105 , \AES_ENC/us12/n1104 ,\AES_ENC/us12/n1103 , \AES_ENC/us12/n1102 , \AES_ENC/us12/n1101 ,\AES_ENC/us12/n1100 , \AES_ENC/us12/n1099 , \AES_ENC/us12/n1098 ,\AES_ENC/us12/n1097 , \AES_ENC/us12/n1096 , \AES_ENC/us12/n1095 ,\AES_ENC/us12/n1094 , \AES_ENC/us12/n1093 , \AES_ENC/us12/n1092 ,\AES_ENC/us12/n1091 , \AES_ENC/us12/n1090 , \AES_ENC/us12/n1089 ,\AES_ENC/us12/n1088 , \AES_ENC/us12/n1087 , \AES_ENC/us12/n1086 ,\AES_ENC/us12/n1085 , \AES_ENC/us12/n1084 , \AES_ENC/us12/n1083 ,\AES_ENC/us12/n1082 , \AES_ENC/us12/n1081 , \AES_ENC/us12/n1080 ,\AES_ENC/us12/n1079 , \AES_ENC/us12/n1078 , \AES_ENC/us12/n1077 ,\AES_ENC/us12/n1076 , \AES_ENC/us12/n1075 , \AES_ENC/us12/n1074 ,\AES_ENC/us12/n1073 , \AES_ENC/us12/n1072 , \AES_ENC/us12/n1071 ,\AES_ENC/us12/n1070 , \AES_ENC/us12/n1069 , \AES_ENC/us12/n1068 ,\AES_ENC/us12/n1067 , \AES_ENC/us12/n1066 , \AES_ENC/us12/n1065 ,\AES_ENC/us12/n1064 , \AES_ENC/us12/n1063 , \AES_ENC/us12/n1062 ,\AES_ENC/us12/n1061 , \AES_ENC/us12/n1060 , \AES_ENC/us12/n1059 ,\AES_ENC/us12/n1058 , \AES_ENC/us12/n1057 , \AES_ENC/us12/n1056 ,\AES_ENC/us12/n1055 , \AES_ENC/us12/n1054 , \AES_ENC/us12/n1053 ,\AES_ENC/us12/n1052 , \AES_ENC/us12/n1051 , \AES_ENC/us12/n1050 ,\AES_ENC/us12/n1049 , \AES_ENC/us12/n1048 , \AES_ENC/us12/n1047 ,\AES_ENC/us12/n1046 , \AES_ENC/us12/n1045 , \AES_ENC/us12/n1044 ,\AES_ENC/us12/n1043 , \AES_ENC/us12/n1042 , \AES_ENC/us12/n1041 ,\AES_ENC/us12/n1040 , \AES_ENC/us12/n1039 , \AES_ENC/us12/n1038 ,\AES_ENC/us12/n1037 , \AES_ENC/us12/n1036 , \AES_ENC/us12/n1035 ,\AES_ENC/us12/n1034 , \AES_ENC/us12/n1033 , \AES_ENC/us12/n1032 ,\AES_ENC/us12/n1031 , \AES_ENC/us12/n1030 , \AES_ENC/us12/n1029 ,\AES_ENC/us12/n1028 , \AES_ENC/us12/n1027 , \AES_ENC/us12/n1026 ,\AES_ENC/us12/n1025 , \AES_ENC/us12/n1024 , \AES_ENC/us12/n1023 ,\AES_ENC/us12/n1022 , \AES_ENC/us12/n1021 , \AES_ENC/us12/n1020 ,\AES_ENC/us12/n1019 , \AES_ENC/us12/n1018 , \AES_ENC/us12/n1017 ,\AES_ENC/us12/n1016 , \AES_ENC/us12/n1015 , \AES_ENC/us12/n1014 ,\AES_ENC/us12/n1013 , \AES_ENC/us12/n1012 , \AES_ENC/us12/n1011 ,\AES_ENC/us12/n1010 , \AES_ENC/us12/n1009 , \AES_ENC/us12/n1008 ,\AES_ENC/us12/n1007 , \AES_ENC/us12/n1006 , \AES_ENC/us12/n1005 ,\AES_ENC/us12/n1004 , \AES_ENC/us12/n1003 , \AES_ENC/us12/n1002 ,\AES_ENC/us12/n1001 , \AES_ENC/us12/n1000 , \AES_ENC/us12/n999 ,\AES_ENC/us12/n998 , \AES_ENC/us12/n997 , \AES_ENC/us12/n996 ,\AES_ENC/us12/n995 , \AES_ENC/us12/n994 , \AES_ENC/us12/n993 ,\AES_ENC/us12/n992 , \AES_ENC/us12/n991 , \AES_ENC/us12/n990 ,\AES_ENC/us12/n989 , \AES_ENC/us12/n988 , \AES_ENC/us12/n987 ,\AES_ENC/us12/n986 , \AES_ENC/us12/n985 , \AES_ENC/us12/n984 ,\AES_ENC/us12/n983 , \AES_ENC/us12/n982 , \AES_ENC/us12/n981 ,\AES_ENC/us12/n980 , \AES_ENC/us12/n979 , \AES_ENC/us12/n978 ,\AES_ENC/us12/n977 , \AES_ENC/us12/n976 , \AES_ENC/us12/n975 ,\AES_ENC/us12/n974 , \AES_ENC/us12/n973 , \AES_ENC/us12/n972 ,\AES_ENC/us12/n971 , \AES_ENC/us12/n970 , \AES_ENC/us12/n969 ,\AES_ENC/us12/n968 , \AES_ENC/us12/n967 , \AES_ENC/us12/n966 ,\AES_ENC/us12/n965 , \AES_ENC/us12/n964 , \AES_ENC/us12/n963 ,\AES_ENC/us12/n962 , \AES_ENC/us12/n961 , \AES_ENC/us12/n960 ,\AES_ENC/us12/n959 , \AES_ENC/us12/n958 , \AES_ENC/us12/n957 ,\AES_ENC/us12/n956 , \AES_ENC/us12/n955 , \AES_ENC/us12/n954 ,\AES_ENC/us12/n953 , \AES_ENC/us12/n952 , \AES_ENC/us12/n951 ,\AES_ENC/us12/n950 , \AES_ENC/us12/n949 , \AES_ENC/us12/n948 ,\AES_ENC/us12/n947 , \AES_ENC/us12/n946 , \AES_ENC/us12/n945 ,\AES_ENC/us12/n944 , \AES_ENC/us12/n943 , \AES_ENC/us12/n942 ,\AES_ENC/us12/n941 , \AES_ENC/us12/n940 , \AES_ENC/us12/n939 ,\AES_ENC/us12/n938 , \AES_ENC/us12/n937 , \AES_ENC/us12/n936 ,\AES_ENC/us12/n935 , \AES_ENC/us12/n934 , \AES_ENC/us12/n933 ,\AES_ENC/us12/n932 , \AES_ENC/us12/n931 , \AES_ENC/us12/n930 ,\AES_ENC/us12/n929 , \AES_ENC/us12/n928 , \AES_ENC/us12/n927 ,\AES_ENC/us12/n926 , \AES_ENC/us12/n925 , \AES_ENC/us12/n924 ,\AES_ENC/us12/n923 , \AES_ENC/us12/n922 , \AES_ENC/us12/n921 ,\AES_ENC/us12/n920 , \AES_ENC/us12/n919 , \AES_ENC/us12/n918 ,\AES_ENC/us12/n917 , \AES_ENC/us12/n916 , \AES_ENC/us12/n915 ,\AES_ENC/us12/n914 , \AES_ENC/us12/n913 , \AES_ENC/us12/n912 ,\AES_ENC/us12/n911 , \AES_ENC/us12/n910 , \AES_ENC/us12/n909 ,\AES_ENC/us12/n908 , \AES_ENC/us12/n907 , \AES_ENC/us12/n906 ,\AES_ENC/us12/n905 , \AES_ENC/us12/n904 , \AES_ENC/us12/n903 ,\AES_ENC/us12/n902 , \AES_ENC/us12/n901 , \AES_ENC/us12/n900 ,\AES_ENC/us12/n899 , \AES_ENC/us12/n898 , \AES_ENC/us12/n897 ,\AES_ENC/us12/n896 , \AES_ENC/us12/n895 , \AES_ENC/us12/n894 ,\AES_ENC/us12/n893 , \AES_ENC/us12/n892 , \AES_ENC/us12/n891 ,\AES_ENC/us12/n890 , \AES_ENC/us12/n889 , \AES_ENC/us12/n888 ,\AES_ENC/us12/n887 , \AES_ENC/us12/n886 , \AES_ENC/us12/n885 ,\AES_ENC/us12/n884 , \AES_ENC/us12/n883 , \AES_ENC/us12/n882 ,\AES_ENC/us12/n881 , \AES_ENC/us12/n880 , \AES_ENC/us12/n879 ,\AES_ENC/us12/n878 , \AES_ENC/us12/n877 , \AES_ENC/us12/n876 ,\AES_ENC/us12/n875 , \AES_ENC/us12/n874 , \AES_ENC/us12/n873 ,\AES_ENC/us12/n872 , \AES_ENC/us12/n871 , \AES_ENC/us12/n870 ,\AES_ENC/us12/n869 , \AES_ENC/us12/n868 , \AES_ENC/us12/n867 ,\AES_ENC/us12/n866 , \AES_ENC/us12/n865 , \AES_ENC/us12/n864 ,\AES_ENC/us12/n863 , \AES_ENC/us12/n862 , \AES_ENC/us12/n861 ,\AES_ENC/us12/n860 , \AES_ENC/us12/n859 , \AES_ENC/us12/n858 ,\AES_ENC/us12/n857 , \AES_ENC/us12/n856 , \AES_ENC/us12/n855 ,\AES_ENC/us12/n854 , \AES_ENC/us12/n853 , \AES_ENC/us12/n852 ,\AES_ENC/us12/n851 , \AES_ENC/us12/n850 , \AES_ENC/us12/n849 ,\AES_ENC/us12/n848 , \AES_ENC/us12/n847 , \AES_ENC/us12/n846 ,\AES_ENC/us12/n845 , \AES_ENC/us12/n844 , \AES_ENC/us12/n843 ,\AES_ENC/us12/n842 , \AES_ENC/us12/n841 , \AES_ENC/us12/n840 ,\AES_ENC/us12/n839 , \AES_ENC/us12/n838 , \AES_ENC/us12/n837 ,\AES_ENC/us12/n836 , \AES_ENC/us12/n835 , \AES_ENC/us12/n834 ,\AES_ENC/us12/n833 , \AES_ENC/us12/n832 , \AES_ENC/us12/n831 ,\AES_ENC/us12/n830 , \AES_ENC/us12/n829 , \AES_ENC/us12/n828 ,\AES_ENC/us12/n827 , \AES_ENC/us12/n826 , \AES_ENC/us12/n825 ,\AES_ENC/us12/n824 , \AES_ENC/us12/n823 , \AES_ENC/us12/n822 ,\AES_ENC/us12/n821 , \AES_ENC/us12/n820 , \AES_ENC/us12/n819 ,\AES_ENC/us12/n818 , \AES_ENC/us12/n817 , \AES_ENC/us12/n816 ,\AES_ENC/us12/n815 , \AES_ENC/us12/n814 , \AES_ENC/us12/n813 ,\AES_ENC/us12/n812 , \AES_ENC/us12/n811 , \AES_ENC/us12/n810 ,\AES_ENC/us12/n809 , \AES_ENC/us12/n808 , \AES_ENC/us12/n807 ,\AES_ENC/us12/n806 , \AES_ENC/us12/n805 , \AES_ENC/us12/n804 ,\AES_ENC/us12/n803 , \AES_ENC/us12/n802 , \AES_ENC/us12/n801 ,\AES_ENC/us12/n800 , \AES_ENC/us12/n799 , \AES_ENC/us12/n798 ,\AES_ENC/us12/n797 , \AES_ENC/us12/n796 , \AES_ENC/us12/n795 ,\AES_ENC/us12/n794 , \AES_ENC/us12/n793 , \AES_ENC/us12/n792 ,\AES_ENC/us12/n791 , \AES_ENC/us12/n790 , \AES_ENC/us12/n789 ,\AES_ENC/us12/n788 , \AES_ENC/us12/n787 , \AES_ENC/us12/n786 ,\AES_ENC/us12/n785 , \AES_ENC/us12/n784 , \AES_ENC/us12/n783 ,\AES_ENC/us12/n782 , \AES_ENC/us12/n781 , \AES_ENC/us12/n780 ,\AES_ENC/us12/n779 , \AES_ENC/us12/n778 , \AES_ENC/us12/n777 ,\AES_ENC/us12/n776 , \AES_ENC/us12/n775 , \AES_ENC/us12/n774 ,\AES_ENC/us12/n773 , \AES_ENC/us12/n772 , \AES_ENC/us12/n771 ,\AES_ENC/us12/n770 , \AES_ENC/us12/n769 , \AES_ENC/us12/n768 ,\AES_ENC/us12/n767 , \AES_ENC/us12/n766 , \AES_ENC/us12/n765 ,\AES_ENC/us12/n764 , \AES_ENC/us12/n763 , \AES_ENC/us12/n762 ,\AES_ENC/us12/n761 , \AES_ENC/us12/n760 , \AES_ENC/us12/n759 ,\AES_ENC/us12/n758 , \AES_ENC/us12/n757 , \AES_ENC/us12/n756 ,\AES_ENC/us12/n755 , \AES_ENC/us12/n754 , \AES_ENC/us12/n753 ,\AES_ENC/us12/n752 , \AES_ENC/us12/n751 , \AES_ENC/us12/n750 ,\AES_ENC/us12/n749 , \AES_ENC/us12/n748 , \AES_ENC/us12/n747 ,\AES_ENC/us12/n746 , \AES_ENC/us12/n745 , \AES_ENC/us12/n744 ,\AES_ENC/us12/n743 , \AES_ENC/us12/n742 , \AES_ENC/us12/n741 ,\AES_ENC/us12/n740 , \AES_ENC/us12/n739 , \AES_ENC/us12/n738 ,\AES_ENC/us12/n737 , \AES_ENC/us12/n736 , \AES_ENC/us12/n735 ,\AES_ENC/us12/n734 , \AES_ENC/us12/n733 , \AES_ENC/us12/n732 ,\AES_ENC/us12/n731 , \AES_ENC/us12/n730 , \AES_ENC/us12/n729 ,\AES_ENC/us12/n728 , \AES_ENC/us12/n727 , \AES_ENC/us12/n726 ,\AES_ENC/us12/n725 , \AES_ENC/us12/n724 , \AES_ENC/us12/n723 ,\AES_ENC/us12/n722 , \AES_ENC/us12/n721 , \AES_ENC/us12/n720 ,\AES_ENC/us12/n719 , \AES_ENC/us12/n718 , \AES_ENC/us12/n717 ,\AES_ENC/us12/n716 , \AES_ENC/us12/n715 , \AES_ENC/us12/n714 ,\AES_ENC/us12/n713 , \AES_ENC/us12/n712 , \AES_ENC/us12/n711 ,\AES_ENC/us12/n710 , \AES_ENC/us12/n709 , \AES_ENC/us12/n708 ,\AES_ENC/us12/n707 , \AES_ENC/us12/n706 , \AES_ENC/us12/n705 ,\AES_ENC/us12/n704 , \AES_ENC/us12/n703 , \AES_ENC/us12/n702 ,\AES_ENC/us12/n701 , \AES_ENC/us12/n700 , \AES_ENC/us12/n699 ,\AES_ENC/us12/n698 , \AES_ENC/us12/n697 , \AES_ENC/us12/n696 ,\AES_ENC/us12/n695 , \AES_ENC/us12/n694 , \AES_ENC/us12/n693 ,\AES_ENC/us12/n692 , \AES_ENC/us12/n691 , \AES_ENC/us12/n690 ,\AES_ENC/us12/n689 , \AES_ENC/us12/n688 , \AES_ENC/us12/n687 ,\AES_ENC/us12/n686 , \AES_ENC/us12/n685 , \AES_ENC/us12/n684 ,\AES_ENC/us12/n683 , \AES_ENC/us12/n682 , \AES_ENC/us12/n681 ,\AES_ENC/us12/n680 , \AES_ENC/us12/n679 , \AES_ENC/us12/n678 ,\AES_ENC/us12/n677 , \AES_ENC/us12/n676 , \AES_ENC/us12/n675 ,\AES_ENC/us12/n674 , \AES_ENC/us12/n673 , \AES_ENC/us12/n672 ,\AES_ENC/us12/n671 , \AES_ENC/us12/n670 , \AES_ENC/us12/n669 ,\AES_ENC/us12/n668 , \AES_ENC/us12/n667 , \AES_ENC/us12/n666 ,\AES_ENC/us12/n665 , \AES_ENC/us12/n664 , \AES_ENC/us12/n663 ,\AES_ENC/us12/n662 , \AES_ENC/us12/n661 , \AES_ENC/us12/n660 ,\AES_ENC/us12/n659 , \AES_ENC/us12/n658 , \AES_ENC/us12/n657 ,\AES_ENC/us12/n656 , \AES_ENC/us12/n655 , \AES_ENC/us12/n654 ,\AES_ENC/us12/n653 , \AES_ENC/us12/n652 , \AES_ENC/us12/n651 ,\AES_ENC/us12/n650 , \AES_ENC/us12/n649 , \AES_ENC/us12/n648 ,\AES_ENC/us12/n647 , \AES_ENC/us12/n646 , \AES_ENC/us12/n645 ,\AES_ENC/us12/n644 , \AES_ENC/us12/n643 , \AES_ENC/us12/n642 ,\AES_ENC/us12/n641 , \AES_ENC/us12/n640 , \AES_ENC/us12/n639 ,\AES_ENC/us12/n638 , \AES_ENC/us12/n637 , \AES_ENC/us12/n636 ,\AES_ENC/us12/n635 , \AES_ENC/us12/n634 , \AES_ENC/us12/n633 ,\AES_ENC/us12/n632 , \AES_ENC/us12/n631 , \AES_ENC/us12/n630 ,\AES_ENC/us12/n629 , \AES_ENC/us12/n628 , \AES_ENC/us12/n627 ,\AES_ENC/us12/n626 , \AES_ENC/us12/n625 , \AES_ENC/us12/n624 ,\AES_ENC/us12/n623 , \AES_ENC/us12/n622 , \AES_ENC/us12/n621 ,\AES_ENC/us12/n620 , \AES_ENC/us12/n619 , \AES_ENC/us12/n618 ,\AES_ENC/us12/n617 , \AES_ENC/us12/n616 , \AES_ENC/us12/n615 ,\AES_ENC/us12/n614 , \AES_ENC/us12/n613 , \AES_ENC/us12/n612 ,\AES_ENC/us12/n611 , \AES_ENC/us12/n610 , \AES_ENC/us12/n609 ,\AES_ENC/us12/n608 , \AES_ENC/us12/n607 , \AES_ENC/us12/n606 ,\AES_ENC/us12/n605 , \AES_ENC/us12/n604 , \AES_ENC/us12/n603 ,\AES_ENC/us12/n602 , \AES_ENC/us12/n601 , \AES_ENC/us12/n600 ,\AES_ENC/us12/n599 , \AES_ENC/us12/n598 , \AES_ENC/us12/n597 ,\AES_ENC/us12/n596 , \AES_ENC/us12/n595 , \AES_ENC/us12/n594 ,\AES_ENC/us12/n593 , \AES_ENC/us12/n592 , \AES_ENC/us12/n591 ,\AES_ENC/us12/n590 , \AES_ENC/us12/n589 , \AES_ENC/us12/n588 ,\AES_ENC/us12/n587 , \AES_ENC/us12/n586 , \AES_ENC/us12/n585 ,\AES_ENC/us12/n584 , \AES_ENC/us12/n583 , \AES_ENC/us12/n582 ,\AES_ENC/us12/n581 , \AES_ENC/us12/n580 , \AES_ENC/us12/n579 ,\AES_ENC/us12/n578 , \AES_ENC/us12/n577 , \AES_ENC/us12/n576 ,\AES_ENC/us12/n575 , \AES_ENC/us12/n574 , \AES_ENC/us12/n573 ,\AES_ENC/us12/n572 , \AES_ENC/us12/n571 , \AES_ENC/us12/n570 ,\AES_ENC/us12/n569 , \AES_ENC/us13/n1135 , \AES_ENC/us13/n1134 ,\AES_ENC/us13/n1133 , \AES_ENC/us13/n1132 , \AES_ENC/us13/n1131 ,\AES_ENC/us13/n1130 , \AES_ENC/us13/n1129 , \AES_ENC/us13/n1128 ,\AES_ENC/us13/n1127 , \AES_ENC/us13/n1126 , \AES_ENC/us13/n1125 ,\AES_ENC/us13/n1124 , \AES_ENC/us13/n1123 , \AES_ENC/us13/n1122 ,\AES_ENC/us13/n1121 , \AES_ENC/us13/n1120 , \AES_ENC/us13/n1119 ,\AES_ENC/us13/n1118 , \AES_ENC/us13/n1117 , \AES_ENC/us13/n1116 ,\AES_ENC/us13/n1115 , \AES_ENC/us13/n1114 , \AES_ENC/us13/n1113 ,\AES_ENC/us13/n1112 , \AES_ENC/us13/n1111 , \AES_ENC/us13/n1110 ,\AES_ENC/us13/n1109 , \AES_ENC/us13/n1108 , \AES_ENC/us13/n1107 ,\AES_ENC/us13/n1106 , \AES_ENC/us13/n1105 , \AES_ENC/us13/n1104 ,\AES_ENC/us13/n1103 , \AES_ENC/us13/n1102 , \AES_ENC/us13/n1101 ,\AES_ENC/us13/n1100 , \AES_ENC/us13/n1099 , \AES_ENC/us13/n1098 ,\AES_ENC/us13/n1097 , \AES_ENC/us13/n1096 , \AES_ENC/us13/n1095 ,\AES_ENC/us13/n1094 , \AES_ENC/us13/n1093 , \AES_ENC/us13/n1092 ,\AES_ENC/us13/n1091 , \AES_ENC/us13/n1090 , \AES_ENC/us13/n1089 ,\AES_ENC/us13/n1088 , \AES_ENC/us13/n1087 , \AES_ENC/us13/n1086 ,\AES_ENC/us13/n1085 , \AES_ENC/us13/n1084 , \AES_ENC/us13/n1083 ,\AES_ENC/us13/n1082 , \AES_ENC/us13/n1081 , \AES_ENC/us13/n1080 ,\AES_ENC/us13/n1079 , \AES_ENC/us13/n1078 , \AES_ENC/us13/n1077 ,\AES_ENC/us13/n1076 , \AES_ENC/us13/n1075 , \AES_ENC/us13/n1074 ,\AES_ENC/us13/n1073 , \AES_ENC/us13/n1072 , \AES_ENC/us13/n1071 ,\AES_ENC/us13/n1070 , \AES_ENC/us13/n1069 , \AES_ENC/us13/n1068 ,\AES_ENC/us13/n1067 , \AES_ENC/us13/n1066 , \AES_ENC/us13/n1065 ,\AES_ENC/us13/n1064 , \AES_ENC/us13/n1063 , \AES_ENC/us13/n1062 ,\AES_ENC/us13/n1061 , \AES_ENC/us13/n1060 , \AES_ENC/us13/n1059 ,\AES_ENC/us13/n1058 , \AES_ENC/us13/n1057 , \AES_ENC/us13/n1056 ,\AES_ENC/us13/n1055 , \AES_ENC/us13/n1054 , \AES_ENC/us13/n1053 ,\AES_ENC/us13/n1052 , \AES_ENC/us13/n1051 , \AES_ENC/us13/n1050 ,\AES_ENC/us13/n1049 , \AES_ENC/us13/n1048 , \AES_ENC/us13/n1047 ,\AES_ENC/us13/n1046 , \AES_ENC/us13/n1045 , \AES_ENC/us13/n1044 ,\AES_ENC/us13/n1043 , \AES_ENC/us13/n1042 , \AES_ENC/us13/n1041 ,\AES_ENC/us13/n1040 , \AES_ENC/us13/n1039 , \AES_ENC/us13/n1038 ,\AES_ENC/us13/n1037 , \AES_ENC/us13/n1036 , \AES_ENC/us13/n1035 ,\AES_ENC/us13/n1034 , \AES_ENC/us13/n1033 , \AES_ENC/us13/n1032 ,\AES_ENC/us13/n1031 , \AES_ENC/us13/n1030 , \AES_ENC/us13/n1029 ,\AES_ENC/us13/n1028 , \AES_ENC/us13/n1027 , \AES_ENC/us13/n1026 ,\AES_ENC/us13/n1025 , \AES_ENC/us13/n1024 , \AES_ENC/us13/n1023 ,\AES_ENC/us13/n1022 , \AES_ENC/us13/n1021 , \AES_ENC/us13/n1020 ,\AES_ENC/us13/n1019 , \AES_ENC/us13/n1018 , \AES_ENC/us13/n1017 ,\AES_ENC/us13/n1016 , \AES_ENC/us13/n1015 , \AES_ENC/us13/n1014 ,\AES_ENC/us13/n1013 , \AES_ENC/us13/n1012 , \AES_ENC/us13/n1011 ,\AES_ENC/us13/n1010 , \AES_ENC/us13/n1009 , \AES_ENC/us13/n1008 ,\AES_ENC/us13/n1007 , \AES_ENC/us13/n1006 , \AES_ENC/us13/n1005 ,\AES_ENC/us13/n1004 , \AES_ENC/us13/n1003 , \AES_ENC/us13/n1002 ,\AES_ENC/us13/n1001 , \AES_ENC/us13/n1000 , \AES_ENC/us13/n999 ,\AES_ENC/us13/n998 , \AES_ENC/us13/n997 , \AES_ENC/us13/n996 ,\AES_ENC/us13/n995 , \AES_ENC/us13/n994 , \AES_ENC/us13/n993 ,\AES_ENC/us13/n992 , \AES_ENC/us13/n991 , \AES_ENC/us13/n990 ,\AES_ENC/us13/n989 , \AES_ENC/us13/n988 , \AES_ENC/us13/n987 ,\AES_ENC/us13/n986 , \AES_ENC/us13/n985 , \AES_ENC/us13/n984 ,\AES_ENC/us13/n983 , \AES_ENC/us13/n982 , \AES_ENC/us13/n981 ,\AES_ENC/us13/n980 , \AES_ENC/us13/n979 , \AES_ENC/us13/n978 ,\AES_ENC/us13/n977 , \AES_ENC/us13/n976 , \AES_ENC/us13/n975 ,\AES_ENC/us13/n974 , \AES_ENC/us13/n973 , \AES_ENC/us13/n972 ,\AES_ENC/us13/n971 , \AES_ENC/us13/n970 , \AES_ENC/us13/n969 ,\AES_ENC/us13/n968 , \AES_ENC/us13/n967 , \AES_ENC/us13/n966 ,\AES_ENC/us13/n965 , \AES_ENC/us13/n964 , \AES_ENC/us13/n963 ,\AES_ENC/us13/n962 , \AES_ENC/us13/n961 , \AES_ENC/us13/n960 ,\AES_ENC/us13/n959 , \AES_ENC/us13/n958 , \AES_ENC/us13/n957 ,\AES_ENC/us13/n956 , \AES_ENC/us13/n955 , \AES_ENC/us13/n954 ,\AES_ENC/us13/n953 , \AES_ENC/us13/n952 , \AES_ENC/us13/n951 ,\AES_ENC/us13/n950 , \AES_ENC/us13/n949 , \AES_ENC/us13/n948 ,\AES_ENC/us13/n947 , \AES_ENC/us13/n946 , \AES_ENC/us13/n945 ,\AES_ENC/us13/n944 , \AES_ENC/us13/n943 , \AES_ENC/us13/n942 ,\AES_ENC/us13/n941 , \AES_ENC/us13/n940 , \AES_ENC/us13/n939 ,\AES_ENC/us13/n938 , \AES_ENC/us13/n937 , \AES_ENC/us13/n936 ,\AES_ENC/us13/n935 , \AES_ENC/us13/n934 , \AES_ENC/us13/n933 ,\AES_ENC/us13/n932 , \AES_ENC/us13/n931 , \AES_ENC/us13/n930 ,\AES_ENC/us13/n929 , \AES_ENC/us13/n928 , \AES_ENC/us13/n927 ,\AES_ENC/us13/n926 , \AES_ENC/us13/n925 , \AES_ENC/us13/n924 ,\AES_ENC/us13/n923 , \AES_ENC/us13/n922 , \AES_ENC/us13/n921 ,\AES_ENC/us13/n920 , \AES_ENC/us13/n919 , \AES_ENC/us13/n918 ,\AES_ENC/us13/n917 , \AES_ENC/us13/n916 , \AES_ENC/us13/n915 ,\AES_ENC/us13/n914 , \AES_ENC/us13/n913 , \AES_ENC/us13/n912 ,\AES_ENC/us13/n911 , \AES_ENC/us13/n910 , \AES_ENC/us13/n909 ,\AES_ENC/us13/n908 , \AES_ENC/us13/n907 , \AES_ENC/us13/n906 ,\AES_ENC/us13/n905 , \AES_ENC/us13/n904 , \AES_ENC/us13/n903 ,\AES_ENC/us13/n902 , \AES_ENC/us13/n901 , \AES_ENC/us13/n900 ,\AES_ENC/us13/n899 , \AES_ENC/us13/n898 , \AES_ENC/us13/n897 ,\AES_ENC/us13/n896 , \AES_ENC/us13/n895 , \AES_ENC/us13/n894 ,\AES_ENC/us13/n893 , \AES_ENC/us13/n892 , \AES_ENC/us13/n891 ,\AES_ENC/us13/n890 , \AES_ENC/us13/n889 , \AES_ENC/us13/n888 ,\AES_ENC/us13/n887 , \AES_ENC/us13/n886 , \AES_ENC/us13/n885 ,\AES_ENC/us13/n884 , \AES_ENC/us13/n883 , \AES_ENC/us13/n882 ,\AES_ENC/us13/n881 , \AES_ENC/us13/n880 , \AES_ENC/us13/n879 ,\AES_ENC/us13/n878 , \AES_ENC/us13/n877 , \AES_ENC/us13/n876 ,\AES_ENC/us13/n875 , \AES_ENC/us13/n874 , \AES_ENC/us13/n873 ,\AES_ENC/us13/n872 , \AES_ENC/us13/n871 , \AES_ENC/us13/n870 ,\AES_ENC/us13/n869 , \AES_ENC/us13/n868 , \AES_ENC/us13/n867 ,\AES_ENC/us13/n866 , \AES_ENC/us13/n865 , \AES_ENC/us13/n864 ,\AES_ENC/us13/n863 , \AES_ENC/us13/n862 , \AES_ENC/us13/n861 ,\AES_ENC/us13/n860 , \AES_ENC/us13/n859 , \AES_ENC/us13/n858 ,\AES_ENC/us13/n857 , \AES_ENC/us13/n856 , \AES_ENC/us13/n855 ,\AES_ENC/us13/n854 , \AES_ENC/us13/n853 , \AES_ENC/us13/n852 ,\AES_ENC/us13/n851 , \AES_ENC/us13/n850 , \AES_ENC/us13/n849 ,\AES_ENC/us13/n848 , \AES_ENC/us13/n847 , \AES_ENC/us13/n846 ,\AES_ENC/us13/n845 , \AES_ENC/us13/n844 , \AES_ENC/us13/n843 ,\AES_ENC/us13/n842 , \AES_ENC/us13/n841 , \AES_ENC/us13/n840 ,\AES_ENC/us13/n839 , \AES_ENC/us13/n838 , \AES_ENC/us13/n837 ,\AES_ENC/us13/n836 , \AES_ENC/us13/n835 , \AES_ENC/us13/n834 ,\AES_ENC/us13/n833 , \AES_ENC/us13/n832 , \AES_ENC/us13/n831 ,\AES_ENC/us13/n830 , \AES_ENC/us13/n829 , \AES_ENC/us13/n828 ,\AES_ENC/us13/n827 , \AES_ENC/us13/n826 , \AES_ENC/us13/n825 ,\AES_ENC/us13/n824 , \AES_ENC/us13/n823 , \AES_ENC/us13/n822 ,\AES_ENC/us13/n821 , \AES_ENC/us13/n820 , \AES_ENC/us13/n819 ,\AES_ENC/us13/n818 , \AES_ENC/us13/n817 , \AES_ENC/us13/n816 ,\AES_ENC/us13/n815 , \AES_ENC/us13/n814 , \AES_ENC/us13/n813 ,\AES_ENC/us13/n812 , \AES_ENC/us13/n811 , \AES_ENC/us13/n810 ,\AES_ENC/us13/n809 , \AES_ENC/us13/n808 , \AES_ENC/us13/n807 ,\AES_ENC/us13/n806 , \AES_ENC/us13/n805 , \AES_ENC/us13/n804 ,\AES_ENC/us13/n803 , \AES_ENC/us13/n802 , \AES_ENC/us13/n801 ,\AES_ENC/us13/n800 , \AES_ENC/us13/n799 , \AES_ENC/us13/n798 ,\AES_ENC/us13/n797 , \AES_ENC/us13/n796 , \AES_ENC/us13/n795 ,\AES_ENC/us13/n794 , \AES_ENC/us13/n793 , \AES_ENC/us13/n792 ,\AES_ENC/us13/n791 , \AES_ENC/us13/n790 , \AES_ENC/us13/n789 ,\AES_ENC/us13/n788 , \AES_ENC/us13/n787 , \AES_ENC/us13/n786 ,\AES_ENC/us13/n785 , \AES_ENC/us13/n784 , \AES_ENC/us13/n783 ,\AES_ENC/us13/n782 , \AES_ENC/us13/n781 , \AES_ENC/us13/n780 ,\AES_ENC/us13/n779 , \AES_ENC/us13/n778 , \AES_ENC/us13/n777 ,\AES_ENC/us13/n776 , \AES_ENC/us13/n775 , \AES_ENC/us13/n774 ,\AES_ENC/us13/n773 , \AES_ENC/us13/n772 , \AES_ENC/us13/n771 ,\AES_ENC/us13/n770 , \AES_ENC/us13/n769 , \AES_ENC/us13/n768 ,\AES_ENC/us13/n767 , \AES_ENC/us13/n766 , \AES_ENC/us13/n765 ,\AES_ENC/us13/n764 , \AES_ENC/us13/n763 , \AES_ENC/us13/n762 ,\AES_ENC/us13/n761 , \AES_ENC/us13/n760 , \AES_ENC/us13/n759 ,\AES_ENC/us13/n758 , \AES_ENC/us13/n757 , \AES_ENC/us13/n756 ,\AES_ENC/us13/n755 , \AES_ENC/us13/n754 , \AES_ENC/us13/n753 ,\AES_ENC/us13/n752 , \AES_ENC/us13/n751 , \AES_ENC/us13/n750 ,\AES_ENC/us13/n749 , \AES_ENC/us13/n748 , \AES_ENC/us13/n747 ,\AES_ENC/us13/n746 , \AES_ENC/us13/n745 , \AES_ENC/us13/n744 ,\AES_ENC/us13/n743 , \AES_ENC/us13/n742 , \AES_ENC/us13/n741 ,\AES_ENC/us13/n740 , \AES_ENC/us13/n739 , \AES_ENC/us13/n738 ,\AES_ENC/us13/n737 , \AES_ENC/us13/n736 , \AES_ENC/us13/n735 ,\AES_ENC/us13/n734 , \AES_ENC/us13/n733 , \AES_ENC/us13/n732 ,\AES_ENC/us13/n731 , \AES_ENC/us13/n730 , \AES_ENC/us13/n729 ,\AES_ENC/us13/n728 , \AES_ENC/us13/n727 , \AES_ENC/us13/n726 ,\AES_ENC/us13/n725 , \AES_ENC/us13/n724 , \AES_ENC/us13/n723 ,\AES_ENC/us13/n722 , \AES_ENC/us13/n721 , \AES_ENC/us13/n720 ,\AES_ENC/us13/n719 , \AES_ENC/us13/n718 , \AES_ENC/us13/n717 ,\AES_ENC/us13/n716 , \AES_ENC/us13/n715 , \AES_ENC/us13/n714 ,\AES_ENC/us13/n713 , \AES_ENC/us13/n712 , \AES_ENC/us13/n711 ,\AES_ENC/us13/n710 , \AES_ENC/us13/n709 , \AES_ENC/us13/n708 ,\AES_ENC/us13/n707 , \AES_ENC/us13/n706 , \AES_ENC/us13/n705 ,\AES_ENC/us13/n704 , \AES_ENC/us13/n703 , \AES_ENC/us13/n702 ,\AES_ENC/us13/n701 , \AES_ENC/us13/n700 , \AES_ENC/us13/n699 ,\AES_ENC/us13/n698 , \AES_ENC/us13/n697 , \AES_ENC/us13/n696 ,\AES_ENC/us13/n695 , \AES_ENC/us13/n694 , \AES_ENC/us13/n693 ,\AES_ENC/us13/n692 , \AES_ENC/us13/n691 , \AES_ENC/us13/n690 ,\AES_ENC/us13/n689 , \AES_ENC/us13/n688 , \AES_ENC/us13/n687 ,\AES_ENC/us13/n686 , \AES_ENC/us13/n685 , \AES_ENC/us13/n684 ,\AES_ENC/us13/n683 , \AES_ENC/us13/n682 , \AES_ENC/us13/n681 ,\AES_ENC/us13/n680 , \AES_ENC/us13/n679 , \AES_ENC/us13/n678 ,\AES_ENC/us13/n677 , \AES_ENC/us13/n676 , \AES_ENC/us13/n675 ,\AES_ENC/us13/n674 , \AES_ENC/us13/n673 , \AES_ENC/us13/n672 ,\AES_ENC/us13/n671 , \AES_ENC/us13/n670 , \AES_ENC/us13/n669 ,\AES_ENC/us13/n668 , \AES_ENC/us13/n667 , \AES_ENC/us13/n666 ,\AES_ENC/us13/n665 , \AES_ENC/us13/n664 , \AES_ENC/us13/n663 ,\AES_ENC/us13/n662 , \AES_ENC/us13/n661 , \AES_ENC/us13/n660 ,\AES_ENC/us13/n659 , \AES_ENC/us13/n658 , \AES_ENC/us13/n657 ,\AES_ENC/us13/n656 , \AES_ENC/us13/n655 , \AES_ENC/us13/n654 ,\AES_ENC/us13/n653 , \AES_ENC/us13/n652 , \AES_ENC/us13/n651 ,\AES_ENC/us13/n650 , \AES_ENC/us13/n649 , \AES_ENC/us13/n648 ,\AES_ENC/us13/n647 , \AES_ENC/us13/n646 , \AES_ENC/us13/n645 ,\AES_ENC/us13/n644 , \AES_ENC/us13/n643 , \AES_ENC/us13/n642 ,\AES_ENC/us13/n641 , \AES_ENC/us13/n640 , \AES_ENC/us13/n639 ,\AES_ENC/us13/n638 , \AES_ENC/us13/n637 , \AES_ENC/us13/n636 ,\AES_ENC/us13/n635 , \AES_ENC/us13/n634 , \AES_ENC/us13/n633 ,\AES_ENC/us13/n632 , \AES_ENC/us13/n631 , \AES_ENC/us13/n630 ,\AES_ENC/us13/n629 , \AES_ENC/us13/n628 , \AES_ENC/us13/n627 ,\AES_ENC/us13/n626 , \AES_ENC/us13/n625 , \AES_ENC/us13/n624 ,\AES_ENC/us13/n623 , \AES_ENC/us13/n622 , \AES_ENC/us13/n621 ,\AES_ENC/us13/n620 , \AES_ENC/us13/n619 , \AES_ENC/us13/n618 ,\AES_ENC/us13/n617 , \AES_ENC/us13/n616 , \AES_ENC/us13/n615 ,\AES_ENC/us13/n614 , \AES_ENC/us13/n613 , \AES_ENC/us13/n612 ,\AES_ENC/us13/n611 , \AES_ENC/us13/n610 , \AES_ENC/us13/n609 ,\AES_ENC/us13/n608 , \AES_ENC/us13/n607 , \AES_ENC/us13/n606 ,\AES_ENC/us13/n605 , \AES_ENC/us13/n604 , \AES_ENC/us13/n603 ,\AES_ENC/us13/n602 , \AES_ENC/us13/n601 , \AES_ENC/us13/n600 ,\AES_ENC/us13/n599 , \AES_ENC/us13/n598 , \AES_ENC/us13/n597 ,\AES_ENC/us13/n596 , \AES_ENC/us13/n595 , \AES_ENC/us13/n594 ,\AES_ENC/us13/n593 , \AES_ENC/us13/n592 , \AES_ENC/us13/n591 ,\AES_ENC/us13/n590 , \AES_ENC/us13/n589 , \AES_ENC/us13/n588 ,\AES_ENC/us13/n587 , \AES_ENC/us13/n586 , \AES_ENC/us13/n585 ,\AES_ENC/us13/n584 , \AES_ENC/us13/n583 , \AES_ENC/us13/n582 ,\AES_ENC/us13/n581 , \AES_ENC/us13/n580 , \AES_ENC/us13/n579 ,\AES_ENC/us13/n578 , \AES_ENC/us13/n577 , \AES_ENC/us13/n576 ,\AES_ENC/us13/n575 , \AES_ENC/us13/n574 , \AES_ENC/us13/n573 ,\AES_ENC/us13/n572 , \AES_ENC/us13/n571 , \AES_ENC/us13/n570 ,\AES_ENC/us13/n569 , \AES_ENC/us20/n1135 , \AES_ENC/us20/n1134 ,\AES_ENC/us20/n1133 , \AES_ENC/us20/n1132 , \AES_ENC/us20/n1131 ,\AES_ENC/us20/n1130 , \AES_ENC/us20/n1129 , \AES_ENC/us20/n1128 ,\AES_ENC/us20/n1127 , \AES_ENC/us20/n1126 , \AES_ENC/us20/n1125 ,\AES_ENC/us20/n1124 , \AES_ENC/us20/n1123 , \AES_ENC/us20/n1122 ,\AES_ENC/us20/n1121 , \AES_ENC/us20/n1120 , \AES_ENC/us20/n1119 ,\AES_ENC/us20/n1118 , \AES_ENC/us20/n1117 , \AES_ENC/us20/n1116 ,\AES_ENC/us20/n1115 , \AES_ENC/us20/n1114 , \AES_ENC/us20/n1113 ,\AES_ENC/us20/n1112 , \AES_ENC/us20/n1111 , \AES_ENC/us20/n1110 ,\AES_ENC/us20/n1109 , \AES_ENC/us20/n1108 , \AES_ENC/us20/n1107 ,\AES_ENC/us20/n1106 , \AES_ENC/us20/n1105 , \AES_ENC/us20/n1104 ,\AES_ENC/us20/n1103 , \AES_ENC/us20/n1102 , \AES_ENC/us20/n1101 ,\AES_ENC/us20/n1100 , \AES_ENC/us20/n1099 , \AES_ENC/us20/n1098 ,\AES_ENC/us20/n1097 , \AES_ENC/us20/n1096 , \AES_ENC/us20/n1095 ,\AES_ENC/us20/n1094 , \AES_ENC/us20/n1093 , \AES_ENC/us20/n1092 ,\AES_ENC/us20/n1091 , \AES_ENC/us20/n1090 , \AES_ENC/us20/n1089 ,\AES_ENC/us20/n1088 , \AES_ENC/us20/n1087 , \AES_ENC/us20/n1086 ,\AES_ENC/us20/n1085 , \AES_ENC/us20/n1084 , \AES_ENC/us20/n1083 ,\AES_ENC/us20/n1082 , \AES_ENC/us20/n1081 , \AES_ENC/us20/n1080 ,\AES_ENC/us20/n1079 , \AES_ENC/us20/n1078 , \AES_ENC/us20/n1077 ,\AES_ENC/us20/n1076 , \AES_ENC/us20/n1075 , \AES_ENC/us20/n1074 ,\AES_ENC/us20/n1073 , \AES_ENC/us20/n1072 , \AES_ENC/us20/n1071 ,\AES_ENC/us20/n1070 , \AES_ENC/us20/n1069 , \AES_ENC/us20/n1068 ,\AES_ENC/us20/n1067 , \AES_ENC/us20/n1066 , \AES_ENC/us20/n1065 ,\AES_ENC/us20/n1064 , \AES_ENC/us20/n1063 , \AES_ENC/us20/n1062 ,\AES_ENC/us20/n1061 , \AES_ENC/us20/n1060 , \AES_ENC/us20/n1059 ,\AES_ENC/us20/n1058 , \AES_ENC/us20/n1057 , \AES_ENC/us20/n1056 ,\AES_ENC/us20/n1055 , \AES_ENC/us20/n1054 , \AES_ENC/us20/n1053 ,\AES_ENC/us20/n1052 , \AES_ENC/us20/n1051 , \AES_ENC/us20/n1050 ,\AES_ENC/us20/n1049 , \AES_ENC/us20/n1048 , \AES_ENC/us20/n1047 ,\AES_ENC/us20/n1046 , \AES_ENC/us20/n1045 , \AES_ENC/us20/n1044 ,\AES_ENC/us20/n1043 , \AES_ENC/us20/n1042 , \AES_ENC/us20/n1041 ,\AES_ENC/us20/n1040 , \AES_ENC/us20/n1039 , \AES_ENC/us20/n1038 ,\AES_ENC/us20/n1037 , \AES_ENC/us20/n1036 , \AES_ENC/us20/n1035 ,\AES_ENC/us20/n1034 , \AES_ENC/us20/n1033 , \AES_ENC/us20/n1032 ,\AES_ENC/us20/n1031 , \AES_ENC/us20/n1030 , \AES_ENC/us20/n1029 ,\AES_ENC/us20/n1028 , \AES_ENC/us20/n1027 , \AES_ENC/us20/n1026 ,\AES_ENC/us20/n1025 , \AES_ENC/us20/n1024 , \AES_ENC/us20/n1023 ,\AES_ENC/us20/n1022 , \AES_ENC/us20/n1021 , \AES_ENC/us20/n1020 ,\AES_ENC/us20/n1019 , \AES_ENC/us20/n1018 , \AES_ENC/us20/n1017 ,\AES_ENC/us20/n1016 , \AES_ENC/us20/n1015 , \AES_ENC/us20/n1014 ,\AES_ENC/us20/n1013 , \AES_ENC/us20/n1012 , \AES_ENC/us20/n1011 ,\AES_ENC/us20/n1010 , \AES_ENC/us20/n1009 , \AES_ENC/us20/n1008 ,\AES_ENC/us20/n1007 , \AES_ENC/us20/n1006 , \AES_ENC/us20/n1005 ,\AES_ENC/us20/n1004 , \AES_ENC/us20/n1003 , \AES_ENC/us20/n1002 ,\AES_ENC/us20/n1001 , \AES_ENC/us20/n1000 , \AES_ENC/us20/n999 ,\AES_ENC/us20/n998 , \AES_ENC/us20/n997 , \AES_ENC/us20/n996 ,\AES_ENC/us20/n995 , \AES_ENC/us20/n994 , \AES_ENC/us20/n993 ,\AES_ENC/us20/n992 , \AES_ENC/us20/n991 , \AES_ENC/us20/n990 ,\AES_ENC/us20/n989 , \AES_ENC/us20/n988 , \AES_ENC/us20/n987 ,\AES_ENC/us20/n986 , \AES_ENC/us20/n985 , \AES_ENC/us20/n984 ,\AES_ENC/us20/n983 , \AES_ENC/us20/n982 , \AES_ENC/us20/n981 ,\AES_ENC/us20/n980 , \AES_ENC/us20/n979 , \AES_ENC/us20/n978 ,\AES_ENC/us20/n977 , \AES_ENC/us20/n976 , \AES_ENC/us20/n975 ,\AES_ENC/us20/n974 , \AES_ENC/us20/n973 , \AES_ENC/us20/n972 ,\AES_ENC/us20/n971 , \AES_ENC/us20/n970 , \AES_ENC/us20/n969 ,\AES_ENC/us20/n968 , \AES_ENC/us20/n967 , \AES_ENC/us20/n966 ,\AES_ENC/us20/n965 , \AES_ENC/us20/n964 , \AES_ENC/us20/n963 ,\AES_ENC/us20/n962 , \AES_ENC/us20/n961 , \AES_ENC/us20/n960 ,\AES_ENC/us20/n959 , \AES_ENC/us20/n958 , \AES_ENC/us20/n957 ,\AES_ENC/us20/n956 , \AES_ENC/us20/n955 , \AES_ENC/us20/n954 ,\AES_ENC/us20/n953 , \AES_ENC/us20/n952 , \AES_ENC/us20/n951 ,\AES_ENC/us20/n950 , \AES_ENC/us20/n949 , \AES_ENC/us20/n948 ,\AES_ENC/us20/n947 , \AES_ENC/us20/n946 , \AES_ENC/us20/n945 ,\AES_ENC/us20/n944 , \AES_ENC/us20/n943 , \AES_ENC/us20/n942 ,\AES_ENC/us20/n941 , \AES_ENC/us20/n940 , \AES_ENC/us20/n939 ,\AES_ENC/us20/n938 , \AES_ENC/us20/n937 , \AES_ENC/us20/n936 ,\AES_ENC/us20/n935 , \AES_ENC/us20/n934 , \AES_ENC/us20/n933 ,\AES_ENC/us20/n932 , \AES_ENC/us20/n931 , \AES_ENC/us20/n930 ,\AES_ENC/us20/n929 , \AES_ENC/us20/n928 , \AES_ENC/us20/n927 ,\AES_ENC/us20/n926 , \AES_ENC/us20/n925 , \AES_ENC/us20/n924 ,\AES_ENC/us20/n923 , \AES_ENC/us20/n922 , \AES_ENC/us20/n921 ,\AES_ENC/us20/n920 , \AES_ENC/us20/n919 , \AES_ENC/us20/n918 ,\AES_ENC/us20/n917 , \AES_ENC/us20/n916 , \AES_ENC/us20/n915 ,\AES_ENC/us20/n914 , \AES_ENC/us20/n913 , \AES_ENC/us20/n912 ,\AES_ENC/us20/n911 , \AES_ENC/us20/n910 , \AES_ENC/us20/n909 ,\AES_ENC/us20/n908 , \AES_ENC/us20/n907 , \AES_ENC/us20/n906 ,\AES_ENC/us20/n905 , \AES_ENC/us20/n904 , \AES_ENC/us20/n903 ,\AES_ENC/us20/n902 , \AES_ENC/us20/n901 , \AES_ENC/us20/n900 ,\AES_ENC/us20/n899 , \AES_ENC/us20/n898 , \AES_ENC/us20/n897 ,\AES_ENC/us20/n896 , \AES_ENC/us20/n895 , \AES_ENC/us20/n894 ,\AES_ENC/us20/n893 , \AES_ENC/us20/n892 , \AES_ENC/us20/n891 ,\AES_ENC/us20/n890 , \AES_ENC/us20/n889 , \AES_ENC/us20/n888 ,\AES_ENC/us20/n887 , \AES_ENC/us20/n886 , \AES_ENC/us20/n885 ,\AES_ENC/us20/n884 , \AES_ENC/us20/n883 , \AES_ENC/us20/n882 ,\AES_ENC/us20/n881 , \AES_ENC/us20/n880 , \AES_ENC/us20/n879 ,\AES_ENC/us20/n878 , \AES_ENC/us20/n877 , \AES_ENC/us20/n876 ,\AES_ENC/us20/n875 , \AES_ENC/us20/n874 , \AES_ENC/us20/n873 ,\AES_ENC/us20/n872 , \AES_ENC/us20/n871 , \AES_ENC/us20/n870 ,\AES_ENC/us20/n869 , \AES_ENC/us20/n868 , \AES_ENC/us20/n867 ,\AES_ENC/us20/n866 , \AES_ENC/us20/n865 , \AES_ENC/us20/n864 ,\AES_ENC/us20/n863 , \AES_ENC/us20/n862 , \AES_ENC/us20/n861 ,\AES_ENC/us20/n860 , \AES_ENC/us20/n859 , \AES_ENC/us20/n858 ,\AES_ENC/us20/n857 , \AES_ENC/us20/n856 , \AES_ENC/us20/n855 ,\AES_ENC/us20/n854 , \AES_ENC/us20/n853 , \AES_ENC/us20/n852 ,\AES_ENC/us20/n851 , \AES_ENC/us20/n850 , \AES_ENC/us20/n849 ,\AES_ENC/us20/n848 , \AES_ENC/us20/n847 , \AES_ENC/us20/n846 ,\AES_ENC/us20/n845 , \AES_ENC/us20/n844 , \AES_ENC/us20/n843 ,\AES_ENC/us20/n842 , \AES_ENC/us20/n841 , \AES_ENC/us20/n840 ,\AES_ENC/us20/n839 , \AES_ENC/us20/n838 , \AES_ENC/us20/n837 ,\AES_ENC/us20/n836 , \AES_ENC/us20/n835 , \AES_ENC/us20/n834 ,\AES_ENC/us20/n833 , \AES_ENC/us20/n832 , \AES_ENC/us20/n831 ,\AES_ENC/us20/n830 , \AES_ENC/us20/n829 , \AES_ENC/us20/n828 ,\AES_ENC/us20/n827 , \AES_ENC/us20/n826 , \AES_ENC/us20/n825 ,\AES_ENC/us20/n824 , \AES_ENC/us20/n823 , \AES_ENC/us20/n822 ,\AES_ENC/us20/n821 , \AES_ENC/us20/n820 , \AES_ENC/us20/n819 ,\AES_ENC/us20/n818 , \AES_ENC/us20/n817 , \AES_ENC/us20/n816 ,\AES_ENC/us20/n815 , \AES_ENC/us20/n814 , \AES_ENC/us20/n813 ,\AES_ENC/us20/n812 , \AES_ENC/us20/n811 , \AES_ENC/us20/n810 ,\AES_ENC/us20/n809 , \AES_ENC/us20/n808 , \AES_ENC/us20/n807 ,\AES_ENC/us20/n806 , \AES_ENC/us20/n805 , \AES_ENC/us20/n804 ,\AES_ENC/us20/n803 , \AES_ENC/us20/n802 , \AES_ENC/us20/n801 ,\AES_ENC/us20/n800 , \AES_ENC/us20/n799 , \AES_ENC/us20/n798 ,\AES_ENC/us20/n797 , \AES_ENC/us20/n796 , \AES_ENC/us20/n795 ,\AES_ENC/us20/n794 , \AES_ENC/us20/n793 , \AES_ENC/us20/n792 ,\AES_ENC/us20/n791 , \AES_ENC/us20/n790 , \AES_ENC/us20/n789 ,\AES_ENC/us20/n788 , \AES_ENC/us20/n787 , \AES_ENC/us20/n786 ,\AES_ENC/us20/n785 , \AES_ENC/us20/n784 , \AES_ENC/us20/n783 ,\AES_ENC/us20/n782 , \AES_ENC/us20/n781 , \AES_ENC/us20/n780 ,\AES_ENC/us20/n779 , \AES_ENC/us20/n778 , \AES_ENC/us20/n777 ,\AES_ENC/us20/n776 , \AES_ENC/us20/n775 , \AES_ENC/us20/n774 ,\AES_ENC/us20/n773 , \AES_ENC/us20/n772 , \AES_ENC/us20/n771 ,\AES_ENC/us20/n770 , \AES_ENC/us20/n769 , \AES_ENC/us20/n768 ,\AES_ENC/us20/n767 , \AES_ENC/us20/n766 , \AES_ENC/us20/n765 ,\AES_ENC/us20/n764 , \AES_ENC/us20/n763 , \AES_ENC/us20/n762 ,\AES_ENC/us20/n761 , \AES_ENC/us20/n760 , \AES_ENC/us20/n759 ,\AES_ENC/us20/n758 , \AES_ENC/us20/n757 , \AES_ENC/us20/n756 ,\AES_ENC/us20/n755 , \AES_ENC/us20/n754 , \AES_ENC/us20/n753 ,\AES_ENC/us20/n752 , \AES_ENC/us20/n751 , \AES_ENC/us20/n750 ,\AES_ENC/us20/n749 , \AES_ENC/us20/n748 , \AES_ENC/us20/n747 ,\AES_ENC/us20/n746 , \AES_ENC/us20/n745 , \AES_ENC/us20/n744 ,\AES_ENC/us20/n743 , \AES_ENC/us20/n742 , \AES_ENC/us20/n741 ,\AES_ENC/us20/n740 , \AES_ENC/us20/n739 , \AES_ENC/us20/n738 ,\AES_ENC/us20/n737 , \AES_ENC/us20/n736 , \AES_ENC/us20/n735 ,\AES_ENC/us20/n734 , \AES_ENC/us20/n733 , \AES_ENC/us20/n732 ,\AES_ENC/us20/n731 , \AES_ENC/us20/n730 , \AES_ENC/us20/n729 ,\AES_ENC/us20/n728 , \AES_ENC/us20/n727 , \AES_ENC/us20/n726 ,\AES_ENC/us20/n725 , \AES_ENC/us20/n724 , \AES_ENC/us20/n723 ,\AES_ENC/us20/n722 , \AES_ENC/us20/n721 , \AES_ENC/us20/n720 ,\AES_ENC/us20/n719 , \AES_ENC/us20/n718 , \AES_ENC/us20/n717 ,\AES_ENC/us20/n716 , \AES_ENC/us20/n715 , \AES_ENC/us20/n714 ,\AES_ENC/us20/n713 , \AES_ENC/us20/n712 , \AES_ENC/us20/n711 ,\AES_ENC/us20/n710 , \AES_ENC/us20/n709 , \AES_ENC/us20/n708 ,\AES_ENC/us20/n707 , \AES_ENC/us20/n706 , \AES_ENC/us20/n705 ,\AES_ENC/us20/n704 , \AES_ENC/us20/n703 , \AES_ENC/us20/n702 ,\AES_ENC/us20/n701 , \AES_ENC/us20/n700 , \AES_ENC/us20/n699 ,\AES_ENC/us20/n698 , \AES_ENC/us20/n697 , \AES_ENC/us20/n696 ,\AES_ENC/us20/n695 , \AES_ENC/us20/n694 , \AES_ENC/us20/n693 ,\AES_ENC/us20/n692 , \AES_ENC/us20/n691 , \AES_ENC/us20/n690 ,\AES_ENC/us20/n689 , \AES_ENC/us20/n688 , \AES_ENC/us20/n687 ,\AES_ENC/us20/n686 , \AES_ENC/us20/n685 , \AES_ENC/us20/n684 ,\AES_ENC/us20/n683 , \AES_ENC/us20/n682 , \AES_ENC/us20/n681 ,\AES_ENC/us20/n680 , \AES_ENC/us20/n679 , \AES_ENC/us20/n678 ,\AES_ENC/us20/n677 , \AES_ENC/us20/n676 , \AES_ENC/us20/n675 ,\AES_ENC/us20/n674 , \AES_ENC/us20/n673 , \AES_ENC/us20/n672 ,\AES_ENC/us20/n671 , \AES_ENC/us20/n670 , \AES_ENC/us20/n669 ,\AES_ENC/us20/n668 , \AES_ENC/us20/n667 , \AES_ENC/us20/n666 ,\AES_ENC/us20/n665 , \AES_ENC/us20/n664 , \AES_ENC/us20/n663 ,\AES_ENC/us20/n662 , \AES_ENC/us20/n661 , \AES_ENC/us20/n660 ,\AES_ENC/us20/n659 , \AES_ENC/us20/n658 , \AES_ENC/us20/n657 ,\AES_ENC/us20/n656 , \AES_ENC/us20/n655 , \AES_ENC/us20/n654 ,\AES_ENC/us20/n653 , \AES_ENC/us20/n652 , \AES_ENC/us20/n651 ,\AES_ENC/us20/n650 , \AES_ENC/us20/n649 , \AES_ENC/us20/n648 ,\AES_ENC/us20/n647 , \AES_ENC/us20/n646 , \AES_ENC/us20/n645 ,\AES_ENC/us20/n644 , \AES_ENC/us20/n643 , \AES_ENC/us20/n642 ,\AES_ENC/us20/n641 , \AES_ENC/us20/n640 , \AES_ENC/us20/n639 ,\AES_ENC/us20/n638 , \AES_ENC/us20/n637 , \AES_ENC/us20/n636 ,\AES_ENC/us20/n635 , \AES_ENC/us20/n634 , \AES_ENC/us20/n633 ,\AES_ENC/us20/n632 , \AES_ENC/us20/n631 , \AES_ENC/us20/n630 ,\AES_ENC/us20/n629 , \AES_ENC/us20/n628 , \AES_ENC/us20/n627 ,\AES_ENC/us20/n626 , \AES_ENC/us20/n625 , \AES_ENC/us20/n624 ,\AES_ENC/us20/n623 , \AES_ENC/us20/n622 , \AES_ENC/us20/n621 ,\AES_ENC/us20/n620 , \AES_ENC/us20/n619 , \AES_ENC/us20/n618 ,\AES_ENC/us20/n617 , \AES_ENC/us20/n616 , \AES_ENC/us20/n615 ,\AES_ENC/us20/n614 , \AES_ENC/us20/n613 , \AES_ENC/us20/n612 ,\AES_ENC/us20/n611 , \AES_ENC/us20/n610 , \AES_ENC/us20/n609 ,\AES_ENC/us20/n608 , \AES_ENC/us20/n607 , \AES_ENC/us20/n606 ,\AES_ENC/us20/n605 , \AES_ENC/us20/n604 , \AES_ENC/us20/n603 ,\AES_ENC/us20/n602 , \AES_ENC/us20/n601 , \AES_ENC/us20/n600 ,\AES_ENC/us20/n599 , \AES_ENC/us20/n598 , \AES_ENC/us20/n597 ,\AES_ENC/us20/n596 , \AES_ENC/us20/n595 , \AES_ENC/us20/n594 ,\AES_ENC/us20/n593 , \AES_ENC/us20/n592 , \AES_ENC/us20/n591 ,\AES_ENC/us20/n590 , \AES_ENC/us20/n589 , \AES_ENC/us20/n588 ,\AES_ENC/us20/n587 , \AES_ENC/us20/n586 , \AES_ENC/us20/n585 ,\AES_ENC/us20/n584 , \AES_ENC/us20/n583 , \AES_ENC/us20/n582 ,\AES_ENC/us20/n581 , \AES_ENC/us20/n580 , \AES_ENC/us20/n579 ,\AES_ENC/us20/n578 , \AES_ENC/us20/n577 , \AES_ENC/us20/n576 ,\AES_ENC/us20/n575 , \AES_ENC/us20/n574 , \AES_ENC/us20/n573 ,\AES_ENC/us20/n572 , \AES_ENC/us20/n571 , \AES_ENC/us20/n570 ,\AES_ENC/us20/n569 , \AES_ENC/us21/n1135 , \AES_ENC/us21/n1134 ,\AES_ENC/us21/n1133 , \AES_ENC/us21/n1132 , \AES_ENC/us21/n1131 ,\AES_ENC/us21/n1130 , \AES_ENC/us21/n1129 , \AES_ENC/us21/n1128 ,\AES_ENC/us21/n1127 , \AES_ENC/us21/n1126 , \AES_ENC/us21/n1125 ,\AES_ENC/us21/n1124 , \AES_ENC/us21/n1123 , \AES_ENC/us21/n1122 ,\AES_ENC/us21/n1121 , \AES_ENC/us21/n1120 , \AES_ENC/us21/n1119 ,\AES_ENC/us21/n1118 , \AES_ENC/us21/n1117 , \AES_ENC/us21/n1116 ,\AES_ENC/us21/n1115 , \AES_ENC/us21/n1114 , \AES_ENC/us21/n1113 ,\AES_ENC/us21/n1112 , \AES_ENC/us21/n1111 , \AES_ENC/us21/n1110 ,\AES_ENC/us21/n1109 , \AES_ENC/us21/n1108 , \AES_ENC/us21/n1107 ,\AES_ENC/us21/n1106 , \AES_ENC/us21/n1105 , \AES_ENC/us21/n1104 ,\AES_ENC/us21/n1103 , \AES_ENC/us21/n1102 , \AES_ENC/us21/n1101 ,\AES_ENC/us21/n1100 , \AES_ENC/us21/n1099 , \AES_ENC/us21/n1098 ,\AES_ENC/us21/n1097 , \AES_ENC/us21/n1096 , \AES_ENC/us21/n1095 ,\AES_ENC/us21/n1094 , \AES_ENC/us21/n1093 , \AES_ENC/us21/n1092 ,\AES_ENC/us21/n1091 , \AES_ENC/us21/n1090 , \AES_ENC/us21/n1089 ,\AES_ENC/us21/n1088 , \AES_ENC/us21/n1087 , \AES_ENC/us21/n1086 ,\AES_ENC/us21/n1085 , \AES_ENC/us21/n1084 , \AES_ENC/us21/n1083 ,\AES_ENC/us21/n1082 , \AES_ENC/us21/n1081 , \AES_ENC/us21/n1080 ,\AES_ENC/us21/n1079 , \AES_ENC/us21/n1078 , \AES_ENC/us21/n1077 ,\AES_ENC/us21/n1076 , \AES_ENC/us21/n1075 , \AES_ENC/us21/n1074 ,\AES_ENC/us21/n1073 , \AES_ENC/us21/n1072 , \AES_ENC/us21/n1071 ,\AES_ENC/us21/n1070 , \AES_ENC/us21/n1069 , \AES_ENC/us21/n1068 ,\AES_ENC/us21/n1067 , \AES_ENC/us21/n1066 , \AES_ENC/us21/n1065 ,\AES_ENC/us21/n1064 , \AES_ENC/us21/n1063 , \AES_ENC/us21/n1062 ,\AES_ENC/us21/n1061 , \AES_ENC/us21/n1060 , \AES_ENC/us21/n1059 ,\AES_ENC/us21/n1058 , \AES_ENC/us21/n1057 , \AES_ENC/us21/n1056 ,\AES_ENC/us21/n1055 , \AES_ENC/us21/n1054 , \AES_ENC/us21/n1053 ,\AES_ENC/us21/n1052 , \AES_ENC/us21/n1051 , \AES_ENC/us21/n1050 ,\AES_ENC/us21/n1049 , \AES_ENC/us21/n1048 , \AES_ENC/us21/n1047 ,\AES_ENC/us21/n1046 , \AES_ENC/us21/n1045 , \AES_ENC/us21/n1044 ,\AES_ENC/us21/n1043 , \AES_ENC/us21/n1042 , \AES_ENC/us21/n1041 ,\AES_ENC/us21/n1040 , \AES_ENC/us21/n1039 , \AES_ENC/us21/n1038 ,\AES_ENC/us21/n1037 , \AES_ENC/us21/n1036 , \AES_ENC/us21/n1035 ,\AES_ENC/us21/n1034 , \AES_ENC/us21/n1033 , \AES_ENC/us21/n1032 ,\AES_ENC/us21/n1031 , \AES_ENC/us21/n1030 , \AES_ENC/us21/n1029 ,\AES_ENC/us21/n1028 , \AES_ENC/us21/n1027 , \AES_ENC/us21/n1026 ,\AES_ENC/us21/n1025 , \AES_ENC/us21/n1024 , \AES_ENC/us21/n1023 ,\AES_ENC/us21/n1022 , \AES_ENC/us21/n1021 , \AES_ENC/us21/n1020 ,\AES_ENC/us21/n1019 , \AES_ENC/us21/n1018 , \AES_ENC/us21/n1017 ,\AES_ENC/us21/n1016 , \AES_ENC/us21/n1015 , \AES_ENC/us21/n1014 ,\AES_ENC/us21/n1013 , \AES_ENC/us21/n1012 , \AES_ENC/us21/n1011 ,\AES_ENC/us21/n1010 , \AES_ENC/us21/n1009 , \AES_ENC/us21/n1008 ,\AES_ENC/us21/n1007 , \AES_ENC/us21/n1006 , \AES_ENC/us21/n1005 ,\AES_ENC/us21/n1004 , \AES_ENC/us21/n1003 , \AES_ENC/us21/n1002 ,\AES_ENC/us21/n1001 , \AES_ENC/us21/n1000 , \AES_ENC/us21/n999 ,\AES_ENC/us21/n998 , \AES_ENC/us21/n997 , \AES_ENC/us21/n996 ,\AES_ENC/us21/n995 , \AES_ENC/us21/n994 , \AES_ENC/us21/n993 ,\AES_ENC/us21/n992 , \AES_ENC/us21/n991 , \AES_ENC/us21/n990 ,\AES_ENC/us21/n989 , \AES_ENC/us21/n988 , \AES_ENC/us21/n987 ,\AES_ENC/us21/n986 , \AES_ENC/us21/n985 , \AES_ENC/us21/n984 ,\AES_ENC/us21/n983 , \AES_ENC/us21/n982 , \AES_ENC/us21/n981 ,\AES_ENC/us21/n980 , \AES_ENC/us21/n979 , \AES_ENC/us21/n978 ,\AES_ENC/us21/n977 , \AES_ENC/us21/n976 , \AES_ENC/us21/n975 ,\AES_ENC/us21/n974 , \AES_ENC/us21/n973 , \AES_ENC/us21/n972 ,\AES_ENC/us21/n971 , \AES_ENC/us21/n970 , \AES_ENC/us21/n969 ,\AES_ENC/us21/n968 , \AES_ENC/us21/n967 , \AES_ENC/us21/n966 ,\AES_ENC/us21/n965 , \AES_ENC/us21/n964 , \AES_ENC/us21/n963 ,\AES_ENC/us21/n962 , \AES_ENC/us21/n961 , \AES_ENC/us21/n960 ,\AES_ENC/us21/n959 , \AES_ENC/us21/n958 , \AES_ENC/us21/n957 ,\AES_ENC/us21/n956 , \AES_ENC/us21/n955 , \AES_ENC/us21/n954 ,\AES_ENC/us21/n953 , \AES_ENC/us21/n952 , \AES_ENC/us21/n951 ,\AES_ENC/us21/n950 , \AES_ENC/us21/n949 , \AES_ENC/us21/n948 ,\AES_ENC/us21/n947 , \AES_ENC/us21/n946 , \AES_ENC/us21/n945 ,\AES_ENC/us21/n944 , \AES_ENC/us21/n943 , \AES_ENC/us21/n942 ,\AES_ENC/us21/n941 , \AES_ENC/us21/n940 , \AES_ENC/us21/n939 ,\AES_ENC/us21/n938 , \AES_ENC/us21/n937 , \AES_ENC/us21/n936 ,\AES_ENC/us21/n935 , \AES_ENC/us21/n934 , \AES_ENC/us21/n933 ,\AES_ENC/us21/n932 , \AES_ENC/us21/n931 , \AES_ENC/us21/n930 ,\AES_ENC/us21/n929 , \AES_ENC/us21/n928 , \AES_ENC/us21/n927 ,\AES_ENC/us21/n926 , \AES_ENC/us21/n925 , \AES_ENC/us21/n924 ,\AES_ENC/us21/n923 , \AES_ENC/us21/n922 , \AES_ENC/us21/n921 ,\AES_ENC/us21/n920 , \AES_ENC/us21/n919 , \AES_ENC/us21/n918 ,\AES_ENC/us21/n917 , \AES_ENC/us21/n916 , \AES_ENC/us21/n915 ,\AES_ENC/us21/n914 , \AES_ENC/us21/n913 , \AES_ENC/us21/n912 ,\AES_ENC/us21/n911 , \AES_ENC/us21/n910 , \AES_ENC/us21/n909 ,\AES_ENC/us21/n908 , \AES_ENC/us21/n907 , \AES_ENC/us21/n906 ,\AES_ENC/us21/n905 , \AES_ENC/us21/n904 , \AES_ENC/us21/n903 ,\AES_ENC/us21/n902 , \AES_ENC/us21/n901 , \AES_ENC/us21/n900 ,\AES_ENC/us21/n899 , \AES_ENC/us21/n898 , \AES_ENC/us21/n897 ,\AES_ENC/us21/n896 , \AES_ENC/us21/n895 , \AES_ENC/us21/n894 ,\AES_ENC/us21/n893 , \AES_ENC/us21/n892 , \AES_ENC/us21/n891 ,\AES_ENC/us21/n890 , \AES_ENC/us21/n889 , \AES_ENC/us21/n888 ,\AES_ENC/us21/n887 , \AES_ENC/us21/n886 , \AES_ENC/us21/n885 ,\AES_ENC/us21/n884 , \AES_ENC/us21/n883 , \AES_ENC/us21/n882 ,\AES_ENC/us21/n881 , \AES_ENC/us21/n880 , \AES_ENC/us21/n879 ,\AES_ENC/us21/n878 , \AES_ENC/us21/n877 , \AES_ENC/us21/n876 ,\AES_ENC/us21/n875 , \AES_ENC/us21/n874 , \AES_ENC/us21/n873 ,\AES_ENC/us21/n872 , \AES_ENC/us21/n871 , \AES_ENC/us21/n870 ,\AES_ENC/us21/n869 , \AES_ENC/us21/n868 , \AES_ENC/us21/n867 ,\AES_ENC/us21/n866 , \AES_ENC/us21/n865 , \AES_ENC/us21/n864 ,\AES_ENC/us21/n863 , \AES_ENC/us21/n862 , \AES_ENC/us21/n861 ,\AES_ENC/us21/n860 , \AES_ENC/us21/n859 , \AES_ENC/us21/n858 ,\AES_ENC/us21/n857 , \AES_ENC/us21/n856 , \AES_ENC/us21/n855 ,\AES_ENC/us21/n854 , \AES_ENC/us21/n853 , \AES_ENC/us21/n852 ,\AES_ENC/us21/n851 , \AES_ENC/us21/n850 , \AES_ENC/us21/n849 ,\AES_ENC/us21/n848 , \AES_ENC/us21/n847 , \AES_ENC/us21/n846 ,\AES_ENC/us21/n845 , \AES_ENC/us21/n844 , \AES_ENC/us21/n843 ,\AES_ENC/us21/n842 , \AES_ENC/us21/n841 , \AES_ENC/us21/n840 ,\AES_ENC/us21/n839 , \AES_ENC/us21/n838 , \AES_ENC/us21/n837 ,\AES_ENC/us21/n836 , \AES_ENC/us21/n835 , \AES_ENC/us21/n834 ,\AES_ENC/us21/n833 , \AES_ENC/us21/n832 , \AES_ENC/us21/n831 ,\AES_ENC/us21/n830 , \AES_ENC/us21/n829 , \AES_ENC/us21/n828 ,\AES_ENC/us21/n827 , \AES_ENC/us21/n826 , \AES_ENC/us21/n825 ,\AES_ENC/us21/n824 , \AES_ENC/us21/n823 , \AES_ENC/us21/n822 ,\AES_ENC/us21/n821 , \AES_ENC/us21/n820 , \AES_ENC/us21/n819 ,\AES_ENC/us21/n818 , \AES_ENC/us21/n817 , \AES_ENC/us21/n816 ,\AES_ENC/us21/n815 , \AES_ENC/us21/n814 , \AES_ENC/us21/n813 ,\AES_ENC/us21/n812 , \AES_ENC/us21/n811 , \AES_ENC/us21/n810 ,\AES_ENC/us21/n809 , \AES_ENC/us21/n808 , \AES_ENC/us21/n807 ,\AES_ENC/us21/n806 , \AES_ENC/us21/n805 , \AES_ENC/us21/n804 ,\AES_ENC/us21/n803 , \AES_ENC/us21/n802 , \AES_ENC/us21/n801 ,\AES_ENC/us21/n800 , \AES_ENC/us21/n799 , \AES_ENC/us21/n798 ,\AES_ENC/us21/n797 , \AES_ENC/us21/n796 , \AES_ENC/us21/n795 ,\AES_ENC/us21/n794 , \AES_ENC/us21/n793 , \AES_ENC/us21/n792 ,\AES_ENC/us21/n791 , \AES_ENC/us21/n790 , \AES_ENC/us21/n789 ,\AES_ENC/us21/n788 , \AES_ENC/us21/n787 , \AES_ENC/us21/n786 ,\AES_ENC/us21/n785 , \AES_ENC/us21/n784 , \AES_ENC/us21/n783 ,\AES_ENC/us21/n782 , \AES_ENC/us21/n781 , \AES_ENC/us21/n780 ,\AES_ENC/us21/n779 , \AES_ENC/us21/n778 , \AES_ENC/us21/n777 ,\AES_ENC/us21/n776 , \AES_ENC/us21/n775 , \AES_ENC/us21/n774 ,\AES_ENC/us21/n773 , \AES_ENC/us21/n772 , \AES_ENC/us21/n771 ,\AES_ENC/us21/n770 , \AES_ENC/us21/n769 , \AES_ENC/us21/n768 ,\AES_ENC/us21/n767 , \AES_ENC/us21/n766 , \AES_ENC/us21/n765 ,\AES_ENC/us21/n764 , \AES_ENC/us21/n763 , \AES_ENC/us21/n762 ,\AES_ENC/us21/n761 , \AES_ENC/us21/n760 , \AES_ENC/us21/n759 ,\AES_ENC/us21/n758 , \AES_ENC/us21/n757 , \AES_ENC/us21/n756 ,\AES_ENC/us21/n755 , \AES_ENC/us21/n754 , \AES_ENC/us21/n753 ,\AES_ENC/us21/n752 , \AES_ENC/us21/n751 , \AES_ENC/us21/n750 ,\AES_ENC/us21/n749 , \AES_ENC/us21/n748 , \AES_ENC/us21/n747 ,\AES_ENC/us21/n746 , \AES_ENC/us21/n745 , \AES_ENC/us21/n744 ,\AES_ENC/us21/n743 , \AES_ENC/us21/n742 , \AES_ENC/us21/n741 ,\AES_ENC/us21/n740 , \AES_ENC/us21/n739 , \AES_ENC/us21/n738 ,\AES_ENC/us21/n737 , \AES_ENC/us21/n736 , \AES_ENC/us21/n735 ,\AES_ENC/us21/n734 , \AES_ENC/us21/n733 , \AES_ENC/us21/n732 ,\AES_ENC/us21/n731 , \AES_ENC/us21/n730 , \AES_ENC/us21/n729 ,\AES_ENC/us21/n728 , \AES_ENC/us21/n727 , \AES_ENC/us21/n726 ,\AES_ENC/us21/n725 , \AES_ENC/us21/n724 , \AES_ENC/us21/n723 ,\AES_ENC/us21/n722 , \AES_ENC/us21/n721 , \AES_ENC/us21/n720 ,\AES_ENC/us21/n719 , \AES_ENC/us21/n718 , \AES_ENC/us21/n717 ,\AES_ENC/us21/n716 , \AES_ENC/us21/n715 , \AES_ENC/us21/n714 ,\AES_ENC/us21/n713 , \AES_ENC/us21/n712 , \AES_ENC/us21/n711 ,\AES_ENC/us21/n710 , \AES_ENC/us21/n709 , \AES_ENC/us21/n708 ,\AES_ENC/us21/n707 , \AES_ENC/us21/n706 , \AES_ENC/us21/n705 ,\AES_ENC/us21/n704 , \AES_ENC/us21/n703 , \AES_ENC/us21/n702 ,\AES_ENC/us21/n701 , \AES_ENC/us21/n700 , \AES_ENC/us21/n699 ,\AES_ENC/us21/n698 , \AES_ENC/us21/n697 , \AES_ENC/us21/n696 ,\AES_ENC/us21/n695 , \AES_ENC/us21/n694 , \AES_ENC/us21/n693 ,\AES_ENC/us21/n692 , \AES_ENC/us21/n691 , \AES_ENC/us21/n690 ,\AES_ENC/us21/n689 , \AES_ENC/us21/n688 , \AES_ENC/us21/n687 ,\AES_ENC/us21/n686 , \AES_ENC/us21/n685 , \AES_ENC/us21/n684 ,\AES_ENC/us21/n683 , \AES_ENC/us21/n682 , \AES_ENC/us21/n681 ,\AES_ENC/us21/n680 , \AES_ENC/us21/n679 , \AES_ENC/us21/n678 ,\AES_ENC/us21/n677 , \AES_ENC/us21/n676 , \AES_ENC/us21/n675 ,\AES_ENC/us21/n674 , \AES_ENC/us21/n673 , \AES_ENC/us21/n672 ,\AES_ENC/us21/n671 , \AES_ENC/us21/n670 , \AES_ENC/us21/n669 ,\AES_ENC/us21/n668 , \AES_ENC/us21/n667 , \AES_ENC/us21/n666 ,\AES_ENC/us21/n665 , \AES_ENC/us21/n664 , \AES_ENC/us21/n663 ,\AES_ENC/us21/n662 , \AES_ENC/us21/n661 , \AES_ENC/us21/n660 ,\AES_ENC/us21/n659 , \AES_ENC/us21/n658 , \AES_ENC/us21/n657 ,\AES_ENC/us21/n656 , \AES_ENC/us21/n655 , \AES_ENC/us21/n654 ,\AES_ENC/us21/n653 , \AES_ENC/us21/n652 , \AES_ENC/us21/n651 ,\AES_ENC/us21/n650 , \AES_ENC/us21/n649 , \AES_ENC/us21/n648 ,\AES_ENC/us21/n647 , \AES_ENC/us21/n646 , \AES_ENC/us21/n645 ,\AES_ENC/us21/n644 , \AES_ENC/us21/n643 , \AES_ENC/us21/n642 ,\AES_ENC/us21/n641 , \AES_ENC/us21/n640 , \AES_ENC/us21/n639 ,\AES_ENC/us21/n638 , \AES_ENC/us21/n637 , \AES_ENC/us21/n636 ,\AES_ENC/us21/n635 , \AES_ENC/us21/n634 , \AES_ENC/us21/n633 ,\AES_ENC/us21/n632 , \AES_ENC/us21/n631 , \AES_ENC/us21/n630 ,\AES_ENC/us21/n629 , \AES_ENC/us21/n628 , \AES_ENC/us21/n627 ,\AES_ENC/us21/n626 , \AES_ENC/us21/n625 , \AES_ENC/us21/n624 ,\AES_ENC/us21/n623 , \AES_ENC/us21/n622 , \AES_ENC/us21/n621 ,\AES_ENC/us21/n620 , \AES_ENC/us21/n619 , \AES_ENC/us21/n618 ,\AES_ENC/us21/n617 , \AES_ENC/us21/n616 , \AES_ENC/us21/n615 ,\AES_ENC/us21/n614 , \AES_ENC/us21/n613 , \AES_ENC/us21/n612 ,\AES_ENC/us21/n611 , \AES_ENC/us21/n610 , \AES_ENC/us21/n609 ,\AES_ENC/us21/n608 , \AES_ENC/us21/n607 , \AES_ENC/us21/n606 ,\AES_ENC/us21/n605 , \AES_ENC/us21/n604 , \AES_ENC/us21/n603 ,\AES_ENC/us21/n602 , \AES_ENC/us21/n601 , \AES_ENC/us21/n600 ,\AES_ENC/us21/n599 , \AES_ENC/us21/n598 , \AES_ENC/us21/n597 ,\AES_ENC/us21/n596 , \AES_ENC/us21/n595 , \AES_ENC/us21/n594 ,\AES_ENC/us21/n593 , \AES_ENC/us21/n592 , \AES_ENC/us21/n591 ,\AES_ENC/us21/n590 , \AES_ENC/us21/n589 , \AES_ENC/us21/n588 ,\AES_ENC/us21/n587 , \AES_ENC/us21/n586 , \AES_ENC/us21/n585 ,\AES_ENC/us21/n584 , \AES_ENC/us21/n583 , \AES_ENC/us21/n582 ,\AES_ENC/us21/n581 , \AES_ENC/us21/n580 , \AES_ENC/us21/n579 ,\AES_ENC/us21/n578 , \AES_ENC/us21/n577 , \AES_ENC/us21/n576 ,\AES_ENC/us21/n575 , \AES_ENC/us21/n574 , \AES_ENC/us21/n573 ,\AES_ENC/us21/n572 , \AES_ENC/us21/n571 , \AES_ENC/us21/n570 ,\AES_ENC/us21/n569 , \AES_ENC/us22/n1135 , \AES_ENC/us22/n1134 ,\AES_ENC/us22/n1133 , \AES_ENC/us22/n1132 , \AES_ENC/us22/n1131 ,\AES_ENC/us22/n1130 , \AES_ENC/us22/n1129 , \AES_ENC/us22/n1128 ,\AES_ENC/us22/n1127 , \AES_ENC/us22/n1126 , \AES_ENC/us22/n1125 ,\AES_ENC/us22/n1124 , \AES_ENC/us22/n1123 , \AES_ENC/us22/n1122 ,\AES_ENC/us22/n1121 , \AES_ENC/us22/n1120 , \AES_ENC/us22/n1119 ,\AES_ENC/us22/n1118 , \AES_ENC/us22/n1117 , \AES_ENC/us22/n1116 ,\AES_ENC/us22/n1115 , \AES_ENC/us22/n1114 , \AES_ENC/us22/n1113 ,\AES_ENC/us22/n1112 , \AES_ENC/us22/n1111 , \AES_ENC/us22/n1110 ,\AES_ENC/us22/n1109 , \AES_ENC/us22/n1108 , \AES_ENC/us22/n1107 ,\AES_ENC/us22/n1106 , \AES_ENC/us22/n1105 , \AES_ENC/us22/n1104 ,\AES_ENC/us22/n1103 , \AES_ENC/us22/n1102 , \AES_ENC/us22/n1101 ,\AES_ENC/us22/n1100 , \AES_ENC/us22/n1099 , \AES_ENC/us22/n1098 ,\AES_ENC/us22/n1097 , \AES_ENC/us22/n1096 , \AES_ENC/us22/n1095 ,\AES_ENC/us22/n1094 , \AES_ENC/us22/n1093 , \AES_ENC/us22/n1092 ,\AES_ENC/us22/n1091 , \AES_ENC/us22/n1090 , \AES_ENC/us22/n1089 ,\AES_ENC/us22/n1088 , \AES_ENC/us22/n1087 , \AES_ENC/us22/n1086 ,\AES_ENC/us22/n1085 , \AES_ENC/us22/n1084 , \AES_ENC/us22/n1083 ,\AES_ENC/us22/n1082 , \AES_ENC/us22/n1081 , \AES_ENC/us22/n1080 ,\AES_ENC/us22/n1079 , \AES_ENC/us22/n1078 , \AES_ENC/us22/n1077 ,\AES_ENC/us22/n1076 , \AES_ENC/us22/n1075 , \AES_ENC/us22/n1074 ,\AES_ENC/us22/n1073 , \AES_ENC/us22/n1072 , \AES_ENC/us22/n1071 ,\AES_ENC/us22/n1070 , \AES_ENC/us22/n1069 , \AES_ENC/us22/n1068 ,\AES_ENC/us22/n1067 , \AES_ENC/us22/n1066 , \AES_ENC/us22/n1065 ,\AES_ENC/us22/n1064 , \AES_ENC/us22/n1063 , \AES_ENC/us22/n1062 ,\AES_ENC/us22/n1061 , \AES_ENC/us22/n1060 , \AES_ENC/us22/n1059 ,\AES_ENC/us22/n1058 , \AES_ENC/us22/n1057 , \AES_ENC/us22/n1056 ,\AES_ENC/us22/n1055 , \AES_ENC/us22/n1054 , \AES_ENC/us22/n1053 ,\AES_ENC/us22/n1052 , \AES_ENC/us22/n1051 , \AES_ENC/us22/n1050 ,\AES_ENC/us22/n1049 , \AES_ENC/us22/n1048 , \AES_ENC/us22/n1047 ,\AES_ENC/us22/n1046 , \AES_ENC/us22/n1045 , \AES_ENC/us22/n1044 ,\AES_ENC/us22/n1043 , \AES_ENC/us22/n1042 , \AES_ENC/us22/n1041 ,\AES_ENC/us22/n1040 , \AES_ENC/us22/n1039 , \AES_ENC/us22/n1038 ,\AES_ENC/us22/n1037 , \AES_ENC/us22/n1036 , \AES_ENC/us22/n1035 ,\AES_ENC/us22/n1034 , \AES_ENC/us22/n1033 , \AES_ENC/us22/n1032 ,\AES_ENC/us22/n1031 , \AES_ENC/us22/n1030 , \AES_ENC/us22/n1029 ,\AES_ENC/us22/n1028 , \AES_ENC/us22/n1027 , \AES_ENC/us22/n1026 ,\AES_ENC/us22/n1025 , \AES_ENC/us22/n1024 , \AES_ENC/us22/n1023 ,\AES_ENC/us22/n1022 , \AES_ENC/us22/n1021 , \AES_ENC/us22/n1020 ,\AES_ENC/us22/n1019 , \AES_ENC/us22/n1018 , \AES_ENC/us22/n1017 ,\AES_ENC/us22/n1016 , \AES_ENC/us22/n1015 , \AES_ENC/us22/n1014 ,\AES_ENC/us22/n1013 , \AES_ENC/us22/n1012 , \AES_ENC/us22/n1011 ,\AES_ENC/us22/n1010 , \AES_ENC/us22/n1009 , \AES_ENC/us22/n1008 ,\AES_ENC/us22/n1007 , \AES_ENC/us22/n1006 , \AES_ENC/us22/n1005 ,\AES_ENC/us22/n1004 , \AES_ENC/us22/n1003 , \AES_ENC/us22/n1002 ,\AES_ENC/us22/n1001 , \AES_ENC/us22/n1000 , \AES_ENC/us22/n999 ,\AES_ENC/us22/n998 , \AES_ENC/us22/n997 , \AES_ENC/us22/n996 ,\AES_ENC/us22/n995 , \AES_ENC/us22/n994 , \AES_ENC/us22/n993 ,\AES_ENC/us22/n992 , \AES_ENC/us22/n991 , \AES_ENC/us22/n990 ,\AES_ENC/us22/n989 , \AES_ENC/us22/n988 , \AES_ENC/us22/n987 ,\AES_ENC/us22/n986 , \AES_ENC/us22/n985 , \AES_ENC/us22/n984 ,\AES_ENC/us22/n983 , \AES_ENC/us22/n982 , \AES_ENC/us22/n981 ,\AES_ENC/us22/n980 , \AES_ENC/us22/n979 , \AES_ENC/us22/n978 ,\AES_ENC/us22/n977 , \AES_ENC/us22/n976 , \AES_ENC/us22/n975 ,\AES_ENC/us22/n974 , \AES_ENC/us22/n973 , \AES_ENC/us22/n972 ,\AES_ENC/us22/n971 , \AES_ENC/us22/n970 , \AES_ENC/us22/n969 ,\AES_ENC/us22/n968 , \AES_ENC/us22/n967 , \AES_ENC/us22/n966 ,\AES_ENC/us22/n965 , \AES_ENC/us22/n964 , \AES_ENC/us22/n963 ,\AES_ENC/us22/n962 , \AES_ENC/us22/n961 , \AES_ENC/us22/n960 ,\AES_ENC/us22/n959 , \AES_ENC/us22/n958 , \AES_ENC/us22/n957 ,\AES_ENC/us22/n956 , \AES_ENC/us22/n955 , \AES_ENC/us22/n954 ,\AES_ENC/us22/n953 , \AES_ENC/us22/n952 , \AES_ENC/us22/n951 ,\AES_ENC/us22/n950 , \AES_ENC/us22/n949 , \AES_ENC/us22/n948 ,\AES_ENC/us22/n947 , \AES_ENC/us22/n946 , \AES_ENC/us22/n945 ,\AES_ENC/us22/n944 , \AES_ENC/us22/n943 , \AES_ENC/us22/n942 ,\AES_ENC/us22/n941 , \AES_ENC/us22/n940 , \AES_ENC/us22/n939 ,\AES_ENC/us22/n938 , \AES_ENC/us22/n937 , \AES_ENC/us22/n936 ,\AES_ENC/us22/n935 , \AES_ENC/us22/n934 , \AES_ENC/us22/n933 ,\AES_ENC/us22/n932 , \AES_ENC/us22/n931 , \AES_ENC/us22/n930 ,\AES_ENC/us22/n929 , \AES_ENC/us22/n928 , \AES_ENC/us22/n927 ,\AES_ENC/us22/n926 , \AES_ENC/us22/n925 , \AES_ENC/us22/n924 ,\AES_ENC/us22/n923 , \AES_ENC/us22/n922 , \AES_ENC/us22/n921 ,\AES_ENC/us22/n920 , \AES_ENC/us22/n919 , \AES_ENC/us22/n918 ,\AES_ENC/us22/n917 , \AES_ENC/us22/n916 , \AES_ENC/us22/n915 ,\AES_ENC/us22/n914 , \AES_ENC/us22/n913 , \AES_ENC/us22/n912 ,\AES_ENC/us22/n911 , \AES_ENC/us22/n910 , \AES_ENC/us22/n909 ,\AES_ENC/us22/n908 , \AES_ENC/us22/n907 , \AES_ENC/us22/n906 ,\AES_ENC/us22/n905 , \AES_ENC/us22/n904 , \AES_ENC/us22/n903 ,\AES_ENC/us22/n902 , \AES_ENC/us22/n901 , \AES_ENC/us22/n900 ,\AES_ENC/us22/n899 , \AES_ENC/us22/n898 , \AES_ENC/us22/n897 ,\AES_ENC/us22/n896 , \AES_ENC/us22/n895 , \AES_ENC/us22/n894 ,\AES_ENC/us22/n893 , \AES_ENC/us22/n892 , \AES_ENC/us22/n891 ,\AES_ENC/us22/n890 , \AES_ENC/us22/n889 , \AES_ENC/us22/n888 ,\AES_ENC/us22/n887 , \AES_ENC/us22/n886 , \AES_ENC/us22/n885 ,\AES_ENC/us22/n884 , \AES_ENC/us22/n883 , \AES_ENC/us22/n882 ,\AES_ENC/us22/n881 , \AES_ENC/us22/n880 , \AES_ENC/us22/n879 ,\AES_ENC/us22/n878 , \AES_ENC/us22/n877 , \AES_ENC/us22/n876 ,\AES_ENC/us22/n875 , \AES_ENC/us22/n874 , \AES_ENC/us22/n873 ,\AES_ENC/us22/n872 , \AES_ENC/us22/n871 , \AES_ENC/us22/n870 ,\AES_ENC/us22/n869 , \AES_ENC/us22/n868 , \AES_ENC/us22/n867 ,\AES_ENC/us22/n866 , \AES_ENC/us22/n865 , \AES_ENC/us22/n864 ,\AES_ENC/us22/n863 , \AES_ENC/us22/n862 , \AES_ENC/us22/n861 ,\AES_ENC/us22/n860 , \AES_ENC/us22/n859 , \AES_ENC/us22/n858 ,\AES_ENC/us22/n857 , \AES_ENC/us22/n856 , \AES_ENC/us22/n855 ,\AES_ENC/us22/n854 , \AES_ENC/us22/n853 , \AES_ENC/us22/n852 ,\AES_ENC/us22/n851 , \AES_ENC/us22/n850 , \AES_ENC/us22/n849 ,\AES_ENC/us22/n848 , \AES_ENC/us22/n847 , \AES_ENC/us22/n846 ,\AES_ENC/us22/n845 , \AES_ENC/us22/n844 , \AES_ENC/us22/n843 ,\AES_ENC/us22/n842 , \AES_ENC/us22/n841 , \AES_ENC/us22/n840 ,\AES_ENC/us22/n839 , \AES_ENC/us22/n838 , \AES_ENC/us22/n837 ,\AES_ENC/us22/n836 , \AES_ENC/us22/n835 , \AES_ENC/us22/n834 ,\AES_ENC/us22/n833 , \AES_ENC/us22/n832 , \AES_ENC/us22/n831 ,\AES_ENC/us22/n830 , \AES_ENC/us22/n829 , \AES_ENC/us22/n828 ,\AES_ENC/us22/n827 , \AES_ENC/us22/n826 , \AES_ENC/us22/n825 ,\AES_ENC/us22/n824 , \AES_ENC/us22/n823 , \AES_ENC/us22/n822 ,\AES_ENC/us22/n821 , \AES_ENC/us22/n820 , \AES_ENC/us22/n819 ,\AES_ENC/us22/n818 , \AES_ENC/us22/n817 , \AES_ENC/us22/n816 ,\AES_ENC/us22/n815 , \AES_ENC/us22/n814 , \AES_ENC/us22/n813 ,\AES_ENC/us22/n812 , \AES_ENC/us22/n811 , \AES_ENC/us22/n810 ,\AES_ENC/us22/n809 , \AES_ENC/us22/n808 , \AES_ENC/us22/n807 ,\AES_ENC/us22/n806 , \AES_ENC/us22/n805 , \AES_ENC/us22/n804 ,\AES_ENC/us22/n803 , \AES_ENC/us22/n802 , \AES_ENC/us22/n801 ,\AES_ENC/us22/n800 , \AES_ENC/us22/n799 , \AES_ENC/us22/n798 ,\AES_ENC/us22/n797 , \AES_ENC/us22/n796 , \AES_ENC/us22/n795 ,\AES_ENC/us22/n794 , \AES_ENC/us22/n793 , \AES_ENC/us22/n792 ,\AES_ENC/us22/n791 , \AES_ENC/us22/n790 , \AES_ENC/us22/n789 ,\AES_ENC/us22/n788 , \AES_ENC/us22/n787 , \AES_ENC/us22/n786 ,\AES_ENC/us22/n785 , \AES_ENC/us22/n784 , \AES_ENC/us22/n783 ,\AES_ENC/us22/n782 , \AES_ENC/us22/n781 , \AES_ENC/us22/n780 ,\AES_ENC/us22/n779 , \AES_ENC/us22/n778 , \AES_ENC/us22/n777 ,\AES_ENC/us22/n776 , \AES_ENC/us22/n775 , \AES_ENC/us22/n774 ,\AES_ENC/us22/n773 , \AES_ENC/us22/n772 , \AES_ENC/us22/n771 ,\AES_ENC/us22/n770 , \AES_ENC/us22/n769 , \AES_ENC/us22/n768 ,\AES_ENC/us22/n767 , \AES_ENC/us22/n766 , \AES_ENC/us22/n765 ,\AES_ENC/us22/n764 , \AES_ENC/us22/n763 , \AES_ENC/us22/n762 ,\AES_ENC/us22/n761 , \AES_ENC/us22/n760 , \AES_ENC/us22/n759 ,\AES_ENC/us22/n758 , \AES_ENC/us22/n757 , \AES_ENC/us22/n756 ,\AES_ENC/us22/n755 , \AES_ENC/us22/n754 , \AES_ENC/us22/n753 ,\AES_ENC/us22/n752 , \AES_ENC/us22/n751 , \AES_ENC/us22/n750 ,\AES_ENC/us22/n749 , \AES_ENC/us22/n748 , \AES_ENC/us22/n747 ,\AES_ENC/us22/n746 , \AES_ENC/us22/n745 , \AES_ENC/us22/n744 ,\AES_ENC/us22/n743 , \AES_ENC/us22/n742 , \AES_ENC/us22/n741 ,\AES_ENC/us22/n740 , \AES_ENC/us22/n739 , \AES_ENC/us22/n738 ,\AES_ENC/us22/n737 , \AES_ENC/us22/n736 , \AES_ENC/us22/n735 ,\AES_ENC/us22/n734 , \AES_ENC/us22/n733 , \AES_ENC/us22/n732 ,\AES_ENC/us22/n731 , \AES_ENC/us22/n730 , \AES_ENC/us22/n729 ,\AES_ENC/us22/n728 , \AES_ENC/us22/n727 , \AES_ENC/us22/n726 ,\AES_ENC/us22/n725 , \AES_ENC/us22/n724 , \AES_ENC/us22/n723 ,\AES_ENC/us22/n722 , \AES_ENC/us22/n721 , \AES_ENC/us22/n720 ,\AES_ENC/us22/n719 , \AES_ENC/us22/n718 , \AES_ENC/us22/n717 ,\AES_ENC/us22/n716 , \AES_ENC/us22/n715 , \AES_ENC/us22/n714 ,\AES_ENC/us22/n713 , \AES_ENC/us22/n712 , \AES_ENC/us22/n711 ,\AES_ENC/us22/n710 , \AES_ENC/us22/n709 , \AES_ENC/us22/n708 ,\AES_ENC/us22/n707 , \AES_ENC/us22/n706 , \AES_ENC/us22/n705 ,\AES_ENC/us22/n704 , \AES_ENC/us22/n703 , \AES_ENC/us22/n702 ,\AES_ENC/us22/n701 , \AES_ENC/us22/n700 , \AES_ENC/us22/n699 ,\AES_ENC/us22/n698 , \AES_ENC/us22/n697 , \AES_ENC/us22/n696 ,\AES_ENC/us22/n695 , \AES_ENC/us22/n694 , \AES_ENC/us22/n693 ,\AES_ENC/us22/n692 , \AES_ENC/us22/n691 , \AES_ENC/us22/n690 ,\AES_ENC/us22/n689 , \AES_ENC/us22/n688 , \AES_ENC/us22/n687 ,\AES_ENC/us22/n686 , \AES_ENC/us22/n685 , \AES_ENC/us22/n684 ,\AES_ENC/us22/n683 , \AES_ENC/us22/n682 , \AES_ENC/us22/n681 ,\AES_ENC/us22/n680 , \AES_ENC/us22/n679 , \AES_ENC/us22/n678 ,\AES_ENC/us22/n677 , \AES_ENC/us22/n676 , \AES_ENC/us22/n675 ,\AES_ENC/us22/n674 , \AES_ENC/us22/n673 , \AES_ENC/us22/n672 ,\AES_ENC/us22/n671 , \AES_ENC/us22/n670 , \AES_ENC/us22/n669 ,\AES_ENC/us22/n668 , \AES_ENC/us22/n667 , \AES_ENC/us22/n666 ,\AES_ENC/us22/n665 , \AES_ENC/us22/n664 , \AES_ENC/us22/n663 ,\AES_ENC/us22/n662 , \AES_ENC/us22/n661 , \AES_ENC/us22/n660 ,\AES_ENC/us22/n659 , \AES_ENC/us22/n658 , \AES_ENC/us22/n657 ,\AES_ENC/us22/n656 , \AES_ENC/us22/n655 , \AES_ENC/us22/n654 ,\AES_ENC/us22/n653 , \AES_ENC/us22/n652 , \AES_ENC/us22/n651 ,\AES_ENC/us22/n650 , \AES_ENC/us22/n649 , \AES_ENC/us22/n648 ,\AES_ENC/us22/n647 , \AES_ENC/us22/n646 , \AES_ENC/us22/n645 ,\AES_ENC/us22/n644 , \AES_ENC/us22/n643 , \AES_ENC/us22/n642 ,\AES_ENC/us22/n641 , \AES_ENC/us22/n640 , \AES_ENC/us22/n639 ,\AES_ENC/us22/n638 , \AES_ENC/us22/n637 , \AES_ENC/us22/n636 ,\AES_ENC/us22/n635 , \AES_ENC/us22/n634 , \AES_ENC/us22/n633 ,\AES_ENC/us22/n632 , \AES_ENC/us22/n631 , \AES_ENC/us22/n630 ,\AES_ENC/us22/n629 , \AES_ENC/us22/n628 , \AES_ENC/us22/n627 ,\AES_ENC/us22/n626 , \AES_ENC/us22/n625 , \AES_ENC/us22/n624 ,\AES_ENC/us22/n623 , \AES_ENC/us22/n622 , \AES_ENC/us22/n621 ,\AES_ENC/us22/n620 , \AES_ENC/us22/n619 , \AES_ENC/us22/n618 ,\AES_ENC/us22/n617 , \AES_ENC/us22/n616 , \AES_ENC/us22/n615 ,\AES_ENC/us22/n614 , \AES_ENC/us22/n613 , \AES_ENC/us22/n612 ,\AES_ENC/us22/n611 , \AES_ENC/us22/n610 , \AES_ENC/us22/n609 ,\AES_ENC/us22/n608 , \AES_ENC/us22/n607 , \AES_ENC/us22/n606 ,\AES_ENC/us22/n605 , \AES_ENC/us22/n604 , \AES_ENC/us22/n603 ,\AES_ENC/us22/n602 , \AES_ENC/us22/n601 , \AES_ENC/us22/n600 ,\AES_ENC/us22/n599 , \AES_ENC/us22/n598 , \AES_ENC/us22/n597 ,\AES_ENC/us22/n596 , \AES_ENC/us22/n595 , \AES_ENC/us22/n594 ,\AES_ENC/us22/n593 , \AES_ENC/us22/n592 , \AES_ENC/us22/n591 ,\AES_ENC/us22/n590 , \AES_ENC/us22/n589 , \AES_ENC/us22/n588 ,\AES_ENC/us22/n587 , \AES_ENC/us22/n586 , \AES_ENC/us22/n585 ,\AES_ENC/us22/n584 , \AES_ENC/us22/n583 , \AES_ENC/us22/n582 ,\AES_ENC/us22/n581 , \AES_ENC/us22/n580 , \AES_ENC/us22/n579 ,\AES_ENC/us22/n578 , \AES_ENC/us22/n577 , \AES_ENC/us22/n576 ,\AES_ENC/us22/n575 , \AES_ENC/us22/n574 , \AES_ENC/us22/n573 ,\AES_ENC/us22/n572 , \AES_ENC/us22/n571 , \AES_ENC/us22/n570 ,\AES_ENC/us22/n569 , \AES_ENC/us23/n1135 , \AES_ENC/us23/n1134 ,\AES_ENC/us23/n1133 , \AES_ENC/us23/n1132 , \AES_ENC/us23/n1131 ,\AES_ENC/us23/n1130 , \AES_ENC/us23/n1129 , \AES_ENC/us23/n1128 ,\AES_ENC/us23/n1127 , \AES_ENC/us23/n1126 , \AES_ENC/us23/n1125 ,\AES_ENC/us23/n1124 , \AES_ENC/us23/n1123 , \AES_ENC/us23/n1122 ,\AES_ENC/us23/n1121 , \AES_ENC/us23/n1120 , \AES_ENC/us23/n1119 ,\AES_ENC/us23/n1118 , \AES_ENC/us23/n1117 , \AES_ENC/us23/n1116 ,\AES_ENC/us23/n1115 , \AES_ENC/us23/n1114 , \AES_ENC/us23/n1113 ,\AES_ENC/us23/n1112 , \AES_ENC/us23/n1111 , \AES_ENC/us23/n1110 ,\AES_ENC/us23/n1109 , \AES_ENC/us23/n1108 , \AES_ENC/us23/n1107 ,\AES_ENC/us23/n1106 , \AES_ENC/us23/n1105 , \AES_ENC/us23/n1104 ,\AES_ENC/us23/n1103 , \AES_ENC/us23/n1102 , \AES_ENC/us23/n1101 ,\AES_ENC/us23/n1100 , \AES_ENC/us23/n1099 , \AES_ENC/us23/n1098 ,\AES_ENC/us23/n1097 , \AES_ENC/us23/n1096 , \AES_ENC/us23/n1095 ,\AES_ENC/us23/n1094 , \AES_ENC/us23/n1093 , \AES_ENC/us23/n1092 ,\AES_ENC/us23/n1091 , \AES_ENC/us23/n1090 , \AES_ENC/us23/n1089 ,\AES_ENC/us23/n1088 , \AES_ENC/us23/n1087 , \AES_ENC/us23/n1086 ,\AES_ENC/us23/n1085 , \AES_ENC/us23/n1084 , \AES_ENC/us23/n1083 ,\AES_ENC/us23/n1082 , \AES_ENC/us23/n1081 , \AES_ENC/us23/n1080 ,\AES_ENC/us23/n1079 , \AES_ENC/us23/n1078 , \AES_ENC/us23/n1077 ,\AES_ENC/us23/n1076 , \AES_ENC/us23/n1075 , \AES_ENC/us23/n1074 ,\AES_ENC/us23/n1073 , \AES_ENC/us23/n1072 , \AES_ENC/us23/n1071 ,\AES_ENC/us23/n1070 , \AES_ENC/us23/n1069 , \AES_ENC/us23/n1068 ,\AES_ENC/us23/n1067 , \AES_ENC/us23/n1066 , \AES_ENC/us23/n1065 ,\AES_ENC/us23/n1064 , \AES_ENC/us23/n1063 , \AES_ENC/us23/n1062 ,\AES_ENC/us23/n1061 , \AES_ENC/us23/n1060 , \AES_ENC/us23/n1059 ,\AES_ENC/us23/n1058 , \AES_ENC/us23/n1057 , \AES_ENC/us23/n1056 ,\AES_ENC/us23/n1055 , \AES_ENC/us23/n1054 , \AES_ENC/us23/n1053 ,\AES_ENC/us23/n1052 , \AES_ENC/us23/n1051 , \AES_ENC/us23/n1050 ,\AES_ENC/us23/n1049 , \AES_ENC/us23/n1048 , \AES_ENC/us23/n1047 ,\AES_ENC/us23/n1046 , \AES_ENC/us23/n1045 , \AES_ENC/us23/n1044 ,\AES_ENC/us23/n1043 , \AES_ENC/us23/n1042 , \AES_ENC/us23/n1041 ,\AES_ENC/us23/n1040 , \AES_ENC/us23/n1039 , \AES_ENC/us23/n1038 ,\AES_ENC/us23/n1037 , \AES_ENC/us23/n1036 , \AES_ENC/us23/n1035 ,\AES_ENC/us23/n1034 , \AES_ENC/us23/n1033 , \AES_ENC/us23/n1032 ,\AES_ENC/us23/n1031 , \AES_ENC/us23/n1030 , \AES_ENC/us23/n1029 ,\AES_ENC/us23/n1028 , \AES_ENC/us23/n1027 , \AES_ENC/us23/n1026 ,\AES_ENC/us23/n1025 , \AES_ENC/us23/n1024 , \AES_ENC/us23/n1023 ,\AES_ENC/us23/n1022 , \AES_ENC/us23/n1021 , \AES_ENC/us23/n1020 ,\AES_ENC/us23/n1019 , \AES_ENC/us23/n1018 , \AES_ENC/us23/n1017 ,\AES_ENC/us23/n1016 , \AES_ENC/us23/n1015 , \AES_ENC/us23/n1014 ,\AES_ENC/us23/n1013 , \AES_ENC/us23/n1012 , \AES_ENC/us23/n1011 ,\AES_ENC/us23/n1010 , \AES_ENC/us23/n1009 , \AES_ENC/us23/n1008 ,\AES_ENC/us23/n1007 , \AES_ENC/us23/n1006 , \AES_ENC/us23/n1005 ,\AES_ENC/us23/n1004 , \AES_ENC/us23/n1003 , \AES_ENC/us23/n1002 ,\AES_ENC/us23/n1001 , \AES_ENC/us23/n1000 , \AES_ENC/us23/n999 ,\AES_ENC/us23/n998 , \AES_ENC/us23/n997 , \AES_ENC/us23/n996 ,\AES_ENC/us23/n995 , \AES_ENC/us23/n994 , \AES_ENC/us23/n993 ,\AES_ENC/us23/n992 , \AES_ENC/us23/n991 , \AES_ENC/us23/n990 ,\AES_ENC/us23/n989 , \AES_ENC/us23/n988 , \AES_ENC/us23/n987 ,\AES_ENC/us23/n986 , \AES_ENC/us23/n985 , \AES_ENC/us23/n984 ,\AES_ENC/us23/n983 , \AES_ENC/us23/n982 , \AES_ENC/us23/n981 ,\AES_ENC/us23/n980 , \AES_ENC/us23/n979 , \AES_ENC/us23/n978 ,\AES_ENC/us23/n977 , \AES_ENC/us23/n976 , \AES_ENC/us23/n975 ,\AES_ENC/us23/n974 , \AES_ENC/us23/n973 , \AES_ENC/us23/n972 ,\AES_ENC/us23/n971 , \AES_ENC/us23/n970 , \AES_ENC/us23/n969 ,\AES_ENC/us23/n968 , \AES_ENC/us23/n967 , \AES_ENC/us23/n966 ,\AES_ENC/us23/n965 , \AES_ENC/us23/n964 , \AES_ENC/us23/n963 ,\AES_ENC/us23/n962 , \AES_ENC/us23/n961 , \AES_ENC/us23/n960 ,\AES_ENC/us23/n959 , \AES_ENC/us23/n958 , \AES_ENC/us23/n957 ,\AES_ENC/us23/n956 , \AES_ENC/us23/n955 , \AES_ENC/us23/n954 ,\AES_ENC/us23/n953 , \AES_ENC/us23/n952 , \AES_ENC/us23/n951 ,\AES_ENC/us23/n950 , \AES_ENC/us23/n949 , \AES_ENC/us23/n948 ,\AES_ENC/us23/n947 , \AES_ENC/us23/n946 , \AES_ENC/us23/n945 ,\AES_ENC/us23/n944 , \AES_ENC/us23/n943 , \AES_ENC/us23/n942 ,\AES_ENC/us23/n941 , \AES_ENC/us23/n940 , \AES_ENC/us23/n939 ,\AES_ENC/us23/n938 , \AES_ENC/us23/n937 , \AES_ENC/us23/n936 ,\AES_ENC/us23/n935 , \AES_ENC/us23/n934 , \AES_ENC/us23/n933 ,\AES_ENC/us23/n932 , \AES_ENC/us23/n931 , \AES_ENC/us23/n930 ,\AES_ENC/us23/n929 , \AES_ENC/us23/n928 , \AES_ENC/us23/n927 ,\AES_ENC/us23/n926 , \AES_ENC/us23/n925 , \AES_ENC/us23/n924 ,\AES_ENC/us23/n923 , \AES_ENC/us23/n922 , \AES_ENC/us23/n921 ,\AES_ENC/us23/n920 , \AES_ENC/us23/n919 , \AES_ENC/us23/n918 ,\AES_ENC/us23/n917 , \AES_ENC/us23/n916 , \AES_ENC/us23/n915 ,\AES_ENC/us23/n914 , \AES_ENC/us23/n913 , \AES_ENC/us23/n912 ,\AES_ENC/us23/n911 , \AES_ENC/us23/n910 , \AES_ENC/us23/n909 ,\AES_ENC/us23/n908 , \AES_ENC/us23/n907 , \AES_ENC/us23/n906 ,\AES_ENC/us23/n905 , \AES_ENC/us23/n904 , \AES_ENC/us23/n903 ,\AES_ENC/us23/n902 , \AES_ENC/us23/n901 , \AES_ENC/us23/n900 ,\AES_ENC/us23/n899 , \AES_ENC/us23/n898 , \AES_ENC/us23/n897 ,\AES_ENC/us23/n896 , \AES_ENC/us23/n895 , \AES_ENC/us23/n894 ,\AES_ENC/us23/n893 , \AES_ENC/us23/n892 , \AES_ENC/us23/n891 ,\AES_ENC/us23/n890 , \AES_ENC/us23/n889 , \AES_ENC/us23/n888 ,\AES_ENC/us23/n887 , \AES_ENC/us23/n886 , \AES_ENC/us23/n885 ,\AES_ENC/us23/n884 , \AES_ENC/us23/n883 , \AES_ENC/us23/n882 ,\AES_ENC/us23/n881 , \AES_ENC/us23/n880 , \AES_ENC/us23/n879 ,\AES_ENC/us23/n878 , \AES_ENC/us23/n877 , \AES_ENC/us23/n876 ,\AES_ENC/us23/n875 , \AES_ENC/us23/n874 , \AES_ENC/us23/n873 ,\AES_ENC/us23/n872 , \AES_ENC/us23/n871 , \AES_ENC/us23/n870 ,\AES_ENC/us23/n869 , \AES_ENC/us23/n868 , \AES_ENC/us23/n867 ,\AES_ENC/us23/n866 , \AES_ENC/us23/n865 , \AES_ENC/us23/n864 ,\AES_ENC/us23/n863 , \AES_ENC/us23/n862 , \AES_ENC/us23/n861 ,\AES_ENC/us23/n860 , \AES_ENC/us23/n859 , \AES_ENC/us23/n858 ,\AES_ENC/us23/n857 , \AES_ENC/us23/n856 , \AES_ENC/us23/n855 ,\AES_ENC/us23/n854 , \AES_ENC/us23/n853 , \AES_ENC/us23/n852 ,\AES_ENC/us23/n851 , \AES_ENC/us23/n850 , \AES_ENC/us23/n849 ,\AES_ENC/us23/n848 , \AES_ENC/us23/n847 , \AES_ENC/us23/n846 ,\AES_ENC/us23/n845 , \AES_ENC/us23/n844 , \AES_ENC/us23/n843 ,\AES_ENC/us23/n842 , \AES_ENC/us23/n841 , \AES_ENC/us23/n840 ,\AES_ENC/us23/n839 , \AES_ENC/us23/n838 , \AES_ENC/us23/n837 ,\AES_ENC/us23/n836 , \AES_ENC/us23/n835 , \AES_ENC/us23/n834 ,\AES_ENC/us23/n833 , \AES_ENC/us23/n832 , \AES_ENC/us23/n831 ,\AES_ENC/us23/n830 , \AES_ENC/us23/n829 , \AES_ENC/us23/n828 ,\AES_ENC/us23/n827 , \AES_ENC/us23/n826 , \AES_ENC/us23/n825 ,\AES_ENC/us23/n824 , \AES_ENC/us23/n823 , \AES_ENC/us23/n822 ,\AES_ENC/us23/n821 , \AES_ENC/us23/n820 , \AES_ENC/us23/n819 ,\AES_ENC/us23/n818 , \AES_ENC/us23/n817 , \AES_ENC/us23/n816 ,\AES_ENC/us23/n815 , \AES_ENC/us23/n814 , \AES_ENC/us23/n813 ,\AES_ENC/us23/n812 , \AES_ENC/us23/n811 , \AES_ENC/us23/n810 ,\AES_ENC/us23/n809 , \AES_ENC/us23/n808 , \AES_ENC/us23/n807 ,\AES_ENC/us23/n806 , \AES_ENC/us23/n805 , \AES_ENC/us23/n804 ,\AES_ENC/us23/n803 , \AES_ENC/us23/n802 , \AES_ENC/us23/n801 ,\AES_ENC/us23/n800 , \AES_ENC/us23/n799 , \AES_ENC/us23/n798 ,\AES_ENC/us23/n797 , \AES_ENC/us23/n796 , \AES_ENC/us23/n795 ,\AES_ENC/us23/n794 , \AES_ENC/us23/n793 , \AES_ENC/us23/n792 ,\AES_ENC/us23/n791 , \AES_ENC/us23/n790 , \AES_ENC/us23/n789 ,\AES_ENC/us23/n788 , \AES_ENC/us23/n787 , \AES_ENC/us23/n786 ,\AES_ENC/us23/n785 , \AES_ENC/us23/n784 , \AES_ENC/us23/n783 ,\AES_ENC/us23/n782 , \AES_ENC/us23/n781 , \AES_ENC/us23/n780 ,\AES_ENC/us23/n779 , \AES_ENC/us23/n778 , \AES_ENC/us23/n777 ,\AES_ENC/us23/n776 , \AES_ENC/us23/n775 , \AES_ENC/us23/n774 ,\AES_ENC/us23/n773 , \AES_ENC/us23/n772 , \AES_ENC/us23/n771 ,\AES_ENC/us23/n770 , \AES_ENC/us23/n769 , \AES_ENC/us23/n768 ,\AES_ENC/us23/n767 , \AES_ENC/us23/n766 , \AES_ENC/us23/n765 ,\AES_ENC/us23/n764 , \AES_ENC/us23/n763 , \AES_ENC/us23/n762 ,\AES_ENC/us23/n761 , \AES_ENC/us23/n760 , \AES_ENC/us23/n759 ,\AES_ENC/us23/n758 , \AES_ENC/us23/n757 , \AES_ENC/us23/n756 ,\AES_ENC/us23/n755 , \AES_ENC/us23/n754 , \AES_ENC/us23/n753 ,\AES_ENC/us23/n752 , \AES_ENC/us23/n751 , \AES_ENC/us23/n750 ,\AES_ENC/us23/n749 , \AES_ENC/us23/n748 , \AES_ENC/us23/n747 ,\AES_ENC/us23/n746 , \AES_ENC/us23/n745 , \AES_ENC/us23/n744 ,\AES_ENC/us23/n743 , \AES_ENC/us23/n742 , \AES_ENC/us23/n741 ,\AES_ENC/us23/n740 , \AES_ENC/us23/n739 , \AES_ENC/us23/n738 ,\AES_ENC/us23/n737 , \AES_ENC/us23/n736 , \AES_ENC/us23/n735 ,\AES_ENC/us23/n734 , \AES_ENC/us23/n733 , \AES_ENC/us23/n732 ,\AES_ENC/us23/n731 , \AES_ENC/us23/n730 , \AES_ENC/us23/n729 ,\AES_ENC/us23/n728 , \AES_ENC/us23/n727 , \AES_ENC/us23/n726 ,\AES_ENC/us23/n725 , \AES_ENC/us23/n724 , \AES_ENC/us23/n723 ,\AES_ENC/us23/n722 , \AES_ENC/us23/n721 , \AES_ENC/us23/n720 ,\AES_ENC/us23/n719 , \AES_ENC/us23/n718 , \AES_ENC/us23/n717 ,\AES_ENC/us23/n716 , \AES_ENC/us23/n715 , \AES_ENC/us23/n714 ,\AES_ENC/us23/n713 , \AES_ENC/us23/n712 , \AES_ENC/us23/n711 ,\AES_ENC/us23/n710 , \AES_ENC/us23/n709 , \AES_ENC/us23/n708 ,\AES_ENC/us23/n707 , \AES_ENC/us23/n706 , \AES_ENC/us23/n705 ,\AES_ENC/us23/n704 , \AES_ENC/us23/n703 , \AES_ENC/us23/n702 ,\AES_ENC/us23/n701 , \AES_ENC/us23/n700 , \AES_ENC/us23/n699 ,\AES_ENC/us23/n698 , \AES_ENC/us23/n697 , \AES_ENC/us23/n696 ,\AES_ENC/us23/n695 , \AES_ENC/us23/n694 , \AES_ENC/us23/n693 ,\AES_ENC/us23/n692 , \AES_ENC/us23/n691 , \AES_ENC/us23/n690 ,\AES_ENC/us23/n689 , \AES_ENC/us23/n688 , \AES_ENC/us23/n687 ,\AES_ENC/us23/n686 , \AES_ENC/us23/n685 , \AES_ENC/us23/n684 ,\AES_ENC/us23/n683 , \AES_ENC/us23/n682 , \AES_ENC/us23/n681 ,\AES_ENC/us23/n680 , \AES_ENC/us23/n679 , \AES_ENC/us23/n678 ,\AES_ENC/us23/n677 , \AES_ENC/us23/n676 , \AES_ENC/us23/n675 ,\AES_ENC/us23/n674 , \AES_ENC/us23/n673 , \AES_ENC/us23/n672 ,\AES_ENC/us23/n671 , \AES_ENC/us23/n670 , \AES_ENC/us23/n669 ,\AES_ENC/us23/n668 , \AES_ENC/us23/n667 , \AES_ENC/us23/n666 ,\AES_ENC/us23/n665 , \AES_ENC/us23/n664 , \AES_ENC/us23/n663 ,\AES_ENC/us23/n662 , \AES_ENC/us23/n661 , \AES_ENC/us23/n660 ,\AES_ENC/us23/n659 , \AES_ENC/us23/n658 , \AES_ENC/us23/n657 ,\AES_ENC/us23/n656 , \AES_ENC/us23/n655 , \AES_ENC/us23/n654 ,\AES_ENC/us23/n653 , \AES_ENC/us23/n652 , \AES_ENC/us23/n651 ,\AES_ENC/us23/n650 , \AES_ENC/us23/n649 , \AES_ENC/us23/n648 ,\AES_ENC/us23/n647 , \AES_ENC/us23/n646 , \AES_ENC/us23/n645 ,\AES_ENC/us23/n644 , \AES_ENC/us23/n643 , \AES_ENC/us23/n642 ,\AES_ENC/us23/n641 , \AES_ENC/us23/n640 , \AES_ENC/us23/n639 ,\AES_ENC/us23/n638 , \AES_ENC/us23/n637 , \AES_ENC/us23/n636 ,\AES_ENC/us23/n635 , \AES_ENC/us23/n634 , \AES_ENC/us23/n633 ,\AES_ENC/us23/n632 , \AES_ENC/us23/n631 , \AES_ENC/us23/n630 ,\AES_ENC/us23/n629 , \AES_ENC/us23/n628 , \AES_ENC/us23/n627 ,\AES_ENC/us23/n626 , \AES_ENC/us23/n625 , \AES_ENC/us23/n624 ,\AES_ENC/us23/n623 , \AES_ENC/us23/n622 , \AES_ENC/us23/n621 ,\AES_ENC/us23/n620 , \AES_ENC/us23/n619 , \AES_ENC/us23/n618 ,\AES_ENC/us23/n617 , \AES_ENC/us23/n616 , \AES_ENC/us23/n615 ,\AES_ENC/us23/n614 , \AES_ENC/us23/n613 , \AES_ENC/us23/n612 ,\AES_ENC/us23/n611 , \AES_ENC/us23/n610 , \AES_ENC/us23/n609 ,\AES_ENC/us23/n608 , \AES_ENC/us23/n607 , \AES_ENC/us23/n606 ,\AES_ENC/us23/n605 , \AES_ENC/us23/n604 , \AES_ENC/us23/n603 ,\AES_ENC/us23/n602 , \AES_ENC/us23/n601 , \AES_ENC/us23/n600 ,\AES_ENC/us23/n599 , \AES_ENC/us23/n598 , \AES_ENC/us23/n597 ,\AES_ENC/us23/n596 , \AES_ENC/us23/n595 , \AES_ENC/us23/n594 ,\AES_ENC/us23/n593 , \AES_ENC/us23/n592 , \AES_ENC/us23/n591 ,\AES_ENC/us23/n590 , \AES_ENC/us23/n589 , \AES_ENC/us23/n588 ,\AES_ENC/us23/n587 , \AES_ENC/us23/n586 , \AES_ENC/us23/n585 ,\AES_ENC/us23/n584 , \AES_ENC/us23/n583 , \AES_ENC/us23/n582 ,\AES_ENC/us23/n581 , \AES_ENC/us23/n580 , \AES_ENC/us23/n579 ,\AES_ENC/us23/n578 , \AES_ENC/us23/n577 , \AES_ENC/us23/n576 ,\AES_ENC/us23/n575 , \AES_ENC/us23/n574 , \AES_ENC/us23/n573 ,\AES_ENC/us23/n572 , \AES_ENC/us23/n571 , \AES_ENC/us23/n570 ,\AES_ENC/us23/n569 , \AES_ENC/us30/n1135 , \AES_ENC/us30/n1134 ,\AES_ENC/us30/n1133 , \AES_ENC/us30/n1132 , \AES_ENC/us30/n1131 ,\AES_ENC/us30/n1130 , \AES_ENC/us30/n1129 , \AES_ENC/us30/n1128 ,\AES_ENC/us30/n1127 , \AES_ENC/us30/n1126 , \AES_ENC/us30/n1125 ,\AES_ENC/us30/n1124 , \AES_ENC/us30/n1123 , \AES_ENC/us30/n1122 ,\AES_ENC/us30/n1121 , \AES_ENC/us30/n1120 , \AES_ENC/us30/n1119 ,\AES_ENC/us30/n1118 , \AES_ENC/us30/n1117 , \AES_ENC/us30/n1116 ,\AES_ENC/us30/n1115 , \AES_ENC/us30/n1114 , \AES_ENC/us30/n1113 ,\AES_ENC/us30/n1112 , \AES_ENC/us30/n1111 , \AES_ENC/us30/n1110 ,\AES_ENC/us30/n1109 , \AES_ENC/us30/n1108 , \AES_ENC/us30/n1107 ,\AES_ENC/us30/n1106 , \AES_ENC/us30/n1105 , \AES_ENC/us30/n1104 ,\AES_ENC/us30/n1103 , \AES_ENC/us30/n1102 , \AES_ENC/us30/n1101 ,\AES_ENC/us30/n1100 , \AES_ENC/us30/n1099 , \AES_ENC/us30/n1098 ,\AES_ENC/us30/n1097 , \AES_ENC/us30/n1096 , \AES_ENC/us30/n1095 ,\AES_ENC/us30/n1094 , \AES_ENC/us30/n1093 , \AES_ENC/us30/n1092 ,\AES_ENC/us30/n1091 , \AES_ENC/us30/n1090 , \AES_ENC/us30/n1089 ,\AES_ENC/us30/n1088 , \AES_ENC/us30/n1087 , \AES_ENC/us30/n1086 ,\AES_ENC/us30/n1085 , \AES_ENC/us30/n1084 , \AES_ENC/us30/n1083 ,\AES_ENC/us30/n1082 , \AES_ENC/us30/n1081 , \AES_ENC/us30/n1080 ,\AES_ENC/us30/n1079 , \AES_ENC/us30/n1078 , \AES_ENC/us30/n1077 ,\AES_ENC/us30/n1076 , \AES_ENC/us30/n1075 , \AES_ENC/us30/n1074 ,\AES_ENC/us30/n1073 , \AES_ENC/us30/n1072 , \AES_ENC/us30/n1071 ,\AES_ENC/us30/n1070 , \AES_ENC/us30/n1069 , \AES_ENC/us30/n1068 ,\AES_ENC/us30/n1067 , \AES_ENC/us30/n1066 , \AES_ENC/us30/n1065 ,\AES_ENC/us30/n1064 , \AES_ENC/us30/n1063 , \AES_ENC/us30/n1062 ,\AES_ENC/us30/n1061 , \AES_ENC/us30/n1060 , \AES_ENC/us30/n1059 ,\AES_ENC/us30/n1058 , \AES_ENC/us30/n1057 , \AES_ENC/us30/n1056 ,\AES_ENC/us30/n1055 , \AES_ENC/us30/n1054 , \AES_ENC/us30/n1053 ,\AES_ENC/us30/n1052 , \AES_ENC/us30/n1051 , \AES_ENC/us30/n1050 ,\AES_ENC/us30/n1049 , \AES_ENC/us30/n1048 , \AES_ENC/us30/n1047 ,\AES_ENC/us30/n1046 , \AES_ENC/us30/n1045 , \AES_ENC/us30/n1044 ,\AES_ENC/us30/n1043 , \AES_ENC/us30/n1042 , \AES_ENC/us30/n1041 ,\AES_ENC/us30/n1040 , \AES_ENC/us30/n1039 , \AES_ENC/us30/n1038 ,\AES_ENC/us30/n1037 , \AES_ENC/us30/n1036 , \AES_ENC/us30/n1035 ,\AES_ENC/us30/n1034 , \AES_ENC/us30/n1033 , \AES_ENC/us30/n1032 ,\AES_ENC/us30/n1031 , \AES_ENC/us30/n1030 , \AES_ENC/us30/n1029 ,\AES_ENC/us30/n1028 , \AES_ENC/us30/n1027 , \AES_ENC/us30/n1026 ,\AES_ENC/us30/n1025 , \AES_ENC/us30/n1024 , \AES_ENC/us30/n1023 ,\AES_ENC/us30/n1022 , \AES_ENC/us30/n1021 , \AES_ENC/us30/n1020 ,\AES_ENC/us30/n1019 , \AES_ENC/us30/n1018 , \AES_ENC/us30/n1017 ,\AES_ENC/us30/n1016 , \AES_ENC/us30/n1015 , \AES_ENC/us30/n1014 ,\AES_ENC/us30/n1013 , \AES_ENC/us30/n1012 , \AES_ENC/us30/n1011 ,\AES_ENC/us30/n1010 , \AES_ENC/us30/n1009 , \AES_ENC/us30/n1008 ,\AES_ENC/us30/n1007 , \AES_ENC/us30/n1006 , \AES_ENC/us30/n1005 ,\AES_ENC/us30/n1004 , \AES_ENC/us30/n1003 , \AES_ENC/us30/n1002 ,\AES_ENC/us30/n1001 , \AES_ENC/us30/n1000 , \AES_ENC/us30/n999 ,\AES_ENC/us30/n998 , \AES_ENC/us30/n997 , \AES_ENC/us30/n996 ,\AES_ENC/us30/n995 , \AES_ENC/us30/n994 , \AES_ENC/us30/n993 ,\AES_ENC/us30/n992 , \AES_ENC/us30/n991 , \AES_ENC/us30/n990 ,\AES_ENC/us30/n989 , \AES_ENC/us30/n988 , \AES_ENC/us30/n987 ,\AES_ENC/us30/n986 , \AES_ENC/us30/n985 , \AES_ENC/us30/n984 ,\AES_ENC/us30/n983 , \AES_ENC/us30/n982 , \AES_ENC/us30/n981 ,\AES_ENC/us30/n980 , \AES_ENC/us30/n979 , \AES_ENC/us30/n978 ,\AES_ENC/us30/n977 , \AES_ENC/us30/n976 , \AES_ENC/us30/n975 ,\AES_ENC/us30/n974 , \AES_ENC/us30/n973 , \AES_ENC/us30/n972 ,\AES_ENC/us30/n971 , \AES_ENC/us30/n970 , \AES_ENC/us30/n969 ,\AES_ENC/us30/n968 , \AES_ENC/us30/n967 , \AES_ENC/us30/n966 ,\AES_ENC/us30/n965 , \AES_ENC/us30/n964 , \AES_ENC/us30/n963 ,\AES_ENC/us30/n962 , \AES_ENC/us30/n961 , \AES_ENC/us30/n960 ,\AES_ENC/us30/n959 , \AES_ENC/us30/n958 , \AES_ENC/us30/n957 ,\AES_ENC/us30/n956 , \AES_ENC/us30/n955 , \AES_ENC/us30/n954 ,\AES_ENC/us30/n953 , \AES_ENC/us30/n952 , \AES_ENC/us30/n951 ,\AES_ENC/us30/n950 , \AES_ENC/us30/n949 , \AES_ENC/us30/n948 ,\AES_ENC/us30/n947 , \AES_ENC/us30/n946 , \AES_ENC/us30/n945 ,\AES_ENC/us30/n944 , \AES_ENC/us30/n943 , \AES_ENC/us30/n942 ,\AES_ENC/us30/n941 , \AES_ENC/us30/n940 , \AES_ENC/us30/n939 ,\AES_ENC/us30/n938 , \AES_ENC/us30/n937 , \AES_ENC/us30/n936 ,\AES_ENC/us30/n935 , \AES_ENC/us30/n934 , \AES_ENC/us30/n933 ,\AES_ENC/us30/n932 , \AES_ENC/us30/n931 , \AES_ENC/us30/n930 ,\AES_ENC/us30/n929 , \AES_ENC/us30/n928 , \AES_ENC/us30/n927 ,\AES_ENC/us30/n926 , \AES_ENC/us30/n925 , \AES_ENC/us30/n924 ,\AES_ENC/us30/n923 , \AES_ENC/us30/n922 , \AES_ENC/us30/n921 ,\AES_ENC/us30/n920 , \AES_ENC/us30/n919 , \AES_ENC/us30/n918 ,\AES_ENC/us30/n917 , \AES_ENC/us30/n916 , \AES_ENC/us30/n915 ,\AES_ENC/us30/n914 , \AES_ENC/us30/n913 , \AES_ENC/us30/n912 ,\AES_ENC/us30/n911 , \AES_ENC/us30/n910 , \AES_ENC/us30/n909 ,\AES_ENC/us30/n908 , \AES_ENC/us30/n907 , \AES_ENC/us30/n906 ,\AES_ENC/us30/n905 , \AES_ENC/us30/n904 , \AES_ENC/us30/n903 ,\AES_ENC/us30/n902 , \AES_ENC/us30/n901 , \AES_ENC/us30/n900 ,\AES_ENC/us30/n899 , \AES_ENC/us30/n898 , \AES_ENC/us30/n897 ,\AES_ENC/us30/n896 , \AES_ENC/us30/n895 , \AES_ENC/us30/n894 ,\AES_ENC/us30/n893 , \AES_ENC/us30/n892 , \AES_ENC/us30/n891 ,\AES_ENC/us30/n890 , \AES_ENC/us30/n889 , \AES_ENC/us30/n888 ,\AES_ENC/us30/n887 , \AES_ENC/us30/n886 , \AES_ENC/us30/n885 ,\AES_ENC/us30/n884 , \AES_ENC/us30/n883 , \AES_ENC/us30/n882 ,\AES_ENC/us30/n881 , \AES_ENC/us30/n880 , \AES_ENC/us30/n879 ,\AES_ENC/us30/n878 , \AES_ENC/us30/n877 , \AES_ENC/us30/n876 ,\AES_ENC/us30/n875 , \AES_ENC/us30/n874 , \AES_ENC/us30/n873 ,\AES_ENC/us30/n872 , \AES_ENC/us30/n871 , \AES_ENC/us30/n870 ,\AES_ENC/us30/n869 , \AES_ENC/us30/n868 , \AES_ENC/us30/n867 ,\AES_ENC/us30/n866 , \AES_ENC/us30/n865 , \AES_ENC/us30/n864 ,\AES_ENC/us30/n863 , \AES_ENC/us30/n862 , \AES_ENC/us30/n861 ,\AES_ENC/us30/n860 , \AES_ENC/us30/n859 , \AES_ENC/us30/n858 ,\AES_ENC/us30/n857 , \AES_ENC/us30/n856 , \AES_ENC/us30/n855 ,\AES_ENC/us30/n854 , \AES_ENC/us30/n853 , \AES_ENC/us30/n852 ,\AES_ENC/us30/n851 , \AES_ENC/us30/n850 , \AES_ENC/us30/n849 ,\AES_ENC/us30/n848 , \AES_ENC/us30/n847 , \AES_ENC/us30/n846 ,\AES_ENC/us30/n845 , \AES_ENC/us30/n844 , \AES_ENC/us30/n843 ,\AES_ENC/us30/n842 , \AES_ENC/us30/n841 , \AES_ENC/us30/n840 ,\AES_ENC/us30/n839 , \AES_ENC/us30/n838 , \AES_ENC/us30/n837 ,\AES_ENC/us30/n836 , \AES_ENC/us30/n835 , \AES_ENC/us30/n834 ,\AES_ENC/us30/n833 , \AES_ENC/us30/n832 , \AES_ENC/us30/n831 ,\AES_ENC/us30/n830 , \AES_ENC/us30/n829 , \AES_ENC/us30/n828 ,\AES_ENC/us30/n827 , \AES_ENC/us30/n826 , \AES_ENC/us30/n825 ,\AES_ENC/us30/n824 , \AES_ENC/us30/n823 , \AES_ENC/us30/n822 ,\AES_ENC/us30/n821 , \AES_ENC/us30/n820 , \AES_ENC/us30/n819 ,\AES_ENC/us30/n818 , \AES_ENC/us30/n817 , \AES_ENC/us30/n816 ,\AES_ENC/us30/n815 , \AES_ENC/us30/n814 , \AES_ENC/us30/n813 ,\AES_ENC/us30/n812 , \AES_ENC/us30/n811 , \AES_ENC/us30/n810 ,\AES_ENC/us30/n809 , \AES_ENC/us30/n808 , \AES_ENC/us30/n807 ,\AES_ENC/us30/n806 , \AES_ENC/us30/n805 , \AES_ENC/us30/n804 ,\AES_ENC/us30/n803 , \AES_ENC/us30/n802 , \AES_ENC/us30/n801 ,\AES_ENC/us30/n800 , \AES_ENC/us30/n799 , \AES_ENC/us30/n798 ,\AES_ENC/us30/n797 , \AES_ENC/us30/n796 , \AES_ENC/us30/n795 ,\AES_ENC/us30/n794 , \AES_ENC/us30/n793 , \AES_ENC/us30/n792 ,\AES_ENC/us30/n791 , \AES_ENC/us30/n790 , \AES_ENC/us30/n789 ,\AES_ENC/us30/n788 , \AES_ENC/us30/n787 , \AES_ENC/us30/n786 ,\AES_ENC/us30/n785 , \AES_ENC/us30/n784 , \AES_ENC/us30/n783 ,\AES_ENC/us30/n782 , \AES_ENC/us30/n781 , \AES_ENC/us30/n780 ,\AES_ENC/us30/n779 , \AES_ENC/us30/n778 , \AES_ENC/us30/n777 ,\AES_ENC/us30/n776 , \AES_ENC/us30/n775 , \AES_ENC/us30/n774 ,\AES_ENC/us30/n773 , \AES_ENC/us30/n772 , \AES_ENC/us30/n771 ,\AES_ENC/us30/n770 , \AES_ENC/us30/n769 , \AES_ENC/us30/n768 ,\AES_ENC/us30/n767 , \AES_ENC/us30/n766 , \AES_ENC/us30/n765 ,\AES_ENC/us30/n764 , \AES_ENC/us30/n763 , \AES_ENC/us30/n762 ,\AES_ENC/us30/n761 , \AES_ENC/us30/n760 , \AES_ENC/us30/n759 ,\AES_ENC/us30/n758 , \AES_ENC/us30/n757 , \AES_ENC/us30/n756 ,\AES_ENC/us30/n755 , \AES_ENC/us30/n754 , \AES_ENC/us30/n753 ,\AES_ENC/us30/n752 , \AES_ENC/us30/n751 , \AES_ENC/us30/n750 ,\AES_ENC/us30/n749 , \AES_ENC/us30/n748 , \AES_ENC/us30/n747 ,\AES_ENC/us30/n746 , \AES_ENC/us30/n745 , \AES_ENC/us30/n744 ,\AES_ENC/us30/n743 , \AES_ENC/us30/n742 , \AES_ENC/us30/n741 ,\AES_ENC/us30/n740 , \AES_ENC/us30/n739 , \AES_ENC/us30/n738 ,\AES_ENC/us30/n737 , \AES_ENC/us30/n736 , \AES_ENC/us30/n735 ,\AES_ENC/us30/n734 , \AES_ENC/us30/n733 , \AES_ENC/us30/n732 ,\AES_ENC/us30/n731 , \AES_ENC/us30/n730 , \AES_ENC/us30/n729 ,\AES_ENC/us30/n728 , \AES_ENC/us30/n727 , \AES_ENC/us30/n726 ,\AES_ENC/us30/n725 , \AES_ENC/us30/n724 , \AES_ENC/us30/n723 ,\AES_ENC/us30/n722 , \AES_ENC/us30/n721 , \AES_ENC/us30/n720 ,\AES_ENC/us30/n719 , \AES_ENC/us30/n718 , \AES_ENC/us30/n717 ,\AES_ENC/us30/n716 , \AES_ENC/us30/n715 , \AES_ENC/us30/n714 ,\AES_ENC/us30/n713 , \AES_ENC/us30/n712 , \AES_ENC/us30/n711 ,\AES_ENC/us30/n710 , \AES_ENC/us30/n709 , \AES_ENC/us30/n708 ,\AES_ENC/us30/n707 , \AES_ENC/us30/n706 , \AES_ENC/us30/n705 ,\AES_ENC/us30/n704 , \AES_ENC/us30/n703 , \AES_ENC/us30/n702 ,\AES_ENC/us30/n701 , \AES_ENC/us30/n700 , \AES_ENC/us30/n699 ,\AES_ENC/us30/n698 , \AES_ENC/us30/n697 , \AES_ENC/us30/n696 ,\AES_ENC/us30/n695 , \AES_ENC/us30/n694 , \AES_ENC/us30/n693 ,\AES_ENC/us30/n692 , \AES_ENC/us30/n691 , \AES_ENC/us30/n690 ,\AES_ENC/us30/n689 , \AES_ENC/us30/n688 , \AES_ENC/us30/n687 ,\AES_ENC/us30/n686 , \AES_ENC/us30/n685 , \AES_ENC/us30/n684 ,\AES_ENC/us30/n683 , \AES_ENC/us30/n682 , \AES_ENC/us30/n681 ,\AES_ENC/us30/n680 , \AES_ENC/us30/n679 , \AES_ENC/us30/n678 ,\AES_ENC/us30/n677 , \AES_ENC/us30/n676 , \AES_ENC/us30/n675 ,\AES_ENC/us30/n674 , \AES_ENC/us30/n673 , \AES_ENC/us30/n672 ,\AES_ENC/us30/n671 , \AES_ENC/us30/n670 , \AES_ENC/us30/n669 ,\AES_ENC/us30/n668 , \AES_ENC/us30/n667 , \AES_ENC/us30/n666 ,\AES_ENC/us30/n665 , \AES_ENC/us30/n664 , \AES_ENC/us30/n663 ,\AES_ENC/us30/n662 , \AES_ENC/us30/n661 , \AES_ENC/us30/n660 ,\AES_ENC/us30/n659 , \AES_ENC/us30/n658 , \AES_ENC/us30/n657 ,\AES_ENC/us30/n656 , \AES_ENC/us30/n655 , \AES_ENC/us30/n654 ,\AES_ENC/us30/n653 , \AES_ENC/us30/n652 , \AES_ENC/us30/n651 ,\AES_ENC/us30/n650 , \AES_ENC/us30/n649 , \AES_ENC/us30/n648 ,\AES_ENC/us30/n647 , \AES_ENC/us30/n646 , \AES_ENC/us30/n645 ,\AES_ENC/us30/n644 , \AES_ENC/us30/n643 , \AES_ENC/us30/n642 ,\AES_ENC/us30/n641 , \AES_ENC/us30/n640 , \AES_ENC/us30/n639 ,\AES_ENC/us30/n638 , \AES_ENC/us30/n637 , \AES_ENC/us30/n636 ,\AES_ENC/us30/n635 , \AES_ENC/us30/n634 , \AES_ENC/us30/n633 ,\AES_ENC/us30/n632 , \AES_ENC/us30/n631 , \AES_ENC/us30/n630 ,\AES_ENC/us30/n629 , \AES_ENC/us30/n628 , \AES_ENC/us30/n627 ,\AES_ENC/us30/n626 , \AES_ENC/us30/n625 , \AES_ENC/us30/n624 ,\AES_ENC/us30/n623 , \AES_ENC/us30/n622 , \AES_ENC/us30/n621 ,\AES_ENC/us30/n620 , \AES_ENC/us30/n619 , \AES_ENC/us30/n618 ,\AES_ENC/us30/n617 , \AES_ENC/us30/n616 , \AES_ENC/us30/n615 ,\AES_ENC/us30/n614 , \AES_ENC/us30/n613 , \AES_ENC/us30/n612 ,\AES_ENC/us30/n611 , \AES_ENC/us30/n610 , \AES_ENC/us30/n609 ,\AES_ENC/us30/n608 , \AES_ENC/us30/n607 , \AES_ENC/us30/n606 ,\AES_ENC/us30/n605 , \AES_ENC/us30/n604 , \AES_ENC/us30/n603 ,\AES_ENC/us30/n602 , \AES_ENC/us30/n601 , \AES_ENC/us30/n600 ,\AES_ENC/us30/n599 , \AES_ENC/us30/n598 , \AES_ENC/us30/n597 ,\AES_ENC/us30/n596 , \AES_ENC/us30/n595 , \AES_ENC/us30/n594 ,\AES_ENC/us30/n593 , \AES_ENC/us30/n592 , \AES_ENC/us30/n591 ,\AES_ENC/us30/n590 , \AES_ENC/us30/n589 , \AES_ENC/us30/n588 ,\AES_ENC/us30/n587 , \AES_ENC/us30/n586 , \AES_ENC/us30/n585 ,\AES_ENC/us30/n584 , \AES_ENC/us30/n583 , \AES_ENC/us30/n582 ,\AES_ENC/us30/n581 , \AES_ENC/us30/n580 , \AES_ENC/us30/n579 ,\AES_ENC/us30/n578 , \AES_ENC/us30/n577 , \AES_ENC/us30/n576 ,\AES_ENC/us30/n575 , \AES_ENC/us30/n574 , \AES_ENC/us30/n573 ,\AES_ENC/us30/n572 , \AES_ENC/us30/n571 , \AES_ENC/us30/n570 ,\AES_ENC/us30/n569 , \AES_ENC/us31/n1135 , \AES_ENC/us31/n1134 ,\AES_ENC/us31/n1133 , \AES_ENC/us31/n1132 , \AES_ENC/us31/n1131 ,\AES_ENC/us31/n1130 , \AES_ENC/us31/n1129 , \AES_ENC/us31/n1128 ,\AES_ENC/us31/n1127 , \AES_ENC/us31/n1126 , \AES_ENC/us31/n1125 ,\AES_ENC/us31/n1124 , \AES_ENC/us31/n1123 , \AES_ENC/us31/n1122 ,\AES_ENC/us31/n1121 , \AES_ENC/us31/n1120 , \AES_ENC/us31/n1119 ,\AES_ENC/us31/n1118 , \AES_ENC/us31/n1117 , \AES_ENC/us31/n1116 ,\AES_ENC/us31/n1115 , \AES_ENC/us31/n1114 , \AES_ENC/us31/n1113 ,\AES_ENC/us31/n1112 , \AES_ENC/us31/n1111 , \AES_ENC/us31/n1110 ,\AES_ENC/us31/n1109 , \AES_ENC/us31/n1108 , \AES_ENC/us31/n1107 ,\AES_ENC/us31/n1106 , \AES_ENC/us31/n1105 , \AES_ENC/us31/n1104 ,\AES_ENC/us31/n1103 , \AES_ENC/us31/n1102 , \AES_ENC/us31/n1101 ,\AES_ENC/us31/n1100 , \AES_ENC/us31/n1099 , \AES_ENC/us31/n1098 ,\AES_ENC/us31/n1097 , \AES_ENC/us31/n1096 , \AES_ENC/us31/n1095 ,\AES_ENC/us31/n1094 , \AES_ENC/us31/n1093 , \AES_ENC/us31/n1092 ,\AES_ENC/us31/n1091 , \AES_ENC/us31/n1090 , \AES_ENC/us31/n1089 ,\AES_ENC/us31/n1088 , \AES_ENC/us31/n1087 , \AES_ENC/us31/n1086 ,\AES_ENC/us31/n1085 , \AES_ENC/us31/n1084 , \AES_ENC/us31/n1083 ,\AES_ENC/us31/n1082 , \AES_ENC/us31/n1081 , \AES_ENC/us31/n1080 ,\AES_ENC/us31/n1079 , \AES_ENC/us31/n1078 , \AES_ENC/us31/n1077 ,\AES_ENC/us31/n1076 , \AES_ENC/us31/n1075 , \AES_ENC/us31/n1074 ,\AES_ENC/us31/n1073 , \AES_ENC/us31/n1072 , \AES_ENC/us31/n1071 ,\AES_ENC/us31/n1070 , \AES_ENC/us31/n1069 , \AES_ENC/us31/n1068 ,\AES_ENC/us31/n1067 , \AES_ENC/us31/n1066 , \AES_ENC/us31/n1065 ,\AES_ENC/us31/n1064 , \AES_ENC/us31/n1063 , \AES_ENC/us31/n1062 ,\AES_ENC/us31/n1061 , \AES_ENC/us31/n1060 , \AES_ENC/us31/n1059 ,\AES_ENC/us31/n1058 , \AES_ENC/us31/n1057 , \AES_ENC/us31/n1056 ,\AES_ENC/us31/n1055 , \AES_ENC/us31/n1054 , \AES_ENC/us31/n1053 ,\AES_ENC/us31/n1052 , \AES_ENC/us31/n1051 , \AES_ENC/us31/n1050 ,\AES_ENC/us31/n1049 , \AES_ENC/us31/n1048 , \AES_ENC/us31/n1047 ,\AES_ENC/us31/n1046 , \AES_ENC/us31/n1045 , \AES_ENC/us31/n1044 ,\AES_ENC/us31/n1043 , \AES_ENC/us31/n1042 , \AES_ENC/us31/n1041 ,\AES_ENC/us31/n1040 , \AES_ENC/us31/n1039 , \AES_ENC/us31/n1038 ,\AES_ENC/us31/n1037 , \AES_ENC/us31/n1036 , \AES_ENC/us31/n1035 ,\AES_ENC/us31/n1034 , \AES_ENC/us31/n1033 , \AES_ENC/us31/n1032 ,\AES_ENC/us31/n1031 , \AES_ENC/us31/n1030 , \AES_ENC/us31/n1029 ,\AES_ENC/us31/n1028 , \AES_ENC/us31/n1027 , \AES_ENC/us31/n1026 ,\AES_ENC/us31/n1025 , \AES_ENC/us31/n1024 , \AES_ENC/us31/n1023 ,\AES_ENC/us31/n1022 , \AES_ENC/us31/n1021 , \AES_ENC/us31/n1020 ,\AES_ENC/us31/n1019 , \AES_ENC/us31/n1018 , \AES_ENC/us31/n1017 ,\AES_ENC/us31/n1016 , \AES_ENC/us31/n1015 , \AES_ENC/us31/n1014 ,\AES_ENC/us31/n1013 , \AES_ENC/us31/n1012 , \AES_ENC/us31/n1011 ,\AES_ENC/us31/n1010 , \AES_ENC/us31/n1009 , \AES_ENC/us31/n1008 ,\AES_ENC/us31/n1007 , \AES_ENC/us31/n1006 , \AES_ENC/us31/n1005 ,\AES_ENC/us31/n1004 , \AES_ENC/us31/n1003 , \AES_ENC/us31/n1002 ,\AES_ENC/us31/n1001 , \AES_ENC/us31/n1000 , \AES_ENC/us31/n999 ,\AES_ENC/us31/n998 , \AES_ENC/us31/n997 , \AES_ENC/us31/n996 ,\AES_ENC/us31/n995 , \AES_ENC/us31/n994 , \AES_ENC/us31/n993 ,\AES_ENC/us31/n992 , \AES_ENC/us31/n991 , \AES_ENC/us31/n990 ,\AES_ENC/us31/n989 , \AES_ENC/us31/n988 , \AES_ENC/us31/n987 ,\AES_ENC/us31/n986 , \AES_ENC/us31/n985 , \AES_ENC/us31/n984 ,\AES_ENC/us31/n983 , \AES_ENC/us31/n982 , \AES_ENC/us31/n981 ,\AES_ENC/us31/n980 , \AES_ENC/us31/n979 , \AES_ENC/us31/n978 ,\AES_ENC/us31/n977 , \AES_ENC/us31/n976 , \AES_ENC/us31/n975 ,\AES_ENC/us31/n974 , \AES_ENC/us31/n973 , \AES_ENC/us31/n972 ,\AES_ENC/us31/n971 , \AES_ENC/us31/n970 , \AES_ENC/us31/n969 ,\AES_ENC/us31/n968 , \AES_ENC/us31/n967 , \AES_ENC/us31/n966 ,\AES_ENC/us31/n965 , \AES_ENC/us31/n964 , \AES_ENC/us31/n963 ,\AES_ENC/us31/n962 , \AES_ENC/us31/n961 , \AES_ENC/us31/n960 ,\AES_ENC/us31/n959 , \AES_ENC/us31/n958 , \AES_ENC/us31/n957 ,\AES_ENC/us31/n956 , \AES_ENC/us31/n955 , \AES_ENC/us31/n954 ,\AES_ENC/us31/n953 , \AES_ENC/us31/n952 , \AES_ENC/us31/n951 ,\AES_ENC/us31/n950 , \AES_ENC/us31/n949 , \AES_ENC/us31/n948 ,\AES_ENC/us31/n947 , \AES_ENC/us31/n946 , \AES_ENC/us31/n945 ,\AES_ENC/us31/n944 , \AES_ENC/us31/n943 , \AES_ENC/us31/n942 ,\AES_ENC/us31/n941 , \AES_ENC/us31/n940 , \AES_ENC/us31/n939 ,\AES_ENC/us31/n938 , \AES_ENC/us31/n937 , \AES_ENC/us31/n936 ,\AES_ENC/us31/n935 , \AES_ENC/us31/n934 , \AES_ENC/us31/n933 ,\AES_ENC/us31/n932 , \AES_ENC/us31/n931 , \AES_ENC/us31/n930 ,\AES_ENC/us31/n929 , \AES_ENC/us31/n928 , \AES_ENC/us31/n927 ,\AES_ENC/us31/n926 , \AES_ENC/us31/n925 , \AES_ENC/us31/n924 ,\AES_ENC/us31/n923 , \AES_ENC/us31/n922 , \AES_ENC/us31/n921 ,\AES_ENC/us31/n920 , \AES_ENC/us31/n919 , \AES_ENC/us31/n918 ,\AES_ENC/us31/n917 , \AES_ENC/us31/n916 , \AES_ENC/us31/n915 ,\AES_ENC/us31/n914 , \AES_ENC/us31/n913 , \AES_ENC/us31/n912 ,\AES_ENC/us31/n911 , \AES_ENC/us31/n910 , \AES_ENC/us31/n909 ,\AES_ENC/us31/n908 , \AES_ENC/us31/n907 , \AES_ENC/us31/n906 ,\AES_ENC/us31/n905 , \AES_ENC/us31/n904 , \AES_ENC/us31/n903 ,\AES_ENC/us31/n902 , \AES_ENC/us31/n901 , \AES_ENC/us31/n900 ,\AES_ENC/us31/n899 , \AES_ENC/us31/n898 , \AES_ENC/us31/n897 ,\AES_ENC/us31/n896 , \AES_ENC/us31/n895 , \AES_ENC/us31/n894 ,\AES_ENC/us31/n893 , \AES_ENC/us31/n892 , \AES_ENC/us31/n891 ,\AES_ENC/us31/n890 , \AES_ENC/us31/n889 , \AES_ENC/us31/n888 ,\AES_ENC/us31/n887 , \AES_ENC/us31/n886 , \AES_ENC/us31/n885 ,\AES_ENC/us31/n884 , \AES_ENC/us31/n883 , \AES_ENC/us31/n882 ,\AES_ENC/us31/n881 , \AES_ENC/us31/n880 , \AES_ENC/us31/n879 ,\AES_ENC/us31/n878 , \AES_ENC/us31/n877 , \AES_ENC/us31/n876 ,\AES_ENC/us31/n875 , \AES_ENC/us31/n874 , \AES_ENC/us31/n873 ,\AES_ENC/us31/n872 , \AES_ENC/us31/n871 , \AES_ENC/us31/n870 ,\AES_ENC/us31/n869 , \AES_ENC/us31/n868 , \AES_ENC/us31/n867 ,\AES_ENC/us31/n866 , \AES_ENC/us31/n865 , \AES_ENC/us31/n864 ,\AES_ENC/us31/n863 , \AES_ENC/us31/n862 , \AES_ENC/us31/n861 ,\AES_ENC/us31/n860 , \AES_ENC/us31/n859 , \AES_ENC/us31/n858 ,\AES_ENC/us31/n857 , \AES_ENC/us31/n856 , \AES_ENC/us31/n855 ,\AES_ENC/us31/n854 , \AES_ENC/us31/n853 , \AES_ENC/us31/n852 ,\AES_ENC/us31/n851 , \AES_ENC/us31/n850 , \AES_ENC/us31/n849 ,\AES_ENC/us31/n848 , \AES_ENC/us31/n847 , \AES_ENC/us31/n846 ,\AES_ENC/us31/n845 , \AES_ENC/us31/n844 , \AES_ENC/us31/n843 ,\AES_ENC/us31/n842 , \AES_ENC/us31/n841 , \AES_ENC/us31/n840 ,\AES_ENC/us31/n839 , \AES_ENC/us31/n838 , \AES_ENC/us31/n837 ,\AES_ENC/us31/n836 , \AES_ENC/us31/n835 , \AES_ENC/us31/n834 ,\AES_ENC/us31/n833 , \AES_ENC/us31/n832 , \AES_ENC/us31/n831 ,\AES_ENC/us31/n830 , \AES_ENC/us31/n829 , \AES_ENC/us31/n828 ,\AES_ENC/us31/n827 , \AES_ENC/us31/n826 , \AES_ENC/us31/n825 ,\AES_ENC/us31/n824 , \AES_ENC/us31/n823 , \AES_ENC/us31/n822 ,\AES_ENC/us31/n821 , \AES_ENC/us31/n820 , \AES_ENC/us31/n819 ,\AES_ENC/us31/n818 , \AES_ENC/us31/n817 , \AES_ENC/us31/n816 ,\AES_ENC/us31/n815 , \AES_ENC/us31/n814 , \AES_ENC/us31/n813 ,\AES_ENC/us31/n812 , \AES_ENC/us31/n811 , \AES_ENC/us31/n810 ,\AES_ENC/us31/n809 , \AES_ENC/us31/n808 , \AES_ENC/us31/n807 ,\AES_ENC/us31/n806 , \AES_ENC/us31/n805 , \AES_ENC/us31/n804 ,\AES_ENC/us31/n803 , \AES_ENC/us31/n802 , \AES_ENC/us31/n801 ,\AES_ENC/us31/n800 , \AES_ENC/us31/n799 , \AES_ENC/us31/n798 ,\AES_ENC/us31/n797 , \AES_ENC/us31/n796 , \AES_ENC/us31/n795 ,\AES_ENC/us31/n794 , \AES_ENC/us31/n793 , \AES_ENC/us31/n792 ,\AES_ENC/us31/n791 , \AES_ENC/us31/n790 , \AES_ENC/us31/n789 ,\AES_ENC/us31/n788 , \AES_ENC/us31/n787 , \AES_ENC/us31/n786 ,\AES_ENC/us31/n785 , \AES_ENC/us31/n784 , \AES_ENC/us31/n783 ,\AES_ENC/us31/n782 , \AES_ENC/us31/n781 , \AES_ENC/us31/n780 ,\AES_ENC/us31/n779 , \AES_ENC/us31/n778 , \AES_ENC/us31/n777 ,\AES_ENC/us31/n776 , \AES_ENC/us31/n775 , \AES_ENC/us31/n774 ,\AES_ENC/us31/n773 , \AES_ENC/us31/n772 , \AES_ENC/us31/n771 ,\AES_ENC/us31/n770 , \AES_ENC/us31/n769 , \AES_ENC/us31/n768 ,\AES_ENC/us31/n767 , \AES_ENC/us31/n766 , \AES_ENC/us31/n765 ,\AES_ENC/us31/n764 , \AES_ENC/us31/n763 , \AES_ENC/us31/n762 ,\AES_ENC/us31/n761 , \AES_ENC/us31/n760 , \AES_ENC/us31/n759 ,\AES_ENC/us31/n758 , \AES_ENC/us31/n757 , \AES_ENC/us31/n756 ,\AES_ENC/us31/n755 , \AES_ENC/us31/n754 , \AES_ENC/us31/n753 ,\AES_ENC/us31/n752 , \AES_ENC/us31/n751 , \AES_ENC/us31/n750 ,\AES_ENC/us31/n749 , \AES_ENC/us31/n748 , \AES_ENC/us31/n747 ,\AES_ENC/us31/n746 , \AES_ENC/us31/n745 , \AES_ENC/us31/n744 ,\AES_ENC/us31/n743 , \AES_ENC/us31/n742 , \AES_ENC/us31/n741 ,\AES_ENC/us31/n740 , \AES_ENC/us31/n739 , \AES_ENC/us31/n738 ,\AES_ENC/us31/n737 , \AES_ENC/us31/n736 , \AES_ENC/us31/n735 ,\AES_ENC/us31/n734 , \AES_ENC/us31/n733 , \AES_ENC/us31/n732 ,\AES_ENC/us31/n731 , \AES_ENC/us31/n730 , \AES_ENC/us31/n729 ,\AES_ENC/us31/n728 , \AES_ENC/us31/n727 , \AES_ENC/us31/n726 ,\AES_ENC/us31/n725 , \AES_ENC/us31/n724 , \AES_ENC/us31/n723 ,\AES_ENC/us31/n722 , \AES_ENC/us31/n721 , \AES_ENC/us31/n720 ,\AES_ENC/us31/n719 , \AES_ENC/us31/n718 , \AES_ENC/us31/n717 ,\AES_ENC/us31/n716 , \AES_ENC/us31/n715 , \AES_ENC/us31/n714 ,\AES_ENC/us31/n713 , \AES_ENC/us31/n712 , \AES_ENC/us31/n711 ,\AES_ENC/us31/n710 , \AES_ENC/us31/n709 , \AES_ENC/us31/n708 ,\AES_ENC/us31/n707 , \AES_ENC/us31/n706 , \AES_ENC/us31/n705 ,\AES_ENC/us31/n704 , \AES_ENC/us31/n703 , \AES_ENC/us31/n702 ,\AES_ENC/us31/n701 , \AES_ENC/us31/n700 , \AES_ENC/us31/n699 ,\AES_ENC/us31/n698 , \AES_ENC/us31/n697 , \AES_ENC/us31/n696 ,\AES_ENC/us31/n695 , \AES_ENC/us31/n694 , \AES_ENC/us31/n693 ,\AES_ENC/us31/n692 , \AES_ENC/us31/n691 , \AES_ENC/us31/n690 ,\AES_ENC/us31/n689 , \AES_ENC/us31/n688 , \AES_ENC/us31/n687 ,\AES_ENC/us31/n686 , \AES_ENC/us31/n685 , \AES_ENC/us31/n684 ,\AES_ENC/us31/n683 , \AES_ENC/us31/n682 , \AES_ENC/us31/n681 ,\AES_ENC/us31/n680 , \AES_ENC/us31/n679 , \AES_ENC/us31/n678 ,\AES_ENC/us31/n677 , \AES_ENC/us31/n676 , \AES_ENC/us31/n675 ,\AES_ENC/us31/n674 , \AES_ENC/us31/n673 , \AES_ENC/us31/n672 ,\AES_ENC/us31/n671 , \AES_ENC/us31/n670 , \AES_ENC/us31/n669 ,\AES_ENC/us31/n668 , \AES_ENC/us31/n667 , \AES_ENC/us31/n666 ,\AES_ENC/us31/n665 , \AES_ENC/us31/n664 , \AES_ENC/us31/n663 ,\AES_ENC/us31/n662 , \AES_ENC/us31/n661 , \AES_ENC/us31/n660 ,\AES_ENC/us31/n659 , \AES_ENC/us31/n658 , \AES_ENC/us31/n657 ,\AES_ENC/us31/n656 , \AES_ENC/us31/n655 , \AES_ENC/us31/n654 ,\AES_ENC/us31/n653 , \AES_ENC/us31/n652 , \AES_ENC/us31/n651 ,\AES_ENC/us31/n650 , \AES_ENC/us31/n649 , \AES_ENC/us31/n648 ,\AES_ENC/us31/n647 , \AES_ENC/us31/n646 , \AES_ENC/us31/n645 ,\AES_ENC/us31/n644 , \AES_ENC/us31/n643 , \AES_ENC/us31/n642 ,\AES_ENC/us31/n641 , \AES_ENC/us31/n640 , \AES_ENC/us31/n639 ,\AES_ENC/us31/n638 , \AES_ENC/us31/n637 , \AES_ENC/us31/n636 ,\AES_ENC/us31/n635 , \AES_ENC/us31/n634 , \AES_ENC/us31/n633 ,\AES_ENC/us31/n632 , \AES_ENC/us31/n631 , \AES_ENC/us31/n630 ,\AES_ENC/us31/n629 , \AES_ENC/us31/n628 , \AES_ENC/us31/n627 ,\AES_ENC/us31/n626 , \AES_ENC/us31/n625 , \AES_ENC/us31/n624 ,\AES_ENC/us31/n623 , \AES_ENC/us31/n622 , \AES_ENC/us31/n621 ,\AES_ENC/us31/n620 , \AES_ENC/us31/n619 , \AES_ENC/us31/n618 ,\AES_ENC/us31/n617 , \AES_ENC/us31/n616 , \AES_ENC/us31/n615 ,\AES_ENC/us31/n614 , \AES_ENC/us31/n613 , \AES_ENC/us31/n612 ,\AES_ENC/us31/n611 , \AES_ENC/us31/n610 , \AES_ENC/us31/n609 ,\AES_ENC/us31/n608 , \AES_ENC/us31/n607 , \AES_ENC/us31/n606 ,\AES_ENC/us31/n605 , \AES_ENC/us31/n604 , \AES_ENC/us31/n603 ,\AES_ENC/us31/n602 , \AES_ENC/us31/n601 , \AES_ENC/us31/n600 ,\AES_ENC/us31/n599 , \AES_ENC/us31/n598 , \AES_ENC/us31/n597 ,\AES_ENC/us31/n596 , \AES_ENC/us31/n595 , \AES_ENC/us31/n594 ,\AES_ENC/us31/n593 , \AES_ENC/us31/n592 , \AES_ENC/us31/n591 ,\AES_ENC/us31/n590 , \AES_ENC/us31/n589 , \AES_ENC/us31/n588 ,\AES_ENC/us31/n587 , \AES_ENC/us31/n586 , \AES_ENC/us31/n585 ,\AES_ENC/us31/n584 , \AES_ENC/us31/n583 , \AES_ENC/us31/n582 ,\AES_ENC/us31/n581 , \AES_ENC/us31/n580 , \AES_ENC/us31/n579 ,\AES_ENC/us31/n578 , \AES_ENC/us31/n577 , \AES_ENC/us31/n576 ,\AES_ENC/us31/n575 , \AES_ENC/us31/n574 , \AES_ENC/us31/n573 ,\AES_ENC/us31/n572 , \AES_ENC/us31/n571 , \AES_ENC/us31/n570 ,\AES_ENC/us31/n569 , \AES_ENC/us32/n1135 , \AES_ENC/us32/n1134 ,\AES_ENC/us32/n1133 , \AES_ENC/us32/n1132 , \AES_ENC/us32/n1131 ,\AES_ENC/us32/n1130 , \AES_ENC/us32/n1129 , \AES_ENC/us32/n1128 ,\AES_ENC/us32/n1127 , \AES_ENC/us32/n1126 , \AES_ENC/us32/n1125 ,\AES_ENC/us32/n1124 , \AES_ENC/us32/n1123 , \AES_ENC/us32/n1122 ,\AES_ENC/us32/n1121 , \AES_ENC/us32/n1120 , \AES_ENC/us32/n1119 ,\AES_ENC/us32/n1118 , \AES_ENC/us32/n1117 , \AES_ENC/us32/n1116 ,\AES_ENC/us32/n1115 , \AES_ENC/us32/n1114 , \AES_ENC/us32/n1113 ,\AES_ENC/us32/n1112 , \AES_ENC/us32/n1111 , \AES_ENC/us32/n1110 ,\AES_ENC/us32/n1109 , \AES_ENC/us32/n1108 , \AES_ENC/us32/n1107 ,\AES_ENC/us32/n1106 , \AES_ENC/us32/n1105 , \AES_ENC/us32/n1104 ,\AES_ENC/us32/n1103 , \AES_ENC/us32/n1102 , \AES_ENC/us32/n1101 ,\AES_ENC/us32/n1100 , \AES_ENC/us32/n1099 , \AES_ENC/us32/n1098 ,\AES_ENC/us32/n1097 , \AES_ENC/us32/n1096 , \AES_ENC/us32/n1095 ,\AES_ENC/us32/n1094 , \AES_ENC/us32/n1093 , \AES_ENC/us32/n1092 ,\AES_ENC/us32/n1091 , \AES_ENC/us32/n1090 , \AES_ENC/us32/n1089 ,\AES_ENC/us32/n1088 , \AES_ENC/us32/n1087 , \AES_ENC/us32/n1086 ,\AES_ENC/us32/n1085 , \AES_ENC/us32/n1084 , \AES_ENC/us32/n1083 ,\AES_ENC/us32/n1082 , \AES_ENC/us32/n1081 , \AES_ENC/us32/n1080 ,\AES_ENC/us32/n1079 , \AES_ENC/us32/n1078 , \AES_ENC/us32/n1077 ,\AES_ENC/us32/n1076 , \AES_ENC/us32/n1075 , \AES_ENC/us32/n1074 ,\AES_ENC/us32/n1073 , \AES_ENC/us32/n1072 , \AES_ENC/us32/n1071 ,\AES_ENC/us32/n1070 , \AES_ENC/us32/n1069 , \AES_ENC/us32/n1068 ,\AES_ENC/us32/n1067 , \AES_ENC/us32/n1066 , \AES_ENC/us32/n1065 ,\AES_ENC/us32/n1064 , \AES_ENC/us32/n1063 , \AES_ENC/us32/n1062 ,\AES_ENC/us32/n1061 , \AES_ENC/us32/n1060 , \AES_ENC/us32/n1059 ,\AES_ENC/us32/n1058 , \AES_ENC/us32/n1057 , \AES_ENC/us32/n1056 ,\AES_ENC/us32/n1055 , \AES_ENC/us32/n1054 , \AES_ENC/us32/n1053 ,\AES_ENC/us32/n1052 , \AES_ENC/us32/n1051 , \AES_ENC/us32/n1050 ,\AES_ENC/us32/n1049 , \AES_ENC/us32/n1048 , \AES_ENC/us32/n1047 ,\AES_ENC/us32/n1046 , \AES_ENC/us32/n1045 , \AES_ENC/us32/n1044 ,\AES_ENC/us32/n1043 , \AES_ENC/us32/n1042 , \AES_ENC/us32/n1041 ,\AES_ENC/us32/n1040 , \AES_ENC/us32/n1039 , \AES_ENC/us32/n1038 ,\AES_ENC/us32/n1037 , \AES_ENC/us32/n1036 , \AES_ENC/us32/n1035 ,\AES_ENC/us32/n1034 , \AES_ENC/us32/n1033 , \AES_ENC/us32/n1032 ,\AES_ENC/us32/n1031 , \AES_ENC/us32/n1030 , \AES_ENC/us32/n1029 ,\AES_ENC/us32/n1028 , \AES_ENC/us32/n1027 , \AES_ENC/us32/n1026 ,\AES_ENC/us32/n1025 , \AES_ENC/us32/n1024 , \AES_ENC/us32/n1023 ,\AES_ENC/us32/n1022 , \AES_ENC/us32/n1021 , \AES_ENC/us32/n1020 ,\AES_ENC/us32/n1019 , \AES_ENC/us32/n1018 , \AES_ENC/us32/n1017 ,\AES_ENC/us32/n1016 , \AES_ENC/us32/n1015 , \AES_ENC/us32/n1014 ,\AES_ENC/us32/n1013 , \AES_ENC/us32/n1012 , \AES_ENC/us32/n1011 ,\AES_ENC/us32/n1010 , \AES_ENC/us32/n1009 , \AES_ENC/us32/n1008 ,\AES_ENC/us32/n1007 , \AES_ENC/us32/n1006 , \AES_ENC/us32/n1005 ,\AES_ENC/us32/n1004 , \AES_ENC/us32/n1003 , \AES_ENC/us32/n1002 ,\AES_ENC/us32/n1001 , \AES_ENC/us32/n1000 , \AES_ENC/us32/n999 ,\AES_ENC/us32/n998 , \AES_ENC/us32/n997 , \AES_ENC/us32/n996 ,\AES_ENC/us32/n995 , \AES_ENC/us32/n994 , \AES_ENC/us32/n993 ,\AES_ENC/us32/n992 , \AES_ENC/us32/n991 , \AES_ENC/us32/n990 ,\AES_ENC/us32/n989 , \AES_ENC/us32/n988 , \AES_ENC/us32/n987 ,\AES_ENC/us32/n986 , \AES_ENC/us32/n985 , \AES_ENC/us32/n984 ,\AES_ENC/us32/n983 , \AES_ENC/us32/n982 , \AES_ENC/us32/n981 ,\AES_ENC/us32/n980 , \AES_ENC/us32/n979 , \AES_ENC/us32/n978 ,\AES_ENC/us32/n977 , \AES_ENC/us32/n976 , \AES_ENC/us32/n975 ,\AES_ENC/us32/n974 , \AES_ENC/us32/n973 , \AES_ENC/us32/n972 ,\AES_ENC/us32/n971 , \AES_ENC/us32/n970 , \AES_ENC/us32/n969 ,\AES_ENC/us32/n968 , \AES_ENC/us32/n967 , \AES_ENC/us32/n966 ,\AES_ENC/us32/n965 , \AES_ENC/us32/n964 , \AES_ENC/us32/n963 ,\AES_ENC/us32/n962 , \AES_ENC/us32/n961 , \AES_ENC/us32/n960 ,\AES_ENC/us32/n959 , \AES_ENC/us32/n958 , \AES_ENC/us32/n957 ,\AES_ENC/us32/n956 , \AES_ENC/us32/n955 , \AES_ENC/us32/n954 ,\AES_ENC/us32/n953 , \AES_ENC/us32/n952 , \AES_ENC/us32/n951 ,\AES_ENC/us32/n950 , \AES_ENC/us32/n949 , \AES_ENC/us32/n948 ,\AES_ENC/us32/n947 , \AES_ENC/us32/n946 , \AES_ENC/us32/n945 ,\AES_ENC/us32/n944 , \AES_ENC/us32/n943 , \AES_ENC/us32/n942 ,\AES_ENC/us32/n941 , \AES_ENC/us32/n940 , \AES_ENC/us32/n939 ,\AES_ENC/us32/n938 , \AES_ENC/us32/n937 , \AES_ENC/us32/n936 ,\AES_ENC/us32/n935 , \AES_ENC/us32/n934 , \AES_ENC/us32/n933 ,\AES_ENC/us32/n932 , \AES_ENC/us32/n931 , \AES_ENC/us32/n930 ,\AES_ENC/us32/n929 , \AES_ENC/us32/n928 , \AES_ENC/us32/n927 ,\AES_ENC/us32/n926 , \AES_ENC/us32/n925 , \AES_ENC/us32/n924 ,\AES_ENC/us32/n923 , \AES_ENC/us32/n922 , \AES_ENC/us32/n921 ,\AES_ENC/us32/n920 , \AES_ENC/us32/n919 , \AES_ENC/us32/n918 ,\AES_ENC/us32/n917 , \AES_ENC/us32/n916 , \AES_ENC/us32/n915 ,\AES_ENC/us32/n914 , \AES_ENC/us32/n913 , \AES_ENC/us32/n912 ,\AES_ENC/us32/n911 , \AES_ENC/us32/n910 , \AES_ENC/us32/n909 ,\AES_ENC/us32/n908 , \AES_ENC/us32/n907 , \AES_ENC/us32/n906 ,\AES_ENC/us32/n905 , \AES_ENC/us32/n904 , \AES_ENC/us32/n903 ,\AES_ENC/us32/n902 , \AES_ENC/us32/n901 , \AES_ENC/us32/n900 ,\AES_ENC/us32/n899 , \AES_ENC/us32/n898 , \AES_ENC/us32/n897 ,\AES_ENC/us32/n896 , \AES_ENC/us32/n895 , \AES_ENC/us32/n894 ,\AES_ENC/us32/n893 , \AES_ENC/us32/n892 , \AES_ENC/us32/n891 ,\AES_ENC/us32/n890 , \AES_ENC/us32/n889 , \AES_ENC/us32/n888 ,\AES_ENC/us32/n887 , \AES_ENC/us32/n886 , \AES_ENC/us32/n885 ,\AES_ENC/us32/n884 , \AES_ENC/us32/n883 , \AES_ENC/us32/n882 ,\AES_ENC/us32/n881 , \AES_ENC/us32/n880 , \AES_ENC/us32/n879 ,\AES_ENC/us32/n878 , \AES_ENC/us32/n877 , \AES_ENC/us32/n876 ,\AES_ENC/us32/n875 , \AES_ENC/us32/n874 , \AES_ENC/us32/n873 ,\AES_ENC/us32/n872 , \AES_ENC/us32/n871 , \AES_ENC/us32/n870 ,\AES_ENC/us32/n869 , \AES_ENC/us32/n868 , \AES_ENC/us32/n867 ,\AES_ENC/us32/n866 , \AES_ENC/us32/n865 , \AES_ENC/us32/n864 ,\AES_ENC/us32/n863 , \AES_ENC/us32/n862 , \AES_ENC/us32/n861 ,\AES_ENC/us32/n860 , \AES_ENC/us32/n859 , \AES_ENC/us32/n858 ,\AES_ENC/us32/n857 , \AES_ENC/us32/n856 , \AES_ENC/us32/n855 ,\AES_ENC/us32/n854 , \AES_ENC/us32/n853 , \AES_ENC/us32/n852 ,\AES_ENC/us32/n851 , \AES_ENC/us32/n850 , \AES_ENC/us32/n849 ,\AES_ENC/us32/n848 , \AES_ENC/us32/n847 , \AES_ENC/us32/n846 ,\AES_ENC/us32/n845 , \AES_ENC/us32/n844 , \AES_ENC/us32/n843 ,\AES_ENC/us32/n842 , \AES_ENC/us32/n841 , \AES_ENC/us32/n840 ,\AES_ENC/us32/n839 , \AES_ENC/us32/n838 , \AES_ENC/us32/n837 ,\AES_ENC/us32/n836 , \AES_ENC/us32/n835 , \AES_ENC/us32/n834 ,\AES_ENC/us32/n833 , \AES_ENC/us32/n832 , \AES_ENC/us32/n831 ,\AES_ENC/us32/n830 , \AES_ENC/us32/n829 , \AES_ENC/us32/n828 ,\AES_ENC/us32/n827 , \AES_ENC/us32/n826 , \AES_ENC/us32/n825 ,\AES_ENC/us32/n824 , \AES_ENC/us32/n823 , \AES_ENC/us32/n822 ,\AES_ENC/us32/n821 , \AES_ENC/us32/n820 , \AES_ENC/us32/n819 ,\AES_ENC/us32/n818 , \AES_ENC/us32/n817 , \AES_ENC/us32/n816 ,\AES_ENC/us32/n815 , \AES_ENC/us32/n814 , \AES_ENC/us32/n813 ,\AES_ENC/us32/n812 , \AES_ENC/us32/n811 , \AES_ENC/us32/n810 ,\AES_ENC/us32/n809 , \AES_ENC/us32/n808 , \AES_ENC/us32/n807 ,\AES_ENC/us32/n806 , \AES_ENC/us32/n805 , \AES_ENC/us32/n804 ,\AES_ENC/us32/n803 , \AES_ENC/us32/n802 , \AES_ENC/us32/n801 ,\AES_ENC/us32/n800 , \AES_ENC/us32/n799 , \AES_ENC/us32/n798 ,\AES_ENC/us32/n797 , \AES_ENC/us32/n796 , \AES_ENC/us32/n795 ,\AES_ENC/us32/n794 , \AES_ENC/us32/n793 , \AES_ENC/us32/n792 ,\AES_ENC/us32/n791 , \AES_ENC/us32/n790 , \AES_ENC/us32/n789 ,\AES_ENC/us32/n788 , \AES_ENC/us32/n787 , \AES_ENC/us32/n786 ,\AES_ENC/us32/n785 , \AES_ENC/us32/n784 , \AES_ENC/us32/n783 ,\AES_ENC/us32/n782 , \AES_ENC/us32/n781 , \AES_ENC/us32/n780 ,\AES_ENC/us32/n779 , \AES_ENC/us32/n778 , \AES_ENC/us32/n777 ,\AES_ENC/us32/n776 , \AES_ENC/us32/n775 , \AES_ENC/us32/n774 ,\AES_ENC/us32/n773 , \AES_ENC/us32/n772 , \AES_ENC/us32/n771 ,\AES_ENC/us32/n770 , \AES_ENC/us32/n769 , \AES_ENC/us32/n768 ,\AES_ENC/us32/n767 , \AES_ENC/us32/n766 , \AES_ENC/us32/n765 ,\AES_ENC/us32/n764 , \AES_ENC/us32/n763 , \AES_ENC/us32/n762 ,\AES_ENC/us32/n761 , \AES_ENC/us32/n760 , \AES_ENC/us32/n759 ,\AES_ENC/us32/n758 , \AES_ENC/us32/n757 , \AES_ENC/us32/n756 ,\AES_ENC/us32/n755 , \AES_ENC/us32/n754 , \AES_ENC/us32/n753 ,\AES_ENC/us32/n752 , \AES_ENC/us32/n751 , \AES_ENC/us32/n750 ,\AES_ENC/us32/n749 , \AES_ENC/us32/n748 , \AES_ENC/us32/n747 ,\AES_ENC/us32/n746 , \AES_ENC/us32/n745 , \AES_ENC/us32/n744 ,\AES_ENC/us32/n743 , \AES_ENC/us32/n742 , \AES_ENC/us32/n741 ,\AES_ENC/us32/n740 , \AES_ENC/us32/n739 , \AES_ENC/us32/n738 ,\AES_ENC/us32/n737 , \AES_ENC/us32/n736 , \AES_ENC/us32/n735 ,\AES_ENC/us32/n734 , \AES_ENC/us32/n733 , \AES_ENC/us32/n732 ,\AES_ENC/us32/n731 , \AES_ENC/us32/n730 , \AES_ENC/us32/n729 ,\AES_ENC/us32/n728 , \AES_ENC/us32/n727 , \AES_ENC/us32/n726 ,\AES_ENC/us32/n725 , \AES_ENC/us32/n724 , \AES_ENC/us32/n723 ,\AES_ENC/us32/n722 , \AES_ENC/us32/n721 , \AES_ENC/us32/n720 ,\AES_ENC/us32/n719 , \AES_ENC/us32/n718 , \AES_ENC/us32/n717 ,\AES_ENC/us32/n716 , \AES_ENC/us32/n715 , \AES_ENC/us32/n714 ,\AES_ENC/us32/n713 , \AES_ENC/us32/n712 , \AES_ENC/us32/n711 ,\AES_ENC/us32/n710 , \AES_ENC/us32/n709 , \AES_ENC/us32/n708 ,\AES_ENC/us32/n707 , \AES_ENC/us32/n706 , \AES_ENC/us32/n705 ,\AES_ENC/us32/n704 , \AES_ENC/us32/n703 , \AES_ENC/us32/n702 ,\AES_ENC/us32/n701 , \AES_ENC/us32/n700 , \AES_ENC/us32/n699 ,\AES_ENC/us32/n698 , \AES_ENC/us32/n697 , \AES_ENC/us32/n696 ,\AES_ENC/us32/n695 , \AES_ENC/us32/n694 , \AES_ENC/us32/n693 ,\AES_ENC/us32/n692 , \AES_ENC/us32/n691 , \AES_ENC/us32/n690 ,\AES_ENC/us32/n689 , \AES_ENC/us32/n688 , \AES_ENC/us32/n687 ,\AES_ENC/us32/n686 , \AES_ENC/us32/n685 , \AES_ENC/us32/n684 ,\AES_ENC/us32/n683 , \AES_ENC/us32/n682 , \AES_ENC/us32/n681 ,\AES_ENC/us32/n680 , \AES_ENC/us32/n679 , \AES_ENC/us32/n678 ,\AES_ENC/us32/n677 , \AES_ENC/us32/n676 , \AES_ENC/us32/n675 ,\AES_ENC/us32/n674 , \AES_ENC/us32/n673 , \AES_ENC/us32/n672 ,\AES_ENC/us32/n671 , \AES_ENC/us32/n670 , \AES_ENC/us32/n669 ,\AES_ENC/us32/n668 , \AES_ENC/us32/n667 , \AES_ENC/us32/n666 ,\AES_ENC/us32/n665 , \AES_ENC/us32/n664 , \AES_ENC/us32/n663 ,\AES_ENC/us32/n662 , \AES_ENC/us32/n661 , \AES_ENC/us32/n660 ,\AES_ENC/us32/n659 , \AES_ENC/us32/n658 , \AES_ENC/us32/n657 ,\AES_ENC/us32/n656 , \AES_ENC/us32/n655 , \AES_ENC/us32/n654 ,\AES_ENC/us32/n653 , \AES_ENC/us32/n652 , \AES_ENC/us32/n651 ,\AES_ENC/us32/n650 , \AES_ENC/us32/n649 , \AES_ENC/us32/n648 ,\AES_ENC/us32/n647 , \AES_ENC/us32/n646 , \AES_ENC/us32/n645 ,\AES_ENC/us32/n644 , \AES_ENC/us32/n643 , \AES_ENC/us32/n642 ,\AES_ENC/us32/n641 , \AES_ENC/us32/n640 , \AES_ENC/us32/n639 ,\AES_ENC/us32/n638 , \AES_ENC/us32/n637 , \AES_ENC/us32/n636 ,\AES_ENC/us32/n635 , \AES_ENC/us32/n634 , \AES_ENC/us32/n633 ,\AES_ENC/us32/n632 , \AES_ENC/us32/n631 , \AES_ENC/us32/n630 ,\AES_ENC/us32/n629 , \AES_ENC/us32/n628 , \AES_ENC/us32/n627 ,\AES_ENC/us32/n626 , \AES_ENC/us32/n625 , \AES_ENC/us32/n624 ,\AES_ENC/us32/n623 , \AES_ENC/us32/n622 , \AES_ENC/us32/n621 ,\AES_ENC/us32/n620 , \AES_ENC/us32/n619 , \AES_ENC/us32/n618 ,\AES_ENC/us32/n617 , \AES_ENC/us32/n616 , \AES_ENC/us32/n615 ,\AES_ENC/us32/n614 , \AES_ENC/us32/n613 , \AES_ENC/us32/n612 ,\AES_ENC/us32/n611 , \AES_ENC/us32/n610 , \AES_ENC/us32/n609 ,\AES_ENC/us32/n608 , \AES_ENC/us32/n607 , \AES_ENC/us32/n606 ,\AES_ENC/us32/n605 , \AES_ENC/us32/n604 , \AES_ENC/us32/n603 ,\AES_ENC/us32/n602 , \AES_ENC/us32/n601 , \AES_ENC/us32/n600 ,\AES_ENC/us32/n599 , \AES_ENC/us32/n598 , \AES_ENC/us32/n597 ,\AES_ENC/us32/n596 , \AES_ENC/us32/n595 , \AES_ENC/us32/n594 ,\AES_ENC/us32/n593 , \AES_ENC/us32/n592 , \AES_ENC/us32/n591 ,\AES_ENC/us32/n590 , \AES_ENC/us32/n589 , \AES_ENC/us32/n588 ,\AES_ENC/us32/n587 , \AES_ENC/us32/n586 , \AES_ENC/us32/n585 ,\AES_ENC/us32/n584 , \AES_ENC/us32/n583 , \AES_ENC/us32/n582 ,\AES_ENC/us32/n581 , \AES_ENC/us32/n580 , \AES_ENC/us32/n579 ,\AES_ENC/us32/n578 , \AES_ENC/us32/n577 , \AES_ENC/us32/n576 ,\AES_ENC/us32/n575 , \AES_ENC/us32/n574 , \AES_ENC/us32/n573 ,\AES_ENC/us32/n572 , \AES_ENC/us32/n571 , \AES_ENC/us32/n570 ,\AES_ENC/us32/n569 , \AES_ENC/us33/n1135 , \AES_ENC/us33/n1134 ,\AES_ENC/us33/n1133 , \AES_ENC/us33/n1132 , \AES_ENC/us33/n1131 ,\AES_ENC/us33/n1130 , \AES_ENC/us33/n1129 , \AES_ENC/us33/n1128 ,\AES_ENC/us33/n1127 , \AES_ENC/us33/n1126 , \AES_ENC/us33/n1125 ,\AES_ENC/us33/n1124 , \AES_ENC/us33/n1123 , \AES_ENC/us33/n1122 ,\AES_ENC/us33/n1121 , \AES_ENC/us33/n1120 , \AES_ENC/us33/n1119 ,\AES_ENC/us33/n1118 , \AES_ENC/us33/n1117 , \AES_ENC/us33/n1116 ,\AES_ENC/us33/n1115 , \AES_ENC/us33/n1114 , \AES_ENC/us33/n1113 ,\AES_ENC/us33/n1112 , \AES_ENC/us33/n1111 , \AES_ENC/us33/n1110 ,\AES_ENC/us33/n1109 , \AES_ENC/us33/n1108 , \AES_ENC/us33/n1107 ,\AES_ENC/us33/n1106 , \AES_ENC/us33/n1105 , \AES_ENC/us33/n1104 ,\AES_ENC/us33/n1103 , \AES_ENC/us33/n1102 , \AES_ENC/us33/n1101 ,\AES_ENC/us33/n1100 , \AES_ENC/us33/n1099 , \AES_ENC/us33/n1098 ,\AES_ENC/us33/n1097 , \AES_ENC/us33/n1096 , \AES_ENC/us33/n1095 ,\AES_ENC/us33/n1094 , \AES_ENC/us33/n1093 , \AES_ENC/us33/n1092 ,\AES_ENC/us33/n1091 , \AES_ENC/us33/n1090 , \AES_ENC/us33/n1089 ,\AES_ENC/us33/n1088 , \AES_ENC/us33/n1087 , \AES_ENC/us33/n1086 ,\AES_ENC/us33/n1085 , \AES_ENC/us33/n1084 , \AES_ENC/us33/n1083 ,\AES_ENC/us33/n1082 , \AES_ENC/us33/n1081 , \AES_ENC/us33/n1080 ,\AES_ENC/us33/n1079 , \AES_ENC/us33/n1078 , \AES_ENC/us33/n1077 ,\AES_ENC/us33/n1076 , \AES_ENC/us33/n1075 , \AES_ENC/us33/n1074 ,\AES_ENC/us33/n1073 , \AES_ENC/us33/n1072 , \AES_ENC/us33/n1071 ,\AES_ENC/us33/n1070 , \AES_ENC/us33/n1069 , \AES_ENC/us33/n1068 ,\AES_ENC/us33/n1067 , \AES_ENC/us33/n1066 , \AES_ENC/us33/n1065 ,\AES_ENC/us33/n1064 , \AES_ENC/us33/n1063 , \AES_ENC/us33/n1062 ,\AES_ENC/us33/n1061 , \AES_ENC/us33/n1060 , \AES_ENC/us33/n1059 ,\AES_ENC/us33/n1058 , \AES_ENC/us33/n1057 , \AES_ENC/us33/n1056 ,\AES_ENC/us33/n1055 , \AES_ENC/us33/n1054 , \AES_ENC/us33/n1053 ,\AES_ENC/us33/n1052 , \AES_ENC/us33/n1051 , \AES_ENC/us33/n1050 ,\AES_ENC/us33/n1049 , \AES_ENC/us33/n1048 , \AES_ENC/us33/n1047 ,\AES_ENC/us33/n1046 , \AES_ENC/us33/n1045 , \AES_ENC/us33/n1044 ,\AES_ENC/us33/n1043 , \AES_ENC/us33/n1042 , \AES_ENC/us33/n1041 ,\AES_ENC/us33/n1040 , \AES_ENC/us33/n1039 , \AES_ENC/us33/n1038 ,\AES_ENC/us33/n1037 , \AES_ENC/us33/n1036 , \AES_ENC/us33/n1035 ,\AES_ENC/us33/n1034 , \AES_ENC/us33/n1033 , \AES_ENC/us33/n1032 ,\AES_ENC/us33/n1031 , \AES_ENC/us33/n1030 , \AES_ENC/us33/n1029 ,\AES_ENC/us33/n1028 , \AES_ENC/us33/n1027 , \AES_ENC/us33/n1026 ,\AES_ENC/us33/n1025 , \AES_ENC/us33/n1024 , \AES_ENC/us33/n1023 ,\AES_ENC/us33/n1022 , \AES_ENC/us33/n1021 , \AES_ENC/us33/n1020 ,\AES_ENC/us33/n1019 , \AES_ENC/us33/n1018 , \AES_ENC/us33/n1017 ,\AES_ENC/us33/n1016 , \AES_ENC/us33/n1015 , \AES_ENC/us33/n1014 ,\AES_ENC/us33/n1013 , \AES_ENC/us33/n1012 , \AES_ENC/us33/n1011 ,\AES_ENC/us33/n1010 , \AES_ENC/us33/n1009 , \AES_ENC/us33/n1008 ,\AES_ENC/us33/n1007 , \AES_ENC/us33/n1006 , \AES_ENC/us33/n1005 ,\AES_ENC/us33/n1004 , \AES_ENC/us33/n1003 , \AES_ENC/us33/n1002 ,\AES_ENC/us33/n1001 , \AES_ENC/us33/n1000 , \AES_ENC/us33/n999 ,\AES_ENC/us33/n998 , \AES_ENC/us33/n997 , \AES_ENC/us33/n996 ,\AES_ENC/us33/n995 , \AES_ENC/us33/n994 , \AES_ENC/us33/n993 ,\AES_ENC/us33/n992 , \AES_ENC/us33/n991 , \AES_ENC/us33/n990 ,\AES_ENC/us33/n989 , \AES_ENC/us33/n988 , \AES_ENC/us33/n987 ,\AES_ENC/us33/n986 , \AES_ENC/us33/n985 , \AES_ENC/us33/n984 ,\AES_ENC/us33/n983 , \AES_ENC/us33/n982 , \AES_ENC/us33/n981 ,\AES_ENC/us33/n980 , \AES_ENC/us33/n979 , \AES_ENC/us33/n978 ,\AES_ENC/us33/n977 , \AES_ENC/us33/n976 , \AES_ENC/us33/n975 ,\AES_ENC/us33/n974 , \AES_ENC/us33/n973 , \AES_ENC/us33/n972 ,\AES_ENC/us33/n971 , \AES_ENC/us33/n970 , \AES_ENC/us33/n969 ,\AES_ENC/us33/n968 , \AES_ENC/us33/n967 , \AES_ENC/us33/n966 ,\AES_ENC/us33/n965 , \AES_ENC/us33/n964 , \AES_ENC/us33/n963 ,\AES_ENC/us33/n962 , \AES_ENC/us33/n961 , \AES_ENC/us33/n960 ,\AES_ENC/us33/n959 , \AES_ENC/us33/n958 , \AES_ENC/us33/n957 ,\AES_ENC/us33/n956 , \AES_ENC/us33/n955 , \AES_ENC/us33/n954 ,\AES_ENC/us33/n953 , \AES_ENC/us33/n952 , \AES_ENC/us33/n951 ,\AES_ENC/us33/n950 , \AES_ENC/us33/n949 , \AES_ENC/us33/n948 ,\AES_ENC/us33/n947 , \AES_ENC/us33/n946 , \AES_ENC/us33/n945 ,\AES_ENC/us33/n944 , \AES_ENC/us33/n943 , \AES_ENC/us33/n942 ,\AES_ENC/us33/n941 , \AES_ENC/us33/n940 , \AES_ENC/us33/n939 ,\AES_ENC/us33/n938 , \AES_ENC/us33/n937 , \AES_ENC/us33/n936 ,\AES_ENC/us33/n935 , \AES_ENC/us33/n934 , \AES_ENC/us33/n933 ,\AES_ENC/us33/n932 , \AES_ENC/us33/n931 , \AES_ENC/us33/n930 ,\AES_ENC/us33/n929 , \AES_ENC/us33/n928 , \AES_ENC/us33/n927 ,\AES_ENC/us33/n926 , \AES_ENC/us33/n925 , \AES_ENC/us33/n924 ,\AES_ENC/us33/n923 , \AES_ENC/us33/n922 , \AES_ENC/us33/n921 ,\AES_ENC/us33/n920 , \AES_ENC/us33/n919 , \AES_ENC/us33/n918 ,\AES_ENC/us33/n917 , \AES_ENC/us33/n916 , \AES_ENC/us33/n915 ,\AES_ENC/us33/n914 , \AES_ENC/us33/n913 , \AES_ENC/us33/n912 ,\AES_ENC/us33/n911 , \AES_ENC/us33/n910 , \AES_ENC/us33/n909 ,\AES_ENC/us33/n908 , \AES_ENC/us33/n907 , \AES_ENC/us33/n906 ,\AES_ENC/us33/n905 , \AES_ENC/us33/n904 , \AES_ENC/us33/n903 ,\AES_ENC/us33/n902 , \AES_ENC/us33/n901 , \AES_ENC/us33/n900 ,\AES_ENC/us33/n899 , \AES_ENC/us33/n898 , \AES_ENC/us33/n897 ,\AES_ENC/us33/n896 , \AES_ENC/us33/n895 , \AES_ENC/us33/n894 ,\AES_ENC/us33/n893 , \AES_ENC/us33/n892 , \AES_ENC/us33/n891 ,\AES_ENC/us33/n890 , \AES_ENC/us33/n889 , \AES_ENC/us33/n888 ,\AES_ENC/us33/n887 , \AES_ENC/us33/n886 , \AES_ENC/us33/n885 ,\AES_ENC/us33/n884 , \AES_ENC/us33/n883 , \AES_ENC/us33/n882 ,\AES_ENC/us33/n881 , \AES_ENC/us33/n880 , \AES_ENC/us33/n879 ,\AES_ENC/us33/n878 , \AES_ENC/us33/n877 , \AES_ENC/us33/n876 ,\AES_ENC/us33/n875 , \AES_ENC/us33/n874 , \AES_ENC/us33/n873 ,\AES_ENC/us33/n872 , \AES_ENC/us33/n871 , \AES_ENC/us33/n870 ,\AES_ENC/us33/n869 , \AES_ENC/us33/n868 , \AES_ENC/us33/n867 ,\AES_ENC/us33/n866 , \AES_ENC/us33/n865 , \AES_ENC/us33/n864 ,\AES_ENC/us33/n863 , \AES_ENC/us33/n862 , \AES_ENC/us33/n861 ,\AES_ENC/us33/n860 , \AES_ENC/us33/n859 , \AES_ENC/us33/n858 ,\AES_ENC/us33/n857 , \AES_ENC/us33/n856 , \AES_ENC/us33/n855 ,\AES_ENC/us33/n854 , \AES_ENC/us33/n853 , \AES_ENC/us33/n852 ,\AES_ENC/us33/n851 , \AES_ENC/us33/n850 , \AES_ENC/us33/n849 ,\AES_ENC/us33/n848 , \AES_ENC/us33/n847 , \AES_ENC/us33/n846 ,\AES_ENC/us33/n845 , \AES_ENC/us33/n844 , \AES_ENC/us33/n843 ,\AES_ENC/us33/n842 , \AES_ENC/us33/n841 , \AES_ENC/us33/n840 ,\AES_ENC/us33/n839 , \AES_ENC/us33/n838 , \AES_ENC/us33/n837 ,\AES_ENC/us33/n836 , \AES_ENC/us33/n835 , \AES_ENC/us33/n834 ,\AES_ENC/us33/n833 , \AES_ENC/us33/n832 , \AES_ENC/us33/n831 ,\AES_ENC/us33/n830 , \AES_ENC/us33/n829 , \AES_ENC/us33/n828 ,\AES_ENC/us33/n827 , \AES_ENC/us33/n826 , \AES_ENC/us33/n825 ,\AES_ENC/us33/n824 , \AES_ENC/us33/n823 , \AES_ENC/us33/n822 ,\AES_ENC/us33/n821 , \AES_ENC/us33/n820 , \AES_ENC/us33/n819 ,\AES_ENC/us33/n818 , \AES_ENC/us33/n817 , \AES_ENC/us33/n816 ,\AES_ENC/us33/n815 , \AES_ENC/us33/n814 , \AES_ENC/us33/n813 ,\AES_ENC/us33/n812 , \AES_ENC/us33/n811 , \AES_ENC/us33/n810 ,\AES_ENC/us33/n809 , \AES_ENC/us33/n808 , \AES_ENC/us33/n807 ,\AES_ENC/us33/n806 , \AES_ENC/us33/n805 , \AES_ENC/us33/n804 ,\AES_ENC/us33/n803 , \AES_ENC/us33/n802 , \AES_ENC/us33/n801 ,\AES_ENC/us33/n800 , \AES_ENC/us33/n799 , \AES_ENC/us33/n798 ,\AES_ENC/us33/n797 , \AES_ENC/us33/n796 , \AES_ENC/us33/n795 ,\AES_ENC/us33/n794 , \AES_ENC/us33/n793 , \AES_ENC/us33/n792 ,\AES_ENC/us33/n791 , \AES_ENC/us33/n790 , \AES_ENC/us33/n789 ,\AES_ENC/us33/n788 , \AES_ENC/us33/n787 , \AES_ENC/us33/n786 ,\AES_ENC/us33/n785 , \AES_ENC/us33/n784 , \AES_ENC/us33/n783 ,\AES_ENC/us33/n782 , \AES_ENC/us33/n781 , \AES_ENC/us33/n780 ,\AES_ENC/us33/n779 , \AES_ENC/us33/n778 , \AES_ENC/us33/n777 ,\AES_ENC/us33/n776 , \AES_ENC/us33/n775 , \AES_ENC/us33/n774 ,\AES_ENC/us33/n773 , \AES_ENC/us33/n772 , \AES_ENC/us33/n771 ,\AES_ENC/us33/n770 , \AES_ENC/us33/n769 , \AES_ENC/us33/n768 ,\AES_ENC/us33/n767 , \AES_ENC/us33/n766 , \AES_ENC/us33/n765 ,\AES_ENC/us33/n764 , \AES_ENC/us33/n763 , \AES_ENC/us33/n762 ,\AES_ENC/us33/n761 , \AES_ENC/us33/n760 , \AES_ENC/us33/n759 ,\AES_ENC/us33/n758 , \AES_ENC/us33/n757 , \AES_ENC/us33/n756 ,\AES_ENC/us33/n755 , \AES_ENC/us33/n754 , \AES_ENC/us33/n753 ,\AES_ENC/us33/n752 , \AES_ENC/us33/n751 , \AES_ENC/us33/n750 ,\AES_ENC/us33/n749 , \AES_ENC/us33/n748 , \AES_ENC/us33/n747 ,\AES_ENC/us33/n746 , \AES_ENC/us33/n745 , \AES_ENC/us33/n744 ,\AES_ENC/us33/n743 , \AES_ENC/us33/n742 , \AES_ENC/us33/n741 ,\AES_ENC/us33/n740 , \AES_ENC/us33/n739 , \AES_ENC/us33/n738 ,\AES_ENC/us33/n737 , \AES_ENC/us33/n736 , \AES_ENC/us33/n735 ,\AES_ENC/us33/n734 , \AES_ENC/us33/n733 , \AES_ENC/us33/n732 ,\AES_ENC/us33/n731 , \AES_ENC/us33/n730 , \AES_ENC/us33/n729 ,\AES_ENC/us33/n728 , \AES_ENC/us33/n727 , \AES_ENC/us33/n726 ,\AES_ENC/us33/n725 , \AES_ENC/us33/n724 , \AES_ENC/us33/n723 ,\AES_ENC/us33/n722 , \AES_ENC/us33/n721 , \AES_ENC/us33/n720 ,\AES_ENC/us33/n719 , \AES_ENC/us33/n718 , \AES_ENC/us33/n717 ,\AES_ENC/us33/n716 , \AES_ENC/us33/n715 , \AES_ENC/us33/n714 ,\AES_ENC/us33/n713 , \AES_ENC/us33/n712 , \AES_ENC/us33/n711 ,\AES_ENC/us33/n710 , \AES_ENC/us33/n709 , \AES_ENC/us33/n708 ,\AES_ENC/us33/n707 , \AES_ENC/us33/n706 , \AES_ENC/us33/n705 ,\AES_ENC/us33/n704 , \AES_ENC/us33/n703 , \AES_ENC/us33/n702 ,\AES_ENC/us33/n701 , \AES_ENC/us33/n700 , \AES_ENC/us33/n699 ,\AES_ENC/us33/n698 , \AES_ENC/us33/n697 , \AES_ENC/us33/n696 ,\AES_ENC/us33/n695 , \AES_ENC/us33/n694 , \AES_ENC/us33/n693 ,\AES_ENC/us33/n692 , \AES_ENC/us33/n691 , \AES_ENC/us33/n690 ,\AES_ENC/us33/n689 , \AES_ENC/us33/n688 , \AES_ENC/us33/n687 ,\AES_ENC/us33/n686 , \AES_ENC/us33/n685 , \AES_ENC/us33/n684 ,\AES_ENC/us33/n683 , \AES_ENC/us33/n682 , \AES_ENC/us33/n681 ,\AES_ENC/us33/n680 , \AES_ENC/us33/n679 , \AES_ENC/us33/n678 ,\AES_ENC/us33/n677 , \AES_ENC/us33/n676 , \AES_ENC/us33/n675 ,\AES_ENC/us33/n674 , \AES_ENC/us33/n673 , \AES_ENC/us33/n672 ,\AES_ENC/us33/n671 , \AES_ENC/us33/n670 , \AES_ENC/us33/n669 ,\AES_ENC/us33/n668 , \AES_ENC/us33/n667 , \AES_ENC/us33/n666 ,\AES_ENC/us33/n665 , \AES_ENC/us33/n664 , \AES_ENC/us33/n663 ,\AES_ENC/us33/n662 , \AES_ENC/us33/n661 , \AES_ENC/us33/n660 ,\AES_ENC/us33/n659 , \AES_ENC/us33/n658 , \AES_ENC/us33/n657 ,\AES_ENC/us33/n656 , \AES_ENC/us33/n655 , \AES_ENC/us33/n654 ,\AES_ENC/us33/n653 , \AES_ENC/us33/n652 , \AES_ENC/us33/n651 ,\AES_ENC/us33/n650 , \AES_ENC/us33/n649 , \AES_ENC/us33/n648 ,\AES_ENC/us33/n647 , \AES_ENC/us33/n646 , \AES_ENC/us33/n645 ,\AES_ENC/us33/n644 , \AES_ENC/us33/n643 , \AES_ENC/us33/n642 ,\AES_ENC/us33/n641 , \AES_ENC/us33/n640 , \AES_ENC/us33/n639 ,\AES_ENC/us33/n638 , \AES_ENC/us33/n637 , \AES_ENC/us33/n636 ,\AES_ENC/us33/n635 , \AES_ENC/us33/n634 , \AES_ENC/us33/n633 ,\AES_ENC/us33/n632 , \AES_ENC/us33/n631 , \AES_ENC/us33/n630 ,\AES_ENC/us33/n629 , \AES_ENC/us33/n628 , \AES_ENC/us33/n627 ,\AES_ENC/us33/n626 , \AES_ENC/us33/n625 , \AES_ENC/us33/n624 ,\AES_ENC/us33/n623 , \AES_ENC/us33/n622 , \AES_ENC/us33/n621 ,\AES_ENC/us33/n620 , \AES_ENC/us33/n619 , \AES_ENC/us33/n618 ,\AES_ENC/us33/n617 , \AES_ENC/us33/n616 , \AES_ENC/us33/n615 ,\AES_ENC/us33/n614 , \AES_ENC/us33/n613 , \AES_ENC/us33/n612 ,\AES_ENC/us33/n611 , \AES_ENC/us33/n610 , \AES_ENC/us33/n609 ,\AES_ENC/us33/n608 , \AES_ENC/us33/n607 , \AES_ENC/us33/n606 ,\AES_ENC/us33/n605 , \AES_ENC/us33/n604 , \AES_ENC/us33/n603 ,\AES_ENC/us33/n602 , \AES_ENC/us33/n601 , \AES_ENC/us33/n600 ,\AES_ENC/us33/n599 , \AES_ENC/us33/n598 , \AES_ENC/us33/n597 ,\AES_ENC/us33/n596 , \AES_ENC/us33/n595 , \AES_ENC/us33/n594 ,\AES_ENC/us33/n593 , \AES_ENC/us33/n592 , \AES_ENC/us33/n591 ,\AES_ENC/us33/n590 , \AES_ENC/us33/n589 , \AES_ENC/us33/n588 ,\AES_ENC/us33/n587 , \AES_ENC/us33/n586 , \AES_ENC/us33/n585 ,\AES_ENC/us33/n584 , \AES_ENC/us33/n583 , \AES_ENC/us33/n582 ,\AES_ENC/us33/n581 , \AES_ENC/us33/n580 , \AES_ENC/us33/n579 ,\AES_ENC/us33/n578 , \AES_ENC/us33/n577 , \AES_ENC/us33/n576 ,\AES_ENC/us33/n575 , \AES_ENC/us33/n574 , \AES_ENC/us33/n573 ,\AES_ENC/us33/n572 , \AES_ENC/us33/n571 , \AES_ENC/us33/n570 ,\AES_ENC/us33/n569 , \add_506/n647 , \add_506/n646 , \add_506/n645 ,\add_506/n644 , \add_506/n643 , \add_506/n642 , \add_506/n641 ,\add_506/n640 , \add_506/n639 , \add_506/n638 , \add_506/n637 ,\add_506/n636 , \add_506/n635 , \add_506/n634 , \add_506/n633 ,\add_506/n632 , \add_506/n631 , \add_506/n630 , \add_506/n629 ,\add_506/n628 , \add_506/n627 , \add_506/n626 , \add_506/n625 ,\add_506/n624 , \add_506/n623 , \add_506/n622 , \add_506/n621 ,\add_506/n620 , \add_506/n619 , \add_506/n618 , \add_506/n617 ,\add_506/n616 , \add_506/n615 , \add_506/n614 , \add_506/n613 ,\add_506/n612 , \add_506/n611 , \add_506/n610 , \add_506/n609 ,\add_506/n608 , \add_506/n607 , \add_506/n606 , \add_506/n605 ,\add_506/n604 , \add_506/n603 , \add_506/n602 , \add_506/n601 ,\add_506/n600 , \add_506/n599 , \add_506/n598 , \add_506/n597 ,\add_506/n596 , \add_506/n595 , \add_506/n594 , \add_506/n593 ,\add_506/n592 , \add_506/n591 , \add_506/n590 , \add_506/n589 ,\add_506/n588 , \add_506/n587 , \add_506/n586 , \add_506/n585 ,\add_506/n584 , \add_506/n583 , \add_506/n582 , \add_506/n581 ,\add_506/n580 , \add_506/n579 , \add_506/n578 , \add_506/n577 ,\add_506/n576 , \add_506/n575 , \add_506/n574 , \add_506/n573 ,\add_506/n572 , \add_506/n571 , \add_506/n570 , \add_506/n569 ,\add_506/n568 , \add_506/n567 , \add_506/n566 , \add_506/n565 ,\add_506/n564 , \add_506/n563 , \add_506/n562 , \add_506/n561 ,\add_506/n560 , \add_506/n559 , \add_506/n558 , \add_506/n557 ,\add_506/n556 , \add_506/n555 , \add_506/n554 , \add_506/n553 ,\add_506/n552 , \add_506/n551 , \add_506/n550 , \add_506/n549 ,\add_506/n548 , \add_506/n547 , \add_506/n546 , \add_506/n545 ,\add_506/n544 , \add_506/n543 , \add_506/n542 , \add_506/n541 ,\add_506/n540 , \add_506/n539 , \add_506/n538 , \add_506/n537 ,\add_506/n536 , \add_506/n535 , \add_506/n534 , \add_506/n533 ,\add_506/n532 , \add_506/n531 , \add_506/n530 , \add_506/n529 ,\add_506/n528 , \add_506/n527 , \add_506/n526 , \add_506/n525 ,\add_506/n524 , \add_506/n523 , \add_506/n522 , \add_506/n521 ,\add_506/n520 , \add_506/n519 , \add_506/n518 , \add_506/n517 ,\add_506/n516 , \add_506/n515 , \add_506/n514 , \add_506/n513 ,\add_506/n512 , \add_506/n511 , \add_506/n510 , \add_506/n509 ,\add_506/n508 , \add_506/n507 , \add_506/n506 , \add_506/n505 ,\add_506/n504 , \add_506/n503 , \add_506/n502 , \add_506/n501 ,\add_506/n500 , \add_506/n499 , \add_506/n498 , \add_506/n497 ,\add_506/n496 , \add_506/n495 , \add_506/n494 , \add_506/n493 ,\add_506/n492 , \add_506/n491 , \add_506/n490 , \add_506/n489 ,\add_506/n488 , \add_506/n487 , \add_506/n486 , \add_506/n485 ,\add_506/n484 , \add_506/n483 , \add_506/n482 , \add_506/n481 ,\add_506/n480 , \add_506/n479 , \add_506/n478 , \add_506/n477 ,\add_506/n476 , \add_506/n475 , \add_506/n474 , \add_506/n473 ,\add_506/n472 , \add_506/n471 , \add_506/n470 , \add_506/n469 ,\add_506/n468 , \add_506/n467 , \add_506/n466 , \add_506/n465 ,\add_506/n464 , \add_506/n463 , \add_506/n462 , \add_506/n461 ,\add_506/n460 , \add_506/n459 , \add_506/n458 , \add_506/n457 ,\add_506/n456 , \add_506/n455 , \add_506/n454 , \add_506/n453 ,\add_506/n452 , \add_506/n451 , \add_506/n450 , \add_506/n449 ,\add_506/n448 , \add_506/n447 , \add_506/n446 , \add_506/n445 ,\add_506/n444 , \add_506/n443 , \add_506/n442 , \add_506/n441 ,\add_506/n440 , \add_506/n439 , \add_506/n438 , \add_506/n437 ,\add_506/n436 , \add_506/n435 , \add_506/n434 , \add_506/n433 ,\add_506/n432 , \add_506/n431 , \add_506/n430 , \add_506/n429 ,\add_506/n428 , \add_506/n427 , \add_506/n426 , \add_506/n425 ,\add_506/n424 , \add_506/n423 , \add_506/n422 , \add_506/n421 ,\add_506/n420 , \add_506/n419 , \add_506/n418 , \add_506/n417 ,\add_506/n416 , \add_506/n415 , \add_506/n414 , \add_506/n413 ,\add_506/n412 , \add_506/n411 , \add_506/n410 , \add_506/n409 ,\add_506/n408 , \add_506/n407 , \add_506/n406 , \add_506/n405 ,\add_506/n404 , \add_506/n403 , \add_506/n402 , \add_506/n401 ,\add_506/n400 , \add_506/n399 , \add_506/n398 , \add_506/n397 ,\add_506/n396 , \add_506/n395 , \add_506/n394 , \add_506/n393 ,\add_506/n392 , \add_506/n391 , \add_506/n390 , \add_506/n389 ,\add_506/n388 , \add_506/n387 , \add_506/n386 , \add_506/n385 ,\add_506/n384 , \add_506/n383 , \add_506/n382 , \add_506/n381 ,\add_506/n380 , \add_506/n379 , \add_506/n378 , \add_506/n377 ,\add_506/n376 , \add_506/n375 , \add_506/n374 , \add_506/n373 ,\add_506/n372 , \add_506/n371 , \add_506/n370 , \add_506/n369 ,\add_506/n368 , \add_506/n367 , \add_506/n366 , \add_506/n365 ,\add_506/n364 , \add_506/n363 , \add_506/n362 , \add_506/n361 ,\add_506/n360 , \add_506/n359 , \add_506/n358 , \add_506/n357 ,\add_506/n356 , \add_506/n355 , \add_506/n354 , \add_506/n353 ,\add_506/n352 , \add_506/n351 , \add_506/n350 , \add_506/n349 ,\add_506/n348 , \add_506/n347 , \add_506/n346 , \add_506/n345 ,\add_506/n344 , \add_506/n343 , \add_506/n342 , \add_506/n341 ,\add_506/n340 , \add_506/n339 , \add_506/n338 , \add_506/n337 ,\add_506/n336 , \add_506/n335 , \add_506/n334 , \add_506/n333 ,\add_506/n332 , \add_506/n331 , \add_506/n330 , \add_506/n329 ,\add_506/n328 , \add_506/n327 , \add_506/n326 , \add_506/n325 ,\add_506/n324 , \add_506/n323 , \add_506/n322 , \add_506/n321 ,\add_506/n320 , \add_506/n319 , \add_506/n318 , \add_506/n317 ,\add_506/n316 , \add_506/n315 , \add_506/n314 , \add_506/n313 ,\add_506/n312 , \add_506/n311 , \add_506/n310 , \add_506/n309 ,\add_506/n308 , \add_506/n307 , \add_506/n306 , \add_506/n305 ,\add_506/n304 , \add_506/n303 , \add_506/n302 , \add_506/n301 ,\add_506/n300 , \add_506/n299 , \add_506/n298 , \add_506/n297 ,\add_506/n296 , \add_506/n295 , \add_506/n294 , \add_506/n293 ,\add_506/n292 , \add_506/n291 , \add_506/n290 , \add_506/n289 ,\add_506/n288 , \add_506/n287 , \add_506/n286 , \add_506/n285 ,\add_506/n284 , \add_506/n283 , \add_506/n282 , \add_506/n281 ,\add_506/n280 , \add_506/n279 , \add_506/n278 , \add_506/n277 ,\add_506/n276 , \add_506/n275 , \add_506/n274 , \add_506/n273 ,\add_506/n272 , \add_506/n271 , \add_506/n270 , \add_506/n269 ,\add_506/n268 , \add_506/n267 , \add_506/n266 , \add_506/n265 ,\add_506/n264 , \add_506/n263 , \add_506/n262 , \add_506/n261 ,\add_506/n260 , \add_506/n259 , \add_506/n258 , \add_506/n257 ,\add_506/n256 , \add_506/n255 , \add_506/n254 , \add_506/n253 ,\add_506/n252 , \add_506/n251 , \add_506/n250 , \add_506/n249 ,\add_506/n248 , \add_506/n247 , \add_506/n246 , \add_506/n245 ,\add_506/n244 , \add_506/n243 , \add_506/n242 , \add_506/n241 ,\add_506/n240 , \add_506/n239 , \add_506/n238 , \add_506/n237 ,\add_506/n236 , \add_506/n235 , \add_506/n234 , \add_506/n233 ,\add_506/n232 , \add_506/n231 , \add_506/n230 , \add_506/n229 ,\add_506/n228 , \add_506/n227 , \add_506/n226 , \add_506/n225 ,\add_506/n224 , \add_506/n223 , \add_506/n222 , \add_506/n221 ,\add_506/n220 , \add_506/n219 , \add_506/n218 , \add_506/n217 ,\add_506/n216 , \add_506/n215 , \add_506/n214 , \add_506/n213 ,\add_506/n212 , \add_506/n211 , \add_506/n210 , \add_506/n209 ,\add_506/n208 , \add_506/n207 , \add_506/n206 , \add_506/n205 ,\add_506/n204 , \add_506/n203 , \add_506/n202 , \add_506/n201 ,\add_506/n200 , \add_506/n199 , \add_506/n198 , \add_506/n197 ,\add_506/n196 , \add_506/n195 , \add_506/n194 , \add_506/n193 ,\add_506/n192 , \add_506/n191 , \add_506/n190 , \add_506/n189 ,\add_506/n188 , \add_506/n187 , \add_506/n186 , \add_506/n185 ,\add_506/n184 , \add_506/n183 , \add_506/n182 , \add_506/n181 ,\add_506/n180 , \add_506/n179 , \add_506/n178 , \add_506/n177 ,\add_506/n176 , \add_506/n175 , \add_506/n174 , \add_506/n173 ,\add_506/n172 , \add_506/n171 , \add_506/n170 , \add_506/n169 ,\add_506/n168 , \add_506/n167 , \add_506/n166 , \add_506/n165 ,\add_506/n164 , \add_506/n163 , \add_506/n162 , \add_506/n161 ,\add_506/n160 , \add_506/n159 , \add_506/n158 , \add_506/n157 ,\add_506/n156 , \add_506/n155 , \add_506/n154 , \add_506/n153 ,\add_506/n152 , \add_506/n151 , \add_506/n150 , \add_506/n149 ,\add_506/n148 , \add_506/n147 , \add_506/n146 , \add_506/n145 ,\add_506/n144 , \add_506/n143 , \add_506/n142 , \add_506/n141 ,\add_506/n140 , \add_506/n139 , \add_506/n138 , \add_506/n137 ,\add_506/n136 , \add_506/n135 , \add_506/n134 , \add_506/n133 ,\add_506/n132 , \add_506/n131 , \add_506/n130 , \add_506/n129 ,\add_506/n128 , \add_506/n127 , \add_506/n126 , \add_506/n125 ,\add_506/n124 , \add_506/n123 , \add_506/n122 , \add_506/n121 ,\add_506/n120 , \add_506/n119 , \add_506/n118 , \add_506/n117 ,\add_506/n116 , \add_506/n115 , \add_506/n114 , \add_506/n113 ,\add_506/n112 , \add_506/n111 , \add_506/n110 , \add_506/n109 ,\add_506/n108 , \add_506/n107 , \add_506/n106 , \add_506/n105 ,\add_506/n104 , \add_506/n103 , \add_506/n102 , \add_506/n101 ,\add_506/n100 , \add_506/n99 , \add_506/n98 , \add_506/n97 ,\add_506/n96 , \add_506/n95 , \add_506/n94 , \add_506/n93 ,\add_506/n92 , \add_506/n91 , \add_506/n90 , \add_506/n89 ,\add_506/n88 , \add_506/n87 , \add_506/n86 , \add_506/n85 ,\add_506/n84 , \add_506/n83 , \add_506/n82 , \add_506/n81 ,\add_506/n80 , \add_506/n79 , \add_506/n78 , \add_506/n77 ,\add_506/n76 , \add_506/n75 , \add_506/n74 , \add_506/n73 ,\add_506/n72 , \add_506/n71 , \add_506/n70 , \add_506/n69 ,\add_506/n68 , \add_506/n67 , \add_506/n66 , \add_506/n65 ,\add_506/n64 , \add_506/n63 , \add_506/n62 , \add_506/n61 ,\add_506/n60 , \add_506/n59 , \add_506/n58 , \add_506/n57 ,\add_506/n56 , \add_506/n55 , \add_506/n54 , \add_506/n53 ,\add_506/n52 , \add_506/n51 , \add_506/n50 , \add_506/n49 ,\add_506/n48 , \add_506/n47 , \add_506/n46 , \add_506/n45 ,\add_506/n44 , \add_506/n43 , \add_506/n42 , \add_506/n41 ,\add_506/n40 , \add_506/n39 , \add_506/n38 , \add_506/n37 ,\add_506/n36 , \add_506/n35 , \add_506/n34 , \add_506/n33 ,\add_506/n32 , \add_506/n31 , \add_506/n30 , \add_506/n29 ,\add_506/n28 , \add_506/n27 , \add_506/n26 , \add_506/n25 ,\add_506/n24 , \add_506/n23 , \add_506/n22 , \add_506/n21 ,\add_506/n20 , \add_506/n19 , \add_506/n18 , \add_506/n17 ,\add_506/n16 , \add_506/n15 , \add_506/n14 , \add_506/n13 ,\add_506/n12 , \add_506/n11 , \add_506/n10 , \add_506/n9 ,\add_506/n8 , \add_506/n7 , \add_506/n6 , \add_506/n4 , \add_506/n3 ,\add_506/n2 , \add_506/n1 , \add_1_root_add_519_2/n224 ,\add_1_root_add_519_2/n223 , \add_1_root_add_519_2/n222 ,\add_1_root_add_519_2/n221 , \add_1_root_add_519_2/n220 ,\add_1_root_add_519_2/n219 , \add_1_root_add_519_2/n218 ,\add_1_root_add_519_2/n217 , \add_1_root_add_519_2/n216 ,\add_1_root_add_519_2/n215 , \add_1_root_add_519_2/n214 ,\add_1_root_add_519_2/n213 , \add_1_root_add_519_2/n212 ,\add_1_root_add_519_2/n211 , \add_1_root_add_519_2/n210 ,\add_1_root_add_519_2/n209 , \add_1_root_add_519_2/n208 ,\add_1_root_add_519_2/n207 , \add_1_root_add_519_2/n206 ,\add_1_root_add_519_2/n205 , \add_1_root_add_519_2/n204 ,\add_1_root_add_519_2/n203 , \add_1_root_add_519_2/n202 ,\add_1_root_add_519_2/n201 , \add_1_root_add_519_2/n200 ,\add_1_root_add_519_2/n199 , \add_1_root_add_519_2/n198 ,\add_1_root_add_519_2/n197 , \add_1_root_add_519_2/n196 ,\add_1_root_add_519_2/n195 , \add_1_root_add_519_2/n194 ,\add_1_root_add_519_2/n193 , \add_1_root_add_519_2/n192 ,\add_1_root_add_519_2/n191 , \add_1_root_add_519_2/n190 ,\add_1_root_add_519_2/n189 , \add_1_root_add_519_2/n188 ,\add_1_root_add_519_2/n187 , \add_1_root_add_519_2/n186 ,\add_1_root_add_519_2/n185 , \add_1_root_add_519_2/n184 ,\add_1_root_add_519_2/n183 , \add_1_root_add_519_2/n182 ,\add_1_root_add_519_2/n181 , \add_1_root_add_519_2/n180 ,\add_1_root_add_519_2/n179 , \add_1_root_add_519_2/n178 ,\add_1_root_add_519_2/n177 , \add_1_root_add_519_2/n176 ,\add_1_root_add_519_2/n175 , \add_1_root_add_519_2/n174 ,\add_1_root_add_519_2/n173 , \add_1_root_add_519_2/n172 ,\add_1_root_add_519_2/n171 , \add_1_root_add_519_2/n170 ,\add_1_root_add_519_2/n169 , \add_1_root_add_519_2/n168 ,\add_1_root_add_519_2/n167 , \add_1_root_add_519_2/n166 ,\add_1_root_add_519_2/n165 , \add_1_root_add_519_2/n164 ,\add_1_root_add_519_2/n163 , \add_1_root_add_519_2/n162 ,\add_1_root_add_519_2/n161 , \add_1_root_add_519_2/n160 ,\add_1_root_add_519_2/n159 , \add_1_root_add_519_2/n158 ,\add_1_root_add_519_2/n157 , \add_1_root_add_519_2/n156 ,\add_1_root_add_519_2/n155 , \add_1_root_add_519_2/n154 ,\add_1_root_add_519_2/n153 , \add_1_root_add_519_2/n152 ,\add_1_root_add_519_2/n151 , \add_1_root_add_519_2/n150 ,\add_1_root_add_519_2/n149 , \add_1_root_add_519_2/n148 ,\add_1_root_add_519_2/n147 , \add_1_root_add_519_2/n146 ,\add_1_root_add_519_2/n145 , \add_1_root_add_519_2/n144 ,\add_1_root_add_519_2/n143 , \add_1_root_add_519_2/n142 ,\add_1_root_add_519_2/n141 , \add_1_root_add_519_2/n140 ,\add_1_root_add_519_2/n139 , \add_1_root_add_519_2/n138 ,\add_1_root_add_519_2/n137 , \add_1_root_add_519_2/n136 ,\add_1_root_add_519_2/n135 , \add_1_root_add_519_2/n134 ,\add_1_root_add_519_2/n133 , \add_1_root_add_519_2/n132 ,\add_1_root_add_519_2/n131 , \add_1_root_add_519_2/n130 ,\add_1_root_add_519_2/n129 , \add_1_root_add_519_2/n128 ,\add_1_root_add_519_2/n127 , \add_1_root_add_519_2/n126 ,\add_1_root_add_519_2/n125 , \add_1_root_add_519_2/n124 ,\add_1_root_add_519_2/n123 , \add_1_root_add_519_2/n122 ,\add_1_root_add_519_2/n121 , \add_1_root_add_519_2/n120 ,\add_1_root_add_519_2/n119 , \add_1_root_add_519_2/n118 ,\add_1_root_add_519_2/n117 , \add_1_root_add_519_2/n116 ,\add_1_root_add_519_2/n115 , \add_1_root_add_519_2/n114 ,\add_1_root_add_519_2/n113 , \add_1_root_add_519_2/n112 ,\add_1_root_add_519_2/n111 , \add_1_root_add_519_2/n110 ,\add_1_root_add_519_2/n109 , \add_1_root_add_519_2/n108 ,\add_1_root_add_519_2/n107 , \add_1_root_add_519_2/n106 ,\add_1_root_add_519_2/n105 , \add_1_root_add_519_2/n104 ,\add_1_root_add_519_2/n103 , \add_1_root_add_519_2/n102 ,\add_1_root_add_519_2/n101 , \add_1_root_add_519_2/n100 ,\add_1_root_add_519_2/n99 , \add_1_root_add_519_2/n98 ,\add_1_root_add_519_2/n97 , \add_1_root_add_519_2/n96 ,\add_1_root_add_519_2/n95 , \add_1_root_add_519_2/n94 ,\add_1_root_add_519_2/n93 , \add_1_root_add_519_2/n92 ,\add_1_root_add_519_2/n91 , \add_1_root_add_519_2/n90 ,\add_1_root_add_519_2/n89 , \add_1_root_add_519_2/n88 ,\add_1_root_add_519_2/n87 , \add_1_root_add_519_2/n86 ,\add_1_root_add_519_2/n85 , \add_1_root_add_519_2/n84 ,\add_1_root_add_519_2/n83 , \add_1_root_add_519_2/n82 ,\add_1_root_add_519_2/n81 , \add_1_root_add_519_2/n80 ,\add_1_root_add_519_2/n79 , \add_1_root_add_519_2/n78 ,\add_1_root_add_519_2/n77 , \add_1_root_add_519_2/n76 ,\add_1_root_add_519_2/n75 , \add_1_root_add_519_2/n74 ,\add_1_root_add_519_2/n73 , \add_1_root_add_519_2/n72 ,\add_1_root_add_519_2/n71 , \add_1_root_add_519_2/n70 ,\add_1_root_add_519_2/n69 , \add_1_root_add_519_2/n68 ,\add_1_root_add_519_2/n67 , \add_1_root_add_519_2/n66 ,\add_1_root_add_519_2/n65 , \add_1_root_add_519_2/n64 ,\add_1_root_add_519_2/n63 , \add_1_root_add_519_2/n62 ,\add_1_root_add_519_2/n61 , \add_1_root_add_519_2/n60 ,\add_1_root_add_519_2/n59 , \add_1_root_add_519_2/n58 ,\add_1_root_add_519_2/n57 , \add_1_root_add_519_2/n56 ,\add_1_root_add_519_2/n55 , \add_1_root_add_519_2/n54 ,\add_1_root_add_519_2/n53 , \add_1_root_add_519_2/n52 ,\add_1_root_add_519_2/n51 , \add_1_root_add_519_2/n50 ,\add_1_root_add_519_2/n49 , \add_1_root_add_519_2/n48 ,\add_1_root_add_519_2/n47 , \add_1_root_add_519_2/n46 ,\add_1_root_add_519_2/n45 , \add_1_root_add_519_2/n44 ,\add_1_root_add_519_2/n43 , \add_1_root_add_519_2/n42 ,\add_1_root_add_519_2/n41 , \add_1_root_add_519_2/n40 ,\add_1_root_add_519_2/n39 , \add_1_root_add_519_2/n38 ,\add_1_root_add_519_2/n37 , \add_1_root_add_519_2/n36 ,\add_1_root_add_519_2/n35 , \add_1_root_add_519_2/n34 ,\add_1_root_add_519_2/n33 , \add_1_root_add_519_2/n32 ,\add_1_root_add_519_2/n31 , \add_1_root_add_519_2/n30 ,\add_1_root_add_519_2/n29 , \add_1_root_add_519_2/n28 ,\add_1_root_add_519_2/n27 , \add_1_root_add_519_2/n26 ,\add_1_root_add_519_2/n25 , \add_1_root_add_519_2/n24 ,\add_1_root_add_519_2/n23 , \add_1_root_add_519_2/n22 ,\add_1_root_add_519_2/n21 , \add_1_root_add_519_2/n20 ,\add_1_root_add_519_2/n19 , \add_1_root_add_519_2/n18 ,\add_1_root_add_519_2/n17 , \add_1_root_add_519_2/n16 ,\add_1_root_add_519_2/n15 , \add_1_root_add_519_2/n14 ,\add_1_root_add_519_2/n13 , \add_1_root_add_519_2/n12 ,\add_1_root_add_519_2/n11 , \add_1_root_add_519_2/n10 ,\add_1_root_add_519_2/n9 , \add_1_root_add_519_2/n8 ,\add_1_root_add_519_2/n7 , \add_1_root_add_519_2/n6 ,\add_1_root_add_519_2/n5 , \add_1_root_add_519_2/n4 ,\add_1_root_add_519_2/n3 , \add_1_root_add_519_2/n2 ,\add_1_root_add_519_2/n1 , \add_1_root_add_513_2/n224 ,\add_1_root_add_513_2/n223 , \add_1_root_add_513_2/n222 ,\add_1_root_add_513_2/n221 , \add_1_root_add_513_2/n220 ,\add_1_root_add_513_2/n219 , \add_1_root_add_513_2/n218 ,\add_1_root_add_513_2/n217 , \add_1_root_add_513_2/n216 ,\add_1_root_add_513_2/n215 , \add_1_root_add_513_2/n214 ,\add_1_root_add_513_2/n213 , \add_1_root_add_513_2/n212 ,\add_1_root_add_513_2/n211 , \add_1_root_add_513_2/n210 ,\add_1_root_add_513_2/n209 , \add_1_root_add_513_2/n208 ,\add_1_root_add_513_2/n207 , \add_1_root_add_513_2/n206 ,\add_1_root_add_513_2/n205 , \add_1_root_add_513_2/n204 ,\add_1_root_add_513_2/n203 , \add_1_root_add_513_2/n202 ,\add_1_root_add_513_2/n201 , \add_1_root_add_513_2/n200 ,\add_1_root_add_513_2/n199 , \add_1_root_add_513_2/n198 ,\add_1_root_add_513_2/n197 , \add_1_root_add_513_2/n196 ,\add_1_root_add_513_2/n195 , \add_1_root_add_513_2/n194 ,\add_1_root_add_513_2/n193 , \add_1_root_add_513_2/n192 ,\add_1_root_add_513_2/n191 , \add_1_root_add_513_2/n190 ,\add_1_root_add_513_2/n189 , \add_1_root_add_513_2/n188 ,\add_1_root_add_513_2/n187 , \add_1_root_add_513_2/n186 ,\add_1_root_add_513_2/n185 , \add_1_root_add_513_2/n184 ,\add_1_root_add_513_2/n183 , \add_1_root_add_513_2/n182 ,\add_1_root_add_513_2/n181 , \add_1_root_add_513_2/n180 ,\add_1_root_add_513_2/n179 , \add_1_root_add_513_2/n178 ,\add_1_root_add_513_2/n177 , \add_1_root_add_513_2/n176 ,\add_1_root_add_513_2/n175 , \add_1_root_add_513_2/n174 ,\add_1_root_add_513_2/n173 , \add_1_root_add_513_2/n172 ,\add_1_root_add_513_2/n171 , \add_1_root_add_513_2/n170 ,\add_1_root_add_513_2/n169 , \add_1_root_add_513_2/n168 ,\add_1_root_add_513_2/n167 , \add_1_root_add_513_2/n166 ,\add_1_root_add_513_2/n165 , \add_1_root_add_513_2/n164 ,\add_1_root_add_513_2/n163 , \add_1_root_add_513_2/n162 ,\add_1_root_add_513_2/n161 , \add_1_root_add_513_2/n160 ,\add_1_root_add_513_2/n159 , \add_1_root_add_513_2/n158 ,\add_1_root_add_513_2/n157 , \add_1_root_add_513_2/n156 ,\add_1_root_add_513_2/n155 , \add_1_root_add_513_2/n154 ,\add_1_root_add_513_2/n153 , \add_1_root_add_513_2/n152 ,\add_1_root_add_513_2/n151 , \add_1_root_add_513_2/n150 ,\add_1_root_add_513_2/n149 , \add_1_root_add_513_2/n148 ,\add_1_root_add_513_2/n147 , \add_1_root_add_513_2/n146 ,\add_1_root_add_513_2/n145 , \add_1_root_add_513_2/n144 ,\add_1_root_add_513_2/n143 , \add_1_root_add_513_2/n142 ,\add_1_root_add_513_2/n141 , \add_1_root_add_513_2/n140 ,\add_1_root_add_513_2/n139 , \add_1_root_add_513_2/n138 ,\add_1_root_add_513_2/n137 , \add_1_root_add_513_2/n136 ,\add_1_root_add_513_2/n135 , \add_1_root_add_513_2/n134 ,\add_1_root_add_513_2/n133 , \add_1_root_add_513_2/n132 ,\add_1_root_add_513_2/n131 , \add_1_root_add_513_2/n130 ,\add_1_root_add_513_2/n129 , \add_1_root_add_513_2/n128 ,\add_1_root_add_513_2/n127 , \add_1_root_add_513_2/n126 ,\add_1_root_add_513_2/n125 , \add_1_root_add_513_2/n124 ,\add_1_root_add_513_2/n123 , \add_1_root_add_513_2/n122 ,\add_1_root_add_513_2/n121 , \add_1_root_add_513_2/n120 ,\add_1_root_add_513_2/n119 , \add_1_root_add_513_2/n118 ,\add_1_root_add_513_2/n117 , \add_1_root_add_513_2/n116 ,\add_1_root_add_513_2/n115 , \add_1_root_add_513_2/n114 ,\add_1_root_add_513_2/n113 , \add_1_root_add_513_2/n112 ,\add_1_root_add_513_2/n111 , \add_1_root_add_513_2/n110 ,\add_1_root_add_513_2/n109 , \add_1_root_add_513_2/n108 ,\add_1_root_add_513_2/n107 , \add_1_root_add_513_2/n106 ,\add_1_root_add_513_2/n105 , \add_1_root_add_513_2/n104 ,\add_1_root_add_513_2/n103 , \add_1_root_add_513_2/n102 ,\add_1_root_add_513_2/n101 , \add_1_root_add_513_2/n100 ,\add_1_root_add_513_2/n99 , \add_1_root_add_513_2/n98 ,\add_1_root_add_513_2/n97 , \add_1_root_add_513_2/n96 ,\add_1_root_add_513_2/n95 , \add_1_root_add_513_2/n94 ,\add_1_root_add_513_2/n93 , \add_1_root_add_513_2/n92 ,\add_1_root_add_513_2/n91 , \add_1_root_add_513_2/n90 ,\add_1_root_add_513_2/n89 , \add_1_root_add_513_2/n88 ,\add_1_root_add_513_2/n87 , \add_1_root_add_513_2/n86 ,\add_1_root_add_513_2/n85 , \add_1_root_add_513_2/n84 ,\add_1_root_add_513_2/n83 , \add_1_root_add_513_2/n82 ,\add_1_root_add_513_2/n81 , \add_1_root_add_513_2/n80 ,\add_1_root_add_513_2/n79 , \add_1_root_add_513_2/n78 ,\add_1_root_add_513_2/n77 , \add_1_root_add_513_2/n76 ,\add_1_root_add_513_2/n75 , \add_1_root_add_513_2/n74 ,\add_1_root_add_513_2/n73 , \add_1_root_add_513_2/n72 ,\add_1_root_add_513_2/n71 , \add_1_root_add_513_2/n70 ,\add_1_root_add_513_2/n69 , \add_1_root_add_513_2/n68 ,\add_1_root_add_513_2/n67 , \add_1_root_add_513_2/n66 ,\add_1_root_add_513_2/n65 , \add_1_root_add_513_2/n64 ,\add_1_root_add_513_2/n63 , \add_1_root_add_513_2/n62 ,\add_1_root_add_513_2/n61 , \add_1_root_add_513_2/n60 ,\add_1_root_add_513_2/n59 , \add_1_root_add_513_2/n58 ,\add_1_root_add_513_2/n57 , \add_1_root_add_513_2/n56 ,\add_1_root_add_513_2/n55 , \add_1_root_add_513_2/n54 ,\add_1_root_add_513_2/n53 , \add_1_root_add_513_2/n52 ,\add_1_root_add_513_2/n51 , \add_1_root_add_513_2/n50 ,\add_1_root_add_513_2/n49 , \add_1_root_add_513_2/n48 ,\add_1_root_add_513_2/n47 , \add_1_root_add_513_2/n46 ,\add_1_root_add_513_2/n45 , \add_1_root_add_513_2/n44 ,\add_1_root_add_513_2/n43 , \add_1_root_add_513_2/n42 ,\add_1_root_add_513_2/n41 , \add_1_root_add_513_2/n40 ,\add_1_root_add_513_2/n39 , \add_1_root_add_513_2/n38 ,\add_1_root_add_513_2/n37 , \add_1_root_add_513_2/n36 ,\add_1_root_add_513_2/n35 , \add_1_root_add_513_2/n34 ,\add_1_root_add_513_2/n33 , \add_1_root_add_513_2/n32 ,\add_1_root_add_513_2/n31 , \add_1_root_add_513_2/n30 ,\add_1_root_add_513_2/n29 , \add_1_root_add_513_2/n28 ,\add_1_root_add_513_2/n27 , \add_1_root_add_513_2/n26 ,\add_1_root_add_513_2/n25 , \add_1_root_add_513_2/n24 ,\add_1_root_add_513_2/n23 , \add_1_root_add_513_2/n22 ,\add_1_root_add_513_2/n21 , \add_1_root_add_513_2/n20 ,\add_1_root_add_513_2/n19 , \add_1_root_add_513_2/n18 ,\add_1_root_add_513_2/n17 , \add_1_root_add_513_2/n16 ,\add_1_root_add_513_2/n15 , \add_1_root_add_513_2/n14 ,\add_1_root_add_513_2/n13 , \add_1_root_add_513_2/n12 ,\add_1_root_add_513_2/n11 , \add_1_root_add_513_2/n10 ,\add_1_root_add_513_2/n9 , \add_1_root_add_513_2/n8 ,\add_1_root_add_513_2/n7 , \add_1_root_add_513_2/n6 ,\add_1_root_add_513_2/n5 , \add_1_root_add_513_2/n4 ,\add_1_root_add_513_2/n3 , \add_1_root_add_513_2/n2 ,\add_1_root_add_513_2/n1 ;
wire   [9:0] state;
wire   [127:0] aes_text_in;
wire   [127:0] aes_text_out;
wire   [63:0] aad_byte_cnt;
wire   [63:0] enc_byte_cnt;
wire   [127:0] z_out;
wire   [127:0] v_in;
wire   [127:0] z_in;
wire   [127:0] b_in;
wire   [127:0] v_out;
wire   [7:0] \AES_ENC/sa00_next ;
wire   [7:0] \AES_ENC/sa00 ;
wire   [7:0] \AES_ENC/sa10_next ;
wire   [7:0] \AES_ENC/sa10 ;
wire   [7:0] \AES_ENC/sa20_next ;
wire   [7:0] \AES_ENC/sa20 ;
wire   [7:0] \AES_ENC/sa30_next ;
wire   [7:0] \AES_ENC/sa30 ;
wire   [7:0] \AES_ENC/sa01_next ;
wire   [7:0] \AES_ENC/sa01 ;
wire   [7:0] \AES_ENC/sa11_next ;
wire   [7:0] \AES_ENC/sa11 ;
wire   [7:0] \AES_ENC/sa21_next ;
wire   [7:0] \AES_ENC/sa21 ;
wire   [7:0] \AES_ENC/sa31_next ;
wire   [7:0] \AES_ENC/sa31 ;
wire   [7:0] \AES_ENC/sa02_next ;
wire   [7:0] \AES_ENC/sa02 ;
wire   [7:0] \AES_ENC/sa12_next ;
wire   [7:0] \AES_ENC/sa12 ;
wire   [7:0] \AES_ENC/sa22_next ;
wire   [7:0] \AES_ENC/sa22 ;
wire   [7:0] \AES_ENC/sa32_next ;
wire   [7:0] \AES_ENC/sa32 ;
wire   [7:0] \AES_ENC/sa03_next ;
wire   [7:0] \AES_ENC/sa03 ;
wire   [7:0] \AES_ENC/sa13_next ;
wire   [7:0] \AES_ENC/sa13 ;
wire   [7:0] \AES_ENC/sa23_next ;
wire   [7:0] \AES_ENC/sa23 ;
wire   [7:0] \AES_ENC/sa33_next ;
wire   [7:0] \AES_ENC/sa33 ;
wire   [31:24] \AES_ENC/u0/rcon ;
DFFR_X1 H_reg_127_ ( .D(n6027), .CK(clk), .RN(n17825), .Q(n17292), .QN() );
DFFR_X1 H_reg_126_ ( .D(n6028), .CK(clk), .RN(n17825), .Q(n17293), .QN() );
DFFR_X1 H_reg_125_ ( .D(n6029), .CK(clk), .RN(n17825), .Q(n17294), .QN() );
DFFR_X1 H_reg_124_ ( .D(n6030), .CK(clk), .RN(n17825), .Q(n17295), .QN() );
DFFR_X1 H_reg_123_ ( .D(n6031), .CK(clk), .RN(n17825), .Q(n17296), .QN() );
DFFR_X1 H_reg_122_ ( .D(n6032), .CK(clk), .RN(n17825), .Q(n17297), .QN() );
DFFR_X1 H_reg_121_ ( .D(n6033), .CK(clk), .RN(n17825), .Q(n17298), .QN() );
DFFR_X1 H_reg_120_ ( .D(n6034), .CK(clk), .RN(n17825), .Q(n17299), .QN() );
DFFR_X1 H_reg_119_ ( .D(n6035), .CK(clk), .RN(n17825), .Q(n17300), .QN() );
DFFR_X1 H_reg_118_ ( .D(n6036), .CK(clk), .RN(n17825), .Q(n17301), .QN() );
DFFR_X1 H_reg_117_ ( .D(n6037), .CK(clk), .RN(n17825), .Q(n17302), .QN() );
DFFR_X1 H_reg_116_ ( .D(n6038), .CK(clk), .RN(n17826), .Q(n17303), .QN() );
DFFR_X1 H_reg_115_ ( .D(n6039), .CK(clk), .RN(n17826), .Q(n17304), .QN() );
DFFR_X1 H_reg_114_ ( .D(n6040), .CK(clk), .RN(n17826), .Q(n17305), .QN() );
DFFR_X1 H_reg_113_ ( .D(n6041), .CK(clk), .RN(n17826), .Q(n17306), .QN() );
DFFR_X1 H_reg_112_ ( .D(n6042), .CK(clk), .RN(n17826), .Q(n17307), .QN() );
DFFR_X1 H_reg_111_ ( .D(n6043), .CK(clk), .RN(n17826), .Q(n17308), .QN() );
DFFR_X1 H_reg_110_ ( .D(n6044), .CK(clk), .RN(n17826), .Q(n17309), .QN() );
DFFR_X1 H_reg_109_ ( .D(n6045), .CK(clk), .RN(n17826), .Q(n17310), .QN() );
DFFR_X1 H_reg_108_ ( .D(n6046), .CK(clk), .RN(n17826), .Q(n17311), .QN() );
DFFR_X1 H_reg_107_ ( .D(n6047), .CK(clk), .RN(n17826), .Q(n17312), .QN() );
DFFR_X1 H_reg_106_ ( .D(n6048), .CK(clk), .RN(n17826), .Q(n17313), .QN() );
DFFR_X1 H_reg_105_ ( .D(n6049), .CK(clk), .RN(n17826), .Q(n17314), .QN() );
DFFR_X1 H_reg_104_ ( .D(n6050), .CK(clk), .RN(n17827), .Q(n17315), .QN() );
DFFR_X1 H_reg_103_ ( .D(n6051), .CK(clk), .RN(n17827), .Q(n17316), .QN() );
DFFR_X1 H_reg_102_ ( .D(n6052), .CK(clk), .RN(n17827), .Q(n17317), .QN() );
DFFR_X1 H_reg_101_ ( .D(n6053), .CK(clk), .RN(n17827), .Q(n17318), .QN() );
DFFR_X1 H_reg_100_ ( .D(n6054), .CK(clk), .RN(n17827), .Q(n17319), .QN() );
DFFR_X1 H_reg_99_ ( .D(n6055), .CK(clk), .RN(n17827), .Q(n17320), .QN() );
DFFR_X1 H_reg_98_ ( .D(n6056), .CK(clk), .RN(n17827), .Q(n17321), .QN() );
DFFR_X1 H_reg_97_ ( .D(n6057), .CK(clk), .RN(n17827), .Q(n17322), .QN() );
DFFR_X1 H_reg_96_ ( .D(n6058), .CK(clk), .RN(n17827), .Q(n17323), .QN() );
DFFR_X1 H_reg_95_ ( .D(n6059), .CK(clk), .RN(n17827), .Q(n17324), .QN() );
DFFR_X1 H_reg_94_ ( .D(n6060), .CK(clk), .RN(n17827), .Q(n17325), .QN() );
DFFR_X1 H_reg_93_ ( .D(n6061), .CK(clk), .RN(n17827), .Q(n17326), .QN() );
DFFR_X1 H_reg_92_ ( .D(n6062), .CK(clk), .RN(n17828), .Q(n17327), .QN() );
DFFR_X1 H_reg_91_ ( .D(n6063), .CK(clk), .RN(n17828), .Q(n17328), .QN() );
DFFR_X1 H_reg_90_ ( .D(n6064), .CK(clk), .RN(n17828), .Q(n17329), .QN() );
DFFR_X1 H_reg_89_ ( .D(n6065), .CK(clk), .RN(n17828), .Q(n17330), .QN() );
DFFR_X1 H_reg_88_ ( .D(n6066), .CK(clk), .RN(n17828), .Q(n17331), .QN() );
DFFR_X1 H_reg_87_ ( .D(n6067), .CK(clk), .RN(n17828), .Q(n17332), .QN() );
DFFR_X1 H_reg_86_ ( .D(n6068), .CK(clk), .RN(n17828), .Q(n17333), .QN() );
DFFR_X1 H_reg_85_ ( .D(n6069), .CK(clk), .RN(n17828), .Q(n17334), .QN() );
DFFR_X1 H_reg_84_ ( .D(n6070), .CK(clk), .RN(n17828), .Q(n17335), .QN() );
DFFR_X1 H_reg_83_ ( .D(n6071), .CK(clk), .RN(n17828), .Q(n17336), .QN() );
DFFR_X1 H_reg_82_ ( .D(n6072), .CK(clk), .RN(n17828), .Q(n17337), .QN() );
DFFR_X1 H_reg_81_ ( .D(n6073), .CK(clk), .RN(n17828), .Q(n17338), .QN() );
DFFR_X1 H_reg_80_ ( .D(n6074), .CK(clk), .RN(n17829), .Q(n17339), .QN() );
DFFR_X1 H_reg_79_ ( .D(n6075), .CK(clk), .RN(n17829), .Q(n17340), .QN() );
DFFR_X1 H_reg_78_ ( .D(n6076), .CK(clk), .RN(n17829), .Q(n17341), .QN() );
DFFR_X1 H_reg_77_ ( .D(n6077), .CK(clk), .RN(n17829), .Q(n17342), .QN() );
DFFR_X1 H_reg_76_ ( .D(n6078), .CK(clk), .RN(n17829), .Q(n17343), .QN() );
DFFR_X1 H_reg_75_ ( .D(n6079), .CK(clk), .RN(n17829), .Q(n17344), .QN() );
DFFR_X1 H_reg_74_ ( .D(n6080), .CK(clk), .RN(n17829), .Q(n17345), .QN() );
DFFR_X1 H_reg_73_ ( .D(n6081), .CK(clk), .RN(n17829), .Q(n17346), .QN() );
DFFR_X1 H_reg_72_ ( .D(n6082), .CK(clk), .RN(n17829), .Q(n17347), .QN() );
DFFR_X1 H_reg_71_ ( .D(n6083), .CK(clk), .RN(n17829), .Q(n17348), .QN() );
DFFR_X1 H_reg_70_ ( .D(n6084), .CK(clk), .RN(n17829), .Q(n17349), .QN() );
DFFR_X1 H_reg_69_ ( .D(n6085), .CK(clk), .RN(n17829), .Q(n17350), .QN() );
DFFR_X1 H_reg_68_ ( .D(n6086), .CK(clk), .RN(n17830), .Q(n17351), .QN() );
DFFR_X1 H_reg_67_ ( .D(n6087), .CK(clk), .RN(n17830), .Q(n17352), .QN() );
DFFR_X1 H_reg_66_ ( .D(n6088), .CK(clk), .RN(n17830), .Q(n17353), .QN() );
DFFR_X1 H_reg_65_ ( .D(n6089), .CK(clk), .RN(n17830), .Q(n17354), .QN() );
DFFR_X1 H_reg_64_ ( .D(n6090), .CK(clk), .RN(n17830), .Q(n17355), .QN() );
DFFR_X1 H_reg_63_ ( .D(n6091), .CK(clk), .RN(n17830), .Q(n17356), .QN() );
DFFR_X1 H_reg_62_ ( .D(n6092), .CK(clk), .RN(n17830), .Q(n17357), .QN() );
DFFR_X1 H_reg_61_ ( .D(n6093), .CK(clk), .RN(n17830), .Q(n17358), .QN() );
DFFR_X1 H_reg_60_ ( .D(n6094), .CK(clk), .RN(n17830), .Q(n17359), .QN() );
DFFR_X1 H_reg_59_ ( .D(n6095), .CK(clk), .RN(n17830), .Q(n17360), .QN() );
DFFR_X1 H_reg_58_ ( .D(n6096), .CK(clk), .RN(n17830), .Q(n17361), .QN() );
DFFR_X1 H_reg_57_ ( .D(n6097), .CK(clk), .RN(n17830), .Q(n17362), .QN() );
DFFR_X1 H_reg_56_ ( .D(n6098), .CK(clk), .RN(n17831), .Q(n17363), .QN() );
DFFR_X1 H_reg_55_ ( .D(n6099), .CK(clk), .RN(n17831), .Q(n17364), .QN() );
DFFR_X1 H_reg_54_ ( .D(n6100), .CK(clk), .RN(n17831), .Q(n17365), .QN() );
DFFR_X1 H_reg_53_ ( .D(n6101), .CK(clk), .RN(n17831), .Q(n17366), .QN() );
DFFR_X1 H_reg_52_ ( .D(n6102), .CK(clk), .RN(n17831), .Q(n17367), .QN() );
DFFR_X1 H_reg_51_ ( .D(n6103), .CK(clk), .RN(n17831), .Q(n17368), .QN() );
DFFR_X1 H_reg_50_ ( .D(n6104), .CK(clk), .RN(n17831), .Q(n17369), .QN() );
DFFR_X1 H_reg_49_ ( .D(n6105), .CK(clk), .RN(n17831), .Q(n17370), .QN() );
DFFR_X1 H_reg_48_ ( .D(n6106), .CK(clk), .RN(n17831), .Q(n17371), .QN() );
DFFR_X1 H_reg_47_ ( .D(n6107), .CK(clk), .RN(n17831), .Q(n17372), .QN() );
DFFR_X1 H_reg_46_ ( .D(n6108), .CK(clk), .RN(n17831), .Q(n17373), .QN() );
DFFR_X1 H_reg_45_ ( .D(n6109), .CK(clk), .RN(n17831), .Q(n17374), .QN() );
DFFR_X1 EkY0_reg_126_ ( .D(n6156), .CK(clk), .RN(n17832), .Q(), .QN(n17027));
DFFR_X1 EkY0_reg_125_ ( .D(n6157), .CK(clk), .RN(n17832), .Q(), .QN(n17029));
DFFR_X1 EkY0_reg_123_ ( .D(n6159), .CK(clk), .RN(n17832), .Q(), .QN(n17033));
DFFR_X1 EkY0_reg_121_ ( .D(n6161), .CK(clk), .RN(n17832), .Q(), .QN(n17037));
DFFR_X1 EkY0_reg_120_ ( .D(n6162), .CK(clk), .RN(n17832), .Q(), .QN(n17039));
DFFR_X1 EkY0_reg_119_ ( .D(n6163), .CK(clk), .RN(n17832), .Q(), .QN(n17041));
DFFR_X1 EkY0_reg_118_ ( .D(n6164), .CK(clk), .RN(n17832), .Q(), .QN(n17043));
DFFR_X1 EkY0_reg_117_ ( .D(n6165), .CK(clk), .RN(n17832), .Q(), .QN(n17045));
DFFR_X1 EkY0_reg_116_ ( .D(n6166), .CK(clk), .RN(n17832), .Q(), .QN(n17047));
DFFR_X1 EkY0_reg_115_ ( .D(n6167), .CK(clk), .RN(n17832), .Q(), .QN(n17049));
DFFR_X1 EkY0_reg_114_ ( .D(n6168), .CK(clk), .RN(n17833), .Q(), .QN(n17051));
DFFR_X1 EkY0_reg_113_ ( .D(n6169), .CK(clk), .RN(n17833), .Q(), .QN(n17053));
DFFR_X1 EkY0_reg_112_ ( .D(n6170), .CK(clk), .RN(n17833), .Q(), .QN(n17055));
DFFR_X1 EkY0_reg_111_ ( .D(n6171), .CK(clk), .RN(n17833), .Q(), .QN(n17057));
DFFR_X1 EkY0_reg_110_ ( .D(n6172), .CK(clk), .RN(n17833), .Q(), .QN(n17059));
DFFR_X1 EkY0_reg_109_ ( .D(n6173), .CK(clk), .RN(n17833), .Q(), .QN(n17061));
DFFR_X1 EkY0_reg_108_ ( .D(n6174), .CK(clk), .RN(n17833), .Q(), .QN(n17063));
DFFR_X1 EkY0_reg_107_ ( .D(n6175), .CK(clk), .RN(n17833), .Q(), .QN(n17065));
DFFR_X1 EkY0_reg_106_ ( .D(n6176), .CK(clk), .RN(n17833), .Q(), .QN(n17067));
DFFR_X1 EkY0_reg_105_ ( .D(n6177), .CK(clk), .RN(n17833), .Q(), .QN(n17069));
DFFR_X1 EkY0_reg_104_ ( .D(n6178), .CK(clk), .RN(n17833), .Q(), .QN(n17071));
DFFR_X1 EkY0_reg_103_ ( .D(n6179), .CK(clk), .RN(n17833), .Q(), .QN(n17073));
DFFR_X1 EkY0_reg_102_ ( .D(n6180), .CK(clk), .RN(n17834), .Q(), .QN(n17075));
DFFR_X1 EkY0_reg_101_ ( .D(n6181), .CK(clk), .RN(n17834), .Q(), .QN(n17077));
DFFR_X1 EkY0_reg_100_ ( .D(n6182), .CK(clk), .RN(n17834), .Q(), .QN(n17079));
DFFR_X1 EkY0_reg_99_ ( .D(n6183), .CK(clk), .RN(n17834), .Q(), .QN(n17081));
DFFR_X1 EkY0_reg_98_ ( .D(n6184), .CK(clk), .RN(n17834), .Q(), .QN(n17083));
DFFR_X1 EkY0_reg_97_ ( .D(n6185), .CK(clk), .RN(n17834), .Q(), .QN(n17085));
DFFR_X1 EkY0_reg_96_ ( .D(n6186), .CK(clk), .RN(n17834), .Q(), .QN(n17087));
DFFR_X1 EkY0_reg_95_ ( .D(n6187), .CK(clk), .RN(n17834), .Q(), .QN(n17089));
DFFR_X1 EkY0_reg_94_ ( .D(n6188), .CK(clk), .RN(n17834), .Q(), .QN(n17091));
DFFR_X1 EkY0_reg_93_ ( .D(n6189), .CK(clk), .RN(n17834), .Q(), .QN(n17093));
DFFR_X1 EkY0_reg_92_ ( .D(n6190), .CK(clk), .RN(n17834), .Q(), .QN(n17095));
DFFR_X1 EkY0_reg_91_ ( .D(n6191), .CK(clk), .RN(n17834), .Q(), .QN(n17097));
DFFR_X1 EkY0_reg_90_ ( .D(n6192), .CK(clk), .RN(n17835), .Q(), .QN(n17099));
DFFR_X1 EkY0_reg_89_ ( .D(n6193), .CK(clk), .RN(n17835), .Q(), .QN(n17101));
DFFR_X1 EkY0_reg_88_ ( .D(n6194), .CK(clk), .RN(n17835), .Q(), .QN(n17103));
DFFR_X1 EkY0_reg_87_ ( .D(n6195), .CK(clk), .RN(n17835), .Q(), .QN(n17105));
DFFR_X1 EkY0_reg_86_ ( .D(n6196), .CK(clk), .RN(n17835), .Q(), .QN(n17107));
DFFR_X1 EkY0_reg_85_ ( .D(n6197), .CK(clk), .RN(n17835), .Q(), .QN(n17109));
DFFR_X1 EkY0_reg_84_ ( .D(n6198), .CK(clk), .RN(n17835), .Q(), .QN(n17111));
DFFR_X1 EkY0_reg_83_ ( .D(n6199), .CK(clk), .RN(n17835), .Q(), .QN(n17113));
DFFR_X1 EkY0_reg_82_ ( .D(n6200), .CK(clk), .RN(n17835), .Q(), .QN(n17115));
DFFR_X1 EkY0_reg_81_ ( .D(n6201), .CK(clk), .RN(n17835), .Q(), .QN(n17117));
DFFR_X1 EkY0_reg_80_ ( .D(n6202), .CK(clk), .RN(n17835), .Q(), .QN(n17119));
DFFR_X1 EkY0_reg_79_ ( .D(n6203), .CK(clk), .RN(n17835), .Q(), .QN(n17121));
DFFR_X1 EkY0_reg_78_ ( .D(n6204), .CK(clk), .RN(n17836), .Q(), .QN(n17123));
DFFR_X1 EkY0_reg_77_ ( .D(n6205), .CK(clk), .RN(n17836), .Q(), .QN(n17125));
DFFR_X1 EkY0_reg_76_ ( .D(n6206), .CK(clk), .RN(n17836), .Q(), .QN(n17127));
DFFR_X1 EkY0_reg_75_ ( .D(n6207), .CK(clk), .RN(n17836), .Q(), .QN(n17129));
DFFR_X1 EkY0_reg_74_ ( .D(n6208), .CK(clk), .RN(n17836), .Q(), .QN(n17131));
DFFR_X1 EkY0_reg_73_ ( .D(n6209), .CK(clk), .RN(n17836), .Q(), .QN(n17133));
DFFR_X1 EkY0_reg_72_ ( .D(n6210), .CK(clk), .RN(n17836), .Q(), .QN(n17135));
DFFR_X1 EkY0_reg_71_ ( .D(n6211), .CK(clk), .RN(n17836), .Q(), .QN(n17137));
DFFR_X1 EkY0_reg_70_ ( .D(n6212), .CK(clk), .RN(n17836), .Q(), .QN(n17139));
DFFR_X1 EkY0_reg_69_ ( .D(n6213), .CK(clk), .RN(n17751), .Q(), .QN(n17141));
DFFR_X1 EkY0_reg_68_ ( .D(n6214), .CK(clk), .RN(n17818), .Q(), .QN(n17143));
DFFR_X1 EkY0_reg_67_ ( .D(n6215), .CK(clk), .RN(n17818), .Q(), .QN(n17145));
DFFR_X1 EkY0_reg_66_ ( .D(n6216), .CK(clk), .RN(n17818), .Q(), .QN(n17147));
DFFR_X1 EkY0_reg_65_ ( .D(n6217), .CK(clk), .RN(n17818), .Q(), .QN(n17149));
DFFR_X1 EkY0_reg_64_ ( .D(n6218), .CK(clk), .RN(n17818), .Q(), .QN(n17151));
DFFR_X1 EkY0_reg_63_ ( .D(n6219), .CK(clk), .RN(n17818), .Q(), .QN(n17153));
DFFR_X1 EkY0_reg_62_ ( .D(n6220), .CK(clk), .RN(n17818), .Q(), .QN(n17155));
DFFR_X1 EkY0_reg_61_ ( .D(n6221), .CK(clk), .RN(n17818), .Q(), .QN(n17157));
DFFR_X1 EkY0_reg_60_ ( .D(n6222), .CK(clk), .RN(n17818), .Q(), .QN(n17159));
DFFR_X1 EkY0_reg_59_ ( .D(n6223), .CK(clk), .RN(n17818), .Q(), .QN(n17161));
DFFR_X1 EkY0_reg_58_ ( .D(n6224), .CK(clk), .RN(n17818), .Q(), .QN(n17163));
DFFR_X1 EkY0_reg_57_ ( .D(n6225), .CK(clk), .RN(n17819), .Q(), .QN(n17165));
DFFR_X1 EkY0_reg_56_ ( .D(n6226), .CK(clk), .RN(n17819), .Q(), .QN(n17167));
DFFR_X1 EkY0_reg_55_ ( .D(n6227), .CK(clk), .RN(n17819), .Q(), .QN(n17169));
DFFR_X1 EkY0_reg_54_ ( .D(n6228), .CK(clk), .RN(n17819), .Q(), .QN(n17171));
DFFR_X1 EkY0_reg_53_ ( .D(n6229), .CK(clk), .RN(n17819), .Q(), .QN(n17173));
DFFR_X1 EkY0_reg_52_ ( .D(n6230), .CK(clk), .RN(n17819), .Q(), .QN(n17175));
DFFR_X1 EkY0_reg_51_ ( .D(n6231), .CK(clk), .RN(n17819), .Q(), .QN(n17177));
DFFR_X1 EkY0_reg_43_ ( .D(n6239), .CK(clk), .RN(n17820), .Q(), .QN(n17193));
DFFR_X1 EkY0_reg_38_ ( .D(n6244), .CK(clk), .RN(n17820), .Q(), .QN(n17203));
DFFR_X1 EkY0_reg_37_ ( .D(n6245), .CK(clk), .RN(n17820), .Q(), .QN(n17205));
DFFR_X1 EkY0_reg_36_ ( .D(n6246), .CK(clk), .RN(n17820), .Q(), .QN(n17207));
DFFR_X1 EkY0_reg_35_ ( .D(n6247), .CK(clk), .RN(n17820), .Q(), .QN(n17209));
DFFR_X1 EkY0_reg_34_ ( .D(n6248), .CK(clk), .RN(n17820), .Q(), .QN(n17211));
DFFR_X1 EkY0_reg_33_ ( .D(n6249), .CK(clk), .RN(n17821), .Q(), .QN(n17213));
DFFR_X1 EkY0_reg_32_ ( .D(n6250), .CK(clk), .RN(n17821), .Q(), .QN(n17215));
DFFR_X1 EkY0_reg_31_ ( .D(n6251), .CK(clk), .RN(n17821), .Q(), .QN(n17217));
DFFR_X1 EkY0_reg_30_ ( .D(n6252), .CK(clk), .RN(n17821), .Q(), .QN(n17219));
DFFR_X1 EkY0_reg_29_ ( .D(n6253), .CK(clk), .RN(n17821), .Q(), .QN(n17221));
DFFR_X1 EkY0_reg_28_ ( .D(n6254), .CK(clk), .RN(n17821), .Q(), .QN(n17223));
DFFR_X1 EkY0_reg_27_ ( .D(n6255), .CK(clk), .RN(n17821), .Q(), .QN(n17225));
DFFR_X1 EkY0_reg_26_ ( .D(n6256), .CK(clk), .RN(n17821), .Q(), .QN(n17227));
DFFR_X1 EkY0_reg_25_ ( .D(n6257), .CK(clk), .RN(n17821), .Q(), .QN(n17229));
DFFR_X1 EkY0_reg_24_ ( .D(n6258), .CK(clk), .RN(n17821), .Q(), .QN(n17231));
DFFR_X1 EkY0_reg_23_ ( .D(n6259), .CK(clk), .RN(n17821), .Q(), .QN(n17233));
DFFR_X1 EkY0_reg_20_ ( .D(n6262), .CK(clk), .RN(n17822), .Q(), .QN(n17239));
DFFR_X1 EkY0_reg_17_ ( .D(n6265), .CK(clk), .RN(n17822), .Q(), .QN(n17245));
DFFR_X1 EkY0_reg_16_ ( .D(n6266), .CK(clk), .RN(n17822), .Q(), .QN(n17247));
DFFR_X1 EkY0_reg_15_ ( .D(n6267), .CK(clk), .RN(n17822), .Q(), .QN(n17249));
DFFR_X1 EkY0_reg_14_ ( .D(n6268), .CK(clk), .RN(n17822), .Q(), .QN(n17251));
DFFR_X1 EkY0_reg_13_ ( .D(n6269), .CK(clk), .RN(n17822), .Q(), .QN(n17253));
DFFR_X1 EkY0_reg_12_ ( .D(n6270), .CK(clk), .RN(n17822), .Q(), .QN(n17255));
DFFR_X1 EkY0_reg_11_ ( .D(n6271), .CK(clk), .RN(n17822), .Q(), .QN(n17257));
DFFR_X1 EkY0_reg_10_ ( .D(n6272), .CK(clk), .RN(n17822), .Q(), .QN(n17259));
DFFR_X1 EkY0_reg_9_ ( .D(n6273), .CK(clk), .RN(n17823), .Q(), .QN(n17261) );
DFFR_X1 EkY0_reg_8_ ( .D(n6274), .CK(clk), .RN(n17823), .Q(), .QN(n17263) );
DFFR_X1 EkY0_reg_7_ ( .D(n6275), .CK(clk), .RN(n17823), .Q(), .QN(n17265) );
DFFR_X1 EkY0_reg_6_ ( .D(n6276), .CK(clk), .RN(n17823), .Q(), .QN(n17267) );
DFFR_X1 EkY0_reg_5_ ( .D(n6277), .CK(clk), .RN(n17823), .Q(), .QN(n17269) );
DFFR_X1 EkY0_reg_4_ ( .D(n6278), .CK(clk), .RN(n17823), .Q(), .QN(n17271) );
DFFR_X1 EkY0_reg_3_ ( .D(n6279), .CK(clk), .RN(n17823), .Q(), .QN(n17273) );
DFFR_X1 EkY0_reg_0_ ( .D(n6282), .CK(clk), .RN(n17823), .Q(), .QN(n17279) );
DFF_X2 Yi_reg_98_ ( .D(n17744), .CK(clk), .Q(n18197), .QN(n5473) );
DFF_X2 Yi_reg_0_ ( .D(n5956), .CK(clk), .Q(n18589), .QN(n5571) );
DFF_X2 Yi_reg_1_ ( .D(n5955), .CK(clk), .Q(n18585), .QN(n5570) );
DFF_X2 Yi_reg_2_ ( .D(n5954), .CK(clk), .Q(n18581), .QN(n5569) );
DFF_X2 Yi_reg_3_ ( .D(n5953), .CK(clk), .Q(n18577), .QN(n5568) );
DFF_X2 Yi_reg_4_ ( .D(n5952), .CK(clk), .Q(n18573), .QN(n5567) );
DFF_X2 Yi_reg_5_ ( .D(n5951), .CK(clk), .Q(n18569), .QN(n5566) );
DFF_X2 Yi_reg_6_ ( .D(n5950), .CK(clk), .Q(n18565), .QN(n5565) );
DFF_X2 Yi_reg_7_ ( .D(n5949), .CK(clk), .Q(n18561), .QN(n5564) );
DFF_X2 Yi_reg_8_ ( .D(n5948), .CK(clk), .Q(n18557), .QN(n5563) );
DFF_X2 Yi_reg_9_ ( .D(n5947), .CK(clk), .Q(n18553), .QN(n5562) );
DFF_X2 Yi_reg_10_ ( .D(n5946), .CK(clk), .Q(n18549), .QN(n5561) );
DFF_X2 Yi_reg_11_ ( .D(n5945), .CK(clk), .Q(n18545), .QN(n5560) );
DFF_X2 Yi_reg_12_ ( .D(n5944), .CK(clk), .Q(n18541), .QN(n5559) );
DFF_X2 Yi_reg_13_ ( .D(n5943), .CK(clk), .Q(n18537), .QN(n5558) );
DFF_X2 Yi_reg_14_ ( .D(n5942), .CK(clk), .Q(n18533), .QN(n5557) );
DFF_X2 Yi_reg_15_ ( .D(n5941), .CK(clk), .Q(n18529), .QN(n5556) );
DFF_X2 Yi_reg_16_ ( .D(n17726), .CK(clk), .Q(n18525), .QN(n5555) );
DFF_X2 Yi_reg_17_ ( .D(n17724), .CK(clk), .Q(n18521), .QN(n5554) );
DFF_X2 Yi_reg_18_ ( .D(n17722), .CK(clk), .Q(n18517), .QN(n5553) );
DFF_X2 Yi_reg_19_ ( .D(n17720), .CK(clk), .Q(n18513), .QN(n5552) );
DFF_X2 Yi_reg_20_ ( .D(n17718), .CK(clk), .Q(n18509), .QN(n5551) );
DFF_X2 Yi_reg_21_ ( .D(n17716), .CK(clk), .Q(n18505), .QN(n5550) );
DFF_X2 Yi_reg_22_ ( .D(n17714), .CK(clk), .Q(n18501), .QN(n5549) );
DFF_X2 Yi_reg_23_ ( .D(n17712), .CK(clk), .Q(n18497), .QN(n5548) );
DFF_X2 Yi_reg_24_ ( .D(n17710), .CK(clk), .Q(n18493), .QN(n5547) );
DFF_X2 Yi_reg_25_ ( .D(n17708), .CK(clk), .Q(n18489), .QN(n5546) );
DFF_X2 Yi_reg_26_ ( .D(n17706), .CK(clk), .Q(n18485), .QN(n5545) );
DFF_X2 Yi_reg_27_ ( .D(n17704), .CK(clk), .Q(n18481), .QN(n5544) );
DFF_X2 Yi_reg_28_ ( .D(n17702), .CK(clk), .Q(n18477), .QN(n5543) );
DFF_X2 Yi_reg_29_ ( .D(n17700), .CK(clk), .Q(n18473), .QN(n5542) );
DFF_X2 Yi_reg_30_ ( .D(n17698), .CK(clk), .Q(n18469), .QN(n5541) );
DFF_X2 Yi_reg_31_ ( .D(n17696), .CK(clk), .Q(n18465), .QN(n5540) );
DFF_X2 Yi_reg_32_ ( .D(n17694), .CK(clk), .Q(n18461), .QN(n5539) );
DFF_X2 Yi_reg_33_ ( .D(n17692), .CK(clk), .Q(n18457), .QN(n5538) );
DFF_X2 Yi_reg_34_ ( .D(n17690), .CK(clk), .Q(n18453), .QN(n5537) );
DFF_X2 Yi_reg_35_ ( .D(n17688), .CK(clk), .Q(n18449), .QN(n5536) );
DFF_X2 Yi_reg_36_ ( .D(n17686), .CK(clk), .Q(n18445), .QN(n5535) );
DFF_X2 Yi_reg_37_ ( .D(n17684), .CK(clk), .Q(n18441), .QN(n5534) );
DFF_X2 Yi_reg_38_ ( .D(n17682), .CK(clk), .Q(n18437), .QN(n5533) );
DFF_X2 Yi_reg_39_ ( .D(n17680), .CK(clk), .Q(n18433), .QN(n5532) );
DFF_X2 Yi_reg_40_ ( .D(n17678), .CK(clk), .Q(n18429), .QN(n5531) );
DFF_X2 Yi_reg_41_ ( .D(n17676), .CK(clk), .Q(n18425), .QN(n5530) );
DFF_X2 Yi_reg_42_ ( .D(n17674), .CK(clk), .Q(n18421), .QN(n5529) );
DFF_X2 Yi_reg_43_ ( .D(n17672), .CK(clk), .Q(n18417), .QN(n5528) );
DFF_X2 Yi_reg_44_ ( .D(n17670), .CK(clk), .Q(n18413), .QN(n5527) );
DFF_X2 Yi_reg_45_ ( .D(n17668), .CK(clk), .Q(n18409), .QN(n5526) );
DFF_X2 Yi_reg_46_ ( .D(n17666), .CK(clk), .Q(n18405), .QN(n5525) );
DFF_X2 Yi_reg_47_ ( .D(n17664), .CK(clk), .Q(n18401), .QN(n5524) );
DFF_X2 Yi_reg_48_ ( .D(n17662), .CK(clk), .Q(n18397), .QN(n5523) );
DFF_X2 Yi_reg_49_ ( .D(n17660), .CK(clk), .Q(n18393), .QN(n5522) );
DFF_X2 Yi_reg_50_ ( .D(n17658), .CK(clk), .Q(n18389), .QN(n5521) );
DFF_X2 Yi_reg_51_ ( .D(n17656), .CK(clk), .Q(n18385), .QN(n5520) );
DFF_X2 Yi_reg_52_ ( .D(n17654), .CK(clk), .Q(n18381), .QN(n5519) );
DFF_X2 Yi_reg_53_ ( .D(n17652), .CK(clk), .Q(n18377), .QN(n5518) );
DFF_X2 Yi_reg_54_ ( .D(n17650), .CK(clk), .Q(n18373), .QN(n5517) );
DFF_X2 Yi_reg_55_ ( .D(n17648), .CK(clk), .Q(n18369), .QN(n5516) );
DFF_X2 Yi_reg_56_ ( .D(n17646), .CK(clk), .Q(n18365), .QN(n5515) );
DFF_X2 Yi_reg_57_ ( .D(n17644), .CK(clk), .Q(n18361), .QN(n5514) );
DFF_X2 Yi_reg_58_ ( .D(n17642), .CK(clk), .Q(n18357), .QN(n5513) );
DFF_X2 Yi_reg_59_ ( .D(n17640), .CK(clk), .Q(n18353), .QN(n5512) );
DFF_X2 Yi_reg_60_ ( .D(n17638), .CK(clk), .Q(n18349), .QN(n5511) );
DFF_X2 Yi_reg_61_ ( .D(n17636), .CK(clk), .Q(n18345), .QN(n5510) );
DFF_X2 Yi_reg_62_ ( .D(n17634), .CK(clk), .Q(n18341), .QN(n5509) );
DFF_X2 Yi_reg_63_ ( .D(n17632), .CK(clk), .Q(n18337), .QN(n5508) );
DFF_X2 Yi_reg_64_ ( .D(n17630), .CK(clk), .Q(n18333), .QN(n5507) );
DFF_X2 Yi_reg_65_ ( .D(n17628), .CK(clk), .Q(n18329), .QN(n5506) );
DFF_X2 Yi_reg_66_ ( .D(n17626), .CK(clk), .Q(n18325), .QN(n5505) );
DFF_X2 Yi_reg_67_ ( .D(n5889), .CK(clk), .Q(n18321), .QN(n5504) );
DFF_X2 Yi_reg_68_ ( .D(n5888), .CK(clk), .Q(n18317), .QN(n5503) );
DFF_X2 Yi_reg_69_ ( .D(n5887), .CK(clk), .Q(n18313), .QN(n5502) );
DFF_X2 Yi_reg_70_ ( .D(n5886), .CK(clk), .Q(n18309), .QN(n5501) );
DFF_X2 Yi_reg_71_ ( .D(n5885), .CK(clk), .Q(n18305), .QN(n5500) );
DFF_X2 Yi_reg_72_ ( .D(n17614), .CK(clk), .Q(n18301), .QN(n5499) );
DFF_X2 Yi_reg_73_ ( .D(n17612), .CK(clk), .Q(n18297), .QN(n5498) );
DFF_X2 Yi_reg_74_ ( .D(n17610), .CK(clk), .Q(n18293), .QN(n5497) );
DFF_X2 Yi_reg_75_ ( .D(n17608), .CK(clk), .Q(n18289), .QN(n5496) );
DFF_X2 Yi_reg_76_ ( .D(n17606), .CK(clk), .Q(n18285), .QN(n5495) );
DFF_X2 Yi_reg_77_ ( .D(n17604), .CK(clk), .Q(n18281), .QN(n5494) );
DFF_X2 Yi_reg_78_ ( .D(n17602), .CK(clk), .Q(n18277), .QN(n5493) );
DFF_X2 Yi_reg_79_ ( .D(n17600), .CK(clk), .Q(n18273), .QN(n5492) );
DFF_X2 Yi_reg_80_ ( .D(n17598), .CK(clk), .Q(n18269), .QN(n5491) );
DFF_X2 Yi_reg_81_ ( .D(n17596), .CK(clk), .Q(n18265), .QN(n5490) );
DFF_X2 Yi_reg_82_ ( .D(n17594), .CK(clk), .Q(n18261), .QN(n5489) );
DFF_X2 Yi_reg_83_ ( .D(n17592), .CK(clk), .Q(n18257), .QN(n5488) );
DFF_X2 Yi_reg_84_ ( .D(n17590), .CK(clk), .Q(n18253), .QN(n5487) );
DFF_X2 Yi_reg_85_ ( .D(n17588), .CK(clk), .Q(n18249), .QN(n5486) );
DFF_X2 Yi_reg_86_ ( .D(n17586), .CK(clk), .Q(n18245), .QN(n5485) );
DFF_X2 Yi_reg_87_ ( .D(n17584), .CK(clk), .Q(n18241), .QN(n5484) );
DFF_X2 Yi_reg_88_ ( .D(n17582), .CK(clk), .Q(n18237), .QN(n5483) );
DFF_X2 Yi_reg_89_ ( .D(n17580), .CK(clk), .Q(n18233), .QN(n5482) );
DFF_X2 Yi_reg_90_ ( .D(n17578), .CK(clk), .Q(n18229), .QN(n5481) );
DFF_X2 Yi_reg_91_ ( .D(n17576), .CK(clk), .Q(n18225), .QN(n5480) );
DFF_X2 Yi_reg_92_ ( .D(n17574), .CK(clk), .Q(n18221), .QN(n5479) );
DFF_X2 Yi_reg_93_ ( .D(n17572), .CK(clk), .Q(n18217), .QN(n5478) );
DFF_X2 Yi_reg_94_ ( .D(n17570), .CK(clk), .Q(n18213), .QN(n5477) );
DFF_X2 Yi_reg_95_ ( .D(n17568), .CK(clk), .Q(n18209), .QN(n5476) );
DFF_X2 Yi_reg_96_ ( .D(n17566), .CK(clk), .Q(n18205), .QN(n5475) );
DFF_X2 Yi_reg_97_ ( .D(n17564), .CK(clk), .Q(n18201), .QN(n5474) );
DFF_X2 Yi_reg_99_ ( .D(n17562), .CK(clk), .Q(n18193), .QN(n5472) );
DFF_X2 Yi_reg_100_ ( .D(n17560), .CK(clk), .Q(n18189), .QN(n5471) );
DFF_X2 Yi_reg_101_ ( .D(n17558), .CK(clk), .Q(n18185), .QN(n5470) );
DFF_X2 Yi_reg_102_ ( .D(n17556), .CK(clk), .Q(n18181), .QN(n5469) );
DFF_X2 Yi_reg_103_ ( .D(n17554), .CK(clk), .Q(n18177), .QN(n5468) );
DFF_X2 Yi_reg_104_ ( .D(n17552), .CK(clk), .Q(n18173), .QN(n5467) );
DFF_X2 Yi_reg_105_ ( .D(n17550), .CK(clk), .Q(n18169), .QN(n5466) );
DFF_X2 Yi_reg_106_ ( .D(n17548), .CK(clk), .Q(n18165), .QN(n5465) );
DFF_X2 Yi_reg_107_ ( .D(n17546), .CK(clk), .Q(n18161), .QN(n5464) );
DFF_X2 Yi_reg_108_ ( .D(n17544), .CK(clk), .Q(n18157), .QN(n5463) );
DFF_X2 Yi_reg_109_ ( .D(n17542), .CK(clk), .Q(n18153), .QN(n5462) );
DFF_X2 Yi_reg_110_ ( .D(n17540), .CK(clk), .Q(n18149), .QN(n5461) );
DFF_X2 Yi_reg_111_ ( .D(n17538), .CK(clk), .Q(n18145), .QN(n5460) );
DFF_X2 Yi_reg_112_ ( .D(n5845), .CK(clk), .Q(n18141), .QN(n5459) );
DFF_X2 Yi_reg_113_ ( .D(n5844), .CK(clk), .Q(n18137), .QN(n5458) );
DFF_X2 Yi_reg_114_ ( .D(n5843), .CK(clk), .Q(n18133), .QN(n5457) );
DFF_X2 Yi_reg_115_ ( .D(n5842), .CK(clk), .Q(n18129), .QN(n5456) );
DFF_X2 Yi_reg_116_ ( .D(n5841), .CK(clk), .Q(n18125), .QN(n5455) );
DFF_X2 Yi_reg_117_ ( .D(n5840), .CK(clk), .Q(n18121), .QN(n5454) );
DFF_X2 Yi_reg_118_ ( .D(n5839), .CK(clk), .Q(n18117), .QN(n5453) );
DFF_X2 Yi_reg_119_ ( .D(n5838), .CK(clk), .Q(n18113), .QN(n5452) );
DFF_X2 Yi_reg_120_ ( .D(n17521), .CK(clk), .Q(n18109), .QN(n5451) );
DFF_X2 Yi_reg_121_ ( .D(n17519), .CK(clk), .Q(n18105), .QN(n5450) );
DFF_X2 Yi_reg_122_ ( .D(n17517), .CK(clk), .Q(n18101), .QN(n5449) );
DFF_X2 Yi_reg_123_ ( .D(n17515), .CK(clk), .Q(n18097), .QN(n5448) );
DFF_X2 Yi_reg_124_ ( .D(n17513), .CK(clk), .Q(n18093), .QN(n5447) );
DFF_X2 Yi_reg_125_ ( .D(n17511), .CK(clk), .Q(n18089), .QN(n5446) );
DFF_X2 Yi_reg_126_ ( .D(n17509), .CK(clk), .Q(n18082), .QN(n5445) );
DFF_X2 Yi_reg_127_ ( .D(n17507), .CK(clk), .Q(n18593), .QN(n5444) );
DFF_X2 Tag_vld_reg ( .D(n17847), .CK(clk), .Q(Tag_vld), .QN() );
DFF_X2 Out_vld_reg ( .D(n17505), .CK(clk), .Q(Out_vld), .QN() );
DFF_X2 Out_last_word_reg ( .D(n6022), .CK(clk), .Q(Out_last_word), .QN() );
DFF_X2 Out_data_size_reg_3_ ( .D(n6023), .CK(clk), .Q(Out_data_size[3]),.QN() );
DFF_X2 Out_data_size_reg_2_ ( .D(n17504), .CK(clk), .Q(Out_data_size[2]),.QN() );
DFF_X2 Out_data_size_reg_1_ ( .D(n17503), .CK(clk), .Q(Out_data_size[1]),.QN() );
DFF_X2 Out_data_size_reg_0_ ( .D(n6026), .CK(clk), .Q(Out_data_size[0]),.QN() );
DFF_X2 gfm_cnt_reg_3_ ( .D(n6295), .CK(clk), .Q(n16839), .QN() );
DFF_X2 v_in_reg_0_ ( .D(N2815), .CK(clk), .Q(v_in[0]), .QN() );
DFF_X2 Out_data_reg_0_ ( .D(n5701), .CK(clk), .Q(Out_data[0]), .QN() );
DFF_X2 b_in_reg_0_ ( .D(N3071), .CK(clk), .Q(b_in[0]), .QN() );
DFF_X2 z_in_reg_0_ ( .D(N2943), .CK(clk), .Q(z_in[0]), .QN() );
DFF_X2 Out_data_reg_1_ ( .D(n5700), .CK(clk), .Q(Out_data[1]), .QN() );
DFF_X2 b_in_reg_1_ ( .D(N3072), .CK(clk), .Q(b_in[1]), .QN() );
DFF_X2 z_in_reg_1_ ( .D(N2944), .CK(clk), .Q(z_in[1]), .QN() );
DFF_X2 Out_data_reg_2_ ( .D(n5699), .CK(clk), .Q(Out_data[2]), .QN() );
DFF_X2 b_in_reg_2_ ( .D(N3073), .CK(clk), .Q(b_in[2]), .QN() );
DFF_X2 z_in_reg_2_ ( .D(N2945), .CK(clk), .Q(z_in[2]), .QN() );
DFF_X2 Out_data_reg_3_ ( .D(n5698), .CK(clk), .Q(Out_data[3]), .QN() );
DFF_X2 b_in_reg_3_ ( .D(N3074), .CK(clk), .Q(b_in[3]), .QN() );
DFF_X2 z_in_reg_3_ ( .D(N2946), .CK(clk), .Q(z_in[3]), .QN() );
DFF_X2 Out_data_reg_4_ ( .D(n5697), .CK(clk), .Q(Out_data[4]), .QN() );
DFF_X2 b_in_reg_4_ ( .D(N3075), .CK(clk), .Q(b_in[4]), .QN() );
DFF_X2 z_in_reg_4_ ( .D(N2947), .CK(clk), .Q(z_in[4]), .QN() );
DFF_X2 Out_data_reg_5_ ( .D(n5696), .CK(clk), .Q(Out_data[5]), .QN() );
DFF_X2 b_in_reg_5_ ( .D(N3076), .CK(clk), .Q(b_in[5]), .QN() );
DFF_X2 z_in_reg_5_ ( .D(N2948), .CK(clk), .Q(z_in[5]), .QN() );
DFF_X2 Out_data_reg_6_ ( .D(n5695), .CK(clk), .Q(Out_data[6]), .QN() );
DFF_X2 b_in_reg_6_ ( .D(N3077), .CK(clk), .Q(b_in[6]), .QN() );
DFF_X2 z_in_reg_6_ ( .D(N2949), .CK(clk), .Q(z_in[6]), .QN() );
DFF_X2 Out_data_reg_7_ ( .D(n5694), .CK(clk), .Q(Out_data[7]), .QN() );
DFF_X2 b_in_reg_7_ ( .D(N3078), .CK(clk), .Q(b_in[7]), .QN() );
DFF_X2 z_in_reg_7_ ( .D(N2950), .CK(clk), .Q(z_in[7]), .QN() );
DFF_X2 Out_data_reg_8_ ( .D(n5693), .CK(clk), .Q(Out_data[8]), .QN() );
DFF_X2 b_in_reg_8_ ( .D(N3079), .CK(clk), .Q(b_in[8]), .QN() );
DFF_X2 z_in_reg_8_ ( .D(N2951), .CK(clk), .Q(z_in[8]), .QN() );
DFF_X2 Out_data_reg_9_ ( .D(n5692), .CK(clk), .Q(Out_data[9]), .QN() );
DFF_X2 b_in_reg_9_ ( .D(N3080), .CK(clk), .Q(b_in[9]), .QN() );
DFF_X2 z_in_reg_9_ ( .D(N2952), .CK(clk), .Q(z_in[9]), .QN() );
DFF_X2 Out_data_reg_10_ ( .D(n5691), .CK(clk), .Q(Out_data[10]), .QN() );
DFF_X2 b_in_reg_10_ ( .D(N3081), .CK(clk), .Q(b_in[10]), .QN() );
DFF_X2 z_in_reg_10_ ( .D(N2953), .CK(clk), .Q(z_in[10]), .QN() );
DFF_X2 Out_data_reg_11_ ( .D(n5690), .CK(clk), .Q(Out_data[11]), .QN() );
DFF_X2 b_in_reg_11_ ( .D(N3082), .CK(clk), .Q(b_in[11]), .QN() );
DFF_X2 z_in_reg_11_ ( .D(N2954), .CK(clk), .Q(z_in[11]), .QN() );
DFF_X2 Out_data_reg_12_ ( .D(n5689), .CK(clk), .Q(Out_data[12]), .QN() );
DFF_X2 b_in_reg_12_ ( .D(N3083), .CK(clk), .Q(b_in[12]), .QN() );
DFF_X2 z_in_reg_12_ ( .D(N2955), .CK(clk), .Q(z_in[12]), .QN() );
DFF_X2 Out_data_reg_13_ ( .D(n5688), .CK(clk), .Q(Out_data[13]), .QN() );
DFF_X2 b_in_reg_13_ ( .D(N3084), .CK(clk), .Q(b_in[13]), .QN() );
DFF_X2 z_in_reg_13_ ( .D(N2956), .CK(clk), .Q(z_in[13]), .QN() );
DFF_X2 Out_data_reg_14_ ( .D(n5687), .CK(clk), .Q(Out_data[14]), .QN() );
DFF_X2 b_in_reg_14_ ( .D(N3085), .CK(clk), .Q(b_in[14]), .QN() );
DFF_X2 z_in_reg_14_ ( .D(N2957), .CK(clk), .Q(z_in[14]), .QN() );
DFF_X2 Out_data_reg_15_ ( .D(n5686), .CK(clk), .Q(Out_data[15]), .QN() );
DFF_X2 b_in_reg_15_ ( .D(N3086), .CK(clk), .Q(b_in[15]), .QN() );
DFF_X2 z_in_reg_15_ ( .D(N2958), .CK(clk), .Q(z_in[15]), .QN() );
DFF_X2 Out_data_reg_16_ ( .D(n5685), .CK(clk), .Q(Out_data[16]), .QN() );
DFF_X2 b_in_reg_16_ ( .D(N3087), .CK(clk), .Q(b_in[16]), .QN() );
DFF_X2 z_in_reg_16_ ( .D(N2959), .CK(clk), .Q(z_in[16]), .QN() );
DFF_X2 Out_data_reg_17_ ( .D(n5684), .CK(clk), .Q(Out_data[17]), .QN() );
DFF_X2 b_in_reg_17_ ( .D(N3088), .CK(clk), .Q(b_in[17]), .QN() );
DFF_X2 z_in_reg_17_ ( .D(N2960), .CK(clk), .Q(z_in[17]), .QN() );
DFF_X2 Out_data_reg_18_ ( .D(n5683), .CK(clk), .Q(Out_data[18]), .QN() );
DFF_X2 b_in_reg_18_ ( .D(N3089), .CK(clk), .Q(b_in[18]), .QN() );
DFF_X2 z_in_reg_18_ ( .D(N2961), .CK(clk), .Q(z_in[18]), .QN() );
DFF_X2 Out_data_reg_19_ ( .D(n5682), .CK(clk), .Q(Out_data[19]), .QN() );
DFF_X2 b_in_reg_19_ ( .D(N3090), .CK(clk), .Q(b_in[19]), .QN() );
DFF_X2 z_in_reg_19_ ( .D(N2962), .CK(clk), .Q(z_in[19]), .QN() );
DFF_X2 Out_data_reg_20_ ( .D(n5681), .CK(clk), .Q(Out_data[20]), .QN() );
DFF_X2 b_in_reg_20_ ( .D(N3091), .CK(clk), .Q(b_in[20]), .QN() );
DFF_X2 z_in_reg_20_ ( .D(N2963), .CK(clk), .Q(z_in[20]), .QN() );
DFF_X2 Out_data_reg_21_ ( .D(n5680), .CK(clk), .Q(Out_data[21]), .QN() );
DFF_X2 b_in_reg_21_ ( .D(N3092), .CK(clk), .Q(b_in[21]), .QN() );
DFF_X2 z_in_reg_21_ ( .D(N2964), .CK(clk), .Q(z_in[21]), .QN() );
DFF_X2 Out_data_reg_22_ ( .D(n5679), .CK(clk), .Q(Out_data[22]), .QN() );
DFF_X2 b_in_reg_22_ ( .D(N3093), .CK(clk), .Q(b_in[22]), .QN() );
DFF_X2 z_in_reg_22_ ( .D(N2965), .CK(clk), .Q(z_in[22]), .QN() );
DFF_X2 Out_data_reg_23_ ( .D(n5678), .CK(clk), .Q(Out_data[23]), .QN() );
DFF_X2 b_in_reg_23_ ( .D(N3094), .CK(clk), .Q(b_in[23]), .QN() );
DFF_X2 z_in_reg_23_ ( .D(N2966), .CK(clk), .Q(z_in[23]), .QN() );
DFF_X2 Out_data_reg_24_ ( .D(n5677), .CK(clk), .Q(Out_data[24]), .QN() );
DFF_X2 b_in_reg_24_ ( .D(N3095), .CK(clk), .Q(b_in[24]), .QN() );
DFF_X2 z_in_reg_24_ ( .D(N2967), .CK(clk), .Q(z_in[24]), .QN() );
DFF_X2 Out_data_reg_25_ ( .D(n5676), .CK(clk), .Q(Out_data[25]), .QN() );
DFF_X2 b_in_reg_25_ ( .D(N3096), .CK(clk), .Q(b_in[25]), .QN() );
DFF_X2 z_in_reg_25_ ( .D(N2968), .CK(clk), .Q(z_in[25]), .QN() );
DFF_X2 Out_data_reg_26_ ( .D(n5675), .CK(clk), .Q(Out_data[26]), .QN() );
DFF_X2 b_in_reg_26_ ( .D(N3097), .CK(clk), .Q(b_in[26]), .QN() );
DFF_X2 z_in_reg_26_ ( .D(N2969), .CK(clk), .Q(z_in[26]), .QN() );
DFF_X2 Out_data_reg_27_ ( .D(n5674), .CK(clk), .Q(Out_data[27]), .QN() );
DFF_X2 b_in_reg_27_ ( .D(N3098), .CK(clk), .Q(b_in[27]), .QN() );
DFF_X2 z_in_reg_27_ ( .D(N2970), .CK(clk), .Q(z_in[27]), .QN() );
DFF_X2 Out_data_reg_28_ ( .D(n5673), .CK(clk), .Q(Out_data[28]), .QN() );
DFF_X2 b_in_reg_28_ ( .D(N3099), .CK(clk), .Q(b_in[28]), .QN() );
DFF_X2 z_in_reg_28_ ( .D(N2971), .CK(clk), .Q(z_in[28]), .QN() );
DFF_X2 Out_data_reg_29_ ( .D(n5672), .CK(clk), .Q(Out_data[29]), .QN() );
DFF_X2 b_in_reg_29_ ( .D(N3100), .CK(clk), .Q(b_in[29]), .QN() );
DFF_X2 z_in_reg_29_ ( .D(N2972), .CK(clk), .Q(z_in[29]), .QN() );
DFF_X2 Out_data_reg_30_ ( .D(n5671), .CK(clk), .Q(Out_data[30]), .QN() );
DFF_X2 b_in_reg_30_ ( .D(N3101), .CK(clk), .Q(b_in[30]), .QN() );
DFF_X2 z_in_reg_30_ ( .D(N2973), .CK(clk), .Q(z_in[30]), .QN() );
DFF_X2 Out_data_reg_31_ ( .D(n5670), .CK(clk), .Q(Out_data[31]), .QN() );
DFF_X2 b_in_reg_31_ ( .D(N3102), .CK(clk), .Q(b_in[31]), .QN() );
DFF_X2 z_in_reg_31_ ( .D(N2974), .CK(clk), .Q(z_in[31]), .QN() );
DFF_X2 Out_data_reg_32_ ( .D(n5669), .CK(clk), .Q(Out_data[32]), .QN() );
DFF_X2 b_in_reg_32_ ( .D(N3103), .CK(clk), .Q(b_in[32]), .QN() );
DFF_X2 z_in_reg_32_ ( .D(N2975), .CK(clk), .Q(z_in[32]), .QN() );
DFF_X2 Out_data_reg_33_ ( .D(n5668), .CK(clk), .Q(Out_data[33]), .QN() );
DFF_X2 b_in_reg_33_ ( .D(N3104), .CK(clk), .Q(b_in[33]), .QN() );
DFF_X2 z_in_reg_33_ ( .D(N2976), .CK(clk), .Q(z_in[33]), .QN() );
DFF_X2 Out_data_reg_34_ ( .D(n5667), .CK(clk), .Q(Out_data[34]), .QN() );
DFF_X2 b_in_reg_34_ ( .D(N3105), .CK(clk), .Q(b_in[34]), .QN() );
DFF_X2 z_in_reg_34_ ( .D(N2977), .CK(clk), .Q(z_in[34]), .QN() );
DFF_X2 Out_data_reg_35_ ( .D(n5666), .CK(clk), .Q(Out_data[35]), .QN() );
DFF_X2 b_in_reg_35_ ( .D(N3106), .CK(clk), .Q(b_in[35]), .QN() );
DFF_X2 z_in_reg_35_ ( .D(N2978), .CK(clk), .Q(z_in[35]), .QN() );
DFF_X2 Out_data_reg_36_ ( .D(n5665), .CK(clk), .Q(Out_data[36]), .QN() );
DFF_X2 b_in_reg_36_ ( .D(N3107), .CK(clk), .Q(b_in[36]), .QN() );
DFF_X2 z_in_reg_36_ ( .D(N2979), .CK(clk), .Q(z_in[36]), .QN() );
DFF_X2 Out_data_reg_37_ ( .D(n5664), .CK(clk), .Q(Out_data[37]), .QN() );
DFF_X2 b_in_reg_37_ ( .D(N3108), .CK(clk), .Q(b_in[37]), .QN() );
DFF_X2 z_in_reg_37_ ( .D(N2980), .CK(clk), .Q(z_in[37]), .QN() );
DFF_X2 Out_data_reg_38_ ( .D(n5663), .CK(clk), .Q(Out_data[38]), .QN() );
DFF_X2 b_in_reg_38_ ( .D(N3109), .CK(clk), .Q(b_in[38]), .QN() );
DFF_X2 z_in_reg_38_ ( .D(N2981), .CK(clk), .Q(z_in[38]), .QN() );
DFF_X2 Out_data_reg_39_ ( .D(n5662), .CK(clk), .Q(Out_data[39]), .QN() );
DFF_X2 b_in_reg_39_ ( .D(N3110), .CK(clk), .Q(b_in[39]), .QN() );
DFF_X2 z_in_reg_39_ ( .D(N2982), .CK(clk), .Q(z_in[39]), .QN() );
DFF_X2 Out_data_reg_40_ ( .D(n5661), .CK(clk), .Q(Out_data[40]), .QN() );
DFF_X2 b_in_reg_40_ ( .D(N3111), .CK(clk), .Q(b_in[40]), .QN() );
DFF_X2 z_in_reg_40_ ( .D(N2983), .CK(clk), .Q(z_in[40]), .QN() );
DFF_X2 Out_data_reg_41_ ( .D(n5660), .CK(clk), .Q(Out_data[41]), .QN() );
DFF_X2 b_in_reg_41_ ( .D(N3112), .CK(clk), .Q(b_in[41]), .QN() );
DFF_X2 z_in_reg_41_ ( .D(N2984), .CK(clk), .Q(z_in[41]), .QN() );
DFF_X2 Out_data_reg_42_ ( .D(n5659), .CK(clk), .Q(Out_data[42]), .QN() );
DFF_X2 b_in_reg_42_ ( .D(N3113), .CK(clk), .Q(b_in[42]), .QN() );
DFF_X2 z_in_reg_42_ ( .D(N2985), .CK(clk), .Q(z_in[42]), .QN() );
DFF_X2 Out_data_reg_43_ ( .D(n5658), .CK(clk), .Q(Out_data[43]), .QN() );
DFF_X2 b_in_reg_43_ ( .D(N3114), .CK(clk), .Q(b_in[43]), .QN() );
DFF_X2 z_in_reg_43_ ( .D(N2986), .CK(clk), .Q(z_in[43]), .QN() );
DFF_X2 Out_data_reg_44_ ( .D(n5657), .CK(clk), .Q(Out_data[44]), .QN() );
DFF_X2 b_in_reg_44_ ( .D(N3115), .CK(clk), .Q(b_in[44]), .QN() );
DFF_X2 z_in_reg_44_ ( .D(N2987), .CK(clk), .Q(z_in[44]), .QN() );
DFF_X2 Out_data_reg_45_ ( .D(n5656), .CK(clk), .Q(Out_data[45]), .QN() );
DFF_X2 b_in_reg_45_ ( .D(N3116), .CK(clk), .Q(b_in[45]), .QN() );
DFF_X2 z_in_reg_45_ ( .D(N2988), .CK(clk), .Q(z_in[45]), .QN() );
DFF_X2 Out_data_reg_46_ ( .D(n5655), .CK(clk), .Q(Out_data[46]), .QN() );
DFF_X2 b_in_reg_46_ ( .D(N3117), .CK(clk), .Q(b_in[46]), .QN() );
DFF_X2 z_in_reg_46_ ( .D(N2989), .CK(clk), .Q(z_in[46]), .QN() );
DFF_X2 Out_data_reg_47_ ( .D(n5654), .CK(clk), .Q(Out_data[47]), .QN() );
DFF_X2 b_in_reg_47_ ( .D(N3118), .CK(clk), .Q(b_in[47]), .QN() );
DFF_X2 z_in_reg_47_ ( .D(N2990), .CK(clk), .Q(z_in[47]), .QN() );
DFF_X2 Out_data_reg_48_ ( .D(n5653), .CK(clk), .Q(Out_data[48]), .QN() );
DFF_X2 b_in_reg_48_ ( .D(N3119), .CK(clk), .Q(b_in[48]), .QN() );
DFF_X2 z_in_reg_48_ ( .D(N2991), .CK(clk), .Q(z_in[48]), .QN() );
DFF_X2 Out_data_reg_49_ ( .D(n5652), .CK(clk), .Q(Out_data[49]), .QN() );
DFF_X2 b_in_reg_49_ ( .D(N3120), .CK(clk), .Q(b_in[49]), .QN() );
DFF_X2 z_in_reg_49_ ( .D(N2992), .CK(clk), .Q(z_in[49]), .QN() );
DFF_X2 Out_data_reg_50_ ( .D(n5651), .CK(clk), .Q(Out_data[50]), .QN() );
DFF_X2 b_in_reg_50_ ( .D(N3121), .CK(clk), .Q(b_in[50]), .QN() );
DFF_X2 z_in_reg_50_ ( .D(N2993), .CK(clk), .Q(z_in[50]), .QN() );
DFF_X2 Out_data_reg_51_ ( .D(n5650), .CK(clk), .Q(Out_data[51]), .QN() );
DFF_X2 b_in_reg_51_ ( .D(N3122), .CK(clk), .Q(b_in[51]), .QN() );
DFF_X2 z_in_reg_51_ ( .D(N2994), .CK(clk), .Q(z_in[51]), .QN() );
DFF_X2 Out_data_reg_52_ ( .D(n5649), .CK(clk), .Q(Out_data[52]), .QN() );
DFF_X2 b_in_reg_52_ ( .D(N3123), .CK(clk), .Q(b_in[52]), .QN() );
DFF_X2 z_in_reg_52_ ( .D(N2995), .CK(clk), .Q(z_in[52]), .QN() );
DFF_X2 Out_data_reg_53_ ( .D(n5648), .CK(clk), .Q(Out_data[53]), .QN() );
DFF_X2 b_in_reg_53_ ( .D(N3124), .CK(clk), .Q(b_in[53]), .QN() );
DFF_X2 z_in_reg_53_ ( .D(N2996), .CK(clk), .Q(z_in[53]), .QN() );
DFF_X2 Out_data_reg_54_ ( .D(n5647), .CK(clk), .Q(Out_data[54]), .QN() );
DFF_X2 b_in_reg_54_ ( .D(N3125), .CK(clk), .Q(b_in[54]), .QN() );
DFF_X2 z_in_reg_54_ ( .D(N2997), .CK(clk), .Q(z_in[54]), .QN() );
DFF_X2 Out_data_reg_55_ ( .D(n5646), .CK(clk), .Q(Out_data[55]), .QN() );
DFF_X2 b_in_reg_55_ ( .D(N3126), .CK(clk), .Q(b_in[55]), .QN() );
DFF_X2 z_in_reg_55_ ( .D(N2998), .CK(clk), .Q(z_in[55]), .QN() );
DFF_X2 Out_data_reg_56_ ( .D(n5645), .CK(clk), .Q(Out_data[56]), .QN() );
DFF_X2 b_in_reg_56_ ( .D(N3127), .CK(clk), .Q(b_in[56]), .QN() );
DFF_X2 z_in_reg_56_ ( .D(N2999), .CK(clk), .Q(z_in[56]), .QN() );
DFF_X2 Out_data_reg_57_ ( .D(n5644), .CK(clk), .Q(Out_data[57]), .QN() );
DFF_X2 b_in_reg_57_ ( .D(N3128), .CK(clk), .Q(b_in[57]), .QN() );
DFF_X2 z_in_reg_57_ ( .D(N3000), .CK(clk), .Q(z_in[57]), .QN() );
DFF_X2 Out_data_reg_58_ ( .D(n5643), .CK(clk), .Q(Out_data[58]), .QN() );
DFF_X2 b_in_reg_58_ ( .D(N3129), .CK(clk), .Q(b_in[58]), .QN() );
DFF_X2 z_in_reg_58_ ( .D(N3001), .CK(clk), .Q(z_in[58]), .QN() );
DFF_X2 Out_data_reg_59_ ( .D(n5642), .CK(clk), .Q(Out_data[59]), .QN() );
DFF_X2 b_in_reg_59_ ( .D(N3130), .CK(clk), .Q(b_in[59]), .QN() );
DFF_X2 z_in_reg_59_ ( .D(N3002), .CK(clk), .Q(z_in[59]), .QN() );
DFF_X2 Out_data_reg_60_ ( .D(n5641), .CK(clk), .Q(Out_data[60]), .QN() );
DFF_X2 b_in_reg_60_ ( .D(N3131), .CK(clk), .Q(b_in[60]), .QN() );
DFF_X2 z_in_reg_60_ ( .D(N3003), .CK(clk), .Q(z_in[60]), .QN() );
DFF_X2 Out_data_reg_61_ ( .D(n5640), .CK(clk), .Q(Out_data[61]), .QN() );
DFF_X2 b_in_reg_61_ ( .D(N3132), .CK(clk), .Q(b_in[61]), .QN() );
DFF_X2 z_in_reg_61_ ( .D(N3004), .CK(clk), .Q(z_in[61]), .QN() );
DFF_X2 Out_data_reg_62_ ( .D(n5639), .CK(clk), .Q(Out_data[62]), .QN() );
DFF_X2 b_in_reg_62_ ( .D(N3133), .CK(clk), .Q(b_in[62]), .QN() );
DFF_X2 z_in_reg_62_ ( .D(N3005), .CK(clk), .Q(z_in[62]), .QN() );
DFF_X2 Out_data_reg_63_ ( .D(n5638), .CK(clk), .Q(Out_data[63]), .QN() );
DFF_X2 b_in_reg_63_ ( .D(N3134), .CK(clk), .Q(b_in[63]), .QN() );
DFF_X2 z_in_reg_63_ ( .D(N3006), .CK(clk), .Q(z_in[63]), .QN() );
DFF_X2 Out_data_reg_64_ ( .D(n5637), .CK(clk), .Q(Out_data[64]), .QN() );
DFF_X2 b_in_reg_64_ ( .D(N3135), .CK(clk), .Q(b_in[64]), .QN() );
DFF_X2 z_in_reg_64_ ( .D(N3007), .CK(clk), .Q(z_in[64]), .QN() );
DFF_X2 Out_data_reg_65_ ( .D(n5636), .CK(clk), .Q(Out_data[65]), .QN() );
DFF_X2 b_in_reg_65_ ( .D(N3136), .CK(clk), .Q(b_in[65]), .QN() );
DFF_X2 z_in_reg_65_ ( .D(N3008), .CK(clk), .Q(z_in[65]), .QN() );
DFF_X2 Out_data_reg_66_ ( .D(n5635), .CK(clk), .Q(Out_data[66]), .QN() );
DFF_X2 b_in_reg_66_ ( .D(N3137), .CK(clk), .Q(b_in[66]), .QN() );
DFF_X2 z_in_reg_66_ ( .D(N3009), .CK(clk), .Q(z_in[66]), .QN() );
DFF_X2 Out_data_reg_67_ ( .D(n5634), .CK(clk), .Q(Out_data[67]), .QN() );
DFF_X2 b_in_reg_67_ ( .D(N3138), .CK(clk), .Q(b_in[67]), .QN() );
DFF_X2 z_in_reg_67_ ( .D(N3010), .CK(clk), .Q(z_in[67]), .QN() );
DFF_X2 Out_data_reg_68_ ( .D(n5633), .CK(clk), .Q(Out_data[68]), .QN() );
DFF_X2 b_in_reg_68_ ( .D(N3139), .CK(clk), .Q(b_in[68]), .QN() );
DFF_X2 z_in_reg_68_ ( .D(N3011), .CK(clk), .Q(z_in[68]), .QN() );
DFF_X2 Out_data_reg_69_ ( .D(n5632), .CK(clk), .Q(Out_data[69]), .QN() );
DFF_X2 b_in_reg_69_ ( .D(N3140), .CK(clk), .Q(b_in[69]), .QN() );
DFF_X2 z_in_reg_69_ ( .D(N3012), .CK(clk), .Q(z_in[69]), .QN() );
DFF_X2 Out_data_reg_70_ ( .D(n5631), .CK(clk), .Q(Out_data[70]), .QN() );
DFF_X2 b_in_reg_70_ ( .D(N3141), .CK(clk), .Q(b_in[70]), .QN() );
DFF_X2 z_in_reg_70_ ( .D(N3013), .CK(clk), .Q(z_in[70]), .QN() );
DFF_X2 Out_data_reg_71_ ( .D(n5630), .CK(clk), .Q(Out_data[71]), .QN() );
DFF_X2 b_in_reg_71_ ( .D(N3142), .CK(clk), .Q(b_in[71]), .QN() );
DFF_X2 z_in_reg_71_ ( .D(N3014), .CK(clk), .Q(z_in[71]), .QN() );
DFF_X2 Out_data_reg_72_ ( .D(n5629), .CK(clk), .Q(Out_data[72]), .QN() );
DFF_X2 b_in_reg_72_ ( .D(N3143), .CK(clk), .Q(b_in[72]), .QN() );
DFF_X2 z_in_reg_72_ ( .D(N3015), .CK(clk), .Q(z_in[72]), .QN() );
DFF_X2 Out_data_reg_73_ ( .D(n5628), .CK(clk), .Q(Out_data[73]), .QN() );
DFF_X2 b_in_reg_73_ ( .D(N3144), .CK(clk), .Q(b_in[73]), .QN() );
DFF_X2 z_in_reg_73_ ( .D(N3016), .CK(clk), .Q(z_in[73]), .QN() );
DFF_X2 Out_data_reg_74_ ( .D(n5627), .CK(clk), .Q(Out_data[74]), .QN() );
DFF_X2 b_in_reg_74_ ( .D(N3145), .CK(clk), .Q(b_in[74]), .QN() );
DFF_X2 z_in_reg_74_ ( .D(N3017), .CK(clk), .Q(z_in[74]), .QN() );
DFF_X2 Out_data_reg_75_ ( .D(n5626), .CK(clk), .Q(Out_data[75]), .QN() );
DFF_X2 b_in_reg_75_ ( .D(N3146), .CK(clk), .Q(b_in[75]), .QN() );
DFF_X2 z_in_reg_75_ ( .D(N3018), .CK(clk), .Q(z_in[75]), .QN() );
DFF_X2 Out_data_reg_76_ ( .D(n5625), .CK(clk), .Q(Out_data[76]), .QN() );
DFF_X2 b_in_reg_76_ ( .D(N3147), .CK(clk), .Q(b_in[76]), .QN() );
DFF_X2 z_in_reg_76_ ( .D(N3019), .CK(clk), .Q(z_in[76]), .QN() );
DFF_X2 Out_data_reg_77_ ( .D(n5624), .CK(clk), .Q(Out_data[77]), .QN() );
DFF_X2 b_in_reg_77_ ( .D(N3148), .CK(clk), .Q(b_in[77]), .QN() );
DFF_X2 z_in_reg_77_ ( .D(N3020), .CK(clk), .Q(z_in[77]), .QN() );
DFF_X2 Out_data_reg_78_ ( .D(n5623), .CK(clk), .Q(Out_data[78]), .QN() );
DFF_X2 b_in_reg_78_ ( .D(N3149), .CK(clk), .Q(b_in[78]), .QN() );
DFF_X2 z_in_reg_78_ ( .D(N3021), .CK(clk), .Q(z_in[78]), .QN() );
DFF_X2 Out_data_reg_79_ ( .D(n5622), .CK(clk), .Q(Out_data[79]), .QN() );
DFF_X2 b_in_reg_79_ ( .D(N3150), .CK(clk), .Q(b_in[79]), .QN() );
DFF_X2 z_in_reg_79_ ( .D(N3022), .CK(clk), .Q(z_in[79]), .QN() );
DFF_X2 Out_data_reg_80_ ( .D(n5621), .CK(clk), .Q(Out_data[80]), .QN() );
DFF_X2 b_in_reg_80_ ( .D(N3151), .CK(clk), .Q(b_in[80]), .QN() );
DFF_X2 z_in_reg_80_ ( .D(N3023), .CK(clk), .Q(z_in[80]), .QN() );
DFF_X2 Out_data_reg_81_ ( .D(n5620), .CK(clk), .Q(Out_data[81]), .QN() );
DFF_X2 b_in_reg_81_ ( .D(N3152), .CK(clk), .Q(b_in[81]), .QN() );
DFF_X2 z_in_reg_81_ ( .D(N3024), .CK(clk), .Q(z_in[81]), .QN() );
DFF_X2 Out_data_reg_82_ ( .D(n5619), .CK(clk), .Q(Out_data[82]), .QN() );
DFF_X2 b_in_reg_82_ ( .D(N3153), .CK(clk), .Q(b_in[82]), .QN() );
DFF_X2 z_in_reg_82_ ( .D(N3025), .CK(clk), .Q(z_in[82]), .QN() );
DFF_X2 Out_data_reg_83_ ( .D(n5618), .CK(clk), .Q(Out_data[83]), .QN() );
DFF_X2 b_in_reg_83_ ( .D(N3154), .CK(clk), .Q(b_in[83]), .QN() );
DFF_X2 z_in_reg_83_ ( .D(N3026), .CK(clk), .Q(z_in[83]), .QN() );
DFF_X2 Out_data_reg_84_ ( .D(n5617), .CK(clk), .Q(Out_data[84]), .QN() );
DFF_X2 b_in_reg_84_ ( .D(N3155), .CK(clk), .Q(b_in[84]), .QN() );
DFF_X2 z_in_reg_84_ ( .D(N3027), .CK(clk), .Q(z_in[84]), .QN() );
DFF_X2 Out_data_reg_85_ ( .D(n5616), .CK(clk), .Q(Out_data[85]), .QN() );
DFF_X2 b_in_reg_85_ ( .D(N3156), .CK(clk), .Q(b_in[85]), .QN() );
DFF_X2 z_in_reg_85_ ( .D(N3028), .CK(clk), .Q(z_in[85]), .QN() );
DFF_X2 Out_data_reg_86_ ( .D(n5615), .CK(clk), .Q(Out_data[86]), .QN() );
DFF_X2 b_in_reg_86_ ( .D(N3157), .CK(clk), .Q(b_in[86]), .QN() );
DFF_X2 z_in_reg_86_ ( .D(N3029), .CK(clk), .Q(z_in[86]), .QN() );
DFF_X2 Out_data_reg_87_ ( .D(n5614), .CK(clk), .Q(Out_data[87]), .QN() );
DFF_X2 b_in_reg_87_ ( .D(N3158), .CK(clk), .Q(b_in[87]), .QN() );
DFF_X2 z_in_reg_87_ ( .D(N3030), .CK(clk), .Q(z_in[87]), .QN() );
DFF_X2 Out_data_reg_88_ ( .D(n5613), .CK(clk), .Q(Out_data[88]), .QN() );
DFF_X2 b_in_reg_88_ ( .D(N3159), .CK(clk), .Q(b_in[88]), .QN() );
DFF_X2 z_in_reg_88_ ( .D(N3031), .CK(clk), .Q(z_in[88]), .QN() );
DFF_X2 Out_data_reg_89_ ( .D(n5612), .CK(clk), .Q(Out_data[89]), .QN() );
DFF_X2 b_in_reg_89_ ( .D(N3160), .CK(clk), .Q(b_in[89]), .QN() );
DFF_X2 z_in_reg_89_ ( .D(N3032), .CK(clk), .Q(z_in[89]), .QN() );
DFF_X2 Out_data_reg_90_ ( .D(n5611), .CK(clk), .Q(Out_data[90]), .QN() );
DFF_X2 b_in_reg_90_ ( .D(N3161), .CK(clk), .Q(b_in[90]), .QN() );
DFF_X2 z_in_reg_90_ ( .D(N3033), .CK(clk), .Q(z_in[90]), .QN() );
DFF_X2 Out_data_reg_91_ ( .D(n5610), .CK(clk), .Q(Out_data[91]), .QN() );
DFF_X2 b_in_reg_91_ ( .D(N3162), .CK(clk), .Q(b_in[91]), .QN() );
DFF_X2 z_in_reg_91_ ( .D(N3034), .CK(clk), .Q(z_in[91]), .QN() );
DFF_X2 Out_data_reg_92_ ( .D(n5609), .CK(clk), .Q(Out_data[92]), .QN() );
DFF_X2 b_in_reg_92_ ( .D(N3163), .CK(clk), .Q(b_in[92]), .QN() );
DFF_X2 z_in_reg_92_ ( .D(N3035), .CK(clk), .Q(z_in[92]), .QN() );
DFF_X2 Out_data_reg_93_ ( .D(n5608), .CK(clk), .Q(Out_data[93]), .QN() );
DFF_X2 b_in_reg_93_ ( .D(N3164), .CK(clk), .Q(b_in[93]), .QN() );
DFF_X2 z_in_reg_93_ ( .D(N3036), .CK(clk), .Q(z_in[93]), .QN() );
DFF_X2 Out_data_reg_94_ ( .D(n5607), .CK(clk), .Q(Out_data[94]), .QN() );
DFF_X2 b_in_reg_94_ ( .D(N3165), .CK(clk), .Q(b_in[94]), .QN() );
DFF_X2 z_in_reg_94_ ( .D(N3037), .CK(clk), .Q(z_in[94]), .QN() );
DFF_X2 Out_data_reg_95_ ( .D(n5606), .CK(clk), .Q(Out_data[95]), .QN() );
DFF_X2 b_in_reg_95_ ( .D(N3166), .CK(clk), .Q(b_in[95]), .QN() );
DFF_X2 z_in_reg_95_ ( .D(N3038), .CK(clk), .Q(z_in[95]), .QN() );
DFF_X2 Out_data_reg_96_ ( .D(n5605), .CK(clk), .Q(Out_data[96]), .QN() );
DFF_X2 b_in_reg_96_ ( .D(N3167), .CK(clk), .Q(b_in[96]), .QN() );
DFF_X2 z_in_reg_96_ ( .D(N3039), .CK(clk), .Q(z_in[96]), .QN() );
DFF_X2 Out_data_reg_97_ ( .D(n5604), .CK(clk), .Q(Out_data[97]), .QN() );
DFF_X2 b_in_reg_97_ ( .D(N3168), .CK(clk), .Q(b_in[97]), .QN() );
DFF_X2 z_in_reg_97_ ( .D(N3040), .CK(clk), .Q(z_in[97]), .QN() );
DFF_X2 Out_data_reg_98_ ( .D(n5603), .CK(clk), .Q(Out_data[98]), .QN() );
DFF_X2 b_in_reg_98_ ( .D(N3169), .CK(clk), .Q(b_in[98]), .QN() );
DFF_X2 z_in_reg_98_ ( .D(N3041), .CK(clk), .Q(z_in[98]), .QN() );
DFF_X2 Out_data_reg_99_ ( .D(n5602), .CK(clk), .Q(Out_data[99]), .QN() );
DFF_X2 b_in_reg_99_ ( .D(N3170), .CK(clk), .Q(b_in[99]), .QN() );
DFF_X2 z_in_reg_99_ ( .D(N3042), .CK(clk), .Q(z_in[99]), .QN() );
DFF_X2 Out_data_reg_100_ ( .D(n5601), .CK(clk), .Q(Out_data[100]), .QN() );
DFF_X2 b_in_reg_100_ ( .D(N3171), .CK(clk), .Q(b_in[100]), .QN() );
DFF_X2 z_in_reg_100_ ( .D(N3043), .CK(clk), .Q(z_in[100]), .QN() );
DFF_X2 Out_data_reg_101_ ( .D(n5600), .CK(clk), .Q(Out_data[101]), .QN() );
DFF_X2 b_in_reg_101_ ( .D(N3172), .CK(clk), .Q(b_in[101]), .QN() );
DFF_X2 z_in_reg_101_ ( .D(N3044), .CK(clk), .Q(z_in[101]), .QN() );
DFF_X2 Out_data_reg_102_ ( .D(n5599), .CK(clk), .Q(Out_data[102]), .QN() );
DFF_X2 b_in_reg_102_ ( .D(N3173), .CK(clk), .Q(b_in[102]), .QN() );
DFF_X2 z_in_reg_102_ ( .D(N3045), .CK(clk), .Q(z_in[102]), .QN() );
DFF_X2 Out_data_reg_103_ ( .D(n5598), .CK(clk), .Q(Out_data[103]), .QN() );
DFF_X2 b_in_reg_103_ ( .D(N3174), .CK(clk), .Q(b_in[103]), .QN() );
DFF_X2 z_in_reg_103_ ( .D(N3046), .CK(clk), .Q(z_in[103]), .QN() );
DFF_X2 Out_data_reg_104_ ( .D(n5597), .CK(clk), .Q(Out_data[104]), .QN() );
DFF_X2 b_in_reg_104_ ( .D(N3175), .CK(clk), .Q(b_in[104]), .QN() );
DFF_X2 z_in_reg_104_ ( .D(N3047), .CK(clk), .Q(z_in[104]), .QN() );
DFF_X2 Out_data_reg_105_ ( .D(n5596), .CK(clk), .Q(Out_data[105]), .QN() );
DFF_X2 b_in_reg_105_ ( .D(N3176), .CK(clk), .Q(b_in[105]), .QN() );
DFF_X2 z_in_reg_105_ ( .D(N3048), .CK(clk), .Q(z_in[105]), .QN() );
DFF_X2 Out_data_reg_106_ ( .D(n5595), .CK(clk), .Q(Out_data[106]), .QN() );
DFF_X2 b_in_reg_106_ ( .D(N3177), .CK(clk), .Q(b_in[106]), .QN() );
DFF_X2 z_in_reg_106_ ( .D(N3049), .CK(clk), .Q(z_in[106]), .QN() );
DFF_X2 Out_data_reg_107_ ( .D(n5594), .CK(clk), .Q(Out_data[107]), .QN() );
DFF_X2 b_in_reg_107_ ( .D(N3178), .CK(clk), .Q(b_in[107]), .QN() );
DFF_X2 z_in_reg_107_ ( .D(N3050), .CK(clk), .Q(z_in[107]), .QN() );
DFF_X2 Out_data_reg_108_ ( .D(n5593), .CK(clk), .Q(Out_data[108]), .QN() );
DFF_X2 b_in_reg_108_ ( .D(N3179), .CK(clk), .Q(b_in[108]), .QN() );
DFF_X2 z_in_reg_108_ ( .D(N3051), .CK(clk), .Q(z_in[108]), .QN() );
DFF_X2 Out_data_reg_109_ ( .D(n5592), .CK(clk), .Q(Out_data[109]), .QN() );
DFF_X2 b_in_reg_109_ ( .D(N3180), .CK(clk), .Q(b_in[109]), .QN() );
DFF_X2 z_in_reg_109_ ( .D(N3052), .CK(clk), .Q(z_in[109]), .QN() );
DFF_X2 Out_data_reg_110_ ( .D(n5591), .CK(clk), .Q(Out_data[110]), .QN() );
DFF_X2 b_in_reg_110_ ( .D(N3181), .CK(clk), .Q(b_in[110]), .QN() );
DFF_X2 z_in_reg_110_ ( .D(N3053), .CK(clk), .Q(z_in[110]), .QN() );
DFF_X2 Out_data_reg_111_ ( .D(n5590), .CK(clk), .Q(Out_data[111]), .QN() );
DFF_X2 b_in_reg_111_ ( .D(N3182), .CK(clk), .Q(b_in[111]), .QN() );
DFF_X2 z_in_reg_111_ ( .D(N3054), .CK(clk), .Q(z_in[111]), .QN() );
DFF_X2 Out_data_reg_112_ ( .D(n5589), .CK(clk), .Q(Out_data[112]), .QN() );
DFF_X2 b_in_reg_112_ ( .D(N3183), .CK(clk), .Q(b_in[112]), .QN() );
DFF_X2 z_in_reg_112_ ( .D(N3055), .CK(clk), .Q(z_in[112]), .QN() );
DFF_X2 Out_data_reg_113_ ( .D(n5588), .CK(clk), .Q(Out_data[113]), .QN() );
DFF_X2 b_in_reg_113_ ( .D(N3184), .CK(clk), .Q(b_in[113]), .QN() );
DFF_X2 z_in_reg_113_ ( .D(N3056), .CK(clk), .Q(z_in[113]), .QN() );
DFF_X2 Out_data_reg_114_ ( .D(n5587), .CK(clk), .Q(Out_data[114]), .QN() );
DFF_X2 b_in_reg_114_ ( .D(N3185), .CK(clk), .Q(b_in[114]), .QN() );
DFF_X2 z_in_reg_114_ ( .D(N3057), .CK(clk), .Q(z_in[114]), .QN() );
DFF_X2 Out_data_reg_115_ ( .D(n5586), .CK(clk), .Q(Out_data[115]), .QN() );
DFF_X2 b_in_reg_115_ ( .D(N3186), .CK(clk), .Q(b_in[115]), .QN() );
DFF_X2 z_in_reg_115_ ( .D(N3058), .CK(clk), .Q(z_in[115]), .QN() );
DFF_X2 Out_data_reg_116_ ( .D(n5585), .CK(clk), .Q(Out_data[116]), .QN() );
DFF_X2 b_in_reg_116_ ( .D(N3187), .CK(clk), .Q(b_in[116]), .QN() );
DFF_X2 z_in_reg_116_ ( .D(N3059), .CK(clk), .Q(z_in[116]), .QN() );
DFF_X2 Out_data_reg_117_ ( .D(n5584), .CK(clk), .Q(Out_data[117]), .QN() );
DFF_X2 b_in_reg_117_ ( .D(N3188), .CK(clk), .Q(b_in[117]), .QN() );
DFF_X2 z_in_reg_117_ ( .D(N3060), .CK(clk), .Q(z_in[117]), .QN() );
DFF_X2 Out_data_reg_118_ ( .D(n5583), .CK(clk), .Q(Out_data[118]), .QN() );
DFF_X2 b_in_reg_118_ ( .D(N3189), .CK(clk), .Q(b_in[118]), .QN() );
DFF_X2 z_in_reg_118_ ( .D(N3061), .CK(clk), .Q(z_in[118]), .QN() );
DFF_X2 Out_data_reg_119_ ( .D(n5582), .CK(clk), .Q(Out_data[119]), .QN() );
DFF_X2 b_in_reg_119_ ( .D(N3190), .CK(clk), .Q(b_in[119]), .QN() );
DFF_X2 z_in_reg_119_ ( .D(N3062), .CK(clk), .Q(z_in[119]), .QN() );
DFF_X2 Out_data_reg_120_ ( .D(n5581), .CK(clk), .Q(Out_data[120]), .QN() );
DFF_X2 b_in_reg_120_ ( .D(N3191), .CK(clk), .Q(b_in[120]), .QN() );
DFF_X2 z_in_reg_120_ ( .D(N3063), .CK(clk), .Q(z_in[120]), .QN() );
DFF_X2 Out_data_reg_121_ ( .D(n5580), .CK(clk), .Q(Out_data[121]), .QN() );
DFF_X2 b_in_reg_121_ ( .D(N3192), .CK(clk), .Q(b_in[121]), .QN() );
DFF_X2 z_in_reg_121_ ( .D(N3064), .CK(clk), .Q(z_in[121]), .QN() );
DFF_X2 Out_data_reg_122_ ( .D(n5579), .CK(clk), .Q(Out_data[122]), .QN() );
DFF_X2 b_in_reg_122_ ( .D(N3193), .CK(clk), .Q(b_in[122]), .QN() );
DFF_X2 z_in_reg_122_ ( .D(N3065), .CK(clk), .Q(z_in[122]), .QN() );
DFF_X2 Out_data_reg_123_ ( .D(n5578), .CK(clk), .Q(Out_data[123]), .QN() );
DFF_X2 b_in_reg_123_ ( .D(N3194), .CK(clk), .Q(b_in[123]), .QN() );
DFF_X2 z_in_reg_123_ ( .D(N3066), .CK(clk), .Q(z_in[123]), .QN() );
DFF_X2 Out_data_reg_124_ ( .D(n5577), .CK(clk), .Q(Out_data[124]), .QN() );
DFF_X2 b_in_reg_124_ ( .D(N3195), .CK(clk), .Q(b_in[124]), .QN() );
DFF_X2 z_in_reg_124_ ( .D(N3067), .CK(clk), .Q(z_in[124]), .QN() );
DFF_X2 Out_data_reg_125_ ( .D(n5576), .CK(clk), .Q(Out_data[125]), .QN() );
DFF_X2 b_in_reg_125_ ( .D(N3196), .CK(clk), .Q(b_in[125]), .QN() );
DFF_X2 z_in_reg_125_ ( .D(N3068), .CK(clk), .Q(z_in[125]), .QN() );
DFF_X2 Out_data_reg_126_ ( .D(n5575), .CK(clk), .Q(Out_data[126]), .QN() );
DFF_X2 b_in_reg_126_ ( .D(N3197), .CK(clk), .Q(b_in[126]), .QN() );
DFF_X2 z_in_reg_126_ ( .D(N3069), .CK(clk), .Q(z_in[126]), .QN() );
DFF_X2 Out_data_reg_127_ ( .D(n5574), .CK(clk), .Q(Out_data[127]), .QN() );
DFF_X2 b_in_reg_127_ ( .D(N3198), .CK(clk), .Q(b_in[127]), .QN() );
DFF_X2 z_in_reg_127_ ( .D(N3070), .CK(clk), .Q(z_in[127]), .QN() );
DFF_X2 v_in_reg_1_ ( .D(N2816), .CK(clk), .Q(v_in[1]), .QN() );
DFF_X2 v_in_reg_2_ ( .D(N2817), .CK(clk), .Q(v_in[2]), .QN() );
DFF_X2 v_in_reg_3_ ( .D(N2818), .CK(clk), .Q(v_in[3]), .QN() );
DFF_X2 v_in_reg_4_ ( .D(N2819), .CK(clk), .Q(v_in[4]), .QN() );
DFF_X2 v_in_reg_5_ ( .D(N2820), .CK(clk), .Q(v_in[5]), .QN() );
DFF_X2 v_in_reg_6_ ( .D(N2821), .CK(clk), .Q(v_in[6]), .QN() );
DFF_X2 v_in_reg_7_ ( .D(N2822), .CK(clk), .Q(v_in[7]), .QN() );
DFF_X2 v_in_reg_8_ ( .D(N2823), .CK(clk), .Q(v_in[8]), .QN() );
DFF_X2 v_in_reg_9_ ( .D(N2824), .CK(clk), .Q(v_in[9]), .QN() );
DFF_X2 v_in_reg_10_ ( .D(N2825), .CK(clk), .Q(v_in[10]), .QN() );
DFF_X2 v_in_reg_11_ ( .D(N2826), .CK(clk), .Q(v_in[11]), .QN() );
DFF_X2 v_in_reg_12_ ( .D(N2827), .CK(clk), .Q(v_in[12]), .QN() );
DFF_X2 v_in_reg_13_ ( .D(N2828), .CK(clk), .Q(v_in[13]), .QN() );
DFF_X2 v_in_reg_14_ ( .D(N2829), .CK(clk), .Q(v_in[14]), .QN() );
DFF_X2 v_in_reg_15_ ( .D(N2830), .CK(clk), .Q(v_in[15]), .QN() );
DFF_X2 v_in_reg_16_ ( .D(N2831), .CK(clk), .Q(v_in[16]), .QN() );
DFF_X2 v_in_reg_17_ ( .D(N2832), .CK(clk), .Q(v_in[17]), .QN() );
DFF_X2 v_in_reg_18_ ( .D(N2833), .CK(clk), .Q(v_in[18]), .QN() );
DFF_X2 v_in_reg_19_ ( .D(N2834), .CK(clk), .Q(v_in[19]), .QN() );
DFF_X2 v_in_reg_20_ ( .D(N2835), .CK(clk), .Q(v_in[20]), .QN() );
DFF_X2 v_in_reg_21_ ( .D(N2836), .CK(clk), .Q(v_in[21]), .QN() );
DFF_X2 v_in_reg_22_ ( .D(N2837), .CK(clk), .Q(v_in[22]), .QN() );
DFF_X2 v_in_reg_23_ ( .D(N2838), .CK(clk), .Q(v_in[23]), .QN() );
DFF_X2 v_in_reg_24_ ( .D(N2839), .CK(clk), .Q(v_in[24]), .QN() );
DFF_X2 v_in_reg_25_ ( .D(N2840), .CK(clk), .Q(v_in[25]), .QN() );
DFF_X2 v_in_reg_26_ ( .D(N2841), .CK(clk), .Q(v_in[26]), .QN() );
DFF_X2 v_in_reg_27_ ( .D(N2842), .CK(clk), .Q(v_in[27]), .QN() );
DFF_X2 v_in_reg_28_ ( .D(N2843), .CK(clk), .Q(v_in[28]), .QN() );
DFF_X2 v_in_reg_29_ ( .D(N2844), .CK(clk), .Q(v_in[29]), .QN() );
DFF_X2 v_in_reg_30_ ( .D(N2845), .CK(clk), .Q(v_in[30]), .QN() );
DFF_X2 v_in_reg_31_ ( .D(N2846), .CK(clk), .Q(v_in[31]), .QN() );
DFF_X2 v_in_reg_32_ ( .D(N2847), .CK(clk), .Q(v_in[32]), .QN() );
DFF_X2 v_in_reg_33_ ( .D(N2848), .CK(clk), .Q(v_in[33]), .QN() );
DFF_X2 v_in_reg_34_ ( .D(N2849), .CK(clk), .Q(v_in[34]), .QN() );
DFF_X2 v_in_reg_35_ ( .D(N2850), .CK(clk), .Q(v_in[35]), .QN() );
DFF_X2 v_in_reg_36_ ( .D(N2851), .CK(clk), .Q(v_in[36]), .QN() );
DFF_X2 v_in_reg_37_ ( .D(N2852), .CK(clk), .Q(v_in[37]), .QN() );
DFF_X2 v_in_reg_38_ ( .D(N2853), .CK(clk), .Q(v_in[38]), .QN() );
DFF_X2 v_in_reg_39_ ( .D(N2854), .CK(clk), .Q(v_in[39]), .QN() );
DFF_X2 v_in_reg_40_ ( .D(N2855), .CK(clk), .Q(v_in[40]), .QN() );
DFF_X2 v_in_reg_41_ ( .D(N2856), .CK(clk), .Q(v_in[41]), .QN() );
DFF_X2 v_in_reg_42_ ( .D(N2857), .CK(clk), .Q(v_in[42]), .QN() );
DFF_X2 v_in_reg_43_ ( .D(N2858), .CK(clk), .Q(v_in[43]), .QN() );
DFF_X2 v_in_reg_44_ ( .D(N2859), .CK(clk), .Q(v_in[44]), .QN() );
DFF_X2 v_in_reg_45_ ( .D(N2860), .CK(clk), .Q(v_in[45]), .QN() );
DFF_X2 v_in_reg_46_ ( .D(N2861), .CK(clk), .Q(v_in[46]), .QN() );
DFF_X2 v_in_reg_47_ ( .D(N2862), .CK(clk), .Q(v_in[47]), .QN() );
DFF_X2 v_in_reg_48_ ( .D(N2863), .CK(clk), .Q(v_in[48]), .QN() );
DFF_X2 v_in_reg_49_ ( .D(N2864), .CK(clk), .Q(v_in[49]), .QN() );
DFF_X2 v_in_reg_50_ ( .D(N2865), .CK(clk), .Q(v_in[50]), .QN() );
DFF_X2 v_in_reg_51_ ( .D(N2866), .CK(clk), .Q(v_in[51]), .QN() );
DFF_X2 v_in_reg_52_ ( .D(N2867), .CK(clk), .Q(v_in[52]), .QN() );
DFF_X2 v_in_reg_53_ ( .D(N2868), .CK(clk), .Q(v_in[53]), .QN() );
DFF_X2 v_in_reg_54_ ( .D(N2869), .CK(clk), .Q(v_in[54]), .QN() );
DFF_X2 v_in_reg_55_ ( .D(N2870), .CK(clk), .Q(v_in[55]), .QN() );
DFF_X2 v_in_reg_56_ ( .D(N2871), .CK(clk), .Q(v_in[56]), .QN() );
DFF_X2 v_in_reg_57_ ( .D(N2872), .CK(clk), .Q(v_in[57]), .QN() );
DFF_X2 v_in_reg_58_ ( .D(N2873), .CK(clk), .Q(v_in[58]), .QN() );
DFF_X2 v_in_reg_59_ ( .D(N2874), .CK(clk), .Q(v_in[59]), .QN() );
DFF_X2 v_in_reg_60_ ( .D(N2875), .CK(clk), .Q(v_in[60]), .QN() );
DFF_X2 v_in_reg_61_ ( .D(N2876), .CK(clk), .Q(v_in[61]), .QN() );
DFF_X2 v_in_reg_62_ ( .D(N2877), .CK(clk), .Q(v_in[62]), .QN() );
DFF_X2 v_in_reg_63_ ( .D(N2878), .CK(clk), .Q(v_in[63]), .QN() );
DFF_X2 v_in_reg_64_ ( .D(N2879), .CK(clk), .Q(v_in[64]), .QN() );
DFF_X2 v_in_reg_65_ ( .D(N2880), .CK(clk), .Q(v_in[65]), .QN() );
DFF_X2 v_in_reg_66_ ( .D(N2881), .CK(clk), .Q(v_in[66]), .QN() );
DFF_X2 v_in_reg_67_ ( .D(N2882), .CK(clk), .Q(v_in[67]), .QN() );
DFF_X2 v_in_reg_68_ ( .D(N2883), .CK(clk), .Q(v_in[68]), .QN() );
DFF_X2 v_in_reg_69_ ( .D(N2884), .CK(clk), .Q(v_in[69]), .QN() );
DFF_X2 v_in_reg_70_ ( .D(N2885), .CK(clk), .Q(v_in[70]), .QN() );
DFF_X2 v_in_reg_71_ ( .D(N2886), .CK(clk), .Q(v_in[71]), .QN() );
DFF_X2 v_in_reg_72_ ( .D(N2887), .CK(clk), .Q(v_in[72]), .QN() );
DFF_X2 v_in_reg_73_ ( .D(N2888), .CK(clk), .Q(v_in[73]), .QN() );
DFF_X2 v_in_reg_74_ ( .D(N2889), .CK(clk), .Q(v_in[74]), .QN() );
DFF_X2 v_in_reg_75_ ( .D(N2890), .CK(clk), .Q(v_in[75]), .QN() );
DFF_X2 v_in_reg_76_ ( .D(N2891), .CK(clk), .Q(v_in[76]), .QN() );
DFF_X2 v_in_reg_77_ ( .D(N2892), .CK(clk), .Q(v_in[77]), .QN() );
DFF_X2 v_in_reg_78_ ( .D(N2893), .CK(clk), .Q(v_in[78]), .QN() );
DFF_X2 v_in_reg_79_ ( .D(N2894), .CK(clk), .Q(v_in[79]), .QN() );
DFF_X2 v_in_reg_80_ ( .D(N2895), .CK(clk), .Q(v_in[80]), .QN() );
DFF_X2 v_in_reg_81_ ( .D(N2896), .CK(clk), .Q(v_in[81]), .QN() );
DFF_X2 v_in_reg_82_ ( .D(N2897), .CK(clk), .Q(v_in[82]), .QN() );
DFF_X2 v_in_reg_83_ ( .D(N2898), .CK(clk), .Q(v_in[83]), .QN() );
DFF_X2 v_in_reg_84_ ( .D(N2899), .CK(clk), .Q(v_in[84]), .QN() );
DFF_X2 v_in_reg_85_ ( .D(N2900), .CK(clk), .Q(v_in[85]), .QN() );
DFF_X2 v_in_reg_86_ ( .D(N2901), .CK(clk), .Q(v_in[86]), .QN() );
DFF_X2 v_in_reg_87_ ( .D(N2902), .CK(clk), .Q(v_in[87]), .QN() );
DFF_X2 v_in_reg_88_ ( .D(N2903), .CK(clk), .Q(v_in[88]), .QN() );
DFF_X2 v_in_reg_89_ ( .D(N2904), .CK(clk), .Q(v_in[89]), .QN() );
DFF_X2 v_in_reg_90_ ( .D(N2905), .CK(clk), .Q(v_in[90]), .QN() );
DFF_X2 v_in_reg_91_ ( .D(N2906), .CK(clk), .Q(v_in[91]), .QN() );
DFF_X2 v_in_reg_92_ ( .D(N2907), .CK(clk), .Q(v_in[92]), .QN() );
DFF_X2 v_in_reg_93_ ( .D(N2908), .CK(clk), .Q(v_in[93]), .QN() );
DFF_X2 v_in_reg_94_ ( .D(N2909), .CK(clk), .Q(v_in[94]), .QN() );
DFF_X2 v_in_reg_95_ ( .D(N2910), .CK(clk), .Q(v_in[95]), .QN() );
DFF_X2 v_in_reg_96_ ( .D(N2911), .CK(clk), .Q(v_in[96]), .QN() );
DFF_X2 v_in_reg_97_ ( .D(N2912), .CK(clk), .Q(v_in[97]), .QN() );
DFF_X2 v_in_reg_98_ ( .D(N2913), .CK(clk), .Q(v_in[98]), .QN() );
DFF_X2 v_in_reg_99_ ( .D(N2914), .CK(clk), .Q(v_in[99]), .QN() );
DFF_X2 v_in_reg_100_ ( .D(N2915), .CK(clk), .Q(v_in[100]), .QN() );
DFF_X2 v_in_reg_101_ ( .D(N2916), .CK(clk), .Q(v_in[101]), .QN() );
DFF_X2 v_in_reg_102_ ( .D(N2917), .CK(clk), .Q(v_in[102]), .QN() );
DFF_X2 v_in_reg_103_ ( .D(N2918), .CK(clk), .Q(v_in[103]), .QN() );
DFF_X2 v_in_reg_104_ ( .D(N2919), .CK(clk), .Q(v_in[104]), .QN() );
DFF_X2 v_in_reg_105_ ( .D(N2920), .CK(clk), .Q(v_in[105]), .QN() );
DFF_X2 v_in_reg_106_ ( .D(N2921), .CK(clk), .Q(v_in[106]), .QN() );
DFF_X2 v_in_reg_107_ ( .D(N2922), .CK(clk), .Q(v_in[107]), .QN() );
DFF_X2 v_in_reg_108_ ( .D(N2923), .CK(clk), .Q(v_in[108]), .QN() );
DFF_X2 v_in_reg_109_ ( .D(N2924), .CK(clk), .Q(v_in[109]), .QN() );
DFF_X2 v_in_reg_110_ ( .D(N2925), .CK(clk), .Q(v_in[110]), .QN() );
DFF_X2 v_in_reg_111_ ( .D(N2926), .CK(clk), .Q(v_in[111]), .QN() );
DFF_X2 v_in_reg_112_ ( .D(N2927), .CK(clk), .Q(v_in[112]), .QN() );
DFF_X2 v_in_reg_113_ ( .D(N2928), .CK(clk), .Q(v_in[113]), .QN() );
DFF_X2 v_in_reg_114_ ( .D(N2929), .CK(clk), .Q(v_in[114]), .QN() );
DFF_X2 v_in_reg_115_ ( .D(N2930), .CK(clk), .Q(v_in[115]), .QN() );
DFF_X2 v_in_reg_116_ ( .D(N2931), .CK(clk), .Q(v_in[116]), .QN() );
DFF_X2 v_in_reg_117_ ( .D(N2932), .CK(clk), .Q(v_in[117]), .QN() );
DFF_X2 v_in_reg_118_ ( .D(N2933), .CK(clk), .Q(v_in[118]), .QN() );
DFF_X2 v_in_reg_119_ ( .D(N2934), .CK(clk), .Q(v_in[119]), .QN() );
DFF_X2 v_in_reg_120_ ( .D(N2935), .CK(clk), .Q(v_in[120]), .QN() );
DFF_X2 v_in_reg_121_ ( .D(N2936), .CK(clk), .Q(v_in[121]), .QN() );
DFF_X2 v_in_reg_122_ ( .D(N2937), .CK(clk), .Q(v_in[122]), .QN() );
DFF_X2 v_in_reg_123_ ( .D(N2938), .CK(clk), .Q(v_in[123]), .QN() );
DFF_X2 v_in_reg_124_ ( .D(N2939), .CK(clk), .Q(v_in[124]), .QN() );
DFF_X2 v_in_reg_125_ ( .D(N2940), .CK(clk), .Q(v_in[125]), .QN() );
DFF_X2 v_in_reg_126_ ( .D(N2941), .CK(clk), .Q(v_in[126]), .QN() );
DFF_X2 v_in_reg_127_ ( .D(N2942), .CK(clk), .Q(v_in[127]), .QN() );
NAND2_X2 U6736 ( .A1(n17747), .A2(n11931), .ZN(n6292) );
NAND2_X2 U6741 ( .A1(n11935), .A2(n11936), .ZN(n6290) );
NAND2_X2 U6743 ( .A1(n11923), .A2(n18893), .ZN(n11935) );
NAND2_X2 U6744 ( .A1(n18745), .A2(n11937), .ZN(n11923) );
NAND2_X2 U6749 ( .A1(n11939), .A2(n11940), .ZN(n6289) );
NAND2_X2 U6752 ( .A1(state[6]), .A2(n11926), .ZN(n11941) );
NAND2_X2 U6753 ( .A1(n11942), .A2(n11943), .ZN(n6287) );
NAND2_X2 U6755 ( .A1(n18747), .A2(n11944), .ZN(n11926) );
NAND2_X2 U6762 ( .A1(n11953), .A2(n11954), .ZN(n11948) );
NAND2_X2 U6763 ( .A1(n11955), .A2(n18892), .ZN(n11954) );
NAND2_X2 U6767 ( .A1(n11961), .A2(n11962), .ZN(n6283) );
NAND2_X2 U6768 ( .A1(state[0]), .A2(n11963), .ZN(n11962) );
NAND2_X2 U6769 ( .A1(n17375), .A2(n11953), .ZN(n11963) );
AND3_X2 U6770 ( .A1(n11964), .A2(n11965), .A3(n11966), .ZN(n11953) );
NAND2_X2 U6773 ( .A1(cii_IV_vld), .A2(aes_done), .ZN(n11968) );
NAND2_X2 U6774 ( .A1(n11960), .A2(dii_data_not_ready), .ZN(n11964) );
AND4_X2 U6775 ( .A1(n18844), .A2(n11957), .A3(n18014), .A4(n11970), .ZN(n11960) );
NAND4_X2 U6777 ( .A1(state[5]), .A2(n11973), .A3(n18627), .A4(n18601), .ZN(n11957) );
NAND2_X2 U6782 ( .A1(n11979), .A2(n11980), .ZN(n6282) );
OR2_X2 U6783 ( .A1(n18030), .A2(n17279), .ZN(n11980) );
NAND2_X2 U6784 ( .A1(aes_text_out[0]), .A2(n18022), .ZN(n11979) );
NAND2_X2 U6785 ( .A1(n11981), .A2(n11982), .ZN(n6281) );
OR2_X2 U6786 ( .A1(n18026), .A2(n17277), .ZN(n11982) );
NAND2_X2 U6787 ( .A1(aes_text_out[1]), .A2(n18022), .ZN(n11981) );
NAND2_X2 U6788 ( .A1(n11983), .A2(n11984), .ZN(n6280) );
OR2_X2 U6789 ( .A1(n18026), .A2(n17275), .ZN(n11984) );
NAND2_X2 U6790 ( .A1(aes_text_out[2]), .A2(n18023), .ZN(n11983) );
NAND2_X2 U6791 ( .A1(n11985), .A2(n11986), .ZN(n6279) );
OR2_X2 U6792 ( .A1(n18028), .A2(n17273), .ZN(n11986) );
NAND2_X2 U6793 ( .A1(aes_text_out[3]), .A2(n18023), .ZN(n11985) );
NAND2_X2 U6794 ( .A1(n11987), .A2(n11988), .ZN(n6278) );
OR2_X2 U6795 ( .A1(n18027), .A2(n17271), .ZN(n11988) );
NAND2_X2 U6796 ( .A1(aes_text_out[4]), .A2(n18023), .ZN(n11987) );
NAND2_X2 U6797 ( .A1(n11989), .A2(n11990), .ZN(n6277) );
OR2_X2 U6798 ( .A1(n18027), .A2(n17269), .ZN(n11990) );
NAND2_X2 U6799 ( .A1(aes_text_out[5]), .A2(n18024), .ZN(n11989) );
NAND2_X2 U6800 ( .A1(n11991), .A2(n11992), .ZN(n6276) );
OR2_X2 U6801 ( .A1(n18028), .A2(n17267), .ZN(n11992) );
NAND2_X2 U6802 ( .A1(aes_text_out[6]), .A2(n18024), .ZN(n11991) );
NAND2_X2 U6803 ( .A1(n11993), .A2(n11994), .ZN(n6275) );
OR2_X2 U6804 ( .A1(n18027), .A2(n17265), .ZN(n11994) );
NAND2_X2 U6805 ( .A1(aes_text_out[7]), .A2(n18023), .ZN(n11993) );
NAND2_X2 U6806 ( .A1(n11995), .A2(n11996), .ZN(n6274) );
OR2_X2 U6807 ( .A1(n18029), .A2(n17263), .ZN(n11996) );
NAND2_X2 U6808 ( .A1(aes_text_out[8]), .A2(n18025), .ZN(n11995) );
NAND2_X2 U6809 ( .A1(n11997), .A2(n11998), .ZN(n6273) );
OR2_X2 U6810 ( .A1(n18028), .A2(n17261), .ZN(n11998) );
NAND2_X2 U6811 ( .A1(aes_text_out[9]), .A2(n18025), .ZN(n11997) );
NAND2_X2 U6812 ( .A1(n11999), .A2(n12000), .ZN(n6272) );
OR2_X2 U6813 ( .A1(n18028), .A2(n17259), .ZN(n12000) );
NAND2_X2 U6814 ( .A1(aes_text_out[10]), .A2(n18023), .ZN(n11999) );
NAND2_X2 U6815 ( .A1(n12001), .A2(n12002), .ZN(n6271) );
OR2_X2 U6816 ( .A1(n18028), .A2(n17257), .ZN(n12002) );
NAND2_X2 U6817 ( .A1(aes_text_out[11]), .A2(n18025), .ZN(n12001) );
NAND2_X2 U6818 ( .A1(n12003), .A2(n12004), .ZN(n6270) );
OR2_X2 U6819 ( .A1(n18029), .A2(n17255), .ZN(n12004) );
NAND2_X2 U6820 ( .A1(aes_text_out[12]), .A2(n18025), .ZN(n12003) );
NAND2_X2 U6821 ( .A1(n12005), .A2(n12006), .ZN(n6269) );
OR2_X2 U6822 ( .A1(n18029), .A2(n17253), .ZN(n12006) );
NAND2_X2 U6823 ( .A1(aes_text_out[13]), .A2(n18023), .ZN(n12005) );
NAND2_X2 U6824 ( .A1(n12007), .A2(n12008), .ZN(n6268) );
OR2_X2 U6825 ( .A1(n18029), .A2(n17251), .ZN(n12008) );
NAND2_X2 U6826 ( .A1(aes_text_out[14]), .A2(n18026), .ZN(n12007) );
NAND2_X2 U6827 ( .A1(n12009), .A2(n12010), .ZN(n6267) );
OR2_X2 U6828 ( .A1(n18029), .A2(n17249), .ZN(n12010) );
NAND2_X2 U6829 ( .A1(aes_text_out[15]), .A2(n18026), .ZN(n12009) );
NAND2_X2 U6830 ( .A1(n12011), .A2(n12012), .ZN(n6266) );
OR2_X2 U6831 ( .A1(n18029), .A2(n17247), .ZN(n12012) );
NAND2_X2 U6832 ( .A1(aes_text_out[16]), .A2(n18024), .ZN(n12011) );
NAND2_X2 U6833 ( .A1(n12013), .A2(n12014), .ZN(n6265) );
OR2_X2 U6834 ( .A1(n18030), .A2(n17245), .ZN(n12014) );
NAND2_X2 U6835 ( .A1(aes_text_out[17]), .A2(n18026), .ZN(n12013) );
NAND2_X2 U6836 ( .A1(n12015), .A2(n12016), .ZN(n6264) );
OR2_X2 U6837 ( .A1(n18030), .A2(n17243), .ZN(n12016) );
NAND2_X2 U6838 ( .A1(aes_text_out[18]), .A2(n18026), .ZN(n12015) );
NAND2_X2 U6839 ( .A1(n12017), .A2(n12018), .ZN(n6263) );
OR2_X2 U6840 ( .A1(n18030), .A2(n17241), .ZN(n12018) );
NAND2_X2 U6841 ( .A1(aes_text_out[19]), .A2(n18026), .ZN(n12017) );
NAND2_X2 U6842 ( .A1(n12019), .A2(n12020), .ZN(n6262) );
OR2_X2 U6843 ( .A1(n18031), .A2(n17239), .ZN(n12020) );
NAND2_X2 U6844 ( .A1(aes_text_out[20]), .A2(n18024), .ZN(n12019) );
NAND2_X2 U6845 ( .A1(n12021), .A2(n12022), .ZN(n6261) );
OR2_X2 U6846 ( .A1(n18031), .A2(n17237), .ZN(n12022) );
NAND2_X2 U6847 ( .A1(aes_text_out[21]), .A2(n18026), .ZN(n12021) );
NAND2_X2 U6848 ( .A1(n12023), .A2(n12024), .ZN(n6260) );
OR2_X2 U6849 ( .A1(n18031), .A2(n17235), .ZN(n12024) );
NAND2_X2 U6850 ( .A1(aes_text_out[22]), .A2(n18026), .ZN(n12023) );
NAND2_X2 U6851 ( .A1(n12025), .A2(n12026), .ZN(n6259) );
OR2_X2 U6852 ( .A1(n18031), .A2(n17233), .ZN(n12026) );
NAND2_X2 U6853 ( .A1(aes_text_out[23]), .A2(n18025), .ZN(n12025) );
NAND2_X2 U6854 ( .A1(n12027), .A2(n12028), .ZN(n6258) );
OR2_X2 U6855 ( .A1(n18031), .A2(n17231), .ZN(n12028) );
NAND2_X2 U6856 ( .A1(aes_text_out[24]), .A2(n18025), .ZN(n12027) );
NAND2_X2 U6857 ( .A1(n12029), .A2(n12030), .ZN(n6257) );
OR2_X2 U6858 ( .A1(n18032), .A2(n17229), .ZN(n12030) );
NAND2_X2 U6859 ( .A1(aes_text_out[25]), .A2(n18025), .ZN(n12029) );
NAND2_X2 U6860 ( .A1(n12031), .A2(n12032), .ZN(n6256) );
OR2_X2 U6861 ( .A1(n18032), .A2(n17227), .ZN(n12032) );
NAND2_X2 U6862 ( .A1(aes_text_out[26]), .A2(n18025), .ZN(n12031) );
NAND2_X2 U6863 ( .A1(n12033), .A2(n12034), .ZN(n6255) );
OR2_X2 U6864 ( .A1(n18032), .A2(n17225), .ZN(n12034) );
NAND2_X2 U6865 ( .A1(aes_text_out[27]), .A2(n18025), .ZN(n12033) );
NAND2_X2 U6866 ( .A1(n12035), .A2(n12036), .ZN(n6254) );
OR2_X2 U6867 ( .A1(n18032), .A2(n17223), .ZN(n12036) );
NAND2_X2 U6868 ( .A1(aes_text_out[28]), .A2(n18025), .ZN(n12035) );
NAND2_X2 U6869 ( .A1(n12037), .A2(n12038), .ZN(n6253) );
OR2_X2 U6870 ( .A1(n18032), .A2(n17221), .ZN(n12038) );
NAND2_X2 U6871 ( .A1(aes_text_out[29]), .A2(n18023), .ZN(n12037) );
NAND2_X2 U6872 ( .A1(n12039), .A2(n12040), .ZN(n6252) );
OR2_X2 U6873 ( .A1(n18033), .A2(n17219), .ZN(n12040) );
NAND2_X2 U6874 ( .A1(aes_text_out[30]), .A2(n18025), .ZN(n12039) );
NAND2_X2 U6875 ( .A1(n12041), .A2(n12042), .ZN(n6251) );
OR2_X2 U6876 ( .A1(n18033), .A2(n17217), .ZN(n12042) );
NAND2_X2 U6877 ( .A1(aes_text_out[31]), .A2(n18024), .ZN(n12041) );
NAND2_X2 U6878 ( .A1(n12043), .A2(n12044), .ZN(n6250) );
OR2_X2 U6879 ( .A1(n18033), .A2(n17215), .ZN(n12044) );
NAND2_X2 U6880 ( .A1(aes_text_out[32]), .A2(n18024), .ZN(n12043) );
NAND2_X2 U6881 ( .A1(n12045), .A2(n12046), .ZN(n6249) );
OR2_X2 U6882 ( .A1(n18033), .A2(n17213), .ZN(n12046) );
NAND2_X2 U6883 ( .A1(aes_text_out[33]), .A2(n18024), .ZN(n12045) );
NAND2_X2 U6884 ( .A1(n12047), .A2(n12048), .ZN(n6248) );
OR2_X2 U6885 ( .A1(n18034), .A2(n17211), .ZN(n12048) );
NAND2_X2 U6886 ( .A1(aes_text_out[34]), .A2(n18024), .ZN(n12047) );
NAND2_X2 U6887 ( .A1(n12049), .A2(n12050), .ZN(n6247) );
OR2_X2 U6888 ( .A1(n18034), .A2(n17209), .ZN(n12050) );
NAND2_X2 U6889 ( .A1(aes_text_out[35]), .A2(n18024), .ZN(n12049) );
NAND2_X2 U6890 ( .A1(n12051), .A2(n12052), .ZN(n6246) );
OR2_X2 U6891 ( .A1(n18034), .A2(n17207), .ZN(n12052) );
NAND2_X2 U6892 ( .A1(aes_text_out[36]), .A2(n18024), .ZN(n12051) );
NAND2_X2 U6893 ( .A1(n12053), .A2(n12054), .ZN(n6245) );
OR2_X2 U6894 ( .A1(n18034), .A2(n17205), .ZN(n12054) );
NAND2_X2 U6895 ( .A1(aes_text_out[37]), .A2(n18024), .ZN(n12053) );
NAND2_X2 U6896 ( .A1(n12055), .A2(n12056), .ZN(n6244) );
OR2_X2 U6897 ( .A1(n18034), .A2(n17203), .ZN(n12056) );
NAND2_X2 U6898 ( .A1(aes_text_out[38]), .A2(n18023), .ZN(n12055) );
NAND2_X2 U6899 ( .A1(n12057), .A2(n12058), .ZN(n6243) );
OR2_X2 U6900 ( .A1(n18035), .A2(n17201), .ZN(n12058) );
NAND2_X2 U6901 ( .A1(aes_text_out[39]), .A2(n18023), .ZN(n12057) );
NAND2_X2 U6902 ( .A1(n12059), .A2(n12060), .ZN(n6242) );
OR2_X2 U6903 ( .A1(n18035), .A2(n17199), .ZN(n12060) );
NAND2_X2 U6904 ( .A1(aes_text_out[40]), .A2(n18023), .ZN(n12059) );
NAND2_X2 U6905 ( .A1(n12061), .A2(n12062), .ZN(n6241) );
OR2_X2 U6906 ( .A1(n18035), .A2(n17197), .ZN(n12062) );
NAND2_X2 U6907 ( .A1(aes_text_out[41]), .A2(n18023), .ZN(n12061) );
NAND2_X2 U6908 ( .A1(n12063), .A2(n12064), .ZN(n6240) );
OR2_X2 U6909 ( .A1(n18035), .A2(n17195), .ZN(n12064) );
NAND2_X2 U6910 ( .A1(aes_text_out[42]), .A2(n18022), .ZN(n12063) );
NAND2_X2 U6911 ( .A1(n12065), .A2(n12066), .ZN(n6239) );
OR2_X2 U6912 ( .A1(n18027), .A2(n17193), .ZN(n12066) );
NAND2_X2 U6913 ( .A1(aes_text_out[43]), .A2(n18022), .ZN(n12065) );
NAND2_X2 U6914 ( .A1(n12067), .A2(n12068), .ZN(n6238) );
OR2_X2 U6915 ( .A1(n18035), .A2(n17191), .ZN(n12068) );
NAND2_X2 U6916 ( .A1(aes_text_out[44]), .A2(n18022), .ZN(n12067) );
NAND2_X2 U6917 ( .A1(n12069), .A2(n12070), .ZN(n6237) );
OR2_X2 U6918 ( .A1(n18035), .A2(n17189), .ZN(n12070) );
NAND2_X2 U6919 ( .A1(aes_text_out[45]), .A2(n18022), .ZN(n12069) );
NAND2_X2 U6920 ( .A1(n12071), .A2(n12072), .ZN(n6236) );
OR2_X2 U6921 ( .A1(n18035), .A2(n17187), .ZN(n12072) );
NAND2_X2 U6922 ( .A1(aes_text_out[46]), .A2(n18022), .ZN(n12071) );
NAND2_X2 U6923 ( .A1(n12073), .A2(n12074), .ZN(n6235) );
OR2_X2 U6924 ( .A1(n18035), .A2(n17185), .ZN(n12074) );
NAND2_X2 U6925 ( .A1(aes_text_out[47]), .A2(n18022), .ZN(n12073) );
NAND2_X2 U6926 ( .A1(n12075), .A2(n12076), .ZN(n6234) );
OR2_X2 U6927 ( .A1(n18035), .A2(n17183), .ZN(n12076) );
NAND2_X2 U6928 ( .A1(aes_text_out[48]), .A2(n18022), .ZN(n12075) );
NAND2_X2 U6929 ( .A1(n12077), .A2(n12078), .ZN(n6233) );
OR2_X2 U6930 ( .A1(n18035), .A2(n17181), .ZN(n12078) );
NAND2_X2 U6931 ( .A1(aes_text_out[49]), .A2(n18022), .ZN(n12077) );
NAND2_X2 U6932 ( .A1(n12079), .A2(n12080), .ZN(n6232) );
OR2_X2 U6933 ( .A1(n18035), .A2(n17179), .ZN(n12080) );
NAND2_X2 U6934 ( .A1(aes_text_out[50]), .A2(n18021), .ZN(n12079) );
NAND2_X2 U6935 ( .A1(n12081), .A2(n12082), .ZN(n6231) );
OR2_X2 U6936 ( .A1(n18034), .A2(n17177), .ZN(n12082) );
NAND2_X2 U6937 ( .A1(aes_text_out[51]), .A2(n18021), .ZN(n12081) );
NAND2_X2 U6938 ( .A1(n12083), .A2(n12084), .ZN(n6230) );
OR2_X2 U6939 ( .A1(n18034), .A2(n17175), .ZN(n12084) );
NAND2_X2 U6940 ( .A1(aes_text_out[52]), .A2(n18021), .ZN(n12083) );
NAND2_X2 U6941 ( .A1(n12085), .A2(n12086), .ZN(n6229) );
OR2_X2 U6942 ( .A1(n18034), .A2(n17173), .ZN(n12086) );
NAND2_X2 U6943 ( .A1(aes_text_out[53]), .A2(n18021), .ZN(n12085) );
NAND2_X2 U6944 ( .A1(n12087), .A2(n12088), .ZN(n6228) );
OR2_X2 U6945 ( .A1(n18034), .A2(n17171), .ZN(n12088) );
NAND2_X2 U6946 ( .A1(aes_text_out[54]), .A2(n18021), .ZN(n12087) );
NAND2_X2 U6947 ( .A1(n12089), .A2(n12090), .ZN(n6227) );
OR2_X2 U6948 ( .A1(n18034), .A2(n17169), .ZN(n12090) );
NAND2_X2 U6949 ( .A1(aes_text_out[55]), .A2(n18021), .ZN(n12089) );
NAND2_X2 U6950 ( .A1(n12091), .A2(n12092), .ZN(n6226) );
OR2_X2 U6951 ( .A1(n18034), .A2(n17167), .ZN(n12092) );
NAND2_X2 U6952 ( .A1(aes_text_out[56]), .A2(n18021), .ZN(n12091) );
NAND2_X2 U6953 ( .A1(n12093), .A2(n12094), .ZN(n6225) );
OR2_X2 U6954 ( .A1(n18034), .A2(n17165), .ZN(n12094) );
NAND2_X2 U6955 ( .A1(aes_text_out[57]), .A2(n18021), .ZN(n12093) );
NAND2_X2 U6956 ( .A1(n12095), .A2(n12096), .ZN(n6224) );
OR2_X2 U6957 ( .A1(n18034), .A2(n17163), .ZN(n12096) );
NAND2_X2 U6958 ( .A1(aes_text_out[58]), .A2(n18021), .ZN(n12095) );
NAND2_X2 U6959 ( .A1(n12097), .A2(n12098), .ZN(n6223) );
OR2_X2 U6960 ( .A1(n18034), .A2(n17161), .ZN(n12098) );
NAND2_X2 U6961 ( .A1(aes_text_out[59]), .A2(n18021), .ZN(n12097) );
NAND2_X2 U6962 ( .A1(n12099), .A2(n12100), .ZN(n6222) );
OR2_X2 U6963 ( .A1(n18033), .A2(n17159), .ZN(n12100) );
NAND2_X2 U6964 ( .A1(aes_text_out[60]), .A2(n18021), .ZN(n12099) );
NAND2_X2 U6965 ( .A1(n12101), .A2(n12102), .ZN(n6221) );
OR2_X2 U6966 ( .A1(n18033), .A2(n17157), .ZN(n12102) );
NAND2_X2 U6967 ( .A1(aes_text_out[61]), .A2(n18020), .ZN(n12101) );
NAND2_X2 U6968 ( .A1(n12103), .A2(n12104), .ZN(n6220) );
OR2_X2 U6969 ( .A1(n18033), .A2(n17155), .ZN(n12104) );
NAND2_X2 U6970 ( .A1(aes_text_out[62]), .A2(n18020), .ZN(n12103) );
NAND2_X2 U6971 ( .A1(n12105), .A2(n12106), .ZN(n6219) );
OR2_X2 U6972 ( .A1(n18033), .A2(n17153), .ZN(n12106) );
NAND2_X2 U6973 ( .A1(aes_text_out[63]), .A2(n18022), .ZN(n12105) );
NAND2_X2 U6974 ( .A1(n12107), .A2(n12108), .ZN(n6218) );
OR2_X2 U6975 ( .A1(n18033), .A2(n17151), .ZN(n12108) );
NAND2_X2 U6976 ( .A1(aes_text_out[64]), .A2(n18020), .ZN(n12107) );
NAND2_X2 U6977 ( .A1(n12109), .A2(n12110), .ZN(n6217) );
OR2_X2 U6978 ( .A1(n18033), .A2(n17149), .ZN(n12110) );
NAND2_X2 U6979 ( .A1(aes_text_out[65]), .A2(n18020), .ZN(n12109) );
NAND2_X2 U6980 ( .A1(n12111), .A2(n12112), .ZN(n6216) );
OR2_X2 U6981 ( .A1(n18033), .A2(n17147), .ZN(n12112) );
NAND2_X2 U6982 ( .A1(aes_text_out[66]), .A2(n18020), .ZN(n12111) );
NAND2_X2 U6983 ( .A1(n12113), .A2(n12114), .ZN(n6215) );
OR2_X2 U6984 ( .A1(n18033), .A2(n17145), .ZN(n12114) );
NAND2_X2 U6985 ( .A1(aes_text_out[67]), .A2(n18020), .ZN(n12113) );
NAND2_X2 U6986 ( .A1(n12115), .A2(n12116), .ZN(n6214) );
OR2_X2 U6987 ( .A1(n18033), .A2(n17143), .ZN(n12116) );
NAND2_X2 U6988 ( .A1(aes_text_out[68]), .A2(n18020), .ZN(n12115) );
NAND2_X2 U6989 ( .A1(n12117), .A2(n12118), .ZN(n6213) );
OR2_X2 U6990 ( .A1(n18033), .A2(n17141), .ZN(n12118) );
NAND2_X2 U6991 ( .A1(aes_text_out[69]), .A2(n18020), .ZN(n12117) );
NAND2_X2 U6992 ( .A1(n12119), .A2(n12120), .ZN(n6212) );
OR2_X2 U6993 ( .A1(n18032), .A2(n17139), .ZN(n12120) );
NAND2_X2 U6994 ( .A1(aes_text_out[70]), .A2(n18020), .ZN(n12119) );
NAND2_X2 U6995 ( .A1(n12121), .A2(n12122), .ZN(n6211) );
OR2_X2 U6996 ( .A1(n18032), .A2(n17137), .ZN(n12122) );
NAND2_X2 U6997 ( .A1(aes_text_out[71]), .A2(n18020), .ZN(n12121) );
NAND2_X2 U6998 ( .A1(n12123), .A2(n12124), .ZN(n6210) );
OR2_X2 U6999 ( .A1(n18032), .A2(n17135), .ZN(n12124) );
NAND2_X2 U7000 ( .A1(aes_text_out[72]), .A2(n18019), .ZN(n12123) );
NAND2_X2 U7001 ( .A1(n12125), .A2(n12126), .ZN(n6209) );
OR2_X2 U7002 ( .A1(n18032), .A2(n17133), .ZN(n12126) );
NAND2_X2 U7003 ( .A1(aes_text_out[73]), .A2(n18019), .ZN(n12125) );
NAND2_X2 U7004 ( .A1(n12127), .A2(n12128), .ZN(n6208) );
OR2_X2 U7005 ( .A1(n18032), .A2(n17131), .ZN(n12128) );
NAND2_X2 U7006 ( .A1(aes_text_out[74]), .A2(n18019), .ZN(n12127) );
NAND2_X2 U7007 ( .A1(n12129), .A2(n12130), .ZN(n6207) );
OR2_X2 U7008 ( .A1(n18032), .A2(n17129), .ZN(n12130) );
NAND2_X2 U7009 ( .A1(aes_text_out[75]), .A2(n18019), .ZN(n12129) );
NAND2_X2 U7010 ( .A1(n12131), .A2(n12132), .ZN(n6206) );
OR2_X2 U7011 ( .A1(n18032), .A2(n17127), .ZN(n12132) );
NAND2_X2 U7012 ( .A1(aes_text_out[76]), .A2(n18019), .ZN(n12131) );
NAND2_X2 U7013 ( .A1(n12133), .A2(n12134), .ZN(n6205) );
OR2_X2 U7014 ( .A1(n18032), .A2(n17125), .ZN(n12134) );
NAND2_X2 U7015 ( .A1(aes_text_out[77]), .A2(n18019), .ZN(n12133) );
NAND2_X2 U7016 ( .A1(n12135), .A2(n12136), .ZN(n6204) );
OR2_X2 U7017 ( .A1(n18032), .A2(n17123), .ZN(n12136) );
NAND2_X2 U7018 ( .A1(aes_text_out[78]), .A2(n18019), .ZN(n12135) );
NAND2_X2 U7019 ( .A1(n12137), .A2(n12138), .ZN(n6203) );
OR2_X2 U7020 ( .A1(n18031), .A2(n17121), .ZN(n12138) );
NAND2_X2 U7021 ( .A1(aes_text_out[79]), .A2(n18019), .ZN(n12137) );
NAND2_X2 U7022 ( .A1(n12139), .A2(n12140), .ZN(n6202) );
OR2_X2 U7023 ( .A1(n18031), .A2(n17119), .ZN(n12140) );
NAND2_X2 U7024 ( .A1(aes_text_out[80]), .A2(n18019), .ZN(n12139) );
NAND2_X2 U7025 ( .A1(n12141), .A2(n12142), .ZN(n6201) );
OR2_X2 U7026 ( .A1(n18031), .A2(n17117), .ZN(n12142) );
NAND2_X2 U7027 ( .A1(aes_text_out[81]), .A2(n18019), .ZN(n12141) );
NAND2_X2 U7028 ( .A1(n12143), .A2(n12144), .ZN(n6200) );
OR2_X2 U7029 ( .A1(n18031), .A2(n17115), .ZN(n12144) );
NAND2_X2 U7030 ( .A1(aes_text_out[82]), .A2(n18019), .ZN(n12143) );
NAND2_X2 U7031 ( .A1(n12145), .A2(n12146), .ZN(n6199) );
OR2_X2 U7032 ( .A1(n18031), .A2(n17113), .ZN(n12146) );
NAND2_X2 U7033 ( .A1(aes_text_out[83]), .A2(n18018), .ZN(n12145) );
NAND2_X2 U7034 ( .A1(n12147), .A2(n12148), .ZN(n6198) );
OR2_X2 U7035 ( .A1(n18031), .A2(n17111), .ZN(n12148) );
NAND2_X2 U7036 ( .A1(aes_text_out[84]), .A2(n18018), .ZN(n12147) );
NAND2_X2 U7037 ( .A1(n12149), .A2(n12150), .ZN(n6197) );
OR2_X2 U7038 ( .A1(n18031), .A2(n17109), .ZN(n12150) );
NAND2_X2 U7039 ( .A1(aes_text_out[85]), .A2(n18018), .ZN(n12149) );
NAND2_X2 U7040 ( .A1(n12151), .A2(n12152), .ZN(n6196) );
OR2_X2 U7041 ( .A1(n18031), .A2(n17107), .ZN(n12152) );
NAND2_X2 U7042 ( .A1(aes_text_out[86]), .A2(n18018), .ZN(n12151) );
NAND2_X2 U7043 ( .A1(n12153), .A2(n12154), .ZN(n6195) );
OR2_X2 U7044 ( .A1(n18031), .A2(n17105), .ZN(n12154) );
NAND2_X2 U7045 ( .A1(aes_text_out[87]), .A2(n18018), .ZN(n12153) );
NAND2_X2 U7046 ( .A1(n12155), .A2(n12156), .ZN(n6194) );
OR2_X2 U7047 ( .A1(n18030), .A2(n17103), .ZN(n12156) );
NAND2_X2 U7048 ( .A1(aes_text_out[88]), .A2(n18018), .ZN(n12155) );
NAND2_X2 U7049 ( .A1(n12157), .A2(n12158), .ZN(n6193) );
OR2_X2 U7050 ( .A1(n18030), .A2(n17101), .ZN(n12158) );
NAND2_X2 U7051 ( .A1(aes_text_out[89]), .A2(n18018), .ZN(n12157) );
NAND2_X2 U7052 ( .A1(n12159), .A2(n12160), .ZN(n6192) );
OR2_X2 U7053 ( .A1(n18030), .A2(n17099), .ZN(n12160) );
NAND2_X2 U7054 ( .A1(aes_text_out[90]), .A2(n18018), .ZN(n12159) );
NAND2_X2 U7055 ( .A1(n12161), .A2(n12162), .ZN(n6191) );
OR2_X2 U7056 ( .A1(n18030), .A2(n17097), .ZN(n12162) );
NAND2_X2 U7057 ( .A1(aes_text_out[91]), .A2(n18018), .ZN(n12161) );
NAND2_X2 U7058 ( .A1(n12163), .A2(n12164), .ZN(n6190) );
OR2_X2 U7059 ( .A1(n18030), .A2(n17095), .ZN(n12164) );
NAND2_X2 U7060 ( .A1(aes_text_out[92]), .A2(n18018), .ZN(n12163) );
NAND2_X2 U7061 ( .A1(n12165), .A2(n12166), .ZN(n6189) );
OR2_X2 U7062 ( .A1(n18030), .A2(n17093), .ZN(n12166) );
NAND2_X2 U7063 ( .A1(aes_text_out[93]), .A2(n18018), .ZN(n12165) );
NAND2_X2 U7064 ( .A1(n12167), .A2(n12168), .ZN(n6188) );
OR2_X2 U7065 ( .A1(n18030), .A2(n17091), .ZN(n12168) );
NAND2_X2 U7066 ( .A1(aes_text_out[94]), .A2(n18017), .ZN(n12167) );
NAND2_X2 U7067 ( .A1(n12169), .A2(n12170), .ZN(n6187) );
OR2_X2 U7068 ( .A1(n18030), .A2(n17089), .ZN(n12170) );
NAND2_X2 U7069 ( .A1(aes_text_out[95]), .A2(n18017), .ZN(n12169) );
NAND2_X2 U7070 ( .A1(n12171), .A2(n12172), .ZN(n6186) );
OR2_X2 U7071 ( .A1(n18030), .A2(n17087), .ZN(n12172) );
NAND2_X2 U7072 ( .A1(aes_text_out[96]), .A2(n18017), .ZN(n12171) );
NAND2_X2 U7073 ( .A1(n12173), .A2(n12174), .ZN(n6185) );
OR2_X2 U7074 ( .A1(n18029), .A2(n17085), .ZN(n12174) );
NAND2_X2 U7075 ( .A1(aes_text_out[97]), .A2(n18017), .ZN(n12173) );
NAND2_X2 U7076 ( .A1(n12175), .A2(n12176), .ZN(n6184) );
OR2_X2 U7077 ( .A1(n18030), .A2(n17083), .ZN(n12176) );
NAND2_X2 U7078 ( .A1(aes_text_out[98]), .A2(n18017), .ZN(n12175) );
NAND2_X2 U7079 ( .A1(n12177), .A2(n12178), .ZN(n6183) );
OR2_X2 U7080 ( .A1(n18029), .A2(n17081), .ZN(n12178) );
NAND2_X2 U7081 ( .A1(aes_text_out[99]), .A2(n18017), .ZN(n12177) );
NAND2_X2 U7082 ( .A1(n12179), .A2(n12180), .ZN(n6182) );
OR2_X2 U7083 ( .A1(n18029), .A2(n17079), .ZN(n12180) );
NAND2_X2 U7084 ( .A1(aes_text_out[100]), .A2(n18017), .ZN(n12179) );
NAND2_X2 U7085 ( .A1(n12181), .A2(n12182), .ZN(n6181) );
OR2_X2 U7086 ( .A1(n18029), .A2(n17077), .ZN(n12182) );
NAND2_X2 U7087 ( .A1(aes_text_out[101]), .A2(n18017), .ZN(n12181) );
NAND2_X2 U7088 ( .A1(n12183), .A2(n12184), .ZN(n6180) );
OR2_X2 U7089 ( .A1(n18029), .A2(n17075), .ZN(n12184) );
NAND2_X2 U7090 ( .A1(aes_text_out[102]), .A2(n18017), .ZN(n12183) );
NAND2_X2 U7091 ( .A1(n12185), .A2(n12186), .ZN(n6179) );
OR2_X2 U7092 ( .A1(n18029), .A2(n17073), .ZN(n12186) );
NAND2_X2 U7093 ( .A1(aes_text_out[103]), .A2(n18017), .ZN(n12185) );
NAND2_X2 U7094 ( .A1(n12187), .A2(n12188), .ZN(n6178) );
OR2_X2 U7095 ( .A1(n18028), .A2(n17071), .ZN(n12188) );
NAND2_X2 U7096 ( .A1(aes_text_out[104]), .A2(n18017), .ZN(n12187) );
NAND2_X2 U7097 ( .A1(n12189), .A2(n12190), .ZN(n6177) );
OR2_X2 U7098 ( .A1(n18029), .A2(n17069), .ZN(n12190) );
NAND2_X2 U7099 ( .A1(aes_text_out[105]), .A2(n18016), .ZN(n12189) );
NAND2_X2 U7100 ( .A1(n12191), .A2(n12192), .ZN(n6176) );
OR2_X2 U7101 ( .A1(n18028), .A2(n17067), .ZN(n12192) );
NAND2_X2 U7102 ( .A1(aes_text_out[106]), .A2(n18016), .ZN(n12191) );
NAND2_X2 U7103 ( .A1(n12193), .A2(n12194), .ZN(n6175) );
OR2_X2 U7104 ( .A1(n18028), .A2(n17065), .ZN(n12194) );
NAND2_X2 U7105 ( .A1(aes_text_out[107]), .A2(n18016), .ZN(n12193) );
NAND2_X2 U7106 ( .A1(n12195), .A2(n12196), .ZN(n6174) );
OR2_X2 U7107 ( .A1(n18028), .A2(n17063), .ZN(n12196) );
NAND2_X2 U7108 ( .A1(aes_text_out[108]), .A2(n18016), .ZN(n12195) );
NAND2_X2 U7109 ( .A1(n12197), .A2(n12198), .ZN(n6173) );
OR2_X2 U7110 ( .A1(n18028), .A2(n17061), .ZN(n12198) );
NAND2_X2 U7111 ( .A1(aes_text_out[109]), .A2(n18016), .ZN(n12197) );
NAND2_X2 U7112 ( .A1(n12199), .A2(n12200), .ZN(n6172) );
OR2_X2 U7113 ( .A1(n18028), .A2(n17059), .ZN(n12200) );
NAND2_X2 U7114 ( .A1(aes_text_out[110]), .A2(n18016), .ZN(n12199) );
NAND2_X2 U7115 ( .A1(n12201), .A2(n12202), .ZN(n6171) );
OR2_X2 U7116 ( .A1(n18028), .A2(n17057), .ZN(n12202) );
NAND2_X2 U7117 ( .A1(aes_text_out[111]), .A2(n18016), .ZN(n12201) );
NAND2_X2 U7118 ( .A1(n12203), .A2(n12204), .ZN(n6170) );
OR2_X2 U7119 ( .A1(n18027), .A2(n17055), .ZN(n12204) );
NAND2_X2 U7120 ( .A1(aes_text_out[112]), .A2(n18016), .ZN(n12203) );
NAND2_X2 U7121 ( .A1(n12205), .A2(n12206), .ZN(n6169) );
OR2_X2 U7122 ( .A1(n18027), .A2(n17053), .ZN(n12206) );
NAND2_X2 U7123 ( .A1(aes_text_out[113]), .A2(n18016), .ZN(n12205) );
NAND2_X2 U7124 ( .A1(n12207), .A2(n12208), .ZN(n6168) );
OR2_X2 U7125 ( .A1(n18029), .A2(n17051), .ZN(n12208) );
NAND2_X2 U7126 ( .A1(aes_text_out[114]), .A2(n18016), .ZN(n12207) );
NAND2_X2 U7127 ( .A1(n12209), .A2(n12210), .ZN(n6167) );
OR2_X2 U7128 ( .A1(n18028), .A2(n17049), .ZN(n12210) );
NAND2_X2 U7129 ( .A1(aes_text_out[115]), .A2(n18016), .ZN(n12209) );
NAND2_X2 U7130 ( .A1(n12211), .A2(n12212), .ZN(n6166) );
OR2_X2 U7131 ( .A1(n18027), .A2(n17047), .ZN(n12212) );
NAND2_X2 U7132 ( .A1(aes_text_out[116]), .A2(n18015), .ZN(n12211) );
NAND2_X2 U7133 ( .A1(n12213), .A2(n12214), .ZN(n6165) );
OR2_X2 U7134 ( .A1(n18027), .A2(n17045), .ZN(n12214) );
NAND2_X2 U7135 ( .A1(aes_text_out[117]), .A2(n18015), .ZN(n12213) );
NAND2_X2 U7136 ( .A1(n12215), .A2(n12216), .ZN(n6164) );
OR2_X2 U7137 ( .A1(n18027), .A2(n17043), .ZN(n12216) );
NAND2_X2 U7138 ( .A1(aes_text_out[118]), .A2(n18015), .ZN(n12215) );
NAND2_X2 U7139 ( .A1(n12217), .A2(n12218), .ZN(n6163) );
OR2_X2 U7140 ( .A1(n18027), .A2(n17041), .ZN(n12218) );
NAND2_X2 U7141 ( .A1(aes_text_out[119]), .A2(n18015), .ZN(n12217) );
NAND2_X2 U7142 ( .A1(n12219), .A2(n12220), .ZN(n6162) );
OR2_X2 U7143 ( .A1(n18027), .A2(n17039), .ZN(n12220) );
NAND2_X2 U7144 ( .A1(aes_text_out[120]), .A2(n18015), .ZN(n12219) );
NAND2_X2 U7145 ( .A1(n12221), .A2(n12222), .ZN(n6161) );
OR2_X2 U7146 ( .A1(n18027), .A2(n17037), .ZN(n12222) );
NAND2_X2 U7147 ( .A1(aes_text_out[121]), .A2(n18015), .ZN(n12221) );
NAND2_X2 U7148 ( .A1(n12223), .A2(n12224), .ZN(n6160) );
OR2_X2 U7149 ( .A1(n18026), .A2(n17035), .ZN(n12224) );
NAND2_X2 U7150 ( .A1(aes_text_out[122]), .A2(n18015), .ZN(n12223) );
NAND2_X2 U7151 ( .A1(n12225), .A2(n12226), .ZN(n6159) );
OR2_X2 U7152 ( .A1(n18027), .A2(n17033), .ZN(n12226) );
NAND2_X2 U7153 ( .A1(aes_text_out[123]), .A2(n18015), .ZN(n12225) );
NAND2_X2 U7154 ( .A1(n12227), .A2(n12228), .ZN(n6158) );
OR2_X2 U7155 ( .A1(n18026), .A2(n17031), .ZN(n12228) );
NAND2_X2 U7156 ( .A1(aes_text_out[124]), .A2(n18015), .ZN(n12227) );
NAND2_X2 U7157 ( .A1(n12229), .A2(n12230), .ZN(n6157) );
OR2_X2 U7158 ( .A1(n18028), .A2(n17029), .ZN(n12230) );
NAND2_X2 U7159 ( .A1(aes_text_out[125]), .A2(n18015), .ZN(n12229) );
NAND2_X2 U7160 ( .A1(n12231), .A2(n12232), .ZN(n6156) );
OR2_X2 U7161 ( .A1(n18027), .A2(n17027), .ZN(n12232) );
NAND2_X2 U7162 ( .A1(aes_text_out[126]), .A2(n18015), .ZN(n12231) );
NAND2_X2 U7163 ( .A1(n12233), .A2(n12234), .ZN(n6155) );
OR2_X2 U7164 ( .A1(n18026), .A2(n17025), .ZN(n12234) );
NAND2_X2 U7165 ( .A1(aes_text_out[127]), .A2(n18020), .ZN(n12233) );
NAND2_X2 U7168 ( .A1(n12236), .A2(n12237), .ZN(n6154) );
NAND2_X2 U7169 ( .A1(aes_text_out[0]), .A2(n17989), .ZN(n12237) );
NAND2_X2 U7170 ( .A1(n17988), .A2(n18891), .ZN(n12236) );
NAND2_X2 U7171 ( .A1(n12239), .A2(n12240), .ZN(n6153) );
NAND2_X2 U7172 ( .A1(aes_text_out[1]), .A2(n17989), .ZN(n12240) );
NAND2_X2 U7173 ( .A1(n17988), .A2(n18890), .ZN(n12239) );
NAND2_X2 U7174 ( .A1(n12241), .A2(n12242), .ZN(n6152) );
NAND2_X2 U7175 ( .A1(aes_text_out[2]), .A2(n17989), .ZN(n12242) );
NAND2_X2 U7176 ( .A1(n17988), .A2(n18889), .ZN(n12241) );
NAND2_X2 U7177 ( .A1(n12243), .A2(n12244), .ZN(n6151) );
NAND2_X2 U7178 ( .A1(aes_text_out[3]), .A2(n17995), .ZN(n12244) );
NAND2_X2 U7179 ( .A1(n17988), .A2(n18888), .ZN(n12243) );
NAND2_X2 U7180 ( .A1(n12245), .A2(n12246), .ZN(n6150) );
NAND2_X2 U7181 ( .A1(aes_text_out[4]), .A2(n17995), .ZN(n12246) );
NAND2_X2 U7182 ( .A1(n17988), .A2(n18887), .ZN(n12245) );
NAND2_X2 U7183 ( .A1(n12247), .A2(n12248), .ZN(n6149) );
NAND2_X2 U7184 ( .A1(aes_text_out[5]), .A2(n17995), .ZN(n12248) );
NAND2_X2 U7185 ( .A1(n17988), .A2(n18886), .ZN(n12247) );
NAND2_X2 U7186 ( .A1(n12249), .A2(n12250), .ZN(n6148) );
NAND2_X2 U7187 ( .A1(aes_text_out[6]), .A2(n17995), .ZN(n12250) );
NAND2_X2 U7188 ( .A1(n17988), .A2(n18885), .ZN(n12249) );
NAND2_X2 U7189 ( .A1(n12251), .A2(n12252), .ZN(n6147) );
NAND2_X2 U7190 ( .A1(aes_text_out[7]), .A2(n17995), .ZN(n12252) );
NAND2_X2 U7191 ( .A1(n17987), .A2(n18884), .ZN(n12251) );
NAND2_X2 U7192 ( .A1(n12253), .A2(n12254), .ZN(n6146) );
NAND2_X2 U7193 ( .A1(aes_text_out[8]), .A2(n17995), .ZN(n12254) );
NAND2_X2 U7194 ( .A1(n17987), .A2(n18883), .ZN(n12253) );
NAND2_X2 U7195 ( .A1(n12255), .A2(n12256), .ZN(n6145) );
NAND2_X2 U7196 ( .A1(aes_text_out[9]), .A2(n17995), .ZN(n12256) );
NAND2_X2 U7197 ( .A1(n17987), .A2(n18882), .ZN(n12255) );
NAND2_X2 U7198 ( .A1(n12257), .A2(n12258), .ZN(n6144) );
NAND2_X2 U7199 ( .A1(aes_text_out[10]), .A2(n17995), .ZN(n12258) );
NAND2_X2 U7200 ( .A1(n17987), .A2(n18881), .ZN(n12257) );
NAND2_X2 U7201 ( .A1(n12259), .A2(n12260), .ZN(n6143) );
NAND2_X2 U7202 ( .A1(aes_text_out[11]), .A2(n17995), .ZN(n12260) );
NAND2_X2 U7203 ( .A1(n17987), .A2(n18880), .ZN(n12259) );
NAND2_X2 U7204 ( .A1(n12261), .A2(n12262), .ZN(n6142) );
NAND2_X2 U7205 ( .A1(aes_text_out[12]), .A2(n17995), .ZN(n12262) );
NAND2_X2 U7206 ( .A1(n17987), .A2(n18879), .ZN(n12261) );
NAND2_X2 U7207 ( .A1(n12263), .A2(n12264), .ZN(n6141) );
NAND2_X2 U7208 ( .A1(aes_text_out[13]), .A2(n17995), .ZN(n12264) );
NAND2_X2 U7209 ( .A1(n17987), .A2(n18878), .ZN(n12263) );
NAND2_X2 U7210 ( .A1(n12265), .A2(n12266), .ZN(n6140) );
NAND2_X2 U7211 ( .A1(aes_text_out[14]), .A2(n17995), .ZN(n12266) );
NAND2_X2 U7212 ( .A1(n17987), .A2(n18877), .ZN(n12265) );
NAND2_X2 U7213 ( .A1(n12267), .A2(n12268), .ZN(n6139) );
NAND2_X2 U7214 ( .A1(aes_text_out[15]), .A2(n17995), .ZN(n12268) );
NAND2_X2 U7215 ( .A1(n17987), .A2(n18876), .ZN(n12267) );
NAND2_X2 U7216 ( .A1(n12269), .A2(n12270), .ZN(n6138) );
NAND2_X2 U7217 ( .A1(aes_text_out[16]), .A2(n17995), .ZN(n12270) );
NAND2_X2 U7218 ( .A1(n17987), .A2(n18875), .ZN(n12269) );
NAND2_X2 U7219 ( .A1(n12271), .A2(n12272), .ZN(n6137) );
NAND2_X2 U7220 ( .A1(aes_text_out[17]), .A2(n17995), .ZN(n12272) );
NAND2_X2 U7221 ( .A1(n17987), .A2(n18874), .ZN(n12271) );
NAND2_X2 U7222 ( .A1(n12273), .A2(n12274), .ZN(n6136) );
NAND2_X2 U7223 ( .A1(aes_text_out[18]), .A2(n17995), .ZN(n12274) );
NAND2_X2 U7224 ( .A1(n17986), .A2(n18873), .ZN(n12273) );
NAND2_X2 U7225 ( .A1(n12275), .A2(n12276), .ZN(n6135) );
NAND2_X2 U7226 ( .A1(aes_text_out[19]), .A2(n17995), .ZN(n12276) );
NAND2_X2 U7227 ( .A1(n17986), .A2(n18872), .ZN(n12275) );
NAND2_X2 U7228 ( .A1(n12277), .A2(n12278), .ZN(n6134) );
NAND2_X2 U7229 ( .A1(aes_text_out[20]), .A2(n17995), .ZN(n12278) );
NAND2_X2 U7230 ( .A1(n17986), .A2(n18871), .ZN(n12277) );
NAND2_X2 U7231 ( .A1(n12279), .A2(n12280), .ZN(n6133) );
NAND2_X2 U7232 ( .A1(aes_text_out[21]), .A2(n17995), .ZN(n12280) );
NAND2_X2 U7233 ( .A1(n17986), .A2(n18870), .ZN(n12279) );
NAND2_X2 U7234 ( .A1(n12281), .A2(n12282), .ZN(n6132) );
NAND2_X2 U7235 ( .A1(aes_text_out[22]), .A2(n17995), .ZN(n12282) );
NAND2_X2 U7236 ( .A1(n17986), .A2(n18869), .ZN(n12281) );
NAND2_X2 U7237 ( .A1(n12283), .A2(n12284), .ZN(n6131) );
NAND2_X2 U7238 ( .A1(aes_text_out[23]), .A2(n17995), .ZN(n12284) );
NAND2_X2 U7239 ( .A1(n17986), .A2(n18868), .ZN(n12283) );
NAND2_X2 U7240 ( .A1(n12285), .A2(n12286), .ZN(n6130) );
NAND2_X2 U7241 ( .A1(aes_text_out[24]), .A2(n17994), .ZN(n12286) );
NAND2_X2 U7242 ( .A1(n17986), .A2(n18867), .ZN(n12285) );
NAND2_X2 U7243 ( .A1(n12287), .A2(n12288), .ZN(n6129) );
NAND2_X2 U7244 ( .A1(aes_text_out[25]), .A2(n17994), .ZN(n12288) );
NAND2_X2 U7245 ( .A1(n17986), .A2(n18866), .ZN(n12287) );
NAND2_X2 U7246 ( .A1(n12289), .A2(n12290), .ZN(n6128) );
NAND2_X2 U7247 ( .A1(aes_text_out[26]), .A2(n17994), .ZN(n12290) );
NAND2_X2 U7248 ( .A1(n17986), .A2(n18865), .ZN(n12289) );
NAND2_X2 U7249 ( .A1(n12291), .A2(n12292), .ZN(n6127) );
NAND2_X2 U7250 ( .A1(aes_text_out[27]), .A2(n17994), .ZN(n12292) );
NAND2_X2 U7251 ( .A1(n17986), .A2(n18864), .ZN(n12291) );
NAND2_X2 U7252 ( .A1(n12293), .A2(n12294), .ZN(n6126) );
NAND2_X2 U7253 ( .A1(aes_text_out[28]), .A2(n17994), .ZN(n12294) );
NAND2_X2 U7254 ( .A1(n17986), .A2(n18863), .ZN(n12293) );
NAND2_X2 U7255 ( .A1(n12295), .A2(n12296), .ZN(n6125) );
NAND2_X2 U7256 ( .A1(aes_text_out[29]), .A2(n17994), .ZN(n12296) );
NAND2_X2 U7257 ( .A1(n17985), .A2(n18862), .ZN(n12295) );
NAND2_X2 U7258 ( .A1(n12297), .A2(n12298), .ZN(n6124) );
NAND2_X2 U7259 ( .A1(aes_text_out[30]), .A2(n17994), .ZN(n12298) );
NAND2_X2 U7260 ( .A1(n17985), .A2(n18861), .ZN(n12297) );
NAND2_X2 U7261 ( .A1(n12299), .A2(n12300), .ZN(n6123) );
NAND2_X2 U7262 ( .A1(aes_text_out[31]), .A2(n17994), .ZN(n12300) );
NAND2_X2 U7263 ( .A1(n17985), .A2(n18860), .ZN(n12299) );
NAND2_X2 U7264 ( .A1(n12301), .A2(n12302), .ZN(n6122) );
NAND2_X2 U7265 ( .A1(aes_text_out[32]), .A2(n17994), .ZN(n12302) );
NAND2_X2 U7266 ( .A1(n17985), .A2(n18859), .ZN(n12301) );
NAND2_X2 U7267 ( .A1(n12303), .A2(n12304), .ZN(n6121) );
NAND2_X2 U7268 ( .A1(aes_text_out[33]), .A2(n17994), .ZN(n12304) );
NAND2_X2 U7269 ( .A1(n17985), .A2(n18858), .ZN(n12303) );
NAND2_X2 U7270 ( .A1(n12305), .A2(n12306), .ZN(n6120) );
NAND2_X2 U7271 ( .A1(aes_text_out[34]), .A2(n17994), .ZN(n12306) );
NAND2_X2 U7272 ( .A1(n17985), .A2(n18857), .ZN(n12305) );
NAND2_X2 U7273 ( .A1(n12307), .A2(n12308), .ZN(n6119) );
NAND2_X2 U7274 ( .A1(aes_text_out[35]), .A2(n17994), .ZN(n12308) );
NAND2_X2 U7275 ( .A1(n17985), .A2(n18856), .ZN(n12307) );
NAND2_X2 U7276 ( .A1(n12309), .A2(n12310), .ZN(n6118) );
NAND2_X2 U7277 ( .A1(aes_text_out[36]), .A2(n17994), .ZN(n12310) );
NAND2_X2 U7278 ( .A1(n17985), .A2(n18855), .ZN(n12309) );
NAND2_X2 U7279 ( .A1(n12311), .A2(n12312), .ZN(n6117) );
NAND2_X2 U7280 ( .A1(aes_text_out[37]), .A2(n17994), .ZN(n12312) );
NAND2_X2 U7281 ( .A1(n17985), .A2(n18854), .ZN(n12311) );
NAND2_X2 U7282 ( .A1(n12313), .A2(n12314), .ZN(n6116) );
NAND2_X2 U7283 ( .A1(aes_text_out[38]), .A2(n17994), .ZN(n12314) );
NAND2_X2 U7284 ( .A1(n17985), .A2(n18853), .ZN(n12313) );
NAND2_X2 U7285 ( .A1(n12315), .A2(n12316), .ZN(n6115) );
NAND2_X2 U7286 ( .A1(aes_text_out[39]), .A2(n17994), .ZN(n12316) );
NAND2_X2 U7287 ( .A1(n17985), .A2(n18852), .ZN(n12315) );
NAND2_X2 U7288 ( .A1(n12317), .A2(n12318), .ZN(n6114) );
NAND2_X2 U7289 ( .A1(aes_text_out[40]), .A2(n17994), .ZN(n12318) );
NAND2_X2 U7290 ( .A1(n17984), .A2(n18851), .ZN(n12317) );
NAND2_X2 U7291 ( .A1(n12319), .A2(n12320), .ZN(n6113) );
NAND2_X2 U7292 ( .A1(aes_text_out[41]), .A2(n17994), .ZN(n12320) );
NAND2_X2 U7293 ( .A1(n17984), .A2(n18850), .ZN(n12319) );
NAND2_X2 U7294 ( .A1(n12321), .A2(n12322), .ZN(n6112) );
NAND2_X2 U7295 ( .A1(aes_text_out[42]), .A2(n17994), .ZN(n12322) );
NAND2_X2 U7296 ( .A1(n17984), .A2(n18849), .ZN(n12321) );
NAND2_X2 U7297 ( .A1(n12323), .A2(n12324), .ZN(n6111) );
NAND2_X2 U7298 ( .A1(aes_text_out[43]), .A2(n17994), .ZN(n12324) );
NAND2_X2 U7299 ( .A1(n17984), .A2(n18848), .ZN(n12323) );
NAND2_X2 U7300 ( .A1(n12325), .A2(n12326), .ZN(n6110) );
NAND2_X2 U7301 ( .A1(aes_text_out[44]), .A2(n17994), .ZN(n12326) );
NAND2_X2 U7302 ( .A1(n17984), .A2(n18847), .ZN(n12325) );
NAND2_X2 U7303 ( .A1(n12327), .A2(n12328), .ZN(n6109) );
NAND2_X2 U7304 ( .A1(aes_text_out[45]), .A2(n17993), .ZN(n12328) );
NAND2_X2 U7305 ( .A1(n17984), .A2(n17374), .ZN(n12327) );
NAND2_X2 U7306 ( .A1(n12329), .A2(n12330), .ZN(n6108) );
NAND2_X2 U7307 ( .A1(aes_text_out[46]), .A2(n17993), .ZN(n12330) );
NAND2_X2 U7308 ( .A1(n17984), .A2(n17373), .ZN(n12329) );
NAND2_X2 U7309 ( .A1(n12331), .A2(n12332), .ZN(n6107) );
NAND2_X2 U7310 ( .A1(aes_text_out[47]), .A2(n17993), .ZN(n12332) );
NAND2_X2 U7311 ( .A1(n17984), .A2(n17372), .ZN(n12331) );
NAND2_X2 U7312 ( .A1(n12333), .A2(n12334), .ZN(n6106) );
NAND2_X2 U7313 ( .A1(aes_text_out[48]), .A2(n17993), .ZN(n12334) );
NAND2_X2 U7314 ( .A1(n17984), .A2(n17371), .ZN(n12333) );
NAND2_X2 U7315 ( .A1(n12335), .A2(n12336), .ZN(n6105) );
NAND2_X2 U7316 ( .A1(aes_text_out[49]), .A2(n17993), .ZN(n12336) );
NAND2_X2 U7317 ( .A1(n17984), .A2(n17370), .ZN(n12335) );
NAND2_X2 U7318 ( .A1(n12337), .A2(n12338), .ZN(n6104) );
NAND2_X2 U7319 ( .A1(aes_text_out[50]), .A2(n17993), .ZN(n12338) );
NAND2_X2 U7320 ( .A1(n17984), .A2(n17369), .ZN(n12337) );
NAND2_X2 U7321 ( .A1(n12339), .A2(n12340), .ZN(n6103) );
NAND2_X2 U7322 ( .A1(aes_text_out[51]), .A2(n17993), .ZN(n12340) );
NAND2_X2 U7323 ( .A1(n17983), .A2(n17368), .ZN(n12339) );
NAND2_X2 U7324 ( .A1(n12341), .A2(n12342), .ZN(n6102) );
NAND2_X2 U7325 ( .A1(aes_text_out[52]), .A2(n17993), .ZN(n12342) );
NAND2_X2 U7326 ( .A1(n17983), .A2(n17367), .ZN(n12341) );
NAND2_X2 U7327 ( .A1(n12343), .A2(n12344), .ZN(n6101) );
NAND2_X2 U7328 ( .A1(aes_text_out[53]), .A2(n17993), .ZN(n12344) );
NAND2_X2 U7329 ( .A1(n17983), .A2(n17366), .ZN(n12343) );
NAND2_X2 U7330 ( .A1(n12345), .A2(n12346), .ZN(n6100) );
NAND2_X2 U7331 ( .A1(aes_text_out[54]), .A2(n17993), .ZN(n12346) );
NAND2_X2 U7332 ( .A1(n17983), .A2(n17365), .ZN(n12345) );
NAND2_X2 U7333 ( .A1(n12347), .A2(n12348), .ZN(n6099) );
NAND2_X2 U7334 ( .A1(aes_text_out[55]), .A2(n17993), .ZN(n12348) );
NAND2_X2 U7335 ( .A1(n17983), .A2(n17364), .ZN(n12347) );
NAND2_X2 U7336 ( .A1(n12349), .A2(n12350), .ZN(n6098) );
NAND2_X2 U7337 ( .A1(aes_text_out[56]), .A2(n17993), .ZN(n12350) );
NAND2_X2 U7338 ( .A1(n17983), .A2(n17363), .ZN(n12349) );
NAND2_X2 U7339 ( .A1(n12351), .A2(n12352), .ZN(n6097) );
NAND2_X2 U7340 ( .A1(aes_text_out[57]), .A2(n17993), .ZN(n12352) );
NAND2_X2 U7341 ( .A1(n17983), .A2(n17362), .ZN(n12351) );
NAND2_X2 U7342 ( .A1(n12353), .A2(n12354), .ZN(n6096) );
NAND2_X2 U7343 ( .A1(aes_text_out[58]), .A2(n17993), .ZN(n12354) );
NAND2_X2 U7344 ( .A1(n17983), .A2(n17361), .ZN(n12353) );
NAND2_X2 U7345 ( .A1(n12355), .A2(n12356), .ZN(n6095) );
NAND2_X2 U7346 ( .A1(aes_text_out[59]), .A2(n17993), .ZN(n12356) );
NAND2_X2 U7347 ( .A1(n17983), .A2(n17360), .ZN(n12355) );
NAND2_X2 U7348 ( .A1(n12357), .A2(n12358), .ZN(n6094) );
NAND2_X2 U7349 ( .A1(aes_text_out[60]), .A2(n17993), .ZN(n12358) );
NAND2_X2 U7350 ( .A1(n17983), .A2(n17359), .ZN(n12357) );
NAND2_X2 U7351 ( .A1(n12359), .A2(n12360), .ZN(n6093) );
NAND2_X2 U7352 ( .A1(aes_text_out[61]), .A2(n17993), .ZN(n12360) );
NAND2_X2 U7353 ( .A1(n17983), .A2(n17358), .ZN(n12359) );
NAND2_X2 U7354 ( .A1(n12361), .A2(n12362), .ZN(n6092) );
NAND2_X2 U7355 ( .A1(aes_text_out[62]), .A2(n17993), .ZN(n12362) );
NAND2_X2 U7356 ( .A1(n17982), .A2(n17357), .ZN(n12361) );
NAND2_X2 U7357 ( .A1(n12363), .A2(n12364), .ZN(n6091) );
NAND2_X2 U7358 ( .A1(aes_text_out[63]), .A2(n17993), .ZN(n12364) );
NAND2_X2 U7359 ( .A1(n17982), .A2(n17356), .ZN(n12363) );
NAND2_X2 U7360 ( .A1(n12365), .A2(n12366), .ZN(n6090) );
NAND2_X2 U7361 ( .A1(aes_text_out[64]), .A2(n17993), .ZN(n12366) );
NAND2_X2 U7362 ( .A1(n17982), .A2(n17355), .ZN(n12365) );
NAND2_X2 U7363 ( .A1(n12367), .A2(n12368), .ZN(n6089) );
NAND2_X2 U7364 ( .A1(aes_text_out[65]), .A2(n17993), .ZN(n12368) );
NAND2_X2 U7365 ( .A1(n17982), .A2(n17354), .ZN(n12367) );
NAND2_X2 U7366 ( .A1(n12369), .A2(n12370), .ZN(n6088) );
NAND2_X2 U7367 ( .A1(aes_text_out[66]), .A2(n17992), .ZN(n12370) );
NAND2_X2 U7368 ( .A1(n17982), .A2(n17353), .ZN(n12369) );
NAND2_X2 U7369 ( .A1(n12371), .A2(n12372), .ZN(n6087) );
NAND2_X2 U7370 ( .A1(aes_text_out[67]), .A2(n17992), .ZN(n12372) );
NAND2_X2 U7371 ( .A1(n17982), .A2(n17352), .ZN(n12371) );
NAND2_X2 U7372 ( .A1(n12373), .A2(n12374), .ZN(n6086) );
NAND2_X2 U7373 ( .A1(aes_text_out[68]), .A2(n17992), .ZN(n12374) );
NAND2_X2 U7374 ( .A1(n17982), .A2(n17351), .ZN(n12373) );
NAND2_X2 U7375 ( .A1(n12375), .A2(n12376), .ZN(n6085) );
NAND2_X2 U7376 ( .A1(aes_text_out[69]), .A2(n17992), .ZN(n12376) );
NAND2_X2 U7377 ( .A1(n17982), .A2(n17350), .ZN(n12375) );
NAND2_X2 U7378 ( .A1(n12377), .A2(n12378), .ZN(n6084) );
NAND2_X2 U7379 ( .A1(aes_text_out[70]), .A2(n17992), .ZN(n12378) );
NAND2_X2 U7380 ( .A1(n17982), .A2(n17349), .ZN(n12377) );
NAND2_X2 U7381 ( .A1(n12379), .A2(n12380), .ZN(n6083) );
NAND2_X2 U7382 ( .A1(aes_text_out[71]), .A2(n17992), .ZN(n12380) );
NAND2_X2 U7383 ( .A1(n17982), .A2(n17348), .ZN(n12379) );
NAND2_X2 U7384 ( .A1(n12381), .A2(n12382), .ZN(n6082) );
NAND2_X2 U7385 ( .A1(aes_text_out[72]), .A2(n17992), .ZN(n12382) );
NAND2_X2 U7386 ( .A1(n17982), .A2(n17347), .ZN(n12381) );
NAND2_X2 U7387 ( .A1(n12383), .A2(n12384), .ZN(n6081) );
NAND2_X2 U7388 ( .A1(aes_text_out[73]), .A2(n17992), .ZN(n12384) );
NAND2_X2 U7389 ( .A1(n17981), .A2(n17346), .ZN(n12383) );
NAND2_X2 U7390 ( .A1(n12385), .A2(n12386), .ZN(n6080) );
NAND2_X2 U7391 ( .A1(aes_text_out[74]), .A2(n17992), .ZN(n12386) );
NAND2_X2 U7392 ( .A1(n17981), .A2(n17345), .ZN(n12385) );
NAND2_X2 U7393 ( .A1(n12387), .A2(n12388), .ZN(n6079) );
NAND2_X2 U7394 ( .A1(aes_text_out[75]), .A2(n17992), .ZN(n12388) );
NAND2_X2 U7395 ( .A1(n17981), .A2(n17344), .ZN(n12387) );
NAND2_X2 U7396 ( .A1(n12389), .A2(n12390), .ZN(n6078) );
NAND2_X2 U7397 ( .A1(aes_text_out[76]), .A2(n17992), .ZN(n12390) );
NAND2_X2 U7398 ( .A1(n17981), .A2(n17343), .ZN(n12389) );
NAND2_X2 U7399 ( .A1(n12391), .A2(n12392), .ZN(n6077) );
NAND2_X2 U7400 ( .A1(aes_text_out[77]), .A2(n17992), .ZN(n12392) );
NAND2_X2 U7401 ( .A1(n17981), .A2(n17342), .ZN(n12391) );
NAND2_X2 U7402 ( .A1(n12393), .A2(n12394), .ZN(n6076) );
NAND2_X2 U7403 ( .A1(aes_text_out[78]), .A2(n17992), .ZN(n12394) );
NAND2_X2 U7404 ( .A1(n17981), .A2(n17341), .ZN(n12393) );
NAND2_X2 U7405 ( .A1(n12395), .A2(n12396), .ZN(n6075) );
NAND2_X2 U7406 ( .A1(aes_text_out[79]), .A2(n17992), .ZN(n12396) );
NAND2_X2 U7407 ( .A1(n17981), .A2(n17340), .ZN(n12395) );
NAND2_X2 U7408 ( .A1(n12397), .A2(n12398), .ZN(n6074) );
NAND2_X2 U7409 ( .A1(aes_text_out[80]), .A2(n17992), .ZN(n12398) );
NAND2_X2 U7410 ( .A1(n17981), .A2(n17339), .ZN(n12397) );
NAND2_X2 U7411 ( .A1(n12399), .A2(n12400), .ZN(n6073) );
NAND2_X2 U7412 ( .A1(aes_text_out[81]), .A2(n17992), .ZN(n12400) );
NAND2_X2 U7413 ( .A1(n17981), .A2(n17338), .ZN(n12399) );
NAND2_X2 U7414 ( .A1(n12401), .A2(n12402), .ZN(n6072) );
NAND2_X2 U7415 ( .A1(aes_text_out[82]), .A2(n17992), .ZN(n12402) );
NAND2_X2 U7416 ( .A1(n17981), .A2(n17337), .ZN(n12401) );
NAND2_X2 U7417 ( .A1(n12403), .A2(n12404), .ZN(n6071) );
NAND2_X2 U7418 ( .A1(aes_text_out[83]), .A2(n17992), .ZN(n12404) );
NAND2_X2 U7419 ( .A1(n17981), .A2(n17336), .ZN(n12403) );
NAND2_X2 U7420 ( .A1(n12405), .A2(n12406), .ZN(n6070) );
NAND2_X2 U7421 ( .A1(aes_text_out[84]), .A2(n17992), .ZN(n12406) );
NAND2_X2 U7422 ( .A1(n17980), .A2(n17335), .ZN(n12405) );
NAND2_X2 U7423 ( .A1(n12407), .A2(n12408), .ZN(n6069) );
NAND2_X2 U7424 ( .A1(aes_text_out[85]), .A2(n17992), .ZN(n12408) );
NAND2_X2 U7425 ( .A1(n17980), .A2(n17334), .ZN(n12407) );
NAND2_X2 U7426 ( .A1(n12409), .A2(n12410), .ZN(n6068) );
NAND2_X2 U7427 ( .A1(aes_text_out[86]), .A2(n17992), .ZN(n12410) );
NAND2_X2 U7428 ( .A1(n17980), .A2(n17333), .ZN(n12409) );
NAND2_X2 U7429 ( .A1(n12411), .A2(n12412), .ZN(n6067) );
NAND2_X2 U7430 ( .A1(aes_text_out[87]), .A2(n17991), .ZN(n12412) );
NAND2_X2 U7431 ( .A1(n17980), .A2(n17332), .ZN(n12411) );
NAND2_X2 U7432 ( .A1(n12413), .A2(n12414), .ZN(n6066) );
NAND2_X2 U7433 ( .A1(aes_text_out[88]), .A2(n17991), .ZN(n12414) );
NAND2_X2 U7434 ( .A1(n17980), .A2(n17331), .ZN(n12413) );
NAND2_X2 U7435 ( .A1(n12415), .A2(n12416), .ZN(n6065) );
NAND2_X2 U7436 ( .A1(aes_text_out[89]), .A2(n17991), .ZN(n12416) );
NAND2_X2 U7437 ( .A1(n17980), .A2(n17330), .ZN(n12415) );
NAND2_X2 U7438 ( .A1(n12417), .A2(n12418), .ZN(n6064) );
NAND2_X2 U7439 ( .A1(aes_text_out[90]), .A2(n17991), .ZN(n12418) );
NAND2_X2 U7440 ( .A1(n17980), .A2(n17329), .ZN(n12417) );
NAND2_X2 U7441 ( .A1(n12419), .A2(n12420), .ZN(n6063) );
NAND2_X2 U7442 ( .A1(aes_text_out[91]), .A2(n17991), .ZN(n12420) );
NAND2_X2 U7443 ( .A1(n17980), .A2(n17328), .ZN(n12419) );
NAND2_X2 U7444 ( .A1(n12421), .A2(n12422), .ZN(n6062) );
NAND2_X2 U7445 ( .A1(aes_text_out[92]), .A2(n17991), .ZN(n12422) );
NAND2_X2 U7446 ( .A1(n17980), .A2(n17327), .ZN(n12421) );
NAND2_X2 U7447 ( .A1(n12423), .A2(n12424), .ZN(n6061) );
NAND2_X2 U7448 ( .A1(aes_text_out[93]), .A2(n17991), .ZN(n12424) );
NAND2_X2 U7449 ( .A1(n17980), .A2(n17326), .ZN(n12423) );
NAND2_X2 U7450 ( .A1(n12425), .A2(n12426), .ZN(n6060) );
NAND2_X2 U7451 ( .A1(aes_text_out[94]), .A2(n17991), .ZN(n12426) );
NAND2_X2 U7452 ( .A1(n17980), .A2(n17325), .ZN(n12425) );
NAND2_X2 U7453 ( .A1(n12427), .A2(n12428), .ZN(n6059) );
NAND2_X2 U7454 ( .A1(aes_text_out[95]), .A2(n17991), .ZN(n12428) );
NAND2_X2 U7455 ( .A1(n17979), .A2(n17324), .ZN(n12427) );
NAND2_X2 U7456 ( .A1(n12429), .A2(n12430), .ZN(n6058) );
NAND2_X2 U7457 ( .A1(aes_text_out[96]), .A2(n17991), .ZN(n12430) );
NAND2_X2 U7458 ( .A1(n17979), .A2(n17323), .ZN(n12429) );
NAND2_X2 U7459 ( .A1(n12431), .A2(n12432), .ZN(n6057) );
NAND2_X2 U7460 ( .A1(aes_text_out[97]), .A2(n17991), .ZN(n12432) );
NAND2_X2 U7461 ( .A1(n17979), .A2(n17322), .ZN(n12431) );
NAND2_X2 U7462 ( .A1(n12433), .A2(n12434), .ZN(n6056) );
NAND2_X2 U7463 ( .A1(aes_text_out[98]), .A2(n17991), .ZN(n12434) );
NAND2_X2 U7464 ( .A1(n17979), .A2(n17321), .ZN(n12433) );
NAND2_X2 U7465 ( .A1(n12435), .A2(n12436), .ZN(n6055) );
NAND2_X2 U7466 ( .A1(aes_text_out[99]), .A2(n17991), .ZN(n12436) );
NAND2_X2 U7467 ( .A1(n17979), .A2(n17320), .ZN(n12435) );
NAND2_X2 U7468 ( .A1(n12437), .A2(n12438), .ZN(n6054) );
NAND2_X2 U7469 ( .A1(aes_text_out[100]), .A2(n17991), .ZN(n12438) );
NAND2_X2 U7470 ( .A1(n17979), .A2(n17319), .ZN(n12437) );
NAND2_X2 U7471 ( .A1(n12439), .A2(n12440), .ZN(n6053) );
NAND2_X2 U7472 ( .A1(aes_text_out[101]), .A2(n17991), .ZN(n12440) );
NAND2_X2 U7473 ( .A1(n17979), .A2(n17318), .ZN(n12439) );
NAND2_X2 U7474 ( .A1(n12441), .A2(n12442), .ZN(n6052) );
NAND2_X2 U7475 ( .A1(aes_text_out[102]), .A2(n17991), .ZN(n12442) );
NAND2_X2 U7476 ( .A1(n17979), .A2(n17317), .ZN(n12441) );
NAND2_X2 U7477 ( .A1(n12443), .A2(n12444), .ZN(n6051) );
NAND2_X2 U7478 ( .A1(aes_text_out[103]), .A2(n17991), .ZN(n12444) );
NAND2_X2 U7479 ( .A1(n17979), .A2(n17316), .ZN(n12443) );
NAND2_X2 U7480 ( .A1(n12445), .A2(n12446), .ZN(n6050) );
NAND2_X2 U7481 ( .A1(aes_text_out[104]), .A2(n17991), .ZN(n12446) );
NAND2_X2 U7482 ( .A1(n17979), .A2(n17315), .ZN(n12445) );
NAND2_X2 U7483 ( .A1(n12447), .A2(n12448), .ZN(n6049) );
NAND2_X2 U7484 ( .A1(aes_text_out[105]), .A2(n17991), .ZN(n12448) );
NAND2_X2 U7485 ( .A1(n17979), .A2(n17314), .ZN(n12447) );
NAND2_X2 U7486 ( .A1(n12449), .A2(n12450), .ZN(n6048) );
NAND2_X2 U7487 ( .A1(aes_text_out[106]), .A2(n17991), .ZN(n12450) );
NAND2_X2 U7488 ( .A1(n17978), .A2(n17313), .ZN(n12449) );
NAND2_X2 U7489 ( .A1(n12451), .A2(n12452), .ZN(n6047) );
NAND2_X2 U7490 ( .A1(aes_text_out[107]), .A2(n17991), .ZN(n12452) );
NAND2_X2 U7491 ( .A1(n17978), .A2(n17312), .ZN(n12451) );
NAND2_X2 U7492 ( .A1(n12453), .A2(n12454), .ZN(n6046) );
NAND2_X2 U7493 ( .A1(aes_text_out[108]), .A2(n17990), .ZN(n12454) );
NAND2_X2 U7494 ( .A1(n17978), .A2(n17311), .ZN(n12453) );
NAND2_X2 U7495 ( .A1(n12455), .A2(n12456), .ZN(n6045) );
NAND2_X2 U7496 ( .A1(aes_text_out[109]), .A2(n17990), .ZN(n12456) );
NAND2_X2 U7497 ( .A1(n17978), .A2(n17310), .ZN(n12455) );
NAND2_X2 U7498 ( .A1(n12457), .A2(n12458), .ZN(n6044) );
NAND2_X2 U7499 ( .A1(aes_text_out[110]), .A2(n17990), .ZN(n12458) );
NAND2_X2 U7500 ( .A1(n17978), .A2(n17309), .ZN(n12457) );
NAND2_X2 U7501 ( .A1(n12459), .A2(n12460), .ZN(n6043) );
NAND2_X2 U7502 ( .A1(aes_text_out[111]), .A2(n17990), .ZN(n12460) );
NAND2_X2 U7503 ( .A1(n17978), .A2(n17308), .ZN(n12459) );
NAND2_X2 U7504 ( .A1(n12461), .A2(n12462), .ZN(n6042) );
NAND2_X2 U7505 ( .A1(aes_text_out[112]), .A2(n17990), .ZN(n12462) );
NAND2_X2 U7506 ( .A1(n17978), .A2(n17307), .ZN(n12461) );
NAND2_X2 U7507 ( .A1(n12463), .A2(n12464), .ZN(n6041) );
NAND2_X2 U7508 ( .A1(aes_text_out[113]), .A2(n17990), .ZN(n12464) );
NAND2_X2 U7509 ( .A1(n17978), .A2(n17306), .ZN(n12463) );
NAND2_X2 U7510 ( .A1(n12465), .A2(n12466), .ZN(n6040) );
NAND2_X2 U7511 ( .A1(aes_text_out[114]), .A2(n17990), .ZN(n12466) );
NAND2_X2 U7512 ( .A1(n17978), .A2(n17305), .ZN(n12465) );
NAND2_X2 U7513 ( .A1(n12467), .A2(n12468), .ZN(n6039) );
NAND2_X2 U7514 ( .A1(aes_text_out[115]), .A2(n17990), .ZN(n12468) );
NAND2_X2 U7515 ( .A1(n17978), .A2(n17304), .ZN(n12467) );
NAND2_X2 U7516 ( .A1(n12469), .A2(n12470), .ZN(n6038) );
NAND2_X2 U7517 ( .A1(aes_text_out[116]), .A2(n17990), .ZN(n12470) );
NAND2_X2 U7518 ( .A1(n17978), .A2(n17303), .ZN(n12469) );
NAND2_X2 U7519 ( .A1(n12471), .A2(n12472), .ZN(n6037) );
NAND2_X2 U7520 ( .A1(aes_text_out[117]), .A2(n17990), .ZN(n12472) );
NAND2_X2 U7521 ( .A1(n17977), .A2(n17302), .ZN(n12471) );
NAND2_X2 U7522 ( .A1(n12473), .A2(n12474), .ZN(n6036) );
NAND2_X2 U7523 ( .A1(aes_text_out[118]), .A2(n17990), .ZN(n12474) );
NAND2_X2 U7524 ( .A1(n17977), .A2(n17301), .ZN(n12473) );
NAND2_X2 U7525 ( .A1(n12475), .A2(n12476), .ZN(n6035) );
NAND2_X2 U7526 ( .A1(aes_text_out[119]), .A2(n17990), .ZN(n12476) );
NAND2_X2 U7527 ( .A1(n17977), .A2(n17300), .ZN(n12475) );
NAND2_X2 U7528 ( .A1(n12477), .A2(n12478), .ZN(n6034) );
NAND2_X2 U7529 ( .A1(aes_text_out[120]), .A2(n17990), .ZN(n12478) );
NAND2_X2 U7530 ( .A1(n17977), .A2(n17299), .ZN(n12477) );
NAND2_X2 U7531 ( .A1(n12479), .A2(n12480), .ZN(n6033) );
NAND2_X2 U7532 ( .A1(aes_text_out[121]), .A2(n17990), .ZN(n12480) );
NAND2_X2 U7533 ( .A1(n17977), .A2(n17298), .ZN(n12479) );
NAND2_X2 U7534 ( .A1(n12481), .A2(n12482), .ZN(n6032) );
NAND2_X2 U7535 ( .A1(aes_text_out[122]), .A2(n17990), .ZN(n12482) );
NAND2_X2 U7536 ( .A1(n17977), .A2(n17297), .ZN(n12481) );
NAND2_X2 U7537 ( .A1(n12483), .A2(n12484), .ZN(n6031) );
NAND2_X2 U7538 ( .A1(aes_text_out[123]), .A2(n17990), .ZN(n12484) );
NAND2_X2 U7539 ( .A1(n17977), .A2(n17296), .ZN(n12483) );
NAND2_X2 U7540 ( .A1(n12485), .A2(n12486), .ZN(n6030) );
NAND2_X2 U7541 ( .A1(aes_text_out[124]), .A2(n17990), .ZN(n12486) );
NAND2_X2 U7542 ( .A1(n17977), .A2(n17295), .ZN(n12485) );
NAND2_X2 U7543 ( .A1(n12487), .A2(n12488), .ZN(n6029) );
NAND2_X2 U7544 ( .A1(aes_text_out[125]), .A2(n17990), .ZN(n12488) );
NAND2_X2 U7545 ( .A1(n17977), .A2(n17294), .ZN(n12487) );
NAND2_X2 U7546 ( .A1(n12489), .A2(n12490), .ZN(n6028) );
NAND2_X2 U7547 ( .A1(aes_text_out[126]), .A2(n17990), .ZN(n12490) );
NAND2_X2 U7548 ( .A1(n17977), .A2(n17293), .ZN(n12489) );
NAND2_X2 U7549 ( .A1(n12491), .A2(n12492), .ZN(n6027) );
NAND2_X2 U7550 ( .A1(aes_text_out[127]), .A2(n17990), .ZN(n12492) );
NAND2_X2 U7551 ( .A1(n17977), .A2(n17292), .ZN(n12491) );
NAND2_X2 U7552 ( .A1(n12493), .A2(n12494), .ZN(n6026) );
NAND2_X2 U7553 ( .A1(n17750), .A2(n17281), .ZN(n12494) );
NAND2_X2 U7554 ( .A1(n18744), .A2(Out_data_size[0]), .ZN(n12493) );
NAND2_X2 U7557 ( .A1(n18744), .A2(Out_data_size[1]), .ZN(n12495) );
NAND2_X2 U7560 ( .A1(n18744), .A2(Out_data_size[2]), .ZN(n12497) );
NAND2_X2 U7561 ( .A1(n12499), .A2(n12500), .ZN(n6023) );
NAND2_X2 U7562 ( .A1(n18074), .A2(n17281), .ZN(n12500) );
NAND2_X2 U7563 ( .A1(n18744), .A2(Out_data_size[3]), .ZN(n12499) );
NAND2_X2 U7564 ( .A1(n12501), .A2(n12502), .ZN(n6022) );
NAND2_X2 U7565 ( .A1(n17281), .A2(n17748), .ZN(n12502) );
NAND2_X2 U7566 ( .A1(n18744), .A2(Out_last_word), .ZN(n12501) );
NAND2_X2 U8275 ( .A1(n11967), .A2(aes_done), .ZN(n12238) );
AND4_X2 U8276 ( .A1(state[1]), .A2(n18628), .A3(n18625), .A4(n18629), .ZN(n11967) );
NAND2_X2 U8277 ( .A1(n13019), .A2(n13020), .ZN(n5829) );
NAND2_X2 U8278 ( .A1(n17976), .A2(n18895), .ZN(n13020) );
NAND2_X2 U8279 ( .A1(z_out[0]), .A2(n17961), .ZN(n13019) );
NAND2_X2 U8280 ( .A1(n13023), .A2(n13024), .ZN(n5828) );
NAND2_X2 U8281 ( .A1(n17976), .A2(n18896), .ZN(n13024) );
NAND2_X2 U8282 ( .A1(z_out[1]), .A2(n17958), .ZN(n13023) );
NAND2_X2 U8283 ( .A1(n13025), .A2(n13026), .ZN(n5827) );
NAND2_X2 U8284 ( .A1(n17976), .A2(n18897), .ZN(n13026) );
NAND2_X2 U8285 ( .A1(z_out[2]), .A2(n17958), .ZN(n13025) );
NAND2_X2 U8286 ( .A1(n13027), .A2(n13028), .ZN(n5826) );
NAND2_X2 U8287 ( .A1(n17976), .A2(n18898), .ZN(n13028) );
NAND2_X2 U8288 ( .A1(z_out[3]), .A2(n17958), .ZN(n13027) );
NAND2_X2 U8289 ( .A1(n13029), .A2(n13030), .ZN(n5825) );
NAND2_X2 U8290 ( .A1(n17976), .A2(n18899), .ZN(n13030) );
NAND2_X2 U8291 ( .A1(z_out[4]), .A2(n17958), .ZN(n13029) );
NAND2_X2 U8292 ( .A1(n13031), .A2(n13032), .ZN(n5824) );
NAND2_X2 U8293 ( .A1(n17976), .A2(n18900), .ZN(n13032) );
NAND2_X2 U8294 ( .A1(z_out[5]), .A2(n17958), .ZN(n13031) );
NAND2_X2 U8295 ( .A1(n13033), .A2(n13034), .ZN(n5823) );
NAND2_X2 U8296 ( .A1(n17976), .A2(n18901), .ZN(n13034) );
NAND2_X2 U8297 ( .A1(z_out[6]), .A2(n17958), .ZN(n13033) );
NAND2_X2 U8298 ( .A1(n13035), .A2(n13036), .ZN(n5822) );
NAND2_X2 U8299 ( .A1(n17975), .A2(n18902), .ZN(n13036) );
NAND2_X2 U8300 ( .A1(z_out[7]), .A2(n17958), .ZN(n13035) );
NAND2_X2 U8301 ( .A1(n13037), .A2(n13038), .ZN(n5821) );
NAND2_X2 U8302 ( .A1(n17975), .A2(n18903), .ZN(n13038) );
NAND2_X2 U8303 ( .A1(z_out[8]), .A2(n17958), .ZN(n13037) );
NAND2_X2 U8304 ( .A1(n13039), .A2(n13040), .ZN(n5820) );
NAND2_X2 U8305 ( .A1(n17975), .A2(n18904), .ZN(n13040) );
NAND2_X2 U8306 ( .A1(z_out[9]), .A2(n17958), .ZN(n13039) );
NAND2_X2 U8307 ( .A1(n13041), .A2(n13042), .ZN(n5819) );
NAND2_X2 U8308 ( .A1(n17975), .A2(n18905), .ZN(n13042) );
NAND2_X2 U8309 ( .A1(z_out[10]), .A2(n17958), .ZN(n13041) );
NAND2_X2 U8310 ( .A1(n13043), .A2(n13044), .ZN(n5818) );
NAND2_X2 U8311 ( .A1(n17975), .A2(n18906), .ZN(n13044) );
NAND2_X2 U8312 ( .A1(z_out[11]), .A2(n17958), .ZN(n13043) );
NAND2_X2 U8313 ( .A1(n13045), .A2(n13046), .ZN(n5817) );
NAND2_X2 U8314 ( .A1(n17975), .A2(n18907), .ZN(n13046) );
NAND2_X2 U8315 ( .A1(z_out[12]), .A2(n17958), .ZN(n13045) );
NAND2_X2 U8316 ( .A1(n13047), .A2(n13048), .ZN(n5816) );
NAND2_X2 U8317 ( .A1(n17975), .A2(n18908), .ZN(n13048) );
NAND2_X2 U8318 ( .A1(z_out[13]), .A2(n17958), .ZN(n13047) );
NAND2_X2 U8319 ( .A1(n13049), .A2(n13050), .ZN(n5815) );
NAND2_X2 U8320 ( .A1(n17975), .A2(n18909), .ZN(n13050) );
NAND2_X2 U8321 ( .A1(z_out[14]), .A2(n17958), .ZN(n13049) );
NAND2_X2 U8322 ( .A1(n13051), .A2(n13052), .ZN(n5814) );
NAND2_X2 U8323 ( .A1(n17975), .A2(n18910), .ZN(n13052) );
NAND2_X2 U8324 ( .A1(z_out[15]), .A2(n17958), .ZN(n13051) );
NAND2_X2 U8325 ( .A1(n13053), .A2(n13054), .ZN(n5813) );
NAND2_X2 U8326 ( .A1(n17975), .A2(n18911), .ZN(n13054) );
NAND2_X2 U8327 ( .A1(z_out[16]), .A2(n17958), .ZN(n13053) );
NAND2_X2 U8328 ( .A1(n13055), .A2(n13056), .ZN(n5812) );
NAND2_X2 U8329 ( .A1(n17975), .A2(n18912), .ZN(n13056) );
NAND2_X2 U8330 ( .A1(z_out[17]), .A2(n17958), .ZN(n13055) );
NAND2_X2 U8331 ( .A1(n13057), .A2(n13058), .ZN(n5811) );
NAND2_X2 U8332 ( .A1(n17974), .A2(n18913), .ZN(n13058) );
NAND2_X2 U8333 ( .A1(z_out[18]), .A2(n17959), .ZN(n13057) );
NAND2_X2 U8334 ( .A1(n13059), .A2(n13060), .ZN(n5810) );
NAND2_X2 U8335 ( .A1(n17974), .A2(n18914), .ZN(n13060) );
NAND2_X2 U8336 ( .A1(z_out[19]), .A2(n17959), .ZN(n13059) );
NAND2_X2 U8337 ( .A1(n13061), .A2(n13062), .ZN(n5809) );
NAND2_X2 U8338 ( .A1(n17974), .A2(n18915), .ZN(n13062) );
NAND2_X2 U8339 ( .A1(z_out[20]), .A2(n17959), .ZN(n13061) );
NAND2_X2 U8340 ( .A1(n13063), .A2(n13064), .ZN(n5808) );
NAND2_X2 U8341 ( .A1(n17974), .A2(n18916), .ZN(n13064) );
NAND2_X2 U8342 ( .A1(z_out[21]), .A2(n17959), .ZN(n13063) );
NAND2_X2 U8343 ( .A1(n13065), .A2(n13066), .ZN(n5807) );
NAND2_X2 U8344 ( .A1(n17974), .A2(n18917), .ZN(n13066) );
NAND2_X2 U8345 ( .A1(z_out[22]), .A2(n17959), .ZN(n13065) );
NAND2_X2 U8346 ( .A1(n13067), .A2(n13068), .ZN(n5806) );
NAND2_X2 U8347 ( .A1(n17974), .A2(n18918), .ZN(n13068) );
NAND2_X2 U8348 ( .A1(z_out[23]), .A2(n17959), .ZN(n13067) );
NAND2_X2 U8349 ( .A1(n13069), .A2(n13070), .ZN(n5805) );
NAND2_X2 U8350 ( .A1(n17974), .A2(n18919), .ZN(n13070) );
NAND2_X2 U8351 ( .A1(z_out[24]), .A2(n17959), .ZN(n13069) );
NAND2_X2 U8352 ( .A1(n13071), .A2(n13072), .ZN(n5804) );
NAND2_X2 U8353 ( .A1(n17974), .A2(n18920), .ZN(n13072) );
NAND2_X2 U8354 ( .A1(z_out[25]), .A2(n17959), .ZN(n13071) );
NAND2_X2 U8355 ( .A1(n13073), .A2(n13074), .ZN(n5803) );
NAND2_X2 U8356 ( .A1(n17974), .A2(n18921), .ZN(n13074) );
NAND2_X2 U8357 ( .A1(z_out[26]), .A2(n17959), .ZN(n13073) );
NAND2_X2 U8358 ( .A1(n13075), .A2(n13076), .ZN(n5802) );
NAND2_X2 U8359 ( .A1(n17974), .A2(n18922), .ZN(n13076) );
NAND2_X2 U8360 ( .A1(z_out[27]), .A2(n17959), .ZN(n13075) );
NAND2_X2 U8361 ( .A1(n13077), .A2(n13078), .ZN(n5801) );
NAND2_X2 U8362 ( .A1(n17974), .A2(n18923), .ZN(n13078) );
NAND2_X2 U8363 ( .A1(z_out[28]), .A2(n17959), .ZN(n13077) );
NAND2_X2 U8364 ( .A1(n13079), .A2(n13080), .ZN(n5800) );
NAND2_X2 U8365 ( .A1(n17973), .A2(n18924), .ZN(n13080) );
NAND2_X2 U8366 ( .A1(z_out[29]), .A2(n17959), .ZN(n13079) );
NAND2_X2 U8367 ( .A1(n13081), .A2(n13082), .ZN(n5799) );
NAND2_X2 U8368 ( .A1(n17973), .A2(n18925), .ZN(n13082) );
NAND2_X2 U8369 ( .A1(z_out[30]), .A2(n17959), .ZN(n13081) );
NAND2_X2 U8370 ( .A1(n13083), .A2(n13084), .ZN(n5798) );
NAND2_X2 U8371 ( .A1(n17973), .A2(n18926), .ZN(n13084) );
NAND2_X2 U8372 ( .A1(z_out[31]), .A2(n17959), .ZN(n13083) );
NAND2_X2 U8373 ( .A1(n13085), .A2(n13086), .ZN(n5797) );
NAND2_X2 U8374 ( .A1(n17973), .A2(n18927), .ZN(n13086) );
NAND2_X2 U8375 ( .A1(z_out[32]), .A2(n17959), .ZN(n13085) );
NAND2_X2 U8376 ( .A1(n13087), .A2(n13088), .ZN(n5796) );
NAND2_X2 U8377 ( .A1(n17973), .A2(n18928), .ZN(n13088) );
NAND2_X2 U8378 ( .A1(z_out[33]), .A2(n17959), .ZN(n13087) );
NAND2_X2 U8379 ( .A1(n13089), .A2(n13090), .ZN(n5795) );
NAND2_X2 U8380 ( .A1(n17973), .A2(n18929), .ZN(n13090) );
NAND2_X2 U8381 ( .A1(z_out[34]), .A2(n17959), .ZN(n13089) );
NAND2_X2 U8382 ( .A1(n13091), .A2(n13092), .ZN(n5794) );
NAND2_X2 U8383 ( .A1(n17973), .A2(n18930), .ZN(n13092) );
NAND2_X2 U8384 ( .A1(z_out[35]), .A2(n17959), .ZN(n13091) );
NAND2_X2 U8385 ( .A1(n13093), .A2(n13094), .ZN(n5793) );
NAND2_X2 U8386 ( .A1(n17973), .A2(n18931), .ZN(n13094) );
NAND2_X2 U8387 ( .A1(z_out[36]), .A2(n17959), .ZN(n13093) );
NAND2_X2 U8388 ( .A1(n13095), .A2(n13096), .ZN(n5792) );
NAND2_X2 U8389 ( .A1(n17973), .A2(n18932), .ZN(n13096) );
NAND2_X2 U8390 ( .A1(z_out[37]), .A2(n17960), .ZN(n13095) );
NAND2_X2 U8391 ( .A1(n13097), .A2(n13098), .ZN(n5791) );
NAND2_X2 U8392 ( .A1(n17973), .A2(n18933), .ZN(n13098) );
NAND2_X2 U8393 ( .A1(z_out[38]), .A2(n17960), .ZN(n13097) );
NAND2_X2 U8394 ( .A1(n13099), .A2(n13100), .ZN(n5790) );
NAND2_X2 U8395 ( .A1(n17973), .A2(n18934), .ZN(n13100) );
NAND2_X2 U8396 ( .A1(z_out[39]), .A2(n17960), .ZN(n13099) );
NAND2_X2 U8397 ( .A1(n13101), .A2(n13102), .ZN(n5789) );
NAND2_X2 U8398 ( .A1(n17972), .A2(n18935), .ZN(n13102) );
NAND2_X2 U8399 ( .A1(z_out[40]), .A2(n17960), .ZN(n13101) );
NAND2_X2 U8400 ( .A1(n13103), .A2(n13104), .ZN(n5788) );
NAND2_X2 U8401 ( .A1(n17972), .A2(n18936), .ZN(n13104) );
NAND2_X2 U8402 ( .A1(z_out[41]), .A2(n17960), .ZN(n13103) );
NAND2_X2 U8403 ( .A1(n13105), .A2(n13106), .ZN(n5787) );
NAND2_X2 U8404 ( .A1(n17972), .A2(n18937), .ZN(n13106) );
NAND2_X2 U8405 ( .A1(z_out[42]), .A2(n17960), .ZN(n13105) );
NAND2_X2 U8406 ( .A1(n13107), .A2(n13108), .ZN(n5786) );
NAND2_X2 U8407 ( .A1(n17972), .A2(n18938), .ZN(n13108) );
NAND2_X2 U8408 ( .A1(z_out[43]), .A2(n17960), .ZN(n13107) );
NAND2_X2 U8409 ( .A1(n13109), .A2(n13110), .ZN(n5785) );
NAND2_X2 U8410 ( .A1(n17972), .A2(n18939), .ZN(n13110) );
NAND2_X2 U8411 ( .A1(z_out[44]), .A2(n17960), .ZN(n13109) );
NAND2_X2 U8412 ( .A1(n13111), .A2(n13112), .ZN(n5784) );
NAND2_X2 U8413 ( .A1(n17972), .A2(n18940), .ZN(n13112) );
NAND2_X2 U8414 ( .A1(z_out[45]), .A2(n17960), .ZN(n13111) );
NAND2_X2 U8415 ( .A1(n13113), .A2(n13114), .ZN(n5783) );
NAND2_X2 U8416 ( .A1(n17972), .A2(n18941), .ZN(n13114) );
NAND2_X2 U8417 ( .A1(z_out[46]), .A2(n17960), .ZN(n13113) );
NAND2_X2 U8418 ( .A1(n13115), .A2(n13116), .ZN(n5782) );
NAND2_X2 U8419 ( .A1(n17972), .A2(n18942), .ZN(n13116) );
NAND2_X2 U8420 ( .A1(z_out[47]), .A2(n17960), .ZN(n13115) );
NAND2_X2 U8421 ( .A1(n13117), .A2(n13118), .ZN(n5781) );
NAND2_X2 U8422 ( .A1(n17972), .A2(n18943), .ZN(n13118) );
NAND2_X2 U8423 ( .A1(z_out[48]), .A2(n17960), .ZN(n13117) );
NAND2_X2 U8424 ( .A1(n13119), .A2(n13120), .ZN(n5780) );
NAND2_X2 U8425 ( .A1(n17972), .A2(n18944), .ZN(n13120) );
NAND2_X2 U8426 ( .A1(z_out[49]), .A2(n17960), .ZN(n13119) );
NAND2_X2 U8427 ( .A1(n13121), .A2(n13122), .ZN(n5779) );
NAND2_X2 U8428 ( .A1(n17972), .A2(n18945), .ZN(n13122) );
NAND2_X2 U8429 ( .A1(z_out[50]), .A2(n17960), .ZN(n13121) );
NAND2_X2 U8430 ( .A1(n13123), .A2(n13124), .ZN(n5778) );
NAND2_X2 U8431 ( .A1(n17971), .A2(n18946), .ZN(n13124) );
NAND2_X2 U8432 ( .A1(z_out[51]), .A2(n17960), .ZN(n13123) );
NAND2_X2 U8433 ( .A1(n13125), .A2(n13126), .ZN(n5777) );
NAND2_X2 U8434 ( .A1(n17971), .A2(n18947), .ZN(n13126) );
NAND2_X2 U8435 ( .A1(z_out[52]), .A2(n17960), .ZN(n13125) );
NAND2_X2 U8436 ( .A1(n13127), .A2(n13128), .ZN(n5776) );
NAND2_X2 U8437 ( .A1(n17971), .A2(n18948), .ZN(n13128) );
NAND2_X2 U8438 ( .A1(z_out[53]), .A2(n17960), .ZN(n13127) );
NAND2_X2 U8439 ( .A1(n13129), .A2(n13130), .ZN(n5775) );
NAND2_X2 U8440 ( .A1(n17971), .A2(n18949), .ZN(n13130) );
NAND2_X2 U8441 ( .A1(z_out[54]), .A2(n17960), .ZN(n13129) );
NAND2_X2 U8442 ( .A1(n13131), .A2(n13132), .ZN(n5774) );
NAND2_X2 U8443 ( .A1(n17971), .A2(n18950), .ZN(n13132) );
NAND2_X2 U8444 ( .A1(z_out[55]), .A2(n17960), .ZN(n13131) );
NAND2_X2 U8445 ( .A1(n13133), .A2(n13134), .ZN(n5773) );
NAND2_X2 U8446 ( .A1(n17971), .A2(n18951), .ZN(n13134) );
NAND2_X2 U8447 ( .A1(z_out[56]), .A2(n17961), .ZN(n13133) );
NAND2_X2 U8448 ( .A1(n13135), .A2(n13136), .ZN(n5772) );
NAND2_X2 U8449 ( .A1(n17971), .A2(n18952), .ZN(n13136) );
NAND2_X2 U8450 ( .A1(z_out[57]), .A2(n17961), .ZN(n13135) );
NAND2_X2 U8451 ( .A1(n13137), .A2(n13138), .ZN(n5771) );
NAND2_X2 U8452 ( .A1(n17971), .A2(n18953), .ZN(n13138) );
NAND2_X2 U8453 ( .A1(z_out[58]), .A2(n17961), .ZN(n13137) );
NAND2_X2 U8454 ( .A1(n13139), .A2(n13140), .ZN(n5770) );
NAND2_X2 U8455 ( .A1(n17971), .A2(n18954), .ZN(n13140) );
NAND2_X2 U8456 ( .A1(z_out[59]), .A2(n17961), .ZN(n13139) );
NAND2_X2 U8457 ( .A1(n13141), .A2(n13142), .ZN(n5769) );
NAND2_X2 U8458 ( .A1(n17971), .A2(n18955), .ZN(n13142) );
NAND2_X2 U8459 ( .A1(z_out[60]), .A2(n17961), .ZN(n13141) );
NAND2_X2 U8460 ( .A1(n13143), .A2(n13144), .ZN(n5768) );
NAND2_X2 U8461 ( .A1(n17971), .A2(n18956), .ZN(n13144) );
NAND2_X2 U8462 ( .A1(z_out[61]), .A2(n17961), .ZN(n13143) );
NAND2_X2 U8463 ( .A1(n13145), .A2(n13146), .ZN(n5767) );
NAND2_X2 U8464 ( .A1(n17970), .A2(n18957), .ZN(n13146) );
NAND2_X2 U8465 ( .A1(z_out[62]), .A2(n17961), .ZN(n13145) );
NAND2_X2 U8466 ( .A1(n13147), .A2(n13148), .ZN(n5766) );
NAND2_X2 U8467 ( .A1(n17970), .A2(n18958), .ZN(n13148) );
NAND2_X2 U8468 ( .A1(z_out[63]), .A2(n17961), .ZN(n13147) );
NAND2_X2 U8469 ( .A1(n13149), .A2(n13150), .ZN(n5765) );
NAND2_X2 U8470 ( .A1(n17970), .A2(n18959), .ZN(n13150) );
NAND2_X2 U8471 ( .A1(z_out[64]), .A2(n17961), .ZN(n13149) );
NAND2_X2 U8472 ( .A1(n13151), .A2(n13152), .ZN(n5764) );
NAND2_X2 U8473 ( .A1(n17970), .A2(n18960), .ZN(n13152) );
NAND2_X2 U8474 ( .A1(z_out[65]), .A2(n17961), .ZN(n13151) );
NAND2_X2 U8475 ( .A1(n13153), .A2(n13154), .ZN(n5763) );
NAND2_X2 U8476 ( .A1(n17970), .A2(n18961), .ZN(n13154) );
NAND2_X2 U8477 ( .A1(z_out[66]), .A2(n17961), .ZN(n13153) );
NAND2_X2 U8478 ( .A1(n13155), .A2(n13156), .ZN(n5762) );
NAND2_X2 U8479 ( .A1(n17970), .A2(n18962), .ZN(n13156) );
NAND2_X2 U8480 ( .A1(z_out[67]), .A2(n17961), .ZN(n13155) );
NAND2_X2 U8481 ( .A1(n13157), .A2(n13158), .ZN(n5761) );
NAND2_X2 U8482 ( .A1(n17970), .A2(n18963), .ZN(n13158) );
NAND2_X2 U8483 ( .A1(z_out[68]), .A2(n17961), .ZN(n13157) );
NAND2_X2 U8484 ( .A1(n13159), .A2(n13160), .ZN(n5760) );
NAND2_X2 U8485 ( .A1(n17970), .A2(n18964), .ZN(n13160) );
NAND2_X2 U8486 ( .A1(z_out[69]), .A2(n17961), .ZN(n13159) );
NAND2_X2 U8487 ( .A1(n13161), .A2(n13162), .ZN(n5759) );
NAND2_X2 U8488 ( .A1(n17970), .A2(n18965), .ZN(n13162) );
NAND2_X2 U8489 ( .A1(z_out[70]), .A2(n17961), .ZN(n13161) );
NAND2_X2 U8490 ( .A1(n13163), .A2(n13164), .ZN(n5758) );
NAND2_X2 U8491 ( .A1(n17970), .A2(n18966), .ZN(n13164) );
NAND2_X2 U8492 ( .A1(z_out[71]), .A2(n17961), .ZN(n13163) );
NAND2_X2 U8493 ( .A1(n13165), .A2(n13166), .ZN(n5757) );
NAND2_X2 U8494 ( .A1(n17970), .A2(n18967), .ZN(n13166) );
NAND2_X2 U8495 ( .A1(z_out[72]), .A2(n17961), .ZN(n13165) );
NAND2_X2 U8496 ( .A1(n13167), .A2(n13168), .ZN(n5756) );
NAND2_X2 U8497 ( .A1(n17969), .A2(n18968), .ZN(n13168) );
NAND2_X2 U8498 ( .A1(z_out[73]), .A2(n17961), .ZN(n13167) );
NAND2_X2 U8499 ( .A1(n13169), .A2(n13170), .ZN(n5755) );
NAND2_X2 U8500 ( .A1(n17969), .A2(n18969), .ZN(n13170) );
NAND2_X2 U8501 ( .A1(z_out[74]), .A2(n17962), .ZN(n13169) );
NAND2_X2 U8502 ( .A1(n13171), .A2(n13172), .ZN(n5754) );
NAND2_X2 U8503 ( .A1(n17969), .A2(n18970), .ZN(n13172) );
NAND2_X2 U8504 ( .A1(z_out[75]), .A2(n17962), .ZN(n13171) );
NAND2_X2 U8505 ( .A1(n13173), .A2(n13174), .ZN(n5753) );
NAND2_X2 U8506 ( .A1(n17969), .A2(n18971), .ZN(n13174) );
NAND2_X2 U8507 ( .A1(z_out[76]), .A2(n17962), .ZN(n13173) );
NAND2_X2 U8508 ( .A1(n13175), .A2(n13176), .ZN(n5752) );
NAND2_X2 U8509 ( .A1(n17969), .A2(n18972), .ZN(n13176) );
NAND2_X2 U8510 ( .A1(z_out[77]), .A2(n17962), .ZN(n13175) );
NAND2_X2 U8511 ( .A1(n13177), .A2(n13178), .ZN(n5751) );
NAND2_X2 U8512 ( .A1(n17969), .A2(n18973), .ZN(n13178) );
NAND2_X2 U8513 ( .A1(z_out[78]), .A2(n17962), .ZN(n13177) );
NAND2_X2 U8514 ( .A1(n13179), .A2(n13180), .ZN(n5750) );
NAND2_X2 U8515 ( .A1(n17969), .A2(n18974), .ZN(n13180) );
NAND2_X2 U8516 ( .A1(z_out[79]), .A2(n17962), .ZN(n13179) );
NAND2_X2 U8517 ( .A1(n13181), .A2(n13182), .ZN(n5749) );
NAND2_X2 U8518 ( .A1(n17969), .A2(n18975), .ZN(n13182) );
NAND2_X2 U8519 ( .A1(z_out[80]), .A2(n17962), .ZN(n13181) );
NAND2_X2 U8520 ( .A1(n13183), .A2(n13184), .ZN(n5748) );
NAND2_X2 U8521 ( .A1(n17969), .A2(n18976), .ZN(n13184) );
NAND2_X2 U8522 ( .A1(z_out[81]), .A2(n17962), .ZN(n13183) );
NAND2_X2 U8523 ( .A1(n13185), .A2(n13186), .ZN(n5747) );
NAND2_X2 U8524 ( .A1(n17969), .A2(n18977), .ZN(n13186) );
NAND2_X2 U8525 ( .A1(z_out[82]), .A2(n17962), .ZN(n13185) );
NAND2_X2 U8526 ( .A1(n13187), .A2(n13188), .ZN(n5746) );
NAND2_X2 U8527 ( .A1(n17969), .A2(n18978), .ZN(n13188) );
NAND2_X2 U8528 ( .A1(z_out[83]), .A2(n17962), .ZN(n13187) );
NAND2_X2 U8529 ( .A1(n13189), .A2(n13190), .ZN(n5745) );
NAND2_X2 U8530 ( .A1(n17968), .A2(n18979), .ZN(n13190) );
NAND2_X2 U8531 ( .A1(z_out[84]), .A2(n17962), .ZN(n13189) );
NAND2_X2 U8532 ( .A1(n13191), .A2(n13192), .ZN(n5744) );
NAND2_X2 U8533 ( .A1(n17968), .A2(n18980), .ZN(n13192) );
NAND2_X2 U8534 ( .A1(z_out[85]), .A2(n17962), .ZN(n13191) );
NAND2_X2 U8535 ( .A1(n13193), .A2(n13194), .ZN(n5743) );
NAND2_X2 U8536 ( .A1(n17968), .A2(n18981), .ZN(n13194) );
NAND2_X2 U8537 ( .A1(z_out[86]), .A2(n17962), .ZN(n13193) );
NAND2_X2 U8538 ( .A1(n13195), .A2(n13196), .ZN(n5742) );
NAND2_X2 U8539 ( .A1(n17968), .A2(n18982), .ZN(n13196) );
NAND2_X2 U8540 ( .A1(z_out[87]), .A2(n17962), .ZN(n13195) );
NAND2_X2 U8541 ( .A1(n13197), .A2(n13198), .ZN(n5741) );
NAND2_X2 U8542 ( .A1(n17968), .A2(n18983), .ZN(n13198) );
NAND2_X2 U8543 ( .A1(z_out[88]), .A2(n17962), .ZN(n13197) );
NAND2_X2 U8544 ( .A1(n13199), .A2(n13200), .ZN(n5740) );
NAND2_X2 U8545 ( .A1(n17968), .A2(n18984), .ZN(n13200) );
NAND2_X2 U8546 ( .A1(z_out[89]), .A2(n17962), .ZN(n13199) );
NAND2_X2 U8547 ( .A1(n13201), .A2(n13202), .ZN(n5739) );
NAND2_X2 U8548 ( .A1(n17968), .A2(n18985), .ZN(n13202) );
NAND2_X2 U8549 ( .A1(z_out[90]), .A2(n17962), .ZN(n13201) );
NAND2_X2 U8550 ( .A1(n13203), .A2(n13204), .ZN(n5738) );
NAND2_X2 U8551 ( .A1(n17968), .A2(n18986), .ZN(n13204) );
NAND2_X2 U8552 ( .A1(z_out[91]), .A2(n17962), .ZN(n13203) );
NAND2_X2 U8553 ( .A1(n13205), .A2(n13206), .ZN(n5737) );
NAND2_X2 U8554 ( .A1(n17968), .A2(n18987), .ZN(n13206) );
NAND2_X2 U8555 ( .A1(z_out[92]), .A2(n17962), .ZN(n13205) );
NAND2_X2 U8556 ( .A1(n13207), .A2(n13208), .ZN(n5736) );
NAND2_X2 U8557 ( .A1(n17968), .A2(n18988), .ZN(n13208) );
NAND2_X2 U8558 ( .A1(z_out[93]), .A2(n17963), .ZN(n13207) );
NAND2_X2 U8559 ( .A1(n13209), .A2(n13210), .ZN(n5735) );
NAND2_X2 U8560 ( .A1(n17968), .A2(n18989), .ZN(n13210) );
NAND2_X2 U8561 ( .A1(z_out[94]), .A2(n17963), .ZN(n13209) );
NAND2_X2 U8562 ( .A1(n13211), .A2(n13212), .ZN(n5734) );
NAND2_X2 U8563 ( .A1(n17967), .A2(n18990), .ZN(n13212) );
NAND2_X2 U8564 ( .A1(z_out[95]), .A2(n17963), .ZN(n13211) );
NAND2_X2 U8565 ( .A1(n13213), .A2(n13214), .ZN(n5733) );
NAND2_X2 U8566 ( .A1(n17967), .A2(n18991), .ZN(n13214) );
NAND2_X2 U8567 ( .A1(z_out[96]), .A2(n17963), .ZN(n13213) );
NAND2_X2 U8568 ( .A1(n13215), .A2(n13216), .ZN(n5732) );
NAND2_X2 U8569 ( .A1(n17967), .A2(n18992), .ZN(n13216) );
NAND2_X2 U8570 ( .A1(z_out[97]), .A2(n17963), .ZN(n13215) );
NAND2_X2 U8571 ( .A1(n13217), .A2(n13218), .ZN(n5731) );
NAND2_X2 U8572 ( .A1(n17967), .A2(n18993), .ZN(n13218) );
NAND2_X2 U8573 ( .A1(z_out[98]), .A2(n17963), .ZN(n13217) );
NAND2_X2 U8574 ( .A1(n13219), .A2(n13220), .ZN(n5730) );
NAND2_X2 U8575 ( .A1(n17967), .A2(n18994), .ZN(n13220) );
NAND2_X2 U8576 ( .A1(z_out[99]), .A2(n17963), .ZN(n13219) );
NAND2_X2 U8577 ( .A1(n13221), .A2(n13222), .ZN(n5729) );
NAND2_X2 U8578 ( .A1(n17967), .A2(n18995), .ZN(n13222) );
NAND2_X2 U8579 ( .A1(z_out[100]), .A2(n17963), .ZN(n13221) );
NAND2_X2 U8580 ( .A1(n13223), .A2(n13224), .ZN(n5728) );
NAND2_X2 U8581 ( .A1(n17967), .A2(n18996), .ZN(n13224) );
NAND2_X2 U8582 ( .A1(z_out[101]), .A2(n17963), .ZN(n13223) );
NAND2_X2 U8583 ( .A1(n13225), .A2(n13226), .ZN(n5727) );
NAND2_X2 U8584 ( .A1(n17967), .A2(n18997), .ZN(n13226) );
NAND2_X2 U8585 ( .A1(z_out[102]), .A2(n17963), .ZN(n13225) );
NAND2_X2 U8586 ( .A1(n13227), .A2(n13228), .ZN(n5726) );
NAND2_X2 U8587 ( .A1(n17967), .A2(n18998), .ZN(n13228) );
NAND2_X2 U8588 ( .A1(z_out[103]), .A2(n17963), .ZN(n13227) );
NAND2_X2 U8589 ( .A1(n13229), .A2(n13230), .ZN(n5725) );
NAND2_X2 U8590 ( .A1(n17967), .A2(n18999), .ZN(n13230) );
NAND2_X2 U8591 ( .A1(z_out[104]), .A2(n17963), .ZN(n13229) );
NAND2_X2 U8592 ( .A1(n13231), .A2(n13232), .ZN(n5724) );
NAND2_X2 U8593 ( .A1(n17967), .A2(n19000), .ZN(n13232) );
NAND2_X2 U8594 ( .A1(z_out[105]), .A2(n17963), .ZN(n13231) );
NAND2_X2 U8595 ( .A1(n13233), .A2(n13234), .ZN(n5723) );
NAND2_X2 U8596 ( .A1(n17966), .A2(n19001), .ZN(n13234) );
NAND2_X2 U8597 ( .A1(z_out[106]), .A2(n17963), .ZN(n13233) );
NAND2_X2 U8598 ( .A1(n13235), .A2(n13236), .ZN(n5722) );
NAND2_X2 U8599 ( .A1(n17966), .A2(n19002), .ZN(n13236) );
NAND2_X2 U8600 ( .A1(z_out[107]), .A2(n17963), .ZN(n13235) );
NAND2_X2 U8601 ( .A1(n13237), .A2(n13238), .ZN(n5721) );
NAND2_X2 U8602 ( .A1(n17966), .A2(n19003), .ZN(n13238) );
NAND2_X2 U8603 ( .A1(z_out[108]), .A2(n17963), .ZN(n13237) );
NAND2_X2 U8604 ( .A1(n13239), .A2(n13240), .ZN(n5720) );
NAND2_X2 U8605 ( .A1(n17966), .A2(n19004), .ZN(n13240) );
NAND2_X2 U8606 ( .A1(z_out[109]), .A2(n17963), .ZN(n13239) );
NAND2_X2 U8607 ( .A1(n13241), .A2(n13242), .ZN(n5719) );
NAND2_X2 U8608 ( .A1(n17966), .A2(n19005), .ZN(n13242) );
NAND2_X2 U8609 ( .A1(z_out[110]), .A2(n17963), .ZN(n13241) );
NAND2_X2 U8610 ( .A1(n13243), .A2(n13244), .ZN(n5718) );
NAND2_X2 U8611 ( .A1(n17966), .A2(n19006), .ZN(n13244) );
NAND2_X2 U8612 ( .A1(z_out[111]), .A2(n17963), .ZN(n13243) );
NAND2_X2 U8613 ( .A1(n13245), .A2(n13246), .ZN(n5717) );
NAND2_X2 U8614 ( .A1(n17966), .A2(n19007), .ZN(n13246) );
NAND2_X2 U8615 ( .A1(z_out[112]), .A2(n17964), .ZN(n13245) );
NAND2_X2 U8616 ( .A1(n13247), .A2(n13248), .ZN(n5716) );
NAND2_X2 U8617 ( .A1(n17966), .A2(n19008), .ZN(n13248) );
NAND2_X2 U8618 ( .A1(z_out[113]), .A2(n17964), .ZN(n13247) );
NAND2_X2 U8619 ( .A1(n13249), .A2(n13250), .ZN(n5715) );
NAND2_X2 U8620 ( .A1(n17966), .A2(n19009), .ZN(n13250) );
NAND2_X2 U8621 ( .A1(z_out[114]), .A2(n17964), .ZN(n13249) );
NAND2_X2 U8622 ( .A1(n13251), .A2(n13252), .ZN(n5714) );
NAND2_X2 U8623 ( .A1(n17966), .A2(n19010), .ZN(n13252) );
NAND2_X2 U8624 ( .A1(z_out[115]), .A2(n17964), .ZN(n13251) );
NAND2_X2 U8625 ( .A1(n13253), .A2(n13254), .ZN(n5713) );
NAND2_X2 U8626 ( .A1(n17966), .A2(n19011), .ZN(n13254) );
NAND2_X2 U8627 ( .A1(z_out[116]), .A2(n17964), .ZN(n13253) );
NAND2_X2 U8628 ( .A1(n13255), .A2(n13256), .ZN(n5712) );
NAND2_X2 U8629 ( .A1(n17965), .A2(n19012), .ZN(n13256) );
NAND2_X2 U8630 ( .A1(z_out[117]), .A2(n17964), .ZN(n13255) );
NAND2_X2 U8631 ( .A1(n13257), .A2(n13258), .ZN(n5711) );
NAND2_X2 U8632 ( .A1(n17965), .A2(n19013), .ZN(n13258) );
NAND2_X2 U8633 ( .A1(z_out[118]), .A2(n17964), .ZN(n13257) );
NAND2_X2 U8634 ( .A1(n13259), .A2(n13260), .ZN(n5710) );
NAND2_X2 U8635 ( .A1(n17965), .A2(n19014), .ZN(n13260) );
NAND2_X2 U8636 ( .A1(z_out[119]), .A2(n17964), .ZN(n13259) );
NAND2_X2 U8637 ( .A1(n13261), .A2(n13262), .ZN(n5709) );
NAND2_X2 U8638 ( .A1(n17965), .A2(n19015), .ZN(n13262) );
NAND2_X2 U8639 ( .A1(z_out[120]), .A2(n17964), .ZN(n13261) );
NAND2_X2 U8640 ( .A1(n13263), .A2(n13264), .ZN(n5708) );
NAND2_X2 U8641 ( .A1(n17965), .A2(n19016), .ZN(n13264) );
NAND2_X2 U8642 ( .A1(z_out[121]), .A2(n17964), .ZN(n13263) );
NAND2_X2 U8643 ( .A1(n13265), .A2(n13266), .ZN(n5707) );
NAND2_X2 U8644 ( .A1(n17965), .A2(n19017), .ZN(n13266) );
NAND2_X2 U8645 ( .A1(z_out[122]), .A2(n17964), .ZN(n13265) );
NAND2_X2 U8646 ( .A1(n13267), .A2(n13268), .ZN(n5706) );
NAND2_X2 U8647 ( .A1(n17965), .A2(n19018), .ZN(n13268) );
NAND2_X2 U8648 ( .A1(z_out[123]), .A2(n17964), .ZN(n13267) );
NAND2_X2 U8649 ( .A1(n13269), .A2(n13270), .ZN(n5705) );
NAND2_X2 U8650 ( .A1(n17965), .A2(n19019), .ZN(n13270) );
NAND2_X2 U8651 ( .A1(z_out[124]), .A2(n17964), .ZN(n13269) );
NAND2_X2 U8652 ( .A1(n13271), .A2(n13272), .ZN(n5704) );
NAND2_X2 U8653 ( .A1(n17965), .A2(n19020), .ZN(n13272) );
NAND2_X2 U8654 ( .A1(z_out[125]), .A2(n17964), .ZN(n13271) );
NAND2_X2 U8655 ( .A1(n13273), .A2(n13274), .ZN(n5703) );
NAND2_X2 U8656 ( .A1(n17965), .A2(n19021), .ZN(n13274) );
NAND2_X2 U8657 ( .A1(z_out[126]), .A2(n17964), .ZN(n13273) );
NAND2_X2 U8658 ( .A1(n13275), .A2(n13276), .ZN(n5702) );
NAND2_X2 U8659 ( .A1(n17965), .A2(n19022), .ZN(n13276) );
NAND2_X2 U8661 ( .A1(z_out[127]), .A2(n17958), .ZN(n13275) );
NAND4_X2 U8663 ( .A1(n13277), .A2(n13278), .A3(n13279), .A4(n13280), .ZN(n5701) );
NAND2_X2 U8664 ( .A1(n13281), .A2(n17847), .ZN(n13279) );
XNOR2_X2 U8665 ( .A(n17279), .B(z_out[0]), .ZN(n13281) );
NAND2_X2 U8666 ( .A1(n17957), .A2(Out_data[0]), .ZN(n13278) );
NAND2_X2 U8667 ( .A1(n17935), .A2(aes_text_out[0]), .ZN(n13277) );
NAND4_X2 U8668 ( .A1(n13284), .A2(n13285), .A3(n13286), .A4(n13287), .ZN(n5700) );
NAND2_X2 U8669 ( .A1(n13288), .A2(n17847), .ZN(n13286) );
XNOR2_X2 U8670 ( .A(n17277), .B(z_out[1]), .ZN(n13288) );
NAND2_X2 U8671 ( .A1(n17957), .A2(Out_data[1]), .ZN(n13285) );
NAND2_X2 U8672 ( .A1(n17933), .A2(aes_text_out[1]), .ZN(n13284) );
NAND4_X2 U8673 ( .A1(n13289), .A2(n13290), .A3(n13291), .A4(n13292), .ZN(n5699) );
NAND2_X2 U8674 ( .A1(n13293), .A2(n17847), .ZN(n13291) );
XNOR2_X2 U8675 ( .A(n17275), .B(z_out[2]), .ZN(n13293) );
NAND2_X2 U8676 ( .A1(n17957), .A2(Out_data[2]), .ZN(n13290) );
NAND2_X2 U8677 ( .A1(n17934), .A2(aes_text_out[2]), .ZN(n13289) );
NAND4_X2 U8678 ( .A1(n13294), .A2(n13295), .A3(n13296), .A4(n13297), .ZN(n5698) );
NAND2_X2 U8679 ( .A1(n13298), .A2(n17847), .ZN(n13296) );
XNOR2_X2 U8680 ( .A(n17273), .B(z_out[3]), .ZN(n13298) );
NAND2_X2 U8681 ( .A1(n17957), .A2(Out_data[3]), .ZN(n13295) );
NAND2_X2 U8682 ( .A1(n17933), .A2(aes_text_out[3]), .ZN(n13294) );
NAND4_X2 U8683 ( .A1(n13299), .A2(n13300), .A3(n13301), .A4(n13302), .ZN(n5697) );
NAND2_X2 U8684 ( .A1(n13303), .A2(n17847), .ZN(n13301) );
XNOR2_X2 U8685 ( .A(n17271), .B(z_out[4]), .ZN(n13303) );
NAND2_X2 U8686 ( .A1(n17957), .A2(Out_data[4]), .ZN(n13300) );
NAND2_X2 U8687 ( .A1(n17934), .A2(aes_text_out[4]), .ZN(n13299) );
NAND4_X2 U8688 ( .A1(n13304), .A2(n13305), .A3(n13306), .A4(n13307), .ZN(n5696) );
NAND2_X2 U8689 ( .A1(n13308), .A2(n17847), .ZN(n13306) );
XNOR2_X2 U8690 ( .A(n17269), .B(z_out[5]), .ZN(n13308) );
NAND2_X2 U8691 ( .A1(n17957), .A2(Out_data[5]), .ZN(n13305) );
NAND2_X2 U8692 ( .A1(n17934), .A2(aes_text_out[5]), .ZN(n13304) );
NAND4_X2 U8693 ( .A1(n13309), .A2(n13310), .A3(n13311), .A4(n13312), .ZN(n5695) );
NAND2_X2 U8694 ( .A1(n13313), .A2(n17847), .ZN(n13311) );
XNOR2_X2 U8695 ( .A(n17267), .B(z_out[6]), .ZN(n13313) );
NAND2_X2 U8696 ( .A1(n17957), .A2(Out_data[6]), .ZN(n13310) );
NAND2_X2 U8697 ( .A1(n17935), .A2(aes_text_out[6]), .ZN(n13309) );
NAND4_X2 U8698 ( .A1(n13314), .A2(n13315), .A3(n13316), .A4(n13317), .ZN(n5694) );
NAND2_X2 U8699 ( .A1(n13318), .A2(n17847), .ZN(n13316) );
XNOR2_X2 U8700 ( .A(n17265), .B(z_out[7]), .ZN(n13318) );
NAND2_X2 U8701 ( .A1(n17956), .A2(Out_data[7]), .ZN(n13315) );
NAND2_X2 U8702 ( .A1(n17935), .A2(aes_text_out[7]), .ZN(n13314) );
NAND4_X2 U8703 ( .A1(n13319), .A2(n13320), .A3(n13321), .A4(n13322), .ZN(n5693) );
NAND2_X2 U8704 ( .A1(aes_text_out[8]), .A2(n13323), .ZN(n13321) );
NAND2_X2 U8705 ( .A1(n13324), .A2(n17847), .ZN(n13320) );
XNOR2_X2 U8706 ( .A(n17263), .B(z_out[8]), .ZN(n13324) );
NAND2_X2 U8707 ( .A1(n17956), .A2(Out_data[8]), .ZN(n13319) );
NAND4_X2 U8708 ( .A1(n13325), .A2(n13326), .A3(n13327), .A4(n13328), .ZN(n5692) );
NAND2_X2 U8709 ( .A1(aes_text_out[9]), .A2(n13329), .ZN(n13327) );
NAND2_X2 U8710 ( .A1(n13330), .A2(n17847), .ZN(n13326) );
XNOR2_X2 U8711 ( .A(n17261), .B(z_out[9]), .ZN(n13330) );
NAND2_X2 U8712 ( .A1(n17956), .A2(Out_data[9]), .ZN(n13325) );
NAND4_X2 U8713 ( .A1(n13331), .A2(n13332), .A3(n13333), .A4(n13334), .ZN(n5691) );
NAND2_X2 U8714 ( .A1(aes_text_out[10]), .A2(n13335), .ZN(n13333) );
NAND2_X2 U8715 ( .A1(n13336), .A2(n17847), .ZN(n13332) );
XNOR2_X2 U8716 ( .A(n17259), .B(z_out[10]), .ZN(n13336) );
NAND2_X2 U8717 ( .A1(n17956), .A2(Out_data[10]), .ZN(n13331) );
NAND4_X2 U8718 ( .A1(n13337), .A2(n13338), .A3(n13339), .A4(n13340), .ZN(n5690) );
NAND2_X2 U8719 ( .A1(aes_text_out[11]), .A2(n13341), .ZN(n13339) );
NAND2_X2 U8720 ( .A1(n13342), .A2(n17847), .ZN(n13338) );
XNOR2_X2 U8721 ( .A(n17257), .B(z_out[11]), .ZN(n13342) );
NAND2_X2 U8722 ( .A1(n17956), .A2(Out_data[11]), .ZN(n13337) );
NAND4_X2 U8723 ( .A1(n13343), .A2(n13344), .A3(n13345), .A4(n13346), .ZN(n5689) );
NAND2_X2 U8724 ( .A1(aes_text_out[12]), .A2(n13347), .ZN(n13345) );
NAND2_X2 U8725 ( .A1(n13348), .A2(n17847), .ZN(n13344) );
XNOR2_X2 U8726 ( .A(n17255), .B(z_out[12]), .ZN(n13348) );
NAND2_X2 U8727 ( .A1(n17956), .A2(Out_data[12]), .ZN(n13343) );
NAND4_X2 U8728 ( .A1(n13349), .A2(n13350), .A3(n13351), .A4(n13352), .ZN(n5688) );
NAND2_X2 U8729 ( .A1(aes_text_out[13]), .A2(n13353), .ZN(n13351) );
NAND2_X2 U8730 ( .A1(n13354), .A2(n17847), .ZN(n13350) );
XNOR2_X2 U8731 ( .A(n17253), .B(z_out[13]), .ZN(n13354) );
NAND2_X2 U8732 ( .A1(n17956), .A2(Out_data[13]), .ZN(n13349) );
NAND4_X2 U8733 ( .A1(n13355), .A2(n13356), .A3(n13357), .A4(n13358), .ZN(n5687) );
NAND2_X2 U8734 ( .A1(aes_text_out[14]), .A2(n13359), .ZN(n13357) );
NAND2_X2 U8735 ( .A1(n13360), .A2(n17847), .ZN(n13356) );
XNOR2_X2 U8736 ( .A(n17251), .B(z_out[14]), .ZN(n13360) );
NAND2_X2 U8737 ( .A1(n17956), .A2(Out_data[14]), .ZN(n13355) );
NAND4_X2 U8738 ( .A1(n13361), .A2(n13362), .A3(n13363), .A4(n13364), .ZN(n5686) );
NAND2_X2 U8739 ( .A1(aes_text_out[15]), .A2(n13365), .ZN(n13363) );
NAND2_X2 U8740 ( .A1(n13366), .A2(n17846), .ZN(n13362) );
XNOR2_X2 U8741 ( .A(n17249), .B(z_out[15]), .ZN(n13366) );
NAND2_X2 U8742 ( .A1(n17956), .A2(Out_data[15]), .ZN(n13361) );
NAND4_X2 U8743 ( .A1(n13367), .A2(n13368), .A3(n13369), .A4(n13370), .ZN(n5685) );
NAND2_X2 U8744 ( .A1(n13371), .A2(n17846), .ZN(n13369) );
XNOR2_X2 U8745 ( .A(n17247), .B(z_out[16]), .ZN(n13371) );
NAND2_X2 U8746 ( .A1(n17956), .A2(Out_data[16]), .ZN(n13368) );
NAND2_X2 U8747 ( .A1(n13372), .A2(n17936), .ZN(n13367) );
NAND4_X2 U8748 ( .A1(n13373), .A2(n13374), .A3(n13375), .A4(n13376), .ZN(n5684) );
NAND2_X2 U8749 ( .A1(n13377), .A2(n17846), .ZN(n13375) );
XNOR2_X2 U8750 ( .A(n17245), .B(z_out[17]), .ZN(n13377) );
NAND2_X2 U8751 ( .A1(n17956), .A2(Out_data[17]), .ZN(n13374) );
NAND2_X2 U8752 ( .A1(n13378), .A2(n17936), .ZN(n13373) );
NAND4_X2 U8753 ( .A1(n13379), .A2(n13380), .A3(n13381), .A4(n13382), .ZN(n5683) );
NAND2_X2 U8754 ( .A1(n13383), .A2(n17846), .ZN(n13381) );
XNOR2_X2 U8755 ( .A(n17243), .B(z_out[18]), .ZN(n13383) );
NAND2_X2 U8756 ( .A1(n17955), .A2(Out_data[18]), .ZN(n13380) );
NAND2_X2 U8757 ( .A1(n13384), .A2(n17936), .ZN(n13379) );
NAND4_X2 U8758 ( .A1(n13385), .A2(n13386), .A3(n13387), .A4(n13388), .ZN(n5682) );
NAND2_X2 U8759 ( .A1(n13389), .A2(n17846), .ZN(n13387) );
XNOR2_X2 U8760 ( .A(n17241), .B(z_out[19]), .ZN(n13389) );
NAND2_X2 U8761 ( .A1(n17955), .A2(Out_data[19]), .ZN(n13386) );
NAND2_X2 U8762 ( .A1(n13390), .A2(n17936), .ZN(n13385) );
NAND4_X2 U8763 ( .A1(n13391), .A2(n13392), .A3(n13393), .A4(n13394), .ZN(n5681) );
NAND2_X2 U8764 ( .A1(n13395), .A2(n17846), .ZN(n13393) );
XNOR2_X2 U8765 ( .A(n17239), .B(z_out[20]), .ZN(n13395) );
NAND2_X2 U8766 ( .A1(n17955), .A2(Out_data[20]), .ZN(n13392) );
NAND2_X2 U8767 ( .A1(n13396), .A2(n17936), .ZN(n13391) );
NAND4_X2 U8768 ( .A1(n13397), .A2(n13398), .A3(n13399), .A4(n13400), .ZN(n5680) );
NAND2_X2 U8769 ( .A1(n13401), .A2(n17846), .ZN(n13399) );
XNOR2_X2 U8770 ( .A(n17237), .B(z_out[21]), .ZN(n13401) );
NAND2_X2 U8771 ( .A1(n17955), .A2(Out_data[21]), .ZN(n13398) );
NAND2_X2 U8772 ( .A1(n13402), .A2(n17936), .ZN(n13397) );
NAND4_X2 U8773 ( .A1(n13403), .A2(n13404), .A3(n13405), .A4(n13406), .ZN(n5679) );
NAND2_X2 U8774 ( .A1(n13407), .A2(n17846), .ZN(n13405) );
XNOR2_X2 U8775 ( .A(n17235), .B(z_out[22]), .ZN(n13407) );
NAND2_X2 U8776 ( .A1(n17955), .A2(Out_data[22]), .ZN(n13404) );
NAND2_X2 U8777 ( .A1(n13408), .A2(n17936), .ZN(n13403) );
NAND4_X2 U8778 ( .A1(n13409), .A2(n13410), .A3(n13411), .A4(n13412), .ZN(n5678) );
NAND2_X2 U8779 ( .A1(n13413), .A2(n17846), .ZN(n13411) );
XNOR2_X2 U8780 ( .A(n17233), .B(z_out[23]), .ZN(n13413) );
NAND2_X2 U8781 ( .A1(n17955), .A2(Out_data[23]), .ZN(n13410) );
NAND2_X2 U8782 ( .A1(n13414), .A2(n17936), .ZN(n13409) );
NAND4_X2 U8783 ( .A1(n13415), .A2(n13416), .A3(n13417), .A4(n13418), .ZN(n5677) );
NAND2_X2 U8784 ( .A1(n13419), .A2(n17846), .ZN(n13417) );
XNOR2_X2 U8785 ( .A(n17231), .B(z_out[24]), .ZN(n13419) );
NAND2_X2 U8786 ( .A1(n17955), .A2(Out_data[24]), .ZN(n13416) );
NAND2_X2 U8787 ( .A1(n18835), .A2(n17936), .ZN(n13415) );
NAND4_X2 U8788 ( .A1(n13421), .A2(n13422), .A3(n13423), .A4(n13424), .ZN(n5676) );
NAND2_X2 U8789 ( .A1(n13425), .A2(n17846), .ZN(n13423) );
XNOR2_X2 U8790 ( .A(n17229), .B(z_out[25]), .ZN(n13425) );
NAND2_X2 U8791 ( .A1(n17955), .A2(Out_data[25]), .ZN(n13422) );
NAND2_X2 U8792 ( .A1(n18834), .A2(n17936), .ZN(n13421) );
NAND4_X2 U8793 ( .A1(n13427), .A2(n13428), .A3(n13429), .A4(n13430), .ZN(n5675) );
NAND2_X2 U8794 ( .A1(n13431), .A2(n17846), .ZN(n13429) );
XNOR2_X2 U8795 ( .A(n17227), .B(z_out[26]), .ZN(n13431) );
NAND2_X2 U8796 ( .A1(n17955), .A2(Out_data[26]), .ZN(n13428) );
NAND2_X2 U8797 ( .A1(n18833), .A2(n17936), .ZN(n13427) );
NAND4_X2 U8798 ( .A1(n13433), .A2(n13434), .A3(n13435), .A4(n13436), .ZN(n5674) );
NAND2_X2 U8799 ( .A1(n13437), .A2(n17846), .ZN(n13435) );
XNOR2_X2 U8800 ( .A(n17225), .B(z_out[27]), .ZN(n13437) );
NAND2_X2 U8801 ( .A1(n17955), .A2(Out_data[27]), .ZN(n13434) );
NAND2_X2 U8802 ( .A1(n18832), .A2(n17937), .ZN(n13433) );
NAND4_X2 U8803 ( .A1(n13439), .A2(n13440), .A3(n13441), .A4(n13442), .ZN(n5673) );
NAND2_X2 U8804 ( .A1(n13443), .A2(n17846), .ZN(n13441) );
XNOR2_X2 U8805 ( .A(n17223), .B(z_out[28]), .ZN(n13443) );
NAND2_X2 U8806 ( .A1(n17955), .A2(Out_data[28]), .ZN(n13440) );
NAND2_X2 U8807 ( .A1(n18831), .A2(n17937), .ZN(n13439) );
NAND4_X2 U8808 ( .A1(n13445), .A2(n13446), .A3(n13447), .A4(n13448), .ZN(n5672) );
NAND2_X2 U8809 ( .A1(n13449), .A2(n17846), .ZN(n13447) );
XNOR2_X2 U8810 ( .A(n17221), .B(z_out[29]), .ZN(n13449) );
NAND2_X2 U8811 ( .A1(n17954), .A2(Out_data[29]), .ZN(n13446) );
NAND2_X2 U8812 ( .A1(n18830), .A2(n17937), .ZN(n13445) );
NAND4_X2 U8813 ( .A1(n13451), .A2(n13452), .A3(n13453), .A4(n13454), .ZN(n5671) );
NAND2_X2 U8814 ( .A1(n13455), .A2(n17846), .ZN(n13453) );
XNOR2_X2 U8815 ( .A(n17219), .B(z_out[30]), .ZN(n13455) );
NAND2_X2 U8816 ( .A1(n17954), .A2(Out_data[30]), .ZN(n13452) );
NAND2_X2 U8817 ( .A1(n18829), .A2(n17937), .ZN(n13451) );
NAND4_X2 U8818 ( .A1(n13457), .A2(n13458), .A3(n13459), .A4(n13460), .ZN(n5670) );
NAND2_X2 U8819 ( .A1(n13461), .A2(n17846), .ZN(n13459) );
XNOR2_X2 U8820 ( .A(n17217), .B(z_out[31]), .ZN(n13461) );
NAND2_X2 U8821 ( .A1(n17954), .A2(Out_data[31]), .ZN(n13458) );
NAND2_X2 U8822 ( .A1(n18828), .A2(n17937), .ZN(n13457) );
NAND4_X2 U8823 ( .A1(n13463), .A2(n13464), .A3(n13465), .A4(n13466), .ZN(n5669) );
NAND2_X2 U8824 ( .A1(n13467), .A2(n17846), .ZN(n13465) );
XNOR2_X2 U8825 ( .A(n17215), .B(z_out[32]), .ZN(n13467) );
NAND2_X2 U8826 ( .A1(n17954), .A2(Out_data[32]), .ZN(n13464) );
NAND2_X2 U8827 ( .A1(n13468), .A2(n17937), .ZN(n13463) );
NAND4_X2 U8828 ( .A1(n13469), .A2(n13470), .A3(n13471), .A4(n13472), .ZN(n5668) );
NAND2_X2 U8829 ( .A1(n13473), .A2(n17846), .ZN(n13471) );
XNOR2_X2 U8830 ( .A(n17213), .B(z_out[33]), .ZN(n13473) );
NAND2_X2 U8831 ( .A1(n17954), .A2(Out_data[33]), .ZN(n13470) );
NAND2_X2 U8832 ( .A1(n13474), .A2(n17937), .ZN(n13469) );
NAND4_X2 U8833 ( .A1(n13475), .A2(n13476), .A3(n13477), .A4(n13478), .ZN(n5667) );
NAND2_X2 U8834 ( .A1(n13479), .A2(n17845), .ZN(n13477) );
XNOR2_X2 U8835 ( .A(n17211), .B(z_out[34]), .ZN(n13479) );
NAND2_X2 U8836 ( .A1(n17954), .A2(Out_data[34]), .ZN(n13476) );
NAND2_X2 U8837 ( .A1(n13480), .A2(n17937), .ZN(n13475) );
NAND4_X2 U8838 ( .A1(n13481), .A2(n13482), .A3(n13483), .A4(n13484), .ZN(n5666) );
NAND2_X2 U8839 ( .A1(n13485), .A2(n17845), .ZN(n13483) );
XNOR2_X2 U8840 ( .A(n17209), .B(z_out[35]), .ZN(n13485) );
NAND2_X2 U8841 ( .A1(n17954), .A2(Out_data[35]), .ZN(n13482) );
NAND2_X2 U8842 ( .A1(n13486), .A2(n17937), .ZN(n13481) );
NAND4_X2 U8843 ( .A1(n13487), .A2(n13488), .A3(n13489), .A4(n13490), .ZN(n5665) );
NAND2_X2 U8844 ( .A1(n13491), .A2(n17845), .ZN(n13489) );
XNOR2_X2 U8845 ( .A(n17207), .B(z_out[36]), .ZN(n13491) );
NAND2_X2 U8846 ( .A1(n17954), .A2(Out_data[36]), .ZN(n13488) );
NAND2_X2 U8847 ( .A1(n13492), .A2(n17937), .ZN(n13487) );
NAND4_X2 U8848 ( .A1(n13493), .A2(n13494), .A3(n13495), .A4(n13496), .ZN(n5664) );
NAND2_X2 U8849 ( .A1(n13497), .A2(n17845), .ZN(n13495) );
XNOR2_X2 U8850 ( .A(n17205), .B(z_out[37]), .ZN(n13497) );
NAND2_X2 U8851 ( .A1(n17954), .A2(Out_data[37]), .ZN(n13494) );
NAND2_X2 U8852 ( .A1(n13498), .A2(n17937), .ZN(n13493) );
NAND4_X2 U8853 ( .A1(n13499), .A2(n13500), .A3(n13501), .A4(n13502), .ZN(n5663) );
NAND2_X2 U8854 ( .A1(n13503), .A2(n17845), .ZN(n13501) );
XNOR2_X2 U8855 ( .A(n17203), .B(z_out[38]), .ZN(n13503) );
NAND2_X2 U8856 ( .A1(n17954), .A2(Out_data[38]), .ZN(n13500) );
NAND2_X2 U8857 ( .A1(n13504), .A2(n17937), .ZN(n13499) );
NAND4_X2 U8858 ( .A1(n13505), .A2(n13506), .A3(n13507), .A4(n13508), .ZN(n5662) );
NAND2_X2 U8859 ( .A1(n13509), .A2(n17845), .ZN(n13507) );
XNOR2_X2 U8860 ( .A(n17201), .B(z_out[39]), .ZN(n13509) );
NAND2_X2 U8861 ( .A1(n17954), .A2(Out_data[39]), .ZN(n13506) );
NAND2_X2 U8862 ( .A1(n13510), .A2(n17938), .ZN(n13505) );
NAND4_X2 U8863 ( .A1(n13511), .A2(n13512), .A3(n13513), .A4(n13514), .ZN(n5661) );
NAND2_X2 U8864 ( .A1(n13515), .A2(n17845), .ZN(n13513) );
XNOR2_X2 U8865 ( .A(n17199), .B(z_out[40]), .ZN(n13515) );
NAND2_X2 U8866 ( .A1(n17953), .A2(Out_data[40]), .ZN(n13512) );
NAND2_X2 U8867 ( .A1(n18827), .A2(n17938), .ZN(n13511) );
NAND4_X2 U8868 ( .A1(n13517), .A2(n13518), .A3(n13519), .A4(n13520), .ZN(n5660) );
NAND2_X2 U8869 ( .A1(n13521), .A2(n17845), .ZN(n13519) );
XNOR2_X2 U8870 ( .A(n17197), .B(z_out[41]), .ZN(n13521) );
NAND2_X2 U8871 ( .A1(n17953), .A2(Out_data[41]), .ZN(n13518) );
NAND2_X2 U8872 ( .A1(n18826), .A2(n17938), .ZN(n13517) );
NAND4_X2 U8873 ( .A1(n13523), .A2(n13524), .A3(n13525), .A4(n13526), .ZN(n5659) );
NAND2_X2 U8874 ( .A1(n13527), .A2(n17845), .ZN(n13525) );
XNOR2_X2 U8875 ( .A(n17195), .B(z_out[42]), .ZN(n13527) );
NAND2_X2 U8876 ( .A1(n17953), .A2(Out_data[42]), .ZN(n13524) );
NAND2_X2 U8877 ( .A1(n18825), .A2(n17938), .ZN(n13523) );
NAND4_X2 U8878 ( .A1(n13529), .A2(n13530), .A3(n13531), .A4(n13532), .ZN(n5658) );
NAND2_X2 U8879 ( .A1(n13533), .A2(n17845), .ZN(n13531) );
XNOR2_X2 U8880 ( .A(n17193), .B(z_out[43]), .ZN(n13533) );
NAND2_X2 U8881 ( .A1(n17953), .A2(Out_data[43]), .ZN(n13530) );
NAND2_X2 U8882 ( .A1(n18824), .A2(n17938), .ZN(n13529) );
NAND4_X2 U8883 ( .A1(n13535), .A2(n13536), .A3(n13537), .A4(n13538), .ZN(n5657) );
NAND2_X2 U8884 ( .A1(n13539), .A2(n17845), .ZN(n13537) );
XNOR2_X2 U8885 ( .A(n17191), .B(z_out[44]), .ZN(n13539) );
NAND2_X2 U8886 ( .A1(n17953), .A2(Out_data[44]), .ZN(n13536) );
NAND2_X2 U8887 ( .A1(n18823), .A2(n17940), .ZN(n13535) );
NAND4_X2 U8888 ( .A1(n13541), .A2(n13542), .A3(n13543), .A4(n13544), .ZN(n5656) );
NAND2_X2 U8889 ( .A1(n13545), .A2(n17845), .ZN(n13543) );
XNOR2_X2 U8890 ( .A(n17189), .B(z_out[45]), .ZN(n13545) );
NAND2_X2 U8891 ( .A1(n17953), .A2(Out_data[45]), .ZN(n13542) );
NAND2_X2 U8892 ( .A1(n18822), .A2(n17938), .ZN(n13541) );
NAND4_X2 U8893 ( .A1(n13547), .A2(n13548), .A3(n13549), .A4(n13550), .ZN(n5655) );
NAND2_X2 U8894 ( .A1(n13551), .A2(n17845), .ZN(n13549) );
XNOR2_X2 U8895 ( .A(n17187), .B(z_out[46]), .ZN(n13551) );
NAND2_X2 U8896 ( .A1(n17953), .A2(Out_data[46]), .ZN(n13548) );
NAND2_X2 U8897 ( .A1(n18821), .A2(n17938), .ZN(n13547) );
NAND4_X2 U8898 ( .A1(n13553), .A2(n13554), .A3(n13555), .A4(n13556), .ZN(n5654) );
NAND2_X2 U8899 ( .A1(n13557), .A2(n17845), .ZN(n13555) );
XNOR2_X2 U8900 ( .A(n17185), .B(z_out[47]), .ZN(n13557) );
NAND2_X2 U8901 ( .A1(n17953), .A2(Out_data[47]), .ZN(n13554) );
NAND2_X2 U8902 ( .A1(n18820), .A2(n17938), .ZN(n13553) );
NAND4_X2 U8903 ( .A1(n13559), .A2(n13560), .A3(n13561), .A4(n13562), .ZN(n5653) );
NAND2_X2 U8904 ( .A1(n13563), .A2(n17845), .ZN(n13561) );
XNOR2_X2 U8905 ( .A(n17183), .B(z_out[48]), .ZN(n13563) );
NAND2_X2 U8906 ( .A1(n17953), .A2(Out_data[48]), .ZN(n13560) );
NAND2_X2 U8907 ( .A1(n13564), .A2(n17938), .ZN(n13559) );
NAND4_X2 U8908 ( .A1(n13565), .A2(n13566), .A3(n13567), .A4(n13568), .ZN(n5652) );
NAND2_X2 U8909 ( .A1(n13569), .A2(n17845), .ZN(n13567) );
XNOR2_X2 U8910 ( .A(n17181), .B(z_out[49]), .ZN(n13569) );
NAND2_X2 U8911 ( .A1(n17953), .A2(Out_data[49]), .ZN(n13566) );
NAND2_X2 U8912 ( .A1(n13570), .A2(n17938), .ZN(n13565) );
NAND4_X2 U8913 ( .A1(n13571), .A2(n13572), .A3(n13573), .A4(n13574), .ZN(n5651) );
NAND2_X2 U8914 ( .A1(n13575), .A2(n17845), .ZN(n13573) );
XNOR2_X2 U8915 ( .A(n17179), .B(z_out[50]), .ZN(n13575) );
NAND2_X2 U8916 ( .A1(n17953), .A2(Out_data[50]), .ZN(n13572) );
NAND2_X2 U8917 ( .A1(n13576), .A2(n17938), .ZN(n13571) );
NAND4_X2 U8918 ( .A1(n13577), .A2(n13578), .A3(n13579), .A4(n13580), .ZN(n5650) );
NAND2_X2 U8919 ( .A1(n13581), .A2(n17845), .ZN(n13579) );
XNOR2_X2 U8920 ( .A(n17177), .B(z_out[51]), .ZN(n13581) );
NAND2_X2 U8921 ( .A1(n17952), .A2(Out_data[51]), .ZN(n13578) );
NAND2_X2 U8922 ( .A1(n13582), .A2(n17938), .ZN(n13577) );
NAND4_X2 U8923 ( .A1(n13583), .A2(n13584), .A3(n13585), .A4(n13586), .ZN(n5649) );
NAND2_X2 U8924 ( .A1(n13587), .A2(n17845), .ZN(n13585) );
XNOR2_X2 U8925 ( .A(n17175), .B(z_out[52]), .ZN(n13587) );
NAND2_X2 U8926 ( .A1(n17952), .A2(Out_data[52]), .ZN(n13584) );
NAND2_X2 U8927 ( .A1(n13588), .A2(n17939), .ZN(n13583) );
NAND4_X2 U8928 ( .A1(n13589), .A2(n13590), .A3(n13591), .A4(n13592), .ZN(n5648) );
NAND2_X2 U8929 ( .A1(n13593), .A2(n17844), .ZN(n13591) );
XNOR2_X2 U8930 ( .A(n17173), .B(z_out[53]), .ZN(n13593) );
NAND2_X2 U8931 ( .A1(n17952), .A2(Out_data[53]), .ZN(n13590) );
NAND2_X2 U8932 ( .A1(n13594), .A2(n17939), .ZN(n13589) );
NAND4_X2 U8933 ( .A1(n13595), .A2(n13596), .A3(n13597), .A4(n13598), .ZN(n5647) );
NAND2_X2 U8934 ( .A1(n13599), .A2(n17844), .ZN(n13597) );
XNOR2_X2 U8935 ( .A(n17171), .B(z_out[54]), .ZN(n13599) );
NAND2_X2 U8936 ( .A1(n17952), .A2(Out_data[54]), .ZN(n13596) );
NAND2_X2 U8937 ( .A1(n13600), .A2(n17939), .ZN(n13595) );
NAND4_X2 U8938 ( .A1(n13601), .A2(n13602), .A3(n13603), .A4(n13604), .ZN(n5646) );
NAND2_X2 U8939 ( .A1(n13605), .A2(n17844), .ZN(n13603) );
XNOR2_X2 U8940 ( .A(n17169), .B(z_out[55]), .ZN(n13605) );
NAND2_X2 U8941 ( .A1(n17952), .A2(Out_data[55]), .ZN(n13602) );
NAND2_X2 U8942 ( .A1(n13606), .A2(n17939), .ZN(n13601) );
NAND4_X2 U8943 ( .A1(n13607), .A2(n13608), .A3(n13609), .A4(n13610), .ZN(n5645) );
NAND2_X2 U8944 ( .A1(n13611), .A2(n17844), .ZN(n13609) );
XNOR2_X2 U8945 ( .A(n17167), .B(z_out[56]), .ZN(n13611) );
NAND2_X2 U8946 ( .A1(n17952), .A2(Out_data[56]), .ZN(n13608) );
NAND2_X2 U8947 ( .A1(n18819), .A2(n17939), .ZN(n13607) );
NAND4_X2 U8948 ( .A1(n13613), .A2(n13614), .A3(n13615), .A4(n13616), .ZN(n5644) );
NAND2_X2 U8949 ( .A1(n13617), .A2(n17844), .ZN(n13615) );
XNOR2_X2 U8950 ( .A(n17165), .B(z_out[57]), .ZN(n13617) );
NAND2_X2 U8951 ( .A1(n17952), .A2(Out_data[57]), .ZN(n13614) );
NAND2_X2 U8952 ( .A1(n18818), .A2(n17939), .ZN(n13613) );
NAND4_X2 U8953 ( .A1(n13619), .A2(n13620), .A3(n13621), .A4(n13622), .ZN(n5643) );
NAND2_X2 U8954 ( .A1(n13623), .A2(n17844), .ZN(n13621) );
XNOR2_X2 U8955 ( .A(n17163), .B(z_out[58]), .ZN(n13623) );
NAND2_X2 U8956 ( .A1(n17952), .A2(Out_data[58]), .ZN(n13620) );
NAND2_X2 U8957 ( .A1(n18817), .A2(n17939), .ZN(n13619) );
NAND4_X2 U8958 ( .A1(n13625), .A2(n13626), .A3(n13627), .A4(n13628), .ZN(n5642) );
NAND2_X2 U8959 ( .A1(n13629), .A2(n17844), .ZN(n13627) );
XNOR2_X2 U8960 ( .A(n17161), .B(z_out[59]), .ZN(n13629) );
NAND2_X2 U8961 ( .A1(n17952), .A2(Out_data[59]), .ZN(n13626) );
NAND2_X2 U8962 ( .A1(n18816), .A2(n17939), .ZN(n13625) );
NAND4_X2 U8963 ( .A1(n13631), .A2(n13632), .A3(n13633), .A4(n13634), .ZN(n5641) );
NAND2_X2 U8964 ( .A1(n13635), .A2(n17844), .ZN(n13633) );
XNOR2_X2 U8965 ( .A(n17159), .B(z_out[60]), .ZN(n13635) );
NAND2_X2 U8966 ( .A1(n17952), .A2(Out_data[60]), .ZN(n13632) );
NAND2_X2 U8967 ( .A1(n18815), .A2(n17939), .ZN(n13631) );
NAND4_X2 U8968 ( .A1(n13637), .A2(n13638), .A3(n13639), .A4(n13640), .ZN(n5640) );
NAND2_X2 U8969 ( .A1(n13641), .A2(n17844), .ZN(n13639) );
XNOR2_X2 U8970 ( .A(n17157), .B(z_out[61]), .ZN(n13641) );
NAND2_X2 U8971 ( .A1(n17952), .A2(Out_data[61]), .ZN(n13638) );
NAND2_X2 U8972 ( .A1(n18814), .A2(n17939), .ZN(n13637) );
NAND4_X2 U8973 ( .A1(n13643), .A2(n13644), .A3(n13645), .A4(n13646), .ZN(n5639) );
NAND2_X2 U8974 ( .A1(n13647), .A2(n17844), .ZN(n13645) );
XNOR2_X2 U8975 ( .A(n17155), .B(z_out[62]), .ZN(n13647) );
NAND2_X2 U8976 ( .A1(n17951), .A2(Out_data[62]), .ZN(n13644) );
NAND2_X2 U8977 ( .A1(n18813), .A2(n17939), .ZN(n13643) );
NAND4_X2 U8978 ( .A1(n13649), .A2(n13650), .A3(n13651), .A4(n13652), .ZN(n5638) );
NAND2_X2 U8979 ( .A1(n13653), .A2(n17844), .ZN(n13651) );
XNOR2_X2 U8980 ( .A(n17153), .B(z_out[63]), .ZN(n13653) );
NAND2_X2 U8981 ( .A1(n17951), .A2(Out_data[63]), .ZN(n13650) );
NAND2_X2 U8982 ( .A1(n18812), .A2(n17939), .ZN(n13649) );
NAND4_X2 U8983 ( .A1(n13655), .A2(n13656), .A3(n13657), .A4(n13658), .ZN(n5637) );
NAND2_X2 U8984 ( .A1(n13659), .A2(n17844), .ZN(n13658) );
XNOR2_X2 U8985 ( .A(n17151), .B(z_out[64]), .ZN(n13659) );
NAND2_X2 U8986 ( .A1(n17951), .A2(Out_data[64]), .ZN(n13657) );
NAND2_X2 U8988 ( .A1(n18811), .A2(n17940), .ZN(n13655) );
NAND4_X2 U8989 ( .A1(n13663), .A2(n13664), .A3(n13665), .A4(n13666), .ZN(n5636) );
NAND2_X2 U8990 ( .A1(n13667), .A2(n17844), .ZN(n13666) );
XNOR2_X2 U8991 ( .A(n17149), .B(z_out[65]), .ZN(n13667) );
NAND2_X2 U8992 ( .A1(n17951), .A2(Out_data[65]), .ZN(n13665) );
NAND2_X2 U8993 ( .A1(n17930), .A2(n13668), .ZN(n13664) );
NAND2_X2 U8994 ( .A1(n18810), .A2(n17940), .ZN(n13663) );
NAND4_X2 U8995 ( .A1(n13670), .A2(n13671), .A3(n13672), .A4(n13673), .ZN(n5635) );
NAND2_X2 U8996 ( .A1(n13674), .A2(n17844), .ZN(n13673) );
XNOR2_X2 U8997 ( .A(n17147), .B(z_out[66]), .ZN(n13674) );
NAND2_X2 U8998 ( .A1(n17951), .A2(Out_data[66]), .ZN(n13672) );
NAND2_X2 U9000 ( .A1(n18809), .A2(n17940), .ZN(n13670) );
NAND4_X2 U9001 ( .A1(n13677), .A2(n13678), .A3(n13679), .A4(n13680), .ZN(n5634) );
NAND2_X2 U9002 ( .A1(n13681), .A2(n17844), .ZN(n13679) );
XNOR2_X2 U9003 ( .A(n17145), .B(z_out[67]), .ZN(n13681) );
NAND2_X2 U9004 ( .A1(n17951), .A2(Out_data[67]), .ZN(n13678) );
NAND2_X2 U9005 ( .A1(n18808), .A2(n17940), .ZN(n13677) );
NAND4_X2 U9006 ( .A1(n13683), .A2(n13684), .A3(n13685), .A4(n13686), .ZN(n5633) );
NAND2_X2 U9007 ( .A1(n13687), .A2(n17844), .ZN(n13685) );
XNOR2_X2 U9008 ( .A(n17143), .B(z_out[68]), .ZN(n13687) );
NAND2_X2 U9009 ( .A1(n17951), .A2(Out_data[68]), .ZN(n13684) );
NAND2_X2 U9010 ( .A1(n18807), .A2(n17940), .ZN(n13683) );
NAND4_X2 U9011 ( .A1(n13689), .A2(n13690), .A3(n13691), .A4(n13692), .ZN(n5632) );
NAND2_X2 U9012 ( .A1(n13693), .A2(n17844), .ZN(n13691) );
XNOR2_X2 U9013 ( .A(n17141), .B(z_out[69]), .ZN(n13693) );
NAND2_X2 U9014 ( .A1(n17951), .A2(Out_data[69]), .ZN(n13690) );
NAND2_X2 U9015 ( .A1(n18806), .A2(n17940), .ZN(n13689) );
NAND4_X2 U9016 ( .A1(n13695), .A2(n13696), .A3(n13697), .A4(n13698), .ZN(n5631) );
NAND2_X2 U9017 ( .A1(n13699), .A2(n17844), .ZN(n13697) );
XNOR2_X2 U9018 ( .A(n17139), .B(z_out[70]), .ZN(n13699) );
NAND2_X2 U9019 ( .A1(n17951), .A2(Out_data[70]), .ZN(n13696) );
NAND2_X2 U9020 ( .A1(n18805), .A2(n17940), .ZN(n13695) );
NAND4_X2 U9021 ( .A1(n13701), .A2(n13702), .A3(n13703), .A4(n13704), .ZN(n5630) );
NAND2_X2 U9022 ( .A1(n13705), .A2(n17844), .ZN(n13703) );
XNOR2_X2 U9023 ( .A(n17137), .B(z_out[71]), .ZN(n13705) );
NAND2_X2 U9024 ( .A1(n17951), .A2(Out_data[71]), .ZN(n13702) );
NAND2_X2 U9025 ( .A1(n18804), .A2(n17940), .ZN(n13701) );
NAND4_X2 U9026 ( .A1(n13707), .A2(n13708), .A3(n13709), .A4(n13710), .ZN(n5629) );
NAND2_X2 U9027 ( .A1(n13711), .A2(n17843), .ZN(n13709) );
XNOR2_X2 U9028 ( .A(n17135), .B(z_out[72]), .ZN(n13711) );
NAND2_X2 U9029 ( .A1(n17951), .A2(Out_data[72]), .ZN(n13708) );
NAND2_X2 U9030 ( .A1(n18803), .A2(n17940), .ZN(n13707) );
NAND4_X2 U9031 ( .A1(n13713), .A2(n13714), .A3(n13715), .A4(n13716), .ZN(n5628) );
NAND2_X2 U9032 ( .A1(n13717), .A2(n17843), .ZN(n13715) );
XNOR2_X2 U9033 ( .A(n17133), .B(z_out[73]), .ZN(n13717) );
NAND2_X2 U9034 ( .A1(n17950), .A2(Out_data[73]), .ZN(n13714) );
NAND2_X2 U9035 ( .A1(n18802), .A2(n17940), .ZN(n13713) );
NAND4_X2 U9036 ( .A1(n13719), .A2(n13720), .A3(n13721), .A4(n13722), .ZN(n5627) );
NAND2_X2 U9037 ( .A1(n13723), .A2(n17843), .ZN(n13721) );
XNOR2_X2 U9038 ( .A(n17131), .B(z_out[74]), .ZN(n13723) );
NAND2_X2 U9039 ( .A1(n17950), .A2(Out_data[74]), .ZN(n13720) );
NAND2_X2 U9040 ( .A1(n18801), .A2(n17940), .ZN(n13719) );
NAND4_X2 U9041 ( .A1(n13725), .A2(n13726), .A3(n13727), .A4(n13728), .ZN(n5626) );
NAND2_X2 U9042 ( .A1(n13729), .A2(n17843), .ZN(n13727) );
XNOR2_X2 U9043 ( .A(n17129), .B(z_out[75]), .ZN(n13729) );
NAND2_X2 U9044 ( .A1(n17950), .A2(Out_data[75]), .ZN(n13726) );
NAND2_X2 U9045 ( .A1(n18800), .A2(n17941), .ZN(n13725) );
NAND4_X2 U9046 ( .A1(n13731), .A2(n13732), .A3(n13733), .A4(n13734), .ZN(n5625) );
NAND2_X2 U9047 ( .A1(n13735), .A2(n17843), .ZN(n13733) );
XNOR2_X2 U9048 ( .A(n17127), .B(z_out[76]), .ZN(n13735) );
NAND2_X2 U9049 ( .A1(n17950), .A2(Out_data[76]), .ZN(n13732) );
NAND2_X2 U9050 ( .A1(n18799), .A2(n17941), .ZN(n13731) );
NAND4_X2 U9051 ( .A1(n13737), .A2(n13738), .A3(n13739), .A4(n13740), .ZN(n5624) );
NAND2_X2 U9052 ( .A1(n13741), .A2(n17843), .ZN(n13739) );
XNOR2_X2 U9053 ( .A(n17125), .B(z_out[77]), .ZN(n13741) );
NAND2_X2 U9054 ( .A1(n17950), .A2(Out_data[77]), .ZN(n13738) );
NAND2_X2 U9055 ( .A1(n18798), .A2(n17941), .ZN(n13737) );
NAND4_X2 U9056 ( .A1(n13743), .A2(n13744), .A3(n13745), .A4(n13746), .ZN(n5623) );
NAND2_X2 U9057 ( .A1(n13747), .A2(n17843), .ZN(n13745) );
XNOR2_X2 U9058 ( .A(n17123), .B(z_out[78]), .ZN(n13747) );
NAND2_X2 U9059 ( .A1(n17950), .A2(Out_data[78]), .ZN(n13744) );
NAND2_X2 U9060 ( .A1(n18797), .A2(n17941), .ZN(n13743) );
NAND4_X2 U9061 ( .A1(n13749), .A2(n13750), .A3(n13751), .A4(n13752), .ZN(n5622) );
NAND2_X2 U9062 ( .A1(n13753), .A2(n17843), .ZN(n13751) );
XNOR2_X2 U9063 ( .A(n17121), .B(z_out[79]), .ZN(n13753) );
NAND2_X2 U9064 ( .A1(n17950), .A2(Out_data[79]), .ZN(n13750) );
NAND2_X2 U9065 ( .A1(n18796), .A2(n17941), .ZN(n13749) );
NAND4_X2 U9066 ( .A1(n13755), .A2(n13756), .A3(n13757), .A4(n13758), .ZN(n5621) );
NAND2_X2 U9067 ( .A1(n13759), .A2(n17843), .ZN(n13757) );
XNOR2_X2 U9068 ( .A(n17119), .B(z_out[80]), .ZN(n13759) );
NAND2_X2 U9069 ( .A1(n17950), .A2(Out_data[80]), .ZN(n13756) );
NAND2_X2 U9070 ( .A1(n18795), .A2(n17941), .ZN(n13755) );
NAND4_X2 U9071 ( .A1(n13761), .A2(n13762), .A3(n13763), .A4(n13764), .ZN(n5620) );
NAND2_X2 U9072 ( .A1(n13765), .A2(n17843), .ZN(n13763) );
XNOR2_X2 U9073 ( .A(n17117), .B(z_out[81]), .ZN(n13765) );
NAND2_X2 U9074 ( .A1(n17950), .A2(Out_data[81]), .ZN(n13762) );
NAND2_X2 U9075 ( .A1(n18794), .A2(n17941), .ZN(n13761) );
NAND4_X2 U9076 ( .A1(n13767), .A2(n13768), .A3(n13769), .A4(n13770), .ZN(n5619) );
NAND2_X2 U9077 ( .A1(n13771), .A2(n17843), .ZN(n13769) );
XNOR2_X2 U9078 ( .A(n17115), .B(z_out[82]), .ZN(n13771) );
NAND2_X2 U9079 ( .A1(n17950), .A2(Out_data[82]), .ZN(n13768) );
NAND2_X2 U9080 ( .A1(n18793), .A2(n17941), .ZN(n13767) );
NAND4_X2 U9081 ( .A1(n13773), .A2(n13774), .A3(n13775), .A4(n13776), .ZN(n5618) );
NAND2_X2 U9082 ( .A1(n13777), .A2(n17843), .ZN(n13775) );
XNOR2_X2 U9083 ( .A(n17113), .B(z_out[83]), .ZN(n13777) );
NAND2_X2 U9084 ( .A1(n17950), .A2(Out_data[83]), .ZN(n13774) );
NAND2_X2 U9085 ( .A1(n18792), .A2(n17941), .ZN(n13773) );
NAND4_X2 U9086 ( .A1(n13779), .A2(n13780), .A3(n13781), .A4(n13782), .ZN(n5617) );
NAND2_X2 U9087 ( .A1(n13783), .A2(n17843), .ZN(n13781) );
XNOR2_X2 U9088 ( .A(n17111), .B(z_out[84]), .ZN(n13783) );
NAND2_X2 U9089 ( .A1(n17949), .A2(Out_data[84]), .ZN(n13780) );
NAND2_X2 U9090 ( .A1(n18791), .A2(n17941), .ZN(n13779) );
NAND4_X2 U9091 ( .A1(n13785), .A2(n13786), .A3(n13787), .A4(n13788), .ZN(n5616) );
NAND2_X2 U9092 ( .A1(n13789), .A2(n17843), .ZN(n13787) );
XNOR2_X2 U9093 ( .A(n17109), .B(z_out[85]), .ZN(n13789) );
NAND2_X2 U9094 ( .A1(n17949), .A2(Out_data[85]), .ZN(n13786) );
NAND2_X2 U9095 ( .A1(n18790), .A2(n17941), .ZN(n13785) );
NAND4_X2 U9096 ( .A1(n13791), .A2(n13792), .A3(n13793), .A4(n13794), .ZN(n5615) );
NAND2_X2 U9097 ( .A1(n13795), .A2(n17843), .ZN(n13793) );
XNOR2_X2 U9098 ( .A(n17107), .B(z_out[86]), .ZN(n13795) );
NAND2_X2 U9099 ( .A1(n17949), .A2(Out_data[86]), .ZN(n13792) );
NAND2_X2 U9100 ( .A1(n18789), .A2(n17941), .ZN(n13791) );
NAND4_X2 U9101 ( .A1(n13797), .A2(n13798), .A3(n13799), .A4(n13800), .ZN(n5614) );
NAND2_X2 U9102 ( .A1(n13801), .A2(n17843), .ZN(n13799) );
XNOR2_X2 U9103 ( .A(n17105), .B(z_out[87]), .ZN(n13801) );
NAND2_X2 U9104 ( .A1(n17949), .A2(Out_data[87]), .ZN(n13798) );
NAND2_X2 U9105 ( .A1(n18788), .A2(n17942), .ZN(n13797) );
NAND4_X2 U9106 ( .A1(n13803), .A2(n13804), .A3(n13805), .A4(n13806), .ZN(n5613) );
NAND2_X2 U9107 ( .A1(n13807), .A2(n17843), .ZN(n13805) );
XNOR2_X2 U9108 ( .A(n17103), .B(z_out[88]), .ZN(n13807) );
NAND2_X2 U9109 ( .A1(n17949), .A2(Out_data[88]), .ZN(n13804) );
NAND2_X2 U9110 ( .A1(n18787), .A2(n17942), .ZN(n13803) );
NAND4_X2 U9111 ( .A1(n13809), .A2(n13810), .A3(n13811), .A4(n13812), .ZN(n5612) );
NAND2_X2 U9112 ( .A1(n13813), .A2(n17843), .ZN(n13811) );
XNOR2_X2 U9113 ( .A(n17101), .B(z_out[89]), .ZN(n13813) );
NAND2_X2 U9114 ( .A1(n17949), .A2(Out_data[89]), .ZN(n13810) );
NAND2_X2 U9115 ( .A1(n18786), .A2(n17942), .ZN(n13809) );
NAND4_X2 U9116 ( .A1(n13815), .A2(n13816), .A3(n13817), .A4(n13818), .ZN(n5611) );
NAND2_X2 U9117 ( .A1(n13819), .A2(n17843), .ZN(n13817) );
XNOR2_X2 U9118 ( .A(n17099), .B(z_out[90]), .ZN(n13819) );
NAND2_X2 U9119 ( .A1(n17949), .A2(Out_data[90]), .ZN(n13816) );
NAND2_X2 U9120 ( .A1(n18785), .A2(n17942), .ZN(n13815) );
NAND4_X2 U9121 ( .A1(n13821), .A2(n13822), .A3(n13823), .A4(n13824), .ZN(n5610) );
NAND2_X2 U9122 ( .A1(n13825), .A2(n17842), .ZN(n13823) );
XNOR2_X2 U9123 ( .A(n17097), .B(z_out[91]), .ZN(n13825) );
NAND2_X2 U9124 ( .A1(n17949), .A2(Out_data[91]), .ZN(n13822) );
NAND2_X2 U9125 ( .A1(n18784), .A2(n17942), .ZN(n13821) );
NAND4_X2 U9126 ( .A1(n13827), .A2(n13828), .A3(n13829), .A4(n13830), .ZN(n5609) );
NAND2_X2 U9127 ( .A1(n13831), .A2(n17842), .ZN(n13829) );
XNOR2_X2 U9128 ( .A(n17095), .B(z_out[92]), .ZN(n13831) );
NAND2_X2 U9129 ( .A1(n17949), .A2(Out_data[92]), .ZN(n13828) );
NAND2_X2 U9130 ( .A1(n18783), .A2(n17942), .ZN(n13827) );
NAND4_X2 U9131 ( .A1(n13833), .A2(n13834), .A3(n13835), .A4(n13836), .ZN(n5608) );
NAND2_X2 U9132 ( .A1(n13837), .A2(n17842), .ZN(n13835) );
XNOR2_X2 U9133 ( .A(n17093), .B(z_out[93]), .ZN(n13837) );
NAND2_X2 U9134 ( .A1(n17949), .A2(Out_data[93]), .ZN(n13834) );
NAND2_X2 U9135 ( .A1(n18782), .A2(n17942), .ZN(n13833) );
NAND4_X2 U9136 ( .A1(n13839), .A2(n13840), .A3(n13841), .A4(n13842), .ZN(n5607) );
NAND2_X2 U9137 ( .A1(n13843), .A2(n17842), .ZN(n13841) );
XNOR2_X2 U9138 ( .A(n17091), .B(z_out[94]), .ZN(n13843) );
NAND2_X2 U9139 ( .A1(n17949), .A2(Out_data[94]), .ZN(n13840) );
NAND2_X2 U9140 ( .A1(n18781), .A2(n17942), .ZN(n13839) );
NAND4_X2 U9141 ( .A1(n13845), .A2(n13846), .A3(n13847), .A4(n13848), .ZN(n5606) );
NAND2_X2 U9142 ( .A1(n13849), .A2(n17842), .ZN(n13847) );
XNOR2_X2 U9143 ( .A(n17089), .B(z_out[95]), .ZN(n13849) );
NAND2_X2 U9144 ( .A1(n17948), .A2(Out_data[95]), .ZN(n13846) );
NAND2_X2 U9145 ( .A1(n18780), .A2(n17942), .ZN(n13845) );
NAND4_X2 U9146 ( .A1(n13851), .A2(n13852), .A3(n13853), .A4(n13854), .ZN(n5605) );
NAND2_X2 U9147 ( .A1(n13855), .A2(n17842), .ZN(n13853) );
XNOR2_X2 U9148 ( .A(n17087), .B(z_out[96]), .ZN(n13855) );
NAND2_X2 U9149 ( .A1(n17948), .A2(Out_data[96]), .ZN(n13852) );
NAND2_X2 U9150 ( .A1(n18779), .A2(n17942), .ZN(n13851) );
NAND4_X2 U9151 ( .A1(n13857), .A2(n13858), .A3(n13859), .A4(n13860), .ZN(n5604) );
NAND2_X2 U9152 ( .A1(n13861), .A2(n17842), .ZN(n13859) );
XNOR2_X2 U9153 ( .A(n17085), .B(z_out[97]), .ZN(n13861) );
NAND2_X2 U9154 ( .A1(n17948), .A2(Out_data[97]), .ZN(n13858) );
NAND2_X2 U9155 ( .A1(n18778), .A2(n17942), .ZN(n13857) );
NAND4_X2 U9156 ( .A1(n13863), .A2(n13864), .A3(n13865), .A4(n13866), .ZN(n5603) );
NAND2_X2 U9157 ( .A1(n13867), .A2(n17842), .ZN(n13865) );
XNOR2_X2 U9158 ( .A(n17083), .B(z_out[98]), .ZN(n13867) );
NAND2_X2 U9159 ( .A1(n17948), .A2(Out_data[98]), .ZN(n13864) );
NAND2_X2 U9160 ( .A1(n18777), .A2(n17942), .ZN(n13863) );
NAND4_X2 U9161 ( .A1(n13869), .A2(n13870), .A3(n13871), .A4(n13872), .ZN(n5602) );
NAND2_X2 U9162 ( .A1(n13873), .A2(n17842), .ZN(n13871) );
XNOR2_X2 U9163 ( .A(n17081), .B(z_out[99]), .ZN(n13873) );
NAND2_X2 U9164 ( .A1(n17948), .A2(Out_data[99]), .ZN(n13870) );
NAND2_X2 U9165 ( .A1(n18776), .A2(n17943), .ZN(n13869) );
NAND4_X2 U9166 ( .A1(n13875), .A2(n13876), .A3(n13877), .A4(n13878), .ZN(n5601) );
NAND2_X2 U9167 ( .A1(n13879), .A2(n17842), .ZN(n13877) );
XNOR2_X2 U9168 ( .A(n17079), .B(z_out[100]), .ZN(n13879) );
NAND2_X2 U9169 ( .A1(n17948), .A2(Out_data[100]), .ZN(n13876) );
NAND2_X2 U9170 ( .A1(n18775), .A2(n17943), .ZN(n13875) );
NAND4_X2 U9171 ( .A1(n13881), .A2(n13882), .A3(n13883), .A4(n13884), .ZN(n5600) );
NAND2_X2 U9172 ( .A1(n13885), .A2(n17842), .ZN(n13883) );
XNOR2_X2 U9173 ( .A(n17077), .B(z_out[101]), .ZN(n13885) );
NAND2_X2 U9174 ( .A1(n17948), .A2(Out_data[101]), .ZN(n13882) );
NAND2_X2 U9175 ( .A1(n18774), .A2(n17943), .ZN(n13881) );
NAND4_X2 U9176 ( .A1(n13887), .A2(n13888), .A3(n13889), .A4(n13890), .ZN(n5599) );
NAND2_X2 U9177 ( .A1(n13891), .A2(n17842), .ZN(n13889) );
XNOR2_X2 U9178 ( .A(n17075), .B(z_out[102]), .ZN(n13891) );
NAND2_X2 U9179 ( .A1(n17948), .A2(Out_data[102]), .ZN(n13888) );
NAND2_X2 U9180 ( .A1(n18773), .A2(n17943), .ZN(n13887) );
NAND4_X2 U9181 ( .A1(n13893), .A2(n13894), .A3(n13895), .A4(n13896), .ZN(n5598) );
NAND2_X2 U9182 ( .A1(n13897), .A2(n17842), .ZN(n13895) );
XNOR2_X2 U9183 ( .A(n17073), .B(z_out[103]), .ZN(n13897) );
NAND2_X2 U9184 ( .A1(n17948), .A2(Out_data[103]), .ZN(n13894) );
NAND2_X2 U9185 ( .A1(n18772), .A2(n17943), .ZN(n13893) );
NAND4_X2 U9186 ( .A1(n13899), .A2(n13900), .A3(n13901), .A4(n13902), .ZN(n5597) );
NAND2_X2 U9187 ( .A1(n13903), .A2(n17842), .ZN(n13901) );
XNOR2_X2 U9188 ( .A(n17071), .B(z_out[104]), .ZN(n13903) );
NAND2_X2 U9189 ( .A1(n17948), .A2(Out_data[104]), .ZN(n13900) );
NAND2_X2 U9190 ( .A1(n18771), .A2(n17943), .ZN(n13899) );
NAND4_X2 U9191 ( .A1(n13905), .A2(n13906), .A3(n13907), .A4(n13908), .ZN(n5596) );
NAND2_X2 U9192 ( .A1(n13909), .A2(n17842), .ZN(n13907) );
XNOR2_X2 U9193 ( .A(n17069), .B(z_out[105]), .ZN(n13909) );
NAND2_X2 U9194 ( .A1(n17948), .A2(Out_data[105]), .ZN(n13906) );
NAND2_X2 U9195 ( .A1(n18770), .A2(n17943), .ZN(n13905) );
NAND4_X2 U9196 ( .A1(n13911), .A2(n13912), .A3(n13913), .A4(n13914), .ZN(n5595) );
NAND2_X2 U9197 ( .A1(n13915), .A2(n17842), .ZN(n13913) );
XNOR2_X2 U9198 ( .A(n17067), .B(z_out[106]), .ZN(n13915) );
NAND2_X2 U9199 ( .A1(n17947), .A2(Out_data[106]), .ZN(n13912) );
NAND2_X2 U9200 ( .A1(n18769), .A2(n17943), .ZN(n13911) );
NAND4_X2 U9201 ( .A1(n13917), .A2(n13918), .A3(n13919), .A4(n13920), .ZN(n5594) );
NAND2_X2 U9202 ( .A1(n13921), .A2(n17842), .ZN(n13919) );
XNOR2_X2 U9203 ( .A(n17065), .B(z_out[107]), .ZN(n13921) );
NAND2_X2 U9204 ( .A1(n17947), .A2(Out_data[107]), .ZN(n13918) );
NAND2_X2 U9205 ( .A1(n18768), .A2(n17943), .ZN(n13917) );
NAND4_X2 U9206 ( .A1(n13923), .A2(n13924), .A3(n13925), .A4(n13926), .ZN(n5593) );
NAND2_X2 U9207 ( .A1(n13927), .A2(n17842), .ZN(n13925) );
XNOR2_X2 U9208 ( .A(n17063), .B(z_out[108]), .ZN(n13927) );
NAND2_X2 U9209 ( .A1(n17947), .A2(Out_data[108]), .ZN(n13924) );
NAND2_X2 U9210 ( .A1(n18767), .A2(n17943), .ZN(n13923) );
NAND4_X2 U9211 ( .A1(n13929), .A2(n13930), .A3(n13931), .A4(n13932), .ZN(n5592) );
NAND2_X2 U9212 ( .A1(n13933), .A2(n17842), .ZN(n13931) );
XNOR2_X2 U9213 ( .A(n17061), .B(z_out[109]), .ZN(n13933) );
NAND2_X2 U9214 ( .A1(n17947), .A2(Out_data[109]), .ZN(n13930) );
NAND2_X2 U9215 ( .A1(n18766), .A2(n17943), .ZN(n13929) );
NAND4_X2 U9216 ( .A1(n13935), .A2(n13936), .A3(n13937), .A4(n13938), .ZN(n5591) );
NAND2_X2 U9217 ( .A1(n13939), .A2(n17841), .ZN(n13937) );
XNOR2_X2 U9218 ( .A(n17059), .B(z_out[110]), .ZN(n13939) );
NAND2_X2 U9219 ( .A1(n17947), .A2(Out_data[110]), .ZN(n13936) );
NAND2_X2 U9220 ( .A1(n18765), .A2(n17943), .ZN(n13935) );
NAND4_X2 U9221 ( .A1(n13941), .A2(n13942), .A3(n13943), .A4(n13944), .ZN(n5590) );
NAND2_X2 U9222 ( .A1(n13945), .A2(n17841), .ZN(n13943) );
XNOR2_X2 U9223 ( .A(n17057), .B(z_out[111]), .ZN(n13945) );
NAND2_X2 U9224 ( .A1(n17947), .A2(Out_data[111]), .ZN(n13942) );
NAND2_X2 U9225 ( .A1(n18764), .A2(n17944), .ZN(n13941) );
NAND4_X2 U9226 ( .A1(n13947), .A2(n13948), .A3(n13949), .A4(n13950), .ZN(n5589) );
NAND2_X2 U9227 ( .A1(n13951), .A2(n17841), .ZN(n13949) );
XNOR2_X2 U9228 ( .A(n17055), .B(z_out[112]), .ZN(n13951) );
NAND2_X2 U9229 ( .A1(n17947), .A2(Out_data[112]), .ZN(n13948) );
NAND2_X2 U9230 ( .A1(n18763), .A2(n17944), .ZN(n13947) );
NAND4_X2 U9231 ( .A1(n13953), .A2(n13954), .A3(n13955), .A4(n13956), .ZN(n5588) );
NAND2_X2 U9232 ( .A1(n13957), .A2(n17841), .ZN(n13955) );
XNOR2_X2 U9233 ( .A(n17053), .B(z_out[113]), .ZN(n13957) );
NAND2_X2 U9234 ( .A1(n17947), .A2(Out_data[113]), .ZN(n13954) );
NAND2_X2 U9235 ( .A1(n18762), .A2(n17944), .ZN(n13953) );
NAND4_X2 U9236 ( .A1(n13959), .A2(n13960), .A3(n13961), .A4(n13962), .ZN(n5587) );
NAND2_X2 U9237 ( .A1(n13963), .A2(n17841), .ZN(n13961) );
XNOR2_X2 U9238 ( .A(n17051), .B(z_out[114]), .ZN(n13963) );
NAND2_X2 U9239 ( .A1(n17947), .A2(Out_data[114]), .ZN(n13960) );
NAND2_X2 U9240 ( .A1(n18761), .A2(n17944), .ZN(n13959) );
NAND4_X2 U9241 ( .A1(n13965), .A2(n13966), .A3(n13967), .A4(n13968), .ZN(n5586) );
NAND2_X2 U9242 ( .A1(n13969), .A2(n17841), .ZN(n13967) );
XNOR2_X2 U9243 ( .A(n17049), .B(z_out[115]), .ZN(n13969) );
NAND2_X2 U9244 ( .A1(n17947), .A2(Out_data[115]), .ZN(n13966) );
NAND2_X2 U9245 ( .A1(n18760), .A2(n17944), .ZN(n13965) );
NAND4_X2 U9246 ( .A1(n13971), .A2(n13972), .A3(n13973), .A4(n13974), .ZN(n5585) );
NAND2_X2 U9247 ( .A1(n13975), .A2(n17841), .ZN(n13973) );
XNOR2_X2 U9248 ( .A(n17047), .B(z_out[116]), .ZN(n13975) );
NAND2_X2 U9249 ( .A1(n17947), .A2(Out_data[116]), .ZN(n13972) );
NAND2_X2 U9250 ( .A1(n18759), .A2(n17944), .ZN(n13971) );
NAND4_X2 U9251 ( .A1(n13977), .A2(n13978), .A3(n13979), .A4(n13980), .ZN(n5584) );
NAND2_X2 U9252 ( .A1(n13981), .A2(n17841), .ZN(n13979) );
XNOR2_X2 U9253 ( .A(n17045), .B(z_out[117]), .ZN(n13981) );
NAND2_X2 U9254 ( .A1(n17946), .A2(Out_data[117]), .ZN(n13978) );
NAND2_X2 U9255 ( .A1(n18758), .A2(n17944), .ZN(n13977) );
NAND4_X2 U9256 ( .A1(n13983), .A2(n13984), .A3(n13985), .A4(n13986), .ZN(n5583) );
NAND2_X2 U9257 ( .A1(n13987), .A2(n17841), .ZN(n13985) );
XNOR2_X2 U9258 ( .A(n17043), .B(z_out[118]), .ZN(n13987) );
NAND2_X2 U9259 ( .A1(n17946), .A2(Out_data[118]), .ZN(n13984) );
NAND2_X2 U9260 ( .A1(n18757), .A2(n17944), .ZN(n13983) );
NAND4_X2 U9261 ( .A1(n13989), .A2(n13990), .A3(n13991), .A4(n13992), .ZN(n5582) );
NAND2_X2 U9262 ( .A1(n13993), .A2(n17841), .ZN(n13991) );
XNOR2_X2 U9263 ( .A(n17041), .B(z_out[119]), .ZN(n13993) );
NAND2_X2 U9264 ( .A1(n17946), .A2(Out_data[119]), .ZN(n13990) );
NAND2_X2 U9265 ( .A1(n18756), .A2(n17944), .ZN(n13989) );
NAND2_X2 U9267 ( .A1(n13998), .A2(n17841), .ZN(n13996) );
XNOR2_X2 U9268 ( .A(n17039), .B(z_out[120]), .ZN(n13998) );
NAND2_X2 U9269 ( .A1(n17946), .A2(Out_data[120]), .ZN(n13995) );
NAND2_X2 U9271 ( .A1(n14002), .A2(n17841), .ZN(n14000) );
XNOR2_X2 U9272 ( .A(n17037), .B(z_out[121]), .ZN(n14002) );
NAND2_X2 U9273 ( .A1(n17946), .A2(Out_data[121]), .ZN(n13999) );
NAND2_X2 U9275 ( .A1(n14006), .A2(n17841), .ZN(n14004) );
XNOR2_X2 U9276 ( .A(n17035), .B(z_out[122]), .ZN(n14006) );
NAND2_X2 U9277 ( .A1(n17946), .A2(Out_data[122]), .ZN(n14003) );
NAND2_X2 U9279 ( .A1(n14010), .A2(n17841), .ZN(n14008) );
XNOR2_X2 U9280 ( .A(n17033), .B(z_out[123]), .ZN(n14010) );
NAND2_X2 U9281 ( .A1(n17946), .A2(Out_data[123]), .ZN(n14007) );
NAND2_X2 U9283 ( .A1(n14014), .A2(n17841), .ZN(n14012) );
XNOR2_X2 U9284 ( .A(n17031), .B(z_out[124]), .ZN(n14014) );
NAND2_X2 U9285 ( .A1(n17946), .A2(Out_data[124]), .ZN(n14011) );
NAND2_X2 U9287 ( .A1(n14018), .A2(n17841), .ZN(n14016) );
XNOR2_X2 U9288 ( .A(n17029), .B(z_out[125]), .ZN(n14018) );
NAND2_X2 U9289 ( .A1(n17946), .A2(Out_data[125]), .ZN(n14015) );
NAND2_X2 U9291 ( .A1(n14022), .A2(n17841), .ZN(n14020) );
XNOR2_X2 U9292 ( .A(n17027), .B(z_out[126]), .ZN(n14022) );
NAND2_X2 U9293 ( .A1(n17946), .A2(Out_data[126]), .ZN(n14019) );
NAND2_X2 U9295 ( .A1(n14026), .A2(n17841), .ZN(n14024) );
XNOR2_X2 U9296 ( .A(n17025), .B(z_out[127]), .ZN(n14026) );
NAND2_X2 U9297 ( .A1(n17946), .A2(Out_data[127]), .ZN(n14023) );
AND4_X2 U9301 ( .A1(state[9]), .A2(n18845), .A3(n18601), .A4(n18079), .ZN(n11955) );
NAND2_X2 U9622 ( .A1(n18014), .A2(n17747), .ZN(aes_kld) );
AND4_X2 U9624 ( .A1(n18078), .A2(n18629), .A3(n18630), .A4(n14155), .ZN(n11971) );
NAND2_X2 U9631 ( .A1(n14158), .A2(n14159), .ZN(N3198) );
NAND2_X2 U9632 ( .A1(n14160), .A2(n18064), .ZN(n14159) );
XNOR2_X2 U9633 ( .A(n17024), .B(n14161), .ZN(n14160) );
NAND4_X2 U9634 ( .A1(n14025), .A2(n14162), .A3(n14163), .A4(n14164), .ZN(n14161) );
NAND2_X2 U9635 ( .A1(n17916), .A2(n14166), .ZN(n14164) );
NAND2_X2 U9636 ( .A1(n17906), .A2(dii_data[127]), .ZN(n14163) );
AND2_X2 U9638 ( .A1(n14168), .A2(n14169), .ZN(n14025) );
NAND2_X2 U9639 ( .A1(n14170), .A2(n18748), .ZN(n14169) );
NAND2_X2 U9640 ( .A1(n14171), .A2(n14172), .ZN(n14170) );
NAND2_X2 U9641 ( .A1(n17935), .A2(n14166), .ZN(n14172) );
NAND2_X2 U9642 ( .A1(n17288), .A2(dii_data[127]), .ZN(n14171) );
NAND2_X2 U9643 ( .A1(aes_text_out[127]), .A2(n14173), .ZN(n14168) );
NAND2_X2 U9644 ( .A1(n14174), .A2(n14175), .ZN(n14173) );
NAND2_X2 U9645 ( .A1(n19023), .A2(n17944), .ZN(n14175) );
NAND4_X2 U9646 ( .A1(n14176), .A2(n14177), .A3(n14178), .A4(n14179), .ZN(n14166) );
NAND2_X2 U9655 ( .A1(n17877), .A2(dii_data[95]), .ZN(n14177) );
NAND2_X2 U9656 ( .A1(n17849), .A2(dii_data[119]), .ZN(n14176) );
OR2_X2 U9657 ( .A1(n17932), .A2(dii_data[127]), .ZN(n14174) );
NAND2_X2 U9658 ( .A1(n18037), .A2(b_in[111]), .ZN(n14158) );
NAND2_X2 U9659 ( .A1(n14192), .A2(n14193), .ZN(N3197) );
NAND2_X2 U9660 ( .A1(n14194), .A2(n18064), .ZN(n14193) );
XNOR2_X2 U9661 ( .A(n17026), .B(n14195), .ZN(n14194) );
NAND4_X2 U9662 ( .A1(n14021), .A2(n14196), .A3(n14197), .A4(n14198), .ZN(n14195) );
NAND2_X2 U9663 ( .A1(n17916), .A2(n14199), .ZN(n14198) );
NAND2_X2 U9664 ( .A1(n17906), .A2(dii_data[126]), .ZN(n14197) );
AND2_X2 U9666 ( .A1(n14200), .A2(n14201), .ZN(n14021) );
NAND2_X2 U9667 ( .A1(n14202), .A2(n18749), .ZN(n14201) );
NAND2_X2 U9668 ( .A1(n14203), .A2(n14204), .ZN(n14202) );
NAND2_X2 U9669 ( .A1(n17935), .A2(n14199), .ZN(n14204) );
NAND2_X2 U9670 ( .A1(n17288), .A2(dii_data[126]), .ZN(n14203) );
NAND2_X2 U9671 ( .A1(aes_text_out[126]), .A2(n14205), .ZN(n14200) );
NAND2_X2 U9672 ( .A1(n14206), .A2(n14207), .ZN(n14205) );
NAND2_X2 U9673 ( .A1(n19024), .A2(n17944), .ZN(n14207) );
NAND4_X2 U9674 ( .A1(n14208), .A2(n14209), .A3(n14210), .A4(n14211), .ZN(n14199) );
NAND2_X2 U9683 ( .A1(n17873), .A2(dii_data[94]), .ZN(n14209) );
NAND2_X2 U9684 ( .A1(n17848), .A2(dii_data[118]), .ZN(n14208) );
OR2_X2 U9685 ( .A1(n17932), .A2(dii_data[126]), .ZN(n14206) );
NAND2_X2 U9686 ( .A1(n18043), .A2(b_in[110]), .ZN(n14192) );
NAND2_X2 U9687 ( .A1(n14221), .A2(n14222), .ZN(N3196) );
NAND2_X2 U9688 ( .A1(n14223), .A2(n18064), .ZN(n14222) );
XNOR2_X2 U9689 ( .A(n17028), .B(n14224), .ZN(n14223) );
NAND4_X2 U9690 ( .A1(n14017), .A2(n14225), .A3(n14226), .A4(n14227), .ZN(n14224) );
NAND2_X2 U9691 ( .A1(n17916), .A2(n14228), .ZN(n14227) );
NAND2_X2 U9692 ( .A1(n17906), .A2(dii_data[125]), .ZN(n14226) );
AND2_X2 U9694 ( .A1(n14229), .A2(n14230), .ZN(n14017) );
NAND2_X2 U9695 ( .A1(n14231), .A2(n18750), .ZN(n14230) );
NAND2_X2 U9696 ( .A1(n14232), .A2(n14233), .ZN(n14231) );
NAND2_X2 U9697 ( .A1(n17935), .A2(n14228), .ZN(n14233) );
NAND2_X2 U9698 ( .A1(n17288), .A2(dii_data[125]), .ZN(n14232) );
NAND2_X2 U9699 ( .A1(aes_text_out[125]), .A2(n14234), .ZN(n14229) );
NAND2_X2 U9700 ( .A1(n14235), .A2(n14236), .ZN(n14234) );
NAND2_X2 U9701 ( .A1(n19025), .A2(n17944), .ZN(n14236) );
NAND4_X2 U9702 ( .A1(n14237), .A2(n14238), .A3(n14239), .A4(n14240), .ZN(n14228) );
NAND2_X2 U9711 ( .A1(n17873), .A2(dii_data[93]), .ZN(n14238) );
NAND2_X2 U9712 ( .A1(n17848), .A2(dii_data[117]), .ZN(n14237) );
OR2_X2 U9713 ( .A1(n17932), .A2(dii_data[125]), .ZN(n14235) );
NAND2_X2 U9714 ( .A1(n18043), .A2(b_in[109]), .ZN(n14221) );
NAND2_X2 U9715 ( .A1(n14250), .A2(n14251), .ZN(N3195) );
NAND2_X2 U9716 ( .A1(n14252), .A2(n18064), .ZN(n14251) );
XNOR2_X2 U9717 ( .A(n17030), .B(n14253), .ZN(n14252) );
NAND4_X2 U9718 ( .A1(n14013), .A2(n14254), .A3(n14255), .A4(n14256), .ZN(n14253) );
NAND2_X2 U9719 ( .A1(n17916), .A2(n14257), .ZN(n14256) );
NAND2_X2 U9720 ( .A1(n17906), .A2(dii_data[124]), .ZN(n14255) );
AND2_X2 U9722 ( .A1(n14258), .A2(n14259), .ZN(n14013) );
NAND2_X2 U9723 ( .A1(n14260), .A2(n18751), .ZN(n14259) );
NAND2_X2 U9724 ( .A1(n14261), .A2(n14262), .ZN(n14260) );
NAND2_X2 U9725 ( .A1(n17935), .A2(n14257), .ZN(n14262) );
NAND2_X2 U9726 ( .A1(n17288), .A2(dii_data[124]), .ZN(n14261) );
NAND2_X2 U9727 ( .A1(aes_text_out[124]), .A2(n14263), .ZN(n14258) );
NAND2_X2 U9728 ( .A1(n14264), .A2(n14265), .ZN(n14263) );
NAND2_X2 U9729 ( .A1(n19026), .A2(n17945), .ZN(n14265) );
NAND4_X2 U9730 ( .A1(n14266), .A2(n14267), .A3(n14268), .A4(n14269), .ZN(n14257) );
NAND2_X2 U9739 ( .A1(n17873), .A2(dii_data[92]), .ZN(n14267) );
NAND2_X2 U9740 ( .A1(n17848), .A2(dii_data[116]), .ZN(n14266) );
OR2_X2 U9741 ( .A1(n17932), .A2(dii_data[124]), .ZN(n14264) );
NAND2_X2 U9742 ( .A1(n18043), .A2(b_in[108]), .ZN(n14250) );
NAND2_X2 U9743 ( .A1(n14279), .A2(n14280), .ZN(N3194) );
NAND2_X2 U9744 ( .A1(n14281), .A2(n18064), .ZN(n14280) );
XNOR2_X2 U9745 ( .A(n17032), .B(n14282), .ZN(n14281) );
NAND4_X2 U9746 ( .A1(n14009), .A2(n14283), .A3(n14284), .A4(n14285), .ZN(n14282) );
NAND2_X2 U9747 ( .A1(n17915), .A2(n14286), .ZN(n14285) );
NAND2_X2 U9748 ( .A1(n17906), .A2(dii_data[123]), .ZN(n14284) );
AND2_X2 U9750 ( .A1(n14287), .A2(n14288), .ZN(n14009) );
NAND2_X2 U9751 ( .A1(n14289), .A2(n18752), .ZN(n14288) );
NAND2_X2 U9752 ( .A1(n14290), .A2(n14291), .ZN(n14289) );
NAND2_X2 U9753 ( .A1(n17935), .A2(n14286), .ZN(n14291) );
NAND2_X2 U9754 ( .A1(n17288), .A2(dii_data[123]), .ZN(n14290) );
NAND2_X2 U9755 ( .A1(aes_text_out[123]), .A2(n14292), .ZN(n14287) );
NAND2_X2 U9756 ( .A1(n14293), .A2(n14294), .ZN(n14292) );
NAND2_X2 U9757 ( .A1(n19027), .A2(n17945), .ZN(n14294) );
NAND4_X2 U9758 ( .A1(n14295), .A2(n14296), .A3(n14297), .A4(n14298), .ZN(n14286) );
NAND2_X2 U9767 ( .A1(n17873), .A2(dii_data[91]), .ZN(n14296) );
NAND2_X2 U9768 ( .A1(n17848), .A2(dii_data[115]), .ZN(n14295) );
OR2_X2 U9769 ( .A1(n17932), .A2(dii_data[123]), .ZN(n14293) );
NAND2_X2 U9770 ( .A1(n18043), .A2(b_in[107]), .ZN(n14279) );
NAND2_X2 U9771 ( .A1(n14308), .A2(n14309), .ZN(N3193) );
NAND2_X2 U9772 ( .A1(n14310), .A2(n18064), .ZN(n14309) );
XNOR2_X2 U9773 ( .A(n17034), .B(n14311), .ZN(n14310) );
NAND4_X2 U9774 ( .A1(n14005), .A2(n14312), .A3(n14313), .A4(n14314), .ZN(n14311) );
NAND2_X2 U9775 ( .A1(n17915), .A2(n14315), .ZN(n14314) );
NAND2_X2 U9776 ( .A1(n17906), .A2(dii_data[122]), .ZN(n14313) );
AND2_X2 U9778 ( .A1(n14316), .A2(n14317), .ZN(n14005) );
NAND2_X2 U9779 ( .A1(n14318), .A2(n18753), .ZN(n14317) );
NAND2_X2 U9780 ( .A1(n14319), .A2(n14320), .ZN(n14318) );
NAND2_X2 U9781 ( .A1(n17935), .A2(n14315), .ZN(n14320) );
NAND2_X2 U9782 ( .A1(n17288), .A2(dii_data[122]), .ZN(n14319) );
NAND2_X2 U9783 ( .A1(aes_text_out[122]), .A2(n14321), .ZN(n14316) );
NAND2_X2 U9784 ( .A1(n14322), .A2(n14323), .ZN(n14321) );
NAND2_X2 U9785 ( .A1(n19028), .A2(n17945), .ZN(n14323) );
NAND4_X2 U9786 ( .A1(n14324), .A2(n14325), .A3(n14326), .A4(n14327), .ZN(n14315) );
NAND2_X2 U9795 ( .A1(n17873), .A2(dii_data[90]), .ZN(n14325) );
NAND2_X2 U9796 ( .A1(n17848), .A2(dii_data[114]), .ZN(n14324) );
OR2_X2 U9797 ( .A1(n17932), .A2(dii_data[122]), .ZN(n14322) );
NAND2_X2 U9798 ( .A1(n18043), .A2(b_in[106]), .ZN(n14308) );
NAND2_X2 U9799 ( .A1(n14337), .A2(n14338), .ZN(N3192) );
NAND2_X2 U9800 ( .A1(n14339), .A2(n18064), .ZN(n14338) );
XNOR2_X2 U9801 ( .A(n17036), .B(n14340), .ZN(n14339) );
NAND4_X2 U9802 ( .A1(n14001), .A2(n14341), .A3(n14342), .A4(n14343), .ZN(n14340) );
NAND2_X2 U9803 ( .A1(n17915), .A2(n14344), .ZN(n14343) );
NAND2_X2 U9804 ( .A1(n17906), .A2(dii_data[121]), .ZN(n14342) );
AND2_X2 U9806 ( .A1(n14345), .A2(n14346), .ZN(n14001) );
NAND2_X2 U9807 ( .A1(n14347), .A2(n18754), .ZN(n14346) );
NAND2_X2 U9808 ( .A1(n14348), .A2(n14349), .ZN(n14347) );
NAND2_X2 U9809 ( .A1(n17935), .A2(n14344), .ZN(n14349) );
NAND2_X2 U9810 ( .A1(n17288), .A2(dii_data[121]), .ZN(n14348) );
NAND2_X2 U9811 ( .A1(aes_text_out[121]), .A2(n14350), .ZN(n14345) );
NAND2_X2 U9812 ( .A1(n14351), .A2(n14352), .ZN(n14350) );
NAND2_X2 U9813 ( .A1(n19029), .A2(n17945), .ZN(n14352) );
NAND4_X2 U9814 ( .A1(n14353), .A2(n14354), .A3(n14355), .A4(n14356), .ZN(n14344) );
NAND2_X2 U9823 ( .A1(n17873), .A2(dii_data[89]), .ZN(n14354) );
NAND2_X2 U9824 ( .A1(n17848), .A2(dii_data[113]), .ZN(n14353) );
OR2_X2 U9825 ( .A1(n17932), .A2(dii_data[121]), .ZN(n14351) );
NAND2_X2 U9826 ( .A1(n18043), .A2(b_in[105]), .ZN(n14337) );
NAND2_X2 U9827 ( .A1(n14366), .A2(n14367), .ZN(N3191) );
NAND2_X2 U9828 ( .A1(n14368), .A2(n18064), .ZN(n14367) );
XNOR2_X2 U9829 ( .A(n17038), .B(n14369), .ZN(n14368) );
NAND4_X2 U9830 ( .A1(n13997), .A2(n14370), .A3(n14371), .A4(n14372), .ZN(n14369) );
NAND2_X2 U9831 ( .A1(n17915), .A2(n14373), .ZN(n14372) );
NAND2_X2 U9832 ( .A1(n17907), .A2(dii_data[120]), .ZN(n14371) );
AND2_X2 U9834 ( .A1(n14374), .A2(n14375), .ZN(n13997) );
NAND2_X2 U9835 ( .A1(n14376), .A2(n18755), .ZN(n14375) );
NAND2_X2 U9836 ( .A1(n14377), .A2(n14378), .ZN(n14376) );
NAND2_X2 U9837 ( .A1(n17934), .A2(n14373), .ZN(n14378) );
NAND2_X2 U9838 ( .A1(n17288), .A2(dii_data[120]), .ZN(n14377) );
NAND2_X2 U9839 ( .A1(aes_text_out[120]), .A2(n14379), .ZN(n14374) );
NAND2_X2 U9840 ( .A1(n14380), .A2(n14381), .ZN(n14379) );
NAND2_X2 U9841 ( .A1(n19030), .A2(n17945), .ZN(n14381) );
NAND4_X2 U9842 ( .A1(n14382), .A2(n14383), .A3(n14384), .A4(n14385), .ZN(n14373) );
NAND2_X2 U9846 ( .A1(n17897), .A2(n18076), .ZN(n14184) );
NAND2_X2 U9848 ( .A1(n17892), .A2(n18072), .ZN(n14186) );
NAND2_X2 U9850 ( .A1(n14393), .A2(n17892), .ZN(n14187) );
NAND2_X2 U9854 ( .A1(n17873), .A2(dii_data[88]), .ZN(n14383) );
NAND2_X2 U9855 ( .A1(n17848), .A2(dii_data[112]), .ZN(n14382) );
OR2_X2 U9856 ( .A1(n17932), .A2(dii_data[120]), .ZN(n14380) );
NAND2_X2 U9857 ( .A1(n18043), .A2(b_in[104]), .ZN(n14366) );
NAND2_X2 U9858 ( .A1(n14398), .A2(n14399), .ZN(N3190) );
NAND2_X2 U9859 ( .A1(n14400), .A2(n18064), .ZN(n14399) );
XNOR2_X2 U9860 ( .A(n19014), .B(n14401), .ZN(n14400) );
NAND2_X2 U9862 ( .A1(n17919), .A2(n14405), .ZN(n13992) );
XOR2_X2 U9863 ( .A(n17523), .B(aes_text_out[119]), .Z(n14405) );
XNOR2_X2 U9865 ( .A(n14407), .B(aes_text_out[119]), .ZN(n13994) );
AND2_X2 U9866 ( .A1(dii_data[119]), .A2(n17908), .ZN(n14403) );
NAND2_X2 U9867 ( .A1(n14408), .A2(n14409), .ZN(n14402) );
NAND2_X2 U9869 ( .A1(n17915), .A2(n14407), .ZN(n14408) );
NAND4_X2 U9870 ( .A1(n14410), .A2(n14411), .A3(n14412), .A4(n14413), .ZN(n14407) );
NAND2_X2 U9871 ( .A1(n19047), .A2(n17890), .ZN(n14413) );
NAND2_X2 U9875 ( .A1(n19031), .A2(n17896), .ZN(n14411) );
NAND2_X2 U9877 ( .A1(n14421), .A2(n18071), .ZN(n14420) );
NAND2_X2 U9878 ( .A1(n14393), .A2(n19151), .ZN(n14419) );
NAND2_X2 U9879 ( .A1(n17882), .A2(n19032), .ZN(n14418) );
NAND2_X2 U9880 ( .A1(n19079), .A2(n17898), .ZN(n14410) );
NAND2_X2 U9881 ( .A1(n18043), .A2(b_in[103]), .ZN(n14398) );
NAND2_X2 U9882 ( .A1(n14423), .A2(n14424), .ZN(N3189) );
NAND2_X2 U9883 ( .A1(n14425), .A2(n18064), .ZN(n14424) );
XNOR2_X2 U9884 ( .A(n19013), .B(n14426), .ZN(n14425) );
NAND2_X2 U9886 ( .A1(n17919), .A2(n14430), .ZN(n13986) );
XOR2_X2 U9887 ( .A(n17525), .B(aes_text_out[118]), .Z(n14430) );
XNOR2_X2 U9889 ( .A(n14431), .B(aes_text_out[118]), .ZN(n13988) );
AND2_X2 U9890 ( .A1(dii_data[118]), .A2(n17908), .ZN(n14428) );
NAND2_X2 U9891 ( .A1(n14432), .A2(n14433), .ZN(n14427) );
NAND2_X2 U9893 ( .A1(n17915), .A2(n14431), .ZN(n14432) );
NAND4_X2 U9894 ( .A1(n14434), .A2(n14435), .A3(n14436), .A4(n14437), .ZN(n14431) );
NAND2_X2 U9895 ( .A1(n19049), .A2(n17890), .ZN(n14437) );
NAND2_X2 U9899 ( .A1(n19033), .A2(n17896), .ZN(n14435) );
NAND2_X2 U9901 ( .A1(n14444), .A2(n18071), .ZN(n14443) );
NAND2_X2 U9902 ( .A1(n14393), .A2(n19152), .ZN(n14442) );
NAND2_X2 U9903 ( .A1(n17884), .A2(n19034), .ZN(n14441) );
NAND2_X2 U9904 ( .A1(n19082), .A2(n17899), .ZN(n14434) );
NAND2_X2 U9905 ( .A1(n18043), .A2(b_in[102]), .ZN(n14423) );
NAND2_X2 U9906 ( .A1(n14445), .A2(n14446), .ZN(N3188) );
NAND2_X2 U9907 ( .A1(n14447), .A2(n18064), .ZN(n14446) );
XNOR2_X2 U9908 ( .A(n19012), .B(n14448), .ZN(n14447) );
NAND2_X2 U9910 ( .A1(n17919), .A2(n14452), .ZN(n13980) );
XOR2_X2 U9911 ( .A(n17527), .B(aes_text_out[117]), .Z(n14452) );
XNOR2_X2 U9913 ( .A(n14453), .B(aes_text_out[117]), .ZN(n13982) );
AND2_X2 U9914 ( .A1(dii_data[117]), .A2(n17908), .ZN(n14450) );
NAND2_X2 U9915 ( .A1(n14454), .A2(n14455), .ZN(n14449) );
NAND2_X2 U9917 ( .A1(n17915), .A2(n14453), .ZN(n14454) );
NAND4_X2 U9918 ( .A1(n14456), .A2(n14457), .A3(n14458), .A4(n14459), .ZN(n14453) );
NAND2_X2 U9919 ( .A1(n19051), .A2(n17890), .ZN(n14459) );
NAND2_X2 U9923 ( .A1(n19035), .A2(n17896), .ZN(n14457) );
NAND2_X2 U9925 ( .A1(n14466), .A2(n18071), .ZN(n14465) );
NAND2_X2 U9926 ( .A1(n14393), .A2(n19153), .ZN(n14464) );
NAND2_X2 U9927 ( .A1(n17884), .A2(n19036), .ZN(n14463) );
NAND2_X2 U9928 ( .A1(n19085), .A2(n17899), .ZN(n14456) );
NAND2_X2 U9929 ( .A1(n18043), .A2(b_in[101]), .ZN(n14445) );
NAND2_X2 U9930 ( .A1(n14467), .A2(n14468), .ZN(N3187) );
NAND2_X2 U9931 ( .A1(n14469), .A2(n18064), .ZN(n14468) );
XNOR2_X2 U9932 ( .A(n19011), .B(n14470), .ZN(n14469) );
NAND2_X2 U9934 ( .A1(n17919), .A2(n14474), .ZN(n13974) );
XOR2_X2 U9935 ( .A(n17529), .B(aes_text_out[116]), .Z(n14474) );
XNOR2_X2 U9937 ( .A(n14475), .B(aes_text_out[116]), .ZN(n13976) );
AND2_X2 U9938 ( .A1(dii_data[116]), .A2(n17908), .ZN(n14472) );
NAND2_X2 U9939 ( .A1(n14476), .A2(n14477), .ZN(n14471) );
NAND2_X2 U9940 ( .A1(n17998), .A2(aad_byte_cnt[49]), .ZN(n14477) );
NAND2_X2 U9941 ( .A1(n17915), .A2(n14475), .ZN(n14476) );
NAND4_X2 U9942 ( .A1(n14478), .A2(n14479), .A3(n14480), .A4(n14481), .ZN(n14475) );
NAND2_X2 U9943 ( .A1(n19053), .A2(n17890), .ZN(n14481) );
NAND2_X2 U9947 ( .A1(n19037), .A2(n17896), .ZN(n14479) );
NAND2_X2 U9949 ( .A1(n14488), .A2(n18071), .ZN(n14487) );
NAND2_X2 U9950 ( .A1(n14393), .A2(n19154), .ZN(n14486) );
NAND2_X2 U9951 ( .A1(n17884), .A2(n19038), .ZN(n14485) );
NAND2_X2 U9952 ( .A1(n19088), .A2(n17899), .ZN(n14478) );
NAND2_X2 U9953 ( .A1(n18043), .A2(b_in[100]), .ZN(n14467) );
NAND2_X2 U9954 ( .A1(n14489), .A2(n14490), .ZN(N3186) );
NAND2_X2 U9955 ( .A1(n14491), .A2(n18064), .ZN(n14490) );
XNOR2_X2 U9956 ( .A(n19010), .B(n14492), .ZN(n14491) );
NAND2_X2 U9958 ( .A1(n17919), .A2(n14496), .ZN(n13968) );
XOR2_X2 U9959 ( .A(n17531), .B(aes_text_out[115]), .Z(n14496) );
XNOR2_X2 U9961 ( .A(n14497), .B(aes_text_out[115]), .ZN(n13970) );
AND2_X2 U9962 ( .A1(dii_data[115]), .A2(n17908), .ZN(n14494) );
NAND2_X2 U9963 ( .A1(n14498), .A2(n14499), .ZN(n14493) );
NAND2_X2 U9964 ( .A1(n17996), .A2(aad_byte_cnt[48]), .ZN(n14499) );
NAND2_X2 U9965 ( .A1(n17915), .A2(n14497), .ZN(n14498) );
NAND4_X2 U9966 ( .A1(n14500), .A2(n14501), .A3(n14502), .A4(n14503), .ZN(n14497) );
NAND2_X2 U9967 ( .A1(n19055), .A2(n17890), .ZN(n14503) );
NAND2_X2 U9971 ( .A1(n19039), .A2(n17896), .ZN(n14501) );
NAND2_X2 U9973 ( .A1(n14510), .A2(n18071), .ZN(n14509) );
NAND2_X2 U9974 ( .A1(n14393), .A2(n19155), .ZN(n14508) );
NAND2_X2 U9975 ( .A1(n17884), .A2(n19040), .ZN(n14507) );
NAND2_X2 U9976 ( .A1(n19091), .A2(n17899), .ZN(n14500) );
NAND2_X2 U9977 ( .A1(n18043), .A2(b_in[99]), .ZN(n14489) );
NAND2_X2 U9978 ( .A1(n14511), .A2(n14512), .ZN(N3185) );
NAND2_X2 U9979 ( .A1(n14513), .A2(n18064), .ZN(n14512) );
XNOR2_X2 U9980 ( .A(n19009), .B(n14514), .ZN(n14513) );
NAND2_X2 U9982 ( .A1(n17919), .A2(n14518), .ZN(n13962) );
XOR2_X2 U9983 ( .A(n17533), .B(aes_text_out[114]), .Z(n14518) );
XNOR2_X2 U9985 ( .A(n14519), .B(aes_text_out[114]), .ZN(n13964) );
AND2_X2 U9986 ( .A1(dii_data[114]), .A2(n17908), .ZN(n14516) );
NAND2_X2 U9987 ( .A1(n14520), .A2(n14521), .ZN(n14515) );
NAND2_X2 U9988 ( .A1(n17996), .A2(aad_byte_cnt[47]), .ZN(n14521) );
NAND2_X2 U9989 ( .A1(n17915), .A2(n14519), .ZN(n14520) );
NAND4_X2 U9990 ( .A1(n14522), .A2(n14523), .A3(n14524), .A4(n14525), .ZN(n14519) );
NAND2_X2 U9991 ( .A1(n19057), .A2(n17890), .ZN(n14525) );
NAND2_X2 U9995 ( .A1(n19041), .A2(n17896), .ZN(n14523) );
NAND2_X2 U9997 ( .A1(n14532), .A2(n18071), .ZN(n14531) );
NAND2_X2 U9998 ( .A1(n14393), .A2(n19156), .ZN(n14530) );
NAND2_X2 U9999 ( .A1(n17884), .A2(n19042), .ZN(n14529) );
NAND2_X2 U10000 ( .A1(n19094), .A2(n17898), .ZN(n14522) );
NAND2_X2 U10001 ( .A1(n18043), .A2(b_in[98]), .ZN(n14511) );
NAND2_X2 U10002 ( .A1(n14533), .A2(n14534), .ZN(N3184) );
NAND2_X2 U10003 ( .A1(n14535), .A2(n18064), .ZN(n14534) );
XNOR2_X2 U10004 ( .A(n19008), .B(n14536), .ZN(n14535) );
NAND2_X2 U10006 ( .A1(n17919), .A2(n14540), .ZN(n13956) );
XOR2_X2 U10007 ( .A(n17535), .B(aes_text_out[113]), .Z(n14540) );
XNOR2_X2 U10009 ( .A(n14541), .B(aes_text_out[113]), .ZN(n13958) );
AND2_X2 U10010 ( .A1(dii_data[113]), .A2(n17908), .ZN(n14538) );
NAND2_X2 U10011 ( .A1(n14542), .A2(n14543), .ZN(n14537) );
NAND2_X2 U10012 ( .A1(n17996), .A2(aad_byte_cnt[46]), .ZN(n14543) );
NAND2_X2 U10013 ( .A1(n17915), .A2(n14541), .ZN(n14542) );
NAND4_X2 U10014 ( .A1(n14544), .A2(n14545), .A3(n14546), .A4(n14547), .ZN(n14541) );
NAND2_X2 U10015 ( .A1(n19059), .A2(n17889), .ZN(n14547) );
NAND2_X2 U10019 ( .A1(n19043), .A2(n17895), .ZN(n14545) );
NAND2_X2 U10021 ( .A1(n14554), .A2(n18071), .ZN(n14553) );
NAND2_X2 U10022 ( .A1(n14393), .A2(n19157), .ZN(n14552) );
NAND2_X2 U10023 ( .A1(n17884), .A2(n19044), .ZN(n14551) );
NAND2_X2 U10024 ( .A1(n19097), .A2(n17898), .ZN(n14544) );
NAND2_X2 U10025 ( .A1(n18043), .A2(b_in[97]), .ZN(n14533) );
NAND2_X2 U10026 ( .A1(n14555), .A2(n14556), .ZN(N3183) );
NAND2_X2 U10027 ( .A1(n14557), .A2(n18064), .ZN(n14556) );
XNOR2_X2 U10028 ( .A(n19007), .B(n14558), .ZN(n14557) );
NAND2_X2 U10030 ( .A1(n17919), .A2(n14562), .ZN(n13950) );
XOR2_X2 U10031 ( .A(n17537), .B(aes_text_out[112]), .Z(n14562) );
NAND2_X2 U10033 ( .A1(n17935), .A2(n14563), .ZN(n14406) );
NAND2_X2 U10034 ( .A1(n19200), .A2(n14564), .ZN(n14563) );
XNOR2_X2 U10035 ( .A(n14565), .B(aes_text_out[112]), .ZN(n13952) );
AND2_X2 U10036 ( .A1(dii_data[112]), .A2(n17908), .ZN(n14560) );
NAND2_X2 U10037 ( .A1(n14566), .A2(n14567), .ZN(n14559) );
NAND2_X2 U10038 ( .A1(n17996), .A2(aad_byte_cnt[45]), .ZN(n14567) );
NAND2_X2 U10039 ( .A1(n17914), .A2(n14565), .ZN(n14566) );
NAND4_X2 U10040 ( .A1(n14568), .A2(n14569), .A3(n14570), .A4(n14571), .ZN(n14565) );
NAND2_X2 U10041 ( .A1(n19061), .A2(n17889), .ZN(n14571) );
NAND2_X2 U10045 ( .A1(n19045), .A2(n17895), .ZN(n14569) );
NAND2_X2 U10047 ( .A1(n14578), .A2(n18071), .ZN(n14577) );
NAND2_X2 U10048 ( .A1(n14393), .A2(n19158), .ZN(n14576) );
NAND2_X2 U10049 ( .A1(n17884), .A2(n19046), .ZN(n14575) );
NAND2_X2 U10050 ( .A1(n19100), .A2(n17898), .ZN(n14568) );
NAND2_X2 U10051 ( .A1(n18043), .A2(b_in[96]), .ZN(n14555) );
NAND2_X2 U10052 ( .A1(n14579), .A2(n14580), .ZN(N3182) );
NAND2_X2 U10053 ( .A1(n14581), .A2(n18065), .ZN(n14580) );
XNOR2_X2 U10054 ( .A(n19006), .B(n14582), .ZN(n14581) );
NAND2_X2 U10056 ( .A1(n17919), .A2(n14586), .ZN(n13944) );
XNOR2_X2 U10057 ( .A(n19032), .B(aes_text_out[111]), .ZN(n14586) );
XNOR2_X2 U10059 ( .A(n14588), .B(aes_text_out[111]), .ZN(n13946) );
NAND2_X2 U10061 ( .A1(n14589), .A2(n14590), .ZN(n14583) );
NAND2_X2 U10062 ( .A1(n17996), .A2(aad_byte_cnt[44]), .ZN(n14590) );
NAND2_X2 U10063 ( .A1(n17914), .A2(n14588), .ZN(n14589) );
NAND4_X2 U10064 ( .A1(n14591), .A2(n14592), .A3(n14593), .A4(n14594), .ZN(n14588) );
NAND2_X2 U10065 ( .A1(n19063), .A2(n17889), .ZN(n14594) );
NAND2_X2 U10069 ( .A1(n19047), .A2(n17895), .ZN(n14592) );
NAND2_X2 U10071 ( .A1(n19127), .A2(n18071), .ZN(n14600) );
NAND2_X2 U10072 ( .A1(n14393), .A2(n19159), .ZN(n14599) );
NAND2_X2 U10073 ( .A1(n17884), .A2(n19048), .ZN(n14598) );
NAND2_X2 U10074 ( .A1(n19103), .A2(n17898), .ZN(n14591) );
NAND2_X2 U10075 ( .A1(n18043), .A2(b_in[95]), .ZN(n14579) );
NAND2_X2 U10076 ( .A1(n14601), .A2(n14602), .ZN(N3181) );
NAND2_X2 U10077 ( .A1(n14603), .A2(n18065), .ZN(n14602) );
XNOR2_X2 U10078 ( .A(n19005), .B(n14604), .ZN(n14603) );
NAND2_X2 U10080 ( .A1(n17919), .A2(n14608), .ZN(n13938) );
XNOR2_X2 U10081 ( .A(n19034), .B(aes_text_out[110]), .ZN(n14608) );
XNOR2_X2 U10083 ( .A(n14609), .B(aes_text_out[110]), .ZN(n13940) );
NAND2_X2 U10085 ( .A1(n14610), .A2(n14611), .ZN(n14605) );
NAND2_X2 U10086 ( .A1(n17996), .A2(aad_byte_cnt[43]), .ZN(n14611) );
NAND2_X2 U10087 ( .A1(n17914), .A2(n14609), .ZN(n14610) );
NAND4_X2 U10088 ( .A1(n14612), .A2(n14613), .A3(n14614), .A4(n14615), .ZN(n14609) );
NAND2_X2 U10089 ( .A1(n19065), .A2(n17889), .ZN(n14615) );
NAND2_X2 U10093 ( .A1(n19049), .A2(n17895), .ZN(n14613) );
NAND2_X2 U10095 ( .A1(n19128), .A2(n18071), .ZN(n14621) );
NAND2_X2 U10096 ( .A1(n14393), .A2(n19160), .ZN(n14620) );
NAND2_X2 U10097 ( .A1(n17884), .A2(n19050), .ZN(n14619) );
NAND2_X2 U10098 ( .A1(n19106), .A2(n17898), .ZN(n14612) );
NAND2_X2 U10099 ( .A1(n18042), .A2(b_in[94]), .ZN(n14601) );
NAND2_X2 U10100 ( .A1(n14622), .A2(n14623), .ZN(N3180) );
NAND2_X2 U10101 ( .A1(n14624), .A2(n18065), .ZN(n14623) );
XNOR2_X2 U10102 ( .A(n19004), .B(n14625), .ZN(n14624) );
NAND2_X2 U10104 ( .A1(n17919), .A2(n14629), .ZN(n13932) );
XNOR2_X2 U10105 ( .A(n19036), .B(aes_text_out[109]), .ZN(n14629) );
XNOR2_X2 U10107 ( .A(n14630), .B(aes_text_out[109]), .ZN(n13934) );
NAND2_X2 U10109 ( .A1(n14631), .A2(n14632), .ZN(n14626) );
NAND2_X2 U10110 ( .A1(n17996), .A2(aad_byte_cnt[42]), .ZN(n14632) );
NAND2_X2 U10111 ( .A1(n17914), .A2(n14630), .ZN(n14631) );
NAND4_X2 U10112 ( .A1(n14633), .A2(n14634), .A3(n14635), .A4(n14636), .ZN(n14630) );
NAND2_X2 U10113 ( .A1(n19067), .A2(n17889), .ZN(n14636) );
NAND2_X2 U10117 ( .A1(n19051), .A2(n17895), .ZN(n14634) );
NAND2_X2 U10119 ( .A1(n19129), .A2(n18071), .ZN(n14642) );
NAND2_X2 U10120 ( .A1(n14393), .A2(n19161), .ZN(n14641) );
NAND2_X2 U10121 ( .A1(n17884), .A2(n19052), .ZN(n14640) );
NAND2_X2 U10122 ( .A1(n19109), .A2(n17898), .ZN(n14633) );
NAND2_X2 U10123 ( .A1(n18042), .A2(b_in[93]), .ZN(n14622) );
NAND2_X2 U10124 ( .A1(n14643), .A2(n14644), .ZN(N3179) );
NAND2_X2 U10125 ( .A1(n14645), .A2(n18065), .ZN(n14644) );
XNOR2_X2 U10126 ( .A(n19003), .B(n14646), .ZN(n14645) );
NAND2_X2 U10128 ( .A1(n17920), .A2(n14650), .ZN(n13926) );
XNOR2_X2 U10129 ( .A(n19038), .B(aes_text_out[108]), .ZN(n14650) );
XNOR2_X2 U10131 ( .A(n14651), .B(aes_text_out[108]), .ZN(n13928) );
NAND2_X2 U10133 ( .A1(n14652), .A2(n14653), .ZN(n14647) );
NAND2_X2 U10134 ( .A1(n17996), .A2(aad_byte_cnt[41]), .ZN(n14653) );
NAND2_X2 U10135 ( .A1(n17914), .A2(n14651), .ZN(n14652) );
NAND4_X2 U10136 ( .A1(n14654), .A2(n14655), .A3(n14656), .A4(n14657), .ZN(n14651) );
NAND2_X2 U10137 ( .A1(n19069), .A2(n17889), .ZN(n14657) );
NAND2_X2 U10141 ( .A1(n19053), .A2(n17895), .ZN(n14655) );
NAND2_X2 U10143 ( .A1(n19130), .A2(n18071), .ZN(n14663) );
NAND2_X2 U10144 ( .A1(n14393), .A2(n19162), .ZN(n14662) );
NAND2_X2 U10145 ( .A1(n17884), .A2(n19054), .ZN(n14661) );
NAND2_X2 U10146 ( .A1(n19112), .A2(n17898), .ZN(n14654) );
NAND2_X2 U10147 ( .A1(n18042), .A2(b_in[92]), .ZN(n14643) );
NAND2_X2 U10148 ( .A1(n14664), .A2(n14665), .ZN(N3178) );
NAND2_X2 U10149 ( .A1(n14666), .A2(n18065), .ZN(n14665) );
XNOR2_X2 U10150 ( .A(n19002), .B(n14667), .ZN(n14666) );
NAND2_X2 U10152 ( .A1(n17920), .A2(n14671), .ZN(n13920) );
XNOR2_X2 U10153 ( .A(n19040), .B(aes_text_out[107]), .ZN(n14671) );
XNOR2_X2 U10155 ( .A(n14672), .B(aes_text_out[107]), .ZN(n13922) );
NAND2_X2 U10157 ( .A1(n14673), .A2(n14674), .ZN(n14668) );
NAND2_X2 U10158 ( .A1(n17996), .A2(aad_byte_cnt[40]), .ZN(n14674) );
NAND2_X2 U10159 ( .A1(n17914), .A2(n14672), .ZN(n14673) );
NAND4_X2 U10160 ( .A1(n14675), .A2(n14676), .A3(n14677), .A4(n14678), .ZN(n14672) );
NAND2_X2 U10161 ( .A1(n19071), .A2(n17889), .ZN(n14678) );
NAND2_X2 U10165 ( .A1(n19055), .A2(n17895), .ZN(n14676) );
NAND2_X2 U10167 ( .A1(n19131), .A2(n18072), .ZN(n14684) );
NAND2_X2 U10168 ( .A1(n14393), .A2(n19163), .ZN(n14683) );
NAND2_X2 U10169 ( .A1(n17883), .A2(n19056), .ZN(n14682) );
NAND2_X2 U10170 ( .A1(n19115), .A2(n17898), .ZN(n14675) );
NAND2_X2 U10171 ( .A1(n18042), .A2(b_in[91]), .ZN(n14664) );
NAND2_X2 U10172 ( .A1(n14685), .A2(n14686), .ZN(N3177) );
NAND2_X2 U10173 ( .A1(n14687), .A2(n18065), .ZN(n14686) );
XNOR2_X2 U10174 ( .A(n19001), .B(n14688), .ZN(n14687) );
NAND2_X2 U10176 ( .A1(n17920), .A2(n14692), .ZN(n13914) );
XNOR2_X2 U10177 ( .A(n19042), .B(aes_text_out[106]), .ZN(n14692) );
XNOR2_X2 U10179 ( .A(n14693), .B(aes_text_out[106]), .ZN(n13916) );
NAND2_X2 U10181 ( .A1(n14694), .A2(n14695), .ZN(n14689) );
NAND2_X2 U10182 ( .A1(n17996), .A2(aad_byte_cnt[39]), .ZN(n14695) );
NAND2_X2 U10183 ( .A1(n17914), .A2(n14693), .ZN(n14694) );
NAND4_X2 U10184 ( .A1(n14696), .A2(n14697), .A3(n14698), .A4(n14699), .ZN(n14693) );
NAND2_X2 U10185 ( .A1(n19073), .A2(n17889), .ZN(n14699) );
NAND2_X2 U10189 ( .A1(n19057), .A2(n17895), .ZN(n14697) );
NAND2_X2 U10191 ( .A1(n19132), .A2(n18071), .ZN(n14705) );
NAND2_X2 U10192 ( .A1(n14393), .A2(n19164), .ZN(n14704) );
NAND2_X2 U10193 ( .A1(n17883), .A2(n19058), .ZN(n14703) );
NAND2_X2 U10194 ( .A1(n19118), .A2(n17898), .ZN(n14696) );
NAND2_X2 U10195 ( .A1(n18042), .A2(b_in[90]), .ZN(n14685) );
NAND2_X2 U10196 ( .A1(n14706), .A2(n14707), .ZN(N3176) );
NAND2_X2 U10197 ( .A1(n14708), .A2(n18065), .ZN(n14707) );
XNOR2_X2 U10198 ( .A(n19000), .B(n14709), .ZN(n14708) );
NAND2_X2 U10200 ( .A1(n17920), .A2(n14713), .ZN(n13908) );
XNOR2_X2 U10201 ( .A(n19044), .B(aes_text_out[105]), .ZN(n14713) );
XNOR2_X2 U10203 ( .A(n14714), .B(aes_text_out[105]), .ZN(n13910) );
NAND2_X2 U10205 ( .A1(n14715), .A2(n14716), .ZN(n14710) );
NAND2_X2 U10206 ( .A1(n17996), .A2(aad_byte_cnt[38]), .ZN(n14716) );
NAND2_X2 U10207 ( .A1(n17914), .A2(n14714), .ZN(n14715) );
NAND4_X2 U10208 ( .A1(n14717), .A2(n14718), .A3(n14719), .A4(n14720), .ZN(n14714) );
NAND2_X2 U10209 ( .A1(n19075), .A2(n17889), .ZN(n14720) );
NAND2_X2 U10213 ( .A1(n19059), .A2(n17895), .ZN(n14718) );
NAND2_X2 U10215 ( .A1(n19133), .A2(n18071), .ZN(n14726) );
NAND2_X2 U10216 ( .A1(n14393), .A2(n19165), .ZN(n14725) );
NAND2_X2 U10217 ( .A1(n17883), .A2(n19060), .ZN(n14724) );
NAND2_X2 U10218 ( .A1(n19121), .A2(n17898), .ZN(n14717) );
NAND2_X2 U10219 ( .A1(n18042), .A2(b_in[89]), .ZN(n14706) );
NAND2_X2 U10220 ( .A1(n14727), .A2(n14728), .ZN(N3175) );
NAND2_X2 U10221 ( .A1(n14729), .A2(n18065), .ZN(n14728) );
XNOR2_X2 U10222 ( .A(n18999), .B(n14730), .ZN(n14729) );
NAND2_X2 U10224 ( .A1(n17920), .A2(n14734), .ZN(n13902) );
XNOR2_X2 U10225 ( .A(n19046), .B(aes_text_out[104]), .ZN(n14734) );
NAND2_X2 U10227 ( .A1(n17934), .A2(n14735), .ZN(n14587) );
NAND2_X2 U10228 ( .A1(n19200), .A2(n19204), .ZN(n14735) );
XNOR2_X2 U10229 ( .A(n14737), .B(aes_text_out[104]), .ZN(n13904) );
NAND2_X2 U10231 ( .A1(n14738), .A2(n14739), .ZN(n14731) );
NAND2_X2 U10232 ( .A1(n17996), .A2(aad_byte_cnt[37]), .ZN(n14739) );
NAND2_X2 U10233 ( .A1(n17914), .A2(n14737), .ZN(n14738) );
NAND4_X2 U10234 ( .A1(n14740), .A2(n14741), .A3(n14742), .A4(n14743), .ZN(n14737) );
NAND2_X2 U10235 ( .A1(n19077), .A2(n17889), .ZN(n14743) );
NAND2_X2 U10239 ( .A1(n19061), .A2(n17895), .ZN(n14741) );
NAND2_X2 U10241 ( .A1(n19134), .A2(n18071), .ZN(n14749) );
NAND2_X2 U10242 ( .A1(n14393), .A2(n19166), .ZN(n14748) );
NAND2_X2 U10244 ( .A1(n17883), .A2(n19062), .ZN(n14747) );
NAND2_X2 U10245 ( .A1(n19124), .A2(n17898), .ZN(n14740) );
NAND2_X2 U10246 ( .A1(n18042), .A2(b_in[88]), .ZN(n14727) );
NAND2_X2 U10247 ( .A1(n14750), .A2(n14751), .ZN(N3174) );
NAND2_X2 U10248 ( .A1(n14752), .A2(n18065), .ZN(n14751) );
XNOR2_X2 U10249 ( .A(n18998), .B(n14753), .ZN(n14752) );
NAND2_X2 U10251 ( .A1(n17920), .A2(n14757), .ZN(n13896) );
XNOR2_X2 U10252 ( .A(n19048), .B(aes_text_out[103]), .ZN(n14757) );
XNOR2_X2 U10254 ( .A(n14759), .B(aes_text_out[103]), .ZN(n13898) );
NAND2_X2 U10256 ( .A1(n14760), .A2(n14761), .ZN(n14754) );
NAND2_X2 U10257 ( .A1(n17996), .A2(aad_byte_cnt[36]), .ZN(n14761) );
NAND2_X2 U10258 ( .A1(n17914), .A2(n14759), .ZN(n14760) );
NAND4_X2 U10259 ( .A1(n14762), .A2(n14763), .A3(n14764), .A4(n14765), .ZN(n14759) );
NAND2_X2 U10260 ( .A1(n19080), .A2(n17889), .ZN(n14765) );
NAND2_X2 U10264 ( .A1(n19063), .A2(n17895), .ZN(n14763) );
NAND4_X2 U10265 ( .A1(n14769), .A2(n14770), .A3(n14771), .A4(n17881), .ZN(n14417) );
NAND2_X2 U10266 ( .A1(n17883), .A2(n19064), .ZN(n14771) );
NAND2_X2 U10267 ( .A1(n19167), .A2(n18076), .ZN(n14770) );
NAND2_X2 U10268 ( .A1(n19135), .A2(n18071), .ZN(n14769) );
NAND2_X2 U10269 ( .A1(n17897), .A2(n14773), .ZN(n14762) );
NAND2_X2 U10270 ( .A1(n18042), .A2(b_in[87]), .ZN(n14750) );
NAND2_X2 U10271 ( .A1(n14774), .A2(n14775), .ZN(N3173) );
NAND2_X2 U10272 ( .A1(n14776), .A2(n18065), .ZN(n14775) );
XNOR2_X2 U10273 ( .A(n18997), .B(n14777), .ZN(n14776) );
NAND2_X2 U10275 ( .A1(n17920), .A2(n14781), .ZN(n13890) );
XNOR2_X2 U10276 ( .A(n19050), .B(aes_text_out[102]), .ZN(n14781) );
XNOR2_X2 U10278 ( .A(n14782), .B(aes_text_out[102]), .ZN(n13892) );
NAND2_X2 U10280 ( .A1(n14783), .A2(n14784), .ZN(n14778) );
NAND2_X2 U10281 ( .A1(n17996), .A2(aad_byte_cnt[35]), .ZN(n14784) );
NAND2_X2 U10282 ( .A1(n17914), .A2(n14782), .ZN(n14783) );
NAND4_X2 U10283 ( .A1(n14785), .A2(n14786), .A3(n14787), .A4(n14788), .ZN(n14782) );
NAND2_X2 U10284 ( .A1(n19083), .A2(n17889), .ZN(n14788) );
NAND2_X2 U10288 ( .A1(n19065), .A2(n17895), .ZN(n14786) );
NAND4_X2 U10289 ( .A1(n14792), .A2(n14793), .A3(n14794), .A4(n17881), .ZN(n14440) );
NAND2_X2 U10290 ( .A1(n17883), .A2(n19066), .ZN(n14794) );
NAND2_X2 U10291 ( .A1(n19168), .A2(n18076), .ZN(n14793) );
NAND2_X2 U10292 ( .A1(n19136), .A2(n18072), .ZN(n14792) );
NAND2_X2 U10293 ( .A1(n17897), .A2(n14795), .ZN(n14785) );
NAND2_X2 U10294 ( .A1(n18042), .A2(b_in[86]), .ZN(n14774) );
NAND2_X2 U10295 ( .A1(n14796), .A2(n14797), .ZN(N3172) );
NAND2_X2 U10296 ( .A1(n14798), .A2(n18065), .ZN(n14797) );
XNOR2_X2 U10297 ( .A(n18996), .B(n14799), .ZN(n14798) );
NAND2_X2 U10299 ( .A1(n17920), .A2(n14803), .ZN(n13884) );
XNOR2_X2 U10300 ( .A(n19052), .B(aes_text_out[101]), .ZN(n14803) );
XNOR2_X2 U10302 ( .A(n14804), .B(aes_text_out[101]), .ZN(n13886) );
NAND2_X2 U10304 ( .A1(n14805), .A2(n14806), .ZN(n14800) );
NAND2_X2 U10305 ( .A1(n17997), .A2(aad_byte_cnt[34]), .ZN(n14806) );
NAND2_X2 U10306 ( .A1(n17913), .A2(n14804), .ZN(n14805) );
NAND4_X2 U10307 ( .A1(n14807), .A2(n14808), .A3(n14809), .A4(n14810), .ZN(n14804) );
NAND2_X2 U10308 ( .A1(n19086), .A2(n17888), .ZN(n14810) );
NAND2_X2 U10312 ( .A1(n19067), .A2(n17894), .ZN(n14808) );
NAND4_X2 U10313 ( .A1(n14814), .A2(n14815), .A3(n14816), .A4(n17881), .ZN(n14462) );
NAND2_X2 U10314 ( .A1(n17883), .A2(n19068), .ZN(n14816) );
NAND2_X2 U10315 ( .A1(n19169), .A2(n18076), .ZN(n14815) );
NAND2_X2 U10316 ( .A1(n19137), .A2(n18072), .ZN(n14814) );
NAND2_X2 U10317 ( .A1(n17897), .A2(n14817), .ZN(n14807) );
NAND2_X2 U10318 ( .A1(n18042), .A2(b_in[85]), .ZN(n14796) );
NAND2_X2 U10319 ( .A1(n14818), .A2(n14819), .ZN(N3171) );
NAND2_X2 U10320 ( .A1(n14820), .A2(n18065), .ZN(n14819) );
XNOR2_X2 U10321 ( .A(n18995), .B(n14821), .ZN(n14820) );
NAND2_X2 U10323 ( .A1(n17920), .A2(n14825), .ZN(n13878) );
XNOR2_X2 U10324 ( .A(n19054), .B(aes_text_out[100]), .ZN(n14825) );
XNOR2_X2 U10326 ( .A(n14826), .B(aes_text_out[100]), .ZN(n13880) );
NAND2_X2 U10328 ( .A1(n14827), .A2(n14828), .ZN(n14822) );
NAND2_X2 U10329 ( .A1(n17996), .A2(aad_byte_cnt[33]), .ZN(n14828) );
NAND2_X2 U10330 ( .A1(n17913), .A2(n14826), .ZN(n14827) );
NAND4_X2 U10331 ( .A1(n14829), .A2(n14830), .A3(n14831), .A4(n14832), .ZN(n14826) );
NAND2_X2 U10332 ( .A1(n19089), .A2(n17888), .ZN(n14832) );
NAND2_X2 U10336 ( .A1(n19069), .A2(n17894), .ZN(n14830) );
NAND4_X2 U10337 ( .A1(n14836), .A2(n14837), .A3(n14838), .A4(n17881), .ZN(n14484) );
NAND2_X2 U10338 ( .A1(n17883), .A2(n19070), .ZN(n14838) );
NAND2_X2 U10339 ( .A1(n19170), .A2(n18076), .ZN(n14837) );
NAND2_X2 U10340 ( .A1(n19138), .A2(n18072), .ZN(n14836) );
NAND2_X2 U10341 ( .A1(n17897), .A2(n14839), .ZN(n14829) );
NAND2_X2 U10342 ( .A1(n18042), .A2(b_in[84]), .ZN(n14818) );
NAND2_X2 U10343 ( .A1(n14840), .A2(n14841), .ZN(N3170) );
NAND2_X2 U10344 ( .A1(n14842), .A2(n18065), .ZN(n14841) );
XNOR2_X2 U10345 ( .A(n18994), .B(n14843), .ZN(n14842) );
NAND2_X2 U10347 ( .A1(n17920), .A2(n14847), .ZN(n13872) );
XNOR2_X2 U10348 ( .A(n19056), .B(aes_text_out[99]), .ZN(n14847) );
XNOR2_X2 U10350 ( .A(n14848), .B(aes_text_out[99]), .ZN(n13874) );
NAND2_X2 U10352 ( .A1(n14849), .A2(n14850), .ZN(n14844) );
NAND2_X2 U10353 ( .A1(n17996), .A2(aad_byte_cnt[32]), .ZN(n14850) );
NAND2_X2 U10354 ( .A1(n17913), .A2(n14848), .ZN(n14849) );
NAND4_X2 U10355 ( .A1(n14851), .A2(n14852), .A3(n14853), .A4(n14854), .ZN(n14848) );
NAND2_X2 U10356 ( .A1(n19092), .A2(n17888), .ZN(n14854) );
NAND2_X2 U10360 ( .A1(n19071), .A2(n17894), .ZN(n14852) );
NAND4_X2 U10361 ( .A1(n14858), .A2(n14859), .A3(n14860), .A4(n17881), .ZN(n14506) );
NAND2_X2 U10362 ( .A1(n17883), .A2(n19072), .ZN(n14860) );
NAND2_X2 U10363 ( .A1(n19171), .A2(n18076), .ZN(n14859) );
NAND2_X2 U10364 ( .A1(n19139), .A2(n18072), .ZN(n14858) );
NAND2_X2 U10365 ( .A1(n17897), .A2(n14861), .ZN(n14851) );
NAND2_X2 U10366 ( .A1(n18042), .A2(b_in[83]), .ZN(n14840) );
NAND2_X2 U10367 ( .A1(n14862), .A2(n14863), .ZN(N3169) );
NAND2_X2 U10368 ( .A1(n14864), .A2(n18065), .ZN(n14863) );
XNOR2_X2 U10369 ( .A(n18993), .B(n14865), .ZN(n14864) );
NAND2_X2 U10371 ( .A1(n17920), .A2(n14869), .ZN(n13866) );
XNOR2_X2 U10372 ( .A(n19058), .B(aes_text_out[98]), .ZN(n14869) );
XNOR2_X2 U10374 ( .A(n14870), .B(aes_text_out[98]), .ZN(n13868) );
NAND2_X2 U10376 ( .A1(n14871), .A2(n14872), .ZN(n14866) );
NAND2_X2 U10377 ( .A1(n17996), .A2(aad_byte_cnt[31]), .ZN(n14872) );
NAND2_X2 U10378 ( .A1(n17913), .A2(n14870), .ZN(n14871) );
NAND4_X2 U10379 ( .A1(n14873), .A2(n14874), .A3(n14875), .A4(n14876), .ZN(n14870) );
NAND2_X2 U10380 ( .A1(n19095), .A2(n17888), .ZN(n14876) );
NAND2_X2 U10384 ( .A1(n19073), .A2(n17894), .ZN(n14874) );
NAND4_X2 U10385 ( .A1(n14880), .A2(n14881), .A3(n14882), .A4(n17881), .ZN(n14528) );
NAND2_X2 U10386 ( .A1(n17883), .A2(n19074), .ZN(n14882) );
NAND2_X2 U10387 ( .A1(n19172), .A2(n18076), .ZN(n14881) );
NAND2_X2 U10388 ( .A1(n19140), .A2(n18072), .ZN(n14880) );
NAND2_X2 U10389 ( .A1(n17897), .A2(n14883), .ZN(n14873) );
NAND2_X2 U10390 ( .A1(n18042), .A2(b_in[82]), .ZN(n14862) );
NAND2_X2 U10391 ( .A1(n14884), .A2(n14885), .ZN(N3168) );
NAND2_X2 U10392 ( .A1(n14886), .A2(n18065), .ZN(n14885) );
XNOR2_X2 U10393 ( .A(n18992), .B(n14887), .ZN(n14886) );
NAND2_X2 U10395 ( .A1(n17921), .A2(n14891), .ZN(n13860) );
XNOR2_X2 U10396 ( .A(n19060), .B(aes_text_out[97]), .ZN(n14891) );
XNOR2_X2 U10398 ( .A(n14892), .B(aes_text_out[97]), .ZN(n13862) );
NAND2_X2 U10400 ( .A1(n14893), .A2(n14894), .ZN(n14888) );
NAND2_X2 U10401 ( .A1(n17997), .A2(aad_byte_cnt[30]), .ZN(n14894) );
NAND2_X2 U10402 ( .A1(n17913), .A2(n14892), .ZN(n14893) );
NAND4_X2 U10403 ( .A1(n14895), .A2(n14896), .A3(n14897), .A4(n14898), .ZN(n14892) );
NAND2_X2 U10404 ( .A1(n19098), .A2(n17888), .ZN(n14898) );
NAND2_X2 U10408 ( .A1(n19075), .A2(n17894), .ZN(n14896) );
NAND4_X2 U10409 ( .A1(n14902), .A2(n14903), .A3(n14904), .A4(n17881), .ZN(n14550) );
NAND2_X2 U10410 ( .A1(n17882), .A2(n19076), .ZN(n14904) );
NAND2_X2 U10411 ( .A1(n19173), .A2(n18076), .ZN(n14903) );
NAND2_X2 U10412 ( .A1(n19141), .A2(n18072), .ZN(n14902) );
NAND2_X2 U10413 ( .A1(n17897), .A2(n14905), .ZN(n14895) );
NAND2_X2 U10414 ( .A1(n18042), .A2(b_in[81]), .ZN(n14884) );
NAND2_X2 U10415 ( .A1(n14906), .A2(n14907), .ZN(N3167) );
NAND2_X2 U10416 ( .A1(n14908), .A2(n18065), .ZN(n14907) );
XNOR2_X2 U10417 ( .A(n18991), .B(n14909), .ZN(n14908) );
NAND2_X2 U10419 ( .A1(n17921), .A2(n14913), .ZN(n13854) );
XNOR2_X2 U10420 ( .A(n19062), .B(aes_text_out[96]), .ZN(n14913) );
NAND2_X2 U10422 ( .A1(n17934), .A2(n14736), .ZN(n14758) );
NAND2_X2 U10424 ( .A1(dii_data_size[1]), .A2(dii_data_size[0]), .ZN(n14914));
XNOR2_X2 U10425 ( .A(n14915), .B(aes_text_out[96]), .ZN(n13856) );
NAND2_X2 U10427 ( .A1(n14916), .A2(n14917), .ZN(n14910) );
NAND2_X2 U10428 ( .A1(n17997), .A2(aad_byte_cnt[29]), .ZN(n14917) );
NAND2_X2 U10429 ( .A1(n17913), .A2(n14915), .ZN(n14916) );
NAND4_X2 U10430 ( .A1(n14918), .A2(n14919), .A3(n14920), .A4(n14921), .ZN(n14915) );
NAND2_X2 U10431 ( .A1(n19101), .A2(n17888), .ZN(n14921) );
NAND2_X2 U10435 ( .A1(n19077), .A2(n17894), .ZN(n14919) );
NAND4_X2 U10436 ( .A1(n14925), .A2(n14926), .A3(n14927), .A4(n17881), .ZN(n14574) );
NAND2_X2 U10437 ( .A1(n17882), .A2(n19078), .ZN(n14927) );
NAND2_X2 U10438 ( .A1(n19174), .A2(n18076), .ZN(n14926) );
NAND2_X2 U10439 ( .A1(n19142), .A2(n18072), .ZN(n14925) );
NAND2_X2 U10440 ( .A1(n17897), .A2(n14928), .ZN(n14918) );
NAND2_X2 U10441 ( .A1(n18042), .A2(b_in[80]), .ZN(n14906) );
NAND2_X2 U10442 ( .A1(n14929), .A2(n14930), .ZN(N3166) );
NAND2_X2 U10443 ( .A1(n14931), .A2(n18065), .ZN(n14930) );
XNOR2_X2 U10444 ( .A(n18990), .B(n14932), .ZN(n14931) );
NAND2_X2 U10446 ( .A1(n17921), .A2(n14936), .ZN(n13848) );
XNOR2_X2 U10447 ( .A(n19064), .B(aes_text_out[95]), .ZN(n14936) );
XNOR2_X2 U10449 ( .A(n14938), .B(aes_text_out[95]), .ZN(n13850) );
NAND2_X2 U10451 ( .A1(n14939), .A2(n14940), .ZN(n14933) );
NAND2_X2 U10452 ( .A1(n17997), .A2(aad_byte_cnt[28]), .ZN(n14940) );
NAND2_X2 U10453 ( .A1(n17913), .A2(n14938), .ZN(n14939) );
NAND4_X2 U10454 ( .A1(n14941), .A2(n14942), .A3(n14943), .A4(n14944), .ZN(n14938) );
NAND2_X2 U10455 ( .A1(n14945), .A2(n14564), .ZN(n14944) );
NAND2_X2 U10459 ( .A1(n19104), .A2(n17888), .ZN(n14942) );
NAND2_X2 U10460 ( .A1(n19080), .A2(n17894), .ZN(n14941) );
NAND2_X2 U10462 ( .A1(n19143), .A2(n18072), .ZN(n14950) );
NAND2_X2 U10463 ( .A1(dii_data_size[2]), .A2(n14185), .ZN(n14949) );
NAND2_X2 U10464 ( .A1(n14951), .A2(n14952), .ZN(n14185) );
NAND2_X2 U10465 ( .A1(n19175), .A2(n18076), .ZN(n14952) );
NAND2_X2 U10466 ( .A1(n18074), .A2(n19081), .ZN(n14951) );
NAND2_X2 U10467 ( .A1(n18042), .A2(b_in[79]), .ZN(n14929) );
NAND2_X2 U10468 ( .A1(n14953), .A2(n14954), .ZN(N3165) );
NAND2_X2 U10469 ( .A1(n14955), .A2(n18065), .ZN(n14954) );
XNOR2_X2 U10470 ( .A(n18989), .B(n14956), .ZN(n14955) );
NAND2_X2 U10472 ( .A1(n17921), .A2(n14960), .ZN(n13842) );
XNOR2_X2 U10473 ( .A(n19066), .B(aes_text_out[94]), .ZN(n14960) );
XNOR2_X2 U10475 ( .A(n14961), .B(aes_text_out[94]), .ZN(n13844) );
NAND2_X2 U10477 ( .A1(n14962), .A2(n14963), .ZN(n14957) );
NAND2_X2 U10478 ( .A1(n17997), .A2(aad_byte_cnt[27]), .ZN(n14963) );
NAND2_X2 U10479 ( .A1(n17913), .A2(n14961), .ZN(n14962) );
NAND4_X2 U10480 ( .A1(n14964), .A2(n14965), .A3(n14966), .A4(n14967), .ZN(n14961) );
NAND2_X2 U10481 ( .A1(n14968), .A2(n14564), .ZN(n14967) );
NAND2_X2 U10485 ( .A1(n19107), .A2(n17888), .ZN(n14965) );
NAND2_X2 U10486 ( .A1(n19083), .A2(n17894), .ZN(n14964) );
NAND2_X2 U10488 ( .A1(n19144), .A2(n18072), .ZN(n14972) );
NAND2_X2 U10489 ( .A1(dii_data_size[2]), .A2(n14216), .ZN(n14971) );
NAND2_X2 U10490 ( .A1(n14973), .A2(n14974), .ZN(n14216) );
NAND2_X2 U10491 ( .A1(n19176), .A2(n18076), .ZN(n14974) );
NAND2_X2 U10492 ( .A1(n18074), .A2(n19084), .ZN(n14973) );
NAND2_X2 U10493 ( .A1(n18042), .A2(b_in[78]), .ZN(n14953) );
NAND2_X2 U10494 ( .A1(n14975), .A2(n14976), .ZN(N3164) );
NAND2_X2 U10495 ( .A1(n14977), .A2(n18065), .ZN(n14976) );
XNOR2_X2 U10496 ( .A(n18988), .B(n14978), .ZN(n14977) );
NAND2_X2 U10498 ( .A1(n17921), .A2(n14982), .ZN(n13836) );
XNOR2_X2 U10499 ( .A(n19068), .B(aes_text_out[93]), .ZN(n14982) );
XNOR2_X2 U10501 ( .A(n14983), .B(aes_text_out[93]), .ZN(n13838) );
NAND2_X2 U10503 ( .A1(n14984), .A2(n14985), .ZN(n14979) );
NAND2_X2 U10504 ( .A1(n17997), .A2(aad_byte_cnt[26]), .ZN(n14985) );
NAND2_X2 U10505 ( .A1(n17913), .A2(n14983), .ZN(n14984) );
NAND4_X2 U10506 ( .A1(n14986), .A2(n14987), .A3(n14988), .A4(n14989), .ZN(n14983) );
NAND2_X2 U10507 ( .A1(n14990), .A2(n14564), .ZN(n14989) );
NAND2_X2 U10511 ( .A1(n19110), .A2(n17888), .ZN(n14987) );
NAND2_X2 U10512 ( .A1(n19086), .A2(n17894), .ZN(n14986) );
NAND2_X2 U10514 ( .A1(n19145), .A2(n18072), .ZN(n14994) );
NAND2_X2 U10515 ( .A1(dii_data_size[2]), .A2(n14245), .ZN(n14993) );
NAND2_X2 U10516 ( .A1(n14995), .A2(n14996), .ZN(n14245) );
NAND2_X2 U10517 ( .A1(n19177), .A2(n18076), .ZN(n14996) );
NAND2_X2 U10518 ( .A1(n18074), .A2(n19087), .ZN(n14995) );
NAND2_X2 U10519 ( .A1(n18041), .A2(b_in[77]), .ZN(n14975) );
NAND2_X2 U10520 ( .A1(n14997), .A2(n14998), .ZN(N3163) );
NAND2_X2 U10521 ( .A1(n14999), .A2(n18065), .ZN(n14998) );
XNOR2_X2 U10522 ( .A(n18987), .B(n15000), .ZN(n14999) );
NAND2_X2 U10524 ( .A1(n17921), .A2(n15004), .ZN(n13830) );
XNOR2_X2 U10525 ( .A(n19070), .B(aes_text_out[92]), .ZN(n15004) );
XNOR2_X2 U10527 ( .A(n15005), .B(aes_text_out[92]), .ZN(n13832) );
NAND2_X2 U10529 ( .A1(n15006), .A2(n15007), .ZN(n15001) );
NAND2_X2 U10530 ( .A1(n17997), .A2(aad_byte_cnt[25]), .ZN(n15007) );
NAND2_X2 U10531 ( .A1(n17913), .A2(n15005), .ZN(n15006) );
NAND4_X2 U10532 ( .A1(n15008), .A2(n15009), .A3(n15010), .A4(n15011), .ZN(n15005) );
NAND2_X2 U10533 ( .A1(n15012), .A2(n14564), .ZN(n15011) );
NAND2_X2 U10537 ( .A1(n19113), .A2(n17888), .ZN(n15009) );
NAND2_X2 U10538 ( .A1(n19089), .A2(n17894), .ZN(n15008) );
NAND2_X2 U10540 ( .A1(n19146), .A2(n18072), .ZN(n15016) );
NAND2_X2 U10541 ( .A1(dii_data_size[2]), .A2(n14274), .ZN(n15015) );
NAND2_X2 U10542 ( .A1(n15017), .A2(n15018), .ZN(n14274) );
NAND2_X2 U10543 ( .A1(n19178), .A2(n18076), .ZN(n15018) );
NAND2_X2 U10544 ( .A1(n18074), .A2(n19090), .ZN(n15017) );
NAND2_X2 U10545 ( .A1(n18041), .A2(b_in[76]), .ZN(n14997) );
NAND2_X2 U10546 ( .A1(n15019), .A2(n15020), .ZN(N3162) );
NAND2_X2 U10547 ( .A1(n15021), .A2(n18065), .ZN(n15020) );
XNOR2_X2 U10548 ( .A(n18986), .B(n15022), .ZN(n15021) );
NAND2_X2 U10550 ( .A1(n17921), .A2(n15026), .ZN(n13824) );
XNOR2_X2 U10551 ( .A(n19072), .B(aes_text_out[91]), .ZN(n15026) );
XNOR2_X2 U10553 ( .A(n15027), .B(aes_text_out[91]), .ZN(n13826) );
NAND2_X2 U10555 ( .A1(n15028), .A2(n15029), .ZN(n15023) );
NAND2_X2 U10556 ( .A1(n17997), .A2(aad_byte_cnt[24]), .ZN(n15029) );
NAND2_X2 U10557 ( .A1(n17913), .A2(n15027), .ZN(n15028) );
NAND4_X2 U10558 ( .A1(n15030), .A2(n15031), .A3(n15032), .A4(n15033), .ZN(n15027) );
NAND2_X2 U10559 ( .A1(n15034), .A2(n14564), .ZN(n15033) );
NAND2_X2 U10563 ( .A1(n19116), .A2(n17888), .ZN(n15031) );
NAND2_X2 U10564 ( .A1(n19092), .A2(n17894), .ZN(n15030) );
NAND2_X2 U10566 ( .A1(n19147), .A2(n18072), .ZN(n15038) );
NAND2_X2 U10567 ( .A1(dii_data_size[2]), .A2(n14303), .ZN(n15037) );
NAND2_X2 U10568 ( .A1(n15039), .A2(n15040), .ZN(n14303) );
NAND2_X2 U10569 ( .A1(n19179), .A2(n18076), .ZN(n15040) );
NAND2_X2 U10570 ( .A1(n18074), .A2(n19093), .ZN(n15039) );
NAND2_X2 U10571 ( .A1(n18041), .A2(b_in[75]), .ZN(n15019) );
NAND2_X2 U10572 ( .A1(n15041), .A2(n15042), .ZN(N3161) );
NAND2_X2 U10573 ( .A1(n15043), .A2(n18066), .ZN(n15042) );
XNOR2_X2 U10574 ( .A(n18985), .B(n15044), .ZN(n15043) );
NAND2_X2 U10576 ( .A1(n17921), .A2(n15048), .ZN(n13818) );
XNOR2_X2 U10577 ( .A(n19074), .B(aes_text_out[90]), .ZN(n15048) );
XNOR2_X2 U10579 ( .A(n15049), .B(aes_text_out[90]), .ZN(n13820) );
NAND2_X2 U10581 ( .A1(n15050), .A2(n15051), .ZN(n15045) );
NAND2_X2 U10582 ( .A1(n17997), .A2(aad_byte_cnt[23]), .ZN(n15051) );
NAND2_X2 U10583 ( .A1(n17912), .A2(n15049), .ZN(n15050) );
NAND4_X2 U10584 ( .A1(n15052), .A2(n15053), .A3(n15054), .A4(n15055), .ZN(n15049) );
NAND2_X2 U10585 ( .A1(n15056), .A2(n14564), .ZN(n15055) );
NAND2_X2 U10589 ( .A1(n19119), .A2(n17888), .ZN(n15053) );
NAND2_X2 U10590 ( .A1(n19095), .A2(n17893), .ZN(n15052) );
NAND2_X2 U10592 ( .A1(n19148), .A2(n18072), .ZN(n15060) );
NAND2_X2 U10593 ( .A1(dii_data_size[2]), .A2(n14332), .ZN(n15059) );
NAND2_X2 U10594 ( .A1(n15061), .A2(n15062), .ZN(n14332) );
NAND2_X2 U10595 ( .A1(n19180), .A2(n18076), .ZN(n15062) );
NAND2_X2 U10596 ( .A1(n18074), .A2(n19096), .ZN(n15061) );
NAND2_X2 U10597 ( .A1(n18041), .A2(b_in[74]), .ZN(n15041) );
NAND2_X2 U10598 ( .A1(n15063), .A2(n15064), .ZN(N3160) );
NAND2_X2 U10599 ( .A1(n15065), .A2(n18066), .ZN(n15064) );
XNOR2_X2 U10600 ( .A(n18984), .B(n15066), .ZN(n15065) );
NAND2_X2 U10602 ( .A1(n17921), .A2(n15070), .ZN(n13812) );
XNOR2_X2 U10603 ( .A(n19076), .B(aes_text_out[89]), .ZN(n15070) );
XNOR2_X2 U10605 ( .A(n15071), .B(aes_text_out[89]), .ZN(n13814) );
NAND2_X2 U10607 ( .A1(n15072), .A2(n15073), .ZN(n15067) );
NAND2_X2 U10608 ( .A1(n17997), .A2(aad_byte_cnt[22]), .ZN(n15073) );
NAND2_X2 U10609 ( .A1(n17912), .A2(n15071), .ZN(n15072) );
NAND4_X2 U10610 ( .A1(n15074), .A2(n15075), .A3(n15076), .A4(n15077), .ZN(n15071) );
NAND2_X2 U10611 ( .A1(n15078), .A2(n14564), .ZN(n15077) );
NAND2_X2 U10615 ( .A1(n19122), .A2(n17887), .ZN(n15075) );
NAND2_X2 U10616 ( .A1(n19098), .A2(n17893), .ZN(n15074) );
NAND2_X2 U10618 ( .A1(n19149), .A2(n18072), .ZN(n15082) );
NAND2_X2 U10619 ( .A1(dii_data_size[2]), .A2(n14361), .ZN(n15081) );
NAND2_X2 U10620 ( .A1(n15083), .A2(n15084), .ZN(n14361) );
NAND2_X2 U10621 ( .A1(n19181), .A2(n18076), .ZN(n15084) );
NAND2_X2 U10622 ( .A1(n18074), .A2(n19099), .ZN(n15083) );
NAND2_X2 U10623 ( .A1(n18041), .A2(b_in[73]), .ZN(n15063) );
NAND2_X2 U10624 ( .A1(n15085), .A2(n15086), .ZN(N3159) );
NAND2_X2 U10625 ( .A1(n15087), .A2(n18066), .ZN(n15086) );
XNOR2_X2 U10626 ( .A(n18983), .B(n15088), .ZN(n15087) );
NAND2_X2 U10628 ( .A1(n17921), .A2(n15092), .ZN(n13806) );
XNOR2_X2 U10629 ( .A(n19078), .B(aes_text_out[88]), .ZN(n15092) );
NAND2_X2 U10631 ( .A1(n17934), .A2(n15093), .ZN(n14937) );
NAND2_X2 U10632 ( .A1(n19201), .A2(n18072), .ZN(n15093) );
XNOR2_X2 U10633 ( .A(n15095), .B(aes_text_out[88]), .ZN(n13808) );
NAND2_X2 U10635 ( .A1(n15096), .A2(n15097), .ZN(n15089) );
NAND2_X2 U10636 ( .A1(n17997), .A2(aad_byte_cnt[21]), .ZN(n15097) );
NAND2_X2 U10637 ( .A1(n17912), .A2(n15095), .ZN(n15096) );
NAND4_X2 U10638 ( .A1(n15098), .A2(n15099), .A3(n15100), .A4(n15101), .ZN(n15095) );
NAND2_X2 U10639 ( .A1(n15102), .A2(n14564), .ZN(n15101) );
NAND2_X2 U10643 ( .A1(n19125), .A2(n17887), .ZN(n15099) );
NAND2_X2 U10644 ( .A1(n19101), .A2(n17893), .ZN(n15098) );
NAND2_X2 U10646 ( .A1(n19150), .A2(n18072), .ZN(n15106) );
NAND2_X2 U10647 ( .A1(dii_data_size[2]), .A2(n14391), .ZN(n15105) );
NAND2_X2 U10648 ( .A1(n15107), .A2(n15108), .ZN(n14391) );
NAND2_X2 U10649 ( .A1(n19182), .A2(n18076), .ZN(n15108) );
NAND2_X2 U10650 ( .A1(n18074), .A2(n19102), .ZN(n15107) );
NAND2_X2 U10651 ( .A1(n18041), .A2(b_in[72]), .ZN(n15085) );
NAND2_X2 U10652 ( .A1(n15109), .A2(n15110), .ZN(N3158) );
NAND2_X2 U10653 ( .A1(n15111), .A2(n18066), .ZN(n15110) );
XNOR2_X2 U10654 ( .A(n18982), .B(n15112), .ZN(n15111) );
NAND2_X2 U10656 ( .A1(n17921), .A2(n15116), .ZN(n13800) );
XNOR2_X2 U10657 ( .A(n19081), .B(aes_text_out[87]), .ZN(n15116) );
XNOR2_X2 U10659 ( .A(n15118), .B(aes_text_out[87]), .ZN(n13802) );
NAND2_X2 U10661 ( .A1(n15119), .A2(n15120), .ZN(n15113) );
NAND2_X2 U10662 ( .A1(n17997), .A2(aad_byte_cnt[20]), .ZN(n15120) );
NAND2_X2 U10663 ( .A1(n17912), .A2(n15118), .ZN(n15119) );
NAND2_X2 U10669 ( .A1(n14945), .A2(n17887), .ZN(n15122) );
NAND2_X2 U10670 ( .A1(n19104), .A2(n17893), .ZN(n15121) );
NAND2_X2 U10672 ( .A1(n19151), .A2(n18072), .ZN(n15129) );
NAND2_X2 U10673 ( .A1(dii_data_size[2]), .A2(n14421), .ZN(n15128) );
NAND2_X2 U10674 ( .A1(n15130), .A2(n15131), .ZN(n14421) );
NAND2_X2 U10675 ( .A1(n19183), .A2(n18076), .ZN(n15131) );
NAND2_X2 U10676 ( .A1(n18074), .A2(n19105), .ZN(n15130) );
NAND2_X2 U10677 ( .A1(n18041), .A2(b_in[71]), .ZN(n15109) );
NAND2_X2 U10678 ( .A1(n15132), .A2(n15133), .ZN(N3157) );
NAND2_X2 U10679 ( .A1(n15134), .A2(n18066), .ZN(n15133) );
XNOR2_X2 U10680 ( .A(n18981), .B(n15135), .ZN(n15134) );
NAND2_X2 U10682 ( .A1(n17922), .A2(n15139), .ZN(n13794) );
XNOR2_X2 U10683 ( .A(n19084), .B(aes_text_out[86]), .ZN(n15139) );
XNOR2_X2 U10685 ( .A(n15140), .B(aes_text_out[86]), .ZN(n13796) );
NAND2_X2 U10687 ( .A1(n15141), .A2(n15142), .ZN(n15136) );
NAND2_X2 U10688 ( .A1(n17997), .A2(aad_byte_cnt[19]), .ZN(n15142) );
NAND2_X2 U10689 ( .A1(n17912), .A2(n15140), .ZN(n15141) );
NAND2_X2 U10695 ( .A1(n14968), .A2(n17887), .ZN(n15144) );
NAND2_X2 U10696 ( .A1(n19107), .A2(n17893), .ZN(n15143) );
NAND2_X2 U10698 ( .A1(n19152), .A2(n18072), .ZN(n15151) );
NAND2_X2 U10699 ( .A1(dii_data_size[2]), .A2(n14444), .ZN(n15150) );
NAND2_X2 U10700 ( .A1(n15152), .A2(n15153), .ZN(n14444) );
NAND2_X2 U10701 ( .A1(n19184), .A2(n18076), .ZN(n15153) );
NAND2_X2 U10702 ( .A1(n18074), .A2(n19108), .ZN(n15152) );
NAND2_X2 U10703 ( .A1(n18041), .A2(b_in[70]), .ZN(n15132) );
NAND2_X2 U10704 ( .A1(n15154), .A2(n15155), .ZN(N3156) );
NAND2_X2 U10705 ( .A1(n15156), .A2(n18066), .ZN(n15155) );
XNOR2_X2 U10706 ( .A(n18980), .B(n15157), .ZN(n15156) );
NAND2_X2 U10708 ( .A1(n17922), .A2(n15161), .ZN(n13788) );
XNOR2_X2 U10709 ( .A(n19087), .B(aes_text_out[85]), .ZN(n15161) );
XNOR2_X2 U10711 ( .A(n15162), .B(aes_text_out[85]), .ZN(n13790) );
NAND2_X2 U10713 ( .A1(n15163), .A2(n15164), .ZN(n15158) );
NAND2_X2 U10714 ( .A1(n17997), .A2(aad_byte_cnt[18]), .ZN(n15164) );
NAND2_X2 U10715 ( .A1(n17912), .A2(n15162), .ZN(n15163) );
NAND2_X2 U10721 ( .A1(n14990), .A2(n17887), .ZN(n15166) );
NAND2_X2 U10722 ( .A1(n19110), .A2(n17893), .ZN(n15165) );
NAND2_X2 U10724 ( .A1(n19153), .A2(n18072), .ZN(n15173) );
NAND2_X2 U10725 ( .A1(dii_data_size[2]), .A2(n14466), .ZN(n15172) );
NAND2_X2 U10726 ( .A1(n15174), .A2(n15175), .ZN(n14466) );
NAND2_X2 U10727 ( .A1(n19185), .A2(n18076), .ZN(n15175) );
NAND2_X2 U10728 ( .A1(n18074), .A2(n19111), .ZN(n15174) );
NAND2_X2 U10729 ( .A1(n18041), .A2(b_in[69]), .ZN(n15154) );
NAND2_X2 U10730 ( .A1(n15176), .A2(n15177), .ZN(N3155) );
NAND2_X2 U10731 ( .A1(n15178), .A2(n18066), .ZN(n15177) );
XNOR2_X2 U10732 ( .A(n18979), .B(n15179), .ZN(n15178) );
NAND2_X2 U10734 ( .A1(n17922), .A2(n15183), .ZN(n13782) );
XNOR2_X2 U10735 ( .A(n19090), .B(aes_text_out[84]), .ZN(n15183) );
XNOR2_X2 U10737 ( .A(n15184), .B(aes_text_out[84]), .ZN(n13784) );
NAND2_X2 U10739 ( .A1(n15185), .A2(n15186), .ZN(n15180) );
NAND2_X2 U10740 ( .A1(n17997), .A2(aad_byte_cnt[17]), .ZN(n15186) );
NAND2_X2 U10741 ( .A1(n17912), .A2(n15184), .ZN(n15185) );
NAND2_X2 U10747 ( .A1(n15012), .A2(n17887), .ZN(n15188) );
NAND2_X2 U10748 ( .A1(n19113), .A2(n17893), .ZN(n15187) );
NAND2_X2 U10750 ( .A1(n19154), .A2(n18072), .ZN(n15195) );
NAND2_X2 U10751 ( .A1(dii_data_size[2]), .A2(n14488), .ZN(n15194) );
NAND2_X2 U10752 ( .A1(n15196), .A2(n15197), .ZN(n14488) );
NAND2_X2 U10753 ( .A1(n19186), .A2(n18076), .ZN(n15197) );
NAND2_X2 U10754 ( .A1(n18074), .A2(n19114), .ZN(n15196) );
NAND2_X2 U10755 ( .A1(n18041), .A2(b_in[68]), .ZN(n15176) );
NAND2_X2 U10756 ( .A1(n15198), .A2(n15199), .ZN(N3154) );
NAND2_X2 U10757 ( .A1(n15200), .A2(n18066), .ZN(n15199) );
XNOR2_X2 U10758 ( .A(n18978), .B(n15201), .ZN(n15200) );
NAND2_X2 U10760 ( .A1(n17922), .A2(n15205), .ZN(n13776) );
XNOR2_X2 U10761 ( .A(n19093), .B(aes_text_out[83]), .ZN(n15205) );
XNOR2_X2 U10763 ( .A(n15206), .B(aes_text_out[83]), .ZN(n13778) );
NAND2_X2 U10765 ( .A1(n15207), .A2(n15208), .ZN(n15202) );
NAND2_X2 U10766 ( .A1(n17997), .A2(aad_byte_cnt[16]), .ZN(n15208) );
NAND2_X2 U10767 ( .A1(n17912), .A2(n15206), .ZN(n15207) );
NAND2_X2 U10773 ( .A1(n15034), .A2(n17887), .ZN(n15210) );
NAND2_X2 U10774 ( .A1(n19116), .A2(n17893), .ZN(n15209) );
NAND2_X2 U10776 ( .A1(n19155), .A2(n18072), .ZN(n15217) );
NAND2_X2 U10777 ( .A1(dii_data_size[2]), .A2(n14510), .ZN(n15216) );
NAND2_X2 U10778 ( .A1(n15218), .A2(n15219), .ZN(n14510) );
NAND2_X2 U10779 ( .A1(n19187), .A2(n18076), .ZN(n15219) );
NAND2_X2 U10780 ( .A1(n18074), .A2(n19117), .ZN(n15218) );
NAND2_X2 U10781 ( .A1(n18041), .A2(b_in[67]), .ZN(n15198) );
NAND2_X2 U10782 ( .A1(n15220), .A2(n15221), .ZN(N3153) );
NAND2_X2 U10783 ( .A1(n15222), .A2(n18066), .ZN(n15221) );
XNOR2_X2 U10784 ( .A(n18977), .B(n15223), .ZN(n15222) );
NAND2_X2 U10786 ( .A1(n17922), .A2(n15227), .ZN(n13770) );
XNOR2_X2 U10787 ( .A(n19096), .B(aes_text_out[82]), .ZN(n15227) );
XNOR2_X2 U10789 ( .A(n15228), .B(aes_text_out[82]), .ZN(n13772) );
NAND2_X2 U10791 ( .A1(n15229), .A2(n15230), .ZN(n15224) );
NAND2_X2 U10792 ( .A1(n17997), .A2(aad_byte_cnt[15]), .ZN(n15230) );
NAND2_X2 U10793 ( .A1(n17912), .A2(n15228), .ZN(n15229) );
NAND2_X2 U10799 ( .A1(n15056), .A2(n17887), .ZN(n15232) );
NAND2_X2 U10800 ( .A1(n19119), .A2(n17893), .ZN(n15231) );
NAND2_X2 U10802 ( .A1(n19156), .A2(n18072), .ZN(n15239) );
NAND2_X2 U10803 ( .A1(dii_data_size[2]), .A2(n14532), .ZN(n15238) );
NAND2_X2 U10804 ( .A1(n15240), .A2(n15241), .ZN(n14532) );
NAND2_X2 U10805 ( .A1(n19188), .A2(n18076), .ZN(n15241) );
NAND2_X2 U10806 ( .A1(n18074), .A2(n19120), .ZN(n15240) );
NAND2_X2 U10807 ( .A1(n18041), .A2(b_in[66]), .ZN(n15220) );
NAND2_X2 U10808 ( .A1(n15242), .A2(n15243), .ZN(N3152) );
NAND2_X2 U10809 ( .A1(n15244), .A2(n18066), .ZN(n15243) );
XNOR2_X2 U10810 ( .A(n18976), .B(n15245), .ZN(n15244) );
NAND2_X2 U10812 ( .A1(n17922), .A2(n15249), .ZN(n13764) );
XNOR2_X2 U10813 ( .A(n19099), .B(aes_text_out[81]), .ZN(n15249) );
XNOR2_X2 U10815 ( .A(n15250), .B(aes_text_out[81]), .ZN(n13766) );
NAND2_X2 U10817 ( .A1(n15251), .A2(n15252), .ZN(n15246) );
NAND2_X2 U10818 ( .A1(n17997), .A2(aad_byte_cnt[14]), .ZN(n15252) );
NAND2_X2 U10819 ( .A1(n17912), .A2(n15250), .ZN(n15251) );
NAND2_X2 U10825 ( .A1(n15078), .A2(n17887), .ZN(n15254) );
NAND2_X2 U10826 ( .A1(n19122), .A2(n17894), .ZN(n15253) );
NAND2_X2 U10828 ( .A1(n19157), .A2(n18072), .ZN(n15261) );
NAND2_X2 U10829 ( .A1(dii_data_size[2]), .A2(n14554), .ZN(n15260) );
NAND2_X2 U10830 ( .A1(n15262), .A2(n15263), .ZN(n14554) );
NAND2_X2 U10831 ( .A1(n18074), .A2(n19123), .ZN(n15263) );
NAND2_X2 U10832 ( .A1(n19189), .A2(n18076), .ZN(n15262) );
NAND2_X2 U10833 ( .A1(n18041), .A2(b_in[65]), .ZN(n15242) );
NAND2_X2 U10834 ( .A1(n15264), .A2(n15265), .ZN(N3151) );
NAND2_X2 U10835 ( .A1(n15266), .A2(n18066), .ZN(n15265) );
XNOR2_X2 U10836 ( .A(n18975), .B(n15267), .ZN(n15266) );
NAND2_X2 U10838 ( .A1(n17922), .A2(n15271), .ZN(n13758) );
XNOR2_X2 U10839 ( .A(n19102), .B(aes_text_out[80]), .ZN(n15271) );
NAND2_X2 U10841 ( .A1(n17934), .A2(n15094), .ZN(n15117) );
NAND2_X2 U10842 ( .A1(n15272), .A2(n15273), .ZN(n15094) );
NAND2_X2 U10843 ( .A1(dii_data_size[2]), .A2(n17865), .ZN(n15273) );
XNOR2_X2 U10844 ( .A(n15274), .B(aes_text_out[80]), .ZN(n13760) );
NAND2_X2 U10846 ( .A1(n15275), .A2(n15276), .ZN(n15268) );
NAND2_X2 U10847 ( .A1(n17997), .A2(aad_byte_cnt[13]), .ZN(n15276) );
NAND2_X2 U10848 ( .A1(n17912), .A2(n15274), .ZN(n15275) );
NAND2_X2 U10854 ( .A1(n15102), .A2(n17887), .ZN(n15278) );
NAND2_X2 U10855 ( .A1(n19125), .A2(n17893), .ZN(n15277) );
NAND2_X2 U10857 ( .A1(n19158), .A2(n18073), .ZN(n15285) );
NAND2_X2 U10858 ( .A1(dii_data_size[2]), .A2(n14578), .ZN(n15284) );
NAND2_X2 U10859 ( .A1(n15286), .A2(n15287), .ZN(n14578) );
NAND2_X2 U10860 ( .A1(n18074), .A2(n19126), .ZN(n15287) );
NAND2_X2 U10861 ( .A1(n19190), .A2(n18075), .ZN(n15286) );
NAND2_X2 U10862 ( .A1(n18041), .A2(b_in[64]), .ZN(n15264) );
NAND2_X2 U10863 ( .A1(n15288), .A2(n15289), .ZN(N3150) );
NAND2_X2 U10864 ( .A1(n15290), .A2(n18066), .ZN(n15289) );
XNOR2_X2 U10865 ( .A(n18974), .B(n15291), .ZN(n15290) );
NAND2_X2 U10867 ( .A1(n17922), .A2(n15295), .ZN(n13752) );
XNOR2_X2 U10868 ( .A(n19105), .B(aes_text_out[79]), .ZN(n15295) );
XNOR2_X2 U10870 ( .A(n15297), .B(aes_text_out[79]), .ZN(n13754) );
NAND2_X2 U10872 ( .A1(n15298), .A2(n15299), .ZN(n15292) );
NAND2_X2 U10873 ( .A1(n17997), .A2(aad_byte_cnt[12]), .ZN(n15299) );
NAND2_X2 U10874 ( .A1(n17911), .A2(n15297), .ZN(n15298) );
NAND4_X2 U10875 ( .A1(n15300), .A2(n15301), .A3(n15302), .A4(n15303), .ZN(n15297) );
AND2_X2 U10880 ( .A1(n15307), .A2(n15308), .ZN(n15127) );
NAND2_X2 U10881 ( .A1(dii_data[31]), .A2(n15309), .ZN(n15308) );
NAND2_X2 U10882 ( .A1(n17882), .A2(dii_data[63]), .ZN(n15307) );
NAND2_X2 U10883 ( .A1(n17857), .A2(dii_data[55]), .ZN(n15302) );
NAND2_X2 U10884 ( .A1(n14945), .A2(n17893), .ZN(n15301) );
AND3_X2 U10885 ( .A1(n15310), .A2(n17881), .A3(n15311), .ZN(n14945) );
NAND2_X2 U10886 ( .A1(n19159), .A2(n18073), .ZN(n15311) );
NAND2_X2 U10887 ( .A1(n19127), .A2(dii_data_size[2]), .ZN(n15310) );
NAND2_X2 U10888 ( .A1(n15312), .A2(n15313), .ZN(n14773) );
NAND2_X2 U10889 ( .A1(dii_data[71]), .A2(n18074), .ZN(n15313) );
NAND2_X2 U10890 ( .A1(dii_data[7]), .A2(n18075), .ZN(n15312) );
NAND2_X2 U10891 ( .A1(n19202), .A2(n17713), .ZN(n15300) );
NAND2_X2 U10892 ( .A1(n18041), .A2(b_in[63]), .ZN(n15288) );
NAND2_X2 U10893 ( .A1(n15314), .A2(n15315), .ZN(N3149) );
NAND2_X2 U10894 ( .A1(n15316), .A2(n18066), .ZN(n15315) );
XNOR2_X2 U10895 ( .A(n18973), .B(n15317), .ZN(n15316) );
NAND2_X2 U10897 ( .A1(n17922), .A2(n15321), .ZN(n13746) );
XNOR2_X2 U10898 ( .A(n19108), .B(aes_text_out[78]), .ZN(n15321) );
XNOR2_X2 U10900 ( .A(n15322), .B(aes_text_out[78]), .ZN(n13748) );
NAND2_X2 U10902 ( .A1(n15323), .A2(n15324), .ZN(n15318) );
NAND2_X2 U10903 ( .A1(n17997), .A2(aad_byte_cnt[11]), .ZN(n15324) );
NAND2_X2 U10904 ( .A1(n17911), .A2(n15322), .ZN(n15323) );
NAND4_X2 U10905 ( .A1(n15325), .A2(n15326), .A3(n15327), .A4(n15328), .ZN(n15322) );
AND2_X2 U10910 ( .A1(n15332), .A2(n15333), .ZN(n15149) );
NAND2_X2 U10911 ( .A1(dii_data[30]), .A2(n15309), .ZN(n15333) );
NAND2_X2 U10912 ( .A1(n17882), .A2(dii_data[62]), .ZN(n15332) );
NAND2_X2 U10913 ( .A1(n17859), .A2(dii_data[54]), .ZN(n15327) );
NAND2_X2 U10914 ( .A1(n14968), .A2(n17893), .ZN(n15326) );
AND3_X2 U10915 ( .A1(n15334), .A2(n17881), .A3(n15335), .ZN(n14968) );
NAND2_X2 U10916 ( .A1(n19160), .A2(n18073), .ZN(n15335) );
NAND2_X2 U10917 ( .A1(n19128), .A2(dii_data_size[2]), .ZN(n15334) );
NAND2_X2 U10918 ( .A1(n15336), .A2(n15337), .ZN(n14795) );
NAND2_X2 U10919 ( .A1(dii_data[6]), .A2(n18075), .ZN(n15337) );
NAND2_X2 U10920 ( .A1(dii_data[70]), .A2(n18074), .ZN(n15336) );
NAND2_X2 U10921 ( .A1(n19202), .A2(n17715), .ZN(n15325) );
NAND2_X2 U10922 ( .A1(n18041), .A2(b_in[62]), .ZN(n15314) );
NAND2_X2 U10923 ( .A1(n15338), .A2(n15339), .ZN(N3148) );
NAND2_X2 U10924 ( .A1(n15340), .A2(n18066), .ZN(n15339) );
XNOR2_X2 U10925 ( .A(n18972), .B(n15341), .ZN(n15340) );
NAND2_X2 U10927 ( .A1(n17922), .A2(n15345), .ZN(n13740) );
XNOR2_X2 U10928 ( .A(n19111), .B(aes_text_out[77]), .ZN(n15345) );
XNOR2_X2 U10930 ( .A(n15346), .B(aes_text_out[77]), .ZN(n13742) );
NAND2_X2 U10932 ( .A1(n15347), .A2(n15348), .ZN(n15342) );
NAND2_X2 U10933 ( .A1(n17998), .A2(aad_byte_cnt[10]), .ZN(n15348) );
NAND2_X2 U10934 ( .A1(n17911), .A2(n15346), .ZN(n15347) );
NAND4_X2 U10935 ( .A1(n15349), .A2(n15350), .A3(n15351), .A4(n15352), .ZN(n15346) );
AND2_X2 U10940 ( .A1(n15356), .A2(n15357), .ZN(n15171) );
NAND2_X2 U10941 ( .A1(dii_data[29]), .A2(n15309), .ZN(n15357) );
NAND2_X2 U10942 ( .A1(n17883), .A2(dii_data[61]), .ZN(n15356) );
NAND2_X2 U10943 ( .A1(n17859), .A2(dii_data[53]), .ZN(n15351) );
NAND2_X2 U10944 ( .A1(n14990), .A2(n17892), .ZN(n15350) );
AND3_X2 U10945 ( .A1(n15358), .A2(n17881), .A3(n15359), .ZN(n14990) );
NAND2_X2 U10946 ( .A1(n19161), .A2(n18073), .ZN(n15359) );
NAND2_X2 U10947 ( .A1(n19129), .A2(dii_data_size[2]), .ZN(n15358) );
NAND2_X2 U10948 ( .A1(n15360), .A2(n15361), .ZN(n14817) );
NAND2_X2 U10949 ( .A1(dii_data[5]), .A2(n18075), .ZN(n15361) );
NAND2_X2 U10950 ( .A1(dii_data[69]), .A2(n18074), .ZN(n15360) );
NAND2_X2 U10951 ( .A1(n19202), .A2(n17717), .ZN(n15349) );
NAND2_X2 U10952 ( .A1(n18041), .A2(b_in[61]), .ZN(n15338) );
NAND2_X2 U10953 ( .A1(n15362), .A2(n15363), .ZN(N3147) );
NAND2_X2 U10954 ( .A1(n15364), .A2(n18066), .ZN(n15363) );
XNOR2_X2 U10955 ( .A(n18971), .B(n15365), .ZN(n15364) );
NAND2_X2 U10957 ( .A1(n17922), .A2(n15369), .ZN(n13734) );
XNOR2_X2 U10958 ( .A(n19114), .B(aes_text_out[76]), .ZN(n15369) );
XNOR2_X2 U10960 ( .A(n15370), .B(aes_text_out[76]), .ZN(n13736) );
NAND2_X2 U10962 ( .A1(n15371), .A2(n15372), .ZN(n15366) );
NAND2_X2 U10963 ( .A1(n17998), .A2(aad_byte_cnt[9]), .ZN(n15372) );
NAND2_X2 U10964 ( .A1(n17911), .A2(n15370), .ZN(n15371) );
NAND4_X2 U10965 ( .A1(n15373), .A2(n15374), .A3(n15375), .A4(n15376), .ZN(n15370) );
AND2_X2 U10970 ( .A1(n15380), .A2(n15381), .ZN(n15193) );
NAND2_X2 U10971 ( .A1(dii_data[28]), .A2(n15309), .ZN(n15381) );
NAND2_X2 U10972 ( .A1(n17882), .A2(dii_data[60]), .ZN(n15380) );
NAND2_X2 U10973 ( .A1(n17859), .A2(dii_data[52]), .ZN(n15375) );
NAND2_X2 U10974 ( .A1(n15012), .A2(n17892), .ZN(n15374) );
AND3_X2 U10975 ( .A1(n15382), .A2(n17881), .A3(n15383), .ZN(n15012) );
NAND2_X2 U10976 ( .A1(n19162), .A2(n18073), .ZN(n15383) );
NAND2_X2 U10977 ( .A1(n19130), .A2(dii_data_size[2]), .ZN(n15382) );
NAND2_X2 U10978 ( .A1(n15384), .A2(n15385), .ZN(n14839) );
NAND2_X2 U10979 ( .A1(dii_data[4]), .A2(n18075), .ZN(n15385) );
NAND2_X2 U10980 ( .A1(dii_data[68]), .A2(n18074), .ZN(n15384) );
NAND2_X2 U10981 ( .A1(n19202), .A2(n17719), .ZN(n15373) );
NAND2_X2 U10982 ( .A1(n18040), .A2(b_in[60]), .ZN(n15362) );
NAND2_X2 U10983 ( .A1(n15386), .A2(n15387), .ZN(N3146) );
NAND2_X2 U10984 ( .A1(n15388), .A2(n18066), .ZN(n15387) );
XNOR2_X2 U10985 ( .A(n18970), .B(n15389), .ZN(n15388) );
NAND2_X2 U10987 ( .A1(n17923), .A2(n15393), .ZN(n13728) );
XNOR2_X2 U10988 ( .A(n19117), .B(aes_text_out[75]), .ZN(n15393) );
XNOR2_X2 U10990 ( .A(n15394), .B(aes_text_out[75]), .ZN(n13730) );
NAND2_X2 U10992 ( .A1(n15395), .A2(n15396), .ZN(n15390) );
NAND2_X2 U10993 ( .A1(n17998), .A2(aad_byte_cnt[8]), .ZN(n15396) );
NAND2_X2 U10994 ( .A1(n17911), .A2(n15394), .ZN(n15395) );
NAND4_X2 U10995 ( .A1(n15397), .A2(n15398), .A3(n15399), .A4(n15400), .ZN(n15394) );
AND2_X2 U11000 ( .A1(n15404), .A2(n15405), .ZN(n15215) );
NAND2_X2 U11001 ( .A1(dii_data[27]), .A2(n15309), .ZN(n15405) );
NAND2_X2 U11002 ( .A1(n17882), .A2(dii_data[59]), .ZN(n15404) );
NAND2_X2 U11003 ( .A1(n17859), .A2(dii_data[51]), .ZN(n15399) );
NAND2_X2 U11004 ( .A1(n15034), .A2(n17892), .ZN(n15398) );
AND3_X2 U11005 ( .A1(n15406), .A2(n17881), .A3(n15407), .ZN(n15034) );
NAND2_X2 U11006 ( .A1(n19163), .A2(n18073), .ZN(n15407) );
NAND2_X2 U11007 ( .A1(n19131), .A2(dii_data_size[2]), .ZN(n15406) );
NAND2_X2 U11008 ( .A1(n15408), .A2(n15409), .ZN(n14861) );
NAND2_X2 U11009 ( .A1(dii_data[3]), .A2(n18075), .ZN(n15409) );
NAND2_X2 U11010 ( .A1(dii_data[67]), .A2(n18074), .ZN(n15408) );
NAND2_X2 U11011 ( .A1(n19202), .A2(n17721), .ZN(n15397) );
NAND2_X2 U11012 ( .A1(n18040), .A2(b_in[59]), .ZN(n15386) );
NAND2_X2 U11013 ( .A1(n15410), .A2(n15411), .ZN(N3145) );
NAND2_X2 U11014 ( .A1(n15412), .A2(n18066), .ZN(n15411) );
XNOR2_X2 U11015 ( .A(n18969), .B(n15413), .ZN(n15412) );
NAND2_X2 U11017 ( .A1(n17923), .A2(n15417), .ZN(n13722) );
XNOR2_X2 U11018 ( .A(n19120), .B(aes_text_out[74]), .ZN(n15417) );
XNOR2_X2 U11020 ( .A(n15418), .B(aes_text_out[74]), .ZN(n13724) );
NAND2_X2 U11022 ( .A1(n15419), .A2(n15420), .ZN(n15414) );
NAND2_X2 U11023 ( .A1(n17998), .A2(aad_byte_cnt[7]), .ZN(n15420) );
NAND2_X2 U11024 ( .A1(n17911), .A2(n15418), .ZN(n15419) );
NAND4_X2 U11025 ( .A1(n15421), .A2(n15422), .A3(n15423), .A4(n15424), .ZN(n15418) );
AND2_X2 U11030 ( .A1(n15428), .A2(n15429), .ZN(n15237) );
NAND2_X2 U11031 ( .A1(dii_data[26]), .A2(n15309), .ZN(n15429) );
NAND2_X2 U11032 ( .A1(n17882), .A2(dii_data[58]), .ZN(n15428) );
NAND2_X2 U11033 ( .A1(n17859), .A2(dii_data[50]), .ZN(n15423) );
NAND2_X2 U11034 ( .A1(n15056), .A2(n17892), .ZN(n15422) );
AND3_X2 U11035 ( .A1(n15430), .A2(n17881), .A3(n15431), .ZN(n15056) );
NAND2_X2 U11036 ( .A1(n19164), .A2(n18073), .ZN(n15431) );
NAND2_X2 U11037 ( .A1(n19132), .A2(dii_data_size[2]), .ZN(n15430) );
NAND2_X2 U11038 ( .A1(n15432), .A2(n15433), .ZN(n14883) );
NAND2_X2 U11039 ( .A1(dii_data[2]), .A2(n18075), .ZN(n15433) );
NAND2_X2 U11040 ( .A1(dii_data[66]), .A2(n18074), .ZN(n15432) );
NAND2_X2 U11041 ( .A1(n19202), .A2(n17723), .ZN(n15421) );
NAND2_X2 U11042 ( .A1(n18040), .A2(b_in[58]), .ZN(n15410) );
NAND2_X2 U11043 ( .A1(n15434), .A2(n15435), .ZN(N3144) );
NAND2_X2 U11044 ( .A1(n15436), .A2(n18066), .ZN(n15435) );
XNOR2_X2 U11045 ( .A(n18968), .B(n15437), .ZN(n15436) );
NAND2_X2 U11047 ( .A1(n17923), .A2(n15441), .ZN(n13716) );
XNOR2_X2 U11048 ( .A(n19123), .B(aes_text_out[73]), .ZN(n15441) );
XNOR2_X2 U11050 ( .A(n15442), .B(aes_text_out[73]), .ZN(n13718) );
NAND2_X2 U11052 ( .A1(n15443), .A2(n15444), .ZN(n15438) );
NAND2_X2 U11053 ( .A1(n17998), .A2(aad_byte_cnt[6]), .ZN(n15444) );
NAND2_X2 U11054 ( .A1(n17911), .A2(n15442), .ZN(n15443) );
NAND4_X2 U11055 ( .A1(n15445), .A2(n15446), .A3(n15447), .A4(n15448), .ZN(n15442) );
AND2_X2 U11060 ( .A1(n15452), .A2(n15453), .ZN(n15259) );
NAND2_X2 U11061 ( .A1(dii_data[25]), .A2(n15309), .ZN(n15453) );
NAND2_X2 U11062 ( .A1(n17882), .A2(dii_data[57]), .ZN(n15452) );
NAND2_X2 U11063 ( .A1(n17859), .A2(dii_data[49]), .ZN(n15447) );
NAND2_X2 U11064 ( .A1(n15078), .A2(n17892), .ZN(n15446) );
AND3_X2 U11065 ( .A1(n15454), .A2(n17881), .A3(n15455), .ZN(n15078) );
NAND2_X2 U11066 ( .A1(n19165), .A2(n18073), .ZN(n15455) );
NAND2_X2 U11067 ( .A1(n19133), .A2(dii_data_size[2]), .ZN(n15454) );
NAND2_X2 U11068 ( .A1(n15456), .A2(n15457), .ZN(n14905) );
NAND2_X2 U11069 ( .A1(dii_data[1]), .A2(n18075), .ZN(n15457) );
NAND2_X2 U11070 ( .A1(dii_data[65]), .A2(n18074), .ZN(n15456) );
NAND2_X2 U11071 ( .A1(n19202), .A2(n17725), .ZN(n15445) );
NAND2_X2 U11072 ( .A1(n18040), .A2(b_in[57]), .ZN(n15434) );
NAND2_X2 U11073 ( .A1(n15458), .A2(n15459), .ZN(N3143) );
NAND2_X2 U11074 ( .A1(n15460), .A2(n18066), .ZN(n15459) );
XNOR2_X2 U11075 ( .A(n18967), .B(n15461), .ZN(n15460) );
NAND2_X2 U11077 ( .A1(n17923), .A2(n15465), .ZN(n13710) );
XNOR2_X2 U11078 ( .A(n19126), .B(aes_text_out[72]), .ZN(n15465) );
NAND2_X2 U11080 ( .A1(n17934), .A2(n15466), .ZN(n15296) );
NAND2_X2 U11081 ( .A1(n15272), .A2(n15467), .ZN(n15466) );
NAND2_X2 U11082 ( .A1(n17892), .A2(dii_data_size[2]), .ZN(n15467) );
XNOR2_X2 U11083 ( .A(n15468), .B(aes_text_out[72]), .ZN(n13712) );
NAND2_X2 U11085 ( .A1(n15469), .A2(n15470), .ZN(n15462) );
NAND2_X2 U11086 ( .A1(n17998), .A2(aad_byte_cnt[5]), .ZN(n15470) );
NAND2_X2 U11087 ( .A1(n17911), .A2(n15468), .ZN(n15469) );
NAND4_X2 U11088 ( .A1(n15471), .A2(n15472), .A3(n15473), .A4(n15474), .ZN(n15468) );
AND2_X2 U11094 ( .A1(n15478), .A2(n15479), .ZN(n15283) );
NAND2_X2 U11095 ( .A1(dii_data[24]), .A2(n15309), .ZN(n15479) );
NAND2_X2 U11096 ( .A1(n17882), .A2(dii_data[56]), .ZN(n15478) );
NAND2_X2 U11097 ( .A1(n17859), .A2(dii_data[48]), .ZN(n15473) );
NAND2_X2 U11098 ( .A1(n15102), .A2(n17892), .ZN(n15472) );
AND3_X2 U11099 ( .A1(n15480), .A2(n17881), .A3(n15481), .ZN(n15102) );
NAND2_X2 U11100 ( .A1(n19166), .A2(n18071), .ZN(n15481) );
NAND2_X2 U11102 ( .A1(n19134), .A2(dii_data_size[2]), .ZN(n15480) );
NAND2_X2 U11103 ( .A1(n15482), .A2(n15483), .ZN(n14928) );
NAND2_X2 U11104 ( .A1(dii_data[0]), .A2(n18075), .ZN(n15483) );
NAND2_X2 U11105 ( .A1(dii_data[64]), .A2(n18074), .ZN(n15482) );
NAND2_X2 U11106 ( .A1(n19202), .A2(n17727), .ZN(n15471) );
NAND2_X2 U11107 ( .A1(n18040), .A2(b_in[56]), .ZN(n15458) );
NAND2_X2 U11108 ( .A1(n15484), .A2(n15485), .ZN(N3142) );
NAND2_X2 U11109 ( .A1(n15486), .A2(n18066), .ZN(n15485) );
XNOR2_X2 U11110 ( .A(n18966), .B(n15487), .ZN(n15486) );
XOR2_X2 U11114 ( .A(aes_text_out[71]), .B(n15491), .Z(n13706) );
AND4_X2 U11115 ( .A1(n15493), .A2(n15494), .A3(n15495), .A4(n15496), .ZN(n15491) );
NAND2_X2 U11124 ( .A1(n17848), .A2(dii_data[63]), .ZN(n15494) );
NAND2_X2 U11125 ( .A1(n15509), .A2(dii_data[7]), .ZN(n15493) );
NAND2_X2 U11126 ( .A1(n15510), .A2(n15511), .ZN(n15488) );
NAND2_X2 U11127 ( .A1(n17906), .A2(dii_data[71]), .ZN(n15511) );
NAND2_X2 U11128 ( .A1(n17998), .A2(aad_byte_cnt[4]), .ZN(n15510) );
NAND2_X2 U11129 ( .A1(n17923), .A2(n15512), .ZN(n13704) );
XOR2_X2 U11130 ( .A(n17617), .B(aes_text_out[71]), .Z(n15512) );
NAND2_X2 U11131 ( .A1(n18040), .A2(b_in[55]), .ZN(n15484) );
NAND2_X2 U11132 ( .A1(n15513), .A2(n15514), .ZN(N3141) );
NAND2_X2 U11133 ( .A1(n15515), .A2(n18066), .ZN(n15514) );
XNOR2_X2 U11134 ( .A(n18965), .B(n15516), .ZN(n15515) );
XOR2_X2 U11138 ( .A(aes_text_out[70]), .B(n15520), .Z(n13700) );
AND4_X2 U11139 ( .A1(n15521), .A2(n15522), .A3(n15523), .A4(n15524), .ZN(n15520) );
NAND2_X2 U11148 ( .A1(n17848), .A2(dii_data[62]), .ZN(n15522) );
NAND2_X2 U11149 ( .A1(n15509), .A2(dii_data[6]), .ZN(n15521) );
NAND2_X2 U11151 ( .A1(n17906), .A2(dii_data[70]), .ZN(n15532) );
NAND2_X2 U11153 ( .A1(n17923), .A2(n15533), .ZN(n13698) );
XOR2_X2 U11154 ( .A(n17619), .B(aes_text_out[70]), .Z(n15533) );
NAND2_X2 U11155 ( .A1(n18040), .A2(b_in[54]), .ZN(n15513) );
NAND2_X2 U11156 ( .A1(n15534), .A2(n15535), .ZN(N3140) );
NAND2_X2 U11157 ( .A1(n15536), .A2(n18067), .ZN(n15535) );
XNOR2_X2 U11158 ( .A(n18964), .B(n15537), .ZN(n15536) );
XOR2_X2 U11162 ( .A(aes_text_out[69]), .B(n15541), .Z(n13694) );
AND4_X2 U11163 ( .A1(n15542), .A2(n15543), .A3(n15544), .A4(n15545), .ZN(n15541) );
NAND2_X2 U11172 ( .A1(n17848), .A2(dii_data[61]), .ZN(n15543) );
NAND2_X2 U11173 ( .A1(n15509), .A2(dii_data[5]), .ZN(n15542) );
NAND2_X2 U11175 ( .A1(n17906), .A2(dii_data[69]), .ZN(n15553) );
NAND2_X2 U11177 ( .A1(n17923), .A2(n15554), .ZN(n13692) );
XOR2_X2 U11178 ( .A(n17621), .B(aes_text_out[69]), .Z(n15554) );
NAND2_X2 U11179 ( .A1(n18040), .A2(b_in[53]), .ZN(n15534) );
NAND2_X2 U11180 ( .A1(n15555), .A2(n15556), .ZN(N3139) );
NAND2_X2 U11181 ( .A1(n15557), .A2(n18067), .ZN(n15556) );
XNOR2_X2 U11182 ( .A(n18963), .B(n15558), .ZN(n15557) );
XOR2_X2 U11186 ( .A(aes_text_out[68]), .B(n15562), .Z(n13688) );
AND4_X2 U11187 ( .A1(n15563), .A2(n15564), .A3(n15565), .A4(n15566), .ZN(n15562) );
NAND2_X2 U11196 ( .A1(n17848), .A2(dii_data[60]), .ZN(n15564) );
NAND2_X2 U11197 ( .A1(n15509), .A2(dii_data[4]), .ZN(n15563) );
NAND2_X2 U11199 ( .A1(n17906), .A2(dii_data[68]), .ZN(n15574) );
NAND2_X2 U11201 ( .A1(n17923), .A2(n15575), .ZN(n13686) );
XOR2_X2 U11202 ( .A(n17623), .B(aes_text_out[68]), .Z(n15575) );
NAND2_X2 U11203 ( .A1(n18040), .A2(b_in[52]), .ZN(n15555) );
NAND2_X2 U11204 ( .A1(n15576), .A2(n15577), .ZN(N3138) );
NAND2_X2 U11205 ( .A1(n15578), .A2(n18067), .ZN(n15577) );
XNOR2_X2 U11206 ( .A(n18962), .B(n15579), .ZN(n15578) );
XOR2_X2 U11210 ( .A(aes_text_out[67]), .B(n15583), .Z(n13682) );
AND4_X2 U11211 ( .A1(n15584), .A2(n15585), .A3(n15586), .A4(n15587), .ZN(n15583) );
NAND2_X2 U11220 ( .A1(n17848), .A2(dii_data[59]), .ZN(n15585) );
NAND2_X2 U11221 ( .A1(n15509), .A2(dii_data[3]), .ZN(n15584) );
NAND2_X2 U11223 ( .A1(n17906), .A2(dii_data[67]), .ZN(n15595) );
NAND2_X2 U11225 ( .A1(n17923), .A2(n15596), .ZN(n13680) );
XOR2_X2 U11226 ( .A(n17625), .B(aes_text_out[67]), .Z(n15596) );
NAND2_X2 U11227 ( .A1(n18040), .A2(b_in[51]), .ZN(n15576) );
NAND2_X2 U11228 ( .A1(n15597), .A2(n15598), .ZN(N3137) );
NAND2_X2 U11229 ( .A1(n15599), .A2(n18067), .ZN(n15598) );
XNOR2_X2 U11230 ( .A(n18961), .B(n15600), .ZN(n15599) );
AND2_X2 U11233 ( .A1(dii_data[66]), .A2(n17908), .ZN(n15603) );
XOR2_X2 U11235 ( .A(aes_text_out[66]), .B(n15605), .Z(n13676) );
AND4_X2 U11236 ( .A1(n15606), .A2(n15607), .A3(n15608), .A4(n15609), .ZN(n15605) );
OR2_X2 U11245 ( .A1(n17872), .A2(n19172), .ZN(n15607) );
NAND2_X2 U11246 ( .A1(n17848), .A2(dii_data[58]), .ZN(n15606) );
AND2_X2 U11247 ( .A1(n13675), .A2(n17930), .ZN(n15601) );
XOR2_X2 U11248 ( .A(aes_text_out[66]), .B(n17627), .Z(n13675) );
NAND2_X2 U11249 ( .A1(n18040), .A2(b_in[50]), .ZN(n15597) );
NAND2_X2 U11250 ( .A1(n15616), .A2(n15617), .ZN(N3136) );
NAND2_X2 U11251 ( .A1(n15618), .A2(n18067), .ZN(n15617) );
XNOR2_X2 U11252 ( .A(n18960), .B(n15619), .ZN(n15618) );
AND2_X2 U11255 ( .A1(dii_data[65]), .A2(n17908), .ZN(n15622) );
XOR2_X2 U11257 ( .A(aes_text_out[65]), .B(n15624), .Z(n13669) );
AND4_X2 U11258 ( .A1(n15625), .A2(n15626), .A3(n15627), .A4(n15628), .ZN(n15624) );
NAND2_X2 U11267 ( .A1(n17848), .A2(dii_data[57]), .ZN(n15626) );
NAND2_X2 U11268 ( .A1(n15509), .A2(dii_data[1]), .ZN(n15625) );
AND2_X2 U11269 ( .A1(n13668), .A2(n17930), .ZN(n15620) );
NAND2_X2 U11271 ( .A1(n18040), .A2(b_in[49]), .ZN(n15616) );
NAND2_X2 U11272 ( .A1(n15635), .A2(n15636), .ZN(N3135) );
NAND2_X2 U11273 ( .A1(n15637), .A2(n18067), .ZN(n15636) );
XNOR2_X2 U11274 ( .A(n18959), .B(n15638), .ZN(n15637) );
AND2_X2 U11277 ( .A1(dii_data[64]), .A2(n17908), .ZN(n15641) );
NAND2_X2 U11279 ( .A1(n17934), .A2(n19199), .ZN(n15492) );
XOR2_X2 U11281 ( .A(aes_text_out[64]), .B(n15643), .Z(n13662) );
AND4_X2 U11282 ( .A1(n15645), .A2(n15646), .A3(n15647), .A4(n15648), .ZN(n15643) );
NAND2_X2 U11291 ( .A1(n17848), .A2(dii_data[56]), .ZN(n15646) );
NAND2_X2 U11292 ( .A1(n15509), .A2(dii_data[0]), .ZN(n15645) );
AND2_X2 U11293 ( .A1(n13661), .A2(n17930), .ZN(n15639) );
XOR2_X2 U11294 ( .A(aes_text_out[64]), .B(n17631), .Z(n13661) );
NAND2_X2 U11295 ( .A1(n18040), .A2(b_in[48]), .ZN(n15635) );
NAND2_X2 U11296 ( .A1(n15655), .A2(n15656), .ZN(N3134) );
NAND2_X2 U11297 ( .A1(n15657), .A2(n18067), .ZN(n15656) );
XNOR2_X2 U11298 ( .A(n18958), .B(n15658), .ZN(n15657) );
XOR2_X2 U11302 ( .A(n15662), .B(aes_text_out[63]), .Z(n13654) );
AND4_X2 U11303 ( .A1(n15664), .A2(n15665), .A3(n15666), .A4(n15667), .ZN(n15662) );
NAND2_X2 U11309 ( .A1(n17848), .A2(dii_data[55]), .ZN(n15666) );
NAND2_X2 U11310 ( .A1(n17859), .A2(dii_data[39]), .ZN(n15665) );
NAND2_X2 U11311 ( .A1(n17852), .A2(dii_data[47]), .ZN(n15664) );
NAND2_X2 U11312 ( .A1(n15672), .A2(n15673), .ZN(n15659) );
NAND2_X2 U11313 ( .A1(n17906), .A2(dii_data[63]), .ZN(n15673) );
NAND2_X2 U11315 ( .A1(n17923), .A2(n15674), .ZN(n13652) );
XNOR2_X2 U11316 ( .A(n19135), .B(aes_text_out[63]), .ZN(n15674) );
NAND2_X2 U11317 ( .A1(n18040), .A2(b_in[47]), .ZN(n15655) );
NAND2_X2 U11318 ( .A1(n15675), .A2(n15676), .ZN(N3133) );
NAND2_X2 U11319 ( .A1(n15677), .A2(n18067), .ZN(n15676) );
XNOR2_X2 U11320 ( .A(n18957), .B(n15678), .ZN(n15677) );
XOR2_X2 U11324 ( .A(n15682), .B(aes_text_out[62]), .Z(n13648) );
AND4_X2 U11325 ( .A1(n15683), .A2(n15684), .A3(n15685), .A4(n15686), .ZN(n15682) );
NAND2_X2 U11331 ( .A1(n17849), .A2(dii_data[54]), .ZN(n15685) );
NAND2_X2 U11332 ( .A1(n17859), .A2(dii_data[38]), .ZN(n15684) );
NAND2_X2 U11333 ( .A1(n17852), .A2(dii_data[46]), .ZN(n15683) );
NAND2_X2 U11334 ( .A1(n15691), .A2(n15692), .ZN(n15679) );
NAND2_X2 U11335 ( .A1(n17906), .A2(dii_data[62]), .ZN(n15692) );
NAND2_X2 U11337 ( .A1(n17923), .A2(n15693), .ZN(n13646) );
XNOR2_X2 U11338 ( .A(n19136), .B(aes_text_out[62]), .ZN(n15693) );
NAND2_X2 U11339 ( .A1(n18040), .A2(b_in[46]), .ZN(n15675) );
NAND2_X2 U11340 ( .A1(n15694), .A2(n15695), .ZN(N3132) );
NAND2_X2 U11341 ( .A1(n15696), .A2(n18067), .ZN(n15695) );
XNOR2_X2 U11342 ( .A(n18956), .B(n15697), .ZN(n15696) );
XOR2_X2 U11346 ( .A(n15701), .B(aes_text_out[61]), .Z(n13642) );
AND4_X2 U11347 ( .A1(n15702), .A2(n15703), .A3(n15704), .A4(n15705), .ZN(n15701) );
NAND2_X2 U11353 ( .A1(n17849), .A2(dii_data[53]), .ZN(n15704) );
NAND2_X2 U11354 ( .A1(n17859), .A2(dii_data[37]), .ZN(n15703) );
NAND2_X2 U11355 ( .A1(n17852), .A2(dii_data[45]), .ZN(n15702) );
NAND2_X2 U11356 ( .A1(n15710), .A2(n15711), .ZN(n15698) );
NAND2_X2 U11357 ( .A1(n17906), .A2(dii_data[61]), .ZN(n15711) );
NAND2_X2 U11359 ( .A1(n17924), .A2(n15712), .ZN(n13640) );
XNOR2_X2 U11360 ( .A(n19137), .B(aes_text_out[61]), .ZN(n15712) );
NAND2_X2 U11361 ( .A1(n18040), .A2(b_in[45]), .ZN(n15694) );
NAND2_X2 U11362 ( .A1(n15713), .A2(n15714), .ZN(N3131) );
NAND2_X2 U11363 ( .A1(n15715), .A2(n18067), .ZN(n15714) );
XNOR2_X2 U11364 ( .A(n18955), .B(n15716), .ZN(n15715) );
XOR2_X2 U11368 ( .A(n15720), .B(aes_text_out[60]), .Z(n13636) );
AND4_X2 U11369 ( .A1(n15721), .A2(n15722), .A3(n15723), .A4(n15724), .ZN(n15720) );
NAND2_X2 U11375 ( .A1(n17849), .A2(dii_data[52]), .ZN(n15723) );
NAND2_X2 U11376 ( .A1(n17859), .A2(dii_data[36]), .ZN(n15722) );
NAND2_X2 U11377 ( .A1(n17852), .A2(dii_data[44]), .ZN(n15721) );
NAND2_X2 U11378 ( .A1(n15729), .A2(n15730), .ZN(n15717) );
NAND2_X2 U11379 ( .A1(n17906), .A2(dii_data[60]), .ZN(n15730) );
NAND2_X2 U11381 ( .A1(n17924), .A2(n15731), .ZN(n13634) );
XNOR2_X2 U11382 ( .A(n19138), .B(aes_text_out[60]), .ZN(n15731) );
NAND2_X2 U11383 ( .A1(n18039), .A2(b_in[44]), .ZN(n15713) );
NAND2_X2 U11384 ( .A1(n15732), .A2(n15733), .ZN(N3130) );
NAND2_X2 U11385 ( .A1(n15734), .A2(n18067), .ZN(n15733) );
XNOR2_X2 U11386 ( .A(n18954), .B(n15735), .ZN(n15734) );
XOR2_X2 U11390 ( .A(n15739), .B(aes_text_out[59]), .Z(n13630) );
AND4_X2 U11391 ( .A1(n15740), .A2(n15741), .A3(n15742), .A4(n15743), .ZN(n15739) );
NAND2_X2 U11397 ( .A1(n17849), .A2(dii_data[51]), .ZN(n15742) );
NAND2_X2 U11398 ( .A1(n17859), .A2(dii_data[35]), .ZN(n15741) );
NAND2_X2 U11399 ( .A1(n17852), .A2(dii_data[43]), .ZN(n15740) );
NAND2_X2 U11400 ( .A1(n15748), .A2(n15749), .ZN(n15736) );
NAND2_X2 U11401 ( .A1(n17906), .A2(dii_data[59]), .ZN(n15749) );
NAND2_X2 U11403 ( .A1(n17924), .A2(n15750), .ZN(n13628) );
XNOR2_X2 U11404 ( .A(n19139), .B(aes_text_out[59]), .ZN(n15750) );
NAND2_X2 U11405 ( .A1(n18039), .A2(b_in[43]), .ZN(n15732) );
NAND2_X2 U11406 ( .A1(n15751), .A2(n15752), .ZN(N3129) );
NAND2_X2 U11407 ( .A1(n15753), .A2(n18067), .ZN(n15752) );
XNOR2_X2 U11408 ( .A(n18953), .B(n15754), .ZN(n15753) );
XOR2_X2 U11412 ( .A(n15758), .B(aes_text_out[58]), .Z(n13624) );
AND4_X2 U11413 ( .A1(n15759), .A2(n15760), .A3(n15761), .A4(n15762), .ZN(n15758) );
NAND2_X2 U11419 ( .A1(n17849), .A2(dii_data[50]), .ZN(n15761) );
NAND2_X2 U11420 ( .A1(n17858), .A2(dii_data[34]), .ZN(n15760) );
NAND2_X2 U11421 ( .A1(n17852), .A2(dii_data[42]), .ZN(n15759) );
NAND2_X2 U11422 ( .A1(n15767), .A2(n15768), .ZN(n15755) );
NAND2_X2 U11423 ( .A1(n17906), .A2(dii_data[58]), .ZN(n15768) );
NAND2_X2 U11425 ( .A1(n17924), .A2(n15769), .ZN(n13622) );
XNOR2_X2 U11426 ( .A(n19140), .B(aes_text_out[58]), .ZN(n15769) );
NAND2_X2 U11427 ( .A1(n18039), .A2(b_in[42]), .ZN(n15751) );
NAND2_X2 U11428 ( .A1(n15770), .A2(n15771), .ZN(N3128) );
NAND2_X2 U11429 ( .A1(n15772), .A2(n18067), .ZN(n15771) );
XNOR2_X2 U11430 ( .A(n18952), .B(n15773), .ZN(n15772) );
XOR2_X2 U11434 ( .A(n15777), .B(aes_text_out[57]), .Z(n13618) );
AND4_X2 U11435 ( .A1(n15778), .A2(n15779), .A3(n15780), .A4(n15781), .ZN(n15777) );
NAND2_X2 U11441 ( .A1(n17849), .A2(dii_data[49]), .ZN(n15780) );
NAND2_X2 U11442 ( .A1(n17858), .A2(dii_data[33]), .ZN(n15779) );
NAND2_X2 U11443 ( .A1(n17852), .A2(dii_data[41]), .ZN(n15778) );
NAND2_X2 U11444 ( .A1(n15786), .A2(n15787), .ZN(n15774) );
NAND2_X2 U11445 ( .A1(n17906), .A2(dii_data[57]), .ZN(n15787) );
NAND2_X2 U11447 ( .A1(n17924), .A2(n15788), .ZN(n13616) );
XNOR2_X2 U11448 ( .A(n19141), .B(aes_text_out[57]), .ZN(n15788) );
NAND2_X2 U11449 ( .A1(n18039), .A2(b_in[41]), .ZN(n15770) );
NAND2_X2 U11450 ( .A1(n15789), .A2(n15790), .ZN(N3127) );
NAND2_X2 U11451 ( .A1(n15791), .A2(n18067), .ZN(n15790) );
XNOR2_X2 U11452 ( .A(n18951), .B(n15792), .ZN(n15791) );
XOR2_X2 U11456 ( .A(n15796), .B(aes_text_out[56]), .Z(n13612) );
AND4_X2 U11457 ( .A1(n15797), .A2(n15798), .A3(n15799), .A4(n15800), .ZN(n15796) );
NAND2_X2 U11463 ( .A1(n17849), .A2(dii_data[48]), .ZN(n15799) );
NAND2_X2 U11464 ( .A1(n17858), .A2(dii_data[32]), .ZN(n15798) );
NAND2_X2 U11465 ( .A1(n17852), .A2(dii_data[40]), .ZN(n15797) );
AND2_X2 U11467 ( .A1(n19202), .A2(n17945), .ZN(n15806) );
NAND2_X2 U11469 ( .A1(n15807), .A2(n15808), .ZN(n15793) );
NAND2_X2 U11470 ( .A1(n17906), .A2(dii_data[56]), .ZN(n15808) );
NAND2_X2 U11472 ( .A1(n17924), .A2(n15809), .ZN(n13610) );
XNOR2_X2 U11473 ( .A(n19142), .B(aes_text_out[56]), .ZN(n15809) );
NAND2_X2 U11474 ( .A1(n18039), .A2(b_in[40]), .ZN(n15789) );
NAND2_X2 U11475 ( .A1(n15810), .A2(n15811), .ZN(N3126) );
NAND2_X2 U11476 ( .A1(n15812), .A2(n18067), .ZN(n15811) );
XNOR2_X2 U11477 ( .A(n18950), .B(n15813), .ZN(n15812) );
NAND2_X2 U11481 ( .A1(n17924), .A2(n15817), .ZN(n13604) );
XNOR2_X2 U11482 ( .A(n19143), .B(aes_text_out[55]), .ZN(n15817) );
NAND2_X2 U11483 ( .A1(n15818), .A2(n15819), .ZN(n15814) );
NAND2_X2 U11484 ( .A1(n13606), .A2(n15805), .ZN(n15819) );
XOR2_X2 U11485 ( .A(n15820), .B(aes_text_out[55]), .Z(n13606) );
NAND2_X2 U11486 ( .A1(n17911), .A2(n15820), .ZN(n15818) );
NAND4_X2 U11487 ( .A1(n15821), .A2(n15822), .A3(n15823), .A4(n15824), .ZN(n15820) );
NAND2_X2 U11492 ( .A1(n17849), .A2(dii_data[47]), .ZN(n15823) );
NAND2_X2 U11493 ( .A1(n17858), .A2(dii_data[31]), .ZN(n15822) );
NAND2_X2 U11494 ( .A1(n17852), .A2(n17681), .ZN(n15821) );
NAND2_X2 U11495 ( .A1(n18039), .A2(b_in[39]), .ZN(n15810) );
NAND2_X2 U11496 ( .A1(n15828), .A2(n15829), .ZN(N3125) );
NAND2_X2 U11497 ( .A1(n15830), .A2(n18067), .ZN(n15829) );
XNOR2_X2 U11498 ( .A(n18949), .B(n15831), .ZN(n15830) );
NAND2_X2 U11502 ( .A1(n17924), .A2(n15835), .ZN(n13598) );
XNOR2_X2 U11503 ( .A(n19144), .B(aes_text_out[54]), .ZN(n15835) );
NAND2_X2 U11504 ( .A1(n15836), .A2(n15837), .ZN(n15832) );
NAND2_X2 U11505 ( .A1(n13600), .A2(n15805), .ZN(n15837) );
XOR2_X2 U11506 ( .A(n15838), .B(aes_text_out[54]), .Z(n13600) );
NAND2_X2 U11507 ( .A1(n17911), .A2(n15838), .ZN(n15836) );
NAND4_X2 U11508 ( .A1(n15839), .A2(n15840), .A3(n15841), .A4(n15842), .ZN(n15838) );
NAND2_X2 U11513 ( .A1(n17849), .A2(dii_data[46]), .ZN(n15841) );
NAND2_X2 U11514 ( .A1(n17858), .A2(dii_data[30]), .ZN(n15840) );
NAND2_X2 U11515 ( .A1(n17852), .A2(n17683), .ZN(n15839) );
NAND2_X2 U11516 ( .A1(n18039), .A2(b_in[38]), .ZN(n15828) );
NAND2_X2 U11517 ( .A1(n15846), .A2(n15847), .ZN(N3124) );
NAND2_X2 U11518 ( .A1(n15848), .A2(n18067), .ZN(n15847) );
XNOR2_X2 U11519 ( .A(n18948), .B(n15849), .ZN(n15848) );
NAND2_X2 U11523 ( .A1(n17924), .A2(n15853), .ZN(n13592) );
XNOR2_X2 U11524 ( .A(n19145), .B(aes_text_out[53]), .ZN(n15853) );
NAND2_X2 U11525 ( .A1(n15854), .A2(n15855), .ZN(n15850) );
NAND2_X2 U11526 ( .A1(n13594), .A2(n15805), .ZN(n15855) );
XOR2_X2 U11527 ( .A(n15856), .B(aes_text_out[53]), .Z(n13594) );
NAND2_X2 U11528 ( .A1(n17911), .A2(n15856), .ZN(n15854) );
NAND4_X2 U11529 ( .A1(n15857), .A2(n15858), .A3(n15859), .A4(n15860), .ZN(n15856) );
NAND2_X2 U11534 ( .A1(n17849), .A2(dii_data[45]), .ZN(n15859) );
NAND2_X2 U11535 ( .A1(n17858), .A2(dii_data[29]), .ZN(n15858) );
NAND2_X2 U11536 ( .A1(n17852), .A2(n17685), .ZN(n15857) );
NAND2_X2 U11537 ( .A1(n18039), .A2(b_in[37]), .ZN(n15846) );
NAND2_X2 U11538 ( .A1(n15864), .A2(n15865), .ZN(N3123) );
NAND2_X2 U11539 ( .A1(n15866), .A2(n18067), .ZN(n15865) );
XNOR2_X2 U11540 ( .A(n18947), .B(n15867), .ZN(n15866) );
NAND2_X2 U11544 ( .A1(n17925), .A2(n15871), .ZN(n13586) );
XNOR2_X2 U11545 ( .A(n19146), .B(aes_text_out[52]), .ZN(n15871) );
NAND2_X2 U11546 ( .A1(n15872), .A2(n15873), .ZN(n15868) );
NAND2_X2 U11547 ( .A1(n13588), .A2(n15805), .ZN(n15873) );
XOR2_X2 U11548 ( .A(n15874), .B(aes_text_out[52]), .Z(n13588) );
NAND2_X2 U11549 ( .A1(n17910), .A2(n15874), .ZN(n15872) );
NAND4_X2 U11550 ( .A1(n15875), .A2(n15876), .A3(n15877), .A4(n15878), .ZN(n15874) );
NAND2_X2 U11555 ( .A1(n17849), .A2(dii_data[44]), .ZN(n15877) );
NAND2_X2 U11556 ( .A1(n17858), .A2(dii_data[28]), .ZN(n15876) );
NAND2_X2 U11557 ( .A1(n17853), .A2(n17687), .ZN(n15875) );
NAND2_X2 U11558 ( .A1(n18039), .A2(b_in[36]), .ZN(n15864) );
NAND2_X2 U11559 ( .A1(n15882), .A2(n15883), .ZN(N3122) );
NAND2_X2 U11560 ( .A1(n15884), .A2(n18067), .ZN(n15883) );
XNOR2_X2 U11561 ( .A(n18946), .B(n15885), .ZN(n15884) );
NAND2_X2 U11565 ( .A1(n17925), .A2(n15889), .ZN(n13580) );
XNOR2_X2 U11566 ( .A(n19147), .B(aes_text_out[51]), .ZN(n15889) );
NAND2_X2 U11567 ( .A1(n15890), .A2(n15891), .ZN(n15886) );
NAND2_X2 U11568 ( .A1(n13582), .A2(n15805), .ZN(n15891) );
XOR2_X2 U11569 ( .A(n15892), .B(aes_text_out[51]), .Z(n13582) );
NAND2_X2 U11570 ( .A1(n17910), .A2(n15892), .ZN(n15890) );
NAND4_X2 U11571 ( .A1(n15893), .A2(n15894), .A3(n15895), .A4(n15896), .ZN(n15892) );
NAND2_X2 U11576 ( .A1(n17849), .A2(dii_data[43]), .ZN(n15895) );
NAND2_X2 U11577 ( .A1(n17858), .A2(dii_data[27]), .ZN(n15894) );
NAND2_X2 U11578 ( .A1(n17853), .A2(n17689), .ZN(n15893) );
NAND2_X2 U11579 ( .A1(n18039), .A2(b_in[35]), .ZN(n15882) );
NAND2_X2 U11580 ( .A1(n15900), .A2(n15901), .ZN(N3121) );
NAND2_X2 U11581 ( .A1(n15902), .A2(n18067), .ZN(n15901) );
XNOR2_X2 U11582 ( .A(n18945), .B(n15903), .ZN(n15902) );
NAND2_X2 U11586 ( .A1(n17925), .A2(n15907), .ZN(n13574) );
XNOR2_X2 U11587 ( .A(n19148), .B(aes_text_out[50]), .ZN(n15907) );
NAND2_X2 U11588 ( .A1(n15908), .A2(n15909), .ZN(n15904) );
NAND2_X2 U11589 ( .A1(n13576), .A2(n15805), .ZN(n15909) );
XOR2_X2 U11590 ( .A(n15910), .B(aes_text_out[50]), .Z(n13576) );
NAND2_X2 U11591 ( .A1(n17910), .A2(n15910), .ZN(n15908) );
NAND4_X2 U11592 ( .A1(n15911), .A2(n15912), .A3(n15913), .A4(n15914), .ZN(n15910) );
NAND2_X2 U11597 ( .A1(n17849), .A2(dii_data[42]), .ZN(n15913) );
NAND2_X2 U11598 ( .A1(n17858), .A2(dii_data[26]), .ZN(n15912) );
NAND2_X2 U11599 ( .A1(n17853), .A2(n17691), .ZN(n15911) );
NAND2_X2 U11600 ( .A1(n18039), .A2(b_in[34]), .ZN(n15900) );
NAND2_X2 U11601 ( .A1(n15918), .A2(n15919), .ZN(N3120) );
NAND2_X2 U11602 ( .A1(n15920), .A2(n18067), .ZN(n15919) );
XNOR2_X2 U11603 ( .A(n18944), .B(n15921), .ZN(n15920) );
NAND2_X2 U11607 ( .A1(n17925), .A2(n15925), .ZN(n13568) );
XNOR2_X2 U11608 ( .A(n19149), .B(aes_text_out[49]), .ZN(n15925) );
NAND2_X2 U11609 ( .A1(n15926), .A2(n15927), .ZN(n15922) );
NAND2_X2 U11610 ( .A1(n13570), .A2(n15805), .ZN(n15927) );
XOR2_X2 U11611 ( .A(n15928), .B(aes_text_out[49]), .Z(n13570) );
NAND2_X2 U11612 ( .A1(n17910), .A2(n15928), .ZN(n15926) );
NAND4_X2 U11613 ( .A1(n15929), .A2(n15930), .A3(n15931), .A4(n15932), .ZN(n15928) );
NAND2_X2 U11618 ( .A1(n17849), .A2(dii_data[41]), .ZN(n15931) );
NAND2_X2 U11619 ( .A1(n17858), .A2(dii_data[25]), .ZN(n15930) );
NAND2_X2 U11620 ( .A1(n17853), .A2(n17693), .ZN(n15929) );
NAND2_X2 U11621 ( .A1(n18039), .A2(b_in[33]), .ZN(n15918) );
NAND2_X2 U11622 ( .A1(n15936), .A2(n15937), .ZN(N3119) );
NAND2_X2 U11623 ( .A1(n15938), .A2(n18068), .ZN(n15937) );
XNOR2_X2 U11624 ( .A(n18943), .B(n15939), .ZN(n15938) );
NAND2_X2 U11628 ( .A1(n17925), .A2(n15943), .ZN(n13562) );
XNOR2_X2 U11629 ( .A(n19150), .B(aes_text_out[48]), .ZN(n15943) );
NAND2_X2 U11630 ( .A1(n15944), .A2(n15945), .ZN(n15940) );
NAND2_X2 U11631 ( .A1(n13564), .A2(n15805), .ZN(n15945) );
NAND2_X2 U11633 ( .A1(n17755), .A2(n17945), .ZN(n15947) );
XOR2_X2 U11634 ( .A(n15948), .B(aes_text_out[48]), .Z(n13564) );
NAND2_X2 U11635 ( .A1(n17910), .A2(n15948), .ZN(n15944) );
NAND4_X2 U11636 ( .A1(n15949), .A2(n15950), .A3(n15951), .A4(n15952), .ZN(n15948) );
NAND2_X2 U11643 ( .A1(n17849), .A2(dii_data[40]), .ZN(n15951) );
NAND2_X2 U11644 ( .A1(n17858), .A2(dii_data[24]), .ZN(n15950) );
NAND2_X2 U11645 ( .A1(n17853), .A2(n17695), .ZN(n15949) );
NAND2_X2 U11646 ( .A1(n18039), .A2(b_in[32]), .ZN(n15936) );
NAND2_X2 U11647 ( .A1(n15956), .A2(n15957), .ZN(N3118) );
NAND2_X2 U11648 ( .A1(n15958), .A2(n18068), .ZN(n15957) );
XNOR2_X2 U11649 ( .A(n18942), .B(n15959), .ZN(n15958) );
XOR2_X2 U11653 ( .A(n15963), .B(aes_text_out[47]), .Z(n13558) );
AND4_X2 U11654 ( .A1(n15964), .A2(n15965), .A3(n15966), .A4(n15967), .ZN(n15963) );
NAND2_X2 U11655 ( .A1(n17858), .A2(dii_data[23]), .ZN(n15967) );
NAND2_X2 U11659 ( .A1(n17853), .A2(dii_data[31]), .ZN(n15965) );
NAND2_X2 U11660 ( .A1(n17849), .A2(dii_data[39]), .ZN(n15964) );
NAND2_X2 U11661 ( .A1(n15970), .A2(n15971), .ZN(n15960) );
NAND2_X2 U11662 ( .A1(n17907), .A2(dii_data[47]), .ZN(n15971) );
NAND2_X2 U11663 ( .A1(n17998), .A2(enc_byte_cnt[44]), .ZN(n15970) );
NAND2_X2 U11664 ( .A1(n17924), .A2(n15972), .ZN(n13556) );
XNOR2_X2 U11665 ( .A(n19151), .B(aes_text_out[47]), .ZN(n15972) );
NAND2_X2 U11666 ( .A1(n18039), .A2(b_in[31]), .ZN(n15956) );
NAND2_X2 U11667 ( .A1(n15973), .A2(n15974), .ZN(N3117) );
NAND2_X2 U11668 ( .A1(n15975), .A2(n18068), .ZN(n15974) );
XNOR2_X2 U11669 ( .A(n18941), .B(n15976), .ZN(n15975) );
XOR2_X2 U11673 ( .A(n15980), .B(aes_text_out[46]), .Z(n13552) );
AND4_X2 U11674 ( .A1(n15981), .A2(n15982), .A3(n15983), .A4(n15984), .ZN(n15980) );
NAND2_X2 U11675 ( .A1(n17858), .A2(dii_data[22]), .ZN(n15984) );
NAND2_X2 U11679 ( .A1(n17853), .A2(dii_data[30]), .ZN(n15982) );
NAND2_X2 U11680 ( .A1(n17850), .A2(dii_data[38]), .ZN(n15981) );
NAND2_X2 U11681 ( .A1(n15987), .A2(n15988), .ZN(n15977) );
NAND2_X2 U11682 ( .A1(n17907), .A2(dii_data[46]), .ZN(n15988) );
NAND2_X2 U11683 ( .A1(n17998), .A2(enc_byte_cnt[43]), .ZN(n15987) );
NAND2_X2 U11684 ( .A1(n17925), .A2(n15989), .ZN(n13550) );
XNOR2_X2 U11685 ( .A(n19152), .B(aes_text_out[46]), .ZN(n15989) );
NAND2_X2 U11686 ( .A1(n18039), .A2(b_in[30]), .ZN(n15973) );
NAND2_X2 U11687 ( .A1(n15990), .A2(n15991), .ZN(N3116) );
NAND2_X2 U11688 ( .A1(n15992), .A2(n18068), .ZN(n15991) );
XNOR2_X2 U11689 ( .A(n18940), .B(n15993), .ZN(n15992) );
XOR2_X2 U11693 ( .A(n15997), .B(aes_text_out[45]), .Z(n13546) );
AND4_X2 U11694 ( .A1(n15998), .A2(n15999), .A3(n16000), .A4(n16001), .ZN(n15997) );
NAND2_X2 U11695 ( .A1(n17858), .A2(dii_data[21]), .ZN(n16001) );
NAND2_X2 U11699 ( .A1(n17853), .A2(dii_data[29]), .ZN(n15999) );
NAND2_X2 U11700 ( .A1(n17850), .A2(dii_data[37]), .ZN(n15998) );
NAND2_X2 U11701 ( .A1(n16004), .A2(n16005), .ZN(n15994) );
NAND2_X2 U11702 ( .A1(n17907), .A2(dii_data[45]), .ZN(n16005) );
NAND2_X2 U11703 ( .A1(n17998), .A2(enc_byte_cnt[42]), .ZN(n16004) );
NAND2_X2 U11704 ( .A1(n17925), .A2(n16006), .ZN(n13544) );
XNOR2_X2 U11705 ( .A(n19153), .B(aes_text_out[45]), .ZN(n16006) );
NAND2_X2 U11706 ( .A1(n18039), .A2(b_in[29]), .ZN(n15990) );
NAND2_X2 U11707 ( .A1(n16007), .A2(n16008), .ZN(N3115) );
NAND2_X2 U11708 ( .A1(n16009), .A2(n18068), .ZN(n16008) );
XNOR2_X2 U11709 ( .A(n18939), .B(n16010), .ZN(n16009) );
XOR2_X2 U11713 ( .A(n16014), .B(aes_text_out[44]), .Z(n13540) );
AND4_X2 U11714 ( .A1(n16015), .A2(n16016), .A3(n16017), .A4(n16018), .ZN(n16014) );
NAND2_X2 U11715 ( .A1(n17858), .A2(dii_data[20]), .ZN(n16018) );
NAND2_X2 U11719 ( .A1(n17853), .A2(dii_data[28]), .ZN(n16016) );
NAND2_X2 U11720 ( .A1(n17850), .A2(dii_data[36]), .ZN(n16015) );
NAND2_X2 U11721 ( .A1(n16021), .A2(n16022), .ZN(n16011) );
NAND2_X2 U11722 ( .A1(n17907), .A2(dii_data[44]), .ZN(n16022) );
NAND2_X2 U11723 ( .A1(n17998), .A2(enc_byte_cnt[41]), .ZN(n16021) );
NAND2_X2 U11724 ( .A1(n17925), .A2(n16023), .ZN(n13538) );
XNOR2_X2 U11725 ( .A(n19154), .B(aes_text_out[44]), .ZN(n16023) );
NAND2_X2 U11726 ( .A1(n18039), .A2(b_in[28]), .ZN(n16007) );
NAND2_X2 U11727 ( .A1(n16024), .A2(n16025), .ZN(N3114) );
NAND2_X2 U11728 ( .A1(n16026), .A2(n18068), .ZN(n16025) );
XNOR2_X2 U11729 ( .A(n18938), .B(n16027), .ZN(n16026) );
XOR2_X2 U11733 ( .A(n16031), .B(aes_text_out[43]), .Z(n13534) );
AND4_X2 U11734 ( .A1(n16032), .A2(n16033), .A3(n16034), .A4(n16035), .ZN(n16031) );
NAND2_X2 U11735 ( .A1(n17858), .A2(dii_data[19]), .ZN(n16035) );
NAND2_X2 U11739 ( .A1(n17853), .A2(dii_data[27]), .ZN(n16033) );
NAND2_X2 U11740 ( .A1(n17850), .A2(dii_data[35]), .ZN(n16032) );
NAND2_X2 U11741 ( .A1(n16038), .A2(n16039), .ZN(n16028) );
NAND2_X2 U11742 ( .A1(n17907), .A2(dii_data[43]), .ZN(n16039) );
NAND2_X2 U11743 ( .A1(n17998), .A2(enc_byte_cnt[40]), .ZN(n16038) );
NAND2_X2 U11744 ( .A1(n17925), .A2(n16040), .ZN(n13532) );
XNOR2_X2 U11745 ( .A(n19155), .B(aes_text_out[43]), .ZN(n16040) );
NAND2_X2 U11746 ( .A1(n18038), .A2(b_in[27]), .ZN(n16024) );
NAND2_X2 U11747 ( .A1(n16041), .A2(n16042), .ZN(N3113) );
NAND2_X2 U11748 ( .A1(n16043), .A2(n18068), .ZN(n16042) );
XNOR2_X2 U11749 ( .A(n18937), .B(n16044), .ZN(n16043) );
XOR2_X2 U11753 ( .A(n16048), .B(aes_text_out[42]), .Z(n13528) );
AND4_X2 U11754 ( .A1(n16049), .A2(n16050), .A3(n16051), .A4(n16052), .ZN(n16048) );
NAND2_X2 U11755 ( .A1(n17858), .A2(dii_data[18]), .ZN(n16052) );
NAND2_X2 U11759 ( .A1(n17853), .A2(dii_data[26]), .ZN(n16050) );
NAND2_X2 U11760 ( .A1(n17850), .A2(dii_data[34]), .ZN(n16049) );
NAND2_X2 U11761 ( .A1(n16055), .A2(n16056), .ZN(n16045) );
NAND2_X2 U11762 ( .A1(n17907), .A2(dii_data[42]), .ZN(n16056) );
NAND2_X2 U11763 ( .A1(n17998), .A2(enc_byte_cnt[39]), .ZN(n16055) );
NAND2_X2 U11764 ( .A1(n17926), .A2(n16057), .ZN(n13526) );
XNOR2_X2 U11765 ( .A(n19156), .B(aes_text_out[42]), .ZN(n16057) );
NAND2_X2 U11766 ( .A1(n18038), .A2(b_in[26]), .ZN(n16041) );
NAND2_X2 U11767 ( .A1(n16058), .A2(n16059), .ZN(N3112) );
NAND2_X2 U11768 ( .A1(n16060), .A2(n18068), .ZN(n16059) );
XNOR2_X2 U11769 ( .A(n18936), .B(n16061), .ZN(n16060) );
XOR2_X2 U11773 ( .A(n16065), .B(aes_text_out[41]), .Z(n13522) );
AND4_X2 U11774 ( .A1(n16066), .A2(n16067), .A3(n16068), .A4(n16069), .ZN(n16065) );
NAND2_X2 U11775 ( .A1(n17858), .A2(dii_data[17]), .ZN(n16069) );
NAND2_X2 U11779 ( .A1(n17854), .A2(dii_data[25]), .ZN(n16067) );
NAND2_X2 U11780 ( .A1(n17850), .A2(dii_data[33]), .ZN(n16066) );
NAND2_X2 U11781 ( .A1(n16072), .A2(n16073), .ZN(n16062) );
NAND2_X2 U11782 ( .A1(n17907), .A2(dii_data[41]), .ZN(n16073) );
NAND2_X2 U11783 ( .A1(n17998), .A2(enc_byte_cnt[38]), .ZN(n16072) );
NAND2_X2 U11784 ( .A1(n17925), .A2(n16074), .ZN(n13520) );
XNOR2_X2 U11785 ( .A(n19157), .B(aes_text_out[41]), .ZN(n16074) );
NAND2_X2 U11786 ( .A1(n18038), .A2(b_in[25]), .ZN(n16058) );
NAND2_X2 U11787 ( .A1(n16075), .A2(n16076), .ZN(N3111) );
NAND2_X2 U11788 ( .A1(n16077), .A2(n18068), .ZN(n16076) );
XNOR2_X2 U11789 ( .A(n18935), .B(n16078), .ZN(n16077) );
NAND4_X2 U11794 ( .A1(n17872), .A2(n17876), .A3(n16083), .A4(n15507), .ZN(n15644) );
XOR2_X2 U11796 ( .A(n16082), .B(aes_text_out[40]), .Z(n13516) );
AND4_X2 U11797 ( .A1(n16084), .A2(n16085), .A3(n16086), .A4(n16087), .ZN(n16082) );
NAND2_X2 U11798 ( .A1(n17857), .A2(dii_data[16]), .ZN(n16087) );
NAND2_X2 U11804 ( .A1(n17854), .A2(dii_data[24]), .ZN(n16085) );
NAND2_X2 U11805 ( .A1(n17850), .A2(dii_data[32]), .ZN(n16084) );
NAND2_X2 U11806 ( .A1(n16090), .A2(n16091), .ZN(n16079) );
NAND2_X2 U11807 ( .A1(n17907), .A2(dii_data[40]), .ZN(n16091) );
NAND2_X2 U11808 ( .A1(n17998), .A2(enc_byte_cnt[37]), .ZN(n16090) );
NAND2_X2 U11809 ( .A1(n17926), .A2(n16092), .ZN(n13514) );
XNOR2_X2 U11810 ( .A(n19158), .B(aes_text_out[40]), .ZN(n16092) );
NAND2_X2 U11811 ( .A1(n18038), .A2(b_in[24]), .ZN(n16075) );
NAND2_X2 U11812 ( .A1(n16093), .A2(n16094), .ZN(N3110) );
NAND2_X2 U11813 ( .A1(n16095), .A2(n18068), .ZN(n16094) );
XNOR2_X2 U11814 ( .A(n18934), .B(n16096), .ZN(n16095) );
NAND2_X2 U11818 ( .A1(n17926), .A2(n16100), .ZN(n13508) );
XNOR2_X2 U11819 ( .A(n19159), .B(aes_text_out[39]), .ZN(n16100) );
NAND2_X2 U11820 ( .A1(n16101), .A2(n16102), .ZN(n16097) );
NAND2_X2 U11821 ( .A1(n13510), .A2(n16103), .ZN(n16102) );
XOR2_X2 U11822 ( .A(n16104), .B(aes_text_out[39]), .Z(n13510) );
NAND2_X2 U11823 ( .A1(n17910), .A2(n16104), .ZN(n16101) );
NAND4_X2 U11824 ( .A1(n16105), .A2(n16106), .A3(n16107), .A4(n16108), .ZN(n16104) );
NAND2_X2 U11825 ( .A1(n17873), .A2(dii_data[7]), .ZN(n16108) );
NAND2_X2 U11826 ( .A1(n17857), .A2(dii_data[15]), .ZN(n16107) );
NAND2_X2 U11827 ( .A1(n17854), .A2(dii_data[23]), .ZN(n16106) );
NAND2_X2 U11828 ( .A1(n17850), .A2(n17697), .ZN(n16105) );
NAND2_X2 U11829 ( .A1(n18038), .A2(b_in[23]), .ZN(n16093) );
NAND2_X2 U11830 ( .A1(n16109), .A2(n16110), .ZN(N3109) );
NAND2_X2 U11831 ( .A1(n16111), .A2(n18068), .ZN(n16110) );
XNOR2_X2 U11832 ( .A(n18933), .B(n16112), .ZN(n16111) );
NAND2_X2 U11836 ( .A1(n17926), .A2(n16116), .ZN(n13502) );
XNOR2_X2 U11837 ( .A(n19160), .B(aes_text_out[38]), .ZN(n16116) );
NAND2_X2 U11838 ( .A1(n16117), .A2(n16118), .ZN(n16113) );
NAND2_X2 U11839 ( .A1(n13504), .A2(n16103), .ZN(n16118) );
XOR2_X2 U11840 ( .A(n16119), .B(aes_text_out[38]), .Z(n13504) );
NAND2_X2 U11841 ( .A1(n17910), .A2(n16119), .ZN(n16117) );
NAND4_X2 U11842 ( .A1(n16120), .A2(n16121), .A3(n16122), .A4(n16123), .ZN(n16119) );
NAND2_X2 U11843 ( .A1(n17873), .A2(dii_data[6]), .ZN(n16123) );
NAND2_X2 U11844 ( .A1(n17857), .A2(dii_data[14]), .ZN(n16122) );
NAND2_X2 U11845 ( .A1(n17854), .A2(dii_data[22]), .ZN(n16121) );
NAND2_X2 U11846 ( .A1(n17850), .A2(n17699), .ZN(n16120) );
NAND2_X2 U11847 ( .A1(n18038), .A2(b_in[22]), .ZN(n16109) );
NAND2_X2 U11848 ( .A1(n16124), .A2(n16125), .ZN(N3108) );
NAND2_X2 U11849 ( .A1(n16126), .A2(n18068), .ZN(n16125) );
XNOR2_X2 U11850 ( .A(n18932), .B(n16127), .ZN(n16126) );
NAND2_X2 U11854 ( .A1(n17926), .A2(n16131), .ZN(n13496) );
XNOR2_X2 U11855 ( .A(n19161), .B(aes_text_out[37]), .ZN(n16131) );
NAND2_X2 U11856 ( .A1(n16132), .A2(n16133), .ZN(n16128) );
NAND2_X2 U11857 ( .A1(n13498), .A2(n16103), .ZN(n16133) );
XOR2_X2 U11858 ( .A(n16134), .B(aes_text_out[37]), .Z(n13498) );
NAND2_X2 U11859 ( .A1(n17910), .A2(n16134), .ZN(n16132) );
NAND4_X2 U11860 ( .A1(n16135), .A2(n16136), .A3(n16137), .A4(n16138), .ZN(n16134) );
NAND2_X2 U11861 ( .A1(n17873), .A2(dii_data[5]), .ZN(n16138) );
NAND2_X2 U11862 ( .A1(n17857), .A2(dii_data[13]), .ZN(n16137) );
NAND2_X2 U11863 ( .A1(n17854), .A2(dii_data[21]), .ZN(n16136) );
NAND2_X2 U11864 ( .A1(n17850), .A2(n17701), .ZN(n16135) );
NAND2_X2 U11865 ( .A1(n18038), .A2(b_in[21]), .ZN(n16124) );
NAND2_X2 U11866 ( .A1(n16139), .A2(n16140), .ZN(N3107) );
NAND2_X2 U11867 ( .A1(n16141), .A2(n18068), .ZN(n16140) );
XNOR2_X2 U11868 ( .A(n18931), .B(n16142), .ZN(n16141) );
NAND2_X2 U11872 ( .A1(n17926), .A2(n16146), .ZN(n13490) );
XNOR2_X2 U11873 ( .A(n19162), .B(aes_text_out[36]), .ZN(n16146) );
NAND2_X2 U11874 ( .A1(n16147), .A2(n16148), .ZN(n16143) );
NAND2_X2 U11875 ( .A1(n13492), .A2(n16103), .ZN(n16148) );
XOR2_X2 U11876 ( .A(n16149), .B(aes_text_out[36]), .Z(n13492) );
NAND2_X2 U11877 ( .A1(n17910), .A2(n16149), .ZN(n16147) );
NAND4_X2 U11878 ( .A1(n16150), .A2(n16151), .A3(n16152), .A4(n16153), .ZN(n16149) );
NAND2_X2 U11879 ( .A1(n17873), .A2(dii_data[4]), .ZN(n16153) );
NAND2_X2 U11880 ( .A1(n17857), .A2(dii_data[12]), .ZN(n16152) );
NAND2_X2 U11881 ( .A1(n17854), .A2(dii_data[20]), .ZN(n16151) );
NAND2_X2 U11882 ( .A1(n17850), .A2(n17703), .ZN(n16150) );
NAND2_X2 U11883 ( .A1(n18038), .A2(b_in[20]), .ZN(n16139) );
NAND2_X2 U11884 ( .A1(n16154), .A2(n16155), .ZN(N3106) );
NAND2_X2 U11885 ( .A1(n16156), .A2(n18068), .ZN(n16155) );
XNOR2_X2 U11886 ( .A(n18930), .B(n16157), .ZN(n16156) );
NAND2_X2 U11890 ( .A1(n17925), .A2(n16161), .ZN(n13484) );
XNOR2_X2 U11891 ( .A(n19163), .B(aes_text_out[35]), .ZN(n16161) );
NAND2_X2 U11892 ( .A1(n16162), .A2(n16163), .ZN(n16158) );
NAND2_X2 U11893 ( .A1(n13486), .A2(n16103), .ZN(n16163) );
XOR2_X2 U11894 ( .A(n16164), .B(aes_text_out[35]), .Z(n13486) );
NAND2_X2 U11895 ( .A1(n17910), .A2(n16164), .ZN(n16162) );
NAND4_X2 U11896 ( .A1(n16165), .A2(n16166), .A3(n16167), .A4(n16168), .ZN(n16164) );
NAND2_X2 U11897 ( .A1(n17873), .A2(dii_data[3]), .ZN(n16168) );
NAND2_X2 U11898 ( .A1(n17858), .A2(dii_data[11]), .ZN(n16167) );
NAND2_X2 U11899 ( .A1(n17854), .A2(dii_data[19]), .ZN(n16166) );
NAND2_X2 U11900 ( .A1(n17850), .A2(n17705), .ZN(n16165) );
NAND2_X2 U11901 ( .A1(n18038), .A2(b_in[19]), .ZN(n16154) );
NAND2_X2 U11902 ( .A1(n16169), .A2(n16170), .ZN(N3105) );
NAND2_X2 U11903 ( .A1(n16171), .A2(n18068), .ZN(n16170) );
XNOR2_X2 U11904 ( .A(n18929), .B(n16172), .ZN(n16171) );
NAND2_X2 U11908 ( .A1(n17926), .A2(n16176), .ZN(n13478) );
XNOR2_X2 U11909 ( .A(n19164), .B(aes_text_out[34]), .ZN(n16176) );
NAND2_X2 U11910 ( .A1(n16177), .A2(n16178), .ZN(n16173) );
NAND2_X2 U11911 ( .A1(n13480), .A2(n16103), .ZN(n16178) );
XOR2_X2 U11912 ( .A(n16179), .B(aes_text_out[34]), .Z(n13480) );
NAND2_X2 U11913 ( .A1(n17910), .A2(n16179), .ZN(n16177) );
NAND4_X2 U11914 ( .A1(n16180), .A2(n16181), .A3(n16182), .A4(n16183), .ZN(n16179) );
NAND2_X2 U11915 ( .A1(n17873), .A2(dii_data[2]), .ZN(n16183) );
NAND2_X2 U11916 ( .A1(n17857), .A2(dii_data[10]), .ZN(n16182) );
NAND2_X2 U11917 ( .A1(n17854), .A2(dii_data[18]), .ZN(n16181) );
NAND2_X2 U11918 ( .A1(n17850), .A2(n17707), .ZN(n16180) );
NAND2_X2 U11919 ( .A1(n18038), .A2(b_in[18]), .ZN(n16169) );
NAND2_X2 U11920 ( .A1(n16184), .A2(n16185), .ZN(N3104) );
NAND2_X2 U11921 ( .A1(n16186), .A2(n18068), .ZN(n16185) );
XNOR2_X2 U11922 ( .A(n18928), .B(n16187), .ZN(n16186) );
NAND2_X2 U11926 ( .A1(n17926), .A2(n16191), .ZN(n13472) );
XNOR2_X2 U11927 ( .A(n19165), .B(aes_text_out[33]), .ZN(n16191) );
NAND2_X2 U11928 ( .A1(n16192), .A2(n16193), .ZN(n16188) );
NAND2_X2 U11929 ( .A1(n13474), .A2(n16103), .ZN(n16193) );
XOR2_X2 U11930 ( .A(n16194), .B(aes_text_out[33]), .Z(n13474) );
NAND2_X2 U11931 ( .A1(n17909), .A2(n16194), .ZN(n16192) );
NAND4_X2 U11932 ( .A1(n16195), .A2(n16196), .A3(n16197), .A4(n16198), .ZN(n16194) );
NAND2_X2 U11933 ( .A1(n17873), .A2(dii_data[1]), .ZN(n16198) );
NAND2_X2 U11934 ( .A1(n17857), .A2(dii_data[9]), .ZN(n16197) );
NAND2_X2 U11935 ( .A1(n17854), .A2(dii_data[17]), .ZN(n16196) );
NAND2_X2 U11936 ( .A1(n17850), .A2(n17709), .ZN(n16195) );
NAND2_X2 U11937 ( .A1(n18038), .A2(b_in[17]), .ZN(n16184) );
NAND2_X2 U11938 ( .A1(n16199), .A2(n16200), .ZN(N3103) );
NAND2_X2 U11939 ( .A1(n16201), .A2(n18068), .ZN(n16200) );
XNOR2_X2 U11940 ( .A(n18927), .B(n16202), .ZN(n16201) );
NAND2_X2 U11944 ( .A1(n17926), .A2(n16206), .ZN(n13466) );
XNOR2_X2 U11945 ( .A(n19166), .B(aes_text_out[32]), .ZN(n16206) );
NAND2_X2 U11946 ( .A1(n16207), .A2(n16208), .ZN(n16203) );
NAND2_X2 U11947 ( .A1(n13468), .A2(n16103), .ZN(n16208) );
NAND2_X2 U11948 ( .A1(n16209), .A2(n16210), .ZN(n16103) );
NAND2_X2 U11949 ( .A1(n17873), .A2(n17945), .ZN(n16210) );
XOR2_X2 U11950 ( .A(n16211), .B(aes_text_out[32]), .Z(n13468) );
NAND2_X2 U11951 ( .A1(n17909), .A2(n16211), .ZN(n16207) );
NAND4_X2 U11952 ( .A1(n16212), .A2(n16213), .A3(n16214), .A4(n16215), .ZN(n16211) );
NAND2_X2 U11953 ( .A1(n17873), .A2(dii_data[0]), .ZN(n16215) );
NAND2_X2 U11954 ( .A1(n17897), .A2(n18074), .ZN(n15501) );
NAND2_X2 U11956 ( .A1(n17857), .A2(dii_data[8]), .ZN(n16214) );
NAND2_X2 U11957 ( .A1(n17854), .A2(dii_data[16]), .ZN(n16213) );
NAND2_X2 U11958 ( .A1(n17850), .A2(n17711), .ZN(n16212) );
NAND2_X2 U11959 ( .A1(n18040), .A2(b_in[16]), .ZN(n16199) );
NAND2_X2 U11960 ( .A1(n16216), .A2(n16217), .ZN(N3102) );
NAND2_X2 U11961 ( .A1(n16218), .A2(n18068), .ZN(n16217) );
XNOR2_X2 U11962 ( .A(n18926), .B(n16219), .ZN(n16218) );
XOR2_X2 U11966 ( .A(n16223), .B(aes_text_out[31]), .Z(n13462) );
AND3_X2 U11967 ( .A1(n16224), .A2(n16225), .A3(n16226), .ZN(n16223) );
NAND2_X2 U11968 ( .A1(n17850), .A2(dii_data[23]), .ZN(n16226) );
NAND2_X2 U11969 ( .A1(n17857), .A2(dii_data[7]), .ZN(n16225) );
NAND2_X2 U11970 ( .A1(n17854), .A2(dii_data[15]), .ZN(n16224) );
NAND2_X2 U11971 ( .A1(n16227), .A2(n16228), .ZN(n16220) );
NAND2_X2 U11972 ( .A1(n17907), .A2(dii_data[31]), .ZN(n16228) );
NAND2_X2 U11973 ( .A1(n17998), .A2(enc_byte_cnt[28]), .ZN(n16227) );
NAND2_X2 U11974 ( .A1(n17926), .A2(n16229), .ZN(n13460) );
XNOR2_X2 U11975 ( .A(n19167), .B(aes_text_out[31]), .ZN(n16229) );
NAND2_X2 U11976 ( .A1(n18038), .A2(b_in[15]), .ZN(n16216) );
NAND2_X2 U11977 ( .A1(n16230), .A2(n16231), .ZN(N3101) );
NAND2_X2 U11978 ( .A1(n16232), .A2(n18068), .ZN(n16231) );
XNOR2_X2 U11979 ( .A(n18925), .B(n16233), .ZN(n16232) );
XOR2_X2 U11983 ( .A(n16237), .B(aes_text_out[30]), .Z(n13456) );
AND3_X2 U11984 ( .A1(n16238), .A2(n16239), .A3(n16240), .ZN(n16237) );
NAND2_X2 U11985 ( .A1(n17850), .A2(dii_data[22]), .ZN(n16240) );
NAND2_X2 U11986 ( .A1(n17857), .A2(dii_data[6]), .ZN(n16239) );
NAND2_X2 U11987 ( .A1(n17855), .A2(dii_data[14]), .ZN(n16238) );
NAND2_X2 U11988 ( .A1(n16241), .A2(n16242), .ZN(n16234) );
NAND2_X2 U11989 ( .A1(n17907), .A2(dii_data[30]), .ZN(n16242) );
NAND2_X2 U11990 ( .A1(n17998), .A2(enc_byte_cnt[27]), .ZN(n16241) );
NAND2_X2 U11991 ( .A1(n17927), .A2(n16243), .ZN(n13454) );
XNOR2_X2 U11992 ( .A(n19168), .B(aes_text_out[30]), .ZN(n16243) );
NAND2_X2 U11993 ( .A1(n18038), .A2(b_in[14]), .ZN(n16230) );
NAND2_X2 U11994 ( .A1(n16244), .A2(n16245), .ZN(N3100) );
NAND2_X2 U11995 ( .A1(n16246), .A2(n18068), .ZN(n16245) );
XNOR2_X2 U11996 ( .A(n18924), .B(n16247), .ZN(n16246) );
XOR2_X2 U12000 ( .A(n16251), .B(aes_text_out[29]), .Z(n13450) );
AND3_X2 U12001 ( .A1(n16252), .A2(n16253), .A3(n16254), .ZN(n16251) );
NAND2_X2 U12002 ( .A1(n17851), .A2(dii_data[21]), .ZN(n16254) );
NAND2_X2 U12003 ( .A1(n17857), .A2(dii_data[5]), .ZN(n16253) );
NAND2_X2 U12004 ( .A1(n17855), .A2(dii_data[13]), .ZN(n16252) );
NAND2_X2 U12005 ( .A1(n16255), .A2(n16256), .ZN(n16248) );
NAND2_X2 U12006 ( .A1(n17907), .A2(dii_data[29]), .ZN(n16256) );
NAND2_X2 U12007 ( .A1(n17998), .A2(enc_byte_cnt[26]), .ZN(n16255) );
NAND2_X2 U12008 ( .A1(n17926), .A2(n16257), .ZN(n13448) );
XNOR2_X2 U12009 ( .A(n19169), .B(aes_text_out[29]), .ZN(n16257) );
NAND2_X2 U12010 ( .A1(n18038), .A2(b_in[13]), .ZN(n16244) );
NAND2_X2 U12011 ( .A1(n16258), .A2(n16259), .ZN(N3099) );
NAND2_X2 U12012 ( .A1(n16260), .A2(n18068), .ZN(n16259) );
XNOR2_X2 U12013 ( .A(n18923), .B(n16261), .ZN(n16260) );
XOR2_X2 U12017 ( .A(n16265), .B(aes_text_out[28]), .Z(n13444) );
AND3_X2 U12018 ( .A1(n16266), .A2(n16267), .A3(n16268), .ZN(n16265) );
NAND2_X2 U12019 ( .A1(n17851), .A2(dii_data[20]), .ZN(n16268) );
NAND2_X2 U12020 ( .A1(n17857), .A2(dii_data[4]), .ZN(n16267) );
NAND2_X2 U12021 ( .A1(n17855), .A2(dii_data[12]), .ZN(n16266) );
NAND2_X2 U12022 ( .A1(n16269), .A2(n16270), .ZN(n16262) );
NAND2_X2 U12023 ( .A1(n17907), .A2(dii_data[28]), .ZN(n16270) );
NAND2_X2 U12024 ( .A1(n17998), .A2(enc_byte_cnt[25]), .ZN(n16269) );
NAND2_X2 U12025 ( .A1(n17927), .A2(n16271), .ZN(n13442) );
XNOR2_X2 U12026 ( .A(n19170), .B(aes_text_out[28]), .ZN(n16271) );
NAND2_X2 U12027 ( .A1(n18038), .A2(b_in[12]), .ZN(n16258) );
NAND2_X2 U12028 ( .A1(n16272), .A2(n16273), .ZN(N3098) );
NAND2_X2 U12029 ( .A1(n16274), .A2(n18069), .ZN(n16273) );
XNOR2_X2 U12030 ( .A(n18922), .B(n16275), .ZN(n16274) );
XOR2_X2 U12034 ( .A(n16279), .B(aes_text_out[27]), .Z(n13438) );
AND3_X2 U12035 ( .A1(n16280), .A2(n16281), .A3(n16282), .ZN(n16279) );
NAND2_X2 U12036 ( .A1(n17851), .A2(dii_data[19]), .ZN(n16282) );
NAND2_X2 U12037 ( .A1(n17857), .A2(dii_data[3]), .ZN(n16281) );
NAND2_X2 U12038 ( .A1(n17855), .A2(dii_data[11]), .ZN(n16280) );
NAND2_X2 U12039 ( .A1(n16283), .A2(n16284), .ZN(n16276) );
NAND2_X2 U12040 ( .A1(n17907), .A2(dii_data[27]), .ZN(n16284) );
NAND2_X2 U12041 ( .A1(n17998), .A2(enc_byte_cnt[24]), .ZN(n16283) );
NAND2_X2 U12042 ( .A1(n17927), .A2(n16285), .ZN(n13436) );
XNOR2_X2 U12043 ( .A(n19171), .B(aes_text_out[27]), .ZN(n16285) );
NAND2_X2 U12044 ( .A1(n18038), .A2(b_in[11]), .ZN(n16272) );
NAND2_X2 U12045 ( .A1(n16286), .A2(n16287), .ZN(N3097) );
NAND2_X2 U12046 ( .A1(n16288), .A2(n18069), .ZN(n16287) );
XNOR2_X2 U12047 ( .A(n18921), .B(n16289), .ZN(n16288) );
XOR2_X2 U12051 ( .A(n16293), .B(aes_text_out[26]), .Z(n13432) );
AND3_X2 U12052 ( .A1(n16294), .A2(n16295), .A3(n16296), .ZN(n16293) );
NAND2_X2 U12053 ( .A1(n17851), .A2(dii_data[18]), .ZN(n16296) );
NAND2_X2 U12054 ( .A1(n17857), .A2(dii_data[2]), .ZN(n16295) );
NAND2_X2 U12055 ( .A1(n17855), .A2(dii_data[10]), .ZN(n16294) );
NAND2_X2 U12056 ( .A1(n16297), .A2(n16298), .ZN(n16290) );
NAND2_X2 U12057 ( .A1(n17907), .A2(dii_data[26]), .ZN(n16298) );
NAND2_X2 U12058 ( .A1(n17999), .A2(enc_byte_cnt[23]), .ZN(n16297) );
NAND2_X2 U12059 ( .A1(n17927), .A2(n16299), .ZN(n13430) );
XNOR2_X2 U12060 ( .A(n19172), .B(aes_text_out[26]), .ZN(n16299) );
NAND2_X2 U12061 ( .A1(n18038), .A2(b_in[10]), .ZN(n16286) );
NAND2_X2 U12062 ( .A1(n16300), .A2(n16301), .ZN(N3096) );
NAND2_X2 U12063 ( .A1(n16302), .A2(n18069), .ZN(n16301) );
XNOR2_X2 U12064 ( .A(n18920), .B(n16303), .ZN(n16302) );
XOR2_X2 U12068 ( .A(n16307), .B(aes_text_out[25]), .Z(n13426) );
AND3_X2 U12069 ( .A1(n16308), .A2(n16309), .A3(n16310), .ZN(n16307) );
NAND2_X2 U12070 ( .A1(n17851), .A2(dii_data[17]), .ZN(n16310) );
NAND2_X2 U12071 ( .A1(n17857), .A2(dii_data[1]), .ZN(n16309) );
NAND2_X2 U12072 ( .A1(n17855), .A2(dii_data[9]), .ZN(n16308) );
NAND2_X2 U12073 ( .A1(n16311), .A2(n16312), .ZN(n16304) );
NAND2_X2 U12074 ( .A1(n17907), .A2(dii_data[25]), .ZN(n16312) );
NAND2_X2 U12075 ( .A1(n17999), .A2(enc_byte_cnt[22]), .ZN(n16311) );
NAND2_X2 U12076 ( .A1(n17927), .A2(n16313), .ZN(n13424) );
XNOR2_X2 U12077 ( .A(n19173), .B(aes_text_out[25]), .ZN(n16313) );
NAND2_X2 U12078 ( .A1(n18037), .A2(b_in[9]), .ZN(n16300) );
NAND2_X2 U12079 ( .A1(n16314), .A2(n16315), .ZN(N3095) );
NAND2_X2 U12080 ( .A1(n16316), .A2(n18069), .ZN(n16315) );
XNOR2_X2 U12081 ( .A(n18919), .B(n16317), .ZN(n16316) );
XOR2_X2 U12085 ( .A(n16321), .B(aes_text_out[24]), .Z(n13420) );
AND3_X2 U12086 ( .A1(n16322), .A2(n16323), .A3(n16324), .ZN(n16321) );
NAND2_X2 U12087 ( .A1(n17851), .A2(dii_data[16]), .ZN(n16324) );
NAND2_X2 U12088 ( .A1(n17857), .A2(dii_data[0]), .ZN(n16323) );
NAND2_X2 U12089 ( .A1(n17855), .A2(dii_data[8]), .ZN(n16322) );
AND2_X2 U12091 ( .A1(n17859), .A2(n17945), .ZN(n16326) );
NAND2_X2 U12094 ( .A1(n16327), .A2(n16328), .ZN(n16318) );
NAND2_X2 U12095 ( .A1(n17907), .A2(dii_data[24]), .ZN(n16328) );
NAND2_X2 U12096 ( .A1(n17999), .A2(enc_byte_cnt[21]), .ZN(n16327) );
NAND2_X2 U12097 ( .A1(n17927), .A2(n16329), .ZN(n13418) );
XNOR2_X2 U12098 ( .A(n19174), .B(aes_text_out[24]), .ZN(n16329) );
NAND2_X2 U12099 ( .A1(n18037), .A2(b_in[8]), .ZN(n16314) );
NAND2_X2 U12100 ( .A1(n16330), .A2(n16331), .ZN(N3094) );
NAND2_X2 U12101 ( .A1(n16332), .A2(n18069), .ZN(n16331) );
XNOR2_X2 U12102 ( .A(n18918), .B(n16333), .ZN(n16332) );
NAND2_X2 U12106 ( .A1(n17927), .A2(n16337), .ZN(n13412) );
XNOR2_X2 U12107 ( .A(n19175), .B(aes_text_out[23]), .ZN(n16337) );
NAND2_X2 U12108 ( .A1(n16338), .A2(n16339), .ZN(n16334) );
NAND2_X2 U12109 ( .A1(n13414), .A2(n16325), .ZN(n16339) );
XOR2_X2 U12110 ( .A(n16340), .B(aes_text_out[23]), .Z(n13414) );
NAND2_X2 U12111 ( .A1(n17909), .A2(n16340), .ZN(n16338) );
NAND2_X2 U12112 ( .A1(n16341), .A2(n16342), .ZN(n16340) );
NAND2_X2 U12113 ( .A1(n17855), .A2(n17736), .ZN(n16342) );
NAND2_X2 U12114 ( .A1(n17851), .A2(n17728), .ZN(n16341) );
NAND2_X2 U12115 ( .A1(n18037), .A2(b_in[7]), .ZN(n16330) );
NAND2_X2 U12116 ( .A1(n16343), .A2(n16344), .ZN(N3093) );
NAND2_X2 U12117 ( .A1(n16345), .A2(n18069), .ZN(n16344) );
XNOR2_X2 U12118 ( .A(n18917), .B(n16346), .ZN(n16345) );
NAND2_X2 U12122 ( .A1(n17927), .A2(n16350), .ZN(n13406) );
XNOR2_X2 U12123 ( .A(n19176), .B(aes_text_out[22]), .ZN(n16350) );
NAND2_X2 U12124 ( .A1(n16351), .A2(n16352), .ZN(n16347) );
NAND2_X2 U12125 ( .A1(n13408), .A2(n16325), .ZN(n16352) );
XOR2_X2 U12126 ( .A(n16353), .B(aes_text_out[22]), .Z(n13408) );
NAND2_X2 U12127 ( .A1(n17909), .A2(n16353), .ZN(n16351) );
NAND2_X2 U12128 ( .A1(n16354), .A2(n16355), .ZN(n16353) );
NAND2_X2 U12129 ( .A1(n17855), .A2(n17737), .ZN(n16355) );
NAND2_X2 U12130 ( .A1(n17851), .A2(n17729), .ZN(n16354) );
NAND2_X2 U12131 ( .A1(n18037), .A2(b_in[6]), .ZN(n16343) );
NAND2_X2 U12132 ( .A1(n16356), .A2(n16357), .ZN(N3092) );
NAND2_X2 U12133 ( .A1(n16358), .A2(n18069), .ZN(n16357) );
XNOR2_X2 U12134 ( .A(n18916), .B(n16359), .ZN(n16358) );
NAND2_X2 U12138 ( .A1(n17927), .A2(n16363), .ZN(n13400) );
XNOR2_X2 U12139 ( .A(n19177), .B(aes_text_out[21]), .ZN(n16363) );
NAND2_X2 U12140 ( .A1(n16364), .A2(n16365), .ZN(n16360) );
NAND2_X2 U12141 ( .A1(n13402), .A2(n16325), .ZN(n16365) );
XOR2_X2 U12142 ( .A(n16366), .B(aes_text_out[21]), .Z(n13402) );
NAND2_X2 U12143 ( .A1(n17909), .A2(n16366), .ZN(n16364) );
NAND2_X2 U12144 ( .A1(n16367), .A2(n16368), .ZN(n16366) );
NAND2_X2 U12145 ( .A1(n17855), .A2(n17738), .ZN(n16368) );
NAND2_X2 U12146 ( .A1(n17851), .A2(n17730), .ZN(n16367) );
NAND2_X2 U12147 ( .A1(n18037), .A2(b_in[5]), .ZN(n16356) );
NAND2_X2 U12148 ( .A1(n16369), .A2(n16370), .ZN(N3091) );
NAND2_X2 U12149 ( .A1(n16371), .A2(n18069), .ZN(n16370) );
XNOR2_X2 U12150 ( .A(n18915), .B(n16372), .ZN(n16371) );
NAND2_X2 U12154 ( .A1(n17928), .A2(n16376), .ZN(n13394) );
XNOR2_X2 U12155 ( .A(n19178), .B(aes_text_out[20]), .ZN(n16376) );
NAND2_X2 U12156 ( .A1(n16377), .A2(n16378), .ZN(n16373) );
NAND2_X2 U12157 ( .A1(n13396), .A2(n16325), .ZN(n16378) );
XOR2_X2 U12158 ( .A(n16379), .B(aes_text_out[20]), .Z(n13396) );
NAND2_X2 U12159 ( .A1(n17909), .A2(n16379), .ZN(n16377) );
NAND2_X2 U12160 ( .A1(n16380), .A2(n16381), .ZN(n16379) );
NAND2_X2 U12161 ( .A1(n17855), .A2(n17739), .ZN(n16381) );
NAND2_X2 U12162 ( .A1(n17851), .A2(n17731), .ZN(n16380) );
NAND2_X2 U12163 ( .A1(n18037), .A2(b_in[4]), .ZN(n16369) );
NAND2_X2 U12164 ( .A1(n16382), .A2(n16383), .ZN(N3090) );
NAND2_X2 U12165 ( .A1(n16384), .A2(n18069), .ZN(n16383) );
XNOR2_X2 U12166 ( .A(n18914), .B(n16385), .ZN(n16384) );
NAND2_X2 U12170 ( .A1(n17927), .A2(n16389), .ZN(n13388) );
XNOR2_X2 U12171 ( .A(n19179), .B(aes_text_out[19]), .ZN(n16389) );
NAND2_X2 U12172 ( .A1(n16390), .A2(n16391), .ZN(n16386) );
NAND2_X2 U12173 ( .A1(n13390), .A2(n16325), .ZN(n16391) );
XOR2_X2 U12174 ( .A(n16392), .B(aes_text_out[19]), .Z(n13390) );
NAND2_X2 U12175 ( .A1(n17909), .A2(n16392), .ZN(n16390) );
NAND2_X2 U12176 ( .A1(n16393), .A2(n16394), .ZN(n16392) );
NAND2_X2 U12177 ( .A1(n17856), .A2(n17740), .ZN(n16394) );
NAND2_X2 U12178 ( .A1(n17851), .A2(n17732), .ZN(n16393) );
NAND2_X2 U12179 ( .A1(n18037), .A2(b_in[3]), .ZN(n16382) );
NAND2_X2 U12180 ( .A1(n16395), .A2(n16396), .ZN(N3089) );
NAND2_X2 U12181 ( .A1(n16397), .A2(n18069), .ZN(n16396) );
XNOR2_X2 U12182 ( .A(n18913), .B(n16398), .ZN(n16397) );
NAND2_X2 U12186 ( .A1(n17928), .A2(n16402), .ZN(n13382) );
XNOR2_X2 U12187 ( .A(n19180), .B(aes_text_out[18]), .ZN(n16402) );
NAND2_X2 U12188 ( .A1(n16403), .A2(n16404), .ZN(n16399) );
NAND2_X2 U12189 ( .A1(n13384), .A2(n16325), .ZN(n16404) );
XOR2_X2 U12190 ( .A(n16405), .B(aes_text_out[18]), .Z(n13384) );
NAND2_X2 U12191 ( .A1(n17909), .A2(n16405), .ZN(n16403) );
NAND2_X2 U12192 ( .A1(n16406), .A2(n16407), .ZN(n16405) );
NAND2_X2 U12193 ( .A1(n17856), .A2(n17741), .ZN(n16407) );
NAND2_X2 U12194 ( .A1(n17851), .A2(n17733), .ZN(n16406) );
NAND2_X2 U12195 ( .A1(n18037), .A2(b_in[2]), .ZN(n16395) );
NAND2_X2 U12196 ( .A1(n16408), .A2(n16409), .ZN(N3088) );
NAND2_X2 U12197 ( .A1(n16410), .A2(n18069), .ZN(n16409) );
XNOR2_X2 U12198 ( .A(n18912), .B(n16411), .ZN(n16410) );
NAND2_X2 U12202 ( .A1(n17927), .A2(n16415), .ZN(n13376) );
XNOR2_X2 U12203 ( .A(n19181), .B(aes_text_out[17]), .ZN(n16415) );
NAND2_X2 U12204 ( .A1(n16416), .A2(n16417), .ZN(n16412) );
NAND2_X2 U12205 ( .A1(n13378), .A2(n16325), .ZN(n16417) );
XOR2_X2 U12206 ( .A(n16418), .B(aes_text_out[17]), .Z(n13378) );
NAND2_X2 U12207 ( .A1(n17909), .A2(n16418), .ZN(n16416) );
NAND2_X2 U12208 ( .A1(n16419), .A2(n16420), .ZN(n16418) );
NAND2_X2 U12209 ( .A1(n17856), .A2(n17742), .ZN(n16420) );
NAND2_X2 U12210 ( .A1(n17851), .A2(n17734), .ZN(n16419) );
NAND2_X2 U12211 ( .A1(n18037), .A2(b_in[1]), .ZN(n16408) );
NAND2_X2 U12212 ( .A1(n16421), .A2(n16422), .ZN(N3087) );
NAND2_X2 U12213 ( .A1(n16423), .A2(n18064), .ZN(n16422) );
XNOR2_X2 U12214 ( .A(n18911), .B(n16424), .ZN(n16423) );
NAND2_X2 U12218 ( .A1(n17928), .A2(n16428), .ZN(n13370) );
XNOR2_X2 U12219 ( .A(n19182), .B(aes_text_out[16]), .ZN(n16428) );
NAND2_X2 U12220 ( .A1(n16429), .A2(n16430), .ZN(n16425) );
NAND2_X2 U12221 ( .A1(n13372), .A2(n16325), .ZN(n16430) );
NAND2_X2 U12223 ( .A1(n17856), .A2(n17945), .ZN(n16432) );
XOR2_X2 U12224 ( .A(n16433), .B(aes_text_out[16]), .Z(n13372) );
NAND2_X2 U12225 ( .A1(n17909), .A2(n16433), .ZN(n16429) );
NAND2_X2 U12226 ( .A1(n16434), .A2(n16435), .ZN(n16433) );
NAND2_X2 U12227 ( .A1(n17856), .A2(n17743), .ZN(n16435) );
NAND2_X2 U12229 ( .A1(n17851), .A2(n17735), .ZN(n16434) );
NAND2_X2 U12230 ( .A1(n18037), .A2(b_in[0]), .ZN(n16421) );
XNOR2_X2 U12232 ( .A(n16437), .B(n18910), .ZN(n16436) );
NAND2_X2 U12236 ( .A1(n16443), .A2(n16444), .ZN(n13365) );
NAND2_X2 U12237 ( .A1(n17933), .A2(n19191), .ZN(n16444) );
NAND2_X2 U12238 ( .A1(n16445), .A2(n16446), .ZN(n13364) );
NAND2_X2 U12240 ( .A1(n18634), .A2(n17736), .ZN(n16448) );
NAND2_X2 U12241 ( .A1(n17928), .A2(n17728), .ZN(n16447) );
NAND2_X2 U12242 ( .A1(aes_text_out[15]), .A2(n16449), .ZN(n16445) );
NAND2_X2 U12243 ( .A1(n17928), .A2(n19183), .ZN(n16449) );
NAND2_X2 U12245 ( .A1(n17907), .A2(n17728), .ZN(n16439) );
NAND2_X2 U12246 ( .A1(n17999), .A2(enc_byte_cnt[12]), .ZN(n16438) );
XNOR2_X2 U12248 ( .A(n16452), .B(n18909), .ZN(n16451) );
NAND2_X2 U12252 ( .A1(n16443), .A2(n16458), .ZN(n13359) );
NAND2_X2 U12253 ( .A1(n17933), .A2(n19192), .ZN(n16458) );
NAND2_X2 U12254 ( .A1(n16459), .A2(n16460), .ZN(n13358) );
NAND2_X2 U12256 ( .A1(n18634), .A2(n17737), .ZN(n16462) );
NAND2_X2 U12257 ( .A1(n17928), .A2(n17729), .ZN(n16461) );
NAND2_X2 U12258 ( .A1(aes_text_out[14]), .A2(n16463), .ZN(n16459) );
NAND2_X2 U12259 ( .A1(n17928), .A2(n19184), .ZN(n16463) );
NAND2_X2 U12261 ( .A1(n17908), .A2(n17729), .ZN(n16454) );
NAND2_X2 U12262 ( .A1(n17999), .A2(enc_byte_cnt[11]), .ZN(n16453) );
XNOR2_X2 U12264 ( .A(n16465), .B(n18908), .ZN(n16464) );
NAND2_X2 U12268 ( .A1(n16443), .A2(n16471), .ZN(n13353) );
NAND2_X2 U12269 ( .A1(n17933), .A2(n19193), .ZN(n16471) );
NAND2_X2 U12270 ( .A1(n16472), .A2(n16473), .ZN(n13352) );
NAND2_X2 U12272 ( .A1(n18634), .A2(n17738), .ZN(n16475) );
NAND2_X2 U12273 ( .A1(n17928), .A2(n17730), .ZN(n16474) );
NAND2_X2 U12274 ( .A1(aes_text_out[13]), .A2(n16476), .ZN(n16472) );
NAND2_X2 U12275 ( .A1(n17928), .A2(n19185), .ZN(n16476) );
NAND2_X2 U12277 ( .A1(n17907), .A2(n17730), .ZN(n16467) );
NAND2_X2 U12278 ( .A1(n17999), .A2(enc_byte_cnt[10]), .ZN(n16466) );
XNOR2_X2 U12280 ( .A(n16478), .B(n18907), .ZN(n16477) );
NAND2_X2 U12284 ( .A1(n16443), .A2(n16484), .ZN(n13347) );
NAND2_X2 U12285 ( .A1(n17933), .A2(n19194), .ZN(n16484) );
NAND2_X2 U12286 ( .A1(n16485), .A2(n16486), .ZN(n13346) );
NAND2_X2 U12288 ( .A1(n18634), .A2(n17739), .ZN(n16488) );
NAND2_X2 U12289 ( .A1(n17928), .A2(n17731), .ZN(n16487) );
NAND2_X2 U12290 ( .A1(aes_text_out[12]), .A2(n16489), .ZN(n16485) );
NAND2_X2 U12291 ( .A1(n17929), .A2(n19186), .ZN(n16489) );
NAND2_X2 U12293 ( .A1(n17908), .A2(n17731), .ZN(n16480) );
NAND2_X2 U12294 ( .A1(n17999), .A2(enc_byte_cnt[9]), .ZN(n16479) );
XNOR2_X2 U12296 ( .A(n16491), .B(n18906), .ZN(n16490) );
NAND2_X2 U12300 ( .A1(n16443), .A2(n16497), .ZN(n13341) );
NAND2_X2 U12301 ( .A1(n17933), .A2(n19195), .ZN(n16497) );
NAND2_X2 U12302 ( .A1(n16498), .A2(n16499), .ZN(n13340) );
NAND2_X2 U12304 ( .A1(n18634), .A2(n17740), .ZN(n16501) );
NAND2_X2 U12305 ( .A1(n17929), .A2(n17732), .ZN(n16500) );
NAND2_X2 U12306 ( .A1(aes_text_out[11]), .A2(n16502), .ZN(n16498) );
NAND2_X2 U12307 ( .A1(n17929), .A2(n19187), .ZN(n16502) );
NAND2_X2 U12309 ( .A1(n17907), .A2(n17732), .ZN(n16493) );
NAND2_X2 U12310 ( .A1(n17999), .A2(enc_byte_cnt[8]), .ZN(n16492) );
XNOR2_X2 U12312 ( .A(n16504), .B(n18905), .ZN(n16503) );
NAND2_X2 U12316 ( .A1(n16443), .A2(n16510), .ZN(n13335) );
NAND2_X2 U12317 ( .A1(n17933), .A2(n19196), .ZN(n16510) );
NAND2_X2 U12318 ( .A1(n16511), .A2(n16512), .ZN(n13334) );
NAND2_X2 U12320 ( .A1(n18634), .A2(n17741), .ZN(n16514) );
NAND2_X2 U12321 ( .A1(n17928), .A2(n17733), .ZN(n16513) );
NAND2_X2 U12322 ( .A1(aes_text_out[10]), .A2(n16515), .ZN(n16511) );
NAND2_X2 U12323 ( .A1(n17929), .A2(n19188), .ZN(n16515) );
NAND2_X2 U12325 ( .A1(n17908), .A2(n17733), .ZN(n16506) );
NAND2_X2 U12326 ( .A1(n17999), .A2(enc_byte_cnt[7]), .ZN(n16505) );
XNOR2_X2 U12328 ( .A(n16517), .B(n18904), .ZN(n16516) );
NAND2_X2 U12332 ( .A1(n16443), .A2(n16523), .ZN(n13329) );
NAND2_X2 U12333 ( .A1(n17933), .A2(n19197), .ZN(n16523) );
NAND2_X2 U12334 ( .A1(n16524), .A2(n16525), .ZN(n13328) );
NAND2_X2 U12336 ( .A1(n18634), .A2(n17742), .ZN(n16527) );
NAND2_X2 U12337 ( .A1(n17929), .A2(n17734), .ZN(n16526) );
NAND2_X2 U12338 ( .A1(aes_text_out[9]), .A2(n16528), .ZN(n16524) );
NAND2_X2 U12339 ( .A1(n17929), .A2(n19189), .ZN(n16528) );
NAND2_X2 U12341 ( .A1(n17907), .A2(n17734), .ZN(n16519) );
NAND2_X2 U12342 ( .A1(n17999), .A2(enc_byte_cnt[6]), .ZN(n16518) );
XNOR2_X2 U12344 ( .A(n16530), .B(n18903), .ZN(n16529) );
NAND2_X2 U12348 ( .A1(n16443), .A2(n16536), .ZN(n13323) );
NAND2_X2 U12349 ( .A1(n17933), .A2(n19198), .ZN(n16536) );
NAND2_X2 U12350 ( .A1(n17933), .A2(n16537), .ZN(n16443) );
NAND2_X2 U12351 ( .A1(n16538), .A2(n16539), .ZN(n13322) );
NAND2_X2 U12353 ( .A1(n18634), .A2(n17743), .ZN(n16541) );
NAND2_X2 U12354 ( .A1(n17851), .A2(n17936), .ZN(n16431) );
NAND2_X2 U12356 ( .A1(n17929), .A2(n17735), .ZN(n16540) );
NAND2_X2 U12357 ( .A1(aes_text_out[8]), .A2(n16543), .ZN(n16538) );
NAND2_X2 U12358 ( .A1(n17929), .A2(n19190), .ZN(n16543) );
NAND2_X2 U12360 ( .A1(n17909), .A2(n17851), .ZN(n16450) );
NAND2_X2 U12361 ( .A1(n17892), .A2(n17882), .ZN(n16537) );
NAND2_X2 U12365 ( .A1(n17906), .A2(n17735), .ZN(n16532) );
NAND2_X2 U12366 ( .A1(n17999), .A2(enc_byte_cnt[5]), .ZN(n16531) );
XNOR2_X2 U12368 ( .A(n17264), .B(n16545), .ZN(n16544) );
NAND2_X2 U12370 ( .A1(n17929), .A2(n16548), .ZN(n13317) );
XNOR2_X2 U12371 ( .A(n19191), .B(aes_text_out[7]), .ZN(n16548) );
XNOR2_X2 U12375 ( .A(n17266), .B(n16550), .ZN(n16549) );
NAND2_X2 U12377 ( .A1(n17930), .A2(n16553), .ZN(n13312) );
XNOR2_X2 U12378 ( .A(n19192), .B(aes_text_out[6]), .ZN(n16553) );
XNOR2_X2 U12382 ( .A(n17268), .B(n16555), .ZN(n16554) );
NAND2_X2 U12384 ( .A1(n17929), .A2(n16558), .ZN(n13307) );
XNOR2_X2 U12385 ( .A(n19193), .B(aes_text_out[5]), .ZN(n16558) );
XNOR2_X2 U12389 ( .A(n17270), .B(n16560), .ZN(n16559) );
NAND2_X2 U12391 ( .A1(n17930), .A2(n16563), .ZN(n13302) );
XNOR2_X2 U12392 ( .A(n19194), .B(aes_text_out[4]), .ZN(n16563) );
XNOR2_X2 U12396 ( .A(n17272), .B(n16565), .ZN(n16564) );
NAND2_X2 U12398 ( .A1(n17930), .A2(n16568), .ZN(n13297) );
XNOR2_X2 U12399 ( .A(n19195), .B(aes_text_out[3]), .ZN(n16568) );
XNOR2_X2 U12403 ( .A(n17274), .B(n16570), .ZN(n16569) );
NAND2_X2 U12406 ( .A1(n17930), .A2(n16572), .ZN(n13292) );
XNOR2_X2 U12407 ( .A(n19196), .B(aes_text_out[2]), .ZN(n16572) );
XNOR2_X2 U12409 ( .A(n17276), .B(n16574), .ZN(n16573) );
NAND2_X2 U12412 ( .A1(n17929), .A2(n16576), .ZN(n13287) );
XNOR2_X2 U12413 ( .A(n19197), .B(aes_text_out[1]), .ZN(n16576) );
XNOR2_X2 U12415 ( .A(n17278), .B(n16578), .ZN(n16577) );
NAND2_X2 U12419 ( .A1(n17930), .A2(n16580), .ZN(n13280) );
XNOR2_X2 U12420 ( .A(n19198), .B(aes_text_out[0]), .ZN(n16580) );
AND2_X2 U12424 ( .A1(n18056), .A2(z_out[127]), .ZN(N3070) );
AND2_X2 U12425 ( .A1(n18056), .A2(z_out[126]), .ZN(N3069) );
AND2_X2 U12426 ( .A1(n18056), .A2(z_out[125]), .ZN(N3068) );
AND2_X2 U12427 ( .A1(n18056), .A2(z_out[124]), .ZN(N3067) );
AND2_X2 U12428 ( .A1(n18056), .A2(z_out[123]), .ZN(N3066) );
AND2_X2 U12429 ( .A1(n18056), .A2(z_out[122]), .ZN(N3065) );
AND2_X2 U12430 ( .A1(n18056), .A2(z_out[121]), .ZN(N3064) );
AND2_X2 U12431 ( .A1(n18056), .A2(z_out[120]), .ZN(N3063) );
AND2_X2 U12432 ( .A1(n18056), .A2(z_out[119]), .ZN(N3062) );
AND2_X2 U12433 ( .A1(n18056), .A2(z_out[118]), .ZN(N3061) );
AND2_X2 U12434 ( .A1(n18056), .A2(z_out[117]), .ZN(N3060) );
AND2_X2 U12435 ( .A1(n18056), .A2(z_out[116]), .ZN(N3059) );
AND2_X2 U12436 ( .A1(n18056), .A2(z_out[115]), .ZN(N3058) );
AND2_X2 U12437 ( .A1(n18056), .A2(z_out[114]), .ZN(N3057) );
AND2_X2 U12438 ( .A1(n18056), .A2(z_out[113]), .ZN(N3056) );
AND2_X2 U12439 ( .A1(n18055), .A2(z_out[112]), .ZN(N3055) );
AND2_X2 U12440 ( .A1(n18055), .A2(z_out[111]), .ZN(N3054) );
AND2_X2 U12441 ( .A1(n18055), .A2(z_out[110]), .ZN(N3053) );
AND2_X2 U12442 ( .A1(n18055), .A2(z_out[109]), .ZN(N3052) );
AND2_X2 U12443 ( .A1(n18055), .A2(z_out[108]), .ZN(N3051) );
AND2_X2 U12444 ( .A1(n18055), .A2(z_out[107]), .ZN(N3050) );
AND2_X2 U12445 ( .A1(n18055), .A2(z_out[106]), .ZN(N3049) );
AND2_X2 U12446 ( .A1(n18055), .A2(z_out[105]), .ZN(N3048) );
AND2_X2 U12447 ( .A1(n18055), .A2(z_out[104]), .ZN(N3047) );
AND2_X2 U12448 ( .A1(n18055), .A2(z_out[103]), .ZN(N3046) );
AND2_X2 U12449 ( .A1(n18055), .A2(z_out[102]), .ZN(N3045) );
AND2_X2 U12450 ( .A1(n18055), .A2(z_out[101]), .ZN(N3044) );
AND2_X2 U12451 ( .A1(n18055), .A2(z_out[100]), .ZN(N3043) );
AND2_X2 U12452 ( .A1(n18055), .A2(z_out[99]), .ZN(N3042) );
AND2_X2 U12453 ( .A1(n18055), .A2(z_out[98]), .ZN(N3041) );
AND2_X2 U12454 ( .A1(n18055), .A2(z_out[97]), .ZN(N3040) );
AND2_X2 U12455 ( .A1(n18055), .A2(z_out[96]), .ZN(N3039) );
AND2_X2 U12456 ( .A1(n18055), .A2(z_out[95]), .ZN(N3038) );
AND2_X2 U12457 ( .A1(n18055), .A2(z_out[94]), .ZN(N3037) );
AND2_X2 U12458 ( .A1(n18055), .A2(z_out[93]), .ZN(N3036) );
AND2_X2 U12459 ( .A1(n18055), .A2(z_out[92]), .ZN(N3035) );
AND2_X2 U12460 ( .A1(n18055), .A2(z_out[91]), .ZN(N3034) );
AND2_X2 U12461 ( .A1(n18055), .A2(z_out[90]), .ZN(N3033) );
AND2_X2 U12462 ( .A1(n18054), .A2(z_out[89]), .ZN(N3032) );
AND2_X2 U12463 ( .A1(n18054), .A2(z_out[88]), .ZN(N3031) );
AND2_X2 U12464 ( .A1(n18054), .A2(z_out[87]), .ZN(N3030) );
AND2_X2 U12465 ( .A1(n18054), .A2(z_out[86]), .ZN(N3029) );
AND2_X2 U12466 ( .A1(n18054), .A2(z_out[85]), .ZN(N3028) );
AND2_X2 U12467 ( .A1(n18054), .A2(z_out[84]), .ZN(N3027) );
AND2_X2 U12468 ( .A1(n18054), .A2(z_out[83]), .ZN(N3026) );
AND2_X2 U12469 ( .A1(n18054), .A2(z_out[82]), .ZN(N3025) );
AND2_X2 U12470 ( .A1(n18054), .A2(z_out[81]), .ZN(N3024) );
AND2_X2 U12471 ( .A1(n18054), .A2(z_out[80]), .ZN(N3023) );
AND2_X2 U12472 ( .A1(n18054), .A2(z_out[79]), .ZN(N3022) );
AND2_X2 U12473 ( .A1(n18054), .A2(z_out[78]), .ZN(N3021) );
AND2_X2 U12474 ( .A1(n18054), .A2(z_out[77]), .ZN(N3020) );
AND2_X2 U12475 ( .A1(n18054), .A2(z_out[76]), .ZN(N3019) );
AND2_X2 U12476 ( .A1(n18054), .A2(z_out[75]), .ZN(N3018) );
AND2_X2 U12477 ( .A1(n18054), .A2(z_out[74]), .ZN(N3017) );
AND2_X2 U12478 ( .A1(n18054), .A2(z_out[73]), .ZN(N3016) );
AND2_X2 U12479 ( .A1(n18054), .A2(z_out[72]), .ZN(N3015) );
AND2_X2 U12480 ( .A1(n18054), .A2(z_out[71]), .ZN(N3014) );
AND2_X2 U12481 ( .A1(n18054), .A2(z_out[70]), .ZN(N3013) );
AND2_X2 U12482 ( .A1(n18054), .A2(z_out[69]), .ZN(N3012) );
AND2_X2 U12483 ( .A1(n18054), .A2(z_out[68]), .ZN(N3011) );
AND2_X2 U12484 ( .A1(n18054), .A2(z_out[67]), .ZN(N3010) );
AND2_X2 U12485 ( .A1(n18053), .A2(z_out[66]), .ZN(N3009) );
AND2_X2 U12486 ( .A1(n18053), .A2(z_out[65]), .ZN(N3008) );
AND2_X2 U12487 ( .A1(n18051), .A2(z_out[64]), .ZN(N3007) );
AND2_X2 U12488 ( .A1(n18053), .A2(z_out[63]), .ZN(N3006) );
AND2_X2 U12489 ( .A1(n18053), .A2(z_out[62]), .ZN(N3005) );
AND2_X2 U12490 ( .A1(n18053), .A2(z_out[61]), .ZN(N3004) );
AND2_X2 U12491 ( .A1(n18053), .A2(z_out[60]), .ZN(N3003) );
AND2_X2 U12492 ( .A1(n18053), .A2(z_out[59]), .ZN(N3002) );
AND2_X2 U12493 ( .A1(n18053), .A2(z_out[58]), .ZN(N3001) );
AND2_X2 U12494 ( .A1(n18053), .A2(z_out[57]), .ZN(N3000) );
AND2_X2 U12495 ( .A1(n18053), .A2(z_out[56]), .ZN(N2999) );
AND2_X2 U12496 ( .A1(n18053), .A2(z_out[55]), .ZN(N2998) );
AND2_X2 U12497 ( .A1(n18053), .A2(z_out[54]), .ZN(N2997) );
AND2_X2 U12498 ( .A1(n18053), .A2(z_out[53]), .ZN(N2996) );
AND2_X2 U12499 ( .A1(n18053), .A2(z_out[52]), .ZN(N2995) );
AND2_X2 U12500 ( .A1(n18053), .A2(z_out[51]), .ZN(N2994) );
AND2_X2 U12501 ( .A1(n18053), .A2(z_out[50]), .ZN(N2993) );
AND2_X2 U12502 ( .A1(n18053), .A2(z_out[49]), .ZN(N2992) );
AND2_X2 U12503 ( .A1(n18053), .A2(z_out[48]), .ZN(N2991) );
AND2_X2 U12504 ( .A1(n18053), .A2(z_out[47]), .ZN(N2990) );
AND2_X2 U12505 ( .A1(n18053), .A2(z_out[46]), .ZN(N2989) );
AND2_X2 U12506 ( .A1(n18053), .A2(z_out[45]), .ZN(N2988) );
AND2_X2 U12507 ( .A1(n18053), .A2(z_out[44]), .ZN(N2987) );
AND2_X2 U12508 ( .A1(n18052), .A2(z_out[43]), .ZN(N2986) );
AND2_X2 U12509 ( .A1(n18052), .A2(z_out[42]), .ZN(N2985) );
AND2_X2 U12510 ( .A1(n18052), .A2(z_out[41]), .ZN(N2984) );
AND2_X2 U12511 ( .A1(n18052), .A2(z_out[40]), .ZN(N2983) );
AND2_X2 U12512 ( .A1(n18052), .A2(z_out[39]), .ZN(N2982) );
AND2_X2 U12513 ( .A1(n18052), .A2(z_out[38]), .ZN(N2981) );
AND2_X2 U12514 ( .A1(n18052), .A2(z_out[37]), .ZN(N2980) );
AND2_X2 U12515 ( .A1(n18052), .A2(z_out[36]), .ZN(N2979) );
AND2_X2 U12516 ( .A1(n18052), .A2(z_out[35]), .ZN(N2978) );
AND2_X2 U12517 ( .A1(n18052), .A2(z_out[34]), .ZN(N2977) );
AND2_X2 U12518 ( .A1(n18052), .A2(z_out[33]), .ZN(N2976) );
AND2_X2 U12519 ( .A1(n18052), .A2(z_out[32]), .ZN(N2975) );
AND2_X2 U12520 ( .A1(n18052), .A2(z_out[31]), .ZN(N2974) );
AND2_X2 U12521 ( .A1(n18052), .A2(z_out[30]), .ZN(N2973) );
AND2_X2 U12522 ( .A1(n18052), .A2(z_out[29]), .ZN(N2972) );
AND2_X2 U12523 ( .A1(n18052), .A2(z_out[28]), .ZN(N2971) );
AND2_X2 U12524 ( .A1(n18052), .A2(z_out[27]), .ZN(N2970) );
AND2_X2 U12525 ( .A1(n18052), .A2(z_out[26]), .ZN(N2969) );
AND2_X2 U12526 ( .A1(n18052), .A2(z_out[25]), .ZN(N2968) );
AND2_X2 U12527 ( .A1(n18052), .A2(z_out[24]), .ZN(N2967) );
AND2_X2 U12528 ( .A1(n18052), .A2(z_out[23]), .ZN(N2966) );
AND2_X2 U12529 ( .A1(n18052), .A2(z_out[22]), .ZN(N2965) );
AND2_X2 U12530 ( .A1(n18052), .A2(z_out[21]), .ZN(N2964) );
AND2_X2 U12531 ( .A1(n18051), .A2(z_out[20]), .ZN(N2963) );
AND2_X2 U12532 ( .A1(n18051), .A2(z_out[19]), .ZN(N2962) );
AND2_X2 U12533 ( .A1(n18051), .A2(z_out[18]), .ZN(N2961) );
AND2_X2 U12534 ( .A1(n18051), .A2(z_out[17]), .ZN(N2960) );
AND2_X2 U12535 ( .A1(n18051), .A2(z_out[16]), .ZN(N2959) );
AND2_X2 U12536 ( .A1(n18051), .A2(z_out[15]), .ZN(N2958) );
AND2_X2 U12537 ( .A1(n18051), .A2(z_out[14]), .ZN(N2957) );
AND2_X2 U12538 ( .A1(n18051), .A2(z_out[13]), .ZN(N2956) );
AND2_X2 U12539 ( .A1(n18051), .A2(z_out[12]), .ZN(N2955) );
AND2_X2 U12540 ( .A1(n18051), .A2(z_out[11]), .ZN(N2954) );
AND2_X2 U12541 ( .A1(n18051), .A2(z_out[10]), .ZN(N2953) );
AND2_X2 U12542 ( .A1(n18051), .A2(z_out[9]), .ZN(N2952) );
AND2_X2 U12543 ( .A1(n18051), .A2(z_out[8]), .ZN(N2951) );
AND2_X2 U12544 ( .A1(n18051), .A2(z_out[7]), .ZN(N2950) );
AND2_X2 U12545 ( .A1(n18051), .A2(z_out[6]), .ZN(N2949) );
AND2_X2 U12546 ( .A1(n18051), .A2(z_out[5]), .ZN(N2948) );
AND2_X2 U12547 ( .A1(n18051), .A2(z_out[4]), .ZN(N2947) );
AND2_X2 U12548 ( .A1(n18051), .A2(z_out[3]), .ZN(N2946) );
AND2_X2 U12549 ( .A1(n18053), .A2(z_out[2]), .ZN(N2945) );
AND2_X2 U12550 ( .A1(n18051), .A2(z_out[1]), .ZN(N2944) );
AND2_X2 U12551 ( .A1(n18056), .A2(z_out[0]), .ZN(N2943) );
NAND2_X2 U12552 ( .A1(n16581), .A2(n16582), .ZN(N2942) );
NAND2_X2 U12553 ( .A1(v_out[127]), .A2(n18047), .ZN(n16582) );
NAND2_X2 U12554 ( .A1(n18059), .A2(n17292), .ZN(n16581) );
NAND2_X2 U12555 ( .A1(n16583), .A2(n16584), .ZN(N2941) );
NAND2_X2 U12556 ( .A1(v_out[126]), .A2(n18044), .ZN(n16584) );
NAND2_X2 U12557 ( .A1(n18059), .A2(n17293), .ZN(n16583) );
NAND2_X2 U12558 ( .A1(n16585), .A2(n16586), .ZN(N2940) );
NAND2_X2 U12559 ( .A1(v_out[125]), .A2(n18044), .ZN(n16586) );
NAND2_X2 U12560 ( .A1(n18059), .A2(n17294), .ZN(n16585) );
NAND2_X2 U12561 ( .A1(n16587), .A2(n16588), .ZN(N2939) );
NAND2_X2 U12562 ( .A1(v_out[124]), .A2(n18044), .ZN(n16588) );
NAND2_X2 U12563 ( .A1(n18059), .A2(n17295), .ZN(n16587) );
NAND2_X2 U12564 ( .A1(n16589), .A2(n16590), .ZN(N2938) );
NAND2_X2 U12565 ( .A1(v_out[123]), .A2(n18044), .ZN(n16590) );
NAND2_X2 U12566 ( .A1(n18059), .A2(n17296), .ZN(n16589) );
NAND2_X2 U12567 ( .A1(n16591), .A2(n16592), .ZN(N2937) );
NAND2_X2 U12568 ( .A1(v_out[122]), .A2(n18044), .ZN(n16592) );
NAND2_X2 U12569 ( .A1(n18059), .A2(n17297), .ZN(n16591) );
NAND2_X2 U12570 ( .A1(n16593), .A2(n16594), .ZN(N2936) );
NAND2_X2 U12571 ( .A1(v_out[121]), .A2(n18044), .ZN(n16594) );
NAND2_X2 U12572 ( .A1(n18059), .A2(n17298), .ZN(n16593) );
NAND2_X2 U12573 ( .A1(n16595), .A2(n16596), .ZN(N2935) );
NAND2_X2 U12574 ( .A1(v_out[120]), .A2(n18044), .ZN(n16596) );
NAND2_X2 U12575 ( .A1(n18059), .A2(n17299), .ZN(n16595) );
NAND2_X2 U12576 ( .A1(n16597), .A2(n16598), .ZN(N2934) );
NAND2_X2 U12577 ( .A1(v_out[119]), .A2(n18044), .ZN(n16598) );
NAND2_X2 U12578 ( .A1(n18059), .A2(n17300), .ZN(n16597) );
NAND2_X2 U12579 ( .A1(n16599), .A2(n16600), .ZN(N2933) );
NAND2_X2 U12580 ( .A1(v_out[118]), .A2(n18044), .ZN(n16600) );
NAND2_X2 U12581 ( .A1(n18059), .A2(n17301), .ZN(n16599) );
NAND2_X2 U12582 ( .A1(n16601), .A2(n16602), .ZN(N2932) );
NAND2_X2 U12583 ( .A1(v_out[117]), .A2(n18044), .ZN(n16602) );
NAND2_X2 U12584 ( .A1(n18059), .A2(n17302), .ZN(n16601) );
NAND2_X2 U12585 ( .A1(n16603), .A2(n16604), .ZN(N2931) );
NAND2_X2 U12586 ( .A1(v_out[116]), .A2(n18044), .ZN(n16604) );
NAND2_X2 U12587 ( .A1(n18059), .A2(n17303), .ZN(n16603) );
NAND2_X2 U12588 ( .A1(n16605), .A2(n16606), .ZN(N2930) );
NAND2_X2 U12589 ( .A1(v_out[115]), .A2(n18044), .ZN(n16606) );
NAND2_X2 U12590 ( .A1(n18059), .A2(n17304), .ZN(n16605) );
NAND2_X2 U12591 ( .A1(n16607), .A2(n16608), .ZN(N2929) );
NAND2_X2 U12592 ( .A1(v_out[114]), .A2(n18044), .ZN(n16608) );
NAND2_X2 U12593 ( .A1(n18059), .A2(n17305), .ZN(n16607) );
NAND2_X2 U12594 ( .A1(n16609), .A2(n16610), .ZN(N2928) );
NAND2_X2 U12595 ( .A1(v_out[113]), .A2(n18044), .ZN(n16610) );
NAND2_X2 U12596 ( .A1(n18060), .A2(n17306), .ZN(n16609) );
NAND2_X2 U12597 ( .A1(n16611), .A2(n16612), .ZN(N2927) );
NAND2_X2 U12598 ( .A1(v_out[112]), .A2(n18044), .ZN(n16612) );
NAND2_X2 U12599 ( .A1(n18059), .A2(n17307), .ZN(n16611) );
NAND2_X2 U12600 ( .A1(n16613), .A2(n16614), .ZN(N2926) );
NAND2_X2 U12601 ( .A1(v_out[111]), .A2(n18044), .ZN(n16614) );
NAND2_X2 U12602 ( .A1(n18059), .A2(n17308), .ZN(n16613) );
NAND2_X2 U12603 ( .A1(n16615), .A2(n16616), .ZN(N2925) );
NAND2_X2 U12604 ( .A1(v_out[110]), .A2(n18044), .ZN(n16616) );
NAND2_X2 U12605 ( .A1(n18059), .A2(n17309), .ZN(n16615) );
NAND2_X2 U12606 ( .A1(n16617), .A2(n16618), .ZN(N2924) );
NAND2_X2 U12607 ( .A1(v_out[109]), .A2(n18045), .ZN(n16618) );
NAND2_X2 U12608 ( .A1(n18059), .A2(n17310), .ZN(n16617) );
NAND2_X2 U12609 ( .A1(n16619), .A2(n16620), .ZN(N2923) );
NAND2_X2 U12610 ( .A1(v_out[108]), .A2(n18045), .ZN(n16620) );
NAND2_X2 U12611 ( .A1(n18060), .A2(n17311), .ZN(n16619) );
NAND2_X2 U12612 ( .A1(n16621), .A2(n16622), .ZN(N2922) );
NAND2_X2 U12613 ( .A1(v_out[107]), .A2(n18045), .ZN(n16622) );
NAND2_X2 U12614 ( .A1(n18060), .A2(n17312), .ZN(n16621) );
NAND2_X2 U12615 ( .A1(n16623), .A2(n16624), .ZN(N2921) );
NAND2_X2 U12616 ( .A1(v_out[106]), .A2(n18045), .ZN(n16624) );
NAND2_X2 U12617 ( .A1(n18060), .A2(n17313), .ZN(n16623) );
NAND2_X2 U12618 ( .A1(n16625), .A2(n16626), .ZN(N2920) );
NAND2_X2 U12619 ( .A1(v_out[105]), .A2(n18045), .ZN(n16626) );
NAND2_X2 U12620 ( .A1(n18060), .A2(n17314), .ZN(n16625) );
NAND2_X2 U12621 ( .A1(n16627), .A2(n16628), .ZN(N2919) );
NAND2_X2 U12622 ( .A1(v_out[104]), .A2(n18045), .ZN(n16628) );
NAND2_X2 U12623 ( .A1(n18060), .A2(n17315), .ZN(n16627) );
NAND2_X2 U12624 ( .A1(n16629), .A2(n16630), .ZN(N2918) );
NAND2_X2 U12625 ( .A1(v_out[103]), .A2(n18045), .ZN(n16630) );
NAND2_X2 U12626 ( .A1(n18060), .A2(n17316), .ZN(n16629) );
NAND2_X2 U12627 ( .A1(n16631), .A2(n16632), .ZN(N2917) );
NAND2_X2 U12628 ( .A1(v_out[102]), .A2(n18045), .ZN(n16632) );
NAND2_X2 U12629 ( .A1(n18060), .A2(n17317), .ZN(n16631) );
NAND2_X2 U12630 ( .A1(n16633), .A2(n16634), .ZN(N2916) );
NAND2_X2 U12631 ( .A1(v_out[101]), .A2(n18045), .ZN(n16634) );
NAND2_X2 U12632 ( .A1(n18060), .A2(n17318), .ZN(n16633) );
NAND2_X2 U12633 ( .A1(n16635), .A2(n16636), .ZN(N2915) );
NAND2_X2 U12634 ( .A1(v_out[100]), .A2(n18045), .ZN(n16636) );
NAND2_X2 U12635 ( .A1(n18060), .A2(n17319), .ZN(n16635) );
NAND2_X2 U12636 ( .A1(n16637), .A2(n16638), .ZN(N2914) );
NAND2_X2 U12637 ( .A1(v_out[99]), .A2(n18045), .ZN(n16638) );
NAND2_X2 U12638 ( .A1(n18060), .A2(n17320), .ZN(n16637) );
NAND2_X2 U12639 ( .A1(n16639), .A2(n16640), .ZN(N2913) );
NAND2_X2 U12640 ( .A1(v_out[98]), .A2(n18045), .ZN(n16640) );
NAND2_X2 U12641 ( .A1(n18060), .A2(n17321), .ZN(n16639) );
NAND2_X2 U12642 ( .A1(n16641), .A2(n16642), .ZN(N2912) );
NAND2_X2 U12643 ( .A1(v_out[97]), .A2(n18045), .ZN(n16642) );
NAND2_X2 U12644 ( .A1(n18060), .A2(n17322), .ZN(n16641) );
NAND2_X2 U12645 ( .A1(n16643), .A2(n16644), .ZN(N2911) );
NAND2_X2 U12646 ( .A1(v_out[96]), .A2(n18045), .ZN(n16644) );
NAND2_X2 U12647 ( .A1(n18060), .A2(n17323), .ZN(n16643) );
NAND2_X2 U12648 ( .A1(n16645), .A2(n16646), .ZN(N2910) );
NAND2_X2 U12649 ( .A1(v_out[95]), .A2(n18045), .ZN(n16646) );
NAND2_X2 U12650 ( .A1(n18060), .A2(n17324), .ZN(n16645) );
NAND2_X2 U12651 ( .A1(n16647), .A2(n16648), .ZN(N2909) );
NAND2_X2 U12652 ( .A1(v_out[94]), .A2(n18045), .ZN(n16648) );
NAND2_X2 U12653 ( .A1(n18060), .A2(n17325), .ZN(n16647) );
NAND2_X2 U12654 ( .A1(n16649), .A2(n16650), .ZN(N2908) );
NAND2_X2 U12655 ( .A1(v_out[93]), .A2(n18045), .ZN(n16650) );
NAND2_X2 U12656 ( .A1(n18060), .A2(n17326), .ZN(n16649) );
NAND2_X2 U12657 ( .A1(n16651), .A2(n16652), .ZN(N2907) );
NAND2_X2 U12658 ( .A1(v_out[92]), .A2(n18045), .ZN(n16652) );
NAND2_X2 U12659 ( .A1(n18058), .A2(n17327), .ZN(n16651) );
NAND2_X2 U12660 ( .A1(n16653), .A2(n16654), .ZN(N2906) );
NAND2_X2 U12661 ( .A1(v_out[91]), .A2(n18046), .ZN(n16654) );
NAND2_X2 U12662 ( .A1(n18060), .A2(n17328), .ZN(n16653) );
NAND2_X2 U12663 ( .A1(n16655), .A2(n16656), .ZN(N2905) );
NAND2_X2 U12664 ( .A1(v_out[90]), .A2(n18046), .ZN(n16656) );
NAND2_X2 U12665 ( .A1(n18060), .A2(n17329), .ZN(n16655) );
NAND2_X2 U12666 ( .A1(n16657), .A2(n16658), .ZN(N2904) );
NAND2_X2 U12667 ( .A1(v_out[89]), .A2(n18046), .ZN(n16658) );
NAND2_X2 U12668 ( .A1(n18060), .A2(n17330), .ZN(n16657) );
NAND2_X2 U12669 ( .A1(n16659), .A2(n16660), .ZN(N2903) );
NAND2_X2 U12670 ( .A1(v_out[88]), .A2(n18046), .ZN(n16660) );
NAND2_X2 U12671 ( .A1(n18060), .A2(n17331), .ZN(n16659) );
NAND2_X2 U12672 ( .A1(n16661), .A2(n16662), .ZN(N2902) );
NAND2_X2 U12673 ( .A1(v_out[87]), .A2(n18046), .ZN(n16662) );
NAND2_X2 U12674 ( .A1(n18058), .A2(n17332), .ZN(n16661) );
NAND2_X2 U12675 ( .A1(n16663), .A2(n16664), .ZN(N2901) );
NAND2_X2 U12676 ( .A1(v_out[86]), .A2(n18046), .ZN(n16664) );
NAND2_X2 U12677 ( .A1(n18057), .A2(n17333), .ZN(n16663) );
NAND2_X2 U12678 ( .A1(n16665), .A2(n16666), .ZN(N2900) );
NAND2_X2 U12679 ( .A1(v_out[85]), .A2(n18046), .ZN(n16666) );
NAND2_X2 U12680 ( .A1(n18064), .A2(n17334), .ZN(n16665) );
NAND2_X2 U12681 ( .A1(n16667), .A2(n16668), .ZN(N2899) );
NAND2_X2 U12682 ( .A1(v_out[84]), .A2(n18046), .ZN(n16668) );
NAND2_X2 U12683 ( .A1(n18066), .A2(n17335), .ZN(n16667) );
NAND2_X2 U12684 ( .A1(n16669), .A2(n16670), .ZN(N2898) );
NAND2_X2 U12685 ( .A1(v_out[83]), .A2(n18046), .ZN(n16670) );
NAND2_X2 U12686 ( .A1(n18068), .A2(n17336), .ZN(n16669) );
NAND2_X2 U12687 ( .A1(n16671), .A2(n16672), .ZN(N2897) );
NAND2_X2 U12688 ( .A1(v_out[82]), .A2(n18046), .ZN(n16672) );
NAND2_X2 U12689 ( .A1(n18067), .A2(n17337), .ZN(n16671) );
NAND2_X2 U12690 ( .A1(n16673), .A2(n16674), .ZN(N2896) );
NAND2_X2 U12691 ( .A1(v_out[81]), .A2(n18046), .ZN(n16674) );
NAND2_X2 U12692 ( .A1(n18065), .A2(n17338), .ZN(n16673) );
NAND2_X2 U12693 ( .A1(n16675), .A2(n16676), .ZN(N2895) );
NAND2_X2 U12694 ( .A1(v_out[80]), .A2(n18046), .ZN(n16676) );
NAND2_X2 U12695 ( .A1(n18069), .A2(n17339), .ZN(n16675) );
NAND2_X2 U12696 ( .A1(n16677), .A2(n16678), .ZN(N2894) );
NAND2_X2 U12697 ( .A1(v_out[79]), .A2(n18046), .ZN(n16678) );
NAND2_X2 U12698 ( .A1(n18057), .A2(n17340), .ZN(n16677) );
NAND2_X2 U12699 ( .A1(n16679), .A2(n16680), .ZN(N2893) );
NAND2_X2 U12700 ( .A1(v_out[78]), .A2(n18046), .ZN(n16680) );
NAND2_X2 U12701 ( .A1(n18064), .A2(n17341), .ZN(n16679) );
NAND2_X2 U12702 ( .A1(n16681), .A2(n16682), .ZN(N2892) );
NAND2_X2 U12703 ( .A1(v_out[77]), .A2(n18046), .ZN(n16682) );
NAND2_X2 U12704 ( .A1(n18066), .A2(n17342), .ZN(n16681) );
NAND2_X2 U12705 ( .A1(n16683), .A2(n16684), .ZN(N2891) );
NAND2_X2 U12706 ( .A1(v_out[76]), .A2(n18046), .ZN(n16684) );
NAND2_X2 U12707 ( .A1(n18068), .A2(n17343), .ZN(n16683) );
NAND2_X2 U12708 ( .A1(n16685), .A2(n16686), .ZN(N2890) );
NAND2_X2 U12709 ( .A1(v_out[75]), .A2(n18046), .ZN(n16686) );
NAND2_X2 U12710 ( .A1(n18067), .A2(n17344), .ZN(n16685) );
NAND2_X2 U12711 ( .A1(n16687), .A2(n16688), .ZN(N2889) );
NAND2_X2 U12712 ( .A1(v_out[74]), .A2(n18046), .ZN(n16688) );
NAND2_X2 U12713 ( .A1(n18065), .A2(n17345), .ZN(n16687) );
NAND2_X2 U12714 ( .A1(n16689), .A2(n16690), .ZN(N2888) );
NAND2_X2 U12715 ( .A1(v_out[73]), .A2(n18047), .ZN(n16690) );
NAND2_X2 U12716 ( .A1(n18069), .A2(n17346), .ZN(n16689) );
NAND2_X2 U12717 ( .A1(n16691), .A2(n16692), .ZN(N2887) );
NAND2_X2 U12718 ( .A1(v_out[72]), .A2(n18047), .ZN(n16692) );
NAND2_X2 U12719 ( .A1(n18069), .A2(n17347), .ZN(n16691) );
NAND2_X2 U12720 ( .A1(n16693), .A2(n16694), .ZN(N2886) );
NAND2_X2 U12721 ( .A1(v_out[71]), .A2(n18047), .ZN(n16694) );
NAND2_X2 U12722 ( .A1(n18069), .A2(n17348), .ZN(n16693) );
NAND2_X2 U12723 ( .A1(n16695), .A2(n16696), .ZN(N2885) );
NAND2_X2 U12724 ( .A1(v_out[70]), .A2(n18047), .ZN(n16696) );
NAND2_X2 U12725 ( .A1(n18069), .A2(n17349), .ZN(n16695) );
NAND2_X2 U12726 ( .A1(n16697), .A2(n16698), .ZN(N2884) );
NAND2_X2 U12727 ( .A1(v_out[69]), .A2(n18047), .ZN(n16698) );
NAND2_X2 U12728 ( .A1(n18069), .A2(n17350), .ZN(n16697) );
NAND2_X2 U12729 ( .A1(n16699), .A2(n16700), .ZN(N2883) );
NAND2_X2 U12730 ( .A1(v_out[68]), .A2(n18047), .ZN(n16700) );
NAND2_X2 U12731 ( .A1(n18069), .A2(n17351), .ZN(n16699) );
NAND2_X2 U12732 ( .A1(n16701), .A2(n16702), .ZN(N2882) );
NAND2_X2 U12733 ( .A1(v_out[67]), .A2(n18047), .ZN(n16702) );
NAND2_X2 U12734 ( .A1(n18061), .A2(n17352), .ZN(n16701) );
NAND2_X2 U12735 ( .A1(n16703), .A2(n16704), .ZN(N2881) );
NAND2_X2 U12736 ( .A1(v_out[66]), .A2(n18047), .ZN(n16704) );
NAND2_X2 U12737 ( .A1(n18061), .A2(n17353), .ZN(n16703) );
NAND2_X2 U12738 ( .A1(n16705), .A2(n16706), .ZN(N2880) );
NAND2_X2 U12739 ( .A1(v_out[65]), .A2(n18047), .ZN(n16706) );
NAND2_X2 U12740 ( .A1(n18061), .A2(n17354), .ZN(n16705) );
NAND2_X2 U12741 ( .A1(n16707), .A2(n16708), .ZN(N2879) );
NAND2_X2 U12742 ( .A1(v_out[64]), .A2(n18047), .ZN(n16708) );
NAND2_X2 U12743 ( .A1(n18064), .A2(n17355), .ZN(n16707) );
NAND2_X2 U12744 ( .A1(n16709), .A2(n16710), .ZN(N2878) );
NAND2_X2 U12745 ( .A1(v_out[63]), .A2(n18047), .ZN(n16710) );
NAND2_X2 U12746 ( .A1(n18064), .A2(n17356), .ZN(n16709) );
NAND2_X2 U12747 ( .A1(n16711), .A2(n16712), .ZN(N2877) );
NAND2_X2 U12748 ( .A1(v_out[62]), .A2(n18047), .ZN(n16712) );
NAND2_X2 U12749 ( .A1(n18064), .A2(n17357), .ZN(n16711) );
NAND2_X2 U12750 ( .A1(n16713), .A2(n16714), .ZN(N2876) );
NAND2_X2 U12751 ( .A1(v_out[61]), .A2(n18047), .ZN(n16714) );
NAND2_X2 U12752 ( .A1(n18064), .A2(n17358), .ZN(n16713) );
NAND2_X2 U12753 ( .A1(n16715), .A2(n16716), .ZN(N2875) );
NAND2_X2 U12754 ( .A1(v_out[60]), .A2(n18047), .ZN(n16716) );
NAND2_X2 U12755 ( .A1(n18063), .A2(n17359), .ZN(n16715) );
NAND2_X2 U12756 ( .A1(n16717), .A2(n16718), .ZN(N2874) );
NAND2_X2 U12757 ( .A1(v_out[59]), .A2(n18047), .ZN(n16718) );
NAND2_X2 U12758 ( .A1(n18063), .A2(n17360), .ZN(n16717) );
NAND2_X2 U12759 ( .A1(n16719), .A2(n16720), .ZN(N2873) );
NAND2_X2 U12760 ( .A1(v_out[58]), .A2(n18047), .ZN(n16720) );
NAND2_X2 U12761 ( .A1(n18063), .A2(n17361), .ZN(n16719) );
NAND2_X2 U12762 ( .A1(n16721), .A2(n16722), .ZN(N2872) );
NAND2_X2 U12763 ( .A1(v_out[57]), .A2(n18048), .ZN(n16722) );
NAND2_X2 U12764 ( .A1(n18063), .A2(n17362), .ZN(n16721) );
NAND2_X2 U12765 ( .A1(n16723), .A2(n16724), .ZN(N2871) );
NAND2_X2 U12766 ( .A1(v_out[56]), .A2(n18048), .ZN(n16724) );
NAND2_X2 U12767 ( .A1(n18063), .A2(n17363), .ZN(n16723) );
NAND2_X2 U12768 ( .A1(n16725), .A2(n16726), .ZN(N2870) );
NAND2_X2 U12769 ( .A1(v_out[55]), .A2(n18048), .ZN(n16726) );
NAND2_X2 U12770 ( .A1(n18063), .A2(n17364), .ZN(n16725) );
NAND2_X2 U12771 ( .A1(n16727), .A2(n16728), .ZN(N2869) );
NAND2_X2 U12772 ( .A1(v_out[54]), .A2(n18048), .ZN(n16728) );
NAND2_X2 U12773 ( .A1(n18063), .A2(n17365), .ZN(n16727) );
NAND2_X2 U12774 ( .A1(n16729), .A2(n16730), .ZN(N2868) );
NAND2_X2 U12775 ( .A1(v_out[53]), .A2(n18048), .ZN(n16730) );
NAND2_X2 U12776 ( .A1(n18063), .A2(n17366), .ZN(n16729) );
NAND2_X2 U12777 ( .A1(n16731), .A2(n16732), .ZN(N2867) );
NAND2_X2 U12778 ( .A1(v_out[52]), .A2(n18048), .ZN(n16732) );
NAND2_X2 U12779 ( .A1(n18063), .A2(n17367), .ZN(n16731) );
NAND2_X2 U12780 ( .A1(n16733), .A2(n16734), .ZN(N2866) );
NAND2_X2 U12781 ( .A1(v_out[51]), .A2(n18048), .ZN(n16734) );
NAND2_X2 U12782 ( .A1(n18063), .A2(n17368), .ZN(n16733) );
NAND2_X2 U12783 ( .A1(n16735), .A2(n16736), .ZN(N2865) );
NAND2_X2 U12784 ( .A1(v_out[50]), .A2(n18048), .ZN(n16736) );
NAND2_X2 U12785 ( .A1(n18063), .A2(n17369), .ZN(n16735) );
NAND2_X2 U12786 ( .A1(n16737), .A2(n16738), .ZN(N2864) );
NAND2_X2 U12787 ( .A1(v_out[49]), .A2(n18048), .ZN(n16738) );
NAND2_X2 U12788 ( .A1(n18063), .A2(n17370), .ZN(n16737) );
NAND2_X2 U12789 ( .A1(n16739), .A2(n16740), .ZN(N2863) );
NAND2_X2 U12790 ( .A1(v_out[48]), .A2(n18048), .ZN(n16740) );
NAND2_X2 U12791 ( .A1(n18063), .A2(n17371), .ZN(n16739) );
NAND2_X2 U12792 ( .A1(n16741), .A2(n16742), .ZN(N2862) );
NAND2_X2 U12793 ( .A1(v_out[47]), .A2(n18048), .ZN(n16742) );
NAND2_X2 U12794 ( .A1(n18063), .A2(n17372), .ZN(n16741) );
NAND2_X2 U12795 ( .A1(n16743), .A2(n16744), .ZN(N2861) );
NAND2_X2 U12796 ( .A1(v_out[46]), .A2(n18048), .ZN(n16744) );
NAND2_X2 U12797 ( .A1(n18063), .A2(n17373), .ZN(n16743) );
NAND2_X2 U12798 ( .A1(n16745), .A2(n16746), .ZN(N2860) );
NAND2_X2 U12799 ( .A1(v_out[45]), .A2(n18048), .ZN(n16746) );
NAND2_X2 U12800 ( .A1(n18063), .A2(n17374), .ZN(n16745) );
NAND2_X2 U12801 ( .A1(n16747), .A2(n16748), .ZN(N2859) );
NAND2_X2 U12802 ( .A1(v_out[44]), .A2(n18048), .ZN(n16748) );
NAND2_X2 U12803 ( .A1(n18063), .A2(n18847), .ZN(n16747) );
NAND2_X2 U12804 ( .A1(n16749), .A2(n16750), .ZN(N2858) );
NAND2_X2 U12805 ( .A1(v_out[43]), .A2(n18048), .ZN(n16750) );
NAND2_X2 U12806 ( .A1(n18062), .A2(n18848), .ZN(n16749) );
NAND2_X2 U12807 ( .A1(n16751), .A2(n16752), .ZN(N2857) );
NAND2_X2 U12808 ( .A1(v_out[42]), .A2(n18048), .ZN(n16752) );
NAND2_X2 U12809 ( .A1(n18063), .A2(n18849), .ZN(n16751) );
NAND2_X2 U12810 ( .A1(n16753), .A2(n16754), .ZN(N2856) );
NAND2_X2 U12811 ( .A1(v_out[41]), .A2(n18048), .ZN(n16754) );
NAND2_X2 U12812 ( .A1(n18063), .A2(n18850), .ZN(n16753) );
NAND2_X2 U12813 ( .A1(n16755), .A2(n16756), .ZN(N2855) );
NAND2_X2 U12814 ( .A1(v_out[40]), .A2(n18048), .ZN(n16756) );
NAND2_X2 U12815 ( .A1(n18063), .A2(n18851), .ZN(n16755) );
NAND2_X2 U12816 ( .A1(n16757), .A2(n16758), .ZN(N2854) );
NAND2_X2 U12817 ( .A1(v_out[39]), .A2(n18049), .ZN(n16758) );
NAND2_X2 U12818 ( .A1(n18063), .A2(n18852), .ZN(n16757) );
NAND2_X2 U12819 ( .A1(n16759), .A2(n16760), .ZN(N2853) );
NAND2_X2 U12820 ( .A1(v_out[38]), .A2(n18049), .ZN(n16760) );
NAND2_X2 U12821 ( .A1(n18062), .A2(n18853), .ZN(n16759) );
NAND2_X2 U12822 ( .A1(n16761), .A2(n16762), .ZN(N2852) );
NAND2_X2 U12823 ( .A1(v_out[37]), .A2(n18049), .ZN(n16762) );
NAND2_X2 U12824 ( .A1(n18062), .A2(n18854), .ZN(n16761) );
NAND2_X2 U12825 ( .A1(n16763), .A2(n16764), .ZN(N2851) );
NAND2_X2 U12826 ( .A1(v_out[36]), .A2(n18049), .ZN(n16764) );
NAND2_X2 U12827 ( .A1(n18062), .A2(n18855), .ZN(n16763) );
NAND2_X2 U12828 ( .A1(n16765), .A2(n16766), .ZN(N2850) );
NAND2_X2 U12829 ( .A1(v_out[35]), .A2(n18049), .ZN(n16766) );
NAND2_X2 U12830 ( .A1(n18062), .A2(n18856), .ZN(n16765) );
NAND2_X2 U12831 ( .A1(n16767), .A2(n16768), .ZN(N2849) );
NAND2_X2 U12832 ( .A1(v_out[34]), .A2(n18049), .ZN(n16768) );
NAND2_X2 U12833 ( .A1(n18062), .A2(n18857), .ZN(n16767) );
NAND2_X2 U12834 ( .A1(n16769), .A2(n16770), .ZN(N2848) );
NAND2_X2 U12835 ( .A1(v_out[33]), .A2(n18049), .ZN(n16770) );
NAND2_X2 U12836 ( .A1(n18062), .A2(n18858), .ZN(n16769) );
NAND2_X2 U12837 ( .A1(n16771), .A2(n16772), .ZN(N2847) );
NAND2_X2 U12838 ( .A1(v_out[32]), .A2(n18049), .ZN(n16772) );
NAND2_X2 U12839 ( .A1(n18062), .A2(n18859), .ZN(n16771) );
NAND2_X2 U12840 ( .A1(n16773), .A2(n16774), .ZN(N2846) );
NAND2_X2 U12841 ( .A1(v_out[31]), .A2(n18049), .ZN(n16774) );
NAND2_X2 U12842 ( .A1(n18062), .A2(n18860), .ZN(n16773) );
NAND2_X2 U12843 ( .A1(n16775), .A2(n16776), .ZN(N2845) );
NAND2_X2 U12844 ( .A1(v_out[30]), .A2(n18049), .ZN(n16776) );
NAND2_X2 U12845 ( .A1(n18062), .A2(n18861), .ZN(n16775) );
NAND2_X2 U12846 ( .A1(n16777), .A2(n16778), .ZN(N2844) );
NAND2_X2 U12847 ( .A1(v_out[29]), .A2(n18049), .ZN(n16778) );
NAND2_X2 U12848 ( .A1(n18062), .A2(n18862), .ZN(n16777) );
NAND2_X2 U12849 ( .A1(n16779), .A2(n16780), .ZN(N2843) );
NAND2_X2 U12850 ( .A1(v_out[28]), .A2(n18049), .ZN(n16780) );
NAND2_X2 U12851 ( .A1(n18062), .A2(n18863), .ZN(n16779) );
NAND2_X2 U12852 ( .A1(n16781), .A2(n16782), .ZN(N2842) );
NAND2_X2 U12853 ( .A1(v_out[27]), .A2(n18049), .ZN(n16782) );
NAND2_X2 U12854 ( .A1(n18062), .A2(n18864), .ZN(n16781) );
NAND2_X2 U12855 ( .A1(n16783), .A2(n16784), .ZN(N2841) );
NAND2_X2 U12856 ( .A1(v_out[26]), .A2(n18049), .ZN(n16784) );
NAND2_X2 U12857 ( .A1(n18062), .A2(n18865), .ZN(n16783) );
NAND2_X2 U12858 ( .A1(n16785), .A2(n16786), .ZN(N2840) );
NAND2_X2 U12859 ( .A1(v_out[25]), .A2(n18049), .ZN(n16786) );
NAND2_X2 U12860 ( .A1(n18062), .A2(n18866), .ZN(n16785) );
NAND2_X2 U12861 ( .A1(n16787), .A2(n16788), .ZN(N2839) );
NAND2_X2 U12862 ( .A1(v_out[24]), .A2(n18049), .ZN(n16788) );
NAND2_X2 U12863 ( .A1(n18062), .A2(n18867), .ZN(n16787) );
NAND2_X2 U12864 ( .A1(n16789), .A2(n16790), .ZN(N2838) );
NAND2_X2 U12865 ( .A1(v_out[23]), .A2(n18049), .ZN(n16790) );
NAND2_X2 U12866 ( .A1(n18062), .A2(n18868), .ZN(n16789) );
NAND2_X2 U12867 ( .A1(n16791), .A2(n16792), .ZN(N2837) );
NAND2_X2 U12868 ( .A1(v_out[22]), .A2(n18049), .ZN(n16792) );
NAND2_X2 U12869 ( .A1(n18062), .A2(n18869), .ZN(n16791) );
NAND2_X2 U12870 ( .A1(n16793), .A2(n16794), .ZN(N2836) );
NAND2_X2 U12871 ( .A1(v_out[21]), .A2(n18050), .ZN(n16794) );
NAND2_X2 U12872 ( .A1(n18062), .A2(n18870), .ZN(n16793) );
NAND2_X2 U12873 ( .A1(n16795), .A2(n16796), .ZN(N2835) );
NAND2_X2 U12874 ( .A1(v_out[20]), .A2(n18050), .ZN(n16796) );
NAND2_X2 U12875 ( .A1(n18062), .A2(n18871), .ZN(n16795) );
NAND2_X2 U12876 ( .A1(n16797), .A2(n16798), .ZN(N2834) );
NAND2_X2 U12877 ( .A1(v_out[19]), .A2(n18050), .ZN(n16798) );
NAND2_X2 U12878 ( .A1(n18062), .A2(n18872), .ZN(n16797) );
NAND2_X2 U12879 ( .A1(n16799), .A2(n16800), .ZN(N2833) );
NAND2_X2 U12880 ( .A1(v_out[18]), .A2(n18050), .ZN(n16800) );
NAND2_X2 U12881 ( .A1(n18061), .A2(n18873), .ZN(n16799) );
NAND2_X2 U12882 ( .A1(n16801), .A2(n16802), .ZN(N2832) );
NAND2_X2 U12883 ( .A1(v_out[17]), .A2(n18050), .ZN(n16802) );
NAND2_X2 U12884 ( .A1(n18061), .A2(n18874), .ZN(n16801) );
NAND2_X2 U12885 ( .A1(n16803), .A2(n16804), .ZN(N2831) );
NAND2_X2 U12886 ( .A1(v_out[16]), .A2(n18050), .ZN(n16804) );
NAND2_X2 U12887 ( .A1(n18061), .A2(n18875), .ZN(n16803) );
NAND2_X2 U12888 ( .A1(n16805), .A2(n16806), .ZN(N2830) );
NAND2_X2 U12889 ( .A1(v_out[15]), .A2(n18050), .ZN(n16806) );
NAND2_X2 U12890 ( .A1(n18061), .A2(n18876), .ZN(n16805) );
NAND2_X2 U12891 ( .A1(n16807), .A2(n16808), .ZN(N2829) );
NAND2_X2 U12892 ( .A1(v_out[14]), .A2(n18050), .ZN(n16808) );
NAND2_X2 U12893 ( .A1(n18061), .A2(n18877), .ZN(n16807) );
NAND2_X2 U12894 ( .A1(n16809), .A2(n16810), .ZN(N2828) );
NAND2_X2 U12895 ( .A1(v_out[13]), .A2(n18050), .ZN(n16810) );
NAND2_X2 U12896 ( .A1(n18061), .A2(n18878), .ZN(n16809) );
NAND2_X2 U12897 ( .A1(n16811), .A2(n16812), .ZN(N2827) );
NAND2_X2 U12898 ( .A1(v_out[12]), .A2(n18050), .ZN(n16812) );
NAND2_X2 U12899 ( .A1(n18061), .A2(n18879), .ZN(n16811) );
NAND2_X2 U12900 ( .A1(n16813), .A2(n16814), .ZN(N2826) );
NAND2_X2 U12901 ( .A1(v_out[11]), .A2(n18050), .ZN(n16814) );
NAND2_X2 U12902 ( .A1(n18061), .A2(n18880), .ZN(n16813) );
NAND2_X2 U12903 ( .A1(n16815), .A2(n16816), .ZN(N2825) );
NAND2_X2 U12904 ( .A1(v_out[10]), .A2(n18050), .ZN(n16816) );
NAND2_X2 U12905 ( .A1(n18061), .A2(n18881), .ZN(n16815) );
NAND2_X2 U12906 ( .A1(n16817), .A2(n16818), .ZN(N2824) );
NAND2_X2 U12907 ( .A1(v_out[9]), .A2(n18050), .ZN(n16818) );
NAND2_X2 U12908 ( .A1(n18061), .A2(n18882), .ZN(n16817) );
NAND2_X2 U12909 ( .A1(n16819), .A2(n16820), .ZN(N2823) );
NAND2_X2 U12910 ( .A1(v_out[8]), .A2(n18050), .ZN(n16820) );
NAND2_X2 U12911 ( .A1(n18061), .A2(n18883), .ZN(n16819) );
NAND2_X2 U12912 ( .A1(n16821), .A2(n16822), .ZN(N2822) );
NAND2_X2 U12913 ( .A1(v_out[7]), .A2(n18050), .ZN(n16822) );
NAND2_X2 U12914 ( .A1(n18061), .A2(n18884), .ZN(n16821) );
NAND2_X2 U12915 ( .A1(n16823), .A2(n16824), .ZN(N2821) );
NAND2_X2 U12916 ( .A1(v_out[6]), .A2(n18050), .ZN(n16824) );
NAND2_X2 U12917 ( .A1(n18061), .A2(n18885), .ZN(n16823) );
NAND2_X2 U12918 ( .A1(n16825), .A2(n16826), .ZN(N2820) );
NAND2_X2 U12919 ( .A1(v_out[5]), .A2(n18050), .ZN(n16826) );
NAND2_X2 U12920 ( .A1(n18061), .A2(n18886), .ZN(n16825) );
NAND2_X2 U12921 ( .A1(n16827), .A2(n16828), .ZN(N2819) );
NAND2_X2 U12922 ( .A1(v_out[4]), .A2(n18050), .ZN(n16828) );
NAND2_X2 U12923 ( .A1(n18061), .A2(n18887), .ZN(n16827) );
NAND2_X2 U12924 ( .A1(n16829), .A2(n16830), .ZN(N2818) );
NAND2_X2 U12925 ( .A1(v_out[3]), .A2(n18051), .ZN(n16830) );
NAND2_X2 U12926 ( .A1(n18061), .A2(n18888), .ZN(n16829) );
NAND2_X2 U12927 ( .A1(n16831), .A2(n16832), .ZN(N2817) );
NAND2_X2 U12928 ( .A1(v_out[2]), .A2(n18051), .ZN(n16832) );
NAND2_X2 U12929 ( .A1(n18061), .A2(n18889), .ZN(n16831) );
NAND2_X2 U12930 ( .A1(n16833), .A2(n16834), .ZN(N2816) );
NAND2_X2 U12931 ( .A1(v_out[1]), .A2(n18047), .ZN(n16834) );
NAND2_X2 U12932 ( .A1(n18061), .A2(n18890), .ZN(n16833) );
NAND2_X2 U12933 ( .A1(n16835), .A2(n16836), .ZN(N2815) );
NAND2_X2 U12934 ( .A1(v_out[0]), .A2(n18043), .ZN(n16836) );
NAND2_X2 U12935 ( .A1(n18059), .A2(n18891), .ZN(n16835) );
NAND2_X2 U12942 ( .A1(n18845), .A2(n18627), .ZN(n11976) );
NAND2_X2 U12944 ( .A1(n11973), .A2(n18600), .ZN(n16837) );
AND4_X2 U12945 ( .A1(n18628), .A2(n18631), .A3(n18629), .A4(n18626), .ZN(n11973) );
DFFR_X1 enc_byte_cnt_reg_4_ ( .D(n5437), .CK(clk), .RN(n18632), .Q(enc_byte_cnt[4]), .QN(n5374) );
DFFR_X1 enc_byte_cnt_reg_2_ ( .D(n5439), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[2]), .QN(n5376) );
DFFR_X1 enc_byte_cnt_reg_1_ ( .D(n5440), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[1]), .QN(n5377) );
DFFR_X1 enc_byte_cnt_reg_3_ ( .D(n5438), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[3]), .QN(n5375) );
DFFR_X1 enc_byte_cnt_reg_5_ ( .D(n5436), .CK(clk), .RN(n18632), .Q(enc_byte_cnt[5]), .QN() );
DFFR_X1 enc_byte_cnt_reg_0_ ( .D(n5441), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[0]), .QN(n5378) );
DFFR_X1 enc_byte_cnt_reg_16_ ( .D(n5425), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[16]), .QN(n5362) );
DFFR_X1 enc_byte_cnt_reg_8_ ( .D(n5433), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[8]), .QN() );
DFFR_X1 enc_byte_cnt_reg_6_ ( .D(n5435), .CK(clk), .RN(n18632), .Q(enc_byte_cnt[6]), .QN() );
DFFR_X1 enc_byte_cnt_reg_9_ ( .D(n5432), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[9]), .QN() );
DFFR_X1 enc_byte_cnt_reg_12_ ( .D(n5429), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[12]), .QN() );
DFFR_X1 enc_byte_cnt_reg_7_ ( .D(n5434), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[7]), .QN() );
DFFR_X1 enc_byte_cnt_reg_24_ ( .D(n5417), .CK(clk), .RN(n18632), .Q(enc_byte_cnt[24]), .QN() );
DFFR_X1 enc_byte_cnt_reg_10_ ( .D(n5431), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[10]), .QN() );
DFFR_X1 enc_byte_cnt_reg_13_ ( .D(n5428), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[13]), .QN(n5365) );
DFFR_X1 enc_byte_cnt_reg_17_ ( .D(n5424), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[17]), .QN(n5361) );
DFFR_X1 enc_byte_cnt_reg_20_ ( .D(n5421), .CK(clk), .RN(n18632), .Q(enc_byte_cnt[20]), .QN(n5358) );
DFFR_X1 enc_byte_cnt_reg_21_ ( .D(n5420), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[21]), .QN() );
DFFR_X1 enc_byte_cnt_reg_18_ ( .D(n5423), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[18]), .QN(n5360) );
DFFR_X1 aad_byte_cnt_reg_4_ ( .D(n6016), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[4]), .QN() );
DFFR_X1 aad_byte_cnt_reg_2_ ( .D(n6018), .CK(clk), .RN(n17820), .Q(aad_byte_cnt[2]), .QN() );
DFFR_X1 aad_byte_cnt_reg_1_ ( .D(n6019), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[1]), .QN() );
DFFR_X1 aad_byte_cnt_reg_3_ ( .D(n6017), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[3]), .QN() );
DFFR_X1 aad_byte_cnt_reg_12_ ( .D(n6008), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[12]), .QN() );
DFFR_X1 aad_byte_cnt_reg_10_ ( .D(n6010), .CK(clk), .RN(n18632), .Q(aad_byte_cnt[10]), .QN() );
DFFR_X1 aad_byte_cnt_reg_9_ ( .D(n6011), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[9]), .QN() );
DFFR_X1 aad_byte_cnt_reg_8_ ( .D(n6012), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[8]), .QN() );
DFFR_X1 aad_byte_cnt_reg_7_ ( .D(n6013), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[7]), .QN() );
DFFR_X1 aad_byte_cnt_reg_6_ ( .D(n6014), .CK(clk), .RN(n17819), .Q(aad_byte_cnt[6]), .QN() );
DFFR_X1 aad_byte_cnt_reg_5_ ( .D(n6015), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[5]), .QN() );
DFFR_X1 aad_byte_cnt_reg_0_ ( .D(n6020), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[0]), .QN() );
DFFR_X1 enc_byte_cnt_reg_14_ ( .D(n5427), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[14]), .QN(n5364) );
DFFR_X1 aad_byte_cnt_reg_16_ ( .D(n6004), .CK(clk), .RN(n17820), .Q(aad_byte_cnt[16]), .QN() );
DFFR_X1 aad_byte_cnt_reg_24_ ( .D(n5996), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[24]), .QN() );
DFFR_X1 aad_byte_cnt_reg_21_ ( .D(n5999), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[21]), .QN() );
DFFR_X1 aad_byte_cnt_reg_20_ ( .D(n6000), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[20]), .QN() );
DFFR_X1 aad_byte_cnt_reg_18_ ( .D(n6002), .CK(clk), .RN(n18632), .Q(aad_byte_cnt[18]), .QN() );
DFFR_X1 aad_byte_cnt_reg_17_ ( .D(n6003), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[17]), .QN() );
DFFR_X1 aad_byte_cnt_reg_14_ ( .D(n6006), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[14]), .QN() );
DFFR_X1 aad_byte_cnt_reg_13_ ( .D(n6007), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[13]), .QN() );
DFFR_X1 enc_byte_cnt_reg_28_ ( .D(n5413), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[28]), .QN() );
DFFR_X1 enc_byte_cnt_reg_11_ ( .D(n5430), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[11]), .QN() );
DFFR_X1 aad_byte_cnt_reg_11_ ( .D(n6009), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[11]), .QN() );
DFFR_X1 aad_byte_cnt_reg_28_ ( .D(n5992), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[28]), .QN() );
DFFR_X1 enc_byte_cnt_reg_25_ ( .D(n5416), .CK(clk), .RN(n17819), .Q(enc_byte_cnt[25]), .QN() );
DFFR_X1 aad_byte_cnt_reg_25_ ( .D(n5995), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[25]), .QN() );
DFFR_X1 enc_byte_cnt_reg_15_ ( .D(n5426), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[15]), .QN(n5363) );
DFFR_X1 aad_byte_cnt_reg_15_ ( .D(n6005), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[15]), .QN() );
DFFR_X1 enc_byte_cnt_reg_36_ ( .D(n5405), .CK(clk), .RN(n17820), .Q(enc_byte_cnt[36]), .QN(n5342) );
DFFR_X1 aad_byte_cnt_reg_36_ ( .D(n5984), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[36]), .QN() );
DFFR_X1 aad_byte_cnt_reg_19_ ( .D(n6001), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[19]), .QN() );
DFFR_X1 enc_byte_cnt_reg_54_ ( .D(n5387), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[54]), .QN() );
DFFR_X1 aad_byte_cnt_reg_54_ ( .D(n5966), .CK(clk), .RN(n18632), .Q(aad_byte_cnt[54]), .QN() );
DFFR_X1 enc_byte_cnt_reg_19_ ( .D(n5422), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[19]), .QN(n5359) );
DFFR_X1 enc_byte_cnt_reg_22_ ( .D(n5419), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[22]), .QN() );
DFFR_X1 aad_byte_cnt_reg_22_ ( .D(n5998), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[22]), .QN() );
DFFR_X1 aad_byte_cnt_reg_29_ ( .D(n5991), .CK(clk), .RN(n17822), .Q(aad_byte_cnt[29]), .QN() );
DFFR_X1 enc_byte_cnt_reg_49_ ( .D(n5392), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[49]), .QN(n5329) );
DFFR_X1 enc_byte_cnt_reg_29_ ( .D(n5412), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[29]), .QN(n5349) );
DFFR_X1 enc_byte_cnt_reg_53_ ( .D(n5388), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[53]), .QN() );
DFFR_X1 enc_byte_cnt_reg_60_ ( .D(n5381), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[60]), .QN() );
DFFR_X1 aad_byte_cnt_reg_60_ ( .D(n5960), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[60]), .QN() );
DFFR_X1 aad_byte_cnt_reg_49_ ( .D(n5971), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[49]), .QN() );
DFFR_X1 aad_byte_cnt_reg_53_ ( .D(n5967), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[53]), .QN() );
DFFR_X1 aad_byte_cnt_reg_52_ ( .D(n5968), .CK(clk), .RN(n17819), .Q(aad_byte_cnt[52]), .QN() );
DFFR_X1 aad_byte_cnt_reg_51_ ( .D(n5969), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[51]), .QN() );
DFFR_X1 enc_byte_cnt_reg_30_ ( .D(n5411), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[30]), .QN(n5348) );
DFFR_X1 enc_byte_cnt_reg_52_ ( .D(n5389), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[52]), .QN(n5326) );
DFFR_X1 enc_byte_cnt_reg_51_ ( .D(n5390), .CK(clk), .RN(n17820), .Q(enc_byte_cnt[51]), .QN(n5327) );
DFFR_X1 enc_byte_cnt_reg_26_ ( .D(n5415), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[26]), .QN() );
DFFR_X1 aad_byte_cnt_reg_26_ ( .D(n5994), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[26]), .QN() );
DFFR_X1 aad_byte_cnt_reg_30_ ( .D(n5990), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[30]), .QN() );
DFFR_X1 enc_byte_cnt_reg_59_ ( .D(n5382), .CK(clk), .RN(n18632), .Q(enc_byte_cnt[59]), .QN() );
DFFR_X1 enc_byte_cnt_reg_58_ ( .D(n5383), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[58]), .QN() );
DFFR_X1 enc_byte_cnt_reg_57_ ( .D(n5384), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[57]), .QN() );
DFFR_X1 enc_byte_cnt_reg_56_ ( .D(n5385), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[56]), .QN() );
DFFR_X1 aad_byte_cnt_reg_59_ ( .D(n5961), .CK(clk), .RN(n17836), .Q(aad_byte_cnt[59]), .QN() );
DFFR_X1 aad_byte_cnt_reg_58_ ( .D(n5962), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[58]), .QN() );
DFFR_X1 aad_byte_cnt_reg_57_ ( .D(n5963), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[57]), .QN() );
DFFR_X1 aad_byte_cnt_reg_56_ ( .D(n5964), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[56]), .QN() );
DFFR_X1 enc_byte_cnt_reg_37_ ( .D(n5404), .CK(clk), .RN(n17822), .Q(enc_byte_cnt[37]), .QN() );
DFFR_X1 aad_byte_cnt_reg_37_ ( .D(n5983), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[37]), .QN() );
DFFR_X1 enc_byte_cnt_reg_32_ ( .D(n5409), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[32]), .QN(n5346) );
DFFR_X1 aad_byte_cnt_reg_32_ ( .D(n5988), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[32]), .QN() );
DFFR_X1 enc_byte_cnt_reg_55_ ( .D(n5386), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[55]), .QN() );
DFFR_X1 aad_byte_cnt_reg_55_ ( .D(n5965), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[55]), .QN() );
DFFR_X1 enc_byte_cnt_reg_34_ ( .D(n5407), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[34]), .QN(n5344) );
DFFR_X1 enc_byte_cnt_reg_33_ ( .D(n5408), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[33]), .QN(n5345) );
DFFR_X1 aad_byte_cnt_reg_34_ ( .D(n5986), .CK(clk), .RN(n17819), .Q(aad_byte_cnt[34]), .QN() );
DFFR_X1 aad_byte_cnt_reg_33_ ( .D(n5987), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[33]), .QN() );
DFFR_X1 enc_byte_cnt_reg_38_ ( .D(n5403), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[38]), .QN() );
DFFR_X1 aad_byte_cnt_reg_38_ ( .D(n5982), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[38]), .QN() );
DFFR_X1 enc_byte_cnt_reg_23_ ( .D(n5418), .CK(clk), .RN(n17823), .Q(enc_byte_cnt[23]), .QN() );
DFFR_X1 aad_byte_cnt_reg_23_ ( .D(n5997), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[23]), .QN() );
DFFR_X1 enc_byte_cnt_reg_50_ ( .D(n5391), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[50]), .QN(n5328) );
DFFR_X1 enc_byte_cnt_reg_31_ ( .D(n5410), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[31]), .QN(n5347) );
DFFR_X1 aad_byte_cnt_reg_50_ ( .D(n5970), .CK(clk), .RN(n17832), .Q(aad_byte_cnt[50]), .QN() );
DFFR_X1 enc_byte_cnt_reg_35_ ( .D(n5406), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[35]), .QN(n5343) );
DFFR_X1 aad_byte_cnt_reg_35_ ( .D(n5985), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[35]), .QN() );
DFFR_X1 aad_byte_cnt_reg_31_ ( .D(n5989), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[31]), .QN() );
DFFR_X1 enc_byte_cnt_reg_27_ ( .D(n5414), .CK(clk), .RN(n17820), .Q(enc_byte_cnt[27]), .QN() );
DFFR_X1 aad_byte_cnt_reg_27_ ( .D(n5993), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[27]), .QN() );
DFFR_X1 aad_byte_cnt_reg_48_ ( .D(n5972), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[48]), .QN() );
DFFR_X1 enc_byte_cnt_reg_46_ ( .D(n5395), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[46]), .QN(n5332) );
DFFR_X1 aad_byte_cnt_reg_46_ ( .D(n5974), .CK(clk), .RN(n18632), .Q(aad_byte_cnt[46]), .QN() );
DFFR_X1 enc_byte_cnt_reg_48_ ( .D(n5393), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[48]), .QN(n5330) );
DFFR_X1 enc_byte_cnt_reg_47_ ( .D(n5394), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[47]), .QN(n5331) );
DFFR_X1 enc_byte_cnt_reg_43_ ( .D(n5398), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[43]), .QN() );
DFFR_X1 aad_byte_cnt_reg_47_ ( .D(n5973), .CK(clk), .RN(n17836), .Q(aad_byte_cnt[47]), .QN() );
DFFR_X1 aad_byte_cnt_reg_43_ ( .D(n5977), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[43]), .QN() );
DFFR_X1 enc_byte_cnt_reg_39_ ( .D(n5402), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[39]), .QN() );
DFFR_X1 aad_byte_cnt_reg_39_ ( .D(n5981), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[39]), .QN() );
DFFR_X1 enc_byte_cnt_reg_42_ ( .D(n5399), .CK(clk), .RN(n17822), .Q(enc_byte_cnt[42]), .QN() );
DFFR_X1 aad_byte_cnt_reg_42_ ( .D(n5978), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[42]), .QN() );
DFFR_X1 enc_byte_cnt_reg_44_ ( .D(n5397), .CK(clk), .RN(n17752), .Q(enc_byte_cnt[44]), .QN() );
DFFR_X1 enc_byte_cnt_reg_41_ ( .D(n5400), .CK(clk), .RN(n17751), .Q(enc_byte_cnt[41]), .QN() );
DFFR_X1 enc_byte_cnt_reg_40_ ( .D(n5401), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[40]), .QN() );
DFFR_X1 aad_byte_cnt_reg_45_ ( .D(n5975), .CK(clk), .RN(n17753), .Q(aad_byte_cnt[45]), .QN() );
DFFR_X1 aad_byte_cnt_reg_44_ ( .D(n5976), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[44]), .QN() );
DFFR_X1 aad_byte_cnt_reg_41_ ( .D(n5979), .CK(clk), .RN(n17751), .Q(aad_byte_cnt[41]), .QN() );
DFFR_X1 aad_byte_cnt_reg_40_ ( .D(n5980), .CK(clk), .RN(n17819), .Q(aad_byte_cnt[40]), .QN() );
DFFR_X1 enc_byte_cnt_reg_45_ ( .D(n5396), .CK(clk), .RN(n17753), .Q(enc_byte_cnt[45]), .QN(n5333) );
DFFS_X1 state_reg_0_ ( .D(n6283), .CK(clk), .SN(n17836), .Q(state[0]), .QN(n18611) );
DFFR_X1 state_reg_2_ ( .D(n6284), .CK(clk), .RN(n17824), .Q(state[2]), .QN(n18630) );
DFFR_X1 enc_byte_cnt_reg_63_ ( .D(n5442), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[63]), .QN() );
DFFR_X1 aad_byte_cnt_reg_63_ ( .D(n6021), .CK(clk), .RN(n17823), .Q(aad_byte_cnt[63]), .QN() );
DFFR_X1 enc_byte_cnt_reg_62_ ( .D(n5379), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[62]), .QN() );
DFFR_X1 enc_byte_cnt_reg_61_ ( .D(n5380), .CK(clk), .RN(n17824), .Q(enc_byte_cnt[61]), .QN() );
DFFR_X1 aad_byte_cnt_reg_62_ ( .D(n5958), .CK(clk), .RN(n17752), .Q(aad_byte_cnt[62]), .QN() );
DFFR_X1 aad_byte_cnt_reg_61_ ( .D(n5959), .CK(clk), .RN(n17823), .Q(aad_byte_cnt[61]), .QN() );
DFFR_X1 state_reg_5_ ( .D(n6286), .CK(clk), .RN(n17818), .Q(state[5]), .QN(n18600) );
DFFR_X1 state_reg_4_ ( .D(n6285), .CK(clk), .RN(n18632), .Q(state[4]), .QN(n18629) );
DFFR_X1 state_reg_1_ ( .D(n6292), .CK(clk), .RN(n17825), .Q(state[1]), .QN(n18631) );
DFFR_X1 state_reg_3_ ( .D(n6287), .CK(clk), .RN(n17753), .Q(state[3]), .QN(n18078) );
DFFR_X1 state_reg_8_ ( .D(n6293), .CK(clk), .RN(n17824), .Q(state[8]), .QN(n18079) );
DFFR_X1 state_reg_6_ ( .D(n6288), .CK(clk), .RN(n17824), .Q(state[6]), .QN(n18626) );
DFFR_X1 state_reg_9_ ( .D(n6294), .CK(clk), .RN(n17824), .Q(state[9]), .QN(n18080) );
DFFR_X1 state_reg_7_ ( .D(n6289), .CK(clk), .RN(n17824), .Q(state[7]), .QN(n18601) );
DFFR_X1 H_reg_2_ ( .D(n6152), .CK(clk), .RN(n17751), .Q(n18889), .QN() );
DFFR_X1 H_reg_1_ ( .D(n6153), .CK(clk), .RN(n17823), .Q(n18890), .QN() );
DFFR_X1 H_reg_0_ ( .D(n6154), .CK(clk), .RN(n17753), .Q(n18891), .QN() );
DFFR_X1 H_reg_44_ ( .D(n6110), .CK(clk), .RN(n17752), .Q(n18847), .QN() );
DFFR_X1 H_reg_43_ ( .D(n6111), .CK(clk), .RN(n17751), .Q(n18848), .QN() );
DFFR_X1 H_reg_42_ ( .D(n6112), .CK(clk), .RN(n17832), .Q(n18849), .QN() );
DFFR_X1 H_reg_41_ ( .D(n6113), .CK(clk), .RN(n17753), .Q(n18850), .QN() );
DFFR_X1 H_reg_40_ ( .D(n6114), .CK(clk), .RN(n17752), .Q(n18851), .QN() );
DFFR_X1 H_reg_39_ ( .D(n6115), .CK(clk), .RN(n17751), .Q(n18852), .QN() );
DFFR_X1 H_reg_38_ ( .D(n6116), .CK(clk), .RN(n17820), .Q(n18853), .QN() );
DFFR_X1 H_reg_37_ ( .D(n6117), .CK(clk), .RN(n17753), .Q(n18854), .QN() );
DFFR_X1 H_reg_36_ ( .D(n6118), .CK(clk), .RN(n17752), .Q(n18855), .QN() );
DFFR_X1 H_reg_35_ ( .D(n6119), .CK(clk), .RN(n17751), .Q(n18856), .QN() );
DFFR_X1 H_reg_34_ ( .D(n6120), .CK(clk), .RN(n18632), .Q(n18857), .QN() );
DFFR_X1 H_reg_33_ ( .D(n6121), .CK(clk), .RN(n17753), .Q(n18858), .QN() );
DFFR_X1 H_reg_32_ ( .D(n6122), .CK(clk), .RN(n17752), .Q(n18859), .QN() );
DFFR_X1 H_reg_31_ ( .D(n6123), .CK(clk), .RN(n17751), .Q(n18860), .QN() );
DFFR_X1 H_reg_30_ ( .D(n6124), .CK(clk), .RN(n17836), .Q(n18861), .QN() );
DFFR_X1 H_reg_29_ ( .D(n6125), .CK(clk), .RN(n17753), .Q(n18862), .QN() );
DFFR_X1 H_reg_28_ ( .D(n6126), .CK(clk), .RN(n17752), .Q(n18863), .QN() );
DFFR_X1 H_reg_27_ ( .D(n6127), .CK(clk), .RN(n17751), .Q(n18864), .QN() );
DFFR_X1 H_reg_26_ ( .D(n6128), .CK(clk), .RN(n17834), .Q(n18865), .QN() );
DFFR_X1 H_reg_25_ ( .D(n6129), .CK(clk), .RN(n17753), .Q(n18866), .QN() );
DFFR_X1 H_reg_24_ ( .D(n6130), .CK(clk), .RN(n17752), .Q(n18867), .QN() );
DFFR_X1 H_reg_23_ ( .D(n6131), .CK(clk), .RN(n17751), .Q(n18868), .QN() );
DFFR_X1 H_reg_22_ ( .D(n6132), .CK(clk), .RN(n17822), .Q(n18869), .QN() );
DFFR_X1 H_reg_21_ ( .D(n6133), .CK(clk), .RN(n17753), .Q(n18870), .QN() );
DFFR_X1 H_reg_20_ ( .D(n6134), .CK(clk), .RN(n17752), .Q(n18871), .QN() );
DFFR_X1 H_reg_19_ ( .D(n6135), .CK(clk), .RN(n17751), .Q(n18872), .QN() );
DFFR_X1 H_reg_18_ ( .D(n6136), .CK(clk), .RN(n17828), .Q(n18873), .QN() );
DFFR_X1 H_reg_17_ ( .D(n6137), .CK(clk), .RN(n17753), .Q(n18874), .QN() );
DFFR_X1 H_reg_16_ ( .D(n6138), .CK(clk), .RN(n17752), .Q(n18875), .QN() );
DFFR_X1 H_reg_15_ ( .D(n6139), .CK(clk), .RN(n17751), .Q(n18876), .QN() );
DFFR_X1 H_reg_14_ ( .D(n6140), .CK(clk), .RN(n17824), .Q(n18877), .QN() );
DFFR_X1 H_reg_13_ ( .D(n6141), .CK(clk), .RN(n17753), .Q(n18878), .QN() );
DFFR_X1 H_reg_12_ ( .D(n6142), .CK(clk), .RN(n17752), .Q(n18879), .QN() );
DFFR_X1 H_reg_11_ ( .D(n6143), .CK(clk), .RN(n17751), .Q(n18880), .QN() );
DFFR_X1 H_reg_10_ ( .D(n6144), .CK(clk), .RN(n17825), .Q(n18881), .QN() );
DFFR_X1 H_reg_9_ ( .D(n6145), .CK(clk), .RN(n17753), .Q(n18882), .QN() );
DFFR_X1 H_reg_8_ ( .D(n6146), .CK(clk), .RN(n17752), .Q(n18883), .QN() );
DFFR_X1 H_reg_7_ ( .D(n6147), .CK(clk), .RN(n17751), .Q(n18884), .QN() );
DFFR_X1 H_reg_6_ ( .D(n6148), .CK(clk), .RN(n17829), .Q(n18885), .QN() );
DFFR_X1 H_reg_5_ ( .D(n6149), .CK(clk), .RN(n17753), .Q(n18886), .QN() );
DFFR_X1 H_reg_4_ ( .D(n6150), .CK(clk), .RN(n17752), .Q(n18887), .QN() );
DFFR_X1 H_reg_3_ ( .D(n6151), .CK(clk), .RN(n17751), .Q(n18888), .QN() );
DFFR_X1 EkY0_reg_50_ ( .D(n6232), .CK(clk), .RN(n17819), .Q(), .QN(n17179));
DFFR_X1 EkY0_reg_49_ ( .D(n6233), .CK(clk), .RN(n17753), .Q(), .QN(n17181));
DFFR_X1 EkY0_reg_48_ ( .D(n6234), .CK(clk), .RN(n17752), .Q(), .QN(n17183));
DFFR_X1 EkY0_reg_47_ ( .D(n6235), .CK(clk), .RN(n17751), .Q(), .QN(n17185));
DFFR_X1 EkY0_reg_46_ ( .D(n6236), .CK(clk), .RN(n17823), .Q(), .QN(n17187));
DFFR_X1 EkY0_reg_45_ ( .D(n6237), .CK(clk), .RN(n17753), .Q(), .QN(n17189));
DFFR_X1 EkY0_reg_44_ ( .D(n6238), .CK(clk), .RN(n17752), .Q(), .QN(n17191));
DFFR_X1 EkY0_reg_42_ ( .D(n6240), .CK(clk), .RN(n17751), .Q(), .QN(n17195));
DFFR_X1 EkY0_reg_41_ ( .D(n6241), .CK(clk), .RN(n17833), .Q(), .QN(n17197));
DFFR_X1 EkY0_reg_40_ ( .D(n6242), .CK(clk), .RN(n17753), .Q(), .QN(n17199));
DFFR_X1 EkY0_reg_39_ ( .D(n6243), .CK(clk), .RN(n17752), .Q(), .QN(n17201));
DFFR_X1 EkY0_reg_127_ ( .D(n6155), .CK(clk), .RN(n17751), .Q(), .QN(n17025));
DFFR_X1 EkY0_reg_124_ ( .D(n6158), .CK(clk), .RN(n17832), .Q(), .QN(n17031));
DFFR_X1 EkY0_reg_122_ ( .D(n6160), .CK(clk), .RN(n17753), .Q(), .QN(n17035));
DFFR_X1 EkY0_reg_2_ ( .D(n6280), .CK(clk), .RN(n17752), .Q(), .QN(n17275) );
DFFR_X1 EkY0_reg_1_ ( .D(n6281), .CK(clk), .RN(n17751), .Q(), .QN(n17277) );
DFFR_X1 EkY0_reg_22_ ( .D(n6260), .CK(clk), .RN(n17820), .Q(), .QN(n17235));
DFFR_X1 EkY0_reg_21_ ( .D(n6261), .CK(clk), .RN(n17753), .Q(), .QN(n17237));
DFFR_X1 EkY0_reg_19_ ( .D(n6263), .CK(clk), .RN(n17752), .Q(), .QN(n17241));
DFFR_X1 EkY0_reg_18_ ( .D(n6264), .CK(clk), .RN(n17751), .Q(), .QN(n17243));
DFF_X1 gfm_result_reg_2_ ( .D(n5827), .CK(clk), .Q(n18897), .QN(n17274) );
DFF_X1 gfm_result_reg_0_ ( .D(n5829), .CK(clk), .Q(n18895), .QN(n17278) );
DFF_X1 gfm_result_reg_3_ ( .D(n5826), .CK(clk), .Q(n18898), .QN(n17272) );
DFF_X1 gfm_result_reg_33_ ( .D(n5796), .CK(clk), .Q(n18928), .QN() );
DFF_X1 gfm_result_reg_14_ ( .D(n5815), .CK(clk), .Q(n18909), .QN() );
DFF_X1 gfm_result_reg_4_ ( .D(n5825), .CK(clk), .Q(n18899), .QN(n17270) );
DFF_X1 gfm_result_reg_36_ ( .D(n5793), .CK(clk), .Q(n18931), .QN() );
DFF_X1 gfm_result_reg_40_ ( .D(n5789), .CK(clk), .Q(n18935), .QN() );
DFF_X1 gfm_result_reg_39_ ( .D(n5790), .CK(clk), .Q(n18934), .QN() );
DFF_X1 gfm_result_reg_41_ ( .D(n5788), .CK(clk), .Q(n18936), .QN() );
DFF_X1 gfm_result_reg_38_ ( .D(n5791), .CK(clk), .Q(n18933), .QN() );
DFF_X1 gfm_result_reg_37_ ( .D(n5792), .CK(clk), .Q(n18932), .QN() );
DFF_X1 gfm_result_reg_43_ ( .D(n5786), .CK(clk), .Q(n18938), .QN() );
DFF_X1 gfm_result_reg_42_ ( .D(n5787), .CK(clk), .Q(n18937), .QN() );
DFF_X1 gfm_result_reg_44_ ( .D(n5785), .CK(clk), .Q(n18939), .QN() );
DFF_X1 gfm_result_reg_45_ ( .D(n5784), .CK(clk), .Q(n18940), .QN() );
DFF_X1 gfm_result_reg_35_ ( .D(n5794), .CK(clk), .Q(n18930), .QN() );
DFF_X1 gfm_result_reg_13_ ( .D(n5816), .CK(clk), .Q(n18908), .QN() );
DFF_X1 gfm_result_reg_1_ ( .D(n5828), .CK(clk), .Q(n18896), .QN(n17276) );
DFF_X1 gfm_result_reg_6_ ( .D(n5823), .CK(clk), .Q(n18901), .QN(n17266) );
DFF_X1 gfm_result_reg_5_ ( .D(n5824), .CK(clk), .Q(n18900), .QN(n17268) );
DFF_X1 gfm_result_reg_7_ ( .D(n5822), .CK(clk), .Q(n18902), .QN(n17264) );
DFF_X1 gfm_result_reg_8_ ( .D(n5821), .CK(clk), .Q(n18903), .QN() );
DFF_X1 gfm_result_reg_9_ ( .D(n5820), .CK(clk), .Q(n18904), .QN() );
DFF_X1 gfm_result_reg_30_ ( .D(n5799), .CK(clk), .Q(n18925), .QN() );
DFF_X1 gfm_result_reg_29_ ( .D(n5800), .CK(clk), .Q(n18924), .QN() );
DFF_X1 gfm_result_reg_28_ ( .D(n5801), .CK(clk), .Q(n18923), .QN() );
DFF_X1 gfm_result_reg_26_ ( .D(n5803), .CK(clk), .Q(n18921), .QN() );
DFF_X1 gfm_result_reg_25_ ( .D(n5804), .CK(clk), .Q(n18920), .QN() );
DFF_X1 gfm_result_reg_24_ ( .D(n5805), .CK(clk), .Q(n18919), .QN() );
DFF_X1 gfm_result_reg_23_ ( .D(n5806), .CK(clk), .Q(n18918), .QN() );
DFF_X1 gfm_result_reg_21_ ( .D(n5808), .CK(clk), .Q(n18916), .QN() );
DFF_X1 gfm_result_reg_20_ ( .D(n5809), .CK(clk), .Q(n18915), .QN() );
DFF_X1 gfm_result_reg_16_ ( .D(n5813), .CK(clk), .Q(n18911), .QN() );
DFF_X1 gfm_result_reg_34_ ( .D(n5795), .CK(clk), .Q(n18929), .QN() );
DFF_X1 gfm_result_reg_10_ ( .D(n5819), .CK(clk), .Q(n18905), .QN() );
DFF_X1 gfm_result_reg_46_ ( .D(n5783), .CK(clk), .Q(n18941), .QN() );
DFF_X1 gfm_result_reg_110_ ( .D(n5719), .CK(clk), .Q(n19005), .QN() );
DFF_X1 gfm_result_reg_109_ ( .D(n5720), .CK(clk), .Q(n19004), .QN() );
DFF_X1 gfm_result_reg_108_ ( .D(n5721), .CK(clk), .Q(n19003), .QN() );
DFF_X1 gfm_result_reg_107_ ( .D(n5722), .CK(clk), .Q(n19002), .QN() );
DFF_X1 gfm_result_reg_106_ ( .D(n5723), .CK(clk), .Q(n19001), .QN() );
DFF_X1 gfm_result_reg_105_ ( .D(n5724), .CK(clk), .Q(n19000), .QN() );
DFF_X1 gfm_result_reg_104_ ( .D(n5725), .CK(clk), .Q(n18999), .QN() );
DFF_X1 gfm_result_reg_103_ ( .D(n5726), .CK(clk), .Q(n18998), .QN() );
DFF_X1 gfm_result_reg_102_ ( .D(n5727), .CK(clk), .Q(n18997), .QN() );
DFF_X1 gfm_result_reg_101_ ( .D(n5728), .CK(clk), .Q(n18996), .QN() );
DFF_X1 gfm_result_reg_100_ ( .D(n5729), .CK(clk), .Q(n18995), .QN() );
DFF_X1 gfm_result_reg_99_ ( .D(n5730), .CK(clk), .Q(n18994), .QN() );
DFF_X1 gfm_result_reg_98_ ( .D(n5731), .CK(clk), .Q(n18993), .QN() );
DFF_X1 gfm_result_reg_97_ ( .D(n5732), .CK(clk), .Q(n18992), .QN() );
DFF_X1 gfm_result_reg_96_ ( .D(n5733), .CK(clk), .Q(n18991), .QN() );
DFF_X1 gfm_result_reg_95_ ( .D(n5734), .CK(clk), .Q(n18990), .QN() );
DFF_X1 gfm_result_reg_94_ ( .D(n5735), .CK(clk), .Q(n18989), .QN() );
DFF_X1 gfm_result_reg_93_ ( .D(n5736), .CK(clk), .Q(n18988), .QN() );
DFF_X1 gfm_result_reg_92_ ( .D(n5737), .CK(clk), .Q(n18987), .QN() );
DFF_X1 gfm_result_reg_91_ ( .D(n5738), .CK(clk), .Q(n18986), .QN() );
DFF_X1 gfm_result_reg_90_ ( .D(n5739), .CK(clk), .Q(n18985), .QN() );
DFF_X1 gfm_result_reg_89_ ( .D(n5740), .CK(clk), .Q(n18984), .QN() );
DFF_X1 gfm_result_reg_88_ ( .D(n5741), .CK(clk), .Q(n18983), .QN() );
DFF_X1 gfm_result_reg_87_ ( .D(n5742), .CK(clk), .Q(n18982), .QN() );
DFF_X1 gfm_result_reg_86_ ( .D(n5743), .CK(clk), .Q(n18981), .QN() );
DFF_X1 gfm_result_reg_85_ ( .D(n5744), .CK(clk), .Q(n18980), .QN() );
DFF_X1 gfm_result_reg_84_ ( .D(n5745), .CK(clk), .Q(n18979), .QN() );
DFF_X1 gfm_result_reg_83_ ( .D(n5746), .CK(clk), .Q(n18978), .QN() );
DFF_X1 gfm_result_reg_82_ ( .D(n5747), .CK(clk), .Q(n18977), .QN() );
DFF_X1 gfm_result_reg_81_ ( .D(n5748), .CK(clk), .Q(n18976), .QN() );
DFF_X1 gfm_result_reg_80_ ( .D(n5749), .CK(clk), .Q(n18975), .QN() );
DFF_X1 gfm_result_reg_79_ ( .D(n5750), .CK(clk), .Q(n18974), .QN() );
DFF_X1 gfm_result_reg_78_ ( .D(n5751), .CK(clk), .Q(n18973), .QN() );
DFF_X1 gfm_result_reg_77_ ( .D(n5752), .CK(clk), .Q(n18972), .QN() );
DFF_X1 gfm_result_reg_76_ ( .D(n5753), .CK(clk), .Q(n18971), .QN() );
DFF_X1 gfm_result_reg_75_ ( .D(n5754), .CK(clk), .Q(n18970), .QN() );
DFF_X1 gfm_result_reg_74_ ( .D(n5755), .CK(clk), .Q(n18969), .QN() );
DFF_X1 gfm_result_reg_73_ ( .D(n5756), .CK(clk), .Q(n18968), .QN() );
DFF_X1 gfm_result_reg_72_ ( .D(n5757), .CK(clk), .Q(n18967), .QN() );
DFF_X1 gfm_result_reg_71_ ( .D(n5758), .CK(clk), .Q(n18966), .QN() );
DFF_X1 gfm_result_reg_70_ ( .D(n5759), .CK(clk), .Q(n18965), .QN() );
DFF_X1 gfm_result_reg_69_ ( .D(n5760), .CK(clk), .Q(n18964), .QN() );
DFF_X1 gfm_result_reg_68_ ( .D(n5761), .CK(clk), .Q(n18963), .QN() );
DFF_X1 gfm_result_reg_67_ ( .D(n5762), .CK(clk), .Q(n18962), .QN() );
DFF_X1 gfm_result_reg_66_ ( .D(n5763), .CK(clk), .Q(n18961), .QN() );
DFF_X1 gfm_result_reg_65_ ( .D(n5764), .CK(clk), .Q(n18960), .QN() );
DFF_X1 gfm_result_reg_64_ ( .D(n5765), .CK(clk), .Q(n18959), .QN() );
DFF_X1 gfm_result_reg_63_ ( .D(n5766), .CK(clk), .Q(n18958), .QN() );
DFF_X1 gfm_result_reg_62_ ( .D(n5767), .CK(clk), .Q(n18957), .QN() );
DFF_X1 gfm_result_reg_61_ ( .D(n5768), .CK(clk), .Q(n18956), .QN() );
DFF_X1 gfm_result_reg_60_ ( .D(n5769), .CK(clk), .Q(n18955), .QN() );
DFF_X1 gfm_result_reg_59_ ( .D(n5770), .CK(clk), .Q(n18954), .QN() );
DFF_X1 gfm_result_reg_58_ ( .D(n5771), .CK(clk), .Q(n18953), .QN() );
DFF_X1 gfm_result_reg_57_ ( .D(n5772), .CK(clk), .Q(n18952), .QN() );
DFF_X1 gfm_result_reg_56_ ( .D(n5773), .CK(clk), .Q(n18951), .QN() );
DFF_X1 gfm_result_reg_55_ ( .D(n5774), .CK(clk), .Q(n18950), .QN() );
DFF_X1 gfm_result_reg_54_ ( .D(n5775), .CK(clk), .Q(n18949), .QN() );
DFF_X1 gfm_result_reg_53_ ( .D(n5776), .CK(clk), .Q(n18948), .QN() );
DFF_X1 gfm_result_reg_52_ ( .D(n5777), .CK(clk), .Q(n18947), .QN() );
DFF_X1 gfm_result_reg_51_ ( .D(n5778), .CK(clk), .Q(n18946), .QN() );
DFF_X1 gfm_result_reg_50_ ( .D(n5779), .CK(clk), .Q(n18945), .QN() );
DFF_X1 gfm_result_reg_49_ ( .D(n5780), .CK(clk), .Q(n18944), .QN() );
DFF_X1 gfm_result_reg_48_ ( .D(n5781), .CK(clk), .Q(n18943), .QN() );
DFF_X1 gfm_result_reg_47_ ( .D(n5782), .CK(clk), .Q(n18942), .QN() );
DFF_X1 gfm_result_reg_27_ ( .D(n5802), .CK(clk), .Q(n18922), .QN() );
DFF_X1 gfm_result_reg_22_ ( .D(n5807), .CK(clk), .Q(n18917), .QN() );
DFF_X1 gfm_result_reg_19_ ( .D(n5810), .CK(clk), .Q(n18914), .QN() );
DFF_X1 gfm_result_reg_18_ ( .D(n5811), .CK(clk), .Q(n18913), .QN() );
DFF_X1 gfm_result_reg_17_ ( .D(n5812), .CK(clk), .Q(n18912), .QN() );
DFF_X1 gfm_result_reg_15_ ( .D(n5814), .CK(clk), .Q(n18910), .QN() );
DFF_X1 gfm_result_reg_11_ ( .D(n5818), .CK(clk), .Q(n18906), .QN() );
DFF_X1 gfm_result_reg_31_ ( .D(n5798), .CK(clk), .Q(n18926), .QN() );
DFF_X1 gfm_result_reg_32_ ( .D(n5797), .CK(clk), .Q(n18927), .QN() );
DFF_X1 gfm_result_reg_12_ ( .D(n5817), .CK(clk), .Q(n18907), .QN() );
DFF_X1 gfm_result_reg_127_ ( .D(n5702), .CK(clk), .Q(n19022), .QN(n17024) );
DFF_X1 gfm_result_reg_124_ ( .D(n5705), .CK(clk), .Q(n19019), .QN(n17030) );
DFF_X1 gfm_result_reg_121_ ( .D(n5708), .CK(clk), .Q(n19016), .QN(n17036) );
DFF_X1 gfm_result_reg_123_ ( .D(n5706), .CK(clk), .Q(n19018), .QN(n17032) );
DFF_X1 gfm_result_reg_122_ ( .D(n5707), .CK(clk), .Q(n19017), .QN(n17034) );
DFF_X1 gfm_result_reg_111_ ( .D(n5718), .CK(clk), .Q(n19006), .QN() );
DFF_X1 gfm_result_reg_126_ ( .D(n5703), .CK(clk), .Q(n19021), .QN(n17026) );
DFF_X1 gfm_result_reg_125_ ( .D(n5704), .CK(clk), .Q(n19020), .QN(n17028) );
DFF_X1 gfm_result_reg_120_ ( .D(n5709), .CK(clk), .Q(n19015), .QN(n17038) );
DFF_X1 gfm_result_reg_116_ ( .D(n5713), .CK(clk), .Q(n19011), .QN() );
DFF_X1 gfm_result_reg_115_ ( .D(n5714), .CK(clk), .Q(n19010), .QN() );
DFF_X1 gfm_result_reg_117_ ( .D(n5712), .CK(clk), .Q(n19012), .QN() );
DFF_X1 gfm_result_reg_112_ ( .D(n5717), .CK(clk), .Q(n19007), .QN() );
DFF_X1 gfm_result_reg_119_ ( .D(n5710), .CK(clk), .Q(n19014), .QN() );
DFF_X1 gfm_result_reg_114_ ( .D(n5715), .CK(clk), .Q(n19009), .QN() );
DFF_X1 gfm_result_reg_118_ ( .D(n5711), .CK(clk), .Q(n19013), .QN() );
DFF_X1 gfm_result_reg_113_ ( .D(n5716), .CK(clk), .Q(n19008), .QN() );
DFF_X1 gfm_cnt_reg_0_ ( .D(n17280), .CK(clk), .Q(n18622), .QN(n6859) );
DFF_X1 gfm_cnt_reg_1_ ( .D(n6291), .CK(clk), .Q(n18624), .QN(n6850) );
DFF_X1 gfm_cnt_reg_2_ ( .D(n6290), .CK(clk), .Q(n18893), .QN(n16838) );
OR3_X4 U13738 ( .A1(n17281), .A2(n17837), .A3(n17996), .ZN(n17282) );
NOR4_X2 U13739 ( .A1(n18079), .A2(n16837), .A3(state[7]), .A4(state[9]),.ZN(n17283) );
OR2_X4 U13740 ( .A1(n11946), .A2(n16542), .ZN(n17284) );
OR2_X4 U13741 ( .A1(n17281), .A2(n17841), .ZN(n17285) );
OR2_X4 U13742 ( .A1(cii_ctl_vld), .A2(n17958), .ZN(n17286) );
NAND3_X2 U13743 ( .A1(dii_data_vld), .A2(n18617), .A3(n18081), .ZN(n18085));
OR2_X4 U13744 ( .A1(n19204), .A2(dii_data_size[0]), .ZN(n17287) );
NOR2_X2 U13745 ( .A1(n19203), .A2(n18744), .ZN(n17288) );
OR2_X4 U13746 ( .A1(n18892), .A2(cii_ctl_vld), .ZN(n17289) );
AND2_X4 U13747 ( .A1(n12235), .A2(state[3]), .ZN(n17290) );
AND2_X4 U13748 ( .A1(n18623), .A2(n18622), .ZN(n17291) );
AND2_X4 U13749 ( .A1(n18619), .A2(n18618), .ZN(n17375) );
BUF_X32 U13750 ( .A(cii_K[64]), .Z(n17376) );
BUF_X32 U13751 ( .A(cii_K[32]), .Z(n17377) );
BUF_X32 U13752 ( .A(cii_K[79]), .Z(n17378) );
BUF_X32 U13753 ( .A(cii_K[47]), .Z(n17379) );
BUF_X32 U13754 ( .A(cii_K[87]), .Z(n17380) );
BUF_X32 U13755 ( .A(cii_K[55]), .Z(n17381) );
BUF_X32 U13756 ( .A(cii_K[95]), .Z(n17382) );
BUF_X32 U13757 ( .A(cii_K[63]), .Z(n17383) );
BUF_X32 U13758 ( .A(cii_K[71]), .Z(n17384) );
BUF_X32 U13759 ( .A(cii_K[39]), .Z(n17385) );
BUF_X32 U13760 ( .A(cii_K[7]), .Z(n17386) );
BUF_X32 U13761 ( .A(cii_K[103]), .Z(n17387) );
BUF_X32 U13762 ( .A(cii_K[70]), .Z(n17388) );
BUF_X32 U13763 ( .A(cii_K[38]), .Z(n17389) );
BUF_X32 U13764 ( .A(cii_K[6]), .Z(n17390) );
BUF_X32 U13765 ( .A(cii_K[102]), .Z(n17391) );
BUF_X32 U13766 ( .A(cii_K[69]), .Z(n17392) );
BUF_X32 U13767 ( .A(cii_K[37]), .Z(n17393) );
BUF_X32 U13768 ( .A(cii_K[5]), .Z(n17394) );
BUF_X32 U13769 ( .A(cii_K[101]), .Z(n17395) );
BUF_X32 U13770 ( .A(cii_K[68]), .Z(n17396) );
BUF_X32 U13771 ( .A(cii_K[36]), .Z(n17397) );
BUF_X32 U13772 ( .A(cii_K[4]), .Z(n17398) );
BUF_X32 U13773 ( .A(cii_K[100]), .Z(n17399) );
BUF_X32 U13774 ( .A(cii_K[67]), .Z(n17400) );
BUF_X32 U13775 ( .A(cii_K[35]), .Z(n17401) );
BUF_X32 U13776 ( .A(cii_K[3]), .Z(n17402) );
BUF_X32 U13777 ( .A(cii_K[99]), .Z(n17403) );
BUF_X32 U13778 ( .A(cii_K[66]), .Z(n17404) );
BUF_X32 U13779 ( .A(cii_K[34]), .Z(n17405) );
BUF_X32 U13780 ( .A(cii_K[2]), .Z(n17406) );
BUF_X32 U13781 ( .A(cii_K[98]), .Z(n17407) );
BUF_X32 U13782 ( .A(cii_K[65]), .Z(n17408) );
BUF_X32 U13783 ( .A(cii_K[33]), .Z(n17409) );
BUF_X32 U13784 ( .A(cii_K[1]), .Z(n17410) );
BUF_X32 U13785 ( .A(cii_K[97]), .Z(n17411) );
BUF_X32 U13786 ( .A(cii_K[31]), .Z(n17412) );
BUF_X32 U13787 ( .A(cii_K[126]), .Z(n17413) );
BUF_X32 U13788 ( .A(cii_K[94]), .Z(n17414) );
BUF_X32 U13789 ( .A(cii_K[62]), .Z(n17415) );
BUF_X32 U13790 ( .A(cii_K[30]), .Z(n17416) );
BUF_X32 U13791 ( .A(cii_K[125]), .Z(n17417) );
BUF_X32 U13792 ( .A(cii_K[93]), .Z(n17418) );
BUF_X32 U13793 ( .A(cii_K[61]), .Z(n17419) );
BUF_X32 U13794 ( .A(cii_K[29]), .Z(n17420) );
BUF_X32 U13795 ( .A(cii_K[124]), .Z(n17421) );
BUF_X32 U13796 ( .A(cii_K[92]), .Z(n17422) );
BUF_X32 U13797 ( .A(cii_K[60]), .Z(n17423) );
BUF_X32 U13798 ( .A(cii_K[28]), .Z(n17424) );
BUF_X32 U13799 ( .A(cii_K[123]), .Z(n17425) );
BUF_X32 U13800 ( .A(cii_K[91]), .Z(n17426) );
BUF_X32 U13801 ( .A(cii_K[59]), .Z(n17427) );
BUF_X32 U13802 ( .A(cii_K[27]), .Z(n17428) );
BUF_X32 U13803 ( .A(cii_K[122]), .Z(n17429) );
BUF_X32 U13804 ( .A(cii_K[90]), .Z(n17430) );
BUF_X32 U13805 ( .A(cii_K[58]), .Z(n17431) );
BUF_X32 U13806 ( .A(cii_K[26]), .Z(n17432) );
BUF_X32 U13807 ( .A(cii_K[121]), .Z(n17433) );
BUF_X32 U13808 ( .A(cii_K[89]), .Z(n17434) );
BUF_X32 U13809 ( .A(cii_K[57]), .Z(n17435) );
BUF_X32 U13810 ( .A(cii_K[25]), .Z(n17436) );
BUF_X32 U13811 ( .A(cii_K[120]), .Z(n17437) );
BUF_X32 U13812 ( .A(cii_K[88]), .Z(n17438) );
BUF_X32 U13813 ( .A(cii_K[56]), .Z(n17439) );
BUF_X32 U13814 ( .A(cii_K[24]), .Z(n17440) );
BUF_X32 U13815 ( .A(cii_K[23]), .Z(n17441) );
BUF_X32 U13816 ( .A(cii_K[119]), .Z(n17442) );
BUF_X32 U13817 ( .A(cii_K[86]), .Z(n17443) );
BUF_X32 U13818 ( .A(cii_K[54]), .Z(n17444) );
BUF_X32 U13819 ( .A(cii_K[22]), .Z(n17445) );
BUF_X32 U13820 ( .A(cii_K[118]), .Z(n17446) );
BUF_X32 U13821 ( .A(cii_K[85]), .Z(n17447) );
BUF_X32 U13822 ( .A(cii_K[53]), .Z(n17448) );
BUF_X32 U13823 ( .A(cii_K[21]), .Z(n17449) );
BUF_X32 U13824 ( .A(cii_K[117]), .Z(n17450) );
BUF_X32 U13825 ( .A(cii_K[84]), .Z(n17451) );
BUF_X32 U13826 ( .A(cii_K[52]), .Z(n17452) );
BUF_X32 U13827 ( .A(cii_K[20]), .Z(n17453) );
BUF_X32 U13828 ( .A(cii_K[116]), .Z(n17454) );
BUF_X32 U13829 ( .A(cii_K[83]), .Z(n17455) );
BUF_X32 U13830 ( .A(cii_K[51]), .Z(n17456) );
BUF_X32 U13831 ( .A(cii_K[19]), .Z(n17457) );
BUF_X32 U13832 ( .A(cii_K[115]), .Z(n17458) );
BUF_X32 U13833 ( .A(cii_K[82]), .Z(n17459) );
BUF_X32 U13834 ( .A(cii_K[50]), .Z(n17460) );
BUF_X32 U13835 ( .A(cii_K[18]), .Z(n17461) );
BUF_X32 U13836 ( .A(cii_K[114]), .Z(n17462) );
BUF_X32 U13837 ( .A(cii_K[81]), .Z(n17463) );
BUF_X32 U13838 ( .A(cii_K[49]), .Z(n17464) );
BUF_X32 U13839 ( .A(cii_K[17]), .Z(n17465) );
BUF_X32 U13840 ( .A(cii_K[113]), .Z(n17466) );
BUF_X32 U13841 ( .A(cii_K[80]), .Z(n17467) );
BUF_X32 U13842 ( .A(cii_K[48]), .Z(n17468) );
BUF_X32 U13843 ( .A(cii_K[16]), .Z(n17469) );
BUF_X32 U13844 ( .A(cii_K[112]), .Z(n17470) );
BUF_X32 U13845 ( .A(cii_K[15]), .Z(n17471) );
BUF_X32 U13846 ( .A(cii_K[111]), .Z(n17472) );
BUF_X32 U13847 ( .A(cii_K[78]), .Z(n17473) );
BUF_X32 U13848 ( .A(cii_K[46]), .Z(n17474) );
BUF_X32 U13849 ( .A(cii_K[14]), .Z(n17475) );
BUF_X32 U13850 ( .A(cii_K[110]), .Z(n17476) );
BUF_X32 U13851 ( .A(cii_K[77]), .Z(n17477) );
BUF_X32 U13852 ( .A(cii_K[45]), .Z(n17478) );
BUF_X32 U13853 ( .A(cii_K[13]), .Z(n17479) );
BUF_X32 U13854 ( .A(cii_K[109]), .Z(n17480) );
BUF_X32 U13855 ( .A(cii_K[76]), .Z(n17481) );
BUF_X32 U13856 ( .A(cii_K[44]), .Z(n17482) );
BUF_X32 U13857 ( .A(cii_K[12]), .Z(n17483) );
BUF_X32 U13858 ( .A(cii_K[108]), .Z(n17484) );
BUF_X32 U13859 ( .A(cii_K[75]), .Z(n17485) );
BUF_X32 U13860 ( .A(cii_K[43]), .Z(n17486) );
BUF_X32 U13861 ( .A(cii_K[11]), .Z(n17487) );
BUF_X32 U13862 ( .A(cii_K[107]), .Z(n17488) );
BUF_X32 U13863 ( .A(cii_K[74]), .Z(n17489) );
BUF_X32 U13864 ( .A(cii_K[42]), .Z(n17490) );
BUF_X32 U13865 ( .A(cii_K[10]), .Z(n17491) );
BUF_X32 U13866 ( .A(cii_K[106]), .Z(n17492) );
BUF_X32 U13867 ( .A(cii_K[73]), .Z(n17493) );
BUF_X32 U13868 ( .A(cii_K[41]), .Z(n17494) );
BUF_X32 U13869 ( .A(cii_K[9]), .Z(n17495) );
BUF_X32 U13870 ( .A(cii_K[105]), .Z(n17496) );
BUF_X32 U13871 ( .A(cii_K[72]), .Z(n17497) );
BUF_X32 U13872 ( .A(cii_K[40]), .Z(n17498) );
BUF_X32 U13873 ( .A(cii_K[8]), .Z(n17499) );
BUF_X32 U13874 ( .A(cii_K[104]), .Z(n17500) );
BUF_X32 U13875 ( .A(cii_K[0]), .Z(n17501) );
BUF_X32 U13876 ( .A(cii_K[96]), .Z(n17502) );
NAND2_X1 U13877 ( .A1(n17930), .A2(n13675), .ZN(n13671) );
XOR2_X1 U13878 ( .A(aes_text_out[65]), .B(n17629), .Z(n13668) );
NAND2_X1 U13879 ( .A1(n17924), .A2(n13661), .ZN(n13656) );
BUF_X32 U13880 ( .A(n6025), .Z(n17503) );
NAND2_X1 U13881 ( .A1(n12495), .A2(n12496), .ZN(n6025) );
NAND2_X1 U13882 ( .A1(dii_data_size[1]), .A2(n17281), .ZN(n12496) );
BUF_X32 U13883 ( .A(n6024), .Z(n17504) );
NAND2_X1 U13884 ( .A1(n12497), .A2(n12498), .ZN(n6024) );
NAND2_X1 U13885 ( .A1(dii_data_size[2]), .A2(n17281), .ZN(n12498) );
NOR3_X1 U13886 ( .A1(n18746), .A2(n11976), .A3(n18601), .ZN(n17281) );
CLKBUF_X2 U13887 ( .A(n17281), .Z(n17505) );
NAND3_X1 U13888 ( .A1(n18596), .A2(n17506), .A3(n18594), .ZN(n5830) );
BUF_X8 U13889 ( .A(n18595), .Z(n17506) );
CLKBUF_X2 U13890 ( .A(n5830), .Z(n17507) );
NAND2_X1 U13891 ( .A1(dii_data[127]), .A2(n17799), .ZN(n18595) );
NAND3_X1 U13892 ( .A1(n18088), .A2(n17508), .A3(n18086), .ZN(n5831) );
BUF_X8 U13893 ( .A(n18087), .Z(n17508) );
CLKBUF_X2 U13894 ( .A(n5831), .Z(n17509) );
NAND2_X1 U13895 ( .A1(dii_data[126]), .A2(n17788), .ZN(n18087) );
NAND3_X1 U13896 ( .A1(n18092), .A2(n17510), .A3(n18090), .ZN(n5832) );
BUF_X8 U13897 ( .A(n18091), .Z(n17510) );
CLKBUF_X2 U13898 ( .A(n5832), .Z(n17511) );
NAND2_X1 U13899 ( .A1(dii_data[125]), .A2(n17788), .ZN(n18091) );
NAND3_X1 U13900 ( .A1(n18096), .A2(n17512), .A3(n18094), .ZN(n5833) );
BUF_X8 U13901 ( .A(n18095), .Z(n17512) );
CLKBUF_X2 U13902 ( .A(n5833), .Z(n17513) );
NAND2_X1 U13903 ( .A1(dii_data[124]), .A2(n17788), .ZN(n18095) );
NAND3_X1 U13904 ( .A1(n18100), .A2(n17514), .A3(n18098), .ZN(n5834) );
BUF_X8 U13905 ( .A(n18099), .Z(n17514) );
CLKBUF_X2 U13906 ( .A(n5834), .Z(n17515) );
NAND2_X1 U13907 ( .A1(dii_data[123]), .A2(n17788), .ZN(n18099) );
NAND3_X1 U13908 ( .A1(n18104), .A2(n17516), .A3(n18102), .ZN(n5835) );
BUF_X8 U13909 ( .A(n18103), .Z(n17516) );
CLKBUF_X2 U13910 ( .A(n5835), .Z(n17517) );
NAND2_X1 U13911 ( .A1(dii_data[122]), .A2(n17788), .ZN(n18103) );
NAND3_X1 U13912 ( .A1(n18108), .A2(n17518), .A3(n18106), .ZN(n5836) );
BUF_X8 U13913 ( .A(n18107), .Z(n17518) );
CLKBUF_X2 U13914 ( .A(n5836), .Z(n17519) );
NAND2_X1 U13915 ( .A1(dii_data[121]), .A2(n17788), .ZN(n18107) );
NAND3_X1 U13916 ( .A1(n18112), .A2(n17520), .A3(n18110), .ZN(n5837) );
BUF_X8 U13917 ( .A(n18111), .Z(n17520) );
CLKBUF_X2 U13918 ( .A(n5837), .Z(n17521) );
NAND2_X1 U13919 ( .A1(dii_data[120]), .A2(n17788), .ZN(n18111) );
CLKBUF_X1 U13920 ( .A(dii_data[119]), .Z(n17523) );
CLKBUF_X2 U13921 ( .A(n17523), .Z(n17522) );
NAND2_X1 U13922 ( .A1(n17522), .A2(n17788), .ZN(n18115) );
CLKBUF_X1 U13923 ( .A(dii_data[118]), .Z(n17525) );
CLKBUF_X2 U13924 ( .A(n17525), .Z(n17524) );
NAND2_X1 U13925 ( .A1(n17524), .A2(n17788), .ZN(n18119) );
CLKBUF_X1 U13926 ( .A(dii_data[117]), .Z(n17527) );
CLKBUF_X2 U13927 ( .A(n17527), .Z(n17526) );
NAND2_X1 U13928 ( .A1(n17526), .A2(n17788), .ZN(n18123) );
CLKBUF_X1 U13929 ( .A(dii_data[116]), .Z(n17529) );
CLKBUF_X2 U13930 ( .A(n17529), .Z(n17528) );
NAND2_X1 U13931 ( .A1(n17528), .A2(n17788), .ZN(n18127) );
CLKBUF_X1 U13932 ( .A(dii_data[115]), .Z(n17531) );
CLKBUF_X2 U13933 ( .A(n17531), .Z(n17530) );
NAND2_X1 U13934 ( .A1(n17530), .A2(n17789), .ZN(n18131) );
CLKBUF_X1 U13935 ( .A(dii_data[114]), .Z(n17533) );
CLKBUF_X2 U13936 ( .A(n17533), .Z(n17532) );
NAND2_X1 U13937 ( .A1(n17532), .A2(n17789), .ZN(n18135) );
CLKBUF_X1 U13938 ( .A(dii_data[113]), .Z(n17535) );
CLKBUF_X2 U13939 ( .A(n17535), .Z(n17534) );
NAND2_X1 U13940 ( .A1(n17534), .A2(n17789), .ZN(n18139) );
CLKBUF_X1 U13941 ( .A(dii_data[112]), .Z(n17537) );
CLKBUF_X2 U13942 ( .A(n17537), .Z(n17536) );
NAND2_X1 U13943 ( .A1(n17536), .A2(n17789), .ZN(n18143) );
NAND3_X1 U13944 ( .A1(n18148), .A2(n18147), .A3(n18146), .ZN(n5846) );
CLKBUF_X2 U13945 ( .A(n5846), .Z(n17538) );
CLKBUF_X2 U13946 ( .A(dii_data[111]), .Z(n17539) );
NAND2_X1 U13947 ( .A1(n17539), .A2(n17789), .ZN(n18147) );
NAND3_X1 U13948 ( .A1(n18152), .A2(n18151), .A3(n18150), .ZN(n5847) );
CLKBUF_X2 U13949 ( .A(n5847), .Z(n17540) );
CLKBUF_X2 U13950 ( .A(dii_data[110]), .Z(n17541) );
NAND2_X1 U13951 ( .A1(n17541), .A2(n17789), .ZN(n18151) );
NAND3_X1 U13952 ( .A1(n18156), .A2(n18155), .A3(n18154), .ZN(n5848) );
CLKBUF_X2 U13953 ( .A(n5848), .Z(n17542) );
CLKBUF_X2 U13954 ( .A(dii_data[109]), .Z(n17543) );
NAND2_X1 U13955 ( .A1(n17543), .A2(n17789), .ZN(n18155) );
NAND3_X1 U13956 ( .A1(n18160), .A2(n18159), .A3(n18158), .ZN(n5849) );
CLKBUF_X2 U13957 ( .A(n5849), .Z(n17544) );
CLKBUF_X2 U13958 ( .A(dii_data[108]), .Z(n17545) );
NAND2_X1 U13959 ( .A1(n17545), .A2(n17789), .ZN(n18159) );
NAND3_X1 U13960 ( .A1(n18164), .A2(n18163), .A3(n18162), .ZN(n5850) );
CLKBUF_X2 U13961 ( .A(n5850), .Z(n17546) );
CLKBUF_X2 U13962 ( .A(dii_data[107]), .Z(n17547) );
NAND2_X1 U13963 ( .A1(n17547), .A2(n17789), .ZN(n18163) );
NAND3_X1 U13964 ( .A1(n18168), .A2(n18167), .A3(n18166), .ZN(n5851) );
CLKBUF_X2 U13965 ( .A(n5851), .Z(n17548) );
CLKBUF_X2 U13966 ( .A(dii_data[106]), .Z(n17549) );
NAND2_X1 U13967 ( .A1(n17549), .A2(n17789), .ZN(n18167) );
NAND3_X1 U13968 ( .A1(n18172), .A2(n18171), .A3(n18170), .ZN(n5852) );
CLKBUF_X2 U13969 ( .A(n5852), .Z(n17550) );
CLKBUF_X2 U13970 ( .A(dii_data[105]), .Z(n17551) );
NAND2_X1 U13971 ( .A1(n17551), .A2(n17789), .ZN(n18171) );
NAND3_X1 U13972 ( .A1(n18176), .A2(n18175), .A3(n18174), .ZN(n5853) );
CLKBUF_X2 U13973 ( .A(n5853), .Z(n17552) );
CLKBUF_X2 U13974 ( .A(dii_data[104]), .Z(n17553) );
NAND2_X1 U13975 ( .A1(n17553), .A2(n17790), .ZN(n18175) );
NAND3_X1 U13976 ( .A1(n18180), .A2(n18179), .A3(n18178), .ZN(n5854) );
CLKBUF_X2 U13977 ( .A(n5854), .Z(n17554) );
CLKBUF_X2 U13978 ( .A(dii_data[103]), .Z(n17555) );
NAND2_X1 U13979 ( .A1(n17555), .A2(n17790), .ZN(n18179) );
NAND3_X1 U13980 ( .A1(n18184), .A2(n18183), .A3(n18182), .ZN(n5855) );
CLKBUF_X2 U13981 ( .A(n5855), .Z(n17556) );
CLKBUF_X2 U13982 ( .A(dii_data[102]), .Z(n17557) );
NAND2_X1 U13983 ( .A1(n17557), .A2(n17790), .ZN(n18183) );
NAND3_X1 U13984 ( .A1(n18188), .A2(n18187), .A3(n18186), .ZN(n5856) );
CLKBUF_X2 U13985 ( .A(n5856), .Z(n17558) );
CLKBUF_X2 U13986 ( .A(dii_data[101]), .Z(n17559) );
NAND2_X1 U13987 ( .A1(n17559), .A2(n17790), .ZN(n18187) );
NAND3_X1 U13988 ( .A1(n18192), .A2(n18191), .A3(n18190), .ZN(n5857) );
CLKBUF_X2 U13989 ( .A(n5857), .Z(n17560) );
CLKBUF_X2 U13990 ( .A(dii_data[100]), .Z(n17561) );
NAND2_X1 U13991 ( .A1(n17561), .A2(n17790), .ZN(n18191) );
NAND3_X1 U13992 ( .A1(n18196), .A2(n18195), .A3(n18194), .ZN(n5858) );
CLKBUF_X2 U13993 ( .A(n5858), .Z(n17562) );
CLKBUF_X2 U13994 ( .A(dii_data[99]), .Z(n17563) );
NAND2_X1 U13995 ( .A1(n17563), .A2(n17790), .ZN(n18195) );
NAND3_X1 U13996 ( .A1(n18204), .A2(n18203), .A3(n18202), .ZN(n5859) );
CLKBUF_X2 U13997 ( .A(n5859), .Z(n17564) );
CLKBUF_X2 U13998 ( .A(dii_data[97]), .Z(n17565) );
NAND2_X1 U13999 ( .A1(n17565), .A2(n17790), .ZN(n18203) );
NAND3_X1 U14000 ( .A1(n18208), .A2(n18207), .A3(n18206), .ZN(n5860) );
CLKBUF_X2 U14001 ( .A(n5860), .Z(n17566) );
CLKBUF_X2 U14002 ( .A(dii_data[96]), .Z(n17567) );
NAND2_X1 U14003 ( .A1(n17567), .A2(n17790), .ZN(n18207) );
NAND3_X1 U14004 ( .A1(n18212), .A2(n18211), .A3(n18210), .ZN(n5861) );
CLKBUF_X2 U14005 ( .A(n5861), .Z(n17568) );
CLKBUF_X2 U14006 ( .A(dii_data[95]), .Z(n17569) );
NAND2_X1 U14007 ( .A1(n17569), .A2(n17790), .ZN(n18211) );
NAND3_X1 U14008 ( .A1(n18216), .A2(n18215), .A3(n18214), .ZN(n5862) );
CLKBUF_X2 U14009 ( .A(n5862), .Z(n17570) );
CLKBUF_X2 U14010 ( .A(dii_data[94]), .Z(n17571) );
NAND2_X1 U14011 ( .A1(n17571), .A2(n17790), .ZN(n18215) );
NAND3_X1 U14012 ( .A1(n18220), .A2(n18219), .A3(n18218), .ZN(n5863) );
CLKBUF_X2 U14013 ( .A(n5863), .Z(n17572) );
CLKBUF_X2 U14014 ( .A(dii_data[93]), .Z(n17573) );
NAND2_X1 U14015 ( .A1(n17573), .A2(n17791), .ZN(n18219) );
NAND3_X1 U14016 ( .A1(n18224), .A2(n18223), .A3(n18222), .ZN(n5864) );
CLKBUF_X2 U14017 ( .A(n5864), .Z(n17574) );
CLKBUF_X2 U14018 ( .A(dii_data[92]), .Z(n17575) );
NAND2_X1 U14019 ( .A1(n17575), .A2(n17791), .ZN(n18223) );
NAND3_X1 U14020 ( .A1(n18228), .A2(n18227), .A3(n18226), .ZN(n5865) );
CLKBUF_X2 U14021 ( .A(n5865), .Z(n17576) );
CLKBUF_X2 U14022 ( .A(dii_data[91]), .Z(n17577) );
NAND2_X1 U14023 ( .A1(n17577), .A2(n17791), .ZN(n18227) );
NAND3_X1 U14024 ( .A1(n18232), .A2(n18231), .A3(n18230), .ZN(n5866) );
CLKBUF_X2 U14025 ( .A(n5866), .Z(n17578) );
CLKBUF_X2 U14026 ( .A(dii_data[90]), .Z(n17579) );
NAND2_X1 U14027 ( .A1(n17579), .A2(n17791), .ZN(n18231) );
NAND3_X1 U14028 ( .A1(n18236), .A2(n18235), .A3(n18234), .ZN(n5867) );
CLKBUF_X2 U14029 ( .A(n5867), .Z(n17580) );
CLKBUF_X2 U14030 ( .A(dii_data[89]), .Z(n17581) );
NAND2_X1 U14031 ( .A1(n17581), .A2(n17791), .ZN(n18235) );
NAND3_X1 U14032 ( .A1(n18240), .A2(n18239), .A3(n18238), .ZN(n5868) );
CLKBUF_X2 U14033 ( .A(n5868), .Z(n17582) );
CLKBUF_X2 U14034 ( .A(dii_data[88]), .Z(n17583) );
NAND2_X1 U14035 ( .A1(n17583), .A2(n17791), .ZN(n18239) );
NAND3_X1 U14036 ( .A1(n18244), .A2(n18243), .A3(n18242), .ZN(n5869) );
CLKBUF_X2 U14037 ( .A(n5869), .Z(n17584) );
CLKBUF_X2 U14038 ( .A(dii_data[87]), .Z(n17585) );
NAND2_X1 U14039 ( .A1(n17585), .A2(n17791), .ZN(n18243) );
NAND3_X1 U14040 ( .A1(n18248), .A2(n18247), .A3(n18246), .ZN(n5870) );
CLKBUF_X2 U14041 ( .A(n5870), .Z(n17586) );
CLKBUF_X2 U14042 ( .A(dii_data[86]), .Z(n17587) );
NAND2_X1 U14043 ( .A1(n17587), .A2(n17791), .ZN(n18247) );
NAND3_X1 U14044 ( .A1(n18252), .A2(n18251), .A3(n18250), .ZN(n5871) );
CLKBUF_X2 U14045 ( .A(n5871), .Z(n17588) );
CLKBUF_X2 U14046 ( .A(dii_data[85]), .Z(n17589) );
NAND2_X1 U14047 ( .A1(n17589), .A2(n17791), .ZN(n18251) );
NAND3_X1 U14048 ( .A1(n18256), .A2(n18255), .A3(n18254), .ZN(n5872) );
CLKBUF_X2 U14049 ( .A(n5872), .Z(n17590) );
CLKBUF_X2 U14050 ( .A(dii_data[84]), .Z(n17591) );
NAND2_X1 U14051 ( .A1(n17591), .A2(n17791), .ZN(n18255) );
NAND3_X1 U14052 ( .A1(n18260), .A2(n18259), .A3(n18258), .ZN(n5873) );
CLKBUF_X2 U14053 ( .A(n5873), .Z(n17592) );
CLKBUF_X2 U14054 ( .A(dii_data[83]), .Z(n17593) );
NAND2_X1 U14055 ( .A1(n17593), .A2(n17791), .ZN(n18259) );
NAND3_X1 U14056 ( .A1(n18264), .A2(n18263), .A3(n18262), .ZN(n5874) );
CLKBUF_X2 U14057 ( .A(n5874), .Z(n17594) );
CLKBUF_X2 U14058 ( .A(dii_data[82]), .Z(n17595) );
NAND2_X1 U14059 ( .A1(n17595), .A2(n17792), .ZN(n18263) );
NAND3_X1 U14060 ( .A1(n18268), .A2(n18267), .A3(n18266), .ZN(n5875) );
CLKBUF_X2 U14061 ( .A(n5875), .Z(n17596) );
CLKBUF_X2 U14062 ( .A(dii_data[81]), .Z(n17597) );
NAND2_X1 U14063 ( .A1(n17597), .A2(n17792), .ZN(n18267) );
NAND3_X1 U14064 ( .A1(n18272), .A2(n18271), .A3(n18270), .ZN(n5876) );
CLKBUF_X2 U14065 ( .A(n5876), .Z(n17598) );
CLKBUF_X2 U14066 ( .A(dii_data[80]), .Z(n17599) );
NAND2_X1 U14067 ( .A1(n17599), .A2(n17792), .ZN(n18271) );
NAND3_X1 U14068 ( .A1(n18276), .A2(n18275), .A3(n18274), .ZN(n5877) );
CLKBUF_X2 U14069 ( .A(n5877), .Z(n17600) );
CLKBUF_X2 U14070 ( .A(dii_data[79]), .Z(n17601) );
NAND2_X1 U14071 ( .A1(n17601), .A2(n17792), .ZN(n18275) );
NAND3_X1 U14072 ( .A1(n18280), .A2(n18279), .A3(n18278), .ZN(n5878) );
CLKBUF_X2 U14073 ( .A(n5878), .Z(n17602) );
CLKBUF_X2 U14074 ( .A(dii_data[78]), .Z(n17603) );
NAND2_X1 U14075 ( .A1(n17603), .A2(n17792), .ZN(n18279) );
NAND3_X1 U14076 ( .A1(n18284), .A2(n18283), .A3(n18282), .ZN(n5879) );
CLKBUF_X2 U14077 ( .A(n5879), .Z(n17604) );
CLKBUF_X2 U14078 ( .A(dii_data[77]), .Z(n17605) );
NAND2_X1 U14079 ( .A1(n17605), .A2(n17792), .ZN(n18283) );
NAND3_X1 U14080 ( .A1(n18288), .A2(n18287), .A3(n18286), .ZN(n5880) );
CLKBUF_X2 U14081 ( .A(n5880), .Z(n17606) );
CLKBUF_X2 U14082 ( .A(dii_data[76]), .Z(n17607) );
NAND2_X1 U14083 ( .A1(n17607), .A2(n17792), .ZN(n18287) );
NAND3_X1 U14084 ( .A1(n18292), .A2(n18291), .A3(n18290), .ZN(n5881) );
CLKBUF_X2 U14085 ( .A(n5881), .Z(n17608) );
CLKBUF_X2 U14086 ( .A(dii_data[75]), .Z(n17609) );
NAND2_X1 U14087 ( .A1(n17609), .A2(n17792), .ZN(n18291) );
NAND3_X1 U14088 ( .A1(n18296), .A2(n18295), .A3(n18294), .ZN(n5882) );
CLKBUF_X2 U14089 ( .A(n5882), .Z(n17610) );
CLKBUF_X2 U14090 ( .A(dii_data[74]), .Z(n17611) );
NAND2_X1 U14091 ( .A1(n17611), .A2(n17792), .ZN(n18295) );
NAND3_X1 U14092 ( .A1(n18300), .A2(n18299), .A3(n18298), .ZN(n5883) );
CLKBUF_X2 U14093 ( .A(n5883), .Z(n17612) );
CLKBUF_X2 U14094 ( .A(dii_data[73]), .Z(n17613) );
NAND2_X1 U14095 ( .A1(n17613), .A2(n17792), .ZN(n18299) );
NAND3_X1 U14096 ( .A1(n18304), .A2(n18303), .A3(n18302), .ZN(n5884) );
CLKBUF_X2 U14097 ( .A(n5884), .Z(n17614) );
CLKBUF_X2 U14098 ( .A(dii_data[72]), .Z(n17615) );
NAND2_X1 U14099 ( .A1(n17615), .A2(n17792), .ZN(n18303) );
CLKBUF_X1 U14100 ( .A(dii_data[71]), .Z(n17617) );
CLKBUF_X2 U14101 ( .A(n17617), .Z(n17616) );
NAND2_X1 U14102 ( .A1(n17616), .A2(n17793), .ZN(n18307) );
CLKBUF_X1 U14103 ( .A(dii_data[70]), .Z(n17619) );
CLKBUF_X2 U14104 ( .A(n17619), .Z(n17618) );
NAND2_X1 U14105 ( .A1(n17618), .A2(n17793), .ZN(n18311) );
CLKBUF_X1 U14106 ( .A(dii_data[69]), .Z(n17621) );
CLKBUF_X2 U14107 ( .A(n17621), .Z(n17620) );
NAND2_X1 U14108 ( .A1(n17620), .A2(n17793), .ZN(n18315) );
CLKBUF_X1 U14109 ( .A(dii_data[68]), .Z(n17623) );
CLKBUF_X2 U14110 ( .A(n17623), .Z(n17622) );
NAND2_X1 U14111 ( .A1(n17622), .A2(n17793), .ZN(n18319) );
CLKBUF_X1 U14112 ( .A(dii_data[67]), .Z(n17625) );
CLKBUF_X2 U14113 ( .A(n17625), .Z(n17624) );
NAND2_X1 U14114 ( .A1(n17624), .A2(n17793), .ZN(n18323) );
CLKBUF_X1 U14115 ( .A(n5890), .Z(n17626) );
NAND3_X1 U14116 ( .A1(n18328), .A2(n18327), .A3(n18326), .ZN(n5890) );
CLKBUF_X2 U14117 ( .A(dii_data[66]), .Z(n17627) );
NAND2_X1 U14118 ( .A1(n17627), .A2(n17793), .ZN(n18327) );
CLKBUF_X1 U14119 ( .A(n5891), .Z(n17628) );
NAND3_X1 U14120 ( .A1(n18332), .A2(n18331), .A3(n18330), .ZN(n5891) );
CLKBUF_X2 U14121 ( .A(dii_data[65]), .Z(n17629) );
NAND2_X1 U14122 ( .A1(n17629), .A2(n17793), .ZN(n18331) );
CLKBUF_X1 U14123 ( .A(n5892), .Z(n17630) );
NAND3_X1 U14124 ( .A1(n18336), .A2(n18335), .A3(n18334), .ZN(n5892) );
CLKBUF_X2 U14125 ( .A(dii_data[64]), .Z(n17631) );
NAND2_X1 U14126 ( .A1(n17631), .A2(n17793), .ZN(n18335) );
NAND3_X1 U14127 ( .A1(n18340), .A2(n18339), .A3(n18338), .ZN(n5893) );
CLKBUF_X2 U14128 ( .A(n5893), .Z(n17632) );
CLKBUF_X2 U14129 ( .A(dii_data[63]), .Z(n17633) );
NAND2_X1 U14130 ( .A1(n17633), .A2(n17793), .ZN(n18339) );
NAND3_X1 U14131 ( .A1(n18344), .A2(n18343), .A3(n18342), .ZN(n5894) );
CLKBUF_X2 U14132 ( .A(n5894), .Z(n17634) );
CLKBUF_X2 U14133 ( .A(dii_data[62]), .Z(n17635) );
NAND2_X1 U14134 ( .A1(n17635), .A2(n17793), .ZN(n18343) );
NAND3_X1 U14135 ( .A1(n18348), .A2(n18347), .A3(n18346), .ZN(n5895) );
CLKBUF_X2 U14136 ( .A(n5895), .Z(n17636) );
CLKBUF_X2 U14137 ( .A(dii_data[61]), .Z(n17637) );
NAND2_X1 U14138 ( .A1(n17637), .A2(n17793), .ZN(n18347) );
NAND3_X1 U14139 ( .A1(n18352), .A2(n18351), .A3(n18350), .ZN(n5896) );
CLKBUF_X2 U14140 ( .A(n5896), .Z(n17638) );
CLKBUF_X2 U14141 ( .A(dii_data[60]), .Z(n17639) );
NAND2_X1 U14142 ( .A1(n17639), .A2(n17794), .ZN(n18351) );
NAND3_X1 U14143 ( .A1(n18356), .A2(n18355), .A3(n18354), .ZN(n5897) );
CLKBUF_X2 U14144 ( .A(n5897), .Z(n17640) );
CLKBUF_X2 U14145 ( .A(dii_data[59]), .Z(n17641) );
NAND2_X1 U14146 ( .A1(n17641), .A2(n17794), .ZN(n18355) );
NAND3_X1 U14147 ( .A1(n18360), .A2(n18359), .A3(n18358), .ZN(n5898) );
CLKBUF_X2 U14148 ( .A(n5898), .Z(n17642) );
CLKBUF_X2 U14149 ( .A(dii_data[58]), .Z(n17643) );
NAND2_X1 U14150 ( .A1(n17643), .A2(n17794), .ZN(n18359) );
NAND3_X1 U14151 ( .A1(n18364), .A2(n18363), .A3(n18362), .ZN(n5899) );
CLKBUF_X2 U14152 ( .A(n5899), .Z(n17644) );
CLKBUF_X2 U14153 ( .A(dii_data[57]), .Z(n17645) );
NAND2_X1 U14154 ( .A1(n17645), .A2(n17794), .ZN(n18363) );
NAND3_X1 U14155 ( .A1(n18368), .A2(n18367), .A3(n18366), .ZN(n5900) );
CLKBUF_X2 U14156 ( .A(n5900), .Z(n17646) );
CLKBUF_X2 U14157 ( .A(dii_data[56]), .Z(n17647) );
NAND2_X1 U14158 ( .A1(n17647), .A2(n17794), .ZN(n18367) );
NAND3_X1 U14159 ( .A1(n18372), .A2(n18371), .A3(n18370), .ZN(n5901) );
CLKBUF_X2 U14160 ( .A(n5901), .Z(n17648) );
CLKBUF_X2 U14161 ( .A(dii_data[55]), .Z(n17649) );
NAND2_X1 U14162 ( .A1(n17649), .A2(n17794), .ZN(n18371) );
NAND3_X1 U14163 ( .A1(n18376), .A2(n18375), .A3(n18374), .ZN(n5902) );
CLKBUF_X2 U14164 ( .A(n5902), .Z(n17650) );
CLKBUF_X2 U14165 ( .A(dii_data[54]), .Z(n17651) );
NAND2_X1 U14166 ( .A1(n17651), .A2(n17794), .ZN(n18375) );
NAND3_X1 U14167 ( .A1(n18380), .A2(n18379), .A3(n18378), .ZN(n5903) );
CLKBUF_X2 U14168 ( .A(n5903), .Z(n17652) );
CLKBUF_X2 U14169 ( .A(dii_data[53]), .Z(n17653) );
NAND2_X1 U14170 ( .A1(n17653), .A2(n17794), .ZN(n18379) );
NAND3_X1 U14171 ( .A1(n18384), .A2(n18383), .A3(n18382), .ZN(n5904) );
CLKBUF_X2 U14172 ( .A(n5904), .Z(n17654) );
CLKBUF_X2 U14173 ( .A(dii_data[52]), .Z(n17655) );
NAND2_X1 U14174 ( .A1(n17655), .A2(n17794), .ZN(n18383) );
NAND3_X1 U14175 ( .A1(n18388), .A2(n18387), .A3(n18386), .ZN(n5905) );
CLKBUF_X2 U14176 ( .A(n5905), .Z(n17656) );
CLKBUF_X2 U14177 ( .A(dii_data[51]), .Z(n17657) );
NAND2_X1 U14178 ( .A1(n17657), .A2(n17794), .ZN(n18387) );
NAND3_X1 U14179 ( .A1(n18392), .A2(n18391), .A3(n18390), .ZN(n5906) );
CLKBUF_X2 U14180 ( .A(n5906), .Z(n17658) );
CLKBUF_X2 U14181 ( .A(dii_data[50]), .Z(n17659) );
NAND2_X1 U14182 ( .A1(n17659), .A2(n17794), .ZN(n18391) );
NAND3_X1 U14183 ( .A1(n18396), .A2(n18395), .A3(n18394), .ZN(n5907) );
CLKBUF_X2 U14184 ( .A(n5907), .Z(n17660) );
CLKBUF_X2 U14185 ( .A(dii_data[49]), .Z(n17661) );
NAND2_X1 U14186 ( .A1(n17661), .A2(n17795), .ZN(n18395) );
NAND3_X1 U14187 ( .A1(n18400), .A2(n18399), .A3(n18398), .ZN(n5908) );
CLKBUF_X2 U14188 ( .A(n5908), .Z(n17662) );
CLKBUF_X2 U14189 ( .A(dii_data[48]), .Z(n17663) );
NAND2_X1 U14190 ( .A1(n17663), .A2(n17795), .ZN(n18399) );
NAND3_X1 U14191 ( .A1(n18404), .A2(n18403), .A3(n18402), .ZN(n5909) );
CLKBUF_X2 U14192 ( .A(n5909), .Z(n17664) );
CLKBUF_X2 U14193 ( .A(dii_data[47]), .Z(n17665) );
NAND2_X1 U14194 ( .A1(n17665), .A2(n17795), .ZN(n18403) );
NAND3_X1 U14195 ( .A1(n18408), .A2(n18407), .A3(n18406), .ZN(n5910) );
CLKBUF_X2 U14196 ( .A(n5910), .Z(n17666) );
CLKBUF_X2 U14197 ( .A(dii_data[46]), .Z(n17667) );
NAND2_X1 U14198 ( .A1(n17667), .A2(n17795), .ZN(n18407) );
NAND3_X1 U14199 ( .A1(n18412), .A2(n18411), .A3(n18410), .ZN(n5911) );
CLKBUF_X2 U14200 ( .A(n5911), .Z(n17668) );
CLKBUF_X2 U14201 ( .A(dii_data[45]), .Z(n17669) );
NAND2_X1 U14202 ( .A1(n17669), .A2(n17795), .ZN(n18411) );
NAND3_X1 U14203 ( .A1(n18416), .A2(n18415), .A3(n18414), .ZN(n5912) );
CLKBUF_X2 U14204 ( .A(n5912), .Z(n17670) );
CLKBUF_X2 U14205 ( .A(dii_data[44]), .Z(n17671) );
NAND2_X1 U14206 ( .A1(n17671), .A2(n17795), .ZN(n18415) );
NAND3_X1 U14207 ( .A1(n18420), .A2(n18419), .A3(n18418), .ZN(n5913) );
CLKBUF_X2 U14208 ( .A(n5913), .Z(n17672) );
CLKBUF_X2 U14209 ( .A(dii_data[43]), .Z(n17673) );
NAND2_X1 U14210 ( .A1(n17673), .A2(n17795), .ZN(n18419) );
NAND3_X1 U14211 ( .A1(n18424), .A2(n18423), .A3(n18422), .ZN(n5914) );
CLKBUF_X2 U14212 ( .A(n5914), .Z(n17674) );
CLKBUF_X2 U14213 ( .A(dii_data[42]), .Z(n17675) );
NAND2_X1 U14214 ( .A1(n17675), .A2(n17795), .ZN(n18423) );
NAND3_X1 U14215 ( .A1(n18428), .A2(n18427), .A3(n18426), .ZN(n5915) );
CLKBUF_X2 U14216 ( .A(n5915), .Z(n17676) );
CLKBUF_X2 U14217 ( .A(dii_data[41]), .Z(n17677) );
NAND2_X1 U14218 ( .A1(n17677), .A2(n17795), .ZN(n18427) );
NAND3_X1 U14219 ( .A1(n18432), .A2(n18431), .A3(n18430), .ZN(n5916) );
CLKBUF_X2 U14220 ( .A(n5916), .Z(n17678) );
CLKBUF_X2 U14221 ( .A(dii_data[40]), .Z(n17679) );
NAND2_X1 U14222 ( .A1(n17679), .A2(n17795), .ZN(n18431) );
CLKBUF_X2 U14223 ( .A(n5917), .Z(n17680) );
CLKBUF_X2 U14224 ( .A(dii_data[39]), .Z(n17681) );
NAND2_X1 U14225 ( .A1(n17681), .A2(n17795), .ZN(n18435) );
CLKBUF_X2 U14226 ( .A(n5918), .Z(n17682) );
CLKBUF_X2 U14227 ( .A(dii_data[38]), .Z(n17683) );
NAND2_X1 U14228 ( .A1(n17683), .A2(n17796), .ZN(n18439) );
CLKBUF_X2 U14229 ( .A(n5919), .Z(n17684) );
CLKBUF_X2 U14230 ( .A(dii_data[37]), .Z(n17685) );
NAND2_X1 U14231 ( .A1(n17685), .A2(n17796), .ZN(n18443) );
CLKBUF_X2 U14232 ( .A(n5920), .Z(n17686) );
CLKBUF_X2 U14233 ( .A(dii_data[36]), .Z(n17687) );
NAND2_X1 U14234 ( .A1(n17687), .A2(n17796), .ZN(n18447) );
CLKBUF_X2 U14235 ( .A(n5921), .Z(n17688) );
CLKBUF_X2 U14236 ( .A(dii_data[35]), .Z(n17689) );
NAND2_X1 U14237 ( .A1(n17689), .A2(n17796), .ZN(n18451) );
CLKBUF_X2 U14238 ( .A(n5922), .Z(n17690) );
CLKBUF_X2 U14239 ( .A(dii_data[34]), .Z(n17691) );
NAND2_X1 U14240 ( .A1(n17691), .A2(n17796), .ZN(n18455) );
CLKBUF_X2 U14241 ( .A(n5923), .Z(n17692) );
CLKBUF_X2 U14242 ( .A(dii_data[33]), .Z(n17693) );
NAND2_X1 U14243 ( .A1(n17693), .A2(n17796), .ZN(n18459) );
CLKBUF_X2 U14244 ( .A(n5924), .Z(n17694) );
CLKBUF_X2 U14245 ( .A(dii_data[32]), .Z(n17695) );
NAND2_X1 U14246 ( .A1(n17695), .A2(n17796), .ZN(n18463) );
CLKBUF_X2 U14247 ( .A(n5925), .Z(n17696) );
CLKBUF_X2 U14248 ( .A(dii_data[31]), .Z(n17697) );
NAND2_X1 U14249 ( .A1(n17697), .A2(n17796), .ZN(n18467) );
CLKBUF_X2 U14250 ( .A(n5926), .Z(n17698) );
CLKBUF_X2 U14251 ( .A(dii_data[30]), .Z(n17699) );
NAND2_X1 U14252 ( .A1(n17699), .A2(n17796), .ZN(n18471) );
CLKBUF_X2 U14253 ( .A(n5927), .Z(n17700) );
CLKBUF_X2 U14254 ( .A(dii_data[29]), .Z(n17701) );
NAND2_X1 U14255 ( .A1(n17701), .A2(n17796), .ZN(n18475) );
CLKBUF_X2 U14256 ( .A(n5928), .Z(n17702) );
CLKBUF_X2 U14257 ( .A(dii_data[28]), .Z(n17703) );
NAND2_X1 U14258 ( .A1(n17703), .A2(n17796), .ZN(n18479) );
CLKBUF_X2 U14259 ( .A(n5929), .Z(n17704) );
CLKBUF_X2 U14260 ( .A(dii_data[27]), .Z(n17705) );
NAND2_X1 U14261 ( .A1(n17705), .A2(n17797), .ZN(n18483) );
CLKBUF_X2 U14262 ( .A(n5930), .Z(n17706) );
CLKBUF_X2 U14263 ( .A(dii_data[26]), .Z(n17707) );
NAND2_X1 U14264 ( .A1(n17707), .A2(n17797), .ZN(n18487) );
CLKBUF_X2 U14265 ( .A(n5931), .Z(n17708) );
CLKBUF_X2 U14266 ( .A(dii_data[25]), .Z(n17709) );
NAND2_X1 U14267 ( .A1(n17709), .A2(n17797), .ZN(n18491) );
CLKBUF_X2 U14268 ( .A(n5932), .Z(n17710) );
CLKBUF_X2 U14269 ( .A(dii_data[24]), .Z(n17711) );
NAND2_X1 U14270 ( .A1(n17711), .A2(n17797), .ZN(n18495) );
CLKBUF_X2 U14271 ( .A(n5933), .Z(n17712) );
CLKBUF_X2 U14272 ( .A(dii_data[23]), .Z(n17713) );
NAND2_X1 U14273 ( .A1(n17713), .A2(n17797), .ZN(n18499) );
CLKBUF_X2 U14274 ( .A(n5934), .Z(n17714) );
CLKBUF_X2 U14275 ( .A(dii_data[22]), .Z(n17715) );
NAND2_X1 U14276 ( .A1(n17715), .A2(n17797), .ZN(n18503) );
CLKBUF_X2 U14277 ( .A(n5935), .Z(n17716) );
CLKBUF_X2 U14278 ( .A(dii_data[21]), .Z(n17717) );
NAND2_X1 U14279 ( .A1(n17717), .A2(n17797), .ZN(n18507) );
CLKBUF_X2 U14280 ( .A(n5936), .Z(n17718) );
CLKBUF_X2 U14281 ( .A(dii_data[20]), .Z(n17719) );
NAND2_X1 U14282 ( .A1(n17719), .A2(n17797), .ZN(n18511) );
CLKBUF_X2 U14283 ( .A(n5937), .Z(n17720) );
CLKBUF_X2 U14284 ( .A(dii_data[19]), .Z(n17721) );
NAND2_X1 U14285 ( .A1(n17721), .A2(n17797), .ZN(n18515) );
CLKBUF_X2 U14286 ( .A(n5938), .Z(n17722) );
CLKBUF_X2 U14287 ( .A(dii_data[18]), .Z(n17723) );
NAND2_X1 U14288 ( .A1(n17723), .A2(n17797), .ZN(n18519) );
CLKBUF_X2 U14289 ( .A(n5939), .Z(n17724) );
CLKBUF_X2 U14290 ( .A(dii_data[17]), .Z(n17725) );
NAND2_X1 U14291 ( .A1(n17725), .A2(n17797), .ZN(n18523) );
CLKBUF_X2 U14292 ( .A(n5940), .Z(n17726) );
CLKBUF_X2 U14293 ( .A(dii_data[16]), .Z(n17727) );
NAND2_X1 U14294 ( .A1(n17727), .A2(n17798), .ZN(n18527) );
CLKBUF_X1 U14295 ( .A(dii_data[15]), .Z(n17728) );
NAND2_X1 U14296 ( .A1(n17728), .A2(n17798), .ZN(n18531) );
CLKBUF_X1 U14297 ( .A(dii_data[14]), .Z(n17729) );
NAND2_X1 U14298 ( .A1(n17729), .A2(n17798), .ZN(n18535) );
CLKBUF_X1 U14299 ( .A(dii_data[13]), .Z(n17730) );
NAND2_X1 U14300 ( .A1(n17730), .A2(n17798), .ZN(n18539) );
CLKBUF_X1 U14301 ( .A(dii_data[12]), .Z(n17731) );
NAND2_X1 U14302 ( .A1(n17731), .A2(n17798), .ZN(n18543) );
CLKBUF_X1 U14303 ( .A(dii_data[11]), .Z(n17732) );
NAND2_X1 U14304 ( .A1(n17732), .A2(n17798), .ZN(n18547) );
CLKBUF_X1 U14305 ( .A(dii_data[10]), .Z(n17733) );
NAND2_X1 U14306 ( .A1(n17733), .A2(n17798), .ZN(n18551) );
CLKBUF_X1 U14307 ( .A(dii_data[9]), .Z(n17734) );
NAND2_X1 U14308 ( .A1(n17734), .A2(n17798), .ZN(n18555) );
CLKBUF_X1 U14309 ( .A(dii_data[8]), .Z(n17735) );
NAND2_X1 U14310 ( .A1(n17735), .A2(n17798), .ZN(n18559) );
CLKBUF_X1 U14311 ( .A(dii_data[7]), .Z(n17736) );
NAND2_X1 U14312 ( .A1(n17736), .A2(n17798), .ZN(n18563) );
CLKBUF_X1 U14313 ( .A(dii_data[6]), .Z(n17737) );
NAND2_X1 U14314 ( .A1(n17737), .A2(n17798), .ZN(n18567) );
CLKBUF_X1 U14315 ( .A(dii_data[5]), .Z(n17738) );
NAND2_X1 U14316 ( .A1(n17738), .A2(n17799), .ZN(n18571) );
CLKBUF_X1 U14317 ( .A(dii_data[4]), .Z(n17739) );
NAND2_X1 U14318 ( .A1(n17739), .A2(n17799), .ZN(n18575) );
CLKBUF_X1 U14319 ( .A(dii_data[3]), .Z(n17740) );
NAND2_X1 U14320 ( .A1(n17740), .A2(n17799), .ZN(n18579) );
CLKBUF_X1 U14321 ( .A(dii_data[2]), .Z(n17741) );
NAND2_X1 U14322 ( .A1(n17741), .A2(n17799), .ZN(n18583) );
CLKBUF_X1 U14323 ( .A(dii_data[1]), .Z(n17742) );
NAND2_X1 U14324 ( .A1(n17742), .A2(n17799), .ZN(n18587) );
CLKBUF_X1 U14325 ( .A(dii_data[0]), .Z(n17743) );
NAND2_X1 U14326 ( .A1(n17743), .A2(n17799), .ZN(n18591) );
NAND3_X1 U14327 ( .A1(n18200), .A2(n18199), .A3(n18198), .ZN(n5957) );
CLKBUF_X2 U14328 ( .A(n5957), .Z(n17744) );
CLKBUF_X2 U14329 ( .A(dii_data[98]), .Z(n17745) );
NAND2_X1 U14330 ( .A1(n17745), .A2(n17790), .ZN(n18199) );
BUF_X16 U14331 ( .A(n11958), .Z(n17746) );
NAND2_X1 U14332 ( .A1(n17746), .A2(n11959), .ZN(n6284) );
NAND2_X1 U14333 ( .A1(n17990), .A2(cii_IV_vld), .ZN(n11958) );
BUF_X32 U14334 ( .A(n11930), .Z(n17747) );
NAND2_X1 U14335 ( .A1(cii_ctl_vld), .A2(n11971), .ZN(n11930) );
BUF_X16 U14336 ( .A(dii_last_word), .Z(n17749) );
NAND2_X1 U14337 ( .A1(n11927), .A2(n11928), .ZN(n6293) );
CLKBUF_X2 U14338 ( .A(n17749), .Z(n17748) );
OR3_X1 U14339 ( .A1(n18892), .A2(n17748), .A3(n11957), .ZN(n11949) );
NAND3_X1 U14340 ( .A1(n18744), .A2(n11946), .A3(n11947), .ZN(n6286) );
NAND3_X1 U14341 ( .A1(dii_data_type), .A2(dii_data_vld), .A3(n18617), .ZN(n11946) );
NAND2_X1 U14342 ( .A1(n11941), .A2(n18085), .ZN(n6288) );
MUX2_X1 U14343 ( .A(aad_byte_cnt[1]), .B(N2480), .S(n17837), .Z(n6019) );
CLKBUF_X1 U14344 ( .A(dii_data_size[0]), .Z(n17750) );
MUX2_X1 U14345 ( .A(enc_byte_cnt[0]), .B(N2349), .S(n17817), .Z(n5441) );
MUX2_X1 U14346 ( .A(enc_byte_cnt[1]), .B(N2350), .S(n17817), .Z(n5440) );
INV_X8 U14347 ( .A(rst), .ZN(n17751) );
INV_X8 U14348 ( .A(rst), .ZN(n17752) );
INV_X8 U14349 ( .A(rst), .ZN(n17753) );
INV_X4 U14350 ( .A(n16431), .ZN(n18634) );
INV_X4 U14351 ( .A(n18057), .ZN(n18036) );
INV_X4 U14352 ( .A(n18057), .ZN(n18037) );
INV_X4 U14353 ( .A(n17282), .ZN(n18044) );
INV_X4 U14354 ( .A(n18058), .ZN(n18045) );
INV_X4 U14355 ( .A(n18058), .ZN(n18046) );
INV_X4 U14356 ( .A(n18058), .ZN(n18048) );
INV_X4 U14357 ( .A(n18058), .ZN(n18049) );
INV_X4 U14358 ( .A(n18058), .ZN(n18050) );
INV_X4 U14359 ( .A(n18058), .ZN(n18047) );
INV_X4 U14360 ( .A(n17282), .ZN(n18042) );
INV_X4 U14361 ( .A(n18058), .ZN(n18041) );
INV_X4 U14362 ( .A(n18057), .ZN(n18039) );
INV_X4 U14363 ( .A(n18058), .ZN(n18040) );
INV_X4 U14364 ( .A(n18058), .ZN(n18038) );
INV_X4 U14365 ( .A(n17282), .ZN(n18043) );
INV_X4 U14366 ( .A(n18057), .ZN(n18052) );
INV_X4 U14367 ( .A(n18057), .ZN(n18053) );
INV_X4 U14368 ( .A(n18057), .ZN(n18051) );
INV_X4 U14369 ( .A(n17931), .ZN(n17928) );
INV_X4 U14370 ( .A(n17931), .ZN(n17922) );
INV_X4 U14371 ( .A(n17931), .ZN(n17923) );
INV_X4 U14372 ( .A(n17931), .ZN(n17924) );
INV_X4 U14373 ( .A(n17931), .ZN(n17925) );
INV_X4 U14374 ( .A(n17931), .ZN(n17926) );
INV_X4 U14375 ( .A(n17931), .ZN(n17927) );
INV_X4 U14376 ( .A(n17931), .ZN(n17929) );
INV_X4 U14377 ( .A(n17931), .ZN(n17919) );
INV_X4 U14378 ( .A(n17931), .ZN(n17920) );
INV_X4 U14379 ( .A(n17931), .ZN(n17921) );
INV_X4 U14380 ( .A(n17931), .ZN(n17930) );
INV_X4 U14381 ( .A(n16537), .ZN(n17849) );
INV_X4 U14382 ( .A(n16537), .ZN(n17850) );
INV_X4 U14383 ( .A(n16537), .ZN(n17851) );
INV_X4 U14384 ( .A(n18070), .ZN(n18058) );
INV_X4 U14385 ( .A(n17288), .ZN(n17931) );
INV_X4 U14386 ( .A(n18042), .ZN(n18060) );
INV_X4 U14387 ( .A(n18042), .ZN(n18063) );
INV_X4 U14388 ( .A(n18043), .ZN(n18062) );
INV_X4 U14389 ( .A(n18042), .ZN(n18061) );
INV_X4 U14390 ( .A(n18070), .ZN(n18059) );
INV_X4 U14391 ( .A(n18070), .ZN(n18064) );
INV_X4 U14392 ( .A(n18070), .ZN(n18065) );
INV_X4 U14393 ( .A(n18070), .ZN(n18066) );
INV_X4 U14394 ( .A(n16537), .ZN(n17848) );
INV_X4 U14395 ( .A(n18057), .ZN(n18055) );
INV_X4 U14396 ( .A(n18057), .ZN(n18054) );
INV_X4 U14397 ( .A(n17288), .ZN(n17932) );
INV_X4 U14398 ( .A(n17754), .ZN(n17944) );
INV_X4 U14399 ( .A(n17754), .ZN(n17943) );
INV_X4 U14400 ( .A(n17754), .ZN(n17942) );
INV_X4 U14401 ( .A(n17754), .ZN(n17941) );
INV_X4 U14402 ( .A(n17754), .ZN(n17939) );
INV_X4 U14403 ( .A(n17754), .ZN(n17940) );
INV_X4 U14404 ( .A(n17754), .ZN(n17938) );
INV_X4 U14405 ( .A(n17754), .ZN(n17937) );
INV_X4 U14406 ( .A(n17754), .ZN(n17936) );
INV_X4 U14407 ( .A(n17754), .ZN(n17934) );
INV_X4 U14408 ( .A(n18057), .ZN(n18056) );
INV_X4 U14409 ( .A(n17285), .ZN(n17949) );
INV_X4 U14410 ( .A(n17285), .ZN(n17950) );
INV_X4 U14411 ( .A(n17285), .ZN(n17951) );
INV_X4 U14412 ( .A(n17285), .ZN(n17952) );
INV_X4 U14413 ( .A(n17285), .ZN(n17953) );
INV_X4 U14414 ( .A(n17285), .ZN(n17954) );
INV_X4 U14415 ( .A(n17285), .ZN(n17955) );
INV_X4 U14416 ( .A(n17285), .ZN(n17956) );
INV_X4 U14417 ( .A(n18083), .ZN(n17779) );
INV_X4 U14418 ( .A(n18083), .ZN(n17780) );
INV_X4 U14419 ( .A(n18083), .ZN(n17781) );
INV_X4 U14420 ( .A(n18083), .ZN(n17782) );
INV_X4 U14421 ( .A(n18083), .ZN(n17783) );
INV_X4 U14422 ( .A(n18083), .ZN(n17784) );
INV_X4 U14423 ( .A(n18083), .ZN(n17785) );
INV_X4 U14424 ( .A(n18083), .ZN(n17786) );
INV_X4 U14425 ( .A(n17754), .ZN(n17935) );
INV_X4 U14426 ( .A(n17754), .ZN(n17945) );
INV_X4 U14427 ( .A(n17285), .ZN(n17957) );
INV_X4 U14428 ( .A(n18083), .ZN(n17787) );
NOR2_X2 U14429 ( .A1(n16325), .A2(n16326), .ZN(n16209) );
NAND2_X2 U14430 ( .A1(n16431), .A2(n16432), .ZN(n16325) );
INV_X4 U14431 ( .A(n17282), .ZN(n18070) );
INV_X4 U14432 ( .A(n18070), .ZN(n18067) );
INV_X4 U14433 ( .A(n18070), .ZN(n18068) );
INV_X4 U14434 ( .A(n14167), .ZN(n17900) );
INV_X4 U14435 ( .A(n14167), .ZN(n17901) );
INV_X4 U14436 ( .A(n14167), .ZN(n17902) );
INV_X4 U14437 ( .A(n14167), .ZN(n17903) );
INV_X4 U14438 ( .A(n14167), .ZN(n17904) );
INV_X4 U14439 ( .A(n14167), .ZN(n17905) );
INV_X4 U14440 ( .A(n15509), .ZN(n17864) );
INV_X4 U14441 ( .A(n17877), .ZN(n17876) );
INV_X4 U14442 ( .A(n17284), .ZN(n17910) );
INV_X4 U14443 ( .A(n17284), .ZN(n17909) );
INV_X4 U14444 ( .A(n17284), .ZN(n17914) );
INV_X4 U14445 ( .A(n17284), .ZN(n17913) );
INV_X4 U14446 ( .A(n17284), .ZN(n17912) );
INV_X4 U14447 ( .A(n17284), .ZN(n17911) );
INV_X4 U14448 ( .A(n17284), .ZN(n17915) );
INV_X4 U14449 ( .A(n17285), .ZN(n17946) );
INV_X4 U14450 ( .A(n17285), .ZN(n17947) );
INV_X4 U14451 ( .A(n17285), .ZN(n17948) );
INV_X4 U14452 ( .A(n18083), .ZN(n17776) );
INV_X4 U14453 ( .A(n18083), .ZN(n17777) );
INV_X4 U14454 ( .A(n18083), .ZN(n17778) );
INV_X4 U14455 ( .A(n18084), .ZN(n17791) );
INV_X4 U14456 ( .A(n18084), .ZN(n17792) );
INV_X4 U14457 ( .A(n18084), .ZN(n17793) );
INV_X4 U14458 ( .A(n18084), .ZN(n17794) );
INV_X4 U14459 ( .A(n18084), .ZN(n17795) );
INV_X4 U14460 ( .A(n18084), .ZN(n17796) );
INV_X4 U14461 ( .A(n18084), .ZN(n17797) );
INV_X4 U14462 ( .A(n18084), .ZN(n17798) );
INV_X4 U14463 ( .A(n18043), .ZN(n18069) );
INV_X4 U14464 ( .A(n17754), .ZN(n17933) );
INV_X4 U14465 ( .A(n18602), .ZN(n18014) );
INV_X4 U14466 ( .A(n18070), .ZN(n18057) );
INV_X4 U14467 ( .A(n18084), .ZN(n17799) );
INV_X4 U14468 ( .A(n17284), .ZN(n17916) );
INV_X4 U14469 ( .A(n17877), .ZN(n17875) );
INV_X4 U14470 ( .A(n17877), .ZN(n17874) );
INV_X4 U14471 ( .A(n15509), .ZN(n17862) );
INV_X4 U14472 ( .A(n15509), .ZN(n17863) );
INV_X4 U14473 ( .A(n15509), .ZN(n17861) );
INV_X4 U14474 ( .A(n15509), .ZN(n17860) );
INV_X4 U14475 ( .A(n11961), .ZN(n17842) );
INV_X4 U14476 ( .A(n11961), .ZN(n17843) );
INV_X4 U14477 ( .A(n11961), .ZN(n17844) );
INV_X4 U14478 ( .A(n11961), .ZN(n17845) );
INV_X4 U14479 ( .A(n11961), .ZN(n17846) );
INV_X4 U14480 ( .A(n11961), .ZN(n17847) );
INV_X4 U14481 ( .A(n17989), .ZN(n17982) );
INV_X4 U14482 ( .A(n17989), .ZN(n17981) );
INV_X4 U14483 ( .A(n17989), .ZN(n17980) );
INV_X4 U14484 ( .A(n17989), .ZN(n17979) );
INV_X4 U14485 ( .A(n17989), .ZN(n17978) );
INV_X4 U14486 ( .A(n17989), .ZN(n17977) );
INV_X4 U14487 ( .A(n18602), .ZN(n18006) );
INV_X4 U14488 ( .A(n18602), .ZN(n18007) );
INV_X4 U14489 ( .A(n18602), .ZN(n18008) );
INV_X4 U14490 ( .A(n18602), .ZN(n18009) );
INV_X4 U14491 ( .A(n18602), .ZN(n18010) );
INV_X4 U14492 ( .A(n18602), .ZN(n18011) );
INV_X4 U14493 ( .A(n18602), .ZN(n18012) );
INV_X4 U14494 ( .A(n18602), .ZN(n18013) );
INV_X4 U14495 ( .A(n17989), .ZN(n17987) );
INV_X4 U14496 ( .A(n17989), .ZN(n17986) );
INV_X4 U14497 ( .A(n17989), .ZN(n17985) );
INV_X4 U14498 ( .A(n17989), .ZN(n17984) );
INV_X4 U14499 ( .A(n17989), .ZN(n17983) );
INV_X4 U14500 ( .A(n18085), .ZN(n17803) );
INV_X4 U14501 ( .A(n18085), .ZN(n17804) );
INV_X4 U14502 ( .A(n18085), .ZN(n17805) );
INV_X4 U14503 ( .A(n18085), .ZN(n17806) );
INV_X4 U14504 ( .A(n18085), .ZN(n17807) );
INV_X4 U14505 ( .A(n18085), .ZN(n17808) );
INV_X4 U14506 ( .A(n18085), .ZN(n17809) );
INV_X4 U14507 ( .A(n18085), .ZN(n17810) );
INV_X4 U14508 ( .A(n18085), .ZN(n17811) );
INV_X4 U14509 ( .A(n17989), .ZN(n17988) );
NOR2_X2 U14510 ( .A1(n15805), .A2(n15806), .ZN(n15663) );
BUF_X4 U14511 ( .A(n11956), .Z(n18026) );
BUF_X4 U14512 ( .A(n11956), .Z(n18034) );
BUF_X4 U14513 ( .A(n11956), .Z(n18033) );
BUF_X4 U14514 ( .A(n11956), .Z(n18032) );
BUF_X4 U14515 ( .A(n11956), .Z(n18031) );
BUF_X4 U14516 ( .A(n11956), .Z(n18030) );
BUF_X4 U14517 ( .A(n11956), .Z(n18029) );
BUF_X4 U14518 ( .A(n11956), .Z(n18028) );
BUF_X4 U14519 ( .A(n11956), .Z(n18027) );
BUF_X4 U14520 ( .A(n11956), .Z(n18035) );
INV_X4 U14521 ( .A(n15501), .ZN(n17877) );
INV_X4 U14522 ( .A(n17916), .ZN(n17918) );
INV_X4 U14523 ( .A(n17916), .ZN(n17917) );
INV_X4 U14524 ( .A(n18000), .ZN(n17996) );
INV_X4 U14525 ( .A(n18001), .ZN(n17999) );
INV_X4 U14526 ( .A(n17905), .ZN(n17906) );
INV_X4 U14527 ( .A(n17903), .ZN(n17907) );
INV_X4 U14528 ( .A(n12238), .ZN(n17990) );
INV_X4 U14529 ( .A(n15508), .ZN(n17857) );
INV_X4 U14530 ( .A(n17904), .ZN(n17908) );
INV_X4 U14531 ( .A(n18084), .ZN(n17788) );
INV_X4 U14532 ( .A(n18084), .ZN(n17789) );
INV_X4 U14533 ( .A(n18084), .ZN(n17790) );
INV_X4 U14534 ( .A(n11961), .ZN(n17841) );
BUF_X4 U14535 ( .A(n11956), .Z(n18025) );
BUF_X4 U14536 ( .A(n11956), .Z(n18024) );
BUF_X4 U14537 ( .A(n11956), .Z(n18023) );
BUF_X4 U14538 ( .A(n11956), .Z(n18021) );
BUF_X4 U14539 ( .A(n11956), .Z(n18022) );
BUF_X4 U14540 ( .A(n11956), .Z(n18019) );
BUF_X4 U14541 ( .A(n11956), .Z(n18018) );
BUF_X4 U14542 ( .A(n11956), .Z(n18017) );
BUF_X4 U14543 ( .A(n11956), .Z(n18016) );
BUF_X4 U14544 ( .A(n11956), .Z(n18015) );
BUF_X4 U14545 ( .A(n11956), .Z(n18020) );
INV_X4 U14546 ( .A(n12238), .ZN(n17989) );
INV_X4 U14547 ( .A(n14564), .ZN(n17867) );
INV_X4 U14548 ( .A(n14564), .ZN(n17866) );
INV_X4 U14549 ( .A(n18000), .ZN(n17997) );
INV_X4 U14550 ( .A(n18001), .ZN(n17998) );
INV_X4 U14551 ( .A(n11946), .ZN(n17839) );
INV_X4 U14552 ( .A(n11946), .ZN(n17838) );
INV_X4 U14553 ( .A(n17988), .ZN(n17993) );
INV_X4 U14554 ( .A(n17988), .ZN(n17992) );
INV_X4 U14555 ( .A(n17988), .ZN(n17991) );
INV_X4 U14556 ( .A(n15508), .ZN(n17858) );
INV_X4 U14557 ( .A(n11946), .ZN(n17840) );
INV_X4 U14558 ( .A(n15508), .ZN(n17859) );
INV_X4 U14559 ( .A(n11939), .ZN(n17812) );
INV_X4 U14560 ( .A(n11939), .ZN(n17813) );
INV_X4 U14561 ( .A(n11939), .ZN(n17814) );
INV_X4 U14562 ( .A(n11939), .ZN(n17815) );
INV_X4 U14563 ( .A(n11939), .ZN(n17816) );
INV_X4 U14564 ( .A(n11939), .ZN(n17817) );
INV_X4 U14565 ( .A(n17286), .ZN(n17968) );
INV_X4 U14566 ( .A(n17286), .ZN(n17969) );
INV_X4 U14567 ( .A(n17286), .ZN(n17970) );
INV_X4 U14568 ( .A(n17286), .ZN(n17971) );
INV_X4 U14569 ( .A(n17286), .ZN(n17972) );
INV_X4 U14570 ( .A(n17286), .ZN(n17973) );
INV_X4 U14571 ( .A(n17286), .ZN(n17974) );
INV_X4 U14572 ( .A(n17286), .ZN(n17975) );
INV_X4 U14573 ( .A(n17885), .ZN(n17884) );
INV_X4 U14574 ( .A(n17885), .ZN(n17883) );
INV_X4 U14575 ( .A(n15507), .ZN(n17854) );
INV_X4 U14576 ( .A(n15507), .ZN(n17855) );
INV_X4 U14577 ( .A(n18602), .ZN(n18004) );
INV_X4 U14578 ( .A(n18602), .ZN(n18005) );
INV_X4 U14579 ( .A(n18602), .ZN(n18003) );
INV_X4 U14580 ( .A(n15507), .ZN(n17852) );
INV_X4 U14581 ( .A(n15507), .ZN(n17853) );
INV_X4 U14582 ( .A(n18085), .ZN(n17800) );
INV_X4 U14583 ( .A(n18085), .ZN(n17801) );
INV_X4 U14584 ( .A(n18085), .ZN(n17802) );
INV_X4 U14585 ( .A(n17286), .ZN(n17976) );
INV_X4 U14586 ( .A(n15507), .ZN(n17856) );
NAND2_X2 U14587 ( .A1(n17934), .A2(n15644), .ZN(n15946) );
OR2_X2 U14588 ( .A1(n18744), .A2(n16542), .ZN(n17754) );
NAND2_X2 U14589 ( .A1(n15946), .A2(n15947), .ZN(n15805) );
NOR4_X2 U14590 ( .A1(n15644), .A2(n19202), .A3(n17755), .A4(n15509), .ZN(n15272) );
INV_X4 U14591 ( .A(n18633), .ZN(n11956) );
NOR2_X2 U14592 ( .A1(n17291), .A2(n18059), .ZN(n17280) );
INV_X4 U14593 ( .A(n17283), .ZN(n18000) );
INV_X4 U14594 ( .A(n14422), .ZN(n17885) );
INV_X4 U14595 ( .A(n11946), .ZN(n17837) );
INV_X4 U14596 ( .A(n17756), .ZN(n17872) );
INV_X4 U14597 ( .A(n15501), .ZN(n17873) );
INV_X4 U14598 ( .A(n17891), .ZN(n17887) );
INV_X4 U14599 ( .A(n17287), .ZN(n17892) );
INV_X4 U14600 ( .A(n17757), .ZN(n17880) );
NOR2_X2 U14601 ( .A1(n17886), .A2(n14190), .ZN(n14189) );
NOR2_X2 U14602 ( .A1(n17886), .A2(n14219), .ZN(n14218) );
NOR2_X2 U14603 ( .A1(n17886), .A2(n14248), .ZN(n14247) );
NOR2_X2 U14604 ( .A1(n17886), .A2(n14277), .ZN(n14276) );
NOR2_X2 U14605 ( .A1(n17886), .A2(n14306), .ZN(n14305) );
NOR2_X2 U14606 ( .A1(n17886), .A2(n14335), .ZN(n14334) );
NOR2_X2 U14607 ( .A1(n17886), .A2(n14364), .ZN(n14363) );
NOR2_X2 U14608 ( .A1(n17891), .A2(n14396), .ZN(n14395) );
NOR2_X2 U14609 ( .A1(n17866), .A2(n14191), .ZN(n14188) );
NOR2_X2 U14610 ( .A1(n17865), .A2(n14220), .ZN(n14217) );
NOR2_X2 U14611 ( .A1(n17865), .A2(n14249), .ZN(n14246) );
NOR2_X2 U14612 ( .A1(n17865), .A2(n14278), .ZN(n14275) );
NOR2_X2 U14613 ( .A1(n17865), .A2(n14307), .ZN(n14304) );
NOR2_X2 U14614 ( .A1(n17866), .A2(n14336), .ZN(n14333) );
NOR2_X2 U14615 ( .A1(n17866), .A2(n14365), .ZN(n14362) );
NOR2_X2 U14616 ( .A1(n17866), .A2(n14397), .ZN(n14394) );
INV_X4 U14617 ( .A(n17757), .ZN(n17881) );
INV_X4 U14618 ( .A(n17756), .ZN(n17871) );
INV_X4 U14619 ( .A(n17756), .ZN(n17870) );
INV_X4 U14620 ( .A(n17755), .ZN(n17869) );
INV_X4 U14621 ( .A(n17755), .ZN(n17868) );
INV_X4 U14622 ( .A(n17758), .ZN(n17879) );
INV_X4 U14623 ( .A(n17758), .ZN(n17878) );
INV_X4 U14624 ( .A(n17283), .ZN(n18001) );
INV_X4 U14625 ( .A(n17988), .ZN(n17995) );
INV_X4 U14626 ( .A(n17985), .ZN(n17994) );
INV_X4 U14627 ( .A(n14564), .ZN(n17865) );
INV_X4 U14628 ( .A(n17289), .ZN(n17963) );
INV_X4 U14629 ( .A(n17289), .ZN(n17962) );
INV_X4 U14630 ( .A(n17289), .ZN(n17960) );
INV_X4 U14631 ( .A(n17289), .ZN(n17959) );
INV_X4 U14632 ( .A(n17289), .ZN(n17961) );
INV_X4 U14633 ( .A(n17289), .ZN(n17964) );
INV_X4 U14634 ( .A(n15504), .ZN(n19202) );
INV_X4 U14635 ( .A(n17891), .ZN(n17889) );
INV_X4 U14636 ( .A(n17886), .ZN(n17888) );
INV_X4 U14637 ( .A(n17287), .ZN(n17895) );
INV_X4 U14638 ( .A(n17287), .ZN(n17894) );
INV_X4 U14639 ( .A(n17287), .ZN(n17893) );
INV_X4 U14640 ( .A(n17286), .ZN(n17965) );
INV_X4 U14641 ( .A(n17286), .ZN(n17966) );
INV_X4 U14642 ( .A(n17286), .ZN(n17967) );
INV_X4 U14643 ( .A(n17885), .ZN(n17882) );
INV_X4 U14644 ( .A(n17886), .ZN(n17890) );
INV_X4 U14645 ( .A(n17287), .ZN(n17896) );
NOR3_X2 U14646 ( .A1(n19204), .A2(n19205), .A3(n18071), .ZN(n15509) );
AND2_X2 U14647 ( .A1(n17887), .A2(n15309), .ZN(n17755) );
NAND2_X2 U14648 ( .A1(n14564), .A2(n14422), .ZN(n15508) );
NOR2_X2 U14649 ( .A1(n17848), .A2(n17857), .ZN(n16083) );
NOR2_X2 U14650 ( .A1(n17864), .A2(n18075), .ZN(n16542) );
NOR4_X2 U14651 ( .A1(n14583), .A2(n14584), .A3(n14585), .A4(n18735), .ZN(n14582) );
NOR2_X2 U14652 ( .A1(n19032), .A2(n17900), .ZN(n14584) );
NOR4_X2 U14653 ( .A1(n14605), .A2(n14606), .A3(n14607), .A4(n18734), .ZN(n14604) );
NOR2_X2 U14654 ( .A1(n19034), .A2(n17900), .ZN(n14606) );
NOR4_X2 U14655 ( .A1(n14626), .A2(n14627), .A3(n14628), .A4(n18733), .ZN(n14625) );
NOR2_X2 U14656 ( .A1(n19036), .A2(n17900), .ZN(n14627) );
NOR4_X2 U14657 ( .A1(n14647), .A2(n14648), .A3(n14649), .A4(n18732), .ZN(n14646) );
NOR2_X2 U14658 ( .A1(n19038), .A2(n17900), .ZN(n14648) );
NOR4_X2 U14659 ( .A1(n14668), .A2(n14669), .A3(n14670), .A4(n18731), .ZN(n14667) );
NOR2_X2 U14660 ( .A1(n19040), .A2(n17900), .ZN(n14669) );
NOR4_X2 U14661 ( .A1(n14689), .A2(n14690), .A3(n14691), .A4(n18730), .ZN(n14688) );
NOR2_X2 U14662 ( .A1(n19042), .A2(n17900), .ZN(n14690) );
NOR4_X2 U14663 ( .A1(n14710), .A2(n14711), .A3(n14712), .A4(n18729), .ZN(n14709) );
NOR2_X2 U14664 ( .A1(n19044), .A2(n17900), .ZN(n14711) );
NOR4_X2 U14665 ( .A1(n14731), .A2(n14732), .A3(n14733), .A4(n18728), .ZN(n14730) );
NOR2_X2 U14666 ( .A1(n19046), .A2(n17900), .ZN(n14732) );
NOR4_X2 U14667 ( .A1(n14754), .A2(n14755), .A3(n14756), .A4(n18727), .ZN(n14753) );
NOR2_X2 U14668 ( .A1(n19048), .A2(n17900), .ZN(n14755) );
NOR4_X2 U14669 ( .A1(n14778), .A2(n14779), .A3(n14780), .A4(n18726), .ZN(n14777) );
NOR2_X2 U14670 ( .A1(n19050), .A2(n17900), .ZN(n14779) );
NOR4_X2 U14671 ( .A1(n14800), .A2(n14801), .A3(n14802), .A4(n18725), .ZN(n14799) );
NOR2_X2 U14672 ( .A1(n19052), .A2(n17900), .ZN(n14801) );
NOR4_X2 U14673 ( .A1(n14822), .A2(n14823), .A3(n14824), .A4(n18724), .ZN(n14821) );
NOR2_X2 U14674 ( .A1(n19054), .A2(n17900), .ZN(n14823) );
NOR4_X2 U14675 ( .A1(n14844), .A2(n14845), .A3(n14846), .A4(n18723), .ZN(n14843) );
NOR2_X2 U14676 ( .A1(n19056), .A2(n17901), .ZN(n14845) );
NOR4_X2 U14677 ( .A1(n14866), .A2(n14867), .A3(n14868), .A4(n18722), .ZN(n14865) );
NOR2_X2 U14678 ( .A1(n19058), .A2(n17901), .ZN(n14867) );
NOR4_X2 U14679 ( .A1(n14888), .A2(n14889), .A3(n14890), .A4(n18721), .ZN(n14887) );
NOR2_X2 U14680 ( .A1(n19060), .A2(n17901), .ZN(n14889) );
NOR4_X2 U14681 ( .A1(n14910), .A2(n14911), .A3(n14912), .A4(n18720), .ZN(n14909) );
NOR2_X2 U14682 ( .A1(n19062), .A2(n17901), .ZN(n14911) );
NOR4_X2 U14683 ( .A1(n14933), .A2(n14934), .A3(n14935), .A4(n18719), .ZN(n14932) );
NOR2_X2 U14684 ( .A1(n19064), .A2(n17901), .ZN(n14934) );
NOR4_X2 U14685 ( .A1(n14957), .A2(n14958), .A3(n14959), .A4(n18718), .ZN(n14956) );
NOR2_X2 U14686 ( .A1(n19066), .A2(n17901), .ZN(n14958) );
NOR4_X2 U14687 ( .A1(n14979), .A2(n14980), .A3(n14981), .A4(n18717), .ZN(n14978) );
NOR2_X2 U14688 ( .A1(n19068), .A2(n17901), .ZN(n14980) );
NOR4_X2 U14689 ( .A1(n15001), .A2(n15002), .A3(n15003), .A4(n18716), .ZN(n15000) );
NOR2_X2 U14690 ( .A1(n19070), .A2(n17901), .ZN(n15002) );
NOR4_X2 U14691 ( .A1(n15023), .A2(n15024), .A3(n15025), .A4(n18715), .ZN(n15022) );
NOR2_X2 U14692 ( .A1(n19072), .A2(n17901), .ZN(n15024) );
NOR4_X2 U14693 ( .A1(n15045), .A2(n15046), .A3(n15047), .A4(n18714), .ZN(n15044) );
NOR2_X2 U14694 ( .A1(n19074), .A2(n17901), .ZN(n15046) );
NOR4_X2 U14695 ( .A1(n15067), .A2(n15068), .A3(n15069), .A4(n18713), .ZN(n15066) );
NOR2_X2 U14696 ( .A1(n19076), .A2(n17901), .ZN(n15068) );
NOR4_X2 U14697 ( .A1(n15089), .A2(n15090), .A3(n15091), .A4(n18712), .ZN(n15088) );
NOR2_X2 U14698 ( .A1(n19078), .A2(n17901), .ZN(n15090) );
NOR4_X2 U14699 ( .A1(n15113), .A2(n15114), .A3(n15115), .A4(n18711), .ZN(n15112) );
NOR2_X2 U14700 ( .A1(n19081), .A2(n17902), .ZN(n15114) );
NOR4_X2 U14701 ( .A1(n15136), .A2(n15137), .A3(n15138), .A4(n18710), .ZN(n15135) );
NOR2_X2 U14702 ( .A1(n19084), .A2(n17902), .ZN(n15137) );
NOR4_X2 U14703 ( .A1(n15158), .A2(n15159), .A3(n15160), .A4(n18709), .ZN(n15157) );
NOR2_X2 U14704 ( .A1(n19087), .A2(n17902), .ZN(n15159) );
NOR4_X2 U14705 ( .A1(n15180), .A2(n15181), .A3(n15182), .A4(n18708), .ZN(n15179) );
NOR2_X2 U14706 ( .A1(n19090), .A2(n17902), .ZN(n15181) );
NOR4_X2 U14707 ( .A1(n15202), .A2(n15203), .A3(n15204), .A4(n18707), .ZN(n15201) );
NOR2_X2 U14708 ( .A1(n19093), .A2(n17902), .ZN(n15203) );
NOR4_X2 U14709 ( .A1(n15224), .A2(n15225), .A3(n15226), .A4(n18706), .ZN(n15223) );
NOR2_X2 U14710 ( .A1(n19096), .A2(n17902), .ZN(n15225) );
NOR4_X2 U14711 ( .A1(n15246), .A2(n15247), .A3(n15248), .A4(n18705), .ZN(n15245) );
NOR2_X2 U14712 ( .A1(n19099), .A2(n17902), .ZN(n15247) );
NOR4_X2 U14713 ( .A1(n15268), .A2(n15269), .A3(n15270), .A4(n18704), .ZN(n15267) );
NOR2_X2 U14714 ( .A1(n19102), .A2(n17902), .ZN(n15269) );
NOR4_X2 U14715 ( .A1(n15292), .A2(n15293), .A3(n15294), .A4(n18703), .ZN(n15291) );
NOR2_X2 U14716 ( .A1(n19105), .A2(n17902), .ZN(n15293) );
NOR4_X2 U14717 ( .A1(n15318), .A2(n15319), .A3(n15320), .A4(n18702), .ZN(n15317) );
NOR2_X2 U14718 ( .A1(n19108), .A2(n17902), .ZN(n15319) );
NOR4_X2 U14719 ( .A1(n15342), .A2(n15343), .A3(n15344), .A4(n18701), .ZN(n15341) );
NOR2_X2 U14720 ( .A1(n19111), .A2(n17902), .ZN(n15343) );
NOR4_X2 U14721 ( .A1(n15366), .A2(n15367), .A3(n15368), .A4(n18700), .ZN(n15365) );
NOR2_X2 U14722 ( .A1(n19114), .A2(n17902), .ZN(n15367) );
NOR4_X2 U14723 ( .A1(n15390), .A2(n15391), .A3(n15392), .A4(n18699), .ZN(n15389) );
NOR2_X2 U14724 ( .A1(n19117), .A2(n17903), .ZN(n15391) );
NOR4_X2 U14725 ( .A1(n15414), .A2(n15415), .A3(n15416), .A4(n18698), .ZN(n15413) );
NOR2_X2 U14726 ( .A1(n19120), .A2(n17903), .ZN(n15415) );
NOR4_X2 U14727 ( .A1(n15438), .A2(n15439), .A3(n15440), .A4(n18697), .ZN(n15437) );
NOR2_X2 U14728 ( .A1(n19123), .A2(n17903), .ZN(n15439) );
NOR4_X2 U14729 ( .A1(n15462), .A2(n15463), .A3(n15464), .A4(n18696), .ZN(n15461) );
NOR2_X2 U14730 ( .A1(n19126), .A2(n17903), .ZN(n15463) );
NOR4_X2 U14731 ( .A1(n18695), .A2(n15488), .A3(n15489), .A4(n15490), .ZN(n15487) );
NOR2_X2 U14732 ( .A1(n15491), .A2(n17284), .ZN(n15490) );
NOR4_X2 U14733 ( .A1(n18694), .A2(n15517), .A3(n15518), .A4(n15519), .ZN(n15516) );
NOR2_X2 U14734 ( .A1(n15520), .A2(n17918), .ZN(n15519) );
NOR4_X2 U14735 ( .A1(n18693), .A2(n15538), .A3(n15539), .A4(n15540), .ZN(n15537) );
NOR2_X2 U14736 ( .A1(n15541), .A2(n17918), .ZN(n15540) );
NOR4_X2 U14737 ( .A1(n18692), .A2(n15559), .A3(n15560), .A4(n15561), .ZN(n15558) );
NOR2_X2 U14738 ( .A1(n15562), .A2(n17918), .ZN(n15561) );
NOR4_X2 U14739 ( .A1(n18691), .A2(n15580), .A3(n15581), .A4(n15582), .ZN(n15579) );
NOR2_X2 U14740 ( .A1(n15583), .A2(n17918), .ZN(n15582) );
NOR4_X2 U14741 ( .A1(n18658), .A2(n16220), .A3(n16221), .A4(n16222), .ZN(n16219) );
NOR2_X2 U14742 ( .A1(n16223), .A2(n17917), .ZN(n16222) );
NOR4_X2 U14743 ( .A1(n18657), .A2(n16234), .A3(n16235), .A4(n16236), .ZN(n16233) );
NOR2_X2 U14744 ( .A1(n16237), .A2(n17917), .ZN(n16236) );
NOR4_X2 U14745 ( .A1(n18656), .A2(n16248), .A3(n16249), .A4(n16250), .ZN(n16247) );
NOR2_X2 U14746 ( .A1(n16251), .A2(n17917), .ZN(n16250) );
NOR4_X2 U14747 ( .A1(n18655), .A2(n16262), .A3(n16263), .A4(n16264), .ZN(n16261) );
NOR2_X2 U14748 ( .A1(n16265), .A2(n17284), .ZN(n16264) );
NOR4_X2 U14749 ( .A1(n18654), .A2(n16276), .A3(n16277), .A4(n16278), .ZN(n16275) );
NOR2_X2 U14750 ( .A1(n16279), .A2(n17284), .ZN(n16278) );
NOR4_X2 U14751 ( .A1(n18653), .A2(n16290), .A3(n16291), .A4(n16292), .ZN(n16289) );
NOR2_X2 U14752 ( .A1(n16293), .A2(n17284), .ZN(n16292) );
NOR4_X2 U14753 ( .A1(n18652), .A2(n16304), .A3(n16305), .A4(n16306), .ZN(n16303) );
NOR2_X2 U14754 ( .A1(n16307), .A2(n17284), .ZN(n16306) );
NOR4_X2 U14755 ( .A1(n18651), .A2(n16318), .A3(n16319), .A4(n16320), .ZN(n16317) );
NOR2_X2 U14756 ( .A1(n16321), .A2(n17284), .ZN(n16320) );
NOR4_X2 U14757 ( .A1(n18690), .A2(n15659), .A3(n15660), .A4(n15661), .ZN(n15658) );
NOR2_X2 U14758 ( .A1(n15662), .A2(n17918), .ZN(n15661) );
NOR4_X2 U14759 ( .A1(n18689), .A2(n15679), .A3(n15680), .A4(n15681), .ZN(n15678) );
NOR2_X2 U14760 ( .A1(n15682), .A2(n17918), .ZN(n15681) );
NOR4_X2 U14761 ( .A1(n18688), .A2(n15698), .A3(n15699), .A4(n15700), .ZN(n15697) );
NOR2_X2 U14762 ( .A1(n15701), .A2(n17918), .ZN(n15700) );
NOR4_X2 U14763 ( .A1(n18687), .A2(n15717), .A3(n15718), .A4(n15719), .ZN(n15716) );
NOR2_X2 U14764 ( .A1(n15720), .A2(n17918), .ZN(n15719) );
NOR4_X2 U14765 ( .A1(n18686), .A2(n15736), .A3(n15737), .A4(n15738), .ZN(n15735) );
NOR2_X2 U14766 ( .A1(n15739), .A2(n17918), .ZN(n15738) );
NOR4_X2 U14767 ( .A1(n18685), .A2(n15755), .A3(n15756), .A4(n15757), .ZN(n15754) );
NOR2_X2 U14768 ( .A1(n15758), .A2(n17918), .ZN(n15757) );
NOR4_X2 U14769 ( .A1(n18684), .A2(n15774), .A3(n15775), .A4(n15776), .ZN(n15773) );
NOR2_X2 U14770 ( .A1(n15777), .A2(n17917), .ZN(n15776) );
NOR4_X2 U14771 ( .A1(n18683), .A2(n15793), .A3(n15794), .A4(n15795), .ZN(n15792) );
NOR2_X2 U14772 ( .A1(n15796), .A2(n17917), .ZN(n15795) );
NOR4_X2 U14773 ( .A1(n18674), .A2(n15960), .A3(n15961), .A4(n15962), .ZN(n15959) );
NOR2_X2 U14774 ( .A1(n15963), .A2(n17917), .ZN(n15962) );
NOR4_X2 U14775 ( .A1(n18673), .A2(n15977), .A3(n15978), .A4(n15979), .ZN(n15976) );
NOR2_X2 U14776 ( .A1(n15980), .A2(n17917), .ZN(n15979) );
NOR4_X2 U14777 ( .A1(n18672), .A2(n15994), .A3(n15995), .A4(n15996), .ZN(n15993) );
NOR2_X2 U14778 ( .A1(n15997), .A2(n17917), .ZN(n15996) );
NOR4_X2 U14779 ( .A1(n18671), .A2(n16011), .A3(n16012), .A4(n16013), .ZN(n16010) );
NOR2_X2 U14780 ( .A1(n16014), .A2(n17917), .ZN(n16013) );
NOR4_X2 U14781 ( .A1(n18670), .A2(n16028), .A3(n16029), .A4(n16030), .ZN(n16027) );
NOR2_X2 U14782 ( .A1(n16031), .A2(n17917), .ZN(n16030) );
NOR4_X2 U14783 ( .A1(n18669), .A2(n16045), .A3(n16046), .A4(n16047), .ZN(n16044) );
NOR2_X2 U14784 ( .A1(n16048), .A2(n17917), .ZN(n16047) );
NOR4_X2 U14785 ( .A1(n18668), .A2(n16062), .A3(n16063), .A4(n16064), .ZN(n16061) );
NOR2_X2 U14786 ( .A1(n16065), .A2(n17917), .ZN(n16064) );
NOR4_X2 U14787 ( .A1(n18667), .A2(n16079), .A3(n16080), .A4(n16081), .ZN(n16078) );
NOR2_X2 U14788 ( .A1(n16082), .A2(n17917), .ZN(n16081) );
NOR2_X2 U14789 ( .A1(n13802), .A2(n15117), .ZN(n15115) );
NOR2_X2 U14790 ( .A1(n13796), .A2(n15117), .ZN(n15138) );
NOR2_X2 U14791 ( .A1(n13790), .A2(n15117), .ZN(n15160) );
NOR2_X2 U14792 ( .A1(n13784), .A2(n15117), .ZN(n15182) );
NOR2_X2 U14793 ( .A1(n13778), .A2(n15117), .ZN(n15204) );
NOR2_X2 U14794 ( .A1(n13772), .A2(n15117), .ZN(n15226) );
NOR2_X2 U14795 ( .A1(n13766), .A2(n15117), .ZN(n15248) );
NOR2_X2 U14796 ( .A1(n13760), .A2(n15117), .ZN(n15270) );
NOR2_X2 U14797 ( .A1(n13898), .A2(n14758), .ZN(n14756) );
NOR2_X2 U14798 ( .A1(n13892), .A2(n14758), .ZN(n14780) );
NOR2_X2 U14799 ( .A1(n13886), .A2(n14758), .ZN(n14802) );
NOR2_X2 U14800 ( .A1(n13880), .A2(n14758), .ZN(n14824) );
NOR2_X2 U14801 ( .A1(n13874), .A2(n14758), .ZN(n14846) );
NOR2_X2 U14802 ( .A1(n13868), .A2(n14758), .ZN(n14868) );
NOR2_X2 U14803 ( .A1(n13862), .A2(n14758), .ZN(n14890) );
NOR2_X2 U14804 ( .A1(n13856), .A2(n14758), .ZN(n14912) );
NOR2_X2 U14805 ( .A1(n13754), .A2(n15296), .ZN(n15294) );
NOR2_X2 U14806 ( .A1(n13748), .A2(n15296), .ZN(n15320) );
NOR2_X2 U14807 ( .A1(n13742), .A2(n15296), .ZN(n15344) );
NOR2_X2 U14808 ( .A1(n13736), .A2(n15296), .ZN(n15368) );
NOR2_X2 U14809 ( .A1(n13730), .A2(n15296), .ZN(n15392) );
NOR2_X2 U14810 ( .A1(n13724), .A2(n15296), .ZN(n15416) );
NOR2_X2 U14811 ( .A1(n13718), .A2(n15296), .ZN(n15440) );
NOR2_X2 U14812 ( .A1(n13712), .A2(n15296), .ZN(n15464) );
NOR2_X2 U14813 ( .A1(n13706), .A2(n15492), .ZN(n15489) );
NOR2_X2 U14814 ( .A1(n13700), .A2(n15492), .ZN(n15518) );
NOR2_X2 U14815 ( .A1(n13694), .A2(n15492), .ZN(n15539) );
NOR2_X2 U14816 ( .A1(n13688), .A2(n15492), .ZN(n15560) );
NOR2_X2 U14817 ( .A1(n13682), .A2(n15492), .ZN(n15581) );
NOR2_X2 U14818 ( .A1(n13946), .A2(n14587), .ZN(n14585) );
NOR2_X2 U14819 ( .A1(n13940), .A2(n14587), .ZN(n14607) );
NOR2_X2 U14820 ( .A1(n13934), .A2(n14587), .ZN(n14628) );
NOR2_X2 U14821 ( .A1(n13928), .A2(n14587), .ZN(n14649) );
NOR2_X2 U14822 ( .A1(n13922), .A2(n14587), .ZN(n14670) );
NOR2_X2 U14823 ( .A1(n13916), .A2(n14587), .ZN(n14691) );
NOR2_X2 U14824 ( .A1(n13910), .A2(n14587), .ZN(n14712) );
NOR2_X2 U14825 ( .A1(n13904), .A2(n14587), .ZN(n14733) );
NOR2_X2 U14826 ( .A1(n13850), .A2(n14937), .ZN(n14935) );
NOR2_X2 U14827 ( .A1(n13844), .A2(n14937), .ZN(n14959) );
NOR2_X2 U14828 ( .A1(n13838), .A2(n14937), .ZN(n14981) );
NOR2_X2 U14829 ( .A1(n13832), .A2(n14937), .ZN(n15003) );
NOR2_X2 U14830 ( .A1(n13826), .A2(n14937), .ZN(n15025) );
NOR2_X2 U14831 ( .A1(n13820), .A2(n14937), .ZN(n15047) );
NOR2_X2 U14832 ( .A1(n13814), .A2(n14937), .ZN(n15069) );
NOR2_X2 U14833 ( .A1(n13808), .A2(n14937), .ZN(n15091) );
NOR2_X2 U14834 ( .A1(n13994), .A2(n14406), .ZN(n14404) );
NOR2_X2 U14835 ( .A1(n13988), .A2(n14406), .ZN(n14429) );
NOR2_X2 U14836 ( .A1(n13982), .A2(n14406), .ZN(n14451) );
NOR2_X2 U14837 ( .A1(n13976), .A2(n14406), .ZN(n14473) );
NOR2_X2 U14838 ( .A1(n13970), .A2(n14406), .ZN(n14495) );
NOR2_X2 U14839 ( .A1(n13964), .A2(n14406), .ZN(n14517) );
NOR2_X2 U14840 ( .A1(n13958), .A2(n14406), .ZN(n14539) );
NOR2_X2 U14841 ( .A1(n13952), .A2(n14406), .ZN(n14561) );
NOR2_X2 U14842 ( .A1(n13676), .A2(n15492), .ZN(n15602) );
NOR2_X2 U14843 ( .A1(n13669), .A2(n15492), .ZN(n15621) );
NOR2_X2 U14844 ( .A1(n13662), .A2(n15492), .ZN(n15640) );
NOR2_X2 U14845 ( .A1(n16209), .A2(n13462), .ZN(n16221) );
NOR2_X2 U14846 ( .A1(n16209), .A2(n13456), .ZN(n16235) );
NOR2_X2 U14847 ( .A1(n16209), .A2(n13450), .ZN(n16249) );
NOR2_X2 U14848 ( .A1(n16209), .A2(n13444), .ZN(n16263) );
NOR2_X2 U14849 ( .A1(n16209), .A2(n13438), .ZN(n16277) );
NOR2_X2 U14850 ( .A1(n16209), .A2(n13432), .ZN(n16291) );
NOR2_X2 U14851 ( .A1(n16209), .A2(n13426), .ZN(n16305) );
NOR2_X2 U14852 ( .A1(n16209), .A2(n13420), .ZN(n16319) );
NOR2_X2 U14853 ( .A1(n15663), .A2(n13654), .ZN(n15660) );
NOR2_X2 U14854 ( .A1(n15663), .A2(n13648), .ZN(n15680) );
NOR2_X2 U14855 ( .A1(n15663), .A2(n13642), .ZN(n15699) );
NOR2_X2 U14856 ( .A1(n15663), .A2(n13636), .ZN(n15718) );
NOR2_X2 U14857 ( .A1(n15663), .A2(n13630), .ZN(n15737) );
NOR2_X2 U14858 ( .A1(n15663), .A2(n13624), .ZN(n15756) );
NOR2_X2 U14859 ( .A1(n15663), .A2(n13618), .ZN(n15775) );
NOR2_X2 U14860 ( .A1(n15663), .A2(n13612), .ZN(n15794) );
NOR2_X2 U14861 ( .A1(n13558), .A2(n15946), .ZN(n15961) );
NOR2_X2 U14862 ( .A1(n13552), .A2(n15946), .ZN(n15978) );
NOR2_X2 U14863 ( .A1(n13546), .A2(n15946), .ZN(n15995) );
NOR2_X2 U14864 ( .A1(n13540), .A2(n15946), .ZN(n16012) );
NOR2_X2 U14865 ( .A1(n13534), .A2(n15946), .ZN(n16029) );
NOR2_X2 U14866 ( .A1(n13528), .A2(n15946), .ZN(n16046) );
NOR2_X2 U14867 ( .A1(n13522), .A2(n15946), .ZN(n16063) );
NOR2_X2 U14868 ( .A1(n13516), .A2(n15946), .ZN(n16080) );
AND2_X2 U14869 ( .A1(n17892), .A2(n15309), .ZN(n17756) );
NOR2_X2 U14870 ( .A1(n19191), .A2(n17905), .ZN(n16546) );
NOR2_X2 U14871 ( .A1(n19192), .A2(n17905), .ZN(n16551) );
NOR2_X2 U14872 ( .A1(n19193), .A2(n17905), .ZN(n16556) );
NOR2_X2 U14873 ( .A1(n19194), .A2(n17905), .ZN(n16561) );
NOR2_X2 U14874 ( .A1(n19195), .A2(n17905), .ZN(n16566) );
INV_X4 U14875 ( .A(n14414), .ZN(n17891) );
NOR2_X2 U14876 ( .A1(n18037), .A2(n16436), .ZN(N3086) );
NAND3_X2 U14877 ( .A1(n16438), .A2(n16439), .A3(n16440), .ZN(n16437) );
NOR2_X2 U14878 ( .A1(n18037), .A2(n16451), .ZN(N3085) );
NAND3_X2 U14879 ( .A1(n16453), .A2(n16454), .A3(n16455), .ZN(n16452) );
NOR2_X2 U14880 ( .A1(n18037), .A2(n16464), .ZN(N3084) );
NAND3_X2 U14881 ( .A1(n16466), .A2(n16467), .A3(n16468), .ZN(n16465) );
NOR2_X2 U14882 ( .A1(n18036), .A2(n16477), .ZN(N3083) );
NAND3_X2 U14883 ( .A1(n16479), .A2(n16480), .A3(n16481), .ZN(n16478) );
NOR2_X2 U14884 ( .A1(n18036), .A2(n16490), .ZN(N3082) );
NAND3_X2 U14885 ( .A1(n16492), .A2(n16493), .A3(n16494), .ZN(n16491) );
NOR2_X2 U14886 ( .A1(n18036), .A2(n16503), .ZN(N3081) );
NAND3_X2 U14887 ( .A1(n16505), .A2(n16506), .A3(n16507), .ZN(n16504) );
NOR2_X2 U14888 ( .A1(n18036), .A2(n16516), .ZN(N3080) );
NAND3_X2 U14889 ( .A1(n16518), .A2(n16519), .A3(n16520), .ZN(n16517) );
NOR2_X2 U14890 ( .A1(n18036), .A2(n16529), .ZN(N3079) );
NAND3_X2 U14891 ( .A1(n16531), .A2(n16532), .A3(n16533), .ZN(n16530) );
NOR2_X2 U14892 ( .A1(n19203), .A2(n11946), .ZN(n14167) );
NOR2_X2 U14893 ( .A1(n18075), .A2(n18071), .ZN(n14422) );
INV_X4 U14894 ( .A(n17775), .ZN(n17897) );
NOR4_X2 U14895 ( .A1(n14180), .A2(n14181), .A3(n14182), .A4(n14183), .ZN(n14179) );
NOR2_X2 U14896 ( .A1(n19135), .A2(n17860), .ZN(n14183) );
NOR2_X2 U14897 ( .A1(n19143), .A2(n14187), .ZN(n14180) );
NOR2_X2 U14898 ( .A1(n14185), .A2(n14186), .ZN(n14181) );
NOR4_X2 U14899 ( .A1(n14212), .A2(n14213), .A3(n14214), .A4(n14215), .ZN(n14211) );
NOR2_X2 U14900 ( .A1(n19136), .A2(n17860), .ZN(n14215) );
NOR2_X2 U14901 ( .A1(n19144), .A2(n14187), .ZN(n14212) );
NOR2_X2 U14902 ( .A1(n14216), .A2(n14186), .ZN(n14213) );
NOR4_X2 U14903 ( .A1(n14241), .A2(n14242), .A3(n14243), .A4(n14244), .ZN(n14240) );
NOR2_X2 U14904 ( .A1(n19137), .A2(n17860), .ZN(n14244) );
NOR2_X2 U14905 ( .A1(n19145), .A2(n14187), .ZN(n14241) );
NOR2_X2 U14906 ( .A1(n14245), .A2(n14186), .ZN(n14242) );
NOR4_X2 U14907 ( .A1(n14270), .A2(n14271), .A3(n14272), .A4(n14273), .ZN(n14269) );
NOR2_X2 U14908 ( .A1(n19138), .A2(n17860), .ZN(n14273) );
NOR2_X2 U14909 ( .A1(n19146), .A2(n14187), .ZN(n14270) );
NOR2_X2 U14910 ( .A1(n14274), .A2(n14186), .ZN(n14271) );
NOR4_X2 U14911 ( .A1(n14299), .A2(n14300), .A3(n14301), .A4(n14302), .ZN(n14298) );
NOR2_X2 U14912 ( .A1(n19139), .A2(n17860), .ZN(n14302) );
NOR2_X2 U14913 ( .A1(n19147), .A2(n14187), .ZN(n14299) );
NOR2_X2 U14914 ( .A1(n14303), .A2(n14186), .ZN(n14300) );
NOR4_X2 U14915 ( .A1(n14328), .A2(n14329), .A3(n14330), .A4(n14331), .ZN(n14327) );
NOR2_X2 U14916 ( .A1(n19140), .A2(n17860), .ZN(n14331) );
NOR2_X2 U14917 ( .A1(n19148), .A2(n14187), .ZN(n14328) );
NOR2_X2 U14918 ( .A1(n14332), .A2(n14186), .ZN(n14329) );
NOR4_X2 U14919 ( .A1(n14357), .A2(n14358), .A3(n14359), .A4(n14360), .ZN(n14356) );
NOR2_X2 U14920 ( .A1(n19141), .A2(n17860), .ZN(n14360) );
NOR2_X2 U14921 ( .A1(n19149), .A2(n14187), .ZN(n14357) );
NOR2_X2 U14922 ( .A1(n14361), .A2(n14186), .ZN(n14358) );
NOR4_X2 U14923 ( .A1(n14386), .A2(n14387), .A3(n14388), .A4(n14389), .ZN(n14385) );
NOR2_X2 U14924 ( .A1(n19142), .A2(n17860), .ZN(n14389) );
NOR2_X2 U14925 ( .A1(n19150), .A2(n14187), .ZN(n14386) );
NOR2_X2 U14926 ( .A1(n14391), .A2(n14186), .ZN(n14387) );
NOR4_X2 U14927 ( .A1(n15610), .A2(n15611), .A3(n15612), .A4(n15613), .ZN(n15609) );
NOR2_X2 U14928 ( .A1(n19148), .A2(n15507), .ZN(n15610) );
NOR2_X2 U14929 ( .A1(n19156), .A2(n15508), .ZN(n15611) );
NOR2_X2 U14930 ( .A1(n19180), .A2(n17869), .ZN(n15612) );
NOR4_X2 U14931 ( .A1(n15629), .A2(n15630), .A3(n15631), .A4(n15632), .ZN(n15628) );
NOR2_X2 U14932 ( .A1(n19149), .A2(n15507), .ZN(n15629) );
NOR2_X2 U14933 ( .A1(n19157), .A2(n15508), .ZN(n15630) );
NOR2_X2 U14934 ( .A1(n19181), .A2(n17869), .ZN(n15631) );
NOR4_X2 U14935 ( .A1(n15649), .A2(n15650), .A3(n15651), .A4(n15652), .ZN(n15648) );
NOR2_X2 U14936 ( .A1(n19150), .A2(n15507), .ZN(n15649) );
NOR2_X2 U14937 ( .A1(n19158), .A2(n15508), .ZN(n15650) );
NOR2_X2 U14938 ( .A1(n19182), .A2(n17869), .ZN(n15651) );
NOR4_X2 U14939 ( .A1(n15668), .A2(n15669), .A3(n15670), .A4(n15671), .ZN(n15667) );
NOR2_X2 U14940 ( .A1(n19191), .A2(n15504), .ZN(n15668) );
NOR2_X2 U14941 ( .A1(n19183), .A2(n17869), .ZN(n15669) );
NOR2_X2 U14942 ( .A1(n19175), .A2(n17870), .ZN(n15670) );
NOR4_X2 U14943 ( .A1(n15687), .A2(n15688), .A3(n15689), .A4(n15690), .ZN(n15686) );
NOR2_X2 U14944 ( .A1(n19192), .A2(n15504), .ZN(n15687) );
NOR2_X2 U14945 ( .A1(n19184), .A2(n17869), .ZN(n15688) );
NOR2_X2 U14946 ( .A1(n19176), .A2(n17870), .ZN(n15689) );
NOR4_X2 U14947 ( .A1(n15706), .A2(n15707), .A3(n15708), .A4(n15709), .ZN(n15705) );
NOR2_X2 U14948 ( .A1(n19193), .A2(n15504), .ZN(n15706) );
NOR2_X2 U14949 ( .A1(n19185), .A2(n17869), .ZN(n15707) );
NOR2_X2 U14950 ( .A1(n19177), .A2(n17870), .ZN(n15708) );
NOR4_X2 U14951 ( .A1(n15725), .A2(n15726), .A3(n15727), .A4(n15728), .ZN(n15724) );
NOR2_X2 U14952 ( .A1(n19194), .A2(n15504), .ZN(n15725) );
NOR2_X2 U14953 ( .A1(n19186), .A2(n17869), .ZN(n15726) );
NOR2_X2 U14954 ( .A1(n19178), .A2(n17870), .ZN(n15727) );
NOR4_X2 U14955 ( .A1(n15744), .A2(n15745), .A3(n15746), .A4(n15747), .ZN(n15743) );
NOR2_X2 U14956 ( .A1(n19195), .A2(n15504), .ZN(n15744) );
NOR2_X2 U14957 ( .A1(n19187), .A2(n17868), .ZN(n15745) );
NOR2_X2 U14958 ( .A1(n19179), .A2(n17870), .ZN(n15746) );
NOR4_X2 U14959 ( .A1(n15763), .A2(n15764), .A3(n15765), .A4(n15766), .ZN(n15762) );
NOR2_X2 U14960 ( .A1(n19196), .A2(n15504), .ZN(n15763) );
NOR2_X2 U14961 ( .A1(n19188), .A2(n17868), .ZN(n15764) );
NOR2_X2 U14962 ( .A1(n19180), .A2(n17871), .ZN(n15765) );
NOR4_X2 U14963 ( .A1(n15782), .A2(n15783), .A3(n15784), .A4(n15785), .ZN(n15781) );
NOR2_X2 U14964 ( .A1(n19197), .A2(n15504), .ZN(n15782) );
NOR2_X2 U14965 ( .A1(n19189), .A2(n17868), .ZN(n15783) );
NOR2_X2 U14966 ( .A1(n19181), .A2(n17871), .ZN(n15784) );
NOR4_X2 U14967 ( .A1(n15801), .A2(n15802), .A3(n15803), .A4(n15804), .ZN(n15800) );
NOR2_X2 U14968 ( .A1(n19198), .A2(n15504), .ZN(n15801) );
NOR2_X2 U14969 ( .A1(n19190), .A2(n17868), .ZN(n15802) );
NOR2_X2 U14970 ( .A1(n19182), .A2(n17871), .ZN(n15803) );
NOR4_X2 U14971 ( .A1(n15497), .A2(n15498), .A3(n15499), .A4(n15500), .ZN(n15496) );
NOR2_X2 U14972 ( .A1(n19183), .A2(n15504), .ZN(n15497) );
NOR2_X2 U14973 ( .A1(n19175), .A2(n17869), .ZN(n15498) );
NOR2_X2 U14974 ( .A1(n19167), .A2(n17871), .ZN(n15499) );
NOR4_X2 U14975 ( .A1(n15525), .A2(n15526), .A3(n15527), .A4(n15528), .ZN(n15524) );
NOR2_X2 U14976 ( .A1(n19184), .A2(n15504), .ZN(n15525) );
NOR2_X2 U14977 ( .A1(n19176), .A2(n17869), .ZN(n15526) );
NOR2_X2 U14978 ( .A1(n19168), .A2(n17870), .ZN(n15527) );
NOR4_X2 U14979 ( .A1(n15546), .A2(n15547), .A3(n15548), .A4(n15549), .ZN(n15545) );
NOR2_X2 U14980 ( .A1(n19185), .A2(n15504), .ZN(n15546) );
NOR2_X2 U14981 ( .A1(n19177), .A2(n17869), .ZN(n15547) );
NOR2_X2 U14982 ( .A1(n19169), .A2(n17870), .ZN(n15548) );
NOR4_X2 U14983 ( .A1(n15567), .A2(n15568), .A3(n15569), .A4(n15570), .ZN(n15566) );
NOR2_X2 U14984 ( .A1(n19186), .A2(n15504), .ZN(n15567) );
NOR2_X2 U14985 ( .A1(n19178), .A2(n17869), .ZN(n15568) );
NOR2_X2 U14986 ( .A1(n19170), .A2(n17870), .ZN(n15569) );
NOR4_X2 U14987 ( .A1(n15588), .A2(n15589), .A3(n15590), .A4(n15591), .ZN(n15587) );
NOR2_X2 U14988 ( .A1(n19187), .A2(n15504), .ZN(n15588) );
NOR2_X2 U14989 ( .A1(n19179), .A2(n17869), .ZN(n15589) );
NOR2_X2 U14990 ( .A1(n19171), .A2(n17870), .ZN(n15590) );
NAND3_X2 U14991 ( .A1(n14418), .A2(n14419), .A3(n14420), .ZN(n14190) );
NAND3_X2 U14992 ( .A1(n14441), .A2(n14442), .A3(n14443), .ZN(n14219) );
NAND3_X2 U14993 ( .A1(n14463), .A2(n14464), .A3(n14465), .ZN(n14248) );
NAND3_X2 U14994 ( .A1(n14485), .A2(n14486), .A3(n14487), .ZN(n14277) );
NAND3_X2 U14995 ( .A1(n14507), .A2(n14508), .A3(n14509), .ZN(n14306) );
NAND3_X2 U14996 ( .A1(n14529), .A2(n14530), .A3(n14531), .ZN(n14335) );
NAND3_X2 U14997 ( .A1(n14551), .A2(n14552), .A3(n14553), .ZN(n14364) );
NAND3_X2 U14998 ( .A1(n14575), .A2(n14576), .A3(n14577), .ZN(n14396) );
NOR2_X2 U14999 ( .A1(n19167), .A2(n14184), .ZN(n14182) );
NOR2_X2 U15000 ( .A1(n19168), .A2(n14184), .ZN(n14214) );
NOR2_X2 U15001 ( .A1(n19169), .A2(n14184), .ZN(n14243) );
NOR2_X2 U15002 ( .A1(n19170), .A2(n14184), .ZN(n14272) );
NOR2_X2 U15003 ( .A1(n19171), .A2(n14184), .ZN(n14301) );
NOR2_X2 U15004 ( .A1(n19172), .A2(n14184), .ZN(n14330) );
NOR2_X2 U15005 ( .A1(n19173), .A2(n14184), .ZN(n14359) );
NOR2_X2 U15006 ( .A1(n19174), .A2(n14184), .ZN(n14388) );
INV_X4 U15007 ( .A(n18075), .ZN(n18074) );
NOR2_X2 U15008 ( .A1(n19159), .A2(n17875), .ZN(n15500) );
NOR2_X2 U15009 ( .A1(n19160), .A2(n17874), .ZN(n15528) );
NOR2_X2 U15010 ( .A1(n19161), .A2(n17874), .ZN(n15549) );
NOR2_X2 U15011 ( .A1(n19162), .A2(n17874), .ZN(n15570) );
NOR2_X2 U15012 ( .A1(n19163), .A2(n17874), .ZN(n15591) );
NOR2_X2 U15013 ( .A1(n19164), .A2(n17874), .ZN(n15613) );
NOR2_X2 U15014 ( .A1(n19165), .A2(n17874), .ZN(n15632) );
NOR2_X2 U15015 ( .A1(n19166), .A2(n17874), .ZN(n15652) );
NOR2_X2 U15016 ( .A1(n19167), .A2(n17874), .ZN(n15671) );
NOR2_X2 U15017 ( .A1(n19168), .A2(n17874), .ZN(n15690) );
NOR2_X2 U15018 ( .A1(n19169), .A2(n17874), .ZN(n15709) );
NOR2_X2 U15019 ( .A1(n19170), .A2(n17874), .ZN(n15728) );
NOR2_X2 U15020 ( .A1(n19171), .A2(n17875), .ZN(n15747) );
NOR2_X2 U15021 ( .A1(n19172), .A2(n17875), .ZN(n15766) );
NOR2_X2 U15022 ( .A1(n19173), .A2(n17875), .ZN(n15785) );
NOR2_X2 U15023 ( .A1(n19174), .A2(n17875), .ZN(n15804) );
NAND2_X2 U15024 ( .A1(n14564), .A2(n15309), .ZN(n15504) );
NOR3_X2 U15025 ( .A1(n15915), .A2(n15916), .A3(n15917), .ZN(n15914) );
NOR2_X2 U15026 ( .A1(n19188), .A2(n17871), .ZN(n15917) );
NOR2_X2 U15027 ( .A1(n19196), .A2(n17868), .ZN(n15916) );
NOR2_X2 U15028 ( .A1(n19180), .A2(n17875), .ZN(n15915) );
NOR3_X2 U15029 ( .A1(n15825), .A2(n15826), .A3(n15827), .ZN(n15824) );
NOR2_X2 U15030 ( .A1(n19183), .A2(n17871), .ZN(n15827) );
NOR2_X2 U15031 ( .A1(n19191), .A2(n17868), .ZN(n15826) );
NOR2_X2 U15032 ( .A1(n19175), .A2(n17875), .ZN(n15825) );
NOR3_X2 U15033 ( .A1(n15843), .A2(n15844), .A3(n15845), .ZN(n15842) );
NOR2_X2 U15034 ( .A1(n19184), .A2(n17871), .ZN(n15845) );
NOR2_X2 U15035 ( .A1(n19192), .A2(n17868), .ZN(n15844) );
NOR2_X2 U15036 ( .A1(n19176), .A2(n17875), .ZN(n15843) );
NOR3_X2 U15037 ( .A1(n15861), .A2(n15862), .A3(n15863), .ZN(n15860) );
NOR2_X2 U15038 ( .A1(n19185), .A2(n17871), .ZN(n15863) );
NOR2_X2 U15039 ( .A1(n19193), .A2(n17868), .ZN(n15862) );
NOR2_X2 U15040 ( .A1(n19177), .A2(n17875), .ZN(n15861) );
NOR3_X2 U15041 ( .A1(n15879), .A2(n15880), .A3(n15881), .ZN(n15878) );
NOR2_X2 U15042 ( .A1(n19186), .A2(n17871), .ZN(n15881) );
NOR2_X2 U15043 ( .A1(n19194), .A2(n17868), .ZN(n15880) );
NOR2_X2 U15044 ( .A1(n19178), .A2(n17875), .ZN(n15879) );
NOR3_X2 U15045 ( .A1(n15897), .A2(n15898), .A3(n15899), .ZN(n15896) );
NOR2_X2 U15046 ( .A1(n19187), .A2(n17871), .ZN(n15899) );
NOR2_X2 U15047 ( .A1(n19195), .A2(n17868), .ZN(n15898) );
NOR2_X2 U15048 ( .A1(n19179), .A2(n17875), .ZN(n15897) );
NOR3_X2 U15049 ( .A1(n15933), .A2(n15934), .A3(n15935), .ZN(n15932) );
NOR2_X2 U15050 ( .A1(n19189), .A2(n17871), .ZN(n15935) );
NOR2_X2 U15051 ( .A1(n19197), .A2(n17868), .ZN(n15934) );
NOR2_X2 U15052 ( .A1(n19181), .A2(n17875), .ZN(n15933) );
NOR3_X2 U15053 ( .A1(n15953), .A2(n15954), .A3(n15955), .ZN(n15952) );
NOR2_X2 U15054 ( .A1(n19190), .A2(n17871), .ZN(n15955) );
NOR2_X2 U15055 ( .A1(n19198), .A2(n17868), .ZN(n15954) );
NOR2_X2 U15056 ( .A1(n19182), .A2(n17876), .ZN(n15953) );
NOR3_X2 U15057 ( .A1(n15304), .A2(n15305), .A3(n15306), .ZN(n15303) );
NOR2_X2 U15058 ( .A1(n15127), .A2(n17891), .ZN(n15304) );
NOR2_X2 U15059 ( .A1(n19183), .A2(n17864), .ZN(n15306) );
NOR2_X2 U15060 ( .A1(n19151), .A2(n17878), .ZN(n15305) );
NOR3_X2 U15061 ( .A1(n15329), .A2(n15330), .A3(n15331), .ZN(n15328) );
NOR2_X2 U15062 ( .A1(n15149), .A2(n17891), .ZN(n15329) );
NOR2_X2 U15063 ( .A1(n19184), .A2(n17864), .ZN(n15331) );
NOR2_X2 U15064 ( .A1(n19152), .A2(n17878), .ZN(n15330) );
NOR3_X2 U15065 ( .A1(n15353), .A2(n15354), .A3(n15355), .ZN(n15352) );
NOR2_X2 U15066 ( .A1(n15171), .A2(n17891), .ZN(n15353) );
NOR2_X2 U15067 ( .A1(n19185), .A2(n17864), .ZN(n15355) );
NOR2_X2 U15068 ( .A1(n19153), .A2(n17878), .ZN(n15354) );
NOR3_X2 U15069 ( .A1(n15377), .A2(n15378), .A3(n15379), .ZN(n15376) );
NOR2_X2 U15070 ( .A1(n15193), .A2(n17891), .ZN(n15377) );
NOR2_X2 U15071 ( .A1(n19186), .A2(n17864), .ZN(n15379) );
NOR2_X2 U15072 ( .A1(n19154), .A2(n17878), .ZN(n15378) );
NOR3_X2 U15073 ( .A1(n15401), .A2(n15402), .A3(n15403), .ZN(n15400) );
NOR2_X2 U15074 ( .A1(n15215), .A2(n17891), .ZN(n15401) );
NOR2_X2 U15075 ( .A1(n19187), .A2(n17864), .ZN(n15403) );
NOR2_X2 U15076 ( .A1(n19155), .A2(n17878), .ZN(n15402) );
NOR3_X2 U15077 ( .A1(n15425), .A2(n15426), .A3(n15427), .ZN(n15424) );
NOR2_X2 U15078 ( .A1(n15237), .A2(n17891), .ZN(n15425) );
NOR2_X2 U15079 ( .A1(n19188), .A2(n17864), .ZN(n15427) );
NOR2_X2 U15080 ( .A1(n19156), .A2(n17878), .ZN(n15426) );
NOR3_X2 U15081 ( .A1(n15449), .A2(n15450), .A3(n15451), .ZN(n15448) );
NOR2_X2 U15082 ( .A1(n15259), .A2(n17891), .ZN(n15449) );
NOR2_X2 U15083 ( .A1(n19189), .A2(n17864), .ZN(n15451) );
NOR2_X2 U15084 ( .A1(n19157), .A2(n17878), .ZN(n15450) );
NOR3_X2 U15085 ( .A1(n15475), .A2(n15476), .A3(n15477), .ZN(n15474) );
NOR2_X2 U15086 ( .A1(n15283), .A2(n17891), .ZN(n15475) );
NOR2_X2 U15087 ( .A1(n19190), .A2(n17864), .ZN(n15477) );
NOR2_X2 U15088 ( .A1(n19158), .A2(n17878), .ZN(n15476) );
NOR2_X2 U15089 ( .A1(n19143), .A2(n17879), .ZN(n15125) );
NOR2_X2 U15090 ( .A1(n19144), .A2(n17879), .ZN(n15147) );
NOR2_X2 U15091 ( .A1(n19145), .A2(n17879), .ZN(n15169) );
NOR2_X2 U15092 ( .A1(n19146), .A2(n17879), .ZN(n15191) );
NOR2_X2 U15093 ( .A1(n19147), .A2(n17878), .ZN(n15213) );
NOR2_X2 U15094 ( .A1(n19148), .A2(n17878), .ZN(n15235) );
NOR2_X2 U15095 ( .A1(n19149), .A2(n17878), .ZN(n15257) );
NOR2_X2 U15096 ( .A1(n19150), .A2(n17878), .ZN(n15281) );
NOR2_X2 U15097 ( .A1(n15127), .A2(n17865), .ZN(n15124) );
NOR2_X2 U15098 ( .A1(n15149), .A2(n17865), .ZN(n15146) );
NOR2_X2 U15099 ( .A1(n15171), .A2(n17865), .ZN(n15168) );
NOR2_X2 U15100 ( .A1(n15193), .A2(n17865), .ZN(n15190) );
NOR2_X2 U15101 ( .A1(n15215), .A2(n17865), .ZN(n15212) );
NOR2_X2 U15102 ( .A1(n15237), .A2(n17865), .ZN(n15234) );
NOR2_X2 U15103 ( .A1(n15259), .A2(n17865), .ZN(n15256) );
NOR2_X2 U15104 ( .A1(n15283), .A2(n17865), .ZN(n15280) );
NOR2_X2 U15105 ( .A1(n19175), .A2(n17863), .ZN(n15126) );
NOR2_X2 U15106 ( .A1(n19176), .A2(n17863), .ZN(n15148) );
NOR2_X2 U15107 ( .A1(n19177), .A2(n17863), .ZN(n15170) );
NOR2_X2 U15108 ( .A1(n19178), .A2(n17863), .ZN(n15192) );
NOR2_X2 U15109 ( .A1(n19179), .A2(n17863), .ZN(n15214) );
NOR2_X2 U15110 ( .A1(n19180), .A2(n17863), .ZN(n15236) );
NOR2_X2 U15111 ( .A1(n19181), .A2(n17863), .ZN(n15258) );
NOR2_X2 U15112 ( .A1(n19182), .A2(n17863), .ZN(n15282) );
NOR2_X2 U15113 ( .A1(n19151), .A2(n15508), .ZN(n15505) );
NOR2_X2 U15114 ( .A1(n19152), .A2(n15508), .ZN(n15529) );
NOR2_X2 U15115 ( .A1(n19153), .A2(n15508), .ZN(n15550) );
NOR2_X2 U15116 ( .A1(n19154), .A2(n15508), .ZN(n15571) );
NOR2_X2 U15117 ( .A1(n19155), .A2(n15508), .ZN(n15592) );
NOR2_X2 U15118 ( .A1(n19196), .A2(n17864), .ZN(n15615) );
AND2_X2 U15119 ( .A1(n18071), .A2(n18075), .ZN(n17757) );
AND2_X2 U15120 ( .A1(n17897), .A2(n15309), .ZN(n17758) );
NOR2_X2 U15121 ( .A1(n19143), .A2(n15507), .ZN(n15506) );
NOR2_X2 U15122 ( .A1(n19144), .A2(n15507), .ZN(n15530) );
NOR2_X2 U15123 ( .A1(n19145), .A2(n15507), .ZN(n15551) );
NOR2_X2 U15124 ( .A1(n19146), .A2(n15507), .ZN(n15572) );
NOR2_X2 U15125 ( .A1(n19147), .A2(n15507), .ZN(n15593) );
NOR2_X2 U15126 ( .A1(n14415), .A2(n14416), .ZN(n14412) );
NOR2_X2 U15127 ( .A1(n17866), .A2(n14417), .ZN(n14416) );
NOR2_X2 U15128 ( .A1(n19143), .A2(n17860), .ZN(n14415) );
NOR2_X2 U15129 ( .A1(n14438), .A2(n14439), .ZN(n14436) );
NOR2_X2 U15130 ( .A1(n17866), .A2(n14440), .ZN(n14439) );
NOR2_X2 U15131 ( .A1(n19144), .A2(n17860), .ZN(n14438) );
NOR2_X2 U15132 ( .A1(n14460), .A2(n14461), .ZN(n14458) );
NOR2_X2 U15133 ( .A1(n17866), .A2(n14462), .ZN(n14461) );
NOR2_X2 U15134 ( .A1(n19145), .A2(n17860), .ZN(n14460) );
NOR2_X2 U15135 ( .A1(n14482), .A2(n14483), .ZN(n14480) );
NOR2_X2 U15136 ( .A1(n17866), .A2(n14484), .ZN(n14483) );
NOR2_X2 U15137 ( .A1(n19146), .A2(n17860), .ZN(n14482) );
NOR2_X2 U15138 ( .A1(n14504), .A2(n14505), .ZN(n14502) );
NOR2_X2 U15139 ( .A1(n17866), .A2(n14506), .ZN(n14505) );
NOR2_X2 U15140 ( .A1(n19147), .A2(n17861), .ZN(n14504) );
NOR2_X2 U15141 ( .A1(n14526), .A2(n14527), .ZN(n14524) );
NOR2_X2 U15142 ( .A1(n17866), .A2(n14528), .ZN(n14527) );
NOR2_X2 U15143 ( .A1(n19148), .A2(n17861), .ZN(n14526) );
NOR2_X2 U15144 ( .A1(n14548), .A2(n14549), .ZN(n14546) );
NOR2_X2 U15145 ( .A1(n17866), .A2(n14550), .ZN(n14549) );
NOR2_X2 U15146 ( .A1(n19149), .A2(n17861), .ZN(n14548) );
NOR2_X2 U15147 ( .A1(n14572), .A2(n14573), .ZN(n14570) );
NOR2_X2 U15148 ( .A1(n17866), .A2(n14574), .ZN(n14573) );
NOR2_X2 U15149 ( .A1(n19150), .A2(n17861), .ZN(n14572) );
NOR2_X2 U15150 ( .A1(n19189), .A2(n15504), .ZN(n15634) );
NOR2_X2 U15151 ( .A1(n19190), .A2(n15504), .ZN(n15654) );
NOR2_X2 U15152 ( .A1(n16088), .A2(n16089), .ZN(n16086) );
NOR2_X2 U15153 ( .A1(n19198), .A2(n17870), .ZN(n16088) );
NOR2_X2 U15154 ( .A1(n19190), .A2(n17874), .ZN(n16089) );
NOR2_X2 U15155 ( .A1(n19188), .A2(n15504), .ZN(n15614) );
NOR2_X2 U15156 ( .A1(n19173), .A2(n17870), .ZN(n15633) );
NOR2_X2 U15157 ( .A1(n19174), .A2(n17870), .ZN(n15653) );
NOR2_X2 U15158 ( .A1(n14595), .A2(n14596), .ZN(n14593) );
NOR2_X2 U15159 ( .A1(n17866), .A2(n14597), .ZN(n14596) );
NOR2_X2 U15160 ( .A1(n19151), .A2(n17861), .ZN(n14595) );
NOR2_X2 U15161 ( .A1(n14616), .A2(n14617), .ZN(n14614) );
NOR2_X2 U15162 ( .A1(n17867), .A2(n14618), .ZN(n14617) );
NOR2_X2 U15163 ( .A1(n19152), .A2(n17861), .ZN(n14616) );
NOR2_X2 U15164 ( .A1(n14637), .A2(n14638), .ZN(n14635) );
NOR2_X2 U15165 ( .A1(n17867), .A2(n14639), .ZN(n14638) );
NOR2_X2 U15166 ( .A1(n19153), .A2(n17861), .ZN(n14637) );
NOR2_X2 U15167 ( .A1(n14658), .A2(n14659), .ZN(n14656) );
NOR2_X2 U15168 ( .A1(n17867), .A2(n14660), .ZN(n14659) );
NOR2_X2 U15169 ( .A1(n19154), .A2(n17861), .ZN(n14658) );
NOR2_X2 U15170 ( .A1(n14679), .A2(n14680), .ZN(n14677) );
NOR2_X2 U15171 ( .A1(n17867), .A2(n14681), .ZN(n14680) );
NOR2_X2 U15172 ( .A1(n19155), .A2(n17861), .ZN(n14679) );
NOR2_X2 U15173 ( .A1(n14700), .A2(n14701), .ZN(n14698) );
NOR2_X2 U15174 ( .A1(n17867), .A2(n14702), .ZN(n14701) );
NOR2_X2 U15175 ( .A1(n19156), .A2(n17861), .ZN(n14700) );
NOR2_X2 U15176 ( .A1(n14721), .A2(n14722), .ZN(n14719) );
NOR2_X2 U15177 ( .A1(n17867), .A2(n14723), .ZN(n14722) );
NOR2_X2 U15178 ( .A1(n19157), .A2(n17861), .ZN(n14721) );
NOR2_X2 U15179 ( .A1(n14744), .A2(n14745), .ZN(n14742) );
NOR2_X2 U15180 ( .A1(n17867), .A2(n14746), .ZN(n14745) );
NOR2_X2 U15181 ( .A1(n19158), .A2(n17861), .ZN(n14744) );
NOR2_X2 U15182 ( .A1(n14766), .A2(n14767), .ZN(n14764) );
NOR2_X2 U15183 ( .A1(n17867), .A2(n14768), .ZN(n14767) );
NOR2_X2 U15184 ( .A1(n19159), .A2(n17862), .ZN(n14766) );
NOR2_X2 U15185 ( .A1(n14789), .A2(n14790), .ZN(n14787) );
NOR2_X2 U15186 ( .A1(n17867), .A2(n14791), .ZN(n14790) );
NOR2_X2 U15187 ( .A1(n19160), .A2(n17862), .ZN(n14789) );
NOR2_X2 U15188 ( .A1(n14811), .A2(n14812), .ZN(n14809) );
NOR2_X2 U15189 ( .A1(n17867), .A2(n14813), .ZN(n14812) );
NOR2_X2 U15190 ( .A1(n19161), .A2(n17862), .ZN(n14811) );
NOR2_X2 U15191 ( .A1(n14833), .A2(n14834), .ZN(n14831) );
NOR2_X2 U15192 ( .A1(n17867), .A2(n14835), .ZN(n14834) );
NOR2_X2 U15193 ( .A1(n19162), .A2(n17862), .ZN(n14833) );
NOR2_X2 U15194 ( .A1(n14855), .A2(n14856), .ZN(n14853) );
NOR2_X2 U15195 ( .A1(n17867), .A2(n14857), .ZN(n14856) );
NOR2_X2 U15196 ( .A1(n19163), .A2(n17862), .ZN(n14855) );
NOR2_X2 U15197 ( .A1(n14877), .A2(n14878), .ZN(n14875) );
NOR2_X2 U15198 ( .A1(n17867), .A2(n14879), .ZN(n14878) );
NOR2_X2 U15199 ( .A1(n19164), .A2(n17862), .ZN(n14877) );
NOR2_X2 U15200 ( .A1(n14899), .A2(n14900), .ZN(n14897) );
NOR2_X2 U15201 ( .A1(n17867), .A2(n14901), .ZN(n14900) );
NOR2_X2 U15202 ( .A1(n19165), .A2(n17862), .ZN(n14899) );
NOR2_X2 U15203 ( .A1(n14922), .A2(n14923), .ZN(n14920) );
NOR2_X2 U15204 ( .A1(n17866), .A2(n14924), .ZN(n14923) );
NOR2_X2 U15205 ( .A1(n19166), .A2(n17862), .ZN(n14922) );
NAND3_X2 U15206 ( .A1(n14598), .A2(n14599), .A3(n14600), .ZN(n14191) );
NAND3_X2 U15207 ( .A1(n14619), .A2(n14620), .A3(n14621), .ZN(n14220) );
NAND3_X2 U15208 ( .A1(n14640), .A2(n14641), .A3(n14642), .ZN(n14249) );
NAND3_X2 U15209 ( .A1(n14661), .A2(n14662), .A3(n14663), .ZN(n14278) );
NAND3_X2 U15210 ( .A1(n14682), .A2(n14683), .A3(n14684), .ZN(n14307) );
NAND3_X2 U15211 ( .A1(n14703), .A2(n14704), .A3(n14705), .ZN(n14336) );
NAND3_X2 U15212 ( .A1(n14724), .A2(n14725), .A3(n14726), .ZN(n14365) );
NAND3_X2 U15213 ( .A1(n14747), .A2(n14748), .A3(n14749), .ZN(n14397) );
NAND3_X2 U15214 ( .A1(n15121), .A2(n15122), .A3(n15123), .ZN(n15118) );
NOR3_X2 U15215 ( .A1(n15124), .A2(n15125), .A3(n15126), .ZN(n15123) );
NAND3_X2 U15216 ( .A1(n15143), .A2(n15144), .A3(n15145), .ZN(n15140) );
NOR3_X2 U15217 ( .A1(n15146), .A2(n15147), .A3(n15148), .ZN(n15145) );
NAND3_X2 U15218 ( .A1(n15165), .A2(n15166), .A3(n15167), .ZN(n15162) );
NOR3_X2 U15219 ( .A1(n15168), .A2(n15169), .A3(n15170), .ZN(n15167) );
NAND3_X2 U15220 ( .A1(n15187), .A2(n15188), .A3(n15189), .ZN(n15184) );
NOR3_X2 U15221 ( .A1(n15190), .A2(n15191), .A3(n15192), .ZN(n15189) );
NAND3_X2 U15222 ( .A1(n15209), .A2(n15210), .A3(n15211), .ZN(n15206) );
NOR3_X2 U15223 ( .A1(n15212), .A2(n15213), .A3(n15214), .ZN(n15211) );
NAND3_X2 U15224 ( .A1(n15231), .A2(n15232), .A3(n15233), .ZN(n15228) );
NOR3_X2 U15225 ( .A1(n15234), .A2(n15235), .A3(n15236), .ZN(n15233) );
NAND3_X2 U15226 ( .A1(n15253), .A2(n15254), .A3(n15255), .ZN(n15250) );
NOR3_X2 U15227 ( .A1(n15256), .A2(n15257), .A3(n15258), .ZN(n15255) );
NAND3_X2 U15228 ( .A1(n15277), .A2(n15278), .A3(n15279), .ZN(n15274) );
NOR3_X2 U15229 ( .A1(n15280), .A2(n15281), .A3(n15282), .ZN(n15279) );
NOR2_X2 U15230 ( .A1(n14946), .A2(n14947), .ZN(n14943) );
NOR2_X2 U15231 ( .A1(n19167), .A2(n17862), .ZN(n14947) );
NOR2_X2 U15232 ( .A1(n19135), .A2(n17879), .ZN(n14946) );
NOR2_X2 U15233 ( .A1(n14969), .A2(n14970), .ZN(n14966) );
NOR2_X2 U15234 ( .A1(n19168), .A2(n17862), .ZN(n14970) );
NOR2_X2 U15235 ( .A1(n19136), .A2(n17879), .ZN(n14969) );
NOR2_X2 U15236 ( .A1(n14991), .A2(n14992), .ZN(n14988) );
NOR2_X2 U15237 ( .A1(n19169), .A2(n17862), .ZN(n14992) );
NOR2_X2 U15238 ( .A1(n19137), .A2(n17879), .ZN(n14991) );
NOR2_X2 U15239 ( .A1(n15013), .A2(n15014), .ZN(n15010) );
NOR2_X2 U15240 ( .A1(n19170), .A2(n17862), .ZN(n15014) );
NOR2_X2 U15241 ( .A1(n19138), .A2(n17879), .ZN(n15013) );
NOR2_X2 U15242 ( .A1(n15035), .A2(n15036), .ZN(n15032) );
NOR2_X2 U15243 ( .A1(n19171), .A2(n17863), .ZN(n15036) );
NOR2_X2 U15244 ( .A1(n19139), .A2(n17879), .ZN(n15035) );
NOR2_X2 U15245 ( .A1(n15079), .A2(n15080), .ZN(n15076) );
NOR2_X2 U15246 ( .A1(n19173), .A2(n17863), .ZN(n15080) );
NOR2_X2 U15247 ( .A1(n19141), .A2(n17879), .ZN(n15079) );
NOR2_X2 U15248 ( .A1(n15103), .A2(n15104), .ZN(n15100) );
NOR2_X2 U15249 ( .A1(n19174), .A2(n17863), .ZN(n15104) );
NOR2_X2 U15250 ( .A1(n19142), .A2(n17879), .ZN(n15103) );
NOR2_X2 U15251 ( .A1(n15057), .A2(n15058), .ZN(n15054) );
NOR2_X2 U15252 ( .A1(n19172), .A2(n17863), .ZN(n15058) );
NOR2_X2 U15253 ( .A1(n19140), .A2(n17879), .ZN(n15057) );
INV_X4 U15254 ( .A(n17289), .ZN(n17958) );
NOR2_X2 U15255 ( .A1(n16053), .A2(n16054), .ZN(n16051) );
NOR2_X2 U15256 ( .A1(n19196), .A2(n17872), .ZN(n16053) );
NOR2_X2 U15257 ( .A1(n19188), .A2(n17876), .ZN(n16054) );
NOR2_X2 U15258 ( .A1(n15968), .A2(n15969), .ZN(n15966) );
NOR2_X2 U15259 ( .A1(n19191), .A2(n17872), .ZN(n15968) );
NOR2_X2 U15260 ( .A1(n19183), .A2(n17876), .ZN(n15969) );
NOR2_X2 U15261 ( .A1(n15985), .A2(n15986), .ZN(n15983) );
NOR2_X2 U15262 ( .A1(n19192), .A2(n17872), .ZN(n15985) );
NOR2_X2 U15263 ( .A1(n19184), .A2(n17876), .ZN(n15986) );
NOR2_X2 U15264 ( .A1(n16002), .A2(n16003), .ZN(n16000) );
NOR2_X2 U15265 ( .A1(n19193), .A2(n17872), .ZN(n16002) );
NOR2_X2 U15266 ( .A1(n19185), .A2(n17876), .ZN(n16003) );
NOR2_X2 U15267 ( .A1(n16019), .A2(n16020), .ZN(n16017) );
NOR2_X2 U15268 ( .A1(n19194), .A2(n17872), .ZN(n16019) );
NOR2_X2 U15269 ( .A1(n19186), .A2(n17876), .ZN(n16020) );
NOR2_X2 U15270 ( .A1(n16036), .A2(n16037), .ZN(n16034) );
NOR2_X2 U15271 ( .A1(n19195), .A2(n17872), .ZN(n16036) );
NOR2_X2 U15272 ( .A1(n19187), .A2(n17876), .ZN(n16037) );
NOR2_X2 U15273 ( .A1(n16070), .A2(n16071), .ZN(n16068) );
NOR2_X2 U15274 ( .A1(n19197), .A2(n17872), .ZN(n16070) );
NOR2_X2 U15275 ( .A1(n19189), .A2(n17876), .ZN(n16071) );
NOR2_X2 U15276 ( .A1(n18071), .A2(n18074), .ZN(n14393) );
INV_X4 U15277 ( .A(n17775), .ZN(n17898) );
INV_X4 U15278 ( .A(n17283), .ZN(n18002) );
INV_X4 U15279 ( .A(n17775), .ZN(n17899) );
BUF_X4 U15280 ( .A(n17752), .Z(n17823) );
BUF_X4 U15281 ( .A(n17753), .Z(n17822) );
BUF_X4 U15282 ( .A(n17818), .Z(n17821) );
BUF_X4 U15283 ( .A(n17751), .Z(n17820) );
BUF_X4 U15284 ( .A(n17752), .Z(n17819) );
BUF_X4 U15285 ( .A(n18632), .Z(n17835) );
BUF_X4 U15286 ( .A(n17753), .Z(n17834) );
BUF_X4 U15287 ( .A(n17752), .Z(n17833) );
BUF_X4 U15288 ( .A(n17751), .Z(n17832) );
BUF_X4 U15289 ( .A(n17826), .Z(n17831) );
BUF_X4 U15290 ( .A(n17751), .Z(n17830) );
BUF_X4 U15291 ( .A(n17752), .Z(n17829) );
BUF_X4 U15292 ( .A(n17753), .Z(n17828) );
BUF_X4 U15293 ( .A(n17830), .Z(n17827) );
BUF_X4 U15294 ( .A(n17751), .Z(n17826) );
BUF_X4 U15295 ( .A(n17752), .Z(n17825) );
BUF_X4 U15296 ( .A(n17753), .Z(n17824) );
BUF_X4 U15297 ( .A(n17751), .Z(n17818) );
BUF_X4 U15298 ( .A(n17752), .Z(n17836) );
NOR4_X2 U15299 ( .A1(n14157), .A2(state[0]), .A3(state[1]), .A4(state[4]),.ZN(n12235) );
NOR4_X2 U15300 ( .A1(n14402), .A2(n14403), .A3(n14404), .A4(n18743), .ZN(n14401) );
NOR4_X2 U15301 ( .A1(n14427), .A2(n14428), .A3(n14429), .A4(n18742), .ZN(n14426) );
NOR4_X2 U15302 ( .A1(n14449), .A2(n14450), .A3(n14451), .A4(n18741), .ZN(n14448) );
NOR4_X2 U15303 ( .A1(n14471), .A2(n14472), .A3(n14473), .A4(n18740), .ZN(n14470) );
NOR4_X2 U15304 ( .A1(n14493), .A2(n14494), .A3(n14495), .A4(n18739), .ZN(n14492) );
NOR4_X2 U15305 ( .A1(n14515), .A2(n14516), .A3(n14517), .A4(n18738), .ZN(n14514) );
NOR4_X2 U15306 ( .A1(n14537), .A2(n14538), .A3(n14539), .A4(n18737), .ZN(n14536) );
NOR4_X2 U15307 ( .A1(n14559), .A2(n14560), .A3(n14561), .A4(n18736), .ZN(n14558) );
NOR4_X2 U15308 ( .A1(n15814), .A2(n18682), .A3(n15815), .A4(n15816), .ZN(n15813) );
NOR2_X2 U15309 ( .A1(n19143), .A2(n17903), .ZN(n15815) );
NOR4_X2 U15310 ( .A1(n15832), .A2(n18681), .A3(n15833), .A4(n15834), .ZN(n15831) );
NOR2_X2 U15311 ( .A1(n19144), .A2(n17903), .ZN(n15833) );
NOR4_X2 U15312 ( .A1(n15850), .A2(n18680), .A3(n15851), .A4(n15852), .ZN(n15849) );
NOR2_X2 U15313 ( .A1(n19145), .A2(n17903), .ZN(n15851) );
NOR4_X2 U15314 ( .A1(n15868), .A2(n18679), .A3(n15869), .A4(n15870), .ZN(n15867) );
NOR2_X2 U15315 ( .A1(n5329), .A2(n18001), .ZN(n15870) );
NOR2_X2 U15316 ( .A1(n19146), .A2(n17903), .ZN(n15869) );
NOR4_X2 U15317 ( .A1(n15886), .A2(n18678), .A3(n15887), .A4(n15888), .ZN(n15885) );
NOR2_X2 U15318 ( .A1(n5330), .A2(n18000), .ZN(n15888) );
NOR2_X2 U15319 ( .A1(n19147), .A2(n17903), .ZN(n15887) );
NOR4_X2 U15320 ( .A1(n15904), .A2(n18677), .A3(n15905), .A4(n15906), .ZN(n15903) );
NOR2_X2 U15321 ( .A1(n5331), .A2(n18000), .ZN(n15906) );
NOR2_X2 U15322 ( .A1(n19148), .A2(n17903), .ZN(n15905) );
NOR4_X2 U15323 ( .A1(n15922), .A2(n18676), .A3(n15923), .A4(n15924), .ZN(n15921) );
NOR2_X2 U15324 ( .A1(n5332), .A2(n18000), .ZN(n15924) );
NOR2_X2 U15325 ( .A1(n19149), .A2(n17903), .ZN(n15923) );
NOR4_X2 U15326 ( .A1(n15940), .A2(n18675), .A3(n15941), .A4(n15942), .ZN(n15939) );
NOR2_X2 U15327 ( .A1(n5333), .A2(n18000), .ZN(n15942) );
NOR2_X2 U15328 ( .A1(n19150), .A2(n17903), .ZN(n15941) );
NOR4_X2 U15329 ( .A1(n16334), .A2(n18650), .A3(n16335), .A4(n16336), .ZN(n16333) );
NOR2_X2 U15330 ( .A1(n5358), .A2(n18001), .ZN(n16336) );
NOR2_X2 U15331 ( .A1(n19175), .A2(n17904), .ZN(n16335) );
NOR4_X2 U15332 ( .A1(n16347), .A2(n18649), .A3(n16348), .A4(n16349), .ZN(n16346) );
NOR2_X2 U15333 ( .A1(n5359), .A2(n18001), .ZN(n16349) );
NOR2_X2 U15334 ( .A1(n19176), .A2(n17904), .ZN(n16348) );
NOR4_X2 U15335 ( .A1(n16360), .A2(n18648), .A3(n16361), .A4(n16362), .ZN(n16359) );
NOR2_X2 U15336 ( .A1(n5360), .A2(n18001), .ZN(n16362) );
NOR2_X2 U15337 ( .A1(n19177), .A2(n17904), .ZN(n16361) );
NOR4_X2 U15338 ( .A1(n16373), .A2(n18647), .A3(n16374), .A4(n16375), .ZN(n16372) );
NOR2_X2 U15339 ( .A1(n5361), .A2(n18001), .ZN(n16375) );
NOR2_X2 U15340 ( .A1(n19178), .A2(n17904), .ZN(n16374) );
NOR4_X2 U15341 ( .A1(n16386), .A2(n18646), .A3(n16387), .A4(n16388), .ZN(n16385) );
NOR2_X2 U15342 ( .A1(n5362), .A2(n18001), .ZN(n16388) );
NOR2_X2 U15343 ( .A1(n19179), .A2(n17905), .ZN(n16387) );
NOR4_X2 U15344 ( .A1(n16399), .A2(n18645), .A3(n16400), .A4(n16401), .ZN(n16398) );
NOR2_X2 U15345 ( .A1(n5363), .A2(n18002), .ZN(n16401) );
NOR2_X2 U15346 ( .A1(n19180), .A2(n17905), .ZN(n16400) );
NOR4_X2 U15347 ( .A1(n16412), .A2(n18644), .A3(n16413), .A4(n16414), .ZN(n16411) );
NOR2_X2 U15348 ( .A1(n5364), .A2(n18002), .ZN(n16414) );
NOR2_X2 U15349 ( .A1(n19181), .A2(n17905), .ZN(n16413) );
NOR4_X2 U15350 ( .A1(n16425), .A2(n18643), .A3(n16426), .A4(n16427), .ZN(n16424) );
NOR2_X2 U15351 ( .A1(n5365), .A2(n18002), .ZN(n16427) );
NOR2_X2 U15352 ( .A1(n19182), .A2(n17905), .ZN(n16426) );
NOR4_X2 U15353 ( .A1(n15601), .A2(n15602), .A3(n15603), .A4(n15604), .ZN(n15600) );
NOR2_X2 U15354 ( .A1(n15605), .A2(n17918), .ZN(n15604) );
NOR4_X2 U15355 ( .A1(n15620), .A2(n15621), .A3(n15622), .A4(n15623), .ZN(n15619) );
NOR2_X2 U15356 ( .A1(n15624), .A2(n17918), .ZN(n15623) );
NOR4_X2 U15357 ( .A1(n15639), .A2(n15640), .A3(n15641), .A4(n15642), .ZN(n15638) );
NOR2_X2 U15358 ( .A1(n15643), .A2(n17918), .ZN(n15642) );
NOR4_X2 U15359 ( .A1(n16097), .A2(n18666), .A3(n16098), .A4(n16099), .ZN(n16096) );
NOR2_X2 U15360 ( .A1(n5342), .A2(n18000), .ZN(n16099) );
NOR2_X2 U15361 ( .A1(n19159), .A2(n17904), .ZN(n16098) );
NOR4_X2 U15362 ( .A1(n16113), .A2(n18665), .A3(n16114), .A4(n16115), .ZN(n16112) );
NOR2_X2 U15363 ( .A1(n5343), .A2(n18001), .ZN(n16115) );
NOR2_X2 U15364 ( .A1(n19160), .A2(n17904), .ZN(n16114) );
NOR4_X2 U15365 ( .A1(n16128), .A2(n18664), .A3(n16129), .A4(n16130), .ZN(n16127) );
NOR2_X2 U15366 ( .A1(n5344), .A2(n18001), .ZN(n16130) );
NOR2_X2 U15367 ( .A1(n19161), .A2(n17904), .ZN(n16129) );
NOR4_X2 U15368 ( .A1(n16143), .A2(n18663), .A3(n16144), .A4(n16145), .ZN(n16142) );
NOR2_X2 U15369 ( .A1(n5345), .A2(n18001), .ZN(n16145) );
NOR2_X2 U15370 ( .A1(n19162), .A2(n17904), .ZN(n16144) );
NOR4_X2 U15371 ( .A1(n16158), .A2(n18662), .A3(n16159), .A4(n16160), .ZN(n16157) );
NOR2_X2 U15372 ( .A1(n5346), .A2(n18001), .ZN(n16160) );
NOR2_X2 U15373 ( .A1(n19163), .A2(n17904), .ZN(n16159) );
NOR4_X2 U15374 ( .A1(n16173), .A2(n18661), .A3(n16174), .A4(n16175), .ZN(n16172) );
NOR2_X2 U15375 ( .A1(n5347), .A2(n18001), .ZN(n16175) );
NOR2_X2 U15376 ( .A1(n19164), .A2(n17904), .ZN(n16174) );
NOR4_X2 U15377 ( .A1(n16188), .A2(n18660), .A3(n16189), .A4(n16190), .ZN(n16187) );
NOR2_X2 U15378 ( .A1(n5348), .A2(n18001), .ZN(n16190) );
NOR2_X2 U15379 ( .A1(n19165), .A2(n17904), .ZN(n16189) );
NOR4_X2 U15380 ( .A1(n16203), .A2(n18659), .A3(n16204), .A4(n16205), .ZN(n16202) );
NOR2_X2 U15381 ( .A1(n5349), .A2(n18001), .ZN(n16205) );
NOR2_X2 U15382 ( .A1(n19166), .A2(n17904), .ZN(n16204) );
NOR2_X2 U15383 ( .A1(n18036), .A2(n16549), .ZN(N3077) );
NOR2_X2 U15384 ( .A1(n18036), .A2(n16554), .ZN(N3076) );
NOR2_X2 U15385 ( .A1(n18036), .A2(n16559), .ZN(N3075) );
NOR2_X2 U15386 ( .A1(n18036), .A2(n16564), .ZN(N3074) );
AND3_X2 U15387 ( .A1(n17759), .A2(n13364), .A3(n17760), .ZN(n16440) );
OR2_X4 U15388 ( .A1(n19191), .A2(n16450), .ZN(n17759) );
NAND3_X2 U15389 ( .A1(n18634), .A2(n13365), .A3(aes_text_out[15]), .ZN(n17760) );
AND3_X2 U15390 ( .A1(n17761), .A2(n13358), .A3(n17762), .ZN(n16455) );
OR2_X4 U15391 ( .A1(n19192), .A2(n16450), .ZN(n17761) );
NAND3_X2 U15392 ( .A1(n18634), .A2(n13359), .A3(aes_text_out[14]), .ZN(n17762) );
AND3_X2 U15393 ( .A1(n17763), .A2(n13352), .A3(n17764), .ZN(n16468) );
OR2_X4 U15394 ( .A1(n19193), .A2(n16450), .ZN(n17763) );
NAND3_X2 U15395 ( .A1(n18634), .A2(n13353), .A3(aes_text_out[13]), .ZN(n17764) );
AND3_X2 U15396 ( .A1(n17765), .A2(n13346), .A3(n17766), .ZN(n16481) );
OR2_X4 U15397 ( .A1(n19194), .A2(n16450), .ZN(n17765) );
NAND3_X2 U15398 ( .A1(n18634), .A2(n13347), .A3(aes_text_out[12]), .ZN(n17766) );
AND3_X2 U15399 ( .A1(n17767), .A2(n13340), .A3(n17768), .ZN(n16494) );
OR2_X4 U15400 ( .A1(n19195), .A2(n16450), .ZN(n17767) );
NAND3_X2 U15401 ( .A1(n18634), .A2(n13341), .A3(aes_text_out[11]), .ZN(n17768) );
AND3_X2 U15402 ( .A1(n17769), .A2(n13334), .A3(n17770), .ZN(n16507) );
OR2_X4 U15403 ( .A1(n19196), .A2(n16450), .ZN(n17769) );
NAND3_X2 U15404 ( .A1(n18634), .A2(n13335), .A3(aes_text_out[10]), .ZN(n17770) );
AND3_X2 U15405 ( .A1(n17771), .A2(n13328), .A3(n17772), .ZN(n16520) );
OR2_X4 U15406 ( .A1(n19197), .A2(n16450), .ZN(n17771) );
NAND3_X2 U15407 ( .A1(n18634), .A2(n13329), .A3(aes_text_out[9]), .ZN(n17772) );
AND3_X2 U15408 ( .A1(n17773), .A2(n13322), .A3(n17774), .ZN(n16533) );
OR2_X4 U15409 ( .A1(n19198), .A2(n16450), .ZN(n17773) );
NAND3_X2 U15410 ( .A1(n18634), .A2(n13323), .A3(aes_text_out[8]), .ZN(n17774) );
NAND3_X2 U15411 ( .A1(n16447), .A2(n18836), .A3(n16448), .ZN(n16446) );
NAND3_X2 U15412 ( .A1(n16461), .A2(n18837), .A3(n16462), .ZN(n16460) );
NAND3_X2 U15413 ( .A1(n16474), .A2(n18838), .A3(n16475), .ZN(n16473) );
NAND3_X2 U15414 ( .A1(n16487), .A2(n18839), .A3(n16488), .ZN(n16486) );
NAND3_X2 U15415 ( .A1(n16500), .A2(n18840), .A3(n16501), .ZN(n16499) );
NAND3_X2 U15416 ( .A1(n16513), .A2(n18841), .A3(n16514), .ZN(n16512) );
NAND3_X2 U15417 ( .A1(n16526), .A2(n18842), .A3(n16527), .ZN(n16525) );
NAND3_X2 U15418 ( .A1(n16540), .A2(n18843), .A3(n16541), .ZN(n16539) );
NOR2_X2 U15419 ( .A1(n18036), .A2(n16544), .ZN(N3078) );
NOR3_X2 U15420 ( .A1(n16546), .A2(n16547), .A3(n18642), .ZN(n16545) );
NOR2_X2 U15421 ( .A1(n5374), .A2(n18002), .ZN(n16547) );
OR3_X2 U15422 ( .A1(n19205), .A2(dii_data_size[2]), .A3(n19204), .ZN(n17775));
NAND3_X2 U15423 ( .A1(n12235), .A2(n18078), .A3(state[2]), .ZN(n11942) );
INV_X4 U15424 ( .A(dii_data_size[2]), .ZN(n18071) );
NOR2_X2 U15425 ( .A1(n18036), .A2(n16573), .ZN(N3072) );
NOR2_X2 U15426 ( .A1(n18636), .A2(n16575), .ZN(n16574) );
NOR2_X2 U15427 ( .A1(n19197), .A2(n17905), .ZN(n16575) );
NOR2_X2 U15428 ( .A1(n18037), .A2(n16577), .ZN(N3071) );
NOR2_X2 U15429 ( .A1(n18635), .A2(n16579), .ZN(n16578) );
NOR2_X2 U15430 ( .A1(n19198), .A2(n17905), .ZN(n16579) );
NAND3_X2 U15431 ( .A1(n11949), .A2(n18633), .A3(n11950), .ZN(n6285) );
INV_X4 U15432 ( .A(n14414), .ZN(n17886) );
NOR2_X2 U15433 ( .A1(n19205), .A2(dii_data_size[1]), .ZN(n14414) );
NAND3_X2 U15434 ( .A1(n14914), .A2(n18071), .A3(n19201), .ZN(n14736) );
NAND3_X2 U15435 ( .A1(n18846), .A2(n11929), .A3(n17748), .ZN(n11928) );
INV_X4 U15436 ( .A(dii_data_size[3]), .ZN(n18075) );
NOR2_X2 U15437 ( .A1(n11921), .A2(n18894), .ZN(n6295) );
NOR2_X2 U15438 ( .A1(n11922), .A2(n11923), .ZN(n11921) );
NOR2_X2 U15439 ( .A1(n11924), .A2(n18893), .ZN(n11922) );
NOR2_X2 U15440 ( .A1(n18036), .A2(n16569), .ZN(N3073) );
NOR2_X2 U15441 ( .A1(n18637), .A2(n16571), .ZN(n16570) );
NOR2_X2 U15442 ( .A1(n19196), .A2(n17905), .ZN(n16571) );
NAND3_X2 U15443 ( .A1(n14023), .A2(n14024), .A3(n14025), .ZN(n5574) );
NAND3_X2 U15444 ( .A1(n14019), .A2(n14020), .A3(n14021), .ZN(n5575) );
NAND3_X2 U15445 ( .A1(n14015), .A2(n14016), .A3(n14017), .ZN(n5576) );
NAND3_X2 U15446 ( .A1(n14011), .A2(n14012), .A3(n14013), .ZN(n5577) );
NAND3_X2 U15447 ( .A1(n14007), .A2(n14008), .A3(n14009), .ZN(n5578) );
NAND3_X2 U15448 ( .A1(n14003), .A2(n14004), .A3(n14005), .ZN(n5579) );
NAND3_X2 U15449 ( .A1(n13999), .A2(n14000), .A3(n14001), .ZN(n5580) );
NAND3_X2 U15450 ( .A1(n13995), .A2(n13996), .A3(n13997), .ZN(n5581) );
NOR2_X2 U15451 ( .A1(dii_data_size[0]), .A2(dii_data_size[1]), .ZN(n14564));
NOR2_X2 U15452 ( .A1(n18075), .A2(dii_data_size[2]), .ZN(n15309) );
NOR4_X2 U15453 ( .A1(n6850), .A2(n6859), .A3(n16839), .A4(n16838), .ZN(n11929) );
NOR2_X2 U15454 ( .A1(n14188), .A2(n14189), .ZN(n14178) );
NOR2_X2 U15455 ( .A1(n14217), .A2(n14218), .ZN(n14210) );
NOR2_X2 U15456 ( .A1(n14246), .A2(n14247), .ZN(n14239) );
NOR2_X2 U15457 ( .A1(n14275), .A2(n14276), .ZN(n14268) );
NOR2_X2 U15458 ( .A1(n14304), .A2(n14305), .ZN(n14297) );
NOR2_X2 U15459 ( .A1(n14333), .A2(n14334), .ZN(n14326) );
NOR2_X2 U15460 ( .A1(n14362), .A2(n14363), .ZN(n14355) );
NOR2_X2 U15461 ( .A1(n14394), .A2(n14395), .ZN(n14384) );
NOR2_X2 U15462 ( .A1(n15505), .A2(n15506), .ZN(n15495) );
NOR2_X2 U15463 ( .A1(n15529), .A2(n15530), .ZN(n15523) );
NOR2_X2 U15464 ( .A1(n15550), .A2(n15551), .ZN(n15544) );
NOR2_X2 U15465 ( .A1(n15571), .A2(n15572), .ZN(n15565) );
NOR2_X2 U15466 ( .A1(n15592), .A2(n15593), .ZN(n15586) );
NOR2_X2 U15467 ( .A1(n15614), .A2(n15615), .ZN(n15608) );
NOR2_X2 U15468 ( .A1(n15633), .A2(n15634), .ZN(n15627) );
NOR2_X2 U15469 ( .A1(n15653), .A2(n15654), .ZN(n15647) );
NAND3_X2 U15470 ( .A1(n14949), .A2(n17880), .A3(n14950), .ZN(n14597) );
NAND3_X2 U15471 ( .A1(n14971), .A2(n17880), .A3(n14972), .ZN(n14618) );
NAND3_X2 U15472 ( .A1(n14993), .A2(n17881), .A3(n14994), .ZN(n14639) );
NAND3_X2 U15473 ( .A1(n15015), .A2(n17881), .A3(n15016), .ZN(n14660) );
NAND3_X2 U15474 ( .A1(n15037), .A2(n17881), .A3(n15038), .ZN(n14681) );
NAND3_X2 U15475 ( .A1(n15059), .A2(n17880), .A3(n15060), .ZN(n14702) );
NAND3_X2 U15476 ( .A1(n15081), .A2(n17881), .A3(n15082), .ZN(n14723) );
NAND3_X2 U15477 ( .A1(n15105), .A2(n17880), .A3(n15106), .ZN(n14746) );
NAND3_X2 U15478 ( .A1(n15128), .A2(n17880), .A3(n15129), .ZN(n14768) );
NAND3_X2 U15479 ( .A1(n15150), .A2(n17880), .A3(n15151), .ZN(n14791) );
NAND3_X2 U15480 ( .A1(n15172), .A2(n17880), .A3(n15173), .ZN(n14813) );
NAND3_X2 U15481 ( .A1(n15194), .A2(n17880), .A3(n15195), .ZN(n14835) );
NAND3_X2 U15482 ( .A1(n15216), .A2(n17880), .A3(n15217), .ZN(n14857) );
NAND3_X2 U15483 ( .A1(n15238), .A2(n17880), .A3(n15239), .ZN(n14879) );
NAND3_X2 U15484 ( .A1(n15260), .A2(n17880), .A3(n15261), .ZN(n14901) );
NAND3_X2 U15485 ( .A1(n15284), .A2(n17880), .A3(n15285), .ZN(n14924) );
INV_X4 U15486 ( .A(dii_data_size[2]), .ZN(n18072) );
INV_X4 U15487 ( .A(dii_data_size[3]), .ZN(n18076) );
NAND2_X2 U15488 ( .A1(n17882), .A2(dii_data_size[0]), .ZN(n15507) );
INV_X4 U15489 ( .A(dii_data_size[2]), .ZN(n18073) );
INV_X4 U15490 ( .A(rst), .ZN(n18632) );
NAND2_X2 U15491 ( .A1(state[9]), .A2(n11926), .ZN(n18077) );
NAND2_X2 U15492 ( .A1(n18002), .A2(n18077), .ZN(n6294) );
NAND3_X2 U15493 ( .A1(n18630), .A2(n18078), .A3(n18611), .ZN(n18598) );
INV_X4 U15494 ( .A(n18598), .ZN(n18628) );
NAND2_X2 U15495 ( .A1(n18080), .A2(n18079), .ZN(n18597) );
INV_X4 U15496 ( .A(n18597), .ZN(n18627) );
NAND4_X2 U15497 ( .A1(n18600), .A2(n18601), .A3(n18627), .A4(n18626), .ZN(n14157) );
INV_X4 U15498 ( .A(n14157), .ZN(n18625) );
NAND4_X2 U15499 ( .A1(n18628), .A2(state[4]), .A3(n18625), .A4(n18631), .ZN(dii_data_not_ready) );
INV_X4 U15500 ( .A(dii_data_not_ready), .ZN(n18617) );
INV_X4 U15501 ( .A(dii_data_type), .ZN(n18081) );
NAND2_X2 U15502 ( .A1(n11958), .A2(n18085), .ZN(n18083) );
NAND2_X2 U15503 ( .A1(n17776), .A2(n18082), .ZN(n18088) );
NAND2_X2 U15504 ( .A1(n18083), .A2(n18085), .ZN(n18084) );
NAND2_X2 U15505 ( .A1(N2153), .A2(n17800), .ZN(n18086) );
NAND2_X2 U15506 ( .A1(n17776), .A2(n18089), .ZN(n18092) );
NAND2_X2 U15507 ( .A1(N2152), .A2(n17800), .ZN(n18090) );
NAND2_X2 U15508 ( .A1(n17776), .A2(n18093), .ZN(n18096) );
NAND2_X2 U15509 ( .A1(N2151), .A2(n17800), .ZN(n18094) );
NAND2_X2 U15510 ( .A1(n17776), .A2(n18097), .ZN(n18100) );
NAND2_X2 U15511 ( .A1(N2150), .A2(n17800), .ZN(n18098) );
NAND2_X2 U15512 ( .A1(n17776), .A2(n18101), .ZN(n18104) );
NAND2_X2 U15513 ( .A1(N2149), .A2(n17800), .ZN(n18102) );
NAND2_X2 U15514 ( .A1(n17776), .A2(n18105), .ZN(n18108) );
NAND2_X2 U15515 ( .A1(N2148), .A2(n17800), .ZN(n18106) );
NAND2_X2 U15516 ( .A1(n17776), .A2(n18109), .ZN(n18112) );
NAND2_X2 U15517 ( .A1(N2147), .A2(n17800), .ZN(n18110) );
NAND2_X2 U15518 ( .A1(n17776), .A2(n18113), .ZN(n18116) );
NAND2_X2 U15519 ( .A1(N2146), .A2(n17800), .ZN(n18114) );
NAND3_X2 U15520 ( .A1(n18116), .A2(n18115), .A3(n18114), .ZN(n5838) );
NAND2_X2 U15521 ( .A1(n17776), .A2(n18117), .ZN(n18120) );
NAND2_X2 U15522 ( .A1(N2145), .A2(n17800), .ZN(n18118) );
NAND3_X2 U15523 ( .A1(n18120), .A2(n18119), .A3(n18118), .ZN(n5839) );
NAND2_X2 U15524 ( .A1(n17776), .A2(n18121), .ZN(n18124) );
NAND2_X2 U15525 ( .A1(N2144), .A2(n17800), .ZN(n18122) );
NAND3_X2 U15526 ( .A1(n18124), .A2(n18123), .A3(n18122), .ZN(n5840) );
NAND2_X2 U15527 ( .A1(n17776), .A2(n18125), .ZN(n18128) );
NAND2_X2 U15528 ( .A1(N2143), .A2(n17800), .ZN(n18126) );
NAND3_X2 U15529 ( .A1(n18128), .A2(n18127), .A3(n18126), .ZN(n5841) );
NAND2_X2 U15530 ( .A1(n17777), .A2(n18129), .ZN(n18132) );
NAND2_X2 U15531 ( .A1(N2142), .A2(n17801), .ZN(n18130) );
NAND3_X2 U15532 ( .A1(n18132), .A2(n18131), .A3(n18130), .ZN(n5842) );
NAND2_X2 U15533 ( .A1(n17777), .A2(n18133), .ZN(n18136) );
NAND2_X2 U15534 ( .A1(N2141), .A2(n17801), .ZN(n18134) );
NAND3_X2 U15535 ( .A1(n18136), .A2(n18135), .A3(n18134), .ZN(n5843) );
NAND2_X2 U15536 ( .A1(n17777), .A2(n18137), .ZN(n18140) );
NAND2_X2 U15537 ( .A1(N2140), .A2(n17801), .ZN(n18138) );
NAND3_X2 U15538 ( .A1(n18140), .A2(n18139), .A3(n18138), .ZN(n5844) );
NAND2_X2 U15539 ( .A1(n17777), .A2(n18141), .ZN(n18144) );
NAND2_X2 U15540 ( .A1(N2139), .A2(n17801), .ZN(n18142) );
NAND3_X2 U15541 ( .A1(n18144), .A2(n18143), .A3(n18142), .ZN(n5845) );
NAND2_X2 U15542 ( .A1(n17777), .A2(n18145), .ZN(n18148) );
NAND2_X2 U15543 ( .A1(N2138), .A2(n17801), .ZN(n18146) );
NAND2_X2 U15544 ( .A1(n17777), .A2(n18149), .ZN(n18152) );
NAND2_X2 U15545 ( .A1(N2137), .A2(n17801), .ZN(n18150) );
NAND2_X2 U15546 ( .A1(n17777), .A2(n18153), .ZN(n18156) );
NAND2_X2 U15547 ( .A1(N2136), .A2(n17801), .ZN(n18154) );
NAND2_X2 U15548 ( .A1(n17777), .A2(n18157), .ZN(n18160) );
NAND2_X2 U15549 ( .A1(N2135), .A2(n17801), .ZN(n18158) );
NAND2_X2 U15550 ( .A1(n17777), .A2(n18161), .ZN(n18164) );
NAND2_X2 U15551 ( .A1(N2134), .A2(n17801), .ZN(n18162) );
NAND2_X2 U15552 ( .A1(n17777), .A2(n18165), .ZN(n18168) );
NAND2_X2 U15553 ( .A1(N2133), .A2(n17801), .ZN(n18166) );
NAND2_X2 U15554 ( .A1(n17777), .A2(n18169), .ZN(n18172) );
NAND2_X2 U15555 ( .A1(N2132), .A2(n17801), .ZN(n18170) );
NAND2_X2 U15556 ( .A1(n17778), .A2(n18173), .ZN(n18176) );
NAND2_X2 U15557 ( .A1(N2131), .A2(n17802), .ZN(n18174) );
NAND2_X2 U15558 ( .A1(n17778), .A2(n18177), .ZN(n18180) );
NAND2_X2 U15559 ( .A1(N2130), .A2(n17802), .ZN(n18178) );
NAND2_X2 U15560 ( .A1(n17778), .A2(n18181), .ZN(n18184) );
NAND2_X2 U15561 ( .A1(N2129), .A2(n17802), .ZN(n18182) );
NAND2_X2 U15562 ( .A1(n17778), .A2(n18185), .ZN(n18188) );
NAND2_X2 U15563 ( .A1(N2128), .A2(n17802), .ZN(n18186) );
NAND2_X2 U15564 ( .A1(n17778), .A2(n18189), .ZN(n18192) );
NAND2_X2 U15565 ( .A1(N2127), .A2(n17802), .ZN(n18190) );
NAND2_X2 U15566 ( .A1(n17778), .A2(n18193), .ZN(n18196) );
NAND2_X2 U15567 ( .A1(N2126), .A2(n17802), .ZN(n18194) );
NAND2_X2 U15568 ( .A1(n17778), .A2(n18197), .ZN(n18200) );
NAND2_X2 U15569 ( .A1(N2125), .A2(n17802), .ZN(n18198) );
NAND2_X2 U15570 ( .A1(n17778), .A2(n18201), .ZN(n18204) );
NAND2_X2 U15571 ( .A1(N2124), .A2(n17802), .ZN(n18202) );
NAND2_X2 U15572 ( .A1(n17778), .A2(n18205), .ZN(n18208) );
NAND2_X2 U15573 ( .A1(N2123), .A2(n17802), .ZN(n18206) );
NAND2_X2 U15574 ( .A1(n17778), .A2(n18209), .ZN(n18212) );
NAND2_X2 U15575 ( .A1(N2122), .A2(n17802), .ZN(n18210) );
NAND2_X2 U15576 ( .A1(n17778), .A2(n18213), .ZN(n18216) );
NAND2_X2 U15577 ( .A1(N2121), .A2(n17802), .ZN(n18214) );
NAND2_X2 U15578 ( .A1(n17779), .A2(n18217), .ZN(n18220) );
NAND2_X2 U15579 ( .A1(N2120), .A2(n17803), .ZN(n18218) );
NAND2_X2 U15580 ( .A1(n17779), .A2(n18221), .ZN(n18224) );
NAND2_X2 U15581 ( .A1(N2119), .A2(n17803), .ZN(n18222) );
NAND2_X2 U15582 ( .A1(n17779), .A2(n18225), .ZN(n18228) );
NAND2_X2 U15583 ( .A1(N2118), .A2(n17803), .ZN(n18226) );
NAND2_X2 U15584 ( .A1(n17779), .A2(n18229), .ZN(n18232) );
NAND2_X2 U15585 ( .A1(N2117), .A2(n17803), .ZN(n18230) );
NAND2_X2 U15586 ( .A1(n17779), .A2(n18233), .ZN(n18236) );
NAND2_X2 U15587 ( .A1(N2116), .A2(n17803), .ZN(n18234) );
NAND2_X2 U15588 ( .A1(n17779), .A2(n18237), .ZN(n18240) );
NAND2_X2 U15589 ( .A1(N2115), .A2(n17803), .ZN(n18238) );
NAND2_X2 U15590 ( .A1(n17779), .A2(n18241), .ZN(n18244) );
NAND2_X2 U15591 ( .A1(N2114), .A2(n17803), .ZN(n18242) );
NAND2_X2 U15592 ( .A1(n17779), .A2(n18245), .ZN(n18248) );
NAND2_X2 U15593 ( .A1(N2113), .A2(n17803), .ZN(n18246) );
NAND2_X2 U15594 ( .A1(n17779), .A2(n18249), .ZN(n18252) );
NAND2_X2 U15595 ( .A1(N2112), .A2(n17803), .ZN(n18250) );
NAND2_X2 U15596 ( .A1(n17779), .A2(n18253), .ZN(n18256) );
NAND2_X2 U15597 ( .A1(N2111), .A2(n17803), .ZN(n18254) );
NAND2_X2 U15598 ( .A1(n17779), .A2(n18257), .ZN(n18260) );
NAND2_X2 U15599 ( .A1(N2110), .A2(n17803), .ZN(n18258) );
NAND2_X2 U15600 ( .A1(n17780), .A2(n18261), .ZN(n18264) );
NAND2_X2 U15601 ( .A1(N2109), .A2(n17804), .ZN(n18262) );
NAND2_X2 U15602 ( .A1(n17780), .A2(n18265), .ZN(n18268) );
NAND2_X2 U15603 ( .A1(N2108), .A2(n17804), .ZN(n18266) );
NAND2_X2 U15604 ( .A1(n17780), .A2(n18269), .ZN(n18272) );
NAND2_X2 U15605 ( .A1(N2107), .A2(n17804), .ZN(n18270) );
NAND2_X2 U15606 ( .A1(n17780), .A2(n18273), .ZN(n18276) );
NAND2_X2 U15607 ( .A1(N2106), .A2(n17804), .ZN(n18274) );
NAND2_X2 U15608 ( .A1(n17780), .A2(n18277), .ZN(n18280) );
NAND2_X2 U15609 ( .A1(N2105), .A2(n17804), .ZN(n18278) );
NAND2_X2 U15610 ( .A1(n17780), .A2(n18281), .ZN(n18284) );
NAND2_X2 U15611 ( .A1(N2104), .A2(n17804), .ZN(n18282) );
NAND2_X2 U15612 ( .A1(n17780), .A2(n18285), .ZN(n18288) );
NAND2_X2 U15613 ( .A1(N2103), .A2(n17804), .ZN(n18286) );
NAND2_X2 U15614 ( .A1(n17780), .A2(n18289), .ZN(n18292) );
NAND2_X2 U15615 ( .A1(N2102), .A2(n17804), .ZN(n18290) );
NAND2_X2 U15616 ( .A1(n17780), .A2(n18293), .ZN(n18296) );
NAND2_X2 U15617 ( .A1(N2101), .A2(n17804), .ZN(n18294) );
NAND2_X2 U15618 ( .A1(n17780), .A2(n18297), .ZN(n18300) );
NAND2_X2 U15619 ( .A1(N2100), .A2(n17804), .ZN(n18298) );
NAND2_X2 U15620 ( .A1(n17780), .A2(n18301), .ZN(n18304) );
NAND2_X2 U15621 ( .A1(N2099), .A2(n17804), .ZN(n18302) );
NAND2_X2 U15622 ( .A1(n17781), .A2(n18305), .ZN(n18308) );
NAND2_X2 U15623 ( .A1(N2098), .A2(n17805), .ZN(n18306) );
NAND3_X2 U15624 ( .A1(n18308), .A2(n18307), .A3(n18306), .ZN(n5885) );
NAND2_X2 U15625 ( .A1(n17781), .A2(n18309), .ZN(n18312) );
NAND2_X2 U15626 ( .A1(N2097), .A2(n17805), .ZN(n18310) );
NAND3_X2 U15627 ( .A1(n18312), .A2(n18311), .A3(n18310), .ZN(n5886) );
NAND2_X2 U15628 ( .A1(n17781), .A2(n18313), .ZN(n18316) );
NAND2_X2 U15629 ( .A1(N2096), .A2(n17805), .ZN(n18314) );
NAND3_X2 U15630 ( .A1(n18316), .A2(n18315), .A3(n18314), .ZN(n5887) );
NAND2_X2 U15631 ( .A1(n17781), .A2(n18317), .ZN(n18320) );
NAND2_X2 U15632 ( .A1(N2095), .A2(n17805), .ZN(n18318) );
NAND3_X2 U15633 ( .A1(n18320), .A2(n18319), .A3(n18318), .ZN(n5888) );
NAND2_X2 U15634 ( .A1(n17781), .A2(n18321), .ZN(n18324) );
NAND2_X2 U15635 ( .A1(N2094), .A2(n17805), .ZN(n18322) );
NAND3_X2 U15636 ( .A1(n18324), .A2(n18323), .A3(n18322), .ZN(n5889) );
NAND2_X2 U15637 ( .A1(n17781), .A2(n18325), .ZN(n18328) );
NAND2_X2 U15638 ( .A1(N2093), .A2(n17805), .ZN(n18326) );
NAND2_X2 U15639 ( .A1(n17781), .A2(n18329), .ZN(n18332) );
NAND2_X2 U15640 ( .A1(N2092), .A2(n17805), .ZN(n18330) );
NAND2_X2 U15641 ( .A1(n17781), .A2(n18333), .ZN(n18336) );
NAND2_X2 U15642 ( .A1(N2091), .A2(n17805), .ZN(n18334) );
NAND2_X2 U15643 ( .A1(n17781), .A2(n18337), .ZN(n18340) );
NAND2_X2 U15644 ( .A1(N2090), .A2(n17805), .ZN(n18338) );
NAND2_X2 U15645 ( .A1(n17781), .A2(n18341), .ZN(n18344) );
NAND2_X2 U15646 ( .A1(N2089), .A2(n17805), .ZN(n18342) );
NAND2_X2 U15647 ( .A1(n17781), .A2(n18345), .ZN(n18348) );
NAND2_X2 U15648 ( .A1(N2088), .A2(n17805), .ZN(n18346) );
NAND2_X2 U15649 ( .A1(n17782), .A2(n18349), .ZN(n18352) );
NAND2_X2 U15650 ( .A1(N2087), .A2(n17806), .ZN(n18350) );
NAND2_X2 U15651 ( .A1(n17782), .A2(n18353), .ZN(n18356) );
NAND2_X2 U15652 ( .A1(N2086), .A2(n17806), .ZN(n18354) );
NAND2_X2 U15653 ( .A1(n17782), .A2(n18357), .ZN(n18360) );
NAND2_X2 U15654 ( .A1(N2085), .A2(n17806), .ZN(n18358) );
NAND2_X2 U15655 ( .A1(n17782), .A2(n18361), .ZN(n18364) );
NAND2_X2 U15656 ( .A1(N2084), .A2(n17806), .ZN(n18362) );
NAND2_X2 U15657 ( .A1(n17782), .A2(n18365), .ZN(n18368) );
NAND2_X2 U15658 ( .A1(N2083), .A2(n17806), .ZN(n18366) );
NAND2_X2 U15659 ( .A1(n17782), .A2(n18369), .ZN(n18372) );
NAND2_X2 U15660 ( .A1(N2082), .A2(n17806), .ZN(n18370) );
NAND2_X2 U15661 ( .A1(n17782), .A2(n18373), .ZN(n18376) );
NAND2_X2 U15662 ( .A1(N2081), .A2(n17806), .ZN(n18374) );
NAND2_X2 U15663 ( .A1(n17782), .A2(n18377), .ZN(n18380) );
NAND2_X2 U15664 ( .A1(N2080), .A2(n17806), .ZN(n18378) );
NAND2_X2 U15665 ( .A1(n17782), .A2(n18381), .ZN(n18384) );
NAND2_X2 U15666 ( .A1(N2079), .A2(n17806), .ZN(n18382) );
NAND2_X2 U15667 ( .A1(n17782), .A2(n18385), .ZN(n18388) );
NAND2_X2 U15668 ( .A1(N2078), .A2(n17806), .ZN(n18386) );
NAND2_X2 U15669 ( .A1(n17782), .A2(n18389), .ZN(n18392) );
NAND2_X2 U15670 ( .A1(N2077), .A2(n17806), .ZN(n18390) );
NAND2_X2 U15671 ( .A1(n17783), .A2(n18393), .ZN(n18396) );
NAND2_X2 U15672 ( .A1(N2076), .A2(n17807), .ZN(n18394) );
NAND2_X2 U15673 ( .A1(n17783), .A2(n18397), .ZN(n18400) );
NAND2_X2 U15674 ( .A1(N2075), .A2(n17807), .ZN(n18398) );
NAND2_X2 U15675 ( .A1(n17783), .A2(n18401), .ZN(n18404) );
NAND2_X2 U15676 ( .A1(N2074), .A2(n17807), .ZN(n18402) );
NAND2_X2 U15677 ( .A1(n17783), .A2(n18405), .ZN(n18408) );
NAND2_X2 U15678 ( .A1(N2073), .A2(n17807), .ZN(n18406) );
NAND2_X2 U15679 ( .A1(n17783), .A2(n18409), .ZN(n18412) );
NAND2_X2 U15680 ( .A1(N2072), .A2(n17807), .ZN(n18410) );
NAND2_X2 U15681 ( .A1(n17783), .A2(n18413), .ZN(n18416) );
NAND2_X2 U15682 ( .A1(N2071), .A2(n17807), .ZN(n18414) );
NAND2_X2 U15683 ( .A1(n17783), .A2(n18417), .ZN(n18420) );
NAND2_X2 U15684 ( .A1(N2070), .A2(n17807), .ZN(n18418) );
NAND2_X2 U15685 ( .A1(n17783), .A2(n18421), .ZN(n18424) );
NAND2_X2 U15686 ( .A1(N2069), .A2(n17807), .ZN(n18422) );
NAND2_X2 U15687 ( .A1(n17783), .A2(n18425), .ZN(n18428) );
NAND2_X2 U15688 ( .A1(N2068), .A2(n17807), .ZN(n18426) );
NAND2_X2 U15689 ( .A1(n17783), .A2(n18429), .ZN(n18432) );
NAND2_X2 U15690 ( .A1(N2067), .A2(n17807), .ZN(n18430) );
NAND2_X2 U15691 ( .A1(n17783), .A2(n18433), .ZN(n18436) );
NAND2_X2 U15692 ( .A1(N2066), .A2(n17807), .ZN(n18434) );
NAND3_X2 U15693 ( .A1(n18436), .A2(n18435), .A3(n18434), .ZN(n5917) );
NAND2_X2 U15694 ( .A1(n17784), .A2(n18437), .ZN(n18440) );
NAND2_X2 U15695 ( .A1(N2065), .A2(n17808), .ZN(n18438) );
NAND3_X2 U15696 ( .A1(n18440), .A2(n18439), .A3(n18438), .ZN(n5918) );
NAND2_X2 U15697 ( .A1(n17784), .A2(n18441), .ZN(n18444) );
NAND2_X2 U15698 ( .A1(N2064), .A2(n17808), .ZN(n18442) );
NAND3_X2 U15699 ( .A1(n18444), .A2(n18443), .A3(n18442), .ZN(n5919) );
NAND2_X2 U15700 ( .A1(n17784), .A2(n18445), .ZN(n18448) );
NAND2_X2 U15701 ( .A1(N2063), .A2(n17808), .ZN(n18446) );
NAND3_X2 U15702 ( .A1(n18448), .A2(n18447), .A3(n18446), .ZN(n5920) );
NAND2_X2 U15703 ( .A1(n17784), .A2(n18449), .ZN(n18452) );
NAND2_X2 U15704 ( .A1(N2062), .A2(n17808), .ZN(n18450) );
NAND3_X2 U15705 ( .A1(n18452), .A2(n18451), .A3(n18450), .ZN(n5921) );
NAND2_X2 U15706 ( .A1(n17784), .A2(n18453), .ZN(n18456) );
NAND2_X2 U15707 ( .A1(N2061), .A2(n17808), .ZN(n18454) );
NAND3_X2 U15708 ( .A1(n18456), .A2(n18455), .A3(n18454), .ZN(n5922) );
NAND2_X2 U15709 ( .A1(n17784), .A2(n18457), .ZN(n18460) );
NAND2_X2 U15710 ( .A1(N2060), .A2(n17808), .ZN(n18458) );
NAND3_X2 U15711 ( .A1(n18460), .A2(n18459), .A3(n18458), .ZN(n5923) );
NAND2_X2 U15712 ( .A1(n17784), .A2(n18461), .ZN(n18464) );
NAND2_X2 U15713 ( .A1(N2059), .A2(n17808), .ZN(n18462) );
NAND3_X2 U15714 ( .A1(n18464), .A2(n18463), .A3(n18462), .ZN(n5924) );
NAND2_X2 U15715 ( .A1(n17784), .A2(n18465), .ZN(n18468) );
NAND2_X2 U15716 ( .A1(N2058), .A2(n17808), .ZN(n18466) );
NAND3_X2 U15717 ( .A1(n18468), .A2(n18467), .A3(n18466), .ZN(n5925) );
NAND2_X2 U15718 ( .A1(n17784), .A2(n18469), .ZN(n18472) );
NAND2_X2 U15719 ( .A1(N2057), .A2(n17808), .ZN(n18470) );
NAND3_X2 U15720 ( .A1(n18472), .A2(n18471), .A3(n18470), .ZN(n5926) );
NAND2_X2 U15721 ( .A1(n17784), .A2(n18473), .ZN(n18476) );
NAND2_X2 U15722 ( .A1(N2056), .A2(n17808), .ZN(n18474) );
NAND3_X2 U15723 ( .A1(n18476), .A2(n18475), .A3(n18474), .ZN(n5927) );
NAND2_X2 U15724 ( .A1(n17784), .A2(n18477), .ZN(n18480) );
NAND2_X2 U15725 ( .A1(N2055), .A2(n17808), .ZN(n18478) );
NAND3_X2 U15726 ( .A1(n18480), .A2(n18479), .A3(n18478), .ZN(n5928) );
NAND2_X2 U15727 ( .A1(n17785), .A2(n18481), .ZN(n18484) );
NAND2_X2 U15728 ( .A1(N2054), .A2(n17809), .ZN(n18482) );
NAND3_X2 U15729 ( .A1(n18484), .A2(n18483), .A3(n18482), .ZN(n5929) );
NAND2_X2 U15730 ( .A1(n17785), .A2(n18485), .ZN(n18488) );
NAND2_X2 U15731 ( .A1(N2053), .A2(n17809), .ZN(n18486) );
NAND3_X2 U15732 ( .A1(n18488), .A2(n18487), .A3(n18486), .ZN(n5930) );
NAND2_X2 U15733 ( .A1(n17785), .A2(n18489), .ZN(n18492) );
NAND2_X2 U15734 ( .A1(N2052), .A2(n17809), .ZN(n18490) );
NAND3_X2 U15735 ( .A1(n18492), .A2(n18491), .A3(n18490), .ZN(n5931) );
NAND2_X2 U15736 ( .A1(n17785), .A2(n18493), .ZN(n18496) );
NAND2_X2 U15737 ( .A1(N2051), .A2(n17809), .ZN(n18494) );
NAND3_X2 U15738 ( .A1(n18496), .A2(n18495), .A3(n18494), .ZN(n5932) );
NAND2_X2 U15739 ( .A1(n17785), .A2(n18497), .ZN(n18500) );
NAND2_X2 U15740 ( .A1(N2050), .A2(n17809), .ZN(n18498) );
NAND3_X2 U15741 ( .A1(n18500), .A2(n18499), .A3(n18498), .ZN(n5933) );
NAND2_X2 U15742 ( .A1(n17785), .A2(n18501), .ZN(n18504) );
NAND2_X2 U15743 ( .A1(N2049), .A2(n17809), .ZN(n18502) );
NAND3_X2 U15744 ( .A1(n18504), .A2(n18503), .A3(n18502), .ZN(n5934) );
NAND2_X2 U15745 ( .A1(n17785), .A2(n18505), .ZN(n18508) );
NAND2_X2 U15746 ( .A1(N2048), .A2(n17809), .ZN(n18506) );
NAND3_X2 U15747 ( .A1(n18508), .A2(n18507), .A3(n18506), .ZN(n5935) );
NAND2_X2 U15748 ( .A1(n17785), .A2(n18509), .ZN(n18512) );
NAND2_X2 U15749 ( .A1(N2047), .A2(n17809), .ZN(n18510) );
NAND3_X2 U15750 ( .A1(n18512), .A2(n18511), .A3(n18510), .ZN(n5936) );
NAND2_X2 U15751 ( .A1(n17785), .A2(n18513), .ZN(n18516) );
NAND2_X2 U15752 ( .A1(N2046), .A2(n17809), .ZN(n18514) );
NAND3_X2 U15753 ( .A1(n18516), .A2(n18515), .A3(n18514), .ZN(n5937) );
NAND2_X2 U15754 ( .A1(n17785), .A2(n18517), .ZN(n18520) );
NAND2_X2 U15755 ( .A1(N2045), .A2(n17809), .ZN(n18518) );
NAND3_X2 U15756 ( .A1(n18520), .A2(n18519), .A3(n18518), .ZN(n5938) );
NAND2_X2 U15757 ( .A1(n17785), .A2(n18521), .ZN(n18524) );
NAND2_X2 U15758 ( .A1(N2044), .A2(n17809), .ZN(n18522) );
NAND3_X2 U15759 ( .A1(n18524), .A2(n18523), .A3(n18522), .ZN(n5939) );
NAND2_X2 U15760 ( .A1(n17786), .A2(n18525), .ZN(n18528) );
NAND2_X2 U15761 ( .A1(N2043), .A2(n17810), .ZN(n18526) );
NAND3_X2 U15762 ( .A1(n18528), .A2(n18527), .A3(n18526), .ZN(n5940) );
NAND2_X2 U15763 ( .A1(n17786), .A2(n18529), .ZN(n18532) );
NAND2_X2 U15764 ( .A1(N2042), .A2(n17810), .ZN(n18530) );
NAND3_X2 U15765 ( .A1(n18532), .A2(n18531), .A3(n18530), .ZN(n5941) );
NAND2_X2 U15766 ( .A1(n17786), .A2(n18533), .ZN(n18536) );
NAND2_X2 U15767 ( .A1(N2041), .A2(n17810), .ZN(n18534) );
NAND3_X2 U15768 ( .A1(n18536), .A2(n18535), .A3(n18534), .ZN(n5942) );
NAND2_X2 U15769 ( .A1(n17786), .A2(n18537), .ZN(n18540) );
NAND2_X2 U15770 ( .A1(N2040), .A2(n17810), .ZN(n18538) );
NAND3_X2 U15771 ( .A1(n18540), .A2(n18539), .A3(n18538), .ZN(n5943) );
NAND2_X2 U15772 ( .A1(n17786), .A2(n18541), .ZN(n18544) );
NAND2_X2 U15773 ( .A1(N2039), .A2(n17810), .ZN(n18542) );
NAND3_X2 U15774 ( .A1(n18544), .A2(n18543), .A3(n18542), .ZN(n5944) );
NAND2_X2 U15775 ( .A1(n17786), .A2(n18545), .ZN(n18548) );
NAND2_X2 U15776 ( .A1(N2038), .A2(n17810), .ZN(n18546) );
NAND3_X2 U15777 ( .A1(n18548), .A2(n18547), .A3(n18546), .ZN(n5945) );
NAND2_X2 U15778 ( .A1(n17786), .A2(n18549), .ZN(n18552) );
NAND2_X2 U15779 ( .A1(N2037), .A2(n17810), .ZN(n18550) );
NAND3_X2 U15780 ( .A1(n18552), .A2(n18551), .A3(n18550), .ZN(n5946) );
NAND2_X2 U15781 ( .A1(n17786), .A2(n18553), .ZN(n18556) );
NAND2_X2 U15782 ( .A1(N2036), .A2(n17810), .ZN(n18554) );
NAND3_X2 U15783 ( .A1(n18556), .A2(n18555), .A3(n18554), .ZN(n5947) );
NAND2_X2 U15784 ( .A1(n17786), .A2(n18557), .ZN(n18560) );
NAND2_X2 U15785 ( .A1(N2035), .A2(n17810), .ZN(n18558) );
NAND3_X2 U15786 ( .A1(n18560), .A2(n18559), .A3(n18558), .ZN(n5948) );
NAND2_X2 U15787 ( .A1(n17786), .A2(n18561), .ZN(n18564) );
NAND2_X2 U15788 ( .A1(N2034), .A2(n17810), .ZN(n18562) );
NAND3_X2 U15789 ( .A1(n18564), .A2(n18563), .A3(n18562), .ZN(n5949) );
NAND2_X2 U15790 ( .A1(n17786), .A2(n18565), .ZN(n18568) );
NAND2_X2 U15791 ( .A1(N2033), .A2(n17810), .ZN(n18566) );
NAND3_X2 U15792 ( .A1(n18568), .A2(n18567), .A3(n18566), .ZN(n5950) );
NAND2_X2 U15793 ( .A1(n17787), .A2(n18569), .ZN(n18572) );
NAND2_X2 U15794 ( .A1(N2032), .A2(n17811), .ZN(n18570) );
NAND3_X2 U15795 ( .A1(n18572), .A2(n18571), .A3(n18570), .ZN(n5951) );
NAND2_X2 U15796 ( .A1(n17787), .A2(n18573), .ZN(n18576) );
NAND2_X2 U15797 ( .A1(N2031), .A2(n17811), .ZN(n18574) );
NAND3_X2 U15798 ( .A1(n18576), .A2(n18575), .A3(n18574), .ZN(n5952) );
NAND2_X2 U15799 ( .A1(n17787), .A2(n18577), .ZN(n18580) );
NAND2_X2 U15800 ( .A1(N2030), .A2(n17811), .ZN(n18578) );
NAND3_X2 U15801 ( .A1(n18580), .A2(n18579), .A3(n18578), .ZN(n5953) );
NAND2_X2 U15802 ( .A1(n17787), .A2(n18581), .ZN(n18584) );
NAND2_X2 U15803 ( .A1(N2029), .A2(n17811), .ZN(n18582) );
NAND3_X2 U15804 ( .A1(n18584), .A2(n18583), .A3(n18582), .ZN(n5954) );
NAND2_X2 U15805 ( .A1(n17787), .A2(n18585), .ZN(n18588) );
NAND2_X2 U15806 ( .A1(N2028), .A2(n17811), .ZN(n18586) );
NAND3_X2 U15807 ( .A1(n18588), .A2(n18587), .A3(n18586), .ZN(n5955) );
NAND2_X2 U15808 ( .A1(n17787), .A2(n18589), .ZN(n18592) );
NAND2_X2 U15809 ( .A1(N2027), .A2(n17811), .ZN(n18590) );
NAND3_X2 U15810 ( .A1(n18592), .A2(n18591), .A3(n18590), .ZN(n5956) );
NAND2_X2 U15811 ( .A1(n17787), .A2(n18593), .ZN(n18596) );
NAND2_X2 U15812 ( .A1(N2154), .A2(n17811), .ZN(n18594) );
NOR4_X2 U15813 ( .A1(state[4]), .A2(n18598), .A3(n18626), .A4(n18597), .ZN(n18599) );
NAND4_X2 U15814 ( .A1(n18631), .A2(n18601), .A3(n18600), .A4(n18599), .ZN(n11939) );
NAND2_X2 U15815 ( .A1(n11942), .A2(n11939), .ZN(n18602) );
NOR2_X2 U15816 ( .A1(n5444), .A2(n18003), .ZN(aes_text_in[127]) );
NOR2_X2 U15817 ( .A1(n5445), .A2(n18014), .ZN(aes_text_in[126]) );
NOR2_X2 U15818 ( .A1(n5446), .A2(n18014), .ZN(aes_text_in[125]) );
NOR2_X2 U15819 ( .A1(n5447), .A2(n18014), .ZN(aes_text_in[124]) );
NOR2_X2 U15820 ( .A1(n5448), .A2(n18014), .ZN(aes_text_in[123]) );
NOR2_X2 U15821 ( .A1(n5449), .A2(n18014), .ZN(aes_text_in[122]) );
NOR2_X2 U15822 ( .A1(n5450), .A2(n18014), .ZN(aes_text_in[121]) );
NOR2_X2 U15823 ( .A1(n5451), .A2(n18014), .ZN(aes_text_in[120]) );
NOR2_X2 U15824 ( .A1(n5452), .A2(n18013), .ZN(aes_text_in[119]) );
NOR2_X2 U15825 ( .A1(n5453), .A2(n18013), .ZN(aes_text_in[118]) );
NOR2_X2 U15826 ( .A1(n5454), .A2(n18013), .ZN(aes_text_in[117]) );
NOR2_X2 U15827 ( .A1(n5455), .A2(n18013), .ZN(aes_text_in[116]) );
NOR2_X2 U15828 ( .A1(n5456), .A2(n18013), .ZN(aes_text_in[115]) );
NOR2_X2 U15829 ( .A1(n5457), .A2(n18013), .ZN(aes_text_in[114]) );
NOR2_X2 U15830 ( .A1(n5458), .A2(n18013), .ZN(aes_text_in[113]) );
NOR2_X2 U15831 ( .A1(n5459), .A2(n18013), .ZN(aes_text_in[112]) );
NOR2_X2 U15832 ( .A1(n5460), .A2(n18013), .ZN(aes_text_in[111]) );
NOR2_X2 U15833 ( .A1(n5461), .A2(n18013), .ZN(aes_text_in[110]) );
NOR2_X2 U15834 ( .A1(n5462), .A2(n18012), .ZN(aes_text_in[109]) );
NOR2_X2 U15835 ( .A1(n5463), .A2(n18013), .ZN(aes_text_in[108]) );
NOR2_X2 U15836 ( .A1(n5464), .A2(n18012), .ZN(aes_text_in[107]) );
NOR2_X2 U15837 ( .A1(n5465), .A2(n18012), .ZN(aes_text_in[106]) );
NOR2_X2 U15838 ( .A1(n5466), .A2(n18012), .ZN(aes_text_in[105]) );
NOR2_X2 U15839 ( .A1(n5467), .A2(n18012), .ZN(aes_text_in[104]) );
NOR2_X2 U15840 ( .A1(n5468), .A2(n18012), .ZN(aes_text_in[103]) );
NOR2_X2 U15841 ( .A1(n5469), .A2(n18012), .ZN(aes_text_in[102]) );
NOR2_X2 U15842 ( .A1(n5470), .A2(n18012), .ZN(aes_text_in[101]) );
NOR2_X2 U15843 ( .A1(n5471), .A2(n18012), .ZN(aes_text_in[100]) );
NOR2_X2 U15844 ( .A1(n5472), .A2(n18012), .ZN(aes_text_in[99]) );
NOR2_X2 U15845 ( .A1(n5473), .A2(n18012), .ZN(aes_text_in[98]) );
NOR2_X2 U15846 ( .A1(n5474), .A2(n18011), .ZN(aes_text_in[97]) );
NOR2_X2 U15847 ( .A1(n5475), .A2(n18011), .ZN(aes_text_in[96]) );
NOR2_X2 U15848 ( .A1(n5476), .A2(n18011), .ZN(aes_text_in[95]) );
NOR2_X2 U15849 ( .A1(n5477), .A2(n18011), .ZN(aes_text_in[94]) );
NOR2_X2 U15850 ( .A1(n5478), .A2(n18011), .ZN(aes_text_in[93]) );
NOR2_X2 U15851 ( .A1(n5479), .A2(n18011), .ZN(aes_text_in[92]) );
NOR2_X2 U15852 ( .A1(n5480), .A2(n18011), .ZN(aes_text_in[91]) );
NOR2_X2 U15853 ( .A1(n5481), .A2(n18011), .ZN(aes_text_in[90]) );
NOR2_X2 U15854 ( .A1(n5482), .A2(n18011), .ZN(aes_text_in[89]) );
NOR2_X2 U15855 ( .A1(n5483), .A2(n18011), .ZN(aes_text_in[88]) );
NOR2_X2 U15856 ( .A1(n5484), .A2(n18011), .ZN(aes_text_in[87]) );
NOR2_X2 U15857 ( .A1(n5485), .A2(n18010), .ZN(aes_text_in[86]) );
NOR2_X2 U15858 ( .A1(n5486), .A2(n18010), .ZN(aes_text_in[85]) );
NOR2_X2 U15859 ( .A1(n5487), .A2(n18010), .ZN(aes_text_in[84]) );
NOR2_X2 U15860 ( .A1(n5488), .A2(n18010), .ZN(aes_text_in[83]) );
NOR2_X2 U15861 ( .A1(n5489), .A2(n18010), .ZN(aes_text_in[82]) );
NOR2_X2 U15862 ( .A1(n5490), .A2(n18010), .ZN(aes_text_in[81]) );
NOR2_X2 U15863 ( .A1(n5491), .A2(n18010), .ZN(aes_text_in[80]) );
NOR2_X2 U15864 ( .A1(n5492), .A2(n18010), .ZN(aes_text_in[79]) );
NOR2_X2 U15865 ( .A1(n5493), .A2(n18010), .ZN(aes_text_in[78]) );
NOR2_X2 U15866 ( .A1(n5494), .A2(n18010), .ZN(aes_text_in[77]) );
NOR2_X2 U15867 ( .A1(n5495), .A2(n18010), .ZN(aes_text_in[76]) );
NOR2_X2 U15868 ( .A1(n5496), .A2(n18009), .ZN(aes_text_in[75]) );
NOR2_X2 U15869 ( .A1(n5497), .A2(n18009), .ZN(aes_text_in[74]) );
NOR2_X2 U15870 ( .A1(n5498), .A2(n18009), .ZN(aes_text_in[73]) );
NOR2_X2 U15871 ( .A1(n5499), .A2(n18009), .ZN(aes_text_in[72]) );
NOR2_X2 U15872 ( .A1(n5500), .A2(n18009), .ZN(aes_text_in[71]) );
NOR2_X2 U15873 ( .A1(n5501), .A2(n18009), .ZN(aes_text_in[70]) );
NOR2_X2 U15874 ( .A1(n5502), .A2(n18009), .ZN(aes_text_in[69]) );
NOR2_X2 U15875 ( .A1(n5503), .A2(n18009), .ZN(aes_text_in[68]) );
NOR2_X2 U15876 ( .A1(n5504), .A2(n18009), .ZN(aes_text_in[67]) );
NOR2_X2 U15877 ( .A1(n5505), .A2(n18009), .ZN(aes_text_in[66]) );
NOR2_X2 U15878 ( .A1(n5506), .A2(n18009), .ZN(aes_text_in[65]) );
NOR2_X2 U15879 ( .A1(n5507), .A2(n18008), .ZN(aes_text_in[64]) );
NOR2_X2 U15880 ( .A1(n5508), .A2(n18008), .ZN(aes_text_in[63]) );
NOR2_X2 U15881 ( .A1(n5509), .A2(n18008), .ZN(aes_text_in[62]) );
NOR2_X2 U15882 ( .A1(n5510), .A2(n18008), .ZN(aes_text_in[61]) );
NOR2_X2 U15883 ( .A1(n5511), .A2(n18008), .ZN(aes_text_in[60]) );
NOR2_X2 U15884 ( .A1(n5512), .A2(n18008), .ZN(aes_text_in[59]) );
NOR2_X2 U15885 ( .A1(n5513), .A2(n18008), .ZN(aes_text_in[58]) );
NOR2_X2 U15886 ( .A1(n5514), .A2(n18008), .ZN(aes_text_in[57]) );
NOR2_X2 U15887 ( .A1(n5515), .A2(n18008), .ZN(aes_text_in[56]) );
NOR2_X2 U15888 ( .A1(n5516), .A2(n18008), .ZN(aes_text_in[55]) );
NOR2_X2 U15889 ( .A1(n5517), .A2(n18007), .ZN(aes_text_in[54]) );
NOR2_X2 U15890 ( .A1(n5518), .A2(n18007), .ZN(aes_text_in[53]) );
NOR2_X2 U15891 ( .A1(n5519), .A2(n18007), .ZN(aes_text_in[52]) );
NOR2_X2 U15892 ( .A1(n5520), .A2(n18007), .ZN(aes_text_in[51]) );
NOR2_X2 U15893 ( .A1(n5521), .A2(n18007), .ZN(aes_text_in[50]) );
NOR2_X2 U15894 ( .A1(n5522), .A2(n18007), .ZN(aes_text_in[49]) );
NOR2_X2 U15895 ( .A1(n5523), .A2(n18007), .ZN(aes_text_in[48]) );
NOR2_X2 U15896 ( .A1(n5524), .A2(n18007), .ZN(aes_text_in[47]) );
NOR2_X2 U15897 ( .A1(n5525), .A2(n18007), .ZN(aes_text_in[46]) );
NOR2_X2 U15898 ( .A1(n5526), .A2(n18007), .ZN(aes_text_in[45]) );
NOR2_X2 U15899 ( .A1(n5527), .A2(n18007), .ZN(aes_text_in[44]) );
NOR2_X2 U15900 ( .A1(n5528), .A2(n18006), .ZN(aes_text_in[43]) );
NOR2_X2 U15901 ( .A1(n5529), .A2(n18006), .ZN(aes_text_in[42]) );
NOR2_X2 U15902 ( .A1(n5530), .A2(n18006), .ZN(aes_text_in[41]) );
NOR2_X2 U15903 ( .A1(n5531), .A2(n18006), .ZN(aes_text_in[40]) );
NOR2_X2 U15904 ( .A1(n5532), .A2(n18006), .ZN(aes_text_in[39]) );
NOR2_X2 U15905 ( .A1(n5533), .A2(n18006), .ZN(aes_text_in[38]) );
NOR2_X2 U15906 ( .A1(n5534), .A2(n18006), .ZN(aes_text_in[37]) );
NOR2_X2 U15907 ( .A1(n5535), .A2(n18006), .ZN(aes_text_in[36]) );
NOR2_X2 U15908 ( .A1(n5536), .A2(n18006), .ZN(aes_text_in[35]) );
NOR2_X2 U15909 ( .A1(n5537), .A2(n18006), .ZN(aes_text_in[34]) );
NOR2_X2 U15910 ( .A1(n5538), .A2(n18006), .ZN(aes_text_in[33]) );
NOR2_X2 U15911 ( .A1(n5539), .A2(n18005), .ZN(aes_text_in[32]) );
NOR2_X2 U15912 ( .A1(n5540), .A2(n18005), .ZN(aes_text_in[31]) );
NOR2_X2 U15913 ( .A1(n5541), .A2(n18008), .ZN(aes_text_in[30]) );
NOR2_X2 U15914 ( .A1(n5542), .A2(n18005), .ZN(aes_text_in[29]) );
NOR2_X2 U15915 ( .A1(n5543), .A2(n18005), .ZN(aes_text_in[28]) );
NOR2_X2 U15916 ( .A1(n5544), .A2(n18005), .ZN(aes_text_in[27]) );
NOR2_X2 U15917 ( .A1(n5545), .A2(n18005), .ZN(aes_text_in[26]) );
NOR2_X2 U15918 ( .A1(n5546), .A2(n18005), .ZN(aes_text_in[25]) );
NOR2_X2 U15919 ( .A1(n5547), .A2(n18005), .ZN(aes_text_in[24]) );
NOR2_X2 U15920 ( .A1(n5548), .A2(n18005), .ZN(aes_text_in[23]) );
NOR2_X2 U15921 ( .A1(n5549), .A2(n18005), .ZN(aes_text_in[22]) );
NOR2_X2 U15922 ( .A1(n5550), .A2(n18005), .ZN(aes_text_in[21]) );
NOR2_X2 U15923 ( .A1(n5551), .A2(n18004), .ZN(aes_text_in[20]) );
NOR2_X2 U15924 ( .A1(n5552), .A2(n18004), .ZN(aes_text_in[19]) );
NOR2_X2 U15925 ( .A1(n5553), .A2(n18004), .ZN(aes_text_in[18]) );
NOR2_X2 U15926 ( .A1(n5554), .A2(n18004), .ZN(aes_text_in[17]) );
NOR2_X2 U15927 ( .A1(n5555), .A2(n18004), .ZN(aes_text_in[16]) );
NOR2_X2 U15928 ( .A1(n5556), .A2(n18004), .ZN(aes_text_in[15]) );
NOR2_X2 U15929 ( .A1(n5557), .A2(n18004), .ZN(aes_text_in[14]) );
NOR2_X2 U15930 ( .A1(n5558), .A2(n18004), .ZN(aes_text_in[13]) );
NOR2_X2 U15931 ( .A1(n5559), .A2(n18004), .ZN(aes_text_in[12]) );
NOR2_X2 U15932 ( .A1(n5560), .A2(n18004), .ZN(aes_text_in[11]) );
NOR2_X2 U15933 ( .A1(n5561), .A2(n18004), .ZN(aes_text_in[10]) );
NOR2_X2 U15934 ( .A1(n5562), .A2(n18003), .ZN(aes_text_in[9]) );
NOR2_X2 U15935 ( .A1(n5563), .A2(n18003), .ZN(aes_text_in[8]) );
NOR2_X2 U15936 ( .A1(n5564), .A2(n18003), .ZN(aes_text_in[7]) );
NOR2_X2 U15937 ( .A1(n5565), .A2(n18003), .ZN(aes_text_in[6]) );
NOR2_X2 U15938 ( .A1(n5566), .A2(n18003), .ZN(aes_text_in[5]) );
NOR2_X2 U15939 ( .A1(n5567), .A2(n18003), .ZN(aes_text_in[4]) );
NOR2_X2 U15940 ( .A1(n5568), .A2(n18003), .ZN(aes_text_in[3]) );
NOR2_X2 U15941 ( .A1(n5569), .A2(n18003), .ZN(aes_text_in[2]) );
NOR2_X2 U15942 ( .A1(n5570), .A2(n18003), .ZN(aes_text_in[1]) );
NOR2_X2 U15943 ( .A1(n5571), .A2(n18003), .ZN(aes_text_in[0]) );
NAND2_X2 U15944 ( .A1(n11955), .A2(n11929), .ZN(n11961) );
MUX2_X2 U15945 ( .A(enc_byte_cnt[60]), .B(N2409), .S(n17812), .Z(n5381) );
MUX2_X2 U15946 ( .A(enc_byte_cnt[59]), .B(N2408), .S(n17812), .Z(n5382) );
MUX2_X2 U15947 ( .A(enc_byte_cnt[58]), .B(N2407), .S(n17812), .Z(n5383) );
MUX2_X2 U15948 ( .A(enc_byte_cnt[57]), .B(N2406), .S(n17812), .Z(n5384) );
MUX2_X2 U15949 ( .A(enc_byte_cnt[56]), .B(N2405), .S(n17812), .Z(n5385) );
MUX2_X2 U15950 ( .A(enc_byte_cnt[55]), .B(N2404), .S(n17812), .Z(n5386) );
MUX2_X2 U15951 ( .A(enc_byte_cnt[54]), .B(N2403), .S(n17812), .Z(n5387) );
MUX2_X2 U15952 ( .A(enc_byte_cnt[53]), .B(N2402), .S(n17812), .Z(n5388) );
MUX2_X2 U15953 ( .A(enc_byte_cnt[52]), .B(N2401), .S(n17812), .Z(n5389) );
MUX2_X2 U15954 ( .A(enc_byte_cnt[51]), .B(N2400), .S(n17812), .Z(n5390) );
MUX2_X2 U15955 ( .A(enc_byte_cnt[50]), .B(N2399), .S(n17812), .Z(n5391) );
MUX2_X2 U15956 ( .A(enc_byte_cnt[49]), .B(N2398), .S(n17813), .Z(n5392) );
MUX2_X2 U15957 ( .A(enc_byte_cnt[48]), .B(N2397), .S(n17813), .Z(n5393) );
MUX2_X2 U15958 ( .A(enc_byte_cnt[47]), .B(N2396), .S(n17813), .Z(n5394) );
MUX2_X2 U15959 ( .A(enc_byte_cnt[46]), .B(N2395), .S(n17813), .Z(n5395) );
MUX2_X2 U15960 ( .A(enc_byte_cnt[45]), .B(N2394), .S(n17813), .Z(n5396) );
MUX2_X2 U15961 ( .A(enc_byte_cnt[44]), .B(N2393), .S(n17813), .Z(n5397) );
MUX2_X2 U15962 ( .A(enc_byte_cnt[43]), .B(N2392), .S(n17813), .Z(n5398) );
MUX2_X2 U15963 ( .A(enc_byte_cnt[42]), .B(N2391), .S(n17813), .Z(n5399) );
MUX2_X2 U15964 ( .A(enc_byte_cnt[41]), .B(N2390), .S(n17813), .Z(n5400) );
MUX2_X2 U15965 ( .A(enc_byte_cnt[40]), .B(N2389), .S(n17813), .Z(n5401) );
MUX2_X2 U15966 ( .A(enc_byte_cnt[39]), .B(N2388), .S(n17813), .Z(n5402) );
MUX2_X2 U15967 ( .A(enc_byte_cnt[38]), .B(N2387), .S(n17814), .Z(n5403) );
MUX2_X2 U15968 ( .A(enc_byte_cnt[37]), .B(N2386), .S(n17814), .Z(n5404) );
MUX2_X2 U15969 ( .A(enc_byte_cnt[36]), .B(N2385), .S(n17814), .Z(n5405) );
MUX2_X2 U15970 ( .A(enc_byte_cnt[35]), .B(N2384), .S(n17814), .Z(n5406) );
MUX2_X2 U15971 ( .A(enc_byte_cnt[34]), .B(N2383), .S(n17814), .Z(n5407) );
MUX2_X2 U15972 ( .A(enc_byte_cnt[33]), .B(N2382), .S(n17814), .Z(n5408) );
MUX2_X2 U15973 ( .A(enc_byte_cnt[32]), .B(N2381), .S(n17814), .Z(n5409) );
MUX2_X2 U15974 ( .A(enc_byte_cnt[31]), .B(N2380), .S(n17814), .Z(n5410) );
MUX2_X2 U15975 ( .A(enc_byte_cnt[30]), .B(N2379), .S(n17814), .Z(n5411) );
MUX2_X2 U15976 ( .A(enc_byte_cnt[29]), .B(N2378), .S(n17814), .Z(n5412) );
MUX2_X2 U15977 ( .A(enc_byte_cnt[28]), .B(N2377), .S(n17814), .Z(n5413) );
MUX2_X2 U15978 ( .A(enc_byte_cnt[27]), .B(N2376), .S(n17815), .Z(n5414) );
MUX2_X2 U15979 ( .A(enc_byte_cnt[26]), .B(N2375), .S(n17815), .Z(n5415) );
MUX2_X2 U15980 ( .A(enc_byte_cnt[25]), .B(N2374), .S(n17815), .Z(n5416) );
MUX2_X2 U15981 ( .A(enc_byte_cnt[24]), .B(N2373), .S(n17815), .Z(n5417) );
MUX2_X2 U15982 ( .A(enc_byte_cnt[23]), .B(N2372), .S(n17815), .Z(n5418) );
MUX2_X2 U15983 ( .A(enc_byte_cnt[22]), .B(N2371), .S(n17815), .Z(n5419) );
MUX2_X2 U15984 ( .A(enc_byte_cnt[21]), .B(N2370), .S(n17815), .Z(n5420) );
MUX2_X2 U15985 ( .A(enc_byte_cnt[20]), .B(N2369), .S(n17815), .Z(n5421) );
MUX2_X2 U15986 ( .A(enc_byte_cnt[19]), .B(N2368), .S(n17815), .Z(n5422) );
MUX2_X2 U15987 ( .A(enc_byte_cnt[18]), .B(N2367), .S(n17815), .Z(n5423) );
MUX2_X2 U15988 ( .A(enc_byte_cnt[17]), .B(N2366), .S(n17815), .Z(n5424) );
MUX2_X2 U15989 ( .A(enc_byte_cnt[16]), .B(N2365), .S(n17816), .Z(n5425) );
MUX2_X2 U15990 ( .A(enc_byte_cnt[15]), .B(N2364), .S(n17816), .Z(n5426) );
MUX2_X2 U15991 ( .A(enc_byte_cnt[14]), .B(N2363), .S(n17816), .Z(n5427) );
MUX2_X2 U15992 ( .A(enc_byte_cnt[13]), .B(N2362), .S(n17816), .Z(n5428) );
MUX2_X2 U15993 ( .A(enc_byte_cnt[12]), .B(N2361), .S(n17816), .Z(n5429) );
MUX2_X2 U15994 ( .A(enc_byte_cnt[11]), .B(N2360), .S(n17816), .Z(n5430) );
MUX2_X2 U15995 ( .A(enc_byte_cnt[10]), .B(N2359), .S(n17816), .Z(n5431) );
MUX2_X2 U15996 ( .A(enc_byte_cnt[9]), .B(N2358), .S(n17816), .Z(n5432) );
MUX2_X2 U15997 ( .A(enc_byte_cnt[8]), .B(N2357), .S(n17816), .Z(n5433) );
MUX2_X2 U15998 ( .A(enc_byte_cnt[7]), .B(N2356), .S(n17816), .Z(n5434) );
MUX2_X2 U15999 ( .A(enc_byte_cnt[6]), .B(N2355), .S(n17816), .Z(n5435) );
MUX2_X2 U16000 ( .A(enc_byte_cnt[5]), .B(N2354), .S(n17817), .Z(n5436) );
MUX2_X2 U16001 ( .A(enc_byte_cnt[4]), .B(N2353), .S(n17817), .Z(n5437) );
MUX2_X2 U16002 ( .A(enc_byte_cnt[3]), .B(N2352), .S(n17817), .Z(n5438) );
MUX2_X2 U16003 ( .A(enc_byte_cnt[2]), .B(N2351), .S(n17817), .Z(n5439) );
NOR2_X2 U16004 ( .A1(n5378), .A2(n18002), .ZN(n18603) );
NOR3_X2 U16005 ( .A1(n16566), .A2(n18638), .A3(n18603), .ZN(n16565) );
NOR2_X2 U16006 ( .A1(n5377), .A2(n18002), .ZN(n18604) );
NOR3_X2 U16007 ( .A1(n16561), .A2(n18639), .A3(n18604), .ZN(n16560) );
NOR2_X2 U16008 ( .A1(n5376), .A2(n18002), .ZN(n18605) );
NOR3_X2 U16009 ( .A1(n16556), .A2(n18640), .A3(n18605), .ZN(n16555) );
NOR2_X2 U16010 ( .A1(n5375), .A2(n18002), .ZN(n18606) );
NOR3_X2 U16011 ( .A1(n16551), .A2(n18641), .A3(n18606), .ZN(n16550) );
NOR2_X2 U16012 ( .A1(n5328), .A2(n18002), .ZN(n15852) );
NOR2_X2 U16013 ( .A1(n5327), .A2(n18002), .ZN(n15834) );
NOR2_X2 U16014 ( .A1(n5326), .A2(n18002), .ZN(n15816) );
NAND2_X2 U16015 ( .A1(n17996), .A2(enc_byte_cnt[53]), .ZN(n15807) );
NAND2_X2 U16016 ( .A1(n17999), .A2(enc_byte_cnt[54]), .ZN(n15786) );
NAND2_X2 U16017 ( .A1(n17283), .A2(enc_byte_cnt[55]), .ZN(n15767) );
NAND2_X2 U16018 ( .A1(n17999), .A2(enc_byte_cnt[56]), .ZN(n15748) );
NAND2_X2 U16019 ( .A1(n17999), .A2(enc_byte_cnt[57]), .ZN(n15729) );
NAND2_X2 U16020 ( .A1(n17999), .A2(enc_byte_cnt[58]), .ZN(n15710) );
NAND2_X2 U16021 ( .A1(n17999), .A2(enc_byte_cnt[59]), .ZN(n15691) );
NAND2_X2 U16022 ( .A1(n17999), .A2(enc_byte_cnt[60]), .ZN(n15672) );
MUX2_X2 U16023 ( .A(aad_byte_cnt[60]), .B(N2539), .S(n17840), .Z(n5960) );
MUX2_X2 U16024 ( .A(aad_byte_cnt[59]), .B(N2538), .S(n17840), .Z(n5961) );
MUX2_X2 U16025 ( .A(aad_byte_cnt[58]), .B(N2537), .S(n17840), .Z(n5962) );
MUX2_X2 U16026 ( .A(aad_byte_cnt[57]), .B(N2536), .S(n17840), .Z(n5963) );
MUX2_X2 U16027 ( .A(aad_byte_cnt[56]), .B(N2535), .S(n17840), .Z(n5964) );
MUX2_X2 U16028 ( .A(aad_byte_cnt[55]), .B(N2534), .S(n17840), .Z(n5965) );
MUX2_X2 U16029 ( .A(aad_byte_cnt[54]), .B(N2533), .S(n17840), .Z(n5966) );
MUX2_X2 U16030 ( .A(aad_byte_cnt[53]), .B(N2532), .S(n17840), .Z(n5967) );
MUX2_X2 U16031 ( .A(aad_byte_cnt[52]), .B(N2531), .S(n17840), .Z(n5968) );
MUX2_X2 U16032 ( .A(aad_byte_cnt[51]), .B(N2530), .S(n17840), .Z(n5969) );
MUX2_X2 U16033 ( .A(aad_byte_cnt[50]), .B(N2529), .S(n17840), .Z(n5970) );
MUX2_X2 U16034 ( .A(aad_byte_cnt[49]), .B(N2528), .S(n17840), .Z(n5971) );
MUX2_X2 U16035 ( .A(aad_byte_cnt[48]), .B(N2527), .S(n17840), .Z(n5972) );
MUX2_X2 U16036 ( .A(aad_byte_cnt[47]), .B(N2526), .S(n17840), .Z(n5973) );
MUX2_X2 U16037 ( .A(aad_byte_cnt[46]), .B(N2525), .S(n17839), .Z(n5974) );
MUX2_X2 U16038 ( .A(aad_byte_cnt[45]), .B(N2524), .S(n17839), .Z(n5975) );
MUX2_X2 U16039 ( .A(aad_byte_cnt[44]), .B(N2523), .S(n17839), .Z(n5976) );
MUX2_X2 U16040 ( .A(aad_byte_cnt[43]), .B(N2522), .S(n17839), .Z(n5977) );
MUX2_X2 U16041 ( .A(aad_byte_cnt[42]), .B(N2521), .S(n17839), .Z(n5978) );
MUX2_X2 U16042 ( .A(aad_byte_cnt[41]), .B(N2520), .S(n17839), .Z(n5979) );
MUX2_X2 U16043 ( .A(aad_byte_cnt[40]), .B(N2519), .S(n17839), .Z(n5980) );
MUX2_X2 U16044 ( .A(aad_byte_cnt[39]), .B(N2518), .S(n17839), .Z(n5981) );
MUX2_X2 U16045 ( .A(aad_byte_cnt[38]), .B(N2517), .S(n17839), .Z(n5982) );
MUX2_X2 U16046 ( .A(aad_byte_cnt[37]), .B(N2516), .S(n17839), .Z(n5983) );
MUX2_X2 U16047 ( .A(aad_byte_cnt[36]), .B(N2515), .S(n17839), .Z(n5984) );
MUX2_X2 U16048 ( .A(aad_byte_cnt[35]), .B(N2514), .S(n17839), .Z(n5985) );
MUX2_X2 U16049 ( .A(aad_byte_cnt[34]), .B(N2513), .S(n17839), .Z(n5986) );
MUX2_X2 U16050 ( .A(aad_byte_cnt[33]), .B(N2512), .S(n17839), .Z(n5987) );
MUX2_X2 U16051 ( .A(aad_byte_cnt[32]), .B(N2511), .S(n17839), .Z(n5988) );
MUX2_X2 U16052 ( .A(aad_byte_cnt[31]), .B(N2510), .S(n17839), .Z(n5989) );
MUX2_X2 U16053 ( .A(aad_byte_cnt[30]), .B(N2509), .S(n17839), .Z(n5990) );
MUX2_X2 U16054 ( .A(aad_byte_cnt[29]), .B(N2508), .S(n17838), .Z(n5991) );
MUX2_X2 U16055 ( .A(aad_byte_cnt[28]), .B(N2507), .S(n17838), .Z(n5992) );
MUX2_X2 U16056 ( .A(aad_byte_cnt[27]), .B(N2506), .S(n17838), .Z(n5993) );
MUX2_X2 U16057 ( .A(aad_byte_cnt[26]), .B(N2505), .S(n17838), .Z(n5994) );
MUX2_X2 U16058 ( .A(aad_byte_cnt[25]), .B(N2504), .S(n17838), .Z(n5995) );
MUX2_X2 U16059 ( .A(aad_byte_cnt[24]), .B(N2503), .S(n17838), .Z(n5996) );
MUX2_X2 U16060 ( .A(aad_byte_cnt[23]), .B(N2502), .S(n17838), .Z(n5997) );
MUX2_X2 U16061 ( .A(aad_byte_cnt[22]), .B(N2501), .S(n17838), .Z(n5998) );
MUX2_X2 U16062 ( .A(aad_byte_cnt[21]), .B(N2500), .S(n17838), .Z(n5999) );
MUX2_X2 U16063 ( .A(aad_byte_cnt[20]), .B(N2499), .S(n17838), .Z(n6000) );
MUX2_X2 U16064 ( .A(aad_byte_cnt[19]), .B(N2498), .S(n17838), .Z(n6001) );
MUX2_X2 U16065 ( .A(aad_byte_cnt[18]), .B(N2497), .S(n17838), .Z(n6002) );
MUX2_X2 U16066 ( .A(aad_byte_cnt[17]), .B(N2496), .S(n17838), .Z(n6003) );
MUX2_X2 U16067 ( .A(aad_byte_cnt[16]), .B(N2495), .S(n17838), .Z(n6004) );
MUX2_X2 U16068 ( .A(aad_byte_cnt[15]), .B(N2494), .S(n17838), .Z(n6005) );
MUX2_X2 U16069 ( .A(aad_byte_cnt[14]), .B(N2493), .S(n17838), .Z(n6006) );
MUX2_X2 U16070 ( .A(aad_byte_cnt[13]), .B(N2492), .S(n17838), .Z(n6007) );
MUX2_X2 U16071 ( .A(aad_byte_cnt[12]), .B(N2491), .S(n17837), .Z(n6008) );
MUX2_X2 U16072 ( .A(aad_byte_cnt[11]), .B(N2490), .S(n17837), .Z(n6009) );
MUX2_X2 U16073 ( .A(aad_byte_cnt[10]), .B(N2489), .S(n17837), .Z(n6010) );
MUX2_X2 U16074 ( .A(aad_byte_cnt[9]), .B(N2488), .S(n17837), .Z(n6011) );
MUX2_X2 U16075 ( .A(aad_byte_cnt[8]), .B(N2487), .S(n17837), .Z(n6012) );
MUX2_X2 U16076 ( .A(aad_byte_cnt[7]), .B(N2486), .S(n17837), .Z(n6013) );
MUX2_X2 U16077 ( .A(aad_byte_cnt[6]), .B(N2485), .S(n17837), .Z(n6014) );
MUX2_X2 U16078 ( .A(aad_byte_cnt[5]), .B(N2484), .S(n17837), .Z(n6015) );
MUX2_X2 U16079 ( .A(aad_byte_cnt[4]), .B(N2483), .S(n17837), .Z(n6016) );
MUX2_X2 U16080 ( .A(aad_byte_cnt[3]), .B(N2482), .S(n17837), .Z(n6017) );
MUX2_X2 U16081 ( .A(aad_byte_cnt[2]), .B(N2481), .S(n17837), .Z(n6018) );
MUX2_X2 U16082 ( .A(aad_byte_cnt[0]), .B(N2479), .S(n17837), .Z(n6020) );
NAND2_X2 U16083 ( .A1(n17999), .A2(aad_byte_cnt[0]), .ZN(n18607) );
NAND2_X2 U16084 ( .A1(n15595), .A2(n18607), .ZN(n15580) );
NAND2_X2 U16085 ( .A1(n17999), .A2(aad_byte_cnt[1]), .ZN(n18608) );
NAND2_X2 U16086 ( .A1(n15574), .A2(n18608), .ZN(n15559) );
NAND2_X2 U16087 ( .A1(n17999), .A2(aad_byte_cnt[2]), .ZN(n18609) );
NAND2_X2 U16088 ( .A1(n15553), .A2(n18609), .ZN(n15538) );
NAND2_X2 U16089 ( .A1(n17999), .A2(aad_byte_cnt[3]), .ZN(n18610) );
NAND2_X2 U16090 ( .A1(n15532), .A2(n18610), .ZN(n15517) );
NAND2_X2 U16091 ( .A1(aad_byte_cnt[50]), .A2(n17283), .ZN(n14455) );
NAND2_X2 U16092 ( .A1(aad_byte_cnt[51]), .A2(n17283), .ZN(n14433) );
NAND2_X2 U16093 ( .A1(aad_byte_cnt[52]), .A2(n17283), .ZN(n14409) );
NAND2_X2 U16094 ( .A1(aad_byte_cnt[53]), .A2(n17283), .ZN(n14370) );
NAND2_X2 U16095 ( .A1(aad_byte_cnt[54]), .A2(n17283), .ZN(n14341) );
NAND2_X2 U16096 ( .A1(aad_byte_cnt[55]), .A2(n17283), .ZN(n14312) );
NAND2_X2 U16097 ( .A1(aad_byte_cnt[56]), .A2(n17283), .ZN(n14283) );
NAND2_X2 U16098 ( .A1(aad_byte_cnt[57]), .A2(n17283), .ZN(n14254) );
NAND2_X2 U16099 ( .A1(aad_byte_cnt[58]), .A2(n17283), .ZN(n14225) );
NAND2_X2 U16100 ( .A1(aad_byte_cnt[59]), .A2(n17283), .ZN(n14196) );
NAND2_X2 U16101 ( .A1(aad_byte_cnt[60]), .A2(n17283), .ZN(n14162) );
NOR3_X2 U16102 ( .A1(n14157), .A2(state[1]), .A3(n18611), .ZN(n14155) );
NAND2_X2 U16103 ( .A1(n18892), .A2(n18044), .ZN(n11924) );
INV_X4 U16104 ( .A(n11924), .ZN(n18623) );
NAND2_X2 U16105 ( .A1(n6850), .A2(n18623), .ZN(n11937) );
INV_X4 U16106 ( .A(n11937), .ZN(n18612) );
NAND2_X2 U16107 ( .A1(n18612), .A2(n18622), .ZN(n18614) );
NAND2_X2 U16108 ( .A1(n17280), .A2(n18624), .ZN(n18613) );
NAND2_X2 U16109 ( .A1(n18614), .A2(n18613), .ZN(n6291) );
NAND3_X2 U16110 ( .A1(n18630), .A2(aes_done), .A3(n17290), .ZN(n18633) );
NAND2_X2 U16111 ( .A1(n17290), .A2(n18630), .ZN(n18615) );
NAND2_X2 U16112 ( .A1(n11976), .A2(n18615), .ZN(n18621) );
INV_X4 U16113 ( .A(n18621), .ZN(n18844) );
NOR4_X2 U16114 ( .A1(n11967), .A2(n11955), .A3(n11971), .A4(n17996), .ZN(n11970) );
NAND2_X2 U16115 ( .A1(n11968), .A2(n11967), .ZN(n11965) );
NAND2_X2 U16116 ( .A1(n18846), .A2(n18892), .ZN(n11966) );
INV_X4 U16117 ( .A(dii_data_vld), .ZN(n18616) );
NAND2_X2 U16118 ( .A1(n18617), .A2(n18616), .ZN(n18619) );
NAND2_X2 U16119 ( .A1(n19206), .A2(n11971), .ZN(n18618) );
NAND2_X2 U16120 ( .A1(n11960), .A2(state[2]), .ZN(n11959) );
NAND2_X2 U16121 ( .A1(n18747), .A2(n17375), .ZN(n18620) );
NAND2_X2 U16122 ( .A1(state[4]), .A2(n18620), .ZN(n11950) );
NAND2_X2 U16123 ( .A1(n11948), .A2(state[5]), .ZN(n11947) );
NAND2_X2 U16124 ( .A1(n18746), .A2(n18621), .ZN(n11944) );
NAND2_X2 U16125 ( .A1(n11926), .A2(state[3]), .ZN(n11943) );
NAND2_X2 U16126 ( .A1(state[7]), .A2(n11926), .ZN(n11940) );
NAND3_X2 U16127 ( .A1(n16838), .A2(n17291), .A3(n18624), .ZN(n11936) );
NAND2_X2 U16128 ( .A1(n11926), .A2(state[1]), .ZN(n11931) );
NAND2_X2 U16129 ( .A1(state[8]), .A2(n11926), .ZN(n11927) );
INV_X4 U16130 ( .A(n16839), .ZN(n18894) );
MUX2_X2 U16131 ( .A(aad_byte_cnt[62]), .B(N2541), .S(n17837), .Z(n5958) );
MUX2_X2 U16132 ( .A(aad_byte_cnt[61]), .B(N2540), .S(n17837), .Z(n5959) );
MUX2_X2 U16133 ( .A(aad_byte_cnt[63]), .B(N2542), .S(n17837), .Z(n6021) );
MUX2_X2 U16134 ( .A(enc_byte_cnt[62]), .B(N2411), .S(n17817), .Z(n5379) );
MUX2_X2 U16135 ( .A(enc_byte_cnt[61]), .B(N2410), .S(n17817), .Z(n5380) );
MUX2_X2 U16136 ( .A(enc_byte_cnt[63]), .B(N2412), .S(n17817), .Z(n5442) );
INV_X4 U16137 ( .A(n13280), .ZN(n18635) );
INV_X4 U16138 ( .A(n13287), .ZN(n18636) );
INV_X4 U16139 ( .A(n13292), .ZN(n18637) );
INV_X4 U16140 ( .A(n13297), .ZN(n18638) );
INV_X4 U16141 ( .A(n13302), .ZN(n18639) );
INV_X4 U16142 ( .A(n13307), .ZN(n18640) );
INV_X4 U16143 ( .A(n13312), .ZN(n18641) );
INV_X4 U16144 ( .A(n13317), .ZN(n18642) );
INV_X4 U16145 ( .A(n13370), .ZN(n18643) );
INV_X4 U16146 ( .A(n13376), .ZN(n18644) );
INV_X4 U16147 ( .A(n13382), .ZN(n18645) );
INV_X4 U16148 ( .A(n13388), .ZN(n18646) );
INV_X4 U16149 ( .A(n13394), .ZN(n18647) );
INV_X4 U16150 ( .A(n13400), .ZN(n18648) );
INV_X4 U16151 ( .A(n13406), .ZN(n18649) );
INV_X4 U16152 ( .A(n13412), .ZN(n18650) );
INV_X4 U16153 ( .A(n13418), .ZN(n18651) );
INV_X4 U16154 ( .A(n13424), .ZN(n18652) );
INV_X4 U16155 ( .A(n13430), .ZN(n18653) );
INV_X4 U16156 ( .A(n13436), .ZN(n18654) );
INV_X4 U16157 ( .A(n13442), .ZN(n18655) );
INV_X4 U16158 ( .A(n13448), .ZN(n18656) );
INV_X4 U16159 ( .A(n13454), .ZN(n18657) );
INV_X4 U16160 ( .A(n13460), .ZN(n18658) );
INV_X4 U16161 ( .A(n13466), .ZN(n18659) );
INV_X4 U16162 ( .A(n13472), .ZN(n18660) );
INV_X4 U16163 ( .A(n13478), .ZN(n18661) );
INV_X4 U16164 ( .A(n13484), .ZN(n18662) );
INV_X4 U16165 ( .A(n13490), .ZN(n18663) );
INV_X4 U16166 ( .A(n13496), .ZN(n18664) );
INV_X4 U16167 ( .A(n13502), .ZN(n18665) );
INV_X4 U16168 ( .A(n13508), .ZN(n18666) );
INV_X4 U16169 ( .A(n13514), .ZN(n18667) );
INV_X4 U16170 ( .A(n13520), .ZN(n18668) );
INV_X4 U16171 ( .A(n13526), .ZN(n18669) );
INV_X4 U16172 ( .A(n13532), .ZN(n18670) );
INV_X4 U16173 ( .A(n13538), .ZN(n18671) );
INV_X4 U16174 ( .A(n13544), .ZN(n18672) );
INV_X4 U16175 ( .A(n13550), .ZN(n18673) );
INV_X4 U16176 ( .A(n13556), .ZN(n18674) );
INV_X4 U16177 ( .A(n13562), .ZN(n18675) );
INV_X4 U16178 ( .A(n13568), .ZN(n18676) );
INV_X4 U16179 ( .A(n13574), .ZN(n18677) );
INV_X4 U16180 ( .A(n13580), .ZN(n18678) );
INV_X4 U16181 ( .A(n13586), .ZN(n18679) );
INV_X4 U16182 ( .A(n13592), .ZN(n18680) );
INV_X4 U16183 ( .A(n13598), .ZN(n18681) );
INV_X4 U16184 ( .A(n13604), .ZN(n18682) );
INV_X4 U16185 ( .A(n13610), .ZN(n18683) );
INV_X4 U16186 ( .A(n13616), .ZN(n18684) );
INV_X4 U16187 ( .A(n13622), .ZN(n18685) );
INV_X4 U16188 ( .A(n13628), .ZN(n18686) );
INV_X4 U16189 ( .A(n13634), .ZN(n18687) );
INV_X4 U16190 ( .A(n13640), .ZN(n18688) );
INV_X4 U16191 ( .A(n13646), .ZN(n18689) );
INV_X4 U16192 ( .A(n13652), .ZN(n18690) );
INV_X4 U16193 ( .A(n13680), .ZN(n18691) );
INV_X4 U16194 ( .A(n13686), .ZN(n18692) );
INV_X4 U16195 ( .A(n13692), .ZN(n18693) );
INV_X4 U16196 ( .A(n13698), .ZN(n18694) );
INV_X4 U16197 ( .A(n13704), .ZN(n18695) );
INV_X4 U16198 ( .A(n13710), .ZN(n18696) );
INV_X4 U16199 ( .A(n13716), .ZN(n18697) );
INV_X4 U16200 ( .A(n13722), .ZN(n18698) );
INV_X4 U16201 ( .A(n13728), .ZN(n18699) );
INV_X4 U16202 ( .A(n13734), .ZN(n18700) );
INV_X4 U16203 ( .A(n13740), .ZN(n18701) );
INV_X4 U16204 ( .A(n13746), .ZN(n18702) );
INV_X4 U16205 ( .A(n13752), .ZN(n18703) );
INV_X4 U16206 ( .A(n13758), .ZN(n18704) );
INV_X4 U16207 ( .A(n13764), .ZN(n18705) );
INV_X4 U16208 ( .A(n13770), .ZN(n18706) );
INV_X4 U16209 ( .A(n13776), .ZN(n18707) );
INV_X4 U16210 ( .A(n13782), .ZN(n18708) );
INV_X4 U16211 ( .A(n13788), .ZN(n18709) );
INV_X4 U16212 ( .A(n13794), .ZN(n18710) );
INV_X4 U16213 ( .A(n13800), .ZN(n18711) );
INV_X4 U16214 ( .A(n13806), .ZN(n18712) );
INV_X4 U16215 ( .A(n13812), .ZN(n18713) );
INV_X4 U16216 ( .A(n13818), .ZN(n18714) );
INV_X4 U16217 ( .A(n13824), .ZN(n18715) );
INV_X4 U16218 ( .A(n13830), .ZN(n18716) );
INV_X4 U16219 ( .A(n13836), .ZN(n18717) );
INV_X4 U16220 ( .A(n13842), .ZN(n18718) );
INV_X4 U16221 ( .A(n13848), .ZN(n18719) );
INV_X4 U16222 ( .A(n13854), .ZN(n18720) );
INV_X4 U16223 ( .A(n13860), .ZN(n18721) );
INV_X4 U16224 ( .A(n13866), .ZN(n18722) );
INV_X4 U16225 ( .A(n13872), .ZN(n18723) );
INV_X4 U16226 ( .A(n13878), .ZN(n18724) );
INV_X4 U16227 ( .A(n13884), .ZN(n18725) );
INV_X4 U16228 ( .A(n13890), .ZN(n18726) );
INV_X4 U16229 ( .A(n13896), .ZN(n18727) );
INV_X4 U16230 ( .A(n13902), .ZN(n18728) );
INV_X4 U16231 ( .A(n13908), .ZN(n18729) );
INV_X4 U16232 ( .A(n13914), .ZN(n18730) );
INV_X4 U16233 ( .A(n13920), .ZN(n18731) );
INV_X4 U16234 ( .A(n13926), .ZN(n18732) );
INV_X4 U16235 ( .A(n13932), .ZN(n18733) );
INV_X4 U16236 ( .A(n13938), .ZN(n18734) );
INV_X4 U16237 ( .A(n13944), .ZN(n18735) );
INV_X4 U16238 ( .A(n13950), .ZN(n18736) );
INV_X4 U16239 ( .A(n13956), .ZN(n18737) );
INV_X4 U16240 ( .A(n13962), .ZN(n18738) );
INV_X4 U16241 ( .A(n13968), .ZN(n18739) );
INV_X4 U16242 ( .A(n13974), .ZN(n18740) );
INV_X4 U16243 ( .A(n13980), .ZN(n18741) );
INV_X4 U16244 ( .A(n13986), .ZN(n18742) );
INV_X4 U16245 ( .A(n13992), .ZN(n18743) );
INV_X4 U16246 ( .A(n17281), .ZN(n18744) );
INV_X4 U16247 ( .A(n17280), .ZN(n18745) );
INV_X4 U16248 ( .A(aes_done), .ZN(n18746) );
INV_X4 U16249 ( .A(n11948), .ZN(n18747) );
INV_X4 U16250 ( .A(aes_text_out[127]), .ZN(n18748) );
INV_X4 U16251 ( .A(aes_text_out[126]), .ZN(n18749) );
INV_X4 U16252 ( .A(aes_text_out[125]), .ZN(n18750) );
INV_X4 U16253 ( .A(aes_text_out[124]), .ZN(n18751) );
INV_X4 U16254 ( .A(aes_text_out[123]), .ZN(n18752) );
INV_X4 U16255 ( .A(aes_text_out[122]), .ZN(n18753) );
INV_X4 U16256 ( .A(aes_text_out[121]), .ZN(n18754) );
INV_X4 U16257 ( .A(aes_text_out[120]), .ZN(n18755) );
INV_X4 U16258 ( .A(n13994), .ZN(n18756) );
INV_X4 U16259 ( .A(n13988), .ZN(n18757) );
INV_X4 U16260 ( .A(n13982), .ZN(n18758) );
INV_X4 U16261 ( .A(n13976), .ZN(n18759) );
INV_X4 U16262 ( .A(n13970), .ZN(n18760) );
INV_X4 U16263 ( .A(n13964), .ZN(n18761) );
INV_X4 U16264 ( .A(n13958), .ZN(n18762) );
INV_X4 U16265 ( .A(n13952), .ZN(n18763) );
INV_X4 U16266 ( .A(n13946), .ZN(n18764) );
INV_X4 U16267 ( .A(n13940), .ZN(n18765) );
INV_X4 U16268 ( .A(n13934), .ZN(n18766) );
INV_X4 U16269 ( .A(n13928), .ZN(n18767) );
INV_X4 U16270 ( .A(n13922), .ZN(n18768) );
INV_X4 U16271 ( .A(n13916), .ZN(n18769) );
INV_X4 U16272 ( .A(n13910), .ZN(n18770) );
INV_X4 U16273 ( .A(n13904), .ZN(n18771) );
INV_X4 U16274 ( .A(n13898), .ZN(n18772) );
INV_X4 U16275 ( .A(n13892), .ZN(n18773) );
INV_X4 U16276 ( .A(n13886), .ZN(n18774) );
INV_X4 U16277 ( .A(n13880), .ZN(n18775) );
INV_X4 U16278 ( .A(n13874), .ZN(n18776) );
INV_X4 U16279 ( .A(n13868), .ZN(n18777) );
INV_X4 U16280 ( .A(n13862), .ZN(n18778) );
INV_X4 U16281 ( .A(n13856), .ZN(n18779) );
INV_X4 U16282 ( .A(n13850), .ZN(n18780) );
INV_X4 U16283 ( .A(n13844), .ZN(n18781) );
INV_X4 U16284 ( .A(n13838), .ZN(n18782) );
INV_X4 U16285 ( .A(n13832), .ZN(n18783) );
INV_X4 U16286 ( .A(n13826), .ZN(n18784) );
INV_X4 U16287 ( .A(n13820), .ZN(n18785) );
INV_X4 U16288 ( .A(n13814), .ZN(n18786) );
INV_X4 U16289 ( .A(n13808), .ZN(n18787) );
INV_X4 U16290 ( .A(n13802), .ZN(n18788) );
INV_X4 U16291 ( .A(n13796), .ZN(n18789) );
INV_X4 U16292 ( .A(n13790), .ZN(n18790) );
INV_X4 U16293 ( .A(n13784), .ZN(n18791) );
INV_X4 U16294 ( .A(n13778), .ZN(n18792) );
INV_X4 U16295 ( .A(n13772), .ZN(n18793) );
INV_X4 U16296 ( .A(n13766), .ZN(n18794) );
INV_X4 U16297 ( .A(n13760), .ZN(n18795) );
INV_X4 U16298 ( .A(n13754), .ZN(n18796) );
INV_X4 U16299 ( .A(n13748), .ZN(n18797) );
INV_X4 U16300 ( .A(n13742), .ZN(n18798) );
INV_X4 U16301 ( .A(n13736), .ZN(n18799) );
INV_X4 U16302 ( .A(n13730), .ZN(n18800) );
INV_X4 U16303 ( .A(n13724), .ZN(n18801) );
INV_X4 U16304 ( .A(n13718), .ZN(n18802) );
INV_X4 U16305 ( .A(n13712), .ZN(n18803) );
INV_X4 U16306 ( .A(n13706), .ZN(n18804) );
INV_X4 U16307 ( .A(n13700), .ZN(n18805) );
INV_X4 U16308 ( .A(n13694), .ZN(n18806) );
INV_X4 U16309 ( .A(n13688), .ZN(n18807) );
INV_X4 U16310 ( .A(n13682), .ZN(n18808) );
INV_X4 U16311 ( .A(n13676), .ZN(n18809) );
INV_X4 U16312 ( .A(n13669), .ZN(n18810) );
INV_X4 U16313 ( .A(n13662), .ZN(n18811) );
INV_X4 U16314 ( .A(n13654), .ZN(n18812) );
INV_X4 U16315 ( .A(n13648), .ZN(n18813) );
INV_X4 U16316 ( .A(n13642), .ZN(n18814) );
INV_X4 U16317 ( .A(n13636), .ZN(n18815) );
INV_X4 U16318 ( .A(n13630), .ZN(n18816) );
INV_X4 U16319 ( .A(n13624), .ZN(n18817) );
INV_X4 U16320 ( .A(n13618), .ZN(n18818) );
INV_X4 U16321 ( .A(n13612), .ZN(n18819) );
INV_X4 U16322 ( .A(n13558), .ZN(n18820) );
INV_X4 U16323 ( .A(n13552), .ZN(n18821) );
INV_X4 U16324 ( .A(n13546), .ZN(n18822) );
INV_X4 U16325 ( .A(n13540), .ZN(n18823) );
INV_X4 U16326 ( .A(n13534), .ZN(n18824) );
INV_X4 U16327 ( .A(n13528), .ZN(n18825) );
INV_X4 U16328 ( .A(n13522), .ZN(n18826) );
INV_X4 U16329 ( .A(n13516), .ZN(n18827) );
INV_X4 U16330 ( .A(n13462), .ZN(n18828) );
INV_X4 U16331 ( .A(n13456), .ZN(n18829) );
INV_X4 U16332 ( .A(n13450), .ZN(n18830) );
INV_X4 U16333 ( .A(n13444), .ZN(n18831) );
INV_X4 U16334 ( .A(n13438), .ZN(n18832) );
INV_X4 U16335 ( .A(n13432), .ZN(n18833) );
INV_X4 U16336 ( .A(n13426), .ZN(n18834) );
INV_X4 U16337 ( .A(n13420), .ZN(n18835) );
INV_X4 U16338 ( .A(aes_text_out[15]), .ZN(n18836) );
INV_X4 U16339 ( .A(aes_text_out[14]), .ZN(n18837) );
INV_X4 U16340 ( .A(aes_text_out[13]), .ZN(n18838) );
INV_X4 U16341 ( .A(aes_text_out[12]), .ZN(n18839) );
INV_X4 U16342 ( .A(aes_text_out[11]), .ZN(n18840) );
INV_X4 U16343 ( .A(aes_text_out[10]), .ZN(n18841) );
INV_X4 U16344 ( .A(aes_text_out[9]), .ZN(n18842) );
INV_X4 U16345 ( .A(aes_text_out[8]), .ZN(n18843) );
INV_X4 U16346 ( .A(n16837), .ZN(n18845) );
INV_X4 U16347 ( .A(n11957), .ZN(n18846) );
INV_X4 U16348 ( .A(n11929), .ZN(n18892) );
INV_X4 U16349 ( .A(n14166), .ZN(n19023) );
INV_X4 U16350 ( .A(n14199), .ZN(n19024) );
INV_X4 U16351 ( .A(n14228), .ZN(n19025) );
INV_X4 U16352 ( .A(n14257), .ZN(n19026) );
INV_X4 U16353 ( .A(n14286), .ZN(n19027) );
INV_X4 U16354 ( .A(n14315), .ZN(n19028) );
INV_X4 U16355 ( .A(n14344), .ZN(n19029) );
INV_X4 U16356 ( .A(n14373), .ZN(n19030) );
INV_X4 U16357 ( .A(n14190), .ZN(n19031) );
INV_X4 U16358 ( .A(n17539), .ZN(n19032) );
INV_X4 U16359 ( .A(n14219), .ZN(n19033) );
INV_X4 U16360 ( .A(n17541), .ZN(n19034) );
INV_X4 U16361 ( .A(n14248), .ZN(n19035) );
INV_X4 U16362 ( .A(n17543), .ZN(n19036) );
INV_X4 U16363 ( .A(n14277), .ZN(n19037) );
INV_X4 U16364 ( .A(n17545), .ZN(n19038) );
INV_X4 U16365 ( .A(n14306), .ZN(n19039) );
INV_X4 U16366 ( .A(n17547), .ZN(n19040) );
INV_X4 U16367 ( .A(n14335), .ZN(n19041) );
INV_X4 U16368 ( .A(n17549), .ZN(n19042) );
INV_X4 U16369 ( .A(n14364), .ZN(n19043) );
INV_X4 U16370 ( .A(n17551), .ZN(n19044) );
INV_X4 U16371 ( .A(n14396), .ZN(n19045) );
INV_X4 U16372 ( .A(n17553), .ZN(n19046) );
INV_X4 U16373 ( .A(n14191), .ZN(n19047) );
INV_X4 U16374 ( .A(n17555), .ZN(n19048) );
INV_X4 U16375 ( .A(n14220), .ZN(n19049) );
INV_X4 U16376 ( .A(n17557), .ZN(n19050) );
INV_X4 U16377 ( .A(n14249), .ZN(n19051) );
INV_X4 U16378 ( .A(n17559), .ZN(n19052) );
INV_X4 U16379 ( .A(n14278), .ZN(n19053) );
INV_X4 U16380 ( .A(n17561), .ZN(n19054) );
INV_X4 U16381 ( .A(n14307), .ZN(n19055) );
INV_X4 U16382 ( .A(n17563), .ZN(n19056) );
INV_X4 U16383 ( .A(n14336), .ZN(n19057) );
INV_X4 U16384 ( .A(n17745), .ZN(n19058) );
INV_X4 U16385 ( .A(n14365), .ZN(n19059) );
INV_X4 U16386 ( .A(n17565), .ZN(n19060) );
INV_X4 U16387 ( .A(n14397), .ZN(n19061) );
INV_X4 U16388 ( .A(n17567), .ZN(n19062) );
INV_X4 U16389 ( .A(n14417), .ZN(n19063) );
INV_X4 U16390 ( .A(n17569), .ZN(n19064) );
INV_X4 U16391 ( .A(n14440), .ZN(n19065) );
INV_X4 U16392 ( .A(n17571), .ZN(n19066) );
INV_X4 U16393 ( .A(n14462), .ZN(n19067) );
INV_X4 U16394 ( .A(n17573), .ZN(n19068) );
INV_X4 U16395 ( .A(n14484), .ZN(n19069) );
INV_X4 U16396 ( .A(n17575), .ZN(n19070) );
INV_X4 U16397 ( .A(n14506), .ZN(n19071) );
INV_X4 U16398 ( .A(n17577), .ZN(n19072) );
INV_X4 U16399 ( .A(n14528), .ZN(n19073) );
INV_X4 U16400 ( .A(n17579), .ZN(n19074) );
INV_X4 U16401 ( .A(n14550), .ZN(n19075) );
INV_X4 U16402 ( .A(n17581), .ZN(n19076) );
INV_X4 U16403 ( .A(n14574), .ZN(n19077) );
INV_X4 U16404 ( .A(n17583), .ZN(n19078) );
INV_X4 U16405 ( .A(n14185), .ZN(n19079) );
INV_X4 U16406 ( .A(n14597), .ZN(n19080) );
INV_X4 U16407 ( .A(n17585), .ZN(n19081) );
INV_X4 U16408 ( .A(n14216), .ZN(n19082) );
INV_X4 U16409 ( .A(n14618), .ZN(n19083) );
INV_X4 U16410 ( .A(n17587), .ZN(n19084) );
INV_X4 U16411 ( .A(n14245), .ZN(n19085) );
INV_X4 U16412 ( .A(n14639), .ZN(n19086) );
INV_X4 U16413 ( .A(n17589), .ZN(n19087) );
INV_X4 U16414 ( .A(n14274), .ZN(n19088) );
INV_X4 U16415 ( .A(n14660), .ZN(n19089) );
INV_X4 U16416 ( .A(n17591), .ZN(n19090) );
INV_X4 U16417 ( .A(n14303), .ZN(n19091) );
INV_X4 U16418 ( .A(n14681), .ZN(n19092) );
INV_X4 U16419 ( .A(n17593), .ZN(n19093) );
INV_X4 U16420 ( .A(n14332), .ZN(n19094) );
INV_X4 U16421 ( .A(n14702), .ZN(n19095) );
INV_X4 U16422 ( .A(n17595), .ZN(n19096) );
INV_X4 U16423 ( .A(n14361), .ZN(n19097) );
INV_X4 U16424 ( .A(n14723), .ZN(n19098) );
INV_X4 U16425 ( .A(n17597), .ZN(n19099) );
INV_X4 U16426 ( .A(n14391), .ZN(n19100) );
INV_X4 U16427 ( .A(n14746), .ZN(n19101) );
INV_X4 U16428 ( .A(n17599), .ZN(n19102) );
INV_X4 U16429 ( .A(n14421), .ZN(n19103) );
INV_X4 U16430 ( .A(n14768), .ZN(n19104) );
INV_X4 U16431 ( .A(n17601), .ZN(n19105) );
INV_X4 U16432 ( .A(n14444), .ZN(n19106) );
INV_X4 U16433 ( .A(n14791), .ZN(n19107) );
INV_X4 U16434 ( .A(n17603), .ZN(n19108) );
INV_X4 U16435 ( .A(n14466), .ZN(n19109) );
INV_X4 U16436 ( .A(n14813), .ZN(n19110) );
INV_X4 U16437 ( .A(n17605), .ZN(n19111) );
INV_X4 U16438 ( .A(n14488), .ZN(n19112) );
INV_X4 U16439 ( .A(n14835), .ZN(n19113) );
INV_X4 U16440 ( .A(n17607), .ZN(n19114) );
INV_X4 U16441 ( .A(n14510), .ZN(n19115) );
INV_X4 U16442 ( .A(n14857), .ZN(n19116) );
INV_X4 U16443 ( .A(n17609), .ZN(n19117) );
INV_X4 U16444 ( .A(n14532), .ZN(n19118) );
INV_X4 U16445 ( .A(n14879), .ZN(n19119) );
INV_X4 U16446 ( .A(n17611), .ZN(n19120) );
INV_X4 U16447 ( .A(n14554), .ZN(n19121) );
INV_X4 U16448 ( .A(n14901), .ZN(n19122) );
INV_X4 U16449 ( .A(n17613), .ZN(n19123) );
INV_X4 U16450 ( .A(n14578), .ZN(n19124) );
INV_X4 U16451 ( .A(n14924), .ZN(n19125) );
INV_X4 U16452 ( .A(n17615), .ZN(n19126) );
INV_X4 U16453 ( .A(n14773), .ZN(n19127) );
INV_X4 U16454 ( .A(n14795), .ZN(n19128) );
INV_X4 U16455 ( .A(n14817), .ZN(n19129) );
INV_X4 U16456 ( .A(n14839), .ZN(n19130) );
INV_X4 U16457 ( .A(n14861), .ZN(n19131) );
INV_X4 U16458 ( .A(n14883), .ZN(n19132) );
INV_X4 U16459 ( .A(n14905), .ZN(n19133) );
INV_X4 U16460 ( .A(n14928), .ZN(n19134) );
INV_X4 U16461 ( .A(n17633), .ZN(n19135) );
INV_X4 U16462 ( .A(n17635), .ZN(n19136) );
INV_X4 U16463 ( .A(n17637), .ZN(n19137) );
INV_X4 U16464 ( .A(n17639), .ZN(n19138) );
INV_X4 U16465 ( .A(n17641), .ZN(n19139) );
INV_X4 U16466 ( .A(n17643), .ZN(n19140) );
INV_X4 U16467 ( .A(n17645), .ZN(n19141) );
INV_X4 U16468 ( .A(n17647), .ZN(n19142) );
INV_X4 U16469 ( .A(n17649), .ZN(n19143) );
INV_X4 U16470 ( .A(n17651), .ZN(n19144) );
INV_X4 U16471 ( .A(n17653), .ZN(n19145) );
INV_X4 U16472 ( .A(n17655), .ZN(n19146) );
INV_X4 U16473 ( .A(n17657), .ZN(n19147) );
INV_X4 U16474 ( .A(n17659), .ZN(n19148) );
INV_X4 U16475 ( .A(n17661), .ZN(n19149) );
INV_X4 U16476 ( .A(n17663), .ZN(n19150) );
INV_X4 U16477 ( .A(n17665), .ZN(n19151) );
INV_X4 U16478 ( .A(n17667), .ZN(n19152) );
INV_X4 U16479 ( .A(n17669), .ZN(n19153) );
INV_X4 U16480 ( .A(n17671), .ZN(n19154) );
INV_X4 U16481 ( .A(n17673), .ZN(n19155) );
INV_X4 U16482 ( .A(n17675), .ZN(n19156) );
INV_X4 U16483 ( .A(n17677), .ZN(n19157) );
INV_X4 U16484 ( .A(n17679), .ZN(n19158) );
INV_X4 U16485 ( .A(n17681), .ZN(n19159) );
INV_X4 U16486 ( .A(n17683), .ZN(n19160) );
INV_X4 U16487 ( .A(n17685), .ZN(n19161) );
INV_X4 U16488 ( .A(n17687), .ZN(n19162) );
INV_X4 U16489 ( .A(n17689), .ZN(n19163) );
INV_X4 U16490 ( .A(n17691), .ZN(n19164) );
INV_X4 U16491 ( .A(n17693), .ZN(n19165) );
INV_X4 U16492 ( .A(n17695), .ZN(n19166) );
INV_X4 U16493 ( .A(n17697), .ZN(n19167) );
INV_X4 U16494 ( .A(n17699), .ZN(n19168) );
INV_X4 U16495 ( .A(n17701), .ZN(n19169) );
INV_X4 U16496 ( .A(n17703), .ZN(n19170) );
INV_X4 U16497 ( .A(n17705), .ZN(n19171) );
INV_X4 U16498 ( .A(n17707), .ZN(n19172) );
INV_X4 U16499 ( .A(n17709), .ZN(n19173) );
INV_X4 U16500 ( .A(n17711), .ZN(n19174) );
INV_X4 U16501 ( .A(n17713), .ZN(n19175) );
INV_X4 U16502 ( .A(n17715), .ZN(n19176) );
INV_X4 U16503 ( .A(n17717), .ZN(n19177) );
INV_X4 U16504 ( .A(n17719), .ZN(n19178) );
INV_X4 U16505 ( .A(n17721), .ZN(n19179) );
INV_X4 U16506 ( .A(n17723), .ZN(n19180) );
INV_X4 U16507 ( .A(n17725), .ZN(n19181) );
INV_X4 U16508 ( .A(n17727), .ZN(n19182) );
INV_X4 U16509 ( .A(n17728), .ZN(n19183) );
INV_X4 U16510 ( .A(n17729), .ZN(n19184) );
INV_X4 U16511 ( .A(n17730), .ZN(n19185) );
INV_X4 U16512 ( .A(n17731), .ZN(n19186) );
INV_X4 U16513 ( .A(n17732), .ZN(n19187) );
INV_X4 U16514 ( .A(n17733), .ZN(n19188) );
INV_X4 U16515 ( .A(n17734), .ZN(n19189) );
INV_X4 U16516 ( .A(n17735), .ZN(n19190) );
INV_X4 U16517 ( .A(n17736), .ZN(n19191) );
INV_X4 U16518 ( .A(n17737), .ZN(n19192) );
INV_X4 U16519 ( .A(n17738), .ZN(n19193) );
INV_X4 U16520 ( .A(n17739), .ZN(n19194) );
INV_X4 U16521 ( .A(n17740), .ZN(n19195) );
INV_X4 U16522 ( .A(n17741), .ZN(n19196) );
INV_X4 U16523 ( .A(n17742), .ZN(n19197) );
INV_X4 U16524 ( .A(n17743), .ZN(n19198) );
INV_X4 U16525 ( .A(n15272), .ZN(n19199) );
INV_X4 U16526 ( .A(n14736), .ZN(n19200) );
INV_X4 U16527 ( .A(n15094), .ZN(n19201) );
INV_X4 U16528 ( .A(n16542), .ZN(n19203) );
INV_X4 U16529 ( .A(dii_data_size[1]), .ZN(n19204) );
INV_X4 U16530 ( .A(dii_data_size[0]), .ZN(n19205) );
INV_X4 U16531 ( .A(cii_ctl_vld), .ZN(n19206) );
INV_X4 \GFM/U4594  ( .A(v_in[127]), .ZN(\GFM/n2699 ) );
INV_X4 \GFM/U4593  ( .A(v_in[125]), .ZN(\GFM/n26980 ) );
INV_X4 \GFM/U4592  ( .A(v_in[124]), .ZN(\GFM/n2697 ) );
INV_X4 \GFM/U4591  ( .A(v_in[123]), .ZN(\GFM/n2696 ) );
INV_X4 \GFM/U4590  ( .A(v_in[122]), .ZN(\GFM/n2695 ) );
INV_X4 \GFM/U4589  ( .A(v_out[123]), .ZN(\GFM/n2585 ) );
INV_X4 \GFM/U4588  ( .A(v_out[122]), .ZN(\GFM/n25830 ) );
INV_X4 \GFM/U4587  ( .A(v_out[121]), .ZN(\GFM/n25810 ) );
INV_X4 \GFM/U4586  ( .A(\GFM/N4250 ), .ZN(\GFM/n2579 ) );
INV_X4 \GFM/U4585  ( .A(\GFM/N4248 ), .ZN(\GFM/n25770 ) );
INV_X4 \GFM/U4584  ( .A(v_out[118]), .ZN(\GFM/n2575 ) );
INV_X4 \GFM/U4583  ( .A(\GFM/N4254 ), .ZN(\GFM/n25740 ) );
INV_X4 \GFM/U4582  ( .A(v_out[117]), .ZN(\GFM/n2572 ) );
INV_X4 \GFM/U4581  ( .A(\GFM/N4257 ), .ZN(\GFM/n2571 ) );
INV_X4 \GFM/U4580  ( .A(v_out[116]), .ZN(\GFM/n25690 ) );
INV_X4 \GFM/U4579  ( .A(\GFM/N4242 ), .ZN(\GFM/n2568 ) );
INV_X4 \GFM/U4578  ( .A(v_in[4]), .ZN(\GFM/n25660 ) );
INV_X4 \GFM/U4577  ( .A(v_out[115]), .ZN(\GFM/n2565 ) );
INV_X4 \GFM/U4576  ( .A(\GFM/N4239 ), .ZN(\GFM/n2564 ) );
INV_X4 \GFM/U4575  ( .A(v_in[3]), .ZN(\GFM/n25620 ) );
INV_X4 \GFM/U4574  ( .A(v_out[114]), .ZN(\GFM/n25611 ) );
INV_X4 \GFM/U4573  ( .A(\GFM/N4232 ), .ZN(\GFM/n25600 ) );
INV_X4 \GFM/U4572  ( .A(v_in[2]), .ZN(\GFM/n25580 ) );
INV_X4 \GFM/U4571  ( .A(v_out[113]), .ZN(\GFM/n25570 ) );
INV_X4 \GFM/U4570  ( .A(\GFM/N4235 ), .ZN(\GFM/n2556 ) );
INV_X4 \GFM/U4569  ( .A(v_in[1]), .ZN(\GFM/n2554 ) );
INV_X4 \GFM/U4568  ( .A(b_in[115]), .ZN(\GFM/n25530 ) );
INV_X4 \GFM/U4567  ( .A(\GFM/N4224 ), .ZN(\GFM/n25500 ) );
INV_X4 \GFM/U4566  ( .A(v_out[112]), .ZN(\GFM/n25490 ) );
INV_X4 \GFM/U4565  ( .A(\GFM/N4227 ), .ZN(\GFM/n2548 ) );
INV_X4 \GFM/U4564  ( .A(v_in[0]), .ZN(\GFM/n25460 ) );
BUF_X4 \GFM/U4563  ( .A(v_in[98]), .Z(v_out[82]) );
BUF_X4 \GFM/U4562  ( .A(v_in[99]), .Z(v_out[83]) );
BUF_X4 \GFM/U4561  ( .A(v_in[100]), .Z(v_out[84]) );
BUF_X4 \GFM/U4560  ( .A(v_in[101]), .Z(v_out[85]) );
BUF_X4 \GFM/U4559  ( .A(v_in[102]), .Z(v_out[86]) );
BUF_X4 \GFM/U4558  ( .A(v_in[103]), .Z(v_out[87]) );
BUF_X4 \GFM/U4557  ( .A(v_in[104]), .Z(v_out[88]) );
BUF_X4 \GFM/U4556  ( .A(v_in[105]), .Z(v_out[89]) );
BUF_X4 \GFM/U4555  ( .A(v_in[106]), .Z(v_out[90]) );
BUF_X4 \GFM/U4554  ( .A(v_in[107]), .Z(v_out[91]) );
BUF_X4 \GFM/U4553  ( .A(v_in[108]), .Z(v_out[92]) );
BUF_X4 \GFM/U4552  ( .A(v_in[109]), .Z(v_out[93]) );
BUF_X4 \GFM/U4551  ( .A(v_in[110]), .Z(v_out[94]) );
BUF_X4 \GFM/U4550  ( .A(v_in[111]), .Z(v_out[95]) );
BUF_X4 \GFM/U4549  ( .A(v_in[112]), .Z(v_out[96]) );
BUF_X4 \GFM/U4548  ( .A(v_in[113]), .Z(v_out[97]) );
BUF_X4 \GFM/U4547  ( .A(v_in[114]), .Z(v_out[98]) );
BUF_X4 \GFM/U4546  ( .A(v_in[115]), .Z(v_out[99]) );
BUF_X4 \GFM/U4545  ( .A(v_in[116]), .Z(v_out[100]) );
BUF_X4 \GFM/U4544  ( .A(v_in[117]), .Z(v_out[101]) );
BUF_X4 \GFM/U4543  ( .A(v_in[118]), .Z(v_out[102]) );
BUF_X4 \GFM/U4542  ( .A(v_in[119]), .Z(v_out[103]) );
BUF_X4 \GFM/U4541  ( .A(v_in[120]), .Z(v_out[104]) );
INV_X4 \GFM/U4540  ( .A(v_in[36]), .ZN(\GFM/n2610 ) );
INV_X4 \GFM/U4539  ( .A(v_in[34]), .ZN(\GFM/n26080 ) );
INV_X4 \GFM/U4538  ( .A(v_in[33]), .ZN(\GFM/n26070 ) );
INV_X4 \GFM/U4537  ( .A(v_in[32]), .ZN(\GFM/n2606 ) );
INV_X4 \GFM/U4536  ( .A(v_in[46]), .ZN(\GFM/n26200 ) );
INV_X4 \GFM/U4535  ( .A(v_in[45]), .ZN(\GFM/n26190 ) );
INV_X4 \GFM/U4534  ( .A(v_in[43]), .ZN(\GFM/n2617 ) );
INV_X4 \GFM/U4533  ( .A(v_in[44]), .ZN(\GFM/n2618 ) );
INV_X4 \GFM/U4532  ( .A(v_in[38]), .ZN(\GFM/n26120 ) );
INV_X4 \GFM/U4531  ( .A(v_in[39]), .ZN(\GFM/n2613 ) );
INV_X4 \GFM/U4530  ( .A(v_in[42]), .ZN(\GFM/n2616 ) );
INV_X4 \GFM/U4529  ( .A(v_in[40]), .ZN(\GFM/n26140 ) );
INV_X4 \GFM/U4528  ( .A(v_in[41]), .ZN(\GFM/n26150 ) );
INV_X4 \GFM/U4527  ( .A(v_in[37]), .ZN(\GFM/n26110 ) );
INV_X4 \GFM/U4526  ( .A(v_in[16]), .ZN(\GFM/n25901 ) );
INV_X4 \GFM/U4525  ( .A(v_in[17]), .ZN(\GFM/n25910 ) );
INV_X4 \GFM/U4524  ( .A(v_in[18]), .ZN(\GFM/n2592 ) );
INV_X4 \GFM/U4523  ( .A(v_in[19]), .ZN(\GFM/n25930 ) );
INV_X4 \GFM/U4522  ( .A(v_in[20]), .ZN(\GFM/n25940 ) );
INV_X4 \GFM/U4521  ( .A(v_in[21]), .ZN(\GFM/n2595 ) );
INV_X4 \GFM/U4520  ( .A(v_in[22]), .ZN(\GFM/n2596 ) );
INV_X4 \GFM/U4519  ( .A(v_in[23]), .ZN(\GFM/n25970 ) );
INV_X4 \GFM/U4518  ( .A(v_in[24]), .ZN(\GFM/n25980 ) );
INV_X4 \GFM/U4517  ( .A(v_in[25]), .ZN(\GFM/n2599 ) );
INV_X4 \GFM/U4516  ( .A(v_in[26]), .ZN(\GFM/n26000 ) );
INV_X4 \GFM/U4515  ( .A(v_in[27]), .ZN(\GFM/n26010 ) );
INV_X4 \GFM/U4514  ( .A(v_in[28]), .ZN(\GFM/n2602 ) );
INV_X4 \GFM/U4513  ( .A(v_in[29]), .ZN(\GFM/n2603 ) );
INV_X4 \GFM/U4512  ( .A(v_in[30]), .ZN(\GFM/n2604 ) );
INV_X4 \GFM/U4511  ( .A(v_in[31]), .ZN(\GFM/n26050 ) );
INV_X4 \GFM/U4510  ( .A(v_in[35]), .ZN(\GFM/n2609 ) );
INV_X4 \GFM/U4509  ( .A(v_in[47]), .ZN(\GFM/n2621 ) );
INV_X4 \GFM/U4508  ( .A(v_in[48]), .ZN(\GFM/n26220 ) );
INV_X4 \GFM/U4507  ( .A(v_in[49]), .ZN(\GFM/n2623 ) );
INV_X4 \GFM/U4506  ( .A(v_in[50]), .ZN(\GFM/n26240 ) );
INV_X4 \GFM/U4505  ( .A(v_in[51]), .ZN(\GFM/n26250 ) );
INV_X4 \GFM/U4504  ( .A(v_in[52]), .ZN(\GFM/n2626 ) );
INV_X4 \GFM/U4503  ( .A(v_in[53]), .ZN(\GFM/n2627 ) );
INV_X4 \GFM/U4502  ( .A(v_in[54]), .ZN(\GFM/n26280 ) );
INV_X4 \GFM/U4501  ( .A(v_in[55]), .ZN(\GFM/n26290 ) );
INV_X4 \GFM/U4500  ( .A(v_in[56]), .ZN(\GFM/n26301 ) );
INV_X4 \GFM/U4499  ( .A(v_in[57]), .ZN(\GFM/n26310 ) );
INV_X4 \GFM/U4498  ( .A(v_in[58]), .ZN(\GFM/n26320 ) );
INV_X4 \GFM/U4497  ( .A(v_in[59]), .ZN(\GFM/n2633 ) );
INV_X4 \GFM/U4496  ( .A(v_in[60]), .ZN(\GFM/n2634 ) );
INV_X4 \GFM/U4495  ( .A(v_in[61]), .ZN(\GFM/n2635 ) );
INV_X4 \GFM/U4494  ( .A(v_in[62]), .ZN(\GFM/n26360 ) );
INV_X4 \GFM/U4493  ( .A(v_in[63]), .ZN(\GFM/n2637 ) );
INV_X4 \GFM/U4492  ( .A(v_in[64]), .ZN(\GFM/n26380 ) );
INV_X4 \GFM/U4491  ( .A(v_in[68]), .ZN(\GFM/n26420 ) );
INV_X4 \GFM/U4490  ( .A(v_in[69]), .ZN(\GFM/n26430 ) );
INV_X4 \GFM/U4489  ( .A(v_in[70]), .ZN(\GFM/n2644 ) );
INV_X4 \GFM/U4488  ( .A(v_in[71]), .ZN(\GFM/n26450 ) );
INV_X4 \GFM/U4487  ( .A(v_in[72]), .ZN(\GFM/n26460 ) );
INV_X4 \GFM/U4486  ( .A(v_in[73]), .ZN(\GFM/n2647 ) );
INV_X4 \GFM/U4485  ( .A(v_in[74]), .ZN(\GFM/n2648 ) );
INV_X4 \GFM/U4484  ( .A(v_in[75]), .ZN(\GFM/n2649 ) );
INV_X4 \GFM/U4483  ( .A(v_in[76]), .ZN(\GFM/n26500 ) );
INV_X4 \GFM/U4482  ( .A(v_in[77]), .ZN(\GFM/n26510 ) );
INV_X4 \GFM/U4481  ( .A(v_in[78]), .ZN(\GFM/n2652 ) );
INV_X4 \GFM/U4480  ( .A(v_in[79]), .ZN(\GFM/n26530 ) );
INV_X4 \GFM/U4479  ( .A(v_in[80]), .ZN(\GFM/n2654 ) );
INV_X4 \GFM/U4478  ( .A(v_in[81]), .ZN(\GFM/n26550 ) );
INV_X4 \GFM/U4477  ( .A(v_in[82]), .ZN(\GFM/n26560 ) );
INV_X4 \GFM/U4476  ( .A(v_in[83]), .ZN(\GFM/n2657 ) );
INV_X4 \GFM/U4475  ( .A(v_in[84]), .ZN(\GFM/n2658 ) );
INV_X4 \GFM/U4474  ( .A(v_in[85]), .ZN(\GFM/n26590 ) );
INV_X4 \GFM/U4473  ( .A(v_in[86]), .ZN(\GFM/n26600 ) );
INV_X4 \GFM/U4472  ( .A(v_in[87]), .ZN(\GFM/n26611 ) );
INV_X4 \GFM/U4471  ( .A(v_in[88]), .ZN(\GFM/n26620 ) );
INV_X4 \GFM/U4470  ( .A(v_in[89]), .ZN(\GFM/n26630 ) );
INV_X4 \GFM/U4469  ( .A(v_in[90]), .ZN(\GFM/n2664 ) );
INV_X4 \GFM/U4468  ( .A(v_in[91]), .ZN(\GFM/n2665 ) );
INV_X4 \GFM/U4467  ( .A(v_in[92]), .ZN(\GFM/n2666 ) );
INV_X4 \GFM/U4466  ( .A(v_in[93]), .ZN(\GFM/n26670 ) );
INV_X4 \GFM/U4465  ( .A(v_in[94]), .ZN(\GFM/n2668 ) );
INV_X4 \GFM/U4464  ( .A(v_in[95]), .ZN(\GFM/n26690 ) );
INV_X4 \GFM/U4463  ( .A(v_in[96]), .ZN(\GFM/n26700 ) );
INV_X4 \GFM/U4462  ( .A(v_in[97]), .ZN(\GFM/n2671 ) );
INV_X4 \GFM/U4461  ( .A(v_in[98]), .ZN(\GFM/n2672 ) );
INV_X4 \GFM/U4460  ( .A(v_in[99]), .ZN(\GFM/n26730 ) );
INV_X4 \GFM/U4459  ( .A(v_in[100]), .ZN(\GFM/n26740 ) );
INV_X4 \GFM/U4458  ( .A(v_in[101]), .ZN(\GFM/n2675 ) );
INV_X4 \GFM/U4457  ( .A(v_in[102]), .ZN(\GFM/n26760 ) );
INV_X4 \GFM/U4456  ( .A(v_in[103]), .ZN(\GFM/n26770 ) );
INV_X4 \GFM/U4455  ( .A(v_in[104]), .ZN(\GFM/n2678 ) );
INV_X4 \GFM/U4454  ( .A(v_in[105]), .ZN(\GFM/n2679 ) );
INV_X4 \GFM/U4453  ( .A(v_in[106]), .ZN(\GFM/n26801 ) );
INV_X4 \GFM/U4452  ( .A(v_in[107]), .ZN(\GFM/n26810 ) );
INV_X4 \GFM/U4451  ( .A(v_in[108]), .ZN(\GFM/n26820 ) );
INV_X4 \GFM/U4450  ( .A(v_in[109]), .ZN(\GFM/n2683 ) );
INV_X4 \GFM/U4449  ( .A(v_in[110]), .ZN(\GFM/n26840 ) );
INV_X4 \GFM/U4448  ( .A(v_in[111]), .ZN(\GFM/n2685 ) );
INV_X4 \GFM/U4447  ( .A(v_in[112]), .ZN(\GFM/n26860 ) );
INV_X4 \GFM/U4446  ( .A(v_in[113]), .ZN(\GFM/n26870 ) );
INV_X4 \GFM/U4445  ( .A(v_in[114]), .ZN(\GFM/n2688 ) );
INV_X4 \GFM/U4444  ( .A(v_in[115]), .ZN(\GFM/n2689 ) );
INV_X4 \GFM/U4443  ( .A(v_in[116]), .ZN(\GFM/n26900 ) );
INV_X4 \GFM/U4442  ( .A(v_in[117]), .ZN(\GFM/n26910 ) );
INV_X4 \GFM/U4441  ( .A(v_in[118]), .ZN(\GFM/n26921 ) );
INV_X4 \GFM/U4440  ( .A(v_in[119]), .ZN(\GFM/n26930 ) );
INV_X4 \GFM/U4439  ( .A(v_in[120]), .ZN(\GFM/n26940 ) );
BUF_X4 \GFM/U4438  ( .A(v_in[16]), .Z(v_out[0]) );
BUF_X4 \GFM/U4437  ( .A(v_in[17]), .Z(v_out[1]) );
BUF_X4 \GFM/U4436  ( .A(v_in[18]), .Z(v_out[2]) );
BUF_X4 \GFM/U4435  ( .A(v_in[19]), .Z(v_out[3]) );
BUF_X4 \GFM/U4434  ( .A(v_in[20]), .Z(v_out[4]) );
BUF_X4 \GFM/U4433  ( .A(v_in[21]), .Z(v_out[5]) );
BUF_X4 \GFM/U4432  ( .A(v_in[22]), .Z(v_out[6]) );
BUF_X4 \GFM/U4431  ( .A(v_in[23]), .Z(v_out[7]) );
BUF_X4 \GFM/U4430  ( .A(v_in[24]), .Z(v_out[8]) );
BUF_X4 \GFM/U4429  ( .A(v_in[25]), .Z(v_out[9]) );
BUF_X4 \GFM/U4428  ( .A(v_in[26]), .Z(v_out[10]) );
BUF_X4 \GFM/U4427  ( .A(v_in[27]), .Z(v_out[11]) );
BUF_X4 \GFM/U4426  ( .A(v_in[28]), .Z(v_out[12]) );
BUF_X4 \GFM/U4425  ( .A(v_in[29]), .Z(v_out[13]) );
BUF_X4 \GFM/U4424  ( .A(v_in[30]), .Z(v_out[14]) );
BUF_X4 \GFM/U4423  ( .A(v_in[31]), .Z(v_out[15]) );
BUF_X4 \GFM/U4422  ( .A(v_in[32]), .Z(v_out[16]) );
BUF_X4 \GFM/U4421  ( .A(v_in[33]), .Z(v_out[17]) );
BUF_X4 \GFM/U4420  ( .A(v_in[34]), .Z(v_out[18]) );
BUF_X4 \GFM/U4419  ( .A(v_in[35]), .Z(v_out[19]) );
BUF_X4 \GFM/U4418  ( .A(v_in[36]), .Z(v_out[20]) );
BUF_X4 \GFM/U4417  ( .A(v_in[37]), .Z(v_out[21]) );
BUF_X4 \GFM/U4416  ( .A(v_in[38]), .Z(v_out[22]) );
BUF_X4 \GFM/U4415  ( .A(v_in[39]), .Z(v_out[23]) );
BUF_X4 \GFM/U4414  ( .A(v_in[40]), .Z(v_out[24]) );
BUF_X4 \GFM/U4413  ( .A(v_in[41]), .Z(v_out[25]) );
BUF_X4 \GFM/U4412  ( .A(v_in[42]), .Z(v_out[26]) );
BUF_X4 \GFM/U4411  ( .A(v_in[43]), .Z(v_out[27]) );
BUF_X4 \GFM/U4410  ( .A(v_in[44]), .Z(v_out[28]) );
BUF_X4 \GFM/U4409  ( .A(v_in[45]), .Z(v_out[29]) );
BUF_X4 \GFM/U4408  ( .A(v_in[46]), .Z(v_out[30]) );
BUF_X4 \GFM/U4407  ( .A(v_in[47]), .Z(v_out[31]) );
BUF_X4 \GFM/U4406  ( .A(v_in[48]), .Z(v_out[32]) );
BUF_X4 \GFM/U4405  ( .A(v_in[49]), .Z(v_out[33]) );
BUF_X4 \GFM/U4404  ( .A(v_in[50]), .Z(v_out[34]) );
BUF_X4 \GFM/U4403  ( .A(v_in[51]), .Z(v_out[35]) );
BUF_X4 \GFM/U4402  ( .A(v_in[52]), .Z(v_out[36]) );
BUF_X4 \GFM/U4401  ( .A(v_in[53]), .Z(v_out[37]) );
BUF_X4 \GFM/U4400  ( .A(v_in[54]), .Z(v_out[38]) );
BUF_X4 \GFM/U4399  ( .A(v_in[55]), .Z(v_out[39]) );
BUF_X4 \GFM/U4398  ( .A(v_in[56]), .Z(v_out[40]) );
BUF_X4 \GFM/U4397  ( .A(v_in[57]), .Z(v_out[41]) );
BUF_X4 \GFM/U4396  ( .A(v_in[58]), .Z(v_out[42]) );
BUF_X4 \GFM/U4395  ( .A(v_in[59]), .Z(v_out[43]) );
BUF_X4 \GFM/U4394  ( .A(v_in[60]), .Z(v_out[44]) );
BUF_X4 \GFM/U4393  ( .A(v_in[61]), .Z(v_out[45]) );
BUF_X4 \GFM/U4392  ( .A(v_in[62]), .Z(v_out[46]) );
BUF_X4 \GFM/U4391  ( .A(v_in[63]), .Z(v_out[47]) );
BUF_X4 \GFM/U4390  ( .A(v_in[64]), .Z(v_out[48]) );
BUF_X4 \GFM/U4389  ( .A(v_in[65]), .Z(v_out[49]) );
BUF_X4 \GFM/U4388  ( .A(v_in[66]), .Z(v_out[50]) );
BUF_X4 \GFM/U4387  ( .A(v_in[67]), .Z(v_out[51]) );
BUF_X4 \GFM/U4386  ( .A(v_in[68]), .Z(v_out[52]) );
BUF_X4 \GFM/U4385  ( .A(v_in[69]), .Z(v_out[53]) );
BUF_X4 \GFM/U4384  ( .A(v_in[70]), .Z(v_out[54]) );
BUF_X4 \GFM/U4383  ( .A(v_in[71]), .Z(v_out[55]) );
BUF_X4 \GFM/U4382  ( .A(v_in[72]), .Z(v_out[56]) );
BUF_X4 \GFM/U4381  ( .A(v_in[73]), .Z(v_out[57]) );
BUF_X4 \GFM/U4380  ( .A(v_in[74]), .Z(v_out[58]) );
BUF_X4 \GFM/U4379  ( .A(v_in[75]), .Z(v_out[59]) );
BUF_X4 \GFM/U4378  ( .A(v_in[76]), .Z(v_out[60]) );
BUF_X4 \GFM/U4377  ( .A(v_in[77]), .Z(v_out[61]) );
BUF_X4 \GFM/U4376  ( .A(v_in[78]), .Z(v_out[62]) );
BUF_X4 \GFM/U4375  ( .A(v_in[79]), .Z(v_out[63]) );
BUF_X4 \GFM/U4374  ( .A(v_in[80]), .Z(v_out[64]) );
BUF_X4 \GFM/U4373  ( .A(v_in[81]), .Z(v_out[65]) );
BUF_X4 \GFM/U4372  ( .A(v_in[82]), .Z(v_out[66]) );
BUF_X4 \GFM/U4371  ( .A(v_in[83]), .Z(v_out[67]) );
BUF_X4 \GFM/U4370  ( .A(v_in[84]), .Z(v_out[68]) );
BUF_X4 \GFM/U4369  ( .A(v_in[85]), .Z(v_out[69]) );
BUF_X4 \GFM/U4368  ( .A(v_in[86]), .Z(v_out[70]) );
BUF_X4 \GFM/U4367  ( .A(v_in[87]), .Z(v_out[71]) );
BUF_X4 \GFM/U4366  ( .A(v_in[88]), .Z(v_out[72]) );
BUF_X4 \GFM/U4365  ( .A(v_in[89]), .Z(v_out[73]) );
BUF_X4 \GFM/U4364  ( .A(v_in[90]), .Z(v_out[74]) );
BUF_X4 \GFM/U4363  ( .A(v_in[91]), .Z(v_out[75]) );
BUF_X4 \GFM/U4362  ( .A(v_in[92]), .Z(v_out[76]) );
BUF_X4 \GFM/U4361  ( .A(v_in[93]), .Z(v_out[77]) );
BUF_X4 \GFM/U4360  ( .A(v_in[94]), .Z(v_out[78]) );
BUF_X4 \GFM/U4359  ( .A(v_in[95]), .Z(v_out[79]) );
BUF_X4 \GFM/U4358  ( .A(v_in[96]), .Z(v_out[80]) );
BUF_X4 \GFM/U4357  ( .A(v_in[97]), .Z(v_out[81]) );
NOR2_X2 \GFM/U4356  ( .A1(\GFM/n2409 ), .A2(\GFM/n2572 ), .ZN(\GFM/N3985 ));
NOR2_X2 \GFM/U4355  ( .A1(\GFM/n2697 ), .A2(\GFM/n2516 ), .ZN(\GFM/N4049 ));
NOR2_X2 \GFM/U4354  ( .A1(\GFM/n2695 ), .A2(\GFM/n25360 ), .ZN(\GFM/N4047 ));
NAND3_X2 \GFM/U4353  ( .A1(b_in[119]), .A2(\GFM/n25760 ), .A3(v_in[6]), .ZN(\GFM/n17911 ) );
BUF_X4 \GFM/U4352  ( .A(v_in[15]), .Z(v_out[127]) );
NAND3_X2 \GFM/U4351  ( .A1(b_in[115]), .A2(\GFM/n25840 ), .A3(v_in[10]),.ZN(\GFM/n17511 ) );
NAND3_X2 \GFM/U4350  ( .A1(b_in[116]), .A2(\GFM/n25821 ), .A3(v_in[9]), .ZN(\GFM/n18310 ) );
NAND3_X2 \GFM/U4349  ( .A1(b_in[117]), .A2(\GFM/n25800 ), .A3(v_in[8]), .ZN(\GFM/n2121 ) );
NAND3_X2 \GFM/U4348  ( .A1(b_in[118]), .A2(\GFM/n2578 ), .A3(v_in[7]), .ZN(\GFM/n181 ) );
NAND3_X2 \GFM/U4347  ( .A1(b_in[113]), .A2(\GFM/n2587 ), .A3(v_in[12]), .ZN(\GFM/n17310 ) );
NAND3_X2 \GFM/U4346  ( .A1(b_in[120]), .A2(\GFM/n2573 ), .A3(v_in[5]), .ZN(\GFM/n21230 ) );
NAND3_X2 \GFM/U4345  ( .A1(b_in[114]), .A2(\GFM/n2586 ), .A3(v_in[11]), .ZN(\GFM/n177 ) );
NAND3_X2 \GFM/U4344  ( .A1(b_in[126]), .A2(\GFM/n25460 ), .A3(v_in[127]),.ZN(\GFM/n21350 ) );
NAND3_X2 \GFM/U4343  ( .A1(v_in[3]), .A2(\GFM/n25660 ), .A3(b_in[122]), .ZN(\GFM/n21290 ) );
NAND3_X2 \GFM/U4342  ( .A1(b_in[112]), .A2(\GFM/n25880 ), .A3(v_in[13]),.ZN(\GFM/n17110 ) );
NAND3_X2 \GFM/U4341  ( .A1(v_in[4]), .A2(\GFM/n25700 ), .A3(b_in[121]), .ZN(\GFM/n2125 ) );
NAND3_X2 \GFM/U4340  ( .A1(v_in[2]), .A2(\GFM/n25620 ), .A3(b_in[123]), .ZN(\GFM/n2127 ) );
NAND3_X2 \GFM/U4339  ( .A1(v_in[1]), .A2(\GFM/n25580 ), .A3(b_in[124]), .ZN(\GFM/n2131 ) );
NAND3_X2 \GFM/U4338  ( .A1(v_in[0]), .A2(\GFM/n2554 ), .A3(b_in[125]), .ZN(\GFM/n21330 ) );
INV_X4 \GFM/U4337  ( .A(v_in[5]), .ZN(\GFM/n25700 ) );
INV_X4 \GFM/U4336  ( .A(v_in[6]), .ZN(\GFM/n2573 ) );
INV_X4 \GFM/U4335  ( .A(v_in[7]), .ZN(\GFM/n25760 ) );
INV_X4 \GFM/U4334  ( .A(v_in[8]), .ZN(\GFM/n2578 ) );
INV_X4 \GFM/U4333  ( .A(v_in[9]), .ZN(\GFM/n25800 ) );
INV_X4 \GFM/U4332  ( .A(v_in[65]), .ZN(\GFM/n26390 ) );
INV_X4 \GFM/U4331  ( .A(v_in[66]), .ZN(\GFM/n26401 ) );
INV_X4 \GFM/U4330  ( .A(v_in[67]), .ZN(\GFM/n2641 ) );
INV_X4 \GFM/U4329  ( .A(v_in[10]), .ZN(\GFM/n25821 ) );
INV_X4 \GFM/U2238  ( .A(v_in[15]), .ZN(\GFM/n25890 ) );
INV_X4 \GFM/U2237  ( .A(v_in[11]), .ZN(\GFM/n25840 ) );
NOR2_X2 \GFM/U2236  ( .A1(\GFM/n25890 ), .A2(\GFM/n2387 ), .ZN(\GFM/N28 ) );
NOR2_X2 \GFM/U2235  ( .A1(\GFM/n25890 ), .A2(\GFM/n23970 ), .ZN(\GFM/N58 ));
NOR2_X2 \GFM/U2234  ( .A1(\GFM/n23980 ), .A2(\GFM/n25901 ), .ZN(\GFM/N89 ));
NOR2_X2 \GFM/U2233  ( .A1(\GFM/n2406 ), .A2(\GFM/n25910 ), .ZN(\GFM/N120 ));
NOR2_X2 \GFM/U2232  ( .A1(\GFM/n24050 ), .A2(\GFM/n2592 ), .ZN(\GFM/N151 ));
NOR2_X2 \GFM/U2231  ( .A1(\GFM/n2404 ), .A2(\GFM/n25930 ), .ZN(\GFM/N182 ));
NOR2_X2 \GFM/U2230  ( .A1(\GFM/n24030 ), .A2(\GFM/n25940 ), .ZN(\GFM/N213 ));
NOR2_X2 \GFM/U2229  ( .A1(\GFM/n24030 ), .A2(\GFM/n2595 ), .ZN(\GFM/N244 ));
NOR2_X2 \GFM/U2228  ( .A1(\GFM/n24020 ), .A2(\GFM/n2596 ), .ZN(\GFM/N275 ));
NOR2_X2 \GFM/U2227  ( .A1(\GFM/n2401 ), .A2(\GFM/n25970 ), .ZN(\GFM/N306 ));
NOR2_X2 \GFM/U2226  ( .A1(\GFM/n2400 ), .A2(\GFM/n25980 ), .ZN(\GFM/N337 ));
NOR2_X2 \GFM/U2225  ( .A1(\GFM/n2400 ), .A2(\GFM/n2599 ), .ZN(\GFM/N368 ) );
NOR2_X2 \GFM/U2224  ( .A1(\GFM/n2399 ), .A2(\GFM/n26000 ), .ZN(\GFM/N399 ));
NOR2_X2 \GFM/U2223  ( .A1(\GFM/n2399 ), .A2(\GFM/n26010 ), .ZN(\GFM/N430 ));
NOR2_X2 \GFM/U2222  ( .A1(\GFM/n23980 ), .A2(\GFM/n2602 ), .ZN(\GFM/N461 ));
NOR2_X2 \GFM/U2221  ( .A1(\GFM/n2399 ), .A2(\GFM/n2603 ), .ZN(\GFM/N492 ) );
NOR2_X2 \GFM/U2220  ( .A1(\GFM/n23980 ), .A2(\GFM/n2604 ), .ZN(\GFM/N523 ));
NOR2_X2 \GFM/U2219  ( .A1(\GFM/n2606 ), .A2(\GFM/n2387 ), .ZN(\GFM/N555 ) );
NOR2_X2 \GFM/U2218  ( .A1(\GFM/n2606 ), .A2(\GFM/n23970 ), .ZN(\GFM/N585 ));
NOR2_X2 \GFM/U2217  ( .A1(\GFM/n26070 ), .A2(\GFM/n23970 ), .ZN(\GFM/N616 ));
NOR2_X2 \GFM/U2216  ( .A1(\GFM/n26080 ), .A2(\GFM/n23970 ), .ZN(\GFM/N647 ));
NOR2_X2 \GFM/U2215  ( .A1(\GFM/n2610 ), .A2(\GFM/n2387 ), .ZN(\GFM/N679 ) );
NOR2_X2 \GFM/U2214  ( .A1(\GFM/n2610 ), .A2(\GFM/n23970 ), .ZN(\GFM/N709 ));
NOR2_X2 \GFM/U2213  ( .A1(\GFM/n23980 ), .A2(\GFM/n26110 ), .ZN(\GFM/N740 ));
NOR2_X2 \GFM/U2212  ( .A1(\GFM/n23980 ), .A2(\GFM/n26120 ), .ZN(\GFM/N771 ));
NOR2_X2 \GFM/U2211  ( .A1(\GFM/n23980 ), .A2(\GFM/n2613 ), .ZN(\GFM/N802 ));
NOR2_X2 \GFM/U2210  ( .A1(\GFM/n23980 ), .A2(\GFM/n26140 ), .ZN(\GFM/N833 ));
NOR2_X2 \GFM/U2209  ( .A1(\GFM/n23980 ), .A2(\GFM/n26150 ), .ZN(\GFM/N864 ));
NOR2_X2 \GFM/U2208  ( .A1(\GFM/n23980 ), .A2(\GFM/n2616 ), .ZN(\GFM/N895 ));
NOR2_X2 \GFM/U2207  ( .A1(\GFM/n2387 ), .A2(\GFM/n2618 ), .ZN(\GFM/N927 ) );
NOR2_X2 \GFM/U2206  ( .A1(\GFM/n23980 ), .A2(\GFM/n2618 ), .ZN(\GFM/N957 ));
NOR2_X2 \GFM/U2205  ( .A1(\GFM/n24020 ), .A2(\GFM/n26190 ), .ZN(\GFM/N988 ));
NOR2_X2 \GFM/U2204  ( .A1(\GFM/n26200 ), .A2(\GFM/n23970 ), .ZN(\GFM/N1019 ));
NOR2_X2 \GFM/U2203  ( .A1(\GFM/n23980 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1050 ));
NOR2_X2 \GFM/U2202  ( .A1(\GFM/n2406 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1081 ));
NOR2_X2 \GFM/U2201  ( .A1(\GFM/n2406 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1112 ));
NOR2_X2 \GFM/U2200  ( .A1(\GFM/n2406 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1143 ));
NOR2_X2 \GFM/U2199  ( .A1(\GFM/n2406 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1174 ));
NOR2_X2 \GFM/U2198  ( .A1(\GFM/n2406 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1205 ));
NOR2_X2 \GFM/U2197  ( .A1(\GFM/n2406 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1236 ));
NOR2_X2 \GFM/U2196  ( .A1(\GFM/n2406 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1267 ));
NOR2_X2 \GFM/U2195  ( .A1(\GFM/n2406 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1298 ));
NOR2_X2 \GFM/U2194  ( .A1(\GFM/n2406 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1329 ));
NOR2_X2 \GFM/U2193  ( .A1(\GFM/n2406 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1360 ));
NOR2_X2 \GFM/U2192  ( .A1(\GFM/n24050 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1391 ));
NOR2_X2 \GFM/U2191  ( .A1(\GFM/n24050 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1422 ));
NOR2_X2 \GFM/U2190  ( .A1(\GFM/n24050 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1453 ));
NOR2_X2 \GFM/U2189  ( .A1(\GFM/n24050 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1484 ));
NOR2_X2 \GFM/U2188  ( .A1(\GFM/n24050 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1515 ));
NOR2_X2 \GFM/U2187  ( .A1(\GFM/n24050 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1546 ));
NOR2_X2 \GFM/U2186  ( .A1(\GFM/n24050 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1577 ));
NOR2_X2 \GFM/U2185  ( .A1(\GFM/n24050 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1608 ));
NOR2_X2 \GFM/U2184  ( .A1(\GFM/n24050 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1639 ));
NOR2_X2 \GFM/U2183  ( .A1(\GFM/n24050 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1670 ));
NOR2_X2 \GFM/U2182  ( .A1(\GFM/n24050 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1701 ));
NOR2_X2 \GFM/U2181  ( .A1(\GFM/n24050 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1732 ));
NOR2_X2 \GFM/U2180  ( .A1(\GFM/n2404 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1763 ));
NOR2_X2 \GFM/U2179  ( .A1(\GFM/n2404 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1794 ));
NOR2_X2 \GFM/U2178  ( .A1(\GFM/n2404 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1825 ));
NOR2_X2 \GFM/U2177  ( .A1(\GFM/n2404 ), .A2(\GFM/n2647 ), .ZN(\GFM/N1856 ));
NOR2_X2 \GFM/U2176  ( .A1(\GFM/n2404 ), .A2(\GFM/n2648 ), .ZN(\GFM/N1887 ));
NOR2_X2 \GFM/U2175  ( .A1(\GFM/n2404 ), .A2(\GFM/n2649 ), .ZN(\GFM/N1918 ));
NOR2_X2 \GFM/U2174  ( .A1(\GFM/n2404 ), .A2(\GFM/n26500 ), .ZN(\GFM/N1949 ));
NOR2_X2 \GFM/U2173  ( .A1(\GFM/n2404 ), .A2(\GFM/n26510 ), .ZN(\GFM/N1980 ));
NOR2_X2 \GFM/U2172  ( .A1(\GFM/n2404 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2011 ));
NOR2_X2 \GFM/U2171  ( .A1(\GFM/n2404 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2042 ));
NOR2_X2 \GFM/U2170  ( .A1(\GFM/n2404 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2073 ));
NOR2_X2 \GFM/U2169  ( .A1(\GFM/n2404 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2104 ));
NOR2_X2 \GFM/U2168  ( .A1(\GFM/n24030 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2135 ));
NOR2_X2 \GFM/U2167  ( .A1(\GFM/n24030 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2166 ));
NOR2_X2 \GFM/U2166  ( .A1(\GFM/n24030 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2197 ));
NOR2_X2 \GFM/U2165  ( .A1(\GFM/n24030 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2228 ));
NOR2_X2 \GFM/U2164  ( .A1(\GFM/n24030 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2259 ));
NOR2_X2 \GFM/U2163  ( .A1(\GFM/n24030 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2290 ));
NOR2_X2 \GFM/U2162  ( .A1(\GFM/n24030 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2321 ));
NOR2_X2 \GFM/U2161  ( .A1(\GFM/n24030 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2352 ));
NOR2_X2 \GFM/U2160  ( .A1(\GFM/n24030 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2383 ));
NOR2_X2 \GFM/U2159  ( .A1(\GFM/n24030 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2414 ));
NOR2_X2 \GFM/U2158  ( .A1(\GFM/n24030 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2445 ));
NOR2_X2 \GFM/U2157  ( .A1(\GFM/n24020 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2476 ));
NOR2_X2 \GFM/U2156  ( .A1(\GFM/n24020 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2507 ));
NOR2_X2 \GFM/U2155  ( .A1(\GFM/n24020 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2538 ));
NOR2_X2 \GFM/U2154  ( .A1(\GFM/n24020 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2569 ));
NOR2_X2 \GFM/U2153  ( .A1(\GFM/n24020 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2600 ));
NOR2_X2 \GFM/U2152  ( .A1(\GFM/n24020 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2631 ));
NOR2_X2 \GFM/U2151  ( .A1(\GFM/n24020 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2662 ));
NOR2_X2 \GFM/U2150  ( .A1(\GFM/n24020 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2693 ));
NOR2_X2 \GFM/U2149  ( .A1(\GFM/n24020 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2724 ));
NOR2_X2 \GFM/U2148  ( .A1(\GFM/n24020 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2755 ));
NOR2_X2 \GFM/U2147  ( .A1(\GFM/n24020 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2786 ));
NOR2_X2 \GFM/U2146  ( .A1(\GFM/n2401 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2817 ));
NOR2_X2 \GFM/U2145  ( .A1(\GFM/n2401 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2848 ));
NOR2_X2 \GFM/U2144  ( .A1(\GFM/n2401 ), .A2(\GFM/n26801 ), .ZN(\GFM/N2879 ));
NOR2_X2 \GFM/U2143  ( .A1(\GFM/n2401 ), .A2(\GFM/n26810 ), .ZN(\GFM/N2910 ));
NOR2_X2 \GFM/U2142  ( .A1(\GFM/n2401 ), .A2(\GFM/n26820 ), .ZN(\GFM/N2941 ));
NOR2_X2 \GFM/U2141  ( .A1(\GFM/n2401 ), .A2(\GFM/n2683 ), .ZN(\GFM/N2972 ));
NOR2_X2 \GFM/U2140  ( .A1(\GFM/n2401 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3003 ));
NOR2_X2 \GFM/U2139  ( .A1(\GFM/n2401 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3034 ));
NOR2_X2 \GFM/U2138  ( .A1(\GFM/n2401 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3065 ));
NOR2_X2 \GFM/U2137  ( .A1(\GFM/n2401 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3096 ));
NOR2_X2 \GFM/U2136  ( .A1(\GFM/n2401 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3127 ));
NOR2_X2 \GFM/U2135  ( .A1(\GFM/n2401 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3158 ));
NOR2_X2 \GFM/U2134  ( .A1(\GFM/n2400 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3189 ));
NOR2_X2 \GFM/U2133  ( .A1(\GFM/n2400 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3220 ));
NOR2_X2 \GFM/U2132  ( .A1(\GFM/n2400 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3251 ));
NOR2_X2 \GFM/U2131  ( .A1(\GFM/n2400 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3282 ));
NOR2_X2 \GFM/U2130  ( .A1(\GFM/n25180 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3747 ));
NOR2_X2 \GFM/U2129  ( .A1(\GFM/n25380 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3745 ));
NOR2_X2 \GFM/U2128  ( .A1(\GFM/n2547 ), .A2(\GFM/n25270 ), .ZN(\GFM/N3931 ));
NOR2_X2 \GFM/U2127  ( .A1(\GFM/n25380 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3928 ));
INV_X4 \GFM/U2126  ( .A(v_in[12]), .ZN(\GFM/n2586 ) );
INV_X4 \GFM/U2125  ( .A(v_in[14]), .ZN(\GFM/n25880 ) );
INV_X4 \GFM/U2124  ( .A(v_in[13]), .ZN(\GFM/n2587 ) );
INV_X4 \GFM/U2123  ( .A(b_in[123]), .ZN(\GFM/n24960 ) );
INV_X4 \GFM/U2122  ( .A(b_in[112]), .ZN(\GFM/n2387 ) );
INV_X4 \GFM/U2121  ( .A(b_in[114]), .ZN(\GFM/n24070 ) );
INV_X4 \GFM/U2120  ( .A(b_in[113]), .ZN(\GFM/n23970 ) );
INV_X4 \GFM/U2119  ( .A(b_in[117]), .ZN(\GFM/n24360 ) );
INV_X4 \GFM/U2118  ( .A(b_in[118]), .ZN(\GFM/n24460 ) );
INV_X4 \GFM/U2117  ( .A(b_in[120]), .ZN(\GFM/n2466 ) );
INV_X4 \GFM/U2116  ( .A(b_in[119]), .ZN(\GFM/n24560 ) );
INV_X4 \GFM/U2115  ( .A(b_in[122]), .ZN(\GFM/n2486 ) );
INV_X4 \GFM/U2114  ( .A(b_in[121]), .ZN(\GFM/n24760 ) );
INV_X4 \GFM/U2113  ( .A(b_in[124]), .ZN(\GFM/n2506 ) );
NOR2_X2 \GFM/U2112  ( .A1(\GFM/n25210 ), .A2(\GFM/n26080 ), .ZN(\GFM/N996 ));
NOR2_X2 \GFM/U2111  ( .A1(\GFM/n25180 ), .A2(\GFM/n26070 ), .ZN(\GFM/N965 ));
NOR2_X2 \GFM/U2110  ( .A1(\GFM/n2525 ), .A2(\GFM/n26200 ), .ZN(\GFM/N1368 ));
NOR2_X2 \GFM/U2109  ( .A1(\GFM/n2525 ), .A2(\GFM/n26190 ), .ZN(\GFM/N1337 ));
NOR2_X2 \GFM/U2108  ( .A1(\GFM/n2399 ), .A2(\GFM/n2617 ), .ZN(\GFM/N926 ) );
NOR2_X2 \GFM/U2107  ( .A1(\GFM/n24120 ), .A2(\GFM/n2618 ), .ZN(\GFM/N985 ));
NOR2_X2 \GFM/U2106  ( .A1(\GFM/n24080 ), .A2(\GFM/n26120 ), .ZN(\GFM/N799 ));
NOR2_X2 \GFM/U2105  ( .A1(\GFM/n2409 ), .A2(\GFM/n2613 ), .ZN(\GFM/N830 ) );
NOR2_X2 \GFM/U2104  ( .A1(\GFM/n24080 ), .A2(\GFM/n2616 ), .ZN(\GFM/N923 ));
NOR2_X2 \GFM/U2103  ( .A1(\GFM/n24650 ), .A2(\GFM/n2616 ), .ZN(\GFM/N1074 ));
NOR2_X2 \GFM/U2102  ( .A1(\GFM/n24080 ), .A2(\GFM/n26140 ), .ZN(\GFM/N861 ));
NOR2_X2 \GFM/U2101  ( .A1(\GFM/n24080 ), .A2(\GFM/n26150 ), .ZN(\GFM/N892 ));
NOR2_X2 \GFM/U2100  ( .A1(\GFM/n24650 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1043 ));
NOR2_X2 \GFM/U2099  ( .A1(\GFM/n24080 ), .A2(\GFM/n26110 ), .ZN(\GFM/N768 ));
NOR2_X2 \GFM/U2098  ( .A1(\GFM/n24570 ), .A2(\GFM/n26110 ), .ZN(\GFM/N919 ));
NOR2_X2 \GFM/U2097  ( .A1(\GFM/n2525 ), .A2(\GFM/n26110 ), .ZN(\GFM/N1089 ));
NOR2_X2 \GFM/U2096  ( .A1(\GFM/n2416 ), .A2(\GFM/n25901 ), .ZN(\GFM/N117 ));
NOR2_X2 \GFM/U2095  ( .A1(\GFM/n2461 ), .A2(\GFM/n25901 ), .ZN(\GFM/N268 ));
NOR2_X2 \GFM/U2094  ( .A1(\GFM/n24120 ), .A2(\GFM/n2595 ), .ZN(\GFM/N272 ));
NOR2_X2 \GFM/U2093  ( .A1(\GFM/n24110 ), .A2(\GFM/n2596 ), .ZN(\GFM/N303 ));
NOR2_X2 \GFM/U2092  ( .A1(\GFM/n24101 ), .A2(\GFM/n25970 ), .ZN(\GFM/N334 ));
NOR2_X2 \GFM/U2091  ( .A1(\GFM/n24101 ), .A2(\GFM/n25980 ), .ZN(\GFM/N365 ));
NOR2_X2 \GFM/U2090  ( .A1(\GFM/n2409 ), .A2(\GFM/n2599 ), .ZN(\GFM/N396 ) );
NOR2_X2 \GFM/U2089  ( .A1(\GFM/n2509 ), .A2(\GFM/n25901 ), .ZN(\GFM/N411 ));
NOR2_X2 \GFM/U2088  ( .A1(\GFM/n2409 ), .A2(\GFM/n26000 ), .ZN(\GFM/N427 ));
NOR2_X2 \GFM/U2087  ( .A1(\GFM/n25080 ), .A2(\GFM/n25910 ), .ZN(\GFM/N442 ));
NOR2_X2 \GFM/U2086  ( .A1(\GFM/n2409 ), .A2(\GFM/n26010 ), .ZN(\GFM/N458 ));
NOR2_X2 \GFM/U2085  ( .A1(\GFM/n2509 ), .A2(\GFM/n2592 ), .ZN(\GFM/N473 ) );
NOR2_X2 \GFM/U2084  ( .A1(\GFM/n24080 ), .A2(\GFM/n2602 ), .ZN(\GFM/N489 ));
NOR2_X2 \GFM/U2083  ( .A1(\GFM/n2509 ), .A2(\GFM/n25930 ), .ZN(\GFM/N504 ));
NOR2_X2 \GFM/U2082  ( .A1(\GFM/n2409 ), .A2(\GFM/n2603 ), .ZN(\GFM/N520 ) );
NOR2_X2 \GFM/U2081  ( .A1(\GFM/n2509 ), .A2(\GFM/n25940 ), .ZN(\GFM/N535 ));
NOR2_X2 \GFM/U2080  ( .A1(\GFM/n24080 ), .A2(\GFM/n2604 ), .ZN(\GFM/N551 ));
NOR2_X2 \GFM/U2079  ( .A1(\GFM/n2399 ), .A2(\GFM/n26050 ), .ZN(\GFM/N554 ));
NOR2_X2 \GFM/U2078  ( .A1(\GFM/n25080 ), .A2(\GFM/n2595 ), .ZN(\GFM/N566 ));
NOR2_X2 \GFM/U2077  ( .A1(\GFM/n24080 ), .A2(\GFM/n26050 ), .ZN(\GFM/N582 ));
NOR2_X2 \GFM/U2076  ( .A1(\GFM/n2509 ), .A2(\GFM/n2596 ), .ZN(\GFM/N597 ) );
NOR2_X2 \GFM/U2075  ( .A1(\GFM/n25080 ), .A2(\GFM/n25970 ), .ZN(\GFM/N628 ));
NOR2_X2 \GFM/U2074  ( .A1(\GFM/n24570 ), .A2(\GFM/n2602 ), .ZN(\GFM/N640 ));
NOR2_X2 \GFM/U2073  ( .A1(\GFM/n25080 ), .A2(\GFM/n25980 ), .ZN(\GFM/N659 ));
NOR2_X2 \GFM/U2072  ( .A1(\GFM/n2458 ), .A2(\GFM/n2603 ), .ZN(\GFM/N671 ) );
NOR2_X2 \GFM/U2071  ( .A1(\GFM/n23980 ), .A2(\GFM/n2609 ), .ZN(\GFM/N678 ));
NOR2_X2 \GFM/U2070  ( .A1(\GFM/n25080 ), .A2(\GFM/n2599 ), .ZN(\GFM/N690 ));
NOR2_X2 \GFM/U2069  ( .A1(\GFM/n24080 ), .A2(\GFM/n2609 ), .ZN(\GFM/N706 ));
NOR2_X2 \GFM/U2068  ( .A1(\GFM/n24570 ), .A2(\GFM/n2604 ), .ZN(\GFM/N702 ));
NOR2_X2 \GFM/U2067  ( .A1(\GFM/n25080 ), .A2(\GFM/n26000 ), .ZN(\GFM/N721 ));
NOR2_X2 \GFM/U2066  ( .A1(\GFM/n2517 ), .A2(\GFM/n26000 ), .ZN(\GFM/N748 ));
NOR2_X2 \GFM/U2065  ( .A1(\GFM/n25080 ), .A2(\GFM/n2602 ), .ZN(\GFM/N783 ));
NOR2_X2 \GFM/U2064  ( .A1(\GFM/n25180 ), .A2(\GFM/n2602 ), .ZN(\GFM/N810 ));
NOR2_X2 \GFM/U2063  ( .A1(\GFM/n24570 ), .A2(\GFM/n2609 ), .ZN(\GFM/N857 ));
NOR2_X2 \GFM/U2062  ( .A1(\GFM/n25080 ), .A2(\GFM/n26050 ), .ZN(\GFM/N876 ));
NOR2_X2 \GFM/U2061  ( .A1(\GFM/n24770 ), .A2(\GFM/n2609 ), .ZN(\GFM/N910 ));
NOR2_X2 \GFM/U2060  ( .A1(\GFM/n2511 ), .A2(\GFM/n2609 ), .ZN(\GFM/N1000 ));
NOR2_X2 \GFM/U2059  ( .A1(\GFM/n2517 ), .A2(\GFM/n2609 ), .ZN(\GFM/N1027 ));
NOR2_X2 \GFM/U2058  ( .A1(\GFM/n24080 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1078 ));
NOR2_X2 \GFM/U2057  ( .A1(\GFM/n2416 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1109 ));
NOR2_X2 \GFM/U2056  ( .A1(\GFM/n2416 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1140 ));
NOR2_X2 \GFM/U2055  ( .A1(\GFM/n2416 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1171 ));
NOR2_X2 \GFM/U2054  ( .A1(\GFM/n2455 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1194 ));
NOR2_X2 \GFM/U2053  ( .A1(\GFM/n2416 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1202 ));
NOR2_X2 \GFM/U2052  ( .A1(\GFM/n2455 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1225 ));
NOR2_X2 \GFM/U2051  ( .A1(\GFM/n24650 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1229 ));
NOR2_X2 \GFM/U2050  ( .A1(\GFM/n2416 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1233 ));
NOR2_X2 \GFM/U2049  ( .A1(\GFM/n2455 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1256 ));
NOR2_X2 \GFM/U2048  ( .A1(\GFM/n2416 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1264 ));
NOR2_X2 \GFM/U2047  ( .A1(\GFM/n2455 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1287 ));
NOR2_X2 \GFM/U2046  ( .A1(\GFM/n2416 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1295 ));
NOR2_X2 \GFM/U2045  ( .A1(\GFM/n2416 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1326 ));
NOR2_X2 \GFM/U2044  ( .A1(\GFM/n2416 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1357 ));
NOR2_X2 \GFM/U2043  ( .A1(\GFM/n2416 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1388 ));
NOR2_X2 \GFM/U2042  ( .A1(\GFM/n2524 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1399 ));
NOR2_X2 \GFM/U2041  ( .A1(\GFM/n24150 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1419 ));
NOR2_X2 \GFM/U2040  ( .A1(\GFM/n2524 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1430 ));
NOR2_X2 \GFM/U2039  ( .A1(\GFM/n24150 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1450 ));
NOR2_X2 \GFM/U2038  ( .A1(\GFM/n2524 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1461 ));
NOR2_X2 \GFM/U2037  ( .A1(\GFM/n24150 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1481 ));
NOR2_X2 \GFM/U2036  ( .A1(\GFM/n2524 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1492 ));
NOR2_X2 \GFM/U2035  ( .A1(\GFM/n24150 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1512 ));
NOR2_X2 \GFM/U2034  ( .A1(\GFM/n2524 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1523 ));
NOR2_X2 \GFM/U2033  ( .A1(\GFM/n24150 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1543 ));
NOR2_X2 \GFM/U2032  ( .A1(\GFM/n2524 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1554 ));
NOR2_X2 \GFM/U2031  ( .A1(\GFM/n24150 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1574 ));
NOR2_X2 \GFM/U2030  ( .A1(\GFM/n2524 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1585 ));
NOR2_X2 \GFM/U2029  ( .A1(\GFM/n24150 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1605 ));
NOR2_X2 \GFM/U2028  ( .A1(\GFM/n25150 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1620 ));
NOR2_X2 \GFM/U2027  ( .A1(\GFM/n24150 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1636 ));
NOR2_X2 \GFM/U2026  ( .A1(\GFM/n25150 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1651 ));
NOR2_X2 \GFM/U2025  ( .A1(\GFM/n24150 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1667 ));
NOR2_X2 \GFM/U2024  ( .A1(\GFM/n25140 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1682 ));
NOR2_X2 \GFM/U2023  ( .A1(\GFM/n24150 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1698 ));
NOR2_X2 \GFM/U2022  ( .A1(\GFM/n25140 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1713 ));
NOR2_X2 \GFM/U2021  ( .A1(\GFM/n24150 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1729 ));
NOR2_X2 \GFM/U2020  ( .A1(\GFM/n25140 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1744 ));
NOR2_X2 \GFM/U2019  ( .A1(\GFM/n24150 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1760 ));
NOR2_X2 \GFM/U2018  ( .A1(\GFM/n25140 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1775 ));
NOR2_X2 \GFM/U2017  ( .A1(\GFM/n24140 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1791 ));
NOR2_X2 \GFM/U2016  ( .A1(\GFM/n25140 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1806 ));
NOR2_X2 \GFM/U2015  ( .A1(\GFM/n24140 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1822 ));
NOR2_X2 \GFM/U2014  ( .A1(\GFM/n25140 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1837 ));
NOR2_X2 \GFM/U2013  ( .A1(\GFM/n24140 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1853 ));
NOR2_X2 \GFM/U2012  ( .A1(\GFM/n25140 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1868 ));
NOR2_X2 \GFM/U2011  ( .A1(\GFM/n24140 ), .A2(\GFM/n2647 ), .ZN(\GFM/N1884 ));
NOR2_X2 \GFM/U2010  ( .A1(\GFM/n25140 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1899 ));
NOR2_X2 \GFM/U2009  ( .A1(\GFM/n24140 ), .A2(\GFM/n2648 ), .ZN(\GFM/N1915 ));
NOR2_X2 \GFM/U2008  ( .A1(\GFM/n25140 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1930 ));
NOR2_X2 \GFM/U2007  ( .A1(\GFM/n24140 ), .A2(\GFM/n2649 ), .ZN(\GFM/N1946 ));
NOR2_X2 \GFM/U2006  ( .A1(\GFM/n25140 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1961 ));
NOR2_X2 \GFM/U2005  ( .A1(\GFM/n24140 ), .A2(\GFM/n26500 ), .ZN(\GFM/N1977 ));
NOR2_X2 \GFM/U2004  ( .A1(\GFM/n25140 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1992 ));
NOR2_X2 \GFM/U2003  ( .A1(\GFM/n24140 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2008 ));
NOR2_X2 \GFM/U2002  ( .A1(\GFM/n25140 ), .A2(\GFM/n26420 ), .ZN(\GFM/N2023 ));
NOR2_X2 \GFM/U2001  ( .A1(\GFM/n24140 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2039 ));
NOR2_X2 \GFM/U2000  ( .A1(\GFM/n2513 ), .A2(\GFM/n26430 ), .ZN(\GFM/N2054 ));
NOR2_X2 \GFM/U1999  ( .A1(\GFM/n24140 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2070 ));
NOR2_X2 \GFM/U1998  ( .A1(\GFM/n2513 ), .A2(\GFM/n2644 ), .ZN(\GFM/N2085 ));
NOR2_X2 \GFM/U1997  ( .A1(\GFM/n24140 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2101 ));
NOR2_X2 \GFM/U1996  ( .A1(\GFM/n2513 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2116 ));
NOR2_X2 \GFM/U1995  ( .A1(\GFM/n2413 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2132 ));
NOR2_X2 \GFM/U1994  ( .A1(\GFM/n2513 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2147 ));
NOR2_X2 \GFM/U1993  ( .A1(\GFM/n2413 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2163 ));
NOR2_X2 \GFM/U1992  ( .A1(\GFM/n2513 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2178 ));
NOR2_X2 \GFM/U1991  ( .A1(\GFM/n2413 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2194 ));
NOR2_X2 \GFM/U1990  ( .A1(\GFM/n2513 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2209 ));
NOR2_X2 \GFM/U1989  ( .A1(\GFM/n2413 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2225 ));
NOR2_X2 \GFM/U1988  ( .A1(\GFM/n2513 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2240 ));
NOR2_X2 \GFM/U1987  ( .A1(\GFM/n2413 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2256 ));
NOR2_X2 \GFM/U1986  ( .A1(\GFM/n2513 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2271 ));
NOR2_X2 \GFM/U1985  ( .A1(\GFM/n2413 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2287 ));
NOR2_X2 \GFM/U1984  ( .A1(\GFM/n2513 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2302 ));
NOR2_X2 \GFM/U1983  ( .A1(\GFM/n2413 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2318 ));
NOR2_X2 \GFM/U1982  ( .A1(\GFM/n2513 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2333 ));
NOR2_X2 \GFM/U1981  ( .A1(\GFM/n2413 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2349 ));
NOR2_X2 \GFM/U1980  ( .A1(\GFM/n2513 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2364 ));
NOR2_X2 \GFM/U1979  ( .A1(\GFM/n2413 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2380 ));
NOR2_X2 \GFM/U1978  ( .A1(\GFM/n2513 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2395 ));
NOR2_X2 \GFM/U1977  ( .A1(\GFM/n2413 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2411 ));
NOR2_X2 \GFM/U1976  ( .A1(\GFM/n25120 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2426 ));
NOR2_X2 \GFM/U1975  ( .A1(\GFM/n2413 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2442 ));
NOR2_X2 \GFM/U1974  ( .A1(\GFM/n25120 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2457 ));
NOR2_X2 \GFM/U1973  ( .A1(\GFM/n24120 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2473 ));
NOR2_X2 \GFM/U1972  ( .A1(\GFM/n25120 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2488 ));
NOR2_X2 \GFM/U1971  ( .A1(\GFM/n24120 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2504 ));
NOR2_X2 \GFM/U1970  ( .A1(\GFM/n25120 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2519 ));
NOR2_X2 \GFM/U1969  ( .A1(\GFM/n24120 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2535 ));
NOR2_X2 \GFM/U1968  ( .A1(\GFM/n25120 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2550 ));
NOR2_X2 \GFM/U1967  ( .A1(\GFM/n24120 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2566 ));
NOR2_X2 \GFM/U1966  ( .A1(\GFM/n25120 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2581 ));
NOR2_X2 \GFM/U1965  ( .A1(\GFM/n24120 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2597 ));
NOR2_X2 \GFM/U1964  ( .A1(\GFM/n25120 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2612 ));
NOR2_X2 \GFM/U1963  ( .A1(\GFM/n24120 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2628 ));
NOR2_X2 \GFM/U1962  ( .A1(\GFM/n25120 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2643 ));
NOR2_X2 \GFM/U1961  ( .A1(\GFM/n25120 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2674 ));
NOR2_X2 \GFM/U1960  ( .A1(\GFM/n25120 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2705 ));
NOR2_X2 \GFM/U1959  ( .A1(\GFM/n25120 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2736 ));
NOR2_X2 \GFM/U1958  ( .A1(\GFM/n25120 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2767 ));
NOR2_X2 \GFM/U1957  ( .A1(\GFM/n2511 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2798 ));
NOR2_X2 \GFM/U1956  ( .A1(\GFM/n2511 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2829 ));
NOR2_X2 \GFM/U1955  ( .A1(\GFM/n2511 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2860 ));
NOR2_X2 \GFM/U1954  ( .A1(\GFM/n2511 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2891 ));
NOR2_X2 \GFM/U1953  ( .A1(\GFM/n2511 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2922 ));
NOR2_X2 \GFM/U1952  ( .A1(\GFM/n24120 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2659 ));
NOR2_X2 \GFM/U1951  ( .A1(\GFM/n24120 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2690 ));
NOR2_X2 \GFM/U1950  ( .A1(\GFM/n24120 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2721 ));
NOR2_X2 \GFM/U1949  ( .A1(\GFM/n24120 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2752 ));
NOR2_X2 \GFM/U1948  ( .A1(\GFM/n24120 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2783 ));
NOR2_X2 \GFM/U1947  ( .A1(\GFM/n24110 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2814 ));
NOR2_X2 \GFM/U1946  ( .A1(\GFM/n24110 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2845 ));
NOR2_X2 \GFM/U1945  ( .A1(\GFM/n24110 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2876 ));
NOR2_X2 \GFM/U1944  ( .A1(\GFM/n24110 ), .A2(\GFM/n26801 ), .ZN(\GFM/N2907 ));
NOR2_X2 \GFM/U1943  ( .A1(\GFM/n24110 ), .A2(\GFM/n26810 ), .ZN(\GFM/N2938 ));
NOR2_X2 \GFM/U1942  ( .A1(\GFM/n2511 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2953 ));
NOR2_X2 \GFM/U1941  ( .A1(\GFM/n24110 ), .A2(\GFM/n26820 ), .ZN(\GFM/N2969 ));
NOR2_X2 \GFM/U1940  ( .A1(\GFM/n2511 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2984 ));
NOR2_X2 \GFM/U1939  ( .A1(\GFM/n24110 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3000 ));
NOR2_X2 \GFM/U1938  ( .A1(\GFM/n2511 ), .A2(\GFM/n26740 ), .ZN(\GFM/N3015 ));
NOR2_X2 \GFM/U1937  ( .A1(\GFM/n24110 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3031 ));
NOR2_X2 \GFM/U1936  ( .A1(\GFM/n2511 ), .A2(\GFM/n2675 ), .ZN(\GFM/N3046 ));
NOR2_X2 \GFM/U1935  ( .A1(\GFM/n24110 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3062 ));
NOR2_X2 \GFM/U1934  ( .A1(\GFM/n2511 ), .A2(\GFM/n26760 ), .ZN(\GFM/N3077 ));
NOR2_X2 \GFM/U1933  ( .A1(\GFM/n24110 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3093 ));
NOR2_X2 \GFM/U1932  ( .A1(\GFM/n2511 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3108 ));
NOR2_X2 \GFM/U1931  ( .A1(\GFM/n24110 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3124 ));
NOR2_X2 \GFM/U1930  ( .A1(\GFM/n25101 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3139 ));
NOR2_X2 \GFM/U1929  ( .A1(\GFM/n24110 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3155 ));
NOR2_X2 \GFM/U1928  ( .A1(\GFM/n25101 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3170 ));
NOR2_X2 \GFM/U1927  ( .A1(\GFM/n24101 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3186 ));
NOR2_X2 \GFM/U1926  ( .A1(\GFM/n25101 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3201 ));
NOR2_X2 \GFM/U1925  ( .A1(\GFM/n24101 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3217 ));
NOR2_X2 \GFM/U1924  ( .A1(\GFM/n25101 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3232 ));
NOR2_X2 \GFM/U1923  ( .A1(\GFM/n24101 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3248 ));
NOR2_X2 \GFM/U1922  ( .A1(\GFM/n25101 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3263 ));
NOR2_X2 \GFM/U1921  ( .A1(\GFM/n24101 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3279 ));
NOR2_X2 \GFM/U1920  ( .A1(\GFM/n24900 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3294 ));
NOR2_X2 \GFM/U1919  ( .A1(\GFM/n24590 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3309 ));
NOR2_X2 \GFM/U1918  ( .A1(\GFM/n24101 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3313 ));
NOR2_X2 \GFM/U1917  ( .A1(\GFM/n24900 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3326 ));
NOR2_X2 \GFM/U1916  ( .A1(\GFM/n24101 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3346 ));
NOR2_X2 \GFM/U1915  ( .A1(\GFM/n24590 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3341 ));
NOR2_X2 \GFM/U1914  ( .A1(\GFM/n24900 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3359 ));
NOR2_X2 \GFM/U1913  ( .A1(\GFM/n24590 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3374 ));
NOR2_X2 \GFM/U1912  ( .A1(\GFM/n24900 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3393 ));
NOR2_X2 \GFM/U1911  ( .A1(\GFM/n24290 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3402 ));
NOR2_X2 \GFM/U1910  ( .A1(\GFM/n24900 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3429 ));
NOR2_X2 \GFM/U1909  ( .A1(\GFM/n24590 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3514 ));
NOR2_X2 \GFM/U1908  ( .A1(\GFM/n25000 ), .A2(\GFM/n2610 ), .ZN(\GFM/N999 ));
NOR2_X2 \GFM/U1907  ( .A1(\GFM/n2497 ), .A2(\GFM/n26080 ), .ZN(\GFM/N937 ));
NOR2_X2 \GFM/U1906  ( .A1(\GFM/n2497 ), .A2(\GFM/n2606 ), .ZN(\GFM/N875 ) );
NOR2_X2 \GFM/U1905  ( .A1(\GFM/n25050 ), .A2(\GFM/n26200 ), .ZN(\GFM/N1309 ));
NOR2_X2 \GFM/U1904  ( .A1(\GFM/n25050 ), .A2(\GFM/n26190 ), .ZN(\GFM/N1278 ));
NOR2_X2 \GFM/U1903  ( .A1(\GFM/n2525 ), .A2(\GFM/n2617 ), .ZN(\GFM/N1275 ));
NOR2_X2 \GFM/U1902  ( .A1(\GFM/n25050 ), .A2(\GFM/n2617 ), .ZN(\GFM/N1216 ));
NOR2_X2 \GFM/U1901  ( .A1(\GFM/n2525 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1213 ));
NOR2_X2 \GFM/U1900  ( .A1(\GFM/n24210 ), .A2(\GFM/n2617 ), .ZN(\GFM/N986 ));
NOR2_X2 \GFM/U1899  ( .A1(\GFM/n2417 ), .A2(\GFM/n2618 ), .ZN(\GFM/N1017 ));
NOR2_X2 \GFM/U1898  ( .A1(\GFM/n2417 ), .A2(\GFM/n26120 ), .ZN(\GFM/N831 ));
NOR2_X2 \GFM/U1897  ( .A1(\GFM/n2471 ), .A2(\GFM/n26120 ), .ZN(\GFM/N982 ));
NOR2_X2 \GFM/U1896  ( .A1(\GFM/n25050 ), .A2(\GFM/n26120 ), .ZN(\GFM/N1061 ));
NOR2_X2 \GFM/U1895  ( .A1(\GFM/n2417 ), .A2(\GFM/n2613 ), .ZN(\GFM/N862 ) );
NOR2_X2 \GFM/U1894  ( .A1(\GFM/n24670 ), .A2(\GFM/n2613 ), .ZN(\GFM/N1013 ));
NOR2_X2 \GFM/U1893  ( .A1(\GFM/n25050 ), .A2(\GFM/n2613 ), .ZN(\GFM/N1092 ));
NOR2_X2 \GFM/U1892  ( .A1(\GFM/n2431 ), .A2(\GFM/n2616 ), .ZN(\GFM/N979 ) );
NOR2_X2 \GFM/U1891  ( .A1(\GFM/n24511 ), .A2(\GFM/n26140 ), .ZN(\GFM/N977 ));
NOR2_X2 \GFM/U1890  ( .A1(\GFM/n25050 ), .A2(\GFM/n2616 ), .ZN(\GFM/N1185 ));
NOR2_X2 \GFM/U1889  ( .A1(\GFM/n2525 ), .A2(\GFM/n26140 ), .ZN(\GFM/N1182 ));
NOR2_X2 \GFM/U1888  ( .A1(\GFM/n2417 ), .A2(\GFM/n2616 ), .ZN(\GFM/N955 ) );
NOR2_X2 \GFM/U1887  ( .A1(\GFM/n2475 ), .A2(\GFM/n2616 ), .ZN(\GFM/N1106 ));
NOR2_X2 \GFM/U1886  ( .A1(\GFM/n25050 ), .A2(\GFM/n26140 ), .ZN(\GFM/N1123 ));
NOR2_X2 \GFM/U1885  ( .A1(\GFM/n2525 ), .A2(\GFM/n26120 ), .ZN(\GFM/N1120 ));
NOR2_X2 \GFM/U1884  ( .A1(\GFM/n2417 ), .A2(\GFM/n26140 ), .ZN(\GFM/N893 ));
NOR2_X2 \GFM/U1883  ( .A1(\GFM/n2427 ), .A2(\GFM/n26140 ), .ZN(\GFM/N917 ));
NOR2_X2 \GFM/U1882  ( .A1(\GFM/n2475 ), .A2(\GFM/n26140 ), .ZN(\GFM/N1044 ));
NOR2_X2 \GFM/U1881  ( .A1(\GFM/n26980 ), .A2(\GFM/n25070 ), .ZN(\GFM/N4052 ));
NOR2_X2 \GFM/U1880  ( .A1(\GFM/n2427 ), .A2(\GFM/n26150 ), .ZN(\GFM/N948 ));
NOR2_X2 \GFM/U1879  ( .A1(\GFM/n2613 ), .A2(\GFM/n24460 ), .ZN(\GFM/N946 ));
NOR2_X2 \GFM/U1878  ( .A1(\GFM/n25050 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1154 ));
NOR2_X2 \GFM/U1877  ( .A1(\GFM/n2525 ), .A2(\GFM/n2613 ), .ZN(\GFM/N1151 ));
NOR2_X2 \GFM/U1876  ( .A1(\GFM/n2417 ), .A2(\GFM/n26150 ), .ZN(\GFM/N924 ));
NOR2_X2 \GFM/U1875  ( .A1(\GFM/n2475 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1075 ));
NOR2_X2 \GFM/U1874  ( .A1(\GFM/n2417 ), .A2(\GFM/n26110 ), .ZN(\GFM/N800 ));
NOR2_X2 \GFM/U1873  ( .A1(\GFM/n2437 ), .A2(\GFM/n26110 ), .ZN(\GFM/N852 ));
NOR2_X2 \GFM/U1872  ( .A1(\GFM/n24670 ), .A2(\GFM/n26110 ), .ZN(\GFM/N951 ));
NOR2_X2 \GFM/U1871  ( .A1(\GFM/n25050 ), .A2(\GFM/n26110 ), .ZN(\GFM/N1030 ));
NOR2_X2 \GFM/U1870  ( .A1(\GFM/n24330 ), .A2(\GFM/n25910 ), .ZN(\GFM/N204 ));
NOR2_X2 \GFM/U1869  ( .A1(\GFM/n25890 ), .A2(\GFM/n2447 ), .ZN(\GFM/N202 ));
NOR2_X2 \GFM/U1868  ( .A1(\GFM/n2427 ), .A2(\GFM/n2604 ), .ZN(\GFM/N607 ) );
NOR2_X2 \GFM/U1867  ( .A1(\GFM/n2448 ), .A2(\GFM/n2602 ), .ZN(\GFM/N605 ) );
NOR2_X2 \GFM/U1866  ( .A1(\GFM/n2427 ), .A2(\GFM/n26050 ), .ZN(\GFM/N638 ));
NOR2_X2 \GFM/U1865  ( .A1(\GFM/n2447 ), .A2(\GFM/n2603 ), .ZN(\GFM/N636 ) );
NOR2_X2 \GFM/U1864  ( .A1(\GFM/n2435 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1320 ));
NOR2_X2 \GFM/U1863  ( .A1(\GFM/n2455 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1318 ));
NOR2_X2 \GFM/U1862  ( .A1(\GFM/n2435 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1351 ));
NOR2_X2 \GFM/U1861  ( .A1(\GFM/n2455 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1349 ));
NOR2_X2 \GFM/U1860  ( .A1(\GFM/n2435 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1382 ));
NOR2_X2 \GFM/U1859  ( .A1(\GFM/n2455 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1380 ));
NOR2_X2 \GFM/U1858  ( .A1(\GFM/n2435 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1413 ));
NOR2_X2 \GFM/U1857  ( .A1(\GFM/n2455 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1411 ));
NOR2_X2 \GFM/U1856  ( .A1(\GFM/n2435 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1444 ));
NOR2_X2 \GFM/U1855  ( .A1(\GFM/n2455 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1442 ));
NOR2_X2 \GFM/U1854  ( .A1(\GFM/n2435 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1475 ));
NOR2_X2 \GFM/U1853  ( .A1(\GFM/n2455 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1473 ));
NOR2_X2 \GFM/U1852  ( .A1(\GFM/n2435 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1506 ));
NOR2_X2 \GFM/U1851  ( .A1(\GFM/n2454 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1504 ));
NOR2_X2 \GFM/U1850  ( .A1(\GFM/n24330 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2002 ));
NOR2_X2 \GFM/U1849  ( .A1(\GFM/n24530 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2000 ));
NOR2_X2 \GFM/U1848  ( .A1(\GFM/n24330 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2033 ));
NOR2_X2 \GFM/U1847  ( .A1(\GFM/n24530 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2031 ));
NOR2_X2 \GFM/U1846  ( .A1(\GFM/n24330 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2064 ));
NOR2_X2 \GFM/U1845  ( .A1(\GFM/n24530 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2062 ));
NOR2_X2 \GFM/U1844  ( .A1(\GFM/n2396 ), .A2(\GFM/n2592 ), .ZN(\GFM/N121 ) );
NOR2_X2 \GFM/U1843  ( .A1(\GFM/n2424 ), .A2(\GFM/n25901 ), .ZN(\GFM/N149 ));
NOR2_X2 \GFM/U1842  ( .A1(\GFM/n2423 ), .A2(\GFM/n25910 ), .ZN(\GFM/N180 ));
NOR2_X2 \GFM/U1841  ( .A1(\GFM/n2423 ), .A2(\GFM/n2592 ), .ZN(\GFM/N211 ) );
NOR2_X2 \GFM/U1840  ( .A1(\GFM/n24220 ), .A2(\GFM/n25930 ), .ZN(\GFM/N242 ));
NOR2_X2 \GFM/U1839  ( .A1(\GFM/n24210 ), .A2(\GFM/n25940 ), .ZN(\GFM/N273 ));
NOR2_X2 \GFM/U1838  ( .A1(\GFM/n23910 ), .A2(\GFM/n25970 ), .ZN(\GFM/N276 ));
NOR2_X2 \GFM/U1837  ( .A1(\GFM/n24700 ), .A2(\GFM/n25901 ), .ZN(\GFM/N300 ));
NOR2_X2 \GFM/U1836  ( .A1(\GFM/n24201 ), .A2(\GFM/n2595 ), .ZN(\GFM/N304 ));
NOR2_X2 \GFM/U1835  ( .A1(\GFM/n23910 ), .A2(\GFM/n25980 ), .ZN(\GFM/N307 ));
NOR2_X2 \GFM/U1834  ( .A1(\GFM/n24690 ), .A2(\GFM/n25910 ), .ZN(\GFM/N331 ));
NOR2_X2 \GFM/U1833  ( .A1(\GFM/n24190 ), .A2(\GFM/n2596 ), .ZN(\GFM/N335 ));
NOR2_X2 \GFM/U1832  ( .A1(\GFM/n23900 ), .A2(\GFM/n2599 ), .ZN(\GFM/N338 ));
NOR2_X2 \GFM/U1831  ( .A1(\GFM/n2489 ), .A2(\GFM/n25901 ), .ZN(\GFM/N351 ));
NOR2_X2 \GFM/U1830  ( .A1(\GFM/n24690 ), .A2(\GFM/n2592 ), .ZN(\GFM/N362 ));
NOR2_X2 \GFM/U1829  ( .A1(\GFM/n24190 ), .A2(\GFM/n25970 ), .ZN(\GFM/N366 ));
NOR2_X2 \GFM/U1828  ( .A1(\GFM/n23900 ), .A2(\GFM/n26000 ), .ZN(\GFM/N369 ));
NOR2_X2 \GFM/U1827  ( .A1(\GFM/n24980 ), .A2(\GFM/n25901 ), .ZN(\GFM/N379 ));
NOR2_X2 \GFM/U1826  ( .A1(\GFM/n24910 ), .A2(\GFM/n25910 ), .ZN(\GFM/N382 ));
NOR2_X2 \GFM/U1825  ( .A1(\GFM/n2468 ), .A2(\GFM/n25930 ), .ZN(\GFM/N393 ));
NOR2_X2 \GFM/U1824  ( .A1(\GFM/n2418 ), .A2(\GFM/n25980 ), .ZN(\GFM/N397 ));
NOR2_X2 \GFM/U1823  ( .A1(\GFM/n2389 ), .A2(\GFM/n26010 ), .ZN(\GFM/N400 ));
NOR2_X2 \GFM/U1822  ( .A1(\GFM/n24980 ), .A2(\GFM/n25910 ), .ZN(\GFM/N410 ));
NOR2_X2 \GFM/U1821  ( .A1(\GFM/n2489 ), .A2(\GFM/n2592 ), .ZN(\GFM/N413 ) );
NOR2_X2 \GFM/U1820  ( .A1(\GFM/n24690 ), .A2(\GFM/n25940 ), .ZN(\GFM/N424 ));
NOR2_X2 \GFM/U1819  ( .A1(\GFM/n2418 ), .A2(\GFM/n2599 ), .ZN(\GFM/N428 ) );
NOR2_X2 \GFM/U1818  ( .A1(\GFM/n2389 ), .A2(\GFM/n2602 ), .ZN(\GFM/N431 ) );
NOR2_X2 \GFM/U1817  ( .A1(\GFM/n24980 ), .A2(\GFM/n2592 ), .ZN(\GFM/N441 ));
NOR2_X2 \GFM/U1816  ( .A1(\GFM/n2489 ), .A2(\GFM/n25930 ), .ZN(\GFM/N444 ));
NOR2_X2 \GFM/U1815  ( .A1(\GFM/n2468 ), .A2(\GFM/n2595 ), .ZN(\GFM/N455 ) );
NOR2_X2 \GFM/U1814  ( .A1(\GFM/n2418 ), .A2(\GFM/n26000 ), .ZN(\GFM/N459 ));
NOR2_X2 \GFM/U1813  ( .A1(\GFM/n23880 ), .A2(\GFM/n2603 ), .ZN(\GFM/N462 ));
NOR2_X2 \GFM/U1812  ( .A1(\GFM/n2497 ), .A2(\GFM/n25930 ), .ZN(\GFM/N472 ));
NOR2_X2 \GFM/U1811  ( .A1(\GFM/n24880 ), .A2(\GFM/n25940 ), .ZN(\GFM/N475 ));
NOR2_X2 \GFM/U1810  ( .A1(\GFM/n2468 ), .A2(\GFM/n2596 ), .ZN(\GFM/N486 ) );
NOR2_X2 \GFM/U1809  ( .A1(\GFM/n2417 ), .A2(\GFM/n26010 ), .ZN(\GFM/N490 ));
NOR2_X2 \GFM/U1808  ( .A1(\GFM/n23880 ), .A2(\GFM/n2604 ), .ZN(\GFM/N493 ));
NOR2_X2 \GFM/U1807  ( .A1(\GFM/n24980 ), .A2(\GFM/n25940 ), .ZN(\GFM/N503 ));
NOR2_X2 \GFM/U1806  ( .A1(\GFM/n24880 ), .A2(\GFM/n2595 ), .ZN(\GFM/N506 ));
NOR2_X2 \GFM/U1805  ( .A1(\GFM/n2468 ), .A2(\GFM/n25970 ), .ZN(\GFM/N517 ));
NOR2_X2 \GFM/U1804  ( .A1(\GFM/n2418 ), .A2(\GFM/n2602 ), .ZN(\GFM/N521 ) );
NOR2_X2 \GFM/U1803  ( .A1(\GFM/n24980 ), .A2(\GFM/n2595 ), .ZN(\GFM/N534 ));
NOR2_X2 \GFM/U1802  ( .A1(\GFM/n24880 ), .A2(\GFM/n2596 ), .ZN(\GFM/N537 ));
NOR2_X2 \GFM/U1801  ( .A1(\GFM/n2468 ), .A2(\GFM/n25980 ), .ZN(\GFM/N548 ));
NOR2_X2 \GFM/U1800  ( .A1(\GFM/n2418 ), .A2(\GFM/n2603 ), .ZN(\GFM/N552 ) );
NOR2_X2 \GFM/U1799  ( .A1(\GFM/n2497 ), .A2(\GFM/n2596 ), .ZN(\GFM/N565 ) );
NOR2_X2 \GFM/U1798  ( .A1(\GFM/n24880 ), .A2(\GFM/n25970 ), .ZN(\GFM/N568 ));
NOR2_X2 \GFM/U1797  ( .A1(\GFM/n24670 ), .A2(\GFM/n2599 ), .ZN(\GFM/N579 ));
NOR2_X2 \GFM/U1796  ( .A1(\GFM/n2417 ), .A2(\GFM/n2604 ), .ZN(\GFM/N583 ) );
NOR2_X2 \GFM/U1795  ( .A1(\GFM/n2497 ), .A2(\GFM/n25970 ), .ZN(\GFM/N596 ));
NOR2_X2 \GFM/U1794  ( .A1(\GFM/n24880 ), .A2(\GFM/n25980 ), .ZN(\GFM/N599 ));
NOR2_X2 \GFM/U1793  ( .A1(\GFM/n24670 ), .A2(\GFM/n26000 ), .ZN(\GFM/N610 ));
NOR2_X2 \GFM/U1792  ( .A1(\GFM/n2417 ), .A2(\GFM/n26050 ), .ZN(\GFM/N614 ));
NOR2_X2 \GFM/U1791  ( .A1(\GFM/n24980 ), .A2(\GFM/n25980 ), .ZN(\GFM/N627 ));
NOR2_X2 \GFM/U1790  ( .A1(\GFM/n24880 ), .A2(\GFM/n2599 ), .ZN(\GFM/N630 ));
NOR2_X2 \GFM/U1789  ( .A1(\GFM/n24670 ), .A2(\GFM/n26010 ), .ZN(\GFM/N641 ));
NOR2_X2 \GFM/U1788  ( .A1(\GFM/n2497 ), .A2(\GFM/n2599 ), .ZN(\GFM/N658 ) );
NOR2_X2 \GFM/U1787  ( .A1(\GFM/n24880 ), .A2(\GFM/n26000 ), .ZN(\GFM/N661 ));
NOR2_X2 \GFM/U1786  ( .A1(\GFM/n2468 ), .A2(\GFM/n2602 ), .ZN(\GFM/N672 ) );
NOR2_X2 \GFM/U1785  ( .A1(\GFM/n2497 ), .A2(\GFM/n26000 ), .ZN(\GFM/N689 ));
NOR2_X2 \GFM/U1784  ( .A1(\GFM/n24880 ), .A2(\GFM/n26010 ), .ZN(\GFM/N692 ));
NOR2_X2 \GFM/U1783  ( .A1(\GFM/n24670 ), .A2(\GFM/n2603 ), .ZN(\GFM/N703 ));
NOR2_X2 \GFM/U1782  ( .A1(\GFM/n2497 ), .A2(\GFM/n26010 ), .ZN(\GFM/N720 ));
NOR2_X2 \GFM/U1781  ( .A1(\GFM/n24880 ), .A2(\GFM/n2602 ), .ZN(\GFM/N723 ));
NOR2_X2 \GFM/U1780  ( .A1(\GFM/n2468 ), .A2(\GFM/n2604 ), .ZN(\GFM/N734 ) );
NOR2_X2 \GFM/U1779  ( .A1(\GFM/n2417 ), .A2(\GFM/n2609 ), .ZN(\GFM/N738 ) );
NOR2_X2 \GFM/U1778  ( .A1(\GFM/n24870 ), .A2(\GFM/n2603 ), .ZN(\GFM/N754 ));
NOR2_X2 \GFM/U1777  ( .A1(\GFM/n2497 ), .A2(\GFM/n2602 ), .ZN(\GFM/N751 ) );
NOR2_X2 \GFM/U1776  ( .A1(\GFM/n24670 ), .A2(\GFM/n26050 ), .ZN(\GFM/N765 ));
NOR2_X2 \GFM/U1775  ( .A1(\GFM/n2497 ), .A2(\GFM/n2603 ), .ZN(\GFM/N782 ) );
NOR2_X2 \GFM/U1774  ( .A1(\GFM/n2489 ), .A2(\GFM/n2604 ), .ZN(\GFM/N785 ) );
NOR2_X2 \GFM/U1773  ( .A1(\GFM/n24870 ), .A2(\GFM/n26050 ), .ZN(\GFM/N816 ));
NOR2_X2 \GFM/U1772  ( .A1(\GFM/n2497 ), .A2(\GFM/n2604 ), .ZN(\GFM/N813 ) );
NOR2_X2 \GFM/U1771  ( .A1(\GFM/n24670 ), .A2(\GFM/n2609 ), .ZN(\GFM/N889 ));
NOR2_X2 \GFM/U1770  ( .A1(\GFM/n24880 ), .A2(\GFM/n2609 ), .ZN(\GFM/N940 ));
NOR2_X2 \GFM/U1769  ( .A1(\GFM/n2387 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1020 ));
NOR2_X2 \GFM/U1768  ( .A1(\GFM/n2396 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1051 ));
NOR2_X2 \GFM/U1767  ( .A1(\GFM/n2396 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1082 ));
NOR2_X2 \GFM/U1766  ( .A1(\GFM/n24250 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1110 ));
NOR2_X2 \GFM/U1765  ( .A1(\GFM/n2396 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1113 ));
NOR2_X2 \GFM/U1764  ( .A1(\GFM/n2427 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1134 ));
NOR2_X2 \GFM/U1763  ( .A1(\GFM/n24250 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1141 ));
NOR2_X2 \GFM/U1762  ( .A1(\GFM/n2396 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1144 ));
NOR2_X2 \GFM/U1761  ( .A1(\GFM/n24450 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1162 ));
NOR2_X2 \GFM/U1760  ( .A1(\GFM/n2435 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1165 ));
NOR2_X2 \GFM/U1759  ( .A1(\GFM/n24250 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1172 ));
NOR2_X2 \GFM/U1758  ( .A1(\GFM/n2396 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1175 ));
NOR2_X2 \GFM/U1757  ( .A1(\GFM/n24450 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1193 ));
NOR2_X2 \GFM/U1756  ( .A1(\GFM/n2435 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1196 ));
NOR2_X2 \GFM/U1755  ( .A1(\GFM/n24250 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1203 ));
NOR2_X2 \GFM/U1754  ( .A1(\GFM/n2396 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1206 ));
NOR2_X2 \GFM/U1753  ( .A1(\GFM/n24450 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1224 ));
NOR2_X2 \GFM/U1752  ( .A1(\GFM/n2435 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1227 ));
NOR2_X2 \GFM/U1751  ( .A1(\GFM/n24250 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1234 ));
NOR2_X2 \GFM/U1750  ( .A1(\GFM/n2396 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1237 ));
NOR2_X2 \GFM/U1749  ( .A1(\GFM/n24450 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1255 ));
NOR2_X2 \GFM/U1748  ( .A1(\GFM/n2435 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1258 ));
NOR2_X2 \GFM/U1747  ( .A1(\GFM/n2475 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1261 ));
NOR2_X2 \GFM/U1746  ( .A1(\GFM/n24250 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1265 ));
NOR2_X2 \GFM/U1745  ( .A1(\GFM/n2396 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1268 ));
NOR2_X2 \GFM/U1744  ( .A1(\GFM/n24450 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1286 ));
NOR2_X2 \GFM/U1743  ( .A1(\GFM/n2435 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1289 ));
NOR2_X2 \GFM/U1742  ( .A1(\GFM/n2475 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1292 ));
NOR2_X2 \GFM/U1741  ( .A1(\GFM/n24250 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1296 ));
NOR2_X2 \GFM/U1740  ( .A1(\GFM/n24950 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1312 ));
NOR2_X2 \GFM/U1739  ( .A1(\GFM/n2475 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1323 ));
NOR2_X2 \GFM/U1738  ( .A1(\GFM/n24250 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1327 ));
NOR2_X2 \GFM/U1737  ( .A1(\GFM/n24950 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1343 ));
NOR2_X2 \GFM/U1736  ( .A1(\GFM/n25040 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1340 ));
NOR2_X2 \GFM/U1735  ( .A1(\GFM/n2475 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1354 ));
NOR2_X2 \GFM/U1734  ( .A1(\GFM/n24250 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1358 ));
NOR2_X2 \GFM/U1733  ( .A1(\GFM/n24950 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1374 ));
NOR2_X2 \GFM/U1732  ( .A1(\GFM/n25040 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1371 ));
NOR2_X2 \GFM/U1731  ( .A1(\GFM/n2475 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1385 ));
NOR2_X2 \GFM/U1730  ( .A1(\GFM/n24250 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1389 ));
NOR2_X2 \GFM/U1729  ( .A1(\GFM/n24950 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1405 ));
NOR2_X2 \GFM/U1728  ( .A1(\GFM/n25040 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1402 ));
NOR2_X2 \GFM/U1727  ( .A1(\GFM/n2475 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1416 ));
NOR2_X2 \GFM/U1726  ( .A1(\GFM/n24250 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1420 ));
NOR2_X2 \GFM/U1725  ( .A1(\GFM/n24950 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1436 ));
NOR2_X2 \GFM/U1724  ( .A1(\GFM/n25040 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1433 ));
NOR2_X2 \GFM/U1723  ( .A1(\GFM/n2475 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1447 ));
NOR2_X2 \GFM/U1722  ( .A1(\GFM/n2424 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1451 ));
NOR2_X2 \GFM/U1721  ( .A1(\GFM/n24950 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1467 ));
NOR2_X2 \GFM/U1720  ( .A1(\GFM/n25040 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1464 ));
NOR2_X2 \GFM/U1719  ( .A1(\GFM/n24740 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1478 ));
NOR2_X2 \GFM/U1718  ( .A1(\GFM/n2424 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1482 ));
NOR2_X2 \GFM/U1717  ( .A1(\GFM/n24950 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1498 ));
NOR2_X2 \GFM/U1716  ( .A1(\GFM/n25040 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1495 ));
NOR2_X2 \GFM/U1715  ( .A1(\GFM/n24740 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1509 ));
NOR2_X2 \GFM/U1714  ( .A1(\GFM/n2424 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1513 ));
NOR2_X2 \GFM/U1713  ( .A1(\GFM/n24950 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1529 ));
NOR2_X2 \GFM/U1712  ( .A1(\GFM/n25040 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1526 ));
NOR2_X2 \GFM/U1711  ( .A1(\GFM/n24740 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1540 ));
NOR2_X2 \GFM/U1710  ( .A1(\GFM/n2424 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1544 ));
NOR2_X2 \GFM/U1709  ( .A1(\GFM/n24950 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1560 ));
NOR2_X2 \GFM/U1708  ( .A1(\GFM/n25040 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1557 ));
NOR2_X2 \GFM/U1707  ( .A1(\GFM/n24740 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1571 ));
NOR2_X2 \GFM/U1706  ( .A1(\GFM/n2424 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1575 ));
NOR2_X2 \GFM/U1705  ( .A1(\GFM/n24950 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1591 ));
NOR2_X2 \GFM/U1704  ( .A1(\GFM/n25040 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1588 ));
NOR2_X2 \GFM/U1703  ( .A1(\GFM/n24740 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1602 ));
NOR2_X2 \GFM/U1702  ( .A1(\GFM/n2424 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1606 ));
NOR2_X2 \GFM/U1701  ( .A1(\GFM/n25040 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1619 ));
NOR2_X2 \GFM/U1700  ( .A1(\GFM/n2494 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1622 ));
NOR2_X2 \GFM/U1699  ( .A1(\GFM/n24740 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1633 ));
NOR2_X2 \GFM/U1698  ( .A1(\GFM/n2424 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1637 ));
NOR2_X2 \GFM/U1697  ( .A1(\GFM/n25040 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1650 ));
NOR2_X2 \GFM/U1696  ( .A1(\GFM/n2494 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1653 ));
NOR2_X2 \GFM/U1695  ( .A1(\GFM/n24740 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1664 ));
NOR2_X2 \GFM/U1694  ( .A1(\GFM/n2424 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1668 ));
NOR2_X2 \GFM/U1693  ( .A1(\GFM/n25040 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1681 ));
NOR2_X2 \GFM/U1692  ( .A1(\GFM/n2494 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1684 ));
NOR2_X2 \GFM/U1691  ( .A1(\GFM/n24740 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1695 ));
NOR2_X2 \GFM/U1690  ( .A1(\GFM/n2424 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1699 ));
NOR2_X2 \GFM/U1689  ( .A1(\GFM/n2503 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1712 ));
NOR2_X2 \GFM/U1688  ( .A1(\GFM/n2494 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1715 ));
NOR2_X2 \GFM/U1687  ( .A1(\GFM/n24740 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1726 ));
NOR2_X2 \GFM/U1686  ( .A1(\GFM/n2424 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1730 ));
NOR2_X2 \GFM/U1685  ( .A1(\GFM/n2503 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1743 ));
NOR2_X2 \GFM/U1684  ( .A1(\GFM/n2494 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1746 ));
NOR2_X2 \GFM/U1683  ( .A1(\GFM/n24740 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1757 ));
NOR2_X2 \GFM/U1682  ( .A1(\GFM/n2424 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1761 ));
NOR2_X2 \GFM/U1681  ( .A1(\GFM/n2503 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1774 ));
NOR2_X2 \GFM/U1680  ( .A1(\GFM/n2494 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1777 ));
NOR2_X2 \GFM/U1679  ( .A1(\GFM/n24740 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1788 ));
NOR2_X2 \GFM/U1678  ( .A1(\GFM/n2424 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1792 ));
NOR2_X2 \GFM/U1677  ( .A1(\GFM/n2503 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1805 ));
NOR2_X2 \GFM/U1676  ( .A1(\GFM/n2494 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1808 ));
NOR2_X2 \GFM/U1675  ( .A1(\GFM/n24730 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1819 ));
NOR2_X2 \GFM/U1674  ( .A1(\GFM/n2423 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1823 ));
NOR2_X2 \GFM/U1673  ( .A1(\GFM/n2503 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1836 ));
NOR2_X2 \GFM/U1672  ( .A1(\GFM/n2494 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1839 ));
NOR2_X2 \GFM/U1671  ( .A1(\GFM/n24730 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1850 ));
NOR2_X2 \GFM/U1670  ( .A1(\GFM/n2423 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1854 ));
NOR2_X2 \GFM/U1669  ( .A1(\GFM/n2503 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1867 ));
NOR2_X2 \GFM/U1668  ( .A1(\GFM/n2494 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1870 ));
NOR2_X2 \GFM/U1667  ( .A1(\GFM/n24730 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1881 ));
NOR2_X2 \GFM/U1666  ( .A1(\GFM/n2423 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1885 ));
NOR2_X2 \GFM/U1665  ( .A1(\GFM/n2503 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1898 ));
NOR2_X2 \GFM/U1664  ( .A1(\GFM/n2494 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1901 ));
NOR2_X2 \GFM/U1663  ( .A1(\GFM/n24730 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1912 ));
NOR2_X2 \GFM/U1662  ( .A1(\GFM/n2423 ), .A2(\GFM/n2647 ), .ZN(\GFM/N1916 ));
NOR2_X2 \GFM/U1661  ( .A1(\GFM/n2503 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1929 ));
NOR2_X2 \GFM/U1660  ( .A1(\GFM/n2494 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1932 ));
NOR2_X2 \GFM/U1659  ( .A1(\GFM/n24730 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1943 ));
NOR2_X2 \GFM/U1658  ( .A1(\GFM/n2423 ), .A2(\GFM/n2648 ), .ZN(\GFM/N1947 ));
NOR2_X2 \GFM/U1657  ( .A1(\GFM/n2503 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1960 ));
NOR2_X2 \GFM/U1656  ( .A1(\GFM/n2493 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1963 ));
NOR2_X2 \GFM/U1655  ( .A1(\GFM/n24730 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1974 ));
NOR2_X2 \GFM/U1654  ( .A1(\GFM/n2423 ), .A2(\GFM/n2649 ), .ZN(\GFM/N1978 ));
NOR2_X2 \GFM/U1653  ( .A1(\GFM/n2503 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1991 ));
NOR2_X2 \GFM/U1652  ( .A1(\GFM/n2493 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1994 ));
NOR2_X2 \GFM/U1651  ( .A1(\GFM/n24730 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2005 ));
NOR2_X2 \GFM/U1650  ( .A1(\GFM/n2423 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2009 ));
NOR2_X2 \GFM/U1649  ( .A1(\GFM/n2503 ), .A2(\GFM/n26430 ), .ZN(\GFM/N2022 ));
NOR2_X2 \GFM/U1648  ( .A1(\GFM/n2493 ), .A2(\GFM/n2644 ), .ZN(\GFM/N2025 ));
NOR2_X2 \GFM/U1647  ( .A1(\GFM/n24730 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2036 ));
NOR2_X2 \GFM/U1646  ( .A1(\GFM/n2423 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2040 ));
NOR2_X2 \GFM/U1645  ( .A1(\GFM/n2503 ), .A2(\GFM/n2644 ), .ZN(\GFM/N2053 ));
NOR2_X2 \GFM/U1644  ( .A1(\GFM/n2493 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2056 ));
NOR2_X2 \GFM/U1643  ( .A1(\GFM/n24730 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2067 ));
NOR2_X2 \GFM/U1642  ( .A1(\GFM/n2423 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2071 ));
NOR2_X2 \GFM/U1641  ( .A1(\GFM/n2502 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2084 ));
NOR2_X2 \GFM/U1640  ( .A1(\GFM/n2493 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2087 ));
NOR2_X2 \GFM/U1639  ( .A1(\GFM/n24730 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2098 ));
NOR2_X2 \GFM/U1638  ( .A1(\GFM/n2423 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2102 ));
NOR2_X2 \GFM/U1637  ( .A1(\GFM/n2502 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2115 ));
NOR2_X2 \GFM/U1636  ( .A1(\GFM/n2493 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2118 ));
NOR2_X2 \GFM/U1635  ( .A1(\GFM/n24730 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2129 ));
NOR2_X2 \GFM/U1634  ( .A1(\GFM/n2423 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2133 ));
NOR2_X2 \GFM/U1633  ( .A1(\GFM/n2502 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2146 ));
NOR2_X2 \GFM/U1632  ( .A1(\GFM/n2493 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2149 ));
NOR2_X2 \GFM/U1631  ( .A1(\GFM/n2472 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2160 ));
NOR2_X2 \GFM/U1630  ( .A1(\GFM/n24220 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2164 ));
NOR2_X2 \GFM/U1629  ( .A1(\GFM/n2502 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2177 ));
NOR2_X2 \GFM/U1628  ( .A1(\GFM/n2493 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2180 ));
NOR2_X2 \GFM/U1627  ( .A1(\GFM/n2472 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2191 ));
NOR2_X2 \GFM/U1626  ( .A1(\GFM/n24220 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2195 ));
NOR2_X2 \GFM/U1625  ( .A1(\GFM/n2502 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2208 ));
NOR2_X2 \GFM/U1624  ( .A1(\GFM/n2493 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2211 ));
NOR2_X2 \GFM/U1623  ( .A1(\GFM/n2472 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2222 ));
NOR2_X2 \GFM/U1622  ( .A1(\GFM/n24220 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2226 ));
NOR2_X2 \GFM/U1621  ( .A1(\GFM/n2502 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2239 ));
NOR2_X2 \GFM/U1620  ( .A1(\GFM/n2493 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2242 ));
NOR2_X2 \GFM/U1619  ( .A1(\GFM/n2472 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2253 ));
NOR2_X2 \GFM/U1618  ( .A1(\GFM/n24220 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2257 ));
NOR2_X2 \GFM/U1617  ( .A1(\GFM/n2502 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2270 ));
NOR2_X2 \GFM/U1616  ( .A1(\GFM/n2493 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2273 ));
NOR2_X2 \GFM/U1615  ( .A1(\GFM/n2472 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2284 ));
NOR2_X2 \GFM/U1614  ( .A1(\GFM/n24220 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2288 ));
NOR2_X2 \GFM/U1613  ( .A1(\GFM/n2502 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2301 ));
NOR2_X2 \GFM/U1612  ( .A1(\GFM/n2493 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2304 ));
NOR2_X2 \GFM/U1611  ( .A1(\GFM/n2472 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2315 ));
NOR2_X2 \GFM/U1610  ( .A1(\GFM/n24220 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2319 ));
NOR2_X2 \GFM/U1609  ( .A1(\GFM/n2502 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2332 ));
NOR2_X2 \GFM/U1608  ( .A1(\GFM/n24921 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2335 ));
NOR2_X2 \GFM/U1607  ( .A1(\GFM/n2472 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2346 ));
NOR2_X2 \GFM/U1606  ( .A1(\GFM/n24220 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2350 ));
NOR2_X2 \GFM/U1605  ( .A1(\GFM/n2502 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2363 ));
NOR2_X2 \GFM/U1604  ( .A1(\GFM/n24921 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2366 ));
NOR2_X2 \GFM/U1603  ( .A1(\GFM/n2472 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2377 ));
NOR2_X2 \GFM/U1602  ( .A1(\GFM/n24220 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2381 ));
NOR2_X2 \GFM/U1601  ( .A1(\GFM/n2502 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2394 ));
NOR2_X2 \GFM/U1600  ( .A1(\GFM/n24921 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2397 ));
NOR2_X2 \GFM/U1599  ( .A1(\GFM/n2472 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2408 ));
NOR2_X2 \GFM/U1598  ( .A1(\GFM/n24220 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2412 ));
NOR2_X2 \GFM/U1597  ( .A1(\GFM/n2502 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2425 ));
NOR2_X2 \GFM/U1596  ( .A1(\GFM/n24921 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2428 ));
NOR2_X2 \GFM/U1595  ( .A1(\GFM/n2472 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2439 ));
NOR2_X2 \GFM/U1594  ( .A1(\GFM/n24220 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2443 ));
NOR2_X2 \GFM/U1593  ( .A1(\GFM/n25010 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2456 ));
NOR2_X2 \GFM/U1592  ( .A1(\GFM/n24921 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2459 ));
NOR2_X2 \GFM/U1591  ( .A1(\GFM/n2472 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2470 ));
NOR2_X2 \GFM/U1590  ( .A1(\GFM/n24220 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2474 ));
NOR2_X2 \GFM/U1589  ( .A1(\GFM/n25010 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2487 ));
NOR2_X2 \GFM/U1588  ( .A1(\GFM/n24921 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2490 ));
NOR2_X2 \GFM/U1587  ( .A1(\GFM/n2472 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2501 ));
NOR2_X2 \GFM/U1586  ( .A1(\GFM/n24210 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2505 ));
NOR2_X2 \GFM/U1585  ( .A1(\GFM/n25010 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2518 ));
NOR2_X2 \GFM/U1584  ( .A1(\GFM/n24921 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2521 ));
NOR2_X2 \GFM/U1583  ( .A1(\GFM/n2472 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2532 ));
NOR2_X2 \GFM/U1582  ( .A1(\GFM/n24210 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2536 ));
NOR2_X2 \GFM/U1581  ( .A1(\GFM/n25010 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2549 ));
NOR2_X2 \GFM/U1580  ( .A1(\GFM/n24921 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2552 ));
NOR2_X2 \GFM/U1579  ( .A1(\GFM/n2471 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2563 ));
NOR2_X2 \GFM/U1578  ( .A1(\GFM/n24210 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2567 ));
NOR2_X2 \GFM/U1577  ( .A1(\GFM/n25010 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2580 ));
NOR2_X2 \GFM/U1576  ( .A1(\GFM/n24921 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2583 ));
NOR2_X2 \GFM/U1575  ( .A1(\GFM/n2471 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2594 ));
NOR2_X2 \GFM/U1574  ( .A1(\GFM/n24210 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2598 ));
NOR2_X2 \GFM/U1573  ( .A1(\GFM/n25010 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2611 ));
NOR2_X2 \GFM/U1572  ( .A1(\GFM/n24921 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2614 ));
NOR2_X2 \GFM/U1571  ( .A1(\GFM/n2471 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2625 ));
NOR2_X2 \GFM/U1570  ( .A1(\GFM/n24210 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2629 ));
NOR2_X2 \GFM/U1569  ( .A1(\GFM/n25010 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2642 ));
NOR2_X2 \GFM/U1568  ( .A1(\GFM/n24921 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2645 ));
NOR2_X2 \GFM/U1567  ( .A1(\GFM/n2471 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2656 ));
NOR2_X2 \GFM/U1566  ( .A1(\GFM/n24210 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2660 ));
NOR2_X2 \GFM/U1565  ( .A1(\GFM/n25010 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2673 ));
NOR2_X2 \GFM/U1564  ( .A1(\GFM/n24921 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2676 ));
NOR2_X2 \GFM/U1563  ( .A1(\GFM/n2471 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2687 ));
NOR2_X2 \GFM/U1562  ( .A1(\GFM/n25010 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2704 ));
NOR2_X2 \GFM/U1561  ( .A1(\GFM/n24910 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2707 ));
NOR2_X2 \GFM/U1560  ( .A1(\GFM/n2471 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2718 ));
NOR2_X2 \GFM/U1559  ( .A1(\GFM/n25010 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2735 ));
NOR2_X2 \GFM/U1558  ( .A1(\GFM/n24910 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2738 ));
NOR2_X2 \GFM/U1557  ( .A1(\GFM/n2471 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2749 ));
NOR2_X2 \GFM/U1556  ( .A1(\GFM/n25010 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2766 ));
NOR2_X2 \GFM/U1555  ( .A1(\GFM/n24910 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2769 ));
NOR2_X2 \GFM/U1554  ( .A1(\GFM/n2471 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2780 ));
NOR2_X2 \GFM/U1553  ( .A1(\GFM/n25010 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2797 ));
NOR2_X2 \GFM/U1552  ( .A1(\GFM/n24910 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2800 ));
NOR2_X2 \GFM/U1551  ( .A1(\GFM/n2471 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2811 ));
NOR2_X2 \GFM/U1550  ( .A1(\GFM/n25000 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2828 ));
NOR2_X2 \GFM/U1549  ( .A1(\GFM/n24910 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2831 ));
NOR2_X2 \GFM/U1548  ( .A1(\GFM/n25000 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2859 ));
NOR2_X2 \GFM/U1547  ( .A1(\GFM/n24910 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2862 ));
NOR2_X2 \GFM/U1546  ( .A1(\GFM/n25000 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2890 ));
NOR2_X2 \GFM/U1545  ( .A1(\GFM/n24210 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2691 ));
NOR2_X2 \GFM/U1544  ( .A1(\GFM/n24210 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2722 ));
NOR2_X2 \GFM/U1543  ( .A1(\GFM/n24210 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2753 ));
NOR2_X2 \GFM/U1542  ( .A1(\GFM/n24210 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2784 ));
NOR2_X2 \GFM/U1541  ( .A1(\GFM/n24210 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2815 ));
NOR2_X2 \GFM/U1540  ( .A1(\GFM/n2471 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2842 ));
NOR2_X2 \GFM/U1539  ( .A1(\GFM/n24201 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2846 ));
NOR2_X2 \GFM/U1538  ( .A1(\GFM/n2471 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2873 ));
NOR2_X2 \GFM/U1537  ( .A1(\GFM/n24201 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2877 ));
NOR2_X2 \GFM/U1536  ( .A1(\GFM/n24910 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2893 ));
NOR2_X2 \GFM/U1535  ( .A1(\GFM/n2471 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2904 ));
NOR2_X2 \GFM/U1534  ( .A1(\GFM/n24201 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2908 ));
NOR2_X2 \GFM/U1533  ( .A1(\GFM/n25000 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2921 ));
NOR2_X2 \GFM/U1532  ( .A1(\GFM/n24910 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2924 ));
NOR2_X2 \GFM/U1531  ( .A1(\GFM/n24700 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2935 ));
NOR2_X2 \GFM/U1530  ( .A1(\GFM/n24201 ), .A2(\GFM/n26801 ), .ZN(\GFM/N2939 ));
NOR2_X2 \GFM/U1529  ( .A1(\GFM/n25000 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2952 ));
NOR2_X2 \GFM/U1528  ( .A1(\GFM/n24910 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2955 ));
NOR2_X2 \GFM/U1527  ( .A1(\GFM/n24700 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2966 ));
NOR2_X2 \GFM/U1526  ( .A1(\GFM/n24201 ), .A2(\GFM/n26810 ), .ZN(\GFM/N2970 ));
NOR2_X2 \GFM/U1525  ( .A1(\GFM/n25000 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2983 ));
NOR2_X2 \GFM/U1524  ( .A1(\GFM/n24910 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2986 ));
NOR2_X2 \GFM/U1523  ( .A1(\GFM/n24700 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2997 ));
NOR2_X2 \GFM/U1522  ( .A1(\GFM/n24201 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3001 ));
NOR2_X2 \GFM/U1521  ( .A1(\GFM/n25000 ), .A2(\GFM/n2675 ), .ZN(\GFM/N3014 ));
NOR2_X2 \GFM/U1520  ( .A1(\GFM/n24910 ), .A2(\GFM/n26760 ), .ZN(\GFM/N3017 ));
NOR2_X2 \GFM/U1519  ( .A1(\GFM/n24700 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3028 ));
NOR2_X2 \GFM/U1518  ( .A1(\GFM/n24201 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3032 ));
NOR2_X2 \GFM/U1517  ( .A1(\GFM/n25000 ), .A2(\GFM/n26760 ), .ZN(\GFM/N3045 ));
NOR2_X2 \GFM/U1516  ( .A1(\GFM/n24900 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3048 ));
NOR2_X2 \GFM/U1515  ( .A1(\GFM/n24700 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3059 ));
NOR2_X2 \GFM/U1514  ( .A1(\GFM/n24201 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3063 ));
NOR2_X2 \GFM/U1513  ( .A1(\GFM/n25000 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3076 ));
NOR2_X2 \GFM/U1512  ( .A1(\GFM/n24900 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3079 ));
NOR2_X2 \GFM/U1511  ( .A1(\GFM/n24700 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3090 ));
NOR2_X2 \GFM/U1510  ( .A1(\GFM/n24201 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3094 ));
NOR2_X2 \GFM/U1509  ( .A1(\GFM/n25000 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3107 ));
NOR2_X2 \GFM/U1508  ( .A1(\GFM/n24900 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3110 ));
NOR2_X2 \GFM/U1507  ( .A1(\GFM/n24700 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3121 ));
NOR2_X2 \GFM/U1506  ( .A1(\GFM/n24201 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3125 ));
NOR2_X2 \GFM/U1505  ( .A1(\GFM/n25000 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3138 ));
NOR2_X2 \GFM/U1504  ( .A1(\GFM/n24900 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3141 ));
NOR2_X2 \GFM/U1503  ( .A1(\GFM/n24700 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3152 ));
NOR2_X2 \GFM/U1502  ( .A1(\GFM/n24201 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3156 ));
NOR2_X2 \GFM/U1501  ( .A1(\GFM/n2499 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3169 ));
NOR2_X2 \GFM/U1500  ( .A1(\GFM/n24900 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3172 ));
NOR2_X2 \GFM/U1499  ( .A1(\GFM/n24700 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3183 ));
NOR2_X2 \GFM/U1498  ( .A1(\GFM/n24201 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3187 ));
NOR2_X2 \GFM/U1497  ( .A1(\GFM/n2499 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3200 ));
NOR2_X2 \GFM/U1496  ( .A1(\GFM/n24900 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3203 ));
NOR2_X2 \GFM/U1495  ( .A1(\GFM/n24700 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3214 ));
NOR2_X2 \GFM/U1494  ( .A1(\GFM/n24190 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3218 ));
NOR2_X2 \GFM/U1493  ( .A1(\GFM/n2499 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3231 ));
NOR2_X2 \GFM/U1492  ( .A1(\GFM/n24910 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3234 ));
NOR2_X2 \GFM/U1491  ( .A1(\GFM/n24700 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3245 ));
NOR2_X2 \GFM/U1490  ( .A1(\GFM/n24190 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3249 ));
NOR2_X2 \GFM/U1489  ( .A1(\GFM/n2499 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3262 ));
NOR2_X2 \GFM/U1488  ( .A1(\GFM/n24900 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3265 ));
NOR2_X2 \GFM/U1487  ( .A1(\GFM/n24700 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3276 ));
NOR2_X2 \GFM/U1486  ( .A1(\GFM/n24190 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3280 ));
NOR2_X2 \GFM/U1485  ( .A1(\GFM/n2499 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3293 ));
NOR2_X2 \GFM/U1484  ( .A1(\GFM/n25101 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3296 ));
NOR2_X2 \GFM/U1483  ( .A1(\GFM/n24500 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3308 ));
NOR2_X2 \GFM/U1482  ( .A1(\GFM/n2400 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3312 ));
NOR2_X2 \GFM/U1481  ( .A1(\GFM/n2499 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3325 ));
NOR2_X2 \GFM/U1480  ( .A1(\GFM/n25101 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3328 ));
NOR2_X2 \GFM/U1479  ( .A1(\GFM/n2449 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3340 ));
NOR2_X2 \GFM/U1478  ( .A1(\GFM/n2499 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3358 ));
NOR2_X2 \GFM/U1477  ( .A1(\GFM/n25101 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3361 ));
NOR2_X2 \GFM/U1476  ( .A1(\GFM/n2449 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3373 ));
NOR2_X2 \GFM/U1475  ( .A1(\GFM/n2499 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3392 ));
NOR2_X2 \GFM/U1474  ( .A1(\GFM/n25101 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3395 ));
NOR2_X2 \GFM/U1473  ( .A1(\GFM/n24690 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3398 ));
NOR2_X2 \GFM/U1472  ( .A1(\GFM/n2499 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3428 ));
NOR2_X2 \GFM/U1471  ( .A1(\GFM/n25101 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3431 ));
NOR2_X2 \GFM/U1470  ( .A1(\GFM/n24690 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3434 ));
NOR2_X2 \GFM/U1469  ( .A1(\GFM/n24690 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3472 ));
NOR2_X2 \GFM/U1468  ( .A1(\GFM/n2449 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3483 ));
NOR2_X2 \GFM/U1467  ( .A1(\GFM/n24690 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3513 ));
NOR2_X2 \GFM/U1466  ( .A1(\GFM/n24690 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3556 ));
NOR2_X2 \GFM/U1465  ( .A1(\GFM/n2509 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3750 ));
NOR2_X2 \GFM/U1464  ( .A1(\GFM/n2610 ), .A2(\GFM/n24070 ), .ZN(\GFM/N737 ));
NOR2_X2 \GFM/U1463  ( .A1(\GFM/n2610 ), .A2(\GFM/n2516 ), .ZN(\GFM/N1058 ));
NOR2_X2 \GFM/U1462  ( .A1(\GFM/n26080 ), .A2(\GFM/n2506 ), .ZN(\GFM/N969 ));
NOR2_X2 \GFM/U1461  ( .A1(\GFM/n26070 ), .A2(\GFM/n24760 ), .ZN(\GFM/N848 ));
NOR2_X2 \GFM/U1460  ( .A1(\GFM/n26070 ), .A2(\GFM/n2506 ), .ZN(\GFM/N938 ));
NOR2_X2 \GFM/U1459  ( .A1(\GFM/n2606 ), .A2(\GFM/n24070 ), .ZN(\GFM/N613 ));
NOR2_X2 \GFM/U1458  ( .A1(\GFM/n2606 ), .A2(\GFM/n24560 ), .ZN(\GFM/N764 ));
NOR2_X2 \GFM/U1457  ( .A1(\GFM/n26200 ), .A2(\GFM/n24460 ), .ZN(\GFM/N1163 ));
NOR2_X2 \GFM/U1456  ( .A1(\GFM/n26190 ), .A2(\GFM/n24070 ), .ZN(\GFM/N1016 ));
NOR2_X2 \GFM/U1455  ( .A1(\GFM/n26190 ), .A2(\GFM/n24460 ), .ZN(\GFM/N1132 ));
NOR2_X2 \GFM/U1454  ( .A1(\GFM/n26190 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1310 ));
NOR2_X2 \GFM/U1453  ( .A1(\GFM/n2617 ), .A2(\GFM/n24070 ), .ZN(\GFM/N954 ));
NOR2_X2 \GFM/U1452  ( .A1(\GFM/n26120 ), .A2(\GFM/n24460 ), .ZN(\GFM/N915 ));
NOR2_X2 \GFM/U1451  ( .A1(\GFM/n2517 ), .A2(\GFM/n25700 ), .ZN(\GFM/N97 ) );
NOR2_X2 \GFM/U1450  ( .A1(\GFM/n25150 ), .A2(\GFM/n25760 ), .ZN(\GFM/N132 ));
NOR2_X2 \GFM/U1449  ( .A1(\GFM/n25150 ), .A2(\GFM/n2578 ), .ZN(\GFM/N163 ));
NOR2_X2 \GFM/U1448  ( .A1(\GFM/n2610 ), .A2(\GFM/n24870 ), .ZN(\GFM/N971 ));
NOR2_X2 \GFM/U1447  ( .A1(\GFM/n26080 ), .A2(\GFM/n2427 ), .ZN(\GFM/N731 ));
NOR2_X2 \GFM/U1446  ( .A1(\GFM/n2606 ), .A2(\GFM/n24460 ), .ZN(\GFM/N729 ));
NOR2_X2 \GFM/U1445  ( .A1(\GFM/n26080 ), .A2(\GFM/n2387 ), .ZN(\GFM/N617 ));
NOR2_X2 \GFM/U1444  ( .A1(\GFM/n26070 ), .A2(\GFM/n2437 ), .ZN(\GFM/N728 ));
NOR2_X2 \GFM/U1443  ( .A1(\GFM/n24770 ), .A2(\GFM/n2603 ), .ZN(\GFM/N724 ));
NOR2_X2 \GFM/U1442  ( .A1(\GFM/n26070 ), .A2(\GFM/n2387 ), .ZN(\GFM/N586 ));
NOR2_X2 \GFM/U1441  ( .A1(\GFM/n26070 ), .A2(\GFM/n25530 ), .ZN(\GFM/N676 ));
NOR2_X2 \GFM/U1440  ( .A1(\GFM/n26070 ), .A2(\GFM/n2466 ), .ZN(\GFM/N827 ));
NOR2_X2 \GFM/U1439  ( .A1(\GFM/n26070 ), .A2(\GFM/n24870 ), .ZN(\GFM/N878 ));
NOR2_X2 \GFM/U1438  ( .A1(\GFM/n2606 ), .A2(\GFM/n2427 ), .ZN(\GFM/N669 ) );
NOR2_X2 \GFM/U1437  ( .A1(\GFM/n2448 ), .A2(\GFM/n2604 ), .ZN(\GFM/N667 ) );
NOR2_X2 \GFM/U1436  ( .A1(\GFM/n2606 ), .A2(\GFM/n25530 ), .ZN(\GFM/N645 ));
NOR2_X2 \GFM/U1435  ( .A1(\GFM/n2606 ), .A2(\GFM/n2466 ), .ZN(\GFM/N796 ) );
NOR2_X2 \GFM/U1434  ( .A1(\GFM/n26200 ), .A2(\GFM/n24360 ), .ZN(\GFM/N1131 ));
NOR2_X2 \GFM/U1433  ( .A1(\GFM/n26190 ), .A2(\GFM/n24260 ), .ZN(\GFM/N1072 ));
NOR2_X2 \GFM/U1432  ( .A1(\GFM/n2617 ), .A2(\GFM/n24460 ), .ZN(\GFM/N1070 ));
NOR2_X2 \GFM/U1431  ( .A1(\GFM/n26190 ), .A2(\GFM/n24360 ), .ZN(\GFM/N1100 ));
NOR2_X2 \GFM/U1430  ( .A1(\GFM/n26150 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1096 ));
NOR2_X2 \GFM/U1429  ( .A1(\GFM/n26190 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1250 ));
NOR2_X2 \GFM/U1428  ( .A1(\GFM/n2617 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1248 ));
NOR2_X2 \GFM/U1427  ( .A1(\GFM/n26190 ), .A2(\GFM/n25530 ), .ZN(\GFM/N1048 ));
NOR2_X2 \GFM/U1426  ( .A1(\GFM/n26190 ), .A2(\GFM/n2466 ), .ZN(\GFM/N1199 ));
NOR2_X2 \GFM/U1425  ( .A1(\GFM/n2617 ), .A2(\GFM/n2466 ), .ZN(\GFM/N1137 ));
NOR2_X2 \GFM/U1424  ( .A1(\GFM/n2618 ), .A2(\GFM/n2466 ), .ZN(\GFM/N1168 ));
NOR2_X2 \GFM/U1423  ( .A1(\GFM/n26120 ), .A2(\GFM/n24260 ), .ZN(\GFM/N855 ));
NOR2_X2 \GFM/U1422  ( .A1(\GFM/n26120 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1033 ));
NOR2_X2 \GFM/U1421  ( .A1(\GFM/n2613 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1064 ));
NOR2_X2 \GFM/U1420  ( .A1(\GFM/n26140 ), .A2(\GFM/n24360 ), .ZN(\GFM/N945 ));
NOR2_X2 \GFM/U1419  ( .A1(\GFM/n2610 ), .A2(\GFM/n24760 ), .ZN(\GFM/N941 ));
NOR2_X2 \GFM/U1418  ( .A1(\GFM/n26140 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1095 ));
NOR2_X2 \GFM/U1417  ( .A1(\GFM/n26150 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1126 ));
NOR2_X2 \GFM/U1416  ( .A1(\GFM/n2613 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1124 ));
NOR2_X2 \GFM/U1415  ( .A1(\GFM/n25140 ), .A2(\GFM/n25800 ), .ZN(\GFM/N194 ));
NOR2_X2 \GFM/U1414  ( .A1(\GFM/n24880 ), .A2(\GFM/n25700 ), .ZN(\GFM/N10 ));
NOR2_X2 \GFM/U1413  ( .A1(\GFM/n24980 ), .A2(\GFM/n25700 ), .ZN(\GFM/N38 ));
NOR2_X2 \GFM/U1412  ( .A1(\GFM/n24570 ), .A2(\GFM/n25821 ), .ZN(\GFM/N82 ));
NOR2_X2 \GFM/U1411  ( .A1(\GFM/n2513 ), .A2(\GFM/n25821 ), .ZN(\GFM/N225 ));
NOR2_X2 \GFM/U1410  ( .A1(\GFM/n2489 ), .A2(\GFM/n2573 ), .ZN(\GFM/N41 ) );
NOR2_X2 \GFM/U1409  ( .A1(\GFM/n2497 ), .A2(\GFM/n2573 ), .ZN(\GFM/N69 ) );
NOR2_X2 \GFM/U1408  ( .A1(\GFM/n24730 ), .A2(\GFM/n25760 ), .ZN(\GFM/N21 ));
NOR2_X2 \GFM/U1407  ( .A1(\GFM/n24880 ), .A2(\GFM/n25760 ), .ZN(\GFM/N72 ));
NOR2_X2 \GFM/U1406  ( .A1(\GFM/n2497 ), .A2(\GFM/n25760 ), .ZN(\GFM/N100 ));
NOR2_X2 \GFM/U1405  ( .A1(\GFM/n24650 ), .A2(\GFM/n25840 ), .ZN(\GFM/N113 ));
NOR2_X2 \GFM/U1404  ( .A1(\GFM/n25120 ), .A2(\GFM/n25840 ), .ZN(\GFM/N256 ));
NOR2_X2 \GFM/U1403  ( .A1(\GFM/n2468 ), .A2(\GFM/n2578 ), .ZN(\GFM/N52 ) );
NOR2_X2 \GFM/U1402  ( .A1(\GFM/n24950 ), .A2(\GFM/n2578 ), .ZN(\GFM/N103 ));
NOR2_X2 \GFM/U1401  ( .A1(\GFM/n25050 ), .A2(\GFM/n2578 ), .ZN(\GFM/N131 ));
NOR2_X2 \GFM/U1400  ( .A1(\GFM/n24650 ), .A2(\GFM/n2586 ), .ZN(\GFM/N144 ));
NOR2_X2 \GFM/U1399  ( .A1(\GFM/n2511 ), .A2(\GFM/n2586 ), .ZN(\GFM/N287 ) );
NOR2_X2 \GFM/U1398  ( .A1(\GFM/n25201 ), .A2(\GFM/n2586 ), .ZN(\GFM/N314 ));
NOR2_X2 \GFM/U1397  ( .A1(\GFM/n24670 ), .A2(\GFM/n25800 ), .ZN(\GFM/N83 ));
NOR2_X2 \GFM/U1396  ( .A1(\GFM/n24950 ), .A2(\GFM/n25800 ), .ZN(\GFM/N134 ));
NOR2_X2 \GFM/U1395  ( .A1(\GFM/n25040 ), .A2(\GFM/n25800 ), .ZN(\GFM/N162 ));
NOR2_X2 \GFM/U1394  ( .A1(\GFM/n2475 ), .A2(\GFM/n25821 ), .ZN(\GFM/N114 ));
NOR2_X2 \GFM/U1393  ( .A1(\GFM/n2494 ), .A2(\GFM/n25821 ), .ZN(\GFM/N165 ));
NOR2_X2 \GFM/U1392  ( .A1(\GFM/n2503 ), .A2(\GFM/n25821 ), .ZN(\GFM/N193 ));
NOR2_X2 \GFM/U1391  ( .A1(\GFM/n2413 ), .A2(\GFM/n2587 ), .ZN(\GFM/N24 ) );
NOR2_X2 \GFM/U1390  ( .A1(\GFM/n24640 ), .A2(\GFM/n2587 ), .ZN(\GFM/N175 ));
NOR2_X2 \GFM/U1389  ( .A1(\GFM/n25101 ), .A2(\GFM/n2587 ), .ZN(\GFM/N318 ));
NOR2_X2 \GFM/U1388  ( .A1(\GFM/n25190 ), .A2(\GFM/n2587 ), .ZN(\GFM/N345 ));
NOR2_X2 \GFM/U1387  ( .A1(\GFM/n24340 ), .A2(\GFM/n25840 ), .ZN(\GFM/N18 ));
NOR2_X2 \GFM/U1386  ( .A1(\GFM/n2454 ), .A2(\GFM/n25800 ), .ZN(\GFM/N16 ) );
NOR2_X2 \GFM/U1385  ( .A1(\GFM/n24740 ), .A2(\GFM/n25840 ), .ZN(\GFM/N145 ));
NOR2_X2 \GFM/U1384  ( .A1(\GFM/n2494 ), .A2(\GFM/n25840 ), .ZN(\GFM/N196 ));
NOR2_X2 \GFM/U1383  ( .A1(\GFM/n2502 ), .A2(\GFM/n25840 ), .ZN(\GFM/N224 ));
NOR2_X2 \GFM/U1382  ( .A1(\GFM/n24380 ), .A2(\GFM/n2586 ), .ZN(\GFM/N77 ) );
NOR2_X2 \GFM/U1381  ( .A1(\GFM/n2478 ), .A2(\GFM/n2578 ), .ZN(\GFM/N73 ) );
NOR2_X2 \GFM/U1380  ( .A1(\GFM/n24220 ), .A2(\GFM/n2586 ), .ZN(\GFM/N25 ) );
NOR2_X2 \GFM/U1379  ( .A1(\GFM/n24740 ), .A2(\GFM/n2586 ), .ZN(\GFM/N176 ));
NOR2_X2 \GFM/U1378  ( .A1(\GFM/n2493 ), .A2(\GFM/n2586 ), .ZN(\GFM/N227 ) );
NOR2_X2 \GFM/U1377  ( .A1(\GFM/n25010 ), .A2(\GFM/n2586 ), .ZN(\GFM/N255 ));
NOR2_X2 \GFM/U1376  ( .A1(\GFM/n2427 ), .A2(\GFM/n2587 ), .ZN(\GFM/N80 ) );
NOR2_X2 \GFM/U1375  ( .A1(\GFM/n2448 ), .A2(\GFM/n25840 ), .ZN(\GFM/N78 ) );
NOR2_X2 \GFM/U1374  ( .A1(\GFM/n2418 ), .A2(\GFM/n2587 ), .ZN(\GFM/N56 ) );
NOR2_X2 \GFM/U1373  ( .A1(\GFM/n24730 ), .A2(\GFM/n2587 ), .ZN(\GFM/N207 ));
NOR2_X2 \GFM/U1372  ( .A1(\GFM/n24921 ), .A2(\GFM/n2587 ), .ZN(\GFM/N258 ));
NOR2_X2 \GFM/U1371  ( .A1(\GFM/n25000 ), .A2(\GFM/n2587 ), .ZN(\GFM/N286 ));
NOR2_X2 \GFM/U1370  ( .A1(\GFM/n25890 ), .A2(\GFM/n24570 ), .ZN(\GFM/N237 ));
NOR2_X2 \GFM/U1369  ( .A1(\GFM/n25890 ), .A2(\GFM/n25070 ), .ZN(\GFM/N380 ));
NOR2_X2 \GFM/U1368  ( .A1(\GFM/n25700 ), .A2(\GFM/n25070 ), .ZN(\GFM/N70 ));
NOR2_X2 \GFM/U1367  ( .A1(\GFM/n25890 ), .A2(\GFM/n24870 ), .ZN(\GFM/N320 ));
NOR2_X2 \GFM/U1366  ( .A1(\GFM/n25880 ), .A2(\GFM/n23980 ), .ZN(\GFM/N27 ));
NOR2_X2 \GFM/U1365  ( .A1(\GFM/n25880 ), .A2(\GFM/n24070 ), .ZN(\GFM/N55 ));
NOR2_X2 \GFM/U1364  ( .A1(\GFM/n25880 ), .A2(\GFM/n24570 ), .ZN(\GFM/N206 ));
NOR2_X2 \GFM/U1363  ( .A1(\GFM/n25880 ), .A2(\GFM/n25070 ), .ZN(\GFM/N349 ));
NOR2_X2 \GFM/U1362  ( .A1(\GFM/n25880 ), .A2(\GFM/n25530 ), .ZN(\GFM/N87 ));
NOR2_X2 \GFM/U1361  ( .A1(\GFM/n25880 ), .A2(\GFM/n24670 ), .ZN(\GFM/N238 ));
NOR2_X2 \GFM/U1360  ( .A1(\GFM/n25880 ), .A2(\GFM/n24870 ), .ZN(\GFM/N289 ));
NOR2_X2 \GFM/U1359  ( .A1(\GFM/n25620 ), .A2(\GFM/n25070 ), .ZN(\GFM/N8 ) );
NOR2_X2 \GFM/U1358  ( .A1(\GFM/n25660 ), .A2(\GFM/n25070 ), .ZN(\GFM/N39 ));
NOR2_X2 \GFM/U1357  ( .A1(\GFM/n25660 ), .A2(\GFM/n24960 ), .ZN(\GFM/N7 ) );
NOR2_X2 \GFM/U1356  ( .A1(\GFM/n25700 ), .A2(\GFM/n24760 ), .ZN(\GFM/N4332 ));
NOR2_X2 \GFM/U1355  ( .A1(\GFM/n25580 ), .A2(\GFM/n2516 ), .ZN(\GFM/N4 ) );
NOR2_X2 \GFM/U1354  ( .A1(\GFM/n25620 ), .A2(\GFM/n2516 ), .ZN(\GFM/N35 ) );
NOR2_X2 \GFM/U1353  ( .A1(\GFM/n26070 ), .A2(\GFM/n24070 ), .ZN(\GFM/N644 ));
NOR2_X2 \GFM/U1352  ( .A1(\GFM/n26080 ), .A2(\GFM/n24070 ), .ZN(\GFM/N675 ));
NOR2_X2 \GFM/U1351  ( .A1(\GFM/n26080 ), .A2(\GFM/n24250 ), .ZN(\GFM/N707 ));
NOR2_X2 \GFM/U1350  ( .A1(\GFM/n25080 ), .A2(\GFM/n26010 ), .ZN(\GFM/N752 ));
NOR2_X2 \GFM/U1349  ( .A1(\GFM/n2610 ), .A2(\GFM/n24250 ), .ZN(\GFM/N769 ));
NOR2_X2 \GFM/U1348  ( .A1(\GFM/n25080 ), .A2(\GFM/n2603 ), .ZN(\GFM/N814 ));
NOR2_X2 \GFM/U1347  ( .A1(\GFM/n2610 ), .A2(\GFM/n24460 ), .ZN(\GFM/N853 ));
NOR2_X2 \GFM/U1346  ( .A1(\GFM/n26110 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1002 ));
NOR2_X2 \GFM/U1345  ( .A1(\GFM/n2610 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1031 ));
NOR2_X2 \GFM/U1344  ( .A1(\GFM/n26200 ), .A2(\GFM/n24070 ), .ZN(\GFM/N1047 ));
NOR2_X2 \GFM/U1343  ( .A1(\GFM/n26110 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1062 ));
NOR2_X2 \GFM/U1342  ( .A1(\GFM/n26200 ), .A2(\GFM/n25530 ), .ZN(\GFM/N1079 ));
NOR2_X2 \GFM/U1341  ( .A1(\GFM/n26120 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1093 ));
NOR2_X2 \GFM/U1340  ( .A1(\GFM/n26200 ), .A2(\GFM/n25070 ), .ZN(\GFM/N1341 ));
NOR2_X2 \GFM/U1339  ( .A1(\GFM/n25150 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1372 ));
NOR2_X2 \GFM/U1338  ( .A1(\GFM/n25150 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1403 ));
NOR2_X2 \GFM/U1337  ( .A1(\GFM/n25150 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1434 ));
NOR2_X2 \GFM/U1336  ( .A1(\GFM/n25150 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1465 ));
NOR2_X2 \GFM/U1335  ( .A1(\GFM/n25150 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1496 ));
NOR2_X2 \GFM/U1334  ( .A1(\GFM/n25150 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1527 ));
NOR2_X2 \GFM/U1333  ( .A1(\GFM/n25150 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1558 ));
NOR2_X2 \GFM/U1332  ( .A1(\GFM/n25150 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1589 ));
NOR2_X2 \GFM/U1331  ( .A1(\GFM/n24401 ), .A2(\GFM/n25940 ), .ZN(\GFM/N325 ));
NOR2_X2 \GFM/U1330  ( .A1(\GFM/n2480 ), .A2(\GFM/n25901 ), .ZN(\GFM/N321 ));
NOR2_X2 \GFM/U1329  ( .A1(\GFM/n24390 ), .A2(\GFM/n2595 ), .ZN(\GFM/N356 ));
NOR2_X2 \GFM/U1328  ( .A1(\GFM/n2479 ), .A2(\GFM/n25910 ), .ZN(\GFM/N352 ));
NOR2_X2 \GFM/U1327  ( .A1(\GFM/n24390 ), .A2(\GFM/n2596 ), .ZN(\GFM/N387 ));
NOR2_X2 \GFM/U1326  ( .A1(\GFM/n2479 ), .A2(\GFM/n2592 ), .ZN(\GFM/N383 ) );
NOR2_X2 \GFM/U1325  ( .A1(\GFM/n24390 ), .A2(\GFM/n25970 ), .ZN(\GFM/N418 ));
NOR2_X2 \GFM/U1324  ( .A1(\GFM/n2479 ), .A2(\GFM/n25930 ), .ZN(\GFM/N414 ));
NOR2_X2 \GFM/U1323  ( .A1(\GFM/n24380 ), .A2(\GFM/n25980 ), .ZN(\GFM/N449 ));
NOR2_X2 \GFM/U1322  ( .A1(\GFM/n2479 ), .A2(\GFM/n25940 ), .ZN(\GFM/N445 ));
NOR2_X2 \GFM/U1321  ( .A1(\GFM/n24380 ), .A2(\GFM/n2599 ), .ZN(\GFM/N480 ));
NOR2_X2 \GFM/U1320  ( .A1(\GFM/n2478 ), .A2(\GFM/n2595 ), .ZN(\GFM/N476 ) );
NOR2_X2 \GFM/U1319  ( .A1(\GFM/n24380 ), .A2(\GFM/n26000 ), .ZN(\GFM/N511 ));
NOR2_X2 \GFM/U1318  ( .A1(\GFM/n2478 ), .A2(\GFM/n2596 ), .ZN(\GFM/N507 ) );
NOR2_X2 \GFM/U1317  ( .A1(\GFM/n24380 ), .A2(\GFM/n26010 ), .ZN(\GFM/N542 ));
NOR2_X2 \GFM/U1316  ( .A1(\GFM/n2478 ), .A2(\GFM/n25970 ), .ZN(\GFM/N538 ));
NOR2_X2 \GFM/U1315  ( .A1(\GFM/n24380 ), .A2(\GFM/n2602 ), .ZN(\GFM/N573 ));
NOR2_X2 \GFM/U1314  ( .A1(\GFM/n2478 ), .A2(\GFM/n25980 ), .ZN(\GFM/N569 ));
NOR2_X2 \GFM/U1313  ( .A1(\GFM/n2437 ), .A2(\GFM/n2603 ), .ZN(\GFM/N604 ) );
NOR2_X2 \GFM/U1312  ( .A1(\GFM/n2478 ), .A2(\GFM/n2599 ), .ZN(\GFM/N600 ) );
NOR2_X2 \GFM/U1311  ( .A1(\GFM/n24380 ), .A2(\GFM/n2604 ), .ZN(\GFM/N635 ));
NOR2_X2 \GFM/U1310  ( .A1(\GFM/n2478 ), .A2(\GFM/n26000 ), .ZN(\GFM/N631 ));
NOR2_X2 \GFM/U1309  ( .A1(\GFM/n2437 ), .A2(\GFM/n26050 ), .ZN(\GFM/N666 ));
NOR2_X2 \GFM/U1308  ( .A1(\GFM/n2478 ), .A2(\GFM/n26010 ), .ZN(\GFM/N662 ));
NOR2_X2 \GFM/U1307  ( .A1(\GFM/n2478 ), .A2(\GFM/n2602 ), .ZN(\GFM/N693 ) );
NOR2_X2 \GFM/U1306  ( .A1(\GFM/n2606 ), .A2(\GFM/n24360 ), .ZN(\GFM/N697 ));
NOR2_X2 \GFM/U1305  ( .A1(\GFM/n24770 ), .A2(\GFM/n2604 ), .ZN(\GFM/N755 ));
NOR2_X2 \GFM/U1304  ( .A1(\GFM/n26080 ), .A2(\GFM/n24360 ), .ZN(\GFM/N759 ));
NOR2_X2 \GFM/U1303  ( .A1(\GFM/n24380 ), .A2(\GFM/n2609 ), .ZN(\GFM/N790 ));
NOR2_X2 \GFM/U1302  ( .A1(\GFM/n2480 ), .A2(\GFM/n26050 ), .ZN(\GFM/N786 ));
NOR2_X2 \GFM/U1301  ( .A1(\GFM/n2606 ), .A2(\GFM/n24770 ), .ZN(\GFM/N817 ));
NOR2_X2 \GFM/U1300  ( .A1(\GFM/n2610 ), .A2(\GFM/n24360 ), .ZN(\GFM/N821 ));
NOR2_X2 \GFM/U1299  ( .A1(\GFM/n2517 ), .A2(\GFM/n2603 ), .ZN(\GFM/N841 ) );
NOR2_X2 \GFM/U1298  ( .A1(\GFM/n24960 ), .A2(\GFM/n26050 ), .ZN(\GFM/N844 ));
NOR2_X2 \GFM/U1297  ( .A1(\GFM/n26080 ), .A2(\GFM/n24770 ), .ZN(\GFM/N879 ));
NOR2_X2 \GFM/U1296  ( .A1(\GFM/n26120 ), .A2(\GFM/n24360 ), .ZN(\GFM/N883 ));
NOR2_X2 \GFM/U1295  ( .A1(\GFM/n2517 ), .A2(\GFM/n26050 ), .ZN(\GFM/N903 ));
NOR2_X2 \GFM/U1294  ( .A1(\GFM/n24960 ), .A2(\GFM/n26070 ), .ZN(\GFM/N906 ));
NOR2_X2 \GFM/U1293  ( .A1(\GFM/n2441 ), .A2(\GFM/n26150 ), .ZN(\GFM/N976 ));
NOR2_X2 \GFM/U1292  ( .A1(\GFM/n24810 ), .A2(\GFM/n26110 ), .ZN(\GFM/N972 ));
NOR2_X2 \GFM/U1291  ( .A1(\GFM/n24450 ), .A2(\GFM/n25821 ), .ZN(\GFM/N15 ));
NOR2_X2 \GFM/U1290  ( .A1(\GFM/n2485 ), .A2(\GFM/n2573 ), .ZN(\GFM/N11 ) );
NOR2_X2 \GFM/U1289  ( .A1(\GFM/n24380 ), .A2(\GFM/n25840 ), .ZN(\GFM/N46 ));
NOR2_X2 \GFM/U1288  ( .A1(\GFM/n2478 ), .A2(\GFM/n25760 ), .ZN(\GFM/N42 ) );
NOR2_X2 \GFM/U1287  ( .A1(\GFM/n2437 ), .A2(\GFM/n2587 ), .ZN(\GFM/N108 ) );
NOR2_X2 \GFM/U1286  ( .A1(\GFM/n2479 ), .A2(\GFM/n25800 ), .ZN(\GFM/N104 ));
NOR2_X2 \GFM/U1285  ( .A1(\GFM/n2485 ), .A2(\GFM/n25821 ), .ZN(\GFM/N135 ));
NOR2_X2 \GFM/U1284  ( .A1(\GFM/n25880 ), .A2(\GFM/n24360 ), .ZN(\GFM/N139 ));
NOR2_X2 \GFM/U1283  ( .A1(\GFM/n25890 ), .A2(\GFM/n2437 ), .ZN(\GFM/N170 ));
NOR2_X2 \GFM/U1282  ( .A1(\GFM/n24840 ), .A2(\GFM/n25840 ), .ZN(\GFM/N166 ));
NOR2_X2 \GFM/U1281  ( .A1(\GFM/n2616 ), .A2(\GFM/n24360 ), .ZN(\GFM/N1007 ));
NOR2_X2 \GFM/U1280  ( .A1(\GFM/n26120 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1003 ));
NOR2_X2 \GFM/U1279  ( .A1(\GFM/n2617 ), .A2(\GFM/n24360 ), .ZN(\GFM/N1038 ));
NOR2_X2 \GFM/U1278  ( .A1(\GFM/n2613 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1034 ));
NOR2_X2 \GFM/U1277  ( .A1(\GFM/n2618 ), .A2(\GFM/n24360 ), .ZN(\GFM/N1069 ));
NOR2_X2 \GFM/U1276  ( .A1(\GFM/n26140 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1065 ));
NOR2_X2 \GFM/U1275  ( .A1(\GFM/n25050 ), .A2(\GFM/n2618 ), .ZN(\GFM/N1247 ));
NOR2_X2 \GFM/U1274  ( .A1(\GFM/n2525 ), .A2(\GFM/n2616 ), .ZN(\GFM/N1244 ));
NOR2_X2 \GFM/U1273  ( .A1(\GFM/n24450 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1317 ));
NOR2_X2 \GFM/U1272  ( .A1(\GFM/n2485 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1313 ));
NOR2_X2 \GFM/U1271  ( .A1(\GFM/n24450 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1348 ));
NOR2_X2 \GFM/U1270  ( .A1(\GFM/n2485 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1344 ));
NOR2_X2 \GFM/U1269  ( .A1(\GFM/n24450 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1379 ));
NOR2_X2 \GFM/U1268  ( .A1(\GFM/n2485 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1375 ));
NOR2_X2 \GFM/U1267  ( .A1(\GFM/n24450 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1410 ));
NOR2_X2 \GFM/U1266  ( .A1(\GFM/n2485 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1406 ));
NOR2_X2 \GFM/U1265  ( .A1(\GFM/n24450 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1441 ));
NOR2_X2 \GFM/U1264  ( .A1(\GFM/n2485 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1437 ));
NOR2_X2 \GFM/U1263  ( .A1(\GFM/n24450 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1472 ));
NOR2_X2 \GFM/U1262  ( .A1(\GFM/n2485 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1468 ));
NOR2_X2 \GFM/U1261  ( .A1(\GFM/n2444 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1503 ));
NOR2_X2 \GFM/U1260  ( .A1(\GFM/n2485 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1499 ));
NOR2_X2 \GFM/U1259  ( .A1(\GFM/n2444 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1534 ));
NOR2_X2 \GFM/U1258  ( .A1(\GFM/n2485 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1530 ));
NOR2_X2 \GFM/U1257  ( .A1(\GFM/n2444 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1565 ));
NOR2_X2 \GFM/U1256  ( .A1(\GFM/n2485 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1561 ));
NOR2_X2 \GFM/U1255  ( .A1(\GFM/n2444 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1596 ));
NOR2_X2 \GFM/U1254  ( .A1(\GFM/n24840 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1592 ));
NOR2_X2 \GFM/U1253  ( .A1(\GFM/n2444 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1627 ));
NOR2_X2 \GFM/U1252  ( .A1(\GFM/n24840 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1623 ));
NOR2_X2 \GFM/U1251  ( .A1(\GFM/n2444 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1658 ));
NOR2_X2 \GFM/U1250  ( .A1(\GFM/n24840 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1654 ));
NOR2_X2 \GFM/U1249  ( .A1(\GFM/n2444 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1689 ));
NOR2_X2 \GFM/U1248  ( .A1(\GFM/n24840 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1685 ));
NOR2_X2 \GFM/U1247  ( .A1(\GFM/n2444 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1720 ));
NOR2_X2 \GFM/U1246  ( .A1(\GFM/n24840 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1716 ));
NOR2_X2 \GFM/U1245  ( .A1(\GFM/n2444 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1751 ));
NOR2_X2 \GFM/U1244  ( .A1(\GFM/n24840 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1747 ));
NOR2_X2 \GFM/U1243  ( .A1(\GFM/n2444 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1782 ));
NOR2_X2 \GFM/U1242  ( .A1(\GFM/n24840 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1778 ));
NOR2_X2 \GFM/U1241  ( .A1(\GFM/n2444 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1813 ));
NOR2_X2 \GFM/U1240  ( .A1(\GFM/n24840 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1809 ));
NOR2_X2 \GFM/U1239  ( .A1(\GFM/n2444 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1844 ));
NOR2_X2 \GFM/U1238  ( .A1(\GFM/n24840 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1840 ));
NOR2_X2 \GFM/U1237  ( .A1(\GFM/n2444 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1875 ));
NOR2_X2 \GFM/U1236  ( .A1(\GFM/n24840 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1871 ));
NOR2_X2 \GFM/U1235  ( .A1(\GFM/n24430 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1906 ));
NOR2_X2 \GFM/U1234  ( .A1(\GFM/n24840 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1902 ));
NOR2_X2 \GFM/U1233  ( .A1(\GFM/n24430 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1937 ));
NOR2_X2 \GFM/U1232  ( .A1(\GFM/n24840 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1933 ));
NOR2_X2 \GFM/U1231  ( .A1(\GFM/n24430 ), .A2(\GFM/n2647 ), .ZN(\GFM/N1968 ));
NOR2_X2 \GFM/U1230  ( .A1(\GFM/n24830 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1964 ));
NOR2_X2 \GFM/U1229  ( .A1(\GFM/n24430 ), .A2(\GFM/n2648 ), .ZN(\GFM/N1999 ));
NOR2_X2 \GFM/U1228  ( .A1(\GFM/n24830 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1995 ));
NOR2_X2 \GFM/U1227  ( .A1(\GFM/n24430 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2030 ));
NOR2_X2 \GFM/U1226  ( .A1(\GFM/n24830 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2026 ));
NOR2_X2 \GFM/U1225  ( .A1(\GFM/n24430 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2061 ));
NOR2_X2 \GFM/U1224  ( .A1(\GFM/n24830 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2057 ));
NOR2_X2 \GFM/U1223  ( .A1(\GFM/n24430 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2092 ));
NOR2_X2 \GFM/U1222  ( .A1(\GFM/n24830 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2088 ));
NOR2_X2 \GFM/U1221  ( .A1(\GFM/n24430 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2123 ));
NOR2_X2 \GFM/U1220  ( .A1(\GFM/n24830 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2119 ));
NOR2_X2 \GFM/U1219  ( .A1(\GFM/n24430 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2154 ));
NOR2_X2 \GFM/U1218  ( .A1(\GFM/n24830 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2150 ));
NOR2_X2 \GFM/U1217  ( .A1(\GFM/n24430 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2185 ));
NOR2_X2 \GFM/U1216  ( .A1(\GFM/n24830 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2181 ));
NOR2_X2 \GFM/U1215  ( .A1(\GFM/n24430 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2216 ));
NOR2_X2 \GFM/U1214  ( .A1(\GFM/n24830 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2212 ));
NOR2_X2 \GFM/U1213  ( .A1(\GFM/n24430 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2247 ));
NOR2_X2 \GFM/U1212  ( .A1(\GFM/n24830 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2243 ));
NOR2_X2 \GFM/U1211  ( .A1(\GFM/n24420 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2278 ));
NOR2_X2 \GFM/U1210  ( .A1(\GFM/n24830 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2274 ));
NOR2_X2 \GFM/U1209  ( .A1(\GFM/n24420 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2309 ));
NOR2_X2 \GFM/U1208  ( .A1(\GFM/n2482 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2305 ));
NOR2_X2 \GFM/U1207  ( .A1(\GFM/n24420 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2340 ));
NOR2_X2 \GFM/U1206  ( .A1(\GFM/n2482 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2336 ));
NOR2_X2 \GFM/U1205  ( .A1(\GFM/n24420 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2371 ));
NOR2_X2 \GFM/U1204  ( .A1(\GFM/n2482 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2367 ));
NOR2_X2 \GFM/U1203  ( .A1(\GFM/n24420 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2402 ));
NOR2_X2 \GFM/U1202  ( .A1(\GFM/n2482 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2398 ));
NOR2_X2 \GFM/U1201  ( .A1(\GFM/n24420 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2433 ));
NOR2_X2 \GFM/U1200  ( .A1(\GFM/n2482 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2429 ));
NOR2_X2 \GFM/U1199  ( .A1(\GFM/n24420 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2464 ));
NOR2_X2 \GFM/U1198  ( .A1(\GFM/n2482 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2460 ));
NOR2_X2 \GFM/U1197  ( .A1(\GFM/n24420 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2495 ));
NOR2_X2 \GFM/U1196  ( .A1(\GFM/n2482 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2491 ));
NOR2_X2 \GFM/U1195  ( .A1(\GFM/n24420 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2526 ));
NOR2_X2 \GFM/U1194  ( .A1(\GFM/n2482 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2522 ));
NOR2_X2 \GFM/U1193  ( .A1(\GFM/n24420 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2557 ));
NOR2_X2 \GFM/U1192  ( .A1(\GFM/n2482 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2553 ));
NOR2_X2 \GFM/U1191  ( .A1(\GFM/n24420 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2588 ));
NOR2_X2 \GFM/U1190  ( .A1(\GFM/n2482 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2584 ));
NOR2_X2 \GFM/U1189  ( .A1(\GFM/n24420 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2619 ));
NOR2_X2 \GFM/U1188  ( .A1(\GFM/n2482 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2615 ));
NOR2_X2 \GFM/U1187  ( .A1(\GFM/n2441 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2650 ));
NOR2_X2 \GFM/U1186  ( .A1(\GFM/n2482 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2646 ));
NOR2_X2 \GFM/U1185  ( .A1(\GFM/n2441 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2681 ));
NOR2_X2 \GFM/U1184  ( .A1(\GFM/n2482 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2677 ));
NOR2_X2 \GFM/U1183  ( .A1(\GFM/n2441 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2712 ));
NOR2_X2 \GFM/U1182  ( .A1(\GFM/n24810 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2708 ));
NOR2_X2 \GFM/U1181  ( .A1(\GFM/n2441 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2743 ));
NOR2_X2 \GFM/U1180  ( .A1(\GFM/n24810 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2739 ));
NOR2_X2 \GFM/U1179  ( .A1(\GFM/n2441 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2774 ));
NOR2_X2 \GFM/U1178  ( .A1(\GFM/n24810 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2770 ));
NOR2_X2 \GFM/U1177  ( .A1(\GFM/n2441 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2805 ));
NOR2_X2 \GFM/U1176  ( .A1(\GFM/n24810 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2801 ));
NOR2_X2 \GFM/U1175  ( .A1(\GFM/n2441 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2836 ));
NOR2_X2 \GFM/U1174  ( .A1(\GFM/n24810 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2832 ));
NOR2_X2 \GFM/U1173  ( .A1(\GFM/n2441 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2867 ));
NOR2_X2 \GFM/U1172  ( .A1(\GFM/n24810 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2863 ));
NOR2_X2 \GFM/U1171  ( .A1(\GFM/n2441 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2898 ));
NOR2_X2 \GFM/U1170  ( .A1(\GFM/n24810 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2894 ));
NOR2_X2 \GFM/U1169  ( .A1(\GFM/n2441 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2929 ));
NOR2_X2 \GFM/U1168  ( .A1(\GFM/n24810 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2925 ));
NOR2_X2 \GFM/U1167  ( .A1(\GFM/n24401 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2960 ));
NOR2_X2 \GFM/U1166  ( .A1(\GFM/n24810 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2956 ));
NOR2_X2 \GFM/U1165  ( .A1(\GFM/n24401 ), .A2(\GFM/n26801 ), .ZN(\GFM/N2991 ));
NOR2_X2 \GFM/U1164  ( .A1(\GFM/n24810 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2987 ));
NOR2_X2 \GFM/U1163  ( .A1(\GFM/n24401 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3022 ));
NOR2_X2 \GFM/U1162  ( .A1(\GFM/n24810 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3018 ));
NOR2_X2 \GFM/U1161  ( .A1(\GFM/n24401 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3053 ));
NOR2_X2 \GFM/U1160  ( .A1(\GFM/n2480 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3049 ));
NOR2_X2 \GFM/U1159  ( .A1(\GFM/n24401 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3084 ));
NOR2_X2 \GFM/U1158  ( .A1(\GFM/n2480 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3080 ));
NOR2_X2 \GFM/U1157  ( .A1(\GFM/n24401 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3115 ));
NOR2_X2 \GFM/U1156  ( .A1(\GFM/n2480 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3111 ));
NOR2_X2 \GFM/U1155  ( .A1(\GFM/n24401 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3146 ));
NOR2_X2 \GFM/U1154  ( .A1(\GFM/n2480 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3142 ));
NOR2_X2 \GFM/U1153  ( .A1(\GFM/n24401 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3177 ));
NOR2_X2 \GFM/U1152  ( .A1(\GFM/n2480 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3173 ));
NOR2_X2 \GFM/U1151  ( .A1(\GFM/n24401 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3208 ));
NOR2_X2 \GFM/U1150  ( .A1(\GFM/n2480 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3204 ));
NOR2_X2 \GFM/U1149  ( .A1(\GFM/n24401 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3239 ));
NOR2_X2 \GFM/U1148  ( .A1(\GFM/n24810 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3235 ));
NOR2_X2 \GFM/U1147  ( .A1(\GFM/n24401 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3270 ));
NOR2_X2 \GFM/U1146  ( .A1(\GFM/n2480 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3266 ));
NOR2_X2 \GFM/U1145  ( .A1(\GFM/n24690 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3299 ));
NOR2_X2 \GFM/U1144  ( .A1(\GFM/n2480 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3298 ));
NOR2_X2 \GFM/U1143  ( .A1(\GFM/n24690 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3331 ));
NOR2_X2 \GFM/U1142  ( .A1(\GFM/n2480 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3330 ));
NOR2_X2 \GFM/U1141  ( .A1(\GFM/n24690 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3364 ));
NOR2_X2 \GFM/U1140  ( .A1(\GFM/n2480 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3363 ));
NOR2_X2 \GFM/U1139  ( .A1(\GFM/n24390 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3407 ));
NOR2_X2 \GFM/U1138  ( .A1(\GFM/n2449 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3406 ));
NOR2_X2 \GFM/U1137  ( .A1(\GFM/n24390 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3444 ));
NOR2_X2 \GFM/U1136  ( .A1(\GFM/n2449 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3443 ));
NOR2_X2 \GFM/U1135  ( .A1(\GFM/n2499 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3466 ));
NOR2_X2 \GFM/U1134  ( .A1(\GFM/n25190 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3463 ));
NOR2_X2 \GFM/U1133  ( .A1(\GFM/n2509 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3505 ));
NOR2_X2 \GFM/U1132  ( .A1(\GFM/n25290 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3503 ));
NOR2_X2 \GFM/U1131  ( .A1(\GFM/n25101 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3548 ));
NOR2_X2 \GFM/U1130  ( .A1(\GFM/n25290 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3546 ));
NOR2_X2 \GFM/U1129  ( .A1(\GFM/n2509 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3594 ));
NOR2_X2 \GFM/U1128  ( .A1(\GFM/n2528 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3592 ));
NOR2_X2 \GFM/U1127  ( .A1(\GFM/n2509 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3643 ));
NOR2_X2 \GFM/U1126  ( .A1(\GFM/n2528 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3641 ));
NOR2_X2 \GFM/U1125  ( .A1(\GFM/n2509 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3695 ));
NOR2_X2 \GFM/U1124  ( .A1(\GFM/n2528 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3693 ));
NOR2_X2 \GFM/U1123  ( .A1(\GFM/n2697 ), .A2(\GFM/n25070 ), .ZN(\GFM/N3999 ));
NOR2_X2 \GFM/U1122  ( .A1(\GFM/n2695 ), .A2(\GFM/n25260 ), .ZN(\GFM/N3997 ));
NOR2_X2 \GFM/U1121  ( .A1(\GFM/n25890 ), .A2(\GFM/n24070 ), .ZN(\GFM/N86 ));
NOR2_X2 \GFM/U1120  ( .A1(\GFM/n25080 ), .A2(\GFM/n2573 ), .ZN(\GFM/N101 ));
NOR2_X2 \GFM/U1119  ( .A1(\GFM/n25890 ), .A2(\GFM/n25530 ), .ZN(\GFM/N118 ));
NOR2_X2 \GFM/U1118  ( .A1(\GFM/n24150 ), .A2(\GFM/n25910 ), .ZN(\GFM/N148 ));
NOR2_X2 \GFM/U1117  ( .A1(\GFM/n24140 ), .A2(\GFM/n2592 ), .ZN(\GFM/N179 ));
NOR2_X2 \GFM/U1116  ( .A1(\GFM/n24140 ), .A2(\GFM/n25930 ), .ZN(\GFM/N210 ));
NOR2_X2 \GFM/U1115  ( .A1(\GFM/n2413 ), .A2(\GFM/n25940 ), .ZN(\GFM/N241 ));
NOR2_X2 \GFM/U1114  ( .A1(\GFM/n24430 ), .A2(\GFM/n25901 ), .ZN(\GFM/N201 ));
NOR2_X2 \GFM/U1113  ( .A1(\GFM/n24830 ), .A2(\GFM/n2586 ), .ZN(\GFM/N197 ));
NOR2_X2 \GFM/U1112  ( .A1(\GFM/n24420 ), .A2(\GFM/n25910 ), .ZN(\GFM/N232 ));
NOR2_X2 \GFM/U1111  ( .A1(\GFM/n24830 ), .A2(\GFM/n2587 ), .ZN(\GFM/N228 ));
NOR2_X2 \GFM/U1110  ( .A1(\GFM/n2441 ), .A2(\GFM/n2592 ), .ZN(\GFM/N263 ) );
NOR2_X2 \GFM/U1109  ( .A1(\GFM/n25880 ), .A2(\GFM/n24770 ), .ZN(\GFM/N259 ));
NOR2_X2 \GFM/U1108  ( .A1(\GFM/n2441 ), .A2(\GFM/n25930 ), .ZN(\GFM/N294 ));
NOR2_X2 \GFM/U1107  ( .A1(\GFM/n25890 ), .A2(\GFM/n24770 ), .ZN(\GFM/N290 ));
NOR2_X2 \GFM/U1106  ( .A1(\GFM/n25890 ), .A2(\GFM/n2466 ), .ZN(\GFM/N269 ));
NOR2_X2 \GFM/U1105  ( .A1(\GFM/n24600 ), .A2(\GFM/n25910 ), .ZN(\GFM/N299 ));
NOR2_X2 \GFM/U1104  ( .A1(\GFM/n24600 ), .A2(\GFM/n2592 ), .ZN(\GFM/N330 ));
NOR2_X2 \GFM/U1103  ( .A1(\GFM/n24590 ), .A2(\GFM/n25930 ), .ZN(\GFM/N361 ));
NOR2_X2 \GFM/U1102  ( .A1(\GFM/n2458 ), .A2(\GFM/n25940 ), .ZN(\GFM/N392 ));
NOR2_X2 \GFM/U1101  ( .A1(\GFM/n25890 ), .A2(\GFM/n2516 ), .ZN(\GFM/N407 ));
NOR2_X2 \GFM/U1100  ( .A1(\GFM/n2458 ), .A2(\GFM/n2595 ), .ZN(\GFM/N423 ) );
NOR2_X2 \GFM/U1099  ( .A1(\GFM/n25180 ), .A2(\GFM/n25901 ), .ZN(\GFM/N438 ));
NOR2_X2 \GFM/U1098  ( .A1(\GFM/n2458 ), .A2(\GFM/n2596 ), .ZN(\GFM/N454 ) );
NOR2_X2 \GFM/U1097  ( .A1(\GFM/n2517 ), .A2(\GFM/n25910 ), .ZN(\GFM/N469 ));
NOR2_X2 \GFM/U1096  ( .A1(\GFM/n2458 ), .A2(\GFM/n25970 ), .ZN(\GFM/N485 ));
NOR2_X2 \GFM/U1095  ( .A1(\GFM/n25180 ), .A2(\GFM/n2592 ), .ZN(\GFM/N500 ));
NOR2_X2 \GFM/U1094  ( .A1(\GFM/n2458 ), .A2(\GFM/n25980 ), .ZN(\GFM/N516 ));
NOR2_X2 \GFM/U1093  ( .A1(\GFM/n25180 ), .A2(\GFM/n25930 ), .ZN(\GFM/N531 ));
NOR2_X2 \GFM/U1092  ( .A1(\GFM/n2458 ), .A2(\GFM/n2599 ), .ZN(\GFM/N547 ) );
NOR2_X2 \GFM/U1091  ( .A1(\GFM/n25180 ), .A2(\GFM/n25940 ), .ZN(\GFM/N562 ));
NOR2_X2 \GFM/U1090  ( .A1(\GFM/n24570 ), .A2(\GFM/n26000 ), .ZN(\GFM/N578 ));
NOR2_X2 \GFM/U1089  ( .A1(\GFM/n2517 ), .A2(\GFM/n2595 ), .ZN(\GFM/N593 ) );
NOR2_X2 \GFM/U1088  ( .A1(\GFM/n2458 ), .A2(\GFM/n26010 ), .ZN(\GFM/N609 ));
NOR2_X2 \GFM/U1087  ( .A1(\GFM/n25180 ), .A2(\GFM/n2596 ), .ZN(\GFM/N624 ));
NOR2_X2 \GFM/U1086  ( .A1(\GFM/n2517 ), .A2(\GFM/n25970 ), .ZN(\GFM/N655 ));
NOR2_X2 \GFM/U1085  ( .A1(\GFM/n2517 ), .A2(\GFM/n25980 ), .ZN(\GFM/N686 ));
NOR2_X2 \GFM/U1084  ( .A1(\GFM/n2517 ), .A2(\GFM/n2599 ), .ZN(\GFM/N717 ) );
NOR2_X2 \GFM/U1083  ( .A1(\GFM/n24570 ), .A2(\GFM/n26050 ), .ZN(\GFM/N733 ));
NOR2_X2 \GFM/U1082  ( .A1(\GFM/n2517 ), .A2(\GFM/n26010 ), .ZN(\GFM/N779 ));
NOR2_X2 \GFM/U1081  ( .A1(\GFM/n26070 ), .A2(\GFM/n24560 ), .ZN(\GFM/N795 ));
NOR2_X2 \GFM/U1080  ( .A1(\GFM/n26080 ), .A2(\GFM/n24560 ), .ZN(\GFM/N826 ));
NOR2_X2 \GFM/U1079  ( .A1(\GFM/n26080 ), .A2(\GFM/n2466 ), .ZN(\GFM/N858 ));
NOR2_X2 \GFM/U1078  ( .A1(\GFM/n2517 ), .A2(\GFM/n2604 ), .ZN(\GFM/N872 ) );
NOR2_X2 \GFM/U1077  ( .A1(\GFM/n2610 ), .A2(\GFM/n24560 ), .ZN(\GFM/N888 ));
NOR2_X2 \GFM/U1076  ( .A1(\GFM/n2610 ), .A2(\GFM/n2466 ), .ZN(\GFM/N920 ) );
NOR2_X2 \GFM/U1075  ( .A1(\GFM/n2525 ), .A2(\GFM/n2573 ), .ZN(\GFM/N128 ) );
NOR2_X2 \GFM/U1074  ( .A1(\GFM/n2524 ), .A2(\GFM/n25760 ), .ZN(\GFM/N159 ));
NOR2_X2 \GFM/U1073  ( .A1(\GFM/n2523 ), .A2(\GFM/n2578 ), .ZN(\GFM/N190 ) );
NOR2_X2 \GFM/U1072  ( .A1(\GFM/n25220 ), .A2(\GFM/n25800 ), .ZN(\GFM/N221 ));
NOR2_X2 \GFM/U1071  ( .A1(\GFM/n2613 ), .A2(\GFM/n24360 ), .ZN(\GFM/N914 ));
NOR2_X2 \GFM/U1070  ( .A1(\GFM/n2517 ), .A2(\GFM/n2606 ), .ZN(\GFM/N934 ) );
NOR2_X2 \GFM/U1069  ( .A1(\GFM/n26120 ), .A2(\GFM/n24560 ), .ZN(\GFM/N950 ));
NOR2_X2 \GFM/U1068  ( .A1(\GFM/n24960 ), .A2(\GFM/n2609 ), .ZN(\GFM/N968 ));
NOR2_X2 \GFM/U1067  ( .A1(\GFM/n2461 ), .A2(\GFM/n2613 ), .ZN(\GFM/N981 ) );
NOR2_X2 \GFM/U1066  ( .A1(\GFM/n2458 ), .A2(\GFM/n26140 ), .ZN(\GFM/N1012 ));
NOR2_X2 \GFM/U1065  ( .A1(\GFM/n2617 ), .A2(\GFM/n24560 ), .ZN(\GFM/N1105 ));
NOR2_X2 \GFM/U1064  ( .A1(\GFM/n2616 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1127 ));
NOR2_X2 \GFM/U1063  ( .A1(\GFM/n2618 ), .A2(\GFM/n24560 ), .ZN(\GFM/N1136 ));
NOR2_X2 \GFM/U1062  ( .A1(\GFM/n2617 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1158 ));
NOR2_X2 \GFM/U1061  ( .A1(\GFM/n26190 ), .A2(\GFM/n24560 ), .ZN(\GFM/N1167 ));
NOR2_X2 \GFM/U1060  ( .A1(\GFM/n2618 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1189 ));
NOR2_X2 \GFM/U1059  ( .A1(\GFM/n26200 ), .A2(\GFM/n24560 ), .ZN(\GFM/N1198 ));
NOR2_X2 \GFM/U1058  ( .A1(\GFM/n26190 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1220 ));
NOR2_X2 \GFM/U1057  ( .A1(\GFM/n26200 ), .A2(\GFM/n2466 ), .ZN(\GFM/N1230 ));
NOR2_X2 \GFM/U1056  ( .A1(\GFM/n26200 ), .A2(\GFM/n24760 ), .ZN(\GFM/N1251 ));
NOR2_X2 \GFM/U1055  ( .A1(\GFM/n24650 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1260 ));
NOR2_X2 \GFM/U1054  ( .A1(\GFM/n2485 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1282 ));
NOR2_X2 \GFM/U1053  ( .A1(\GFM/n24650 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1291 ));
NOR2_X2 \GFM/U1052  ( .A1(\GFM/n2525 ), .A2(\GFM/n2618 ), .ZN(\GFM/N1306 ));
NOR2_X2 \GFM/U1051  ( .A1(\GFM/n24650 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1322 ));
NOR2_X2 \GFM/U1050  ( .A1(\GFM/n24650 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1353 ));
NOR2_X2 \GFM/U1049  ( .A1(\GFM/n24650 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1384 ));
NOR2_X2 \GFM/U1048  ( .A1(\GFM/n24650 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1415 ));
NOR2_X2 \GFM/U1047  ( .A1(\GFM/n24650 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1446 ));
NOR2_X2 \GFM/U1046  ( .A1(\GFM/n24640 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1477 ));
NOR2_X2 \GFM/U1045  ( .A1(\GFM/n24640 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1508 ));
NOR2_X2 \GFM/U1044  ( .A1(\GFM/n24640 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1539 ));
NOR2_X2 \GFM/U1043  ( .A1(\GFM/n24640 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1570 ));
NOR2_X2 \GFM/U1042  ( .A1(\GFM/n24640 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1601 ));
NOR2_X2 \GFM/U1041  ( .A1(\GFM/n2524 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1616 ));
NOR2_X2 \GFM/U1040  ( .A1(\GFM/n24640 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1632 ));
NOR2_X2 \GFM/U1039  ( .A1(\GFM/n2524 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1647 ));
NOR2_X2 \GFM/U1038  ( .A1(\GFM/n24640 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1663 ));
NOR2_X2 \GFM/U1037  ( .A1(\GFM/n2524 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1678 ));
NOR2_X2 \GFM/U1036  ( .A1(\GFM/n24640 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1694 ));
NOR2_X2 \GFM/U1035  ( .A1(\GFM/n2524 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1709 ));
NOR2_X2 \GFM/U1034  ( .A1(\GFM/n24640 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1725 ));
NOR2_X2 \GFM/U1033  ( .A1(\GFM/n2524 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1740 ));
NOR2_X2 \GFM/U1032  ( .A1(\GFM/n24640 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1756 ));
NOR2_X2 \GFM/U1031  ( .A1(\GFM/n2523 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1771 ));
NOR2_X2 \GFM/U1030  ( .A1(\GFM/n24640 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1787 ));
NOR2_X2 \GFM/U1029  ( .A1(\GFM/n2523 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1802 ));
NOR2_X2 \GFM/U1028  ( .A1(\GFM/n24640 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1818 ));
NOR2_X2 \GFM/U1027  ( .A1(\GFM/n2523 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1833 ));
NOR2_X2 \GFM/U1026  ( .A1(\GFM/n2463 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1849 ));
NOR2_X2 \GFM/U1025  ( .A1(\GFM/n2523 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1864 ));
NOR2_X2 \GFM/U1024  ( .A1(\GFM/n2463 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1880 ));
NOR2_X2 \GFM/U1023  ( .A1(\GFM/n2523 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1895 ));
NOR2_X2 \GFM/U1022  ( .A1(\GFM/n2463 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1911 ));
NOR2_X2 \GFM/U1021  ( .A1(\GFM/n2523 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1926 ));
NOR2_X2 \GFM/U1020  ( .A1(\GFM/n2463 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1942 ));
NOR2_X2 \GFM/U1019  ( .A1(\GFM/n2523 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1957 ));
NOR2_X2 \GFM/U1018  ( .A1(\GFM/n2463 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1973 ));
NOR2_X2 \GFM/U1017  ( .A1(\GFM/n2523 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1988 ));
NOR2_X2 \GFM/U1016  ( .A1(\GFM/n2463 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2004 ));
NOR2_X2 \GFM/U1015  ( .A1(\GFM/n2523 ), .A2(\GFM/n2641 ), .ZN(\GFM/N2019 ));
NOR2_X2 \GFM/U1014  ( .A1(\GFM/n2463 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2035 ));
NOR2_X2 \GFM/U1013  ( .A1(\GFM/n2523 ), .A2(\GFM/n26420 ), .ZN(\GFM/N2050 ));
NOR2_X2 \GFM/U1012  ( .A1(\GFM/n2463 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2066 ));
NOR2_X2 \GFM/U1011  ( .A1(\GFM/n2523 ), .A2(\GFM/n26430 ), .ZN(\GFM/N2081 ));
NOR2_X2 \GFM/U1010  ( .A1(\GFM/n2463 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2097 ));
NOR2_X2 \GFM/U1009  ( .A1(\GFM/n2523 ), .A2(\GFM/n2644 ), .ZN(\GFM/N2112 ));
NOR2_X2 \GFM/U1008  ( .A1(\GFM/n2463 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2128 ));
NOR2_X2 \GFM/U1007  ( .A1(\GFM/n25220 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2143 ));
NOR2_X2 \GFM/U1006  ( .A1(\GFM/n2463 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2159 ));
NOR2_X2 \GFM/U1005  ( .A1(\GFM/n25220 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2174 ));
NOR2_X2 \GFM/U1004  ( .A1(\GFM/n2463 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2190 ));
NOR2_X2 \GFM/U1003  ( .A1(\GFM/n25220 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2205 ));
NOR2_X2 \GFM/U1002  ( .A1(\GFM/n2462 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2221 ));
NOR2_X2 \GFM/U1001  ( .A1(\GFM/n25220 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2236 ));
NOR2_X2 \GFM/U1000  ( .A1(\GFM/n2462 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2252 ));
NOR2_X2 \GFM/U999  ( .A1(\GFM/n25220 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2267 ));
NOR2_X2 \GFM/U998  ( .A1(\GFM/n2462 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2283 ));
NOR2_X2 \GFM/U997  ( .A1(\GFM/n25220 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2298 ));
NOR2_X2 \GFM/U996  ( .A1(\GFM/n2462 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2314 ));
NOR2_X2 \GFM/U995  ( .A1(\GFM/n25220 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2329 ));
NOR2_X2 \GFM/U994  ( .A1(\GFM/n2462 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2345 ) );
NOR2_X2 \GFM/U993  ( .A1(\GFM/n25220 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2360 ));
NOR2_X2 \GFM/U992  ( .A1(\GFM/n2462 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2376 ) );
NOR2_X2 \GFM/U991  ( .A1(\GFM/n25220 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2391 ));
NOR2_X2 \GFM/U990  ( .A1(\GFM/n2462 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2407 ));
NOR2_X2 \GFM/U989  ( .A1(\GFM/n25220 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2422 ));
NOR2_X2 \GFM/U988  ( .A1(\GFM/n2462 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2438 ));
NOR2_X2 \GFM/U987  ( .A1(\GFM/n25220 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2453 ));
NOR2_X2 \GFM/U986  ( .A1(\GFM/n2462 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2469 ));
NOR2_X2 \GFM/U985  ( .A1(\GFM/n25220 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2484 ));
NOR2_X2 \GFM/U984  ( .A1(\GFM/n2462 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2500 ));
NOR2_X2 \GFM/U983  ( .A1(\GFM/n25210 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2515 ));
NOR2_X2 \GFM/U982  ( .A1(\GFM/n2462 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2531 ));
NOR2_X2 \GFM/U981  ( .A1(\GFM/n25210 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2546 ));
NOR2_X2 \GFM/U980  ( .A1(\GFM/n2462 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2562 ) );
NOR2_X2 \GFM/U979  ( .A1(\GFM/n25210 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2577 ));
NOR2_X2 \GFM/U978  ( .A1(\GFM/n2462 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2593 ) );
NOR2_X2 \GFM/U977  ( .A1(\GFM/n25210 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2608 ));
NOR2_X2 \GFM/U976  ( .A1(\GFM/n2461 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2624 ) );
NOR2_X2 \GFM/U975  ( .A1(\GFM/n25210 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2639 ));
NOR2_X2 \GFM/U974  ( .A1(\GFM/n2461 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2655 ));
NOR2_X2 \GFM/U973  ( .A1(\GFM/n25210 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2670 ));
NOR2_X2 \GFM/U972  ( .A1(\GFM/n2461 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2686 ) );
NOR2_X2 \GFM/U971  ( .A1(\GFM/n25210 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2701 ));
NOR2_X2 \GFM/U970  ( .A1(\GFM/n2461 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2717 ));
NOR2_X2 \GFM/U969  ( .A1(\GFM/n25210 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2732 ));
NOR2_X2 \GFM/U968  ( .A1(\GFM/n2461 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2748 ));
NOR2_X2 \GFM/U967  ( .A1(\GFM/n25210 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2763 ));
NOR2_X2 \GFM/U966  ( .A1(\GFM/n2461 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2779 ) );
NOR2_X2 \GFM/U965  ( .A1(\GFM/n25210 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2794 ));
NOR2_X2 \GFM/U964  ( .A1(\GFM/n2461 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2810 ) );
NOR2_X2 \GFM/U963  ( .A1(\GFM/n25210 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2825 ));
NOR2_X2 \GFM/U962  ( .A1(\GFM/n2461 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2841 ));
NOR2_X2 \GFM/U961  ( .A1(\GFM/n25201 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2856 ));
NOR2_X2 \GFM/U960  ( .A1(\GFM/n2461 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2872 ));
NOR2_X2 \GFM/U959  ( .A1(\GFM/n25201 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2887 ));
NOR2_X2 \GFM/U958  ( .A1(\GFM/n2461 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2903 ) );
NOR2_X2 \GFM/U957  ( .A1(\GFM/n25201 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2918 ));
NOR2_X2 \GFM/U956  ( .A1(\GFM/n2461 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2934 ));
NOR2_X2 \GFM/U955  ( .A1(\GFM/n25201 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2949 ));
NOR2_X2 \GFM/U954  ( .A1(\GFM/n24600 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2965 ));
NOR2_X2 \GFM/U953  ( .A1(\GFM/n25201 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2980 ));
NOR2_X2 \GFM/U952  ( .A1(\GFM/n24600 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2996 ));
NOR2_X2 \GFM/U951  ( .A1(\GFM/n25201 ), .A2(\GFM/n26730 ), .ZN(\GFM/N3011 ));
NOR2_X2 \GFM/U950  ( .A1(\GFM/n24600 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3027 ));
NOR2_X2 \GFM/U949  ( .A1(\GFM/n25201 ), .A2(\GFM/n26740 ), .ZN(\GFM/N3042 ));
NOR2_X2 \GFM/U948  ( .A1(\GFM/n24600 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3058 ));
NOR2_X2 \GFM/U947  ( .A1(\GFM/n25201 ), .A2(\GFM/n2675 ), .ZN(\GFM/N3073 ));
NOR2_X2 \GFM/U946  ( .A1(\GFM/n24600 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3089 ));
NOR2_X2 \GFM/U945  ( .A1(\GFM/n25201 ), .A2(\GFM/n26760 ), .ZN(\GFM/N3104 ));
NOR2_X2 \GFM/U944  ( .A1(\GFM/n24600 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3120 ));
NOR2_X2 \GFM/U943  ( .A1(\GFM/n25201 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3135 ));
NOR2_X2 \GFM/U942  ( .A1(\GFM/n24600 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3151 ));
NOR2_X2 \GFM/U941  ( .A1(\GFM/n25201 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3166 ));
NOR2_X2 \GFM/U940  ( .A1(\GFM/n24600 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3182 ));
NOR2_X2 \GFM/U939  ( .A1(\GFM/n25190 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3197 ));
NOR2_X2 \GFM/U938  ( .A1(\GFM/n24600 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3213 ));
NOR2_X2 \GFM/U937  ( .A1(\GFM/n25190 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3228 ));
NOR2_X2 \GFM/U936  ( .A1(\GFM/n24600 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3244 ));
NOR2_X2 \GFM/U935  ( .A1(\GFM/n25190 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3259 ));
NOR2_X2 \GFM/U934  ( .A1(\GFM/n24600 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3275 ));
NOR2_X2 \GFM/U933  ( .A1(\GFM/n25190 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3290 ));
NOR2_X2 \GFM/U932  ( .A1(\GFM/n24190 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3306 ));
NOR2_X2 \GFM/U931  ( .A1(\GFM/n25190 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3322 ));
NOR2_X2 \GFM/U930  ( .A1(\GFM/n25190 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3355 ));
NOR2_X2 \GFM/U929  ( .A1(\GFM/n25190 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3389 ));
NOR2_X2 \GFM/U928  ( .A1(\GFM/n25190 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3425 ));
NOR2_X2 \GFM/U927  ( .A1(\GFM/n2432 ), .A2(\GFM/n2592 ), .ZN(\GFM/N235 ) );
NOR2_X2 \GFM/U926  ( .A1(\GFM/n24520 ), .A2(\GFM/n25901 ), .ZN(\GFM/N233 ));
NOR2_X2 \GFM/U925  ( .A1(\GFM/n2431 ), .A2(\GFM/n25930 ), .ZN(\GFM/N266 ) );
NOR2_X2 \GFM/U924  ( .A1(\GFM/n24511 ), .A2(\GFM/n25910 ), .ZN(\GFM/N264 ));
NOR2_X2 \GFM/U923  ( .A1(\GFM/n2430 ), .A2(\GFM/n25940 ), .ZN(\GFM/N297 ) );
NOR2_X2 \GFM/U922  ( .A1(\GFM/n24511 ), .A2(\GFM/n2592 ), .ZN(\GFM/N295 ) );
NOR2_X2 \GFM/U921  ( .A1(\GFM/n2430 ), .A2(\GFM/n2595 ), .ZN(\GFM/N328 ) );
NOR2_X2 \GFM/U920  ( .A1(\GFM/n24500 ), .A2(\GFM/n25930 ), .ZN(\GFM/N326 ));
NOR2_X2 \GFM/U919  ( .A1(\GFM/n24290 ), .A2(\GFM/n2596 ), .ZN(\GFM/N359 ) );
NOR2_X2 \GFM/U918  ( .A1(\GFM/n2449 ), .A2(\GFM/n25940 ), .ZN(\GFM/N357 ) );
NOR2_X2 \GFM/U917  ( .A1(\GFM/n24280 ), .A2(\GFM/n25970 ), .ZN(\GFM/N390 ));
NOR2_X2 \GFM/U916  ( .A1(\GFM/n2449 ), .A2(\GFM/n2595 ), .ZN(\GFM/N388 ) );
NOR2_X2 \GFM/U915  ( .A1(\GFM/n24280 ), .A2(\GFM/n25980 ), .ZN(\GFM/N421 ));
NOR2_X2 \GFM/U914  ( .A1(\GFM/n2448 ), .A2(\GFM/n2596 ), .ZN(\GFM/N419 ) );
NOR2_X2 \GFM/U913  ( .A1(\GFM/n24290 ), .A2(\GFM/n2599 ), .ZN(\GFM/N452 ) );
NOR2_X2 \GFM/U912  ( .A1(\GFM/n2448 ), .A2(\GFM/n25970 ), .ZN(\GFM/N450 ) );
NOR2_X2 \GFM/U911  ( .A1(\GFM/n24280 ), .A2(\GFM/n26000 ), .ZN(\GFM/N483 ));
NOR2_X2 \GFM/U910  ( .A1(\GFM/n2448 ), .A2(\GFM/n25980 ), .ZN(\GFM/N481 ) );
NOR2_X2 \GFM/U909  ( .A1(\GFM/n24280 ), .A2(\GFM/n26010 ), .ZN(\GFM/N514 ));
NOR2_X2 \GFM/U908  ( .A1(\GFM/n2448 ), .A2(\GFM/n2599 ), .ZN(\GFM/N512 ) );
NOR2_X2 \GFM/U907  ( .A1(\GFM/n24280 ), .A2(\GFM/n2602 ), .ZN(\GFM/N545 ) );
NOR2_X2 \GFM/U906  ( .A1(\GFM/n2448 ), .A2(\GFM/n26000 ), .ZN(\GFM/N543 ) );
NOR2_X2 \GFM/U905  ( .A1(\GFM/n24280 ), .A2(\GFM/n2603 ), .ZN(\GFM/N576 ) );
NOR2_X2 \GFM/U904  ( .A1(\GFM/n2448 ), .A2(\GFM/n26010 ), .ZN(\GFM/N574 ) );
NOR2_X2 \GFM/U903  ( .A1(\GFM/n26070 ), .A2(\GFM/n2427 ), .ZN(\GFM/N700 ) );
NOR2_X2 \GFM/U902  ( .A1(\GFM/n2447 ), .A2(\GFM/n26050 ), .ZN(\GFM/N698 ) );
NOR2_X2 \GFM/U901  ( .A1(\GFM/n24280 ), .A2(\GFM/n2609 ), .ZN(\GFM/N762 ) );
NOR2_X2 \GFM/U900  ( .A1(\GFM/n26070 ), .A2(\GFM/n2447 ), .ZN(\GFM/N760 ) );
NOR2_X2 \GFM/U899  ( .A1(\GFM/n2610 ), .A2(\GFM/n24260 ), .ZN(\GFM/N793 ) );
NOR2_X2 \GFM/U898  ( .A1(\GFM/n26080 ), .A2(\GFM/n24460 ), .ZN(\GFM/N791 ));
NOR2_X2 \GFM/U897  ( .A1(\GFM/n24280 ), .A2(\GFM/n26110 ), .ZN(\GFM/N824 ));
NOR2_X2 \GFM/U896  ( .A1(\GFM/n2447 ), .A2(\GFM/n2609 ), .ZN(\GFM/N822 ) );
NOR2_X2 \GFM/U895  ( .A1(\GFM/n25080 ), .A2(\GFM/n2604 ), .ZN(\GFM/N845 ) );
NOR2_X2 \GFM/U894  ( .A1(\GFM/n2606 ), .A2(\GFM/n2486 ), .ZN(\GFM/N847 ) );
NOR2_X2 \GFM/U893  ( .A1(\GFM/n2447 ), .A2(\GFM/n26110 ), .ZN(\GFM/N884 ) );
NOR2_X2 \GFM/U892  ( .A1(\GFM/n2613 ), .A2(\GFM/n24260 ), .ZN(\GFM/N886 ) );
NOR2_X2 \GFM/U891  ( .A1(\GFM/n2606 ), .A2(\GFM/n25070 ), .ZN(\GFM/N907 ) );
NOR2_X2 \GFM/U890  ( .A1(\GFM/n26080 ), .A2(\GFM/n2486 ), .ZN(\GFM/N909 ) );
NOR2_X2 \GFM/U889  ( .A1(\GFM/n2447 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1008 ));
NOR2_X2 \GFM/U888  ( .A1(\GFM/n2617 ), .A2(\GFM/n24260 ), .ZN(\GFM/N1010 ));
NOR2_X2 \GFM/U887  ( .A1(\GFM/n2618 ), .A2(\GFM/n24260 ), .ZN(\GFM/N1041 ));
NOR2_X2 \GFM/U886  ( .A1(\GFM/n2616 ), .A2(\GFM/n24460 ), .ZN(\GFM/N1039 ));
NOR2_X2 \GFM/U885  ( .A1(\GFM/n26200 ), .A2(\GFM/n24260 ), .ZN(\GFM/N1103 ));
NOR2_X2 \GFM/U884  ( .A1(\GFM/n2618 ), .A2(\GFM/n24460 ), .ZN(\GFM/N1101 ));
NOR2_X2 \GFM/U883  ( .A1(\GFM/n2616 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1157 ) );
NOR2_X2 \GFM/U882  ( .A1(\GFM/n26140 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1155 ));
NOR2_X2 \GFM/U881  ( .A1(\GFM/n2618 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1219 ) );
NOR2_X2 \GFM/U880  ( .A1(\GFM/n2616 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1217 ) );
NOR2_X2 \GFM/U879  ( .A1(\GFM/n26200 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1281 ));
NOR2_X2 \GFM/U878  ( .A1(\GFM/n2618 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1279 ) );
NOR2_X2 \GFM/U877  ( .A1(\GFM/n24340 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1537 ));
NOR2_X2 \GFM/U876  ( .A1(\GFM/n2454 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1535 ));
NOR2_X2 \GFM/U875  ( .A1(\GFM/n24340 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1568 ));
NOR2_X2 \GFM/U874  ( .A1(\GFM/n2454 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1566 ) );
NOR2_X2 \GFM/U873  ( .A1(\GFM/n24340 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1599 ));
NOR2_X2 \GFM/U872  ( .A1(\GFM/n2454 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1597 ) );
NOR2_X2 \GFM/U871  ( .A1(\GFM/n24340 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1630 ));
NOR2_X2 \GFM/U870  ( .A1(\GFM/n2454 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1628 ) );
NOR2_X2 \GFM/U869  ( .A1(\GFM/n24340 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1661 ));
NOR2_X2 \GFM/U868  ( .A1(\GFM/n2454 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1659 ));
NOR2_X2 \GFM/U867  ( .A1(\GFM/n24340 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1692 ));
NOR2_X2 \GFM/U866  ( .A1(\GFM/n2454 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1690 ) );
NOR2_X2 \GFM/U865  ( .A1(\GFM/n24340 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1723 ));
NOR2_X2 \GFM/U864  ( .A1(\GFM/n2454 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1721 ));
NOR2_X2 \GFM/U863  ( .A1(\GFM/n24340 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1754 ));
NOR2_X2 \GFM/U862  ( .A1(\GFM/n2454 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1752 ));
NOR2_X2 \GFM/U861  ( .A1(\GFM/n24340 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1785 ));
NOR2_X2 \GFM/U860  ( .A1(\GFM/n2454 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1783 ));
NOR2_X2 \GFM/U859  ( .A1(\GFM/n24340 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1816 ));
NOR2_X2 \GFM/U858  ( .A1(\GFM/n2454 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1814 ) );
NOR2_X2 \GFM/U857  ( .A1(\GFM/n24340 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1847 ));
NOR2_X2 \GFM/U856  ( .A1(\GFM/n2454 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1845 ));
NOR2_X2 \GFM/U855  ( .A1(\GFM/n24330 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1878 ));
NOR2_X2 \GFM/U854  ( .A1(\GFM/n24530 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1876 ));
NOR2_X2 \GFM/U853  ( .A1(\GFM/n24330 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1909 ));
NOR2_X2 \GFM/U852  ( .A1(\GFM/n24530 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1907 ));
NOR2_X2 \GFM/U851  ( .A1(\GFM/n24330 ), .A2(\GFM/n2647 ), .ZN(\GFM/N1940 ));
NOR2_X2 \GFM/U850  ( .A1(\GFM/n24530 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1938 ));
NOR2_X2 \GFM/U849  ( .A1(\GFM/n24330 ), .A2(\GFM/n2648 ), .ZN(\GFM/N1971 ));
NOR2_X2 \GFM/U848  ( .A1(\GFM/n24530 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1969 ));
NOR2_X2 \GFM/U847  ( .A1(\GFM/n24330 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2095 ));
NOR2_X2 \GFM/U846  ( .A1(\GFM/n24530 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2093 ));
NOR2_X2 \GFM/U845  ( .A1(\GFM/n24330 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2126 ));
NOR2_X2 \GFM/U844  ( .A1(\GFM/n24530 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2124 ));
NOR2_X2 \GFM/U843  ( .A1(\GFM/n24330 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2157 ));
NOR2_X2 \GFM/U842  ( .A1(\GFM/n24530 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2155 ));
NOR2_X2 \GFM/U841  ( .A1(\GFM/n24330 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2188 ));
NOR2_X2 \GFM/U840  ( .A1(\GFM/n24530 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2186 ));
NOR2_X2 \GFM/U839  ( .A1(\GFM/n24330 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2219 ));
NOR2_X2 \GFM/U838  ( .A1(\GFM/n24530 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2217 ));
NOR2_X2 \GFM/U837  ( .A1(\GFM/n2432 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2250 ) );
NOR2_X2 \GFM/U836  ( .A1(\GFM/n24530 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2248 ));
NOR2_X2 \GFM/U835  ( .A1(\GFM/n2432 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2281 ) );
NOR2_X2 \GFM/U834  ( .A1(\GFM/n24520 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2279 ));
NOR2_X2 \GFM/U833  ( .A1(\GFM/n2432 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2312 ));
NOR2_X2 \GFM/U832  ( .A1(\GFM/n24520 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2310 ));
NOR2_X2 \GFM/U831  ( .A1(\GFM/n2432 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2343 ));
NOR2_X2 \GFM/U830  ( .A1(\GFM/n24520 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2341 ));
NOR2_X2 \GFM/U829  ( .A1(\GFM/n2432 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2374 ));
NOR2_X2 \GFM/U828  ( .A1(\GFM/n24520 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2372 ));
NOR2_X2 \GFM/U827  ( .A1(\GFM/n2432 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2405 ));
NOR2_X2 \GFM/U826  ( .A1(\GFM/n24520 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2403 ));
NOR2_X2 \GFM/U825  ( .A1(\GFM/n2432 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2436 ));
NOR2_X2 \GFM/U824  ( .A1(\GFM/n24520 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2434 ));
NOR2_X2 \GFM/U823  ( .A1(\GFM/n2432 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2467 ) );
NOR2_X2 \GFM/U822  ( .A1(\GFM/n24520 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2465 ));
NOR2_X2 \GFM/U821  ( .A1(\GFM/n2432 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2498 ) );
NOR2_X2 \GFM/U820  ( .A1(\GFM/n24520 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2496 ));
NOR2_X2 \GFM/U819  ( .A1(\GFM/n2432 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2529 ) );
NOR2_X2 \GFM/U818  ( .A1(\GFM/n24520 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2527 ));
NOR2_X2 \GFM/U817  ( .A1(\GFM/n2432 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2560 ));
NOR2_X2 \GFM/U816  ( .A1(\GFM/n24520 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2558 ));
NOR2_X2 \GFM/U815  ( .A1(\GFM/n2432 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2591 ) );
NOR2_X2 \GFM/U814  ( .A1(\GFM/n24520 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2589 ));
NOR2_X2 \GFM/U813  ( .A1(\GFM/n2431 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2622 ));
NOR2_X2 \GFM/U812  ( .A1(\GFM/n24520 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2620 ));
NOR2_X2 \GFM/U811  ( .A1(\GFM/n2431 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2653 ));
NOR2_X2 \GFM/U810  ( .A1(\GFM/n24511 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2651 ));
NOR2_X2 \GFM/U809  ( .A1(\GFM/n2431 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2684 ) );
NOR2_X2 \GFM/U808  ( .A1(\GFM/n24511 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2682 ));
NOR2_X2 \GFM/U807  ( .A1(\GFM/n2431 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2715 ) );
NOR2_X2 \GFM/U806  ( .A1(\GFM/n24511 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2713 ));
NOR2_X2 \GFM/U805  ( .A1(\GFM/n2431 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2746 ));
NOR2_X2 \GFM/U804  ( .A1(\GFM/n24511 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2744 ));
NOR2_X2 \GFM/U803  ( .A1(\GFM/n2463 ), .A2(\GFM/n2578 ), .ZN(\GFM/N20 ) );
NOR2_X2 \GFM/U802  ( .A1(\GFM/n25210 ), .A2(\GFM/n25821 ), .ZN(\GFM/N252 ));
NOR2_X2 \GFM/U801  ( .A1(\GFM/n2617 ), .A2(\GFM/n2486 ), .ZN(\GFM/N1188 ) );
NOR2_X2 \GFM/U800  ( .A1(\GFM/n26150 ), .A2(\GFM/n2506 ), .ZN(\GFM/N1186 ));
NOR2_X2 \GFM/U799  ( .A1(\GFM/n2431 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2777 ));
NOR2_X2 \GFM/U798  ( .A1(\GFM/n24511 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2775 ));
NOR2_X2 \GFM/U797  ( .A1(\GFM/n2431 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2808 ) );
NOR2_X2 \GFM/U796  ( .A1(\GFM/n24511 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2806 ));
NOR2_X2 \GFM/U795  ( .A1(\GFM/n2431 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2839 ));
NOR2_X2 \GFM/U794  ( .A1(\GFM/n24511 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2837 ));
NOR2_X2 \GFM/U793  ( .A1(\GFM/n2431 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2870 ));
NOR2_X2 \GFM/U792  ( .A1(\GFM/n24511 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2868 ));
NOR2_X2 \GFM/U791  ( .A1(\GFM/n2431 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2901 ) );
NOR2_X2 \GFM/U790  ( .A1(\GFM/n24511 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2899 ));
NOR2_X2 \GFM/U789  ( .A1(\GFM/n2431 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2932 ) );
NOR2_X2 \GFM/U788  ( .A1(\GFM/n24511 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2930 ));
NOR2_X2 \GFM/U787  ( .A1(\GFM/n2430 ), .A2(\GFM/n26801 ), .ZN(\GFM/N2963 ));
NOR2_X2 \GFM/U786  ( .A1(\GFM/n24500 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2961 ));
NOR2_X2 \GFM/U785  ( .A1(\GFM/n2430 ), .A2(\GFM/n26810 ), .ZN(\GFM/N2994 ));
NOR2_X2 \GFM/U784  ( .A1(\GFM/n24500 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2992 ));
NOR2_X2 \GFM/U783  ( .A1(\GFM/n2430 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3025 ));
NOR2_X2 \GFM/U782  ( .A1(\GFM/n24500 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3023 ));
NOR2_X2 \GFM/U781  ( .A1(\GFM/n2430 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3056 ) );
NOR2_X2 \GFM/U780  ( .A1(\GFM/n24500 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3054 ));
NOR2_X2 \GFM/U779  ( .A1(\GFM/n2430 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3087 ));
NOR2_X2 \GFM/U778  ( .A1(\GFM/n24500 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3085 ));
NOR2_X2 \GFM/U777  ( .A1(\GFM/n2430 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3118 ) );
NOR2_X2 \GFM/U776  ( .A1(\GFM/n24500 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3116 ));
NOR2_X2 \GFM/U775  ( .A1(\GFM/n2430 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3149 ));
NOR2_X2 \GFM/U774  ( .A1(\GFM/n24500 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3147 ));
NOR2_X2 \GFM/U773  ( .A1(\GFM/n2430 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3180 ));
NOR2_X2 \GFM/U772  ( .A1(\GFM/n24500 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3178 ));
NOR2_X2 \GFM/U771  ( .A1(\GFM/n2430 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3211 ) );
NOR2_X2 \GFM/U770  ( .A1(\GFM/n24500 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3209 ));
NOR2_X2 \GFM/U769  ( .A1(\GFM/n2430 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3242 ) );
NOR2_X2 \GFM/U768  ( .A1(\GFM/n24500 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3240 ));
NOR2_X2 \GFM/U767  ( .A1(\GFM/n2430 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3273 ));
NOR2_X2 \GFM/U766  ( .A1(\GFM/n24500 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3271 ));
NOR2_X2 \GFM/U765  ( .A1(\GFM/n24401 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3304 ));
NOR2_X2 \GFM/U764  ( .A1(\GFM/n24290 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3303 ));
NOR2_X2 \GFM/U763  ( .A1(\GFM/n24390 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3336 ));
NOR2_X2 \GFM/U762  ( .A1(\GFM/n24290 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3335 ));
NOR2_X2 \GFM/U761  ( .A1(\GFM/n24390 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3369 ));
NOR2_X2 \GFM/U760  ( .A1(\GFM/n24290 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3368 ));
NOR2_X2 \GFM/U759  ( .A1(\GFM/n25101 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3469 ));
NOR2_X2 \GFM/U758  ( .A1(\GFM/n2489 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3467 ));
NOR2_X2 \GFM/U757  ( .A1(\GFM/n2479 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3509 ));
NOR2_X2 \GFM/U756  ( .A1(\GFM/n2489 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3508 ));
NOR2_X2 \GFM/U754  ( .A1(\GFM/n2479 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3552 ));
NOR2_X2 \GFM/U753  ( .A1(\GFM/n2489 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3551 ));
NOR2_X2 \GFM/U752  ( .A1(\GFM/n2479 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3598 ));
NOR2_X2 \GFM/U751  ( .A1(\GFM/n2489 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3597 ));
NOR2_X2 \GFM/U750  ( .A1(\GFM/n25201 ), .A2(\GFM/n25840 ), .ZN(\GFM/N283 ));
NOR2_X2 \GFM/U749  ( .A1(\GFM/n2458 ), .A2(\GFM/n25800 ), .ZN(\GFM/N51 ) );
NOR2_X2 \GFM/U748  ( .A1(\GFM/n25660 ), .A2(\GFM/n2516 ), .ZN(\GFM/N66 ) );
NOR2_X2 \GFM/U747  ( .A1(\GFM/n25880 ), .A2(\GFM/n24960 ), .ZN(\GFM/N317 ));
NOR2_X2 \GFM/U746  ( .A1(\GFM/n24280 ), .A2(\GFM/n2586 ), .ZN(\GFM/N49 ) );
NOR2_X2 \GFM/U745  ( .A1(\GFM/n2448 ), .A2(\GFM/n25821 ), .ZN(\GFM/N47 ) );
NOR2_X2 \GFM/U744  ( .A1(\GFM/n2455 ), .A2(\GFM/n2586 ), .ZN(\GFM/N109 ) );
NOR2_X2 \GFM/U743  ( .A1(\GFM/n25880 ), .A2(\GFM/n24260 ), .ZN(\GFM/N111 ));
NOR2_X2 \GFM/U742  ( .A1(\GFM/n25890 ), .A2(\GFM/n24960 ), .ZN(\GFM/N348 ));
NOR2_X2 \GFM/U741  ( .A1(\GFM/n25880 ), .A2(\GFM/n2516 ), .ZN(\GFM/N376 ) );
NOR2_X2 \GFM/U740  ( .A1(\GFM/n2455 ), .A2(\GFM/n2587 ), .ZN(\GFM/N140 ) );
NOR2_X2 \GFM/U739  ( .A1(\GFM/n25890 ), .A2(\GFM/n24260 ), .ZN(\GFM/N142 ));
NOR2_X2 \GFM/U738  ( .A1(\GFM/n24340 ), .A2(\GFM/n25901 ), .ZN(\GFM/N173 ));
NOR2_X2 \GFM/U736  ( .A1(\GFM/n25880 ), .A2(\GFM/n24460 ), .ZN(\GFM/N171 ));
INV_X4 \GFM/U735  ( .A(b_in[127]), .ZN(\GFM/n25360 ) );
INV_X4 \GFM/U734  ( .A(b_in[125]), .ZN(\GFM/n2516 ) );
INV_X4 \GFM/U733  ( .A(b_in[116]), .ZN(\GFM/n24260 ) );
INV_X4 \GFM/U732  ( .A(b_in[126]), .ZN(\GFM/n25260 ) );
NOR2_X2 \GFM/U731  ( .A1(\GFM/n25380 ), .A2(\GFM/n2699 ), .ZN(\GFM/N4322 ));
NOR2_X2 \GFM/U730  ( .A1(\GFM/n2696 ), .A2(\GFM/n25360 ), .ZN(\GFM/N4102 ));
NOR2_X2 \GFM/U729  ( .A1(\GFM/n2697 ), .A2(\GFM/n25360 ), .ZN(\GFM/N4159 ));
NOR2_X2 \GFM/U728  ( .A1(\GFM/n2696 ), .A2(\GFM/n2516 ), .ZN(\GFM/N3996 ) );
NOR2_X2 \GFM/U727  ( .A1(\GFM/n25390 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3287 ));
NOR2_X2 \GFM/U726  ( .A1(\GFM/n25390 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3319 ));
NOR2_X2 \GFM/U725  ( .A1(\GFM/n25390 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3352 ));
NOR2_X2 \GFM/U724  ( .A1(\GFM/n25390 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3386 ));
NOR2_X2 \GFM/U723  ( .A1(\GFM/n25390 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3422 ));
NOR2_X2 \GFM/U722  ( .A1(\GFM/n25390 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3460 ));
NOR2_X2 \GFM/U721  ( .A1(\GFM/n25390 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3500 ));
NOR2_X2 \GFM/U720  ( .A1(\GFM/n25390 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3543 ));
NOR2_X2 \GFM/U719  ( .A1(\GFM/n25390 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3589 ));
NOR2_X2 \GFM/U718  ( .A1(\GFM/n2540 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3638 ) );
NOR2_X2 \GFM/U716  ( .A1(\GFM/n25380 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3690 ));
NOR2_X2 \GFM/U715  ( .A1(\GFM/n25380 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3803 ));
NOR2_X2 \GFM/U714  ( .A1(\GFM/n25380 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3864 ));
NOR2_X2 \GFM/U713  ( .A1(\GFM/n2697 ), .A2(\GFM/n25270 ), .ZN(\GFM/N4103 ));
NOR2_X2 \GFM/U712  ( .A1(\GFM/n2479 ), .A2(\GFM/n25500 ), .ZN(\GFM/N4004 ));
NOR2_X2 \GFM/U711  ( .A1(\GFM/n21360 ), .A2(\GFM/n24870 ), .ZN(\GFM/N4006 ));
NOR2_X2 \GFM/U710  ( .A1(\GFM/n25310 ), .A2(\GFM/n26070 ), .ZN(\GFM/N995 ));
NOR2_X2 \GFM/U709  ( .A1(\GFM/n2541 ), .A2(\GFM/n2606 ), .ZN(\GFM/N993 ) );
NOR2_X2 \GFM/U708  ( .A1(\GFM/n23910 ), .A2(\GFM/n26200 ), .ZN(\GFM/N989 ));
NOR2_X2 \GFM/U707  ( .A1(\GFM/n25350 ), .A2(\GFM/n26200 ), .ZN(\GFM/N1398 ));
NOR2_X2 \GFM/U706  ( .A1(\GFM/n25450 ), .A2(\GFM/n26190 ), .ZN(\GFM/N1396 ));
NOR2_X2 \GFM/U705  ( .A1(\GFM/n2389 ), .A2(\GFM/n26190 ), .ZN(\GFM/N958 ) );
NOR2_X2 \GFM/U704  ( .A1(\GFM/n23880 ), .A2(\GFM/n2617 ), .ZN(\GFM/N896 ) );
NOR2_X2 \GFM/U703  ( .A1(\GFM/n25350 ), .A2(\GFM/n2617 ), .ZN(\GFM/N1305 ));
NOR2_X2 \GFM/U702  ( .A1(\GFM/n25450 ), .A2(\GFM/n2616 ), .ZN(\GFM/N1303 ));
NOR2_X2 \GFM/U701  ( .A1(\GFM/n23880 ), .A2(\GFM/n26120 ), .ZN(\GFM/N741 ));
NOR2_X2 \GFM/U700  ( .A1(\GFM/n25350 ), .A2(\GFM/n26120 ), .ZN(\GFM/N1150 ));
NOR2_X2 \GFM/U698  ( .A1(\GFM/n25450 ), .A2(\GFM/n26110 ), .ZN(\GFM/N1148 ));
NOR2_X2 \GFM/U697  ( .A1(\GFM/n23880 ), .A2(\GFM/n2613 ), .ZN(\GFM/N772 ) );
NOR2_X2 \GFM/U696  ( .A1(\GFM/n23880 ), .A2(\GFM/n2616 ), .ZN(\GFM/N865 ) );
NOR2_X2 \GFM/U695  ( .A1(\GFM/n25350 ), .A2(\GFM/n2616 ), .ZN(\GFM/N1274 ));
NOR2_X2 \GFM/U694  ( .A1(\GFM/n25450 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1272 ));
NOR2_X2 \GFM/U693  ( .A1(\GFM/n23880 ), .A2(\GFM/n26140 ), .ZN(\GFM/N803 ));
NOR2_X2 \GFM/U692  ( .A1(\GFM/n26980 ), .A2(\GFM/n25260 ), .ZN(\GFM/N4160 ));
NOR2_X2 \GFM/U691  ( .A1(\GFM/n2389 ), .A2(\GFM/n26150 ), .ZN(\GFM/N834 ) );
NOR2_X2 \GFM/U690  ( .A1(\GFM/n25350 ), .A2(\GFM/n26150 ), .ZN(\GFM/N1243 ));
NOR2_X2 \GFM/U689  ( .A1(\GFM/n25450 ), .A2(\GFM/n26140 ), .ZN(\GFM/N1241 ));
NOR2_X2 \GFM/U688  ( .A1(\GFM/n23880 ), .A2(\GFM/n26110 ), .ZN(\GFM/N710 ));
NOR2_X2 \GFM/U687  ( .A1(\GFM/n23880 ), .A2(\GFM/n25901 ), .ZN(\GFM/N59 ) );
NOR2_X2 \GFM/U686  ( .A1(\GFM/n23880 ), .A2(\GFM/n25910 ), .ZN(\GFM/N90 ) );
NOR2_X2 \GFM/U685  ( .A1(\GFM/n23950 ), .A2(\GFM/n25930 ), .ZN(\GFM/N152 ));
NOR2_X2 \GFM/U684  ( .A1(\GFM/n23940 ), .A2(\GFM/n25940 ), .ZN(\GFM/N183 ));
NOR2_X2 \GFM/U683  ( .A1(\GFM/n2393 ), .A2(\GFM/n2595 ), .ZN(\GFM/N214 ) );
NOR2_X2 \GFM/U682  ( .A1(\GFM/n2392 ), .A2(\GFM/n2596 ), .ZN(\GFM/N245 ) );
NOR2_X2 \GFM/U681  ( .A1(\GFM/n2528 ), .A2(\GFM/n25901 ), .ZN(\GFM/N468 ) );
NOR2_X2 \GFM/U680  ( .A1(\GFM/n25890 ), .A2(\GFM/n25360 ), .ZN(\GFM/N466 ));
NOR2_X2 \GFM/U678  ( .A1(\GFM/n23880 ), .A2(\GFM/n26050 ), .ZN(\GFM/N524 ));
NOR2_X2 \GFM/U677  ( .A1(\GFM/n25270 ), .A2(\GFM/n25910 ), .ZN(\GFM/N499 ));
NOR2_X2 \GFM/U676  ( .A1(\GFM/n25380 ), .A2(\GFM/n25901 ), .ZN(\GFM/N497 ));
NOR2_X2 \GFM/U675  ( .A1(\GFM/n2528 ), .A2(\GFM/n2592 ), .ZN(\GFM/N530 ) );
NOR2_X2 \GFM/U674  ( .A1(\GFM/n25380 ), .A2(\GFM/n25910 ), .ZN(\GFM/N528 ));
NOR2_X2 \GFM/U673  ( .A1(\GFM/n2528 ), .A2(\GFM/n25930 ), .ZN(\GFM/N561 ) );
NOR2_X2 \GFM/U672  ( .A1(\GFM/n2537 ), .A2(\GFM/n2592 ), .ZN(\GFM/N559 ) );
NOR2_X2 \GFM/U671  ( .A1(\GFM/n2528 ), .A2(\GFM/n25940 ), .ZN(\GFM/N592 ) );
NOR2_X2 \GFM/U670  ( .A1(\GFM/n25380 ), .A2(\GFM/n25930 ), .ZN(\GFM/N590 ));
NOR2_X2 \GFM/U669  ( .A1(\GFM/n23880 ), .A2(\GFM/n2609 ), .ZN(\GFM/N648 ) );
NOR2_X2 \GFM/U668  ( .A1(\GFM/n25270 ), .A2(\GFM/n2595 ), .ZN(\GFM/N623 ) );
NOR2_X2 \GFM/U667  ( .A1(\GFM/n25380 ), .A2(\GFM/n25940 ), .ZN(\GFM/N621 ));
NOR2_X2 \GFM/U666  ( .A1(\GFM/n25270 ), .A2(\GFM/n2596 ), .ZN(\GFM/N654 ) );
NOR2_X2 \GFM/U665  ( .A1(\GFM/n2537 ), .A2(\GFM/n2595 ), .ZN(\GFM/N652 ) );
NOR2_X2 \GFM/U664  ( .A1(\GFM/n2528 ), .A2(\GFM/n25970 ), .ZN(\GFM/N685 ) );
NOR2_X2 \GFM/U663  ( .A1(\GFM/n2537 ), .A2(\GFM/n2596 ), .ZN(\GFM/N683 ) );
NOR2_X2 \GFM/U662  ( .A1(\GFM/n25270 ), .A2(\GFM/n25980 ), .ZN(\GFM/N716 ));
NOR2_X2 \GFM/U661  ( .A1(\GFM/n2537 ), .A2(\GFM/n25970 ), .ZN(\GFM/N714 ) );
NOR2_X2 \GFM/U660  ( .A1(\GFM/n25270 ), .A2(\GFM/n2599 ), .ZN(\GFM/N747 ) );
NOR2_X2 \GFM/U659  ( .A1(\GFM/n25380 ), .A2(\GFM/n25980 ), .ZN(\GFM/N745 ));
NOR2_X2 \GFM/U658  ( .A1(\GFM/n25270 ), .A2(\GFM/n26000 ), .ZN(\GFM/N778 ));
NOR2_X2 \GFM/U657  ( .A1(\GFM/n2537 ), .A2(\GFM/n2599 ), .ZN(\GFM/N776 ) );
NOR2_X2 \GFM/U656  ( .A1(\GFM/n25270 ), .A2(\GFM/n26010 ), .ZN(\GFM/N809 ));
NOR2_X2 \GFM/U655  ( .A1(\GFM/n25390 ), .A2(\GFM/n26000 ), .ZN(\GFM/N807 ));
NOR2_X2 \GFM/U654  ( .A1(\GFM/n2528 ), .A2(\GFM/n2602 ), .ZN(\GFM/N840 ) );
NOR2_X2 \GFM/U653  ( .A1(\GFM/n2537 ), .A2(\GFM/n26010 ), .ZN(\GFM/N838 ) );
NOR2_X2 \GFM/U652  ( .A1(\GFM/n25270 ), .A2(\GFM/n2603 ), .ZN(\GFM/N871 ) );
NOR2_X2 \GFM/U651  ( .A1(\GFM/n2537 ), .A2(\GFM/n2602 ), .ZN(\GFM/N869 ) );
NOR2_X2 \GFM/U650  ( .A1(\GFM/n25270 ), .A2(\GFM/n2604 ), .ZN(\GFM/N902 ) );
NOR2_X2 \GFM/U649  ( .A1(\GFM/n2537 ), .A2(\GFM/n2603 ), .ZN(\GFM/N900 ) );
NOR2_X2 \GFM/U648  ( .A1(\GFM/n25270 ), .A2(\GFM/n26050 ), .ZN(\GFM/N933 ));
NOR2_X2 \GFM/U647  ( .A1(\GFM/n2537 ), .A2(\GFM/n2604 ), .ZN(\GFM/N931 ) );
NOR2_X2 \GFM/U646  ( .A1(\GFM/n25270 ), .A2(\GFM/n2609 ), .ZN(\GFM/N1057 ));
NOR2_X2 \GFM/U645  ( .A1(\GFM/n26080 ), .A2(\GFM/n25360 ), .ZN(\GFM/N1055 ));
NOR2_X2 \GFM/U644  ( .A1(\GFM/n23950 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1299 ));
NOR2_X2 \GFM/U643  ( .A1(\GFM/n23950 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1330 ));
NOR2_X2 \GFM/U642  ( .A1(\GFM/n23950 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1361 ));
NOR2_X2 \GFM/U641  ( .A1(\GFM/n23950 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1392 ));
NOR2_X2 \GFM/U640  ( .A1(\GFM/n23950 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1423 ));
NOR2_X2 \GFM/U639  ( .A1(\GFM/n23950 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1454 ));
NOR2_X2 \GFM/U638  ( .A1(\GFM/n2534 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1429 ) );
NOR2_X2 \GFM/U637  ( .A1(\GFM/n25450 ), .A2(\GFM/n26200 ), .ZN(\GFM/N1427 ));
NOR2_X2 \GFM/U636  ( .A1(\GFM/n23950 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1485 ));
NOR2_X2 \GFM/U635  ( .A1(\GFM/n2534 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1460 ));
NOR2_X2 \GFM/U634  ( .A1(\GFM/n2544 ), .A2(\GFM/n2621 ), .ZN(\GFM/N1458 ) );
NOR2_X2 \GFM/U633  ( .A1(\GFM/n23950 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1516 ));
NOR2_X2 \GFM/U632  ( .A1(\GFM/n2534 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1491 ) );
NOR2_X2 \GFM/U631  ( .A1(\GFM/n2544 ), .A2(\GFM/n26220 ), .ZN(\GFM/N1489 ));
NOR2_X2 \GFM/U630  ( .A1(\GFM/n23950 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1547 ));
NOR2_X2 \GFM/U629  ( .A1(\GFM/n2534 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1522 ));
NOR2_X2 \GFM/U628  ( .A1(\GFM/n2544 ), .A2(\GFM/n2623 ), .ZN(\GFM/N1520 ) );
NOR2_X2 \GFM/U627  ( .A1(\GFM/n23950 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1578 ));
NOR2_X2 \GFM/U626  ( .A1(\GFM/n2534 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1553 ));
NOR2_X2 \GFM/U625  ( .A1(\GFM/n2544 ), .A2(\GFM/n26240 ), .ZN(\GFM/N1551 ));
NOR2_X2 \GFM/U624  ( .A1(\GFM/n23950 ), .A2(\GFM/n26401 ), .ZN(\GFM/N1609 ));
NOR2_X2 \GFM/U623  ( .A1(\GFM/n2534 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1584 ) );
NOR2_X2 \GFM/U622  ( .A1(\GFM/n2544 ), .A2(\GFM/n26250 ), .ZN(\GFM/N1582 ));
NOR2_X2 \GFM/U621  ( .A1(\GFM/n23950 ), .A2(\GFM/n2641 ), .ZN(\GFM/N1640 ));
NOR2_X2 \GFM/U620  ( .A1(\GFM/n2534 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1615 ) );
NOR2_X2 \GFM/U619  ( .A1(\GFM/n2544 ), .A2(\GFM/n2626 ), .ZN(\GFM/N1613 ) );
NOR2_X2 \GFM/U618  ( .A1(\GFM/n23940 ), .A2(\GFM/n26420 ), .ZN(\GFM/N1671 ));
NOR2_X2 \GFM/U617  ( .A1(\GFM/n2534 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1646 ));
NOR2_X2 \GFM/U616  ( .A1(\GFM/n2544 ), .A2(\GFM/n2627 ), .ZN(\GFM/N1644 ) );
NOR2_X2 \GFM/U615  ( .A1(\GFM/n23940 ), .A2(\GFM/n26430 ), .ZN(\GFM/N1702 ));
NOR2_X2 \GFM/U614  ( .A1(\GFM/n2534 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1677 ));
NOR2_X2 \GFM/U613  ( .A1(\GFM/n2544 ), .A2(\GFM/n26280 ), .ZN(\GFM/N1675 ));
NOR2_X2 \GFM/U612  ( .A1(\GFM/n23940 ), .A2(\GFM/n2644 ), .ZN(\GFM/N1733 ));
NOR2_X2 \GFM/U611  ( .A1(\GFM/n2534 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1708 ));
NOR2_X2 \GFM/U610  ( .A1(\GFM/n2544 ), .A2(\GFM/n26290 ), .ZN(\GFM/N1706 ));
NOR2_X2 \GFM/U609  ( .A1(\GFM/n23940 ), .A2(\GFM/n26450 ), .ZN(\GFM/N1764 ));
NOR2_X2 \GFM/U608  ( .A1(\GFM/n2534 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1739 ));
NOR2_X2 \GFM/U607  ( .A1(\GFM/n2544 ), .A2(\GFM/n26301 ), .ZN(\GFM/N1737 ));
NOR2_X2 \GFM/U606  ( .A1(\GFM/n23940 ), .A2(\GFM/n26460 ), .ZN(\GFM/N1795 ));
NOR2_X2 \GFM/U605  ( .A1(\GFM/n2534 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1770 ));
NOR2_X2 \GFM/U604  ( .A1(\GFM/n2544 ), .A2(\GFM/n26310 ), .ZN(\GFM/N1768 ));
NOR2_X2 \GFM/U603  ( .A1(\GFM/n23940 ), .A2(\GFM/n2647 ), .ZN(\GFM/N1826 ));
NOR2_X2 \GFM/U602  ( .A1(\GFM/n2533 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1801 ) );
NOR2_X2 \GFM/U601  ( .A1(\GFM/n2544 ), .A2(\GFM/n26320 ), .ZN(\GFM/N1799 ));
NOR2_X2 \GFM/U600  ( .A1(\GFM/n23940 ), .A2(\GFM/n2648 ), .ZN(\GFM/N1857 ));
NOR2_X2 \GFM/U599  ( .A1(\GFM/n2533 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1832 ) );
NOR2_X2 \GFM/U598  ( .A1(\GFM/n25430 ), .A2(\GFM/n2633 ), .ZN(\GFM/N1830 ));
NOR2_X2 \GFM/U597  ( .A1(\GFM/n23940 ), .A2(\GFM/n2649 ), .ZN(\GFM/N1888 ));
NOR2_X2 \GFM/U596  ( .A1(\GFM/n2533 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1863 ) );
NOR2_X2 \GFM/U595  ( .A1(\GFM/n25430 ), .A2(\GFM/n2634 ), .ZN(\GFM/N1861 ));
NOR2_X2 \GFM/U594  ( .A1(\GFM/n23940 ), .A2(\GFM/n26500 ), .ZN(\GFM/N1919 ));
NOR2_X2 \GFM/U593  ( .A1(\GFM/n2533 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1894 ));
NOR2_X2 \GFM/U592  ( .A1(\GFM/n25430 ), .A2(\GFM/n2635 ), .ZN(\GFM/N1892 ));
NOR2_X2 \GFM/U591  ( .A1(\GFM/n23940 ), .A2(\GFM/n26510 ), .ZN(\GFM/N1950 ));
NOR2_X2 \GFM/U590  ( .A1(\GFM/n2533 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1925 ) );
NOR2_X2 \GFM/U589  ( .A1(\GFM/n25430 ), .A2(\GFM/n26360 ), .ZN(\GFM/N1923 ));
NOR2_X2 \GFM/U588  ( .A1(\GFM/n23940 ), .A2(\GFM/n2652 ), .ZN(\GFM/N1981 ));
NOR2_X2 \GFM/U587  ( .A1(\GFM/n2533 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1956 ));
NOR2_X2 \GFM/U586  ( .A1(\GFM/n25430 ), .A2(\GFM/n2637 ), .ZN(\GFM/N1954 ));
NOR2_X2 \GFM/U585  ( .A1(\GFM/n23940 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2012 ));
NOR2_X2 \GFM/U584  ( .A1(\GFM/n2533 ), .A2(\GFM/n26390 ), .ZN(\GFM/N1987 ));
NOR2_X2 \GFM/U583  ( .A1(\GFM/n25430 ), .A2(\GFM/n26380 ), .ZN(\GFM/N1985 ));
NOR2_X2 \GFM/U582  ( .A1(\GFM/n2393 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2043 ) );
NOR2_X2 \GFM/U581  ( .A1(\GFM/n2533 ), .A2(\GFM/n26401 ), .ZN(\GFM/N2018 ));
NOR2_X2 \GFM/U580  ( .A1(\GFM/n25430 ), .A2(\GFM/n26390 ), .ZN(\GFM/N2016 ));
NOR2_X2 \GFM/U579  ( .A1(\GFM/n2393 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2074 ));
NOR2_X2 \GFM/U578  ( .A1(\GFM/n2533 ), .A2(\GFM/n2641 ), .ZN(\GFM/N2049 ) );
NOR2_X2 \GFM/U577  ( .A1(\GFM/n25430 ), .A2(\GFM/n26401 ), .ZN(\GFM/N2047 ));
NOR2_X2 \GFM/U576  ( .A1(\GFM/n2393 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2105 ));
NOR2_X2 \GFM/U575  ( .A1(\GFM/n2533 ), .A2(\GFM/n26420 ), .ZN(\GFM/N2080 ));
NOR2_X2 \GFM/U574  ( .A1(\GFM/n25430 ), .A2(\GFM/n2641 ), .ZN(\GFM/N2078 ));
NOR2_X2 \GFM/U573  ( .A1(\GFM/n2393 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2136 ) );
NOR2_X2 \GFM/U572  ( .A1(\GFM/n2533 ), .A2(\GFM/n26430 ), .ZN(\GFM/N2111 ));
NOR2_X2 \GFM/U571  ( .A1(\GFM/n25430 ), .A2(\GFM/n26420 ), .ZN(\GFM/N2109 ));
NOR2_X2 \GFM/U570  ( .A1(\GFM/n2393 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2167 ) );
NOR2_X2 \GFM/U569  ( .A1(\GFM/n2533 ), .A2(\GFM/n2644 ), .ZN(\GFM/N2142 ) );
NOR2_X2 \GFM/U568  ( .A1(\GFM/n25430 ), .A2(\GFM/n26430 ), .ZN(\GFM/N2140 ));
NOR2_X2 \GFM/U567  ( .A1(\GFM/n2393 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2198 ));
NOR2_X2 \GFM/U566  ( .A1(\GFM/n25320 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2173 ));
NOR2_X2 \GFM/U565  ( .A1(\GFM/n25430 ), .A2(\GFM/n2644 ), .ZN(\GFM/N2171 ));
NOR2_X2 \GFM/U564  ( .A1(\GFM/n2393 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2229 ));
NOR2_X2 \GFM/U563  ( .A1(\GFM/n25320 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2204 ));
NOR2_X2 \GFM/U562  ( .A1(\GFM/n2542 ), .A2(\GFM/n26450 ), .ZN(\GFM/N2202 ));
NOR2_X2 \GFM/U561  ( .A1(\GFM/n2393 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2260 ));
NOR2_X2 \GFM/U560  ( .A1(\GFM/n25320 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2235 ));
NOR2_X2 \GFM/U559  ( .A1(\GFM/n2542 ), .A2(\GFM/n26460 ), .ZN(\GFM/N2233 ));
NOR2_X2 \GFM/U558  ( .A1(\GFM/n2393 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2291 ));
NOR2_X2 \GFM/U557  ( .A1(\GFM/n25320 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2266 ));
NOR2_X2 \GFM/U556  ( .A1(\GFM/n2542 ), .A2(\GFM/n2647 ), .ZN(\GFM/N2264 ) );
NOR2_X2 \GFM/U555  ( .A1(\GFM/n2393 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2322 ));
NOR2_X2 \GFM/U554  ( .A1(\GFM/n25320 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2297 ));
NOR2_X2 \GFM/U553  ( .A1(\GFM/n2542 ), .A2(\GFM/n2648 ), .ZN(\GFM/N2295 ) );
NOR2_X2 \GFM/U552  ( .A1(\GFM/n2393 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2353 ) );
NOR2_X2 \GFM/U551  ( .A1(\GFM/n25320 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2328 ));
NOR2_X2 \GFM/U550  ( .A1(\GFM/n2542 ), .A2(\GFM/n2649 ), .ZN(\GFM/N2326 ) );
NOR2_X2 \GFM/U549  ( .A1(\GFM/n2393 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2384 ) );
NOR2_X2 \GFM/U548  ( .A1(\GFM/n25320 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2359 ));
NOR2_X2 \GFM/U547  ( .A1(\GFM/n2542 ), .A2(\GFM/n26500 ), .ZN(\GFM/N2357 ));
NOR2_X2 \GFM/U546  ( .A1(\GFM/n2392 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2415 ) );
NOR2_X2 \GFM/U545  ( .A1(\GFM/n25320 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2390 ));
NOR2_X2 \GFM/U544  ( .A1(\GFM/n2542 ), .A2(\GFM/n26510 ), .ZN(\GFM/N2388 ));
NOR2_X2 \GFM/U543  ( .A1(\GFM/n2392 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2446 ));
NOR2_X2 \GFM/U542  ( .A1(\GFM/n25320 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2421 ));
NOR2_X2 \GFM/U541  ( .A1(\GFM/n2542 ), .A2(\GFM/n2652 ), .ZN(\GFM/N2419 ) );
NOR2_X2 \GFM/U540  ( .A1(\GFM/n2392 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2477 ) );
NOR2_X2 \GFM/U539  ( .A1(\GFM/n25320 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2452 ));
NOR2_X2 \GFM/U538  ( .A1(\GFM/n2542 ), .A2(\GFM/n26530 ), .ZN(\GFM/N2450 ));
NOR2_X2 \GFM/U537  ( .A1(\GFM/n2392 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2508 ));
NOR2_X2 \GFM/U536  ( .A1(\GFM/n25320 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2483 ));
NOR2_X2 \GFM/U535  ( .A1(\GFM/n2542 ), .A2(\GFM/n2654 ), .ZN(\GFM/N2481 ) );
NOR2_X2 \GFM/U534  ( .A1(\GFM/n2392 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2539 ));
NOR2_X2 \GFM/U533  ( .A1(\GFM/n25310 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2514 ));
NOR2_X2 \GFM/U532  ( .A1(\GFM/n2542 ), .A2(\GFM/n26550 ), .ZN(\GFM/N2512 ));
NOR2_X2 \GFM/U531  ( .A1(\GFM/n2392 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2570 ) );
NOR2_X2 \GFM/U530  ( .A1(\GFM/n25310 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2545 ));
NOR2_X2 \GFM/U529  ( .A1(\GFM/n2541 ), .A2(\GFM/n26560 ), .ZN(\GFM/N2543 ));
NOR2_X2 \GFM/U528  ( .A1(\GFM/n25310 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2576 ));
NOR2_X2 \GFM/U527  ( .A1(\GFM/n2541 ), .A2(\GFM/n2657 ), .ZN(\GFM/N2574 ) );
NOR2_X2 \GFM/U526  ( .A1(\GFM/n25310 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2607 ));
NOR2_X2 \GFM/U525  ( .A1(\GFM/n2541 ), .A2(\GFM/n2658 ), .ZN(\GFM/N2605 ) );
NOR2_X2 \GFM/U524  ( .A1(\GFM/n25310 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2638 ));
NOR2_X2 \GFM/U523  ( .A1(\GFM/n2541 ), .A2(\GFM/n26590 ), .ZN(\GFM/N2636 ));
NOR2_X2 \GFM/U522  ( .A1(\GFM/n25310 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2669 ));
NOR2_X2 \GFM/U521  ( .A1(\GFM/n2541 ), .A2(\GFM/n26600 ), .ZN(\GFM/N2667 ));
NOR2_X2 \GFM/U520  ( .A1(\GFM/n25310 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2700 ));
NOR2_X2 \GFM/U519  ( .A1(\GFM/n2541 ), .A2(\GFM/n26611 ), .ZN(\GFM/N2698 ));
NOR2_X2 \GFM/U518  ( .A1(\GFM/n25310 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2731 ));
NOR2_X2 \GFM/U517  ( .A1(\GFM/n2541 ), .A2(\GFM/n26620 ), .ZN(\GFM/N2729 ));
NOR2_X2 \GFM/U516  ( .A1(\GFM/n25310 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2762 ));
NOR2_X2 \GFM/U515  ( .A1(\GFM/n2541 ), .A2(\GFM/n26630 ), .ZN(\GFM/N2760 ));
NOR2_X2 \GFM/U514  ( .A1(\GFM/n25310 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2793 ));
NOR2_X2 \GFM/U513  ( .A1(\GFM/n2541 ), .A2(\GFM/n2664 ), .ZN(\GFM/N2791 ) );
NOR2_X2 \GFM/U512  ( .A1(\GFM/n25310 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2824 ));
NOR2_X2 \GFM/U511  ( .A1(\GFM/n2541 ), .A2(\GFM/n2665 ), .ZN(\GFM/N2822 ) );
NOR2_X2 \GFM/U510  ( .A1(\GFM/n2530 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2855 ));
NOR2_X2 \GFM/U509  ( .A1(\GFM/n2541 ), .A2(\GFM/n2666 ), .ZN(\GFM/N2853 ) );
NOR2_X2 \GFM/U508  ( .A1(\GFM/n2530 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2886 ) );
NOR2_X2 \GFM/U507  ( .A1(\GFM/n2540 ), .A2(\GFM/n26670 ), .ZN(\GFM/N2884 ));
NOR2_X2 \GFM/U506  ( .A1(\GFM/n2530 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2917 ));
NOR2_X2 \GFM/U505  ( .A1(\GFM/n2540 ), .A2(\GFM/n2668 ), .ZN(\GFM/N2915 ) );
NOR2_X2 \GFM/U504  ( .A1(\GFM/n2530 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2948 ));
NOR2_X2 \GFM/U503  ( .A1(\GFM/n2540 ), .A2(\GFM/n26690 ), .ZN(\GFM/N2946 ));
NOR2_X2 \GFM/U502  ( .A1(\GFM/n2530 ), .A2(\GFM/n2671 ), .ZN(\GFM/N2979 ) );
NOR2_X2 \GFM/U501  ( .A1(\GFM/n2540 ), .A2(\GFM/n26700 ), .ZN(\GFM/N2977 ));
NOR2_X2 \GFM/U500  ( .A1(\GFM/n2392 ), .A2(\GFM/n2672 ), .ZN(\GFM/N2601 ) );
NOR2_X2 \GFM/U499  ( .A1(\GFM/n2392 ), .A2(\GFM/n26730 ), .ZN(\GFM/N2632 ));
NOR2_X2 \GFM/U498  ( .A1(\GFM/n2392 ), .A2(\GFM/n26740 ), .ZN(\GFM/N2663 ));
NOR2_X2 \GFM/U497  ( .A1(\GFM/n2392 ), .A2(\GFM/n2675 ), .ZN(\GFM/N2694 ) );
NOR2_X2 \GFM/U496  ( .A1(\GFM/n2392 ), .A2(\GFM/n26760 ), .ZN(\GFM/N2725 ));
NOR2_X2 \GFM/U495  ( .A1(\GFM/n2392 ), .A2(\GFM/n26770 ), .ZN(\GFM/N2756 ));
NOR2_X2 \GFM/U494  ( .A1(\GFM/n23910 ), .A2(\GFM/n2678 ), .ZN(\GFM/N2787 ));
NOR2_X2 \GFM/U493  ( .A1(\GFM/n23910 ), .A2(\GFM/n2679 ), .ZN(\GFM/N2818 ));
NOR2_X2 \GFM/U492  ( .A1(\GFM/n23910 ), .A2(\GFM/n26801 ), .ZN(\GFM/N2849 ));
NOR2_X2 \GFM/U491  ( .A1(\GFM/n23910 ), .A2(\GFM/n26810 ), .ZN(\GFM/N2880 ));
NOR2_X2 \GFM/U490  ( .A1(\GFM/n23910 ), .A2(\GFM/n26820 ), .ZN(\GFM/N2911 ));
NOR2_X2 \GFM/U489  ( .A1(\GFM/n23910 ), .A2(\GFM/n2683 ), .ZN(\GFM/N2942 ));
NOR2_X2 \GFM/U488  ( .A1(\GFM/n23910 ), .A2(\GFM/n26840 ), .ZN(\GFM/N2973 ));
NOR2_X2 \GFM/U485  ( .A1(\GFM/n23910 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3004 ));
NOR2_X2 \GFM/U484  ( .A1(\GFM/n23910 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3035 ));
NOR2_X2 \GFM/U483  ( .A1(\GFM/n23910 ), .A2(\GFM/n26870 ), .ZN(\GFM/N3066 ));
NOR2_X2 \GFM/U482  ( .A1(\GFM/n23900 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3097 ));
NOR2_X2 \GFM/U481  ( .A1(\GFM/n23900 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3128 ));
NOR2_X2 \GFM/U480  ( .A1(\GFM/n23900 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3159 ));
NOR2_X2 \GFM/U478  ( .A1(\GFM/n23900 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3190 ));
NOR2_X2 \GFM/U477  ( .A1(\GFM/n23900 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3221 ));
NOR2_X2 \GFM/U476  ( .A1(\GFM/n23900 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3252 ));
NOR2_X2 \GFM/U475  ( .A1(\GFM/n23900 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3283 ));
NOR2_X2 \GFM/U474  ( .A1(\GFM/n25290 ), .A2(\GFM/n26810 ), .ZN(\GFM/N3289 ));
NOR2_X2 \GFM/U473  ( .A1(\GFM/n25290 ), .A2(\GFM/n26820 ), .ZN(\GFM/N3321 ));
NOR2_X2 \GFM/U472  ( .A1(\GFM/n25290 ), .A2(\GFM/n2683 ), .ZN(\GFM/N3354 ));
NOR2_X2 \GFM/U471  ( .A1(\GFM/n25290 ), .A2(\GFM/n26840 ), .ZN(\GFM/N3388 ));
NOR2_X2 \GFM/U470  ( .A1(\GFM/n25290 ), .A2(\GFM/n2685 ), .ZN(\GFM/N3424 ));
NOR2_X2 \GFM/U469  ( .A1(\GFM/n25290 ), .A2(\GFM/n26860 ), .ZN(\GFM/N3462 ));
NOR2_X2 \GFM/U468  ( .A1(\GFM/n25190 ), .A2(\GFM/n2688 ), .ZN(\GFM/N3502 ));
NOR2_X2 \GFM/U467  ( .A1(\GFM/n25190 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3545 ));
NOR2_X2 \GFM/U466  ( .A1(\GFM/n25190 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3591 ));
NOR2_X2 \GFM/U465  ( .A1(\GFM/n25180 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3640 ));
NOR2_X2 \GFM/U464  ( .A1(\GFM/n25180 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3692 ));
NOR2_X2 \GFM/U463  ( .A1(\GFM/n2528 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3804 ));
NOR2_X2 \GFM/U462  ( .A1(\GFM/n2528 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3865 ));
NOR2_X2 \GFM/U461  ( .A1(\GFM/n26080 ), .A2(\GFM/n25260 ), .ZN(\GFM/N1026 ));
NOR2_X2 \GFM/U460  ( .A1(\GFM/n26070 ), .A2(\GFM/n25360 ), .ZN(\GFM/N1024 ));
NOR2_X2 \GFM/U459  ( .A1(\GFM/n2534 ), .A2(\GFM/n2573 ), .ZN(\GFM/N158 ) );
NOR2_X2 \GFM/U458  ( .A1(\GFM/n2544 ), .A2(\GFM/n25700 ), .ZN(\GFM/N156 ) );
NOR2_X2 \GFM/U457  ( .A1(\GFM/n25320 ), .A2(\GFM/n2578 ), .ZN(\GFM/N220 ) );
NOR2_X2 \GFM/U456  ( .A1(\GFM/n2542 ), .A2(\GFM/n25760 ), .ZN(\GFM/N218 ) );
NOR2_X2 \GFM/U455  ( .A1(\GFM/n25320 ), .A2(\GFM/n25800 ), .ZN(\GFM/N251 ));
NOR2_X2 \GFM/U454  ( .A1(\GFM/n2542 ), .A2(\GFM/n2578 ), .ZN(\GFM/N249 ) );
NOR2_X2 \GFM/U453  ( .A1(\GFM/n2530 ), .A2(\GFM/n25840 ), .ZN(\GFM/N313 ) );
NOR2_X2 \GFM/U452  ( .A1(\GFM/n2540 ), .A2(\GFM/n25821 ), .ZN(\GFM/N311 ) );
NOR2_X2 \GFM/U451  ( .A1(\GFM/n25290 ), .A2(\GFM/n2586 ), .ZN(\GFM/N344 ) );
NOR2_X2 \GFM/U450  ( .A1(\GFM/n25390 ), .A2(\GFM/n25840 ), .ZN(\GFM/N342 ));
NOR2_X2 \GFM/U449  ( .A1(\GFM/n25290 ), .A2(\GFM/n2587 ), .ZN(\GFM/N375 ) );
NOR2_X2 \GFM/U448  ( .A1(\GFM/n25380 ), .A2(\GFM/n2586 ), .ZN(\GFM/N373 ) );
NOR2_X2 \GFM/U447  ( .A1(\GFM/n2547 ), .A2(\GFM/n24770 ), .ZN(\GFM/N3647 ));
NOR2_X2 \GFM/U446  ( .A1(\GFM/n2489 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3648 ));
NOR2_X2 \GFM/U445  ( .A1(\GFM/n25890 ), .A2(\GFM/n25260 ), .ZN(\GFM/N437 ));
NOR2_X2 \GFM/U444  ( .A1(\GFM/n25880 ), .A2(\GFM/n25360 ), .ZN(\GFM/N435 ));
NOR2_X2 \GFM/U443  ( .A1(\GFM/n2554 ), .A2(\GFM/n25260 ), .ZN(\GFM/N3 ) );
NOR2_X2 \GFM/U442  ( .A1(\GFM/n25460 ), .A2(\GFM/n25360 ), .ZN(\GFM/N1 ) );
NOR2_X2 \GFM/U441  ( .A1(\GFM/n25620 ), .A2(\GFM/n25260 ), .ZN(\GFM/N65 ) );
NOR2_X2 \GFM/U440  ( .A1(\GFM/n25580 ), .A2(\GFM/n25360 ), .ZN(\GFM/N63 ) );
NOR2_X2 \GFM/U439  ( .A1(\GFM/n25660 ), .A2(\GFM/n25260 ), .ZN(\GFM/N96 ) );
NOR2_X2 \GFM/U438  ( .A1(\GFM/n25620 ), .A2(\GFM/n25360 ), .ZN(\GFM/N94 ) );
NOR2_X2 \GFM/U437  ( .A1(\GFM/n25180 ), .A2(\GFM/n2554 ), .ZN(\GFM/N4325 ));
NOR2_X2 \GFM/U436  ( .A1(\GFM/n2509 ), .A2(\GFM/n25580 ), .ZN(\GFM/N4329 ));
NOR2_X2 \GFM/U435  ( .A1(\GFM/n25290 ), .A2(\GFM/n25460 ), .ZN(\GFM/N4324 ));
NOR2_X2 \GFM/U434  ( .A1(\GFM/n23880 ), .A2(\GFM/n25880 ), .ZN(\GFM/N4349 ));
NOR2_X2 \GFM/U433  ( .A1(\GFM/n24980 ), .A2(\GFM/n25620 ), .ZN(\GFM/N4328 ));
NOR2_X2 \GFM/U432  ( .A1(\GFM/n25760 ), .A2(\GFM/n24570 ), .ZN(\GFM/N4341 ));
NOR2_X2 \GFM/U431  ( .A1(\GFM/n2578 ), .A2(\GFM/n2447 ), .ZN(\GFM/N4337 ) );
NOR2_X2 \GFM/U430  ( .A1(\GFM/n2573 ), .A2(\GFM/n24670 ), .ZN(\GFM/N4342 ));
NOR2_X2 \GFM/U429  ( .A1(\GFM/n24900 ), .A2(\GFM/n25660 ), .ZN(\GFM/N4331 ));
NOR2_X2 \GFM/U428  ( .A1(\GFM/n25800 ), .A2(\GFM/n2437 ), .ZN(\GFM/N4336 ));
NOR2_X2 \GFM/U427  ( .A1(\GFM/n25821 ), .A2(\GFM/n24260 ), .ZN(\GFM/N4339 ));
NOR2_X2 \GFM/U426  ( .A1(\GFM/n2586 ), .A2(\GFM/n24080 ), .ZN(\GFM/N4345 ));
NOR2_X2 \GFM/U425  ( .A1(\GFM/n25840 ), .A2(\GFM/n25530 ), .ZN(\GFM/N4346 ));
NOR2_X2 \GFM/U424  ( .A1(\GFM/n2587 ), .A2(\GFM/n23970 ), .ZN(\GFM/N4348 ));
NOR2_X2 \GFM/U423  ( .A1(\GFM/n21360 ), .A2(\GFM/n25070 ), .ZN(\GFM/N4108 ));
NOR2_X2 \GFM/U422  ( .A1(\GFM/n26980 ), .A2(\GFM/n2516 ), .ZN(\GFM/N4106 ));
NOR2_X2 \GFM/U421  ( .A1(\GFM/n21360 ), .A2(\GFM/n24960 ), .ZN(\GFM/N4059 ));
INV_X4 \GFM/U420  ( .A(v_out[109]), .ZN(\GFM/n25670 ) );
INV_X4 \GFM/U419  ( .A(v_out[108]), .ZN(\GFM/n25630 ) );
INV_X4 \GFM/U418  ( .A(v_out[107]), .ZN(\GFM/n2559 ) );
INV_X4 \GFM/U417  ( .A(v_out[106]), .ZN(\GFM/n2555 ) );
INV_X4 \GFM/U416  ( .A(v_out[105]), .ZN(\GFM/n2547 ) );
NOR2_X2 \GFM/U415  ( .A1(\GFM/n2696 ), .A2(\GFM/n25260 ), .ZN(\GFM/N4050 ));
NOR2_X2 \GFM/U414  ( .A1(\GFM/n24590 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3484 ));
NOR2_X2 \GFM/U413  ( .A1(\GFM/n2547 ), .A2(\GFM/n25070 ), .ZN(\GFM/N3808 ));
NOR2_X2 \GFM/U412  ( .A1(\GFM/n25180 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3809 ));
NOR2_X2 \GFM/U411  ( .A1(\GFM/n2509 ), .A2(\GFM/n25500 ), .ZN(\GFM/N4167 ));
NOR2_X2 \GFM/U410  ( .A1(\GFM/n21360 ), .A2(\GFM/n2516 ), .ZN(\GFM/N4164 ));
NOR2_X2 \GFM/U409  ( .A1(\GFM/n26980 ), .A2(\GFM/n24960 ), .ZN(\GFM/N4007 ));
NOR2_X2 \GFM/U408  ( .A1(\GFM/n24190 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3338 ));
NOR2_X2 \GFM/U407  ( .A1(\GFM/n24190 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3371 ));
NOR2_X2 \GFM/U406  ( .A1(\GFM/n2480 ), .A2(\GFM/n2689 ), .ZN(\GFM/N3397 ) );
NOR2_X2 \GFM/U405  ( .A1(\GFM/n2499 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3511 ));
NOR2_X2 \GFM/U404  ( .A1(\GFM/n2559 ), .A2(\GFM/n23970 ), .ZN(\GFM/N3413 ));
NOR2_X2 \GFM/U403  ( .A1(\GFM/n24590 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3409 ));
NOR2_X2 \GFM/U402  ( .A1(\GFM/n25630 ), .A2(\GFM/n23970 ), .ZN(\GFM/N3450 ));
NOR2_X2 \GFM/U401  ( .A1(\GFM/n24590 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3446 ));
NOR2_X2 \GFM/U400  ( .A1(\GFM/n2528 ), .A2(\GFM/n2606 ), .ZN(\GFM/N964 ) );
NOR2_X2 \GFM/U399  ( .A1(\GFM/n2537 ), .A2(\GFM/n26050 ), .ZN(\GFM/N962 ) );
NOR2_X2 \GFM/U398  ( .A1(\GFM/n2537 ), .A2(\GFM/n2609 ), .ZN(\GFM/N1086 ) );
NOR2_X2 \GFM/U397  ( .A1(\GFM/n2610 ), .A2(\GFM/n25260 ), .ZN(\GFM/N1088 ));
NOR2_X2 \GFM/U396  ( .A1(\GFM/n25350 ), .A2(\GFM/n26110 ), .ZN(\GFM/N1119 ));
NOR2_X2 \GFM/U395  ( .A1(\GFM/n2610 ), .A2(\GFM/n25360 ), .ZN(\GFM/N1117 ));
NOR2_X2 \GFM/U394  ( .A1(\GFM/n25350 ), .A2(\GFM/n2613 ), .ZN(\GFM/N1181 ));
NOR2_X2 \GFM/U393  ( .A1(\GFM/n25450 ), .A2(\GFM/n26120 ), .ZN(\GFM/N1179 ));
NOR2_X2 \GFM/U392  ( .A1(\GFM/n25350 ), .A2(\GFM/n26140 ), .ZN(\GFM/N1212 ));
NOR2_X2 \GFM/U391  ( .A1(\GFM/n25450 ), .A2(\GFM/n2613 ), .ZN(\GFM/N1210 ));
NOR2_X2 \GFM/U390  ( .A1(\GFM/n25350 ), .A2(\GFM/n2618 ), .ZN(\GFM/N1336 ));
NOR2_X2 \GFM/U387  ( .A1(\GFM/n25450 ), .A2(\GFM/n2617 ), .ZN(\GFM/N1334 ));
NOR2_X2 \GFM/U385  ( .A1(\GFM/n25350 ), .A2(\GFM/n26190 ), .ZN(\GFM/N1367 ));
NOR2_X2 \GFM/U383  ( .A1(\GFM/n25450 ), .A2(\GFM/n2618 ), .ZN(\GFM/N1365 ));
NOR2_X2 \GFM/U382  ( .A1(\GFM/n2530 ), .A2(\GFM/n2672 ), .ZN(\GFM/N3010 ) );
NOR2_X2 \GFM/U380  ( .A1(\GFM/n2540 ), .A2(\GFM/n2671 ), .ZN(\GFM/N3008 ) );
NOR2_X2 \GFM/U378  ( .A1(\GFM/n2530 ), .A2(\GFM/n26730 ), .ZN(\GFM/N3041 ));
NOR2_X2 \GFM/U376  ( .A1(\GFM/n2540 ), .A2(\GFM/n2672 ), .ZN(\GFM/N3039 ) );
NOR2_X2 \GFM/U374  ( .A1(\GFM/n2530 ), .A2(\GFM/n26740 ), .ZN(\GFM/N3072 ));
NOR2_X2 \GFM/U372  ( .A1(\GFM/n2540 ), .A2(\GFM/n26730 ), .ZN(\GFM/N3070 ));
NOR2_X2 \GFM/U370  ( .A1(\GFM/n2530 ), .A2(\GFM/n2675 ), .ZN(\GFM/N3103 ) );
NOR2_X2 \GFM/U368  ( .A1(\GFM/n2540 ), .A2(\GFM/n26740 ), .ZN(\GFM/N3101 ));
NOR2_X2 \GFM/U366  ( .A1(\GFM/n2530 ), .A2(\GFM/n26760 ), .ZN(\GFM/N3134 ));
NOR2_X2 \GFM/U364  ( .A1(\GFM/n2540 ), .A2(\GFM/n2675 ), .ZN(\GFM/N3132 ) );
NOR2_X2 \GFM/U362  ( .A1(\GFM/n2530 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3165 ));
NOR2_X2 \GFM/U360  ( .A1(\GFM/n2540 ), .A2(\GFM/n26760 ), .ZN(\GFM/N3163 ));
NOR2_X2 \GFM/U358  ( .A1(\GFM/n25290 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3196 ));
NOR2_X2 \GFM/U357  ( .A1(\GFM/n2540 ), .A2(\GFM/n26770 ), .ZN(\GFM/N3194 ));
NOR2_X2 \GFM/U355  ( .A1(\GFM/n25290 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3227 ));
NOR2_X2 \GFM/U353  ( .A1(\GFM/n25390 ), .A2(\GFM/n2678 ), .ZN(\GFM/N3225 ));
NOR2_X2 \GFM/U351  ( .A1(\GFM/n2530 ), .A2(\GFM/n26801 ), .ZN(\GFM/N3258 ));
NOR2_X2 \GFM/U349  ( .A1(\GFM/n25390 ), .A2(\GFM/n2679 ), .ZN(\GFM/N3256 ));
NOR2_X2 \GFM/U347  ( .A1(\GFM/n21360 ), .A2(\GFM/n25260 ), .ZN(\GFM/N4221 ));
NOR2_X2 \GFM/U345  ( .A1(\GFM/n26980 ), .A2(\GFM/n2537 ), .ZN(\GFM/N4218 ));
NOR2_X2 \GFM/U343  ( .A1(\GFM/n2479 ), .A2(\GFM/n26900 ), .ZN(\GFM/N3433 ));
NOR2_X2 \GFM/U341  ( .A1(\GFM/n2479 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3471 ));
NOR2_X2 \GFM/U340  ( .A1(\GFM/n2499 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3600 ));
NOR2_X2 \GFM/U338  ( .A1(\GFM/n24980 ), .A2(\GFM/n26930 ), .ZN(\GFM/N3649 ));
NOR2_X2 \GFM/U336  ( .A1(\GFM/n24980 ), .A2(\GFM/n26940 ), .ZN(\GFM/N3703 ));
NOR2_X2 \GFM/U334  ( .A1(\GFM/n2499 ), .A2(\GFM/n26910 ), .ZN(\GFM/N3554 ));
NOR2_X2 \GFM/U332  ( .A1(\GFM/n2528 ), .A2(\GFM/n26921 ), .ZN(\GFM/N3748 ));
NOR2_X2 \GFM/U330  ( .A1(\GFM/n2533 ), .A2(\GFM/n25760 ), .ZN(\GFM/N189 ) );
NOR2_X2 \GFM/U328  ( .A1(\GFM/n25430 ), .A2(\GFM/n2573 ), .ZN(\GFM/N187 ) );
NOR2_X2 \GFM/U326  ( .A1(\GFM/n25310 ), .A2(\GFM/n25821 ), .ZN(\GFM/N282 ));
NOR2_X2 \GFM/U324  ( .A1(\GFM/n2541 ), .A2(\GFM/n25800 ), .ZN(\GFM/N280 ) );
NOR2_X2 \GFM/U323  ( .A1(\GFM/n25380 ), .A2(\GFM/n2587 ), .ZN(\GFM/N404 ) );
NOR2_X2 \GFM/U322  ( .A1(\GFM/n25880 ), .A2(\GFM/n25260 ), .ZN(\GFM/N406 ));
NOR2_X2 \GFM/U321  ( .A1(\GFM/n2554 ), .A2(\GFM/n2537 ), .ZN(\GFM/N32 ) );
NOR2_X2 \GFM/U320  ( .A1(\GFM/n25580 ), .A2(\GFM/n25260 ), .ZN(\GFM/N34 ) );
NOR2_X2 \GFM/U319  ( .A1(\GFM/n25350 ), .A2(\GFM/n25700 ), .ZN(\GFM/N127 ));
NOR2_X2 \GFM/U318  ( .A1(\GFM/n25660 ), .A2(\GFM/n25360 ), .ZN(\GFM/N125 ));
INV_X4 \GFM/U317  ( .A(v_out[111]), .ZN(\GFM/n25511 ) );
INV_X4 \GFM/U316  ( .A(v_out[110]), .ZN(\GFM/n25520 ) );
NOR2_X2 \GFM/U315  ( .A1(\GFM/n2399 ), .A2(\GFM/n2585 ), .ZN(\GFM/N4269 ) );
NOR2_X2 \GFM/U314  ( .A1(\GFM/n2399 ), .A2(\GFM/n25830 ), .ZN(\GFM/N4210 ));
NOR2_X2 \GFM/U313  ( .A1(\GFM/n2389 ), .A2(\GFM/n2575 ), .ZN(\GFM/N3923 ) );
NOR2_X2 \GFM/U312  ( .A1(\GFM/n2389 ), .A2(\GFM/n2585 ), .ZN(\GFM/N4213 ) );
NOR2_X2 \GFM/U311  ( .A1(\GFM/n2409 ), .A2(\GFM/n25690 ), .ZN(\GFM/N3918 ));
NOR2_X2 \GFM/U310  ( .A1(\GFM/n2418 ), .A2(\GFM/n25690 ), .ZN(\GFM/N3966 ));
NOR2_X2 \GFM/U309  ( .A1(\GFM/n2399 ), .A2(\GFM/n25810 ), .ZN(\GFM/N4151 ));
NOR2_X2 \GFM/U308  ( .A1(\GFM/n2409 ), .A2(\GFM/n25810 ), .ZN(\GFM/N4203 ));
NOR2_X2 \GFM/U307  ( .A1(\GFM/n2389 ), .A2(\GFM/n25830 ), .ZN(\GFM/N4154 ));
NOR2_X2 \GFM/U306  ( .A1(\GFM/n2389 ), .A2(\GFM/n2572 ), .ZN(\GFM/N3859 ) );
NOR2_X2 \GFM/U305  ( .A1(\GFM/n2399 ), .A2(\GFM/n2572 ), .ZN(\GFM/N3914 ) );
NOR2_X2 \GFM/U304  ( .A1(\GFM/n2409 ), .A2(\GFM/n2565 ), .ZN(\GFM/N3854 ) );
NOR2_X2 \GFM/U303  ( .A1(\GFM/n24190 ), .A2(\GFM/n2565 ), .ZN(\GFM/N3899 ));
NOR2_X2 \GFM/U302  ( .A1(\GFM/n2399 ), .A2(\GFM/n2579 ), .ZN(\GFM/N4094 ) );
NOR2_X2 \GFM/U301  ( .A1(\GFM/n2389 ), .A2(\GFM/n25810 ), .ZN(\GFM/N4097 ));
NOR2_X2 \GFM/U300  ( .A1(\GFM/n2489 ), .A2(\GFM/n2548 ), .ZN(\GFM/N4113 ) );
NOR2_X2 \GFM/U299  ( .A1(\GFM/n24980 ), .A2(\GFM/n25500 ), .ZN(\GFM/N4116 ));
NOR2_X2 \GFM/U298  ( .A1(\GFM/n24880 ), .A2(\GFM/n2556 ), .ZN(\GFM/N4172 ));
NOR2_X2 \GFM/U297  ( .A1(\GFM/n24980 ), .A2(\GFM/n2548 ), .ZN(\GFM/N4175 ));
NOR2_X2 \GFM/U296  ( .A1(\GFM/n2489 ), .A2(\GFM/n25600 ), .ZN(\GFM/N4233 ));
NOR2_X2 \GFM/U295  ( .A1(\GFM/n24980 ), .A2(\GFM/n2556 ), .ZN(\GFM/N4236 ));
NOR2_X2 \GFM/U294  ( .A1(\GFM/n24380 ), .A2(\GFM/n2564 ), .ZN(\GFM/N4017 ));
NOR2_X2 \GFM/U293  ( .A1(\GFM/n2400 ), .A2(\GFM/n25770 ), .ZN(\GFM/N4039 ));
NOR2_X2 \GFM/U292  ( .A1(\GFM/n2449 ), .A2(\GFM/n25600 ), .ZN(\GFM/N4024 ));
NOR2_X2 \GFM/U291  ( .A1(\GFM/n2409 ), .A2(\GFM/n25740 ), .ZN(\GFM/N4032 ));
NOR2_X2 \GFM/U290  ( .A1(\GFM/n2449 ), .A2(\GFM/n2564 ), .ZN(\GFM/N4079 ) );
NOR2_X2 \GFM/U289  ( .A1(\GFM/n24101 ), .A2(\GFM/n25770 ), .ZN(\GFM/N4087 ));
NOR2_X2 \GFM/U288  ( .A1(\GFM/n2478 ), .A2(\GFM/n2548 ), .ZN(\GFM/N4063 ) );
NOR2_X2 \GFM/U287  ( .A1(\GFM/n24390 ), .A2(\GFM/n2568 ), .ZN(\GFM/N4072 ));
NOR2_X2 \GFM/U286  ( .A1(\GFM/n2479 ), .A2(\GFM/n2556 ), .ZN(\GFM/N4120 ) );
NOR2_X2 \GFM/U285  ( .A1(\GFM/n24390 ), .A2(\GFM/n2571 ), .ZN(\GFM/N4129 ));
NOR2_X2 \GFM/U284  ( .A1(\GFM/n2448 ), .A2(\GFM/n2568 ), .ZN(\GFM/N4136 ) );
NOR2_X2 \GFM/U283  ( .A1(\GFM/n2409 ), .A2(\GFM/n2579 ), .ZN(\GFM/N4144 ) );
NOR2_X2 \GFM/U282  ( .A1(\GFM/n24380 ), .A2(\GFM/n25740 ), .ZN(\GFM/N4188 ));
NOR2_X2 \GFM/U281  ( .A1(\GFM/n2448 ), .A2(\GFM/n2571 ), .ZN(\GFM/N4195 ) );
NOR2_X2 \GFM/U280  ( .A1(\GFM/n24380 ), .A2(\GFM/n25770 ), .ZN(\GFM/N4249 ));
NOR2_X2 \GFM/U279  ( .A1(\GFM/n2449 ), .A2(\GFM/n25740 ), .ZN(\GFM/N4255 ));
NOR2_X2 \GFM/U278  ( .A1(\GFM/n25180 ), .A2(\GFM/n25500 ), .ZN(\GFM/N4225 ));
NOR2_X2 \GFM/U277  ( .A1(\GFM/n2509 ), .A2(\GFM/n2548 ), .ZN(\GFM/N4228 ) );
NOR2_X2 \GFM/U276  ( .A1(\GFM/n2489 ), .A2(\GFM/n25500 ), .ZN(\GFM/N4057 ));
NOR2_X2 \GFM/U275  ( .A1(\GFM/n2418 ), .A2(\GFM/n25810 ), .ZN(\GFM/N4265 ));
NOR2_X2 \GFM/U274  ( .A1(\GFM/n2400 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3580 ));
NOR2_X2 \GFM/U273  ( .A1(\GFM/n24101 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3615 ));
NOR2_X2 \GFM/U272  ( .A1(\GFM/n2449 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3844 ));
NOR2_X2 \GFM/U271  ( .A1(\GFM/n24590 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3889 ));
NOR2_X2 \GFM/U270  ( .A1(\GFM/n2418 ), .A2(\GFM/n25611 ), .ZN(\GFM/N3835 ));
NOR2_X2 \GFM/U269  ( .A1(\GFM/n2400 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3534 ));
NOR2_X2 \GFM/U268  ( .A1(\GFM/n24101 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3566 ));
NOR2_X2 \GFM/U267  ( .A1(\GFM/n2449 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3783 ));
NOR2_X2 \GFM/U266  ( .A1(\GFM/n2458 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3825 ));
NOR2_X2 \GFM/U265  ( .A1(\GFM/n2389 ), .A2(\GFM/n2565 ), .ZN(\GFM/N3740 ) );
NOR2_X2 \GFM/U264  ( .A1(\GFM/n2399 ), .A2(\GFM/n2565 ), .ZN(\GFM/N3789 ) );
NOR2_X2 \GFM/U263  ( .A1(\GFM/n24290 ), .A2(\GFM/n2565 ), .ZN(\GFM/N3962 ));
NOR2_X2 \GFM/U262  ( .A1(\GFM/n2400 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3681 ));
NOR2_X2 \GFM/U261  ( .A1(\GFM/n2409 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3735 ));
NOR2_X2 \GFM/U260  ( .A1(\GFM/n2448 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3975 ));
NOR2_X2 \GFM/U259  ( .A1(\GFM/n24690 ), .A2(\GFM/n2548 ), .ZN(\GFM/N4012 ));
NOR2_X2 \GFM/U258  ( .A1(\GFM/n24280 ), .A2(\GFM/n2568 ), .ZN(\GFM/N4020 ));
NOR2_X2 \GFM/U257  ( .A1(\GFM/n23900 ), .A2(\GFM/n2579 ), .ZN(\GFM/N4042 ));
NOR2_X2 \GFM/U256  ( .A1(\GFM/n24190 ), .A2(\GFM/n2571 ), .ZN(\GFM/N4035 ));
NOR2_X2 \GFM/U255  ( .A1(\GFM/n2418 ), .A2(\GFM/n25740 ), .ZN(\GFM/N4090 ));
NOR2_X2 \GFM/U254  ( .A1(\GFM/n24280 ), .A2(\GFM/n2571 ), .ZN(\GFM/N4075 ));
NOR2_X2 \GFM/U253  ( .A1(\GFM/n24290 ), .A2(\GFM/n25740 ), .ZN(\GFM/N4132 ));
NOR2_X2 \GFM/U252  ( .A1(\GFM/n2418 ), .A2(\GFM/n25770 ), .ZN(\GFM/N4147 ));
NOR2_X2 \GFM/U251  ( .A1(\GFM/n2468 ), .A2(\GFM/n2564 ), .ZN(\GFM/N4182 ) );
NOR2_X2 \GFM/U250  ( .A1(\GFM/n24280 ), .A2(\GFM/n25770 ), .ZN(\GFM/N4191 ));
NOR2_X2 \GFM/U249  ( .A1(\GFM/n2418 ), .A2(\GFM/n2579 ), .ZN(\GFM/N4206 ) );
NOR2_X2 \GFM/U248  ( .A1(\GFM/n24690 ), .A2(\GFM/n2568 ), .ZN(\GFM/N4243 ));
NOR2_X2 \GFM/U247  ( .A1(\GFM/n24280 ), .A2(\GFM/n2579 ), .ZN(\GFM/N4251 ));
NOR2_X2 \GFM/U246  ( .A1(\GFM/n24590 ), .A2(\GFM/n2571 ), .ZN(\GFM/N4258 ));
NOR2_X2 \GFM/U245  ( .A1(\GFM/n23900 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3538 ));
NOR2_X2 \GFM/U244  ( .A1(\GFM/n24190 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3662 ));
NOR2_X2 \GFM/U243  ( .A1(\GFM/n24290 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3715 ));
NOR2_X2 \GFM/U242  ( .A1(\GFM/n24390 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3780 ));
NOR2_X2 \GFM/U241  ( .A1(\GFM/n2468 ), .A2(\GFM/n25511 ), .ZN(\GFM/N3951 ));
NOR2_X2 \GFM/U240  ( .A1(\GFM/n2389 ), .A2(\GFM/n25611 ), .ZN(\GFM/N3685 ));
NOR2_X2 \GFM/U239  ( .A1(\GFM/n2400 ), .A2(\GFM/n25611 ), .ZN(\GFM/N3731 ));
NOR2_X2 \GFM/U238  ( .A1(\GFM/n24290 ), .A2(\GFM/n25611 ), .ZN(\GFM/N3895 ));
NOR2_X2 \GFM/U237  ( .A1(\GFM/n24390 ), .A2(\GFM/n25611 ), .ZN(\GFM/N3971 ));
NOR2_X2 \GFM/U236  ( .A1(\GFM/n23900 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3495 ));
NOR2_X2 \GFM/U235  ( .A1(\GFM/n24190 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3611 ));
NOR2_X2 \GFM/U234  ( .A1(\GFM/n24290 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3670 ));
NOR2_X2 \GFM/U233  ( .A1(\GFM/n24390 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3723 ));
NOR2_X2 \GFM/U232  ( .A1(\GFM/n2479 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3944 ));
NOR2_X2 \GFM/U231  ( .A1(\GFM/n2400 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3629 ));
NOR2_X2 \GFM/U230  ( .A1(\GFM/n24101 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3666 ));
NOR2_X2 \GFM/U229  ( .A1(\GFM/n2418 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3719 ));
NOR2_X2 \GFM/U228  ( .A1(\GFM/n2449 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3908 ));
NOR2_X2 \GFM/U227  ( .A1(\GFM/n24590 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3955 ));
NOR2_X2 \GFM/U226  ( .A1(\GFM/n23900 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3633 ));
NOR2_X2 \GFM/U225  ( .A1(\GFM/n24290 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3831 ));
NOR2_X2 \GFM/U224  ( .A1(\GFM/n25670 ), .A2(\GFM/n24260 ), .ZN(\GFM/N3620 ));
NOR2_X2 \GFM/U223  ( .A1(\GFM/n25670 ), .A2(\GFM/n2437 ), .ZN(\GFM/N3672 ));
NOR2_X2 \GFM/U222  ( .A1(\GFM/n25670 ), .A2(\GFM/n24560 ), .ZN(\GFM/N3764 ));
NOR2_X2 \GFM/U221  ( .A1(\GFM/n25670 ), .A2(\GFM/n24670 ), .ZN(\GFM/N3818 ));
NOR2_X2 \GFM/U220  ( .A1(\GFM/n25670 ), .A2(\GFM/n24770 ), .ZN(\GFM/N3881 ));
NOR2_X2 \GFM/U219  ( .A1(\GFM/n2389 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3584 ));
NOR2_X2 \GFM/U218  ( .A1(\GFM/n24290 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3771 ));
NOR2_X2 \GFM/U217  ( .A1(\GFM/n24390 ), .A2(\GFM/n25490 ), .ZN(\GFM/N3840 ));
NOR2_X2 \GFM/U216  ( .A1(\GFM/n25630 ), .A2(\GFM/n24080 ), .ZN(\GFM/N3491 ));
NOR2_X2 \GFM/U215  ( .A1(\GFM/n25630 ), .A2(\GFM/n24570 ), .ZN(\GFM/N3708 ));
NOR2_X2 \GFM/U214  ( .A1(\GFM/n25630 ), .A2(\GFM/n24960 ), .ZN(\GFM/N3939 ));
NOR2_X2 \GFM/U213  ( .A1(\GFM/n2559 ), .A2(\GFM/n24070 ), .ZN(\GFM/N3452 ));
NOR2_X2 \GFM/U212  ( .A1(\GFM/n2559 ), .A2(\GFM/n2427 ), .ZN(\GFM/N3521 ) );
NOR2_X2 \GFM/U211  ( .A1(\GFM/n2559 ), .A2(\GFM/n24560 ), .ZN(\GFM/N3655 ));
NOR2_X2 \GFM/U210  ( .A1(\GFM/n25670 ), .A2(\GFM/n2387 ), .ZN(\GFM/N3455 ));
NOR2_X2 \GFM/U209  ( .A1(\GFM/n25670 ), .A2(\GFM/n23970 ), .ZN(\GFM/N3489 ));
NOR2_X2 \GFM/U208  ( .A1(\GFM/n25670 ), .A2(\GFM/n25530 ), .ZN(\GFM/N3563 ));
NOR2_X2 \GFM/U207  ( .A1(\GFM/n2555 ), .A2(\GFM/n24080 ), .ZN(\GFM/N3415 ));
NOR2_X2 \GFM/U206  ( .A1(\GFM/n2555 ), .A2(\GFM/n2427 ), .ZN(\GFM/N3477 ) );
NOR2_X2 \GFM/U205  ( .A1(\GFM/n2555 ), .A2(\GFM/n2437 ), .ZN(\GFM/N3527 ) );
NOR2_X2 \GFM/U204  ( .A1(\GFM/n2555 ), .A2(\GFM/n24560 ), .ZN(\GFM/N3605 ));
NOR2_X2 \GFM/U203  ( .A1(\GFM/n2555 ), .A2(\GFM/n24870 ), .ZN(\GFM/N3754 ));
NOR2_X2 \GFM/U202  ( .A1(\GFM/n25630 ), .A2(\GFM/n2387 ), .ZN(\GFM/N3418 ));
NOR2_X2 \GFM/U201  ( .A1(\GFM/n25630 ), .A2(\GFM/n25530 ), .ZN(\GFM/N3519 ));
NOR2_X2 \GFM/U200  ( .A1(\GFM/n25630 ), .A2(\GFM/n2437 ), .ZN(\GFM/N3618 ));
NOR2_X2 \GFM/U199  ( .A1(\GFM/n2559 ), .A2(\GFM/n2387 ), .ZN(\GFM/N3383 ) );
NOR2_X2 \GFM/U198  ( .A1(\GFM/n2559 ), .A2(\GFM/n2417 ), .ZN(\GFM/N3479 ) );
NOR2_X2 \GFM/U197  ( .A1(\GFM/n2559 ), .A2(\GFM/n2437 ), .ZN(\GFM/N3569 ) );
NOR2_X2 \GFM/U196  ( .A1(\GFM/n2559 ), .A2(\GFM/n24670 ), .ZN(\GFM/N3706 ));
NOR2_X2 \GFM/U195  ( .A1(\GFM/n2559 ), .A2(\GFM/n24770 ), .ZN(\GFM/N3756 ));
NOR2_X2 \GFM/U194  ( .A1(\GFM/n2547 ), .A2(\GFM/n24870 ), .ZN(\GFM/N3699 ));
NOR2_X2 \GFM/U193  ( .A1(\GFM/n2555 ), .A2(\GFM/n24770 ), .ZN(\GFM/N3701 ));
NOR2_X2 \GFM/U192  ( .A1(\GFM/n2547 ), .A2(\GFM/n24070 ), .ZN(\GFM/N3380 ));
NOR2_X2 \GFM/U191  ( .A1(\GFM/n2547 ), .A2(\GFM/n24260 ), .ZN(\GFM/N3439 ));
NOR2_X2 \GFM/U190  ( .A1(\GFM/n2547 ), .A2(\GFM/n2437 ), .ZN(\GFM/N3482 ) );
NOR2_X2 \GFM/U189  ( .A1(\GFM/n2547 ), .A2(\GFM/n24570 ), .ZN(\GFM/N3558 ));
NOR2_X2 \GFM/U188  ( .A1(\GFM/n2547 ), .A2(\GFM/n24960 ), .ZN(\GFM/N3759 ));
NOR2_X2 \GFM/U187  ( .A1(\GFM/n2555 ), .A2(\GFM/n2387 ), .ZN(\GFM/N3349 ) );
NOR2_X2 \GFM/U186  ( .A1(\GFM/n2555 ), .A2(\GFM/n23970 ), .ZN(\GFM/N3378 ));
NOR2_X2 \GFM/U185  ( .A1(\GFM/n2555 ), .A2(\GFM/n25530 ), .ZN(\GFM/N3441 ));
NOR2_X2 \GFM/U184  ( .A1(\GFM/n2555 ), .A2(\GFM/n24460 ), .ZN(\GFM/N3574 ));
NOR2_X2 \GFM/U183  ( .A1(\GFM/n2555 ), .A2(\GFM/n2466 ), .ZN(\GFM/N3653 ) );
NOR2_X2 \GFM/U182  ( .A1(\GFM/n2555 ), .A2(\GFM/n2516 ), .ZN(\GFM/N3936 ) );
NOR2_X2 \GFM/U181  ( .A1(\GFM/n2547 ), .A2(\GFM/n2387 ), .ZN(\GFM/N3316 ) );
NOR2_X2 \GFM/U180  ( .A1(\GFM/n2547 ), .A2(\GFM/n23970 ), .ZN(\GFM/N3345 ));
NOR2_X2 \GFM/U179  ( .A1(\GFM/n2547 ), .A2(\GFM/n2417 ), .ZN(\GFM/N3404 ) );
NOR2_X2 \GFM/U178  ( .A1(\GFM/n2547 ), .A2(\GFM/n2447 ), .ZN(\GFM/N3529 ) );
NOR2_X2 \GFM/U177  ( .A1(\GFM/n2547 ), .A2(\GFM/n2466 ), .ZN(\GFM/N3603 ) );
NOR2_X2 \GFM/U176  ( .A1(\GFM/n25670 ), .A2(\GFM/n24070 ), .ZN(\GFM/N3524 ));
NOR2_X2 \GFM/U175  ( .A1(\GFM/n25630 ), .A2(\GFM/n2447 ), .ZN(\GFM/N3674 ));
NOR2_X2 \GFM/U174  ( .A1(\GFM/n25670 ), .A2(\GFM/n2447 ), .ZN(\GFM/N3725 ));
NOR2_X2 \GFM/U173  ( .A1(\GFM/n24380 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3904 ));
NOR2_X2 \GFM/U172  ( .A1(\GFM/n2409 ), .A2(\GFM/n25830 ), .ZN(\GFM/N4263 ));
NOR2_X2 \GFM/U171  ( .A1(\GFM/n2399 ), .A2(\GFM/n2575 ), .ZN(\GFM/N3981 ) );
NOR2_X2 \GFM/U170  ( .A1(\GFM/n25630 ), .A2(\GFM/n2427 ), .ZN(\GFM/N3571 ));
NOR2_X2 \GFM/U169  ( .A1(\GFM/n2559 ), .A2(\GFM/n2447 ), .ZN(\GFM/N3623 ) );
NOR2_X2 \GFM/U168  ( .A1(\GFM/n2399 ), .A2(\GFM/n25690 ), .ZN(\GFM/N3850 ));
NOR2_X2 \GFM/U167  ( .A1(\GFM/n2389 ), .A2(\GFM/n25690 ), .ZN(\GFM/N3798 ));
NOR2_X2 \GFM/U166  ( .A1(\GFM/n24101 ), .A2(\GFM/n25611 ), .ZN(\GFM/N3793 ));
NOR2_X2 \GFM/U165  ( .A1(\GFM/n2547 ), .A2(\GFM/n2516 ), .ZN(\GFM/N3871 ) );
NOR2_X2 \GFM/U164  ( .A1(\GFM/n2555 ), .A2(\GFM/n25080 ), .ZN(\GFM/N3869 ));
NOR2_X2 \GFM/U163  ( .A1(\GFM/n25670 ), .A2(\GFM/n24870 ), .ZN(\GFM/N3946 ));
NOR2_X2 \GFM/U162  ( .A1(\GFM/n24190 ), .A2(\GFM/n25570 ), .ZN(\GFM/N3775 ));
NOR2_X2 \GFM/U161  ( .A1(\GFM/n2559 ), .A2(\GFM/n24870 ), .ZN(\GFM/N3821 ));
NOR2_X2 \GFM/U160  ( .A1(\GFM/n25630 ), .A2(\GFM/n24870 ), .ZN(\GFM/N3883 ));
NOR2_X2 \GFM/U159  ( .A1(\GFM/n24590 ), .A2(\GFM/n2556 ), .ZN(\GFM/N4027 ));
NOR2_X2 \GFM/U158  ( .A1(\GFM/n24590 ), .A2(\GFM/n25600 ), .ZN(\GFM/N4082 ));
NOR2_X2 \GFM/U157  ( .A1(\GFM/n2468 ), .A2(\GFM/n2556 ), .ZN(\GFM/N4066 ) );
NOR2_X2 \GFM/U156  ( .A1(\GFM/n2468 ), .A2(\GFM/n25600 ), .ZN(\GFM/N4123 ));
NOR2_X2 \GFM/U155  ( .A1(\GFM/n2458 ), .A2(\GFM/n2564 ), .ZN(\GFM/N4139 ) );
NOR2_X2 \GFM/U154  ( .A1(\GFM/n2478 ), .A2(\GFM/n25600 ), .ZN(\GFM/N4179 ));
NOR2_X2 \GFM/U153  ( .A1(\GFM/n2458 ), .A2(\GFM/n2568 ), .ZN(\GFM/N4198 ) );
NOR2_X2 \GFM/U152  ( .A1(\GFM/n2478 ), .A2(\GFM/n2564 ), .ZN(\GFM/N4240 ) );
NOR2_X2 \GFM/U151  ( .A1(\GFM/n25630 ), .A2(\GFM/n2466 ), .ZN(\GFM/N3762 ));
NOR2_X2 \GFM/U150  ( .A1(\GFM/n2559 ), .A2(\GFM/n25070 ), .ZN(\GFM/N3934 ));
NOR2_X2 \GFM/U149  ( .A1(\GFM/n2555 ), .A2(\GFM/n24960 ), .ZN(\GFM/N3812 ));
NOR2_X2 \GFM/U148  ( .A1(\GFM/n25630 ), .A2(\GFM/n24770 ), .ZN(\GFM/N3816 ));
NOR2_X2 \GFM/U147  ( .A1(\GFM/n2468 ), .A2(\GFM/n25520 ), .ZN(\GFM/N3879 ));
NOR2_X2 \GFM/U146  ( .A1(\GFM/n2559 ), .A2(\GFM/n24960 ), .ZN(\GFM/N3874 ));
INV_X4 \GFM/U145  ( .A(b_in[112]), .ZN(\GFM/n2396 ) );
INV_X4 \GFM/U144  ( .A(b_in[114]), .ZN(\GFM/n2416 ) );
INV_X4 \GFM/U143  ( .A(b_in[120]), .ZN(\GFM/n2475 ) );
INV_X4 \GFM/U142  ( .A(b_in[113]), .ZN(\GFM/n2406 ) );
INV_X4 \GFM/U141  ( .A(b_in[125]), .ZN(\GFM/n2525 ) );
INV_X4 \GFM/U140  ( .A(b_in[123]), .ZN(\GFM/n25050 ) );
INV_X4 \GFM/U139  ( .A(b_in[115]), .ZN(\GFM/n24250 ) );
INV_X4 \GFM/U138  ( .A(b_in[121]), .ZN(\GFM/n2485 ) );
INV_X4 \GFM/U137  ( .A(b_in[117]), .ZN(\GFM/n24450 ) );
INV_X4 \GFM/U136  ( .A(b_in[118]), .ZN(\GFM/n2455 ) );
INV_X4 \GFM/U135  ( .A(b_in[122]), .ZN(\GFM/n24950 ) );
INV_X4 \GFM/U134  ( .A(b_in[119]), .ZN(\GFM/n24650 ) );
INV_X4 \GFM/U133  ( .A(b_in[124]), .ZN(\GFM/n25150 ) );
INV_X4 \GFM/U132  ( .A(b_in[116]), .ZN(\GFM/n2435 ) );
INV_X4 \GFM/U131  ( .A(b_in[116]), .ZN(\GFM/n2427 ) );
INV_X4 \GFM/U130  ( .A(b_in[121]), .ZN(\GFM/n24770 ) );
INV_X4 \GFM/U129  ( .A(b_in[122]), .ZN(\GFM/n24870 ) );
INV_X4 \GFM/U128  ( .A(b_in[124]), .ZN(\GFM/n25070 ) );
INV_X4 \GFM/U127  ( .A(b_in[118]), .ZN(\GFM/n2454 ) );
INV_X4 \GFM/U126  ( .A(b_in[116]), .ZN(\GFM/n24340 ) );
INV_X4 \GFM/U125  ( .A(b_in[122]), .ZN(\GFM/n24880 ) );
INV_X4 \GFM/U124  ( .A(b_in[119]), .ZN(\GFM/n2463 ) );
INV_X4 \GFM/U123  ( .A(b_in[120]), .ZN(\GFM/n24730 ) );
INV_X4 \GFM/U122  ( .A(b_in[114]), .ZN(\GFM/n2413 ) );
INV_X4 \GFM/U121  ( .A(b_in[115]), .ZN(\GFM/n24220 ) );
INV_X4 \GFM/U120  ( .A(b_in[121]), .ZN(\GFM/n2478 ) );
INV_X4 \GFM/U119  ( .A(b_in[117]), .ZN(\GFM/n24380 ) );
INV_X4 \GFM/U118  ( .A(b_in[118]), .ZN(\GFM/n2448 ) );
INV_X4 \GFM/U117  ( .A(b_in[116]), .ZN(\GFM/n24280 ) );
INV_X4 \GFM/U116  ( .A(b_in[122]), .ZN(\GFM/n2489 ) );
INV_X4 \GFM/U115  ( .A(b_in[119]), .ZN(\GFM/n2458 ) );
INV_X4 \GFM/U114  ( .A(b_in[120]), .ZN(\GFM/n2468 ) );
INV_X4 \GFM/U113  ( .A(b_in[115]), .ZN(\GFM/n2418 ) );
INV_X4 \GFM/U112  ( .A(b_in[123]), .ZN(\GFM/n2497 ) );
INV_X4 \GFM/U111  ( .A(b_in[121]), .ZN(\GFM/n2479 ) );
INV_X4 \GFM/U110  ( .A(b_in[125]), .ZN(\GFM/n2517 ) );
INV_X4 \GFM/U109  ( .A(b_in[114]), .ZN(\GFM/n24150 ) );
INV_X4 \GFM/U108  ( .A(b_in[115]), .ZN(\GFM/n2424 ) );
INV_X4 \GFM/U107  ( .A(b_in[120]), .ZN(\GFM/n24740 ) );
INV_X4 \GFM/U106  ( .A(b_in[113]), .ZN(\GFM/n24050 ) );
INV_X4 \GFM/U105  ( .A(b_in[121]), .ZN(\GFM/n24840 ) );
INV_X4 \GFM/U104  ( .A(b_in[125]), .ZN(\GFM/n2524 ) );
INV_X4 \GFM/U103  ( .A(b_in[123]), .ZN(\GFM/n25040 ) );
INV_X4 \GFM/U102  ( .A(b_in[122]), .ZN(\GFM/n2494 ) );
INV_X4 \GFM/U101  ( .A(b_in[114]), .ZN(\GFM/n24140 ) );
INV_X4 \GFM/U100  ( .A(b_in[115]), .ZN(\GFM/n2423 ) );
INV_X4 \GFM/U99  ( .A(b_in[119]), .ZN(\GFM/n24640 ) );
INV_X4 \GFM/U98  ( .A(b_in[113]), .ZN(\GFM/n2404 ) );
INV_X4 \GFM/U97  ( .A(b_in[121]), .ZN(\GFM/n24830 ) );
INV_X4 \GFM/U96  ( .A(b_in[117]), .ZN(\GFM/n24430 ) );
INV_X4 \GFM/U95  ( .A(b_in[116]), .ZN(\GFM/n24330 ) );
INV_X4 \GFM/U94  ( .A(b_in[125]), .ZN(\GFM/n2523 ) );
INV_X4 \GFM/U93  ( .A(b_in[123]), .ZN(\GFM/n2503 ) );
INV_X4 \GFM/U92  ( .A(b_in[124]), .ZN(\GFM/n25140 ) );
INV_X4 \GFM/U91  ( .A(b_in[113]), .ZN(\GFM/n24030 ) );
INV_X4 \GFM/U90  ( .A(b_in[117]), .ZN(\GFM/n24420 ) );
INV_X4 \GFM/U89  ( .A(b_in[118]), .ZN(\GFM/n24520 ) );
INV_X4 \GFM/U88  ( .A(b_in[116]), .ZN(\GFM/n2432 ) );
INV_X4 \GFM/U87  ( .A(b_in[125]), .ZN(\GFM/n25220 ) );
INV_X4 \GFM/U86  ( .A(b_in[123]), .ZN(\GFM/n2502 ) );
INV_X4 \GFM/U85  ( .A(b_in[124]), .ZN(\GFM/n2513 ) );
INV_X4 \GFM/U84  ( .A(b_in[122]), .ZN(\GFM/n2493 ) );
INV_X4 \GFM/U83  ( .A(b_in[117]), .ZN(\GFM/n2441 ) );
INV_X4 \GFM/U82  ( .A(b_in[118]), .ZN(\GFM/n24511 ) );
INV_X4 \GFM/U81  ( .A(b_in[116]), .ZN(\GFM/n2431 ) );
INV_X4 \GFM/U80  ( .A(b_in[125]), .ZN(\GFM/n25210 ) );
INV_X4 \GFM/U79  ( .A(b_in[123]), .ZN(\GFM/n25010 ) );
INV_X4 \GFM/U78  ( .A(b_in[124]), .ZN(\GFM/n25120 ) );
INV_X4 \GFM/U77  ( .A(b_in[122]), .ZN(\GFM/n24921 ) );
INV_X4 \GFM/U76  ( .A(b_in[119]), .ZN(\GFM/n2461 ) );
INV_X4 \GFM/U75  ( .A(b_in[114]), .ZN(\GFM/n24120 ) );
INV_X4 \GFM/U74  ( .A(b_in[115]), .ZN(\GFM/n24210 ) );
INV_X4 \GFM/U73  ( .A(b_in[113]), .ZN(\GFM/n24020 ) );
INV_X4 \GFM/U72  ( .A(b_in[116]), .ZN(\GFM/n2430 ) );
INV_X4 \GFM/U71  ( .A(b_in[125]), .ZN(\GFM/n25201 ) );
INV_X4 \GFM/U70  ( .A(b_in[123]), .ZN(\GFM/n25000 ) );
INV_X4 \GFM/U69  ( .A(b_in[124]), .ZN(\GFM/n2511 ) );
INV_X4 \GFM/U68  ( .A(b_in[119]), .ZN(\GFM/n24600 ) );
INV_X4 \GFM/U67  ( .A(b_in[120]), .ZN(\GFM/n24700 ) );
INV_X4 \GFM/U66  ( .A(b_in[114]), .ZN(\GFM/n24110 ) );
INV_X4 \GFM/U65  ( .A(b_in[115]), .ZN(\GFM/n24201 ) );
INV_X4 \GFM/U64  ( .A(b_in[113]), .ZN(\GFM/n2401 ) );
INV_X4 \GFM/U63  ( .A(b_in[121]), .ZN(\GFM/n2480 ) );
INV_X4 \GFM/U62  ( .A(b_in[117]), .ZN(\GFM/n24401 ) );
INV_X4 \GFM/U61  ( .A(b_in[118]), .ZN(\GFM/n24500 ) );
INV_X4 \GFM/U60  ( .A(b_in[124]), .ZN(\GFM/n25101 ) );
INV_X4 \GFM/U59  ( .A(b_in[120]), .ZN(\GFM/n24690 ) );
INV_X4 \GFM/U58  ( .A(b_in[114]), .ZN(\GFM/n24101 ) );
INV_X4 \GFM/U57  ( .A(b_in[115]), .ZN(\GFM/n24190 ) );
INV_X4 \GFM/U56  ( .A(b_in[113]), .ZN(\GFM/n2400 ) );
INV_X4 \GFM/U55  ( .A(b_in[117]), .ZN(\GFM/n24390 ) );
INV_X4 \GFM/U54  ( .A(b_in[118]), .ZN(\GFM/n2449 ) );
INV_X4 \GFM/U53  ( .A(b_in[116]), .ZN(\GFM/n24290 ) );
INV_X4 \GFM/U52  ( .A(b_in[119]), .ZN(\GFM/n24590 ) );
INV_X4 \GFM/U51  ( .A(b_in[122]), .ZN(\GFM/n24910 ) );
INV_X4 \GFM/U50  ( .A(b_in[114]), .ZN(\GFM/n2409 ) );
INV_X4 \GFM/U49  ( .A(b_in[113]), .ZN(\GFM/n2399 ) );
INV_X4 \GFM/U48  ( .A(b_in[121]), .ZN(\GFM/n24810 ) );
INV_X4 \GFM/U47  ( .A(b_in[120]), .ZN(\GFM/n2471 ) );
INV_X4 \GFM/U46  ( .A(b_in[117]), .ZN(\GFM/n2444 ) );
INV_X4 \GFM/U45  ( .A(b_in[118]), .ZN(\GFM/n24530 ) );
INV_X4 \GFM/U44  ( .A(b_in[120]), .ZN(\GFM/n2472 ) );
INV_X4 \GFM/U43  ( .A(b_in[119]), .ZN(\GFM/n2462 ) );
INV_X4 \GFM/U42  ( .A(b_in[121]), .ZN(\GFM/n2482 ) );
INV_X4 \GFM/U41  ( .A(b_in[123]), .ZN(\GFM/n2499 ) );
INV_X4 \GFM/U40  ( .A(b_in[113]), .ZN(\GFM/n23980 ) );
INV_X4 \GFM/U39  ( .A(b_in[124]), .ZN(\GFM/n25080 ) );
INV_X4 \GFM/U38  ( .A(b_in[115]), .ZN(\GFM/n2417 ) );
INV_X4 \GFM/U37  ( .A(b_in[127]), .ZN(\GFM/n25450 ) );
INV_X4 \GFM/U36  ( .A(b_in[126]), .ZN(\GFM/n25350 ) );
INV_X4 \GFM/U35  ( .A(b_in[119]), .ZN(\GFM/n24570 ) );
INV_X4 \GFM/U34  ( .A(b_in[118]), .ZN(\GFM/n2447 ) );
INV_X4 \GFM/U33  ( .A(b_in[117]), .ZN(\GFM/n2437 ) );
INV_X4 \GFM/U32  ( .A(b_in[123]), .ZN(\GFM/n24980 ) );
INV_X4 \GFM/U31  ( .A(b_in[112]), .ZN(\GFM/n23880 ) );
INV_X4 \GFM/U30  ( .A(b_in[112]), .ZN(\GFM/n23950 ) );
INV_X4 \GFM/U29  ( .A(b_in[112]), .ZN(\GFM/n23940 ) );
INV_X4 \GFM/U28  ( .A(b_in[112]), .ZN(\GFM/n2393 ) );
INV_X4 \GFM/U27  ( .A(b_in[112]), .ZN(\GFM/n2392 ) );
INV_X4 \GFM/U26  ( .A(b_in[112]), .ZN(\GFM/n23910 ) );
INV_X4 \GFM/U25  ( .A(b_in[112]), .ZN(\GFM/n23900 ) );
INV_X4 \GFM/U24  ( .A(b_in[125]), .ZN(\GFM/n25190 ) );
INV_X4 \GFM/U23  ( .A(b_in[112]), .ZN(\GFM/n2389 ) );
INV_X4 \GFM/U22  ( .A(b_in[124]), .ZN(\GFM/n2509 ) );
INV_X4 \GFM/U21  ( .A(b_in[125]), .ZN(\GFM/n25180 ) );
INV_X4 \GFM/U20  ( .A(b_in[122]), .ZN(\GFM/n24900 ) );
INV_X4 \GFM/U19  ( .A(b_in[126]), .ZN(\GFM/n25290 ) );
INV_X4 \GFM/U18  ( .A(b_in[126]), .ZN(\GFM/n2528 ) );
INV_X4 \GFM/U17  ( .A(b_in[127]), .ZN(\GFM/n2544 ) );
INV_X4 \GFM/U16  ( .A(b_in[126]), .ZN(\GFM/n2534 ) );
INV_X4 \GFM/U15  ( .A(b_in[127]), .ZN(\GFM/n25430 ) );
INV_X4 \GFM/U14  ( .A(b_in[126]), .ZN(\GFM/n2533 ) );
INV_X4 \GFM/U13  ( .A(b_in[127]), .ZN(\GFM/n2542 ) );
INV_X4 \GFM/U12  ( .A(b_in[126]), .ZN(\GFM/n25320 ) );
INV_X4 \GFM/U11  ( .A(b_in[127]), .ZN(\GFM/n2541 ) );
INV_X4 \GFM/U10  ( .A(b_in[126]), .ZN(\GFM/n25310 ) );
INV_X4 \GFM/U9  ( .A(b_in[127]), .ZN(\GFM/n2540 ) );
INV_X4 \GFM/U8  ( .A(b_in[126]), .ZN(\GFM/n2530 ) );
INV_X4 \GFM/U7  ( .A(b_in[127]), .ZN(\GFM/n25390 ) );
INV_X4 \GFM/U6  ( .A(b_in[127]), .ZN(\GFM/n25380 ) );
INV_X4 \GFM/U5  ( .A(b_in[127]), .ZN(\GFM/n2537 ) );
INV_X4 \GFM/U4  ( .A(b_in[126]), .ZN(\GFM/n25270 ) );
INV_X4 \GFM/U3  ( .A(b_in[114]), .ZN(\GFM/n24080 ) );
INV_X4 \GFM/U2  ( .A(b_in[120]), .ZN(\GFM/n24670 ) );
XOR2_X2 \GFM/U755  ( .A(v_in[121]), .B(v_in[0]), .Z(v_out[105]) );
XNOR2_X2 \GFM/U737  ( .A(\GFM/n2695 ), .B(v_in[1]), .ZN(v_out[106]) );
XNOR2_X2 \GFM/U717  ( .A(\GFM/n2696 ), .B(v_in[2]), .ZN(v_out[107]) );
XNOR2_X2 \GFM/U699  ( .A(\GFM/n2697 ), .B(v_in[3]), .ZN(v_out[108]) );
XNOR2_X2 \GFM/U679  ( .A(\GFM/n26980 ), .B(v_in[4]), .ZN(v_out[109]) );
AND2_X2 \GFM/U487  ( .A1(v_out[119]), .A2(b_in[112]), .ZN(\GFM/N3990 ) );
AND2_X2 \GFM/U486  ( .A1(v_in[121]), .A2(b_in[127]), .ZN(\GFM/N3994 ) );
XOR2_X2 \GFM/U479  ( .A(v_in[126]), .B(\GFM/n25460 ), .Z(\GFM/n21360 ) );
AND2_X2 \GFM/U389  ( .A1(v_out[124]), .A2(b_in[112]), .ZN(\GFM/N4272 ) );
AND2_X2 \GFM/U388  ( .A1(b_in[127]), .A2(v_in[126]), .ZN(\GFM/N4276 ) );
NAND2_X2 \GFM/U386  ( .A1(\GFM/N4324 ), .A2(\GFM/n2699 ), .ZN(\GFM/n2134 ));
NAND2_X2 \GFM/U384  ( .A1(\GFM/n2134 ), .A2(\GFM/n21350 ), .ZN(\GFM/N4279 ));
NAND2_X2 \GFM/U381  ( .A1(\GFM/N4325 ), .A2(\GFM/n25460 ), .ZN(\GFM/n21320 ));
NAND2_X2 \GFM/U379  ( .A1(\GFM/n21320 ), .A2(\GFM/n21330 ), .ZN(\GFM/N4282 ));
NAND2_X2 \GFM/U377  ( .A1(\GFM/N4329 ), .A2(\GFM/n2554 ), .ZN(\GFM/n21301 ));
NAND2_X2 \GFM/U375  ( .A1(\GFM/n21301 ), .A2(\GFM/n2131 ), .ZN(\GFM/N4284 ));
NAND2_X2 \GFM/U373  ( .A1(\GFM/N4331 ), .A2(\GFM/n25620 ), .ZN(\GFM/n21280 ));
NAND2_X2 \GFM/U371  ( .A1(\GFM/n21280 ), .A2(\GFM/n21290 ), .ZN(\GFM/N4288 ));
NAND2_X2 \GFM/U369  ( .A1(\GFM/N4328 ), .A2(\GFM/n25580 ), .ZN(\GFM/n21260 ));
NAND2_X2 \GFM/U367  ( .A1(\GFM/n21260 ), .A2(\GFM/n2127 ), .ZN(\GFM/N4290 ));
NAND2_X2 \GFM/U365  ( .A1(\GFM/N4332 ), .A2(\GFM/n25660 ), .ZN(\GFM/n21240 ));
NAND2_X2 \GFM/U363  ( .A1(\GFM/n21240 ), .A2(\GFM/n2125 ), .ZN(\GFM/N4293 ));
NAND2_X2 \GFM/U361  ( .A1(\GFM/N4342 ), .A2(\GFM/n25700 ), .ZN(\GFM/n2122 ));
NAND2_X2 \GFM/U359  ( .A1(\GFM/n2122 ), .A2(\GFM/n21230 ), .ZN(\GFM/N4295 ));
NAND2_X2 \GFM/U356  ( .A1(\GFM/N4336 ), .A2(\GFM/n2578 ), .ZN(\GFM/n184 ) );
NAND2_X2 \GFM/U354  ( .A1(\GFM/n184 ), .A2(\GFM/n2121 ), .ZN(\GFM/N4300 ) );
NAND2_X2 \GFM/U352  ( .A1(\GFM/N4339 ), .A2(\GFM/n25800 ), .ZN(\GFM/n18210 ));
NAND2_X2 \GFM/U350  ( .A1(\GFM/n18210 ), .A2(\GFM/n18310 ), .ZN(\GFM/N4302 ));
NAND2_X2 \GFM/U348  ( .A1(\GFM/N4337 ), .A2(\GFM/n25760 ), .ZN(\GFM/n18011 ));
NAND2_X2 \GFM/U346  ( .A1(\GFM/n18011 ), .A2(\GFM/n181 ), .ZN(\GFM/N4305 ));
NAND2_X2 \GFM/U344  ( .A1(\GFM/N4341 ), .A2(\GFM/n2573 ), .ZN(\GFM/n178 ) );
NAND2_X2 \GFM/U342  ( .A1(\GFM/n178 ), .A2(\GFM/n17911 ), .ZN(\GFM/N4307 ));
NAND2_X2 \GFM/U339  ( .A1(\GFM/N4345 ), .A2(\GFM/n25840 ), .ZN(\GFM/n17611 ));
NAND2_X2 \GFM/U337  ( .A1(\GFM/n17611 ), .A2(\GFM/n177 ), .ZN(\GFM/N4311 ));
NAND2_X2 \GFM/U335  ( .A1(\GFM/N4346 ), .A2(\GFM/n25821 ), .ZN(\GFM/n174 ));
NAND2_X2 \GFM/U333  ( .A1(\GFM/n174 ), .A2(\GFM/n17511 ), .ZN(\GFM/N4313 ));
NAND2_X2 \GFM/U331  ( .A1(\GFM/N4348 ), .A2(\GFM/n2586 ), .ZN(\GFM/n172 ) );
NAND2_X2 \GFM/U329  ( .A1(\GFM/n172 ), .A2(\GFM/n17310 ), .ZN(\GFM/N4316 ));
NAND2_X2 \GFM/U327  ( .A1(\GFM/N4349 ), .A2(\GFM/n2587 ), .ZN(\GFM/n17011 ));
NAND2_X2 \GFM/U325  ( .A1(\GFM/n17011 ), .A2(\GFM/n17110 ), .ZN(\GFM/N4318 ));
XOR2_X2 \GFM/U1  ( .A(v_in[15]), .B(v_in[14]), .Z(v_out[126]) );
XOR2_X2 \GFM/U4328  ( .A(\GFM/n186 ), .B(\GFM/n185 ), .Z(z_out[0]) );
XOR2_X2 \GFM/U4327  ( .A(\GFM/n188 ), .B(\GFM/n18720 ), .Z(\GFM/n185 ) );
XOR2_X2 \GFM/U4326  ( .A(\GFM/n19000 ), .B(\GFM/n18900 ), .Z(\GFM/n186 ) );
XOR2_X2 \GFM/U4325  ( .A(\GFM/n192 ), .B(\GFM/n191 ), .Z(\GFM/n18720 ) );
XOR2_X2 \GFM/U4324  ( .A(\GFM/n19410 ), .B(\GFM/n19310 ), .Z(\GFM/n188 ) );
XOR2_X2 \GFM/U4323  ( .A(\GFM/n19620 ), .B(\GFM/n195 ), .Z(\GFM/n18900 ) );
XOR2_X2 \GFM/U4322  ( .A(\GFM/n198 ), .B(\GFM/n19700 ), .Z(\GFM/n19000 ) );
XOR2_X2 \GFM/U4321  ( .A(z_in[0]), .B(\GFM/n199 ), .Z(\GFM/n191 ) );
XOR2_X2 \GFM/U4320  ( .A(\GFM/N27 ), .B(\GFM/N28 ), .Z(\GFM/n192 ) );
XOR2_X2 \GFM/U4319  ( .A(\GFM/N24 ), .B(\GFM/N25 ), .Z(\GFM/n19310 ) );
XOR2_X2 \GFM/U4318  ( .A(\GFM/N20 ), .B(\GFM/N21 ), .Z(\GFM/n19410 ) );
XOR2_X2 \GFM/U4317  ( .A(\GFM/N16 ), .B(\GFM/N18 ), .Z(\GFM/n195 ) );
XOR2_X2 \GFM/U4316  ( .A(\GFM/N11 ), .B(\GFM/N15 ), .Z(\GFM/n19620 ) );
XOR2_X2 \GFM/U4315  ( .A(\GFM/N8 ), .B(\GFM/N10 ), .Z(\GFM/n19700 ) );
XOR2_X2 \GFM/U4314  ( .A(\GFM/N4 ), .B(\GFM/N7 ), .Z(\GFM/n198 ) );
XOR2_X2 \GFM/U4313  ( .A(\GFM/N1 ), .B(\GFM/N3 ), .Z(\GFM/n199 ) );
XOR2_X2 \GFM/U4312  ( .A(\GFM/n20100 ), .B(\GFM/n200 ), .Z(z_out[1]) );
XOR2_X2 \GFM/U4311  ( .A(\GFM/n203 ), .B(\GFM/n20200 ), .Z(\GFM/n200 ) );
XOR2_X2 \GFM/U4310  ( .A(\GFM/n205 ), .B(\GFM/n20410 ), .Z(\GFM/n20100 ) );
XOR2_X2 \GFM/U4309  ( .A(\GFM/n20720 ), .B(\GFM/n20600 ), .Z(\GFM/n20200 ));
XOR2_X2 \GFM/U4308  ( .A(\GFM/n209 ), .B(\GFM/n208 ), .Z(\GFM/n203 ) );
XOR2_X2 \GFM/U4307  ( .A(\GFM/n21100 ), .B(\GFM/n21000 ), .Z(\GFM/n20410 ));
XOR2_X2 \GFM/U4306  ( .A(\GFM/n21300 ), .B(\GFM/n212 ), .Z(\GFM/n205 ) );
XOR2_X2 \GFM/U4305  ( .A(z_in[1]), .B(\GFM/n2141 ), .Z(\GFM/n20600 ) );
XOR2_X2 \GFM/U4304  ( .A(\GFM/N58 ), .B(\GFM/N59 ), .Z(\GFM/n20720 ) );
XOR2_X2 \GFM/U4303  ( .A(\GFM/N55 ), .B(\GFM/N56 ), .Z(\GFM/n208 ) );
XOR2_X2 \GFM/U4302  ( .A(\GFM/N51 ), .B(\GFM/N52 ), .Z(\GFM/n209 ) );
XOR2_X2 \GFM/U4301  ( .A(\GFM/N47 ), .B(\GFM/N49 ), .Z(\GFM/n21000 ) );
XOR2_X2 \GFM/U4300  ( .A(\GFM/N42 ), .B(\GFM/N46 ), .Z(\GFM/n21100 ) );
XOR2_X2 \GFM/U4299  ( .A(\GFM/N39 ), .B(\GFM/N41 ), .Z(\GFM/n212 ) );
XOR2_X2 \GFM/U4298  ( .A(\GFM/N35 ), .B(\GFM/N38 ), .Z(\GFM/n21300 ) );
XOR2_X2 \GFM/U4297  ( .A(\GFM/N32 ), .B(\GFM/N34 ), .Z(\GFM/n2141 ) );
XOR2_X2 \GFM/U4296  ( .A(\GFM/n216 ), .B(\GFM/n215 ), .Z(z_out[2]) );
XOR2_X2 \GFM/U4295  ( .A(\GFM/n2182 ), .B(\GFM/n217 ), .Z(\GFM/n215 ) );
XOR2_X2 \GFM/U4294  ( .A(\GFM/n2200 ), .B(\GFM/n219 ), .Z(\GFM/n216 ) );
XOR2_X2 \GFM/U4293  ( .A(\GFM/n222 ), .B(\GFM/n2210 ), .Z(\GFM/n217 ) );
XOR2_X2 \GFM/U4292  ( .A(\GFM/n2241 ), .B(\GFM/n223 ), .Z(\GFM/n2182 ) );
XOR2_X2 \GFM/U4291  ( .A(\GFM/n226 ), .B(\GFM/n2251 ), .Z(\GFM/n219 ) );
XOR2_X2 \GFM/U4290  ( .A(\GFM/n2280 ), .B(\GFM/n2272 ), .Z(\GFM/n2200 ) );
XOR2_X2 \GFM/U4289  ( .A(z_in[2]), .B(\GFM/n229 ), .Z(\GFM/n2210 ) );
XOR2_X2 \GFM/U4288  ( .A(\GFM/N89 ), .B(\GFM/N90 ), .Z(\GFM/n222 ) );
XOR2_X2 \GFM/U4287  ( .A(\GFM/N86 ), .B(\GFM/N87 ), .Z(\GFM/n223 ) );
XOR2_X2 \GFM/U4286  ( .A(\GFM/N82 ), .B(\GFM/N83 ), .Z(\GFM/n2241 ) );
XOR2_X2 \GFM/U4285  ( .A(\GFM/N78 ), .B(\GFM/N80 ), .Z(\GFM/n2251 ) );
XOR2_X2 \GFM/U4284  ( .A(\GFM/N73 ), .B(\GFM/N77 ), .Z(\GFM/n226 ) );
XOR2_X2 \GFM/U4283  ( .A(\GFM/N70 ), .B(\GFM/N72 ), .Z(\GFM/n2272 ) );
XOR2_X2 \GFM/U4282  ( .A(\GFM/N66 ), .B(\GFM/N69 ), .Z(\GFM/n2280 ) );
XOR2_X2 \GFM/U4281  ( .A(\GFM/N63 ), .B(\GFM/N65 ), .Z(\GFM/n229 ) );
XOR2_X2 \GFM/U4280  ( .A(\GFM/n231 ), .B(\GFM/n230 ), .Z(z_out[3]) );
XOR2_X2 \GFM/U4279  ( .A(\GFM/n2330 ), .B(\GFM/n2320 ), .Z(\GFM/n230 ) );
XOR2_X2 \GFM/U4278  ( .A(\GFM/n2351 ), .B(\GFM/n234 ), .Z(\GFM/n231 ) );
XOR2_X2 \GFM/U4277  ( .A(\GFM/n2370 ), .B(\GFM/n236 ), .Z(\GFM/n2320 ) );
XOR2_X2 \GFM/U4276  ( .A(\GFM/n239 ), .B(\GFM/n2382 ), .Z(\GFM/n2330 ) );
XOR2_X2 \GFM/U4275  ( .A(\GFM/n24100 ), .B(\GFM/n240 ), .Z(\GFM/n234 ) );
XOR2_X2 \GFM/U4274  ( .A(\GFM/n243 ), .B(\GFM/n24200 ), .Z(\GFM/n2351 ) );
XOR2_X2 \GFM/U4273  ( .A(z_in[3]), .B(\GFM/n24400 ), .Z(\GFM/n236 ) );
XOR2_X2 \GFM/U4272  ( .A(\GFM/N120 ), .B(\GFM/N121 ), .Z(\GFM/n2370 ) );
XOR2_X2 \GFM/U4271  ( .A(\GFM/N117 ), .B(\GFM/N118 ), .Z(\GFM/n2382 ) );
XOR2_X2 \GFM/U4270  ( .A(\GFM/N113 ), .B(\GFM/N114 ), .Z(\GFM/n239 ) );
XOR2_X2 \GFM/U4269  ( .A(\GFM/N109 ), .B(\GFM/N111 ), .Z(\GFM/n240 ) );
XOR2_X2 \GFM/U4268  ( .A(\GFM/N104 ), .B(\GFM/N108 ), .Z(\GFM/n24100 ) );
XOR2_X2 \GFM/U4267  ( .A(\GFM/N101 ), .B(\GFM/N103 ), .Z(\GFM/n24200 ) );
XOR2_X2 \GFM/U4266  ( .A(\GFM/N97 ), .B(\GFM/N100 ), .Z(\GFM/n243 ) );
XOR2_X2 \GFM/U4265  ( .A(\GFM/N94 ), .B(\GFM/N96 ), .Z(\GFM/n24400 ) );
XOR2_X2 \GFM/U4264  ( .A(\GFM/n246 ), .B(\GFM/n24510 ), .Z(z_out[4]) );
XOR2_X2 \GFM/U4263  ( .A(\GFM/n248 ), .B(\GFM/n247 ), .Z(\GFM/n24510 ) );
XOR2_X2 \GFM/U4262  ( .A(\GFM/n250 ), .B(\GFM/n24920 ), .Z(\GFM/n246 ) );
XOR2_X2 \GFM/U4261  ( .A(\GFM/n25200 ), .B(\GFM/n25100 ), .Z(\GFM/n247 ) );
XOR2_X2 \GFM/U4260  ( .A(\GFM/n254 ), .B(\GFM/n253 ), .Z(\GFM/n248 ) );
XOR2_X2 \GFM/U4259  ( .A(\GFM/n25610 ), .B(\GFM/n25510 ), .Z(\GFM/n24920 ));
XOR2_X2 \GFM/U4258  ( .A(\GFM/n25820 ), .B(\GFM/n257 ), .Z(\GFM/n250 ) );
XOR2_X2 \GFM/U4257  ( .A(z_in[4]), .B(\GFM/n25900 ), .Z(\GFM/n25100 ) );
XOR2_X2 \GFM/U4256  ( .A(\GFM/N151 ), .B(\GFM/N152 ), .Z(\GFM/n25200 ) );
XOR2_X2 \GFM/U4255  ( .A(\GFM/N148 ), .B(\GFM/N149 ), .Z(\GFM/n253 ) );
XOR2_X2 \GFM/U4254  ( .A(\GFM/N144 ), .B(\GFM/N145 ), .Z(\GFM/n254 ) );
XOR2_X2 \GFM/U4253  ( .A(\GFM/N140 ), .B(\GFM/N142 ), .Z(\GFM/n25510 ) );
XOR2_X2 \GFM/U4252  ( .A(\GFM/N135 ), .B(\GFM/N139 ), .Z(\GFM/n25610 ) );
XOR2_X2 \GFM/U4251  ( .A(\GFM/N132 ), .B(\GFM/N134 ), .Z(\GFM/n257 ) );
XOR2_X2 \GFM/U4250  ( .A(\GFM/N128 ), .B(\GFM/N131 ), .Z(\GFM/n25820 ) );
XOR2_X2 \GFM/U4249  ( .A(\GFM/N125 ), .B(\GFM/N127 ), .Z(\GFM/n25900 ) );
XOR2_X2 \GFM/U4248  ( .A(\GFM/n261 ), .B(\GFM/n260 ), .Z(z_out[5]) );
XOR2_X2 \GFM/U4247  ( .A(\GFM/n26300 ), .B(\GFM/n262 ), .Z(\GFM/n260 ) );
XOR2_X2 \GFM/U4246  ( .A(\GFM/n265 ), .B(\GFM/n26400 ), .Z(\GFM/n261 ) );
XOR2_X2 \GFM/U4245  ( .A(\GFM/n267 ), .B(\GFM/n26610 ), .Z(\GFM/n262 ) );
XOR2_X2 \GFM/U4244  ( .A(\GFM/n26920 ), .B(\GFM/n26800 ), .Z(\GFM/n26300 ));
XOR2_X2 \GFM/U4243  ( .A(\GFM/n271 ), .B(\GFM/n270 ), .Z(\GFM/n26400 ) );
XOR2_X2 \GFM/U4242  ( .A(\GFM/n2730 ), .B(\GFM/n2720 ), .Z(\GFM/n265 ) );
XOR2_X2 \GFM/U4241  ( .A(z_in[5]), .B(\GFM/n274 ), .Z(\GFM/n26610 ) );
XOR2_X2 \GFM/U4240  ( .A(\GFM/N182 ), .B(\GFM/N183 ), .Z(\GFM/n267 ) );
XOR2_X2 \GFM/U4239  ( .A(\GFM/N179 ), .B(\GFM/N180 ), .Z(\GFM/n26800 ) );
XOR2_X2 \GFM/U4238  ( .A(\GFM/N175 ), .B(\GFM/N176 ), .Z(\GFM/n26920 ) );
XOR2_X2 \GFM/U4237  ( .A(\GFM/N171 ), .B(\GFM/N173 ), .Z(\GFM/n270 ) );
XOR2_X2 \GFM/U4236  ( .A(\GFM/N166 ), .B(\GFM/N170 ), .Z(\GFM/n271 ) );
XOR2_X2 \GFM/U4235  ( .A(\GFM/N163 ), .B(\GFM/N165 ), .Z(\GFM/n2720 ) );
XOR2_X2 \GFM/U4234  ( .A(\GFM/N159 ), .B(\GFM/N162 ), .Z(\GFM/n2730 ) );
XOR2_X2 \GFM/U4233  ( .A(\GFM/N156 ), .B(\GFM/N158 ), .Z(\GFM/n274 ) );
XOR2_X2 \GFM/U4232  ( .A(\GFM/n2761 ), .B(\GFM/n2750 ), .Z(z_out[6]) );
XOR2_X2 \GFM/U4231  ( .A(\GFM/n278 ), .B(\GFM/n277 ), .Z(\GFM/n2750 ) );
XOR2_X2 \GFM/U4230  ( .A(\GFM/n2802 ), .B(\GFM/n279 ), .Z(\GFM/n2761 ) );
XOR2_X2 \GFM/U4229  ( .A(\GFM/n2820 ), .B(\GFM/n281 ), .Z(\GFM/n277 ) );
XOR2_X2 \GFM/U4228  ( .A(\GFM/n284 ), .B(\GFM/n2830 ), .Z(\GFM/n278 ) );
XOR2_X2 \GFM/U4227  ( .A(\GFM/n2861 ), .B(\GFM/n285 ), .Z(\GFM/n279 ) );
XOR2_X2 \GFM/U4226  ( .A(\GFM/n288 ), .B(\GFM/n2871 ), .Z(\GFM/n2802 ) );
XOR2_X2 \GFM/U4225  ( .A(z_in[6]), .B(\GFM/n2892 ), .Z(\GFM/n281 ) );
XOR2_X2 \GFM/U4224  ( .A(\GFM/N213 ), .B(\GFM/N214 ), .Z(\GFM/n2820 ) );
XOR2_X2 \GFM/U4223  ( .A(\GFM/N210 ), .B(\GFM/N211 ), .Z(\GFM/n2830 ) );
XOR2_X2 \GFM/U4222  ( .A(\GFM/N206 ), .B(\GFM/N207 ), .Z(\GFM/n284 ) );
XOR2_X2 \GFM/U4221  ( .A(\GFM/N202 ), .B(\GFM/N204 ), .Z(\GFM/n285 ) );
XOR2_X2 \GFM/U4220  ( .A(\GFM/N197 ), .B(\GFM/N201 ), .Z(\GFM/n2861 ) );
XOR2_X2 \GFM/U4219  ( .A(\GFM/N194 ), .B(\GFM/N196 ), .Z(\GFM/n2871 ) );
XOR2_X2 \GFM/U4218  ( .A(\GFM/N190 ), .B(\GFM/N193 ), .Z(\GFM/n288 ) );
XOR2_X2 \GFM/U4217  ( .A(\GFM/N187 ), .B(\GFM/N189 ), .Z(\GFM/n2892 ) );
XOR2_X2 \GFM/U4216  ( .A(\GFM/n291 ), .B(\GFM/n2900 ), .Z(z_out[7]) );
XOR2_X2 \GFM/U4215  ( .A(\GFM/n293 ), .B(\GFM/n292 ), .Z(\GFM/n2900 ) );
XOR2_X2 \GFM/U4214  ( .A(\GFM/n2950 ), .B(\GFM/n2940 ), .Z(\GFM/n291 ) );
XOR2_X2 \GFM/U4213  ( .A(\GFM/n2971 ), .B(\GFM/n296 ), .Z(\GFM/n292 ) );
XOR2_X2 \GFM/U4212  ( .A(\GFM/n2990 ), .B(\GFM/n298 ), .Z(\GFM/n293 ) );
XOR2_X2 \GFM/U4211  ( .A(\GFM/n301 ), .B(\GFM/n3002 ), .Z(\GFM/n2940 ) );
XOR2_X2 \GFM/U4210  ( .A(\GFM/n3030 ), .B(\GFM/n302 ), .Z(\GFM/n2950 ) );
XOR2_X2 \GFM/U4209  ( .A(z_in[7]), .B(\GFM/n3040 ), .Z(\GFM/n296 ) );
XOR2_X2 \GFM/U4208  ( .A(\GFM/N244 ), .B(\GFM/N245 ), .Z(\GFM/n2971 ) );
XOR2_X2 \GFM/U4207  ( .A(\GFM/N241 ), .B(\GFM/N242 ), .Z(\GFM/n298 ) );
XOR2_X2 \GFM/U4206  ( .A(\GFM/N237 ), .B(\GFM/N238 ), .Z(\GFM/n2990 ) );
XOR2_X2 \GFM/U4205  ( .A(\GFM/N233 ), .B(\GFM/N235 ), .Z(\GFM/n3002 ) );
XOR2_X2 \GFM/U4204  ( .A(\GFM/N228 ), .B(\GFM/N232 ), .Z(\GFM/n301 ) );
XOR2_X2 \GFM/U4203  ( .A(\GFM/N225 ), .B(\GFM/N227 ), .Z(\GFM/n302 ) );
XOR2_X2 \GFM/U4202  ( .A(\GFM/N221 ), .B(\GFM/N224 ), .Z(\GFM/n3030 ) );
XOR2_X2 \GFM/U4201  ( .A(\GFM/N218 ), .B(\GFM/N220 ), .Z(\GFM/n3040 ) );
XOR2_X2 \GFM/U4200  ( .A(\GFM/n3060 ), .B(\GFM/n305 ), .Z(z_out[8]) );
XOR2_X2 \GFM/U4199  ( .A(\GFM/n308 ), .B(\GFM/n3071 ), .Z(\GFM/n305 ) );
XOR2_X2 \GFM/U4198  ( .A(\GFM/n310 ), .B(\GFM/n309 ), .Z(\GFM/n3060 ) );
XOR2_X2 \GFM/U4197  ( .A(\GFM/n312 ), .B(\GFM/n3112 ), .Z(\GFM/n3071 ) );
XOR2_X2 \GFM/U4196  ( .A(\GFM/n3140 ), .B(\GFM/n3130 ), .Z(\GFM/n308 ) );
XOR2_X2 \GFM/U4195  ( .A(\GFM/n316 ), .B(\GFM/n315 ), .Z(\GFM/n309 ) );
XOR2_X2 \GFM/U4194  ( .A(\GFM/n3181 ), .B(\GFM/n3171 ), .Z(\GFM/n310 ) );
XOR2_X2 \GFM/U4193  ( .A(z_in[8]), .B(\GFM/n319 ), .Z(\GFM/n3112 ) );
XOR2_X2 \GFM/U4192  ( .A(\GFM/N275 ), .B(\GFM/N276 ), .Z(\GFM/n312 ) );
XOR2_X2 \GFM/U4191  ( .A(\GFM/N272 ), .B(\GFM/N273 ), .Z(\GFM/n3130 ) );
XOR2_X2 \GFM/U4190  ( .A(\GFM/N268 ), .B(\GFM/N269 ), .Z(\GFM/n3140 ) );
XOR2_X2 \GFM/U4189  ( .A(\GFM/N264 ), .B(\GFM/N266 ), .Z(\GFM/n315 ) );
XOR2_X2 \GFM/U4188  ( .A(\GFM/N259 ), .B(\GFM/N263 ), .Z(\GFM/n316 ) );
XOR2_X2 \GFM/U4187  ( .A(\GFM/N256 ), .B(\GFM/N258 ), .Z(\GFM/n3171 ) );
XOR2_X2 \GFM/U4186  ( .A(\GFM/N252 ), .B(\GFM/N255 ), .Z(\GFM/n3181 ) );
XOR2_X2 \GFM/U4185  ( .A(\GFM/N249 ), .B(\GFM/N251 ), .Z(\GFM/n319 ) );
XOR2_X2 \GFM/U4184  ( .A(\GFM/n3210 ), .B(\GFM/n3202 ), .Z(z_out[9]) );
XOR2_X2 \GFM/U4183  ( .A(\GFM/n323 ), .B(\GFM/n322 ), .Z(\GFM/n3202 ) );
XOR2_X2 \GFM/U4182  ( .A(\GFM/n3250 ), .B(\GFM/n324 ), .Z(\GFM/n3210 ) );
XOR2_X2 \GFM/U4181  ( .A(\GFM/n327 ), .B(\GFM/n3260 ), .Z(\GFM/n322 ) );
XOR2_X2 \GFM/U4180  ( .A(\GFM/n329 ), .B(\GFM/n3281 ), .Z(\GFM/n323 ) );
XOR2_X2 \GFM/U4179  ( .A(\GFM/n3310 ), .B(\GFM/n3300 ), .Z(\GFM/n324 ) );
XOR2_X2 \GFM/U4178  ( .A(\GFM/n333 ), .B(\GFM/n332 ), .Z(\GFM/n3250 ) );
XOR2_X2 \GFM/U4177  ( .A(z_in[9]), .B(\GFM/n3342 ), .Z(\GFM/n3260 ) );
XOR2_X2 \GFM/U4176  ( .A(\GFM/N306 ), .B(\GFM/N307 ), .Z(\GFM/n327 ) );
XOR2_X2 \GFM/U4175  ( .A(\GFM/N303 ), .B(\GFM/N304 ), .Z(\GFM/n3281 ) );
XOR2_X2 \GFM/U4174  ( .A(\GFM/N299 ), .B(\GFM/N300 ), .Z(\GFM/n329 ) );
XOR2_X2 \GFM/U4173  ( .A(\GFM/N295 ), .B(\GFM/N297 ), .Z(\GFM/n3300 ) );
XOR2_X2 \GFM/U4172  ( .A(\GFM/N290 ), .B(\GFM/N294 ), .Z(\GFM/n3310 ) );
XOR2_X2 \GFM/U4171  ( .A(\GFM/N287 ), .B(\GFM/N289 ), .Z(\GFM/n332 ) );
XOR2_X2 \GFM/U4170  ( .A(\GFM/N283 ), .B(\GFM/N286 ), .Z(\GFM/n333 ) );
XOR2_X2 \GFM/U4169  ( .A(\GFM/N280 ), .B(\GFM/N282 ), .Z(\GFM/n3342 ) );
XOR2_X2 \GFM/U4168  ( .A(\GFM/n336 ), .B(\GFM/n3350 ), .Z(z_out[10]) );
XOR2_X2 \GFM/U4167  ( .A(\GFM/n3381 ), .B(\GFM/n3370 ), .Z(\GFM/n3350 ) );
XOR2_X2 \GFM/U4166  ( .A(\GFM/n340 ), .B(\GFM/n339 ), .Z(\GFM/n336 ) );
XOR2_X2 \GFM/U4165  ( .A(\GFM/n3420 ), .B(\GFM/n341 ), .Z(\GFM/n3370 ) );
XOR2_X2 \GFM/U4164  ( .A(\GFM/n3440 ), .B(\GFM/n343 ), .Z(\GFM/n3381 ) );
XOR2_X2 \GFM/U4163  ( .A(\GFM/n346 ), .B(\GFM/n3451 ), .Z(\GFM/n339 ) );
XOR2_X2 \GFM/U4162  ( .A(\GFM/n3480 ), .B(\GFM/n347 ), .Z(\GFM/n340 ) );
XOR2_X2 \GFM/U4161  ( .A(z_in[10]), .B(\GFM/n3490 ), .Z(\GFM/n341 ) );
XOR2_X2 \GFM/U4160  ( .A(\GFM/N337 ), .B(\GFM/N338 ), .Z(\GFM/n3420 ) );
XOR2_X2 \GFM/U4159  ( .A(\GFM/N334 ), .B(\GFM/N335 ), .Z(\GFM/n343 ) );
XOR2_X2 \GFM/U4158  ( .A(\GFM/N330 ), .B(\GFM/N331 ), .Z(\GFM/n3440 ) );
XOR2_X2 \GFM/U4157  ( .A(\GFM/N326 ), .B(\GFM/N328 ), .Z(\GFM/n3451 ) );
XOR2_X2 \GFM/U4156  ( .A(\GFM/N321 ), .B(\GFM/N325 ), .Z(\GFM/n346 ) );
XOR2_X2 \GFM/U4155  ( .A(\GFM/N318 ), .B(\GFM/N320 ), .Z(\GFM/n347 ) );
XOR2_X2 \GFM/U4154  ( .A(\GFM/N314 ), .B(\GFM/N317 ), .Z(\GFM/n3480 ) );
XOR2_X2 \GFM/U4153  ( .A(\GFM/N311 ), .B(\GFM/N313 ), .Z(\GFM/n3490 ) );
XOR2_X2 \GFM/U4152  ( .A(\GFM/n3510 ), .B(\GFM/n350 ), .Z(z_out[11]) );
XOR2_X2 \GFM/U4151  ( .A(\GFM/n353 ), .B(\GFM/n3520 ), .Z(\GFM/n350 ) );
XOR2_X2 \GFM/U4150  ( .A(\GFM/n355 ), .B(\GFM/n354 ), .Z(\GFM/n3510 ) );
XOR2_X2 \GFM/U4149  ( .A(\GFM/n3570 ), .B(\GFM/n3560 ), .Z(\GFM/n3520 ) );
XOR2_X2 \GFM/U4148  ( .A(\GFM/n3590 ), .B(\GFM/n358 ), .Z(\GFM/n353 ) );
XOR2_X2 \GFM/U4147  ( .A(\GFM/n3610 ), .B(\GFM/n360 ), .Z(\GFM/n354 ) );
XOR2_X2 \GFM/U4146  ( .A(\GFM/n363 ), .B(\GFM/n3621 ), .Z(\GFM/n355 ) );
XOR2_X2 \GFM/U4145  ( .A(z_in[11]), .B(\GFM/n364 ), .Z(\GFM/n3560 ) );
XOR2_X2 \GFM/U4144  ( .A(\GFM/N368 ), .B(\GFM/N369 ), .Z(\GFM/n3570 ) );
XOR2_X2 \GFM/U4143  ( .A(\GFM/N365 ), .B(\GFM/N366 ), .Z(\GFM/n358 ) );
XOR2_X2 \GFM/U4142  ( .A(\GFM/N361 ), .B(\GFM/N362 ), .Z(\GFM/n3590 ) );
XOR2_X2 \GFM/U4141  ( .A(\GFM/N357 ), .B(\GFM/N359 ), .Z(\GFM/n360 ) );
XOR2_X2 \GFM/U4140  ( .A(\GFM/N352 ), .B(\GFM/N356 ), .Z(\GFM/n3610 ) );
XOR2_X2 \GFM/U4139  ( .A(\GFM/N349 ), .B(\GFM/N351 ), .Z(\GFM/n3621 ) );
XOR2_X2 \GFM/U4138  ( .A(\GFM/N345 ), .B(\GFM/N348 ), .Z(\GFM/n363 ) );
XOR2_X2 \GFM/U4137  ( .A(\GFM/N342 ), .B(\GFM/N344 ), .Z(\GFM/n364 ) );
XOR2_X2 \GFM/U4136  ( .A(\GFM/n3660 ), .B(\GFM/n3650 ), .Z(z_out[12]) );
XOR2_X2 \GFM/U4135  ( .A(\GFM/n3680 ), .B(\GFM/n367 ), .Z(\GFM/n3650 ) );
XOR2_X2 \GFM/U4134  ( .A(\GFM/n370 ), .B(\GFM/n3691 ), .Z(\GFM/n3660 ) );
XOR2_X2 \GFM/U4133  ( .A(\GFM/n372 ), .B(\GFM/n371 ), .Z(\GFM/n367 ) );
XOR2_X2 \GFM/U4132  ( .A(\GFM/n374 ), .B(\GFM/n3730 ), .Z(\GFM/n3680 ) );
XOR2_X2 \GFM/U4131  ( .A(\GFM/n3760 ), .B(\GFM/n3751 ), .Z(\GFM/n3691 ) );
XOR2_X2 \GFM/U4130  ( .A(\GFM/n378 ), .B(\GFM/n377 ), .Z(\GFM/n370 ) );
XOR2_X2 \GFM/U4129  ( .A(z_in[12]), .B(\GFM/n3790 ), .Z(\GFM/n371 ) );
XOR2_X2 \GFM/U4128  ( .A(\GFM/N399 ), .B(\GFM/N400 ), .Z(\GFM/n372 ) );
XOR2_X2 \GFM/U4127  ( .A(\GFM/N396 ), .B(\GFM/N397 ), .Z(\GFM/n3730 ) );
XOR2_X2 \GFM/U4126  ( .A(\GFM/N392 ), .B(\GFM/N393 ), .Z(\GFM/n374 ) );
XOR2_X2 \GFM/U4125  ( .A(\GFM/N388 ), .B(\GFM/N390 ), .Z(\GFM/n3751 ) );
XOR2_X2 \GFM/U4124  ( .A(\GFM/N383 ), .B(\GFM/N387 ), .Z(\GFM/n3760 ) );
XOR2_X2 \GFM/U4123  ( .A(\GFM/N380 ), .B(\GFM/N382 ), .Z(\GFM/n377 ) );
XOR2_X2 \GFM/U4122  ( .A(\GFM/N376 ), .B(\GFM/N379 ), .Z(\GFM/n378 ) );
XOR2_X2 \GFM/U4121  ( .A(\GFM/N373 ), .B(\GFM/N375 ), .Z(\GFM/n3790 ) );
XOR2_X2 \GFM/U4120  ( .A(\GFM/n381 ), .B(\GFM/n3800 ), .Z(z_out[13]) );
XOR2_X2 \GFM/U4119  ( .A(\GFM/n3830 ), .B(\GFM/n3820 ), .Z(\GFM/n3800 ) );
XOR2_X2 \GFM/U4118  ( .A(\GFM/n385 ), .B(\GFM/n384 ), .Z(\GFM/n381 ) );
XOR2_X2 \GFM/U4117  ( .A(\GFM/n3870 ), .B(\GFM/n386 ), .Z(\GFM/n3820 ) );
XOR2_X2 \GFM/U4116  ( .A(\GFM/n389 ), .B(\GFM/n3880 ), .Z(\GFM/n3830 ) );
XOR2_X2 \GFM/U4115  ( .A(\GFM/n391 ), .B(\GFM/n3900 ), .Z(\GFM/n384 ) );
XOR2_X2 \GFM/U4114  ( .A(\GFM/n3930 ), .B(\GFM/n3920 ), .Z(\GFM/n385 ) );
XOR2_X2 \GFM/U4113  ( .A(z_in[13]), .B(\GFM/n394 ), .Z(\GFM/n386 ) );
XOR2_X2 \GFM/U4112  ( .A(\GFM/N430 ), .B(\GFM/N431 ), .Z(\GFM/n3870 ) );
XOR2_X2 \GFM/U4111  ( .A(\GFM/N427 ), .B(\GFM/N428 ), .Z(\GFM/n3880 ) );
XOR2_X2 \GFM/U4110  ( .A(\GFM/N423 ), .B(\GFM/N424 ), .Z(\GFM/n389 ) );
XOR2_X2 \GFM/U4109  ( .A(\GFM/N419 ), .B(\GFM/N421 ), .Z(\GFM/n3900 ) );
XOR2_X2 \GFM/U4108  ( .A(\GFM/N414 ), .B(\GFM/N418 ), .Z(\GFM/n391 ) );
XOR2_X2 \GFM/U4107  ( .A(\GFM/N411 ), .B(\GFM/N413 ), .Z(\GFM/n3920 ) );
XOR2_X2 \GFM/U4106  ( .A(\GFM/N407 ), .B(\GFM/N410 ), .Z(\GFM/n3930 ) );
XOR2_X2 \GFM/U4105  ( .A(\GFM/N404 ), .B(\GFM/N406 ), .Z(\GFM/n394 ) );
XOR2_X2 \GFM/U4104  ( .A(\GFM/n3960 ), .B(\GFM/n395 ), .Z(z_out[14]) );
XOR2_X2 \GFM/U4103  ( .A(\GFM/n398 ), .B(\GFM/n3970 ), .Z(\GFM/n395 ) );
XOR2_X2 \GFM/U4102  ( .A(\GFM/n4000 ), .B(\GFM/n3991 ), .Z(\GFM/n3960 ) );
XOR2_X2 \GFM/U4101  ( .A(\GFM/n402 ), .B(\GFM/n401 ), .Z(\GFM/n3970 ) );
XOR2_X2 \GFM/U4100  ( .A(\GFM/n4040 ), .B(\GFM/n403 ), .Z(\GFM/n398 ) );
XOR2_X2 \GFM/U4099  ( .A(\GFM/n4060 ), .B(\GFM/n405 ), .Z(\GFM/n3991 ) );
XOR2_X2 \GFM/U4098  ( .A(\GFM/n408 ), .B(\GFM/n4070 ), .Z(\GFM/n4000 ) );
XOR2_X2 \GFM/U4097  ( .A(z_in[14]), .B(\GFM/n409 ), .Z(\GFM/n401 ) );
XOR2_X2 \GFM/U4096  ( .A(\GFM/N461 ), .B(\GFM/N462 ), .Z(\GFM/n402 ) );
XOR2_X2 \GFM/U4095  ( .A(\GFM/N458 ), .B(\GFM/N459 ), .Z(\GFM/n403 ) );
XOR2_X2 \GFM/U4094  ( .A(\GFM/N454 ), .B(\GFM/N455 ), .Z(\GFM/n4040 ) );
XOR2_X2 \GFM/U4093  ( .A(\GFM/N450 ), .B(\GFM/N452 ), .Z(\GFM/n405 ) );
XOR2_X2 \GFM/U4092  ( .A(\GFM/N445 ), .B(\GFM/N449 ), .Z(\GFM/n4060 ) );
XOR2_X2 \GFM/U4091  ( .A(\GFM/N442 ), .B(\GFM/N444 ), .Z(\GFM/n4070 ) );
XOR2_X2 \GFM/U4090  ( .A(\GFM/N438 ), .B(\GFM/N441 ), .Z(\GFM/n408 ) );
XOR2_X2 \GFM/U4089  ( .A(\GFM/N435 ), .B(\GFM/N437 ), .Z(\GFM/n409 ) );
XOR2_X2 \GFM/U4088  ( .A(\GFM/n4110 ), .B(\GFM/n4100 ), .Z(z_out[15]) );
XOR2_X2 \GFM/U4087  ( .A(\GFM/n4130 ), .B(\GFM/n412 ), .Z(\GFM/n4100 ) );
XOR2_X2 \GFM/U4086  ( .A(\GFM/n415 ), .B(\GFM/n4140 ), .Z(\GFM/n4110 ) );
XOR2_X2 \GFM/U4085  ( .A(\GFM/n417 ), .B(\GFM/n416 ), .Z(\GFM/n412 ) );
XOR2_X2 \GFM/U4084  ( .A(\GFM/n4190 ), .B(\GFM/n4180 ), .Z(\GFM/n4130 ) );
XOR2_X2 \GFM/U4083  ( .A(\GFM/n4211 ), .B(\GFM/n420 ), .Z(\GFM/n4140 ) );
XOR2_X2 \GFM/U4082  ( .A(\GFM/n4230 ), .B(\GFM/n422 ), .Z(\GFM/n415 ) );
XOR2_X2 \GFM/U4081  ( .A(z_in[15]), .B(\GFM/n4241 ), .Z(\GFM/n416 ) );
XOR2_X2 \GFM/U4080  ( .A(\GFM/N492 ), .B(\GFM/N493 ), .Z(\GFM/n417 ) );
XOR2_X2 \GFM/U4079  ( .A(\GFM/N489 ), .B(\GFM/N490 ), .Z(\GFM/n4180 ) );
XOR2_X2 \GFM/U4078  ( .A(\GFM/N485 ), .B(\GFM/N486 ), .Z(\GFM/n4190 ) );
XOR2_X2 \GFM/U4077  ( .A(\GFM/N481 ), .B(\GFM/N483 ), .Z(\GFM/n420 ) );
XOR2_X2 \GFM/U4076  ( .A(\GFM/N476 ), .B(\GFM/N480 ), .Z(\GFM/n4211 ) );
XOR2_X2 \GFM/U4075  ( .A(\GFM/N473 ), .B(\GFM/N475 ), .Z(\GFM/n422 ) );
XOR2_X2 \GFM/U4074  ( .A(\GFM/N469 ), .B(\GFM/N472 ), .Z(\GFM/n4230 ) );
XOR2_X2 \GFM/U4073  ( .A(\GFM/N466 ), .B(\GFM/N468 ), .Z(\GFM/n4241 ) );
XOR2_X2 \GFM/U4072  ( .A(\GFM/n426 ), .B(\GFM/n425 ), .Z(z_out[16]) );
XOR2_X2 \GFM/U4071  ( .A(\GFM/n4280 ), .B(\GFM/n4270 ), .Z(\GFM/n425 ) );
XOR2_X2 \GFM/U4070  ( .A(\GFM/n4301 ), .B(\GFM/n429 ), .Z(\GFM/n426 ) );
XOR2_X2 \GFM/U4069  ( .A(\GFM/n432 ), .B(\GFM/n4310 ), .Z(\GFM/n4270 ) );
XOR2_X2 \GFM/U4068  ( .A(\GFM/n434 ), .B(\GFM/n433 ), .Z(\GFM/n4280 ) );
XOR2_X2 \GFM/U4067  ( .A(\GFM/n436 ), .B(\GFM/n4350 ), .Z(\GFM/n429 ) );
XOR2_X2 \GFM/U4066  ( .A(\GFM/n4380 ), .B(\GFM/n4370 ), .Z(\GFM/n4301 ) );
XOR2_X2 \GFM/U4065  ( .A(z_in[16]), .B(\GFM/n439 ), .Z(\GFM/n4310 ) );
XOR2_X2 \GFM/U4064  ( .A(\GFM/N523 ), .B(\GFM/N524 ), .Z(\GFM/n432 ) );
XOR2_X2 \GFM/U4063  ( .A(\GFM/N520 ), .B(\GFM/N521 ), .Z(\GFM/n433 ) );
XOR2_X2 \GFM/U4062  ( .A(\GFM/N516 ), .B(\GFM/N517 ), .Z(\GFM/n434 ) );
XOR2_X2 \GFM/U4061  ( .A(\GFM/N512 ), .B(\GFM/N514 ), .Z(\GFM/n4350 ) );
XOR2_X2 \GFM/U4060  ( .A(\GFM/N507 ), .B(\GFM/N511 ), .Z(\GFM/n436 ) );
XOR2_X2 \GFM/U4059  ( .A(\GFM/N504 ), .B(\GFM/N506 ), .Z(\GFM/n4370 ) );
XOR2_X2 \GFM/U4058  ( .A(\GFM/N500 ), .B(\GFM/N503 ), .Z(\GFM/n4380 ) );
XOR2_X2 \GFM/U4057  ( .A(\GFM/N497 ), .B(\GFM/N499 ), .Z(\GFM/n439 ) );
XOR2_X2 \GFM/U4056  ( .A(\GFM/n4410 ), .B(\GFM/n440 ), .Z(z_out[17]) );
XOR2_X2 \GFM/U4055  ( .A(\GFM/n443 ), .B(\GFM/n4420 ), .Z(\GFM/n440 ) );
XOR2_X2 \GFM/U4054  ( .A(\GFM/n4450 ), .B(\GFM/n4440 ), .Z(\GFM/n4410 ) );
XOR2_X2 \GFM/U4053  ( .A(\GFM/n447 ), .B(\GFM/n446 ), .Z(\GFM/n4420 ) );
XOR2_X2 \GFM/U4052  ( .A(\GFM/n4490 ), .B(\GFM/n448 ), .Z(\GFM/n443 ) );
XOR2_X2 \GFM/U4051  ( .A(\GFM/n451 ), .B(\GFM/n4500 ), .Z(\GFM/n4440 ) );
XOR2_X2 \GFM/U4050  ( .A(\GFM/n453 ), .B(\GFM/n4520 ), .Z(\GFM/n4450 ) );
XOR2_X2 \GFM/U4049  ( .A(z_in[17]), .B(\GFM/n4540 ), .Z(\GFM/n446 ) );
XOR2_X2 \GFM/U4048  ( .A(\GFM/N554 ), .B(\GFM/N555 ), .Z(\GFM/n447 ) );
XOR2_X2 \GFM/U4047  ( .A(\GFM/N551 ), .B(\GFM/N552 ), .Z(\GFM/n448 ) );
XOR2_X2 \GFM/U4046  ( .A(\GFM/N547 ), .B(\GFM/N548 ), .Z(\GFM/n4490 ) );
XOR2_X2 \GFM/U4045  ( .A(\GFM/N543 ), .B(\GFM/N545 ), .Z(\GFM/n4500 ) );
XOR2_X2 \GFM/U4044  ( .A(\GFM/N538 ), .B(\GFM/N542 ), .Z(\GFM/n451 ) );
XOR2_X2 \GFM/U4043  ( .A(\GFM/N535 ), .B(\GFM/N537 ), .Z(\GFM/n4520 ) );
XOR2_X2 \GFM/U4042  ( .A(\GFM/N531 ), .B(\GFM/N534 ), .Z(\GFM/n453 ) );
XOR2_X2 \GFM/U4041  ( .A(\GFM/N528 ), .B(\GFM/N530 ), .Z(\GFM/n4540 ) );
XOR2_X2 \GFM/U4040  ( .A(\GFM/n456 ), .B(\GFM/n4550 ), .Z(z_out[18]) );
XOR2_X2 \GFM/U4039  ( .A(\GFM/n4580 ), .B(\GFM/n457 ), .Z(\GFM/n4550 ) );
XOR2_X2 \GFM/U4038  ( .A(\GFM/n460 ), .B(\GFM/n4590 ), .Z(\GFM/n456 ) );
XOR2_X2 \GFM/U4037  ( .A(\GFM/n4620 ), .B(\GFM/n4610 ), .Z(\GFM/n457 ) );
XOR2_X2 \GFM/U4036  ( .A(\GFM/n464 ), .B(\GFM/n463 ), .Z(\GFM/n4580 ) );
XOR2_X2 \GFM/U4035  ( .A(\GFM/n4660 ), .B(\GFM/n465 ), .Z(\GFM/n4590 ) );
XOR2_X2 \GFM/U4034  ( .A(\GFM/n4680 ), .B(\GFM/n467 ), .Z(\GFM/n460 ) );
XOR2_X2 \GFM/U4033  ( .A(z_in[18]), .B(\GFM/n4690 ), .Z(\GFM/n4610 ) );
XOR2_X2 \GFM/U4032  ( .A(\GFM/N585 ), .B(\GFM/N586 ), .Z(\GFM/n4620 ) );
XOR2_X2 \GFM/U4031  ( .A(\GFM/N582 ), .B(\GFM/N583 ), .Z(\GFM/n463 ) );
XOR2_X2 \GFM/U4030  ( .A(\GFM/N578 ), .B(\GFM/N579 ), .Z(\GFM/n464 ) );
XOR2_X2 \GFM/U4029  ( .A(\GFM/N574 ), .B(\GFM/N576 ), .Z(\GFM/n465 ) );
XOR2_X2 \GFM/U4028  ( .A(\GFM/N569 ), .B(\GFM/N573 ), .Z(\GFM/n4660 ) );
XOR2_X2 \GFM/U4027  ( .A(\GFM/N566 ), .B(\GFM/N568 ), .Z(\GFM/n467 ) );
XOR2_X2 \GFM/U4026  ( .A(\GFM/N562 ), .B(\GFM/N565 ), .Z(\GFM/n4680 ) );
XOR2_X2 \GFM/U4025  ( .A(\GFM/N559 ), .B(\GFM/N561 ), .Z(\GFM/n4690 ) );
XOR2_X2 \GFM/U4024  ( .A(\GFM/n471 ), .B(\GFM/n470 ), .Z(z_out[19]) );
XOR2_X2 \GFM/U4023  ( .A(\GFM/n4730 ), .B(\GFM/n4720 ), .Z(\GFM/n470 ) );
XOR2_X2 \GFM/U4022  ( .A(\GFM/n4750 ), .B(\GFM/n474 ), .Z(\GFM/n471 ) );
XOR2_X2 \GFM/U4021  ( .A(\GFM/n477 ), .B(\GFM/n4760 ), .Z(\GFM/n4720 ) );
XOR2_X2 \GFM/U4020  ( .A(\GFM/n479 ), .B(\GFM/n478 ), .Z(\GFM/n4730 ) );
XOR2_X2 \GFM/U4019  ( .A(\GFM/n4810 ), .B(\GFM/n4800 ), .Z(\GFM/n474 ) );
XOR2_X2 \GFM/U4018  ( .A(\GFM/n4830 ), .B(\GFM/n482 ), .Z(\GFM/n4750 ) );
XOR2_X2 \GFM/U4017  ( .A(z_in[19]), .B(\GFM/n484 ), .Z(\GFM/n4760 ) );
XOR2_X2 \GFM/U4016  ( .A(\GFM/N616 ), .B(\GFM/N617 ), .Z(\GFM/n477 ) );
XOR2_X2 \GFM/U4015  ( .A(\GFM/N613 ), .B(\GFM/N614 ), .Z(\GFM/n478 ) );
XOR2_X2 \GFM/U4014  ( .A(\GFM/N609 ), .B(\GFM/N610 ), .Z(\GFM/n479 ) );
XOR2_X2 \GFM/U4013  ( .A(\GFM/N605 ), .B(\GFM/N607 ), .Z(\GFM/n4800 ) );
XOR2_X2 \GFM/U4012  ( .A(\GFM/N600 ), .B(\GFM/N604 ), .Z(\GFM/n4810 ) );
XOR2_X2 \GFM/U4011  ( .A(\GFM/N597 ), .B(\GFM/N599 ), .Z(\GFM/n482 ) );
XOR2_X2 \GFM/U4010  ( .A(\GFM/N593 ), .B(\GFM/N596 ), .Z(\GFM/n4830 ) );
XOR2_X2 \GFM/U4009  ( .A(\GFM/N590 ), .B(\GFM/N592 ), .Z(\GFM/n484 ) );
XOR2_X2 \GFM/U4008  ( .A(\GFM/n4860 ), .B(\GFM/n4850 ), .Z(z_out[20]) );
XOR2_X2 \GFM/U4007  ( .A(\GFM/n488 ), .B(\GFM/n487 ), .Z(\GFM/n4850 ) );
XOR2_X2 \GFM/U4006  ( .A(\GFM/n4900 ), .B(\GFM/n4890 ), .Z(\GFM/n4860 ) );
XOR2_X2 \GFM/U4005  ( .A(\GFM/n4920 ), .B(\GFM/n491 ), .Z(\GFM/n487 ) );
XOR2_X2 \GFM/U4004  ( .A(\GFM/n494 ), .B(\GFM/n4930 ), .Z(\GFM/n488 ) );
XOR2_X2 \GFM/U4003  ( .A(\GFM/n496 ), .B(\GFM/n495 ), .Z(\GFM/n4890 ) );
XOR2_X2 \GFM/U4002  ( .A(\GFM/n498 ), .B(\GFM/n4970 ), .Z(\GFM/n4900 ) );
XOR2_X2 \GFM/U4001  ( .A(z_in[20]), .B(\GFM/n4990 ), .Z(\GFM/n491 ) );
XOR2_X2 \GFM/U4000  ( .A(\GFM/N647 ), .B(\GFM/N648 ), .Z(\GFM/n4920 ) );
XOR2_X2 \GFM/U3999  ( .A(\GFM/N644 ), .B(\GFM/N645 ), .Z(\GFM/n4930 ) );
XOR2_X2 \GFM/U3998  ( .A(\GFM/N640 ), .B(\GFM/N641 ), .Z(\GFM/n494 ) );
XOR2_X2 \GFM/U3997  ( .A(\GFM/N636 ), .B(\GFM/N638 ), .Z(\GFM/n495 ) );
XOR2_X2 \GFM/U3996  ( .A(\GFM/N631 ), .B(\GFM/N635 ), .Z(\GFM/n496 ) );
XOR2_X2 \GFM/U3995  ( .A(\GFM/N628 ), .B(\GFM/N630 ), .Z(\GFM/n4970 ) );
XOR2_X2 \GFM/U3994  ( .A(\GFM/N624 ), .B(\GFM/N627 ), .Z(\GFM/n498 ) );
XOR2_X2 \GFM/U3993  ( .A(\GFM/N621 ), .B(\GFM/N623 ), .Z(\GFM/n4990 ) );
XOR2_X2 \GFM/U3992  ( .A(\GFM/n501 ), .B(\GFM/n5000 ), .Z(z_out[21]) );
XOR2_X2 \GFM/U3991  ( .A(\GFM/n5030 ), .B(\GFM/n502 ), .Z(\GFM/n5000 ) );
XOR2_X2 \GFM/U3990  ( .A(\GFM/n505 ), .B(\GFM/n5040 ), .Z(\GFM/n501 ) );
XOR2_X2 \GFM/U3989  ( .A(\GFM/n5070 ), .B(\GFM/n5060 ), .Z(\GFM/n502 ) );
XOR2_X2 \GFM/U3988  ( .A(\GFM/n509 ), .B(\GFM/n508 ), .Z(\GFM/n5030 ) );
XOR2_X2 \GFM/U3987  ( .A(\GFM/n5110 ), .B(\GFM/n510 ), .Z(\GFM/n5040 ) );
XOR2_X2 \GFM/U3986  ( .A(\GFM/n513 ), .B(\GFM/n5120 ), .Z(\GFM/n505 ) );
XOR2_X2 \GFM/U3985  ( .A(z_in[21]), .B(\GFM/n5140 ), .Z(\GFM/n5060 ) );
XOR2_X2 \GFM/U3984  ( .A(\GFM/N678 ), .B(\GFM/N679 ), .Z(\GFM/n5070 ) );
XOR2_X2 \GFM/U3983  ( .A(\GFM/N675 ), .B(\GFM/N676 ), .Z(\GFM/n508 ) );
XOR2_X2 \GFM/U3982  ( .A(\GFM/N671 ), .B(\GFM/N672 ), .Z(\GFM/n509 ) );
XOR2_X2 \GFM/U3981  ( .A(\GFM/N667 ), .B(\GFM/N669 ), .Z(\GFM/n510 ) );
XOR2_X2 \GFM/U3980  ( .A(\GFM/N662 ), .B(\GFM/N666 ), .Z(\GFM/n5110 ) );
XOR2_X2 \GFM/U3979  ( .A(\GFM/N659 ), .B(\GFM/N661 ), .Z(\GFM/n5120 ) );
XOR2_X2 \GFM/U3978  ( .A(\GFM/N655 ), .B(\GFM/N658 ), .Z(\GFM/n513 ) );
XOR2_X2 \GFM/U3977  ( .A(\GFM/N652 ), .B(\GFM/N654 ), .Z(\GFM/n5140 ) );
XOR2_X2 \GFM/U3976  ( .A(\GFM/n5160 ), .B(\GFM/n515 ), .Z(z_out[22]) );
XOR2_X2 \GFM/U3975  ( .A(\GFM/n518 ), .B(\GFM/n5170 ), .Z(\GFM/n515 ) );
XOR2_X2 \GFM/U3974  ( .A(\GFM/n5200 ), .B(\GFM/n519 ), .Z(\GFM/n5160 ) );
XOR2_X2 \GFM/U3973  ( .A(\GFM/n522 ), .B(\GFM/n5210 ), .Z(\GFM/n5170 ) );
XOR2_X2 \GFM/U3972  ( .A(\GFM/n5240 ), .B(\GFM/n5230 ), .Z(\GFM/n518 ) );
XOR2_X2 \GFM/U3971  ( .A(\GFM/n526 ), .B(\GFM/n525 ), .Z(\GFM/n519 ) );
XOR2_X2 \GFM/U3970  ( .A(\GFM/n5280 ), .B(\GFM/n527 ), .Z(\GFM/n5200 ) );
XOR2_X2 \GFM/U3969  ( .A(z_in[22]), .B(\GFM/n529 ), .Z(\GFM/n5210 ) );
XOR2_X2 \GFM/U3968  ( .A(\GFM/N709 ), .B(\GFM/N710 ), .Z(\GFM/n522 ) );
XOR2_X2 \GFM/U3967  ( .A(\GFM/N706 ), .B(\GFM/N707 ), .Z(\GFM/n5230 ) );
XOR2_X2 \GFM/U3966  ( .A(\GFM/N702 ), .B(\GFM/N703 ), .Z(\GFM/n5240 ) );
XOR2_X2 \GFM/U3965  ( .A(\GFM/N698 ), .B(\GFM/N700 ), .Z(\GFM/n525 ) );
XOR2_X2 \GFM/U3964  ( .A(\GFM/N693 ), .B(\GFM/N697 ), .Z(\GFM/n526 ) );
XOR2_X2 \GFM/U3963  ( .A(\GFM/N690 ), .B(\GFM/N692 ), .Z(\GFM/n527 ) );
XOR2_X2 \GFM/U3962  ( .A(\GFM/N686 ), .B(\GFM/N689 ), .Z(\GFM/n5280 ) );
XOR2_X2 \GFM/U3961  ( .A(\GFM/N683 ), .B(\GFM/N685 ), .Z(\GFM/n529 ) );
XOR2_X2 \GFM/U3960  ( .A(\GFM/n5310 ), .B(\GFM/n5300 ), .Z(z_out[23]) );
XOR2_X2 \GFM/U3959  ( .A(\GFM/n533 ), .B(\GFM/n532 ), .Z(\GFM/n5300 ) );
XOR2_X2 \GFM/U3958  ( .A(\GFM/n5350 ), .B(\GFM/n5340 ), .Z(\GFM/n5310 ) );
XOR2_X2 \GFM/U3957  ( .A(\GFM/n5370 ), .B(\GFM/n536 ), .Z(\GFM/n532 ) );
XOR2_X2 \GFM/U3956  ( .A(\GFM/n539 ), .B(\GFM/n5380 ), .Z(\GFM/n533 ) );
XOR2_X2 \GFM/U3955  ( .A(\GFM/n541 ), .B(\GFM/n540 ), .Z(\GFM/n5340 ) );
XOR2_X2 \GFM/U3954  ( .A(\GFM/n5430 ), .B(\GFM/n5420 ), .Z(\GFM/n5350 ) );
XOR2_X2 \GFM/U3953  ( .A(z_in[23]), .B(\GFM/n544 ), .Z(\GFM/n536 ) );
XOR2_X2 \GFM/U3952  ( .A(\GFM/N740 ), .B(\GFM/N741 ), .Z(\GFM/n5370 ) );
XOR2_X2 \GFM/U3951  ( .A(\GFM/N737 ), .B(\GFM/N738 ), .Z(\GFM/n5380 ) );
XOR2_X2 \GFM/U3950  ( .A(\GFM/N733 ), .B(\GFM/N734 ), .Z(\GFM/n539 ) );
XOR2_X2 \GFM/U3949  ( .A(\GFM/N729 ), .B(\GFM/N731 ), .Z(\GFM/n540 ) );
XOR2_X2 \GFM/U3948  ( .A(\GFM/N724 ), .B(\GFM/N728 ), .Z(\GFM/n541 ) );
XOR2_X2 \GFM/U3947  ( .A(\GFM/N721 ), .B(\GFM/N723 ), .Z(\GFM/n5420 ) );
XOR2_X2 \GFM/U3946  ( .A(\GFM/N717 ), .B(\GFM/N720 ), .Z(\GFM/n5430 ) );
XOR2_X2 \GFM/U3945  ( .A(\GFM/N714 ), .B(\GFM/N716 ), .Z(\GFM/n544 ) );
XOR2_X2 \GFM/U3944  ( .A(\GFM/n546 ), .B(\GFM/n5450 ), .Z(z_out[24]) );
XOR2_X2 \GFM/U3943  ( .A(\GFM/n5480 ), .B(\GFM/n5470 ), .Z(\GFM/n5450 ) );
XOR2_X2 \GFM/U3942  ( .A(\GFM/n550 ), .B(\GFM/n549 ), .Z(\GFM/n546 ) );
XOR2_X2 \GFM/U3941  ( .A(\GFM/n5520 ), .B(\GFM/n5510 ), .Z(\GFM/n5470 ) );
XOR2_X2 \GFM/U3940  ( .A(\GFM/n5540 ), .B(\GFM/n553 ), .Z(\GFM/n5480 ) );
XOR2_X2 \GFM/U3939  ( .A(\GFM/n556 ), .B(\GFM/n5550 ), .Z(\GFM/n549 ) );
XOR2_X2 \GFM/U3938  ( .A(\GFM/n558 ), .B(\GFM/n557 ), .Z(\GFM/n550 ) );
XOR2_X2 \GFM/U3937  ( .A(z_in[24]), .B(\GFM/n5590 ), .Z(\GFM/n5510 ) );
XOR2_X2 \GFM/U3936  ( .A(\GFM/N771 ), .B(\GFM/N772 ), .Z(\GFM/n5520 ) );
XOR2_X2 \GFM/U3935  ( .A(\GFM/N768 ), .B(\GFM/N769 ), .Z(\GFM/n553 ) );
XOR2_X2 \GFM/U3934  ( .A(\GFM/N764 ), .B(\GFM/N765 ), .Z(\GFM/n5540 ) );
XOR2_X2 \GFM/U3933  ( .A(\GFM/N760 ), .B(\GFM/N762 ), .Z(\GFM/n5550 ) );
XOR2_X2 \GFM/U3932  ( .A(\GFM/N755 ), .B(\GFM/N759 ), .Z(\GFM/n556 ) );
XOR2_X2 \GFM/U3931  ( .A(\GFM/N752 ), .B(\GFM/N754 ), .Z(\GFM/n557 ) );
XOR2_X2 \GFM/U3930  ( .A(\GFM/N748 ), .B(\GFM/N751 ), .Z(\GFM/n558 ) );
XOR2_X2 \GFM/U3929  ( .A(\GFM/N745 ), .B(\GFM/N747 ), .Z(\GFM/n5590 ) );
XOR2_X2 \GFM/U3928  ( .A(\GFM/n5610 ), .B(\GFM/n560 ), .Z(z_out[25]) );
XOR2_X2 \GFM/U3927  ( .A(\GFM/n563 ), .B(\GFM/n5620 ), .Z(\GFM/n560 ) );
XOR2_X2 \GFM/U3926  ( .A(\GFM/n5650 ), .B(\GFM/n564 ), .Z(\GFM/n5610 ) );
XOR2_X2 \GFM/U3925  ( .A(\GFM/n567 ), .B(\GFM/n5660 ), .Z(\GFM/n5620 ) );
XOR2_X2 \GFM/U3924  ( .A(\GFM/n5690 ), .B(\GFM/n5680 ), .Z(\GFM/n563 ) );
XOR2_X2 \GFM/U3923  ( .A(\GFM/n571 ), .B(\GFM/n570 ), .Z(\GFM/n564 ) );
XOR2_X2 \GFM/U3922  ( .A(\GFM/n5730 ), .B(\GFM/n572 ), .Z(\GFM/n5650 ) );
XOR2_X2 \GFM/U3921  ( .A(z_in[25]), .B(\GFM/n5740 ), .Z(\GFM/n5660 ) );
XOR2_X2 \GFM/U3920  ( .A(\GFM/N802 ), .B(\GFM/N803 ), .Z(\GFM/n567 ) );
XOR2_X2 \GFM/U3919  ( .A(\GFM/N799 ), .B(\GFM/N800 ), .Z(\GFM/n5680 ) );
XOR2_X2 \GFM/U3918  ( .A(\GFM/N795 ), .B(\GFM/N796 ), .Z(\GFM/n5690 ) );
XOR2_X2 \GFM/U3917  ( .A(\GFM/N791 ), .B(\GFM/N793 ), .Z(\GFM/n570 ) );
XOR2_X2 \GFM/U3916  ( .A(\GFM/N786 ), .B(\GFM/N790 ), .Z(\GFM/n571 ) );
XOR2_X2 \GFM/U3915  ( .A(\GFM/N783 ), .B(\GFM/N785 ), .Z(\GFM/n572 ) );
XOR2_X2 \GFM/U3914  ( .A(\GFM/N779 ), .B(\GFM/N782 ), .Z(\GFM/n5730 ) );
XOR2_X2 \GFM/U3913  ( .A(\GFM/N776 ), .B(\GFM/N778 ), .Z(\GFM/n5740 ) );
XOR2_X2 \GFM/U3912  ( .A(\GFM/n5760 ), .B(\GFM/n575 ), .Z(z_out[26]) );
XOR2_X2 \GFM/U3911  ( .A(\GFM/n5780 ), .B(\GFM/n577 ), .Z(\GFM/n575 ) );
XOR2_X2 \GFM/U3910  ( .A(\GFM/n580 ), .B(\GFM/n5790 ), .Z(\GFM/n5760 ) );
XOR2_X2 \GFM/U3909  ( .A(\GFM/n5820 ), .B(\GFM/n581 ), .Z(\GFM/n577 ) );
XOR2_X2 \GFM/U3908  ( .A(\GFM/n584 ), .B(\GFM/n5830 ), .Z(\GFM/n5780 ) );
XOR2_X2 \GFM/U3907  ( .A(\GFM/n5860 ), .B(\GFM/n5850 ), .Z(\GFM/n5790 ) );
XOR2_X2 \GFM/U3906  ( .A(\GFM/n588 ), .B(\GFM/n587 ), .Z(\GFM/n580 ) );
XOR2_X2 \GFM/U3905  ( .A(z_in[26]), .B(\GFM/n589 ), .Z(\GFM/n581 ) );
XOR2_X2 \GFM/U3904  ( .A(\GFM/N833 ), .B(\GFM/N834 ), .Z(\GFM/n5820 ) );
XOR2_X2 \GFM/U3903  ( .A(\GFM/N830 ), .B(\GFM/N831 ), .Z(\GFM/n5830 ) );
XOR2_X2 \GFM/U3902  ( .A(\GFM/N826 ), .B(\GFM/N827 ), .Z(\GFM/n584 ) );
XOR2_X2 \GFM/U3901  ( .A(\GFM/N822 ), .B(\GFM/N824 ), .Z(\GFM/n5850 ) );
XOR2_X2 \GFM/U3900  ( .A(\GFM/N817 ), .B(\GFM/N821 ), .Z(\GFM/n5860 ) );
XOR2_X2 \GFM/U3899  ( .A(\GFM/N814 ), .B(\GFM/N816 ), .Z(\GFM/n587 ) );
XOR2_X2 \GFM/U3898  ( .A(\GFM/N810 ), .B(\GFM/N813 ), .Z(\GFM/n588 ) );
XOR2_X2 \GFM/U3897  ( .A(\GFM/N807 ), .B(\GFM/N809 ), .Z(\GFM/n589 ) );
XOR2_X2 \GFM/U3896  ( .A(\GFM/n591 ), .B(\GFM/n5900 ), .Z(z_out[27]) );
XOR2_X2 \GFM/U3895  ( .A(\GFM/n5930 ), .B(\GFM/n5920 ), .Z(\GFM/n5900 ) );
XOR2_X2 \GFM/U3894  ( .A(\GFM/n595 ), .B(\GFM/n594 ), .Z(\GFM/n591 ) );
XOR2_X2 \GFM/U3893  ( .A(\GFM/n5970 ), .B(\GFM/n5960 ), .Z(\GFM/n5920 ) );
XOR2_X2 \GFM/U3892  ( .A(\GFM/n5990 ), .B(\GFM/n598 ), .Z(\GFM/n5930 ) );
XOR2_X2 \GFM/U3891  ( .A(\GFM/n601 ), .B(\GFM/n6000 ), .Z(\GFM/n594 ) );
XOR2_X2 \GFM/U3890  ( .A(\GFM/n603 ), .B(\GFM/n602 ), .Z(\GFM/n595 ) );
XOR2_X2 \GFM/U3889  ( .A(z_in[27]), .B(\GFM/n6040 ), .Z(\GFM/n5960 ) );
XOR2_X2 \GFM/U3888  ( .A(\GFM/N864 ), .B(\GFM/N865 ), .Z(\GFM/n5970 ) );
XOR2_X2 \GFM/U3887  ( .A(\GFM/N861 ), .B(\GFM/N862 ), .Z(\GFM/n598 ) );
XOR2_X2 \GFM/U3886  ( .A(\GFM/N857 ), .B(\GFM/N858 ), .Z(\GFM/n5990 ) );
XOR2_X2 \GFM/U3885  ( .A(\GFM/N853 ), .B(\GFM/N855 ), .Z(\GFM/n6000 ) );
XOR2_X2 \GFM/U3884  ( .A(\GFM/N848 ), .B(\GFM/N852 ), .Z(\GFM/n601 ) );
XOR2_X2 \GFM/U3883  ( .A(\GFM/N845 ), .B(\GFM/N847 ), .Z(\GFM/n602 ) );
XOR2_X2 \GFM/U3882  ( .A(\GFM/N841 ), .B(\GFM/N844 ), .Z(\GFM/n603 ) );
XOR2_X2 \GFM/U3881  ( .A(\GFM/N838 ), .B(\GFM/N840 ), .Z(\GFM/n6040 ) );
XOR2_X2 \GFM/U3880  ( .A(\GFM/n606 ), .B(\GFM/n6050 ), .Z(z_out[28]) );
XOR2_X2 \GFM/U3879  ( .A(\GFM/n608 ), .B(\GFM/n6070 ), .Z(\GFM/n6050 ) );
XOR2_X2 \GFM/U3878  ( .A(\GFM/n6100 ), .B(\GFM/n6090 ), .Z(\GFM/n606 ) );
XOR2_X2 \GFM/U3877  ( .A(\GFM/n612 ), .B(\GFM/n611 ), .Z(\GFM/n6070 ) );
XOR2_X2 \GFM/U3876  ( .A(\GFM/n6140 ), .B(\GFM/n6130 ), .Z(\GFM/n608 ) );
XOR2_X2 \GFM/U3875  ( .A(\GFM/n6160 ), .B(\GFM/n615 ), .Z(\GFM/n6090 ) );
XOR2_X2 \GFM/U3874  ( .A(\GFM/n618 ), .B(\GFM/n6170 ), .Z(\GFM/n6100 ) );
XOR2_X2 \GFM/U3873  ( .A(z_in[28]), .B(\GFM/n619 ), .Z(\GFM/n611 ) );
XOR2_X2 \GFM/U3872  ( .A(\GFM/N895 ), .B(\GFM/N896 ), .Z(\GFM/n612 ) );
XOR2_X2 \GFM/U3871  ( .A(\GFM/N892 ), .B(\GFM/N893 ), .Z(\GFM/n6130 ) );
XOR2_X2 \GFM/U3870  ( .A(\GFM/N888 ), .B(\GFM/N889 ), .Z(\GFM/n6140 ) );
XOR2_X2 \GFM/U3869  ( .A(\GFM/N884 ), .B(\GFM/N886 ), .Z(\GFM/n615 ) );
XOR2_X2 \GFM/U3868  ( .A(\GFM/N879 ), .B(\GFM/N883 ), .Z(\GFM/n6160 ) );
XOR2_X2 \GFM/U3867  ( .A(\GFM/N876 ), .B(\GFM/N878 ), .Z(\GFM/n6170 ) );
XOR2_X2 \GFM/U3866  ( .A(\GFM/N872 ), .B(\GFM/N875 ), .Z(\GFM/n618 ) );
XOR2_X2 \GFM/U3865  ( .A(\GFM/N869 ), .B(\GFM/N871 ), .Z(\GFM/n619 ) );
XOR2_X2 \GFM/U3864  ( .A(\GFM/n6210 ), .B(\GFM/n620 ), .Z(z_out[29]) );
XOR2_X2 \GFM/U3863  ( .A(\GFM/n6230 ), .B(\GFM/n622 ), .Z(\GFM/n620 ) );
XOR2_X2 \GFM/U3862  ( .A(\GFM/n625 ), .B(\GFM/n6240 ), .Z(\GFM/n6210 ) );
XOR2_X2 \GFM/U3861  ( .A(\GFM/n6270 ), .B(\GFM/n626 ), .Z(\GFM/n622 ) );
XOR2_X2 \GFM/U3860  ( .A(\GFM/n629 ), .B(\GFM/n6280 ), .Z(\GFM/n6230 ) );
XOR2_X2 \GFM/U3859  ( .A(\GFM/n6310 ), .B(\GFM/n6300 ), .Z(\GFM/n6240 ) );
XOR2_X2 \GFM/U3858  ( .A(\GFM/n633 ), .B(\GFM/n632 ), .Z(\GFM/n625 ) );
XOR2_X2 \GFM/U3857  ( .A(z_in[29]), .B(\GFM/n634 ), .Z(\GFM/n626 ) );
XOR2_X2 \GFM/U3856  ( .A(\GFM/N926 ), .B(\GFM/N927 ), .Z(\GFM/n6270 ) );
XOR2_X2 \GFM/U3855  ( .A(\GFM/N923 ), .B(\GFM/N924 ), .Z(\GFM/n6280 ) );
XOR2_X2 \GFM/U3854  ( .A(\GFM/N919 ), .B(\GFM/N920 ), .Z(\GFM/n629 ) );
XOR2_X2 \GFM/U3853  ( .A(\GFM/N915 ), .B(\GFM/N917 ), .Z(\GFM/n6300 ) );
XOR2_X2 \GFM/U3852  ( .A(\GFM/N910 ), .B(\GFM/N914 ), .Z(\GFM/n6310 ) );
XOR2_X2 \GFM/U3851  ( .A(\GFM/N907 ), .B(\GFM/N909 ), .Z(\GFM/n632 ) );
XOR2_X2 \GFM/U3850  ( .A(\GFM/N903 ), .B(\GFM/N906 ), .Z(\GFM/n633 ) );
XOR2_X2 \GFM/U3849  ( .A(\GFM/N900 ), .B(\GFM/N902 ), .Z(\GFM/n634 ) );
XOR2_X2 \GFM/U3848  ( .A(\GFM/n6360 ), .B(\GFM/n6350 ), .Z(z_out[30]) );
XOR2_X2 \GFM/U3847  ( .A(\GFM/n6380 ), .B(\GFM/n637 ), .Z(\GFM/n6350 ) );
XOR2_X2 \GFM/U3846  ( .A(\GFM/n6400 ), .B(\GFM/n639 ), .Z(\GFM/n6360 ) );
XOR2_X2 \GFM/U3845  ( .A(\GFM/n642 ), .B(\GFM/n6410 ), .Z(\GFM/n637 ) );
XOR2_X2 \GFM/U3844  ( .A(\GFM/n6440 ), .B(\GFM/n643 ), .Z(\GFM/n6380 ) );
XOR2_X2 \GFM/U3843  ( .A(\GFM/n646 ), .B(\GFM/n6450 ), .Z(\GFM/n639 ) );
XOR2_X2 \GFM/U3842  ( .A(\GFM/n6480 ), .B(\GFM/n6470 ), .Z(\GFM/n6400 ) );
XOR2_X2 \GFM/U3841  ( .A(z_in[30]), .B(\GFM/n649 ), .Z(\GFM/n6410 ) );
XOR2_X2 \GFM/U3840  ( .A(\GFM/N957 ), .B(\GFM/N958 ), .Z(\GFM/n642 ) );
XOR2_X2 \GFM/U3839  ( .A(\GFM/N954 ), .B(\GFM/N955 ), .Z(\GFM/n643 ) );
XOR2_X2 \GFM/U3838  ( .A(\GFM/N950 ), .B(\GFM/N951 ), .Z(\GFM/n6440 ) );
XOR2_X2 \GFM/U3837  ( .A(\GFM/N946 ), .B(\GFM/N948 ), .Z(\GFM/n6450 ) );
XOR2_X2 \GFM/U3836  ( .A(\GFM/N941 ), .B(\GFM/N945 ), .Z(\GFM/n646 ) );
XOR2_X2 \GFM/U3835  ( .A(\GFM/N938 ), .B(\GFM/N940 ), .Z(\GFM/n6470 ) );
XOR2_X2 \GFM/U3834  ( .A(\GFM/N934 ), .B(\GFM/N937 ), .Z(\GFM/n6480 ) );
XOR2_X2 \GFM/U3833  ( .A(\GFM/N931 ), .B(\GFM/N933 ), .Z(\GFM/n649 ) );
XOR2_X2 \GFM/U3832  ( .A(\GFM/n651 ), .B(\GFM/n650 ), .Z(z_out[31]) );
XOR2_X2 \GFM/U3831  ( .A(\GFM/n653 ), .B(\GFM/n6520 ), .Z(\GFM/n650 ) );
XOR2_X2 \GFM/U3830  ( .A(\GFM/n6550 ), .B(\GFM/n6540 ), .Z(\GFM/n651 ) );
XOR2_X2 \GFM/U3829  ( .A(\GFM/n657 ), .B(\GFM/n656 ), .Z(\GFM/n6520 ) );
XOR2_X2 \GFM/U3828  ( .A(\GFM/n6590 ), .B(\GFM/n6580 ), .Z(\GFM/n653 ) );
XOR2_X2 \GFM/U3827  ( .A(\GFM/n6610 ), .B(\GFM/n660 ), .Z(\GFM/n6540 ) );
XOR2_X2 \GFM/U3826  ( .A(\GFM/n663 ), .B(\GFM/n6620 ), .Z(\GFM/n6550 ) );
XOR2_X2 \GFM/U3825  ( .A(z_in[31]), .B(\GFM/n664 ), .Z(\GFM/n656 ) );
XOR2_X2 \GFM/U3824  ( .A(\GFM/N988 ), .B(\GFM/N989 ), .Z(\GFM/n657 ) );
XOR2_X2 \GFM/U3823  ( .A(\GFM/N985 ), .B(\GFM/N986 ), .Z(\GFM/n6580 ) );
XOR2_X2 \GFM/U3822  ( .A(\GFM/N981 ), .B(\GFM/N982 ), .Z(\GFM/n6590 ) );
XOR2_X2 \GFM/U3821  ( .A(\GFM/N977 ), .B(\GFM/N979 ), .Z(\GFM/n660 ) );
XOR2_X2 \GFM/U3820  ( .A(\GFM/N972 ), .B(\GFM/N976 ), .Z(\GFM/n6610 ) );
XOR2_X2 \GFM/U3819  ( .A(\GFM/N969 ), .B(\GFM/N971 ), .Z(\GFM/n6620 ) );
XOR2_X2 \GFM/U3818  ( .A(\GFM/N965 ), .B(\GFM/N968 ), .Z(\GFM/n663 ) );
XOR2_X2 \GFM/U3817  ( .A(\GFM/N962 ), .B(\GFM/N964 ), .Z(\GFM/n664 ) );
XOR2_X2 \GFM/U3816  ( .A(\GFM/n6660 ), .B(\GFM/n665 ), .Z(z_out[32]) );
XOR2_X2 \GFM/U3815  ( .A(\GFM/n668 ), .B(\GFM/n6670 ), .Z(\GFM/n665 ) );
XOR2_X2 \GFM/U3814  ( .A(\GFM/n670 ), .B(\GFM/n6690 ), .Z(\GFM/n6660 ) );
XOR2_X2 \GFM/U3813  ( .A(\GFM/n6720 ), .B(\GFM/n6710 ), .Z(\GFM/n6670 ) );
XOR2_X2 \GFM/U3812  ( .A(\GFM/n674 ), .B(\GFM/n673 ), .Z(\GFM/n668 ) );
XOR2_X2 \GFM/U3811  ( .A(\GFM/n6760 ), .B(\GFM/n6750 ), .Z(\GFM/n6690 ) );
XOR2_X2 \GFM/U3810  ( .A(\GFM/n6780 ), .B(\GFM/n677 ), .Z(\GFM/n670 ) );
XOR2_X2 \GFM/U3809  ( .A(z_in[32]), .B(\GFM/n6790 ), .Z(\GFM/n6710 ) );
XOR2_X2 \GFM/U3808  ( .A(\GFM/N1019 ), .B(\GFM/N1020 ), .Z(\GFM/n6720 ) );
XOR2_X2 \GFM/U3807  ( .A(\GFM/N1016 ), .B(\GFM/N1017 ), .Z(\GFM/n673 ) );
XOR2_X2 \GFM/U3806  ( .A(\GFM/N1012 ), .B(\GFM/N1013 ), .Z(\GFM/n674 ) );
XOR2_X2 \GFM/U3805  ( .A(\GFM/N1008 ), .B(\GFM/N1010 ), .Z(\GFM/n6750 ) );
XOR2_X2 \GFM/U3804  ( .A(\GFM/N1003 ), .B(\GFM/N1007 ), .Z(\GFM/n6760 ) );
XOR2_X2 \GFM/U3803  ( .A(\GFM/N1000 ), .B(\GFM/N1002 ), .Z(\GFM/n677 ) );
XOR2_X2 \GFM/U3802  ( .A(\GFM/N996 ), .B(\GFM/N999 ), .Z(\GFM/n6780 ) );
XOR2_X2 \GFM/U3801  ( .A(\GFM/N993 ), .B(\GFM/N995 ), .Z(\GFM/n6790 ) );
XOR2_X2 \GFM/U3800  ( .A(\GFM/n681 ), .B(\GFM/n680 ), .Z(z_out[33]) );
XOR2_X2 \GFM/U3799  ( .A(\GFM/n6830 ), .B(\GFM/n682 ), .Z(\GFM/n680 ) );
XOR2_X2 \GFM/U3798  ( .A(\GFM/n6850 ), .B(\GFM/n684 ), .Z(\GFM/n681 ) );
XOR2_X2 \GFM/U3797  ( .A(\GFM/n687 ), .B(\GFM/n6860 ), .Z(\GFM/n682 ) );
XOR2_X2 \GFM/U3796  ( .A(\GFM/n6890 ), .B(\GFM/n688 ), .Z(\GFM/n6830 ) );
XOR2_X2 \GFM/U3795  ( .A(\GFM/n691 ), .B(\GFM/n6900 ), .Z(\GFM/n684 ) );
XOR2_X2 \GFM/U3794  ( .A(\GFM/n6930 ), .B(\GFM/n6920 ), .Z(\GFM/n6850 ) );
XOR2_X2 \GFM/U3793  ( .A(z_in[33]), .B(\GFM/n694 ), .Z(\GFM/n6860 ) );
XOR2_X2 \GFM/U3792  ( .A(\GFM/N1050 ), .B(\GFM/N1051 ), .Z(\GFM/n687 ) );
XOR2_X2 \GFM/U3791  ( .A(\GFM/N1047 ), .B(\GFM/N1048 ), .Z(\GFM/n688 ) );
XOR2_X2 \GFM/U3790  ( .A(\GFM/N1043 ), .B(\GFM/N1044 ), .Z(\GFM/n6890 ) );
XOR2_X2 \GFM/U3789  ( .A(\GFM/N1039 ), .B(\GFM/N1041 ), .Z(\GFM/n6900 ) );
XOR2_X2 \GFM/U3788  ( .A(\GFM/N1034 ), .B(\GFM/N1038 ), .Z(\GFM/n691 ) );
XOR2_X2 \GFM/U3787  ( .A(\GFM/N1031 ), .B(\GFM/N1033 ), .Z(\GFM/n6920 ) );
XOR2_X2 \GFM/U3786  ( .A(\GFM/N1027 ), .B(\GFM/N1030 ), .Z(\GFM/n6930 ) );
XOR2_X2 \GFM/U3785  ( .A(\GFM/N1024 ), .B(\GFM/N1026 ), .Z(\GFM/n694 ) );
XOR2_X2 \GFM/U3784  ( .A(\GFM/n696 ), .B(\GFM/n695 ), .Z(z_out[34]) );
XOR2_X2 \GFM/U3783  ( .A(\GFM/n6980 ), .B(\GFM/n6970 ), .Z(\GFM/n695 ) );
XOR2_X2 \GFM/U3782  ( .A(\GFM/n7000 ), .B(\GFM/n699 ), .Z(\GFM/n696 ) );
XOR2_X2 \GFM/U3781  ( .A(\GFM/n7020 ), .B(\GFM/n701 ), .Z(\GFM/n6970 ) );
XOR2_X2 \GFM/U3780  ( .A(\GFM/n704 ), .B(\GFM/n7030 ), .Z(\GFM/n6980 ) );
XOR2_X2 \GFM/U3779  ( .A(\GFM/n7060 ), .B(\GFM/n705 ), .Z(\GFM/n699 ) );
XOR2_X2 \GFM/U3778  ( .A(\GFM/n708 ), .B(\GFM/n7070 ), .Z(\GFM/n7000 ) );
XOR2_X2 \GFM/U3777  ( .A(z_in[34]), .B(\GFM/n7090 ), .Z(\GFM/n701 ) );
XOR2_X2 \GFM/U3776  ( .A(\GFM/N1081 ), .B(\GFM/N1082 ), .Z(\GFM/n7020 ) );
XOR2_X2 \GFM/U3775  ( .A(\GFM/N1078 ), .B(\GFM/N1079 ), .Z(\GFM/n7030 ) );
XOR2_X2 \GFM/U3774  ( .A(\GFM/N1074 ), .B(\GFM/N1075 ), .Z(\GFM/n704 ) );
XOR2_X2 \GFM/U3773  ( .A(\GFM/N1070 ), .B(\GFM/N1072 ), .Z(\GFM/n705 ) );
XOR2_X2 \GFM/U3772  ( .A(\GFM/N1065 ), .B(\GFM/N1069 ), .Z(\GFM/n7060 ) );
XOR2_X2 \GFM/U3771  ( .A(\GFM/N1062 ), .B(\GFM/N1064 ), .Z(\GFM/n7070 ) );
XOR2_X2 \GFM/U3770  ( .A(\GFM/N1058 ), .B(\GFM/N1061 ), .Z(\GFM/n708 ) );
XOR2_X2 \GFM/U3769  ( .A(\GFM/N1055 ), .B(\GFM/N1057 ), .Z(\GFM/n7090 ) );
XOR2_X2 \GFM/U3768  ( .A(\GFM/n711 ), .B(\GFM/n7100 ), .Z(z_out[35]) );
XOR2_X2 \GFM/U3767  ( .A(\GFM/n713 ), .B(\GFM/n712 ), .Z(\GFM/n7100 ) );
XOR2_X2 \GFM/U3766  ( .A(\GFM/n715 ), .B(\GFM/n7140 ), .Z(\GFM/n711 ) );
XOR2_X2 \GFM/U3765  ( .A(\GFM/n7170 ), .B(\GFM/n7160 ), .Z(\GFM/n712 ) );
XOR2_X2 \GFM/U3764  ( .A(\GFM/n719 ), .B(\GFM/n718 ), .Z(\GFM/n713 ) );
XOR2_X2 \GFM/U3763  ( .A(\GFM/n7210 ), .B(\GFM/n7200 ), .Z(\GFM/n7140 ) );
XOR2_X2 \GFM/U3762  ( .A(\GFM/n7230 ), .B(\GFM/n722 ), .Z(\GFM/n715 ) );
XOR2_X2 \GFM/U3761  ( .A(z_in[35]), .B(\GFM/n7240 ), .Z(\GFM/n7160 ) );
XOR2_X2 \GFM/U3760  ( .A(\GFM/N1112 ), .B(\GFM/N1113 ), .Z(\GFM/n7170 ) );
XOR2_X2 \GFM/U3759  ( .A(\GFM/N1109 ), .B(\GFM/N1110 ), .Z(\GFM/n718 ) );
XOR2_X2 \GFM/U3758  ( .A(\GFM/N1105 ), .B(\GFM/N1106 ), .Z(\GFM/n719 ) );
XOR2_X2 \GFM/U3757  ( .A(\GFM/N1101 ), .B(\GFM/N1103 ), .Z(\GFM/n7200 ) );
XOR2_X2 \GFM/U3756  ( .A(\GFM/N1096 ), .B(\GFM/N1100 ), .Z(\GFM/n7210 ) );
XOR2_X2 \GFM/U3755  ( .A(\GFM/N1093 ), .B(\GFM/N1095 ), .Z(\GFM/n722 ) );
XOR2_X2 \GFM/U3754  ( .A(\GFM/N1089 ), .B(\GFM/N1092 ), .Z(\GFM/n7230 ) );
XOR2_X2 \GFM/U3753  ( .A(\GFM/N1086 ), .B(\GFM/N1088 ), .Z(\GFM/n7240 ) );
XOR2_X2 \GFM/U3752  ( .A(\GFM/n726 ), .B(\GFM/n725 ), .Z(z_out[36]) );
XOR2_X2 \GFM/U3751  ( .A(\GFM/n7280 ), .B(\GFM/n727 ), .Z(\GFM/n725 ) );
XOR2_X2 \GFM/U3750  ( .A(\GFM/n730 ), .B(\GFM/n7290 ), .Z(\GFM/n726 ) );
XOR2_X2 \GFM/U3749  ( .A(\GFM/n732 ), .B(\GFM/n7310 ), .Z(\GFM/n727 ) );
XOR2_X2 \GFM/U3748  ( .A(\GFM/n7340 ), .B(\GFM/n7330 ), .Z(\GFM/n7280 ) );
XOR2_X2 \GFM/U3747  ( .A(\GFM/n736 ), .B(\GFM/n735 ), .Z(\GFM/n7290 ) );
XOR2_X2 \GFM/U3746  ( .A(\GFM/n7380 ), .B(\GFM/n7370 ), .Z(\GFM/n730 ) );
XOR2_X2 \GFM/U3745  ( .A(z_in[36]), .B(\GFM/n739 ), .Z(\GFM/n7310 ) );
XOR2_X2 \GFM/U3744  ( .A(\GFM/N1143 ), .B(\GFM/N1144 ), .Z(\GFM/n732 ) );
XOR2_X2 \GFM/U3743  ( .A(\GFM/N1140 ), .B(\GFM/N1141 ), .Z(\GFM/n7330 ) );
XOR2_X2 \GFM/U3742  ( .A(\GFM/N1136 ), .B(\GFM/N1137 ), .Z(\GFM/n7340 ) );
XOR2_X2 \GFM/U3741  ( .A(\GFM/N1132 ), .B(\GFM/N1134 ), .Z(\GFM/n735 ) );
XOR2_X2 \GFM/U3740  ( .A(\GFM/N1127 ), .B(\GFM/N1131 ), .Z(\GFM/n736 ) );
XOR2_X2 \GFM/U3739  ( .A(\GFM/N1124 ), .B(\GFM/N1126 ), .Z(\GFM/n7370 ) );
XOR2_X2 \GFM/U3738  ( .A(\GFM/N1120 ), .B(\GFM/N1123 ), .Z(\GFM/n7380 ) );
XOR2_X2 \GFM/U3737  ( .A(\GFM/N1117 ), .B(\GFM/N1119 ), .Z(\GFM/n739 ) );
XOR2_X2 \GFM/U3736  ( .A(\GFM/n7410 ), .B(\GFM/n7400 ), .Z(z_out[37]) );
XOR2_X2 \GFM/U3735  ( .A(\GFM/n743 ), .B(\GFM/n742 ), .Z(\GFM/n7400 ) );
XOR2_X2 \GFM/U3734  ( .A(\GFM/n7450 ), .B(\GFM/n744 ), .Z(\GFM/n7410 ) );
XOR2_X2 \GFM/U3733  ( .A(\GFM/n7470 ), .B(\GFM/n746 ), .Z(\GFM/n742 ) );
XOR2_X2 \GFM/U3732  ( .A(\GFM/n749 ), .B(\GFM/n7480 ), .Z(\GFM/n743 ) );
XOR2_X2 \GFM/U3731  ( .A(\GFM/n7510 ), .B(\GFM/n750 ), .Z(\GFM/n744 ) );
XOR2_X2 \GFM/U3730  ( .A(\GFM/n753 ), .B(\GFM/n7520 ), .Z(\GFM/n7450 ) );
XOR2_X2 \GFM/U3729  ( .A(z_in[37]), .B(\GFM/n7540 ), .Z(\GFM/n746 ) );
XOR2_X2 \GFM/U3728  ( .A(\GFM/N1174 ), .B(\GFM/N1175 ), .Z(\GFM/n7470 ) );
XOR2_X2 \GFM/U3727  ( .A(\GFM/N1171 ), .B(\GFM/N1172 ), .Z(\GFM/n7480 ) );
XOR2_X2 \GFM/U3726  ( .A(\GFM/N1167 ), .B(\GFM/N1168 ), .Z(\GFM/n749 ) );
XOR2_X2 \GFM/U3725  ( .A(\GFM/N1163 ), .B(\GFM/N1165 ), .Z(\GFM/n750 ) );
XOR2_X2 \GFM/U3724  ( .A(\GFM/N1158 ), .B(\GFM/N1162 ), .Z(\GFM/n7510 ) );
XOR2_X2 \GFM/U3723  ( .A(\GFM/N1155 ), .B(\GFM/N1157 ), .Z(\GFM/n7520 ) );
XOR2_X2 \GFM/U3722  ( .A(\GFM/N1151 ), .B(\GFM/N1154 ), .Z(\GFM/n753 ) );
XOR2_X2 \GFM/U3721  ( .A(\GFM/N1148 ), .B(\GFM/N1150 ), .Z(\GFM/n7540 ) );
XOR2_X2 \GFM/U3720  ( .A(\GFM/n756 ), .B(\GFM/n7550 ), .Z(z_out[38]) );
XOR2_X2 \GFM/U3719  ( .A(\GFM/n758 ), .B(\GFM/n757 ), .Z(\GFM/n7550 ) );
XOR2_X2 \GFM/U3718  ( .A(\GFM/n7600 ), .B(\GFM/n7590 ), .Z(\GFM/n756 ) );
XOR2_X2 \GFM/U3717  ( .A(\GFM/n7620 ), .B(\GFM/n761 ), .Z(\GFM/n757 ) );
XOR2_X2 \GFM/U3716  ( .A(\GFM/n7640 ), .B(\GFM/n763 ), .Z(\GFM/n758 ) );
XOR2_X2 \GFM/U3715  ( .A(\GFM/n766 ), .B(\GFM/n7650 ), .Z(\GFM/n7590 ) );
XOR2_X2 \GFM/U3714  ( .A(\GFM/n7680 ), .B(\GFM/n767 ), .Z(\GFM/n7600 ) );
XOR2_X2 \GFM/U3713  ( .A(z_in[38]), .B(\GFM/n7690 ), .Z(\GFM/n761 ) );
XOR2_X2 \GFM/U3712  ( .A(\GFM/N1205 ), .B(\GFM/N1206 ), .Z(\GFM/n7620 ) );
XOR2_X2 \GFM/U3711  ( .A(\GFM/N1202 ), .B(\GFM/N1203 ), .Z(\GFM/n763 ) );
XOR2_X2 \GFM/U3710  ( .A(\GFM/N1198 ), .B(\GFM/N1199 ), .Z(\GFM/n7640 ) );
XOR2_X2 \GFM/U3709  ( .A(\GFM/N1194 ), .B(\GFM/N1196 ), .Z(\GFM/n7650 ) );
XOR2_X2 \GFM/U3708  ( .A(\GFM/N1189 ), .B(\GFM/N1193 ), .Z(\GFM/n766 ) );
XOR2_X2 \GFM/U3707  ( .A(\GFM/N1186 ), .B(\GFM/N1188 ), .Z(\GFM/n767 ) );
XOR2_X2 \GFM/U3706  ( .A(\GFM/N1182 ), .B(\GFM/N1185 ), .Z(\GFM/n7680 ) );
XOR2_X2 \GFM/U3705  ( .A(\GFM/N1179 ), .B(\GFM/N1181 ), .Z(\GFM/n7690 ) );
XOR2_X2 \GFM/U3704  ( .A(\GFM/n7710 ), .B(\GFM/n770 ), .Z(z_out[39]) );
XOR2_X2 \GFM/U3703  ( .A(\GFM/n773 ), .B(\GFM/n7720 ), .Z(\GFM/n770 ) );
XOR2_X2 \GFM/U3702  ( .A(\GFM/n775 ), .B(\GFM/n774 ), .Z(\GFM/n7710 ) );
XOR2_X2 \GFM/U3701  ( .A(\GFM/n777 ), .B(\GFM/n7760 ), .Z(\GFM/n7720 ) );
XOR2_X2 \GFM/U3700  ( .A(\GFM/n7790 ), .B(\GFM/n7780 ), .Z(\GFM/n773 ) );
XOR2_X2 \GFM/U3699  ( .A(\GFM/n781 ), .B(\GFM/n780 ), .Z(\GFM/n774 ) );
XOR2_X2 \GFM/U3698  ( .A(\GFM/n7830 ), .B(\GFM/n7820 ), .Z(\GFM/n775 ) );
XOR2_X2 \GFM/U3697  ( .A(z_in[39]), .B(\GFM/n784 ), .Z(\GFM/n7760 ) );
XOR2_X2 \GFM/U3696  ( .A(\GFM/N1236 ), .B(\GFM/N1237 ), .Z(\GFM/n777 ) );
XOR2_X2 \GFM/U3695  ( .A(\GFM/N1233 ), .B(\GFM/N1234 ), .Z(\GFM/n7780 ) );
XOR2_X2 \GFM/U3694  ( .A(\GFM/N1229 ), .B(\GFM/N1230 ), .Z(\GFM/n7790 ) );
XOR2_X2 \GFM/U3693  ( .A(\GFM/N1225 ), .B(\GFM/N1227 ), .Z(\GFM/n780 ) );
XOR2_X2 \GFM/U3692  ( .A(\GFM/N1220 ), .B(\GFM/N1224 ), .Z(\GFM/n781 ) );
XOR2_X2 \GFM/U3691  ( .A(\GFM/N1217 ), .B(\GFM/N1219 ), .Z(\GFM/n7820 ) );
XOR2_X2 \GFM/U3690  ( .A(\GFM/N1213 ), .B(\GFM/N1216 ), .Z(\GFM/n7830 ) );
XOR2_X2 \GFM/U3689  ( .A(\GFM/N1210 ), .B(\GFM/N1212 ), .Z(\GFM/n784 ) );
XOR2_X2 \GFM/U3688  ( .A(\GFM/n7860 ), .B(\GFM/n7850 ), .Z(z_out[40]) );
XOR2_X2 \GFM/U3687  ( .A(\GFM/n788 ), .B(\GFM/n787 ), .Z(\GFM/n7850 ) );
XOR2_X2 \GFM/U3686  ( .A(\GFM/n7900 ), .B(\GFM/n789 ), .Z(\GFM/n7860 ) );
XOR2_X2 \GFM/U3685  ( .A(\GFM/n792 ), .B(\GFM/n7910 ), .Z(\GFM/n787 ) );
XOR2_X2 \GFM/U3684  ( .A(\GFM/n794 ), .B(\GFM/n7930 ), .Z(\GFM/n788 ) );
XOR2_X2 \GFM/U3683  ( .A(\GFM/n7960 ), .B(\GFM/n7950 ), .Z(\GFM/n789 ) );
XOR2_X2 \GFM/U3682  ( .A(\GFM/n798 ), .B(\GFM/n797 ), .Z(\GFM/n7900 ) );
XOR2_X2 \GFM/U3681  ( .A(z_in[40]), .B(\GFM/n7990 ), .Z(\GFM/n7910 ) );
XOR2_X2 \GFM/U3680  ( .A(\GFM/N1267 ), .B(\GFM/N1268 ), .Z(\GFM/n792 ) );
XOR2_X2 \GFM/U3679  ( .A(\GFM/N1264 ), .B(\GFM/N1265 ), .Z(\GFM/n7930 ) );
XOR2_X2 \GFM/U3678  ( .A(\GFM/N1260 ), .B(\GFM/N1261 ), .Z(\GFM/n794 ) );
XOR2_X2 \GFM/U3677  ( .A(\GFM/N1256 ), .B(\GFM/N1258 ), .Z(\GFM/n7950 ) );
XOR2_X2 \GFM/U3676  ( .A(\GFM/N1251 ), .B(\GFM/N1255 ), .Z(\GFM/n7960 ) );
XOR2_X2 \GFM/U3675  ( .A(\GFM/N1248 ), .B(\GFM/N1250 ), .Z(\GFM/n797 ) );
XOR2_X2 \GFM/U3674  ( .A(\GFM/N1244 ), .B(\GFM/N1247 ), .Z(\GFM/n798 ) );
XOR2_X2 \GFM/U3673  ( .A(\GFM/N1241 ), .B(\GFM/N1243 ), .Z(\GFM/n7990 ) );
XOR2_X2 \GFM/U3672  ( .A(\GFM/n801 ), .B(\GFM/n8000 ), .Z(z_out[41]) );
XOR2_X2 \GFM/U3671  ( .A(\GFM/n8030 ), .B(\GFM/n8020 ), .Z(\GFM/n8000 ) );
XOR2_X2 \GFM/U3670  ( .A(\GFM/n805 ), .B(\GFM/n804 ), .Z(\GFM/n801 ) );
XOR2_X2 \GFM/U3669  ( .A(\GFM/n8070 ), .B(\GFM/n806 ), .Z(\GFM/n8020 ) );
XOR2_X2 \GFM/U3668  ( .A(\GFM/n8090 ), .B(\GFM/n808 ), .Z(\GFM/n8030 ) );
XOR2_X2 \GFM/U3667  ( .A(\GFM/n811 ), .B(\GFM/n8100 ), .Z(\GFM/n804 ) );
XOR2_X2 \GFM/U3666  ( .A(\GFM/n8130 ), .B(\GFM/n812 ), .Z(\GFM/n805 ) );
XOR2_X2 \GFM/U3665  ( .A(z_in[41]), .B(\GFM/n8140 ), .Z(\GFM/n806 ) );
XOR2_X2 \GFM/U3664  ( .A(\GFM/N1298 ), .B(\GFM/N1299 ), .Z(\GFM/n8070 ) );
XOR2_X2 \GFM/U3663  ( .A(\GFM/N1295 ), .B(\GFM/N1296 ), .Z(\GFM/n808 ) );
XOR2_X2 \GFM/U3662  ( .A(\GFM/N1291 ), .B(\GFM/N1292 ), .Z(\GFM/n8090 ) );
XOR2_X2 \GFM/U3661  ( .A(\GFM/N1287 ), .B(\GFM/N1289 ), .Z(\GFM/n8100 ) );
XOR2_X2 \GFM/U3660  ( .A(\GFM/N1282 ), .B(\GFM/N1286 ), .Z(\GFM/n811 ) );
XOR2_X2 \GFM/U3659  ( .A(\GFM/N1279 ), .B(\GFM/N1281 ), .Z(\GFM/n812 ) );
XOR2_X2 \GFM/U3658  ( .A(\GFM/N1275 ), .B(\GFM/N1278 ), .Z(\GFM/n8130 ) );
XOR2_X2 \GFM/U3657  ( .A(\GFM/N1272 ), .B(\GFM/N1274 ), .Z(\GFM/n8140 ) );
XOR2_X2 \GFM/U3656  ( .A(\GFM/n8160 ), .B(\GFM/n815 ), .Z(z_out[42]) );
XOR2_X2 \GFM/U3655  ( .A(\GFM/n818 ), .B(\GFM/n8170 ), .Z(\GFM/n815 ) );
XOR2_X2 \GFM/U3654  ( .A(\GFM/n820 ), .B(\GFM/n819 ), .Z(\GFM/n8160 ) );
XOR2_X2 \GFM/U3653  ( .A(\GFM/n8220 ), .B(\GFM/n8210 ), .Z(\GFM/n8170 ) );
XOR2_X2 \GFM/U3652  ( .A(\GFM/n8240 ), .B(\GFM/n823 ), .Z(\GFM/n818 ) );
XOR2_X2 \GFM/U3651  ( .A(\GFM/n8260 ), .B(\GFM/n825 ), .Z(\GFM/n819 ) );
XOR2_X2 \GFM/U3650  ( .A(\GFM/n828 ), .B(\GFM/n8270 ), .Z(\GFM/n820 ) );
XOR2_X2 \GFM/U3649  ( .A(z_in[42]), .B(\GFM/n829 ), .Z(\GFM/n8210 ) );
XOR2_X2 \GFM/U3648  ( .A(\GFM/N1329 ), .B(\GFM/N1330 ), .Z(\GFM/n8220 ) );
XOR2_X2 \GFM/U3647  ( .A(\GFM/N1326 ), .B(\GFM/N1327 ), .Z(\GFM/n823 ) );
XOR2_X2 \GFM/U3646  ( .A(\GFM/N1322 ), .B(\GFM/N1323 ), .Z(\GFM/n8240 ) );
XOR2_X2 \GFM/U3645  ( .A(\GFM/N1318 ), .B(\GFM/N1320 ), .Z(\GFM/n825 ) );
XOR2_X2 \GFM/U3644  ( .A(\GFM/N1313 ), .B(\GFM/N1317 ), .Z(\GFM/n8260 ) );
XOR2_X2 \GFM/U3643  ( .A(\GFM/N1310 ), .B(\GFM/N1312 ), .Z(\GFM/n8270 ) );
XOR2_X2 \GFM/U3642  ( .A(\GFM/N1306 ), .B(\GFM/N1309 ), .Z(\GFM/n828 ) );
XOR2_X2 \GFM/U3641  ( .A(\GFM/N1303 ), .B(\GFM/N1305 ), .Z(\GFM/n829 ) );
XOR2_X2 \GFM/U3640  ( .A(\GFM/n8310 ), .B(\GFM/n8300 ), .Z(z_out[43]) );
XOR2_X2 \GFM/U3639  ( .A(\GFM/n8330 ), .B(\GFM/n832 ), .Z(\GFM/n8300 ) );
XOR2_X2 \GFM/U3638  ( .A(\GFM/n835 ), .B(\GFM/n8340 ), .Z(\GFM/n8310 ) );
XOR2_X2 \GFM/U3637  ( .A(\GFM/n837 ), .B(\GFM/n836 ), .Z(\GFM/n832 ) );
XOR2_X2 \GFM/U3636  ( .A(\GFM/n839 ), .B(\GFM/n8380 ), .Z(\GFM/n8330 ) );
XOR2_X2 \GFM/U3635  ( .A(\GFM/n8410 ), .B(\GFM/n8400 ), .Z(\GFM/n8340 ) );
XOR2_X2 \GFM/U3634  ( .A(\GFM/n843 ), .B(\GFM/n842 ), .Z(\GFM/n835 ) );
XOR2_X2 \GFM/U3633  ( .A(z_in[43]), .B(\GFM/n8440 ), .Z(\GFM/n836 ) );
XOR2_X2 \GFM/U3632  ( .A(\GFM/N1360 ), .B(\GFM/N1361 ), .Z(\GFM/n837 ) );
XOR2_X2 \GFM/U3631  ( .A(\GFM/N1357 ), .B(\GFM/N1358 ), .Z(\GFM/n8380 ) );
XOR2_X2 \GFM/U3630  ( .A(\GFM/N1353 ), .B(\GFM/N1354 ), .Z(\GFM/n839 ) );
XOR2_X2 \GFM/U3629  ( .A(\GFM/N1349 ), .B(\GFM/N1351 ), .Z(\GFM/n8400 ) );
XOR2_X2 \GFM/U3628  ( .A(\GFM/N1344 ), .B(\GFM/N1348 ), .Z(\GFM/n8410 ) );
XOR2_X2 \GFM/U3627  ( .A(\GFM/N1341 ), .B(\GFM/N1343 ), .Z(\GFM/n842 ) );
XOR2_X2 \GFM/U3626  ( .A(\GFM/N1337 ), .B(\GFM/N1340 ), .Z(\GFM/n843 ) );
XOR2_X2 \GFM/U3625  ( .A(\GFM/N1334 ), .B(\GFM/N1336 ), .Z(\GFM/n8440 ) );
XOR2_X2 \GFM/U3624  ( .A(\GFM/n846 ), .B(\GFM/n8450 ), .Z(z_out[44]) );
XOR2_X2 \GFM/U3623  ( .A(\GFM/n8480 ), .B(\GFM/n8470 ), .Z(\GFM/n8450 ) );
XOR2_X2 \GFM/U3622  ( .A(\GFM/n850 ), .B(\GFM/n849 ), .Z(\GFM/n846 ) );
XOR2_X2 \GFM/U3621  ( .A(\GFM/n8520 ), .B(\GFM/n851 ), .Z(\GFM/n8470 ) );
XOR2_X2 \GFM/U3620  ( .A(\GFM/n854 ), .B(\GFM/n8530 ), .Z(\GFM/n8480 ) );
XOR2_X2 \GFM/U3619  ( .A(\GFM/n856 ), .B(\GFM/n8550 ), .Z(\GFM/n849 ) );
XOR2_X2 \GFM/U3618  ( .A(\GFM/n8580 ), .B(\GFM/n8570 ), .Z(\GFM/n850 ) );
XOR2_X2 \GFM/U3617  ( .A(z_in[44]), .B(\GFM/n859 ), .Z(\GFM/n851 ) );
XOR2_X2 \GFM/U3616  ( .A(\GFM/N1391 ), .B(\GFM/N1392 ), .Z(\GFM/n8520 ) );
XOR2_X2 \GFM/U3615  ( .A(\GFM/N1388 ), .B(\GFM/N1389 ), .Z(\GFM/n8530 ) );
XOR2_X2 \GFM/U3614  ( .A(\GFM/N1384 ), .B(\GFM/N1385 ), .Z(\GFM/n854 ) );
XOR2_X2 \GFM/U3613  ( .A(\GFM/N1380 ), .B(\GFM/N1382 ), .Z(\GFM/n8550 ) );
XOR2_X2 \GFM/U3612  ( .A(\GFM/N1375 ), .B(\GFM/N1379 ), .Z(\GFM/n856 ) );
XOR2_X2 \GFM/U3611  ( .A(\GFM/N1372 ), .B(\GFM/N1374 ), .Z(\GFM/n8570 ) );
XOR2_X2 \GFM/U3610  ( .A(\GFM/N1368 ), .B(\GFM/N1371 ), .Z(\GFM/n8580 ) );
XOR2_X2 \GFM/U3609  ( .A(\GFM/N1365 ), .B(\GFM/N1367 ), .Z(\GFM/n859 ) );
XOR2_X2 \GFM/U3608  ( .A(\GFM/n8610 ), .B(\GFM/n860 ), .Z(z_out[45]) );
XOR2_X2 \GFM/U3607  ( .A(\GFM/n863 ), .B(\GFM/n8620 ), .Z(\GFM/n860 ) );
XOR2_X2 \GFM/U3606  ( .A(\GFM/n8650 ), .B(\GFM/n8640 ), .Z(\GFM/n8610 ) );
XOR2_X2 \GFM/U3605  ( .A(\GFM/n867 ), .B(\GFM/n866 ), .Z(\GFM/n8620 ) );
XOR2_X2 \GFM/U3604  ( .A(\GFM/n8690 ), .B(\GFM/n868 ), .Z(\GFM/n863 ) );
XOR2_X2 \GFM/U3603  ( .A(\GFM/n8710 ), .B(\GFM/n870 ), .Z(\GFM/n8640 ) );
XOR2_X2 \GFM/U3602  ( .A(\GFM/n873 ), .B(\GFM/n8720 ), .Z(\GFM/n8650 ) );
XOR2_X2 \GFM/U3601  ( .A(z_in[45]), .B(\GFM/n874 ), .Z(\GFM/n866 ) );
XOR2_X2 \GFM/U3600  ( .A(\GFM/N1422 ), .B(\GFM/N1423 ), .Z(\GFM/n867 ) );
XOR2_X2 \GFM/U3599  ( .A(\GFM/N1419 ), .B(\GFM/N1420 ), .Z(\GFM/n868 ) );
XOR2_X2 \GFM/U3598  ( .A(\GFM/N1415 ), .B(\GFM/N1416 ), .Z(\GFM/n8690 ) );
XOR2_X2 \GFM/U3597  ( .A(\GFM/N1411 ), .B(\GFM/N1413 ), .Z(\GFM/n870 ) );
XOR2_X2 \GFM/U3596  ( .A(\GFM/N1406 ), .B(\GFM/N1410 ), .Z(\GFM/n8710 ) );
XOR2_X2 \GFM/U3595  ( .A(\GFM/N1403 ), .B(\GFM/N1405 ), .Z(\GFM/n8720 ) );
XOR2_X2 \GFM/U3594  ( .A(\GFM/N1399 ), .B(\GFM/N1402 ), .Z(\GFM/n873 ) );
XOR2_X2 \GFM/U3593  ( .A(\GFM/N1396 ), .B(\GFM/N1398 ), .Z(\GFM/n874 ) );
XOR2_X2 \GFM/U3592  ( .A(\GFM/n8760 ), .B(\GFM/n8750 ), .Z(z_out[46]) );
XOR2_X2 \GFM/U3591  ( .A(\GFM/n8780 ), .B(\GFM/n877 ), .Z(\GFM/n8750 ) );
XOR2_X2 \GFM/U3590  ( .A(\GFM/n880 ), .B(\GFM/n8790 ), .Z(\GFM/n8760 ) );
XOR2_X2 \GFM/U3589  ( .A(\GFM/n882 ), .B(\GFM/n881 ), .Z(\GFM/n877 ) );
XOR2_X2 \GFM/U3588  ( .A(\GFM/n8840 ), .B(\GFM/n8830 ), .Z(\GFM/n8780 ) );
XOR2_X2 \GFM/U3587  ( .A(\GFM/n8860 ), .B(\GFM/n885 ), .Z(\GFM/n8790 ) );
XOR2_X2 \GFM/U3586  ( .A(\GFM/n8880 ), .B(\GFM/n887 ), .Z(\GFM/n880 ) );
XOR2_X2 \GFM/U3585  ( .A(z_in[46]), .B(\GFM/n8890 ), .Z(\GFM/n881 ) );
XOR2_X2 \GFM/U3584  ( .A(\GFM/N1453 ), .B(\GFM/N1454 ), .Z(\GFM/n882 ) );
XOR2_X2 \GFM/U3583  ( .A(\GFM/N1450 ), .B(\GFM/N1451 ), .Z(\GFM/n8830 ) );
XOR2_X2 \GFM/U3582  ( .A(\GFM/N1446 ), .B(\GFM/N1447 ), .Z(\GFM/n8840 ) );
XOR2_X2 \GFM/U3581  ( .A(\GFM/N1442 ), .B(\GFM/N1444 ), .Z(\GFM/n885 ) );
XOR2_X2 \GFM/U3580  ( .A(\GFM/N1437 ), .B(\GFM/N1441 ), .Z(\GFM/n8860 ) );
XOR2_X2 \GFM/U3579  ( .A(\GFM/N1434 ), .B(\GFM/N1436 ), .Z(\GFM/n887 ) );
XOR2_X2 \GFM/U3578  ( .A(\GFM/N1430 ), .B(\GFM/N1433 ), .Z(\GFM/n8880 ) );
XOR2_X2 \GFM/U3577  ( .A(\GFM/N1427 ), .B(\GFM/N1429 ), .Z(\GFM/n8890 ) );
XOR2_X2 \GFM/U3576  ( .A(\GFM/n891 ), .B(\GFM/n890 ), .Z(z_out[47]) );
XOR2_X2 \GFM/U3575  ( .A(\GFM/n8930 ), .B(\GFM/n8920 ), .Z(\GFM/n890 ) );
XOR2_X2 \GFM/U3574  ( .A(\GFM/n8950 ), .B(\GFM/n894 ), .Z(\GFM/n891 ) );
XOR2_X2 \GFM/U3573  ( .A(\GFM/n897 ), .B(\GFM/n8960 ), .Z(\GFM/n8920 ) );
XOR2_X2 \GFM/U3572  ( .A(\GFM/n899 ), .B(\GFM/n898 ), .Z(\GFM/n8930 ) );
XOR2_X2 \GFM/U3571  ( .A(\GFM/n901 ), .B(\GFM/n9000 ), .Z(\GFM/n894 ) );
XOR2_X2 \GFM/U3570  ( .A(\GFM/n9030 ), .B(\GFM/n9020 ), .Z(\GFM/n8950 ) );
XOR2_X2 \GFM/U3569  ( .A(z_in[47]), .B(\GFM/n904 ), .Z(\GFM/n8960 ) );
XOR2_X2 \GFM/U3568  ( .A(\GFM/N1484 ), .B(\GFM/N1485 ), .Z(\GFM/n897 ) );
XOR2_X2 \GFM/U3567  ( .A(\GFM/N1481 ), .B(\GFM/N1482 ), .Z(\GFM/n898 ) );
XOR2_X2 \GFM/U3566  ( .A(\GFM/N1477 ), .B(\GFM/N1478 ), .Z(\GFM/n899 ) );
XOR2_X2 \GFM/U3565  ( .A(\GFM/N1473 ), .B(\GFM/N1475 ), .Z(\GFM/n9000 ) );
XOR2_X2 \GFM/U3564  ( .A(\GFM/N1468 ), .B(\GFM/N1472 ), .Z(\GFM/n901 ) );
XOR2_X2 \GFM/U3563  ( .A(\GFM/N1465 ), .B(\GFM/N1467 ), .Z(\GFM/n9020 ) );
XOR2_X2 \GFM/U3562  ( .A(\GFM/N1461 ), .B(\GFM/N1464 ), .Z(\GFM/n9030 ) );
XOR2_X2 \GFM/U3561  ( .A(\GFM/N1458 ), .B(\GFM/N1460 ), .Z(\GFM/n904 ) );
XOR2_X2 \GFM/U3560  ( .A(\GFM/n9060 ), .B(\GFM/n905 ), .Z(z_out[48]) );
XOR2_X2 \GFM/U3559  ( .A(\GFM/n908 ), .B(\GFM/n9070 ), .Z(\GFM/n905 ) );
XOR2_X2 \GFM/U3558  ( .A(\GFM/n9100 ), .B(\GFM/n9090 ), .Z(\GFM/n9060 ) );
XOR2_X2 \GFM/U3557  ( .A(\GFM/n912 ), .B(\GFM/n911 ), .Z(\GFM/n9070 ) );
XOR2_X2 \GFM/U3556  ( .A(\GFM/n9140 ), .B(\GFM/n913 ), .Z(\GFM/n908 ) );
XOR2_X2 \GFM/U3555  ( .A(\GFM/n916 ), .B(\GFM/n9150 ), .Z(\GFM/n9090 ) );
XOR2_X2 \GFM/U3554  ( .A(\GFM/n918 ), .B(\GFM/n9170 ), .Z(\GFM/n9100 ) );
XOR2_X2 \GFM/U3553  ( .A(z_in[48]), .B(\GFM/n9190 ), .Z(\GFM/n911 ) );
XOR2_X2 \GFM/U3552  ( .A(\GFM/N1515 ), .B(\GFM/N1516 ), .Z(\GFM/n912 ) );
XOR2_X2 \GFM/U3551  ( .A(\GFM/N1512 ), .B(\GFM/N1513 ), .Z(\GFM/n913 ) );
XOR2_X2 \GFM/U3550  ( .A(\GFM/N1508 ), .B(\GFM/N1509 ), .Z(\GFM/n9140 ) );
XOR2_X2 \GFM/U3549  ( .A(\GFM/N1504 ), .B(\GFM/N1506 ), .Z(\GFM/n9150 ) );
XOR2_X2 \GFM/U3548  ( .A(\GFM/N1499 ), .B(\GFM/N1503 ), .Z(\GFM/n916 ) );
XOR2_X2 \GFM/U3547  ( .A(\GFM/N1496 ), .B(\GFM/N1498 ), .Z(\GFM/n9170 ) );
XOR2_X2 \GFM/U3546  ( .A(\GFM/N1492 ), .B(\GFM/N1495 ), .Z(\GFM/n918 ) );
XOR2_X2 \GFM/U3545  ( .A(\GFM/N1489 ), .B(\GFM/N1491 ), .Z(\GFM/n9190 ) );
XOR2_X2 \GFM/U3544  ( .A(\GFM/n921 ), .B(\GFM/n9200 ), .Z(z_out[49]) );
XOR2_X2 \GFM/U3543  ( .A(\GFM/n9230 ), .B(\GFM/n922 ), .Z(\GFM/n9200 ) );
XOR2_X2 \GFM/U3542  ( .A(\GFM/n925 ), .B(\GFM/n9240 ), .Z(\GFM/n921 ) );
XOR2_X2 \GFM/U3541  ( .A(\GFM/n9270 ), .B(\GFM/n9260 ), .Z(\GFM/n922 ) );
XOR2_X2 \GFM/U3540  ( .A(\GFM/n929 ), .B(\GFM/n928 ), .Z(\GFM/n9230 ) );
XOR2_X2 \GFM/U3539  ( .A(\GFM/n9310 ), .B(\GFM/n930 ), .Z(\GFM/n9240 ) );
XOR2_X2 \GFM/U3538  ( .A(\GFM/n9330 ), .B(\GFM/n932 ), .Z(\GFM/n925 ) );
XOR2_X2 \GFM/U3537  ( .A(z_in[49]), .B(\GFM/n9340 ), .Z(\GFM/n9260 ) );
XOR2_X2 \GFM/U3536  ( .A(\GFM/N1546 ), .B(\GFM/N1547 ), .Z(\GFM/n9270 ) );
XOR2_X2 \GFM/U3535  ( .A(\GFM/N1543 ), .B(\GFM/N1544 ), .Z(\GFM/n928 ) );
XOR2_X2 \GFM/U3534  ( .A(\GFM/N1539 ), .B(\GFM/N1540 ), .Z(\GFM/n929 ) );
XOR2_X2 \GFM/U3533  ( .A(\GFM/N1535 ), .B(\GFM/N1537 ), .Z(\GFM/n930 ) );
XOR2_X2 \GFM/U3532  ( .A(\GFM/N1530 ), .B(\GFM/N1534 ), .Z(\GFM/n9310 ) );
XOR2_X2 \GFM/U3531  ( .A(\GFM/N1527 ), .B(\GFM/N1529 ), .Z(\GFM/n932 ) );
XOR2_X2 \GFM/U3530  ( .A(\GFM/N1523 ), .B(\GFM/N1526 ), .Z(\GFM/n9330 ) );
XOR2_X2 \GFM/U3529  ( .A(\GFM/N1520 ), .B(\GFM/N1522 ), .Z(\GFM/n9340 ) );
XOR2_X2 \GFM/U3528  ( .A(\GFM/n936 ), .B(\GFM/n935 ), .Z(z_out[50]) );
XOR2_X2 \GFM/U3527  ( .A(\GFM/n9380 ), .B(\GFM/n9370 ), .Z(\GFM/n935 ) );
XOR2_X2 \GFM/U3526  ( .A(\GFM/n9400 ), .B(\GFM/n939 ), .Z(\GFM/n936 ) );
XOR2_X2 \GFM/U3525  ( .A(\GFM/n942 ), .B(\GFM/n9410 ), .Z(\GFM/n9370 ) );
XOR2_X2 \GFM/U3524  ( .A(\GFM/n944 ), .B(\GFM/n943 ), .Z(\GFM/n9380 ) );
XOR2_X2 \GFM/U3523  ( .A(\GFM/n9460 ), .B(\GFM/n9450 ), .Z(\GFM/n939 ) );
XOR2_X2 \GFM/U3522  ( .A(\GFM/n9480 ), .B(\GFM/n947 ), .Z(\GFM/n9400 ) );
XOR2_X2 \GFM/U3521  ( .A(z_in[50]), .B(\GFM/n949 ), .Z(\GFM/n9410 ) );
XOR2_X2 \GFM/U3520  ( .A(\GFM/N1577 ), .B(\GFM/N1578 ), .Z(\GFM/n942 ) );
XOR2_X2 \GFM/U3519  ( .A(\GFM/N1574 ), .B(\GFM/N1575 ), .Z(\GFM/n943 ) );
XOR2_X2 \GFM/U3518  ( .A(\GFM/N1570 ), .B(\GFM/N1571 ), .Z(\GFM/n944 ) );
XOR2_X2 \GFM/U3517  ( .A(\GFM/N1566 ), .B(\GFM/N1568 ), .Z(\GFM/n9450 ) );
XOR2_X2 \GFM/U3516  ( .A(\GFM/N1561 ), .B(\GFM/N1565 ), .Z(\GFM/n9460 ) );
XOR2_X2 \GFM/U3515  ( .A(\GFM/N1558 ), .B(\GFM/N1560 ), .Z(\GFM/n947 ) );
XOR2_X2 \GFM/U3514  ( .A(\GFM/N1554 ), .B(\GFM/N1557 ), .Z(\GFM/n9480 ) );
XOR2_X2 \GFM/U3513  ( .A(\GFM/N1551 ), .B(\GFM/N1553 ), .Z(\GFM/n949 ) );
XOR2_X2 \GFM/U3512  ( .A(\GFM/n9510 ), .B(\GFM/n9500 ), .Z(z_out[51]) );
XOR2_X2 \GFM/U3511  ( .A(\GFM/n953 ), .B(\GFM/n952 ), .Z(\GFM/n9500 ) );
XOR2_X2 \GFM/U3510  ( .A(\GFM/n9550 ), .B(\GFM/n9540 ), .Z(\GFM/n9510 ) );
XOR2_X2 \GFM/U3509  ( .A(\GFM/n9570 ), .B(\GFM/n956 ), .Z(\GFM/n952 ) );
XOR2_X2 \GFM/U3508  ( .A(\GFM/n959 ), .B(\GFM/n9580 ), .Z(\GFM/n953 ) );
XOR2_X2 \GFM/U3507  ( .A(\GFM/n961 ), .B(\GFM/n960 ), .Z(\GFM/n9540 ) );
XOR2_X2 \GFM/U3506  ( .A(\GFM/n963 ), .B(\GFM/n9620 ), .Z(\GFM/n9550 ) );
XOR2_X2 \GFM/U3505  ( .A(z_in[51]), .B(\GFM/n9640 ), .Z(\GFM/n956 ) );
XOR2_X2 \GFM/U3504  ( .A(\GFM/N1608 ), .B(\GFM/N1609 ), .Z(\GFM/n9570 ) );
XOR2_X2 \GFM/U3503  ( .A(\GFM/N1605 ), .B(\GFM/N1606 ), .Z(\GFM/n9580 ) );
XOR2_X2 \GFM/U3502  ( .A(\GFM/N1601 ), .B(\GFM/N1602 ), .Z(\GFM/n959 ) );
XOR2_X2 \GFM/U3501  ( .A(\GFM/N1597 ), .B(\GFM/N1599 ), .Z(\GFM/n960 ) );
XOR2_X2 \GFM/U3500  ( .A(\GFM/N1592 ), .B(\GFM/N1596 ), .Z(\GFM/n961 ) );
XOR2_X2 \GFM/U3499  ( .A(\GFM/N1589 ), .B(\GFM/N1591 ), .Z(\GFM/n9620 ) );
XOR2_X2 \GFM/U3498  ( .A(\GFM/N1585 ), .B(\GFM/N1588 ), .Z(\GFM/n963 ) );
XOR2_X2 \GFM/U3497  ( .A(\GFM/N1582 ), .B(\GFM/N1584 ), .Z(\GFM/n9640 ) );
XOR2_X2 \GFM/U3496  ( .A(\GFM/n966 ), .B(\GFM/n9650 ), .Z(z_out[52]) );
XOR2_X2 \GFM/U3495  ( .A(\GFM/n9680 ), .B(\GFM/n967 ), .Z(\GFM/n9650 ) );
XOR2_X2 \GFM/U3494  ( .A(\GFM/n970 ), .B(\GFM/n9690 ), .Z(\GFM/n966 ) );
XOR2_X2 \GFM/U3493  ( .A(\GFM/n9720 ), .B(\GFM/n9710 ), .Z(\GFM/n967 ) );
XOR2_X2 \GFM/U3492  ( .A(\GFM/n974 ), .B(\GFM/n973 ), .Z(\GFM/n9680 ) );
XOR2_X2 \GFM/U3491  ( .A(\GFM/n9760 ), .B(\GFM/n975 ), .Z(\GFM/n9690 ) );
XOR2_X2 \GFM/U3490  ( .A(\GFM/n978 ), .B(\GFM/n9770 ), .Z(\GFM/n970 ) );
XOR2_X2 \GFM/U3489  ( .A(z_in[52]), .B(\GFM/n9790 ), .Z(\GFM/n9710 ) );
XOR2_X2 \GFM/U3488  ( .A(\GFM/N1639 ), .B(\GFM/N1640 ), .Z(\GFM/n9720 ) );
XOR2_X2 \GFM/U3487  ( .A(\GFM/N1636 ), .B(\GFM/N1637 ), .Z(\GFM/n973 ) );
XOR2_X2 \GFM/U3486  ( .A(\GFM/N1632 ), .B(\GFM/N1633 ), .Z(\GFM/n974 ) );
XOR2_X2 \GFM/U3485  ( .A(\GFM/N1628 ), .B(\GFM/N1630 ), .Z(\GFM/n975 ) );
XOR2_X2 \GFM/U3484  ( .A(\GFM/N1623 ), .B(\GFM/N1627 ), .Z(\GFM/n9760 ) );
XOR2_X2 \GFM/U3483  ( .A(\GFM/N1620 ), .B(\GFM/N1622 ), .Z(\GFM/n9770 ) );
XOR2_X2 \GFM/U3482  ( .A(\GFM/N1616 ), .B(\GFM/N1619 ), .Z(\GFM/n978 ) );
XOR2_X2 \GFM/U3481  ( .A(\GFM/N1613 ), .B(\GFM/N1615 ), .Z(\GFM/n9790 ) );
XOR2_X2 \GFM/U3480  ( .A(\GFM/n9810 ), .B(\GFM/n980 ), .Z(z_out[53]) );
XOR2_X2 \GFM/U3479  ( .A(\GFM/n983 ), .B(\GFM/n9820 ), .Z(\GFM/n980 ) );
XOR2_X2 \GFM/U3478  ( .A(\GFM/n9850 ), .B(\GFM/n984 ), .Z(\GFM/n9810 ) );
XOR2_X2 \GFM/U3477  ( .A(\GFM/n987 ), .B(\GFM/n9860 ), .Z(\GFM/n9820 ) );
XOR2_X2 \GFM/U3476  ( .A(\GFM/n9890 ), .B(\GFM/n9880 ), .Z(\GFM/n983 ) );
XOR2_X2 \GFM/U3475  ( .A(\GFM/n991 ), .B(\GFM/n990 ), .Z(\GFM/n984 ) );
XOR2_X2 \GFM/U3474  ( .A(\GFM/n9930 ), .B(\GFM/n992 ), .Z(\GFM/n9850 ) );
XOR2_X2 \GFM/U3473  ( .A(z_in[53]), .B(\GFM/n994 ), .Z(\GFM/n9860 ) );
XOR2_X2 \GFM/U3472  ( .A(\GFM/N1670 ), .B(\GFM/N1671 ), .Z(\GFM/n987 ) );
XOR2_X2 \GFM/U3471  ( .A(\GFM/N1667 ), .B(\GFM/N1668 ), .Z(\GFM/n9880 ) );
XOR2_X2 \GFM/U3470  ( .A(\GFM/N1663 ), .B(\GFM/N1664 ), .Z(\GFM/n9890 ) );
XOR2_X2 \GFM/U3469  ( .A(\GFM/N1659 ), .B(\GFM/N1661 ), .Z(\GFM/n990 ) );
XOR2_X2 \GFM/U3468  ( .A(\GFM/N1654 ), .B(\GFM/N1658 ), .Z(\GFM/n991 ) );
XOR2_X2 \GFM/U3467  ( .A(\GFM/N1651 ), .B(\GFM/N1653 ), .Z(\GFM/n992 ) );
XOR2_X2 \GFM/U3466  ( .A(\GFM/N1647 ), .B(\GFM/N1650 ), .Z(\GFM/n9930 ) );
XOR2_X2 \GFM/U3465  ( .A(\GFM/N1644 ), .B(\GFM/N1646 ), .Z(\GFM/n994 ) );
XOR2_X2 \GFM/U3464  ( .A(\GFM/n9960 ), .B(\GFM/n9950 ), .Z(z_out[54]) );
XOR2_X2 \GFM/U3463  ( .A(\GFM/n998 ), .B(\GFM/n997 ), .Z(\GFM/n9950 ) );
XOR2_X2 \GFM/U3462  ( .A(\GFM/n10000 ), .B(\GFM/n9990 ), .Z(\GFM/n9960 ) );
XOR2_X2 \GFM/U3461  ( .A(\GFM/n10020 ), .B(\GFM/n1001 ), .Z(\GFM/n997 ) );
XOR2_X2 \GFM/U3460  ( .A(\GFM/n1004 ), .B(\GFM/n10030 ), .Z(\GFM/n998 ) );
XOR2_X2 \GFM/U3459  ( .A(\GFM/n1006 ), .B(\GFM/n1005 ), .Z(\GFM/n9990 ) );
XOR2_X2 \GFM/U3458  ( .A(\GFM/n10080 ), .B(\GFM/n10070 ), .Z(\GFM/n10000 ));
XOR2_X2 \GFM/U3457  ( .A(z_in[54]), .B(\GFM/n1009 ), .Z(\GFM/n1001 ) );
XOR2_X2 \GFM/U3456  ( .A(\GFM/N1701 ), .B(\GFM/N1702 ), .Z(\GFM/n10020 ) );
XOR2_X2 \GFM/U3455  ( .A(\GFM/N1698 ), .B(\GFM/N1699 ), .Z(\GFM/n10030 ) );
XOR2_X2 \GFM/U3454  ( .A(\GFM/N1694 ), .B(\GFM/N1695 ), .Z(\GFM/n1004 ) );
XOR2_X2 \GFM/U3453  ( .A(\GFM/N1690 ), .B(\GFM/N1692 ), .Z(\GFM/n1005 ) );
XOR2_X2 \GFM/U3452  ( .A(\GFM/N1685 ), .B(\GFM/N1689 ), .Z(\GFM/n1006 ) );
XOR2_X2 \GFM/U3451  ( .A(\GFM/N1682 ), .B(\GFM/N1684 ), .Z(\GFM/n10070 ) );
XOR2_X2 \GFM/U3450  ( .A(\GFM/N1678 ), .B(\GFM/N1681 ), .Z(\GFM/n10080 ) );
XOR2_X2 \GFM/U3449  ( .A(\GFM/N1675 ), .B(\GFM/N1677 ), .Z(\GFM/n1009 ) );
XOR2_X2 \GFM/U3448  ( .A(\GFM/n1011 ), .B(\GFM/n10100 ), .Z(z_out[55]) );
XOR2_X2 \GFM/U3447  ( .A(\GFM/n10130 ), .B(\GFM/n10120 ), .Z(\GFM/n10100 ));
XOR2_X2 \GFM/U3446  ( .A(\GFM/n1015 ), .B(\GFM/n1014 ), .Z(\GFM/n1011 ) );
XOR2_X2 \GFM/U3445  ( .A(\GFM/n10170 ), .B(\GFM/n10160 ), .Z(\GFM/n10120 ));
XOR2_X2 \GFM/U3444  ( .A(\GFM/n10190 ), .B(\GFM/n1018 ), .Z(\GFM/n10130 ) );
XOR2_X2 \GFM/U3443  ( .A(\GFM/n1021 ), .B(\GFM/n10200 ), .Z(\GFM/n1014 ) );
XOR2_X2 \GFM/U3442  ( .A(\GFM/n1023 ), .B(\GFM/n1022 ), .Z(\GFM/n1015 ) );
XOR2_X2 \GFM/U3441  ( .A(z_in[55]), .B(\GFM/n10240 ), .Z(\GFM/n10160 ) );
XOR2_X2 \GFM/U3440  ( .A(\GFM/N1732 ), .B(\GFM/N1733 ), .Z(\GFM/n10170 ) );
XOR2_X2 \GFM/U3439  ( .A(\GFM/N1729 ), .B(\GFM/N1730 ), .Z(\GFM/n1018 ) );
XOR2_X2 \GFM/U3438  ( .A(\GFM/N1725 ), .B(\GFM/N1726 ), .Z(\GFM/n10190 ) );
XOR2_X2 \GFM/U3437  ( .A(\GFM/N1721 ), .B(\GFM/N1723 ), .Z(\GFM/n10200 ) );
XOR2_X2 \GFM/U3436  ( .A(\GFM/N1716 ), .B(\GFM/N1720 ), .Z(\GFM/n1021 ) );
XOR2_X2 \GFM/U3435  ( .A(\GFM/N1713 ), .B(\GFM/N1715 ), .Z(\GFM/n1022 ) );
XOR2_X2 \GFM/U3434  ( .A(\GFM/N1709 ), .B(\GFM/N1712 ), .Z(\GFM/n1023 ) );
XOR2_X2 \GFM/U3433  ( .A(\GFM/N1706 ), .B(\GFM/N1708 ), .Z(\GFM/n10240 ) );
XOR2_X2 \GFM/U3432  ( .A(\GFM/n10260 ), .B(\GFM/n1025 ), .Z(z_out[56]) );
XOR2_X2 \GFM/U3431  ( .A(\GFM/n1028 ), .B(\GFM/n10270 ), .Z(\GFM/n1025 ) );
XOR2_X2 \GFM/U3430  ( .A(\GFM/n10300 ), .B(\GFM/n1029 ), .Z(\GFM/n10260 ) );
XOR2_X2 \GFM/U3429  ( .A(\GFM/n1032 ), .B(\GFM/n10310 ), .Z(\GFM/n10270 ) );
XOR2_X2 \GFM/U3428  ( .A(\GFM/n10340 ), .B(\GFM/n10330 ), .Z(\GFM/n1028 ) );
XOR2_X2 \GFM/U3427  ( .A(\GFM/n1036 ), .B(\GFM/n1035 ), .Z(\GFM/n1029 ) );
XOR2_X2 \GFM/U3426  ( .A(\GFM/n10380 ), .B(\GFM/n1037 ), .Z(\GFM/n10300 ) );
XOR2_X2 \GFM/U3425  ( .A(z_in[56]), .B(\GFM/n10390 ), .Z(\GFM/n10310 ) );
XOR2_X2 \GFM/U3424  ( .A(\GFM/N1763 ), .B(\GFM/N1764 ), .Z(\GFM/n1032 ) );
XOR2_X2 \GFM/U3423  ( .A(\GFM/N1760 ), .B(\GFM/N1761 ), .Z(\GFM/n10330 ) );
XOR2_X2 \GFM/U3422  ( .A(\GFM/N1756 ), .B(\GFM/N1757 ), .Z(\GFM/n10340 ) );
XOR2_X2 \GFM/U3421  ( .A(\GFM/N1752 ), .B(\GFM/N1754 ), .Z(\GFM/n1035 ) );
XOR2_X2 \GFM/U3420  ( .A(\GFM/N1747 ), .B(\GFM/N1751 ), .Z(\GFM/n1036 ) );
XOR2_X2 \GFM/U3419  ( .A(\GFM/N1744 ), .B(\GFM/N1746 ), .Z(\GFM/n1037 ) );
XOR2_X2 \GFM/U3418  ( .A(\GFM/N1740 ), .B(\GFM/N1743 ), .Z(\GFM/n10380 ) );
XOR2_X2 \GFM/U3417  ( .A(\GFM/N1737 ), .B(\GFM/N1739 ), .Z(\GFM/n10390 ) );
XOR2_X2 \GFM/U3416  ( .A(\GFM/n10410 ), .B(\GFM/n1040 ), .Z(z_out[57]) );
XOR2_X2 \GFM/U3415  ( .A(\GFM/n10430 ), .B(\GFM/n1042 ), .Z(\GFM/n1040 ) );
XOR2_X2 \GFM/U3414  ( .A(\GFM/n1045 ), .B(\GFM/n10440 ), .Z(\GFM/n10410 ) );
XOR2_X2 \GFM/U3413  ( .A(\GFM/n10470 ), .B(\GFM/n1046 ), .Z(\GFM/n1042 ) );
XOR2_X2 \GFM/U3412  ( .A(\GFM/n1049 ), .B(\GFM/n10480 ), .Z(\GFM/n10430 ) );
XOR2_X2 \GFM/U3411  ( .A(\GFM/n10510 ), .B(\GFM/n10500 ), .Z(\GFM/n10440 ));
XOR2_X2 \GFM/U3410  ( .A(\GFM/n1053 ), .B(\GFM/n1052 ), .Z(\GFM/n1045 ) );
XOR2_X2 \GFM/U3409  ( .A(z_in[57]), .B(\GFM/n1054 ), .Z(\GFM/n1046 ) );
XOR2_X2 \GFM/U3408  ( .A(\GFM/N1794 ), .B(\GFM/N1795 ), .Z(\GFM/n10470 ) );
XOR2_X2 \GFM/U3407  ( .A(\GFM/N1791 ), .B(\GFM/N1792 ), .Z(\GFM/n10480 ) );
XOR2_X2 \GFM/U3406  ( .A(\GFM/N1787 ), .B(\GFM/N1788 ), .Z(\GFM/n1049 ) );
XOR2_X2 \GFM/U3405  ( .A(\GFM/N1783 ), .B(\GFM/N1785 ), .Z(\GFM/n10500 ) );
XOR2_X2 \GFM/U3404  ( .A(\GFM/N1778 ), .B(\GFM/N1782 ), .Z(\GFM/n10510 ) );
XOR2_X2 \GFM/U3403  ( .A(\GFM/N1775 ), .B(\GFM/N1777 ), .Z(\GFM/n1052 ) );
XOR2_X2 \GFM/U3402  ( .A(\GFM/N1771 ), .B(\GFM/N1774 ), .Z(\GFM/n1053 ) );
XOR2_X2 \GFM/U3401  ( .A(\GFM/N1768 ), .B(\GFM/N1770 ), .Z(\GFM/n1054 ) );
XOR2_X2 \GFM/U3400  ( .A(\GFM/n1056 ), .B(\GFM/n10550 ), .Z(z_out[58]) );
XOR2_X2 \GFM/U3399  ( .A(\GFM/n10580 ), .B(\GFM/n10570 ), .Z(\GFM/n10550 ));
XOR2_X2 \GFM/U3398  ( .A(\GFM/n1060 ), .B(\GFM/n1059 ), .Z(\GFM/n1056 ) );
XOR2_X2 \GFM/U3397  ( .A(\GFM/n10620 ), .B(\GFM/n10610 ), .Z(\GFM/n10570 ));
XOR2_X2 \GFM/U3396  ( .A(\GFM/n10640 ), .B(\GFM/n1063 ), .Z(\GFM/n10580 ) );
XOR2_X2 \GFM/U3395  ( .A(\GFM/n1066 ), .B(\GFM/n10650 ), .Z(\GFM/n1059 ) );
XOR2_X2 \GFM/U3394  ( .A(\GFM/n1068 ), .B(\GFM/n1067 ), .Z(\GFM/n1060 ) );
XOR2_X2 \GFM/U3393  ( .A(z_in[58]), .B(\GFM/n10690 ), .Z(\GFM/n10610 ) );
XOR2_X2 \GFM/U3392  ( .A(\GFM/N1825 ), .B(\GFM/N1826 ), .Z(\GFM/n10620 ) );
XOR2_X2 \GFM/U3391  ( .A(\GFM/N1822 ), .B(\GFM/N1823 ), .Z(\GFM/n1063 ) );
XOR2_X2 \GFM/U3390  ( .A(\GFM/N1818 ), .B(\GFM/N1819 ), .Z(\GFM/n10640 ) );
XOR2_X2 \GFM/U3389  ( .A(\GFM/N1814 ), .B(\GFM/N1816 ), .Z(\GFM/n10650 ) );
XOR2_X2 \GFM/U3388  ( .A(\GFM/N1809 ), .B(\GFM/N1813 ), .Z(\GFM/n1066 ) );
XOR2_X2 \GFM/U3387  ( .A(\GFM/N1806 ), .B(\GFM/N1808 ), .Z(\GFM/n1067 ) );
XOR2_X2 \GFM/U3386  ( .A(\GFM/N1802 ), .B(\GFM/N1805 ), .Z(\GFM/n1068 ) );
XOR2_X2 \GFM/U3385  ( .A(\GFM/N1799 ), .B(\GFM/N1801 ), .Z(\GFM/n10690 ) );
XOR2_X2 \GFM/U3384  ( .A(\GFM/n1071 ), .B(\GFM/n10700 ), .Z(z_out[59]) );
XOR2_X2 \GFM/U3383  ( .A(\GFM/n1073 ), .B(\GFM/n10720 ), .Z(\GFM/n10700 ) );
XOR2_X2 \GFM/U3382  ( .A(\GFM/n10750 ), .B(\GFM/n10740 ), .Z(\GFM/n1071 ) );
XOR2_X2 \GFM/U3381  ( .A(\GFM/n1077 ), .B(\GFM/n1076 ), .Z(\GFM/n10720 ) );
XOR2_X2 \GFM/U3380  ( .A(\GFM/n10790 ), .B(\GFM/n10780 ), .Z(\GFM/n1073 ) );
XOR2_X2 \GFM/U3379  ( .A(\GFM/n10810 ), .B(\GFM/n1080 ), .Z(\GFM/n10740 ) );
XOR2_X2 \GFM/U3378  ( .A(\GFM/n1083 ), .B(\GFM/n10820 ), .Z(\GFM/n10750 ) );
XOR2_X2 \GFM/U3377  ( .A(z_in[59]), .B(\GFM/n1084 ), .Z(\GFM/n1076 ) );
XOR2_X2 \GFM/U3376  ( .A(\GFM/N1856 ), .B(\GFM/N1857 ), .Z(\GFM/n1077 ) );
XOR2_X2 \GFM/U3375  ( .A(\GFM/N1853 ), .B(\GFM/N1854 ), .Z(\GFM/n10780 ) );
XOR2_X2 \GFM/U3374  ( .A(\GFM/N1849 ), .B(\GFM/N1850 ), .Z(\GFM/n10790 ) );
XOR2_X2 \GFM/U3373  ( .A(\GFM/N1845 ), .B(\GFM/N1847 ), .Z(\GFM/n1080 ) );
XOR2_X2 \GFM/U3372  ( .A(\GFM/N1840 ), .B(\GFM/N1844 ), .Z(\GFM/n10810 ) );
XOR2_X2 \GFM/U3371  ( .A(\GFM/N1837 ), .B(\GFM/N1839 ), .Z(\GFM/n10820 ) );
XOR2_X2 \GFM/U3370  ( .A(\GFM/N1833 ), .B(\GFM/N1836 ), .Z(\GFM/n1083 ) );
XOR2_X2 \GFM/U3369  ( .A(\GFM/N1830 ), .B(\GFM/N1832 ), .Z(\GFM/n1084 ) );
XOR2_X2 \GFM/U3368  ( .A(\GFM/n10860 ), .B(\GFM/n1085 ), .Z(z_out[60]) );
XOR2_X2 \GFM/U3367  ( .A(\GFM/n10880 ), .B(\GFM/n1087 ), .Z(\GFM/n1085 ) );
XOR2_X2 \GFM/U3366  ( .A(\GFM/n1090 ), .B(\GFM/n10890 ), .Z(\GFM/n10860 ) );
XOR2_X2 \GFM/U3365  ( .A(\GFM/n10920 ), .B(\GFM/n1091 ), .Z(\GFM/n1087 ) );
XOR2_X2 \GFM/U3364  ( .A(\GFM/n1094 ), .B(\GFM/n10930 ), .Z(\GFM/n10880 ) );
XOR2_X2 \GFM/U3363  ( .A(\GFM/n10960 ), .B(\GFM/n10950 ), .Z(\GFM/n10890 ));
XOR2_X2 \GFM/U3362  ( .A(\GFM/n1098 ), .B(\GFM/n1097 ), .Z(\GFM/n1090 ) );
XOR2_X2 \GFM/U3361  ( .A(z_in[60]), .B(\GFM/n1099 ), .Z(\GFM/n1091 ) );
XOR2_X2 \GFM/U3360  ( .A(\GFM/N1887 ), .B(\GFM/N1888 ), .Z(\GFM/n10920 ) );
XOR2_X2 \GFM/U3359  ( .A(\GFM/N1884 ), .B(\GFM/N1885 ), .Z(\GFM/n10930 ) );
XOR2_X2 \GFM/U3358  ( .A(\GFM/N1880 ), .B(\GFM/N1881 ), .Z(\GFM/n1094 ) );
XOR2_X2 \GFM/U3357  ( .A(\GFM/N1876 ), .B(\GFM/N1878 ), .Z(\GFM/n10950 ) );
XOR2_X2 \GFM/U3356  ( .A(\GFM/N1871 ), .B(\GFM/N1875 ), .Z(\GFM/n10960 ) );
XOR2_X2 \GFM/U3355  ( .A(\GFM/N1868 ), .B(\GFM/N1870 ), .Z(\GFM/n1097 ) );
XOR2_X2 \GFM/U3354  ( .A(\GFM/N1864 ), .B(\GFM/N1867 ), .Z(\GFM/n1098 ) );
XOR2_X2 \GFM/U3353  ( .A(\GFM/N1861 ), .B(\GFM/N1863 ), .Z(\GFM/n1099 ) );
XOR2_X2 \GFM/U3352  ( .A(\GFM/n11010 ), .B(\GFM/n11000 ), .Z(z_out[61]) );
XOR2_X2 \GFM/U3351  ( .A(\GFM/n11030 ), .B(\GFM/n1102 ), .Z(\GFM/n11000 ) );
XOR2_X2 \GFM/U3350  ( .A(\GFM/n11050 ), .B(\GFM/n1104 ), .Z(\GFM/n11010 ) );
XOR2_X2 \GFM/U3349  ( .A(\GFM/n1107 ), .B(\GFM/n11060 ), .Z(\GFM/n1102 ) );
XOR2_X2 \GFM/U3348  ( .A(\GFM/n11090 ), .B(\GFM/n1108 ), .Z(\GFM/n11030 ) );
XOR2_X2 \GFM/U3347  ( .A(\GFM/n1111 ), .B(\GFM/n11100 ), .Z(\GFM/n1104 ) );
XOR2_X2 \GFM/U3346  ( .A(\GFM/n11130 ), .B(\GFM/n11120 ), .Z(\GFM/n11050 ));
XOR2_X2 \GFM/U3345  ( .A(z_in[61]), .B(\GFM/n1114 ), .Z(\GFM/n11060 ) );
XOR2_X2 \GFM/U3344  ( .A(\GFM/N1918 ), .B(\GFM/N1919 ), .Z(\GFM/n1107 ) );
XOR2_X2 \GFM/U3343  ( .A(\GFM/N1915 ), .B(\GFM/N1916 ), .Z(\GFM/n1108 ) );
XOR2_X2 \GFM/U3342  ( .A(\GFM/N1911 ), .B(\GFM/N1912 ), .Z(\GFM/n11090 ) );
XOR2_X2 \GFM/U3341  ( .A(\GFM/N1907 ), .B(\GFM/N1909 ), .Z(\GFM/n11100 ) );
XOR2_X2 \GFM/U3340  ( .A(\GFM/N1902 ), .B(\GFM/N1906 ), .Z(\GFM/n1111 ) );
XOR2_X2 \GFM/U3339  ( .A(\GFM/N1899 ), .B(\GFM/N1901 ), .Z(\GFM/n11120 ) );
XOR2_X2 \GFM/U3338  ( .A(\GFM/N1895 ), .B(\GFM/N1898 ), .Z(\GFM/n11130 ) );
XOR2_X2 \GFM/U3337  ( .A(\GFM/N1892 ), .B(\GFM/N1894 ), .Z(\GFM/n1114 ) );
XOR2_X2 \GFM/U3336  ( .A(\GFM/n1116 ), .B(\GFM/n1115 ), .Z(z_out[62]) );
XOR2_X2 \GFM/U3335  ( .A(\GFM/n1118 ), .B(\GFM/n11170 ), .Z(\GFM/n1115 ) );
XOR2_X2 \GFM/U3334  ( .A(\GFM/n11200 ), .B(\GFM/n11190 ), .Z(\GFM/n1116 ) );
XOR2_X2 \GFM/U3333  ( .A(\GFM/n1122 ), .B(\GFM/n1121 ), .Z(\GFM/n11170 ) );
XOR2_X2 \GFM/U3332  ( .A(\GFM/n11240 ), .B(\GFM/n11230 ), .Z(\GFM/n1118 ) );
XOR2_X2 \GFM/U3331  ( .A(\GFM/n11260 ), .B(\GFM/n1125 ), .Z(\GFM/n11190 ) );
XOR2_X2 \GFM/U3330  ( .A(\GFM/n1128 ), .B(\GFM/n11270 ), .Z(\GFM/n11200 ) );
XOR2_X2 \GFM/U3329  ( .A(z_in[62]), .B(\GFM/n1129 ), .Z(\GFM/n1121 ) );
XOR2_X2 \GFM/U3328  ( .A(\GFM/N1949 ), .B(\GFM/N1950 ), .Z(\GFM/n1122 ) );
XOR2_X2 \GFM/U3327  ( .A(\GFM/N1946 ), .B(\GFM/N1947 ), .Z(\GFM/n11230 ) );
XOR2_X2 \GFM/U3326  ( .A(\GFM/N1942 ), .B(\GFM/N1943 ), .Z(\GFM/n11240 ) );
XOR2_X2 \GFM/U3325  ( .A(\GFM/N1938 ), .B(\GFM/N1940 ), .Z(\GFM/n1125 ) );
XOR2_X2 \GFM/U3324  ( .A(\GFM/N1933 ), .B(\GFM/N1937 ), .Z(\GFM/n11260 ) );
XOR2_X2 \GFM/U3323  ( .A(\GFM/N1930 ), .B(\GFM/N1932 ), .Z(\GFM/n11270 ) );
XOR2_X2 \GFM/U3322  ( .A(\GFM/N1926 ), .B(\GFM/N1929 ), .Z(\GFM/n1128 ) );
XOR2_X2 \GFM/U3321  ( .A(\GFM/N1923 ), .B(\GFM/N1925 ), .Z(\GFM/n1129 ) );
XOR2_X2 \GFM/U3320  ( .A(\GFM/n11310 ), .B(\GFM/n1130 ), .Z(z_out[63]) );
XOR2_X2 \GFM/U3319  ( .A(\GFM/n1133 ), .B(\GFM/n11320 ), .Z(\GFM/n1130 ) );
XOR2_X2 \GFM/U3318  ( .A(\GFM/n1135 ), .B(\GFM/n11340 ), .Z(\GFM/n11310 ) );
XOR2_X2 \GFM/U3317  ( .A(\GFM/n11370 ), .B(\GFM/n11360 ), .Z(\GFM/n11320 ));
XOR2_X2 \GFM/U3316  ( .A(\GFM/n1139 ), .B(\GFM/n1138 ), .Z(\GFM/n1133 ) );
XOR2_X2 \GFM/U3315  ( .A(\GFM/n11410 ), .B(\GFM/n11400 ), .Z(\GFM/n11340 ));
XOR2_X2 \GFM/U3314  ( .A(\GFM/n11430 ), .B(\GFM/n1142 ), .Z(\GFM/n1135 ) );
XOR2_X2 \GFM/U3313  ( .A(z_in[63]), .B(\GFM/n11440 ), .Z(\GFM/n11360 ) );
XOR2_X2 \GFM/U3312  ( .A(\GFM/N1980 ), .B(\GFM/N1981 ), .Z(\GFM/n11370 ) );
XOR2_X2 \GFM/U3311  ( .A(\GFM/N1977 ), .B(\GFM/N1978 ), .Z(\GFM/n1138 ) );
XOR2_X2 \GFM/U3310  ( .A(\GFM/N1973 ), .B(\GFM/N1974 ), .Z(\GFM/n1139 ) );
XOR2_X2 \GFM/U3309  ( .A(\GFM/N1969 ), .B(\GFM/N1971 ), .Z(\GFM/n11400 ) );
XOR2_X2 \GFM/U3308  ( .A(\GFM/N1964 ), .B(\GFM/N1968 ), .Z(\GFM/n11410 ) );
XOR2_X2 \GFM/U3307  ( .A(\GFM/N1961 ), .B(\GFM/N1963 ), .Z(\GFM/n1142 ) );
XOR2_X2 \GFM/U3306  ( .A(\GFM/N1957 ), .B(\GFM/N1960 ), .Z(\GFM/n11430 ) );
XOR2_X2 \GFM/U3305  ( .A(\GFM/N1954 ), .B(\GFM/N1956 ), .Z(\GFM/n11440 ) );
XOR2_X2 \GFM/U3304  ( .A(\GFM/n1146 ), .B(\GFM/n1145 ), .Z(z_out[64]) );
XOR2_X2 \GFM/U3303  ( .A(\GFM/n11480 ), .B(\GFM/n1147 ), .Z(\GFM/n1145 ) );
XOR2_X2 \GFM/U3302  ( .A(\GFM/n11500 ), .B(\GFM/n1149 ), .Z(\GFM/n1146 ) );
XOR2_X2 \GFM/U3301  ( .A(\GFM/n1152 ), .B(\GFM/n11510 ), .Z(\GFM/n1147 ) );
XOR2_X2 \GFM/U3300  ( .A(\GFM/n11540 ), .B(\GFM/n1153 ), .Z(\GFM/n11480 ) );
XOR2_X2 \GFM/U3299  ( .A(\GFM/n1156 ), .B(\GFM/n11550 ), .Z(\GFM/n1149 ) );
XOR2_X2 \GFM/U3298  ( .A(\GFM/n11580 ), .B(\GFM/n11570 ), .Z(\GFM/n11500 ));
XOR2_X2 \GFM/U3297  ( .A(z_in[64]), .B(\GFM/n1159 ), .Z(\GFM/n11510 ) );
XOR2_X2 \GFM/U3296  ( .A(\GFM/N2011 ), .B(\GFM/N2012 ), .Z(\GFM/n1152 ) );
XOR2_X2 \GFM/U3295  ( .A(\GFM/N2008 ), .B(\GFM/N2009 ), .Z(\GFM/n1153 ) );
XOR2_X2 \GFM/U3294  ( .A(\GFM/N2004 ), .B(\GFM/N2005 ), .Z(\GFM/n11540 ) );
XOR2_X2 \GFM/U3293  ( .A(\GFM/N2000 ), .B(\GFM/N2002 ), .Z(\GFM/n11550 ) );
XOR2_X2 \GFM/U3292  ( .A(\GFM/N1995 ), .B(\GFM/N1999 ), .Z(\GFM/n1156 ) );
XOR2_X2 \GFM/U3291  ( .A(\GFM/N1992 ), .B(\GFM/N1994 ), .Z(\GFM/n11570 ) );
XOR2_X2 \GFM/U3290  ( .A(\GFM/N1988 ), .B(\GFM/N1991 ), .Z(\GFM/n11580 ) );
XOR2_X2 \GFM/U3289  ( .A(\GFM/N1985 ), .B(\GFM/N1987 ), .Z(\GFM/n1159 ) );
XOR2_X2 \GFM/U3288  ( .A(\GFM/n1161 ), .B(\GFM/n1160 ), .Z(z_out[65]) );
XOR2_X2 \GFM/U3287  ( .A(\GFM/n11630 ), .B(\GFM/n11620 ), .Z(\GFM/n1160 ) );
XOR2_X2 \GFM/U3286  ( .A(\GFM/n11650 ), .B(\GFM/n1164 ), .Z(\GFM/n1161 ) );
XOR2_X2 \GFM/U3285  ( .A(\GFM/n11670 ), .B(\GFM/n1166 ), .Z(\GFM/n11620 ) );
XOR2_X2 \GFM/U3284  ( .A(\GFM/n1169 ), .B(\GFM/n11680 ), .Z(\GFM/n11630 ) );
XOR2_X2 \GFM/U3283  ( .A(\GFM/n11710 ), .B(\GFM/n1170 ), .Z(\GFM/n1164 ) );
XOR2_X2 \GFM/U3282  ( .A(\GFM/n1173 ), .B(\GFM/n11720 ), .Z(\GFM/n11650 ) );
XOR2_X2 \GFM/U3281  ( .A(z_in[65]), .B(\GFM/n11740 ), .Z(\GFM/n1166 ) );
XOR2_X2 \GFM/U3280  ( .A(\GFM/N2042 ), .B(\GFM/N2043 ), .Z(\GFM/n11670 ) );
XOR2_X2 \GFM/U3279  ( .A(\GFM/N2039 ), .B(\GFM/N2040 ), .Z(\GFM/n11680 ) );
XOR2_X2 \GFM/U3278  ( .A(\GFM/N2035 ), .B(\GFM/N2036 ), .Z(\GFM/n1169 ) );
XOR2_X2 \GFM/U3277  ( .A(\GFM/N2031 ), .B(\GFM/N2033 ), .Z(\GFM/n1170 ) );
XOR2_X2 \GFM/U3276  ( .A(\GFM/N2026 ), .B(\GFM/N2030 ), .Z(\GFM/n11710 ) );
XOR2_X2 \GFM/U3275  ( .A(\GFM/N2023 ), .B(\GFM/N2025 ), .Z(\GFM/n11720 ) );
XOR2_X2 \GFM/U3274  ( .A(\GFM/N2019 ), .B(\GFM/N2022 ), .Z(\GFM/n1173 ) );
XOR2_X2 \GFM/U3273  ( .A(\GFM/N2016 ), .B(\GFM/N2018 ), .Z(\GFM/n11740 ) );
XOR2_X2 \GFM/U3272  ( .A(\GFM/n1176 ), .B(\GFM/n11750 ), .Z(z_out[66]) );
XOR2_X2 \GFM/U3271  ( .A(\GFM/n1178 ), .B(\GFM/n1177 ), .Z(\GFM/n11750 ) );
XOR2_X2 \GFM/U3270  ( .A(\GFM/n1180 ), .B(\GFM/n11790 ), .Z(\GFM/n1176 ) );
XOR2_X2 \GFM/U3269  ( .A(\GFM/n11820 ), .B(\GFM/n11810 ), .Z(\GFM/n1177 ) );
XOR2_X2 \GFM/U3268  ( .A(\GFM/n1184 ), .B(\GFM/n1183 ), .Z(\GFM/n1178 ) );
XOR2_X2 \GFM/U3267  ( .A(\GFM/n11860 ), .B(\GFM/n11850 ), .Z(\GFM/n11790 ));
XOR2_X2 \GFM/U3266  ( .A(\GFM/n11880 ), .B(\GFM/n1187 ), .Z(\GFM/n1180 ) );
XOR2_X2 \GFM/U3265  ( .A(z_in[66]), .B(\GFM/n11890 ), .Z(\GFM/n11810 ) );
XOR2_X2 \GFM/U3264  ( .A(\GFM/N2073 ), .B(\GFM/N2074 ), .Z(\GFM/n11820 ) );
XOR2_X2 \GFM/U3263  ( .A(\GFM/N2070 ), .B(\GFM/N2071 ), .Z(\GFM/n1183 ) );
XOR2_X2 \GFM/U3262  ( .A(\GFM/N2066 ), .B(\GFM/N2067 ), .Z(\GFM/n1184 ) );
XOR2_X2 \GFM/U3261  ( .A(\GFM/N2062 ), .B(\GFM/N2064 ), .Z(\GFM/n11850 ) );
XOR2_X2 \GFM/U3260  ( .A(\GFM/N2057 ), .B(\GFM/N2061 ), .Z(\GFM/n11860 ) );
XOR2_X2 \GFM/U3259  ( .A(\GFM/N2054 ), .B(\GFM/N2056 ), .Z(\GFM/n1187 ) );
XOR2_X2 \GFM/U3258  ( .A(\GFM/N2050 ), .B(\GFM/N2053 ), .Z(\GFM/n11880 ) );
XOR2_X2 \GFM/U3257  ( .A(\GFM/N2047 ), .B(\GFM/N2049 ), .Z(\GFM/n11890 ) );
XOR2_X2 \GFM/U3256  ( .A(\GFM/n1191 ), .B(\GFM/n1190 ), .Z(z_out[67]) );
XOR2_X2 \GFM/U3255  ( .A(\GFM/n11930 ), .B(\GFM/n1192 ), .Z(\GFM/n1190 ) );
XOR2_X2 \GFM/U3254  ( .A(\GFM/n1195 ), .B(\GFM/n11940 ), .Z(\GFM/n1191 ) );
XOR2_X2 \GFM/U3253  ( .A(\GFM/n1197 ), .B(\GFM/n11960 ), .Z(\GFM/n1192 ) );
XOR2_X2 \GFM/U3252  ( .A(\GFM/n11990 ), .B(\GFM/n11980 ), .Z(\GFM/n11930 ));
XOR2_X2 \GFM/U3251  ( .A(\GFM/n1201 ), .B(\GFM/n1200 ), .Z(\GFM/n11940 ) );
XOR2_X2 \GFM/U3250  ( .A(\GFM/n12030 ), .B(\GFM/n12020 ), .Z(\GFM/n1195 ) );
XOR2_X2 \GFM/U3249  ( .A(z_in[67]), .B(\GFM/n1204 ), .Z(\GFM/n11960 ) );
XOR2_X2 \GFM/U3248  ( .A(\GFM/N2104 ), .B(\GFM/N2105 ), .Z(\GFM/n1197 ) );
XOR2_X2 \GFM/U3247  ( .A(\GFM/N2101 ), .B(\GFM/N2102 ), .Z(\GFM/n11980 ) );
XOR2_X2 \GFM/U3246  ( .A(\GFM/N2097 ), .B(\GFM/N2098 ), .Z(\GFM/n11990 ) );
XOR2_X2 \GFM/U3245  ( .A(\GFM/N2093 ), .B(\GFM/N2095 ), .Z(\GFM/n1200 ) );
XOR2_X2 \GFM/U3244  ( .A(\GFM/N2088 ), .B(\GFM/N2092 ), .Z(\GFM/n1201 ) );
XOR2_X2 \GFM/U3243  ( .A(\GFM/N2085 ), .B(\GFM/N2087 ), .Z(\GFM/n12020 ) );
XOR2_X2 \GFM/U3242  ( .A(\GFM/N2081 ), .B(\GFM/N2084 ), .Z(\GFM/n12030 ) );
XOR2_X2 \GFM/U3241  ( .A(\GFM/N2078 ), .B(\GFM/N2080 ), .Z(\GFM/n1204 ) );
XOR2_X2 \GFM/U3240  ( .A(\GFM/n12060 ), .B(\GFM/n12050 ), .Z(z_out[68]) );
XOR2_X2 \GFM/U3239  ( .A(\GFM/n1208 ), .B(\GFM/n1207 ), .Z(\GFM/n12050 ) );
XOR2_X2 \GFM/U3238  ( .A(\GFM/n12100 ), .B(\GFM/n1209 ), .Z(\GFM/n12060 ) );
XOR2_X2 \GFM/U3237  ( .A(\GFM/n12120 ), .B(\GFM/n1211 ), .Z(\GFM/n1207 ) );
XOR2_X2 \GFM/U3236  ( .A(\GFM/n1214 ), .B(\GFM/n12130 ), .Z(\GFM/n1208 ) );
XOR2_X2 \GFM/U3235  ( .A(\GFM/n12160 ), .B(\GFM/n1215 ), .Z(\GFM/n1209 ) );
XOR2_X2 \GFM/U3234  ( .A(\GFM/n1218 ), .B(\GFM/n12170 ), .Z(\GFM/n12100 ) );
XOR2_X2 \GFM/U3233  ( .A(z_in[68]), .B(\GFM/n12190 ), .Z(\GFM/n1211 ) );
XOR2_X2 \GFM/U3232  ( .A(\GFM/N2135 ), .B(\GFM/N2136 ), .Z(\GFM/n12120 ) );
XOR2_X2 \GFM/U3231  ( .A(\GFM/N2132 ), .B(\GFM/N2133 ), .Z(\GFM/n12130 ) );
XOR2_X2 \GFM/U3230  ( .A(\GFM/N2128 ), .B(\GFM/N2129 ), .Z(\GFM/n1214 ) );
XOR2_X2 \GFM/U3229  ( .A(\GFM/N2124 ), .B(\GFM/N2126 ), .Z(\GFM/n1215 ) );
XOR2_X2 \GFM/U3228  ( .A(\GFM/N2119 ), .B(\GFM/N2123 ), .Z(\GFM/n12160 ) );
XOR2_X2 \GFM/U3227  ( .A(\GFM/N2116 ), .B(\GFM/N2118 ), .Z(\GFM/n12170 ) );
XOR2_X2 \GFM/U3226  ( .A(\GFM/N2112 ), .B(\GFM/N2115 ), .Z(\GFM/n1218 ) );
XOR2_X2 \GFM/U3225  ( .A(\GFM/N2109 ), .B(\GFM/N2111 ), .Z(\GFM/n12190 ) );
XOR2_X2 \GFM/U3224  ( .A(\GFM/n1221 ), .B(\GFM/n12200 ), .Z(z_out[69]) );
XOR2_X2 \GFM/U3223  ( .A(\GFM/n1223 ), .B(\GFM/n1222 ), .Z(\GFM/n12200 ) );
XOR2_X2 \GFM/U3222  ( .A(\GFM/n12250 ), .B(\GFM/n12240 ), .Z(\GFM/n1221 ) );
XOR2_X2 \GFM/U3221  ( .A(\GFM/n12270 ), .B(\GFM/n1226 ), .Z(\GFM/n1222 ) );
XOR2_X2 \GFM/U3220  ( .A(\GFM/n12290 ), .B(\GFM/n1228 ), .Z(\GFM/n1223 ) );
XOR2_X2 \GFM/U3219  ( .A(\GFM/n1231 ), .B(\GFM/n12300 ), .Z(\GFM/n12240 ) );
XOR2_X2 \GFM/U3218  ( .A(\GFM/n12330 ), .B(\GFM/n1232 ), .Z(\GFM/n12250 ) );
XOR2_X2 \GFM/U3217  ( .A(z_in[69]), .B(\GFM/n12340 ), .Z(\GFM/n1226 ) );
XOR2_X2 \GFM/U3216  ( .A(\GFM/N2166 ), .B(\GFM/N2167 ), .Z(\GFM/n12270 ) );
XOR2_X2 \GFM/U3215  ( .A(\GFM/N2163 ), .B(\GFM/N2164 ), .Z(\GFM/n1228 ) );
XOR2_X2 \GFM/U3214  ( .A(\GFM/N2159 ), .B(\GFM/N2160 ), .Z(\GFM/n12290 ) );
XOR2_X2 \GFM/U3213  ( .A(\GFM/N2155 ), .B(\GFM/N2157 ), .Z(\GFM/n12300 ) );
XOR2_X2 \GFM/U3212  ( .A(\GFM/N2150 ), .B(\GFM/N2154 ), .Z(\GFM/n1231 ) );
XOR2_X2 \GFM/U3211  ( .A(\GFM/N2147 ), .B(\GFM/N2149 ), .Z(\GFM/n1232 ) );
XOR2_X2 \GFM/U3210  ( .A(\GFM/N2143 ), .B(\GFM/N2146 ), .Z(\GFM/n12330 ) );
XOR2_X2 \GFM/U3209  ( .A(\GFM/N2140 ), .B(\GFM/N2142 ), .Z(\GFM/n12340 ) );
XOR2_X2 \GFM/U3208  ( .A(\GFM/n12360 ), .B(\GFM/n1235 ), .Z(z_out[70]) );
XOR2_X2 \GFM/U3207  ( .A(\GFM/n1238 ), .B(\GFM/n12370 ), .Z(\GFM/n1235 ) );
XOR2_X2 \GFM/U3206  ( .A(\GFM/n1240 ), .B(\GFM/n1239 ), .Z(\GFM/n12360 ) );
XOR2_X2 \GFM/U3205  ( .A(\GFM/n1242 ), .B(\GFM/n12410 ), .Z(\GFM/n12370 ) );
XOR2_X2 \GFM/U3204  ( .A(\GFM/n12440 ), .B(\GFM/n12430 ), .Z(\GFM/n1238 ) );
XOR2_X2 \GFM/U3203  ( .A(\GFM/n1246 ), .B(\GFM/n1245 ), .Z(\GFM/n1239 ) );
XOR2_X2 \GFM/U3202  ( .A(\GFM/n12480 ), .B(\GFM/n12470 ), .Z(\GFM/n1240 ) );
XOR2_X2 \GFM/U3201  ( .A(z_in[70]), .B(\GFM/n1249 ), .Z(\GFM/n12410 ) );
XOR2_X2 \GFM/U3200  ( .A(\GFM/N2197 ), .B(\GFM/N2198 ), .Z(\GFM/n1242 ) );
XOR2_X2 \GFM/U3199  ( .A(\GFM/N2194 ), .B(\GFM/N2195 ), .Z(\GFM/n12430 ) );
XOR2_X2 \GFM/U3198  ( .A(\GFM/N2190 ), .B(\GFM/N2191 ), .Z(\GFM/n12440 ) );
XOR2_X2 \GFM/U3197  ( .A(\GFM/N2186 ), .B(\GFM/N2188 ), .Z(\GFM/n1245 ) );
XOR2_X2 \GFM/U3196  ( .A(\GFM/N2181 ), .B(\GFM/N2185 ), .Z(\GFM/n1246 ) );
XOR2_X2 \GFM/U3195  ( .A(\GFM/N2178 ), .B(\GFM/N2180 ), .Z(\GFM/n12470 ) );
XOR2_X2 \GFM/U3194  ( .A(\GFM/N2174 ), .B(\GFM/N2177 ), .Z(\GFM/n12480 ) );
XOR2_X2 \GFM/U3193  ( .A(\GFM/N2171 ), .B(\GFM/N2173 ), .Z(\GFM/n1249 ) );
XOR2_X2 \GFM/U3192  ( .A(\GFM/n12510 ), .B(\GFM/n12500 ), .Z(z_out[71]) );
XOR2_X2 \GFM/U3191  ( .A(\GFM/n1253 ), .B(\GFM/n1252 ), .Z(\GFM/n12500 ) );
XOR2_X2 \GFM/U3190  ( .A(\GFM/n12550 ), .B(\GFM/n1254 ), .Z(\GFM/n12510 ) );
XOR2_X2 \GFM/U3189  ( .A(\GFM/n1257 ), .B(\GFM/n12560 ), .Z(\GFM/n1252 ) );
XOR2_X2 \GFM/U3188  ( .A(\GFM/n1259 ), .B(\GFM/n12580 ), .Z(\GFM/n1253 ) );
XOR2_X2 \GFM/U3187  ( .A(\GFM/n12610 ), .B(\GFM/n12600 ), .Z(\GFM/n1254 ) );
XOR2_X2 \GFM/U3186  ( .A(\GFM/n1263 ), .B(\GFM/n1262 ), .Z(\GFM/n12550 ) );
XOR2_X2 \GFM/U3185  ( .A(z_in[71]), .B(\GFM/n12640 ), .Z(\GFM/n12560 ) );
XOR2_X2 \GFM/U3184  ( .A(\GFM/N2228 ), .B(\GFM/N2229 ), .Z(\GFM/n1257 ) );
XOR2_X2 \GFM/U3183  ( .A(\GFM/N2225 ), .B(\GFM/N2226 ), .Z(\GFM/n12580 ) );
XOR2_X2 \GFM/U3182  ( .A(\GFM/N2221 ), .B(\GFM/N2222 ), .Z(\GFM/n1259 ) );
XOR2_X2 \GFM/U3181  ( .A(\GFM/N2217 ), .B(\GFM/N2219 ), .Z(\GFM/n12600 ) );
XOR2_X2 \GFM/U3180  ( .A(\GFM/N2212 ), .B(\GFM/N2216 ), .Z(\GFM/n12610 ) );
XOR2_X2 \GFM/U3179  ( .A(\GFM/N2209 ), .B(\GFM/N2211 ), .Z(\GFM/n1262 ) );
XOR2_X2 \GFM/U3178  ( .A(\GFM/N2205 ), .B(\GFM/N2208 ), .Z(\GFM/n1263 ) );
XOR2_X2 \GFM/U3177  ( .A(\GFM/N2202 ), .B(\GFM/N2204 ), .Z(\GFM/n12640 ) );
XOR2_X2 \GFM/U3176  ( .A(\GFM/n1266 ), .B(\GFM/n12650 ), .Z(z_out[72]) );
XOR2_X2 \GFM/U3175  ( .A(\GFM/n12680 ), .B(\GFM/n12670 ), .Z(\GFM/n12650 ));
XOR2_X2 \GFM/U3174  ( .A(\GFM/n1270 ), .B(\GFM/n1269 ), .Z(\GFM/n1266 ) );
XOR2_X2 \GFM/U3173  ( .A(\GFM/n12720 ), .B(\GFM/n1271 ), .Z(\GFM/n12670 ) );
XOR2_X2 \GFM/U3172  ( .A(\GFM/n12740 ), .B(\GFM/n1273 ), .Z(\GFM/n12680 ) );
XOR2_X2 \GFM/U3171  ( .A(\GFM/n1276 ), .B(\GFM/n12750 ), .Z(\GFM/n1269 ) );
XOR2_X2 \GFM/U3170  ( .A(\GFM/n12780 ), .B(\GFM/n1277 ), .Z(\GFM/n1270 ) );
XOR2_X2 \GFM/U3169  ( .A(z_in[72]), .B(\GFM/n12790 ), .Z(\GFM/n1271 ) );
XOR2_X2 \GFM/U3168  ( .A(\GFM/N2259 ), .B(\GFM/N2260 ), .Z(\GFM/n12720 ) );
XOR2_X2 \GFM/U3167  ( .A(\GFM/N2256 ), .B(\GFM/N2257 ), .Z(\GFM/n1273 ) );
XOR2_X2 \GFM/U3166  ( .A(\GFM/N2252 ), .B(\GFM/N2253 ), .Z(\GFM/n12740 ) );
XOR2_X2 \GFM/U3165  ( .A(\GFM/N2248 ), .B(\GFM/N2250 ), .Z(\GFM/n12750 ) );
XOR2_X2 \GFM/U3164  ( .A(\GFM/N2243 ), .B(\GFM/N2247 ), .Z(\GFM/n1276 ) );
XOR2_X2 \GFM/U3163  ( .A(\GFM/N2240 ), .B(\GFM/N2242 ), .Z(\GFM/n1277 ) );
XOR2_X2 \GFM/U3162  ( .A(\GFM/N2236 ), .B(\GFM/N2239 ), .Z(\GFM/n12780 ) );
XOR2_X2 \GFM/U3161  ( .A(\GFM/N2233 ), .B(\GFM/N2235 ), .Z(\GFM/n12790 ) );
XOR2_X2 \GFM/U3160  ( .A(\GFM/n12810 ), .B(\GFM/n1280 ), .Z(z_out[73]) );
XOR2_X2 \GFM/U3159  ( .A(\GFM/n1283 ), .B(\GFM/n12820 ), .Z(\GFM/n1280 ) );
XOR2_X2 \GFM/U3158  ( .A(\GFM/n1285 ), .B(\GFM/n1284 ), .Z(\GFM/n12810 ) );
XOR2_X2 \GFM/U3157  ( .A(\GFM/n12870 ), .B(\GFM/n12860 ), .Z(\GFM/n12820 ));
XOR2_X2 \GFM/U3156  ( .A(\GFM/n12890 ), .B(\GFM/n1288 ), .Z(\GFM/n1283 ) );
XOR2_X2 \GFM/U3155  ( .A(\GFM/n12910 ), .B(\GFM/n1290 ), .Z(\GFM/n1284 ) );
XOR2_X2 \GFM/U3154  ( .A(\GFM/n1293 ), .B(\GFM/n12920 ), .Z(\GFM/n1285 ) );
XOR2_X2 \GFM/U3153  ( .A(z_in[73]), .B(\GFM/n1294 ), .Z(\GFM/n12860 ) );
XOR2_X2 \GFM/U3152  ( .A(\GFM/N2290 ), .B(\GFM/N2291 ), .Z(\GFM/n12870 ) );
XOR2_X2 \GFM/U3151  ( .A(\GFM/N2287 ), .B(\GFM/N2288 ), .Z(\GFM/n1288 ) );
XOR2_X2 \GFM/U3150  ( .A(\GFM/N2283 ), .B(\GFM/N2284 ), .Z(\GFM/n12890 ) );
XOR2_X2 \GFM/U3149  ( .A(\GFM/N2279 ), .B(\GFM/N2281 ), .Z(\GFM/n1290 ) );
XOR2_X2 \GFM/U3148  ( .A(\GFM/N2274 ), .B(\GFM/N2278 ), .Z(\GFM/n12910 ) );
XOR2_X2 \GFM/U3147  ( .A(\GFM/N2271 ), .B(\GFM/N2273 ), .Z(\GFM/n12920 ) );
XOR2_X2 \GFM/U3146  ( .A(\GFM/N2267 ), .B(\GFM/N2270 ), .Z(\GFM/n1293 ) );
XOR2_X2 \GFM/U3145  ( .A(\GFM/N2264 ), .B(\GFM/N2266 ), .Z(\GFM/n1294 ) );
XOR2_X2 \GFM/U3144  ( .A(\GFM/n12960 ), .B(\GFM/n12950 ), .Z(z_out[74]) );
XOR2_X2 \GFM/U3143  ( .A(\GFM/n12980 ), .B(\GFM/n1297 ), .Z(\GFM/n12950 ) );
XOR2_X2 \GFM/U3142  ( .A(\GFM/n1300 ), .B(\GFM/n12990 ), .Z(\GFM/n12960 ) );
XOR2_X2 \GFM/U3141  ( .A(\GFM/n1302 ), .B(\GFM/n1301 ), .Z(\GFM/n1297 ) );
XOR2_X2 \GFM/U3140  ( .A(\GFM/n1304 ), .B(\GFM/n13030 ), .Z(\GFM/n12980 ) );
XOR2_X2 \GFM/U3139  ( .A(\GFM/n13060 ), .B(\GFM/n13050 ), .Z(\GFM/n12990 ));
XOR2_X2 \GFM/U3138  ( .A(\GFM/n1308 ), .B(\GFM/n1307 ), .Z(\GFM/n1300 ) );
XOR2_X2 \GFM/U3137  ( .A(z_in[74]), .B(\GFM/n13090 ), .Z(\GFM/n1301 ) );
XOR2_X2 \GFM/U3136  ( .A(\GFM/N2321 ), .B(\GFM/N2322 ), .Z(\GFM/n1302 ) );
XOR2_X2 \GFM/U3135  ( .A(\GFM/N2318 ), .B(\GFM/N2319 ), .Z(\GFM/n13030 ) );
XOR2_X2 \GFM/U3134  ( .A(\GFM/N2314 ), .B(\GFM/N2315 ), .Z(\GFM/n1304 ) );
XOR2_X2 \GFM/U3133  ( .A(\GFM/N2310 ), .B(\GFM/N2312 ), .Z(\GFM/n13050 ) );
XOR2_X2 \GFM/U3132  ( .A(\GFM/N2305 ), .B(\GFM/N2309 ), .Z(\GFM/n13060 ) );
XOR2_X2 \GFM/U3131  ( .A(\GFM/N2302 ), .B(\GFM/N2304 ), .Z(\GFM/n1307 ) );
XOR2_X2 \GFM/U3130  ( .A(\GFM/N2298 ), .B(\GFM/N2301 ), .Z(\GFM/n1308 ) );
XOR2_X2 \GFM/U3129  ( .A(\GFM/N2295 ), .B(\GFM/N2297 ), .Z(\GFM/n13090 ) );
XOR2_X2 \GFM/U3128  ( .A(\GFM/n1311 ), .B(\GFM/n13100 ), .Z(z_out[75]) );
XOR2_X2 \GFM/U3127  ( .A(\GFM/n13130 ), .B(\GFM/n13120 ), .Z(\GFM/n13100 ));
XOR2_X2 \GFM/U3126  ( .A(\GFM/n1315 ), .B(\GFM/n1314 ), .Z(\GFM/n1311 ) );
XOR2_X2 \GFM/U3125  ( .A(\GFM/n13170 ), .B(\GFM/n1316 ), .Z(\GFM/n13120 ) );
XOR2_X2 \GFM/U3124  ( .A(\GFM/n1319 ), .B(\GFM/n13180 ), .Z(\GFM/n13130 ) );
XOR2_X2 \GFM/U3123  ( .A(\GFM/n1321 ), .B(\GFM/n13200 ), .Z(\GFM/n1314 ) );
XOR2_X2 \GFM/U3122  ( .A(\GFM/n13230 ), .B(\GFM/n13220 ), .Z(\GFM/n1315 ) );
XOR2_X2 \GFM/U3121  ( .A(z_in[75]), .B(\GFM/n1324 ), .Z(\GFM/n1316 ) );
XOR2_X2 \GFM/U3120  ( .A(\GFM/N2352 ), .B(\GFM/N2353 ), .Z(\GFM/n13170 ) );
XOR2_X2 \GFM/U3119  ( .A(\GFM/N2349 ), .B(\GFM/N2350 ), .Z(\GFM/n13180 ) );
XOR2_X2 \GFM/U3118  ( .A(\GFM/N2345 ), .B(\GFM/N2346 ), .Z(\GFM/n1319 ) );
XOR2_X2 \GFM/U3117  ( .A(\GFM/N2341 ), .B(\GFM/N2343 ), .Z(\GFM/n13200 ) );
XOR2_X2 \GFM/U3116  ( .A(\GFM/N2336 ), .B(\GFM/N2340 ), .Z(\GFM/n1321 ) );
XOR2_X2 \GFM/U3115  ( .A(\GFM/N2333 ), .B(\GFM/N2335 ), .Z(\GFM/n13220 ) );
XOR2_X2 \GFM/U3114  ( .A(\GFM/N2329 ), .B(\GFM/N2332 ), .Z(\GFM/n13230 ) );
XOR2_X2 \GFM/U3113  ( .A(\GFM/N2326 ), .B(\GFM/N2328 ), .Z(\GFM/n1324 ) );
XOR2_X2 \GFM/U3112  ( .A(\GFM/n13260 ), .B(\GFM/n1325 ), .Z(z_out[76]) );
XOR2_X2 \GFM/U3111  ( .A(\GFM/n1328 ), .B(\GFM/n13270 ), .Z(\GFM/n1325 ) );
XOR2_X2 \GFM/U3110  ( .A(\GFM/n13300 ), .B(\GFM/n13290 ), .Z(\GFM/n13260 ));
XOR2_X2 \GFM/U3109  ( .A(\GFM/n1332 ), .B(\GFM/n1331 ), .Z(\GFM/n13270 ) );
XOR2_X2 \GFM/U3108  ( .A(\GFM/n13340 ), .B(\GFM/n1333 ), .Z(\GFM/n1328 ) );
XOR2_X2 \GFM/U3107  ( .A(\GFM/n13360 ), .B(\GFM/n1335 ), .Z(\GFM/n13290 ) );
XOR2_X2 \GFM/U3106  ( .A(\GFM/n1338 ), .B(\GFM/n13370 ), .Z(\GFM/n13300 ) );
XOR2_X2 \GFM/U3105  ( .A(z_in[76]), .B(\GFM/n1339 ), .Z(\GFM/n1331 ) );
XOR2_X2 \GFM/U3104  ( .A(\GFM/N2383 ), .B(\GFM/N2384 ), .Z(\GFM/n1332 ) );
XOR2_X2 \GFM/U3103  ( .A(\GFM/N2380 ), .B(\GFM/N2381 ), .Z(\GFM/n1333 ) );
XOR2_X2 \GFM/U3102  ( .A(\GFM/N2376 ), .B(\GFM/N2377 ), .Z(\GFM/n13340 ) );
XOR2_X2 \GFM/U3101  ( .A(\GFM/N2372 ), .B(\GFM/N2374 ), .Z(\GFM/n1335 ) );
XOR2_X2 \GFM/U3100  ( .A(\GFM/N2367 ), .B(\GFM/N2371 ), .Z(\GFM/n13360 ) );
XOR2_X2 \GFM/U3099  ( .A(\GFM/N2364 ), .B(\GFM/N2366 ), .Z(\GFM/n13370 ) );
XOR2_X2 \GFM/U3098  ( .A(\GFM/N2360 ), .B(\GFM/N2363 ), .Z(\GFM/n1338 ) );
XOR2_X2 \GFM/U3097  ( .A(\GFM/N2357 ), .B(\GFM/N2359 ), .Z(\GFM/n1339 ) );
XOR2_X2 \GFM/U3096  ( .A(\GFM/n13410 ), .B(\GFM/n13400 ), .Z(z_out[77]) );
XOR2_X2 \GFM/U3095  ( .A(\GFM/n13430 ), .B(\GFM/n1342 ), .Z(\GFM/n13400 ) );
XOR2_X2 \GFM/U3094  ( .A(\GFM/n1345 ), .B(\GFM/n13440 ), .Z(\GFM/n13410 ) );
XOR2_X2 \GFM/U3093  ( .A(\GFM/n1347 ), .B(\GFM/n1346 ), .Z(\GFM/n1342 ) );
XOR2_X2 \GFM/U3092  ( .A(\GFM/n13490 ), .B(\GFM/n13480 ), .Z(\GFM/n13430 ));
XOR2_X2 \GFM/U3091  ( .A(\GFM/n13510 ), .B(\GFM/n1350 ), .Z(\GFM/n13440 ) );
XOR2_X2 \GFM/U3090  ( .A(\GFM/n13530 ), .B(\GFM/n1352 ), .Z(\GFM/n1345 ) );
XOR2_X2 \GFM/U3089  ( .A(z_in[77]), .B(\GFM/n13540 ), .Z(\GFM/n1346 ) );
XOR2_X2 \GFM/U3088  ( .A(\GFM/N2414 ), .B(\GFM/N2415 ), .Z(\GFM/n1347 ) );
XOR2_X2 \GFM/U3087  ( .A(\GFM/N2411 ), .B(\GFM/N2412 ), .Z(\GFM/n13480 ) );
XOR2_X2 \GFM/U3086  ( .A(\GFM/N2407 ), .B(\GFM/N2408 ), .Z(\GFM/n13490 ) );
XOR2_X2 \GFM/U3085  ( .A(\GFM/N2403 ), .B(\GFM/N2405 ), .Z(\GFM/n1350 ) );
XOR2_X2 \GFM/U3084  ( .A(\GFM/N2398 ), .B(\GFM/N2402 ), .Z(\GFM/n13510 ) );
XOR2_X2 \GFM/U3083  ( .A(\GFM/N2395 ), .B(\GFM/N2397 ), .Z(\GFM/n1352 ) );
XOR2_X2 \GFM/U3082  ( .A(\GFM/N2391 ), .B(\GFM/N2394 ), .Z(\GFM/n13530 ) );
XOR2_X2 \GFM/U3081  ( .A(\GFM/N2388 ), .B(\GFM/N2390 ), .Z(\GFM/n13540 ) );
XOR2_X2 \GFM/U3080  ( .A(\GFM/n1356 ), .B(\GFM/n1355 ), .Z(z_out[78]) );
XOR2_X2 \GFM/U3079  ( .A(\GFM/n13580 ), .B(\GFM/n13570 ), .Z(\GFM/n1355 ) );
XOR2_X2 \GFM/U3078  ( .A(\GFM/n13600 ), .B(\GFM/n1359 ), .Z(\GFM/n1356 ) );
XOR2_X2 \GFM/U3077  ( .A(\GFM/n1362 ), .B(\GFM/n13610 ), .Z(\GFM/n13570 ) );
XOR2_X2 \GFM/U3076  ( .A(\GFM/n1364 ), .B(\GFM/n1363 ), .Z(\GFM/n13580 ) );
XOR2_X2 \GFM/U3075  ( .A(\GFM/n1366 ), .B(\GFM/n13650 ), .Z(\GFM/n1359 ) );
XOR2_X2 \GFM/U3074  ( .A(\GFM/n13680 ), .B(\GFM/n13670 ), .Z(\GFM/n13600 ));
XOR2_X2 \GFM/U3073  ( .A(z_in[78]), .B(\GFM/n1369 ), .Z(\GFM/n13610 ) );
XOR2_X2 \GFM/U3072  ( .A(\GFM/N2445 ), .B(\GFM/N2446 ), .Z(\GFM/n1362 ) );
XOR2_X2 \GFM/U3071  ( .A(\GFM/N2442 ), .B(\GFM/N2443 ), .Z(\GFM/n1363 ) );
XOR2_X2 \GFM/U3070  ( .A(\GFM/N2438 ), .B(\GFM/N2439 ), .Z(\GFM/n1364 ) );
XOR2_X2 \GFM/U3069  ( .A(\GFM/N2434 ), .B(\GFM/N2436 ), .Z(\GFM/n13650 ) );
XOR2_X2 \GFM/U3068  ( .A(\GFM/N2429 ), .B(\GFM/N2433 ), .Z(\GFM/n1366 ) );
XOR2_X2 \GFM/U3067  ( .A(\GFM/N2426 ), .B(\GFM/N2428 ), .Z(\GFM/n13670 ) );
XOR2_X2 \GFM/U3066  ( .A(\GFM/N2422 ), .B(\GFM/N2425 ), .Z(\GFM/n13680 ) );
XOR2_X2 \GFM/U3065  ( .A(\GFM/N2419 ), .B(\GFM/N2421 ), .Z(\GFM/n1369 ) );
XOR2_X2 \GFM/U3064  ( .A(\GFM/n13710 ), .B(\GFM/n1370 ), .Z(z_out[79]) );
XOR2_X2 \GFM/U3063  ( .A(\GFM/n1373 ), .B(\GFM/n13720 ), .Z(\GFM/n1370 ) );
XOR2_X2 \GFM/U3062  ( .A(\GFM/n13750 ), .B(\GFM/n13740 ), .Z(\GFM/n13710 ));
XOR2_X2 \GFM/U3061  ( .A(\GFM/n1377 ), .B(\GFM/n1376 ), .Z(\GFM/n13720 ) );
XOR2_X2 \GFM/U3060  ( .A(\GFM/n13790 ), .B(\GFM/n1378 ), .Z(\GFM/n1373 ) );
XOR2_X2 \GFM/U3059  ( .A(\GFM/n1381 ), .B(\GFM/n13800 ), .Z(\GFM/n13740 ) );
XOR2_X2 \GFM/U3058  ( .A(\GFM/n1383 ), .B(\GFM/n13820 ), .Z(\GFM/n13750 ) );
XOR2_X2 \GFM/U3057  ( .A(z_in[79]), .B(\GFM/n13840 ), .Z(\GFM/n1376 ) );
XOR2_X2 \GFM/U3056  ( .A(\GFM/N2476 ), .B(\GFM/N2477 ), .Z(\GFM/n1377 ) );
XOR2_X2 \GFM/U3055  ( .A(\GFM/N2473 ), .B(\GFM/N2474 ), .Z(\GFM/n1378 ) );
XOR2_X2 \GFM/U3054  ( .A(\GFM/N2469 ), .B(\GFM/N2470 ), .Z(\GFM/n13790 ) );
XOR2_X2 \GFM/U3053  ( .A(\GFM/N2465 ), .B(\GFM/N2467 ), .Z(\GFM/n13800 ) );
XOR2_X2 \GFM/U3052  ( .A(\GFM/N2460 ), .B(\GFM/N2464 ), .Z(\GFM/n1381 ) );
XOR2_X2 \GFM/U3051  ( .A(\GFM/N2457 ), .B(\GFM/N2459 ), .Z(\GFM/n13820 ) );
XOR2_X2 \GFM/U3050  ( .A(\GFM/N2453 ), .B(\GFM/N2456 ), .Z(\GFM/n1383 ) );
XOR2_X2 \GFM/U3049  ( .A(\GFM/N2450 ), .B(\GFM/N2452 ), .Z(\GFM/n13840 ) );
XOR2_X2 \GFM/U3048  ( .A(\GFM/n1386 ), .B(\GFM/n13850 ), .Z(z_out[80]) );
XOR2_X2 \GFM/U3047  ( .A(\GFM/n13880 ), .B(\GFM/n1387 ), .Z(\GFM/n13850 ) );
XOR2_X2 \GFM/U3046  ( .A(\GFM/n1390 ), .B(\GFM/n13890 ), .Z(\GFM/n1386 ) );
XOR2_X2 \GFM/U3045  ( .A(\GFM/n13920 ), .B(\GFM/n13910 ), .Z(\GFM/n1387 ) );
XOR2_X2 \GFM/U3044  ( .A(\GFM/n1394 ), .B(\GFM/n1393 ), .Z(\GFM/n13880 ) );
XOR2_X2 \GFM/U3043  ( .A(\GFM/n13960 ), .B(\GFM/n1395 ), .Z(\GFM/n13890 ) );
XOR2_X2 \GFM/U3042  ( .A(\GFM/n13980 ), .B(\GFM/n1397 ), .Z(\GFM/n1390 ) );
XOR2_X2 \GFM/U3041  ( .A(z_in[80]), .B(\GFM/n13990 ), .Z(\GFM/n13910 ) );
XOR2_X2 \GFM/U3040  ( .A(\GFM/N2507 ), .B(\GFM/N2508 ), .Z(\GFM/n13920 ) );
XOR2_X2 \GFM/U3039  ( .A(\GFM/N2504 ), .B(\GFM/N2505 ), .Z(\GFM/n1393 ) );
XOR2_X2 \GFM/U3038  ( .A(\GFM/N2500 ), .B(\GFM/N2501 ), .Z(\GFM/n1394 ) );
XOR2_X2 \GFM/U3037  ( .A(\GFM/N2496 ), .B(\GFM/N2498 ), .Z(\GFM/n1395 ) );
XOR2_X2 \GFM/U3036  ( .A(\GFM/N2491 ), .B(\GFM/N2495 ), .Z(\GFM/n13960 ) );
XOR2_X2 \GFM/U3035  ( .A(\GFM/N2488 ), .B(\GFM/N2490 ), .Z(\GFM/n1397 ) );
XOR2_X2 \GFM/U3034  ( .A(\GFM/N2484 ), .B(\GFM/N2487 ), .Z(\GFM/n13980 ) );
XOR2_X2 \GFM/U3033  ( .A(\GFM/N2481 ), .B(\GFM/N2483 ), .Z(\GFM/n13990 ) );
XOR2_X2 \GFM/U3032  ( .A(\GFM/n1401 ), .B(\GFM/n1400 ), .Z(z_out[81]) );
XOR2_X2 \GFM/U3031  ( .A(\GFM/n14030 ), .B(\GFM/n14020 ), .Z(\GFM/n1400 ) );
XOR2_X2 \GFM/U3030  ( .A(\GFM/n14050 ), .B(\GFM/n1404 ), .Z(\GFM/n1401 ) );
XOR2_X2 \GFM/U3029  ( .A(\GFM/n1407 ), .B(\GFM/n14060 ), .Z(\GFM/n14020 ) );
XOR2_X2 \GFM/U3028  ( .A(\GFM/n1409 ), .B(\GFM/n1408 ), .Z(\GFM/n14030 ) );
XOR2_X2 \GFM/U3027  ( .A(\GFM/n14110 ), .B(\GFM/n14100 ), .Z(\GFM/n1404 ) );
XOR2_X2 \GFM/U3026  ( .A(\GFM/n14130 ), .B(\GFM/n1412 ), .Z(\GFM/n14050 ) );
XOR2_X2 \GFM/U3025  ( .A(z_in[81]), .B(\GFM/n1414 ), .Z(\GFM/n14060 ) );
XOR2_X2 \GFM/U3024  ( .A(\GFM/N2538 ), .B(\GFM/N2539 ), .Z(\GFM/n1407 ) );
XOR2_X2 \GFM/U3023  ( .A(\GFM/N2535 ), .B(\GFM/N2536 ), .Z(\GFM/n1408 ) );
XOR2_X2 \GFM/U3022  ( .A(\GFM/N2531 ), .B(\GFM/N2532 ), .Z(\GFM/n1409 ) );
XOR2_X2 \GFM/U3021  ( .A(\GFM/N2527 ), .B(\GFM/N2529 ), .Z(\GFM/n14100 ) );
XOR2_X2 \GFM/U3020  ( .A(\GFM/N2522 ), .B(\GFM/N2526 ), .Z(\GFM/n14110 ) );
XOR2_X2 \GFM/U3019  ( .A(\GFM/N2519 ), .B(\GFM/N2521 ), .Z(\GFM/n1412 ) );
XOR2_X2 \GFM/U3018  ( .A(\GFM/N2515 ), .B(\GFM/N2518 ), .Z(\GFM/n14130 ) );
XOR2_X2 \GFM/U3017  ( .A(\GFM/N2512 ), .B(\GFM/N2514 ), .Z(\GFM/n1414 ) );
XOR2_X2 \GFM/U3016  ( .A(\GFM/n14160 ), .B(\GFM/n14150 ), .Z(z_out[82]) );
XOR2_X2 \GFM/U3015  ( .A(\GFM/n1418 ), .B(\GFM/n1417 ), .Z(\GFM/n14150 ) );
XOR2_X2 \GFM/U3014  ( .A(\GFM/n14200 ), .B(\GFM/n14190 ), .Z(\GFM/n14160 ));
XOR2_X2 \GFM/U3013  ( .A(\GFM/n14220 ), .B(\GFM/n1421 ), .Z(\GFM/n1417 ) );
XOR2_X2 \GFM/U3012  ( .A(\GFM/n1424 ), .B(\GFM/n14230 ), .Z(\GFM/n1418 ) );
XOR2_X2 \GFM/U3011  ( .A(\GFM/n1426 ), .B(\GFM/n1425 ), .Z(\GFM/n14190 ) );
XOR2_X2 \GFM/U3010  ( .A(\GFM/n1428 ), .B(\GFM/n14270 ), .Z(\GFM/n14200 ) );
XOR2_X2 \GFM/U3009  ( .A(z_in[82]), .B(\GFM/n14290 ), .Z(\GFM/n1421 ) );
XOR2_X2 \GFM/U3008  ( .A(\GFM/N2569 ), .B(\GFM/N2570 ), .Z(\GFM/n14220 ) );
XOR2_X2 \GFM/U3007  ( .A(\GFM/N2566 ), .B(\GFM/N2567 ), .Z(\GFM/n14230 ) );
XOR2_X2 \GFM/U3006  ( .A(\GFM/N2562 ), .B(\GFM/N2563 ), .Z(\GFM/n1424 ) );
XOR2_X2 \GFM/U3005  ( .A(\GFM/N2558 ), .B(\GFM/N2560 ), .Z(\GFM/n1425 ) );
XOR2_X2 \GFM/U3004  ( .A(\GFM/N2553 ), .B(\GFM/N2557 ), .Z(\GFM/n1426 ) );
XOR2_X2 \GFM/U3003  ( .A(\GFM/N2550 ), .B(\GFM/N2552 ), .Z(\GFM/n14270 ) );
XOR2_X2 \GFM/U3002  ( .A(\GFM/N2546 ), .B(\GFM/N2549 ), .Z(\GFM/n1428 ) );
XOR2_X2 \GFM/U3001  ( .A(\GFM/N2543 ), .B(\GFM/N2545 ), .Z(\GFM/n14290 ) );
XOR2_X2 \GFM/U3000  ( .A(\GFM/n1431 ), .B(\GFM/n14300 ), .Z(z_out[83]) );
XOR2_X2 \GFM/U2999  ( .A(\GFM/n14330 ), .B(\GFM/n1432 ), .Z(\GFM/n14300 ) );
XOR2_X2 \GFM/U2998  ( .A(\GFM/n1435 ), .B(\GFM/n14340 ), .Z(\GFM/n1431 ) );
XOR2_X2 \GFM/U2997  ( .A(\GFM/n14370 ), .B(\GFM/n14360 ), .Z(\GFM/n1432 ) );
XOR2_X2 \GFM/U2996  ( .A(\GFM/n1439 ), .B(\GFM/n1438 ), .Z(\GFM/n14330 ) );
XOR2_X2 \GFM/U2995  ( .A(\GFM/n14410 ), .B(\GFM/n1440 ), .Z(\GFM/n14340 ) );
XOR2_X2 \GFM/U2994  ( .A(\GFM/n1443 ), .B(\GFM/n14420 ), .Z(\GFM/n1435 ) );
XOR2_X2 \GFM/U2993  ( .A(z_in[83]), .B(\GFM/n14440 ), .Z(\GFM/n14360 ) );
XOR2_X2 \GFM/U2992  ( .A(\GFM/N2600 ), .B(\GFM/N2601 ), .Z(\GFM/n14370 ) );
XOR2_X2 \GFM/U2991  ( .A(\GFM/N2597 ), .B(\GFM/N2598 ), .Z(\GFM/n1438 ) );
XOR2_X2 \GFM/U2990  ( .A(\GFM/N2593 ), .B(\GFM/N2594 ), .Z(\GFM/n1439 ) );
XOR2_X2 \GFM/U2989  ( .A(\GFM/N2589 ), .B(\GFM/N2591 ), .Z(\GFM/n1440 ) );
XOR2_X2 \GFM/U2988  ( .A(\GFM/N2584 ), .B(\GFM/N2588 ), .Z(\GFM/n14410 ) );
XOR2_X2 \GFM/U2987  ( .A(\GFM/N2581 ), .B(\GFM/N2583 ), .Z(\GFM/n14420 ) );
XOR2_X2 \GFM/U2986  ( .A(\GFM/N2577 ), .B(\GFM/N2580 ), .Z(\GFM/n1443 ) );
XOR2_X2 \GFM/U2985  ( .A(\GFM/N2574 ), .B(\GFM/N2576 ), .Z(\GFM/n14440 ) );
XOR2_X2 \GFM/U2984  ( .A(\GFM/n14460 ), .B(\GFM/n1445 ), .Z(z_out[84]) );
XOR2_X2 \GFM/U2983  ( .A(\GFM/n1448 ), .B(\GFM/n14470 ), .Z(\GFM/n1445 ) );
XOR2_X2 \GFM/U2982  ( .A(\GFM/n14500 ), .B(\GFM/n1449 ), .Z(\GFM/n14460 ) );
XOR2_X2 \GFM/U2981  ( .A(\GFM/n1452 ), .B(\GFM/n14510 ), .Z(\GFM/n14470 ) );
XOR2_X2 \GFM/U2980  ( .A(\GFM/n14540 ), .B(\GFM/n14530 ), .Z(\GFM/n1448 ) );
XOR2_X2 \GFM/U2979  ( .A(\GFM/n1456 ), .B(\GFM/n1455 ), .Z(\GFM/n1449 ) );
XOR2_X2 \GFM/U2978  ( .A(\GFM/n14580 ), .B(\GFM/n1457 ), .Z(\GFM/n14500 ) );
XOR2_X2 \GFM/U2977  ( .A(z_in[84]), .B(\GFM/n1459 ), .Z(\GFM/n14510 ) );
XOR2_X2 \GFM/U2976  ( .A(\GFM/N2631 ), .B(\GFM/N2632 ), .Z(\GFM/n1452 ) );
XOR2_X2 \GFM/U2975  ( .A(\GFM/N2628 ), .B(\GFM/N2629 ), .Z(\GFM/n14530 ) );
XOR2_X2 \GFM/U2974  ( .A(\GFM/N2624 ), .B(\GFM/N2625 ), .Z(\GFM/n14540 ) );
XOR2_X2 \GFM/U2973  ( .A(\GFM/N2620 ), .B(\GFM/N2622 ), .Z(\GFM/n1455 ) );
XOR2_X2 \GFM/U2972  ( .A(\GFM/N2615 ), .B(\GFM/N2619 ), .Z(\GFM/n1456 ) );
XOR2_X2 \GFM/U2971  ( .A(\GFM/N2612 ), .B(\GFM/N2614 ), .Z(\GFM/n1457 ) );
XOR2_X2 \GFM/U2970  ( .A(\GFM/N2608 ), .B(\GFM/N2611 ), .Z(\GFM/n14580 ) );
XOR2_X2 \GFM/U2969  ( .A(\GFM/N2605 ), .B(\GFM/N2607 ), .Z(\GFM/n1459 ) );
XOR2_X2 \GFM/U2968  ( .A(\GFM/n14610 ), .B(\GFM/n14600 ), .Z(z_out[85]) );
XOR2_X2 \GFM/U2967  ( .A(\GFM/n1463 ), .B(\GFM/n1462 ), .Z(\GFM/n14600 ) );
XOR2_X2 \GFM/U2966  ( .A(\GFM/n14650 ), .B(\GFM/n14640 ), .Z(\GFM/n14610 ));
XOR2_X2 \GFM/U2965  ( .A(\GFM/n14670 ), .B(\GFM/n1466 ), .Z(\GFM/n1462 ) );
XOR2_X2 \GFM/U2964  ( .A(\GFM/n1469 ), .B(\GFM/n14680 ), .Z(\GFM/n1463 ) );
XOR2_X2 \GFM/U2963  ( .A(\GFM/n1471 ), .B(\GFM/n1470 ), .Z(\GFM/n14640 ) );
XOR2_X2 \GFM/U2962  ( .A(\GFM/n14730 ), .B(\GFM/n14720 ), .Z(\GFM/n14650 ));
XOR2_X2 \GFM/U2961  ( .A(z_in[85]), .B(\GFM/n1474 ), .Z(\GFM/n1466 ) );
XOR2_X2 \GFM/U2960  ( .A(\GFM/N2662 ), .B(\GFM/N2663 ), .Z(\GFM/n14670 ) );
XOR2_X2 \GFM/U2959  ( .A(\GFM/N2659 ), .B(\GFM/N2660 ), .Z(\GFM/n14680 ) );
XOR2_X2 \GFM/U2958  ( .A(\GFM/N2655 ), .B(\GFM/N2656 ), .Z(\GFM/n1469 ) );
XOR2_X2 \GFM/U2957  ( .A(\GFM/N2651 ), .B(\GFM/N2653 ), .Z(\GFM/n1470 ) );
XOR2_X2 \GFM/U2956  ( .A(\GFM/N2646 ), .B(\GFM/N2650 ), .Z(\GFM/n1471 ) );
XOR2_X2 \GFM/U2955  ( .A(\GFM/N2643 ), .B(\GFM/N2645 ), .Z(\GFM/n14720 ) );
XOR2_X2 \GFM/U2954  ( .A(\GFM/N2639 ), .B(\GFM/N2642 ), .Z(\GFM/n14730 ) );
XOR2_X2 \GFM/U2953  ( .A(\GFM/N2636 ), .B(\GFM/N2638 ), .Z(\GFM/n1474 ) );
XOR2_X2 \GFM/U2952  ( .A(\GFM/n1476 ), .B(\GFM/n14750 ), .Z(z_out[86]) );
XOR2_X2 \GFM/U2951  ( .A(\GFM/n14780 ), .B(\GFM/n14770 ), .Z(\GFM/n14750 ));
XOR2_X2 \GFM/U2950  ( .A(\GFM/n1480 ), .B(\GFM/n1479 ), .Z(\GFM/n1476 ) );
XOR2_X2 \GFM/U2949  ( .A(\GFM/n14820 ), .B(\GFM/n14810 ), .Z(\GFM/n14770 ));
XOR2_X2 \GFM/U2948  ( .A(\GFM/n14840 ), .B(\GFM/n1483 ), .Z(\GFM/n14780 ) );
XOR2_X2 \GFM/U2947  ( .A(\GFM/n1486 ), .B(\GFM/n14850 ), .Z(\GFM/n1479 ) );
XOR2_X2 \GFM/U2946  ( .A(\GFM/n1488 ), .B(\GFM/n1487 ), .Z(\GFM/n1480 ) );
XOR2_X2 \GFM/U2945  ( .A(z_in[86]), .B(\GFM/n14890 ), .Z(\GFM/n14810 ) );
XOR2_X2 \GFM/U2944  ( .A(\GFM/N2693 ), .B(\GFM/N2694 ), .Z(\GFM/n14820 ) );
XOR2_X2 \GFM/U2943  ( .A(\GFM/N2690 ), .B(\GFM/N2691 ), .Z(\GFM/n1483 ) );
XOR2_X2 \GFM/U2942  ( .A(\GFM/N2686 ), .B(\GFM/N2687 ), .Z(\GFM/n14840 ) );
XOR2_X2 \GFM/U2941  ( .A(\GFM/N2682 ), .B(\GFM/N2684 ), .Z(\GFM/n14850 ) );
XOR2_X2 \GFM/U2940  ( .A(\GFM/N2677 ), .B(\GFM/N2681 ), .Z(\GFM/n1486 ) );
XOR2_X2 \GFM/U2939  ( .A(\GFM/N2674 ), .B(\GFM/N2676 ), .Z(\GFM/n1487 ) );
XOR2_X2 \GFM/U2938  ( .A(\GFM/N2670 ), .B(\GFM/N2673 ), .Z(\GFM/n1488 ) );
XOR2_X2 \GFM/U2937  ( .A(\GFM/N2667 ), .B(\GFM/N2669 ), .Z(\GFM/n14890 ) );
XOR2_X2 \GFM/U2936  ( .A(\GFM/n14910 ), .B(\GFM/n1490 ), .Z(z_out[87]) );
XOR2_X2 \GFM/U2935  ( .A(\GFM/n1493 ), .B(\GFM/n14920 ), .Z(\GFM/n1490 ) );
XOR2_X2 \GFM/U2934  ( .A(\GFM/n14950 ), .B(\GFM/n1494 ), .Z(\GFM/n14910 ) );
XOR2_X2 \GFM/U2933  ( .A(\GFM/n1497 ), .B(\GFM/n14960 ), .Z(\GFM/n14920 ) );
XOR2_X2 \GFM/U2932  ( .A(\GFM/n14990 ), .B(\GFM/n14980 ), .Z(\GFM/n1493 ) );
XOR2_X2 \GFM/U2931  ( .A(\GFM/n1501 ), .B(\GFM/n1500 ), .Z(\GFM/n1494 ) );
XOR2_X2 \GFM/U2930  ( .A(\GFM/n15030 ), .B(\GFM/n1502 ), .Z(\GFM/n14950 ) );
XOR2_X2 \GFM/U2929  ( .A(z_in[87]), .B(\GFM/n15040 ), .Z(\GFM/n14960 ) );
XOR2_X2 \GFM/U2928  ( .A(\GFM/N2724 ), .B(\GFM/N2725 ), .Z(\GFM/n1497 ) );
XOR2_X2 \GFM/U2927  ( .A(\GFM/N2721 ), .B(\GFM/N2722 ), .Z(\GFM/n14980 ) );
XOR2_X2 \GFM/U2926  ( .A(\GFM/N2717 ), .B(\GFM/N2718 ), .Z(\GFM/n14990 ) );
XOR2_X2 \GFM/U2925  ( .A(\GFM/N2713 ), .B(\GFM/N2715 ), .Z(\GFM/n1500 ) );
XOR2_X2 \GFM/U2924  ( .A(\GFM/N2708 ), .B(\GFM/N2712 ), .Z(\GFM/n1501 ) );
XOR2_X2 \GFM/U2923  ( .A(\GFM/N2705 ), .B(\GFM/N2707 ), .Z(\GFM/n1502 ) );
XOR2_X2 \GFM/U2922  ( .A(\GFM/N2701 ), .B(\GFM/N2704 ), .Z(\GFM/n15030 ) );
XOR2_X2 \GFM/U2921  ( .A(\GFM/N2698 ), .B(\GFM/N2700 ), .Z(\GFM/n15040 ) );
XOR2_X2 \GFM/U2920  ( .A(\GFM/n15060 ), .B(\GFM/n1505 ), .Z(z_out[88]) );
XOR2_X2 \GFM/U2919  ( .A(\GFM/n15080 ), .B(\GFM/n1507 ), .Z(\GFM/n1505 ) );
XOR2_X2 \GFM/U2918  ( .A(\GFM/n1510 ), .B(\GFM/n15090 ), .Z(\GFM/n15060 ) );
XOR2_X2 \GFM/U2917  ( .A(\GFM/n15120 ), .B(\GFM/n1511 ), .Z(\GFM/n1507 ) );
XOR2_X2 \GFM/U2916  ( .A(\GFM/n1514 ), .B(\GFM/n15130 ), .Z(\GFM/n15080 ) );
XOR2_X2 \GFM/U2915  ( .A(\GFM/n15160 ), .B(\GFM/n15150 ), .Z(\GFM/n15090 ));
XOR2_X2 \GFM/U2914  ( .A(\GFM/n1518 ), .B(\GFM/n1517 ), .Z(\GFM/n1510 ) );
XOR2_X2 \GFM/U2913  ( .A(z_in[88]), .B(\GFM/n1519 ), .Z(\GFM/n1511 ) );
XOR2_X2 \GFM/U2912  ( .A(\GFM/N2755 ), .B(\GFM/N2756 ), .Z(\GFM/n15120 ) );
XOR2_X2 \GFM/U2911  ( .A(\GFM/N2752 ), .B(\GFM/N2753 ), .Z(\GFM/n15130 ) );
XOR2_X2 \GFM/U2910  ( .A(\GFM/N2748 ), .B(\GFM/N2749 ), .Z(\GFM/n1514 ) );
XOR2_X2 \GFM/U2909  ( .A(\GFM/N2744 ), .B(\GFM/N2746 ), .Z(\GFM/n15150 ) );
XOR2_X2 \GFM/U2908  ( .A(\GFM/N2739 ), .B(\GFM/N2743 ), .Z(\GFM/n15160 ) );
XOR2_X2 \GFM/U2907  ( .A(\GFM/N2736 ), .B(\GFM/N2738 ), .Z(\GFM/n1517 ) );
XOR2_X2 \GFM/U2906  ( .A(\GFM/N2732 ), .B(\GFM/N2735 ), .Z(\GFM/n1518 ) );
XOR2_X2 \GFM/U2905  ( .A(\GFM/N2729 ), .B(\GFM/N2731 ), .Z(\GFM/n1519 ) );
XOR2_X2 \GFM/U2904  ( .A(\GFM/n1521 ), .B(\GFM/n15200 ), .Z(z_out[89]) );
XOR2_X2 \GFM/U2903  ( .A(\GFM/n15230 ), .B(\GFM/n15220 ), .Z(\GFM/n15200 ));
XOR2_X2 \GFM/U2902  ( .A(\GFM/n1525 ), .B(\GFM/n1524 ), .Z(\GFM/n1521 ) );
XOR2_X2 \GFM/U2901  ( .A(\GFM/n15270 ), .B(\GFM/n15260 ), .Z(\GFM/n15220 ));
XOR2_X2 \GFM/U2900  ( .A(\GFM/n15290 ), .B(\GFM/n1528 ), .Z(\GFM/n15230 ) );
XOR2_X2 \GFM/U2899  ( .A(\GFM/n1531 ), .B(\GFM/n15300 ), .Z(\GFM/n1524 ) );
XOR2_X2 \GFM/U2898  ( .A(\GFM/n1533 ), .B(\GFM/n1532 ), .Z(\GFM/n1525 ) );
XOR2_X2 \GFM/U2897  ( .A(z_in[89]), .B(\GFM/n15340 ), .Z(\GFM/n15260 ) );
XOR2_X2 \GFM/U2896  ( .A(\GFM/N2786 ), .B(\GFM/N2787 ), .Z(\GFM/n15270 ) );
XOR2_X2 \GFM/U2895  ( .A(\GFM/N2783 ), .B(\GFM/N2784 ), .Z(\GFM/n1528 ) );
XOR2_X2 \GFM/U2894  ( .A(\GFM/N2779 ), .B(\GFM/N2780 ), .Z(\GFM/n15290 ) );
XOR2_X2 \GFM/U2893  ( .A(\GFM/N2775 ), .B(\GFM/N2777 ), .Z(\GFM/n15300 ) );
XOR2_X2 \GFM/U2892  ( .A(\GFM/N2770 ), .B(\GFM/N2774 ), .Z(\GFM/n1531 ) );
XOR2_X2 \GFM/U2891  ( .A(\GFM/N2767 ), .B(\GFM/N2769 ), .Z(\GFM/n1532 ) );
XOR2_X2 \GFM/U2890  ( .A(\GFM/N2763 ), .B(\GFM/N2766 ), .Z(\GFM/n1533 ) );
XOR2_X2 \GFM/U2889  ( .A(\GFM/N2760 ), .B(\GFM/N2762 ), .Z(\GFM/n15340 ) );
XOR2_X2 \GFM/U2888  ( .A(\GFM/n1536 ), .B(\GFM/n15350 ), .Z(z_out[90]) );
XOR2_X2 \GFM/U2887  ( .A(\GFM/n1538 ), .B(\GFM/n15370 ), .Z(\GFM/n15350 ) );
XOR2_X2 \GFM/U2886  ( .A(\GFM/n15400 ), .B(\GFM/n15390 ), .Z(\GFM/n1536 ) );
XOR2_X2 \GFM/U2885  ( .A(\GFM/n1542 ), .B(\GFM/n1541 ), .Z(\GFM/n15370 ) );
XOR2_X2 \GFM/U2884  ( .A(\GFM/n15440 ), .B(\GFM/n15430 ), .Z(\GFM/n1538 ) );
XOR2_X2 \GFM/U2883  ( .A(\GFM/n15460 ), .B(\GFM/n1545 ), .Z(\GFM/n15390 ) );
XOR2_X2 \GFM/U2882  ( .A(\GFM/n1548 ), .B(\GFM/n15470 ), .Z(\GFM/n15400 ) );
XOR2_X2 \GFM/U2881  ( .A(z_in[90]), .B(\GFM/n1549 ), .Z(\GFM/n1541 ) );
XOR2_X2 \GFM/U2880  ( .A(\GFM/N2817 ), .B(\GFM/N2818 ), .Z(\GFM/n1542 ) );
XOR2_X2 \GFM/U2879  ( .A(\GFM/N2814 ), .B(\GFM/N2815 ), .Z(\GFM/n15430 ) );
XOR2_X2 \GFM/U2878  ( .A(\GFM/N2810 ), .B(\GFM/N2811 ), .Z(\GFM/n15440 ) );
XOR2_X2 \GFM/U2877  ( .A(\GFM/N2806 ), .B(\GFM/N2808 ), .Z(\GFM/n1545 ) );
XOR2_X2 \GFM/U2876  ( .A(\GFM/N2801 ), .B(\GFM/N2805 ), .Z(\GFM/n15460 ) );
XOR2_X2 \GFM/U2875  ( .A(\GFM/N2798 ), .B(\GFM/N2800 ), .Z(\GFM/n15470 ) );
XOR2_X2 \GFM/U2874  ( .A(\GFM/N2794 ), .B(\GFM/N2797 ), .Z(\GFM/n1548 ) );
XOR2_X2 \GFM/U2873  ( .A(\GFM/N2791 ), .B(\GFM/N2793 ), .Z(\GFM/n1549 ) );
XOR2_X2 \GFM/U2872  ( .A(\GFM/n15510 ), .B(\GFM/n1550 ), .Z(z_out[91]) );
XOR2_X2 \GFM/U2871  ( .A(\GFM/n15530 ), .B(\GFM/n1552 ), .Z(\GFM/n1550 ) );
XOR2_X2 \GFM/U2870  ( .A(\GFM/n1555 ), .B(\GFM/n15540 ), .Z(\GFM/n15510 ) );
XOR2_X2 \GFM/U2869  ( .A(\GFM/n15570 ), .B(\GFM/n1556 ), .Z(\GFM/n1552 ) );
XOR2_X2 \GFM/U2868  ( .A(\GFM/n1559 ), .B(\GFM/n15580 ), .Z(\GFM/n15530 ) );
XOR2_X2 \GFM/U2867  ( .A(\GFM/n15610 ), .B(\GFM/n15600 ), .Z(\GFM/n15540 ));
XOR2_X2 \GFM/U2866  ( .A(\GFM/n1563 ), .B(\GFM/n1562 ), .Z(\GFM/n1555 ) );
XOR2_X2 \GFM/U2865  ( .A(z_in[91]), .B(\GFM/n1564 ), .Z(\GFM/n1556 ) );
XOR2_X2 \GFM/U2864  ( .A(\GFM/N2848 ), .B(\GFM/N2849 ), .Z(\GFM/n15570 ) );
XOR2_X2 \GFM/U2863  ( .A(\GFM/N2845 ), .B(\GFM/N2846 ), .Z(\GFM/n15580 ) );
XOR2_X2 \GFM/U2862  ( .A(\GFM/N2841 ), .B(\GFM/N2842 ), .Z(\GFM/n1559 ) );
XOR2_X2 \GFM/U2861  ( .A(\GFM/N2837 ), .B(\GFM/N2839 ), .Z(\GFM/n15600 ) );
XOR2_X2 \GFM/U2860  ( .A(\GFM/N2832 ), .B(\GFM/N2836 ), .Z(\GFM/n15610 ) );
XOR2_X2 \GFM/U2859  ( .A(\GFM/N2829 ), .B(\GFM/N2831 ), .Z(\GFM/n1562 ) );
XOR2_X2 \GFM/U2858  ( .A(\GFM/N2825 ), .B(\GFM/N2828 ), .Z(\GFM/n1563 ) );
XOR2_X2 \GFM/U2857  ( .A(\GFM/N2822 ), .B(\GFM/N2824 ), .Z(\GFM/n1564 ) );
XOR2_X2 \GFM/U2856  ( .A(\GFM/n15660 ), .B(\GFM/n15650 ), .Z(z_out[92]) );
XOR2_X2 \GFM/U2855  ( .A(\GFM/n15680 ), .B(\GFM/n1567 ), .Z(\GFM/n15650 ) );
XOR2_X2 \GFM/U2854  ( .A(\GFM/n15700 ), .B(\GFM/n1569 ), .Z(\GFM/n15660 ) );
XOR2_X2 \GFM/U2853  ( .A(\GFM/n1572 ), .B(\GFM/n15710 ), .Z(\GFM/n1567 ) );
XOR2_X2 \GFM/U2852  ( .A(\GFM/n15740 ), .B(\GFM/n1573 ), .Z(\GFM/n15680 ) );
XOR2_X2 \GFM/U2851  ( .A(\GFM/n1576 ), .B(\GFM/n15750 ), .Z(\GFM/n1569 ) );
XOR2_X2 \GFM/U2850  ( .A(\GFM/n15780 ), .B(\GFM/n15770 ), .Z(\GFM/n15700 ));
XOR2_X2 \GFM/U2849  ( .A(z_in[92]), .B(\GFM/n1579 ), .Z(\GFM/n15710 ) );
XOR2_X2 \GFM/U2848  ( .A(\GFM/N2879 ), .B(\GFM/N2880 ), .Z(\GFM/n1572 ) );
XOR2_X2 \GFM/U2847  ( .A(\GFM/N2876 ), .B(\GFM/N2877 ), .Z(\GFM/n1573 ) );
XOR2_X2 \GFM/U2846  ( .A(\GFM/N2872 ), .B(\GFM/N2873 ), .Z(\GFM/n15740 ) );
XOR2_X2 \GFM/U2845  ( .A(\GFM/N2868 ), .B(\GFM/N2870 ), .Z(\GFM/n15750 ) );
XOR2_X2 \GFM/U2844  ( .A(\GFM/N2863 ), .B(\GFM/N2867 ), .Z(\GFM/n1576 ) );
XOR2_X2 \GFM/U2843  ( .A(\GFM/N2860 ), .B(\GFM/N2862 ), .Z(\GFM/n15770 ) );
XOR2_X2 \GFM/U2842  ( .A(\GFM/N2856 ), .B(\GFM/N2859 ), .Z(\GFM/n15780 ) );
XOR2_X2 \GFM/U2841  ( .A(\GFM/N2853 ), .B(\GFM/N2855 ), .Z(\GFM/n1579 ) );
XOR2_X2 \GFM/U2840  ( .A(\GFM/n1581 ), .B(\GFM/n1580 ), .Z(z_out[93]) );
XOR2_X2 \GFM/U2839  ( .A(\GFM/n1583 ), .B(\GFM/n15820 ), .Z(\GFM/n1580 ) );
XOR2_X2 \GFM/U2838  ( .A(\GFM/n15850 ), .B(\GFM/n15840 ), .Z(\GFM/n1581 ) );
XOR2_X2 \GFM/U2837  ( .A(\GFM/n1587 ), .B(\GFM/n1586 ), .Z(\GFM/n15820 ) );
XOR2_X2 \GFM/U2836  ( .A(\GFM/n15890 ), .B(\GFM/n15880 ), .Z(\GFM/n1583 ) );
XOR2_X2 \GFM/U2835  ( .A(\GFM/n15910 ), .B(\GFM/n1590 ), .Z(\GFM/n15840 ) );
XOR2_X2 \GFM/U2834  ( .A(\GFM/n1593 ), .B(\GFM/n15920 ), .Z(\GFM/n15850 ) );
XOR2_X2 \GFM/U2833  ( .A(z_in[93]), .B(\GFM/n1594 ), .Z(\GFM/n1586 ) );
XOR2_X2 \GFM/U2832  ( .A(\GFM/N2910 ), .B(\GFM/N2911 ), .Z(\GFM/n1587 ) );
XOR2_X2 \GFM/U2831  ( .A(\GFM/N2907 ), .B(\GFM/N2908 ), .Z(\GFM/n15880 ) );
XOR2_X2 \GFM/U2830  ( .A(\GFM/N2903 ), .B(\GFM/N2904 ), .Z(\GFM/n15890 ) );
XOR2_X2 \GFM/U2829  ( .A(\GFM/N2899 ), .B(\GFM/N2901 ), .Z(\GFM/n1590 ) );
XOR2_X2 \GFM/U2828  ( .A(\GFM/N2894 ), .B(\GFM/N2898 ), .Z(\GFM/n15910 ) );
XOR2_X2 \GFM/U2827  ( .A(\GFM/N2891 ), .B(\GFM/N2893 ), .Z(\GFM/n15920 ) );
XOR2_X2 \GFM/U2826  ( .A(\GFM/N2887 ), .B(\GFM/N2890 ), .Z(\GFM/n1593 ) );
XOR2_X2 \GFM/U2825  ( .A(\GFM/N2884 ), .B(\GFM/N2886 ), .Z(\GFM/n1594 ) );
XOR2_X2 \GFM/U2824  ( .A(\GFM/n15960 ), .B(\GFM/n1595 ), .Z(z_out[94]) );
XOR2_X2 \GFM/U2823  ( .A(\GFM/n1598 ), .B(\GFM/n15970 ), .Z(\GFM/n1595 ) );
XOR2_X2 \GFM/U2822  ( .A(\GFM/n1600 ), .B(\GFM/n15990 ), .Z(\GFM/n15960 ) );
XOR2_X2 \GFM/U2821  ( .A(\GFM/n16020 ), .B(\GFM/n16010 ), .Z(\GFM/n15970 ));
XOR2_X2 \GFM/U2820  ( .A(\GFM/n1604 ), .B(\GFM/n1603 ), .Z(\GFM/n1598 ) );
XOR2_X2 \GFM/U2819  ( .A(\GFM/n16060 ), .B(\GFM/n16050 ), .Z(\GFM/n15990 ));
XOR2_X2 \GFM/U2818  ( .A(\GFM/n16080 ), .B(\GFM/n1607 ), .Z(\GFM/n1600 ) );
XOR2_X2 \GFM/U2817  ( .A(z_in[94]), .B(\GFM/n16090 ), .Z(\GFM/n16010 ) );
XOR2_X2 \GFM/U2816  ( .A(\GFM/N2941 ), .B(\GFM/N2942 ), .Z(\GFM/n16020 ) );
XOR2_X2 \GFM/U2815  ( .A(\GFM/N2938 ), .B(\GFM/N2939 ), .Z(\GFM/n1603 ) );
XOR2_X2 \GFM/U2814  ( .A(\GFM/N2934 ), .B(\GFM/N2935 ), .Z(\GFM/n1604 ) );
XOR2_X2 \GFM/U2813  ( .A(\GFM/N2930 ), .B(\GFM/N2932 ), .Z(\GFM/n16050 ) );
XOR2_X2 \GFM/U2812  ( .A(\GFM/N2925 ), .B(\GFM/N2929 ), .Z(\GFM/n16060 ) );
XOR2_X2 \GFM/U2811  ( .A(\GFM/N2922 ), .B(\GFM/N2924 ), .Z(\GFM/n1607 ) );
XOR2_X2 \GFM/U2810  ( .A(\GFM/N2918 ), .B(\GFM/N2921 ), .Z(\GFM/n16080 ) );
XOR2_X2 \GFM/U2809  ( .A(\GFM/N2915 ), .B(\GFM/N2917 ), .Z(\GFM/n16090 ) );
XOR2_X2 \GFM/U2808  ( .A(\GFM/n1611 ), .B(\GFM/n1610 ), .Z(z_out[95]) );
XOR2_X2 \GFM/U2807  ( .A(\GFM/n16130 ), .B(\GFM/n1612 ), .Z(\GFM/n1610 ) );
XOR2_X2 \GFM/U2806  ( .A(\GFM/n16150 ), .B(\GFM/n1614 ), .Z(\GFM/n1611 ) );
XOR2_X2 \GFM/U2805  ( .A(\GFM/n1617 ), .B(\GFM/n16160 ), .Z(\GFM/n1612 ) );
XOR2_X2 \GFM/U2804  ( .A(\GFM/n16190 ), .B(\GFM/n1618 ), .Z(\GFM/n16130 ) );
XOR2_X2 \GFM/U2803  ( .A(\GFM/n1621 ), .B(\GFM/n16200 ), .Z(\GFM/n1614 ) );
XOR2_X2 \GFM/U2802  ( .A(\GFM/n16230 ), .B(\GFM/n16220 ), .Z(\GFM/n16150 ));
XOR2_X2 \GFM/U2801  ( .A(z_in[95]), .B(\GFM/n1624 ), .Z(\GFM/n16160 ) );
XOR2_X2 \GFM/U2800  ( .A(\GFM/N2972 ), .B(\GFM/N2973 ), .Z(\GFM/n1617 ) );
XOR2_X2 \GFM/U2799  ( .A(\GFM/N2969 ), .B(\GFM/N2970 ), .Z(\GFM/n1618 ) );
XOR2_X2 \GFM/U2798  ( .A(\GFM/N2965 ), .B(\GFM/N2966 ), .Z(\GFM/n16190 ) );
XOR2_X2 \GFM/U2797  ( .A(\GFM/N2961 ), .B(\GFM/N2963 ), .Z(\GFM/n16200 ) );
XOR2_X2 \GFM/U2796  ( .A(\GFM/N2956 ), .B(\GFM/N2960 ), .Z(\GFM/n1621 ) );
XOR2_X2 \GFM/U2795  ( .A(\GFM/N2953 ), .B(\GFM/N2955 ), .Z(\GFM/n16220 ) );
XOR2_X2 \GFM/U2794  ( .A(\GFM/N2949 ), .B(\GFM/N2952 ), .Z(\GFM/n16230 ) );
XOR2_X2 \GFM/U2793  ( .A(\GFM/N2946 ), .B(\GFM/N2948 ), .Z(\GFM/n1624 ) );
XOR2_X2 \GFM/U2792  ( .A(\GFM/n1626 ), .B(\GFM/n1625 ), .Z(z_out[96]) );
XOR2_X2 \GFM/U2791  ( .A(\GFM/n16280 ), .B(\GFM/n16270 ), .Z(\GFM/n1625 ) );
XOR2_X2 \GFM/U2790  ( .A(\GFM/n16300 ), .B(\GFM/n1629 ), .Z(\GFM/n1626 ) );
XOR2_X2 \GFM/U2789  ( .A(\GFM/n16320 ), .B(\GFM/n1631 ), .Z(\GFM/n16270 ) );
XOR2_X2 \GFM/U2788  ( .A(\GFM/n1634 ), .B(\GFM/n16330 ), .Z(\GFM/n16280 ) );
XOR2_X2 \GFM/U2787  ( .A(\GFM/n16360 ), .B(\GFM/n1635 ), .Z(\GFM/n1629 ) );
XOR2_X2 \GFM/U2786  ( .A(\GFM/n1638 ), .B(\GFM/n16370 ), .Z(\GFM/n16300 ) );
XOR2_X2 \GFM/U2785  ( .A(z_in[96]), .B(\GFM/n16390 ), .Z(\GFM/n1631 ) );
XOR2_X2 \GFM/U2784  ( .A(\GFM/N3003 ), .B(\GFM/N3004 ), .Z(\GFM/n16320 ) );
XOR2_X2 \GFM/U2783  ( .A(\GFM/N3000 ), .B(\GFM/N3001 ), .Z(\GFM/n16330 ) );
XOR2_X2 \GFM/U2782  ( .A(\GFM/N2996 ), .B(\GFM/N2997 ), .Z(\GFM/n1634 ) );
XOR2_X2 \GFM/U2781  ( .A(\GFM/N2992 ), .B(\GFM/N2994 ), .Z(\GFM/n1635 ) );
XOR2_X2 \GFM/U2780  ( .A(\GFM/N2987 ), .B(\GFM/N2991 ), .Z(\GFM/n16360 ) );
XOR2_X2 \GFM/U2779  ( .A(\GFM/N2984 ), .B(\GFM/N2986 ), .Z(\GFM/n16370 ) );
XOR2_X2 \GFM/U2778  ( .A(\GFM/N2980 ), .B(\GFM/N2983 ), .Z(\GFM/n1638 ) );
XOR2_X2 \GFM/U2777  ( .A(\GFM/N2977 ), .B(\GFM/N2979 ), .Z(\GFM/n16390 ) );
XOR2_X2 \GFM/U2776  ( .A(\GFM/n1641 ), .B(\GFM/n16400 ), .Z(z_out[97]) );
XOR2_X2 \GFM/U2775  ( .A(\GFM/n1643 ), .B(\GFM/n1642 ), .Z(\GFM/n16400 ) );
XOR2_X2 \GFM/U2774  ( .A(\GFM/n1645 ), .B(\GFM/n16440 ), .Z(\GFM/n1641 ) );
XOR2_X2 \GFM/U2773  ( .A(\GFM/n16470 ), .B(\GFM/n16460 ), .Z(\GFM/n1642 ) );
XOR2_X2 \GFM/U2772  ( .A(\GFM/n1649 ), .B(\GFM/n1648 ), .Z(\GFM/n1643 ) );
XOR2_X2 \GFM/U2771  ( .A(\GFM/n16510 ), .B(\GFM/n16500 ), .Z(\GFM/n16440 ));
XOR2_X2 \GFM/U2770  ( .A(\GFM/n16530 ), .B(\GFM/n1652 ), .Z(\GFM/n1645 ) );
XOR2_X2 \GFM/U2769  ( .A(z_in[97]), .B(\GFM/n16540 ), .Z(\GFM/n16460 ) );
XOR2_X2 \GFM/U2768  ( .A(\GFM/N3034 ), .B(\GFM/N3035 ), .Z(\GFM/n16470 ) );
XOR2_X2 \GFM/U2767  ( .A(\GFM/N3031 ), .B(\GFM/N3032 ), .Z(\GFM/n1648 ) );
XOR2_X2 \GFM/U2766  ( .A(\GFM/N3027 ), .B(\GFM/N3028 ), .Z(\GFM/n1649 ) );
XOR2_X2 \GFM/U2765  ( .A(\GFM/N3023 ), .B(\GFM/N3025 ), .Z(\GFM/n16500 ) );
XOR2_X2 \GFM/U2764  ( .A(\GFM/N3018 ), .B(\GFM/N3022 ), .Z(\GFM/n16510 ) );
XOR2_X2 \GFM/U2763  ( .A(\GFM/N3015 ), .B(\GFM/N3017 ), .Z(\GFM/n1652 ) );
XOR2_X2 \GFM/U2762  ( .A(\GFM/N3011 ), .B(\GFM/N3014 ), .Z(\GFM/n16530 ) );
XOR2_X2 \GFM/U2761  ( .A(\GFM/N3008 ), .B(\GFM/N3010 ), .Z(\GFM/n16540 ) );
XOR2_X2 \GFM/U2760  ( .A(\GFM/n1656 ), .B(\GFM/n1655 ), .Z(z_out[98]) );
XOR2_X2 \GFM/U2759  ( .A(\GFM/n16580 ), .B(\GFM/n1657 ), .Z(\GFM/n1655 ) );
XOR2_X2 \GFM/U2758  ( .A(\GFM/n1660 ), .B(\GFM/n16590 ), .Z(\GFM/n1656 ) );
XOR2_X2 \GFM/U2757  ( .A(\GFM/n1662 ), .B(\GFM/n16610 ), .Z(\GFM/n1657 ) );
XOR2_X2 \GFM/U2756  ( .A(\GFM/n16640 ), .B(\GFM/n16630 ), .Z(\GFM/n16580 ));
XOR2_X2 \GFM/U2755  ( .A(\GFM/n1666 ), .B(\GFM/n1665 ), .Z(\GFM/n16590 ) );
XOR2_X2 \GFM/U2754  ( .A(\GFM/n16680 ), .B(\GFM/n16670 ), .Z(\GFM/n1660 ) );
XOR2_X2 \GFM/U2753  ( .A(z_in[98]), .B(\GFM/n1669 ), .Z(\GFM/n16610 ) );
XOR2_X2 \GFM/U2752  ( .A(\GFM/N3065 ), .B(\GFM/N3066 ), .Z(\GFM/n1662 ) );
XOR2_X2 \GFM/U2751  ( .A(\GFM/N3062 ), .B(\GFM/N3063 ), .Z(\GFM/n16630 ) );
XOR2_X2 \GFM/U2750  ( .A(\GFM/N3058 ), .B(\GFM/N3059 ), .Z(\GFM/n16640 ) );
XOR2_X2 \GFM/U2749  ( .A(\GFM/N3054 ), .B(\GFM/N3056 ), .Z(\GFM/n1665 ) );
XOR2_X2 \GFM/U2748  ( .A(\GFM/N3049 ), .B(\GFM/N3053 ), .Z(\GFM/n1666 ) );
XOR2_X2 \GFM/U2747  ( .A(\GFM/N3046 ), .B(\GFM/N3048 ), .Z(\GFM/n16670 ) );
XOR2_X2 \GFM/U2746  ( .A(\GFM/N3042 ), .B(\GFM/N3045 ), .Z(\GFM/n16680 ) );
XOR2_X2 \GFM/U2745  ( .A(\GFM/N3039 ), .B(\GFM/N3041 ), .Z(\GFM/n1669 ) );
XOR2_X2 \GFM/U2744  ( .A(\GFM/n16710 ), .B(\GFM/n16700 ), .Z(z_out[99]) );
XOR2_X2 \GFM/U2743  ( .A(\GFM/n1673 ), .B(\GFM/n1672 ), .Z(\GFM/n16700 ) );
XOR2_X2 \GFM/U2742  ( .A(\GFM/n16750 ), .B(\GFM/n1674 ), .Z(\GFM/n16710 ) );
XOR2_X2 \GFM/U2741  ( .A(\GFM/n16770 ), .B(\GFM/n1676 ), .Z(\GFM/n1672 ) );
XOR2_X2 \GFM/U2740  ( .A(\GFM/n1679 ), .B(\GFM/n16780 ), .Z(\GFM/n1673 ) );
XOR2_X2 \GFM/U2739  ( .A(\GFM/n16810 ), .B(\GFM/n1680 ), .Z(\GFM/n1674 ) );
XOR2_X2 \GFM/U2738  ( .A(\GFM/n1683 ), .B(\GFM/n16820 ), .Z(\GFM/n16750 ) );
XOR2_X2 \GFM/U2737  ( .A(z_in[99]), .B(\GFM/n16840 ), .Z(\GFM/n1676 ) );
XOR2_X2 \GFM/U2736  ( .A(\GFM/N3096 ), .B(\GFM/N3097 ), .Z(\GFM/n16770 ) );
XOR2_X2 \GFM/U2735  ( .A(\GFM/N3093 ), .B(\GFM/N3094 ), .Z(\GFM/n16780 ) );
XOR2_X2 \GFM/U2734  ( .A(\GFM/N3089 ), .B(\GFM/N3090 ), .Z(\GFM/n1679 ) );
XOR2_X2 \GFM/U2733  ( .A(\GFM/N3085 ), .B(\GFM/N3087 ), .Z(\GFM/n1680 ) );
XOR2_X2 \GFM/U2732  ( .A(\GFM/N3080 ), .B(\GFM/N3084 ), .Z(\GFM/n16810 ) );
XOR2_X2 \GFM/U2731  ( .A(\GFM/N3077 ), .B(\GFM/N3079 ), .Z(\GFM/n16820 ) );
XOR2_X2 \GFM/U2730  ( .A(\GFM/N3073 ), .B(\GFM/N3076 ), .Z(\GFM/n1683 ) );
XOR2_X2 \GFM/U2729  ( .A(\GFM/N3070 ), .B(\GFM/N3072 ), .Z(\GFM/n16840 ) );
XOR2_X2 \GFM/U2728  ( .A(\GFM/n1686 ), .B(\GFM/n16850 ), .Z(z_out[100]) );
XOR2_X2 \GFM/U2727  ( .A(\GFM/n1688 ), .B(\GFM/n1687 ), .Z(\GFM/n16850 ) );
XOR2_X2 \GFM/U2726  ( .A(\GFM/n16900 ), .B(\GFM/n16890 ), .Z(\GFM/n1686 ) );
XOR2_X2 \GFM/U2725  ( .A(\GFM/n16920 ), .B(\GFM/n1691 ), .Z(\GFM/n1687 ) );
XOR2_X2 \GFM/U2724  ( .A(\GFM/n16940 ), .B(\GFM/n1693 ), .Z(\GFM/n1688 ) );
XOR2_X2 \GFM/U2723  ( .A(\GFM/n1696 ), .B(\GFM/n16950 ), .Z(\GFM/n16890 ) );
XOR2_X2 \GFM/U2722  ( .A(\GFM/n16980 ), .B(\GFM/n1697 ), .Z(\GFM/n16900 ) );
XOR2_X2 \GFM/U2721  ( .A(z_in[100]), .B(\GFM/n16990 ), .Z(\GFM/n1691 ) );
XOR2_X2 \GFM/U2720  ( .A(\GFM/N3127 ), .B(\GFM/N3128 ), .Z(\GFM/n16920 ) );
XOR2_X2 \GFM/U2719  ( .A(\GFM/N3124 ), .B(\GFM/N3125 ), .Z(\GFM/n1693 ) );
XOR2_X2 \GFM/U2718  ( .A(\GFM/N3120 ), .B(\GFM/N3121 ), .Z(\GFM/n16940 ) );
XOR2_X2 \GFM/U2717  ( .A(\GFM/N3116 ), .B(\GFM/N3118 ), .Z(\GFM/n16950 ) );
XOR2_X2 \GFM/U2716  ( .A(\GFM/N3111 ), .B(\GFM/N3115 ), .Z(\GFM/n1696 ) );
XOR2_X2 \GFM/U2715  ( .A(\GFM/N3108 ), .B(\GFM/N3110 ), .Z(\GFM/n1697 ) );
XOR2_X2 \GFM/U2714  ( .A(\GFM/N3104 ), .B(\GFM/N3107 ), .Z(\GFM/n16980 ) );
XOR2_X2 \GFM/U2713  ( .A(\GFM/N3101 ), .B(\GFM/N3103 ), .Z(\GFM/n16990 ) );
XOR2_X2 \GFM/U2712  ( .A(\GFM/n17010 ), .B(\GFM/n1700 ), .Z(z_out[101]) );
XOR2_X2 \GFM/U2711  ( .A(\GFM/n1703 ), .B(\GFM/n17020 ), .Z(\GFM/n1700 ) );
XOR2_X2 \GFM/U2710  ( .A(\GFM/n1705 ), .B(\GFM/n1704 ), .Z(\GFM/n17010 ) );
XOR2_X2 \GFM/U2709  ( .A(\GFM/n1707 ), .B(\GFM/n17060 ), .Z(\GFM/n17020 ) );
XOR2_X2 \GFM/U2708  ( .A(\GFM/n17090 ), .B(\GFM/n17080 ), .Z(\GFM/n1703 ) );
XOR2_X2 \GFM/U2707  ( .A(\GFM/n1711 ), .B(\GFM/n1710 ), .Z(\GFM/n1704 ) );
XOR2_X2 \GFM/U2706  ( .A(\GFM/n17130 ), .B(\GFM/n17120 ), .Z(\GFM/n1705 ) );
XOR2_X2 \GFM/U2705  ( .A(z_in[101]), .B(\GFM/n1714 ), .Z(\GFM/n17060 ) );
XOR2_X2 \GFM/U2704  ( .A(\GFM/N3158 ), .B(\GFM/N3159 ), .Z(\GFM/n1707 ) );
XOR2_X2 \GFM/U2703  ( .A(\GFM/N3155 ), .B(\GFM/N3156 ), .Z(\GFM/n17080 ) );
XOR2_X2 \GFM/U2702  ( .A(\GFM/N3151 ), .B(\GFM/N3152 ), .Z(\GFM/n17090 ) );
XOR2_X2 \GFM/U2701  ( .A(\GFM/N3147 ), .B(\GFM/N3149 ), .Z(\GFM/n1710 ) );
XOR2_X2 \GFM/U2700  ( .A(\GFM/N3142 ), .B(\GFM/N3146 ), .Z(\GFM/n1711 ) );
XOR2_X2 \GFM/U2699  ( .A(\GFM/N3139 ), .B(\GFM/N3141 ), .Z(\GFM/n17120 ) );
XOR2_X2 \GFM/U2698  ( .A(\GFM/N3135 ), .B(\GFM/N3138 ), .Z(\GFM/n17130 ) );
XOR2_X2 \GFM/U2697  ( .A(\GFM/N3132 ), .B(\GFM/N3134 ), .Z(\GFM/n1714 ) );
XOR2_X2 \GFM/U2696  ( .A(\GFM/n17160 ), .B(\GFM/n17150 ), .Z(z_out[102]) );
XOR2_X2 \GFM/U2695  ( .A(\GFM/n1718 ), .B(\GFM/n1717 ), .Z(\GFM/n17150 ) );
XOR2_X2 \GFM/U2694  ( .A(\GFM/n17200 ), .B(\GFM/n1719 ), .Z(\GFM/n17160 ) );
XOR2_X2 \GFM/U2693  ( .A(\GFM/n1722 ), .B(\GFM/n17210 ), .Z(\GFM/n1717 ) );
XOR2_X2 \GFM/U2692  ( .A(\GFM/n1724 ), .B(\GFM/n17230 ), .Z(\GFM/n1718 ) );
XOR2_X2 \GFM/U2691  ( .A(\GFM/n17260 ), .B(\GFM/n17250 ), .Z(\GFM/n1719 ) );
XOR2_X2 \GFM/U2690  ( .A(\GFM/n1728 ), .B(\GFM/n1727 ), .Z(\GFM/n17200 ) );
XOR2_X2 \GFM/U2689  ( .A(z_in[102]), .B(\GFM/n17290 ), .Z(\GFM/n17210 ) );
XOR2_X2 \GFM/U2688  ( .A(\GFM/N3189 ), .B(\GFM/N3190 ), .Z(\GFM/n1722 ) );
XOR2_X2 \GFM/U2687  ( .A(\GFM/N3186 ), .B(\GFM/N3187 ), .Z(\GFM/n17230 ) );
XOR2_X2 \GFM/U2686  ( .A(\GFM/N3182 ), .B(\GFM/N3183 ), .Z(\GFM/n1724 ) );
XOR2_X2 \GFM/U2685  ( .A(\GFM/N3178 ), .B(\GFM/N3180 ), .Z(\GFM/n17250 ) );
XOR2_X2 \GFM/U2684  ( .A(\GFM/N3173 ), .B(\GFM/N3177 ), .Z(\GFM/n17260 ) );
XOR2_X2 \GFM/U2683  ( .A(\GFM/N3170 ), .B(\GFM/N3172 ), .Z(\GFM/n1727 ) );
XOR2_X2 \GFM/U2682  ( .A(\GFM/N3166 ), .B(\GFM/N3169 ), .Z(\GFM/n1728 ) );
XOR2_X2 \GFM/U2681  ( .A(\GFM/N3163 ), .B(\GFM/N3165 ), .Z(\GFM/n17290 ) );
XOR2_X2 \GFM/U2680  ( .A(\GFM/n1731 ), .B(\GFM/n17300 ), .Z(z_out[103]) );
XOR2_X2 \GFM/U2679  ( .A(\GFM/n17330 ), .B(\GFM/n17320 ), .Z(\GFM/n17300 ));
XOR2_X2 \GFM/U2678  ( .A(\GFM/n1735 ), .B(\GFM/n1734 ), .Z(\GFM/n1731 ) );
XOR2_X2 \GFM/U2677  ( .A(\GFM/n17370 ), .B(\GFM/n1736 ), .Z(\GFM/n17320 ) );
XOR2_X2 \GFM/U2676  ( .A(\GFM/n17390 ), .B(\GFM/n1738 ), .Z(\GFM/n17330 ) );
XOR2_X2 \GFM/U2675  ( .A(\GFM/n1741 ), .B(\GFM/n17400 ), .Z(\GFM/n1734 ) );
XOR2_X2 \GFM/U2674  ( .A(\GFM/n17430 ), .B(\GFM/n1742 ), .Z(\GFM/n1735 ) );
XOR2_X2 \GFM/U2673  ( .A(z_in[103]), .B(\GFM/n17440 ), .Z(\GFM/n1736 ) );
XOR2_X2 \GFM/U2672  ( .A(\GFM/N3220 ), .B(\GFM/N3221 ), .Z(\GFM/n17370 ) );
XOR2_X2 \GFM/U2671  ( .A(\GFM/N3217 ), .B(\GFM/N3218 ), .Z(\GFM/n1738 ) );
XOR2_X2 \GFM/U2670  ( .A(\GFM/N3213 ), .B(\GFM/N3214 ), .Z(\GFM/n17390 ) );
XOR2_X2 \GFM/U2669  ( .A(\GFM/N3209 ), .B(\GFM/N3211 ), .Z(\GFM/n17400 ) );
XOR2_X2 \GFM/U2668  ( .A(\GFM/N3204 ), .B(\GFM/N3208 ), .Z(\GFM/n1741 ) );
XOR2_X2 \GFM/U2667  ( .A(\GFM/N3201 ), .B(\GFM/N3203 ), .Z(\GFM/n1742 ) );
XOR2_X2 \GFM/U2666  ( .A(\GFM/N3197 ), .B(\GFM/N3200 ), .Z(\GFM/n17430 ) );
XOR2_X2 \GFM/U2665  ( .A(\GFM/N3194 ), .B(\GFM/N3196 ), .Z(\GFM/n17440 ) );
XOR2_X2 \GFM/U2664  ( .A(\GFM/n17460 ), .B(\GFM/n1745 ), .Z(z_out[104]) );
XOR2_X2 \GFM/U2663  ( .A(\GFM/n1748 ), .B(\GFM/n17470 ), .Z(\GFM/n1745 ) );
XOR2_X2 \GFM/U2662  ( .A(\GFM/n1750 ), .B(\GFM/n1749 ), .Z(\GFM/n17460 ) );
XOR2_X2 \GFM/U2661  ( .A(\GFM/n17520 ), .B(\GFM/n17510 ), .Z(\GFM/n17470 ));
XOR2_X2 \GFM/U2660  ( .A(\GFM/n17540 ), .B(\GFM/n1753 ), .Z(\GFM/n1748 ) );
XOR2_X2 \GFM/U2659  ( .A(\GFM/n17560 ), .B(\GFM/n1755 ), .Z(\GFM/n1749 ) );
XOR2_X2 \GFM/U2658  ( .A(\GFM/n1758 ), .B(\GFM/n17570 ), .Z(\GFM/n1750 ) );
XOR2_X2 \GFM/U2657  ( .A(z_in[104]), .B(\GFM/n1759 ), .Z(\GFM/n17510 ) );
XOR2_X2 \GFM/U2656  ( .A(\GFM/N3251 ), .B(\GFM/N3252 ), .Z(\GFM/n17520 ) );
XOR2_X2 \GFM/U2655  ( .A(\GFM/N3248 ), .B(\GFM/N3249 ), .Z(\GFM/n1753 ) );
XOR2_X2 \GFM/U2654  ( .A(\GFM/N3244 ), .B(\GFM/N3245 ), .Z(\GFM/n17540 ) );
XOR2_X2 \GFM/U2653  ( .A(\GFM/N3240 ), .B(\GFM/N3242 ), .Z(\GFM/n1755 ) );
XOR2_X2 \GFM/U2652  ( .A(\GFM/N3235 ), .B(\GFM/N3239 ), .Z(\GFM/n17560 ) );
XOR2_X2 \GFM/U2651  ( .A(\GFM/N3232 ), .B(\GFM/N3234 ), .Z(\GFM/n17570 ) );
XOR2_X2 \GFM/U2650  ( .A(\GFM/N3228 ), .B(\GFM/N3231 ), .Z(\GFM/n1758 ) );
XOR2_X2 \GFM/U2649  ( .A(\GFM/N3225 ), .B(\GFM/N3227 ), .Z(\GFM/n1759 ) );
XOR2_X2 \GFM/U2648  ( .A(\GFM/n17610 ), .B(\GFM/n17600 ), .Z(z_out[105]) );
XOR2_X2 \GFM/U2647  ( .A(\GFM/n17630 ), .B(\GFM/n1762 ), .Z(\GFM/n17600 ) );
XOR2_X2 \GFM/U2646  ( .A(\GFM/n1765 ), .B(\GFM/n17640 ), .Z(\GFM/n17610 ) );
XOR2_X2 \GFM/U2645  ( .A(\GFM/n1767 ), .B(\GFM/n1766 ), .Z(\GFM/n1762 ) );
XOR2_X2 \GFM/U2644  ( .A(\GFM/n1769 ), .B(\GFM/n17680 ), .Z(\GFM/n17630 ) );
XOR2_X2 \GFM/U2643  ( .A(\GFM/n17710 ), .B(\GFM/n17700 ), .Z(\GFM/n17640 ));
XOR2_X2 \GFM/U2642  ( .A(\GFM/n1773 ), .B(\GFM/n1772 ), .Z(\GFM/n1765 ) );
XOR2_X2 \GFM/U2641  ( .A(z_in[105]), .B(\GFM/n17740 ), .Z(\GFM/n1766 ) );
XOR2_X2 \GFM/U2640  ( .A(\GFM/N3282 ), .B(\GFM/N3283 ), .Z(\GFM/n1767 ) );
XOR2_X2 \GFM/U2639  ( .A(\GFM/N3279 ), .B(\GFM/N3280 ), .Z(\GFM/n17680 ) );
XOR2_X2 \GFM/U2638  ( .A(\GFM/N3275 ), .B(\GFM/N3276 ), .Z(\GFM/n1769 ) );
XOR2_X2 \GFM/U2637  ( .A(\GFM/N3271 ), .B(\GFM/N3273 ), .Z(\GFM/n17700 ) );
XOR2_X2 \GFM/U2636  ( .A(\GFM/N3266 ), .B(\GFM/N3270 ), .Z(\GFM/n17710 ) );
XOR2_X2 \GFM/U2635  ( .A(\GFM/N3263 ), .B(\GFM/N3265 ), .Z(\GFM/n1772 ) );
XOR2_X2 \GFM/U2634  ( .A(\GFM/N3259 ), .B(\GFM/N3262 ), .Z(\GFM/n1773 ) );
XOR2_X2 \GFM/U2633  ( .A(\GFM/N3256 ), .B(\GFM/N3258 ), .Z(\GFM/n17740 ) );
XOR2_X2 \GFM/U2632  ( .A(\GFM/n1776 ), .B(\GFM/n17750 ), .Z(z_out[106]) );
XOR2_X2 \GFM/U2631  ( .A(\GFM/n17780 ), .B(\GFM/n17770 ), .Z(\GFM/n17750 ));
XOR2_X2 \GFM/U2630  ( .A(\GFM/n1780 ), .B(\GFM/n1779 ), .Z(\GFM/n1776 ) );
XOR2_X2 \GFM/U2629  ( .A(\GFM/n17820 ), .B(\GFM/n1781 ), .Z(\GFM/n17770 ) );
XOR2_X2 \GFM/U2628  ( .A(\GFM/n1784 ), .B(\GFM/n17830 ), .Z(\GFM/n17780 ) );
XOR2_X2 \GFM/U2627  ( .A(\GFM/n1786 ), .B(\GFM/n17850 ), .Z(\GFM/n1779 ) );
XOR2_X2 \GFM/U2626  ( .A(\GFM/n17880 ), .B(\GFM/n17870 ), .Z(\GFM/n1780 ) );
XOR2_X2 \GFM/U2625  ( .A(z_in[106]), .B(\GFM/n1789 ), .Z(\GFM/n1781 ) );
XOR2_X2 \GFM/U2624  ( .A(\GFM/N3313 ), .B(\GFM/N3316 ), .Z(\GFM/n17820 ) );
XOR2_X2 \GFM/U2623  ( .A(\GFM/N3309 ), .B(\GFM/N3312 ), .Z(\GFM/n17830 ) );
XOR2_X2 \GFM/U2622  ( .A(\GFM/N3306 ), .B(\GFM/N3308 ), .Z(\GFM/n1784 ) );
XOR2_X2 \GFM/U2621  ( .A(\GFM/N3303 ), .B(\GFM/N3304 ), .Z(\GFM/n17850 ) );
XOR2_X2 \GFM/U2620  ( .A(\GFM/N3298 ), .B(\GFM/N3299 ), .Z(\GFM/n1786 ) );
XOR2_X2 \GFM/U2619  ( .A(\GFM/N3294 ), .B(\GFM/N3296 ), .Z(\GFM/n17870 ) );
XOR2_X2 \GFM/U2618  ( .A(\GFM/N3290 ), .B(\GFM/N3293 ), .Z(\GFM/n17880 ) );
XOR2_X2 \GFM/U2617  ( .A(\GFM/N3287 ), .B(\GFM/N3289 ), .Z(\GFM/n1789 ) );
XOR2_X2 \GFM/U2616  ( .A(\GFM/n17910 ), .B(\GFM/n1790 ), .Z(z_out[107]) );
XOR2_X2 \GFM/U2615  ( .A(\GFM/n1793 ), .B(\GFM/n17920 ), .Z(\GFM/n1790 ) );
XOR2_X2 \GFM/U2614  ( .A(\GFM/n17950 ), .B(\GFM/n17940 ), .Z(\GFM/n17910 ));
XOR2_X2 \GFM/U2613  ( .A(\GFM/n1797 ), .B(\GFM/n1796 ), .Z(\GFM/n17920 ) );
XOR2_X2 \GFM/U2612  ( .A(\GFM/n17990 ), .B(\GFM/n1798 ), .Z(\GFM/n1793 ) );
XOR2_X2 \GFM/U2611  ( .A(\GFM/n18010 ), .B(\GFM/n1800 ), .Z(\GFM/n17940 ) );
XOR2_X2 \GFM/U2610  ( .A(\GFM/n1803 ), .B(\GFM/n18020 ), .Z(\GFM/n17950 ) );
XOR2_X2 \GFM/U2609  ( .A(z_in[107]), .B(\GFM/n1804 ), .Z(\GFM/n1796 ) );
XOR2_X2 \GFM/U2608  ( .A(\GFM/N3346 ), .B(\GFM/N3349 ), .Z(\GFM/n1797 ) );
XOR2_X2 \GFM/U2607  ( .A(\GFM/N3341 ), .B(\GFM/N3345 ), .Z(\GFM/n1798 ) );
XOR2_X2 \GFM/U2606  ( .A(\GFM/N3338 ), .B(\GFM/N3340 ), .Z(\GFM/n17990 ) );
XOR2_X2 \GFM/U2605  ( .A(\GFM/N3335 ), .B(\GFM/N3336 ), .Z(\GFM/n1800 ) );
XOR2_X2 \GFM/U2604  ( .A(\GFM/N3330 ), .B(\GFM/N3331 ), .Z(\GFM/n18010 ) );
XOR2_X2 \GFM/U2603  ( .A(\GFM/N3326 ), .B(\GFM/N3328 ), .Z(\GFM/n18020 ) );
XOR2_X2 \GFM/U2602  ( .A(\GFM/N3322 ), .B(\GFM/N3325 ), .Z(\GFM/n1803 ) );
XOR2_X2 \GFM/U2601  ( .A(\GFM/N3319 ), .B(\GFM/N3321 ), .Z(\GFM/n1804 ) );
XOR2_X2 \GFM/U2600  ( .A(\GFM/n18060 ), .B(\GFM/n18050 ), .Z(z_out[108]) );
XOR2_X2 \GFM/U2599  ( .A(\GFM/n18080 ), .B(\GFM/n1807 ), .Z(\GFM/n18050 ) );
XOR2_X2 \GFM/U2598  ( .A(\GFM/n1810 ), .B(\GFM/n18090 ), .Z(\GFM/n18060 ) );
XOR2_X2 \GFM/U2597  ( .A(\GFM/n1812 ), .B(\GFM/n1811 ), .Z(\GFM/n1807 ) );
XOR2_X2 \GFM/U2596  ( .A(\GFM/n18140 ), .B(\GFM/n18130 ), .Z(\GFM/n18080 ));
XOR2_X2 \GFM/U2595  ( .A(\GFM/n18160 ), .B(\GFM/n1815 ), .Z(\GFM/n18090 ) );
XOR2_X2 \GFM/U2594  ( .A(\GFM/n18180 ), .B(\GFM/n1817 ), .Z(\GFM/n1810 ) );
XOR2_X2 \GFM/U2593  ( .A(z_in[108]), .B(\GFM/n18190 ), .Z(\GFM/n1811 ) );
XOR2_X2 \GFM/U2592  ( .A(\GFM/N3380 ), .B(\GFM/N3383 ), .Z(\GFM/n1812 ) );
XOR2_X2 \GFM/U2591  ( .A(\GFM/N3374 ), .B(\GFM/N3378 ), .Z(\GFM/n18130 ) );
XOR2_X2 \GFM/U2590  ( .A(\GFM/N3371 ), .B(\GFM/N3373 ), .Z(\GFM/n18140 ) );
XOR2_X2 \GFM/U2589  ( .A(\GFM/N3368 ), .B(\GFM/N3369 ), .Z(\GFM/n1815 ) );
XOR2_X2 \GFM/U2588  ( .A(\GFM/N3363 ), .B(\GFM/N3364 ), .Z(\GFM/n18160 ) );
XOR2_X2 \GFM/U2587  ( .A(\GFM/N3359 ), .B(\GFM/N3361 ), .Z(\GFM/n1817 ) );
XOR2_X2 \GFM/U2586  ( .A(\GFM/N3355 ), .B(\GFM/N3358 ), .Z(\GFM/n18180 ) );
XOR2_X2 \GFM/U2585  ( .A(\GFM/N3352 ), .B(\GFM/N3354 ), .Z(\GFM/n18190 ) );
XOR2_X2 \GFM/U2584  ( .A(\GFM/n1821 ), .B(\GFM/n1820 ), .Z(z_out[109]) );
XOR2_X2 \GFM/U2583  ( .A(\GFM/n18230 ), .B(\GFM/n18220 ), .Z(\GFM/n1820 ) );
XOR2_X2 \GFM/U2582  ( .A(\GFM/n18250 ), .B(\GFM/n1824 ), .Z(\GFM/n1821 ) );
XOR2_X2 \GFM/U2581  ( .A(\GFM/n1827 ), .B(\GFM/n18260 ), .Z(\GFM/n18220 ) );
XOR2_X2 \GFM/U2580  ( .A(\GFM/n1829 ), .B(\GFM/n1828 ), .Z(\GFM/n18230 ) );
XOR2_X2 \GFM/U2579  ( .A(\GFM/n1831 ), .B(\GFM/n18300 ), .Z(\GFM/n1824 ) );
XOR2_X2 \GFM/U2578  ( .A(\GFM/n18330 ), .B(\GFM/n18320 ), .Z(\GFM/n18250 ));
XOR2_X2 \GFM/U2577  ( .A(z_in[109]), .B(\GFM/n1834 ), .Z(\GFM/n18260 ) );
XOR2_X2 \GFM/U2576  ( .A(\GFM/N3415 ), .B(\GFM/N3418 ), .Z(\GFM/n1827 ) );
XOR2_X2 \GFM/U2575  ( .A(\GFM/N3409 ), .B(\GFM/N3413 ), .Z(\GFM/n1828 ) );
XOR2_X2 \GFM/U2574  ( .A(\GFM/N3406 ), .B(\GFM/N3407 ), .Z(\GFM/n1829 ) );
XOR2_X2 \GFM/U2573  ( .A(\GFM/N3402 ), .B(\GFM/N3404 ), .Z(\GFM/n18300 ) );
XOR2_X2 \GFM/U2572  ( .A(\GFM/N3397 ), .B(\GFM/N3398 ), .Z(\GFM/n1831 ) );
XOR2_X2 \GFM/U2571  ( .A(\GFM/N3393 ), .B(\GFM/N3395 ), .Z(\GFM/n18320 ) );
XOR2_X2 \GFM/U2570  ( .A(\GFM/N3389 ), .B(\GFM/N3392 ), .Z(\GFM/n18330 ) );
XOR2_X2 \GFM/U2569  ( .A(\GFM/N3386 ), .B(\GFM/N3388 ), .Z(\GFM/n1834 ) );
XOR2_X2 \GFM/U2568  ( .A(\GFM/n18360 ), .B(\GFM/n1835 ), .Z(z_out[110]) );
XOR2_X2 \GFM/U2567  ( .A(\GFM/n1838 ), .B(\GFM/n18370 ), .Z(\GFM/n1835 ) );
XOR2_X2 \GFM/U2566  ( .A(\GFM/n18400 ), .B(\GFM/n18390 ), .Z(\GFM/n18360 ));
XOR2_X2 \GFM/U2565  ( .A(\GFM/n1842 ), .B(\GFM/n1841 ), .Z(\GFM/n18370 ) );
XOR2_X2 \GFM/U2564  ( .A(\GFM/n18440 ), .B(\GFM/n1843 ), .Z(\GFM/n1838 ) );
XOR2_X2 \GFM/U2563  ( .A(\GFM/n1846 ), .B(\GFM/n18450 ), .Z(\GFM/n18390 ) );
XOR2_X2 \GFM/U2562  ( .A(\GFM/n1848 ), .B(\GFM/n18470 ), .Z(\GFM/n18400 ) );
XOR2_X2 \GFM/U2561  ( .A(z_in[110]), .B(\GFM/n18490 ), .Z(\GFM/n1841 ) );
XOR2_X2 \GFM/U2560  ( .A(\GFM/N3452 ), .B(\GFM/N3455 ), .Z(\GFM/n1842 ) );
XOR2_X2 \GFM/U2559  ( .A(\GFM/N3446 ), .B(\GFM/N3450 ), .Z(\GFM/n1843 ) );
XOR2_X2 \GFM/U2558  ( .A(\GFM/N3443 ), .B(\GFM/N3444 ), .Z(\GFM/n18440 ) );
XOR2_X2 \GFM/U2557  ( .A(\GFM/N3439 ), .B(\GFM/N3441 ), .Z(\GFM/n18450 ) );
XOR2_X2 \GFM/U2556  ( .A(\GFM/N3433 ), .B(\GFM/N3434 ), .Z(\GFM/n1846 ) );
XOR2_X2 \GFM/U2555  ( .A(\GFM/N3429 ), .B(\GFM/N3431 ), .Z(\GFM/n18470 ) );
XOR2_X2 \GFM/U2554  ( .A(\GFM/N3425 ), .B(\GFM/N3428 ), .Z(\GFM/n1848 ) );
XOR2_X2 \GFM/U2553  ( .A(\GFM/N3422 ), .B(\GFM/N3424 ), .Z(\GFM/n18490 ) );
XOR2_X2 \GFM/U2552  ( .A(\GFM/n1851 ), .B(\GFM/n18500 ), .Z(z_out[111]) );
XOR2_X2 \GFM/U2551  ( .A(\GFM/n18530 ), .B(\GFM/n1852 ), .Z(\GFM/n18500 ) );
XOR2_X2 \GFM/U2550  ( .A(\GFM/n1855 ), .B(\GFM/n18540 ), .Z(\GFM/n1851 ) );
XOR2_X2 \GFM/U2549  ( .A(\GFM/n18570 ), .B(\GFM/n18560 ), .Z(\GFM/n1852 ) );
XOR2_X2 \GFM/U2548  ( .A(\GFM/n1859 ), .B(\GFM/n1858 ), .Z(\GFM/n18530 ) );
XOR2_X2 \GFM/U2547  ( .A(\GFM/n18610 ), .B(\GFM/n1860 ), .Z(\GFM/n18540 ) );
XOR2_X2 \GFM/U2546  ( .A(\GFM/n18630 ), .B(\GFM/n1862 ), .Z(\GFM/n1855 ) );
XOR2_X2 \GFM/U2545  ( .A(z_in[111]), .B(\GFM/n18640 ), .Z(\GFM/n18560 ) );
XOR2_X2 \GFM/U2544  ( .A(\GFM/N3491 ), .B(\GFM/N3495 ), .Z(\GFM/n18570 ) );
XOR2_X2 \GFM/U2543  ( .A(\GFM/N3484 ), .B(\GFM/N3489 ), .Z(\GFM/n1858 ) );
XOR2_X2 \GFM/U2542  ( .A(\GFM/N3482 ), .B(\GFM/N3483 ), .Z(\GFM/n1859 ) );
XOR2_X2 \GFM/U2541  ( .A(\GFM/N3477 ), .B(\GFM/N3479 ), .Z(\GFM/n1860 ) );
XOR2_X2 \GFM/U2540  ( .A(\GFM/N3471 ), .B(\GFM/N3472 ), .Z(\GFM/n18610 ) );
XOR2_X2 \GFM/U2539  ( .A(\GFM/N3467 ), .B(\GFM/N3469 ), .Z(\GFM/n1862 ) );
XOR2_X2 \GFM/U2538  ( .A(\GFM/N3463 ), .B(\GFM/N3466 ), .Z(\GFM/n18630 ) );
XOR2_X2 \GFM/U2537  ( .A(\GFM/N3460 ), .B(\GFM/N3462 ), .Z(\GFM/n18640 ) );
XOR2_X2 \GFM/U2536  ( .A(\GFM/n1866 ), .B(\GFM/n1865 ), .Z(z_out[112]) );
XOR2_X2 \GFM/U2535  ( .A(\GFM/n18680 ), .B(\GFM/n18670 ), .Z(\GFM/n1865 ) );
XOR2_X2 \GFM/U2534  ( .A(\GFM/n18700 ), .B(\GFM/n1869 ), .Z(\GFM/n1866 ) );
XOR2_X2 \GFM/U2533  ( .A(\GFM/n18721 ), .B(\GFM/n18710 ), .Z(\GFM/n18670 ));
XOR2_X2 \GFM/U2532  ( .A(\GFM/n1874 ), .B(\GFM/n1873 ), .Z(\GFM/n18680 ) );
XOR2_X2 \GFM/U2531  ( .A(\GFM/n18760 ), .B(\GFM/n18750 ), .Z(\GFM/n1869 ) );
XOR2_X2 \GFM/U2530  ( .A(\GFM/n18780 ), .B(\GFM/n1877 ), .Z(\GFM/n18700 ) );
XOR2_X2 \GFM/U2529  ( .A(z_in[112]), .B(\GFM/n1879 ), .Z(\GFM/n18710 ) );
XOR2_X2 \GFM/U2528  ( .A(\GFM/N3534 ), .B(\GFM/N3538 ), .Z(\GFM/n18721 ) );
XOR2_X2 \GFM/U2527  ( .A(\GFM/N3527 ), .B(\GFM/N3529 ), .Z(\GFM/n1873 ) );
XOR2_X2 \GFM/U2526  ( .A(\GFM/N3521 ), .B(\GFM/N3524 ), .Z(\GFM/n1874 ) );
XOR2_X2 \GFM/U2525  ( .A(\GFM/N3514 ), .B(\GFM/N3519 ), .Z(\GFM/n18750 ) );
XOR2_X2 \GFM/U2524  ( .A(\GFM/N3511 ), .B(\GFM/N3513 ), .Z(\GFM/n18760 ) );
XOR2_X2 \GFM/U2523  ( .A(\GFM/N3508 ), .B(\GFM/N3509 ), .Z(\GFM/n1877 ) );
XOR2_X2 \GFM/U2522  ( .A(\GFM/N3503 ), .B(\GFM/N3505 ), .Z(\GFM/n18780 ) );
XOR2_X2 \GFM/U2521  ( .A(\GFM/N3500 ), .B(\GFM/N3502 ), .Z(\GFM/n1879 ) );
XOR2_X2 \GFM/U2520  ( .A(\GFM/n18810 ), .B(\GFM/n18800 ), .Z(z_out[113]) );
XOR2_X2 \GFM/U2519  ( .A(\GFM/n1883 ), .B(\GFM/n1882 ), .Z(\GFM/n18800 ) );
XOR2_X2 \GFM/U2518  ( .A(\GFM/n18850 ), .B(\GFM/n18840 ), .Z(\GFM/n18810 ));
XOR2_X2 \GFM/U2517  ( .A(\GFM/n18870 ), .B(\GFM/n1886 ), .Z(\GFM/n1882 ) );
XOR2_X2 \GFM/U2516  ( .A(\GFM/n1889 ), .B(\GFM/n18880 ), .Z(\GFM/n1883 ) );
XOR2_X2 \GFM/U2515  ( .A(\GFM/n1891 ), .B(\GFM/n18901 ), .Z(\GFM/n18840 ) );
XOR2_X2 \GFM/U2514  ( .A(\GFM/n1893 ), .B(\GFM/n18920 ), .Z(\GFM/n18850 ) );
XOR2_X2 \GFM/U2513  ( .A(z_in[113]), .B(\GFM/n18940 ), .Z(\GFM/n1886 ) );
XOR2_X2 \GFM/U2512  ( .A(\GFM/N3580 ), .B(\GFM/N3584 ), .Z(\GFM/n18870 ) );
XOR2_X2 \GFM/U2511  ( .A(\GFM/N3571 ), .B(\GFM/N3574 ), .Z(\GFM/n18880 ) );
XOR2_X2 \GFM/U2510  ( .A(\GFM/N3566 ), .B(\GFM/N3569 ), .Z(\GFM/n1889 ) );
XOR2_X2 \GFM/U2509  ( .A(\GFM/N3558 ), .B(\GFM/N3563 ), .Z(\GFM/n18901 ) );
XOR2_X2 \GFM/U2508  ( .A(\GFM/N3554 ), .B(\GFM/N3556 ), .Z(\GFM/n1891 ) );
XOR2_X2 \GFM/U2507  ( .A(\GFM/N3551 ), .B(\GFM/N3552 ), .Z(\GFM/n18920 ) );
XOR2_X2 \GFM/U2506  ( .A(\GFM/N3546 ), .B(\GFM/N3548 ), .Z(\GFM/n1893 ) );
XOR2_X2 \GFM/U2505  ( .A(\GFM/N3543 ), .B(\GFM/N3545 ), .Z(\GFM/n18940 ) );
XOR2_X2 \GFM/U2504  ( .A(\GFM/n1896 ), .B(\GFM/n18950 ), .Z(z_out[114]) );
XOR2_X2 \GFM/U2503  ( .A(\GFM/n18980 ), .B(\GFM/n1897 ), .Z(\GFM/n18950 ) );
XOR2_X2 \GFM/U2502  ( .A(\GFM/n19001 ), .B(\GFM/n18990 ), .Z(\GFM/n1896 ) );
XOR2_X2 \GFM/U2501  ( .A(\GFM/n19020 ), .B(\GFM/n19010 ), .Z(\GFM/n1897 ) );
XOR2_X2 \GFM/U2500  ( .A(\GFM/n1904 ), .B(\GFM/n1903 ), .Z(\GFM/n18980 ) );
XOR2_X2 \GFM/U2499  ( .A(\GFM/n19060 ), .B(\GFM/n1905 ), .Z(\GFM/n18990 ) );
XOR2_X2 \GFM/U2498  ( .A(\GFM/n1908 ), .B(\GFM/n19070 ), .Z(\GFM/n19001 ) );
XOR2_X2 \GFM/U2497  ( .A(z_in[114]), .B(\GFM/n19090 ), .Z(\GFM/n19010 ) );
XOR2_X2 \GFM/U2496  ( .A(\GFM/N3629 ), .B(\GFM/N3633 ), .Z(\GFM/n19020 ) );
XOR2_X2 \GFM/U2495  ( .A(\GFM/N3620 ), .B(\GFM/N3623 ), .Z(\GFM/n1903 ) );
XOR2_X2 \GFM/U2494  ( .A(\GFM/N3615 ), .B(\GFM/N3618 ), .Z(\GFM/n1904 ) );
XOR2_X2 \GFM/U2493  ( .A(\GFM/N3605 ), .B(\GFM/N3611 ), .Z(\GFM/n1905 ) );
XOR2_X2 \GFM/U2492  ( .A(\GFM/N3600 ), .B(\GFM/N3603 ), .Z(\GFM/n19060 ) );
XOR2_X2 \GFM/U2491  ( .A(\GFM/N3597 ), .B(\GFM/N3598 ), .Z(\GFM/n19070 ) );
XOR2_X2 \GFM/U2490  ( .A(\GFM/N3592 ), .B(\GFM/N3594 ), .Z(\GFM/n1908 ) );
XOR2_X2 \GFM/U2489  ( .A(\GFM/N3589 ), .B(\GFM/N3591 ), .Z(\GFM/n19090 ) );
XOR2_X2 \GFM/U2488  ( .A(\GFM/n19110 ), .B(\GFM/n1910 ), .Z(z_out[115]) );
XOR2_X2 \GFM/U2487  ( .A(\GFM/n1913 ), .B(\GFM/n19120 ), .Z(\GFM/n1910 ) );
XOR2_X2 \GFM/U2486  ( .A(\GFM/n19150 ), .B(\GFM/n1914 ), .Z(\GFM/n19110 ) );
XOR2_X2 \GFM/U2485  ( .A(\GFM/n1917 ), .B(\GFM/n19160 ), .Z(\GFM/n19120 ) );
XOR2_X2 \GFM/U2484  ( .A(\GFM/n19190 ), .B(\GFM/n19180 ), .Z(\GFM/n1913 ) );
XOR2_X2 \GFM/U2483  ( .A(\GFM/n1921 ), .B(\GFM/n1920 ), .Z(\GFM/n1914 ) );
XOR2_X2 \GFM/U2482  ( .A(\GFM/n19230 ), .B(\GFM/n1922 ), .Z(\GFM/n19150 ) );
XOR2_X2 \GFM/U2481  ( .A(z_in[115]), .B(\GFM/n1924 ), .Z(\GFM/n19160 ) );
XOR2_X2 \GFM/U2480  ( .A(\GFM/N3681 ), .B(\GFM/N3685 ), .Z(\GFM/n1917 ) );
XOR2_X2 \GFM/U2479  ( .A(\GFM/N3672 ), .B(\GFM/N3674 ), .Z(\GFM/n19180 ) );
XOR2_X2 \GFM/U2478  ( .A(\GFM/N3666 ), .B(\GFM/N3670 ), .Z(\GFM/n19190 ) );
XOR2_X2 \GFM/U2477  ( .A(\GFM/N3655 ), .B(\GFM/N3662 ), .Z(\GFM/n1920 ) );
XOR2_X2 \GFM/U2476  ( .A(\GFM/N3649 ), .B(\GFM/N3653 ), .Z(\GFM/n1921 ) );
XOR2_X2 \GFM/U2475  ( .A(\GFM/N3647 ), .B(\GFM/N3648 ), .Z(\GFM/n1922 ) );
XOR2_X2 \GFM/U2474  ( .A(\GFM/N3641 ), .B(\GFM/N3643 ), .Z(\GFM/n19230 ) );
XOR2_X2 \GFM/U2473  ( .A(\GFM/N3638 ), .B(\GFM/N3640 ), .Z(\GFM/n1924 ) );
XOR2_X2 \GFM/U2472  ( .A(\GFM/n19260 ), .B(\GFM/n19250 ), .Z(z_out[116]) );
XOR2_X2 \GFM/U2471  ( .A(\GFM/n1928 ), .B(\GFM/n1927 ), .Z(\GFM/n19250 ) );
XOR2_X2 \GFM/U2470  ( .A(\GFM/n19300 ), .B(\GFM/n19290 ), .Z(\GFM/n19260 ));
XOR2_X2 \GFM/U2469  ( .A(\GFM/n19320 ), .B(\GFM/n19311 ), .Z(\GFM/n1927 ) );
XOR2_X2 \GFM/U2468  ( .A(\GFM/n1934 ), .B(\GFM/n19330 ), .Z(\GFM/n1928 ) );
XOR2_X2 \GFM/U2467  ( .A(\GFM/n1936 ), .B(\GFM/n1935 ), .Z(\GFM/n19290 ) );
XOR2_X2 \GFM/U2466  ( .A(\GFM/n19380 ), .B(\GFM/n19370 ), .Z(\GFM/n19300 ));
XOR2_X2 \GFM/U2465  ( .A(z_in[116]), .B(\GFM/n1939 ), .Z(\GFM/n19311 ) );
XOR2_X2 \GFM/U2464  ( .A(\GFM/N3735 ), .B(\GFM/N3740 ), .Z(\GFM/n19320 ) );
XOR2_X2 \GFM/U2463  ( .A(\GFM/N3725 ), .B(\GFM/N3731 ), .Z(\GFM/n19330 ) );
XOR2_X2 \GFM/U2462  ( .A(\GFM/N3719 ), .B(\GFM/N3723 ), .Z(\GFM/n1934 ) );
XOR2_X2 \GFM/U2461  ( .A(\GFM/N3708 ), .B(\GFM/N3715 ), .Z(\GFM/n1935 ) );
XOR2_X2 \GFM/U2460  ( .A(\GFM/N3703 ), .B(\GFM/N3706 ), .Z(\GFM/n1936 ) );
XOR2_X2 \GFM/U2459  ( .A(\GFM/N3699 ), .B(\GFM/N3701 ), .Z(\GFM/n19370 ) );
XOR2_X2 \GFM/U2458  ( .A(\GFM/N3693 ), .B(\GFM/N3695 ), .Z(\GFM/n19380 ) );
XOR2_X2 \GFM/U2457  ( .A(\GFM/N3690 ), .B(\GFM/N3692 ), .Z(\GFM/n1939 ) );
XOR2_X2 \GFM/U2456  ( .A(\GFM/n19411 ), .B(\GFM/n19400 ), .Z(z_out[117]) );
XOR2_X2 \GFM/U2455  ( .A(\GFM/n19430 ), .B(\GFM/n19420 ), .Z(\GFM/n19400 ));
XOR2_X2 \GFM/U2454  ( .A(\GFM/n1945 ), .B(\GFM/n1944 ), .Z(\GFM/n19411 ) );
XOR2_X2 \GFM/U2453  ( .A(\GFM/n19470 ), .B(\GFM/n19460 ), .Z(\GFM/n19420 ));
XOR2_X2 \GFM/U2452  ( .A(\GFM/n19490 ), .B(\GFM/n1948 ), .Z(\GFM/n19430 ) );
XOR2_X2 \GFM/U2451  ( .A(\GFM/n1951 ), .B(\GFM/n19500 ), .Z(\GFM/n1944 ) );
XOR2_X2 \GFM/U2450  ( .A(\GFM/n1953 ), .B(\GFM/n1952 ), .Z(\GFM/n1945 ) );
XOR2_X2 \GFM/U2449  ( .A(z_in[117]), .B(\GFM/n19540 ), .Z(\GFM/n19460 ) );
XOR2_X2 \GFM/U2448  ( .A(\GFM/N3793 ), .B(\GFM/N3798 ), .Z(\GFM/n19470 ) );
XOR2_X2 \GFM/U2447  ( .A(\GFM/N3783 ), .B(\GFM/N3789 ), .Z(\GFM/n1948 ) );
XOR2_X2 \GFM/U2446  ( .A(\GFM/N3775 ), .B(\GFM/N3780 ), .Z(\GFM/n19490 ) );
XOR2_X2 \GFM/U2445  ( .A(\GFM/N3764 ), .B(\GFM/N3771 ), .Z(\GFM/n19500 ) );
XOR2_X2 \GFM/U2444  ( .A(\GFM/N3759 ), .B(\GFM/N3762 ), .Z(\GFM/n1951 ) );
XOR2_X2 \GFM/U2443  ( .A(\GFM/N3754 ), .B(\GFM/N3756 ), .Z(\GFM/n1952 ) );
XOR2_X2 \GFM/U2442  ( .A(\GFM/N3748 ), .B(\GFM/N3750 ), .Z(\GFM/n1953 ) );
XOR2_X2 \GFM/U2441  ( .A(\GFM/N3745 ), .B(\GFM/N3747 ), .Z(\GFM/n19540 ) );
XOR2_X2 \GFM/U2440  ( .A(\GFM/n19560 ), .B(\GFM/n1955 ), .Z(z_out[118]) );
XOR2_X2 \GFM/U2439  ( .A(\GFM/n1958 ), .B(\GFM/n19570 ), .Z(\GFM/n1955 ) );
XOR2_X2 \GFM/U2438  ( .A(\GFM/n19600 ), .B(\GFM/n1959 ), .Z(\GFM/n19560 ) );
XOR2_X2 \GFM/U2437  ( .A(\GFM/n19621 ), .B(\GFM/n19610 ), .Z(\GFM/n19570 ));
XOR2_X2 \GFM/U2436  ( .A(\GFM/n19640 ), .B(\GFM/n19630 ), .Z(\GFM/n1958 ) );
XOR2_X2 \GFM/U2435  ( .A(\GFM/n1966 ), .B(\GFM/n1965 ), .Z(\GFM/n1959 ) );
XOR2_X2 \GFM/U2434  ( .A(\GFM/n19680 ), .B(\GFM/n1967 ), .Z(\GFM/n19600 ) );
XOR2_X2 \GFM/U2433  ( .A(z_in[118]), .B(\GFM/n19690 ), .Z(\GFM/n19610 ) );
XOR2_X2 \GFM/U2432  ( .A(\GFM/N3854 ), .B(\GFM/N3859 ), .Z(\GFM/n19621 ) );
XOR2_X2 \GFM/U2431  ( .A(\GFM/N3844 ), .B(\GFM/N3850 ), .Z(\GFM/n19630 ) );
XOR2_X2 \GFM/U2430  ( .A(\GFM/N3835 ), .B(\GFM/N3840 ), .Z(\GFM/n19640 ) );
XOR2_X2 \GFM/U2429  ( .A(\GFM/N3825 ), .B(\GFM/N3831 ), .Z(\GFM/n1965 ) );
XOR2_X2 \GFM/U2428  ( .A(\GFM/N3818 ), .B(\GFM/N3821 ), .Z(\GFM/n1966 ) );
XOR2_X2 \GFM/U2427  ( .A(\GFM/N3812 ), .B(\GFM/N3816 ), .Z(\GFM/n1967 ) );
XOR2_X2 \GFM/U2426  ( .A(\GFM/N3808 ), .B(\GFM/N3809 ), .Z(\GFM/n19680 ) );
XOR2_X2 \GFM/U2425  ( .A(\GFM/N3803 ), .B(\GFM/N3804 ), .Z(\GFM/n19690 ) );
XOR2_X2 \GFM/U2424  ( .A(\GFM/n19710 ), .B(\GFM/n19701 ), .Z(z_out[119]) );
XOR2_X2 \GFM/U2423  ( .A(\GFM/n19730 ), .B(\GFM/n1972 ), .Z(\GFM/n19701 ) );
XOR2_X2 \GFM/U2422  ( .A(\GFM/n1975 ), .B(\GFM/n19740 ), .Z(\GFM/n19710 ) );
XOR2_X2 \GFM/U2421  ( .A(\GFM/n19770 ), .B(\GFM/n1976 ), .Z(\GFM/n1972 ) );
XOR2_X2 \GFM/U2420  ( .A(\GFM/n1979 ), .B(\GFM/n19780 ), .Z(\GFM/n19730 ) );
XOR2_X2 \GFM/U2419  ( .A(\GFM/n19810 ), .B(\GFM/n19800 ), .Z(\GFM/n19740 ));
XOR2_X2 \GFM/U2418  ( .A(\GFM/n1983 ), .B(\GFM/n1982 ), .Z(\GFM/n1975 ) );
XOR2_X2 \GFM/U2417  ( .A(z_in[119]), .B(\GFM/n1984 ), .Z(\GFM/n1976 ) );
XOR2_X2 \GFM/U2416  ( .A(\GFM/N3918 ), .B(\GFM/N3923 ), .Z(\GFM/n19770 ) );
XOR2_X2 \GFM/U2415  ( .A(\GFM/N3908 ), .B(\GFM/N3914 ), .Z(\GFM/n19780 ) );
XOR2_X2 \GFM/U2414  ( .A(\GFM/N3899 ), .B(\GFM/N3904 ), .Z(\GFM/n1979 ) );
XOR2_X2 \GFM/U2413  ( .A(\GFM/N3889 ), .B(\GFM/N3895 ), .Z(\GFM/n19800 ) );
XOR2_X2 \GFM/U2412  ( .A(\GFM/N3881 ), .B(\GFM/N3883 ), .Z(\GFM/n19810 ) );
XOR2_X2 \GFM/U2411  ( .A(\GFM/N3874 ), .B(\GFM/N3879 ), .Z(\GFM/n1982 ) );
XOR2_X2 \GFM/U2410  ( .A(\GFM/N3869 ), .B(\GFM/N3871 ), .Z(\GFM/n1983 ) );
XOR2_X2 \GFM/U2409  ( .A(\GFM/N3864 ), .B(\GFM/N3865 ), .Z(\GFM/n1984 ) );
XOR2_X2 \GFM/U2408  ( .A(\GFM/n1986 ), .B(\GFM/n19850 ), .Z(z_out[120]) );
XOR2_X2 \GFM/U2407  ( .A(\GFM/n19880 ), .B(\GFM/n19870 ), .Z(\GFM/n19850 ));
XOR2_X2 \GFM/U2406  ( .A(\GFM/n1990 ), .B(\GFM/n1989 ), .Z(\GFM/n1986 ) );
XOR2_X2 \GFM/U2405  ( .A(\GFM/n19920 ), .B(\GFM/n19910 ), .Z(\GFM/n19870 ));
XOR2_X2 \GFM/U2404  ( .A(\GFM/n19940 ), .B(\GFM/n1993 ), .Z(\GFM/n19880 ) );
XOR2_X2 \GFM/U2403  ( .A(\GFM/n1996 ), .B(\GFM/n19950 ), .Z(\GFM/n1989 ) );
XOR2_X2 \GFM/U2402  ( .A(\GFM/n1998 ), .B(\GFM/n1997 ), .Z(\GFM/n1990 ) );
XOR2_X2 \GFM/U2401  ( .A(z_in[120]), .B(\GFM/n19990 ), .Z(\GFM/n19910 ) );
XOR2_X2 \GFM/U2400  ( .A(\GFM/N3985 ), .B(\GFM/N3990 ), .Z(\GFM/n19920 ) );
XOR2_X2 \GFM/U2399  ( .A(\GFM/N3975 ), .B(\GFM/N3981 ), .Z(\GFM/n1993 ) );
XOR2_X2 \GFM/U2398  ( .A(\GFM/N3966 ), .B(\GFM/N3971 ), .Z(\GFM/n19940 ) );
XOR2_X2 \GFM/U2397  ( .A(\GFM/N3955 ), .B(\GFM/N3962 ), .Z(\GFM/n19950 ) );
XOR2_X2 \GFM/U2396  ( .A(\GFM/N3946 ), .B(\GFM/N3951 ), .Z(\GFM/n1996 ) );
XOR2_X2 \GFM/U2395  ( .A(\GFM/N3939 ), .B(\GFM/N3944 ), .Z(\GFM/n1997 ) );
XOR2_X2 \GFM/U2394  ( .A(\GFM/N3934 ), .B(\GFM/N3936 ), .Z(\GFM/n1998 ) );
XOR2_X2 \GFM/U2393  ( .A(\GFM/N3928 ), .B(\GFM/N3931 ), .Z(\GFM/n19990 ) );
XOR2_X2 \GFM/U2392  ( .A(\GFM/n2001 ), .B(\GFM/n20000 ), .Z(z_out[121]) );
XOR2_X2 \GFM/U2391  ( .A(\GFM/n2003 ), .B(\GFM/n20020 ), .Z(\GFM/n20000 ) );
XOR2_X2 \GFM/U2390  ( .A(\GFM/n20050 ), .B(\GFM/n20040 ), .Z(\GFM/n2001 ) );
XOR2_X2 \GFM/U2389  ( .A(\GFM/n2007 ), .B(\GFM/n2006 ), .Z(\GFM/n20020 ) );
XOR2_X2 \GFM/U2388  ( .A(\GFM/n20090 ), .B(\GFM/n20080 ), .Z(\GFM/n2003 ) );
XOR2_X2 \GFM/U2387  ( .A(\GFM/n20110 ), .B(\GFM/n20101 ), .Z(\GFM/n20040 ));
XOR2_X2 \GFM/U2386  ( .A(\GFM/n2013 ), .B(\GFM/n20120 ), .Z(\GFM/n20050 ) );
XOR2_X2 \GFM/U2385  ( .A(z_in[121]), .B(\GFM/n2014 ), .Z(\GFM/n2006 ) );
XOR2_X2 \GFM/U2384  ( .A(\GFM/N4039 ), .B(\GFM/N4042 ), .Z(\GFM/n2007 ) );
XOR2_X2 \GFM/U2383  ( .A(\GFM/N4032 ), .B(\GFM/N4035 ), .Z(\GFM/n20080 ) );
XOR2_X2 \GFM/U2382  ( .A(\GFM/N4024 ), .B(\GFM/N4027 ), .Z(\GFM/n20090 ) );
XOR2_X2 \GFM/U2381  ( .A(\GFM/N4017 ), .B(\GFM/N4020 ), .Z(\GFM/n20101 ) );
XOR2_X2 \GFM/U2380  ( .A(\GFM/N4007 ), .B(\GFM/N4012 ), .Z(\GFM/n20110 ) );
XOR2_X2 \GFM/U2379  ( .A(\GFM/N4004 ), .B(\GFM/N4006 ), .Z(\GFM/n20120 ) );
XOR2_X2 \GFM/U2378  ( .A(\GFM/N3997 ), .B(\GFM/N3999 ), .Z(\GFM/n2013 ) );
XOR2_X2 \GFM/U2377  ( .A(\GFM/N3994 ), .B(\GFM/N3996 ), .Z(\GFM/n2014 ) );
XOR2_X2 \GFM/U2376  ( .A(\GFM/n20160 ), .B(\GFM/n2015 ), .Z(z_out[122]) );
XOR2_X2 \GFM/U2375  ( .A(\GFM/n20180 ), .B(\GFM/n2017 ), .Z(\GFM/n2015 ) );
XOR2_X2 \GFM/U2374  ( .A(\GFM/n20201 ), .B(\GFM/n20190 ), .Z(\GFM/n20160 ));
XOR2_X2 \GFM/U2373  ( .A(\GFM/n20220 ), .B(\GFM/n2021 ), .Z(\GFM/n2017 ) );
XOR2_X2 \GFM/U2372  ( .A(\GFM/n2024 ), .B(\GFM/n20230 ), .Z(\GFM/n20180 ) );
XOR2_X2 \GFM/U2371  ( .A(\GFM/n20260 ), .B(\GFM/n20250 ), .Z(\GFM/n20190 ));
XOR2_X2 \GFM/U2370  ( .A(\GFM/n2028 ), .B(\GFM/n2027 ), .Z(\GFM/n20201 ) );
XOR2_X2 \GFM/U2369  ( .A(z_in[122]), .B(\GFM/n2029 ), .Z(\GFM/n2021 ) );
XOR2_X2 \GFM/U2368  ( .A(\GFM/N4094 ), .B(\GFM/N4097 ), .Z(\GFM/n20220 ) );
XOR2_X2 \GFM/U2367  ( .A(\GFM/N4087 ), .B(\GFM/N4090 ), .Z(\GFM/n20230 ) );
XOR2_X2 \GFM/U2366  ( .A(\GFM/N4079 ), .B(\GFM/N4082 ), .Z(\GFM/n2024 ) );
XOR2_X2 \GFM/U2365  ( .A(\GFM/N4072 ), .B(\GFM/N4075 ), .Z(\GFM/n20250 ) );
XOR2_X2 \GFM/U2364  ( .A(\GFM/N4063 ), .B(\GFM/N4066 ), .Z(\GFM/n20260 ) );
XOR2_X2 \GFM/U2363  ( .A(\GFM/N4057 ), .B(\GFM/N4059 ), .Z(\GFM/n2027 ) );
XOR2_X2 \GFM/U2362  ( .A(\GFM/N4050 ), .B(\GFM/N4052 ), .Z(\GFM/n2028 ) );
XOR2_X2 \GFM/U2361  ( .A(\GFM/N4047 ), .B(\GFM/N4049 ), .Z(\GFM/n2029 ) );
XOR2_X2 \GFM/U2360  ( .A(\GFM/n20310 ), .B(\GFM/n20300 ), .Z(z_out[123]) );
XOR2_X2 \GFM/U2359  ( .A(\GFM/n20330 ), .B(\GFM/n2032 ), .Z(\GFM/n20300 ) );
XOR2_X2 \GFM/U2358  ( .A(\GFM/n20350 ), .B(\GFM/n2034 ), .Z(\GFM/n20310 ) );
XOR2_X2 \GFM/U2357  ( .A(\GFM/n2037 ), .B(\GFM/n20360 ), .Z(\GFM/n2032 ) );
XOR2_X2 \GFM/U2356  ( .A(\GFM/n20390 ), .B(\GFM/n2038 ), .Z(\GFM/n20330 ) );
XOR2_X2 \GFM/U2355  ( .A(\GFM/n20411 ), .B(\GFM/n20400 ), .Z(\GFM/n2034 ) );
XOR2_X2 \GFM/U2354  ( .A(\GFM/n20430 ), .B(\GFM/n20420 ), .Z(\GFM/n20350 ));
XOR2_X2 \GFM/U2353  ( .A(z_in[123]), .B(\GFM/n2044 ), .Z(\GFM/n20360 ) );
XOR2_X2 \GFM/U2352  ( .A(\GFM/N4151 ), .B(\GFM/N4154 ), .Z(\GFM/n2037 ) );
XOR2_X2 \GFM/U2351  ( .A(\GFM/N4144 ), .B(\GFM/N4147 ), .Z(\GFM/n2038 ) );
XOR2_X2 \GFM/U2350  ( .A(\GFM/N4136 ), .B(\GFM/N4139 ), .Z(\GFM/n20390 ) );
XOR2_X2 \GFM/U2349  ( .A(\GFM/N4129 ), .B(\GFM/N4132 ), .Z(\GFM/n20400 ) );
XOR2_X2 \GFM/U2348  ( .A(\GFM/N4120 ), .B(\GFM/N4123 ), .Z(\GFM/n20411 ) );
XOR2_X2 \GFM/U2347  ( .A(\GFM/N4113 ), .B(\GFM/N4116 ), .Z(\GFM/n20420 ) );
XOR2_X2 \GFM/U2346  ( .A(\GFM/N4106 ), .B(\GFM/N4108 ), .Z(\GFM/n20430 ) );
XOR2_X2 \GFM/U2345  ( .A(\GFM/N4102 ), .B(\GFM/N4103 ), .Z(\GFM/n2044 ) );
XOR2_X2 \GFM/U2344  ( .A(\GFM/n2046 ), .B(\GFM/n2045 ), .Z(z_out[124]) );
XOR2_X2 \GFM/U2343  ( .A(\GFM/n2048 ), .B(\GFM/n20470 ), .Z(\GFM/n2045 ) );
XOR2_X2 \GFM/U2342  ( .A(\GFM/n20500 ), .B(\GFM/n20490 ), .Z(\GFM/n2046 ) );
XOR2_X2 \GFM/U2341  ( .A(\GFM/n2052 ), .B(\GFM/n2051 ), .Z(\GFM/n20470 ) );
XOR2_X2 \GFM/U2340  ( .A(\GFM/n20540 ), .B(\GFM/n20530 ), .Z(\GFM/n2048 ) );
XOR2_X2 \GFM/U2339  ( .A(\GFM/n20560 ), .B(\GFM/n2055 ), .Z(\GFM/n20490 ) );
XOR2_X2 \GFM/U2338  ( .A(\GFM/n2058 ), .B(\GFM/n20570 ), .Z(\GFM/n20500 ) );
XOR2_X2 \GFM/U2337  ( .A(z_in[124]), .B(\GFM/n2059 ), .Z(\GFM/n2051 ) );
XOR2_X2 \GFM/U2336  ( .A(\GFM/N4210 ), .B(\GFM/N4213 ), .Z(\GFM/n2052 ) );
XOR2_X2 \GFM/U2335  ( .A(\GFM/N4203 ), .B(\GFM/N4206 ), .Z(\GFM/n20530 ) );
XOR2_X2 \GFM/U2334  ( .A(\GFM/N4195 ), .B(\GFM/N4198 ), .Z(\GFM/n20540 ) );
XOR2_X2 \GFM/U2333  ( .A(\GFM/N4188 ), .B(\GFM/N4191 ), .Z(\GFM/n2055 ) );
XOR2_X2 \GFM/U2332  ( .A(\GFM/N4179 ), .B(\GFM/N4182 ), .Z(\GFM/n20560 ) );
XOR2_X2 \GFM/U2331  ( .A(\GFM/N4172 ), .B(\GFM/N4175 ), .Z(\GFM/n20570 ) );
XOR2_X2 \GFM/U2330  ( .A(\GFM/N4164 ), .B(\GFM/N4167 ), .Z(\GFM/n2058 ) );
XOR2_X2 \GFM/U2329  ( .A(\GFM/N4159 ), .B(\GFM/N4160 ), .Z(\GFM/n2059 ) );
XOR2_X2 \GFM/U2328  ( .A(\GFM/n20610 ), .B(\GFM/n20601 ), .Z(z_out[125]) );
XOR2_X2 \GFM/U2327  ( .A(\GFM/n2063 ), .B(\GFM/n20620 ), .Z(\GFM/n20601 ) );
XOR2_X2 \GFM/U2326  ( .A(\GFM/n2065 ), .B(\GFM/n20640 ), .Z(\GFM/n20610 ) );
XOR2_X2 \GFM/U2325  ( .A(\GFM/n20670 ), .B(\GFM/n20660 ), .Z(\GFM/n20620 ));
XOR2_X2 \GFM/U2324  ( .A(\GFM/n2069 ), .B(\GFM/n2068 ), .Z(\GFM/n2063 ) );
XOR2_X2 \GFM/U2323  ( .A(\GFM/n20710 ), .B(\GFM/n20700 ), .Z(\GFM/n20640 ));
XOR2_X2 \GFM/U2322  ( .A(\GFM/n20730 ), .B(\GFM/n20721 ), .Z(\GFM/n2065 ) );
XOR2_X2 \GFM/U2321  ( .A(z_in[125]), .B(\GFM/n20740 ), .Z(\GFM/n20660 ) );
XOR2_X2 \GFM/U2320  ( .A(\GFM/N4269 ), .B(\GFM/N4272 ), .Z(\GFM/n20670 ) );
XOR2_X2 \GFM/U2319  ( .A(\GFM/N4263 ), .B(\GFM/N4265 ), .Z(\GFM/n2068 ) );
XOR2_X2 \GFM/U2318  ( .A(\GFM/N4255 ), .B(\GFM/N4258 ), .Z(\GFM/n2069 ) );
XOR2_X2 \GFM/U2317  ( .A(\GFM/N4249 ), .B(\GFM/N4251 ), .Z(\GFM/n20700 ) );
XOR2_X2 \GFM/U2316  ( .A(\GFM/N4240 ), .B(\GFM/N4243 ), .Z(\GFM/n20710 ) );
XOR2_X2 \GFM/U2315  ( .A(\GFM/N4233 ), .B(\GFM/N4236 ), .Z(\GFM/n20721 ) );
XOR2_X2 \GFM/U2314  ( .A(\GFM/N4225 ), .B(\GFM/N4228 ), .Z(\GFM/n20730 ) );
XOR2_X2 \GFM/U2313  ( .A(\GFM/N4218 ), .B(\GFM/N4221 ), .Z(\GFM/n20740 ) );
XOR2_X2 \GFM/U2312  ( .A(\GFM/n2076 ), .B(\GFM/n2075 ), .Z(z_out[126]) );
XOR2_X2 \GFM/U2311  ( .A(\GFM/n20780 ), .B(\GFM/n2077 ), .Z(\GFM/n2075 ) );
XOR2_X2 \GFM/U2310  ( .A(\GFM/n20800 ), .B(\GFM/n2079 ), .Z(\GFM/n2076 ) );
XOR2_X2 \GFM/U2309  ( .A(\GFM/n2082 ), .B(\GFM/n20810 ), .Z(\GFM/n2077 ) );
XOR2_X2 \GFM/U2308  ( .A(\GFM/n20840 ), .B(\GFM/n2083 ), .Z(\GFM/n20780 ) );
XOR2_X2 \GFM/U2307  ( .A(\GFM/n2086 ), .B(\GFM/n20850 ), .Z(\GFM/n2079 ) );
XOR2_X2 \GFM/U2306  ( .A(\GFM/n20880 ), .B(\GFM/n20870 ), .Z(\GFM/n20800 ));
XOR2_X2 \GFM/U2305  ( .A(z_in[126]), .B(\GFM/n2089 ), .Z(\GFM/n20810 ) );
XOR2_X2 \GFM/U2304  ( .A(\GFM/N4316 ), .B(\GFM/N4318 ), .Z(\GFM/n2082 ) );
XOR2_X2 \GFM/U2303  ( .A(\GFM/N4311 ), .B(\GFM/N4313 ), .Z(\GFM/n2083 ) );
XOR2_X2 \GFM/U2302  ( .A(\GFM/N4305 ), .B(\GFM/N4307 ), .Z(\GFM/n20840 ) );
XOR2_X2 \GFM/U2301  ( .A(\GFM/N4300 ), .B(\GFM/N4302 ), .Z(\GFM/n20850 ) );
XOR2_X2 \GFM/U2300  ( .A(\GFM/N4293 ), .B(\GFM/N4295 ), .Z(\GFM/n2086 ) );
XOR2_X2 \GFM/U2299  ( .A(\GFM/N4288 ), .B(\GFM/N4290 ), .Z(\GFM/n20870 ) );
XOR2_X2 \GFM/U2298  ( .A(\GFM/N4282 ), .B(\GFM/N4284 ), .Z(\GFM/n20880 ) );
XOR2_X2 \GFM/U2297  ( .A(\GFM/N4276 ), .B(\GFM/N4279 ), .Z(\GFM/n2089 ) );
XOR2_X2 \GFM/U2296  ( .A(\GFM/n2091 ), .B(\GFM/n2090 ), .Z(z_out[127]) );
XOR2_X2 \GFM/U2295  ( .A(\GFM/n20930 ), .B(\GFM/n20920 ), .Z(\GFM/n2090 ) );
XOR2_X2 \GFM/U2294  ( .A(\GFM/n20950 ), .B(\GFM/n2094 ), .Z(\GFM/n2091 ) );
XOR2_X2 \GFM/U2293  ( .A(\GFM/n20970 ), .B(\GFM/n2096 ), .Z(\GFM/n20920 ) );
XOR2_X2 \GFM/U2292  ( .A(\GFM/n2099 ), .B(\GFM/n20980 ), .Z(\GFM/n20930 ) );
XOR2_X2 \GFM/U2291  ( .A(\GFM/n21010 ), .B(\GFM/n21001 ), .Z(\GFM/n2094 ) );
XOR2_X2 \GFM/U2290  ( .A(\GFM/n2103 ), .B(\GFM/n21020 ), .Z(\GFM/n20950 ) );
XOR2_X2 \GFM/U2289  ( .A(z_in[127]), .B(\GFM/n21040 ), .Z(\GFM/n2096 ) );
XOR2_X2 \GFM/U2288  ( .A(\GFM/N4348 ), .B(\GFM/N4349 ), .Z(\GFM/n20970 ) );
XOR2_X2 \GFM/U2287  ( .A(\GFM/N4345 ), .B(\GFM/N4346 ), .Z(\GFM/n20980 ) );
XOR2_X2 \GFM/U2286  ( .A(\GFM/N4341 ), .B(\GFM/N4342 ), .Z(\GFM/n2099 ) );
XOR2_X2 \GFM/U2285  ( .A(\GFM/N4337 ), .B(\GFM/N4339 ), .Z(\GFM/n21001 ) );
XOR2_X2 \GFM/U2284  ( .A(\GFM/N4332 ), .B(\GFM/N4336 ), .Z(\GFM/n21010 ) );
XOR2_X2 \GFM/U2283  ( .A(\GFM/N4329 ), .B(\GFM/N4331 ), .Z(\GFM/n21020 ) );
XOR2_X2 \GFM/U2282  ( .A(\GFM/N4325 ), .B(\GFM/N4328 ), .Z(\GFM/n2103 ) );
XOR2_X2 \GFM/U2281  ( .A(\GFM/N4322 ), .B(\GFM/N4324 ), .Z(\GFM/n21040 ) );
XOR2_X2 \GFM/U2280  ( .A(v_in[0]), .B(\GFM/n21050 ), .Z(v_out[110]) );
XOR2_X2 \GFM/U2279  ( .A(v_in[126]), .B(v_in[5]), .Z(\GFM/n21050 ) );
XOR2_X2 \GFM/U2278  ( .A(v_in[0]), .B(\GFM/n2106 ), .Z(\GFM/N4224 ) );
XOR2_X2 \GFM/U2277  ( .A(v_in[127]), .B(v_in[1]), .Z(\GFM/n2106 ) );
XOR2_X2 \GFM/U2276  ( .A(v_in[6]), .B(\GFM/N4224 ), .Z(v_out[111]) );
XOR2_X2 \GFM/U2275  ( .A(v_in[0]), .B(\GFM/n2107 ), .Z(\GFM/N4227 ) );
XOR2_X2 \GFM/U2274  ( .A(v_in[2]), .B(v_in[1]), .Z(\GFM/n2107 ) );
XOR2_X2 \GFM/U2273  ( .A(v_in[7]), .B(\GFM/N4227 ), .Z(v_out[112]) );
XOR2_X2 \GFM/U2272  ( .A(v_in[1]), .B(\GFM/n2108 ), .Z(\GFM/N4235 ) );
XOR2_X2 \GFM/U2271  ( .A(v_in[3]), .B(v_in[2]), .Z(\GFM/n2108 ) );
XOR2_X2 \GFM/U2270  ( .A(v_in[8]), .B(\GFM/N4235 ), .Z(v_out[113]) );
XOR2_X2 \GFM/U2269  ( .A(v_in[2]), .B(\GFM/n21090 ), .Z(\GFM/N4232 ) );
XOR2_X2 \GFM/U2268  ( .A(v_in[4]), .B(v_in[3]), .Z(\GFM/n21090 ) );
XOR2_X2 \GFM/U2267  ( .A(v_in[9]), .B(\GFM/N4232 ), .Z(v_out[114]) );
XOR2_X2 \GFM/U2266  ( .A(v_in[3]), .B(\GFM/n21101 ), .Z(\GFM/N4239 ) );
XOR2_X2 \GFM/U2265  ( .A(v_in[5]), .B(v_in[4]), .Z(\GFM/n21101 ) );
XOR2_X2 \GFM/U2264  ( .A(v_in[10]), .B(\GFM/N4239 ), .Z(v_out[115]) );
XOR2_X2 \GFM/U2263  ( .A(v_in[4]), .B(\GFM/n21110 ), .Z(\GFM/N4242 ) );
XOR2_X2 \GFM/U2262  ( .A(v_in[6]), .B(v_in[5]), .Z(\GFM/n21110 ) );
XOR2_X2 \GFM/U2261  ( .A(v_in[11]), .B(\GFM/N4242 ), .Z(v_out[116]) );
XOR2_X2 \GFM/U2260  ( .A(v_in[5]), .B(\GFM/n21120 ), .Z(\GFM/N4257 ) );
XOR2_X2 \GFM/U2259  ( .A(v_in[7]), .B(v_in[6]), .Z(\GFM/n21120 ) );
XOR2_X2 \GFM/U2258  ( .A(v_in[12]), .B(\GFM/N4257 ), .Z(v_out[117]) );
XOR2_X2 \GFM/U2257  ( .A(v_in[6]), .B(\GFM/n2113 ), .Z(\GFM/N4254 ) );
XOR2_X2 \GFM/U2256  ( .A(v_in[8]), .B(v_in[7]), .Z(\GFM/n2113 ) );
XOR2_X2 \GFM/U2255  ( .A(v_in[13]), .B(\GFM/N4254 ), .Z(v_out[118]) );
XOR2_X2 \GFM/U2254  ( .A(v_in[7]), .B(\GFM/n2114 ), .Z(\GFM/N4248 ) );
XOR2_X2 \GFM/U2253  ( .A(v_in[9]), .B(v_in[8]), .Z(\GFM/n2114 ) );
XOR2_X2 \GFM/U2252  ( .A(v_in[14]), .B(\GFM/N4248 ), .Z(v_out[119]) );
XOR2_X2 \GFM/U2251  ( .A(v_in[8]), .B(\GFM/n21150 ), .Z(\GFM/N4250 ) );
XOR2_X2 \GFM/U2250  ( .A(v_in[10]), .B(v_in[9]), .Z(\GFM/n21150 ) );
XOR2_X2 \GFM/U2249  ( .A(v_in[15]), .B(\GFM/N4250 ), .Z(v_out[120]) );
XOR2_X2 \GFM/U2248  ( .A(v_in[9]), .B(\GFM/n21160 ), .Z(v_out[121]) );
XOR2_X2 \GFM/U2247  ( .A(v_in[11]), .B(v_in[10]), .Z(\GFM/n21160 ) );
XOR2_X2 \GFM/U2246  ( .A(v_in[10]), .B(\GFM/n2117 ), .Z(v_out[122]) );
XOR2_X2 \GFM/U2245  ( .A(v_in[12]), .B(v_in[11]), .Z(\GFM/n2117 ) );
XOR2_X2 \GFM/U2244  ( .A(v_in[11]), .B(\GFM/n21180 ), .Z(v_out[123]) );
XOR2_X2 \GFM/U2243  ( .A(v_in[13]), .B(v_in[12]), .Z(\GFM/n21180 ) );
XOR2_X2 \GFM/U2242  ( .A(v_in[12]), .B(\GFM/n21190 ), .Z(v_out[124]) );
XOR2_X2 \GFM/U2241  ( .A(v_in[14]), .B(v_in[13]), .Z(\GFM/n21190 ) );
XOR2_X2 \GFM/U2240  ( .A(v_in[13]), .B(\GFM/n2120 ), .Z(v_out[125]) );
XOR2_X2 \GFM/U2239  ( .A(v_in[15]), .B(v_in[14]), .Z(\GFM/n2120 ) );
INV_X4 \AES_ENC/U1636  ( .A(rst), .ZN(\AES_ENC/n1267 ) );
INV_X4 \AES_ENC/U1635  ( .A(\AES_ENC/n17 ), .ZN(\AES_ENC/n1266 ) );
NAND3_X2 \AES_ENC/U1634  ( .A1(\AES_ENC/n15 ), .A2(\AES_ENC/n1258 ), .A3(\AES_ENC/n16 ), .ZN(\AES_ENC/n796 ) );
NOR2_X2 \AES_ENC/U1633  ( .A1(\AES_ENC/n22 ), .A2(\AES_ENC/n2 ), .ZN(\AES_ENC/n17 ) );
NOR2_X2 \AES_ENC/U1632  ( .A1(\AES_ENC/n1234 ), .A2(\AES_ENC/n1231 ), .ZN(\AES_ENC/n14 ) );
NOR2_X2 \AES_ENC/U1631  ( .A1(\AES_ENC/n1232 ), .A2(\AES_ENC/n22 ), .ZN(\AES_ENC/n11 ) );
INV_X4 \AES_ENC/U1630  ( .A(\AES_ENC/n1258 ), .ZN(\AES_ENC/n1265 ) );
INV_X4 \AES_ENC/U1629  ( .A(\AES_ENC/n1256 ), .ZN(\AES_ENC/n1250 ) );
INV_X4 \AES_ENC/U1628  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1246 ) );
INV_X4 \AES_ENC/U1627  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1247 ) );
INV_X4 \AES_ENC/U1626  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1245 ) );
INV_X4 \AES_ENC/U1625  ( .A(\AES_ENC/n1255 ), .ZN(\AES_ENC/n1248 ) );
INV_X4 \AES_ENC/U1624  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1249 ) );
INV_X4 \AES_ENC/U1623  ( .A(\AES_ENC/n1265 ), .ZN(\AES_ENC/n1259 ) );
INV_X4 \AES_ENC/U1622  ( .A(\AES_ENC/n1238 ), .ZN(\AES_ENC/n1254 ) );
INV_X4 \AES_ENC/U1621  ( .A(\AES_ENC/n1238 ), .ZN(\AES_ENC/n1253 ) );
INV_X4 \AES_ENC/U1620  ( .A(\AES_ENC/n1238 ), .ZN(\AES_ENC/n1252 ) );
INV_X4 \AES_ENC/U1619  ( .A(\AES_ENC/n1238 ), .ZN(\AES_ENC/n1256 ) );
INV_X4 \AES_ENC/U1618  ( .A(\AES_ENC/n1238 ), .ZN(\AES_ENC/n1255 ) );
INV_X4 \AES_ENC/U1617  ( .A(\AES_ENC/n1238 ), .ZN(\AES_ENC/n1251 ) );
INV_X4 \AES_ENC/U1616  ( .A(\AES_ENC/n1265 ), .ZN(\AES_ENC/n12601 ) );
INV_X4 \AES_ENC/U1615  ( .A(\AES_ENC/n1265 ), .ZN(\AES_ENC/n1261 ) );
INV_X4 \AES_ENC/U1614  ( .A(\AES_ENC/n1265 ), .ZN(\AES_ENC/n1262 ) );
INV_X4 \AES_ENC/U1613  ( .A(\AES_ENC/n1265 ), .ZN(\AES_ENC/n1263 ) );
INV_X4 \AES_ENC/U1052  ( .A(\AES_ENC/n1265 ), .ZN(\AES_ENC/n1264 ) );
INV_X4 \AES_ENC/U1051  ( .A(aes_kld), .ZN(\AES_ENC/n1258 ) );
INV_X4 \AES_ENC/U1050  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1244 ) );
INV_X4 \AES_ENC/U1049  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1241 ) );
INV_X4 \AES_ENC/U1048  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1239 ) );
INV_X4 \AES_ENC/U1047  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1242 ) );
INV_X4 \AES_ENC/U1046  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1243 ) );
INV_X4 \AES_ENC/U1045  ( .A(\AES_ENC/n793 ), .ZN(\AES_ENC/n1240 ) );
INV_X4 \AES_ENC/U876  ( .A(\AES_ENC/n1258 ), .ZN(\AES_ENC/n1257 ) );
INV_X4 \AES_ENC/U16  ( .A(\AES_ENC/n1258 ), .ZN(\AES_ENC/n1237 ) );
INV_X4 \AES_ENC/U14  ( .A(\AES_ENC/n1258 ), .ZN(\AES_ENC/n1236 ) );
INV_X4 \AES_ENC/U7  ( .A(\AES_ENC/n1258 ), .ZN(\AES_ENC/n1235 ) );
DFF_X1 \AES_ENC/ld_r_reg  ( .D(aes_kld), .CK(clk), .Q(\AES_ENC/n1238 ), .QN(\AES_ENC/n793 ) );
NAND2_X2 \AES_ENC/U1044  ( .A1(\AES_ENC/sa32_next [6]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n7891 ) );
XOR2_X2 \AES_ENC/U1043  ( .A(\AES_ENC/w2[6] ), .B(\AES_ENC/text_in_r[38] ),.Z(\AES_ENC/n791 ) );
NAND2_X2 \AES_ENC/U1042  ( .A1(\AES_ENC/n791 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n7901 ) );
NAND2_X2 \AES_ENC/U1041  ( .A1(\AES_ENC/n7891 ), .A2(\AES_ENC/n7901 ), .ZN(\AES_ENC/N100 ) );
NAND2_X2 \AES_ENC/U1040  ( .A1(\AES_ENC/sa32_next [7]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n658 ) );
XOR2_X2 \AES_ENC/U1039  ( .A(\AES_ENC/w2[7] ), .B(\AES_ENC/text_in_r[39] ),.Z(\AES_ENC/n6601 ) );
NAND2_X2 \AES_ENC/U1038  ( .A1(\AES_ENC/n6601 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n659 ) );
NAND2_X2 \AES_ENC/U1037  ( .A1(\AES_ENC/n658 ), .A2(\AES_ENC/n659 ), .ZN(\AES_ENC/N101 ) );
NAND2_X2 \AES_ENC/U1036  ( .A1(\AES_ENC/sa22_next [0]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n655 ) );
XOR2_X2 \AES_ENC/U1035  ( .A(\AES_ENC/w2[8] ), .B(\AES_ENC/text_in_r[40] ),.Z(\AES_ENC/n657 ) );
NAND2_X2 \AES_ENC/U1034  ( .A1(\AES_ENC/n657 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n656 ) );
NAND2_X2 \AES_ENC/U1033  ( .A1(\AES_ENC/n655 ), .A2(\AES_ENC/n656 ), .ZN(\AES_ENC/N110 ) );
NAND2_X2 \AES_ENC/U1032  ( .A1(\AES_ENC/sa22_next [1]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n652 ) );
XOR2_X2 \AES_ENC/U1031  ( .A(\AES_ENC/w2[9] ), .B(\AES_ENC/text_in_r[41] ),.Z(\AES_ENC/n654 ) );
NAND2_X2 \AES_ENC/U1030  ( .A1(\AES_ENC/n654 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n653 ) );
NAND2_X2 \AES_ENC/U1029  ( .A1(\AES_ENC/n652 ), .A2(\AES_ENC/n653 ), .ZN(\AES_ENC/N111 ) );
NAND2_X2 \AES_ENC/U1028  ( .A1(\AES_ENC/sa22_next [2]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n649 ) );
XOR2_X2 \AES_ENC/U1027  ( .A(\AES_ENC/w2[10] ), .B(\AES_ENC/text_in_r[42] ),.Z(\AES_ENC/n651 ) );
NAND2_X2 \AES_ENC/U1026  ( .A1(\AES_ENC/n651 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n6501 ) );
NAND2_X2 \AES_ENC/U1025  ( .A1(\AES_ENC/n649 ), .A2(\AES_ENC/n6501 ), .ZN(\AES_ENC/N112 ) );
NAND2_X2 \AES_ENC/U1024  ( .A1(\AES_ENC/sa22_next [3]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n646 ) );
XOR2_X2 \AES_ENC/U1023  ( .A(\AES_ENC/w2[11] ), .B(\AES_ENC/text_in_r[43] ),.Z(\AES_ENC/n648 ) );
NAND2_X2 \AES_ENC/U1022  ( .A1(\AES_ENC/n648 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n647 ) );
NAND2_X2 \AES_ENC/U1021  ( .A1(\AES_ENC/n646 ), .A2(\AES_ENC/n647 ), .ZN(\AES_ENC/N113 ) );
NAND2_X2 \AES_ENC/U1020  ( .A1(\AES_ENC/sa22_next [4]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n643 ) );
XOR2_X2 \AES_ENC/U1019  ( .A(\AES_ENC/w2[12] ), .B(\AES_ENC/text_in_r[44] ),.Z(\AES_ENC/n645 ) );
NAND2_X2 \AES_ENC/U1018  ( .A1(\AES_ENC/n645 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n644 ) );
NAND2_X2 \AES_ENC/U1017  ( .A1(\AES_ENC/n643 ), .A2(\AES_ENC/n644 ), .ZN(\AES_ENC/N114 ) );
NAND2_X2 \AES_ENC/U1016  ( .A1(\AES_ENC/sa22_next [5]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n6401 ) );
XOR2_X2 \AES_ENC/U1015  ( .A(\AES_ENC/w2[13] ), .B(\AES_ENC/text_in_r[45] ),.Z(\AES_ENC/n642 ) );
NAND2_X2 \AES_ENC/U1014  ( .A1(\AES_ENC/n642 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n641 ) );
NAND2_X2 \AES_ENC/U1013  ( .A1(\AES_ENC/n6401 ), .A2(\AES_ENC/n641 ), .ZN(\AES_ENC/N115 ) );
NAND2_X2 \AES_ENC/U1012  ( .A1(\AES_ENC/sa22_next [6]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n637 ) );
XOR2_X2 \AES_ENC/U1011  ( .A(\AES_ENC/w2[14] ), .B(\AES_ENC/text_in_r[46] ),.Z(\AES_ENC/n639 ) );
NAND2_X2 \AES_ENC/U1010  ( .A1(\AES_ENC/n639 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n638 ) );
NAND2_X2 \AES_ENC/U1009  ( .A1(\AES_ENC/n637 ), .A2(\AES_ENC/n638 ), .ZN(\AES_ENC/N116 ) );
NAND2_X2 \AES_ENC/U1008  ( .A1(\AES_ENC/sa22_next [7]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n634 ) );
XOR2_X2 \AES_ENC/U1007  ( .A(\AES_ENC/w2[15] ), .B(\AES_ENC/text_in_r[47] ),.Z(\AES_ENC/n636 ) );
NAND2_X2 \AES_ENC/U1006  ( .A1(\AES_ENC/n636 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n635 ) );
NAND2_X2 \AES_ENC/U1005  ( .A1(\AES_ENC/n634 ), .A2(\AES_ENC/n635 ), .ZN(\AES_ENC/N117 ) );
NAND2_X2 \AES_ENC/U1004  ( .A1(\AES_ENC/sa12_next [0]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n631 ) );
XOR2_X2 \AES_ENC/U1003  ( .A(\AES_ENC/w2[16] ), .B(\AES_ENC/text_in_r[48] ),.Z(\AES_ENC/n633 ) );
NAND2_X2 \AES_ENC/U1002  ( .A1(\AES_ENC/n633 ), .A2(\AES_ENC/n1239 ), .ZN(\AES_ENC/n632 ) );
NAND2_X2 \AES_ENC/U1001  ( .A1(\AES_ENC/n631 ), .A2(\AES_ENC/n632 ), .ZN(\AES_ENC/N126 ) );
NAND2_X2 \AES_ENC/U1000  ( .A1(\AES_ENC/sa12_next [1]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n628 ) );
XOR2_X2 \AES_ENC/U999  ( .A(\AES_ENC/w2[17] ), .B(\AES_ENC/text_in_r[49] ),.Z(\AES_ENC/n6301 ) );
NAND2_X2 \AES_ENC/U998  ( .A1(\AES_ENC/n6301 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n629 ) );
NAND2_X2 \AES_ENC/U997  ( .A1(\AES_ENC/n628 ), .A2(\AES_ENC/n629 ), .ZN(\AES_ENC/N127 ) );
NAND2_X2 \AES_ENC/U996  ( .A1(\AES_ENC/sa12_next [2]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n625 ) );
XOR2_X2 \AES_ENC/U995  ( .A(\AES_ENC/w2[18] ), .B(\AES_ENC/text_in_r[50] ),.Z(\AES_ENC/n627 ) );
NAND2_X2 \AES_ENC/U994  ( .A1(\AES_ENC/n627 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n626 ) );
NAND2_X2 \AES_ENC/U993  ( .A1(\AES_ENC/n625 ), .A2(\AES_ENC/n626 ), .ZN(\AES_ENC/N128 ) );
NAND2_X2 \AES_ENC/U992  ( .A1(\AES_ENC/sa12_next [3]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n622 ) );
XOR2_X2 \AES_ENC/U991  ( .A(\AES_ENC/w2[19] ), .B(\AES_ENC/text_in_r[51] ),.Z(\AES_ENC/n624 ) );
NAND2_X2 \AES_ENC/U990  ( .A1(\AES_ENC/n624 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n623 ) );
NAND2_X2 \AES_ENC/U989  ( .A1(\AES_ENC/n622 ), .A2(\AES_ENC/n623 ), .ZN(\AES_ENC/N129 ) );
NAND2_X2 \AES_ENC/U988  ( .A1(\AES_ENC/sa12_next [4]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n619 ) );
XOR2_X2 \AES_ENC/U987  ( .A(\AES_ENC/w2[20] ), .B(\AES_ENC/text_in_r[52] ),.Z(\AES_ENC/n621 ) );
NAND2_X2 \AES_ENC/U986  ( .A1(\AES_ENC/n621 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n6201 ) );
NAND2_X2 \AES_ENC/U985  ( .A1(\AES_ENC/n619 ), .A2(\AES_ENC/n6201 ), .ZN(\AES_ENC/N130 ) );
NAND2_X2 \AES_ENC/U984  ( .A1(\AES_ENC/sa12_next [5]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n616 ) );
XOR2_X2 \AES_ENC/U983  ( .A(\AES_ENC/w2[21] ), .B(\AES_ENC/text_in_r[53] ),.Z(\AES_ENC/n618 ) );
NAND2_X2 \AES_ENC/U982  ( .A1(\AES_ENC/n618 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n617 ) );
NAND2_X2 \AES_ENC/U981  ( .A1(\AES_ENC/n616 ), .A2(\AES_ENC/n617 ), .ZN(\AES_ENC/N131 ) );
NAND2_X2 \AES_ENC/U980  ( .A1(\AES_ENC/sa12_next [6]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n613 ) );
XOR2_X2 \AES_ENC/U979  ( .A(\AES_ENC/w2[22] ), .B(\AES_ENC/text_in_r[54] ),.Z(\AES_ENC/n615 ) );
NAND2_X2 \AES_ENC/U978  ( .A1(\AES_ENC/n615 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n614 ) );
NAND2_X2 \AES_ENC/U977  ( .A1(\AES_ENC/n613 ), .A2(\AES_ENC/n614 ), .ZN(\AES_ENC/N132 ) );
NAND2_X2 \AES_ENC/U976  ( .A1(\AES_ENC/sa12_next [7]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n610 ) );
XOR2_X2 \AES_ENC/U975  ( .A(\AES_ENC/w2[23] ), .B(\AES_ENC/text_in_r[55] ),.Z(\AES_ENC/n612 ) );
NAND2_X2 \AES_ENC/U974  ( .A1(\AES_ENC/n612 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n611 ) );
NAND2_X2 \AES_ENC/U973  ( .A1(\AES_ENC/n610 ), .A2(\AES_ENC/n611 ), .ZN(\AES_ENC/N133 ) );
NAND2_X2 \AES_ENC/U972  ( .A1(\AES_ENC/sa02_next [0]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n607 ) );
XOR2_X2 \AES_ENC/U971  ( .A(\AES_ENC/w2[24] ), .B(\AES_ENC/text_in_r[56] ),.Z(\AES_ENC/n609 ) );
NAND2_X2 \AES_ENC/U970  ( .A1(\AES_ENC/n609 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n608 ) );
NAND2_X2 \AES_ENC/U969  ( .A1(\AES_ENC/n607 ), .A2(\AES_ENC/n608 ), .ZN(\AES_ENC/N142 ) );
NAND2_X2 \AES_ENC/U968  ( .A1(\AES_ENC/sa02_next [1]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n604 ) );
XOR2_X2 \AES_ENC/U967  ( .A(\AES_ENC/w2[25] ), .B(\AES_ENC/text_in_r[57] ),.Z(\AES_ENC/n606 ) );
NAND2_X2 \AES_ENC/U966  ( .A1(\AES_ENC/n606 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n605 ) );
NAND2_X2 \AES_ENC/U965  ( .A1(\AES_ENC/n604 ), .A2(\AES_ENC/n605 ), .ZN(\AES_ENC/N143 ) );
NAND2_X2 \AES_ENC/U964  ( .A1(\AES_ENC/sa02_next [2]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n601 ) );
XOR2_X2 \AES_ENC/U963  ( .A(\AES_ENC/w2[26] ), .B(\AES_ENC/text_in_r[58] ),.Z(\AES_ENC/n603 ) );
NAND2_X2 \AES_ENC/U962  ( .A1(\AES_ENC/n603 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n602 ) );
NAND2_X2 \AES_ENC/U961  ( .A1(\AES_ENC/n601 ), .A2(\AES_ENC/n602 ), .ZN(\AES_ENC/N144 ) );
NAND2_X2 \AES_ENC/U960  ( .A1(\AES_ENC/sa02_next [3]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n598 ) );
XOR2_X2 \AES_ENC/U959  ( .A(\AES_ENC/w2[27] ), .B(\AES_ENC/text_in_r[59] ),.Z(\AES_ENC/n600 ) );
NAND2_X2 \AES_ENC/U958  ( .A1(\AES_ENC/n600 ), .A2(\AES_ENC/n1240 ), .ZN(\AES_ENC/n599 ) );
NAND2_X2 \AES_ENC/U957  ( .A1(\AES_ENC/n598 ), .A2(\AES_ENC/n599 ), .ZN(\AES_ENC/N145 ) );
NAND2_X2 \AES_ENC/U956  ( .A1(\AES_ENC/sa02_next [4]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n595 ) );
XOR2_X2 \AES_ENC/U955  ( .A(\AES_ENC/w2[28] ), .B(\AES_ENC/text_in_r[60] ),.Z(\AES_ENC/n597 ) );
NAND2_X2 \AES_ENC/U954  ( .A1(\AES_ENC/n597 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n596 ) );
NAND2_X2 \AES_ENC/U953  ( .A1(\AES_ENC/n595 ), .A2(\AES_ENC/n596 ), .ZN(\AES_ENC/N146 ) );
NAND2_X2 \AES_ENC/U952  ( .A1(\AES_ENC/sa02_next [5]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n592 ) );
XOR2_X2 \AES_ENC/U951  ( .A(\AES_ENC/w2[29] ), .B(\AES_ENC/text_in_r[61] ),.Z(\AES_ENC/n594 ) );
NAND2_X2 \AES_ENC/U950  ( .A1(\AES_ENC/n594 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n593 ) );
NAND2_X2 \AES_ENC/U949  ( .A1(\AES_ENC/n592 ), .A2(\AES_ENC/n593 ), .ZN(\AES_ENC/N147 ) );
NAND2_X2 \AES_ENC/U948  ( .A1(\AES_ENC/sa02_next [6]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n589 ) );
XOR2_X2 \AES_ENC/U947  ( .A(\AES_ENC/w2[30] ), .B(\AES_ENC/text_in_r[62] ),.Z(\AES_ENC/n591 ) );
NAND2_X2 \AES_ENC/U946  ( .A1(\AES_ENC/n591 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n590 ) );
NAND2_X2 \AES_ENC/U945  ( .A1(\AES_ENC/n589 ), .A2(\AES_ENC/n590 ), .ZN(\AES_ENC/N148 ) );
NAND2_X2 \AES_ENC/U944  ( .A1(\AES_ENC/sa02_next [7]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n586 ) );
XOR2_X2 \AES_ENC/U943  ( .A(\AES_ENC/w2[31] ), .B(\AES_ENC/text_in_r[63] ),.Z(\AES_ENC/n588 ) );
NAND2_X2 \AES_ENC/U942  ( .A1(\AES_ENC/n588 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n587 ) );
NAND2_X2 \AES_ENC/U941  ( .A1(\AES_ENC/n586 ), .A2(\AES_ENC/n587 ), .ZN(\AES_ENC/N149 ) );
NAND2_X2 \AES_ENC/U940  ( .A1(\AES_ENC/sa31_next [0]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n583 ) );
XOR2_X2 \AES_ENC/U939  ( .A(\AES_ENC/w1[0] ), .B(\AES_ENC/text_in_r[64] ),.Z(\AES_ENC/n585 ) );
NAND2_X2 \AES_ENC/U938  ( .A1(\AES_ENC/n585 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n584 ) );
NAND2_X2 \AES_ENC/U937  ( .A1(\AES_ENC/n583 ), .A2(\AES_ENC/n584 ), .ZN(\AES_ENC/N158 ) );
NAND2_X2 \AES_ENC/U936  ( .A1(\AES_ENC/sa31_next [1]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n580 ) );
XOR2_X2 \AES_ENC/U935  ( .A(\AES_ENC/w1[1] ), .B(\AES_ENC/text_in_r[65] ),.Z(\AES_ENC/n582 ) );
NAND2_X2 \AES_ENC/U934  ( .A1(\AES_ENC/n582 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n581 ) );
NAND2_X2 \AES_ENC/U933  ( .A1(\AES_ENC/n580 ), .A2(\AES_ENC/n581 ), .ZN(\AES_ENC/N159 ) );
NAND2_X2 \AES_ENC/U932  ( .A1(\AES_ENC/sa31_next [2]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n577 ) );
XOR2_X2 \AES_ENC/U931  ( .A(\AES_ENC/w1[2] ), .B(\AES_ENC/text_in_r[66] ),.Z(\AES_ENC/n579 ) );
NAND2_X2 \AES_ENC/U930  ( .A1(\AES_ENC/n579 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n578 ) );
NAND2_X2 \AES_ENC/U929  ( .A1(\AES_ENC/n577 ), .A2(\AES_ENC/n578 ), .ZN(\AES_ENC/N160 ) );
NAND2_X2 \AES_ENC/U928  ( .A1(\AES_ENC/sa31_next [3]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n574 ) );
XOR2_X2 \AES_ENC/U927  ( .A(\AES_ENC/w1[3] ), .B(\AES_ENC/text_in_r[67] ),.Z(\AES_ENC/n576 ) );
NAND2_X2 \AES_ENC/U926  ( .A1(\AES_ENC/n576 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n575 ) );
NAND2_X2 \AES_ENC/U925  ( .A1(\AES_ENC/n574 ), .A2(\AES_ENC/n575 ), .ZN(\AES_ENC/N161 ) );
NAND2_X2 \AES_ENC/U924  ( .A1(\AES_ENC/sa31_next [4]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n571 ) );
XOR2_X2 \AES_ENC/U923  ( .A(\AES_ENC/w1[4] ), .B(\AES_ENC/text_in_r[68] ),.Z(\AES_ENC/n573 ) );
NAND2_X2 \AES_ENC/U922  ( .A1(\AES_ENC/n573 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n572 ) );
NAND2_X2 \AES_ENC/U921  ( .A1(\AES_ENC/n571 ), .A2(\AES_ENC/n572 ), .ZN(\AES_ENC/N162 ) );
NAND2_X2 \AES_ENC/U920  ( .A1(\AES_ENC/sa31_next [5]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n568 ) );
XOR2_X2 \AES_ENC/U919  ( .A(\AES_ENC/w1[5] ), .B(\AES_ENC/text_in_r[69] ),.Z(\AES_ENC/n570 ) );
NAND2_X2 \AES_ENC/U918  ( .A1(\AES_ENC/n570 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n569 ) );
NAND2_X2 \AES_ENC/U917  ( .A1(\AES_ENC/n568 ), .A2(\AES_ENC/n569 ), .ZN(\AES_ENC/N163 ) );
NAND2_X2 \AES_ENC/U916  ( .A1(\AES_ENC/sa31_next [6]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n565 ) );
XOR2_X2 \AES_ENC/U915  ( .A(\AES_ENC/w1[6] ), .B(\AES_ENC/text_in_r[70] ),.Z(\AES_ENC/n567 ) );
NAND2_X2 \AES_ENC/U914  ( .A1(\AES_ENC/n567 ), .A2(\AES_ENC/n1241 ), .ZN(\AES_ENC/n566 ) );
NAND2_X2 \AES_ENC/U913  ( .A1(\AES_ENC/n565 ), .A2(\AES_ENC/n566 ), .ZN(\AES_ENC/N164 ) );
NAND2_X2 \AES_ENC/U912  ( .A1(\AES_ENC/sa31_next [7]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n562 ) );
XOR2_X2 \AES_ENC/U911  ( .A(\AES_ENC/w1[7] ), .B(\AES_ENC/text_in_r[71] ),.Z(\AES_ENC/n564 ) );
NAND2_X2 \AES_ENC/U910  ( .A1(\AES_ENC/n564 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n563 ) );
NAND2_X2 \AES_ENC/U909  ( .A1(\AES_ENC/n562 ), .A2(\AES_ENC/n563 ), .ZN(\AES_ENC/N165 ) );
NAND2_X2 \AES_ENC/U908  ( .A1(\AES_ENC/sa21_next [0]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n559 ) );
XOR2_X2 \AES_ENC/U907  ( .A(\AES_ENC/w1[8] ), .B(\AES_ENC/text_in_r[72] ),.Z(\AES_ENC/n561 ) );
NAND2_X2 \AES_ENC/U906  ( .A1(\AES_ENC/n561 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n560 ) );
NAND2_X2 \AES_ENC/U905  ( .A1(\AES_ENC/n559 ), .A2(\AES_ENC/n560 ), .ZN(\AES_ENC/N174 ) );
NAND2_X2 \AES_ENC/U904  ( .A1(\AES_ENC/sa21_next [1]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n556 ) );
XOR2_X2 \AES_ENC/U903  ( .A(\AES_ENC/w1[9] ), .B(\AES_ENC/text_in_r[73] ),.Z(\AES_ENC/n558 ) );
NAND2_X2 \AES_ENC/U902  ( .A1(\AES_ENC/n558 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n557 ) );
NAND2_X2 \AES_ENC/U901  ( .A1(\AES_ENC/n556 ), .A2(\AES_ENC/n557 ), .ZN(\AES_ENC/N175 ) );
NAND2_X2 \AES_ENC/U900  ( .A1(\AES_ENC/sa21_next [2]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n553 ) );
XOR2_X2 \AES_ENC/U899  ( .A(\AES_ENC/w1[10] ), .B(\AES_ENC/text_in_r[74] ),.Z(\AES_ENC/n555 ) );
NAND2_X2 \AES_ENC/U898  ( .A1(\AES_ENC/n555 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n554 ) );
NAND2_X2 \AES_ENC/U897  ( .A1(\AES_ENC/n553 ), .A2(\AES_ENC/n554 ), .ZN(\AES_ENC/N176 ) );
NAND2_X2 \AES_ENC/U896  ( .A1(\AES_ENC/sa21_next [3]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n550 ) );
XOR2_X2 \AES_ENC/U895  ( .A(\AES_ENC/w1[11] ), .B(\AES_ENC/text_in_r[75] ),.Z(\AES_ENC/n552 ) );
NAND2_X2 \AES_ENC/U894  ( .A1(\AES_ENC/n552 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n551 ) );
NAND2_X2 \AES_ENC/U893  ( .A1(\AES_ENC/n550 ), .A2(\AES_ENC/n551 ), .ZN(\AES_ENC/N177 ) );
NAND2_X2 \AES_ENC/U892  ( .A1(\AES_ENC/sa21_next [4]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n547 ) );
XOR2_X2 \AES_ENC/U891  ( .A(\AES_ENC/w1[12] ), .B(\AES_ENC/text_in_r[76] ),.Z(\AES_ENC/n549 ) );
NAND2_X2 \AES_ENC/U890  ( .A1(\AES_ENC/n549 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n548 ) );
NAND2_X2 \AES_ENC/U889  ( .A1(\AES_ENC/n547 ), .A2(\AES_ENC/n548 ), .ZN(\AES_ENC/N178 ) );
NAND2_X2 \AES_ENC/U888  ( .A1(\AES_ENC/sa21_next [5]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n544 ) );
XOR2_X2 \AES_ENC/U887  ( .A(\AES_ENC/w1[13] ), .B(\AES_ENC/text_in_r[77] ),.Z(\AES_ENC/n546 ) );
NAND2_X2 \AES_ENC/U886  ( .A1(\AES_ENC/n546 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n545 ) );
NAND2_X2 \AES_ENC/U885  ( .A1(\AES_ENC/n544 ), .A2(\AES_ENC/n545 ), .ZN(\AES_ENC/N179 ) );
NAND2_X2 \AES_ENC/U884  ( .A1(\AES_ENC/sa21_next [6]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n541 ) );
XOR2_X2 \AES_ENC/U883  ( .A(\AES_ENC/w1[14] ), .B(\AES_ENC/text_in_r[78] ),.Z(\AES_ENC/n543 ) );
NAND2_X2 \AES_ENC/U882  ( .A1(\AES_ENC/n543 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n542 ) );
NAND2_X2 \AES_ENC/U881  ( .A1(\AES_ENC/n541 ), .A2(\AES_ENC/n542 ), .ZN(\AES_ENC/N180 ) );
NAND2_X2 \AES_ENC/U880  ( .A1(\AES_ENC/sa21_next [7]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n538 ) );
XOR2_X2 \AES_ENC/U879  ( .A(\AES_ENC/w1[15] ), .B(\AES_ENC/text_in_r[79] ),.Z(\AES_ENC/n540 ) );
NAND2_X2 \AES_ENC/U878  ( .A1(\AES_ENC/n540 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n539 ) );
NAND2_X2 \AES_ENC/U877  ( .A1(\AES_ENC/n538 ), .A2(\AES_ENC/n539 ), .ZN(\AES_ENC/N181 ) );
AND4_X2 \AES_ENC/U875  ( .A1(\AES_ENC/n1232 ), .A2(\AES_ENC/n1259 ), .A3(\AES_ENC/n14 ), .A4(\AES_ENC/n792 ), .ZN(\AES_ENC/N19 ) );
NAND2_X2 \AES_ENC/U874  ( .A1(\AES_ENC/sa11_next [0]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n535 ) );
XOR2_X2 \AES_ENC/U873  ( .A(\AES_ENC/w1[16] ), .B(\AES_ENC/text_in_r[80] ),.Z(\AES_ENC/n537 ) );
NAND2_X2 \AES_ENC/U872  ( .A1(\AES_ENC/n537 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n536 ) );
NAND2_X2 \AES_ENC/U871  ( .A1(\AES_ENC/n535 ), .A2(\AES_ENC/n536 ), .ZN(\AES_ENC/N190 ) );
NAND2_X2 \AES_ENC/U870  ( .A1(\AES_ENC/sa11_next [1]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n532 ) );
XOR2_X2 \AES_ENC/U869  ( .A(\AES_ENC/w1[17] ), .B(\AES_ENC/text_in_r[81] ),.Z(\AES_ENC/n534 ) );
NAND2_X2 \AES_ENC/U868  ( .A1(\AES_ENC/n534 ), .A2(\AES_ENC/n1242 ), .ZN(\AES_ENC/n533 ) );
NAND2_X2 \AES_ENC/U867  ( .A1(\AES_ENC/n532 ), .A2(\AES_ENC/n533 ), .ZN(\AES_ENC/N191 ) );
NAND2_X2 \AES_ENC/U866  ( .A1(\AES_ENC/sa11_next [2]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n529 ) );
XOR2_X2 \AES_ENC/U865  ( .A(\AES_ENC/w1[18] ), .B(\AES_ENC/text_in_r[82] ),.Z(\AES_ENC/n531 ) );
NAND2_X2 \AES_ENC/U864  ( .A1(\AES_ENC/n531 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n5301 ) );
NAND2_X2 \AES_ENC/U863  ( .A1(\AES_ENC/n529 ), .A2(\AES_ENC/n5301 ), .ZN(\AES_ENC/N192 ) );
NAND2_X2 \AES_ENC/U862  ( .A1(\AES_ENC/sa11_next [3]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n526 ) );
XOR2_X2 \AES_ENC/U861  ( .A(\AES_ENC/w1[19] ), .B(\AES_ENC/text_in_r[83] ),.Z(\AES_ENC/n528 ) );
NAND2_X2 \AES_ENC/U860  ( .A1(\AES_ENC/n528 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n527 ) );
NAND2_X2 \AES_ENC/U859  ( .A1(\AES_ENC/n526 ), .A2(\AES_ENC/n527 ), .ZN(\AES_ENC/N193 ) );
NAND2_X2 \AES_ENC/U858  ( .A1(\AES_ENC/sa11_next [4]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n523 ) );
XOR2_X2 \AES_ENC/U857  ( .A(\AES_ENC/w1[20] ), .B(\AES_ENC/text_in_r[84] ),.Z(\AES_ENC/n525 ) );
NAND2_X2 \AES_ENC/U856  ( .A1(\AES_ENC/n525 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n524 ) );
NAND2_X2 \AES_ENC/U855  ( .A1(\AES_ENC/n523 ), .A2(\AES_ENC/n524 ), .ZN(\AES_ENC/N194 ) );
NAND2_X2 \AES_ENC/U854  ( .A1(\AES_ENC/sa11_next [5]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n5201 ) );
XOR2_X2 \AES_ENC/U853  ( .A(\AES_ENC/w1[21] ), .B(\AES_ENC/text_in_r[85] ),.Z(\AES_ENC/n522 ) );
NAND2_X2 \AES_ENC/U852  ( .A1(\AES_ENC/n522 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n521 ) );
NAND2_X2 \AES_ENC/U851  ( .A1(\AES_ENC/n5201 ), .A2(\AES_ENC/n521 ), .ZN(\AES_ENC/N195 ) );
NAND2_X2 \AES_ENC/U850  ( .A1(\AES_ENC/sa11_next [6]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n517 ) );
XOR2_X2 \AES_ENC/U849  ( .A(\AES_ENC/w1[22] ), .B(\AES_ENC/text_in_r[86] ),.Z(\AES_ENC/n519 ) );
NAND2_X2 \AES_ENC/U848  ( .A1(\AES_ENC/n519 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n518 ) );
NAND2_X2 \AES_ENC/U847  ( .A1(\AES_ENC/n517 ), .A2(\AES_ENC/n518 ), .ZN(\AES_ENC/N196 ) );
NAND2_X2 \AES_ENC/U846  ( .A1(\AES_ENC/sa11_next [7]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n514 ) );
XOR2_X2 \AES_ENC/U845  ( .A(\AES_ENC/w1[23] ), .B(\AES_ENC/text_in_r[87] ),.Z(\AES_ENC/n516 ) );
NAND2_X2 \AES_ENC/U844  ( .A1(\AES_ENC/n516 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n515 ) );
NAND2_X2 \AES_ENC/U843  ( .A1(\AES_ENC/n514 ), .A2(\AES_ENC/n515 ), .ZN(\AES_ENC/N197 ) );
NAND2_X2 \AES_ENC/U842  ( .A1(\AES_ENC/sa01_next [0]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n511 ) );
XOR2_X2 \AES_ENC/U841  ( .A(\AES_ENC/w1[24] ), .B(\AES_ENC/text_in_r[88] ),.Z(\AES_ENC/n513 ) );
NAND2_X2 \AES_ENC/U840  ( .A1(\AES_ENC/n513 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n512 ) );
NAND2_X2 \AES_ENC/U839  ( .A1(\AES_ENC/n511 ), .A2(\AES_ENC/n512 ), .ZN(\AES_ENC/N206 ) );
NAND2_X2 \AES_ENC/U838  ( .A1(\AES_ENC/sa01_next [1]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n508 ) );
XOR2_X2 \AES_ENC/U837  ( .A(\AES_ENC/w1[25] ), .B(\AES_ENC/text_in_r[89] ),.Z(\AES_ENC/n5101 ) );
NAND2_X2 \AES_ENC/U836  ( .A1(\AES_ENC/n5101 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n509 ) );
NAND2_X2 \AES_ENC/U835  ( .A1(\AES_ENC/n508 ), .A2(\AES_ENC/n509 ), .ZN(\AES_ENC/N207 ) );
NAND2_X2 \AES_ENC/U834  ( .A1(\AES_ENC/sa01_next [2]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n505 ) );
XOR2_X2 \AES_ENC/U833  ( .A(\AES_ENC/w1[26] ), .B(\AES_ENC/text_in_r[90] ),.Z(\AES_ENC/n507 ) );
NAND2_X2 \AES_ENC/U832  ( .A1(\AES_ENC/n507 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n506 ) );
NAND2_X2 \AES_ENC/U831  ( .A1(\AES_ENC/n505 ), .A2(\AES_ENC/n506 ), .ZN(\AES_ENC/N208 ) );
NAND2_X2 \AES_ENC/U830  ( .A1(\AES_ENC/sa01_next [3]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n5021 ) );
XOR2_X2 \AES_ENC/U829  ( .A(\AES_ENC/w1[27] ), .B(\AES_ENC/text_in_r[91] ),.Z(\AES_ENC/n504 ) );
NAND2_X2 \AES_ENC/U828  ( .A1(\AES_ENC/n504 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n503 ) );
NAND2_X2 \AES_ENC/U827  ( .A1(\AES_ENC/n5021 ), .A2(\AES_ENC/n503 ), .ZN(\AES_ENC/N209 ) );
NAND2_X2 \AES_ENC/U826  ( .A1(\AES_ENC/sa01_next [4]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4990 ) );
XOR2_X2 \AES_ENC/U825  ( .A(\AES_ENC/w1[28] ), .B(\AES_ENC/text_in_r[92] ),.Z(\AES_ENC/n5010 ) );
NAND2_X2 \AES_ENC/U824  ( .A1(\AES_ENC/n5010 ), .A2(\AES_ENC/n1243 ), .ZN(\AES_ENC/n5000 ) );
NAND2_X2 \AES_ENC/U823  ( .A1(\AES_ENC/n4990 ), .A2(\AES_ENC/n5000 ), .ZN(\AES_ENC/N210 ) );
NAND2_X2 \AES_ENC/U822  ( .A1(\AES_ENC/sa01_next [5]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4960 ) );
XOR2_X2 \AES_ENC/U821  ( .A(\AES_ENC/w1[29] ), .B(\AES_ENC/text_in_r[93] ),.Z(\AES_ENC/n4980 ) );
NAND2_X2 \AES_ENC/U820  ( .A1(\AES_ENC/n4980 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4970 ) );
NAND2_X2 \AES_ENC/U819  ( .A1(\AES_ENC/n4960 ), .A2(\AES_ENC/n4970 ), .ZN(\AES_ENC/N211 ) );
NAND2_X2 \AES_ENC/U818  ( .A1(\AES_ENC/sa01_next [6]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4930 ) );
XOR2_X2 \AES_ENC/U817  ( .A(\AES_ENC/w1[30] ), .B(\AES_ENC/text_in_r[94] ),.Z(\AES_ENC/n4950 ) );
NAND2_X2 \AES_ENC/U816  ( .A1(\AES_ENC/n4950 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4940 ) );
NAND2_X2 \AES_ENC/U815  ( .A1(\AES_ENC/n4930 ), .A2(\AES_ENC/n4940 ), .ZN(\AES_ENC/N212 ) );
NAND2_X2 \AES_ENC/U814  ( .A1(\AES_ENC/sa01_next [7]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4900 ) );
XOR2_X2 \AES_ENC/U813  ( .A(\AES_ENC/w1[31] ), .B(\AES_ENC/text_in_r[95] ),.Z(\AES_ENC/n4920 ) );
NAND2_X2 \AES_ENC/U812  ( .A1(\AES_ENC/n4920 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4911 ) );
NAND2_X2 \AES_ENC/U811  ( .A1(\AES_ENC/n4900 ), .A2(\AES_ENC/n4911 ), .ZN(\AES_ENC/N213 ) );
NAND2_X2 \AES_ENC/U810  ( .A1(\AES_ENC/sa30_next [0]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4870 ) );
XOR2_X2 \AES_ENC/U809  ( .A(\AES_ENC/w0[0] ), .B(\AES_ENC/text_in_r[96] ),.Z(\AES_ENC/n4890 ) );
NAND2_X2 \AES_ENC/U808  ( .A1(\AES_ENC/n4890 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4880 ) );
NAND2_X2 \AES_ENC/U807  ( .A1(\AES_ENC/n4870 ), .A2(\AES_ENC/n4880 ), .ZN(\AES_ENC/N222 ) );
NAND2_X2 \AES_ENC/U806  ( .A1(\AES_ENC/sa30_next [1]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4840 ) );
XOR2_X2 \AES_ENC/U805  ( .A(\AES_ENC/w0[1] ), .B(\AES_ENC/text_in_r[97] ),.Z(\AES_ENC/n4860 ) );
NAND2_X2 \AES_ENC/U804  ( .A1(\AES_ENC/n4860 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4850 ) );
NAND2_X2 \AES_ENC/U803  ( .A1(\AES_ENC/n4840 ), .A2(\AES_ENC/n4850 ), .ZN(\AES_ENC/N223 ) );
NAND2_X2 \AES_ENC/U802  ( .A1(\AES_ENC/sa30_next [2]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4811 ) );
XOR2_X2 \AES_ENC/U801  ( .A(\AES_ENC/w0[2] ), .B(\AES_ENC/text_in_r[98] ),.Z(\AES_ENC/n4830 ) );
NAND2_X2 \AES_ENC/U800  ( .A1(\AES_ENC/n4830 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4820 ) );
NAND2_X2 \AES_ENC/U799  ( .A1(\AES_ENC/n4811 ), .A2(\AES_ENC/n4820 ), .ZN(\AES_ENC/N224 ) );
NAND2_X2 \AES_ENC/U798  ( .A1(\AES_ENC/sa30_next [3]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4780 ) );
XOR2_X2 \AES_ENC/U797  ( .A(\AES_ENC/w0[3] ), .B(\AES_ENC/text_in_r[99] ),.Z(\AES_ENC/n4800 ) );
NAND2_X2 \AES_ENC/U796  ( .A1(\AES_ENC/n4800 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4790 ) );
NAND2_X2 \AES_ENC/U795  ( .A1(\AES_ENC/n4780 ), .A2(\AES_ENC/n4790 ), .ZN(\AES_ENC/N225 ) );
NAND2_X2 \AES_ENC/U794  ( .A1(\AES_ENC/sa30_next [4]), .A2(\AES_ENC/n1253 ),.ZN(\AES_ENC/n4750 ) );
XOR2_X2 \AES_ENC/U793  ( .A(\AES_ENC/w0[4] ), .B(\AES_ENC/text_in_r[100] ),.Z(\AES_ENC/n4770 ) );
NAND2_X2 \AES_ENC/U792  ( .A1(\AES_ENC/n4770 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4760 ) );
NAND2_X2 \AES_ENC/U791  ( .A1(\AES_ENC/n4750 ), .A2(\AES_ENC/n4760 ), .ZN(\AES_ENC/N226 ) );
NAND2_X2 \AES_ENC/U790  ( .A1(\AES_ENC/sa30_next [5]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4720 ) );
XOR2_X2 \AES_ENC/U789  ( .A(\AES_ENC/w0[5] ), .B(\AES_ENC/text_in_r[101] ),.Z(\AES_ENC/n4740 ) );
NAND2_X2 \AES_ENC/U788  ( .A1(\AES_ENC/n4740 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4730 ) );
NAND2_X2 \AES_ENC/U787  ( .A1(\AES_ENC/n4720 ), .A2(\AES_ENC/n4730 ), .ZN(\AES_ENC/N227 ) );
NAND2_X2 \AES_ENC/U786  ( .A1(\AES_ENC/sa30_next [6]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4690 ) );
XOR2_X2 \AES_ENC/U785  ( .A(\AES_ENC/w0[6] ), .B(\AES_ENC/text_in_r[102] ),.Z(\AES_ENC/n4711 ) );
NAND2_X2 \AES_ENC/U784  ( .A1(\AES_ENC/n4711 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4700 ) );
NAND2_X2 \AES_ENC/U783  ( .A1(\AES_ENC/n4690 ), .A2(\AES_ENC/n4700 ), .ZN(\AES_ENC/N228 ) );
NAND2_X2 \AES_ENC/U782  ( .A1(\AES_ENC/sa30_next [7]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4660 ) );
XOR2_X2 \AES_ENC/U781  ( .A(\AES_ENC/w0[7] ), .B(\AES_ENC/text_in_r[103] ),.Z(\AES_ENC/n4680 ) );
NAND2_X2 \AES_ENC/U780  ( .A1(\AES_ENC/n4680 ), .A2(\AES_ENC/n1244 ), .ZN(\AES_ENC/n4670 ) );
NAND2_X2 \AES_ENC/U779  ( .A1(\AES_ENC/n4660 ), .A2(\AES_ENC/n4670 ), .ZN(\AES_ENC/N229 ) );
NAND2_X2 \AES_ENC/U778  ( .A1(\AES_ENC/sa20_next [0]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4630 ) );
XOR2_X2 \AES_ENC/U777  ( .A(\AES_ENC/w0[8] ), .B(\AES_ENC/text_in_r[104] ),.Z(\AES_ENC/n4650 ) );
NAND2_X2 \AES_ENC/U776  ( .A1(\AES_ENC/n4650 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4640 ) );
NAND2_X2 \AES_ENC/U775  ( .A1(\AES_ENC/n4630 ), .A2(\AES_ENC/n4640 ), .ZN(\AES_ENC/N238 ) );
NAND2_X2 \AES_ENC/U774  ( .A1(\AES_ENC/sa20_next [1]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4600 ) );
XOR2_X2 \AES_ENC/U773  ( .A(\AES_ENC/w0[9] ), .B(\AES_ENC/text_in_r[105] ),.Z(\AES_ENC/n4620 ) );
NAND2_X2 \AES_ENC/U772  ( .A1(\AES_ENC/n4620 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4611 ) );
NAND2_X2 \AES_ENC/U771  ( .A1(\AES_ENC/n4600 ), .A2(\AES_ENC/n4611 ), .ZN(\AES_ENC/N239 ) );
NAND2_X2 \AES_ENC/U770  ( .A1(\AES_ENC/sa20_next [2]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4570 ) );
XOR2_X2 \AES_ENC/U769  ( .A(\AES_ENC/w0[10] ), .B(\AES_ENC/text_in_r[106] ),.Z(\AES_ENC/n4590 ) );
NAND2_X2 \AES_ENC/U768  ( .A1(\AES_ENC/n4590 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4580 ) );
NAND2_X2 \AES_ENC/U767  ( .A1(\AES_ENC/n4570 ), .A2(\AES_ENC/n4580 ), .ZN(\AES_ENC/N240 ) );
NAND2_X2 \AES_ENC/U766  ( .A1(\AES_ENC/sa20_next [3]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4540 ) );
XOR2_X2 \AES_ENC/U765  ( .A(\AES_ENC/w0[11] ), .B(\AES_ENC/text_in_r[107] ),.Z(\AES_ENC/n4560 ) );
NAND2_X2 \AES_ENC/U764  ( .A1(\AES_ENC/n4560 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4550 ) );
NAND2_X2 \AES_ENC/U763  ( .A1(\AES_ENC/n4540 ), .A2(\AES_ENC/n4550 ), .ZN(\AES_ENC/N241 ) );
NAND2_X2 \AES_ENC/U762  ( .A1(\AES_ENC/sa20_next [4]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4510 ) );
XOR2_X2 \AES_ENC/U761  ( .A(\AES_ENC/w0[12] ), .B(\AES_ENC/text_in_r[108] ),.Z(\AES_ENC/n4530 ) );
NAND2_X2 \AES_ENC/U760  ( .A1(\AES_ENC/n4530 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4520 ) );
NAND2_X2 \AES_ENC/U759  ( .A1(\AES_ENC/n4510 ), .A2(\AES_ENC/n4520 ), .ZN(\AES_ENC/N242 ) );
NAND2_X2 \AES_ENC/U758  ( .A1(\AES_ENC/sa20_next [5]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4480 ) );
XOR2_X2 \AES_ENC/U757  ( .A(\AES_ENC/w0[13] ), .B(\AES_ENC/text_in_r[109] ),.Z(\AES_ENC/n4500 ) );
NAND2_X2 \AES_ENC/U756  ( .A1(\AES_ENC/n4500 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4490 ) );
NAND2_X2 \AES_ENC/U755  ( .A1(\AES_ENC/n4480 ), .A2(\AES_ENC/n4490 ), .ZN(\AES_ENC/N243 ) );
NAND2_X2 \AES_ENC/U754  ( .A1(\AES_ENC/sa20_next [6]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4450 ) );
XOR2_X2 \AES_ENC/U753  ( .A(\AES_ENC/w0[14] ), .B(\AES_ENC/text_in_r[110] ),.Z(\AES_ENC/n4470 ) );
NAND2_X2 \AES_ENC/U752  ( .A1(\AES_ENC/n4470 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4460 ) );
NAND2_X2 \AES_ENC/U751  ( .A1(\AES_ENC/n4450 ), .A2(\AES_ENC/n4460 ), .ZN(\AES_ENC/N244 ) );
NAND2_X2 \AES_ENC/U750  ( .A1(\AES_ENC/sa20_next [7]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4420 ) );
XOR2_X2 \AES_ENC/U749  ( .A(\AES_ENC/w0[15] ), .B(\AES_ENC/text_in_r[111] ),.Z(\AES_ENC/n4440 ) );
NAND2_X2 \AES_ENC/U748  ( .A1(\AES_ENC/n4440 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4430 ) );
NAND2_X2 \AES_ENC/U747  ( .A1(\AES_ENC/n4420 ), .A2(\AES_ENC/n4430 ), .ZN(\AES_ENC/N245 ) );
NAND2_X2 \AES_ENC/U746  ( .A1(\AES_ENC/sa10_next [0]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4390 ) );
XOR2_X2 \AES_ENC/U745  ( .A(\AES_ENC/w0[16] ), .B(\AES_ENC/text_in_r[112] ),.Z(\AES_ENC/n4410 ) );
NAND2_X2 \AES_ENC/U744  ( .A1(\AES_ENC/n4410 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4400 ) );
NAND2_X2 \AES_ENC/U743  ( .A1(\AES_ENC/n4390 ), .A2(\AES_ENC/n4400 ), .ZN(\AES_ENC/N254 ) );
NAND2_X2 \AES_ENC/U742  ( .A1(\AES_ENC/sa10_next [1]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4360 ) );
XOR2_X2 \AES_ENC/U741  ( .A(\AES_ENC/w0[17] ), .B(\AES_ENC/text_in_r[113] ),.Z(\AES_ENC/n4380 ) );
NAND2_X2 \AES_ENC/U740  ( .A1(\AES_ENC/n4380 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4370 ) );
NAND2_X2 \AES_ENC/U739  ( .A1(\AES_ENC/n4360 ), .A2(\AES_ENC/n4370 ), .ZN(\AES_ENC/N255 ) );
NAND2_X2 \AES_ENC/U738  ( .A1(\AES_ENC/sa10_next [2]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4330 ) );
XOR2_X2 \AES_ENC/U737  ( .A(\AES_ENC/w0[18] ), .B(\AES_ENC/text_in_r[114] ),.Z(\AES_ENC/n4350 ) );
NAND2_X2 \AES_ENC/U736  ( .A1(\AES_ENC/n4350 ), .A2(\AES_ENC/n1245 ), .ZN(\AES_ENC/n4340 ) );
NAND2_X2 \AES_ENC/U735  ( .A1(\AES_ENC/n4330 ), .A2(\AES_ENC/n4340 ), .ZN(\AES_ENC/N256 ) );
NAND2_X2 \AES_ENC/U734  ( .A1(\AES_ENC/sa10_next [3]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4300 ) );
XOR2_X2 \AES_ENC/U733  ( .A(\AES_ENC/w0[19] ), .B(\AES_ENC/text_in_r[115] ),.Z(\AES_ENC/n4320 ) );
NAND2_X2 \AES_ENC/U732  ( .A1(\AES_ENC/n4320 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4310 ) );
NAND2_X2 \AES_ENC/U731  ( .A1(\AES_ENC/n4300 ), .A2(\AES_ENC/n4310 ), .ZN(\AES_ENC/N257 ) );
NAND2_X2 \AES_ENC/U730  ( .A1(\AES_ENC/sa10_next [4]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4270 ) );
XOR2_X2 \AES_ENC/U729  ( .A(\AES_ENC/w0[20] ), .B(\AES_ENC/text_in_r[116] ),.Z(\AES_ENC/n4290 ) );
NAND2_X2 \AES_ENC/U728  ( .A1(\AES_ENC/n4290 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4280 ) );
NAND2_X2 \AES_ENC/U727  ( .A1(\AES_ENC/n4270 ), .A2(\AES_ENC/n4280 ), .ZN(\AES_ENC/N258 ) );
NAND2_X2 \AES_ENC/U726  ( .A1(\AES_ENC/sa10_next [5]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4240 ) );
XOR2_X2 \AES_ENC/U725  ( .A(\AES_ENC/w0[21] ), .B(\AES_ENC/text_in_r[117] ),.Z(\AES_ENC/n4260 ) );
NAND2_X2 \AES_ENC/U724  ( .A1(\AES_ENC/n4260 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4250 ) );
NAND2_X2 \AES_ENC/U723  ( .A1(\AES_ENC/n4240 ), .A2(\AES_ENC/n4250 ), .ZN(\AES_ENC/N259 ) );
NAND2_X2 \AES_ENC/U722  ( .A1(\AES_ENC/sa10_next [6]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4210 ) );
XOR2_X2 \AES_ENC/U721  ( .A(\AES_ENC/w0[22] ), .B(\AES_ENC/text_in_r[118] ),.Z(\AES_ENC/n4230 ) );
NAND2_X2 \AES_ENC/U720  ( .A1(\AES_ENC/n4230 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4220 ) );
NAND2_X2 \AES_ENC/U719  ( .A1(\AES_ENC/n4210 ), .A2(\AES_ENC/n4220 ), .ZN(\AES_ENC/N260 ) );
NAND2_X2 \AES_ENC/U718  ( .A1(\AES_ENC/sa10_next [7]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4180 ) );
XOR2_X2 \AES_ENC/U717  ( .A(\AES_ENC/w0[23] ), .B(\AES_ENC/text_in_r[119] ),.Z(\AES_ENC/n4200 ) );
NAND2_X2 \AES_ENC/U716  ( .A1(\AES_ENC/n4200 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4190 ) );
NAND2_X2 \AES_ENC/U715  ( .A1(\AES_ENC/n4180 ), .A2(\AES_ENC/n4190 ), .ZN(\AES_ENC/N261 ) );
NAND2_X2 \AES_ENC/U714  ( .A1(\AES_ENC/sa00_next [0]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4150 ) );
XOR2_X2 \AES_ENC/U713  ( .A(\AES_ENC/w0[24] ), .B(\AES_ENC/text_in_r[120] ),.Z(\AES_ENC/n4170 ) );
NAND2_X2 \AES_ENC/U712  ( .A1(\AES_ENC/n4170 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4160 ) );
NAND2_X2 \AES_ENC/U711  ( .A1(\AES_ENC/n4150 ), .A2(\AES_ENC/n4160 ), .ZN(\AES_ENC/N270 ) );
NAND2_X2 \AES_ENC/U710  ( .A1(\AES_ENC/sa00_next [1]), .A2(\AES_ENC/n1254 ),.ZN(\AES_ENC/n4120 ) );
XOR2_X2 \AES_ENC/U709  ( .A(\AES_ENC/w0[25] ), .B(\AES_ENC/text_in_r[121] ),.Z(\AES_ENC/n4140 ) );
NAND2_X2 \AES_ENC/U708  ( .A1(\AES_ENC/n4140 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4130 ) );
NAND2_X2 \AES_ENC/U707  ( .A1(\AES_ENC/n4120 ), .A2(\AES_ENC/n4130 ), .ZN(\AES_ENC/N271 ) );
NAND2_X2 \AES_ENC/U706  ( .A1(\AES_ENC/sa00_next [2]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n4090 ) );
XOR2_X2 \AES_ENC/U705  ( .A(\AES_ENC/w0[26] ), .B(\AES_ENC/text_in_r[122] ),.Z(\AES_ENC/n4110 ) );
NAND2_X2 \AES_ENC/U704  ( .A1(\AES_ENC/n4110 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4100 ) );
NAND2_X2 \AES_ENC/U703  ( .A1(\AES_ENC/n4090 ), .A2(\AES_ENC/n4100 ), .ZN(\AES_ENC/N272 ) );
NAND2_X2 \AES_ENC/U702  ( .A1(\AES_ENC/sa00_next [3]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n4060 ) );
XOR2_X2 \AES_ENC/U701  ( .A(\AES_ENC/w0[27] ), .B(\AES_ENC/text_in_r[123] ),.Z(\AES_ENC/n4080 ) );
NAND2_X2 \AES_ENC/U700  ( .A1(\AES_ENC/n4080 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4070 ) );
NAND2_X2 \AES_ENC/U699  ( .A1(\AES_ENC/n4060 ), .A2(\AES_ENC/n4070 ), .ZN(\AES_ENC/N273 ) );
NAND2_X2 \AES_ENC/U698  ( .A1(\AES_ENC/sa00_next [4]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n4030 ) );
XOR2_X2 \AES_ENC/U697  ( .A(\AES_ENC/w0[28] ), .B(\AES_ENC/text_in_r[124] ),.Z(\AES_ENC/n4050 ) );
NAND2_X2 \AES_ENC/U696  ( .A1(\AES_ENC/n4050 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4040 ) );
NAND2_X2 \AES_ENC/U695  ( .A1(\AES_ENC/n4030 ), .A2(\AES_ENC/n4040 ), .ZN(\AES_ENC/N274 ) );
NAND2_X2 \AES_ENC/U694  ( .A1(\AES_ENC/sa00_next [5]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n4000 ) );
XOR2_X2 \AES_ENC/U693  ( .A(\AES_ENC/w0[29] ), .B(\AES_ENC/text_in_r[125] ),.Z(\AES_ENC/n4020 ) );
NAND2_X2 \AES_ENC/U692  ( .A1(\AES_ENC/n4020 ), .A2(\AES_ENC/n1246 ), .ZN(\AES_ENC/n4010 ) );
NAND2_X2 \AES_ENC/U691  ( .A1(\AES_ENC/n4000 ), .A2(\AES_ENC/n4010 ), .ZN(\AES_ENC/N275 ) );
NAND2_X2 \AES_ENC/U690  ( .A1(\AES_ENC/sa00_next [6]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3970 ) );
XOR2_X2 \AES_ENC/U689  ( .A(\AES_ENC/w0[30] ), .B(\AES_ENC/text_in_r[126] ),.Z(\AES_ENC/n3990 ) );
NAND2_X2 \AES_ENC/U688  ( .A1(\AES_ENC/n3990 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3980 ) );
NAND2_X2 \AES_ENC/U687  ( .A1(\AES_ENC/n3970 ), .A2(\AES_ENC/n3980 ), .ZN(\AES_ENC/N276 ) );
NAND2_X2 \AES_ENC/U686  ( .A1(\AES_ENC/sa00_next [7]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3940 ) );
XOR2_X2 \AES_ENC/U685  ( .A(\AES_ENC/w0[31] ), .B(\AES_ENC/text_in_r[127] ),.Z(\AES_ENC/n3960 ) );
NAND2_X2 \AES_ENC/U684  ( .A1(\AES_ENC/n3960 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3950 ) );
NAND2_X2 \AES_ENC/U683  ( .A1(\AES_ENC/n3940 ), .A2(\AES_ENC/n3950 ), .ZN(\AES_ENC/N277 ) );
NAND2_X2 \AES_ENC/U682  ( .A1(\AES_ENC/sa33_next [0]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3910 ) );
XOR2_X2 \AES_ENC/U681  ( .A(\AES_ENC/w3[0] ), .B(\AES_ENC/text_in_r[0] ),.Z(\AES_ENC/n3930 ) );
NAND2_X2 \AES_ENC/U680  ( .A1(\AES_ENC/n3930 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3920 ) );
NAND2_X2 \AES_ENC/U679  ( .A1(\AES_ENC/n3910 ), .A2(\AES_ENC/n3920 ), .ZN(\AES_ENC/N30 ) );
NAND2_X2 \AES_ENC/U678  ( .A1(\AES_ENC/sa33_next [1]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3880 ) );
XOR2_X2 \AES_ENC/U677  ( .A(\AES_ENC/w3[1] ), .B(\AES_ENC/text_in_r[1] ),.Z(\AES_ENC/n3900 ) );
NAND2_X2 \AES_ENC/U676  ( .A1(\AES_ENC/n3900 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3890 ) );
NAND2_X2 \AES_ENC/U675  ( .A1(\AES_ENC/n3880 ), .A2(\AES_ENC/n3890 ), .ZN(\AES_ENC/N31 ) );
NAND2_X2 \AES_ENC/U674  ( .A1(\AES_ENC/sa33_next [2]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3850 ) );
XOR2_X2 \AES_ENC/U673  ( .A(\AES_ENC/w3[2] ), .B(\AES_ENC/text_in_r[2] ),.Z(\AES_ENC/n3870 ) );
NAND2_X2 \AES_ENC/U672  ( .A1(\AES_ENC/n3870 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3860 ) );
NAND2_X2 \AES_ENC/U671  ( .A1(\AES_ENC/n3850 ), .A2(\AES_ENC/n3860 ), .ZN(\AES_ENC/N32 ) );
NAND2_X2 \AES_ENC/U670  ( .A1(\AES_ENC/sa33_next [3]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3820 ) );
XOR2_X2 \AES_ENC/U669  ( .A(\AES_ENC/w3[3] ), .B(\AES_ENC/text_in_r[3] ),.Z(\AES_ENC/n3840 ) );
NAND2_X2 \AES_ENC/U668  ( .A1(\AES_ENC/n3840 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3830 ) );
NAND2_X2 \AES_ENC/U667  ( .A1(\AES_ENC/n3820 ), .A2(\AES_ENC/n3830 ), .ZN(\AES_ENC/N33 ) );
NAND2_X2 \AES_ENC/U666  ( .A1(\AES_ENC/sa33_next [4]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3790 ) );
XOR2_X2 \AES_ENC/U665  ( .A(\AES_ENC/w3[4] ), .B(\AES_ENC/text_in_r[4] ),.Z(\AES_ENC/n3810 ) );
NAND2_X2 \AES_ENC/U664  ( .A1(\AES_ENC/n3810 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3800 ) );
NAND2_X2 \AES_ENC/U663  ( .A1(\AES_ENC/n3790 ), .A2(\AES_ENC/n3800 ), .ZN(\AES_ENC/N34 ) );
NAND2_X2 \AES_ENC/U662  ( .A1(\AES_ENC/sa33_next [5]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3760 ) );
XOR2_X2 \AES_ENC/U661  ( .A(\AES_ENC/w3[5] ), .B(\AES_ENC/text_in_r[5] ),.Z(\AES_ENC/n3780 ) );
NAND2_X2 \AES_ENC/U660  ( .A1(\AES_ENC/n3780 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3770 ) );
NAND2_X2 \AES_ENC/U659  ( .A1(\AES_ENC/n3760 ), .A2(\AES_ENC/n3770 ), .ZN(\AES_ENC/N35 ) );
NAND2_X2 \AES_ENC/U658  ( .A1(\AES_ENC/sa33_next [6]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n373 ) );
XOR2_X2 \AES_ENC/U657  ( .A(\AES_ENC/w3[6] ), .B(\AES_ENC/text_in_r[6] ),.Z(\AES_ENC/n3750 ) );
NAND2_X2 \AES_ENC/U656  ( .A1(\AES_ENC/n3750 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n3740 ) );
NAND2_X2 \AES_ENC/U655  ( .A1(\AES_ENC/n373 ), .A2(\AES_ENC/n3740 ), .ZN(\AES_ENC/N36 ) );
NAND2_X2 \AES_ENC/U654  ( .A1(\AES_ENC/sa33_next [7]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n3701 ) );
XOR2_X2 \AES_ENC/U653  ( .A(\AES_ENC/w3[7] ), .B(\AES_ENC/text_in_r[7] ),.Z(\AES_ENC/n372 ) );
NAND2_X2 \AES_ENC/U652  ( .A1(\AES_ENC/n372 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n371 ) );
NAND2_X2 \AES_ENC/U651  ( .A1(\AES_ENC/n3701 ), .A2(\AES_ENC/n371 ), .ZN(\AES_ENC/N37 ) );
XOR2_X2 \AES_ENC/U650  ( .A(\AES_ENC/w0[31] ), .B(\AES_ENC/sa00_sub[7] ),.Z(\AES_ENC/N374 ) );
XOR2_X2 \AES_ENC/U649  ( .A(\AES_ENC/w0[30] ), .B(\AES_ENC/sa00_sub[6] ),.Z(\AES_ENC/N375 ) );
XOR2_X2 \AES_ENC/U648  ( .A(\AES_ENC/w0[29] ), .B(\AES_ENC/sa00_sub[5] ),.Z(\AES_ENC/N376 ) );
XOR2_X2 \AES_ENC/U647  ( .A(\AES_ENC/w0[28] ), .B(\AES_ENC/sa00_sub[4] ),.Z(\AES_ENC/N377 ) );
XOR2_X2 \AES_ENC/U646  ( .A(\AES_ENC/w0[27] ), .B(\AES_ENC/sa00_sub[3] ),.Z(\AES_ENC/N378 ) );
XOR2_X2 \AES_ENC/U645  ( .A(\AES_ENC/w0[26] ), .B(\AES_ENC/sa00_sub[2] ),.Z(\AES_ENC/N379 ) );
XOR2_X2 \AES_ENC/U644  ( .A(\AES_ENC/w0[25] ), .B(\AES_ENC/sa00_sub[1] ),.Z(\AES_ENC/N380 ) );
XOR2_X2 \AES_ENC/U643  ( .A(\AES_ENC/w0[24] ), .B(\AES_ENC/sa00_sub[0] ),.Z(\AES_ENC/N381 ) );
XOR2_X2 \AES_ENC/U642  ( .A(\AES_ENC/w1[31] ), .B(\AES_ENC/sa01_sub[7] ),.Z(\AES_ENC/N382 ) );
XOR2_X2 \AES_ENC/U641  ( .A(\AES_ENC/w1[30] ), .B(\AES_ENC/sa01_sub[6] ),.Z(\AES_ENC/N383 ) );
XOR2_X2 \AES_ENC/U640  ( .A(\AES_ENC/w1[29] ), .B(\AES_ENC/sa01_sub[5] ),.Z(\AES_ENC/N384 ) );
XOR2_X2 \AES_ENC/U639  ( .A(\AES_ENC/w1[28] ), .B(\AES_ENC/sa01_sub[4] ),.Z(\AES_ENC/N385 ) );
XOR2_X2 \AES_ENC/U638  ( .A(\AES_ENC/w1[27] ), .B(\AES_ENC/sa01_sub[3] ),.Z(\AES_ENC/N386 ) );
XOR2_X2 \AES_ENC/U637  ( .A(\AES_ENC/w1[26] ), .B(\AES_ENC/sa01_sub[2] ),.Z(\AES_ENC/N387 ) );
XOR2_X2 \AES_ENC/U636  ( .A(\AES_ENC/w1[25] ), .B(\AES_ENC/sa01_sub[1] ),.Z(\AES_ENC/N388 ) );
XOR2_X2 \AES_ENC/U635  ( .A(\AES_ENC/w1[24] ), .B(\AES_ENC/sa01_sub[0] ),.Z(\AES_ENC/N389 ) );
XOR2_X2 \AES_ENC/U634  ( .A(\AES_ENC/w2[31] ), .B(\AES_ENC/sa02_sub[7] ),.Z(\AES_ENC/N390 ) );
XOR2_X2 \AES_ENC/U633  ( .A(\AES_ENC/w2[30] ), .B(\AES_ENC/sa02_sub[6] ),.Z(\AES_ENC/N391 ) );
XOR2_X2 \AES_ENC/U632  ( .A(\AES_ENC/w2[29] ), .B(\AES_ENC/sa02_sub[5] ),.Z(\AES_ENC/N392 ) );
XOR2_X2 \AES_ENC/U631  ( .A(\AES_ENC/w2[28] ), .B(\AES_ENC/sa02_sub[4] ),.Z(\AES_ENC/N393 ) );
XOR2_X2 \AES_ENC/U630  ( .A(\AES_ENC/w2[27] ), .B(\AES_ENC/sa02_sub[3] ),.Z(\AES_ENC/N394 ) );
XOR2_X2 \AES_ENC/U629  ( .A(\AES_ENC/w2[26] ), .B(\AES_ENC/sa02_sub[2] ),.Z(\AES_ENC/N395 ) );
XOR2_X2 \AES_ENC/U628  ( .A(\AES_ENC/w2[25] ), .B(\AES_ENC/sa02_sub[1] ),.Z(\AES_ENC/N396 ) );
XOR2_X2 \AES_ENC/U627  ( .A(\AES_ENC/w2[24] ), .B(\AES_ENC/sa02_sub[0] ),.Z(\AES_ENC/N397 ) );
XOR2_X2 \AES_ENC/U626  ( .A(\AES_ENC/w3[31] ), .B(\AES_ENC/sa03_sub[7] ),.Z(\AES_ENC/N398 ) );
XOR2_X2 \AES_ENC/U625  ( .A(\AES_ENC/w3[30] ), .B(\AES_ENC/sa03_sub[6] ),.Z(\AES_ENC/N399 ) );
XOR2_X2 \AES_ENC/U624  ( .A(\AES_ENC/w3[29] ), .B(\AES_ENC/sa03_sub[5] ),.Z(\AES_ENC/N400 ) );
XOR2_X2 \AES_ENC/U623  ( .A(\AES_ENC/w3[28] ), .B(\AES_ENC/sa03_sub[4] ),.Z(\AES_ENC/N401 ) );
XOR2_X2 \AES_ENC/U622  ( .A(\AES_ENC/w3[27] ), .B(\AES_ENC/sa03_sub[3] ),.Z(\AES_ENC/N402 ) );
XOR2_X2 \AES_ENC/U621  ( .A(\AES_ENC/w3[26] ), .B(\AES_ENC/sa03_sub[2] ),.Z(\AES_ENC/N403 ) );
XOR2_X2 \AES_ENC/U620  ( .A(\AES_ENC/w3[25] ), .B(\AES_ENC/sa03_sub[1] ),.Z(\AES_ENC/N404 ) );
XOR2_X2 \AES_ENC/U619  ( .A(\AES_ENC/w3[24] ), .B(\AES_ENC/sa03_sub[0] ),.Z(\AES_ENC/N405 ) );
XOR2_X2 \AES_ENC/U618  ( .A(\AES_ENC/w0[23] ), .B(\AES_ENC/sa11_sub[7] ),.Z(\AES_ENC/N406 ) );
XOR2_X2 \AES_ENC/U617  ( .A(\AES_ENC/w0[22] ), .B(\AES_ENC/sa11_sub[6] ),.Z(\AES_ENC/N407 ) );
XOR2_X2 \AES_ENC/U616  ( .A(\AES_ENC/w0[21] ), .B(\AES_ENC/sa11_sub[5] ),.Z(\AES_ENC/N408 ) );
XOR2_X2 \AES_ENC/U615  ( .A(\AES_ENC/w0[20] ), .B(\AES_ENC/sa11_sub[4] ),.Z(\AES_ENC/N409 ) );
XOR2_X2 \AES_ENC/U614  ( .A(\AES_ENC/w0[19] ), .B(\AES_ENC/sa11_sub[3] ),.Z(\AES_ENC/N410 ) );
XOR2_X2 \AES_ENC/U613  ( .A(\AES_ENC/w0[18] ), .B(\AES_ENC/sa11_sub[2] ),.Z(\AES_ENC/N411 ) );
XOR2_X2 \AES_ENC/U612  ( .A(\AES_ENC/w0[17] ), .B(\AES_ENC/sa11_sub[1] ),.Z(\AES_ENC/N412 ) );
XOR2_X2 \AES_ENC/U611  ( .A(\AES_ENC/w0[16] ), .B(\AES_ENC/sa11_sub[0] ),.Z(\AES_ENC/N413 ) );
XOR2_X2 \AES_ENC/U610  ( .A(\AES_ENC/w1[23] ), .B(\AES_ENC/sa12_sub[7] ),.Z(\AES_ENC/N414 ) );
XOR2_X2 \AES_ENC/U609  ( .A(\AES_ENC/w1[22] ), .B(\AES_ENC/sa12_sub[6] ),.Z(\AES_ENC/N415 ) );
XOR2_X2 \AES_ENC/U608  ( .A(\AES_ENC/w1[21] ), .B(\AES_ENC/sa12_sub[5] ),.Z(\AES_ENC/N416 ) );
XOR2_X2 \AES_ENC/U607  ( .A(\AES_ENC/w1[20] ), .B(\AES_ENC/sa12_sub[4] ),.Z(\AES_ENC/N417 ) );
XOR2_X2 \AES_ENC/U606  ( .A(\AES_ENC/w1[19] ), .B(\AES_ENC/sa12_sub[3] ),.Z(\AES_ENC/N418 ) );
XOR2_X2 \AES_ENC/U605  ( .A(\AES_ENC/w1[18] ), .B(\AES_ENC/sa12_sub[2] ),.Z(\AES_ENC/N419 ) );
XOR2_X2 \AES_ENC/U604  ( .A(\AES_ENC/w1[17] ), .B(\AES_ENC/sa12_sub[1] ),.Z(\AES_ENC/N420 ) );
XOR2_X2 \AES_ENC/U603  ( .A(\AES_ENC/w1[16] ), .B(\AES_ENC/sa12_sub[0] ),.Z(\AES_ENC/N421 ) );
XOR2_X2 \AES_ENC/U602  ( .A(\AES_ENC/w2[23] ), .B(\AES_ENC/sa13_sub[7] ),.Z(\AES_ENC/N422 ) );
XOR2_X2 \AES_ENC/U601  ( .A(\AES_ENC/w2[22] ), .B(\AES_ENC/sa13_sub[6] ),.Z(\AES_ENC/N423 ) );
XOR2_X2 \AES_ENC/U600  ( .A(\AES_ENC/w2[21] ), .B(\AES_ENC/sa13_sub[5] ),.Z(\AES_ENC/N424 ) );
XOR2_X2 \AES_ENC/U599  ( .A(\AES_ENC/w2[20] ), .B(\AES_ENC/sa13_sub[4] ),.Z(\AES_ENC/N425 ) );
XOR2_X2 \AES_ENC/U598  ( .A(\AES_ENC/w2[19] ), .B(\AES_ENC/sa13_sub[3] ),.Z(\AES_ENC/N426 ) );
XOR2_X2 \AES_ENC/U597  ( .A(\AES_ENC/w2[18] ), .B(\AES_ENC/sa13_sub[2] ),.Z(\AES_ENC/N427 ) );
XOR2_X2 \AES_ENC/U596  ( .A(\AES_ENC/w2[17] ), .B(\AES_ENC/sa13_sub[1] ),.Z(\AES_ENC/N428 ) );
XOR2_X2 \AES_ENC/U595  ( .A(\AES_ENC/w2[16] ), .B(\AES_ENC/sa13_sub[0] ),.Z(\AES_ENC/N429 ) );
XOR2_X2 \AES_ENC/U594  ( .A(\AES_ENC/w3[23] ), .B(\AES_ENC/sa10_sub[7] ),.Z(\AES_ENC/N430 ) );
XOR2_X2 \AES_ENC/U593  ( .A(\AES_ENC/w3[22] ), .B(\AES_ENC/sa10_sub[6] ),.Z(\AES_ENC/N431 ) );
XOR2_X2 \AES_ENC/U592  ( .A(\AES_ENC/w3[21] ), .B(\AES_ENC/sa10_sub[5] ),.Z(\AES_ENC/N432 ) );
XOR2_X2 \AES_ENC/U591  ( .A(\AES_ENC/w3[20] ), .B(\AES_ENC/sa10_sub[4] ),.Z(\AES_ENC/N433 ) );
XOR2_X2 \AES_ENC/U590  ( .A(\AES_ENC/w3[19] ), .B(\AES_ENC/sa10_sub[3] ),.Z(\AES_ENC/N434 ) );
XOR2_X2 \AES_ENC/U589  ( .A(\AES_ENC/w3[18] ), .B(\AES_ENC/sa10_sub[2] ),.Z(\AES_ENC/N435 ) );
XOR2_X2 \AES_ENC/U588  ( .A(\AES_ENC/w3[17] ), .B(\AES_ENC/sa10_sub[1] ),.Z(\AES_ENC/N436 ) );
XOR2_X2 \AES_ENC/U587  ( .A(\AES_ENC/w3[16] ), .B(\AES_ENC/sa10_sub[0] ),.Z(\AES_ENC/N437 ) );
XOR2_X2 \AES_ENC/U586  ( .A(\AES_ENC/w0[15] ), .B(\AES_ENC/sa22_sub[7] ),.Z(\AES_ENC/N438 ) );
XOR2_X2 \AES_ENC/U585  ( .A(\AES_ENC/w0[14] ), .B(\AES_ENC/sa22_sub[6] ),.Z(\AES_ENC/N439 ) );
XOR2_X2 \AES_ENC/U584  ( .A(\AES_ENC/w0[13] ), .B(\AES_ENC/sa22_sub[5] ),.Z(\AES_ENC/N440 ) );
XOR2_X2 \AES_ENC/U583  ( .A(\AES_ENC/w0[12] ), .B(\AES_ENC/sa22_sub[4] ),.Z(\AES_ENC/N441 ) );
XOR2_X2 \AES_ENC/U582  ( .A(\AES_ENC/w0[11] ), .B(\AES_ENC/sa22_sub[3] ),.Z(\AES_ENC/N442 ) );
XOR2_X2 \AES_ENC/U581  ( .A(\AES_ENC/w0[10] ), .B(\AES_ENC/sa22_sub[2] ),.Z(\AES_ENC/N443 ) );
XOR2_X2 \AES_ENC/U580  ( .A(\AES_ENC/w0[9] ), .B(\AES_ENC/sa22_sub[1] ), .Z(\AES_ENC/N444 ) );
XOR2_X2 \AES_ENC/U579  ( .A(\AES_ENC/w0[8] ), .B(\AES_ENC/sa22_sub[0] ), .Z(\AES_ENC/N445 ) );
XOR2_X2 \AES_ENC/U578  ( .A(\AES_ENC/w1[15] ), .B(\AES_ENC/sa23_sub[7] ),.Z(\AES_ENC/N446 ) );
XOR2_X2 \AES_ENC/U577  ( .A(\AES_ENC/w1[14] ), .B(\AES_ENC/sa23_sub[6] ),.Z(\AES_ENC/N447 ) );
XOR2_X2 \AES_ENC/U576  ( .A(\AES_ENC/w1[13] ), .B(\AES_ENC/sa23_sub[5] ),.Z(\AES_ENC/N448 ) );
XOR2_X2 \AES_ENC/U575  ( .A(\AES_ENC/w1[12] ), .B(\AES_ENC/sa23_sub[4] ),.Z(\AES_ENC/N449 ) );
XOR2_X2 \AES_ENC/U574  ( .A(\AES_ENC/w1[11] ), .B(\AES_ENC/sa23_sub[3] ),.Z(\AES_ENC/N450 ) );
XOR2_X2 \AES_ENC/U573  ( .A(\AES_ENC/w1[10] ), .B(\AES_ENC/sa23_sub[2] ),.Z(\AES_ENC/N451 ) );
XOR2_X2 \AES_ENC/U572  ( .A(\AES_ENC/w1[9] ), .B(\AES_ENC/sa23_sub[1] ), .Z(\AES_ENC/N452 ) );
XOR2_X2 \AES_ENC/U571  ( .A(\AES_ENC/w1[8] ), .B(\AES_ENC/sa23_sub[0] ), .Z(\AES_ENC/N453 ) );
XOR2_X2 \AES_ENC/U570  ( .A(\AES_ENC/w2[15] ), .B(\AES_ENC/sa20_sub[7] ),.Z(\AES_ENC/N454 ) );
XOR2_X2 \AES_ENC/U569  ( .A(\AES_ENC/w2[14] ), .B(\AES_ENC/sa20_sub[6] ),.Z(\AES_ENC/N455 ) );
XOR2_X2 \AES_ENC/U568  ( .A(\AES_ENC/w2[13] ), .B(\AES_ENC/sa20_sub[5] ),.Z(\AES_ENC/N456 ) );
XOR2_X2 \AES_ENC/U567  ( .A(\AES_ENC/w2[12] ), .B(\AES_ENC/sa20_sub[4] ),.Z(\AES_ENC/N457 ) );
XOR2_X2 \AES_ENC/U566  ( .A(\AES_ENC/w2[11] ), .B(\AES_ENC/sa20_sub[3] ),.Z(\AES_ENC/N458 ) );
XOR2_X2 \AES_ENC/U565  ( .A(\AES_ENC/w2[10] ), .B(\AES_ENC/sa20_sub[2] ),.Z(\AES_ENC/N459 ) );
NAND2_X2 \AES_ENC/U564  ( .A1(\AES_ENC/sa23_next [0]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n367 ) );
XOR2_X2 \AES_ENC/U563  ( .A(\AES_ENC/w3[8] ), .B(\AES_ENC/text_in_r[8] ),.Z(\AES_ENC/n369 ) );
NAND2_X2 \AES_ENC/U562  ( .A1(\AES_ENC/n369 ), .A2(\AES_ENC/n1247 ), .ZN(\AES_ENC/n368 ) );
NAND2_X2 \AES_ENC/U561  ( .A1(\AES_ENC/n367 ), .A2(\AES_ENC/n368 ), .ZN(\AES_ENC/N46 ) );
XOR2_X2 \AES_ENC/U560  ( .A(\AES_ENC/w2[9] ), .B(\AES_ENC/sa20_sub[1] ), .Z(\AES_ENC/N460 ) );
XOR2_X2 \AES_ENC/U559  ( .A(\AES_ENC/w2[8] ), .B(\AES_ENC/sa20_sub[0] ), .Z(\AES_ENC/N461 ) );
XOR2_X2 \AES_ENC/U558  ( .A(\AES_ENC/w3[15] ), .B(\AES_ENC/sa21_sub[7] ),.Z(\AES_ENC/N462 ) );
XOR2_X2 \AES_ENC/U557  ( .A(\AES_ENC/w3[14] ), .B(\AES_ENC/sa21_sub[6] ),.Z(\AES_ENC/N463 ) );
XOR2_X2 \AES_ENC/U556  ( .A(\AES_ENC/w3[13] ), .B(\AES_ENC/sa21_sub[5] ),.Z(\AES_ENC/N464 ) );
XOR2_X2 \AES_ENC/U555  ( .A(\AES_ENC/w3[12] ), .B(\AES_ENC/sa21_sub[4] ),.Z(\AES_ENC/N465 ) );
XOR2_X2 \AES_ENC/U554  ( .A(\AES_ENC/w3[11] ), .B(\AES_ENC/sa21_sub[3] ),.Z(\AES_ENC/N466 ) );
XOR2_X2 \AES_ENC/U553  ( .A(\AES_ENC/w3[10] ), .B(\AES_ENC/sa21_sub[2] ),.Z(\AES_ENC/N467 ) );
XOR2_X2 \AES_ENC/U552  ( .A(\AES_ENC/w3[9] ), .B(\AES_ENC/sa21_sub[1] ), .Z(\AES_ENC/N468 ) );
XOR2_X2 \AES_ENC/U551  ( .A(\AES_ENC/w3[8] ), .B(\AES_ENC/sa21_sub[0] ), .Z(\AES_ENC/N469 ) );
NAND2_X2 \AES_ENC/U550  ( .A1(\AES_ENC/sa23_next [1]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n364 ) );
XOR2_X2 \AES_ENC/U549  ( .A(\AES_ENC/w3[9] ), .B(\AES_ENC/text_in_r[9] ),.Z(\AES_ENC/n366 ) );
NAND2_X2 \AES_ENC/U548  ( .A1(\AES_ENC/n366 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n365 ) );
NAND2_X2 \AES_ENC/U547  ( .A1(\AES_ENC/n364 ), .A2(\AES_ENC/n365 ), .ZN(\AES_ENC/N47 ) );
XOR2_X2 \AES_ENC/U546  ( .A(\AES_ENC/w0[7] ), .B(\AES_ENC/sa33_sub[7] ), .Z(\AES_ENC/N470 ) );
XOR2_X2 \AES_ENC/U545  ( .A(\AES_ENC/w0[6] ), .B(\AES_ENC/sa33_sub[6] ), .Z(\AES_ENC/N471 ) );
XOR2_X2 \AES_ENC/U544  ( .A(\AES_ENC/w0[5] ), .B(\AES_ENC/sa33_sub[5] ), .Z(\AES_ENC/N472 ) );
XOR2_X2 \AES_ENC/U543  ( .A(\AES_ENC/w0[4] ), .B(\AES_ENC/sa33_sub[4] ), .Z(\AES_ENC/N473 ) );
XOR2_X2 \AES_ENC/U542  ( .A(\AES_ENC/w0[3] ), .B(\AES_ENC/sa33_sub[3] ), .Z(\AES_ENC/N474 ) );
XOR2_X2 \AES_ENC/U541  ( .A(\AES_ENC/w0[2] ), .B(\AES_ENC/sa33_sub[2] ), .Z(\AES_ENC/N475 ) );
XOR2_X2 \AES_ENC/U540  ( .A(\AES_ENC/w0[1] ), .B(\AES_ENC/sa33_sub[1] ), .Z(\AES_ENC/N476 ) );
XOR2_X2 \AES_ENC/U539  ( .A(\AES_ENC/w0[0] ), .B(\AES_ENC/sa33_sub[0] ), .Z(\AES_ENC/N477 ) );
XOR2_X2 \AES_ENC/U538  ( .A(\AES_ENC/w1[7] ), .B(\AES_ENC/sa30_sub[7] ), .Z(\AES_ENC/N478 ) );
XOR2_X2 \AES_ENC/U537  ( .A(\AES_ENC/w1[6] ), .B(\AES_ENC/sa30_sub[6] ), .Z(\AES_ENC/N479 ) );
NAND2_X2 \AES_ENC/U536  ( .A1(\AES_ENC/sa23_next [2]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n361 ) );
XOR2_X2 \AES_ENC/U535  ( .A(\AES_ENC/w3[10] ), .B(\AES_ENC/text_in_r[10] ),.Z(\AES_ENC/n363 ) );
NAND2_X2 \AES_ENC/U534  ( .A1(\AES_ENC/n363 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n362 ) );
NAND2_X2 \AES_ENC/U533  ( .A1(\AES_ENC/n361 ), .A2(\AES_ENC/n362 ), .ZN(\AES_ENC/N48 ) );
XOR2_X2 \AES_ENC/U532  ( .A(\AES_ENC/w1[5] ), .B(\AES_ENC/sa30_sub[5] ), .Z(\AES_ENC/N480 ) );
XOR2_X2 \AES_ENC/U531  ( .A(\AES_ENC/w1[4] ), .B(\AES_ENC/sa30_sub[4] ), .Z(\AES_ENC/N481 ) );
XOR2_X2 \AES_ENC/U530  ( .A(\AES_ENC/w1[3] ), .B(\AES_ENC/sa30_sub[3] ), .Z(\AES_ENC/N482 ) );
XOR2_X2 \AES_ENC/U529  ( .A(\AES_ENC/w1[2] ), .B(\AES_ENC/sa30_sub[2] ), .Z(\AES_ENC/N483 ) );
XOR2_X2 \AES_ENC/U528  ( .A(\AES_ENC/w1[1] ), .B(\AES_ENC/sa30_sub[1] ), .Z(\AES_ENC/N484 ) );
XOR2_X2 \AES_ENC/U527  ( .A(\AES_ENC/w1[0] ), .B(\AES_ENC/sa30_sub[0] ), .Z(\AES_ENC/N485 ) );
XOR2_X2 \AES_ENC/U526  ( .A(\AES_ENC/w2[7] ), .B(\AES_ENC/sa31_sub[7] ), .Z(\AES_ENC/N486 ) );
XOR2_X2 \AES_ENC/U525  ( .A(\AES_ENC/w2[6] ), .B(\AES_ENC/sa31_sub[6] ), .Z(\AES_ENC/N487 ) );
XOR2_X2 \AES_ENC/U524  ( .A(\AES_ENC/w2[5] ), .B(\AES_ENC/sa31_sub[5] ), .Z(\AES_ENC/N488 ) );
XOR2_X2 \AES_ENC/U523  ( .A(\AES_ENC/w2[4] ), .B(\AES_ENC/sa31_sub[4] ), .Z(\AES_ENC/N489 ) );
NAND2_X2 \AES_ENC/U522  ( .A1(\AES_ENC/sa23_next [3]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n358 ) );
XOR2_X2 \AES_ENC/U521  ( .A(\AES_ENC/w3[11] ), .B(\AES_ENC/text_in_r[11] ),.Z(\AES_ENC/n3601 ) );
NAND2_X2 \AES_ENC/U520  ( .A1(\AES_ENC/n3601 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n359 ) );
NAND2_X2 \AES_ENC/U519  ( .A1(\AES_ENC/n358 ), .A2(\AES_ENC/n359 ), .ZN(\AES_ENC/N49 ) );
XOR2_X2 \AES_ENC/U518  ( .A(\AES_ENC/w2[3] ), .B(\AES_ENC/sa31_sub[3] ), .Z(\AES_ENC/N490 ) );
XOR2_X2 \AES_ENC/U517  ( .A(\AES_ENC/w2[2] ), .B(\AES_ENC/sa31_sub[2] ), .Z(\AES_ENC/N491 ) );
XOR2_X2 \AES_ENC/U516  ( .A(\AES_ENC/w2[1] ), .B(\AES_ENC/sa31_sub[1] ), .Z(\AES_ENC/N492 ) );
XOR2_X2 \AES_ENC/U515  ( .A(\AES_ENC/w2[0] ), .B(\AES_ENC/sa31_sub[0] ), .Z(\AES_ENC/N493 ) );
XOR2_X2 \AES_ENC/U514  ( .A(\AES_ENC/w3[7] ), .B(\AES_ENC/sa32_sub[7] ), .Z(\AES_ENC/N494 ) );
XOR2_X2 \AES_ENC/U513  ( .A(\AES_ENC/w3[6] ), .B(\AES_ENC/sa32_sub[6] ), .Z(\AES_ENC/N495 ) );
XOR2_X2 \AES_ENC/U512  ( .A(\AES_ENC/w3[5] ), .B(\AES_ENC/sa32_sub[5] ), .Z(\AES_ENC/N496 ) );
XOR2_X2 \AES_ENC/U511  ( .A(\AES_ENC/w3[4] ), .B(\AES_ENC/sa32_sub[4] ), .Z(\AES_ENC/N497 ) );
XOR2_X2 \AES_ENC/U510  ( .A(\AES_ENC/w3[3] ), .B(\AES_ENC/sa32_sub[3] ), .Z(\AES_ENC/N498 ) );
XOR2_X2 \AES_ENC/U509  ( .A(\AES_ENC/w3[2] ), .B(\AES_ENC/sa32_sub[2] ), .Z(\AES_ENC/N499 ) );
NAND2_X2 \AES_ENC/U508  ( .A1(\AES_ENC/sa23_next [4]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n355 ) );
XOR2_X2 \AES_ENC/U507  ( .A(\AES_ENC/w3[12] ), .B(\AES_ENC/text_in_r[12] ),.Z(\AES_ENC/n357 ) );
NAND2_X2 \AES_ENC/U506  ( .A1(\AES_ENC/n357 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n356 ) );
NAND2_X2 \AES_ENC/U505  ( .A1(\AES_ENC/n355 ), .A2(\AES_ENC/n356 ), .ZN(\AES_ENC/N50 ) );
XOR2_X2 \AES_ENC/U504  ( .A(\AES_ENC/w3[1] ), .B(\AES_ENC/sa32_sub[1] ), .Z(\AES_ENC/N500 ) );
XOR2_X2 \AES_ENC/U503  ( .A(\AES_ENC/w3[0] ), .B(\AES_ENC/sa32_sub[0] ), .Z(\AES_ENC/N501 ) );
NAND2_X2 \AES_ENC/U502  ( .A1(\AES_ENC/sa23_next [5]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n352 ) );
XOR2_X2 \AES_ENC/U501  ( .A(\AES_ENC/w3[13] ), .B(\AES_ENC/text_in_r[13] ),.Z(\AES_ENC/n354 ) );
NAND2_X2 \AES_ENC/U500  ( .A1(\AES_ENC/n354 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n353 ) );
NAND2_X2 \AES_ENC/U499  ( .A1(\AES_ENC/n352 ), .A2(\AES_ENC/n353 ), .ZN(\AES_ENC/N51 ) );
NAND2_X2 \AES_ENC/U498  ( .A1(\AES_ENC/sa23_next [6]), .A2(\AES_ENC/n1255 ),.ZN(\AES_ENC/n349 ) );
XOR2_X2 \AES_ENC/U497  ( .A(\AES_ENC/w3[14] ), .B(\AES_ENC/text_in_r[14] ),.Z(\AES_ENC/n351 ) );
NAND2_X2 \AES_ENC/U496  ( .A1(\AES_ENC/n351 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n3501 ) );
NAND2_X2 \AES_ENC/U495  ( .A1(\AES_ENC/n349 ), .A2(\AES_ENC/n3501 ), .ZN(\AES_ENC/N52 ) );
NAND2_X2 \AES_ENC/U494  ( .A1(\AES_ENC/sa23_next [7]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n346 ) );
XOR2_X2 \AES_ENC/U493  ( .A(\AES_ENC/w3[15] ), .B(\AES_ENC/text_in_r[15] ),.Z(\AES_ENC/n348 ) );
NAND2_X2 \AES_ENC/U492  ( .A1(\AES_ENC/n348 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n347 ) );
NAND2_X2 \AES_ENC/U491  ( .A1(\AES_ENC/n346 ), .A2(\AES_ENC/n347 ), .ZN(\AES_ENC/N53 ) );
NAND2_X2 \AES_ENC/U490  ( .A1(\AES_ENC/sa13_next [0]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n343 ) );
XOR2_X2 \AES_ENC/U489  ( .A(\AES_ENC/w3[16] ), .B(\AES_ENC/text_in_r[16] ),.Z(\AES_ENC/n345 ) );
NAND2_X2 \AES_ENC/U488  ( .A1(\AES_ENC/n345 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n344 ) );
NAND2_X2 \AES_ENC/U487  ( .A1(\AES_ENC/n343 ), .A2(\AES_ENC/n344 ), .ZN(\AES_ENC/N62 ) );
NAND2_X2 \AES_ENC/U486  ( .A1(\AES_ENC/sa13_next [1]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n3401 ) );
XOR2_X2 \AES_ENC/U485  ( .A(\AES_ENC/w3[17] ), .B(\AES_ENC/text_in_r[17] ),.Z(\AES_ENC/n342 ) );
NAND2_X2 \AES_ENC/U484  ( .A1(\AES_ENC/n342 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n341 ) );
NAND2_X2 \AES_ENC/U483  ( .A1(\AES_ENC/n3401 ), .A2(\AES_ENC/n341 ), .ZN(\AES_ENC/N63 ) );
NAND2_X2 \AES_ENC/U482  ( .A1(\AES_ENC/sa13_next [2]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n337 ) );
XOR2_X2 \AES_ENC/U481  ( .A(\AES_ENC/w3[18] ), .B(\AES_ENC/text_in_r[18] ),.Z(\AES_ENC/n339 ) );
NAND2_X2 \AES_ENC/U480  ( .A1(\AES_ENC/n339 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n338 ) );
NAND2_X2 \AES_ENC/U479  ( .A1(\AES_ENC/n337 ), .A2(\AES_ENC/n338 ), .ZN(\AES_ENC/N64 ) );
NAND2_X2 \AES_ENC/U478  ( .A1(\AES_ENC/sa13_next [3]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n334 ) );
XOR2_X2 \AES_ENC/U477  ( .A(\AES_ENC/w3[19] ), .B(\AES_ENC/text_in_r[19] ),.Z(\AES_ENC/n336 ) );
NAND2_X2 \AES_ENC/U476  ( .A1(\AES_ENC/n336 ), .A2(\AES_ENC/n1248 ), .ZN(\AES_ENC/n335 ) );
NAND2_X2 \AES_ENC/U475  ( .A1(\AES_ENC/n334 ), .A2(\AES_ENC/n335 ), .ZN(\AES_ENC/N65 ) );
NAND2_X2 \AES_ENC/U474  ( .A1(\AES_ENC/sa13_next [4]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n331 ) );
XOR2_X2 \AES_ENC/U473  ( .A(\AES_ENC/w3[20] ), .B(\AES_ENC/text_in_r[20] ),.Z(\AES_ENC/n333 ) );
NAND2_X2 \AES_ENC/U472  ( .A1(\AES_ENC/n333 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n332 ) );
NAND2_X2 \AES_ENC/U471  ( .A1(\AES_ENC/n331 ), .A2(\AES_ENC/n332 ), .ZN(\AES_ENC/N66 ) );
NAND2_X2 \AES_ENC/U470  ( .A1(\AES_ENC/sa13_next [5]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n328 ) );
XOR2_X2 \AES_ENC/U469  ( .A(\AES_ENC/w3[21] ), .B(\AES_ENC/text_in_r[21] ),.Z(\AES_ENC/n3301 ) );
NAND2_X2 \AES_ENC/U468  ( .A1(\AES_ENC/n3301 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n329 ) );
NAND2_X2 \AES_ENC/U467  ( .A1(\AES_ENC/n328 ), .A2(\AES_ENC/n329 ), .ZN(\AES_ENC/N67 ) );
NAND2_X2 \AES_ENC/U466  ( .A1(\AES_ENC/sa13_next [6]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n325 ) );
XOR2_X2 \AES_ENC/U465  ( .A(\AES_ENC/w3[22] ), .B(\AES_ENC/text_in_r[22] ),.Z(\AES_ENC/n327 ) );
NAND2_X2 \AES_ENC/U464  ( .A1(\AES_ENC/n327 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n326 ) );
NAND2_X2 \AES_ENC/U463  ( .A1(\AES_ENC/n325 ), .A2(\AES_ENC/n326 ), .ZN(\AES_ENC/N68 ) );
NAND2_X2 \AES_ENC/U462  ( .A1(\AES_ENC/sa13_next [7]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n322 ) );
XOR2_X2 \AES_ENC/U461  ( .A(\AES_ENC/w3[23] ), .B(\AES_ENC/text_in_r[23] ),.Z(\AES_ENC/n324 ) );
NAND2_X2 \AES_ENC/U460  ( .A1(\AES_ENC/n324 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n323 ) );
NAND2_X2 \AES_ENC/U459  ( .A1(\AES_ENC/n322 ), .A2(\AES_ENC/n323 ), .ZN(\AES_ENC/N69 ) );
NAND2_X2 \AES_ENC/U458  ( .A1(\AES_ENC/sa03_next [0]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n319 ) );
XOR2_X2 \AES_ENC/U457  ( .A(\AES_ENC/w3[24] ), .B(\AES_ENC/text_in_r[24] ),.Z(\AES_ENC/n321 ) );
NAND2_X2 \AES_ENC/U456  ( .A1(\AES_ENC/n321 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n3201 ) );
NAND2_X2 \AES_ENC/U455  ( .A1(\AES_ENC/n319 ), .A2(\AES_ENC/n3201 ), .ZN(\AES_ENC/N78 ) );
NAND2_X2 \AES_ENC/U454  ( .A1(\AES_ENC/sa03_next [1]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n316 ) );
XOR2_X2 \AES_ENC/U453  ( .A(\AES_ENC/w3[25] ), .B(\AES_ENC/text_in_r[25] ),.Z(\AES_ENC/n318 ) );
NAND2_X2 \AES_ENC/U452  ( .A1(\AES_ENC/n318 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n317 ) );
NAND2_X2 \AES_ENC/U451  ( .A1(\AES_ENC/n316 ), .A2(\AES_ENC/n317 ), .ZN(\AES_ENC/N79 ) );
NAND2_X2 \AES_ENC/U450  ( .A1(\AES_ENC/sa03_next [2]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n313 ) );
XOR2_X2 \AES_ENC/U449  ( .A(\AES_ENC/w3[26] ), .B(\AES_ENC/text_in_r[26] ),.Z(\AES_ENC/n315 ) );
NAND2_X2 \AES_ENC/U448  ( .A1(\AES_ENC/n315 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n314 ) );
NAND2_X2 \AES_ENC/U447  ( .A1(\AES_ENC/n313 ), .A2(\AES_ENC/n314 ), .ZN(\AES_ENC/N80 ) );
NAND2_X2 \AES_ENC/U446  ( .A1(\AES_ENC/sa03_next [3]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n3101 ) );
XOR2_X2 \AES_ENC/U445  ( .A(\AES_ENC/w3[27] ), .B(\AES_ENC/text_in_r[27] ),.Z(\AES_ENC/n312 ) );
NAND2_X2 \AES_ENC/U444  ( .A1(\AES_ENC/n312 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n311 ) );
NAND2_X2 \AES_ENC/U443  ( .A1(\AES_ENC/n3101 ), .A2(\AES_ENC/n311 ), .ZN(\AES_ENC/N81 ) );
NAND2_X2 \AES_ENC/U442  ( .A1(\AES_ENC/sa03_next [4]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n307 ) );
XOR2_X2 \AES_ENC/U441  ( .A(\AES_ENC/w3[28] ), .B(\AES_ENC/text_in_r[28] ),.Z(\AES_ENC/n309 ) );
NAND2_X2 \AES_ENC/U440  ( .A1(\AES_ENC/n309 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n308 ) );
NAND2_X2 \AES_ENC/U439  ( .A1(\AES_ENC/n307 ), .A2(\AES_ENC/n308 ), .ZN(\AES_ENC/N82 ) );
NAND2_X2 \AES_ENC/U438  ( .A1(\AES_ENC/sa03_next [5]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n304 ) );
XOR2_X2 \AES_ENC/U437  ( .A(\AES_ENC/w3[29] ), .B(\AES_ENC/text_in_r[29] ),.Z(\AES_ENC/n306 ) );
NAND2_X2 \AES_ENC/U436  ( .A1(\AES_ENC/n306 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n305 ) );
NAND2_X2 \AES_ENC/U435  ( .A1(\AES_ENC/n304 ), .A2(\AES_ENC/n305 ), .ZN(\AES_ENC/N83 ) );
NAND2_X2 \AES_ENC/U434  ( .A1(\AES_ENC/sa03_next [6]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n301 ) );
XOR2_X2 \AES_ENC/U433  ( .A(\AES_ENC/w3[30] ), .B(\AES_ENC/text_in_r[30] ),.Z(\AES_ENC/n303 ) );
NAND2_X2 \AES_ENC/U432  ( .A1(\AES_ENC/n303 ), .A2(\AES_ENC/n1249 ), .ZN(\AES_ENC/n302 ) );
NAND2_X2 \AES_ENC/U431  ( .A1(\AES_ENC/n301 ), .A2(\AES_ENC/n302 ), .ZN(\AES_ENC/N84 ) );
NAND2_X2 \AES_ENC/U430  ( .A1(\AES_ENC/sa03_next [7]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n298 ) );
XOR2_X2 \AES_ENC/U429  ( .A(\AES_ENC/w3[31] ), .B(\AES_ENC/text_in_r[31] ),.Z(\AES_ENC/n3001 ) );
NAND2_X2 \AES_ENC/U428  ( .A1(\AES_ENC/n3001 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n299 ) );
NAND2_X2 \AES_ENC/U427  ( .A1(\AES_ENC/n298 ), .A2(\AES_ENC/n299 ), .ZN(\AES_ENC/N85 ) );
NAND2_X2 \AES_ENC/U426  ( .A1(\AES_ENC/sa32_next [0]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n295 ) );
XOR2_X2 \AES_ENC/U425  ( .A(\AES_ENC/w2[0] ), .B(\AES_ENC/text_in_r[32] ),.Z(\AES_ENC/n297 ) );
NAND2_X2 \AES_ENC/U424  ( .A1(\AES_ENC/n297 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n296 ) );
NAND2_X2 \AES_ENC/U423  ( .A1(\AES_ENC/n295 ), .A2(\AES_ENC/n296 ), .ZN(\AES_ENC/N94 ) );
NAND2_X2 \AES_ENC/U422  ( .A1(\AES_ENC/sa32_next [1]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n292 ) );
XOR2_X2 \AES_ENC/U421  ( .A(\AES_ENC/w2[1] ), .B(\AES_ENC/text_in_r[33] ),.Z(\AES_ENC/n294 ) );
NAND2_X2 \AES_ENC/U420  ( .A1(\AES_ENC/n294 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n293 ) );
NAND2_X2 \AES_ENC/U419  ( .A1(\AES_ENC/n292 ), .A2(\AES_ENC/n293 ), .ZN(\AES_ENC/N95 ) );
NAND2_X2 \AES_ENC/U418  ( .A1(\AES_ENC/sa32_next [2]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n289 ) );
XOR2_X2 \AES_ENC/U417  ( .A(\AES_ENC/w2[2] ), .B(\AES_ENC/text_in_r[34] ),.Z(\AES_ENC/n291 ) );
NAND2_X2 \AES_ENC/U416  ( .A1(\AES_ENC/n291 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n290 ) );
NAND2_X2 \AES_ENC/U415  ( .A1(\AES_ENC/n289 ), .A2(\AES_ENC/n290 ), .ZN(\AES_ENC/N96 ) );
NAND2_X2 \AES_ENC/U414  ( .A1(\AES_ENC/sa32_next [3]), .A2(\AES_ENC/n1256 ),.ZN(\AES_ENC/n286 ) );
XOR2_X2 \AES_ENC/U413  ( .A(\AES_ENC/w2[3] ), .B(\AES_ENC/text_in_r[35] ),.Z(\AES_ENC/n288 ) );
NAND2_X2 \AES_ENC/U412  ( .A1(\AES_ENC/n288 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n287 ) );
NAND2_X2 \AES_ENC/U411  ( .A1(\AES_ENC/n286 ), .A2(\AES_ENC/n287 ), .ZN(\AES_ENC/N97 ) );
NAND2_X2 \AES_ENC/U410  ( .A1(\AES_ENC/sa32_next [4]), .A2(\AES_ENC/n1252 ),.ZN(\AES_ENC/n283 ) );
XOR2_X2 \AES_ENC/U409  ( .A(\AES_ENC/w2[4] ), .B(\AES_ENC/text_in_r[36] ),.Z(\AES_ENC/n285 ) );
NAND2_X2 \AES_ENC/U408  ( .A1(\AES_ENC/n285 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n284 ) );
NAND2_X2 \AES_ENC/U407  ( .A1(\AES_ENC/n283 ), .A2(\AES_ENC/n284 ), .ZN(\AES_ENC/N98 ) );
NAND2_X2 \AES_ENC/U406  ( .A1(\AES_ENC/sa32_next [5]), .A2(\AES_ENC/n1251 ),.ZN(\AES_ENC/n280 ) );
XOR2_X2 \AES_ENC/U405  ( .A(\AES_ENC/w2[5] ), .B(\AES_ENC/text_in_r[37] ),.Z(\AES_ENC/n282 ) );
NAND2_X2 \AES_ENC/U404  ( .A1(\AES_ENC/n282 ), .A2(\AES_ENC/n1250 ), .ZN(\AES_ENC/n281 ) );
NAND2_X2 \AES_ENC/U403  ( .A1(\AES_ENC/n280 ), .A2(\AES_ENC/n281 ), .ZN(\AES_ENC/N99 ) );
NAND2_X2 \AES_ENC/U402  ( .A1(aes_text_in[0]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n278 ) );
NAND2_X2 \AES_ENC/U401  ( .A1(\AES_ENC/text_in_r[0] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n279 ) );
NAND2_X2 \AES_ENC/U400  ( .A1(\AES_ENC/n278 ), .A2(\AES_ENC/n279 ), .ZN(\AES_ENC/n661 ) );
NAND2_X2 \AES_ENC/U399  ( .A1(aes_text_in[1]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2760 ) );
NAND2_X2 \AES_ENC/U398  ( .A1(\AES_ENC/text_in_r[1] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2770 ) );
NAND2_X2 \AES_ENC/U397  ( .A1(\AES_ENC/n2760 ), .A2(\AES_ENC/n2770 ), .ZN(\AES_ENC/n662 ) );
NAND2_X2 \AES_ENC/U396  ( .A1(aes_text_in[2]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2740 ) );
NAND2_X2 \AES_ENC/U395  ( .A1(\AES_ENC/text_in_r[2] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2750 ) );
NAND2_X2 \AES_ENC/U394  ( .A1(\AES_ENC/n2740 ), .A2(\AES_ENC/n2750 ), .ZN(\AES_ENC/n663 ) );
NAND2_X2 \AES_ENC/U393  ( .A1(aes_text_in[3]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2720 ) );
NAND2_X2 \AES_ENC/U392  ( .A1(\AES_ENC/text_in_r[3] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2730 ) );
NAND2_X2 \AES_ENC/U391  ( .A1(\AES_ENC/n2720 ), .A2(\AES_ENC/n2730 ), .ZN(\AES_ENC/n664 ) );
NAND2_X2 \AES_ENC/U390  ( .A1(aes_text_in[4]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2700 ) );
NAND2_X2 \AES_ENC/U389  ( .A1(\AES_ENC/text_in_r[4] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2710 ) );
NAND2_X2 \AES_ENC/U388  ( .A1(\AES_ENC/n2700 ), .A2(\AES_ENC/n2710 ), .ZN(\AES_ENC/n665 ) );
NAND2_X2 \AES_ENC/U387  ( .A1(aes_text_in[5]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n268 ) );
NAND2_X2 \AES_ENC/U386  ( .A1(\AES_ENC/text_in_r[5] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n269 ) );
NAND2_X2 \AES_ENC/U385  ( .A1(\AES_ENC/n268 ), .A2(\AES_ENC/n269 ), .ZN(\AES_ENC/n666 ) );
NAND2_X2 \AES_ENC/U384  ( .A1(aes_text_in[6]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n266 ) );
NAND2_X2 \AES_ENC/U383  ( .A1(\AES_ENC/text_in_r[6] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n267 ) );
NAND2_X2 \AES_ENC/U382  ( .A1(\AES_ENC/n266 ), .A2(\AES_ENC/n267 ), .ZN(\AES_ENC/n667 ) );
NAND2_X2 \AES_ENC/U381  ( .A1(aes_text_in[7]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n264 ) );
NAND2_X2 \AES_ENC/U380  ( .A1(\AES_ENC/text_in_r[7] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n265 ) );
NAND2_X2 \AES_ENC/U379  ( .A1(\AES_ENC/n264 ), .A2(\AES_ENC/n265 ), .ZN(\AES_ENC/n668 ) );
NAND2_X2 \AES_ENC/U378  ( .A1(aes_text_in[8]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n262 ) );
NAND2_X2 \AES_ENC/U377  ( .A1(\AES_ENC/text_in_r[8] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n263 ) );
NAND2_X2 \AES_ENC/U376  ( .A1(\AES_ENC/n262 ), .A2(\AES_ENC/n263 ), .ZN(\AES_ENC/n669 ) );
NAND2_X2 \AES_ENC/U375  ( .A1(aes_text_in[9]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2600 ) );
NAND2_X2 \AES_ENC/U374  ( .A1(\AES_ENC/text_in_r[9] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2610 ) );
NAND2_X2 \AES_ENC/U373  ( .A1(\AES_ENC/n2600 ), .A2(\AES_ENC/n2610 ), .ZN(\AES_ENC/n670 ) );
NAND2_X2 \AES_ENC/U372  ( .A1(aes_text_in[10]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2580 ) );
NAND2_X2 \AES_ENC/U371  ( .A1(\AES_ENC/text_in_r[10] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2590 ) );
NAND2_X2 \AES_ENC/U370  ( .A1(\AES_ENC/n2580 ), .A2(\AES_ENC/n2590 ), .ZN(\AES_ENC/n671 ) );
NAND2_X2 \AES_ENC/U369  ( .A1(aes_text_in[11]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2560 ) );
NAND2_X2 \AES_ENC/U368  ( .A1(\AES_ENC/text_in_r[11] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2570 ) );
NAND2_X2 \AES_ENC/U367  ( .A1(\AES_ENC/n2560 ), .A2(\AES_ENC/n2570 ), .ZN(\AES_ENC/n672 ) );
NAND2_X2 \AES_ENC/U366  ( .A1(aes_text_in[12]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2540 ) );
NAND2_X2 \AES_ENC/U365  ( .A1(\AES_ENC/text_in_r[12] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2550 ) );
NAND2_X2 \AES_ENC/U364  ( .A1(\AES_ENC/n2540 ), .A2(\AES_ENC/n2550 ), .ZN(\AES_ENC/n673 ) );
NAND2_X2 \AES_ENC/U363  ( .A1(aes_text_in[13]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n252 ) );
NAND2_X2 \AES_ENC/U362  ( .A1(\AES_ENC/text_in_r[13] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n253 ) );
NAND2_X2 \AES_ENC/U361  ( .A1(\AES_ENC/n252 ), .A2(\AES_ENC/n253 ), .ZN(\AES_ENC/n674 ) );
NAND2_X2 \AES_ENC/U360  ( .A1(aes_text_in[14]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n250 ) );
NAND2_X2 \AES_ENC/U359  ( .A1(\AES_ENC/text_in_r[14] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n251 ) );
NAND2_X2 \AES_ENC/U358  ( .A1(\AES_ENC/n250 ), .A2(\AES_ENC/n251 ), .ZN(\AES_ENC/n675 ) );
NAND2_X2 \AES_ENC/U357  ( .A1(aes_text_in[15]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n248 ) );
NAND2_X2 \AES_ENC/U356  ( .A1(\AES_ENC/text_in_r[15] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n249 ) );
NAND2_X2 \AES_ENC/U355  ( .A1(\AES_ENC/n248 ), .A2(\AES_ENC/n249 ), .ZN(\AES_ENC/n676 ) );
NAND2_X2 \AES_ENC/U354  ( .A1(aes_text_in[16]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n246 ) );
NAND2_X2 \AES_ENC/U353  ( .A1(\AES_ENC/text_in_r[16] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n247 ) );
NAND2_X2 \AES_ENC/U352  ( .A1(\AES_ENC/n246 ), .A2(\AES_ENC/n247 ), .ZN(\AES_ENC/n677 ) );
NAND2_X2 \AES_ENC/U351  ( .A1(aes_text_in[17]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2440 ) );
NAND2_X2 \AES_ENC/U350  ( .A1(\AES_ENC/text_in_r[17] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2450 ) );
NAND2_X2 \AES_ENC/U349  ( .A1(\AES_ENC/n2440 ), .A2(\AES_ENC/n2450 ), .ZN(\AES_ENC/n678 ) );
NAND2_X2 \AES_ENC/U348  ( .A1(aes_text_in[18]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2420 ) );
NAND2_X2 \AES_ENC/U347  ( .A1(\AES_ENC/text_in_r[18] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2430 ) );
NAND2_X2 \AES_ENC/U346  ( .A1(\AES_ENC/n2420 ), .A2(\AES_ENC/n2430 ), .ZN(\AES_ENC/n679 ) );
NAND2_X2 \AES_ENC/U345  ( .A1(aes_text_in[19]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2400 ) );
NAND2_X2 \AES_ENC/U344  ( .A1(\AES_ENC/text_in_r[19] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2410 ) );
NAND2_X2 \AES_ENC/U343  ( .A1(\AES_ENC/n2400 ), .A2(\AES_ENC/n2410 ), .ZN(\AES_ENC/n680 ) );
NAND2_X2 \AES_ENC/U342  ( .A1(aes_text_in[20]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2380 ) );
NAND2_X2 \AES_ENC/U341  ( .A1(\AES_ENC/text_in_r[20] ), .A2(\AES_ENC/n1264 ),.ZN(\AES_ENC/n2390 ) );
NAND2_X2 \AES_ENC/U340  ( .A1(\AES_ENC/n2380 ), .A2(\AES_ENC/n2390 ), .ZN(\AES_ENC/n681 ) );
NAND2_X2 \AES_ENC/U339  ( .A1(aes_text_in[21]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n236 ) );
NAND2_X2 \AES_ENC/U338  ( .A1(\AES_ENC/text_in_r[21] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n237 ) );
NAND2_X2 \AES_ENC/U337  ( .A1(\AES_ENC/n236 ), .A2(\AES_ENC/n237 ), .ZN(\AES_ENC/n682 ) );
NAND2_X2 \AES_ENC/U336  ( .A1(aes_text_in[22]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n234 ) );
NAND2_X2 \AES_ENC/U335  ( .A1(\AES_ENC/text_in_r[22] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n235 ) );
NAND2_X2 \AES_ENC/U334  ( .A1(\AES_ENC/n234 ), .A2(\AES_ENC/n235 ), .ZN(\AES_ENC/n683 ) );
NAND2_X2 \AES_ENC/U333  ( .A1(aes_text_in[23]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n232 ) );
NAND2_X2 \AES_ENC/U332  ( .A1(\AES_ENC/text_in_r[23] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n233 ) );
NAND2_X2 \AES_ENC/U331  ( .A1(\AES_ENC/n232 ), .A2(\AES_ENC/n233 ), .ZN(\AES_ENC/n684 ) );
NAND2_X2 \AES_ENC/U330  ( .A1(aes_text_in[24]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n230 ) );
NAND2_X2 \AES_ENC/U329  ( .A1(\AES_ENC/text_in_r[24] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n231 ) );
NAND2_X2 \AES_ENC/U328  ( .A1(\AES_ENC/n230 ), .A2(\AES_ENC/n231 ), .ZN(\AES_ENC/n685 ) );
NAND2_X2 \AES_ENC/U327  ( .A1(aes_text_in[25]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2280 ) );
NAND2_X2 \AES_ENC/U326  ( .A1(\AES_ENC/text_in_r[25] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2290 ) );
NAND2_X2 \AES_ENC/U325  ( .A1(\AES_ENC/n2280 ), .A2(\AES_ENC/n2290 ), .ZN(\AES_ENC/n686 ) );
NAND2_X2 \AES_ENC/U324  ( .A1(aes_text_in[26]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2260 ) );
NAND2_X2 \AES_ENC/U323  ( .A1(\AES_ENC/text_in_r[26] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2270 ) );
NAND2_X2 \AES_ENC/U322  ( .A1(\AES_ENC/n2260 ), .A2(\AES_ENC/n2270 ), .ZN(\AES_ENC/n687 ) );
NAND2_X2 \AES_ENC/U321  ( .A1(aes_text_in[27]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2240 ) );
NAND2_X2 \AES_ENC/U320  ( .A1(\AES_ENC/text_in_r[27] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2250 ) );
NAND2_X2 \AES_ENC/U319  ( .A1(\AES_ENC/n2240 ), .A2(\AES_ENC/n2250 ), .ZN(\AES_ENC/n688 ) );
NAND2_X2 \AES_ENC/U318  ( .A1(aes_text_in[28]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2220 ) );
NAND2_X2 \AES_ENC/U317  ( .A1(\AES_ENC/text_in_r[28] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2230 ) );
NAND2_X2 \AES_ENC/U316  ( .A1(\AES_ENC/n2220 ), .A2(\AES_ENC/n2230 ), .ZN(\AES_ENC/n689 ) );
NAND2_X2 \AES_ENC/U315  ( .A1(aes_text_in[29]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n220 ) );
NAND2_X2 \AES_ENC/U314  ( .A1(\AES_ENC/text_in_r[29] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n221 ) );
NAND2_X2 \AES_ENC/U313  ( .A1(\AES_ENC/n220 ), .A2(\AES_ENC/n221 ), .ZN(\AES_ENC/n690 ) );
NAND2_X2 \AES_ENC/U312  ( .A1(aes_text_in[30]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n218 ) );
NAND2_X2 \AES_ENC/U311  ( .A1(\AES_ENC/text_in_r[30] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n219 ) );
NAND2_X2 \AES_ENC/U310  ( .A1(\AES_ENC/n218 ), .A2(\AES_ENC/n219 ), .ZN(\AES_ENC/n691 ) );
NAND2_X2 \AES_ENC/U309  ( .A1(aes_text_in[31]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n216 ) );
NAND2_X2 \AES_ENC/U308  ( .A1(\AES_ENC/text_in_r[31] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n217 ) );
NAND2_X2 \AES_ENC/U307  ( .A1(\AES_ENC/n216 ), .A2(\AES_ENC/n217 ), .ZN(\AES_ENC/n692 ) );
NAND2_X2 \AES_ENC/U306  ( .A1(aes_text_in[32]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n214 ) );
NAND2_X2 \AES_ENC/U305  ( .A1(\AES_ENC/text_in_r[32] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n215 ) );
NAND2_X2 \AES_ENC/U304  ( .A1(\AES_ENC/n214 ), .A2(\AES_ENC/n215 ), .ZN(\AES_ENC/n693 ) );
NAND2_X2 \AES_ENC/U303  ( .A1(aes_text_in[33]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2120 ) );
NAND2_X2 \AES_ENC/U302  ( .A1(\AES_ENC/text_in_r[33] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2130 ) );
NAND2_X2 \AES_ENC/U301  ( .A1(\AES_ENC/n2120 ), .A2(\AES_ENC/n2130 ), .ZN(\AES_ENC/n694 ) );
NAND2_X2 \AES_ENC/U300  ( .A1(aes_text_in[34]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2100 ) );
NAND2_X2 \AES_ENC/U299  ( .A1(\AES_ENC/text_in_r[34] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2110 ) );
NAND2_X2 \AES_ENC/U298  ( .A1(\AES_ENC/n2100 ), .A2(\AES_ENC/n2110 ), .ZN(\AES_ENC/n695 ) );
NAND2_X2 \AES_ENC/U297  ( .A1(aes_text_in[35]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2080 ) );
NAND2_X2 \AES_ENC/U296  ( .A1(\AES_ENC/text_in_r[35] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2090 ) );
NAND2_X2 \AES_ENC/U295  ( .A1(\AES_ENC/n2080 ), .A2(\AES_ENC/n2090 ), .ZN(\AES_ENC/n696 ) );
NAND2_X2 \AES_ENC/U294  ( .A1(aes_text_in[36]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n2060 ) );
NAND2_X2 \AES_ENC/U293  ( .A1(\AES_ENC/text_in_r[36] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n2070 ) );
NAND2_X2 \AES_ENC/U292  ( .A1(\AES_ENC/n2060 ), .A2(\AES_ENC/n2070 ), .ZN(\AES_ENC/n697 ) );
NAND2_X2 \AES_ENC/U291  ( .A1(aes_text_in[37]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n204 ) );
NAND2_X2 \AES_ENC/U290  ( .A1(\AES_ENC/text_in_r[37] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n205 ) );
NAND2_X2 \AES_ENC/U289  ( .A1(\AES_ENC/n204 ), .A2(\AES_ENC/n205 ), .ZN(\AES_ENC/n698 ) );
NAND2_X2 \AES_ENC/U288  ( .A1(aes_text_in[38]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n202 ) );
NAND2_X2 \AES_ENC/U287  ( .A1(\AES_ENC/text_in_r[38] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n203 ) );
NAND2_X2 \AES_ENC/U286  ( .A1(\AES_ENC/n202 ), .A2(\AES_ENC/n203 ), .ZN(\AES_ENC/n699 ) );
NAND2_X2 \AES_ENC/U285  ( .A1(aes_text_in[39]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n200 ) );
NAND2_X2 \AES_ENC/U284  ( .A1(\AES_ENC/text_in_r[39] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n201 ) );
NAND2_X2 \AES_ENC/U283  ( .A1(\AES_ENC/n200 ), .A2(\AES_ENC/n201 ), .ZN(\AES_ENC/n700 ) );
NAND2_X2 \AES_ENC/U282  ( .A1(aes_text_in[40]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1981 ) );
NAND2_X2 \AES_ENC/U281  ( .A1(\AES_ENC/text_in_r[40] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n199 ) );
NAND2_X2 \AES_ENC/U280  ( .A1(\AES_ENC/n1981 ), .A2(\AES_ENC/n199 ), .ZN(\AES_ENC/n701 ) );
NAND2_X2 \AES_ENC/U279  ( .A1(aes_text_in[41]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1960 ) );
NAND2_X2 \AES_ENC/U278  ( .A1(\AES_ENC/text_in_r[41] ), .A2(\AES_ENC/n1263 ),.ZN(\AES_ENC/n1970 ) );
NAND2_X2 \AES_ENC/U277  ( .A1(\AES_ENC/n1960 ), .A2(\AES_ENC/n1970 ), .ZN(\AES_ENC/n702 ) );
NAND2_X2 \AES_ENC/U276  ( .A1(aes_text_in[42]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1940 ) );
NAND2_X2 \AES_ENC/U275  ( .A1(\AES_ENC/text_in_r[42] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1950 ) );
NAND2_X2 \AES_ENC/U274  ( .A1(\AES_ENC/n1940 ), .A2(\AES_ENC/n1950 ), .ZN(\AES_ENC/n703 ) );
NAND2_X2 \AES_ENC/U273  ( .A1(aes_text_in[43]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1920 ) );
NAND2_X2 \AES_ENC/U272  ( .A1(\AES_ENC/text_in_r[43] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1930 ) );
NAND2_X2 \AES_ENC/U271  ( .A1(\AES_ENC/n1920 ), .A2(\AES_ENC/n1930 ), .ZN(\AES_ENC/n704 ) );
NAND2_X2 \AES_ENC/U270  ( .A1(aes_text_in[44]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1900 ) );
NAND2_X2 \AES_ENC/U269  ( .A1(\AES_ENC/text_in_r[44] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1910 ) );
NAND2_X2 \AES_ENC/U268  ( .A1(\AES_ENC/n1900 ), .A2(\AES_ENC/n1910 ), .ZN(\AES_ENC/n705 ) );
NAND2_X2 \AES_ENC/U267  ( .A1(aes_text_in[45]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n188 ) );
NAND2_X2 \AES_ENC/U266  ( .A1(\AES_ENC/text_in_r[45] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n189 ) );
NAND2_X2 \AES_ENC/U265  ( .A1(\AES_ENC/n188 ), .A2(\AES_ENC/n189 ), .ZN(\AES_ENC/n706 ) );
NAND2_X2 \AES_ENC/U264  ( .A1(aes_text_in[46]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n186 ) );
NAND2_X2 \AES_ENC/U263  ( .A1(\AES_ENC/text_in_r[46] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n187 ) );
NAND2_X2 \AES_ENC/U262  ( .A1(\AES_ENC/n186 ), .A2(\AES_ENC/n187 ), .ZN(\AES_ENC/n707 ) );
NAND2_X2 \AES_ENC/U261  ( .A1(aes_text_in[47]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n184 ) );
NAND2_X2 \AES_ENC/U260  ( .A1(\AES_ENC/text_in_r[47] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n185 ) );
NAND2_X2 \AES_ENC/U259  ( .A1(\AES_ENC/n184 ), .A2(\AES_ENC/n185 ), .ZN(\AES_ENC/n708 ) );
NAND2_X2 \AES_ENC/U258  ( .A1(aes_text_in[48]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n182 ) );
NAND2_X2 \AES_ENC/U257  ( .A1(\AES_ENC/text_in_r[48] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n183 ) );
NAND2_X2 \AES_ENC/U256  ( .A1(\AES_ENC/n182 ), .A2(\AES_ENC/n183 ), .ZN(\AES_ENC/n709 ) );
NAND2_X2 \AES_ENC/U255  ( .A1(aes_text_in[49]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1800 ) );
NAND2_X2 \AES_ENC/U254  ( .A1(\AES_ENC/text_in_r[49] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1810 ) );
NAND2_X2 \AES_ENC/U253  ( .A1(\AES_ENC/n1800 ), .A2(\AES_ENC/n1810 ), .ZN(\AES_ENC/n710 ) );
NAND2_X2 \AES_ENC/U252  ( .A1(aes_text_in[50]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1780 ) );
NAND2_X2 \AES_ENC/U251  ( .A1(\AES_ENC/text_in_r[50] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1790 ) );
NAND2_X2 \AES_ENC/U250  ( .A1(\AES_ENC/n1780 ), .A2(\AES_ENC/n1790 ), .ZN(\AES_ENC/n711 ) );
NAND2_X2 \AES_ENC/U249  ( .A1(aes_text_in[51]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1760 ) );
NAND2_X2 \AES_ENC/U248  ( .A1(\AES_ENC/text_in_r[51] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1770 ) );
NAND2_X2 \AES_ENC/U247  ( .A1(\AES_ENC/n1760 ), .A2(\AES_ENC/n1770 ), .ZN(\AES_ENC/n712 ) );
NAND2_X2 \AES_ENC/U246  ( .A1(aes_text_in[52]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n1740 ) );
NAND2_X2 \AES_ENC/U245  ( .A1(\AES_ENC/text_in_r[52] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1750 ) );
NAND2_X2 \AES_ENC/U244  ( .A1(\AES_ENC/n1740 ), .A2(\AES_ENC/n1750 ), .ZN(\AES_ENC/n713 ) );
NAND2_X2 \AES_ENC/U243  ( .A1(aes_text_in[53]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n172 ) );
NAND2_X2 \AES_ENC/U242  ( .A1(\AES_ENC/text_in_r[53] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n173 ) );
NAND2_X2 \AES_ENC/U241  ( .A1(\AES_ENC/n172 ), .A2(\AES_ENC/n173 ), .ZN(\AES_ENC/n714 ) );
NAND2_X2 \AES_ENC/U240  ( .A1(aes_text_in[54]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n170 ) );
NAND2_X2 \AES_ENC/U239  ( .A1(\AES_ENC/text_in_r[54] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n171 ) );
NAND2_X2 \AES_ENC/U238  ( .A1(\AES_ENC/n170 ), .A2(\AES_ENC/n171 ), .ZN(\AES_ENC/n715 ) );
NAND2_X2 \AES_ENC/U237  ( .A1(aes_text_in[55]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n168 ) );
NAND2_X2 \AES_ENC/U236  ( .A1(\AES_ENC/text_in_r[55] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n169 ) );
NAND2_X2 \AES_ENC/U235  ( .A1(\AES_ENC/n168 ), .A2(\AES_ENC/n169 ), .ZN(\AES_ENC/n716 ) );
NAND2_X2 \AES_ENC/U234  ( .A1(aes_text_in[56]), .A2(\AES_ENC/n1257 ), .ZN(\AES_ENC/n166 ) );
NAND2_X2 \AES_ENC/U233  ( .A1(\AES_ENC/text_in_r[56] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n167 ) );
NAND2_X2 \AES_ENC/U232  ( .A1(\AES_ENC/n166 ), .A2(\AES_ENC/n167 ), .ZN(\AES_ENC/n717 ) );
NAND2_X2 \AES_ENC/U231  ( .A1(aes_text_in[57]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n1640 ) );
NAND2_X2 \AES_ENC/U230  ( .A1(\AES_ENC/text_in_r[57] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1650 ) );
NAND2_X2 \AES_ENC/U229  ( .A1(\AES_ENC/n1640 ), .A2(\AES_ENC/n1650 ), .ZN(\AES_ENC/n718 ) );
NAND2_X2 \AES_ENC/U228  ( .A1(aes_text_in[58]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n1620 ) );
NAND2_X2 \AES_ENC/U227  ( .A1(\AES_ENC/text_in_r[58] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1630 ) );
NAND2_X2 \AES_ENC/U226  ( .A1(\AES_ENC/n1620 ), .A2(\AES_ENC/n1630 ), .ZN(\AES_ENC/n719 ) );
NAND2_X2 \AES_ENC/U225  ( .A1(aes_text_in[59]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n1600 ) );
NAND2_X2 \AES_ENC/U224  ( .A1(\AES_ENC/text_in_r[59] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1610 ) );
NAND2_X2 \AES_ENC/U223  ( .A1(\AES_ENC/n1600 ), .A2(\AES_ENC/n1610 ), .ZN(\AES_ENC/n720 ) );
NAND2_X2 \AES_ENC/U222  ( .A1(aes_text_in[60]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n1580 ) );
NAND2_X2 \AES_ENC/U221  ( .A1(\AES_ENC/text_in_r[60] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n1590 ) );
NAND2_X2 \AES_ENC/U220  ( .A1(\AES_ENC/n1580 ), .A2(\AES_ENC/n1590 ), .ZN(\AES_ENC/n721 ) );
NAND2_X2 \AES_ENC/U219  ( .A1(aes_text_in[61]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n156 ) );
NAND2_X2 \AES_ENC/U218  ( .A1(\AES_ENC/text_in_r[61] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n157 ) );
NAND2_X2 \AES_ENC/U217  ( .A1(\AES_ENC/n156 ), .A2(\AES_ENC/n157 ), .ZN(\AES_ENC/n722 ) );
NAND2_X2 \AES_ENC/U216  ( .A1(aes_text_in[62]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n154 ) );
NAND2_X2 \AES_ENC/U215  ( .A1(\AES_ENC/text_in_r[62] ), .A2(\AES_ENC/n1262 ),.ZN(\AES_ENC/n155 ) );
NAND2_X2 \AES_ENC/U214  ( .A1(\AES_ENC/n154 ), .A2(\AES_ENC/n155 ), .ZN(\AES_ENC/n723 ) );
NAND2_X2 \AES_ENC/U213  ( .A1(aes_text_in[63]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n152 ) );
NAND2_X2 \AES_ENC/U212  ( .A1(\AES_ENC/text_in_r[63] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n153 ) );
NAND2_X2 \AES_ENC/U211  ( .A1(\AES_ENC/n152 ), .A2(\AES_ENC/n153 ), .ZN(\AES_ENC/n724 ) );
NAND2_X2 \AES_ENC/U210  ( .A1(aes_text_in[64]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n150 ) );
NAND2_X2 \AES_ENC/U209  ( .A1(\AES_ENC/text_in_r[64] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n151 ) );
NAND2_X2 \AES_ENC/U208  ( .A1(\AES_ENC/n150 ), .A2(\AES_ENC/n151 ), .ZN(\AES_ENC/n725 ) );
NAND2_X2 \AES_ENC/U207  ( .A1(aes_text_in[65]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n1480 ) );
NAND2_X2 \AES_ENC/U206  ( .A1(\AES_ENC/text_in_r[65] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1490 ) );
NAND2_X2 \AES_ENC/U205  ( .A1(\AES_ENC/n1480 ), .A2(\AES_ENC/n1490 ), .ZN(\AES_ENC/n726 ) );
NAND2_X2 \AES_ENC/U204  ( .A1(aes_text_in[66]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n1460 ) );
NAND2_X2 \AES_ENC/U203  ( .A1(\AES_ENC/text_in_r[66] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1470 ) );
NAND2_X2 \AES_ENC/U202  ( .A1(\AES_ENC/n1460 ), .A2(\AES_ENC/n1470 ), .ZN(\AES_ENC/n727 ) );
NAND2_X2 \AES_ENC/U201  ( .A1(aes_text_in[67]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n1440 ) );
NAND2_X2 \AES_ENC/U200  ( .A1(\AES_ENC/text_in_r[67] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1450 ) );
NAND2_X2 \AES_ENC/U199  ( .A1(\AES_ENC/n1440 ), .A2(\AES_ENC/n1450 ), .ZN(\AES_ENC/n728 ) );
NAND2_X2 \AES_ENC/U198  ( .A1(aes_text_in[68]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n1420 ) );
NAND2_X2 \AES_ENC/U197  ( .A1(\AES_ENC/text_in_r[68] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1430 ) );
NAND2_X2 \AES_ENC/U196  ( .A1(\AES_ENC/n1420 ), .A2(\AES_ENC/n1430 ), .ZN(\AES_ENC/n729 ) );
NAND2_X2 \AES_ENC/U195  ( .A1(aes_text_in[69]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n140 ) );
NAND2_X2 \AES_ENC/U194  ( .A1(\AES_ENC/text_in_r[69] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n141 ) );
NAND2_X2 \AES_ENC/U193  ( .A1(\AES_ENC/n140 ), .A2(\AES_ENC/n141 ), .ZN(\AES_ENC/n730 ) );
NAND2_X2 \AES_ENC/U192  ( .A1(aes_text_in[70]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n138 ) );
NAND2_X2 \AES_ENC/U191  ( .A1(\AES_ENC/text_in_r[70] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n139 ) );
NAND2_X2 \AES_ENC/U190  ( .A1(\AES_ENC/n138 ), .A2(\AES_ENC/n139 ), .ZN(\AES_ENC/n731 ) );
NAND2_X2 \AES_ENC/U189  ( .A1(aes_text_in[71]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n136 ) );
NAND2_X2 \AES_ENC/U188  ( .A1(\AES_ENC/text_in_r[71] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n137 ) );
NAND2_X2 \AES_ENC/U187  ( .A1(\AES_ENC/n136 ), .A2(\AES_ENC/n137 ), .ZN(\AES_ENC/n732 ) );
NAND2_X2 \AES_ENC/U186  ( .A1(aes_text_in[72]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n134 ) );
NAND2_X2 \AES_ENC/U185  ( .A1(\AES_ENC/text_in_r[72] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n135 ) );
NAND2_X2 \AES_ENC/U184  ( .A1(\AES_ENC/n134 ), .A2(\AES_ENC/n135 ), .ZN(\AES_ENC/n733 ) );
NAND2_X2 \AES_ENC/U183  ( .A1(aes_text_in[73]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n1320 ) );
NAND2_X2 \AES_ENC/U182  ( .A1(\AES_ENC/text_in_r[73] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1330 ) );
NAND2_X2 \AES_ENC/U181  ( .A1(\AES_ENC/n1320 ), .A2(\AES_ENC/n1330 ), .ZN(\AES_ENC/n734 ) );
NAND2_X2 \AES_ENC/U180  ( .A1(aes_text_in[74]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n1300 ) );
NAND2_X2 \AES_ENC/U179  ( .A1(\AES_ENC/text_in_r[74] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1310 ) );
NAND2_X2 \AES_ENC/U178  ( .A1(\AES_ENC/n1300 ), .A2(\AES_ENC/n1310 ), .ZN(\AES_ENC/n735 ) );
NAND2_X2 \AES_ENC/U177  ( .A1(aes_text_in[75]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n1280 ) );
NAND2_X2 \AES_ENC/U176  ( .A1(\AES_ENC/text_in_r[75] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1290 ) );
NAND2_X2 \AES_ENC/U175  ( .A1(\AES_ENC/n1280 ), .A2(\AES_ENC/n1290 ), .ZN(\AES_ENC/n736 ) );
NAND2_X2 \AES_ENC/U174  ( .A1(aes_text_in[76]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n12600 ) );
NAND2_X2 \AES_ENC/U173  ( .A1(\AES_ENC/text_in_r[76] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n1270 ) );
NAND2_X2 \AES_ENC/U172  ( .A1(\AES_ENC/n12600 ), .A2(\AES_ENC/n1270 ), .ZN(\AES_ENC/n737 ) );
NAND2_X2 \AES_ENC/U171  ( .A1(aes_text_in[77]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n124 ) );
NAND2_X2 \AES_ENC/U170  ( .A1(\AES_ENC/text_in_r[77] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n125 ) );
NAND2_X2 \AES_ENC/U169  ( .A1(\AES_ENC/n124 ), .A2(\AES_ENC/n125 ), .ZN(\AES_ENC/n738 ) );
NAND2_X2 \AES_ENC/U168  ( .A1(aes_text_in[78]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n122 ) );
NAND2_X2 \AES_ENC/U167  ( .A1(\AES_ENC/text_in_r[78] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n123 ) );
NAND2_X2 \AES_ENC/U166  ( .A1(\AES_ENC/n122 ), .A2(\AES_ENC/n123 ), .ZN(\AES_ENC/n739 ) );
NAND2_X2 \AES_ENC/U165  ( .A1(aes_text_in[79]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n120 ) );
NAND2_X2 \AES_ENC/U164  ( .A1(\AES_ENC/text_in_r[79] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n121 ) );
NAND2_X2 \AES_ENC/U163  ( .A1(\AES_ENC/n120 ), .A2(\AES_ENC/n121 ), .ZN(\AES_ENC/n740 ) );
NAND2_X2 \AES_ENC/U162  ( .A1(aes_text_in[80]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n118 ) );
NAND2_X2 \AES_ENC/U161  ( .A1(\AES_ENC/text_in_r[80] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n119 ) );
NAND2_X2 \AES_ENC/U160  ( .A1(\AES_ENC/n118 ), .A2(\AES_ENC/n119 ), .ZN(\AES_ENC/n741 ) );
NAND2_X2 \AES_ENC/U159  ( .A1(aes_text_in[81]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n11610 ) );
NAND2_X2 \AES_ENC/U158  ( .A1(\AES_ENC/text_in_r[81] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n11710 ) );
NAND2_X2 \AES_ENC/U157  ( .A1(\AES_ENC/n11610 ), .A2(\AES_ENC/n11710 ), .ZN(\AES_ENC/n742 ) );
NAND2_X2 \AES_ENC/U156  ( .A1(aes_text_in[82]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n11410 ) );
NAND2_X2 \AES_ENC/U155  ( .A1(\AES_ENC/text_in_r[82] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n11510 ) );
NAND2_X2 \AES_ENC/U154  ( .A1(\AES_ENC/n11410 ), .A2(\AES_ENC/n11510 ), .ZN(\AES_ENC/n743 ) );
NAND2_X2 \AES_ENC/U153  ( .A1(aes_text_in[83]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n11210 ) );
NAND2_X2 \AES_ENC/U152  ( .A1(\AES_ENC/text_in_r[83] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n11310 ) );
NAND2_X2 \AES_ENC/U151  ( .A1(\AES_ENC/n11210 ), .A2(\AES_ENC/n11310 ), .ZN(\AES_ENC/n744 ) );
NAND2_X2 \AES_ENC/U150  ( .A1(aes_text_in[84]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n11010 ) );
NAND2_X2 \AES_ENC/U149  ( .A1(\AES_ENC/text_in_r[84] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n11110 ) );
NAND2_X2 \AES_ENC/U148  ( .A1(\AES_ENC/n11010 ), .A2(\AES_ENC/n11110 ), .ZN(\AES_ENC/n745 ) );
NAND2_X2 \AES_ENC/U147  ( .A1(aes_text_in[85]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n108 ) );
NAND2_X2 \AES_ENC/U146  ( .A1(\AES_ENC/text_in_r[85] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n109 ) );
NAND2_X2 \AES_ENC/U145  ( .A1(\AES_ENC/n108 ), .A2(\AES_ENC/n109 ), .ZN(\AES_ENC/n746 ) );
NAND2_X2 \AES_ENC/U144  ( .A1(aes_text_in[86]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n106 ) );
NAND2_X2 \AES_ENC/U143  ( .A1(\AES_ENC/text_in_r[86] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n107 ) );
NAND2_X2 \AES_ENC/U142  ( .A1(\AES_ENC/n106 ), .A2(\AES_ENC/n107 ), .ZN(\AES_ENC/n747 ) );
NAND2_X2 \AES_ENC/U141  ( .A1(aes_text_in[87]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n104 ) );
NAND2_X2 \AES_ENC/U140  ( .A1(\AES_ENC/text_in_r[87] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n105 ) );
NAND2_X2 \AES_ENC/U139  ( .A1(\AES_ENC/n104 ), .A2(\AES_ENC/n105 ), .ZN(\AES_ENC/n748 ) );
NAND2_X2 \AES_ENC/U138  ( .A1(aes_text_in[88]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n102 ) );
NAND2_X2 \AES_ENC/U137  ( .A1(\AES_ENC/text_in_r[88] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n103 ) );
NAND2_X2 \AES_ENC/U136  ( .A1(\AES_ENC/n102 ), .A2(\AES_ENC/n103 ), .ZN(\AES_ENC/n749 ) );
NAND2_X2 \AES_ENC/U135  ( .A1(aes_text_in[89]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n10010 ) );
NAND2_X2 \AES_ENC/U134  ( .A1(\AES_ENC/text_in_r[89] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n10110 ) );
NAND2_X2 \AES_ENC/U133  ( .A1(\AES_ENC/n10010 ), .A2(\AES_ENC/n10110 ), .ZN(\AES_ENC/n750 ) );
NAND2_X2 \AES_ENC/U132  ( .A1(aes_text_in[90]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n9810 ) );
NAND2_X2 \AES_ENC/U131  ( .A1(\AES_ENC/text_in_r[90] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n9910 ) );
NAND2_X2 \AES_ENC/U130  ( .A1(\AES_ENC/n9810 ), .A2(\AES_ENC/n9910 ), .ZN(\AES_ENC/n751 ) );
NAND2_X2 \AES_ENC/U129  ( .A1(aes_text_in[91]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n9610 ) );
NAND2_X2 \AES_ENC/U128  ( .A1(\AES_ENC/text_in_r[91] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n9710 ) );
NAND2_X2 \AES_ENC/U127  ( .A1(\AES_ENC/n9610 ), .A2(\AES_ENC/n9710 ), .ZN(\AES_ENC/n752 ) );
NAND2_X2 \AES_ENC/U126  ( .A1(aes_text_in[92]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n9410 ) );
NAND2_X2 \AES_ENC/U125  ( .A1(\AES_ENC/text_in_r[92] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n9510 ) );
NAND2_X2 \AES_ENC/U124  ( .A1(\AES_ENC/n9410 ), .A2(\AES_ENC/n9510 ), .ZN(\AES_ENC/n753 ) );
NAND2_X2 \AES_ENC/U123  ( .A1(aes_text_in[93]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n92 ) );
NAND2_X2 \AES_ENC/U122  ( .A1(\AES_ENC/text_in_r[93] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n93 ) );
NAND2_X2 \AES_ENC/U121  ( .A1(\AES_ENC/n92 ), .A2(\AES_ENC/n93 ), .ZN(\AES_ENC/n754 ) );
NAND2_X2 \AES_ENC/U120  ( .A1(aes_text_in[94]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n90 ) );
NAND2_X2 \AES_ENC/U119  ( .A1(\AES_ENC/text_in_r[94] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n91 ) );
NAND2_X2 \AES_ENC/U118  ( .A1(\AES_ENC/n90 ), .A2(\AES_ENC/n91 ), .ZN(\AES_ENC/n755 ) );
NAND2_X2 \AES_ENC/U117  ( .A1(aes_text_in[95]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n88 ) );
NAND2_X2 \AES_ENC/U116  ( .A1(\AES_ENC/text_in_r[95] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n89 ) );
NAND2_X2 \AES_ENC/U115  ( .A1(\AES_ENC/n88 ), .A2(\AES_ENC/n89 ), .ZN(\AES_ENC/n756 ) );
NAND2_X2 \AES_ENC/U114  ( .A1(aes_text_in[96]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n86 ) );
NAND2_X2 \AES_ENC/U113  ( .A1(\AES_ENC/text_in_r[96] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n87 ) );
NAND2_X2 \AES_ENC/U112  ( .A1(\AES_ENC/n86 ), .A2(\AES_ENC/n87 ), .ZN(\AES_ENC/n757 ) );
NAND2_X2 \AES_ENC/U111  ( .A1(aes_text_in[97]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n8410 ) );
NAND2_X2 \AES_ENC/U110  ( .A1(\AES_ENC/text_in_r[97] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n8510 ) );
NAND2_X2 \AES_ENC/U109  ( .A1(\AES_ENC/n8410 ), .A2(\AES_ENC/n8510 ), .ZN(\AES_ENC/n758 ) );
NAND2_X2 \AES_ENC/U108  ( .A1(aes_text_in[98]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n8210 ) );
NAND2_X2 \AES_ENC/U107  ( .A1(\AES_ENC/text_in_r[98] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n8310 ) );
NAND2_X2 \AES_ENC/U106  ( .A1(\AES_ENC/n8210 ), .A2(\AES_ENC/n8310 ), .ZN(\AES_ENC/n759 ) );
NAND2_X2 \AES_ENC/U105  ( .A1(aes_text_in[99]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n8010 ) );
NAND2_X2 \AES_ENC/U104  ( .A1(\AES_ENC/text_in_r[99] ), .A2(\AES_ENC/n1261 ),.ZN(\AES_ENC/n8110 ) );
NAND2_X2 \AES_ENC/U103  ( .A1(\AES_ENC/n8010 ), .A2(\AES_ENC/n8110 ), .ZN(\AES_ENC/n760 ) );
NAND2_X2 \AES_ENC/U102  ( .A1(aes_text_in[100]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n7890 ) );
NAND2_X2 \AES_ENC/U101  ( .A1(\AES_ENC/text_in_r[100] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n7900 ) );
NAND2_X2 \AES_ENC/U100  ( .A1(\AES_ENC/n7890 ), .A2(\AES_ENC/n7900 ), .ZN(\AES_ENC/n761 ) );
NAND2_X2 \AES_ENC/U99  ( .A1(aes_text_in[101]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n76 ) );
NAND2_X2 \AES_ENC/U98  ( .A1(\AES_ENC/text_in_r[101] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n77 ) );
NAND2_X2 \AES_ENC/U97  ( .A1(\AES_ENC/n76 ), .A2(\AES_ENC/n77 ), .ZN(\AES_ENC/n762 ) );
NAND2_X2 \AES_ENC/U96  ( .A1(aes_text_in[102]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n74 ) );
NAND2_X2 \AES_ENC/U95  ( .A1(\AES_ENC/text_in_r[102] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n75 ) );
NAND2_X2 \AES_ENC/U94  ( .A1(\AES_ENC/n74 ), .A2(\AES_ENC/n75 ), .ZN(\AES_ENC/n763 ) );
NAND2_X2 \AES_ENC/U93  ( .A1(aes_text_in[103]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n72 ) );
NAND2_X2 \AES_ENC/U92  ( .A1(\AES_ENC/text_in_r[103] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n73 ) );
NAND2_X2 \AES_ENC/U91  ( .A1(\AES_ENC/n72 ), .A2(\AES_ENC/n73 ), .ZN(\AES_ENC/n764 ) );
NAND2_X2 \AES_ENC/U90  ( .A1(aes_text_in[104]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n70 ) );
NAND2_X2 \AES_ENC/U89  ( .A1(\AES_ENC/text_in_r[104] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n71 ) );
NAND2_X2 \AES_ENC/U88  ( .A1(\AES_ENC/n70 ), .A2(\AES_ENC/n71 ), .ZN(\AES_ENC/n765 ) );
NAND2_X2 \AES_ENC/U87  ( .A1(aes_text_in[105]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n6810 ) );
NAND2_X2 \AES_ENC/U86  ( .A1(\AES_ENC/text_in_r[105] ), .A2(\AES_ENC/n12601 ), .ZN(\AES_ENC/n6910 ) );
NAND2_X2 \AES_ENC/U85  ( .A1(\AES_ENC/n6810 ), .A2(\AES_ENC/n6910 ), .ZN(\AES_ENC/n766 ) );
NAND2_X2 \AES_ENC/U84  ( .A1(aes_text_in[106]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n6600 ) );
NAND2_X2 \AES_ENC/U83  ( .A1(\AES_ENC/text_in_r[106] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n6710 ) );
NAND2_X2 \AES_ENC/U82  ( .A1(\AES_ENC/n6600 ), .A2(\AES_ENC/n6710 ), .ZN(\AES_ENC/n767 ) );
NAND2_X2 \AES_ENC/U81  ( .A1(aes_text_in[107]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n6400 ) );
NAND2_X2 \AES_ENC/U80  ( .A1(\AES_ENC/text_in_r[107] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n6500 ) );
NAND2_X2 \AES_ENC/U79  ( .A1(\AES_ENC/n6400 ), .A2(\AES_ENC/n6500 ), .ZN(\AES_ENC/n768 ) );
NAND2_X2 \AES_ENC/U78  ( .A1(aes_text_in[108]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n6200 ) );
NAND2_X2 \AES_ENC/U77  ( .A1(\AES_ENC/text_in_r[108] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n6300 ) );
NAND2_X2 \AES_ENC/U76  ( .A1(\AES_ENC/n6200 ), .A2(\AES_ENC/n6300 ), .ZN(\AES_ENC/n769 ) );
NAND2_X2 \AES_ENC/U75  ( .A1(aes_text_in[109]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n60 ) );
NAND2_X2 \AES_ENC/U74  ( .A1(\AES_ENC/text_in_r[109] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n61 ) );
NAND2_X2 \AES_ENC/U73  ( .A1(\AES_ENC/n60 ), .A2(\AES_ENC/n61 ), .ZN(\AES_ENC/n770 ) );
NAND2_X2 \AES_ENC/U72  ( .A1(aes_text_in[110]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n58 ) );
NAND2_X2 \AES_ENC/U71  ( .A1(\AES_ENC/text_in_r[110] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n59 ) );
NAND2_X2 \AES_ENC/U70  ( .A1(\AES_ENC/n58 ), .A2(\AES_ENC/n59 ), .ZN(\AES_ENC/n771 ) );
NAND2_X2 \AES_ENC/U69  ( .A1(aes_text_in[111]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n56 ) );
NAND2_X2 \AES_ENC/U68  ( .A1(\AES_ENC/text_in_r[111] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n57 ) );
NAND2_X2 \AES_ENC/U67  ( .A1(\AES_ENC/n56 ), .A2(\AES_ENC/n57 ), .ZN(\AES_ENC/n772 ) );
NAND2_X2 \AES_ENC/U66  ( .A1(aes_text_in[112]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n54 ) );
NAND2_X2 \AES_ENC/U65  ( .A1(\AES_ENC/text_in_r[112] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n55 ) );
NAND2_X2 \AES_ENC/U64  ( .A1(\AES_ENC/n54 ), .A2(\AES_ENC/n55 ), .ZN(\AES_ENC/n773 ) );
NAND2_X2 \AES_ENC/U63  ( .A1(aes_text_in[113]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n5200 ) );
NAND2_X2 \AES_ENC/U62  ( .A1(\AES_ENC/text_in_r[113] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n5300 ) );
NAND2_X2 \AES_ENC/U61  ( .A1(\AES_ENC/n5200 ), .A2(\AES_ENC/n5300 ), .ZN(\AES_ENC/n774 ) );
NAND2_X2 \AES_ENC/U60  ( .A1(aes_text_in[114]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n5020 ) );
NAND2_X2 \AES_ENC/U59  ( .A1(\AES_ENC/text_in_r[114] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n5100 ) );
NAND2_X2 \AES_ENC/U58  ( .A1(\AES_ENC/n5020 ), .A2(\AES_ENC/n5100 ), .ZN(\AES_ENC/n775 ) );
NAND2_X2 \AES_ENC/U57  ( .A1(aes_text_in[115]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n4810 ) );
NAND2_X2 \AES_ENC/U56  ( .A1(\AES_ENC/text_in_r[115] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n4910 ) );
NAND2_X2 \AES_ENC/U55  ( .A1(\AES_ENC/n4810 ), .A2(\AES_ENC/n4910 ), .ZN(\AES_ENC/n776 ) );
NAND2_X2 \AES_ENC/U54  ( .A1(aes_text_in[116]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n4610 ) );
NAND2_X2 \AES_ENC/U53  ( .A1(\AES_ENC/text_in_r[116] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n4710 ) );
NAND2_X2 \AES_ENC/U52  ( .A1(\AES_ENC/n4610 ), .A2(\AES_ENC/n4710 ), .ZN(\AES_ENC/n777 ) );
NAND2_X2 \AES_ENC/U51  ( .A1(aes_text_in[117]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n44 ) );
NAND2_X2 \AES_ENC/U50  ( .A1(\AES_ENC/text_in_r[117] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n45 ) );
NAND2_X2 \AES_ENC/U49  ( .A1(\AES_ENC/n44 ), .A2(\AES_ENC/n45 ), .ZN(\AES_ENC/n778 ) );
NAND2_X2 \AES_ENC/U48  ( .A1(aes_text_in[118]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n42 ) );
NAND2_X2 \AES_ENC/U47  ( .A1(\AES_ENC/text_in_r[118] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n43 ) );
NAND2_X2 \AES_ENC/U46  ( .A1(\AES_ENC/n42 ), .A2(\AES_ENC/n43 ), .ZN(\AES_ENC/n779 ) );
NAND2_X2 \AES_ENC/U45  ( .A1(aes_text_in[119]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n40 ) );
NAND2_X2 \AES_ENC/U44  ( .A1(\AES_ENC/text_in_r[119] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n41 ) );
NAND2_X2 \AES_ENC/U43  ( .A1(\AES_ENC/n40 ), .A2(\AES_ENC/n41 ), .ZN(\AES_ENC/n780 ) );
NAND2_X2 \AES_ENC/U42  ( .A1(aes_text_in[120]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n38 ) );
NAND2_X2 \AES_ENC/U41  ( .A1(\AES_ENC/text_in_r[120] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n39 ) );
NAND2_X2 \AES_ENC/U40  ( .A1(\AES_ENC/n38 ), .A2(\AES_ENC/n39 ), .ZN(\AES_ENC/n781 ) );
NAND2_X2 \AES_ENC/U39  ( .A1(aes_text_in[121]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n3600 ) );
NAND2_X2 \AES_ENC/U38  ( .A1(\AES_ENC/text_in_r[121] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n3700 ) );
NAND2_X2 \AES_ENC/U37  ( .A1(\AES_ENC/n3600 ), .A2(\AES_ENC/n3700 ), .ZN(\AES_ENC/n782 ) );
NAND2_X2 \AES_ENC/U36  ( .A1(aes_text_in[122]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n3400 ) );
NAND2_X2 \AES_ENC/U35  ( .A1(\AES_ENC/text_in_r[122] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n3500 ) );
NAND2_X2 \AES_ENC/U34  ( .A1(\AES_ENC/n3400 ), .A2(\AES_ENC/n3500 ), .ZN(\AES_ENC/n783 ) );
NAND2_X2 \AES_ENC/U33  ( .A1(aes_text_in[123]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n3200 ) );
NAND2_X2 \AES_ENC/U32  ( .A1(\AES_ENC/text_in_r[123] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n3300 ) );
NAND2_X2 \AES_ENC/U31  ( .A1(\AES_ENC/n3200 ), .A2(\AES_ENC/n3300 ), .ZN(\AES_ENC/n784 ) );
NAND2_X2 \AES_ENC/U30  ( .A1(aes_text_in[124]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n3000 ) );
NAND2_X2 \AES_ENC/U29  ( .A1(\AES_ENC/text_in_r[124] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n3100 ) );
NAND2_X2 \AES_ENC/U28  ( .A1(\AES_ENC/n3000 ), .A2(\AES_ENC/n3100 ), .ZN(\AES_ENC/n785 ) );
NAND2_X2 \AES_ENC/U27  ( .A1(aes_text_in[125]), .A2(\AES_ENC/n1235 ), .ZN(\AES_ENC/n28 ) );
NAND2_X2 \AES_ENC/U26  ( .A1(\AES_ENC/text_in_r[125] ), .A2(\AES_ENC/n1259 ),.ZN(\AES_ENC/n29 ) );
NAND2_X2 \AES_ENC/U25  ( .A1(\AES_ENC/n28 ), .A2(\AES_ENC/n29 ), .ZN(\AES_ENC/n786 ) );
NAND2_X2 \AES_ENC/U24  ( .A1(aes_text_in[126]), .A2(\AES_ENC/n1236 ), .ZN(\AES_ENC/n26 ) );
NAND2_X2 \AES_ENC/U23  ( .A1(\AES_ENC/text_in_r[126] ), .A2(\AES_ENC/n1258 ),.ZN(\AES_ENC/n27 ) );
NAND2_X2 \AES_ENC/U22  ( .A1(\AES_ENC/n26 ), .A2(\AES_ENC/n27 ), .ZN(\AES_ENC/n787 ) );
NAND2_X2 \AES_ENC/U21  ( .A1(aes_text_in[127]), .A2(\AES_ENC/n1237 ), .ZN(\AES_ENC/n24 ) );
NAND2_X2 \AES_ENC/U20  ( .A1(\AES_ENC/text_in_r[127] ), .A2(\AES_ENC/n1258 ),.ZN(\AES_ENC/n25 ) );
NAND2_X2 \AES_ENC/U19  ( .A1(\AES_ENC/n24 ), .A2(\AES_ENC/n25 ), .ZN(\AES_ENC/n788 ) );
NAND2_X2 \AES_ENC/U18  ( .A1(\AES_ENC/n792 ), .A2(\AES_ENC/n14 ), .ZN(\AES_ENC/n23 ) );
NAND2_X2 \AES_ENC/U17  ( .A1(\AES_ENC/n1258 ), .A2(\AES_ENC/n23 ), .ZN(\AES_ENC/n22 ) );
NAND2_X2 \AES_ENC/U15  ( .A1(\AES_ENC/n11 ), .A2(\AES_ENC/n14 ), .ZN(\AES_ENC/n18 ) );
NAND2_X2 \AES_ENC/U13  ( .A1(\AES_ENC/n1258 ), .A2(\AES_ENC/n1231 ), .ZN(\AES_ENC/n21 ) );
NAND2_X2 \AES_ENC/U12  ( .A1(\AES_ENC/n1266 ), .A2(\AES_ENC/n21 ), .ZN(\AES_ENC/n20 ) );
NAND2_X2 \AES_ENC/U11  ( .A1(\AES_ENC/n20 ), .A2(\AES_ENC/n1234 ), .ZN(\AES_ENC/n1980 ) );
NAND2_X2 \AES_ENC/U10  ( .A1(\AES_ENC/n18 ), .A2(\AES_ENC/n1980 ), .ZN(\AES_ENC/n795 ) );
NAND2_X2 \AES_ENC/U9  ( .A1(\AES_ENC/n17 ), .A2(\AES_ENC/n1231 ), .ZN(\AES_ENC/n15 ) );
NAND2_X2 \AES_ENC/U8  ( .A1(\AES_ENC/n11 ), .A2(\AES_ENC/n794 ), .ZN(\AES_ENC/n16 ) );
NAND2_X2 \AES_ENC/U6  ( .A1(\AES_ENC/n14 ), .A2(\AES_ENC/n1266 ), .ZN(\AES_ENC/n13 ) );
NAND2_X2 \AES_ENC/U5  ( .A1(\AES_ENC/n13 ), .A2(\AES_ENC/n1233 ), .ZN(\AES_ENC/n12 ) );
NAND2_X2 \AES_ENC/U4  ( .A1(\AES_ENC/n1258 ), .A2(\AES_ENC/n12 ), .ZN(\AES_ENC/n797 ) );
OR2_X2 \AES_ENC/U3  ( .A1(\AES_ENC/n1257 ), .A2(\AES_ENC/n11 ), .ZN(\AES_ENC/n798 ) );
DFF_X2 \AES_ENC/text_out_reg_0_  ( .D(\AES_ENC/N501 ), .CK(clk), .Q(aes_text_out[0]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_1_  ( .D(\AES_ENC/N500 ), .CK(clk), .Q(aes_text_out[1]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_2_  ( .D(\AES_ENC/N499 ), .CK(clk), .Q(aes_text_out[2]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_3_  ( .D(\AES_ENC/N498 ), .CK(clk), .Q(aes_text_out[3]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_4_  ( .D(\AES_ENC/N497 ), .CK(clk), .Q(aes_text_out[4]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_5_  ( .D(\AES_ENC/N496 ), .CK(clk), .Q(aes_text_out[5]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_6_  ( .D(\AES_ENC/N495 ), .CK(clk), .Q(aes_text_out[6]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_7_  ( .D(\AES_ENC/N494 ), .CK(clk), .Q(aes_text_out[7]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_8_  ( .D(\AES_ENC/N469 ), .CK(clk), .Q(aes_text_out[8]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_9_  ( .D(\AES_ENC/N468 ), .CK(clk), .Q(aes_text_out[9]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_10_  ( .D(\AES_ENC/N467 ), .CK(clk), .Q(aes_text_out[10]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_11_  ( .D(\AES_ENC/N466 ), .CK(clk), .Q(aes_text_out[11]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_12_  ( .D(\AES_ENC/N465 ), .CK(clk), .Q(aes_text_out[12]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_13_  ( .D(\AES_ENC/N464 ), .CK(clk), .Q(aes_text_out[13]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_14_  ( .D(\AES_ENC/N463 ), .CK(clk), .Q(aes_text_out[14]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_15_  ( .D(\AES_ENC/N462 ), .CK(clk), .Q(aes_text_out[15]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_16_  ( .D(\AES_ENC/N437 ), .CK(clk), .Q(aes_text_out[16]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_17_  ( .D(\AES_ENC/N436 ), .CK(clk), .Q(aes_text_out[17]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_18_  ( .D(\AES_ENC/N435 ), .CK(clk), .Q(aes_text_out[18]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_19_  ( .D(\AES_ENC/N434 ), .CK(clk), .Q(aes_text_out[19]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_20_  ( .D(\AES_ENC/N433 ), .CK(clk), .Q(aes_text_out[20]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_21_  ( .D(\AES_ENC/N432 ), .CK(clk), .Q(aes_text_out[21]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_22_  ( .D(\AES_ENC/N431 ), .CK(clk), .Q(aes_text_out[22]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_23_  ( .D(\AES_ENC/N430 ), .CK(clk), .Q(aes_text_out[23]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_24_  ( .D(\AES_ENC/N405 ), .CK(clk), .Q(aes_text_out[24]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_25_  ( .D(\AES_ENC/N404 ), .CK(clk), .Q(aes_text_out[25]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_26_  ( .D(\AES_ENC/N403 ), .CK(clk), .Q(aes_text_out[26]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_27_  ( .D(\AES_ENC/N402 ), .CK(clk), .Q(aes_text_out[27]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_28_  ( .D(\AES_ENC/N401 ), .CK(clk), .Q(aes_text_out[28]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_29_  ( .D(\AES_ENC/N400 ), .CK(clk), .Q(aes_text_out[29]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_30_  ( .D(\AES_ENC/N399 ), .CK(clk), .Q(aes_text_out[30]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_31_  ( .D(\AES_ENC/N398 ), .CK(clk), .Q(aes_text_out[31]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_32_  ( .D(\AES_ENC/N493 ), .CK(clk), .Q(aes_text_out[32]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_33_  ( .D(\AES_ENC/N492 ), .CK(clk), .Q(aes_text_out[33]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_34_  ( .D(\AES_ENC/N491 ), .CK(clk), .Q(aes_text_out[34]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_35_  ( .D(\AES_ENC/N490 ), .CK(clk), .Q(aes_text_out[35]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_36_  ( .D(\AES_ENC/N489 ), .CK(clk), .Q(aes_text_out[36]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_37_  ( .D(\AES_ENC/N488 ), .CK(clk), .Q(aes_text_out[37]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_38_  ( .D(\AES_ENC/N487 ), .CK(clk), .Q(aes_text_out[38]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_39_  ( .D(\AES_ENC/N486 ), .CK(clk), .Q(aes_text_out[39]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_40_  ( .D(\AES_ENC/N461 ), .CK(clk), .Q(aes_text_out[40]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_41_  ( .D(\AES_ENC/N460 ), .CK(clk), .Q(aes_text_out[41]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_42_  ( .D(\AES_ENC/N459 ), .CK(clk), .Q(aes_text_out[42]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_43_  ( .D(\AES_ENC/N458 ), .CK(clk), .Q(aes_text_out[43]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_44_  ( .D(\AES_ENC/N457 ), .CK(clk), .Q(aes_text_out[44]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_45_  ( .D(\AES_ENC/N456 ), .CK(clk), .Q(aes_text_out[45]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_46_  ( .D(\AES_ENC/N455 ), .CK(clk), .Q(aes_text_out[46]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_47_  ( .D(\AES_ENC/N454 ), .CK(clk), .Q(aes_text_out[47]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_48_  ( .D(\AES_ENC/N429 ), .CK(clk), .Q(aes_text_out[48]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_49_  ( .D(\AES_ENC/N428 ), .CK(clk), .Q(aes_text_out[49]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_50_  ( .D(\AES_ENC/N427 ), .CK(clk), .Q(aes_text_out[50]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_51_  ( .D(\AES_ENC/N426 ), .CK(clk), .Q(aes_text_out[51]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_52_  ( .D(\AES_ENC/N425 ), .CK(clk), .Q(aes_text_out[52]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_53_  ( .D(\AES_ENC/N424 ), .CK(clk), .Q(aes_text_out[53]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_54_  ( .D(\AES_ENC/N423 ), .CK(clk), .Q(aes_text_out[54]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_55_  ( .D(\AES_ENC/N422 ), .CK(clk), .Q(aes_text_out[55]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_56_  ( .D(\AES_ENC/N397 ), .CK(clk), .Q(aes_text_out[56]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_57_  ( .D(\AES_ENC/N396 ), .CK(clk), .Q(aes_text_out[57]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_58_  ( .D(\AES_ENC/N395 ), .CK(clk), .Q(aes_text_out[58]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_59_  ( .D(\AES_ENC/N394 ), .CK(clk), .Q(aes_text_out[59]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_60_  ( .D(\AES_ENC/N393 ), .CK(clk), .Q(aes_text_out[60]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_61_  ( .D(\AES_ENC/N392 ), .CK(clk), .Q(aes_text_out[61]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_62_  ( .D(\AES_ENC/N391 ), .CK(clk), .Q(aes_text_out[62]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_63_  ( .D(\AES_ENC/N390 ), .CK(clk), .Q(aes_text_out[63]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_64_  ( .D(\AES_ENC/N485 ), .CK(clk), .Q(aes_text_out[64]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_65_  ( .D(\AES_ENC/N484 ), .CK(clk), .Q(aes_text_out[65]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_66_  ( .D(\AES_ENC/N483 ), .CK(clk), .Q(aes_text_out[66]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_67_  ( .D(\AES_ENC/N482 ), .CK(clk), .Q(aes_text_out[67]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_68_  ( .D(\AES_ENC/N481 ), .CK(clk), .Q(aes_text_out[68]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_69_  ( .D(\AES_ENC/N480 ), .CK(clk), .Q(aes_text_out[69]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_70_  ( .D(\AES_ENC/N479 ), .CK(clk), .Q(aes_text_out[70]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_71_  ( .D(\AES_ENC/N478 ), .CK(clk), .Q(aes_text_out[71]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_72_  ( .D(\AES_ENC/N453 ), .CK(clk), .Q(aes_text_out[72]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_73_  ( .D(\AES_ENC/N452 ), .CK(clk), .Q(aes_text_out[73]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_74_  ( .D(\AES_ENC/N451 ), .CK(clk), .Q(aes_text_out[74]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_75_  ( .D(\AES_ENC/N450 ), .CK(clk), .Q(aes_text_out[75]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_76_  ( .D(\AES_ENC/N449 ), .CK(clk), .Q(aes_text_out[76]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_77_  ( .D(\AES_ENC/N448 ), .CK(clk), .Q(aes_text_out[77]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_78_  ( .D(\AES_ENC/N447 ), .CK(clk), .Q(aes_text_out[78]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_79_  ( .D(\AES_ENC/N446 ), .CK(clk), .Q(aes_text_out[79]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_80_  ( .D(\AES_ENC/N421 ), .CK(clk), .Q(aes_text_out[80]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_81_  ( .D(\AES_ENC/N420 ), .CK(clk), .Q(aes_text_out[81]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_82_  ( .D(\AES_ENC/N419 ), .CK(clk), .Q(aes_text_out[82]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_83_  ( .D(\AES_ENC/N418 ), .CK(clk), .Q(aes_text_out[83]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_84_  ( .D(\AES_ENC/N417 ), .CK(clk), .Q(aes_text_out[84]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_85_  ( .D(\AES_ENC/N416 ), .CK(clk), .Q(aes_text_out[85]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_86_  ( .D(\AES_ENC/N415 ), .CK(clk), .Q(aes_text_out[86]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_87_  ( .D(\AES_ENC/N414 ), .CK(clk), .Q(aes_text_out[87]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_88_  ( .D(\AES_ENC/N389 ), .CK(clk), .Q(aes_text_out[88]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_89_  ( .D(\AES_ENC/N388 ), .CK(clk), .Q(aes_text_out[89]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_90_  ( .D(\AES_ENC/N387 ), .CK(clk), .Q(aes_text_out[90]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_91_  ( .D(\AES_ENC/N386 ), .CK(clk), .Q(aes_text_out[91]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_92_  ( .D(\AES_ENC/N385 ), .CK(clk), .Q(aes_text_out[92]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_93_  ( .D(\AES_ENC/N384 ), .CK(clk), .Q(aes_text_out[93]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_94_  ( .D(\AES_ENC/N383 ), .CK(clk), .Q(aes_text_out[94]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_95_  ( .D(\AES_ENC/N382 ), .CK(clk), .Q(aes_text_out[95]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_96_  ( .D(\AES_ENC/N477 ), .CK(clk), .Q(aes_text_out[96]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_97_  ( .D(\AES_ENC/N476 ), .CK(clk), .Q(aes_text_out[97]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_98_  ( .D(\AES_ENC/N475 ), .CK(clk), .Q(aes_text_out[98]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_99_  ( .D(\AES_ENC/N474 ), .CK(clk), .Q(aes_text_out[99]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_100_  ( .D(\AES_ENC/N473 ), .CK(clk), .Q(aes_text_out[100]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_101_  ( .D(\AES_ENC/N472 ), .CK(clk), .Q(aes_text_out[101]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_102_  ( .D(\AES_ENC/N471 ), .CK(clk), .Q(aes_text_out[102]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_103_  ( .D(\AES_ENC/N470 ), .CK(clk), .Q(aes_text_out[103]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_104_  ( .D(\AES_ENC/N445 ), .CK(clk), .Q(aes_text_out[104]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_105_  ( .D(\AES_ENC/N444 ), .CK(clk), .Q(aes_text_out[105]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_106_  ( .D(\AES_ENC/N443 ), .CK(clk), .Q(aes_text_out[106]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_107_  ( .D(\AES_ENC/N442 ), .CK(clk), .Q(aes_text_out[107]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_108_  ( .D(\AES_ENC/N441 ), .CK(clk), .Q(aes_text_out[108]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_109_  ( .D(\AES_ENC/N440 ), .CK(clk), .Q(aes_text_out[109]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_110_  ( .D(\AES_ENC/N439 ), .CK(clk), .Q(aes_text_out[110]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_111_  ( .D(\AES_ENC/N438 ), .CK(clk), .Q(aes_text_out[111]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_112_  ( .D(\AES_ENC/N413 ), .CK(clk), .Q(aes_text_out[112]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_113_  ( .D(\AES_ENC/N412 ), .CK(clk), .Q(aes_text_out[113]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_114_  ( .D(\AES_ENC/N411 ), .CK(clk), .Q(aes_text_out[114]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_115_  ( .D(\AES_ENC/N410 ), .CK(clk), .Q(aes_text_out[115]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_116_  ( .D(\AES_ENC/N409 ), .CK(clk), .Q(aes_text_out[116]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_117_  ( .D(\AES_ENC/N408 ), .CK(clk), .Q(aes_text_out[117]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_118_  ( .D(\AES_ENC/N407 ), .CK(clk), .Q(aes_text_out[118]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_119_  ( .D(\AES_ENC/N406 ), .CK(clk), .Q(aes_text_out[119]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_120_  ( .D(\AES_ENC/N381 ), .CK(clk), .Q(aes_text_out[120]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_121_  ( .D(\AES_ENC/N380 ), .CK(clk), .Q(aes_text_out[121]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_122_  ( .D(\AES_ENC/N379 ), .CK(clk), .Q(aes_text_out[122]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_123_  ( .D(\AES_ENC/N378 ), .CK(clk), .Q(aes_text_out[123]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_124_  ( .D(\AES_ENC/N377 ), .CK(clk), .Q(aes_text_out[124]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_125_  ( .D(\AES_ENC/N376 ), .CK(clk), .Q(aes_text_out[125]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_126_  ( .D(\AES_ENC/N375 ), .CK(clk), .Q(aes_text_out[126]), .QN() );
DFF_X2 \AES_ENC/text_out_reg_127_  ( .D(\AES_ENC/N374 ), .CK(clk), .Q(aes_text_out[127]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_7_  ( .D(\AES_ENC/N101 ), .CK(clk), .Q(\AES_ENC/sa32 [7]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_7_  ( .D(\AES_ENC/N229 ), .CK(clk), .Q(\AES_ENC/sa30 [7]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_0_  ( .D(\AES_ENC/N238 ), .CK(clk), .Q(\AES_ENC/sa20 [0]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_1_  ( .D(\AES_ENC/N239 ), .CK(clk), .Q(\AES_ENC/sa20 [1]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_3_  ( .D(\AES_ENC/N241 ), .CK(clk), .Q(\AES_ENC/sa20 [3]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_4_  ( .D(\AES_ENC/N242 ), .CK(clk), .Q(\AES_ENC/sa20 [4]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_7_  ( .D(\AES_ENC/N261 ), .CK(clk), .Q(\AES_ENC/sa10 [7]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_7_  ( .D(\AES_ENC/N277 ), .CK(clk), .Q(\AES_ENC/sa00 [7]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_6_  ( .D(\AES_ENC/N228 ), .CK(clk), .Q(\AES_ENC/sa30 [6]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_6_  ( .D(\AES_ENC/N260 ), .CK(clk), .Q(\AES_ENC/sa10 [6]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_6_  ( .D(\AES_ENC/N276 ), .CK(clk), .Q(\AES_ENC/sa00 [6]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_5_  ( .D(\AES_ENC/N227 ), .CK(clk), .Q(\AES_ENC/sa30 [5]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_6_  ( .D(\AES_ENC/N244 ), .CK(clk), .Q(\AES_ENC/sa20 [6]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_5_  ( .D(\AES_ENC/N259 ), .CK(clk), .Q(\AES_ENC/sa10 [5]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_5_  ( .D(\AES_ENC/N275 ), .CK(clk), .Q(\AES_ENC/sa00 [5]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_4_  ( .D(\AES_ENC/N226 ), .CK(clk), .Q(\AES_ENC/sa30 [4]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_5_  ( .D(\AES_ENC/N243 ), .CK(clk), .Q(\AES_ENC/sa20 [5]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_4_  ( .D(\AES_ENC/N258 ), .CK(clk), .Q(\AES_ENC/sa10 [4]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_4_  ( .D(\AES_ENC/N274 ), .CK(clk), .Q(\AES_ENC/sa00 [4]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_3_  ( .D(\AES_ENC/N225 ), .CK(clk), .Q(\AES_ENC/sa30 [3]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_3_  ( .D(\AES_ENC/N257 ), .CK(clk), .Q(\AES_ENC/sa10 [3]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_3_  ( .D(\AES_ENC/N273 ), .CK(clk), .Q(\AES_ENC/sa00 [3]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_2_  ( .D(\AES_ENC/N224 ), .CK(clk), .Q(\AES_ENC/sa30 [2]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_2_  ( .D(\AES_ENC/N256 ), .CK(clk), .Q(\AES_ENC/sa10 [2]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_2_  ( .D(\AES_ENC/N272 ), .CK(clk), .Q(\AES_ENC/sa00 [2]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_1_  ( .D(\AES_ENC/N223 ), .CK(clk), .Q(\AES_ENC/sa30 [1]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_2_  ( .D(\AES_ENC/N240 ), .CK(clk), .Q(\AES_ENC/sa20 [2]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_1_  ( .D(\AES_ENC/N255 ), .CK(clk), .Q(\AES_ENC/sa10 [1]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_1_  ( .D(\AES_ENC/N271 ), .CK(clk), .Q(\AES_ENC/sa00 [1]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_7_  ( .D(\AES_ENC/N117 ), .CK(clk), .Q(\AES_ENC/sa22 [7]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_7_  ( .D(\AES_ENC/N133 ), .CK(clk), .Q(\AES_ENC/sa12 [7]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_6_  ( .D(\AES_ENC/N132 ), .CK(clk), .Q(\AES_ENC/sa12 [6]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_6_  ( .D(\AES_ENC/N100 ), .CK(clk), .Q(\AES_ENC/sa32 [6]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_6_  ( .D(\AES_ENC/N116 ), .CK(clk), .Q(\AES_ENC/sa22 [6]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_7_  ( .D(\AES_ENC/N149 ), .CK(clk), .Q(\AES_ENC/sa02 [7]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_5_  ( .D(\AES_ENC/N131 ), .CK(clk), .Q(\AES_ENC/sa12 [5]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_5_  ( .D(\AES_ENC/N99 ), .CK(clk), .Q(\AES_ENC/sa32 [5]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_5_  ( .D(\AES_ENC/N115 ), .CK(clk), .Q(\AES_ENC/sa22 [5]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_6_  ( .D(\AES_ENC/N148 ), .CK(clk), .Q(\AES_ENC/sa02 [6]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_4_  ( .D(\AES_ENC/N130 ), .CK(clk), .Q(\AES_ENC/sa12 [4]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_4_  ( .D(\AES_ENC/N98 ), .CK(clk), .Q(\AES_ENC/sa32 [4]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_4_  ( .D(\AES_ENC/N114 ), .CK(clk), .Q(\AES_ENC/sa22 [4]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_5_  ( .D(\AES_ENC/N147 ), .CK(clk), .Q(\AES_ENC/sa02 [5]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_3_  ( .D(\AES_ENC/N129 ), .CK(clk), .Q(\AES_ENC/sa12 [3]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_3_  ( .D(\AES_ENC/N97 ), .CK(clk), .Q(\AES_ENC/sa32 [3]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_3_  ( .D(\AES_ENC/N113 ), .CK(clk), .Q(\AES_ENC/sa22 [3]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_4_  ( .D(\AES_ENC/N146 ), .CK(clk), .Q(\AES_ENC/sa02 [4]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_2_  ( .D(\AES_ENC/N128 ), .CK(clk), .Q(\AES_ENC/sa12 [2]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_2_  ( .D(\AES_ENC/N96 ), .CK(clk), .Q(\AES_ENC/sa32 [2]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_2_  ( .D(\AES_ENC/N112 ), .CK(clk), .Q(\AES_ENC/sa22 [2]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_3_  ( .D(\AES_ENC/N145 ), .CK(clk), .Q(\AES_ENC/sa02 [3]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_1_  ( .D(\AES_ENC/N127 ), .CK(clk), .Q(\AES_ENC/sa12 [1]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_1_  ( .D(\AES_ENC/N95 ), .CK(clk), .Q(\AES_ENC/sa32 [1]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_1_  ( .D(\AES_ENC/N111 ), .CK(clk), .Q(\AES_ENC/sa22 [1]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_2_  ( .D(\AES_ENC/N144 ), .CK(clk), .Q(\AES_ENC/sa02 [2]), .QN() );
DFF_X2 \AES_ENC/sa22_reg_0_  ( .D(\AES_ENC/N110 ), .CK(clk), .Q(\AES_ENC/sa22 [0]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_1_  ( .D(\AES_ENC/N143 ), .CK(clk), .Q(\AES_ENC/sa02 [1]), .QN() );
DFF_X2 \AES_ENC/sa02_reg_0_  ( .D(\AES_ENC/N142 ), .CK(clk), .Q(\AES_ENC/sa02 [0]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_0_  ( .D(\AES_ENC/N62 ), .CK(clk), .Q(\AES_ENC/sa13 [0]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_1_  ( .D(\AES_ENC/N63 ), .CK(clk), .Q(\AES_ENC/sa13 [1]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_3_  ( .D(\AES_ENC/N65 ), .CK(clk), .Q(\AES_ENC/sa13 [3]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_4_  ( .D(\AES_ENC/N66 ), .CK(clk), .Q(\AES_ENC/sa13 [4]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_7_  ( .D(\AES_ENC/N37 ), .CK(clk), .Q(\AES_ENC/sa33 [7]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_7_  ( .D(\AES_ENC/N165 ), .CK(clk), .Q(\AES_ENC/sa31 [7]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_0_  ( .D(\AES_ENC/N46 ), .CK(clk), .Q(\AES_ENC/sa23 [0]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_1_  ( .D(\AES_ENC/N47 ), .CK(clk), .Q(\AES_ENC/sa23 [1]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_3_  ( .D(\AES_ENC/N49 ), .CK(clk), .Q(\AES_ENC/sa23 [3]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_4_  ( .D(\AES_ENC/N50 ), .CK(clk), .Q(\AES_ENC/sa23 [4]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_7_  ( .D(\AES_ENC/N69 ), .CK(clk), .Q(\AES_ENC/sa13 [7]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_6_  ( .D(\AES_ENC/N68 ), .CK(clk), .Q(\AES_ENC/sa13 [6]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_6_  ( .D(\AES_ENC/N36 ), .CK(clk), .Q(\AES_ENC/sa33 [6]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_6_  ( .D(\AES_ENC/N52 ), .CK(clk), .Q(\AES_ENC/sa23 [6]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_5_  ( .D(\AES_ENC/N67 ), .CK(clk), .Q(\AES_ENC/sa13 [5]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_5_  ( .D(\AES_ENC/N35 ), .CK(clk), .Q(\AES_ENC/sa33 [5]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_5_  ( .D(\AES_ENC/N51 ), .CK(clk), .Q(\AES_ENC/sa23 [5]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_6_  ( .D(\AES_ENC/N84 ), .CK(clk), .Q(\AES_ENC/sa03 [6]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_4_  ( .D(\AES_ENC/N34 ), .CK(clk), .Q(\AES_ENC/sa33 [4]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_5_  ( .D(\AES_ENC/N83 ), .CK(clk), .Q(\AES_ENC/sa03 [5]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_3_  ( .D(\AES_ENC/N33 ), .CK(clk), .Q(\AES_ENC/sa33 [3]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_4_  ( .D(\AES_ENC/N82 ), .CK(clk), .Q(\AES_ENC/sa03 [4]), .QN() );
DFF_X2 \AES_ENC/sa13_reg_2_  ( .D(\AES_ENC/N64 ), .CK(clk), .Q(\AES_ENC/sa13 [2]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_2_  ( .D(\AES_ENC/N32 ), .CK(clk), .Q(\AES_ENC/sa33 [2]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_2_  ( .D(\AES_ENC/N48 ), .CK(clk), .Q(\AES_ENC/sa23 [2]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_3_  ( .D(\AES_ENC/N81 ), .CK(clk), .Q(\AES_ENC/sa03 [3]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_1_  ( .D(\AES_ENC/N31 ), .CK(clk), .Q(\AES_ENC/sa33 [1]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_2_  ( .D(\AES_ENC/N80 ), .CK(clk), .Q(\AES_ENC/sa03 [2]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_1_  ( .D(\AES_ENC/N79 ), .CK(clk), .Q(\AES_ENC/sa03 [1]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_7_  ( .D(\AES_ENC/N85 ), .CK(clk), .Q(\AES_ENC/sa03 [7]), .QN() );
DFF_X2 \AES_ENC/sa03_reg_0_  ( .D(\AES_ENC/N78 ), .CK(clk), .Q(\AES_ENC/sa03 [0]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_0_  ( .D(\AES_ENC/N174 ), .CK(clk), .Q(\AES_ENC/sa21 [0]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_1_  ( .D(\AES_ENC/N175 ), .CK(clk), .Q(\AES_ENC/sa21 [1]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_3_  ( .D(\AES_ENC/N177 ), .CK(clk), .Q(\AES_ENC/sa21 [3]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_4_  ( .D(\AES_ENC/N178 ), .CK(clk), .Q(\AES_ENC/sa21 [4]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_7_  ( .D(\AES_ENC/N197 ), .CK(clk), .Q(\AES_ENC/sa11 [7]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_7_  ( .D(\AES_ENC/N181 ), .CK(clk), .Q(\AES_ENC/sa21 [7]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_0_  ( .D(\AES_ENC/N206 ), .CK(clk), .Q(\AES_ENC/sa01 [0]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_1_  ( .D(\AES_ENC/N207 ), .CK(clk), .Q(\AES_ENC/sa01 [1]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_3_  ( .D(\AES_ENC/N209 ), .CK(clk), .Q(\AES_ENC/sa01 [3]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_4_  ( .D(\AES_ENC/N210 ), .CK(clk), .Q(\AES_ENC/sa01 [4]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_6_  ( .D(\AES_ENC/N196 ), .CK(clk), .Q(\AES_ENC/sa11 [6]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_6_  ( .D(\AES_ENC/N164 ), .CK(clk), .Q(\AES_ENC/sa31 [6]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_6_  ( .D(\AES_ENC/N180 ), .CK(clk), .Q(\AES_ENC/sa21 [6]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_5_  ( .D(\AES_ENC/N195 ), .CK(clk), .Q(\AES_ENC/sa11 [5]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_5_  ( .D(\AES_ENC/N163 ), .CK(clk), .Q(\AES_ENC/sa31 [5]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_5_  ( .D(\AES_ENC/N179 ), .CK(clk), .Q(\AES_ENC/sa21 [5]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_6_  ( .D(\AES_ENC/N212 ), .CK(clk), .Q(\AES_ENC/sa01 [6]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_4_  ( .D(\AES_ENC/N194 ), .CK(clk), .Q(\AES_ENC/sa11 [4]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_4_  ( .D(\AES_ENC/N162 ), .CK(clk), .Q(\AES_ENC/sa31 [4]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_5_  ( .D(\AES_ENC/N211 ), .CK(clk), .Q(\AES_ENC/sa01 [5]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_3_  ( .D(\AES_ENC/N193 ), .CK(clk), .Q(\AES_ENC/sa11 [3]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_3_  ( .D(\AES_ENC/N161 ), .CK(clk), .Q(\AES_ENC/sa31 [3]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_2_  ( .D(\AES_ENC/N192 ), .CK(clk), .Q(\AES_ENC/sa11 [2]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_2_  ( .D(\AES_ENC/N160 ), .CK(clk), .Q(\AES_ENC/sa31 [2]), .QN() );
DFF_X2 \AES_ENC/sa21_reg_2_  ( .D(\AES_ENC/N176 ), .CK(clk), .Q(\AES_ENC/sa21 [2]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_1_  ( .D(\AES_ENC/N191 ), .CK(clk), .Q(\AES_ENC/sa11 [1]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_1_  ( .D(\AES_ENC/N159 ), .CK(clk), .Q(\AES_ENC/sa31 [1]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_2_  ( .D(\AES_ENC/N208 ), .CK(clk), .Q(\AES_ENC/sa01 [2]), .QN() );
DFF_X2 \AES_ENC/sa01_reg_7_  ( .D(\AES_ENC/N213 ), .CK(clk), .Q(\AES_ENC/sa01 [7]), .QN() );
DFF_X2 \AES_ENC/sa23_reg_7_  ( .D(\AES_ENC/N53 ), .CK(clk), .Q(\AES_ENC/sa23 [7]), .QN() );
DFF_X2 \AES_ENC/sa10_reg_0_  ( .D(\AES_ENC/N254 ), .CK(clk), .Q(\AES_ENC/sa10 [0]), .QN() );
DFF_X2 \AES_ENC/sa11_reg_0_  ( .D(\AES_ENC/N190 ), .CK(clk), .Q(\AES_ENC/sa11 [0]), .QN() );
DFF_X2 \AES_ENC/sa12_reg_0_  ( .D(\AES_ENC/N126 ), .CK(clk), .Q(\AES_ENC/sa12 [0]), .QN() );
DFF_X2 \AES_ENC/sa20_reg_7_  ( .D(\AES_ENC/N245 ), .CK(clk), .Q(\AES_ENC/sa20 [7]), .QN() );
DFF_X2 \AES_ENC/sa33_reg_0_  ( .D(\AES_ENC/N30 ), .CK(clk), .Q(\AES_ENC/sa33 [0]), .QN() );
DFF_X2 \AES_ENC/sa32_reg_0_  ( .D(\AES_ENC/N94 ), .CK(clk), .Q(\AES_ENC/sa32 [0]), .QN() );
DFF_X2 \AES_ENC/sa31_reg_0_  ( .D(\AES_ENC/N158 ), .CK(clk), .Q(\AES_ENC/sa31 [0]), .QN() );
DFF_X2 \AES_ENC/sa30_reg_0_  ( .D(\AES_ENC/N222 ), .CK(clk), .Q(\AES_ENC/sa30 [0]), .QN() );
DFF_X2 \AES_ENC/sa00_reg_0_  ( .D(\AES_ENC/N270 ), .CK(clk), .Q(\AES_ENC/sa00 [0]), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_0_  ( .D(\AES_ENC/n661 ), .CK(clk), .Q(\AES_ENC/text_in_r[0] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_1_  ( .D(\AES_ENC/n662 ), .CK(clk), .Q(\AES_ENC/text_in_r[1] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_2_  ( .D(\AES_ENC/n663 ), .CK(clk), .Q(\AES_ENC/text_in_r[2] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_3_  ( .D(\AES_ENC/n664 ), .CK(clk), .Q(\AES_ENC/text_in_r[3] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_4_  ( .D(\AES_ENC/n665 ), .CK(clk), .Q(\AES_ENC/text_in_r[4] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_5_  ( .D(\AES_ENC/n666 ), .CK(clk), .Q(\AES_ENC/text_in_r[5] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_6_  ( .D(\AES_ENC/n667 ), .CK(clk), .Q(\AES_ENC/text_in_r[6] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_7_  ( .D(\AES_ENC/n668 ), .CK(clk), .Q(\AES_ENC/text_in_r[7] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_8_  ( .D(\AES_ENC/n669 ), .CK(clk), .Q(\AES_ENC/text_in_r[8] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_9_  ( .D(\AES_ENC/n670 ), .CK(clk), .Q(\AES_ENC/text_in_r[9] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_10_  ( .D(\AES_ENC/n671 ), .CK(clk), .Q(\AES_ENC/text_in_r[10] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_11_  ( .D(\AES_ENC/n672 ), .CK(clk), .Q(\AES_ENC/text_in_r[11] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_12_  ( .D(\AES_ENC/n673 ), .CK(clk), .Q(\AES_ENC/text_in_r[12] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_13_  ( .D(\AES_ENC/n674 ), .CK(clk), .Q(\AES_ENC/text_in_r[13] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_14_  ( .D(\AES_ENC/n675 ), .CK(clk), .Q(\AES_ENC/text_in_r[14] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_15_  ( .D(\AES_ENC/n676 ), .CK(clk), .Q(\AES_ENC/text_in_r[15] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_16_  ( .D(\AES_ENC/n677 ), .CK(clk), .Q(\AES_ENC/text_in_r[16] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_17_  ( .D(\AES_ENC/n678 ), .CK(clk), .Q(\AES_ENC/text_in_r[17] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_18_  ( .D(\AES_ENC/n679 ), .CK(clk), .Q(\AES_ENC/text_in_r[18] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_19_  ( .D(\AES_ENC/n680 ), .CK(clk), .Q(\AES_ENC/text_in_r[19] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_20_  ( .D(\AES_ENC/n681 ), .CK(clk), .Q(\AES_ENC/text_in_r[20] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_21_  ( .D(\AES_ENC/n682 ), .CK(clk), .Q(\AES_ENC/text_in_r[21] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_22_  ( .D(\AES_ENC/n683 ), .CK(clk), .Q(\AES_ENC/text_in_r[22] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_23_  ( .D(\AES_ENC/n684 ), .CK(clk), .Q(\AES_ENC/text_in_r[23] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_24_  ( .D(\AES_ENC/n685 ), .CK(clk), .Q(\AES_ENC/text_in_r[24] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_25_  ( .D(\AES_ENC/n686 ), .CK(clk), .Q(\AES_ENC/text_in_r[25] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_26_  ( .D(\AES_ENC/n687 ), .CK(clk), .Q(\AES_ENC/text_in_r[26] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_27_  ( .D(\AES_ENC/n688 ), .CK(clk), .Q(\AES_ENC/text_in_r[27] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_28_  ( .D(\AES_ENC/n689 ), .CK(clk), .Q(\AES_ENC/text_in_r[28] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_29_  ( .D(\AES_ENC/n690 ), .CK(clk), .Q(\AES_ENC/text_in_r[29] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_30_  ( .D(\AES_ENC/n691 ), .CK(clk), .Q(\AES_ENC/text_in_r[30] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_31_  ( .D(\AES_ENC/n692 ), .CK(clk), .Q(\AES_ENC/text_in_r[31] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_32_  ( .D(\AES_ENC/n693 ), .CK(clk), .Q(\AES_ENC/text_in_r[32] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_33_  ( .D(\AES_ENC/n694 ), .CK(clk), .Q(\AES_ENC/text_in_r[33] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_34_  ( .D(\AES_ENC/n695 ), .CK(clk), .Q(\AES_ENC/text_in_r[34] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_35_  ( .D(\AES_ENC/n696 ), .CK(clk), .Q(\AES_ENC/text_in_r[35] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_36_  ( .D(\AES_ENC/n697 ), .CK(clk), .Q(\AES_ENC/text_in_r[36] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_37_  ( .D(\AES_ENC/n698 ), .CK(clk), .Q(\AES_ENC/text_in_r[37] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_38_  ( .D(\AES_ENC/n699 ), .CK(clk), .Q(\AES_ENC/text_in_r[38] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_39_  ( .D(\AES_ENC/n700 ), .CK(clk), .Q(\AES_ENC/text_in_r[39] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_40_  ( .D(\AES_ENC/n701 ), .CK(clk), .Q(\AES_ENC/text_in_r[40] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_41_  ( .D(\AES_ENC/n702 ), .CK(clk), .Q(\AES_ENC/text_in_r[41] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_42_  ( .D(\AES_ENC/n703 ), .CK(clk), .Q(\AES_ENC/text_in_r[42] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_43_  ( .D(\AES_ENC/n704 ), .CK(clk), .Q(\AES_ENC/text_in_r[43] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_44_  ( .D(\AES_ENC/n705 ), .CK(clk), .Q(\AES_ENC/text_in_r[44] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_45_  ( .D(\AES_ENC/n706 ), .CK(clk), .Q(\AES_ENC/text_in_r[45] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_46_  ( .D(\AES_ENC/n707 ), .CK(clk), .Q(\AES_ENC/text_in_r[46] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_47_  ( .D(\AES_ENC/n708 ), .CK(clk), .Q(\AES_ENC/text_in_r[47] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_48_  ( .D(\AES_ENC/n709 ), .CK(clk), .Q(\AES_ENC/text_in_r[48] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_49_  ( .D(\AES_ENC/n710 ), .CK(clk), .Q(\AES_ENC/text_in_r[49] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_50_  ( .D(\AES_ENC/n711 ), .CK(clk), .Q(\AES_ENC/text_in_r[50] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_51_  ( .D(\AES_ENC/n712 ), .CK(clk), .Q(\AES_ENC/text_in_r[51] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_52_  ( .D(\AES_ENC/n713 ), .CK(clk), .Q(\AES_ENC/text_in_r[52] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_53_  ( .D(\AES_ENC/n714 ), .CK(clk), .Q(\AES_ENC/text_in_r[53] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_54_  ( .D(\AES_ENC/n715 ), .CK(clk), .Q(\AES_ENC/text_in_r[54] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_55_  ( .D(\AES_ENC/n716 ), .CK(clk), .Q(\AES_ENC/text_in_r[55] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_56_  ( .D(\AES_ENC/n717 ), .CK(clk), .Q(\AES_ENC/text_in_r[56] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_57_  ( .D(\AES_ENC/n718 ), .CK(clk), .Q(\AES_ENC/text_in_r[57] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_58_  ( .D(\AES_ENC/n719 ), .CK(clk), .Q(\AES_ENC/text_in_r[58] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_59_  ( .D(\AES_ENC/n720 ), .CK(clk), .Q(\AES_ENC/text_in_r[59] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_60_  ( .D(\AES_ENC/n721 ), .CK(clk), .Q(\AES_ENC/text_in_r[60] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_61_  ( .D(\AES_ENC/n722 ), .CK(clk), .Q(\AES_ENC/text_in_r[61] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_62_  ( .D(\AES_ENC/n723 ), .CK(clk), .Q(\AES_ENC/text_in_r[62] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_63_  ( .D(\AES_ENC/n724 ), .CK(clk), .Q(\AES_ENC/text_in_r[63] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_64_  ( .D(\AES_ENC/n725 ), .CK(clk), .Q(\AES_ENC/text_in_r[64] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_65_  ( .D(\AES_ENC/n726 ), .CK(clk), .Q(\AES_ENC/text_in_r[65] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_66_  ( .D(\AES_ENC/n727 ), .CK(clk), .Q(\AES_ENC/text_in_r[66] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_67_  ( .D(\AES_ENC/n728 ), .CK(clk), .Q(\AES_ENC/text_in_r[67] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_68_  ( .D(\AES_ENC/n729 ), .CK(clk), .Q(\AES_ENC/text_in_r[68] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_69_  ( .D(\AES_ENC/n730 ), .CK(clk), .Q(\AES_ENC/text_in_r[69] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_70_  ( .D(\AES_ENC/n731 ), .CK(clk), .Q(\AES_ENC/text_in_r[70] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_71_  ( .D(\AES_ENC/n732 ), .CK(clk), .Q(\AES_ENC/text_in_r[71] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_72_  ( .D(\AES_ENC/n733 ), .CK(clk), .Q(\AES_ENC/text_in_r[72] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_73_  ( .D(\AES_ENC/n734 ), .CK(clk), .Q(\AES_ENC/text_in_r[73] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_74_  ( .D(\AES_ENC/n735 ), .CK(clk), .Q(\AES_ENC/text_in_r[74] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_75_  ( .D(\AES_ENC/n736 ), .CK(clk), .Q(\AES_ENC/text_in_r[75] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_76_  ( .D(\AES_ENC/n737 ), .CK(clk), .Q(\AES_ENC/text_in_r[76] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_77_  ( .D(\AES_ENC/n738 ), .CK(clk), .Q(\AES_ENC/text_in_r[77] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_78_  ( .D(\AES_ENC/n739 ), .CK(clk), .Q(\AES_ENC/text_in_r[78] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_79_  ( .D(\AES_ENC/n740 ), .CK(clk), .Q(\AES_ENC/text_in_r[79] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_80_  ( .D(\AES_ENC/n741 ), .CK(clk), .Q(\AES_ENC/text_in_r[80] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_81_  ( .D(\AES_ENC/n742 ), .CK(clk), .Q(\AES_ENC/text_in_r[81] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_82_  ( .D(\AES_ENC/n743 ), .CK(clk), .Q(\AES_ENC/text_in_r[82] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_83_  ( .D(\AES_ENC/n744 ), .CK(clk), .Q(\AES_ENC/text_in_r[83] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_84_  ( .D(\AES_ENC/n745 ), .CK(clk), .Q(\AES_ENC/text_in_r[84] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_85_  ( .D(\AES_ENC/n746 ), .CK(clk), .Q(\AES_ENC/text_in_r[85] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_86_  ( .D(\AES_ENC/n747 ), .CK(clk), .Q(\AES_ENC/text_in_r[86] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_87_  ( .D(\AES_ENC/n748 ), .CK(clk), .Q(\AES_ENC/text_in_r[87] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_88_  ( .D(\AES_ENC/n749 ), .CK(clk), .Q(\AES_ENC/text_in_r[88] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_89_  ( .D(\AES_ENC/n750 ), .CK(clk), .Q(\AES_ENC/text_in_r[89] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_90_  ( .D(\AES_ENC/n751 ), .CK(clk), .Q(\AES_ENC/text_in_r[90] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_91_  ( .D(\AES_ENC/n752 ), .CK(clk), .Q(\AES_ENC/text_in_r[91] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_92_  ( .D(\AES_ENC/n753 ), .CK(clk), .Q(\AES_ENC/text_in_r[92] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_93_  ( .D(\AES_ENC/n754 ), .CK(clk), .Q(\AES_ENC/text_in_r[93] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_94_  ( .D(\AES_ENC/n755 ), .CK(clk), .Q(\AES_ENC/text_in_r[94] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_95_  ( .D(\AES_ENC/n756 ), .CK(clk), .Q(\AES_ENC/text_in_r[95] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_96_  ( .D(\AES_ENC/n757 ), .CK(clk), .Q(\AES_ENC/text_in_r[96] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_97_  ( .D(\AES_ENC/n758 ), .CK(clk), .Q(\AES_ENC/text_in_r[97] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_98_  ( .D(\AES_ENC/n759 ), .CK(clk), .Q(\AES_ENC/text_in_r[98] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_99_  ( .D(\AES_ENC/n760 ), .CK(clk), .Q(\AES_ENC/text_in_r[99] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_100_  ( .D(\AES_ENC/n761 ), .CK(clk), .Q(\AES_ENC/text_in_r[100] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_101_  ( .D(\AES_ENC/n762 ), .CK(clk), .Q(\AES_ENC/text_in_r[101] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_102_  ( .D(\AES_ENC/n763 ), .CK(clk), .Q(\AES_ENC/text_in_r[102] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_103_  ( .D(\AES_ENC/n764 ), .CK(clk), .Q(\AES_ENC/text_in_r[103] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_104_  ( .D(\AES_ENC/n765 ), .CK(clk), .Q(\AES_ENC/text_in_r[104] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_105_  ( .D(\AES_ENC/n766 ), .CK(clk), .Q(\AES_ENC/text_in_r[105] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_106_  ( .D(\AES_ENC/n767 ), .CK(clk), .Q(\AES_ENC/text_in_r[106] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_107_  ( .D(\AES_ENC/n768 ), .CK(clk), .Q(\AES_ENC/text_in_r[107] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_108_  ( .D(\AES_ENC/n769 ), .CK(clk), .Q(\AES_ENC/text_in_r[108] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_109_  ( .D(\AES_ENC/n770 ), .CK(clk), .Q(\AES_ENC/text_in_r[109] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_110_  ( .D(\AES_ENC/n771 ), .CK(clk), .Q(\AES_ENC/text_in_r[110] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_111_  ( .D(\AES_ENC/n772 ), .CK(clk), .Q(\AES_ENC/text_in_r[111] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_112_  ( .D(\AES_ENC/n773 ), .CK(clk), .Q(\AES_ENC/text_in_r[112] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_113_  ( .D(\AES_ENC/n774 ), .CK(clk), .Q(\AES_ENC/text_in_r[113] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_114_  ( .D(\AES_ENC/n775 ), .CK(clk), .Q(\AES_ENC/text_in_r[114] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_115_  ( .D(\AES_ENC/n776 ), .CK(clk), .Q(\AES_ENC/text_in_r[115] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_116_  ( .D(\AES_ENC/n777 ), .CK(clk), .Q(\AES_ENC/text_in_r[116] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_117_  ( .D(\AES_ENC/n778 ), .CK(clk), .Q(\AES_ENC/text_in_r[117] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_118_  ( .D(\AES_ENC/n779 ), .CK(clk), .Q(\AES_ENC/text_in_r[118] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_119_  ( .D(\AES_ENC/n780 ), .CK(clk), .Q(\AES_ENC/text_in_r[119] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_120_  ( .D(\AES_ENC/n781 ), .CK(clk), .Q(\AES_ENC/text_in_r[120] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_121_  ( .D(\AES_ENC/n782 ), .CK(clk), .Q(\AES_ENC/text_in_r[121] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_122_  ( .D(\AES_ENC/n783 ), .CK(clk), .Q(\AES_ENC/text_in_r[122] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_123_  ( .D(\AES_ENC/n784 ), .CK(clk), .Q(\AES_ENC/text_in_r[123] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_124_  ( .D(\AES_ENC/n785 ), .CK(clk), .Q(\AES_ENC/text_in_r[124] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_125_  ( .D(\AES_ENC/n786 ), .CK(clk), .Q(\AES_ENC/text_in_r[125] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_126_  ( .D(\AES_ENC/n787 ), .CK(clk), .Q(\AES_ENC/text_in_r[126] ), .QN() );
DFF_X2 \AES_ENC/text_in_r_reg_127_  ( .D(\AES_ENC/n788 ), .CK(clk), .Q(\AES_ENC/text_in_r[127] ), .QN() );
DFF_X2 \AES_ENC/done_reg  ( .D(\AES_ENC/N19 ), .CK(clk), .Q(aes_done), .QN());
XOR2_X2 \AES_ENC/U1612  ( .A(\AES_ENC/sa22_sub[7] ), .B(\AES_ENC/sa33_sub[7] ), .Z(\AES_ENC/n1167 ) );
XOR2_X2 \AES_ENC/U1611  ( .A(\AES_ENC/sa00_sub[6] ), .B(\AES_ENC/sa11_sub[6] ), .Z(\AES_ENC/n1169 ) );
XOR2_X2 \AES_ENC/U1610  ( .A(\AES_ENC/n800 ), .B(\AES_ENC/n799 ), .Z(\AES_ENC/sa00_next [7]) );
XOR2_X2 \AES_ENC/U1609  ( .A(\AES_ENC/n1167 ), .B(\AES_ENC/n1169 ), .Z(\AES_ENC/n799 ) );
XOR2_X2 \AES_ENC/U1608  ( .A(\AES_ENC/w0[31] ), .B(\AES_ENC/sa11_sub[7] ),.Z(\AES_ENC/n800 ) );
XOR2_X2 \AES_ENC/U1607  ( .A(\AES_ENC/sa00_sub[5] ), .B(\AES_ENC/sa11_sub[5] ), .Z(\AES_ENC/n1170 ) );
XOR2_X2 \AES_ENC/U1606  ( .A(\AES_ENC/sa22_sub[6] ), .B(\AES_ENC/sa33_sub[6] ), .Z(\AES_ENC/n1160 ) );
XOR2_X2 \AES_ENC/U1605  ( .A(\AES_ENC/n802 ), .B(\AES_ENC/n801 ), .Z(\AES_ENC/sa00_next [6]) );
XOR2_X2 \AES_ENC/U1604  ( .A(\AES_ENC/n1170 ), .B(\AES_ENC/n1160 ), .Z(\AES_ENC/n801 ) );
XOR2_X2 \AES_ENC/U1603  ( .A(\AES_ENC/w0[30] ), .B(\AES_ENC/sa11_sub[6] ),.Z(\AES_ENC/n802 ) );
XOR2_X2 \AES_ENC/U1602  ( .A(\AES_ENC/sa00_sub[4] ), .B(\AES_ENC/sa11_sub[4] ), .Z(\AES_ENC/n1171 ) );
XOR2_X2 \AES_ENC/U1601  ( .A(\AES_ENC/sa22_sub[5] ), .B(\AES_ENC/sa33_sub[5] ), .Z(\AES_ENC/n1161 ) );
XOR2_X2 \AES_ENC/U1600  ( .A(\AES_ENC/n804 ), .B(\AES_ENC/n803 ), .Z(\AES_ENC/sa00_next [5]) );
XOR2_X2 \AES_ENC/U1599  ( .A(\AES_ENC/n1171 ), .B(\AES_ENC/n1161 ), .Z(\AES_ENC/n803 ) );
XOR2_X2 \AES_ENC/U1598  ( .A(\AES_ENC/w0[29] ), .B(\AES_ENC/sa11_sub[5] ),.Z(\AES_ENC/n804 ) );
XOR2_X2 \AES_ENC/U1597  ( .A(\AES_ENC/sa00_sub[7] ), .B(\AES_ENC/sa11_sub[7] ), .Z(\AES_ENC/n1168 ) );
XOR2_X2 \AES_ENC/U1596  ( .A(\AES_ENC/sa00_sub[3] ), .B(\AES_ENC/sa11_sub[3] ), .Z(\AES_ENC/n1172 ) );
XOR2_X2 \AES_ENC/U1595  ( .A(\AES_ENC/sa22_sub[4] ), .B(\AES_ENC/sa33_sub[4] ), .Z(\AES_ENC/n1162 ) );
XOR2_X2 \AES_ENC/U1594  ( .A(\AES_ENC/n806 ), .B(\AES_ENC/n805 ), .Z(\AES_ENC/sa00_next [4]) );
XOR2_X2 \AES_ENC/U1593  ( .A(\AES_ENC/n1162 ), .B(\AES_ENC/n807 ), .Z(\AES_ENC/n805 ) );
XOR2_X2 \AES_ENC/U1592  ( .A(\AES_ENC/n1168 ), .B(\AES_ENC/n1172 ), .Z(\AES_ENC/n806 ) );
XOR2_X2 \AES_ENC/U1591  ( .A(\AES_ENC/w0[28] ), .B(\AES_ENC/sa11_sub[4] ),.Z(\AES_ENC/n807 ) );
XOR2_X2 \AES_ENC/U1590  ( .A(\AES_ENC/sa00_sub[2] ), .B(\AES_ENC/sa11_sub[2] ), .Z(\AES_ENC/n1173 ) );
XOR2_X2 \AES_ENC/U1589  ( .A(\AES_ENC/sa22_sub[3] ), .B(\AES_ENC/sa33_sub[3] ), .Z(\AES_ENC/n1163 ) );
XOR2_X2 \AES_ENC/U1588  ( .A(\AES_ENC/n809 ), .B(\AES_ENC/n808 ), .Z(\AES_ENC/sa00_next [3]) );
XOR2_X2 \AES_ENC/U1587  ( .A(\AES_ENC/n1163 ), .B(\AES_ENC/n810 ), .Z(\AES_ENC/n808 ) );
XOR2_X2 \AES_ENC/U1586  ( .A(\AES_ENC/n1168 ), .B(\AES_ENC/n1173 ), .Z(\AES_ENC/n809 ) );
XOR2_X2 \AES_ENC/U1585  ( .A(\AES_ENC/w0[27] ), .B(\AES_ENC/sa11_sub[3] ),.Z(\AES_ENC/n810 ) );
XOR2_X2 \AES_ENC/U1584  ( .A(\AES_ENC/sa00_sub[1] ), .B(\AES_ENC/sa11_sub[1] ), .Z(\AES_ENC/n1174 ) );
XOR2_X2 \AES_ENC/U1583  ( .A(\AES_ENC/sa22_sub[2] ), .B(\AES_ENC/sa33_sub[2] ), .Z(\AES_ENC/n1164 ) );
XOR2_X2 \AES_ENC/U1582  ( .A(\AES_ENC/n812 ), .B(\AES_ENC/n811 ), .Z(\AES_ENC/sa00_next [2]) );
XOR2_X2 \AES_ENC/U1581  ( .A(\AES_ENC/n1174 ), .B(\AES_ENC/n1164 ), .Z(\AES_ENC/n811 ) );
XOR2_X2 \AES_ENC/U1580  ( .A(\AES_ENC/w0[26] ), .B(\AES_ENC/sa11_sub[2] ),.Z(\AES_ENC/n812 ) );
XOR2_X2 \AES_ENC/U1579  ( .A(\AES_ENC/sa00_sub[0] ), .B(\AES_ENC/sa11_sub[0] ), .Z(\AES_ENC/n1175 ) );
XOR2_X2 \AES_ENC/U1578  ( .A(\AES_ENC/sa22_sub[1] ), .B(\AES_ENC/sa33_sub[1] ), .Z(\AES_ENC/n1165 ) );
XOR2_X2 \AES_ENC/U1577  ( .A(\AES_ENC/n814 ), .B(\AES_ENC/n813 ), .Z(\AES_ENC/sa00_next [1]) );
XOR2_X2 \AES_ENC/U1576  ( .A(\AES_ENC/n1165 ), .B(\AES_ENC/n815 ), .Z(\AES_ENC/n813 ) );
XOR2_X2 \AES_ENC/U1575  ( .A(\AES_ENC/n1168 ), .B(\AES_ENC/n1175 ), .Z(\AES_ENC/n814 ) );
XOR2_X2 \AES_ENC/U1574  ( .A(\AES_ENC/w0[25] ), .B(\AES_ENC/sa11_sub[1] ),.Z(\AES_ENC/n815 ) );
XOR2_X2 \AES_ENC/U1573  ( .A(\AES_ENC/sa22_sub[0] ), .B(\AES_ENC/sa33_sub[0] ), .Z(\AES_ENC/n1166 ) );
XOR2_X2 \AES_ENC/U1572  ( .A(\AES_ENC/n817 ), .B(\AES_ENC/n816 ), .Z(\AES_ENC/sa00_next [0]) );
XOR2_X2 \AES_ENC/U1571  ( .A(\AES_ENC/n1168 ), .B(\AES_ENC/n1166 ), .Z(\AES_ENC/n816 ) );
XOR2_X2 \AES_ENC/U1570  ( .A(\AES_ENC/w0[24] ), .B(\AES_ENC/sa11_sub[0] ),.Z(\AES_ENC/n817 ) );
XOR2_X2 \AES_ENC/U1569  ( .A(\AES_ENC/n819 ), .B(\AES_ENC/n818 ), .Z(\AES_ENC/sa10_next [7]) );
XOR2_X2 \AES_ENC/U1568  ( .A(\AES_ENC/n1167 ), .B(\AES_ENC/n820 ), .Z(\AES_ENC/n818 ) );
XOR2_X2 \AES_ENC/U1567  ( .A(\AES_ENC/sa11_sub[6] ), .B(\AES_ENC/sa22_sub[6] ), .Z(\AES_ENC/n819 ) );
XOR2_X2 \AES_ENC/U1566  ( .A(\AES_ENC/w0[23] ), .B(\AES_ENC/sa00_sub[7] ),.Z(\AES_ENC/n820 ) );
XOR2_X2 \AES_ENC/U1565  ( .A(\AES_ENC/n822 ), .B(\AES_ENC/n821 ), .Z(\AES_ENC/sa10_next [6]) );
XOR2_X2 \AES_ENC/U1564  ( .A(\AES_ENC/n1160 ), .B(\AES_ENC/n823 ), .Z(\AES_ENC/n821 ) );
XOR2_X2 \AES_ENC/U1563  ( .A(\AES_ENC/sa11_sub[5] ), .B(\AES_ENC/sa22_sub[5] ), .Z(\AES_ENC/n822 ) );
XOR2_X2 \AES_ENC/U1562  ( .A(\AES_ENC/w0[22] ), .B(\AES_ENC/sa00_sub[6] ),.Z(\AES_ENC/n823 ) );
XOR2_X2 \AES_ENC/U1561  ( .A(\AES_ENC/n825 ), .B(\AES_ENC/n824 ), .Z(\AES_ENC/sa10_next [5]) );
XOR2_X2 \AES_ENC/U1560  ( .A(\AES_ENC/n1161 ), .B(\AES_ENC/n826 ), .Z(\AES_ENC/n824 ) );
XOR2_X2 \AES_ENC/U1559  ( .A(\AES_ENC/sa11_sub[4] ), .B(\AES_ENC/sa22_sub[4] ), .Z(\AES_ENC/n825 ) );
XOR2_X2 \AES_ENC/U1558  ( .A(\AES_ENC/w0[21] ), .B(\AES_ENC/sa00_sub[5] ),.Z(\AES_ENC/n826 ) );
XOR2_X2 \AES_ENC/U1557  ( .A(\AES_ENC/sa11_sub[7] ), .B(\AES_ENC/sa22_sub[7] ), .Z(\AES_ENC/n1159 ) );
XOR2_X2 \AES_ENC/U1556  ( .A(\AES_ENC/n828 ), .B(\AES_ENC/n827 ), .Z(\AES_ENC/sa10_next [4]) );
XOR2_X2 \AES_ENC/U1555  ( .A(\AES_ENC/n830 ), .B(\AES_ENC/n829 ), .Z(\AES_ENC/n827 ) );
XOR2_X2 \AES_ENC/U1554  ( .A(\AES_ENC/n1159 ), .B(\AES_ENC/n1162 ), .Z(\AES_ENC/n828 ) );
XOR2_X2 \AES_ENC/U1553  ( .A(\AES_ENC/sa11_sub[3] ), .B(\AES_ENC/sa22_sub[3] ), .Z(\AES_ENC/n829 ) );
XOR2_X2 \AES_ENC/U1552  ( .A(\AES_ENC/w0[20] ), .B(\AES_ENC/sa00_sub[4] ),.Z(\AES_ENC/n830 ) );
XOR2_X2 \AES_ENC/U1551  ( .A(\AES_ENC/n832 ), .B(\AES_ENC/n831 ), .Z(\AES_ENC/sa10_next [3]) );
XOR2_X2 \AES_ENC/U1550  ( .A(\AES_ENC/n834 ), .B(\AES_ENC/n833 ), .Z(\AES_ENC/n831 ) );
XOR2_X2 \AES_ENC/U1549  ( .A(\AES_ENC/n1159 ), .B(\AES_ENC/n1163 ), .Z(\AES_ENC/n832 ) );
XOR2_X2 \AES_ENC/U1548  ( .A(\AES_ENC/sa11_sub[2] ), .B(\AES_ENC/sa22_sub[2] ), .Z(\AES_ENC/n833 ) );
XOR2_X2 \AES_ENC/U1547  ( .A(\AES_ENC/w0[19] ), .B(\AES_ENC/sa00_sub[3] ),.Z(\AES_ENC/n834 ) );
XOR2_X2 \AES_ENC/U1546  ( .A(\AES_ENC/n836 ), .B(\AES_ENC/n835 ), .Z(\AES_ENC/sa10_next [2]) );
XOR2_X2 \AES_ENC/U1545  ( .A(\AES_ENC/n1164 ), .B(\AES_ENC/n837 ), .Z(\AES_ENC/n835 ) );
XOR2_X2 \AES_ENC/U1544  ( .A(\AES_ENC/sa11_sub[1] ), .B(\AES_ENC/sa22_sub[1] ), .Z(\AES_ENC/n836 ) );
XOR2_X2 \AES_ENC/U1543  ( .A(\AES_ENC/w0[18] ), .B(\AES_ENC/sa00_sub[2] ),.Z(\AES_ENC/n837 ) );
XOR2_X2 \AES_ENC/U1542  ( .A(\AES_ENC/n839 ), .B(\AES_ENC/n838 ), .Z(\AES_ENC/sa10_next [1]) );
XOR2_X2 \AES_ENC/U1541  ( .A(\AES_ENC/n841 ), .B(\AES_ENC/n840 ), .Z(\AES_ENC/n838 ) );
XOR2_X2 \AES_ENC/U1540  ( .A(\AES_ENC/n1159 ), .B(\AES_ENC/n1165 ), .Z(\AES_ENC/n839 ) );
XOR2_X2 \AES_ENC/U1539  ( .A(\AES_ENC/sa11_sub[0] ), .B(\AES_ENC/sa22_sub[0] ), .Z(\AES_ENC/n840 ) );
XOR2_X2 \AES_ENC/U1538  ( .A(\AES_ENC/w0[17] ), .B(\AES_ENC/sa00_sub[1] ),.Z(\AES_ENC/n841 ) );
XOR2_X2 \AES_ENC/U1537  ( .A(\AES_ENC/n843 ), .B(\AES_ENC/n842 ), .Z(\AES_ENC/sa10_next [0]) );
XOR2_X2 \AES_ENC/U1536  ( .A(\AES_ENC/n1159 ), .B(\AES_ENC/n1166 ), .Z(\AES_ENC/n842 ) );
XOR2_X2 \AES_ENC/U1535  ( .A(\AES_ENC/w0[16] ), .B(\AES_ENC/sa00_sub[0] ),.Z(\AES_ENC/n843 ) );
XOR2_X2 \AES_ENC/U1534  ( .A(\AES_ENC/n845 ), .B(\AES_ENC/n844 ), .Z(\AES_ENC/sa20_next [7]) );
XOR2_X2 \AES_ENC/U1533  ( .A(\AES_ENC/n1168 ), .B(\AES_ENC/n1160 ), .Z(\AES_ENC/n844 ) );
XOR2_X2 \AES_ENC/U1532  ( .A(\AES_ENC/w0[15] ), .B(\AES_ENC/sa33_sub[7] ),.Z(\AES_ENC/n845 ) );
XOR2_X2 \AES_ENC/U1531  ( .A(\AES_ENC/n847 ), .B(\AES_ENC/n846 ), .Z(\AES_ENC/sa20_next [6]) );
XOR2_X2 \AES_ENC/U1530  ( .A(\AES_ENC/n1169 ), .B(\AES_ENC/n1161 ), .Z(\AES_ENC/n846 ) );
XOR2_X2 \AES_ENC/U1529  ( .A(\AES_ENC/w0[14] ), .B(\AES_ENC/sa33_sub[6] ),.Z(\AES_ENC/n847 ) );
XOR2_X2 \AES_ENC/U1528  ( .A(\AES_ENC/n849 ), .B(\AES_ENC/n848 ), .Z(\AES_ENC/sa20_next [5]) );
XOR2_X2 \AES_ENC/U1527  ( .A(\AES_ENC/n1170 ), .B(\AES_ENC/n1162 ), .Z(\AES_ENC/n848 ) );
XOR2_X2 \AES_ENC/U1526  ( .A(\AES_ENC/w0[13] ), .B(\AES_ENC/sa33_sub[5] ),.Z(\AES_ENC/n849 ) );
XOR2_X2 \AES_ENC/U1525  ( .A(\AES_ENC/n851 ), .B(\AES_ENC/n850 ), .Z(\AES_ENC/sa20_next [4]) );
XOR2_X2 \AES_ENC/U1524  ( .A(\AES_ENC/n1163 ), .B(\AES_ENC/n852 ), .Z(\AES_ENC/n850 ) );
XOR2_X2 \AES_ENC/U1523  ( .A(\AES_ENC/n1167 ), .B(\AES_ENC/n1171 ), .Z(\AES_ENC/n851 ) );
XOR2_X2 \AES_ENC/U1522  ( .A(\AES_ENC/w0[12] ), .B(\AES_ENC/sa33_sub[4] ),.Z(\AES_ENC/n852 ) );
XOR2_X2 \AES_ENC/U1521  ( .A(\AES_ENC/n854 ), .B(\AES_ENC/n853 ), .Z(\AES_ENC/sa20_next [3]) );
XOR2_X2 \AES_ENC/U1520  ( .A(\AES_ENC/n1164 ), .B(\AES_ENC/n855 ), .Z(\AES_ENC/n853 ) );
XOR2_X2 \AES_ENC/U1519  ( .A(\AES_ENC/n1167 ), .B(\AES_ENC/n1172 ), .Z(\AES_ENC/n854 ) );
XOR2_X2 \AES_ENC/U1518  ( .A(\AES_ENC/w0[11] ), .B(\AES_ENC/sa33_sub[3] ),.Z(\AES_ENC/n855 ) );
XOR2_X2 \AES_ENC/U1517  ( .A(\AES_ENC/n857 ), .B(\AES_ENC/n856 ), .Z(\AES_ENC/sa20_next [2]) );
XOR2_X2 \AES_ENC/U1516  ( .A(\AES_ENC/n1173 ), .B(\AES_ENC/n1165 ), .Z(\AES_ENC/n856 ) );
XOR2_X2 \AES_ENC/U1515  ( .A(\AES_ENC/w0[10] ), .B(\AES_ENC/sa33_sub[2] ),.Z(\AES_ENC/n857 ) );
XOR2_X2 \AES_ENC/U1514  ( .A(\AES_ENC/n859 ), .B(\AES_ENC/n858 ), .Z(\AES_ENC/sa20_next [1]) );
XOR2_X2 \AES_ENC/U1513  ( .A(\AES_ENC/n1166 ), .B(\AES_ENC/n860 ), .Z(\AES_ENC/n858 ) );
XOR2_X2 \AES_ENC/U1512  ( .A(\AES_ENC/n1167 ), .B(\AES_ENC/n1174 ), .Z(\AES_ENC/n859 ) );
XOR2_X2 \AES_ENC/U1511  ( .A(\AES_ENC/w0[9] ), .B(\AES_ENC/sa33_sub[1] ),.Z(\AES_ENC/n860 ) );
XOR2_X2 \AES_ENC/U1510  ( .A(\AES_ENC/n862 ), .B(\AES_ENC/n861 ), .Z(\AES_ENC/sa20_next [0]) );
XOR2_X2 \AES_ENC/U1509  ( .A(\AES_ENC/n1167 ), .B(\AES_ENC/n1175 ), .Z(\AES_ENC/n861 ) );
XOR2_X2 \AES_ENC/U1508  ( .A(\AES_ENC/w0[8] ), .B(\AES_ENC/sa33_sub[0] ),.Z(\AES_ENC/n862 ) );
XOR2_X2 \AES_ENC/U1507  ( .A(\AES_ENC/n864 ), .B(\AES_ENC/n863 ), .Z(\AES_ENC/sa30_next [7]) );
XOR2_X2 \AES_ENC/U1506  ( .A(\AES_ENC/n1168 ), .B(\AES_ENC/n865 ), .Z(\AES_ENC/n863 ) );
XOR2_X2 \AES_ENC/U1505  ( .A(\AES_ENC/sa22_sub[7] ), .B(\AES_ENC/sa33_sub[6] ), .Z(\AES_ENC/n864 ) );
XOR2_X2 \AES_ENC/U1504  ( .A(\AES_ENC/w0[7] ), .B(\AES_ENC/sa00_sub[6] ),.Z(\AES_ENC/n865 ) );
XOR2_X2 \AES_ENC/U1503  ( .A(\AES_ENC/n867 ), .B(\AES_ENC/n866 ), .Z(\AES_ENC/sa30_next [6]) );
XOR2_X2 \AES_ENC/U1502  ( .A(\AES_ENC/n1169 ), .B(\AES_ENC/n868 ), .Z(\AES_ENC/n866 ) );
XOR2_X2 \AES_ENC/U1501  ( .A(\AES_ENC/sa22_sub[6] ), .B(\AES_ENC/sa33_sub[5] ), .Z(\AES_ENC/n867 ) );
XOR2_X2 \AES_ENC/U1500  ( .A(\AES_ENC/w0[6] ), .B(\AES_ENC/sa00_sub[5] ),.Z(\AES_ENC/n868 ) );
XOR2_X2 \AES_ENC/U1499  ( .A(\AES_ENC/n870 ), .B(\AES_ENC/n869 ), .Z(\AES_ENC/sa30_next [5]) );
XOR2_X2 \AES_ENC/U1498  ( .A(\AES_ENC/n1170 ), .B(\AES_ENC/n871 ), .Z(\AES_ENC/n869 ) );
XOR2_X2 \AES_ENC/U1497  ( .A(\AES_ENC/sa22_sub[5] ), .B(\AES_ENC/sa33_sub[4] ), .Z(\AES_ENC/n870 ) );
XOR2_X2 \AES_ENC/U1496  ( .A(\AES_ENC/w0[5] ), .B(\AES_ENC/sa00_sub[4] ),.Z(\AES_ENC/n871 ) );
XOR2_X2 \AES_ENC/U1495  ( .A(\AES_ENC/sa00_sub[7] ), .B(\AES_ENC/sa33_sub[7] ), .Z(\AES_ENC/n1176 ) );
XOR2_X2 \AES_ENC/U1494  ( .A(\AES_ENC/n873 ), .B(\AES_ENC/n872 ), .Z(\AES_ENC/sa30_next [4]) );
XOR2_X2 \AES_ENC/U1493  ( .A(\AES_ENC/n875 ), .B(\AES_ENC/n874 ), .Z(\AES_ENC/n872 ) );
XOR2_X2 \AES_ENC/U1492  ( .A(\AES_ENC/n1176 ), .B(\AES_ENC/n1171 ), .Z(\AES_ENC/n873 ) );
XOR2_X2 \AES_ENC/U1491  ( .A(\AES_ENC/sa22_sub[4] ), .B(\AES_ENC/sa33_sub[3] ), .Z(\AES_ENC/n874 ) );
XOR2_X2 \AES_ENC/U1490  ( .A(\AES_ENC/w0[4] ), .B(\AES_ENC/sa00_sub[3] ),.Z(\AES_ENC/n875 ) );
XOR2_X2 \AES_ENC/U1489  ( .A(\AES_ENC/n877 ), .B(\AES_ENC/n876 ), .Z(\AES_ENC/sa30_next [3]) );
XOR2_X2 \AES_ENC/U1488  ( .A(\AES_ENC/n879 ), .B(\AES_ENC/n878 ), .Z(\AES_ENC/n876 ) );
XOR2_X2 \AES_ENC/U1487  ( .A(\AES_ENC/n1176 ), .B(\AES_ENC/n1172 ), .Z(\AES_ENC/n877 ) );
XOR2_X2 \AES_ENC/U1486  ( .A(\AES_ENC/sa22_sub[3] ), .B(\AES_ENC/sa33_sub[2] ), .Z(\AES_ENC/n878 ) );
XOR2_X2 \AES_ENC/U1485  ( .A(\AES_ENC/w0[3] ), .B(\AES_ENC/sa00_sub[2] ),.Z(\AES_ENC/n879 ) );
XOR2_X2 \AES_ENC/U1484  ( .A(\AES_ENC/n881 ), .B(\AES_ENC/n880 ), .Z(\AES_ENC/sa30_next [2]) );
XOR2_X2 \AES_ENC/U1483  ( .A(\AES_ENC/n1173 ), .B(\AES_ENC/n882 ), .Z(\AES_ENC/n880 ) );
XOR2_X2 \AES_ENC/U1482  ( .A(\AES_ENC/sa22_sub[2] ), .B(\AES_ENC/sa33_sub[1] ), .Z(\AES_ENC/n881 ) );
XOR2_X2 \AES_ENC/U1481  ( .A(\AES_ENC/w0[2] ), .B(\AES_ENC/sa00_sub[1] ),.Z(\AES_ENC/n882 ) );
XOR2_X2 \AES_ENC/U1480  ( .A(\AES_ENC/n884 ), .B(\AES_ENC/n883 ), .Z(\AES_ENC/sa30_next [1]) );
XOR2_X2 \AES_ENC/U1479  ( .A(\AES_ENC/n886 ), .B(\AES_ENC/n885 ), .Z(\AES_ENC/n883 ) );
XOR2_X2 \AES_ENC/U1478  ( .A(\AES_ENC/n1176 ), .B(\AES_ENC/n1174 ), .Z(\AES_ENC/n884 ) );
XOR2_X2 \AES_ENC/U1477  ( .A(\AES_ENC/sa22_sub[1] ), .B(\AES_ENC/sa33_sub[0] ), .Z(\AES_ENC/n885 ) );
XOR2_X2 \AES_ENC/U1476  ( .A(\AES_ENC/w0[1] ), .B(\AES_ENC/sa00_sub[0] ),.Z(\AES_ENC/n886 ) );
XOR2_X2 \AES_ENC/U1475  ( .A(\AES_ENC/n888 ), .B(\AES_ENC/n887 ), .Z(\AES_ENC/sa30_next [0]) );
XOR2_X2 \AES_ENC/U1474  ( .A(\AES_ENC/n1176 ), .B(\AES_ENC/n1175 ), .Z(\AES_ENC/n887 ) );
XOR2_X2 \AES_ENC/U1473  ( .A(\AES_ENC/w0[0] ), .B(\AES_ENC/sa22_sub[0] ),.Z(\AES_ENC/n888 ) );
XOR2_X2 \AES_ENC/U1472  ( .A(\AES_ENC/sa23_sub[7] ), .B(\AES_ENC/sa30_sub[7] ), .Z(\AES_ENC/n1185 ) );
XOR2_X2 \AES_ENC/U1471  ( .A(\AES_ENC/sa01_sub[6] ), .B(\AES_ENC/sa12_sub[6] ), .Z(\AES_ENC/n1187 ) );
XOR2_X2 \AES_ENC/U1470  ( .A(\AES_ENC/n890 ), .B(\AES_ENC/n889 ), .Z(\AES_ENC/sa01_next [7]) );
XOR2_X2 \AES_ENC/U1469  ( .A(\AES_ENC/n1185 ), .B(\AES_ENC/n1187 ), .Z(\AES_ENC/n889 ) );
XOR2_X2 \AES_ENC/U1468  ( .A(\AES_ENC/w1[31] ), .B(\AES_ENC/sa12_sub[7] ),.Z(\AES_ENC/n890 ) );
XOR2_X2 \AES_ENC/U1467  ( .A(\AES_ENC/sa01_sub[5] ), .B(\AES_ENC/sa12_sub[5] ), .Z(\AES_ENC/n1188 ) );
XOR2_X2 \AES_ENC/U1466  ( .A(\AES_ENC/sa23_sub[6] ), .B(\AES_ENC/sa30_sub[6] ), .Z(\AES_ENC/n1178 ) );
XOR2_X2 \AES_ENC/U1465  ( .A(\AES_ENC/n892 ), .B(\AES_ENC/n891 ), .Z(\AES_ENC/sa01_next [6]) );
XOR2_X2 \AES_ENC/U1464  ( .A(\AES_ENC/n1188 ), .B(\AES_ENC/n1178 ), .Z(\AES_ENC/n891 ) );
XOR2_X2 \AES_ENC/U1463  ( .A(\AES_ENC/w1[30] ), .B(\AES_ENC/sa12_sub[6] ),.Z(\AES_ENC/n892 ) );
XOR2_X2 \AES_ENC/U1462  ( .A(\AES_ENC/sa01_sub[4] ), .B(\AES_ENC/sa12_sub[4] ), .Z(\AES_ENC/n1189 ) );
XOR2_X2 \AES_ENC/U1461  ( .A(\AES_ENC/sa23_sub[5] ), .B(\AES_ENC/sa30_sub[5] ), .Z(\AES_ENC/n1179 ) );
XOR2_X2 \AES_ENC/U1460  ( .A(\AES_ENC/n894 ), .B(\AES_ENC/n893 ), .Z(\AES_ENC/sa01_next [5]) );
XOR2_X2 \AES_ENC/U1459  ( .A(\AES_ENC/n1189 ), .B(\AES_ENC/n1179 ), .Z(\AES_ENC/n893 ) );
XOR2_X2 \AES_ENC/U1458  ( .A(\AES_ENC/w1[29] ), .B(\AES_ENC/sa12_sub[5] ),.Z(\AES_ENC/n894 ) );
XOR2_X2 \AES_ENC/U1457  ( .A(\AES_ENC/sa01_sub[7] ), .B(\AES_ENC/sa12_sub[7] ), .Z(\AES_ENC/n1186 ) );
XOR2_X2 \AES_ENC/U1456  ( .A(\AES_ENC/sa01_sub[3] ), .B(\AES_ENC/sa12_sub[3] ), .Z(\AES_ENC/n1190 ) );
XOR2_X2 \AES_ENC/U1455  ( .A(\AES_ENC/sa23_sub[4] ), .B(\AES_ENC/sa30_sub[4] ), .Z(\AES_ENC/n1180 ) );
XOR2_X2 \AES_ENC/U1454  ( .A(\AES_ENC/n896 ), .B(\AES_ENC/n895 ), .Z(\AES_ENC/sa01_next [4]) );
XOR2_X2 \AES_ENC/U1453  ( .A(\AES_ENC/n1180 ), .B(\AES_ENC/n897 ), .Z(\AES_ENC/n895 ) );
XOR2_X2 \AES_ENC/U1452  ( .A(\AES_ENC/n1186 ), .B(\AES_ENC/n1190 ), .Z(\AES_ENC/n896 ) );
XOR2_X2 \AES_ENC/U1451  ( .A(\AES_ENC/w1[28] ), .B(\AES_ENC/sa12_sub[4] ),.Z(\AES_ENC/n897 ) );
XOR2_X2 \AES_ENC/U1450  ( .A(\AES_ENC/sa01_sub[2] ), .B(\AES_ENC/sa12_sub[2] ), .Z(\AES_ENC/n1191 ) );
XOR2_X2 \AES_ENC/U1449  ( .A(\AES_ENC/sa23_sub[3] ), .B(\AES_ENC/sa30_sub[3] ), .Z(\AES_ENC/n1181 ) );
XOR2_X2 \AES_ENC/U1448  ( .A(\AES_ENC/n899 ), .B(\AES_ENC/n898 ), .Z(\AES_ENC/sa01_next [3]) );
XOR2_X2 \AES_ENC/U1447  ( .A(\AES_ENC/n1181 ), .B(\AES_ENC/n900 ), .Z(\AES_ENC/n898 ) );
XOR2_X2 \AES_ENC/U1446  ( .A(\AES_ENC/n1186 ), .B(\AES_ENC/n1191 ), .Z(\AES_ENC/n899 ) );
XOR2_X2 \AES_ENC/U1445  ( .A(\AES_ENC/w1[27] ), .B(\AES_ENC/sa12_sub[3] ),.Z(\AES_ENC/n900 ) );
XOR2_X2 \AES_ENC/U1444  ( .A(\AES_ENC/sa01_sub[1] ), .B(\AES_ENC/sa12_sub[1] ), .Z(\AES_ENC/n1192 ) );
XOR2_X2 \AES_ENC/U1443  ( .A(\AES_ENC/sa23_sub[2] ), .B(\AES_ENC/sa30_sub[2] ), .Z(\AES_ENC/n1182 ) );
XOR2_X2 \AES_ENC/U1442  ( .A(\AES_ENC/n902 ), .B(\AES_ENC/n901 ), .Z(\AES_ENC/sa01_next [2]) );
XOR2_X2 \AES_ENC/U1441  ( .A(\AES_ENC/n1192 ), .B(\AES_ENC/n1182 ), .Z(\AES_ENC/n901 ) );
XOR2_X2 \AES_ENC/U1440  ( .A(\AES_ENC/w1[26] ), .B(\AES_ENC/sa12_sub[2] ),.Z(\AES_ENC/n902 ) );
XOR2_X2 \AES_ENC/U1439  ( .A(\AES_ENC/sa01_sub[0] ), .B(\AES_ENC/sa12_sub[0] ), .Z(\AES_ENC/n1193 ) );
XOR2_X2 \AES_ENC/U1438  ( .A(\AES_ENC/sa23_sub[1] ), .B(\AES_ENC/sa30_sub[1] ), .Z(\AES_ENC/n1183 ) );
XOR2_X2 \AES_ENC/U1437  ( .A(\AES_ENC/n904 ), .B(\AES_ENC/n903 ), .Z(\AES_ENC/sa01_next [1]) );
XOR2_X2 \AES_ENC/U1436  ( .A(\AES_ENC/n1183 ), .B(\AES_ENC/n905 ), .Z(\AES_ENC/n903 ) );
XOR2_X2 \AES_ENC/U1435  ( .A(\AES_ENC/n1186 ), .B(\AES_ENC/n1193 ), .Z(\AES_ENC/n904 ) );
XOR2_X2 \AES_ENC/U1434  ( .A(\AES_ENC/w1[25] ), .B(\AES_ENC/sa12_sub[1] ),.Z(\AES_ENC/n905 ) );
XOR2_X2 \AES_ENC/U1433  ( .A(\AES_ENC/sa23_sub[0] ), .B(\AES_ENC/sa30_sub[0] ), .Z(\AES_ENC/n1184 ) );
XOR2_X2 \AES_ENC/U1432  ( .A(\AES_ENC/n907 ), .B(\AES_ENC/n906 ), .Z(\AES_ENC/sa01_next [0]) );
XOR2_X2 \AES_ENC/U1431  ( .A(\AES_ENC/n1186 ), .B(\AES_ENC/n1184 ), .Z(\AES_ENC/n906 ) );
XOR2_X2 \AES_ENC/U1430  ( .A(\AES_ENC/w1[24] ), .B(\AES_ENC/sa12_sub[0] ),.Z(\AES_ENC/n907 ) );
XOR2_X2 \AES_ENC/U1429  ( .A(\AES_ENC/n909 ), .B(\AES_ENC/n908 ), .Z(\AES_ENC/sa11_next [7]) );
XOR2_X2 \AES_ENC/U1428  ( .A(\AES_ENC/n1185 ), .B(\AES_ENC/n910 ), .Z(\AES_ENC/n908 ) );
XOR2_X2 \AES_ENC/U1427  ( .A(\AES_ENC/sa12_sub[6] ), .B(\AES_ENC/sa23_sub[6] ), .Z(\AES_ENC/n909 ) );
XOR2_X2 \AES_ENC/U1426  ( .A(\AES_ENC/w1[23] ), .B(\AES_ENC/sa01_sub[7] ),.Z(\AES_ENC/n910 ) );
XOR2_X2 \AES_ENC/U1425  ( .A(\AES_ENC/n912 ), .B(\AES_ENC/n911 ), .Z(\AES_ENC/sa11_next [6]) );
XOR2_X2 \AES_ENC/U1424  ( .A(\AES_ENC/n1178 ), .B(\AES_ENC/n913 ), .Z(\AES_ENC/n911 ) );
XOR2_X2 \AES_ENC/U1423  ( .A(\AES_ENC/sa12_sub[5] ), .B(\AES_ENC/sa23_sub[5] ), .Z(\AES_ENC/n912 ) );
XOR2_X2 \AES_ENC/U1422  ( .A(\AES_ENC/w1[22] ), .B(\AES_ENC/sa01_sub[6] ),.Z(\AES_ENC/n913 ) );
XOR2_X2 \AES_ENC/U1421  ( .A(\AES_ENC/n915 ), .B(\AES_ENC/n914 ), .Z(\AES_ENC/sa11_next [5]) );
XOR2_X2 \AES_ENC/U1420  ( .A(\AES_ENC/n1179 ), .B(\AES_ENC/n916 ), .Z(\AES_ENC/n914 ) );
XOR2_X2 \AES_ENC/U1419  ( .A(\AES_ENC/sa12_sub[4] ), .B(\AES_ENC/sa23_sub[4] ), .Z(\AES_ENC/n915 ) );
XOR2_X2 \AES_ENC/U1418  ( .A(\AES_ENC/w1[21] ), .B(\AES_ENC/sa01_sub[5] ),.Z(\AES_ENC/n916 ) );
XOR2_X2 \AES_ENC/U1417  ( .A(\AES_ENC/sa12_sub[7] ), .B(\AES_ENC/sa23_sub[7] ), .Z(\AES_ENC/n1177 ) );
XOR2_X2 \AES_ENC/U1416  ( .A(\AES_ENC/n918 ), .B(\AES_ENC/n917 ), .Z(\AES_ENC/sa11_next [4]) );
XOR2_X2 \AES_ENC/U1415  ( .A(\AES_ENC/n920 ), .B(\AES_ENC/n919 ), .Z(\AES_ENC/n917 ) );
XOR2_X2 \AES_ENC/U1414  ( .A(\AES_ENC/n1177 ), .B(\AES_ENC/n1180 ), .Z(\AES_ENC/n918 ) );
XOR2_X2 \AES_ENC/U1413  ( .A(\AES_ENC/sa12_sub[3] ), .B(\AES_ENC/sa23_sub[3] ), .Z(\AES_ENC/n919 ) );
XOR2_X2 \AES_ENC/U1412  ( .A(\AES_ENC/w1[20] ), .B(\AES_ENC/sa01_sub[4] ),.Z(\AES_ENC/n920 ) );
XOR2_X2 \AES_ENC/U1411  ( .A(\AES_ENC/n922 ), .B(\AES_ENC/n921 ), .Z(\AES_ENC/sa11_next [3]) );
XOR2_X2 \AES_ENC/U1410  ( .A(\AES_ENC/n924 ), .B(\AES_ENC/n923 ), .Z(\AES_ENC/n921 ) );
XOR2_X2 \AES_ENC/U1409  ( .A(\AES_ENC/n1177 ), .B(\AES_ENC/n1181 ), .Z(\AES_ENC/n922 ) );
XOR2_X2 \AES_ENC/U1408  ( .A(\AES_ENC/sa12_sub[2] ), .B(\AES_ENC/sa23_sub[2] ), .Z(\AES_ENC/n923 ) );
XOR2_X2 \AES_ENC/U1407  ( .A(\AES_ENC/w1[19] ), .B(\AES_ENC/sa01_sub[3] ),.Z(\AES_ENC/n924 ) );
XOR2_X2 \AES_ENC/U1406  ( .A(\AES_ENC/n926 ), .B(\AES_ENC/n925 ), .Z(\AES_ENC/sa11_next [2]) );
XOR2_X2 \AES_ENC/U1405  ( .A(\AES_ENC/n1182 ), .B(\AES_ENC/n927 ), .Z(\AES_ENC/n925 ) );
XOR2_X2 \AES_ENC/U1404  ( .A(\AES_ENC/sa12_sub[1] ), .B(\AES_ENC/sa23_sub[1] ), .Z(\AES_ENC/n926 ) );
XOR2_X2 \AES_ENC/U1403  ( .A(\AES_ENC/w1[18] ), .B(\AES_ENC/sa01_sub[2] ),.Z(\AES_ENC/n927 ) );
XOR2_X2 \AES_ENC/U1402  ( .A(\AES_ENC/n929 ), .B(\AES_ENC/n928 ), .Z(\AES_ENC/sa11_next [1]) );
XOR2_X2 \AES_ENC/U1401  ( .A(\AES_ENC/n931 ), .B(\AES_ENC/n930 ), .Z(\AES_ENC/n928 ) );
XOR2_X2 \AES_ENC/U1400  ( .A(\AES_ENC/n1177 ), .B(\AES_ENC/n1183 ), .Z(\AES_ENC/n929 ) );
XOR2_X2 \AES_ENC/U1399  ( .A(\AES_ENC/sa12_sub[0] ), .B(\AES_ENC/sa23_sub[0] ), .Z(\AES_ENC/n930 ) );
XOR2_X2 \AES_ENC/U1398  ( .A(\AES_ENC/w1[17] ), .B(\AES_ENC/sa01_sub[1] ),.Z(\AES_ENC/n931 ) );
XOR2_X2 \AES_ENC/U1397  ( .A(\AES_ENC/n933 ), .B(\AES_ENC/n932 ), .Z(\AES_ENC/sa11_next [0]) );
XOR2_X2 \AES_ENC/U1396  ( .A(\AES_ENC/n1177 ), .B(\AES_ENC/n1184 ), .Z(\AES_ENC/n932 ) );
XOR2_X2 \AES_ENC/U1395  ( .A(\AES_ENC/w1[16] ), .B(\AES_ENC/sa01_sub[0] ),.Z(\AES_ENC/n933 ) );
XOR2_X2 \AES_ENC/U1394  ( .A(\AES_ENC/n935 ), .B(\AES_ENC/n934 ), .Z(\AES_ENC/sa21_next [7]) );
XOR2_X2 \AES_ENC/U1393  ( .A(\AES_ENC/n1186 ), .B(\AES_ENC/n1178 ), .Z(\AES_ENC/n934 ) );
XOR2_X2 \AES_ENC/U1392  ( .A(\AES_ENC/w1[15] ), .B(\AES_ENC/sa30_sub[7] ),.Z(\AES_ENC/n935 ) );
XOR2_X2 \AES_ENC/U1391  ( .A(\AES_ENC/n937 ), .B(\AES_ENC/n936 ), .Z(\AES_ENC/sa21_next [6]) );
XOR2_X2 \AES_ENC/U1390  ( .A(\AES_ENC/n1187 ), .B(\AES_ENC/n1179 ), .Z(\AES_ENC/n936 ) );
XOR2_X2 \AES_ENC/U1389  ( .A(\AES_ENC/w1[14] ), .B(\AES_ENC/sa30_sub[6] ),.Z(\AES_ENC/n937 ) );
XOR2_X2 \AES_ENC/U1388  ( .A(\AES_ENC/n939 ), .B(\AES_ENC/n938 ), .Z(\AES_ENC/sa21_next [5]) );
XOR2_X2 \AES_ENC/U1387  ( .A(\AES_ENC/n1188 ), .B(\AES_ENC/n1180 ), .Z(\AES_ENC/n938 ) );
XOR2_X2 \AES_ENC/U1386  ( .A(\AES_ENC/w1[13] ), .B(\AES_ENC/sa30_sub[5] ),.Z(\AES_ENC/n939 ) );
XOR2_X2 \AES_ENC/U1385  ( .A(\AES_ENC/n941 ), .B(\AES_ENC/n940 ), .Z(\AES_ENC/sa21_next [4]) );
XOR2_X2 \AES_ENC/U1384  ( .A(\AES_ENC/n1181 ), .B(\AES_ENC/n942 ), .Z(\AES_ENC/n940 ) );
XOR2_X2 \AES_ENC/U1383  ( .A(\AES_ENC/n1185 ), .B(\AES_ENC/n1189 ), .Z(\AES_ENC/n941 ) );
XOR2_X2 \AES_ENC/U1382  ( .A(\AES_ENC/w1[12] ), .B(\AES_ENC/sa30_sub[4] ),.Z(\AES_ENC/n942 ) );
XOR2_X2 \AES_ENC/U1381  ( .A(\AES_ENC/n944 ), .B(\AES_ENC/n943 ), .Z(\AES_ENC/sa21_next [3]) );
XOR2_X2 \AES_ENC/U1380  ( .A(\AES_ENC/n1182 ), .B(\AES_ENC/n945 ), .Z(\AES_ENC/n943 ) );
XOR2_X2 \AES_ENC/U1379  ( .A(\AES_ENC/n1185 ), .B(\AES_ENC/n1190 ), .Z(\AES_ENC/n944 ) );
XOR2_X2 \AES_ENC/U1378  ( .A(\AES_ENC/w1[11] ), .B(\AES_ENC/sa30_sub[3] ),.Z(\AES_ENC/n945 ) );
XOR2_X2 \AES_ENC/U1377  ( .A(\AES_ENC/n947 ), .B(\AES_ENC/n946 ), .Z(\AES_ENC/sa21_next [2]) );
XOR2_X2 \AES_ENC/U1376  ( .A(\AES_ENC/n1191 ), .B(\AES_ENC/n1183 ), .Z(\AES_ENC/n946 ) );
XOR2_X2 \AES_ENC/U1375  ( .A(\AES_ENC/w1[10] ), .B(\AES_ENC/sa30_sub[2] ),.Z(\AES_ENC/n947 ) );
XOR2_X2 \AES_ENC/U1374  ( .A(\AES_ENC/n949 ), .B(\AES_ENC/n948 ), .Z(\AES_ENC/sa21_next [1]) );
XOR2_X2 \AES_ENC/U1373  ( .A(\AES_ENC/n1184 ), .B(\AES_ENC/n950 ), .Z(\AES_ENC/n948 ) );
XOR2_X2 \AES_ENC/U1372  ( .A(\AES_ENC/n1185 ), .B(\AES_ENC/n1192 ), .Z(\AES_ENC/n949 ) );
XOR2_X2 \AES_ENC/U1371  ( .A(\AES_ENC/w1[9] ), .B(\AES_ENC/sa30_sub[1] ),.Z(\AES_ENC/n950 ) );
XOR2_X2 \AES_ENC/U1370  ( .A(\AES_ENC/n952 ), .B(\AES_ENC/n951 ), .Z(\AES_ENC/sa21_next [0]) );
XOR2_X2 \AES_ENC/U1369  ( .A(\AES_ENC/n1185 ), .B(\AES_ENC/n1193 ), .Z(\AES_ENC/n951 ) );
XOR2_X2 \AES_ENC/U1368  ( .A(\AES_ENC/w1[8] ), .B(\AES_ENC/sa30_sub[0] ),.Z(\AES_ENC/n952 ) );
XOR2_X2 \AES_ENC/U1367  ( .A(\AES_ENC/n954 ), .B(\AES_ENC/n953 ), .Z(\AES_ENC/sa31_next [7]) );
XOR2_X2 \AES_ENC/U1366  ( .A(\AES_ENC/n1186 ), .B(\AES_ENC/n955 ), .Z(\AES_ENC/n953 ) );
XOR2_X2 \AES_ENC/U1365  ( .A(\AES_ENC/sa23_sub[7] ), .B(\AES_ENC/sa30_sub[6] ), .Z(\AES_ENC/n954 ) );
XOR2_X2 \AES_ENC/U1364  ( .A(\AES_ENC/w1[7] ), .B(\AES_ENC/sa01_sub[6] ),.Z(\AES_ENC/n955 ) );
XOR2_X2 \AES_ENC/U1363  ( .A(\AES_ENC/n957 ), .B(\AES_ENC/n956 ), .Z(\AES_ENC/sa31_next [6]) );
XOR2_X2 \AES_ENC/U1362  ( .A(\AES_ENC/n1187 ), .B(\AES_ENC/n958 ), .Z(\AES_ENC/n956 ) );
XOR2_X2 \AES_ENC/U1361  ( .A(\AES_ENC/sa23_sub[6] ), .B(\AES_ENC/sa30_sub[5] ), .Z(\AES_ENC/n957 ) );
XOR2_X2 \AES_ENC/U1360  ( .A(\AES_ENC/w1[6] ), .B(\AES_ENC/sa01_sub[5] ),.Z(\AES_ENC/n958 ) );
XOR2_X2 \AES_ENC/U1359  ( .A(\AES_ENC/n960 ), .B(\AES_ENC/n959 ), .Z(\AES_ENC/sa31_next [5]) );
XOR2_X2 \AES_ENC/U1358  ( .A(\AES_ENC/n1188 ), .B(\AES_ENC/n961 ), .Z(\AES_ENC/n959 ) );
XOR2_X2 \AES_ENC/U1357  ( .A(\AES_ENC/sa23_sub[5] ), .B(\AES_ENC/sa30_sub[4] ), .Z(\AES_ENC/n960 ) );
XOR2_X2 \AES_ENC/U1356  ( .A(\AES_ENC/w1[5] ), .B(\AES_ENC/sa01_sub[4] ),.Z(\AES_ENC/n961 ) );
XOR2_X2 \AES_ENC/U1355  ( .A(\AES_ENC/sa01_sub[7] ), .B(\AES_ENC/sa30_sub[7] ), .Z(\AES_ENC/n1194 ) );
XOR2_X2 \AES_ENC/U1354  ( .A(\AES_ENC/n963 ), .B(\AES_ENC/n962 ), .Z(\AES_ENC/sa31_next [4]) );
XOR2_X2 \AES_ENC/U1353  ( .A(\AES_ENC/n965 ), .B(\AES_ENC/n964 ), .Z(\AES_ENC/n962 ) );
XOR2_X2 \AES_ENC/U1352  ( .A(\AES_ENC/n1194 ), .B(\AES_ENC/n1189 ), .Z(\AES_ENC/n963 ) );
XOR2_X2 \AES_ENC/U1351  ( .A(\AES_ENC/sa23_sub[4] ), .B(\AES_ENC/sa30_sub[3] ), .Z(\AES_ENC/n964 ) );
XOR2_X2 \AES_ENC/U1350  ( .A(\AES_ENC/w1[4] ), .B(\AES_ENC/sa01_sub[3] ),.Z(\AES_ENC/n965 ) );
XOR2_X2 \AES_ENC/U1349  ( .A(\AES_ENC/n967 ), .B(\AES_ENC/n966 ), .Z(\AES_ENC/sa31_next [3]) );
XOR2_X2 \AES_ENC/U1348  ( .A(\AES_ENC/n969 ), .B(\AES_ENC/n968 ), .Z(\AES_ENC/n966 ) );
XOR2_X2 \AES_ENC/U1347  ( .A(\AES_ENC/n1194 ), .B(\AES_ENC/n1190 ), .Z(\AES_ENC/n967 ) );
XOR2_X2 \AES_ENC/U1346  ( .A(\AES_ENC/sa23_sub[3] ), .B(\AES_ENC/sa30_sub[2] ), .Z(\AES_ENC/n968 ) );
XOR2_X2 \AES_ENC/U1345  ( .A(\AES_ENC/w1[3] ), .B(\AES_ENC/sa01_sub[2] ),.Z(\AES_ENC/n969 ) );
XOR2_X2 \AES_ENC/U1344  ( .A(\AES_ENC/n971 ), .B(\AES_ENC/n970 ), .Z(\AES_ENC/sa31_next [2]) );
XOR2_X2 \AES_ENC/U1343  ( .A(\AES_ENC/n1191 ), .B(\AES_ENC/n972 ), .Z(\AES_ENC/n970 ) );
XOR2_X2 \AES_ENC/U1342  ( .A(\AES_ENC/sa23_sub[2] ), .B(\AES_ENC/sa30_sub[1] ), .Z(\AES_ENC/n971 ) );
XOR2_X2 \AES_ENC/U1341  ( .A(\AES_ENC/w1[2] ), .B(\AES_ENC/sa01_sub[1] ),.Z(\AES_ENC/n972 ) );
XOR2_X2 \AES_ENC/U1340  ( .A(\AES_ENC/n974 ), .B(\AES_ENC/n973 ), .Z(\AES_ENC/sa31_next [1]) );
XOR2_X2 \AES_ENC/U1339  ( .A(\AES_ENC/n976 ), .B(\AES_ENC/n975 ), .Z(\AES_ENC/n973 ) );
XOR2_X2 \AES_ENC/U1338  ( .A(\AES_ENC/n1194 ), .B(\AES_ENC/n1192 ), .Z(\AES_ENC/n974 ) );
XOR2_X2 \AES_ENC/U1337  ( .A(\AES_ENC/sa23_sub[1] ), .B(\AES_ENC/sa30_sub[0] ), .Z(\AES_ENC/n975 ) );
XOR2_X2 \AES_ENC/U1336  ( .A(\AES_ENC/w1[1] ), .B(\AES_ENC/sa01_sub[0] ),.Z(\AES_ENC/n976 ) );
XOR2_X2 \AES_ENC/U1335  ( .A(\AES_ENC/n978 ), .B(\AES_ENC/n977 ), .Z(\AES_ENC/sa31_next [0]) );
XOR2_X2 \AES_ENC/U1334  ( .A(\AES_ENC/n1194 ), .B(\AES_ENC/n1193 ), .Z(\AES_ENC/n977 ) );
XOR2_X2 \AES_ENC/U1333  ( .A(\AES_ENC/w1[0] ), .B(\AES_ENC/sa23_sub[0] ),.Z(\AES_ENC/n978 ) );
XOR2_X2 \AES_ENC/U1332  ( .A(\AES_ENC/sa20_sub[7] ), .B(\AES_ENC/sa31_sub[7] ), .Z(\AES_ENC/n1203 ) );
XOR2_X2 \AES_ENC/U1331  ( .A(\AES_ENC/sa02_sub[6] ), .B(\AES_ENC/sa13_sub[6] ), .Z(\AES_ENC/n1205 ) );
XOR2_X2 \AES_ENC/U1330  ( .A(\AES_ENC/n980 ), .B(\AES_ENC/n979 ), .Z(\AES_ENC/sa02_next [7]) );
XOR2_X2 \AES_ENC/U1329  ( .A(\AES_ENC/n1203 ), .B(\AES_ENC/n1205 ), .Z(\AES_ENC/n979 ) );
XOR2_X2 \AES_ENC/U1328  ( .A(\AES_ENC/w2[31] ), .B(\AES_ENC/sa13_sub[7] ),.Z(\AES_ENC/n980 ) );
XOR2_X2 \AES_ENC/U1327  ( .A(\AES_ENC/sa02_sub[5] ), .B(\AES_ENC/sa13_sub[5] ), .Z(\AES_ENC/n1206 ) );
XOR2_X2 \AES_ENC/U1326  ( .A(\AES_ENC/sa20_sub[6] ), .B(\AES_ENC/sa31_sub[6] ), .Z(\AES_ENC/n1196 ) );
XOR2_X2 \AES_ENC/U1325  ( .A(\AES_ENC/n982 ), .B(\AES_ENC/n981 ), .Z(\AES_ENC/sa02_next [6]) );
XOR2_X2 \AES_ENC/U1324  ( .A(\AES_ENC/n1206 ), .B(\AES_ENC/n1196 ), .Z(\AES_ENC/n981 ) );
XOR2_X2 \AES_ENC/U1323  ( .A(\AES_ENC/w2[30] ), .B(\AES_ENC/sa13_sub[6] ),.Z(\AES_ENC/n982 ) );
XOR2_X2 \AES_ENC/U1322  ( .A(\AES_ENC/sa02_sub[4] ), .B(\AES_ENC/sa13_sub[4] ), .Z(\AES_ENC/n1207 ) );
XOR2_X2 \AES_ENC/U1321  ( .A(\AES_ENC/sa20_sub[5] ), .B(\AES_ENC/sa31_sub[5] ), .Z(\AES_ENC/n1197 ) );
XOR2_X2 \AES_ENC/U1320  ( .A(\AES_ENC/n984 ), .B(\AES_ENC/n983 ), .Z(\AES_ENC/sa02_next [5]) );
XOR2_X2 \AES_ENC/U1319  ( .A(\AES_ENC/n1207 ), .B(\AES_ENC/n1197 ), .Z(\AES_ENC/n983 ) );
XOR2_X2 \AES_ENC/U1318  ( .A(\AES_ENC/w2[29] ), .B(\AES_ENC/sa13_sub[5] ),.Z(\AES_ENC/n984 ) );
XOR2_X2 \AES_ENC/U1317  ( .A(\AES_ENC/sa02_sub[7] ), .B(\AES_ENC/sa13_sub[7] ), .Z(\AES_ENC/n1204 ) );
XOR2_X2 \AES_ENC/U1316  ( .A(\AES_ENC/sa02_sub[3] ), .B(\AES_ENC/sa13_sub[3] ), .Z(\AES_ENC/n1208 ) );
XOR2_X2 \AES_ENC/U1315  ( .A(\AES_ENC/sa20_sub[4] ), .B(\AES_ENC/sa31_sub[4] ), .Z(\AES_ENC/n1198 ) );
XOR2_X2 \AES_ENC/U1314  ( .A(\AES_ENC/n986 ), .B(\AES_ENC/n985 ), .Z(\AES_ENC/sa02_next [4]) );
XOR2_X2 \AES_ENC/U1313  ( .A(\AES_ENC/n1198 ), .B(\AES_ENC/n987 ), .Z(\AES_ENC/n985 ) );
XOR2_X2 \AES_ENC/U1312  ( .A(\AES_ENC/n1204 ), .B(\AES_ENC/n1208 ), .Z(\AES_ENC/n986 ) );
XOR2_X2 \AES_ENC/U1311  ( .A(\AES_ENC/w2[28] ), .B(\AES_ENC/sa13_sub[4] ),.Z(\AES_ENC/n987 ) );
XOR2_X2 \AES_ENC/U1310  ( .A(\AES_ENC/sa02_sub[2] ), .B(\AES_ENC/sa13_sub[2] ), .Z(\AES_ENC/n1209 ) );
XOR2_X2 \AES_ENC/U1309  ( .A(\AES_ENC/sa20_sub[3] ), .B(\AES_ENC/sa31_sub[3] ), .Z(\AES_ENC/n1199 ) );
XOR2_X2 \AES_ENC/U1308  ( .A(\AES_ENC/n989 ), .B(\AES_ENC/n988 ), .Z(\AES_ENC/sa02_next [3]) );
XOR2_X2 \AES_ENC/U1307  ( .A(\AES_ENC/n1199 ), .B(\AES_ENC/n990 ), .Z(\AES_ENC/n988 ) );
XOR2_X2 \AES_ENC/U1306  ( .A(\AES_ENC/n1204 ), .B(\AES_ENC/n1209 ), .Z(\AES_ENC/n989 ) );
XOR2_X2 \AES_ENC/U1305  ( .A(\AES_ENC/w2[27] ), .B(\AES_ENC/sa13_sub[3] ),.Z(\AES_ENC/n990 ) );
XOR2_X2 \AES_ENC/U1304  ( .A(\AES_ENC/sa02_sub[1] ), .B(\AES_ENC/sa13_sub[1] ), .Z(\AES_ENC/n1210 ) );
XOR2_X2 \AES_ENC/U1303  ( .A(\AES_ENC/sa20_sub[2] ), .B(\AES_ENC/sa31_sub[2] ), .Z(\AES_ENC/n1200 ) );
XOR2_X2 \AES_ENC/U1302  ( .A(\AES_ENC/n992 ), .B(\AES_ENC/n991 ), .Z(\AES_ENC/sa02_next [2]) );
XOR2_X2 \AES_ENC/U1301  ( .A(\AES_ENC/n1210 ), .B(\AES_ENC/n1200 ), .Z(\AES_ENC/n991 ) );
XOR2_X2 \AES_ENC/U1300  ( .A(\AES_ENC/w2[26] ), .B(\AES_ENC/sa13_sub[2] ),.Z(\AES_ENC/n992 ) );
XOR2_X2 \AES_ENC/U1299  ( .A(\AES_ENC/sa02_sub[0] ), .B(\AES_ENC/sa13_sub[0] ), .Z(\AES_ENC/n1211 ) );
XOR2_X2 \AES_ENC/U1298  ( .A(\AES_ENC/sa20_sub[1] ), .B(\AES_ENC/sa31_sub[1] ), .Z(\AES_ENC/n1201 ) );
XOR2_X2 \AES_ENC/U1297  ( .A(\AES_ENC/n994 ), .B(\AES_ENC/n993 ), .Z(\AES_ENC/sa02_next [1]) );
XOR2_X2 \AES_ENC/U1296  ( .A(\AES_ENC/n1201 ), .B(\AES_ENC/n995 ), .Z(\AES_ENC/n993 ) );
XOR2_X2 \AES_ENC/U1295  ( .A(\AES_ENC/n1204 ), .B(\AES_ENC/n1211 ), .Z(\AES_ENC/n994 ) );
XOR2_X2 \AES_ENC/U1294  ( .A(\AES_ENC/w2[25] ), .B(\AES_ENC/sa13_sub[1] ),.Z(\AES_ENC/n995 ) );
XOR2_X2 \AES_ENC/U1293  ( .A(\AES_ENC/sa20_sub[0] ), .B(\AES_ENC/sa31_sub[0] ), .Z(\AES_ENC/n1202 ) );
XOR2_X2 \AES_ENC/U1292  ( .A(\AES_ENC/n997 ), .B(\AES_ENC/n996 ), .Z(\AES_ENC/sa02_next [0]) );
XOR2_X2 \AES_ENC/U1291  ( .A(\AES_ENC/n1204 ), .B(\AES_ENC/n1202 ), .Z(\AES_ENC/n996 ) );
XOR2_X2 \AES_ENC/U1290  ( .A(\AES_ENC/w2[24] ), .B(\AES_ENC/sa13_sub[0] ),.Z(\AES_ENC/n997 ) );
XOR2_X2 \AES_ENC/U1289  ( .A(\AES_ENC/n999 ), .B(\AES_ENC/n998 ), .Z(\AES_ENC/sa12_next [7]) );
XOR2_X2 \AES_ENC/U1288  ( .A(\AES_ENC/n1203 ), .B(\AES_ENC/n1000 ), .Z(\AES_ENC/n998 ) );
XOR2_X2 \AES_ENC/U1287  ( .A(\AES_ENC/sa13_sub[6] ), .B(\AES_ENC/sa20_sub[6] ), .Z(\AES_ENC/n999 ) );
XOR2_X2 \AES_ENC/U1286  ( .A(\AES_ENC/w2[23] ), .B(\AES_ENC/sa02_sub[7] ),.Z(\AES_ENC/n1000 ) );
XOR2_X2 \AES_ENC/U1285  ( .A(\AES_ENC/n1002 ), .B(\AES_ENC/n1001 ), .Z(\AES_ENC/sa12_next [6]) );
XOR2_X2 \AES_ENC/U1284  ( .A(\AES_ENC/n1196 ), .B(\AES_ENC/n1003 ), .Z(\AES_ENC/n1001 ) );
XOR2_X2 \AES_ENC/U1283  ( .A(\AES_ENC/sa13_sub[5] ), .B(\AES_ENC/sa20_sub[5] ), .Z(\AES_ENC/n1002 ) );
XOR2_X2 \AES_ENC/U1282  ( .A(\AES_ENC/w2[22] ), .B(\AES_ENC/sa02_sub[6] ),.Z(\AES_ENC/n1003 ) );
XOR2_X2 \AES_ENC/U1281  ( .A(\AES_ENC/n1005 ), .B(\AES_ENC/n1004 ), .Z(\AES_ENC/sa12_next [5]) );
XOR2_X2 \AES_ENC/U1280  ( .A(\AES_ENC/n1197 ), .B(\AES_ENC/n1006 ), .Z(\AES_ENC/n1004 ) );
XOR2_X2 \AES_ENC/U1279  ( .A(\AES_ENC/sa13_sub[4] ), .B(\AES_ENC/sa20_sub[4] ), .Z(\AES_ENC/n1005 ) );
XOR2_X2 \AES_ENC/U1278  ( .A(\AES_ENC/w2[21] ), .B(\AES_ENC/sa02_sub[5] ),.Z(\AES_ENC/n1006 ) );
XOR2_X2 \AES_ENC/U1277  ( .A(\AES_ENC/sa13_sub[7] ), .B(\AES_ENC/sa20_sub[7] ), .Z(\AES_ENC/n1195 ) );
XOR2_X2 \AES_ENC/U1276  ( .A(\AES_ENC/n1008 ), .B(\AES_ENC/n1007 ), .Z(\AES_ENC/sa12_next [4]) );
XOR2_X2 \AES_ENC/U1275  ( .A(\AES_ENC/n1010 ), .B(\AES_ENC/n1009 ), .Z(\AES_ENC/n1007 ) );
XOR2_X2 \AES_ENC/U1274  ( .A(\AES_ENC/n1195 ), .B(\AES_ENC/n1198 ), .Z(\AES_ENC/n1008 ) );
XOR2_X2 \AES_ENC/U1273  ( .A(\AES_ENC/sa13_sub[3] ), .B(\AES_ENC/sa20_sub[3] ), .Z(\AES_ENC/n1009 ) );
XOR2_X2 \AES_ENC/U1272  ( .A(\AES_ENC/w2[20] ), .B(\AES_ENC/sa02_sub[4] ),.Z(\AES_ENC/n1010 ) );
XOR2_X2 \AES_ENC/U1271  ( .A(\AES_ENC/n1012 ), .B(\AES_ENC/n1011 ), .Z(\AES_ENC/sa12_next [3]) );
XOR2_X2 \AES_ENC/U1270  ( .A(\AES_ENC/n1014 ), .B(\AES_ENC/n1013 ), .Z(\AES_ENC/n1011 ) );
XOR2_X2 \AES_ENC/U1269  ( .A(\AES_ENC/n1195 ), .B(\AES_ENC/n1199 ), .Z(\AES_ENC/n1012 ) );
XOR2_X2 \AES_ENC/U1268  ( .A(\AES_ENC/sa13_sub[2] ), .B(\AES_ENC/sa20_sub[2] ), .Z(\AES_ENC/n1013 ) );
XOR2_X2 \AES_ENC/U1267  ( .A(\AES_ENC/w2[19] ), .B(\AES_ENC/sa02_sub[3] ),.Z(\AES_ENC/n1014 ) );
XOR2_X2 \AES_ENC/U1266  ( .A(\AES_ENC/n1016 ), .B(\AES_ENC/n1015 ), .Z(\AES_ENC/sa12_next [2]) );
XOR2_X2 \AES_ENC/U1265  ( .A(\AES_ENC/n1200 ), .B(\AES_ENC/n1017 ), .Z(\AES_ENC/n1015 ) );
XOR2_X2 \AES_ENC/U1264  ( .A(\AES_ENC/sa13_sub[1] ), .B(\AES_ENC/sa20_sub[1] ), .Z(\AES_ENC/n1016 ) );
XOR2_X2 \AES_ENC/U1263  ( .A(\AES_ENC/w2[18] ), .B(\AES_ENC/sa02_sub[2] ),.Z(\AES_ENC/n1017 ) );
XOR2_X2 \AES_ENC/U1262  ( .A(\AES_ENC/n1019 ), .B(\AES_ENC/n1018 ), .Z(\AES_ENC/sa12_next [1]) );
XOR2_X2 \AES_ENC/U1261  ( .A(\AES_ENC/n1021 ), .B(\AES_ENC/n1020 ), .Z(\AES_ENC/n1018 ) );
XOR2_X2 \AES_ENC/U1260  ( .A(\AES_ENC/n1195 ), .B(\AES_ENC/n1201 ), .Z(\AES_ENC/n1019 ) );
XOR2_X2 \AES_ENC/U1259  ( .A(\AES_ENC/sa13_sub[0] ), .B(\AES_ENC/sa20_sub[0] ), .Z(\AES_ENC/n1020 ) );
XOR2_X2 \AES_ENC/U1258  ( .A(\AES_ENC/w2[17] ), .B(\AES_ENC/sa02_sub[1] ),.Z(\AES_ENC/n1021 ) );
XOR2_X2 \AES_ENC/U1257  ( .A(\AES_ENC/n1023 ), .B(\AES_ENC/n1022 ), .Z(\AES_ENC/sa12_next [0]) );
XOR2_X2 \AES_ENC/U1256  ( .A(\AES_ENC/n1195 ), .B(\AES_ENC/n1202 ), .Z(\AES_ENC/n1022 ) );
XOR2_X2 \AES_ENC/U1255  ( .A(\AES_ENC/w2[16] ), .B(\AES_ENC/sa02_sub[0] ),.Z(\AES_ENC/n1023 ) );
XOR2_X2 \AES_ENC/U1254  ( .A(\AES_ENC/n1025 ), .B(\AES_ENC/n1024 ), .Z(\AES_ENC/sa22_next [7]) );
XOR2_X2 \AES_ENC/U1253  ( .A(\AES_ENC/n1204 ), .B(\AES_ENC/n1196 ), .Z(\AES_ENC/n1024 ) );
XOR2_X2 \AES_ENC/U1252  ( .A(\AES_ENC/w2[15] ), .B(\AES_ENC/sa31_sub[7] ),.Z(\AES_ENC/n1025 ) );
XOR2_X2 \AES_ENC/U1251  ( .A(\AES_ENC/n1027 ), .B(\AES_ENC/n1026 ), .Z(\AES_ENC/sa22_next [6]) );
XOR2_X2 \AES_ENC/U1250  ( .A(\AES_ENC/n1205 ), .B(\AES_ENC/n1197 ), .Z(\AES_ENC/n1026 ) );
XOR2_X2 \AES_ENC/U1249  ( .A(\AES_ENC/w2[14] ), .B(\AES_ENC/sa31_sub[6] ),.Z(\AES_ENC/n1027 ) );
XOR2_X2 \AES_ENC/U1248  ( .A(\AES_ENC/n1029 ), .B(\AES_ENC/n1028 ), .Z(\AES_ENC/sa22_next [5]) );
XOR2_X2 \AES_ENC/U1247  ( .A(\AES_ENC/n1206 ), .B(\AES_ENC/n1198 ), .Z(\AES_ENC/n1028 ) );
XOR2_X2 \AES_ENC/U1246  ( .A(\AES_ENC/w2[13] ), .B(\AES_ENC/sa31_sub[5] ),.Z(\AES_ENC/n1029 ) );
XOR2_X2 \AES_ENC/U1245  ( .A(\AES_ENC/n1031 ), .B(\AES_ENC/n1030 ), .Z(\AES_ENC/sa22_next [4]) );
XOR2_X2 \AES_ENC/U1244  ( .A(\AES_ENC/n1199 ), .B(\AES_ENC/n1032 ), .Z(\AES_ENC/n1030 ) );
XOR2_X2 \AES_ENC/U1243  ( .A(\AES_ENC/n1203 ), .B(\AES_ENC/n1207 ), .Z(\AES_ENC/n1031 ) );
XOR2_X2 \AES_ENC/U1242  ( .A(\AES_ENC/w2[12] ), .B(\AES_ENC/sa31_sub[4] ),.Z(\AES_ENC/n1032 ) );
XOR2_X2 \AES_ENC/U1241  ( .A(\AES_ENC/n1034 ), .B(\AES_ENC/n1033 ), .Z(\AES_ENC/sa22_next [3]) );
XOR2_X2 \AES_ENC/U1240  ( .A(\AES_ENC/n1200 ), .B(\AES_ENC/n1035 ), .Z(\AES_ENC/n1033 ) );
XOR2_X2 \AES_ENC/U1239  ( .A(\AES_ENC/n1203 ), .B(\AES_ENC/n1208 ), .Z(\AES_ENC/n1034 ) );
XOR2_X2 \AES_ENC/U1238  ( .A(\AES_ENC/w2[11] ), .B(\AES_ENC/sa31_sub[3] ),.Z(\AES_ENC/n1035 ) );
XOR2_X2 \AES_ENC/U1237  ( .A(\AES_ENC/n1037 ), .B(\AES_ENC/n1036 ), .Z(\AES_ENC/sa22_next [2]) );
XOR2_X2 \AES_ENC/U1236  ( .A(\AES_ENC/n1209 ), .B(\AES_ENC/n1201 ), .Z(\AES_ENC/n1036 ) );
XOR2_X2 \AES_ENC/U1235  ( .A(\AES_ENC/w2[10] ), .B(\AES_ENC/sa31_sub[2] ),.Z(\AES_ENC/n1037 ) );
XOR2_X2 \AES_ENC/U1234  ( .A(\AES_ENC/n1039 ), .B(\AES_ENC/n1038 ), .Z(\AES_ENC/sa22_next [1]) );
XOR2_X2 \AES_ENC/U1233  ( .A(\AES_ENC/n1202 ), .B(\AES_ENC/n1040 ), .Z(\AES_ENC/n1038 ) );
XOR2_X2 \AES_ENC/U1232  ( .A(\AES_ENC/n1203 ), .B(\AES_ENC/n1210 ), .Z(\AES_ENC/n1039 ) );
XOR2_X2 \AES_ENC/U1231  ( .A(\AES_ENC/w2[9] ), .B(\AES_ENC/sa31_sub[1] ),.Z(\AES_ENC/n1040 ) );
XOR2_X2 \AES_ENC/U1230  ( .A(\AES_ENC/n1042 ), .B(\AES_ENC/n1041 ), .Z(\AES_ENC/sa22_next [0]) );
XOR2_X2 \AES_ENC/U1229  ( .A(\AES_ENC/n1203 ), .B(\AES_ENC/n1211 ), .Z(\AES_ENC/n1041 ) );
XOR2_X2 \AES_ENC/U1228  ( .A(\AES_ENC/w2[8] ), .B(\AES_ENC/sa31_sub[0] ),.Z(\AES_ENC/n1042 ) );
XOR2_X2 \AES_ENC/U1227  ( .A(\AES_ENC/n1044 ), .B(\AES_ENC/n1043 ), .Z(\AES_ENC/sa32_next [7]) );
XOR2_X2 \AES_ENC/U1226  ( .A(\AES_ENC/n1204 ), .B(\AES_ENC/n1045 ), .Z(\AES_ENC/n1043 ) );
XOR2_X2 \AES_ENC/U1225  ( .A(\AES_ENC/sa20_sub[7] ), .B(\AES_ENC/sa31_sub[6] ), .Z(\AES_ENC/n1044 ) );
XOR2_X2 \AES_ENC/U1224  ( .A(\AES_ENC/w2[7] ), .B(\AES_ENC/sa02_sub[6] ),.Z(\AES_ENC/n1045 ) );
XOR2_X2 \AES_ENC/U1223  ( .A(\AES_ENC/n1047 ), .B(\AES_ENC/n1046 ), .Z(\AES_ENC/sa32_next [6]) );
XOR2_X2 \AES_ENC/U1222  ( .A(\AES_ENC/n1205 ), .B(\AES_ENC/n1048 ), .Z(\AES_ENC/n1046 ) );
XOR2_X2 \AES_ENC/U1221  ( .A(\AES_ENC/sa20_sub[6] ), .B(\AES_ENC/sa31_sub[5] ), .Z(\AES_ENC/n1047 ) );
XOR2_X2 \AES_ENC/U1220  ( .A(\AES_ENC/w2[6] ), .B(\AES_ENC/sa02_sub[5] ),.Z(\AES_ENC/n1048 ) );
XOR2_X2 \AES_ENC/U1219  ( .A(\AES_ENC/n1050 ), .B(\AES_ENC/n1049 ), .Z(\AES_ENC/sa32_next [5]) );
XOR2_X2 \AES_ENC/U1218  ( .A(\AES_ENC/n1206 ), .B(\AES_ENC/n1051 ), .Z(\AES_ENC/n1049 ) );
XOR2_X2 \AES_ENC/U1217  ( .A(\AES_ENC/sa20_sub[5] ), .B(\AES_ENC/sa31_sub[4] ), .Z(\AES_ENC/n1050 ) );
XOR2_X2 \AES_ENC/U1216  ( .A(\AES_ENC/w2[5] ), .B(\AES_ENC/sa02_sub[4] ),.Z(\AES_ENC/n1051 ) );
XOR2_X2 \AES_ENC/U1215  ( .A(\AES_ENC/sa02_sub[7] ), .B(\AES_ENC/sa31_sub[7] ), .Z(\AES_ENC/n1212 ) );
XOR2_X2 \AES_ENC/U1214  ( .A(\AES_ENC/n1053 ), .B(\AES_ENC/n1052 ), .Z(\AES_ENC/sa32_next [4]) );
XOR2_X2 \AES_ENC/U1213  ( .A(\AES_ENC/n1055 ), .B(\AES_ENC/n1054 ), .Z(\AES_ENC/n1052 ) );
XOR2_X2 \AES_ENC/U1212  ( .A(\AES_ENC/n1212 ), .B(\AES_ENC/n1207 ), .Z(\AES_ENC/n1053 ) );
XOR2_X2 \AES_ENC/U1211  ( .A(\AES_ENC/sa20_sub[4] ), .B(\AES_ENC/sa31_sub[3] ), .Z(\AES_ENC/n1054 ) );
XOR2_X2 \AES_ENC/U1210  ( .A(\AES_ENC/w2[4] ), .B(\AES_ENC/sa02_sub[3] ),.Z(\AES_ENC/n1055 ) );
XOR2_X2 \AES_ENC/U1209  ( .A(\AES_ENC/n1057 ), .B(\AES_ENC/n1056 ), .Z(\AES_ENC/sa32_next [3]) );
XOR2_X2 \AES_ENC/U1208  ( .A(\AES_ENC/n1059 ), .B(\AES_ENC/n1058 ), .Z(\AES_ENC/n1056 ) );
XOR2_X2 \AES_ENC/U1207  ( .A(\AES_ENC/n1212 ), .B(\AES_ENC/n1208 ), .Z(\AES_ENC/n1057 ) );
XOR2_X2 \AES_ENC/U1206  ( .A(\AES_ENC/sa20_sub[3] ), .B(\AES_ENC/sa31_sub[2] ), .Z(\AES_ENC/n1058 ) );
XOR2_X2 \AES_ENC/U1205  ( .A(\AES_ENC/w2[3] ), .B(\AES_ENC/sa02_sub[2] ),.Z(\AES_ENC/n1059 ) );
XOR2_X2 \AES_ENC/U1204  ( .A(\AES_ENC/n1061 ), .B(\AES_ENC/n1060 ), .Z(\AES_ENC/sa32_next [2]) );
XOR2_X2 \AES_ENC/U1203  ( .A(\AES_ENC/n1209 ), .B(\AES_ENC/n1062 ), .Z(\AES_ENC/n1060 ) );
XOR2_X2 \AES_ENC/U1202  ( .A(\AES_ENC/sa20_sub[2] ), .B(\AES_ENC/sa31_sub[1] ), .Z(\AES_ENC/n1061 ) );
XOR2_X2 \AES_ENC/U1201  ( .A(\AES_ENC/w2[2] ), .B(\AES_ENC/sa02_sub[1] ),.Z(\AES_ENC/n1062 ) );
XOR2_X2 \AES_ENC/U1200  ( .A(\AES_ENC/n1064 ), .B(\AES_ENC/n1063 ), .Z(\AES_ENC/sa32_next [1]) );
XOR2_X2 \AES_ENC/U1199  ( .A(\AES_ENC/n1066 ), .B(\AES_ENC/n1065 ), .Z(\AES_ENC/n1063 ) );
XOR2_X2 \AES_ENC/U1198  ( .A(\AES_ENC/n1212 ), .B(\AES_ENC/n1210 ), .Z(\AES_ENC/n1064 ) );
XOR2_X2 \AES_ENC/U1197  ( .A(\AES_ENC/sa20_sub[1] ), .B(\AES_ENC/sa31_sub[0] ), .Z(\AES_ENC/n1065 ) );
XOR2_X2 \AES_ENC/U1196  ( .A(\AES_ENC/w2[1] ), .B(\AES_ENC/sa02_sub[0] ),.Z(\AES_ENC/n1066 ) );
XOR2_X2 \AES_ENC/U1195  ( .A(\AES_ENC/n1068 ), .B(\AES_ENC/n1067 ), .Z(\AES_ENC/sa32_next [0]) );
XOR2_X2 \AES_ENC/U1194  ( .A(\AES_ENC/n1212 ), .B(\AES_ENC/n1211 ), .Z(\AES_ENC/n1067 ) );
XOR2_X2 \AES_ENC/U1193  ( .A(\AES_ENC/w2[0] ), .B(\AES_ENC/sa20_sub[0] ),.Z(\AES_ENC/n1068 ) );
XOR2_X2 \AES_ENC/U1192  ( .A(\AES_ENC/sa21_sub[7] ), .B(\AES_ENC/sa32_sub[7] ), .Z(\AES_ENC/n1221 ) );
XOR2_X2 \AES_ENC/U1191  ( .A(\AES_ENC/sa03_sub[6] ), .B(\AES_ENC/sa10_sub[6] ), .Z(\AES_ENC/n1223 ) );
XOR2_X2 \AES_ENC/U1190  ( .A(\AES_ENC/n1070 ), .B(\AES_ENC/n1069 ), .Z(\AES_ENC/sa03_next [7]) );
XOR2_X2 \AES_ENC/U1189  ( .A(\AES_ENC/n1221 ), .B(\AES_ENC/n1223 ), .Z(\AES_ENC/n1069 ) );
XOR2_X2 \AES_ENC/U1188  ( .A(\AES_ENC/w3[31] ), .B(\AES_ENC/sa10_sub[7] ),.Z(\AES_ENC/n1070 ) );
XOR2_X2 \AES_ENC/U1187  ( .A(\AES_ENC/sa03_sub[5] ), .B(\AES_ENC/sa10_sub[5] ), .Z(\AES_ENC/n1224 ) );
XOR2_X2 \AES_ENC/U1186  ( .A(\AES_ENC/sa21_sub[6] ), .B(\AES_ENC/sa32_sub[6] ), .Z(\AES_ENC/n1214 ) );
XOR2_X2 \AES_ENC/U1185  ( .A(\AES_ENC/n1072 ), .B(\AES_ENC/n1071 ), .Z(\AES_ENC/sa03_next [6]) );
XOR2_X2 \AES_ENC/U1184  ( .A(\AES_ENC/n1224 ), .B(\AES_ENC/n1214 ), .Z(\AES_ENC/n1071 ) );
XOR2_X2 \AES_ENC/U1183  ( .A(\AES_ENC/w3[30] ), .B(\AES_ENC/sa10_sub[6] ),.Z(\AES_ENC/n1072 ) );
XOR2_X2 \AES_ENC/U1182  ( .A(\AES_ENC/sa03_sub[4] ), .B(\AES_ENC/sa10_sub[4] ), .Z(\AES_ENC/n1225 ) );
XOR2_X2 \AES_ENC/U1181  ( .A(\AES_ENC/sa21_sub[5] ), .B(\AES_ENC/sa32_sub[5] ), .Z(\AES_ENC/n1215 ) );
XOR2_X2 \AES_ENC/U1180  ( .A(\AES_ENC/n1074 ), .B(\AES_ENC/n1073 ), .Z(\AES_ENC/sa03_next [5]) );
XOR2_X2 \AES_ENC/U1179  ( .A(\AES_ENC/n1225 ), .B(\AES_ENC/n1215 ), .Z(\AES_ENC/n1073 ) );
XOR2_X2 \AES_ENC/U1178  ( .A(\AES_ENC/w3[29] ), .B(\AES_ENC/sa10_sub[5] ),.Z(\AES_ENC/n1074 ) );
XOR2_X2 \AES_ENC/U1177  ( .A(\AES_ENC/sa03_sub[7] ), .B(\AES_ENC/sa10_sub[7] ), .Z(\AES_ENC/n1222 ) );
XOR2_X2 \AES_ENC/U1176  ( .A(\AES_ENC/sa03_sub[3] ), .B(\AES_ENC/sa10_sub[3] ), .Z(\AES_ENC/n1226 ) );
XOR2_X2 \AES_ENC/U1175  ( .A(\AES_ENC/sa21_sub[4] ), .B(\AES_ENC/sa32_sub[4] ), .Z(\AES_ENC/n1216 ) );
XOR2_X2 \AES_ENC/U1174  ( .A(\AES_ENC/n1076 ), .B(\AES_ENC/n1075 ), .Z(\AES_ENC/sa03_next [4]) );
XOR2_X2 \AES_ENC/U1173  ( .A(\AES_ENC/n1216 ), .B(\AES_ENC/n1077 ), .Z(\AES_ENC/n1075 ) );
XOR2_X2 \AES_ENC/U1172  ( .A(\AES_ENC/n1222 ), .B(\AES_ENC/n1226 ), .Z(\AES_ENC/n1076 ) );
XOR2_X2 \AES_ENC/U1171  ( .A(\AES_ENC/w3[28] ), .B(\AES_ENC/sa10_sub[4] ),.Z(\AES_ENC/n1077 ) );
XOR2_X2 \AES_ENC/U1170  ( .A(\AES_ENC/sa03_sub[2] ), .B(\AES_ENC/sa10_sub[2] ), .Z(\AES_ENC/n1227 ) );
XOR2_X2 \AES_ENC/U1169  ( .A(\AES_ENC/sa21_sub[3] ), .B(\AES_ENC/sa32_sub[3] ), .Z(\AES_ENC/n1217 ) );
XOR2_X2 \AES_ENC/U1168  ( .A(\AES_ENC/n1079 ), .B(\AES_ENC/n1078 ), .Z(\AES_ENC/sa03_next [3]) );
XOR2_X2 \AES_ENC/U1167  ( .A(\AES_ENC/n1217 ), .B(\AES_ENC/n1080 ), .Z(\AES_ENC/n1078 ) );
XOR2_X2 \AES_ENC/U1166  ( .A(\AES_ENC/n1222 ), .B(\AES_ENC/n1227 ), .Z(\AES_ENC/n1079 ) );
XOR2_X2 \AES_ENC/U1165  ( .A(\AES_ENC/w3[27] ), .B(\AES_ENC/sa10_sub[3] ),.Z(\AES_ENC/n1080 ) );
XOR2_X2 \AES_ENC/U1164  ( .A(\AES_ENC/sa03_sub[1] ), .B(\AES_ENC/sa10_sub[1] ), .Z(\AES_ENC/n1228 ) );
XOR2_X2 \AES_ENC/U1163  ( .A(\AES_ENC/sa21_sub[2] ), .B(\AES_ENC/sa32_sub[2] ), .Z(\AES_ENC/n1218 ) );
XOR2_X2 \AES_ENC/U1162  ( .A(\AES_ENC/n1082 ), .B(\AES_ENC/n1081 ), .Z(\AES_ENC/sa03_next [2]) );
XOR2_X2 \AES_ENC/U1161  ( .A(\AES_ENC/n1228 ), .B(\AES_ENC/n1218 ), .Z(\AES_ENC/n1081 ) );
XOR2_X2 \AES_ENC/U1160  ( .A(\AES_ENC/w3[26] ), .B(\AES_ENC/sa10_sub[2] ),.Z(\AES_ENC/n1082 ) );
XOR2_X2 \AES_ENC/U1159  ( .A(\AES_ENC/sa03_sub[0] ), .B(\AES_ENC/sa10_sub[0] ), .Z(\AES_ENC/n1229 ) );
XOR2_X2 \AES_ENC/U1158  ( .A(\AES_ENC/sa21_sub[1] ), .B(\AES_ENC/sa32_sub[1] ), .Z(\AES_ENC/n1219 ) );
XOR2_X2 \AES_ENC/U1157  ( .A(\AES_ENC/n1084 ), .B(\AES_ENC/n1083 ), .Z(\AES_ENC/sa03_next [1]) );
XOR2_X2 \AES_ENC/U1156  ( .A(\AES_ENC/n1219 ), .B(\AES_ENC/n1085 ), .Z(\AES_ENC/n1083 ) );
XOR2_X2 \AES_ENC/U1155  ( .A(\AES_ENC/n1222 ), .B(\AES_ENC/n1229 ), .Z(\AES_ENC/n1084 ) );
XOR2_X2 \AES_ENC/U1154  ( .A(\AES_ENC/w3[25] ), .B(\AES_ENC/sa10_sub[1] ),.Z(\AES_ENC/n1085 ) );
XOR2_X2 \AES_ENC/U1153  ( .A(\AES_ENC/sa21_sub[0] ), .B(\AES_ENC/sa32_sub[0] ), .Z(\AES_ENC/n1220 ) );
XOR2_X2 \AES_ENC/U1152  ( .A(\AES_ENC/n1087 ), .B(\AES_ENC/n1086 ), .Z(\AES_ENC/sa03_next [0]) );
XOR2_X2 \AES_ENC/U1151  ( .A(\AES_ENC/n1222 ), .B(\AES_ENC/n1220 ), .Z(\AES_ENC/n1086 ) );
XOR2_X2 \AES_ENC/U1150  ( .A(\AES_ENC/w3[24] ), .B(\AES_ENC/sa10_sub[0] ),.Z(\AES_ENC/n1087 ) );
XOR2_X2 \AES_ENC/U1149  ( .A(\AES_ENC/n1089 ), .B(\AES_ENC/n1088 ), .Z(\AES_ENC/sa13_next [7]) );
XOR2_X2 \AES_ENC/U1148  ( .A(\AES_ENC/n1221 ), .B(\AES_ENC/n1090 ), .Z(\AES_ENC/n1088 ) );
XOR2_X2 \AES_ENC/U1147  ( .A(\AES_ENC/sa10_sub[6] ), .B(\AES_ENC/sa21_sub[6] ), .Z(\AES_ENC/n1089 ) );
XOR2_X2 \AES_ENC/U1146  ( .A(\AES_ENC/w3[23] ), .B(\AES_ENC/sa03_sub[7] ),.Z(\AES_ENC/n1090 ) );
XOR2_X2 \AES_ENC/U1145  ( .A(\AES_ENC/n1092 ), .B(\AES_ENC/n1091 ), .Z(\AES_ENC/sa13_next [6]) );
XOR2_X2 \AES_ENC/U1144  ( .A(\AES_ENC/n1214 ), .B(\AES_ENC/n1093 ), .Z(\AES_ENC/n1091 ) );
XOR2_X2 \AES_ENC/U1143  ( .A(\AES_ENC/sa10_sub[5] ), .B(\AES_ENC/sa21_sub[5] ), .Z(\AES_ENC/n1092 ) );
XOR2_X2 \AES_ENC/U1142  ( .A(\AES_ENC/w3[22] ), .B(\AES_ENC/sa03_sub[6] ),.Z(\AES_ENC/n1093 ) );
XOR2_X2 \AES_ENC/U1141  ( .A(\AES_ENC/n1095 ), .B(\AES_ENC/n1094 ), .Z(\AES_ENC/sa13_next [5]) );
XOR2_X2 \AES_ENC/U1140  ( .A(\AES_ENC/n1215 ), .B(\AES_ENC/n1096 ), .Z(\AES_ENC/n1094 ) );
XOR2_X2 \AES_ENC/U1139  ( .A(\AES_ENC/sa10_sub[4] ), .B(\AES_ENC/sa21_sub[4] ), .Z(\AES_ENC/n1095 ) );
XOR2_X2 \AES_ENC/U1138  ( .A(\AES_ENC/w3[21] ), .B(\AES_ENC/sa03_sub[5] ),.Z(\AES_ENC/n1096 ) );
XOR2_X2 \AES_ENC/U1137  ( .A(\AES_ENC/sa10_sub[7] ), .B(\AES_ENC/sa21_sub[7] ), .Z(\AES_ENC/n1213 ) );
XOR2_X2 \AES_ENC/U1136  ( .A(\AES_ENC/n1098 ), .B(\AES_ENC/n1097 ), .Z(\AES_ENC/sa13_next [4]) );
XOR2_X2 \AES_ENC/U1135  ( .A(\AES_ENC/n1100 ), .B(\AES_ENC/n1099 ), .Z(\AES_ENC/n1097 ) );
XOR2_X2 \AES_ENC/U1134  ( .A(\AES_ENC/n1213 ), .B(\AES_ENC/n1216 ), .Z(\AES_ENC/n1098 ) );
XOR2_X2 \AES_ENC/U1133  ( .A(\AES_ENC/sa10_sub[3] ), .B(\AES_ENC/sa21_sub[3] ), .Z(\AES_ENC/n1099 ) );
XOR2_X2 \AES_ENC/U1132  ( .A(\AES_ENC/w3[20] ), .B(\AES_ENC/sa03_sub[4] ),.Z(\AES_ENC/n1100 ) );
XOR2_X2 \AES_ENC/U1131  ( .A(\AES_ENC/n1102 ), .B(\AES_ENC/n1101 ), .Z(\AES_ENC/sa13_next [3]) );
XOR2_X2 \AES_ENC/U1130  ( .A(\AES_ENC/n1104 ), .B(\AES_ENC/n1103 ), .Z(\AES_ENC/n1101 ) );
XOR2_X2 \AES_ENC/U1129  ( .A(\AES_ENC/n1213 ), .B(\AES_ENC/n1217 ), .Z(\AES_ENC/n1102 ) );
XOR2_X2 \AES_ENC/U1128  ( .A(\AES_ENC/sa10_sub[2] ), .B(\AES_ENC/sa21_sub[2] ), .Z(\AES_ENC/n1103 ) );
XOR2_X2 \AES_ENC/U1127  ( .A(\AES_ENC/w3[19] ), .B(\AES_ENC/sa03_sub[3] ),.Z(\AES_ENC/n1104 ) );
XOR2_X2 \AES_ENC/U1126  ( .A(\AES_ENC/n1106 ), .B(\AES_ENC/n1105 ), .Z(\AES_ENC/sa13_next [2]) );
XOR2_X2 \AES_ENC/U1125  ( .A(\AES_ENC/n1218 ), .B(\AES_ENC/n1107 ), .Z(\AES_ENC/n1105 ) );
XOR2_X2 \AES_ENC/U1124  ( .A(\AES_ENC/sa10_sub[1] ), .B(\AES_ENC/sa21_sub[1] ), .Z(\AES_ENC/n1106 ) );
XOR2_X2 \AES_ENC/U1123  ( .A(\AES_ENC/w3[18] ), .B(\AES_ENC/sa03_sub[2] ),.Z(\AES_ENC/n1107 ) );
XOR2_X2 \AES_ENC/U1122  ( .A(\AES_ENC/n1109 ), .B(\AES_ENC/n1108 ), .Z(\AES_ENC/sa13_next [1]) );
XOR2_X2 \AES_ENC/U1121  ( .A(\AES_ENC/n1111 ), .B(\AES_ENC/n1110 ), .Z(\AES_ENC/n1108 ) );
XOR2_X2 \AES_ENC/U1120  ( .A(\AES_ENC/n1213 ), .B(\AES_ENC/n1219 ), .Z(\AES_ENC/n1109 ) );
XOR2_X2 \AES_ENC/U1119  ( .A(\AES_ENC/sa10_sub[0] ), .B(\AES_ENC/sa21_sub[0] ), .Z(\AES_ENC/n1110 ) );
XOR2_X2 \AES_ENC/U1118  ( .A(\AES_ENC/w3[17] ), .B(\AES_ENC/sa03_sub[1] ),.Z(\AES_ENC/n1111 ) );
XOR2_X2 \AES_ENC/U1117  ( .A(\AES_ENC/n1113 ), .B(\AES_ENC/n1112 ), .Z(\AES_ENC/sa13_next [0]) );
XOR2_X2 \AES_ENC/U1116  ( .A(\AES_ENC/n1213 ), .B(\AES_ENC/n1220 ), .Z(\AES_ENC/n1112 ) );
XOR2_X2 \AES_ENC/U1115  ( .A(\AES_ENC/w3[16] ), .B(\AES_ENC/sa03_sub[0] ),.Z(\AES_ENC/n1113 ) );
XOR2_X2 \AES_ENC/U1114  ( .A(\AES_ENC/n1115 ), .B(\AES_ENC/n1114 ), .Z(\AES_ENC/sa23_next [7]) );
XOR2_X2 \AES_ENC/U1113  ( .A(\AES_ENC/n1222 ), .B(\AES_ENC/n1214 ), .Z(\AES_ENC/n1114 ) );
XOR2_X2 \AES_ENC/U1112  ( .A(\AES_ENC/w3[15] ), .B(\AES_ENC/sa32_sub[7] ),.Z(\AES_ENC/n1115 ) );
XOR2_X2 \AES_ENC/U1111  ( .A(\AES_ENC/n1117 ), .B(\AES_ENC/n1116 ), .Z(\AES_ENC/sa23_next [6]) );
XOR2_X2 \AES_ENC/U1110  ( .A(\AES_ENC/n1223 ), .B(\AES_ENC/n1215 ), .Z(\AES_ENC/n1116 ) );
XOR2_X2 \AES_ENC/U1109  ( .A(\AES_ENC/w3[14] ), .B(\AES_ENC/sa32_sub[6] ),.Z(\AES_ENC/n1117 ) );
XOR2_X2 \AES_ENC/U1108  ( .A(\AES_ENC/n1119 ), .B(\AES_ENC/n1118 ), .Z(\AES_ENC/sa23_next [5]) );
XOR2_X2 \AES_ENC/U1107  ( .A(\AES_ENC/n1224 ), .B(\AES_ENC/n1216 ), .Z(\AES_ENC/n1118 ) );
XOR2_X2 \AES_ENC/U1106  ( .A(\AES_ENC/w3[13] ), .B(\AES_ENC/sa32_sub[5] ),.Z(\AES_ENC/n1119 ) );
XOR2_X2 \AES_ENC/U1105  ( .A(\AES_ENC/n1121 ), .B(\AES_ENC/n1120 ), .Z(\AES_ENC/sa23_next [4]) );
XOR2_X2 \AES_ENC/U1104  ( .A(\AES_ENC/n1217 ), .B(\AES_ENC/n1122 ), .Z(\AES_ENC/n1120 ) );
XOR2_X2 \AES_ENC/U1103  ( .A(\AES_ENC/n1221 ), .B(\AES_ENC/n1225 ), .Z(\AES_ENC/n1121 ) );
XOR2_X2 \AES_ENC/U1102  ( .A(\AES_ENC/w3[12] ), .B(\AES_ENC/sa32_sub[4] ),.Z(\AES_ENC/n1122 ) );
XOR2_X2 \AES_ENC/U1101  ( .A(\AES_ENC/n1124 ), .B(\AES_ENC/n1123 ), .Z(\AES_ENC/sa23_next [3]) );
XOR2_X2 \AES_ENC/U1100  ( .A(\AES_ENC/n1218 ), .B(\AES_ENC/n1125 ), .Z(\AES_ENC/n1123 ) );
XOR2_X2 \AES_ENC/U1099  ( .A(\AES_ENC/n1221 ), .B(\AES_ENC/n1226 ), .Z(\AES_ENC/n1124 ) );
XOR2_X2 \AES_ENC/U1098  ( .A(\AES_ENC/w3[11] ), .B(\AES_ENC/sa32_sub[3] ),.Z(\AES_ENC/n1125 ) );
XOR2_X2 \AES_ENC/U1097  ( .A(\AES_ENC/n1127 ), .B(\AES_ENC/n1126 ), .Z(\AES_ENC/sa23_next [2]) );
XOR2_X2 \AES_ENC/U1096  ( .A(\AES_ENC/n1227 ), .B(\AES_ENC/n1219 ), .Z(\AES_ENC/n1126 ) );
XOR2_X2 \AES_ENC/U1095  ( .A(\AES_ENC/w3[10] ), .B(\AES_ENC/sa32_sub[2] ),.Z(\AES_ENC/n1127 ) );
XOR2_X2 \AES_ENC/U1094  ( .A(\AES_ENC/n1129 ), .B(\AES_ENC/n1128 ), .Z(\AES_ENC/sa23_next [1]) );
XOR2_X2 \AES_ENC/U1093  ( .A(\AES_ENC/n1220 ), .B(\AES_ENC/n1130 ), .Z(\AES_ENC/n1128 ) );
XOR2_X2 \AES_ENC/U1092  ( .A(\AES_ENC/n1221 ), .B(\AES_ENC/n1228 ), .Z(\AES_ENC/n1129 ) );
XOR2_X2 \AES_ENC/U1091  ( .A(\AES_ENC/w3[9] ), .B(\AES_ENC/sa32_sub[1] ),.Z(\AES_ENC/n1130 ) );
XOR2_X2 \AES_ENC/U1090  ( .A(\AES_ENC/n1132 ), .B(\AES_ENC/n1131 ), .Z(\AES_ENC/sa23_next [0]) );
XOR2_X2 \AES_ENC/U1089  ( .A(\AES_ENC/n1221 ), .B(\AES_ENC/n1229 ), .Z(\AES_ENC/n1131 ) );
XOR2_X2 \AES_ENC/U1088  ( .A(\AES_ENC/w3[8] ), .B(\AES_ENC/sa32_sub[0] ),.Z(\AES_ENC/n1132 ) );
XOR2_X2 \AES_ENC/U1087  ( .A(\AES_ENC/n1134 ), .B(\AES_ENC/n1133 ), .Z(\AES_ENC/sa33_next [7]) );
XOR2_X2 \AES_ENC/U1086  ( .A(\AES_ENC/n1222 ), .B(\AES_ENC/n1135 ), .Z(\AES_ENC/n1133 ) );
XOR2_X2 \AES_ENC/U1085  ( .A(\AES_ENC/sa21_sub[7] ), .B(\AES_ENC/sa32_sub[6] ), .Z(\AES_ENC/n1134 ) );
XOR2_X2 \AES_ENC/U1084  ( .A(\AES_ENC/w3[7] ), .B(\AES_ENC/sa03_sub[6] ),.Z(\AES_ENC/n1135 ) );
XOR2_X2 \AES_ENC/U1083  ( .A(\AES_ENC/n1137 ), .B(\AES_ENC/n1136 ), .Z(\AES_ENC/sa33_next [6]) );
XOR2_X2 \AES_ENC/U1082  ( .A(\AES_ENC/n1223 ), .B(\AES_ENC/n1138 ), .Z(\AES_ENC/n1136 ) );
XOR2_X2 \AES_ENC/U1081  ( .A(\AES_ENC/sa21_sub[6] ), .B(\AES_ENC/sa32_sub[5] ), .Z(\AES_ENC/n1137 ) );
XOR2_X2 \AES_ENC/U1080  ( .A(\AES_ENC/w3[6] ), .B(\AES_ENC/sa03_sub[5] ),.Z(\AES_ENC/n1138 ) );
XOR2_X2 \AES_ENC/U1079  ( .A(\AES_ENC/n1140 ), .B(\AES_ENC/n1139 ), .Z(\AES_ENC/sa33_next [5]) );
XOR2_X2 \AES_ENC/U1078  ( .A(\AES_ENC/n1224 ), .B(\AES_ENC/n1141 ), .Z(\AES_ENC/n1139 ) );
XOR2_X2 \AES_ENC/U1077  ( .A(\AES_ENC/sa21_sub[5] ), .B(\AES_ENC/sa32_sub[4] ), .Z(\AES_ENC/n1140 ) );
XOR2_X2 \AES_ENC/U1076  ( .A(\AES_ENC/w3[5] ), .B(\AES_ENC/sa03_sub[4] ),.Z(\AES_ENC/n1141 ) );
XOR2_X2 \AES_ENC/U1075  ( .A(\AES_ENC/sa03_sub[7] ), .B(\AES_ENC/sa32_sub[7] ), .Z(\AES_ENC/n1230 ) );
XOR2_X2 \AES_ENC/U1074  ( .A(\AES_ENC/n1143 ), .B(\AES_ENC/n1142 ), .Z(\AES_ENC/sa33_next [4]) );
XOR2_X2 \AES_ENC/U1073  ( .A(\AES_ENC/n1145 ), .B(\AES_ENC/n1144 ), .Z(\AES_ENC/n1142 ) );
XOR2_X2 \AES_ENC/U1072  ( .A(\AES_ENC/n1230 ), .B(\AES_ENC/n1225 ), .Z(\AES_ENC/n1143 ) );
XOR2_X2 \AES_ENC/U1071  ( .A(\AES_ENC/sa21_sub[4] ), .B(\AES_ENC/sa32_sub[3] ), .Z(\AES_ENC/n1144 ) );
XOR2_X2 \AES_ENC/U1070  ( .A(\AES_ENC/w3[4] ), .B(\AES_ENC/sa03_sub[3] ),.Z(\AES_ENC/n1145 ) );
XOR2_X2 \AES_ENC/U1069  ( .A(\AES_ENC/n1147 ), .B(\AES_ENC/n1146 ), .Z(\AES_ENC/sa33_next [3]) );
XOR2_X2 \AES_ENC/U1068  ( .A(\AES_ENC/n1149 ), .B(\AES_ENC/n1148 ), .Z(\AES_ENC/n1146 ) );
XOR2_X2 \AES_ENC/U1067  ( .A(\AES_ENC/n1230 ), .B(\AES_ENC/n1226 ), .Z(\AES_ENC/n1147 ) );
XOR2_X2 \AES_ENC/U1066  ( .A(\AES_ENC/sa21_sub[3] ), .B(\AES_ENC/sa32_sub[2] ), .Z(\AES_ENC/n1148 ) );
XOR2_X2 \AES_ENC/U1065  ( .A(\AES_ENC/w3[3] ), .B(\AES_ENC/sa03_sub[2] ),.Z(\AES_ENC/n1149 ) );
XOR2_X2 \AES_ENC/U1064  ( .A(\AES_ENC/n1151 ), .B(\AES_ENC/n1150 ), .Z(\AES_ENC/sa33_next [2]) );
XOR2_X2 \AES_ENC/U1063  ( .A(\AES_ENC/n1227 ), .B(\AES_ENC/n1152 ), .Z(\AES_ENC/n1150 ) );
XOR2_X2 \AES_ENC/U1062  ( .A(\AES_ENC/sa21_sub[2] ), .B(\AES_ENC/sa32_sub[1] ), .Z(\AES_ENC/n1151 ) );
XOR2_X2 \AES_ENC/U1061  ( .A(\AES_ENC/w3[2] ), .B(\AES_ENC/sa03_sub[1] ),.Z(\AES_ENC/n1152 ) );
XOR2_X2 \AES_ENC/U1060  ( .A(\AES_ENC/n1154 ), .B(\AES_ENC/n1153 ), .Z(\AES_ENC/sa33_next [1]) );
XOR2_X2 \AES_ENC/U1059  ( .A(\AES_ENC/n1156 ), .B(\AES_ENC/n1155 ), .Z(\AES_ENC/n1153 ) );
XOR2_X2 \AES_ENC/U1058  ( .A(\AES_ENC/n1230 ), .B(\AES_ENC/n1228 ), .Z(\AES_ENC/n1154 ) );
XOR2_X2 \AES_ENC/U1057  ( .A(\AES_ENC/sa21_sub[1] ), .B(\AES_ENC/sa32_sub[0] ), .Z(\AES_ENC/n1155 ) );
XOR2_X2 \AES_ENC/U1056  ( .A(\AES_ENC/w3[1] ), .B(\AES_ENC/sa03_sub[0] ),.Z(\AES_ENC/n1156 ) );
XOR2_X2 \AES_ENC/U1055  ( .A(\AES_ENC/n1158 ), .B(\AES_ENC/n1157 ), .Z(\AES_ENC/sa33_next [0]) );
XOR2_X2 \AES_ENC/U1054  ( .A(\AES_ENC/n1230 ), .B(\AES_ENC/n1229 ), .Z(\AES_ENC/n1157 ) );
XOR2_X2 \AES_ENC/U1053  ( .A(\AES_ENC/w3[0] ), .B(\AES_ENC/sa21_sub[0] ),.Z(\AES_ENC/n1158 ) );
DFFR_X1 \AES_ENC/dcnt_reg_2_  ( .D(\AES_ENC/n795 ), .CK(clk), .RN(\AES_ENC/n1267 ), .Q(\AES_ENC/n1234 ), .QN() );
DFFR_X1 \AES_ENC/dcnt_reg_1_  ( .D(\AES_ENC/n796 ), .CK(clk), .RN(\AES_ENC/n1267 ), .Q(\AES_ENC/n1231 ), .QN(\AES_ENC/n794 ) );
DFFR_X1 \AES_ENC/dcnt_reg_3_  ( .D(\AES_ENC/n797 ), .CK(clk), .RN(\AES_ENC/n1267 ), .Q(\AES_ENC/n1233 ), .QN(\AES_ENC/n792 ) );
DFFR_X1 \AES_ENC/dcnt_reg_0_  ( .D(\AES_ENC/n798 ), .CK(clk), .RN(\AES_ENC/n1267 ), .Q(\AES_ENC/n1232 ), .QN(\AES_ENC/n2 ) );
INV_X4 \AES_ENC/u0/U558  ( .A(\AES_ENC/n1235 ), .ZN(\AES_ENC/u0/n319 ) );
INV_X4 \AES_ENC/u0/U557  ( .A(\AES_ENC/n1235 ), .ZN(\AES_ENC/u0/n325 ) );
INV_X4 \AES_ENC/u0/U556  ( .A(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n324 ) );
INV_X4 \AES_ENC/u0/U555  ( .A(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n322 ) );
INV_X4 \AES_ENC/u0/U554  ( .A(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n323 ) );
INV_X4 \AES_ENC/u0/U553  ( .A(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n321 ) );
INV_X4 \AES_ENC/u0/U552  ( .A(\AES_ENC/n1235 ), .ZN(\AES_ENC/u0/n320 ) );
INV_X4 \AES_ENC/u0/U551  ( .A(\AES_ENC/u0/n319 ), .ZN(\AES_ENC/u0/n318 ) );
INV_X4 \AES_ENC/u0/U550  ( .A(\AES_ENC/u0/n320 ), .ZN(\AES_ENC/u0/n317 ) );
INV_X4 \AES_ENC/u0/U549  ( .A(\AES_ENC/u0/n319 ), .ZN(\AES_ENC/u0/n316 ) );
INV_X4 \AES_ENC/u0/U548  ( .A(\AES_ENC/u0/n319 ), .ZN(\AES_ENC/u0/n315 ) );
NAND2_X1 \AES_ENC/u0/U411  ( .A1(n17502), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n870 ) );
NAND2_X1 \AES_ENC/u0/U410  ( .A1(n17501), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1520 ) );
NAND2_X1 \AES_ENC/u0/U407  ( .A1(n17500), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n630 ) );
NAND2_X1 \AES_ENC/u0/U404  ( .A1(n17499), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1360 ) );
NAND2_X1 \AES_ENC/u0/U401  ( .A1(n17498), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2000 ) );
NAND2_X1 \AES_ENC/u0/U398  ( .A1(n17497), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2640 ) );
NAND2_X1 \AES_ENC/u0/U395  ( .A1(n17496), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n600 ) );
NAND2_X1 \AES_ENC/u0/U392  ( .A1(n17495), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1340 ) );
NAND2_X1 \AES_ENC/u0/U389  ( .A1(n17494), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1980 ) );
NAND2_X1 \AES_ENC/u0/U386  ( .A1(n17493), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2620 ) );
NAND2_X1 \AES_ENC/u0/U383  ( .A1(n17492), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n570 ) );
NAND2_X1 \AES_ENC/u0/U380  ( .A1(n17491), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1320 ) );
NAND2_X1 \AES_ENC/u0/U377  ( .A1(n17490), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1960 ) );
NAND2_X1 \AES_ENC/u0/U374  ( .A1(n17489), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2600 ) );
NAND2_X1 \AES_ENC/u0/U371  ( .A1(n17488), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n540 ) );
NAND2_X1 \AES_ENC/u0/U368  ( .A1(n17487), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1300 ) );
NAND2_X1 \AES_ENC/u0/U365  ( .A1(n17486), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1940 ) );
NAND2_X1 \AES_ENC/u0/U362  ( .A1(n17485), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2580 ) );
NAND2_X1 \AES_ENC/u0/U359  ( .A1(n17484), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n510 ) );
NAND2_X1 \AES_ENC/u0/U356  ( .A1(n17483), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1280 ) );
NAND2_X1 \AES_ENC/u0/U353  ( .A1(n17482), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1920 ) );
NAND2_X1 \AES_ENC/u0/U350  ( .A1(n17481), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2560 ) );
NAND2_X1 \AES_ENC/u0/U347  ( .A1(n17480), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n480 ) );
NAND2_X1 \AES_ENC/u0/U344  ( .A1(n17479), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1260 ) );
NAND2_X1 \AES_ENC/u0/U341  ( .A1(n17478), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1900 ) );
NAND2_X1 \AES_ENC/u0/U338  ( .A1(n17477), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2540 ) );
NAND2_X1 \AES_ENC/u0/U335  ( .A1(n17476), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n450 ) );
NAND2_X1 \AES_ENC/u0/U332  ( .A1(n17475), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1240 ) );
NAND2_X1 \AES_ENC/u0/U329  ( .A1(n17474), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1880 ) );
NAND2_X1 \AES_ENC/u0/U326  ( .A1(n17473), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2520 ) );
NAND2_X1 \AES_ENC/u0/U323  ( .A1(n17472), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n420 ) );
NAND2_X1 \AES_ENC/u0/U320  ( .A1(n17471), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1220 ) );
NAND2_X1 \AES_ENC/u0/U317  ( .A1(n17470), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n39 ) );
NAND2_X1 \AES_ENC/u0/U314  ( .A1(n17469), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1200 ) );
NAND2_X1 \AES_ENC/u0/U311  ( .A1(n17468), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1840 ) );
NAND2_X1 \AES_ENC/u0/U308  ( .A1(n17467), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2480 ) );
NAND2_X1 \AES_ENC/u0/U305  ( .A1(n17466), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n36 ) );
NAND2_X1 \AES_ENC/u0/U30200  ( .A1(n17465), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1180 ) );
NAND2_X1 \AES_ENC/u0/U299  ( .A1(n17464), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1820 ) );
NAND2_X1 \AES_ENC/u0/U296  ( .A1(n17463), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2460 ) );
NAND2_X1 \AES_ENC/u0/U293  ( .A1(n17462), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n33 ) );
NAND2_X1 \AES_ENC/u0/U290  ( .A1(n17461), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1160 ) );
NAND2_X1 \AES_ENC/u0/U287  ( .A1(n17460), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1800 ) );
NAND2_X1 \AES_ENC/u0/U284  ( .A1(n17459), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2440 ) );
NAND2_X1 \AES_ENC/u0/U281  ( .A1(n17458), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n30 ) );
NAND2_X1 \AES_ENC/u0/U278  ( .A1(n17457), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1140 ) );
NAND2_X1 \AES_ENC/u0/U275  ( .A1(n17456), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1780 ) );
NAND2_X1 \AES_ENC/u0/U272  ( .A1(n17455), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2420 ) );
NAND2_X1 \AES_ENC/u0/U269  ( .A1(n17454), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n27 ) );
NAND2_X1 \AES_ENC/u0/U266  ( .A1(n17453), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1120 ) );
NAND2_X1 \AES_ENC/u0/U263  ( .A1(n17452), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1760 ) );
NAND2_X1 \AES_ENC/u0/U260  ( .A1(n17451), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2400 ) );
NAND2_X1 \AES_ENC/u0/U257  ( .A1(n17450), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n24 ) );
NAND2_X1 \AES_ENC/u0/U254  ( .A1(n17449), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1100 ) );
NAND2_X1 \AES_ENC/u0/U251  ( .A1(n17448), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1740 ) );
NAND2_X1 \AES_ENC/u0/U248  ( .A1(n17447), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2380 ) );
NAND2_X1 \AES_ENC/u0/U245  ( .A1(n17446), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n21 ) );
NAND2_X1 \AES_ENC/u0/U242  ( .A1(n17445), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1080 ) );
NAND2_X1 \AES_ENC/u0/U239  ( .A1(n17444), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1720 ) );
NAND2_X1 \AES_ENC/u0/U236  ( .A1(n17443), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2360 ) );
NAND2_X1 \AES_ENC/u0/U233  ( .A1(n17442), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n18 ) );
NAND2_X1 \AES_ENC/u0/U230  ( .A1(n17441), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1060 ) );
NAND2_X1 \AES_ENC/u0/U227  ( .A1(n17440), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1040 ) );
NAND2_X1 \AES_ENC/u0/U224  ( .A1(n17439), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1680 ) );
NAND2_X1 \AES_ENC/u0/U221  ( .A1(n17438), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2320 ) );
NAND2_X1 \AES_ENC/u0/U218  ( .A1(n17437), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1610 ) );
NAND2_X1 \AES_ENC/u0/U215  ( .A1(n17436), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1020 ) );
NAND2_X1 \AES_ENC/u0/U212  ( .A1(n17435), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1660 ) );
NAND2_X1 \AES_ENC/u0/U209  ( .A1(n17434), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2300 ) );
NAND2_X1 \AES_ENC/u0/U206  ( .A1(n17433), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n1400 ) );
NAND2_X1 \AES_ENC/u0/U203  ( .A1(n17432), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1000 ) );
NAND2_X1 \AES_ENC/u0/U200  ( .A1(n17431), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1640 ) );
NAND2_X1 \AES_ENC/u0/U197  ( .A1(n17430), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2280 ) );
NAND2_X1 \AES_ENC/u0/U194  ( .A1(n17429), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1210 ) );
NAND2_X1 \AES_ENC/u0/U191  ( .A1(n17428), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n980 ) );
NAND2_X1 \AES_ENC/u0/U188  ( .A1(n17427), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1620 ) );
NAND2_X1 \AES_ENC/u0/U185  ( .A1(n17426), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2260 ) );
NAND2_X1 \AES_ENC/u0/U182  ( .A1(n17425), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1010 ) );
NAND2_X1 \AES_ENC/u0/U179  ( .A1(n17424), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n960 ) );
NAND2_X1 \AES_ENC/u0/U176  ( .A1(n17423), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1600 ) );
NAND2_X1 \AES_ENC/u0/U173  ( .A1(n17422), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2240 ) );
NAND2_X1 \AES_ENC/u0/U170  ( .A1(n17421), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n8 ) );
NAND2_X1 \AES_ENC/u0/U167  ( .A1(n17420), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n940 ) );
NAND2_X1 \AES_ENC/u0/U164  ( .A1(n17419), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1580 ) );
NAND2_X1 \AES_ENC/u0/U161  ( .A1(n17418), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2220 ) );
NAND2_X1 \AES_ENC/u0/U158  ( .A1(n17417), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n6 ) );
NAND2_X1 \AES_ENC/u0/U155  ( .A1(n17416), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n920 ) );
NAND2_X1 \AES_ENC/u0/U152  ( .A1(n17415), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1560 ) );
NAND2_X1 \AES_ENC/u0/U149  ( .A1(n17414), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2200 ) );
NAND2_X1 \AES_ENC/u0/U146  ( .A1(n17413), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n4 ) );
NAND2_X1 \AES_ENC/u0/U143  ( .A1(n17412), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n900 ) );
NAND2_X1 \AES_ENC/u0/U140  ( .A1(n17411), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n840 ) );
NAND2_X1 \AES_ENC/u0/U137  ( .A1(n17410), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1500 ) );
NAND2_X1 \AES_ENC/u0/U134  ( .A1(n17409), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2140 ) );
NAND2_X1 \AES_ENC/u0/U131  ( .A1(n17408), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n278 ) );
NAND2_X1 \AES_ENC/u0/U128  ( .A1(n17407), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n810 ) );
NAND2_X1 \AES_ENC/u0/U125  ( .A1(n17406), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1480 ) );
NAND2_X1 \AES_ENC/u0/U122  ( .A1(n17405), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2120 ) );
NAND2_X1 \AES_ENC/u0/U118  ( .A1(n17404), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n276 ) );
NAND2_X1 \AES_ENC/u0/U114  ( .A1(n17403), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n780 ) );
NAND2_X1 \AES_ENC/u0/U110  ( .A1(n17402), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1460 ) );
NAND2_X1 \AES_ENC/u0/U106  ( .A1(n17401), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2100 ) );
NAND2_X1 \AES_ENC/u0/U102  ( .A1(n17400), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n274 ) );
NAND2_X1 \AES_ENC/u0/U98  ( .A1(n17399), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n75 ) );
NAND2_X1 \AES_ENC/u0/U94  ( .A1(n17398), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1440 ) );
NAND2_X1 \AES_ENC/u0/U90  ( .A1(n17397), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2080 ) );
NAND2_X1 \AES_ENC/u0/U86  ( .A1(n17396), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n272 ) );
NAND2_X1 \AES_ENC/u0/U82  ( .A1(n17395), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n720 ) );
NAND2_X1 \AES_ENC/u0/U78  ( .A1(n17394), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1420 ) );
NAND2_X1 \AES_ENC/u0/U74  ( .A1(n17393), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n206 ) );
NAND2_X1 \AES_ENC/u0/U70  ( .A1(n17392), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2700 ) );
NAND2_X1 \AES_ENC/u0/U66  ( .A1(n17391), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n690 ) );
NAND2_X1 \AES_ENC/u0/U62  ( .A1(n17390), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1401 ) );
NAND2_X1 \AES_ENC/u0/U58  ( .A1(n17389), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2040 ) );
NAND2_X1 \AES_ENC/u0/U54  ( .A1(n17388), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2680 ) );
NAND2_X1 \AES_ENC/u0/U50  ( .A1(n17387), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n660 ) );
NAND2_X1 \AES_ENC/u0/U46  ( .A1(n17386), .A2(\AES_ENC/u0/n317 ), .ZN(\AES_ENC/u0/n1380 ) );
NAND2_X1 \AES_ENC/u0/U42  ( .A1(n17385), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2020 ) );
NAND2_X1 \AES_ENC/u0/U38  ( .A1(n17384), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2660 ) );
NAND2_X1 \AES_ENC/u0/U34  ( .A1(n17383), .A2(\AES_ENC/u0/n316 ), .ZN(\AES_ENC/u0/n1540 ) );
NAND2_X1 \AES_ENC/u0/U3020  ( .A1(n17382), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2180 ) );
NAND2_X1 \AES_ENC/u0/U26  ( .A1(\AES_ENC/u0/n316 ), .A2(cii_K[127]), .ZN(\AES_ENC/u0/n2 ) );
NAND2_X1 \AES_ENC/u0/U23  ( .A1(\AES_ENC/u0/n2 ), .A2(\AES_ENC/u0/n3 ), .ZN(\AES_ENC/u0/N73 ) );
BUF_X32 \AES_ENC/u0/U20  ( .A(\AES_ENC/u0/N73 ), .Z(\AES_ENC/u0/n314 ) );
NAND2_X1 \AES_ENC/u0/U17  ( .A1(n17381), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1700 ) );
NAND2_X1 \AES_ENC/u0/U14  ( .A1(n17380), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2340 ) );
NAND2_X1 \AES_ENC/u0/U11  ( .A1(n17379), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n1860 ) );
NAND2_X1 \AES_ENC/u0/U8  ( .A1(n17378), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2500 ) );
NAND2_X1 \AES_ENC/u0/U5  ( .A1(n17377), .A2(\AES_ENC/u0/n318 ), .ZN(\AES_ENC/u0/n2160 ) );
NAND2_X1 \AES_ENC/u0/U3010  ( .A1(n17376), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/n280 ) );
NAND2_X2 \AES_ENC/u0/U409  ( .A1(\AES_ENC/u0/N107 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n281 ) );
NAND2_X2 \AES_ENC/u0/U408  ( .A1(\AES_ENC/u0/n280 ), .A2(\AES_ENC/u0/n281 ),.ZN(\AES_ENC/u0/N108 ) );
NAND2_X2 \AES_ENC/u0/U406  ( .A1(\AES_ENC/u0/N106 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n279 ) );
NAND2_X2 \AES_ENC/u0/U405  ( .A1(\AES_ENC/u0/n278 ), .A2(\AES_ENC/u0/n279 ),.ZN(\AES_ENC/u0/N109 ) );
NAND2_X2 \AES_ENC/u0/U403  ( .A1(\AES_ENC/u0/N105 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n277 ) );
NAND2_X2 \AES_ENC/u0/U402  ( .A1(\AES_ENC/u0/n276 ), .A2(\AES_ENC/u0/n277 ),.ZN(\AES_ENC/u0/N110 ) );
NAND2_X2 \AES_ENC/u0/U400  ( .A1(\AES_ENC/u0/N104 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n275 ) );
NAND2_X2 \AES_ENC/u0/U399  ( .A1(\AES_ENC/u0/n274 ), .A2(\AES_ENC/u0/n275 ),.ZN(\AES_ENC/u0/N111 ) );
NAND2_X2 \AES_ENC/u0/U397  ( .A1(\AES_ENC/u0/N103 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n273 ) );
NAND2_X2 \AES_ENC/u0/U396  ( .A1(\AES_ENC/u0/n272 ), .A2(\AES_ENC/u0/n273 ),.ZN(\AES_ENC/u0/N112 ) );
NAND2_X2 \AES_ENC/u0/U394  ( .A1(\AES_ENC/u0/N102 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n2710 ) );
NAND2_X2 \AES_ENC/u0/U393  ( .A1(\AES_ENC/u0/n2700 ), .A2(\AES_ENC/u0/n2710 ), .ZN(\AES_ENC/u0/N113 ) );
NAND2_X2 \AES_ENC/u0/U391  ( .A1(\AES_ENC/u0/N101 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n2690 ) );
NAND2_X2 \AES_ENC/u0/U390  ( .A1(\AES_ENC/u0/n2680 ), .A2(\AES_ENC/u0/n2690 ), .ZN(\AES_ENC/u0/N114 ) );
NAND2_X2 \AES_ENC/u0/U388  ( .A1(\AES_ENC/u0/N100 ), .A2(\AES_ENC/u0/n319 ),.ZN(\AES_ENC/u0/n2670 ) );
NAND2_X2 \AES_ENC/u0/U387  ( .A1(\AES_ENC/u0/n2660 ), .A2(\AES_ENC/u0/n2670 ), .ZN(\AES_ENC/u0/N115 ) );
NAND2_X2 \AES_ENC/u0/U385  ( .A1(\AES_ENC/u0/N99 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2650 ) );
NAND2_X2 \AES_ENC/u0/U384  ( .A1(\AES_ENC/u0/n2640 ), .A2(\AES_ENC/u0/n2650 ), .ZN(\AES_ENC/u0/N116 ) );
NAND2_X2 \AES_ENC/u0/U382  ( .A1(\AES_ENC/u0/N98 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2630 ) );
NAND2_X2 \AES_ENC/u0/U381  ( .A1(\AES_ENC/u0/n2620 ), .A2(\AES_ENC/u0/n2630 ), .ZN(\AES_ENC/u0/N117 ) );
NAND2_X2 \AES_ENC/u0/U379  ( .A1(\AES_ENC/u0/N97 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2610 ) );
NAND2_X2 \AES_ENC/u0/U378  ( .A1(\AES_ENC/u0/n2600 ), .A2(\AES_ENC/u0/n2610 ), .ZN(\AES_ENC/u0/N118 ) );
NAND2_X2 \AES_ENC/u0/U376  ( .A1(\AES_ENC/u0/N96 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2590 ) );
NAND2_X2 \AES_ENC/u0/U375  ( .A1(\AES_ENC/u0/n2580 ), .A2(\AES_ENC/u0/n2590 ), .ZN(\AES_ENC/u0/N119 ) );
NAND2_X2 \AES_ENC/u0/U373  ( .A1(\AES_ENC/u0/N95 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2570 ) );
NAND2_X2 \AES_ENC/u0/U372  ( .A1(\AES_ENC/u0/n2560 ), .A2(\AES_ENC/u0/n2570 ), .ZN(\AES_ENC/u0/N120 ) );
NAND2_X2 \AES_ENC/u0/U370  ( .A1(\AES_ENC/u0/N94 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2550 ) );
NAND2_X2 \AES_ENC/u0/U369  ( .A1(\AES_ENC/u0/n2540 ), .A2(\AES_ENC/u0/n2550 ), .ZN(\AES_ENC/u0/N121 ) );
NAND2_X2 \AES_ENC/u0/U367  ( .A1(\AES_ENC/u0/N93 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2530 ) );
NAND2_X2 \AES_ENC/u0/U366  ( .A1(\AES_ENC/u0/n2520 ), .A2(\AES_ENC/u0/n2530 ), .ZN(\AES_ENC/u0/N122 ) );
NAND2_X2 \AES_ENC/u0/U364  ( .A1(\AES_ENC/u0/N92 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2510 ) );
NAND2_X2 \AES_ENC/u0/U363  ( .A1(\AES_ENC/u0/n2500 ), .A2(\AES_ENC/u0/n2510 ), .ZN(\AES_ENC/u0/N123 ) );
NAND2_X2 \AES_ENC/u0/U361  ( .A1(\AES_ENC/u0/N91 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2490 ) );
NAND2_X2 \AES_ENC/u0/U360  ( .A1(\AES_ENC/u0/n2480 ), .A2(\AES_ENC/u0/n2490 ), .ZN(\AES_ENC/u0/N124 ) );
NAND2_X2 \AES_ENC/u0/U358  ( .A1(\AES_ENC/u0/N90 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2470 ) );
NAND2_X2 \AES_ENC/u0/U357  ( .A1(\AES_ENC/u0/n2460 ), .A2(\AES_ENC/u0/n2470 ), .ZN(\AES_ENC/u0/N125 ) );
NAND2_X2 \AES_ENC/u0/U355  ( .A1(\AES_ENC/u0/N89 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2450 ) );
NAND2_X2 \AES_ENC/u0/U354  ( .A1(\AES_ENC/u0/n2440 ), .A2(\AES_ENC/u0/n2450 ), .ZN(\AES_ENC/u0/N126 ) );
NAND2_X2 \AES_ENC/u0/U352  ( .A1(\AES_ENC/u0/N88 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2430 ) );
NAND2_X2 \AES_ENC/u0/U351  ( .A1(\AES_ENC/u0/n2420 ), .A2(\AES_ENC/u0/n2430 ), .ZN(\AES_ENC/u0/N127 ) );
NAND2_X2 \AES_ENC/u0/U349  ( .A1(\AES_ENC/u0/N87 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2410 ) );
NAND2_X2 \AES_ENC/u0/U348  ( .A1(\AES_ENC/u0/n2400 ), .A2(\AES_ENC/u0/n2410 ), .ZN(\AES_ENC/u0/N128 ) );
NAND2_X2 \AES_ENC/u0/U346  ( .A1(\AES_ENC/u0/N86 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2390 ) );
NAND2_X2 \AES_ENC/u0/U345  ( .A1(\AES_ENC/u0/n2380 ), .A2(\AES_ENC/u0/n2390 ), .ZN(\AES_ENC/u0/N129 ) );
NAND2_X2 \AES_ENC/u0/U343  ( .A1(\AES_ENC/u0/N85 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2370 ) );
NAND2_X2 \AES_ENC/u0/U342  ( .A1(\AES_ENC/u0/n2360 ), .A2(\AES_ENC/u0/n2370 ), .ZN(\AES_ENC/u0/N130 ) );
NAND2_X2 \AES_ENC/u0/U340  ( .A1(\AES_ENC/u0/N84 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2350 ) );
NAND2_X2 \AES_ENC/u0/U339  ( .A1(\AES_ENC/u0/n2340 ), .A2(\AES_ENC/u0/n2350 ), .ZN(\AES_ENC/u0/N131 ) );
NAND2_X2 \AES_ENC/u0/U337  ( .A1(\AES_ENC/u0/N83 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2330 ) );
NAND2_X2 \AES_ENC/u0/U336  ( .A1(\AES_ENC/u0/n2320 ), .A2(\AES_ENC/u0/n2330 ), .ZN(\AES_ENC/u0/N132 ) );
NAND2_X2 \AES_ENC/u0/U334  ( .A1(\AES_ENC/u0/N82 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2310 ) );
NAND2_X2 \AES_ENC/u0/U333  ( .A1(\AES_ENC/u0/n2300 ), .A2(\AES_ENC/u0/n2310 ), .ZN(\AES_ENC/u0/N133 ) );
NAND2_X2 \AES_ENC/u0/U331  ( .A1(\AES_ENC/u0/N81 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2290 ) );
NAND2_X2 \AES_ENC/u0/U330  ( .A1(\AES_ENC/u0/n2280 ), .A2(\AES_ENC/u0/n2290 ), .ZN(\AES_ENC/u0/N134 ) );
NAND2_X2 \AES_ENC/u0/U328  ( .A1(\AES_ENC/u0/N80 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2270 ) );
NAND2_X2 \AES_ENC/u0/U327  ( .A1(\AES_ENC/u0/n2260 ), .A2(\AES_ENC/u0/n2270 ), .ZN(\AES_ENC/u0/N135 ) );
NAND2_X2 \AES_ENC/u0/U325  ( .A1(\AES_ENC/u0/N79 ), .A2(\AES_ENC/u0/n320 ),.ZN(\AES_ENC/u0/n2250 ) );
NAND2_X2 \AES_ENC/u0/U324  ( .A1(\AES_ENC/u0/n2240 ), .A2(\AES_ENC/u0/n2250 ), .ZN(\AES_ENC/u0/N136 ) );
NAND2_X2 \AES_ENC/u0/U322  ( .A1(\AES_ENC/u0/N78 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2230 ) );
NAND2_X2 \AES_ENC/u0/U321  ( .A1(\AES_ENC/u0/n2220 ), .A2(\AES_ENC/u0/n2230 ), .ZN(\AES_ENC/u0/N137 ) );
NAND2_X2 \AES_ENC/u0/U319  ( .A1(\AES_ENC/u0/N77 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2210 ) );
NAND2_X2 \AES_ENC/u0/U318  ( .A1(\AES_ENC/u0/n2200 ), .A2(\AES_ENC/u0/n2210 ), .ZN(\AES_ENC/u0/N138 ) );
NAND2_X2 \AES_ENC/u0/U316  ( .A1(\AES_ENC/u0/N76 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2190 ) );
NAND2_X2 \AES_ENC/u0/U315  ( .A1(\AES_ENC/u0/n2180 ), .A2(\AES_ENC/u0/n2190 ), .ZN(\AES_ENC/u0/N139 ) );
NAND2_X2 \AES_ENC/u0/U313  ( .A1(\AES_ENC/u0/N173 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2170 ) );
NAND2_X2 \AES_ENC/u0/U312  ( .A1(\AES_ENC/u0/n2160 ), .A2(\AES_ENC/u0/n2170 ), .ZN(\AES_ENC/u0/N174 ) );
NAND2_X2 \AES_ENC/u0/U310  ( .A1(\AES_ENC/u0/N172 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2150 ) );
NAND2_X2 \AES_ENC/u0/U309  ( .A1(\AES_ENC/u0/n2140 ), .A2(\AES_ENC/u0/n2150 ), .ZN(\AES_ENC/u0/N175 ) );
NAND2_X2 \AES_ENC/u0/U307  ( .A1(\AES_ENC/u0/N171 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2130 ) );
NAND2_X2 \AES_ENC/u0/U306  ( .A1(\AES_ENC/u0/n2120 ), .A2(\AES_ENC/u0/n2130 ), .ZN(\AES_ENC/u0/N176 ) );
NAND2_X2 \AES_ENC/u0/U304  ( .A1(\AES_ENC/u0/N170 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2110 ) );
NAND2_X2 \AES_ENC/u0/U303  ( .A1(\AES_ENC/u0/n2100 ), .A2(\AES_ENC/u0/n2110 ), .ZN(\AES_ENC/u0/N177 ) );
NAND2_X2 \AES_ENC/u0/U301  ( .A1(\AES_ENC/u0/N169 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2090 ) );
NAND2_X2 \AES_ENC/u0/U300  ( .A1(\AES_ENC/u0/n2080 ), .A2(\AES_ENC/u0/n2090 ), .ZN(\AES_ENC/u0/N178 ) );
NAND2_X2 \AES_ENC/u0/U298  ( .A1(\AES_ENC/u0/N168 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n207 ) );
NAND2_X2 \AES_ENC/u0/U297  ( .A1(\AES_ENC/u0/n206 ), .A2(\AES_ENC/u0/n207 ),.ZN(\AES_ENC/u0/N179 ) );
NAND2_X2 \AES_ENC/u0/U295  ( .A1(\AES_ENC/u0/N167 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2050 ) );
NAND2_X2 \AES_ENC/u0/U294  ( .A1(\AES_ENC/u0/n2040 ), .A2(\AES_ENC/u0/n2050 ), .ZN(\AES_ENC/u0/N180 ) );
NAND2_X2 \AES_ENC/u0/U292  ( .A1(\AES_ENC/u0/N166 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2030 ) );
NAND2_X2 \AES_ENC/u0/U291  ( .A1(\AES_ENC/u0/n2020 ), .A2(\AES_ENC/u0/n2030 ), .ZN(\AES_ENC/u0/N181 ) );
NAND2_X2 \AES_ENC/u0/U289  ( .A1(\AES_ENC/u0/N165 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n2010 ) );
NAND2_X2 \AES_ENC/u0/U288  ( .A1(\AES_ENC/u0/n2000 ), .A2(\AES_ENC/u0/n2010 ), .ZN(\AES_ENC/u0/N182 ) );
NAND2_X2 \AES_ENC/u0/U286  ( .A1(\AES_ENC/u0/N164 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1990 ) );
NAND2_X2 \AES_ENC/u0/U285  ( .A1(\AES_ENC/u0/n1980 ), .A2(\AES_ENC/u0/n1990 ), .ZN(\AES_ENC/u0/N183 ) );
NAND2_X2 \AES_ENC/u0/U283  ( .A1(\AES_ENC/u0/N163 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1970 ) );
NAND2_X2 \AES_ENC/u0/U282  ( .A1(\AES_ENC/u0/n1960 ), .A2(\AES_ENC/u0/n1970 ), .ZN(\AES_ENC/u0/N184 ) );
NAND2_X2 \AES_ENC/u0/U280  ( .A1(\AES_ENC/u0/N162 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1950 ) );
NAND2_X2 \AES_ENC/u0/U279  ( .A1(\AES_ENC/u0/n1940 ), .A2(\AES_ENC/u0/n1950 ), .ZN(\AES_ENC/u0/N185 ) );
NAND2_X2 \AES_ENC/u0/U277  ( .A1(\AES_ENC/u0/N161 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1930 ) );
NAND2_X2 \AES_ENC/u0/U276  ( .A1(\AES_ENC/u0/n1920 ), .A2(\AES_ENC/u0/n1930 ), .ZN(\AES_ENC/u0/N186 ) );
NAND2_X2 \AES_ENC/u0/U274  ( .A1(\AES_ENC/u0/N160 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1910 ) );
NAND2_X2 \AES_ENC/u0/U273  ( .A1(\AES_ENC/u0/n1900 ), .A2(\AES_ENC/u0/n1910 ), .ZN(\AES_ENC/u0/N187 ) );
NAND2_X2 \AES_ENC/u0/U271  ( .A1(\AES_ENC/u0/N159 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1890 ) );
NAND2_X2 \AES_ENC/u0/U270  ( .A1(\AES_ENC/u0/n1880 ), .A2(\AES_ENC/u0/n1890 ), .ZN(\AES_ENC/u0/N188 ) );
NAND2_X2 \AES_ENC/u0/U268  ( .A1(\AES_ENC/u0/N158 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1870 ) );
NAND2_X2 \AES_ENC/u0/U267  ( .A1(\AES_ENC/u0/n1860 ), .A2(\AES_ENC/u0/n1870 ), .ZN(\AES_ENC/u0/N189 ) );
NAND2_X2 \AES_ENC/u0/U265  ( .A1(\AES_ENC/u0/N157 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1850 ) );
NAND2_X2 \AES_ENC/u0/U264  ( .A1(\AES_ENC/u0/n1840 ), .A2(\AES_ENC/u0/n1850 ), .ZN(\AES_ENC/u0/N190 ) );
NAND2_X2 \AES_ENC/u0/U262  ( .A1(\AES_ENC/u0/N156 ), .A2(\AES_ENC/u0/n321 ),.ZN(\AES_ENC/u0/n1830 ) );
NAND2_X2 \AES_ENC/u0/U261  ( .A1(\AES_ENC/u0/n1820 ), .A2(\AES_ENC/u0/n1830 ), .ZN(\AES_ENC/u0/N191 ) );
NAND2_X2 \AES_ENC/u0/U259  ( .A1(\AES_ENC/u0/N155 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1810 ) );
NAND2_X2 \AES_ENC/u0/U258  ( .A1(\AES_ENC/u0/n1800 ), .A2(\AES_ENC/u0/n1810 ), .ZN(\AES_ENC/u0/N192 ) );
NAND2_X2 \AES_ENC/u0/U256  ( .A1(\AES_ENC/u0/N154 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1790 ) );
NAND2_X2 \AES_ENC/u0/U255  ( .A1(\AES_ENC/u0/n1780 ), .A2(\AES_ENC/u0/n1790 ), .ZN(\AES_ENC/u0/N193 ) );
NAND2_X2 \AES_ENC/u0/U253  ( .A1(\AES_ENC/u0/N153 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1770 ) );
NAND2_X2 \AES_ENC/u0/U252  ( .A1(\AES_ENC/u0/n1760 ), .A2(\AES_ENC/u0/n1770 ), .ZN(\AES_ENC/u0/N194 ) );
NAND2_X2 \AES_ENC/u0/U250  ( .A1(\AES_ENC/u0/N152 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1750 ) );
NAND2_X2 \AES_ENC/u0/U249  ( .A1(\AES_ENC/u0/n1740 ), .A2(\AES_ENC/u0/n1750 ), .ZN(\AES_ENC/u0/N195 ) );
NAND2_X2 \AES_ENC/u0/U247  ( .A1(\AES_ENC/u0/N151 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1730 ) );
NAND2_X2 \AES_ENC/u0/U246  ( .A1(\AES_ENC/u0/n1720 ), .A2(\AES_ENC/u0/n1730 ), .ZN(\AES_ENC/u0/N196 ) );
NAND2_X2 \AES_ENC/u0/U244  ( .A1(\AES_ENC/u0/N150 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1711 ) );
NAND2_X2 \AES_ENC/u0/U243  ( .A1(\AES_ENC/u0/n1700 ), .A2(\AES_ENC/u0/n1711 ), .ZN(\AES_ENC/u0/N197 ) );
NAND2_X2 \AES_ENC/u0/U241  ( .A1(\AES_ENC/u0/N149 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1690 ) );
NAND2_X2 \AES_ENC/u0/U240  ( .A1(\AES_ENC/u0/n1680 ), .A2(\AES_ENC/u0/n1690 ), .ZN(\AES_ENC/u0/N198 ) );
NAND2_X2 \AES_ENC/u0/U238  ( .A1(\AES_ENC/u0/N148 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1670 ) );
NAND2_X2 \AES_ENC/u0/U237  ( .A1(\AES_ENC/u0/n1660 ), .A2(\AES_ENC/u0/n1670 ), .ZN(\AES_ENC/u0/N199 ) );
NAND2_X2 \AES_ENC/u0/U235  ( .A1(\AES_ENC/u0/N147 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1650 ) );
NAND2_X2 \AES_ENC/u0/U234  ( .A1(\AES_ENC/u0/n1640 ), .A2(\AES_ENC/u0/n1650 ), .ZN(\AES_ENC/u0/N200 ) );
NAND2_X2 \AES_ENC/u0/U232  ( .A1(\AES_ENC/u0/N146 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1630 ) );
NAND2_X2 \AES_ENC/u0/U231  ( .A1(\AES_ENC/u0/n1620 ), .A2(\AES_ENC/u0/n1630 ), .ZN(\AES_ENC/u0/N201 ) );
NAND2_X2 \AES_ENC/u0/U229  ( .A1(\AES_ENC/u0/N145 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1611 ) );
NAND2_X2 \AES_ENC/u0/U228  ( .A1(\AES_ENC/u0/n1600 ), .A2(\AES_ENC/u0/n1611 ), .ZN(\AES_ENC/u0/N202 ) );
NAND2_X2 \AES_ENC/u0/U226  ( .A1(\AES_ENC/u0/N144 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1590 ) );
NAND2_X2 \AES_ENC/u0/U225  ( .A1(\AES_ENC/u0/n1580 ), .A2(\AES_ENC/u0/n1590 ), .ZN(\AES_ENC/u0/N203 ) );
NAND2_X2 \AES_ENC/u0/U223  ( .A1(\AES_ENC/u0/N143 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1570 ) );
NAND2_X2 \AES_ENC/u0/U222  ( .A1(\AES_ENC/u0/n1560 ), .A2(\AES_ENC/u0/n1570 ), .ZN(\AES_ENC/u0/N204 ) );
NAND2_X2 \AES_ENC/u0/U220  ( .A1(\AES_ENC/u0/N142 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1550 ) );
NAND2_X2 \AES_ENC/u0/U219  ( .A1(\AES_ENC/u0/n1540 ), .A2(\AES_ENC/u0/n1550 ), .ZN(\AES_ENC/u0/N205 ) );
NAND2_X2 \AES_ENC/u0/U217  ( .A1(\AES_ENC/u0/N239 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1530 ) );
NAND2_X2 \AES_ENC/u0/U216  ( .A1(\AES_ENC/u0/n1520 ), .A2(\AES_ENC/u0/n1530 ), .ZN(\AES_ENC/u0/N240 ) );
NAND2_X2 \AES_ENC/u0/U214  ( .A1(\AES_ENC/u0/N238 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1511 ) );
NAND2_X2 \AES_ENC/u0/U213  ( .A1(\AES_ENC/u0/n1500 ), .A2(\AES_ENC/u0/n1511 ), .ZN(\AES_ENC/u0/N241 ) );
NAND2_X2 \AES_ENC/u0/U211  ( .A1(\AES_ENC/u0/N237 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1490 ) );
NAND2_X2 \AES_ENC/u0/U210  ( .A1(\AES_ENC/u0/n1480 ), .A2(\AES_ENC/u0/n1490 ), .ZN(\AES_ENC/u0/N242 ) );
NAND2_X2 \AES_ENC/u0/U208  ( .A1(\AES_ENC/u0/N236 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1470 ) );
NAND2_X2 \AES_ENC/u0/U207  ( .A1(\AES_ENC/u0/n1460 ), .A2(\AES_ENC/u0/n1470 ), .ZN(\AES_ENC/u0/N243 ) );
NAND2_X2 \AES_ENC/u0/U205  ( .A1(\AES_ENC/u0/N235 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1450 ) );
NAND2_X2 \AES_ENC/u0/U204  ( .A1(\AES_ENC/u0/n1440 ), .A2(\AES_ENC/u0/n1450 ), .ZN(\AES_ENC/u0/N244 ) );
NAND2_X2 \AES_ENC/u0/U202  ( .A1(\AES_ENC/u0/N234 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n1430 ) );
NAND2_X2 \AES_ENC/u0/U201  ( .A1(\AES_ENC/u0/n1420 ), .A2(\AES_ENC/u0/n1430 ), .ZN(\AES_ENC/u0/N245 ) );
NAND2_X2 \AES_ENC/u0/U199  ( .A1(\AES_ENC/u0/N233 ), .A2(\AES_ENC/u0/n322 ),.ZN(\AES_ENC/u0/n141 ) );
NAND2_X2 \AES_ENC/u0/U198  ( .A1(\AES_ENC/u0/n1401 ), .A2(\AES_ENC/u0/n141 ),.ZN(\AES_ENC/u0/N246 ) );
NAND2_X2 \AES_ENC/u0/U196  ( .A1(\AES_ENC/u0/N232 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1390 ) );
NAND2_X2 \AES_ENC/u0/U195  ( .A1(\AES_ENC/u0/n1380 ), .A2(\AES_ENC/u0/n1390 ), .ZN(\AES_ENC/u0/N247 ) );
NAND2_X2 \AES_ENC/u0/U193  ( .A1(\AES_ENC/u0/N231 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1370 ) );
NAND2_X2 \AES_ENC/u0/U192  ( .A1(\AES_ENC/u0/n1360 ), .A2(\AES_ENC/u0/n1370 ), .ZN(\AES_ENC/u0/N248 ) );
NAND2_X2 \AES_ENC/u0/U190  ( .A1(\AES_ENC/u0/N230 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1350 ) );
NAND2_X2 \AES_ENC/u0/U189  ( .A1(\AES_ENC/u0/n1340 ), .A2(\AES_ENC/u0/n1350 ), .ZN(\AES_ENC/u0/N249 ) );
NAND2_X2 \AES_ENC/u0/U187  ( .A1(\AES_ENC/u0/N229 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1330 ) );
NAND2_X2 \AES_ENC/u0/U186  ( .A1(\AES_ENC/u0/n1320 ), .A2(\AES_ENC/u0/n1330 ), .ZN(\AES_ENC/u0/N250 ) );
NAND2_X2 \AES_ENC/u0/U184  ( .A1(\AES_ENC/u0/N228 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1311 ) );
NAND2_X2 \AES_ENC/u0/U183  ( .A1(\AES_ENC/u0/n1300 ), .A2(\AES_ENC/u0/n1311 ), .ZN(\AES_ENC/u0/N251 ) );
NAND2_X2 \AES_ENC/u0/U181  ( .A1(\AES_ENC/u0/N227 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1290 ) );
NAND2_X2 \AES_ENC/u0/U180  ( .A1(\AES_ENC/u0/n1280 ), .A2(\AES_ENC/u0/n1290 ), .ZN(\AES_ENC/u0/N252 ) );
NAND2_X2 \AES_ENC/u0/U178  ( .A1(\AES_ENC/u0/N226 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1270 ) );
NAND2_X2 \AES_ENC/u0/U177  ( .A1(\AES_ENC/u0/n1260 ), .A2(\AES_ENC/u0/n1270 ), .ZN(\AES_ENC/u0/N253 ) );
NAND2_X2 \AES_ENC/u0/U175  ( .A1(\AES_ENC/u0/N225 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1250 ) );
NAND2_X2 \AES_ENC/u0/U174  ( .A1(\AES_ENC/u0/n1240 ), .A2(\AES_ENC/u0/n1250 ), .ZN(\AES_ENC/u0/N254 ) );
NAND2_X2 \AES_ENC/u0/U172  ( .A1(\AES_ENC/u0/N224 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1230 ) );
NAND2_X2 \AES_ENC/u0/U171  ( .A1(\AES_ENC/u0/n1220 ), .A2(\AES_ENC/u0/n1230 ), .ZN(\AES_ENC/u0/N255 ) );
NAND2_X2 \AES_ENC/u0/U169  ( .A1(\AES_ENC/u0/N223 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1211 ) );
NAND2_X2 \AES_ENC/u0/U168  ( .A1(\AES_ENC/u0/n1200 ), .A2(\AES_ENC/u0/n1211 ), .ZN(\AES_ENC/u0/N256 ) );
NAND2_X2 \AES_ENC/u0/U166  ( .A1(\AES_ENC/u0/N222 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1190 ) );
NAND2_X2 \AES_ENC/u0/U165  ( .A1(\AES_ENC/u0/n1180 ), .A2(\AES_ENC/u0/n1190 ), .ZN(\AES_ENC/u0/N257 ) );
NAND2_X2 \AES_ENC/u0/U163  ( .A1(\AES_ENC/u0/N221 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1170 ) );
NAND2_X2 \AES_ENC/u0/U162  ( .A1(\AES_ENC/u0/n1160 ), .A2(\AES_ENC/u0/n1170 ), .ZN(\AES_ENC/u0/N258 ) );
NAND2_X2 \AES_ENC/u0/U160  ( .A1(\AES_ENC/u0/N220 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1150 ) );
NAND2_X2 \AES_ENC/u0/U159  ( .A1(\AES_ENC/u0/n1140 ), .A2(\AES_ENC/u0/n1150 ), .ZN(\AES_ENC/u0/N259 ) );
NAND2_X2 \AES_ENC/u0/U157  ( .A1(\AES_ENC/u0/N219 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1130 ) );
NAND2_X2 \AES_ENC/u0/U156  ( .A1(\AES_ENC/u0/n1120 ), .A2(\AES_ENC/u0/n1130 ), .ZN(\AES_ENC/u0/N260 ) );
NAND2_X2 \AES_ENC/u0/U154  ( .A1(\AES_ENC/u0/N218 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1111 ) );
NAND2_X2 \AES_ENC/u0/U153  ( .A1(\AES_ENC/u0/n1100 ), .A2(\AES_ENC/u0/n1111 ), .ZN(\AES_ENC/u0/N261 ) );
NAND2_X2 \AES_ENC/u0/U151  ( .A1(\AES_ENC/u0/N217 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1090 ) );
NAND2_X2 \AES_ENC/u0/U150  ( .A1(\AES_ENC/u0/n1080 ), .A2(\AES_ENC/u0/n1090 ), .ZN(\AES_ENC/u0/N262 ) );
NAND2_X2 \AES_ENC/u0/U148  ( .A1(\AES_ENC/u0/N216 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1070 ) );
NAND2_X2 \AES_ENC/u0/U147  ( .A1(\AES_ENC/u0/n1060 ), .A2(\AES_ENC/u0/n1070 ), .ZN(\AES_ENC/u0/N263 ) );
NAND2_X2 \AES_ENC/u0/U145  ( .A1(\AES_ENC/u0/N215 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1050 ) );
NAND2_X2 \AES_ENC/u0/U144  ( .A1(\AES_ENC/u0/n1040 ), .A2(\AES_ENC/u0/n1050 ), .ZN(\AES_ENC/u0/N264 ) );
NAND2_X2 \AES_ENC/u0/U142  ( .A1(\AES_ENC/u0/N214 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1030 ) );
NAND2_X2 \AES_ENC/u0/U141  ( .A1(\AES_ENC/u0/n1020 ), .A2(\AES_ENC/u0/n1030 ), .ZN(\AES_ENC/u0/N265 ) );
NAND2_X2 \AES_ENC/u0/U139  ( .A1(\AES_ENC/u0/N213 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n1011 ) );
NAND2_X2 \AES_ENC/u0/U138  ( .A1(\AES_ENC/u0/n1000 ), .A2(\AES_ENC/u0/n1011 ), .ZN(\AES_ENC/u0/N266 ) );
NAND2_X2 \AES_ENC/u0/U136  ( .A1(\AES_ENC/u0/N212 ), .A2(\AES_ENC/u0/n323 ),.ZN(\AES_ENC/u0/n990 ) );
NAND2_X2 \AES_ENC/u0/U135  ( .A1(\AES_ENC/u0/n980 ), .A2(\AES_ENC/u0/n990 ),.ZN(\AES_ENC/u0/N267 ) );
NAND2_X2 \AES_ENC/u0/U133  ( .A1(\AES_ENC/u0/N211 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n970 ) );
NAND2_X2 \AES_ENC/u0/U132  ( .A1(\AES_ENC/u0/n960 ), .A2(\AES_ENC/u0/n970 ),.ZN(\AES_ENC/u0/N268 ) );
NAND2_X2 \AES_ENC/u0/U130  ( .A1(\AES_ENC/u0/N210 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n950 ) );
NAND2_X2 \AES_ENC/u0/U129  ( .A1(\AES_ENC/u0/n940 ), .A2(\AES_ENC/u0/n950 ),.ZN(\AES_ENC/u0/N269 ) );
NAND2_X2 \AES_ENC/u0/U127  ( .A1(\AES_ENC/u0/N209 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n930 ) );
NAND2_X2 \AES_ENC/u0/U126  ( .A1(\AES_ENC/u0/n920 ), .A2(\AES_ENC/u0/n930 ),.ZN(\AES_ENC/u0/N270 ) );
NAND2_X2 \AES_ENC/u0/U124  ( .A1(\AES_ENC/u0/N208 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n910 ) );
NAND2_X2 \AES_ENC/u0/U123  ( .A1(\AES_ENC/u0/n900 ), .A2(\AES_ENC/u0/n910 ),.ZN(\AES_ENC/u0/N271 ) );
XOR2_X2 \AES_ENC/u0/U121  ( .A(\AES_ENC/w0[0] ), .B(\AES_ENC/u0/subword[0] ),.Z(\AES_ENC/u0/n890 ) );
NAND2_X2 \AES_ENC/u0/U120  ( .A1(\AES_ENC/u0/n890 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n880 ) );
NAND2_X2 \AES_ENC/u0/U119  ( .A1(\AES_ENC/u0/n870 ), .A2(\AES_ENC/u0/n880 ),.ZN(\AES_ENC/u0/N42 ) );
XOR2_X2 \AES_ENC/u0/U117  ( .A(\AES_ENC/w0[1] ), .B(\AES_ENC/u0/subword[1] ),.Z(\AES_ENC/u0/n860 ) );
NAND2_X2 \AES_ENC/u0/U116  ( .A1(\AES_ENC/u0/n860 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n850 ) );
NAND2_X2 \AES_ENC/u0/U115  ( .A1(\AES_ENC/u0/n840 ), .A2(\AES_ENC/u0/n850 ),.ZN(\AES_ENC/u0/N43 ) );
XOR2_X2 \AES_ENC/u0/U113  ( .A(\AES_ENC/w0[2] ), .B(\AES_ENC/u0/subword[2] ),.Z(\AES_ENC/u0/n830 ) );
NAND2_X2 \AES_ENC/u0/U112  ( .A1(\AES_ENC/u0/n830 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n820 ) );
NAND2_X2 \AES_ENC/u0/U111  ( .A1(\AES_ENC/u0/n810 ), .A2(\AES_ENC/u0/n820 ),.ZN(\AES_ENC/u0/N44 ) );
XOR2_X2 \AES_ENC/u0/U109  ( .A(\AES_ENC/w0[3] ), .B(\AES_ENC/u0/subword[3] ),.Z(\AES_ENC/u0/n800 ) );
NAND2_X2 \AES_ENC/u0/U108  ( .A1(\AES_ENC/u0/n800 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n790 ) );
NAND2_X2 \AES_ENC/u0/U107  ( .A1(\AES_ENC/u0/n780 ), .A2(\AES_ENC/u0/n790 ),.ZN(\AES_ENC/u0/N45 ) );
XOR2_X2 \AES_ENC/u0/U105  ( .A(\AES_ENC/w0[4] ), .B(\AES_ENC/u0/subword[4] ),.Z(\AES_ENC/u0/n770 ) );
NAND2_X2 \AES_ENC/u0/U104  ( .A1(\AES_ENC/u0/n770 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n760 ) );
NAND2_X2 \AES_ENC/u0/U103  ( .A1(\AES_ENC/u0/n75 ), .A2(\AES_ENC/u0/n760 ),.ZN(\AES_ENC/u0/N46 ) );
XOR2_X2 \AES_ENC/u0/U101  ( .A(\AES_ENC/w0[5] ), .B(\AES_ENC/u0/subword[5] ),.Z(\AES_ENC/u0/n74 ) );
NAND2_X2 \AES_ENC/u0/U100  ( .A1(\AES_ENC/u0/n74 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n730 ) );
NAND2_X2 \AES_ENC/u0/U99  ( .A1(\AES_ENC/u0/n720 ), .A2(\AES_ENC/u0/n730 ),.ZN(\AES_ENC/u0/N47 ) );
XOR2_X2 \AES_ENC/u0/U97  ( .A(\AES_ENC/w0[6] ), .B(\AES_ENC/u0/subword[6] ),.Z(\AES_ENC/u0/n710 ) );
NAND2_X2 \AES_ENC/u0/U96  ( .A1(\AES_ENC/u0/n710 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n700 ) );
NAND2_X2 \AES_ENC/u0/U95  ( .A1(\AES_ENC/u0/n690 ), .A2(\AES_ENC/u0/n700 ),.ZN(\AES_ENC/u0/N48 ) );
XOR2_X2 \AES_ENC/u0/U93  ( .A(\AES_ENC/w0[7] ), .B(\AES_ENC/u0/subword[7] ),.Z(\AES_ENC/u0/n680 ) );
NAND2_X2 \AES_ENC/u0/U92  ( .A1(\AES_ENC/u0/n680 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n670 ) );
NAND2_X2 \AES_ENC/u0/U91  ( .A1(\AES_ENC/u0/n660 ), .A2(\AES_ENC/u0/n670 ),.ZN(\AES_ENC/u0/N49 ) );
XOR2_X2 \AES_ENC/u0/U89  ( .A(\AES_ENC/w0[8] ), .B(\AES_ENC/u0/subword[8] ),.Z(\AES_ENC/u0/n650 ) );
NAND2_X2 \AES_ENC/u0/U88  ( .A1(\AES_ENC/u0/n650 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n640 ) );
NAND2_X2 \AES_ENC/u0/U87  ( .A1(\AES_ENC/u0/n630 ), .A2(\AES_ENC/u0/n640 ),.ZN(\AES_ENC/u0/N50 ) );
XOR2_X2 \AES_ENC/u0/U85  ( .A(\AES_ENC/w0[9] ), .B(\AES_ENC/u0/subword[9] ),.Z(\AES_ENC/u0/n620 ) );
NAND2_X2 \AES_ENC/u0/U84  ( .A1(\AES_ENC/u0/n620 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n610 ) );
NAND2_X2 \AES_ENC/u0/U83  ( .A1(\AES_ENC/u0/n600 ), .A2(\AES_ENC/u0/n610 ),.ZN(\AES_ENC/u0/N51 ) );
XOR2_X2 \AES_ENC/u0/U81  ( .A(\AES_ENC/w0[10] ), .B(\AES_ENC/u0/subword[10] ), .Z(\AES_ENC/u0/n590 ) );
NAND2_X2 \AES_ENC/u0/U80  ( .A1(\AES_ENC/u0/n590 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n580 ) );
NAND2_X2 \AES_ENC/u0/U79  ( .A1(\AES_ENC/u0/n570 ), .A2(\AES_ENC/u0/n580 ),.ZN(\AES_ENC/u0/N52 ) );
XOR2_X2 \AES_ENC/u0/U77  ( .A(\AES_ENC/w0[11] ), .B(\AES_ENC/u0/subword[11] ), .Z(\AES_ENC/u0/n560 ) );
NAND2_X2 \AES_ENC/u0/U76  ( .A1(\AES_ENC/u0/n560 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n550 ) );
NAND2_X2 \AES_ENC/u0/U75  ( .A1(\AES_ENC/u0/n540 ), .A2(\AES_ENC/u0/n550 ),.ZN(\AES_ENC/u0/N53 ) );
XOR2_X2 \AES_ENC/u0/U73  ( .A(\AES_ENC/w0[12] ), .B(\AES_ENC/u0/subword[12] ), .Z(\AES_ENC/u0/n530 ) );
NAND2_X2 \AES_ENC/u0/U72  ( .A1(\AES_ENC/u0/n530 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n520 ) );
NAND2_X2 \AES_ENC/u0/U71  ( .A1(\AES_ENC/u0/n510 ), .A2(\AES_ENC/u0/n520 ),.ZN(\AES_ENC/u0/N54 ) );
XOR2_X2 \AES_ENC/u0/U69  ( .A(\AES_ENC/w0[13] ), .B(\AES_ENC/u0/subword[13] ), .Z(\AES_ENC/u0/n500 ) );
NAND2_X2 \AES_ENC/u0/U68  ( .A1(\AES_ENC/u0/n500 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n490 ) );
NAND2_X2 \AES_ENC/u0/U67  ( .A1(\AES_ENC/u0/n480 ), .A2(\AES_ENC/u0/n490 ),.ZN(\AES_ENC/u0/N55 ) );
XOR2_X2 \AES_ENC/u0/U65  ( .A(\AES_ENC/w0[14] ), .B(\AES_ENC/u0/subword[14] ), .Z(\AES_ENC/u0/n470 ) );
NAND2_X2 \AES_ENC/u0/U64  ( .A1(\AES_ENC/u0/n470 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n460 ) );
NAND2_X2 \AES_ENC/u0/U63  ( .A1(\AES_ENC/u0/n450 ), .A2(\AES_ENC/u0/n460 ),.ZN(\AES_ENC/u0/N56 ) );
XOR2_X2 \AES_ENC/u0/U61  ( .A(\AES_ENC/w0[15] ), .B(\AES_ENC/u0/subword[15] ), .Z(\AES_ENC/u0/n440 ) );
NAND2_X2 \AES_ENC/u0/U60  ( .A1(\AES_ENC/u0/n440 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n430 ) );
NAND2_X2 \AES_ENC/u0/U59  ( .A1(\AES_ENC/u0/n420 ), .A2(\AES_ENC/u0/n430 ),.ZN(\AES_ENC/u0/N57 ) );
XOR2_X2 \AES_ENC/u0/U57  ( .A(\AES_ENC/w0[16] ), .B(\AES_ENC/u0/subword[16] ), .Z(\AES_ENC/u0/n41 ) );
NAND2_X2 \AES_ENC/u0/U56  ( .A1(\AES_ENC/u0/n41 ), .A2(\AES_ENC/u0/n324 ),.ZN(\AES_ENC/u0/n40 ) );
NAND2_X2 \AES_ENC/u0/U55  ( .A1(\AES_ENC/u0/n39 ), .A2(\AES_ENC/u0/n40 ),.ZN(\AES_ENC/u0/N58 ) );
XOR2_X2 \AES_ENC/u0/U53  ( .A(\AES_ENC/w0[17] ), .B(\AES_ENC/u0/subword[17] ), .Z(\AES_ENC/u0/n38 ) );
NAND2_X2 \AES_ENC/u0/U52  ( .A1(\AES_ENC/u0/n38 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n37 ) );
NAND2_X2 \AES_ENC/u0/U51  ( .A1(\AES_ENC/u0/n36 ), .A2(\AES_ENC/u0/n37 ),.ZN(\AES_ENC/u0/N59 ) );
XOR2_X2 \AES_ENC/u0/U49  ( .A(\AES_ENC/w0[18] ), .B(\AES_ENC/u0/subword[18] ), .Z(\AES_ENC/u0/n35 ) );
NAND2_X2 \AES_ENC/u0/U48  ( .A1(\AES_ENC/u0/n35 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n34 ) );
NAND2_X2 \AES_ENC/u0/U47  ( .A1(\AES_ENC/u0/n33 ), .A2(\AES_ENC/u0/n34 ),.ZN(\AES_ENC/u0/N60 ) );
XOR2_X2 \AES_ENC/u0/U45  ( .A(\AES_ENC/w0[19] ), .B(\AES_ENC/u0/subword[19] ), .Z(\AES_ENC/u0/n32 ) );
NAND2_X2 \AES_ENC/u0/U44  ( .A1(\AES_ENC/u0/n32 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n31 ) );
NAND2_X2 \AES_ENC/u0/U43  ( .A1(\AES_ENC/u0/n30 ), .A2(\AES_ENC/u0/n31 ),.ZN(\AES_ENC/u0/N61 ) );
XOR2_X2 \AES_ENC/u0/U41  ( .A(\AES_ENC/w0[20] ), .B(\AES_ENC/u0/subword[20] ), .Z(\AES_ENC/u0/n29 ) );
NAND2_X2 \AES_ENC/u0/U40  ( .A1(\AES_ENC/u0/n29 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n28 ) );
NAND2_X2 \AES_ENC/u0/U39  ( .A1(\AES_ENC/u0/n27 ), .A2(\AES_ENC/u0/n28 ),.ZN(\AES_ENC/u0/N62 ) );
XOR2_X2 \AES_ENC/u0/U37  ( .A(\AES_ENC/w0[21] ), .B(\AES_ENC/u0/subword[21] ), .Z(\AES_ENC/u0/n26 ) );
NAND2_X2 \AES_ENC/u0/U36  ( .A1(\AES_ENC/u0/n26 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n25 ) );
NAND2_X2 \AES_ENC/u0/U35  ( .A1(\AES_ENC/u0/n24 ), .A2(\AES_ENC/u0/n25 ),.ZN(\AES_ENC/u0/N63 ) );
XOR2_X2 \AES_ENC/u0/U33  ( .A(\AES_ENC/w0[22] ), .B(\AES_ENC/u0/subword[22] ), .Z(\AES_ENC/u0/n23 ) );
NAND2_X2 \AES_ENC/u0/U32  ( .A1(\AES_ENC/u0/n23 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n22 ) );
NAND2_X2 \AES_ENC/u0/U31  ( .A1(\AES_ENC/u0/n21 ), .A2(\AES_ENC/u0/n22 ),.ZN(\AES_ENC/u0/N64 ) );
XOR2_X2 \AES_ENC/u0/U29  ( .A(\AES_ENC/w0[23] ), .B(\AES_ENC/u0/subword[23] ), .Z(\AES_ENC/u0/n20 ) );
NAND2_X2 \AES_ENC/u0/U28  ( .A1(\AES_ENC/u0/n20 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n19 ) );
NAND2_X2 \AES_ENC/u0/U27  ( .A1(\AES_ENC/u0/n18 ), .A2(\AES_ENC/u0/n19 ),.ZN(\AES_ENC/u0/N65 ) );
NAND2_X2 \AES_ENC/u0/U25  ( .A1(\AES_ENC/u0/N17 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n1710 ) );
NAND2_X2 \AES_ENC/u0/U24  ( .A1(\AES_ENC/u0/n1610 ), .A2(\AES_ENC/u0/n1710 ),.ZN(\AES_ENC/u0/N66 ) );
NAND2_X2 \AES_ENC/u0/U22  ( .A1(\AES_ENC/u0/N16 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n1510 ) );
NAND2_X2 \AES_ENC/u0/U21  ( .A1(\AES_ENC/u0/n1400 ), .A2(\AES_ENC/u0/n1510 ),.ZN(\AES_ENC/u0/N67 ) );
NAND2_X2 \AES_ENC/u0/U19  ( .A1(\AES_ENC/u0/N15 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n1310 ) );
NAND2_X2 \AES_ENC/u0/U18  ( .A1(\AES_ENC/u0/n1210 ), .A2(\AES_ENC/u0/n1310 ),.ZN(\AES_ENC/u0/N68 ) );
NAND2_X2 \AES_ENC/u0/U16  ( .A1(\AES_ENC/u0/N14 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n1110 ) );
NAND2_X2 \AES_ENC/u0/U15  ( .A1(\AES_ENC/u0/n1010 ), .A2(\AES_ENC/u0/n1110 ),.ZN(\AES_ENC/u0/N69 ) );
NAND2_X2 \AES_ENC/u0/U13  ( .A1(\AES_ENC/u0/N13 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n9 ) );
NAND2_X2 \AES_ENC/u0/U12  ( .A1(\AES_ENC/u0/n8 ), .A2(\AES_ENC/u0/n9 ), .ZN(\AES_ENC/u0/N70 ) );
NAND2_X2 \AES_ENC/u0/U10  ( .A1(\AES_ENC/u0/N12 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n7 ) );
NAND2_X2 \AES_ENC/u0/U9  ( .A1(\AES_ENC/u0/n6 ), .A2(\AES_ENC/u0/n7 ), .ZN(\AES_ENC/u0/N71 ) );
NAND2_X2 \AES_ENC/u0/U7  ( .A1(\AES_ENC/u0/N11 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n5 ) );
NAND2_X2 \AES_ENC/u0/U6  ( .A1(\AES_ENC/u0/n4 ), .A2(\AES_ENC/u0/n5 ), .ZN(\AES_ENC/u0/N72 ) );
NAND2_X2 \AES_ENC/u0/U4  ( .A1(\AES_ENC/u0/N10 ), .A2(\AES_ENC/u0/n325 ),.ZN(\AES_ENC/u0/n3 ) );
DFF_X2 \AES_ENC/u0/w_reg_1__0_  ( .D(\AES_ENC/u0/N108 ), .CK(clk), .Q(\AES_ENC/w1[0] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__0_  ( .D(\AES_ENC/u0/N174 ), .CK(clk), .Q(\AES_ENC/w2[0] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__15_  ( .D(\AES_ENC/u0/N123 ), .CK(clk), .Q(\AES_ENC/w1[15] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__15_  ( .D(\AES_ENC/u0/N189 ), .CK(clk), .Q(\AES_ENC/w2[15] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__23_  ( .D(\AES_ENC/u0/N131 ), .CK(clk), .Q(\AES_ENC/w1[23] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__23_  ( .D(\AES_ENC/u0/N197 ), .CK(clk), .Q(\AES_ENC/w2[23] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__31_  ( .D(\AES_ENC/u0/n314 ), .CK(clk), .Q(\AES_ENC/w0[31] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__31_  ( .D(\AES_ENC/u0/N139 ), .CK(clk), .Q(\AES_ENC/w1[31] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__31_  ( .D(\AES_ENC/u0/N205 ), .CK(clk), .Q(\AES_ENC/w2[31] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__7_  ( .D(\AES_ENC/u0/N115 ), .CK(clk), .Q(\AES_ENC/w1[7] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__7_  ( .D(\AES_ENC/u0/N181 ), .CK(clk), .Q(\AES_ENC/w2[7] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__7_  ( .D(\AES_ENC/u0/N247 ), .CK(clk), .Q(\AES_ENC/w3[7] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__7_  ( .D(\AES_ENC/u0/N49 ), .CK(clk), .Q(\AES_ENC/w0[7] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__6_  ( .D(\AES_ENC/u0/N114 ), .CK(clk), .Q(\AES_ENC/w1[6] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__6_  ( .D(\AES_ENC/u0/N180 ), .CK(clk), .Q(\AES_ENC/w2[6] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__6_  ( .D(\AES_ENC/u0/N246 ), .CK(clk), .Q(\AES_ENC/w3[6] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__6_  ( .D(\AES_ENC/u0/N48 ), .CK(clk), .Q(\AES_ENC/w0[6] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__5_  ( .D(\AES_ENC/u0/N113 ), .CK(clk), .Q(\AES_ENC/w1[5] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__5_  ( .D(\AES_ENC/u0/N179 ), .CK(clk), .Q(\AES_ENC/w2[5] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__5_  ( .D(\AES_ENC/u0/N245 ), .CK(clk), .Q(\AES_ENC/w3[5] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__5_  ( .D(\AES_ENC/u0/N47 ), .CK(clk), .Q(\AES_ENC/w0[5] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__4_  ( .D(\AES_ENC/u0/N112 ), .CK(clk), .Q(\AES_ENC/w1[4] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__4_  ( .D(\AES_ENC/u0/N178 ), .CK(clk), .Q(\AES_ENC/w2[4] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__4_  ( .D(\AES_ENC/u0/N244 ), .CK(clk), .Q(\AES_ENC/w3[4] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__4_  ( .D(\AES_ENC/u0/N46 ), .CK(clk), .Q(\AES_ENC/w0[4] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__3_  ( .D(\AES_ENC/u0/N111 ), .CK(clk), .Q(\AES_ENC/w1[3] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__3_  ( .D(\AES_ENC/u0/N177 ), .CK(clk), .Q(\AES_ENC/w2[3] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__3_  ( .D(\AES_ENC/u0/N243 ), .CK(clk), .Q(\AES_ENC/w3[3] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__3_  ( .D(\AES_ENC/u0/N45 ), .CK(clk), .Q(\AES_ENC/w0[3] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__2_  ( .D(\AES_ENC/u0/N110 ), .CK(clk), .Q(\AES_ENC/w1[2] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__2_  ( .D(\AES_ENC/u0/N176 ), .CK(clk), .Q(\AES_ENC/w2[2] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__2_  ( .D(\AES_ENC/u0/N242 ), .CK(clk), .Q(\AES_ENC/w3[2] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__2_  ( .D(\AES_ENC/u0/N44 ), .CK(clk), .Q(\AES_ENC/w0[2] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__1_  ( .D(\AES_ENC/u0/N109 ), .CK(clk), .Q(\AES_ENC/w1[1] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__1_  ( .D(\AES_ENC/u0/N175 ), .CK(clk), .Q(\AES_ENC/w2[1] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__1_  ( .D(\AES_ENC/u0/N241 ), .CK(clk), .Q(\AES_ENC/w3[1] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__1_  ( .D(\AES_ENC/u0/N43 ), .CK(clk), .Q(\AES_ENC/w0[1] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__31_  ( .D(\AES_ENC/u0/N271 ), .CK(clk), .Q(\AES_ENC/w3[31] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__30_  ( .D(\AES_ENC/u0/N72 ), .CK(clk), .Q(\AES_ENC/w0[30] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__30_  ( .D(\AES_ENC/u0/N138 ), .CK(clk), .Q(\AES_ENC/w1[30] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__30_  ( .D(\AES_ENC/u0/N204 ), .CK(clk), .Q(\AES_ENC/w2[30] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__30_  ( .D(\AES_ENC/u0/N270 ), .CK(clk), .Q(\AES_ENC/w3[30] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__29_  ( .D(\AES_ENC/u0/N71 ), .CK(clk), .Q(\AES_ENC/w0[29] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__29_  ( .D(\AES_ENC/u0/N137 ), .CK(clk), .Q(\AES_ENC/w1[29] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__29_  ( .D(\AES_ENC/u0/N203 ), .CK(clk), .Q(\AES_ENC/w2[29] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__29_  ( .D(\AES_ENC/u0/N269 ), .CK(clk), .Q(\AES_ENC/w3[29] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__28_  ( .D(\AES_ENC/u0/N70 ), .CK(clk), .Q(\AES_ENC/w0[28] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__28_  ( .D(\AES_ENC/u0/N136 ), .CK(clk), .Q(\AES_ENC/w1[28] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__28_  ( .D(\AES_ENC/u0/N202 ), .CK(clk), .Q(\AES_ENC/w2[28] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__28_  ( .D(\AES_ENC/u0/N268 ), .CK(clk), .Q(\AES_ENC/w3[28] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__27_  ( .D(\AES_ENC/u0/N69 ), .CK(clk), .Q(\AES_ENC/w0[27] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__27_  ( .D(\AES_ENC/u0/N135 ), .CK(clk), .Q(\AES_ENC/w1[27] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__27_  ( .D(\AES_ENC/u0/N201 ), .CK(clk), .Q(\AES_ENC/w2[27] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__27_  ( .D(\AES_ENC/u0/N267 ), .CK(clk), .Q(\AES_ENC/w3[27] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__26_  ( .D(\AES_ENC/u0/N68 ), .CK(clk), .Q(\AES_ENC/w0[26] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__26_  ( .D(\AES_ENC/u0/N134 ), .CK(clk), .Q(\AES_ENC/w1[26] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__26_  ( .D(\AES_ENC/u0/N200 ), .CK(clk), .Q(\AES_ENC/w2[26] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__26_  ( .D(\AES_ENC/u0/N266 ), .CK(clk), .Q(\AES_ENC/w3[26] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__25_  ( .D(\AES_ENC/u0/N67 ), .CK(clk), .Q(\AES_ENC/w0[25] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__25_  ( .D(\AES_ENC/u0/N133 ), .CK(clk), .Q(\AES_ENC/w1[25] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__25_  ( .D(\AES_ENC/u0/N199 ), .CK(clk), .Q(\AES_ENC/w2[25] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__25_  ( .D(\AES_ENC/u0/N265 ), .CK(clk), .Q(\AES_ENC/w3[25] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__24_  ( .D(\AES_ENC/u0/N66 ), .CK(clk), .Q(\AES_ENC/w0[24] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__24_  ( .D(\AES_ENC/u0/N132 ), .CK(clk), .Q(\AES_ENC/w1[24] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__24_  ( .D(\AES_ENC/u0/N198 ), .CK(clk), .Q(\AES_ENC/w2[24] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__24_  ( .D(\AES_ENC/u0/N264 ), .CK(clk), .Q(\AES_ENC/w3[24] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__23_  ( .D(\AES_ENC/u0/N263 ), .CK(clk), .Q(\AES_ENC/w3[23] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__23_  ( .D(\AES_ENC/u0/N65 ), .CK(clk), .Q(\AES_ENC/w0[23] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__22_  ( .D(\AES_ENC/u0/N130 ), .CK(clk), .Q(\AES_ENC/w1[22] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__22_  ( .D(\AES_ENC/u0/N196 ), .CK(clk), .Q(\AES_ENC/w2[22] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__22_  ( .D(\AES_ENC/u0/N262 ), .CK(clk), .Q(\AES_ENC/w3[22] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__22_  ( .D(\AES_ENC/u0/N64 ), .CK(clk), .Q(\AES_ENC/w0[22] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__21_  ( .D(\AES_ENC/u0/N129 ), .CK(clk), .Q(\AES_ENC/w1[21] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__21_  ( .D(\AES_ENC/u0/N195 ), .CK(clk), .Q(\AES_ENC/w2[21] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__21_  ( .D(\AES_ENC/u0/N261 ), .CK(clk), .Q(\AES_ENC/w3[21] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__21_  ( .D(\AES_ENC/u0/N63 ), .CK(clk), .Q(\AES_ENC/w0[21] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__20_  ( .D(\AES_ENC/u0/N128 ), .CK(clk), .Q(\AES_ENC/w1[20] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__20_  ( .D(\AES_ENC/u0/N194 ), .CK(clk), .Q(\AES_ENC/w2[20] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__20_  ( .D(\AES_ENC/u0/N260 ), .CK(clk), .Q(\AES_ENC/w3[20] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__20_  ( .D(\AES_ENC/u0/N62 ), .CK(clk), .Q(\AES_ENC/w0[20] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__19_  ( .D(\AES_ENC/u0/N127 ), .CK(clk), .Q(\AES_ENC/w1[19] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__19_  ( .D(\AES_ENC/u0/N193 ), .CK(clk), .Q(\AES_ENC/w2[19] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__19_  ( .D(\AES_ENC/u0/N259 ), .CK(clk), .Q(\AES_ENC/w3[19] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__19_  ( .D(\AES_ENC/u0/N61 ), .CK(clk), .Q(\AES_ENC/w0[19] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__18_  ( .D(\AES_ENC/u0/N126 ), .CK(clk), .Q(\AES_ENC/w1[18] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__18_  ( .D(\AES_ENC/u0/N192 ), .CK(clk), .Q(\AES_ENC/w2[18] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__18_  ( .D(\AES_ENC/u0/N258 ), .CK(clk), .Q(\AES_ENC/w3[18] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__18_  ( .D(\AES_ENC/u0/N60 ), .CK(clk), .Q(\AES_ENC/w0[18] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__17_  ( .D(\AES_ENC/u0/N125 ), .CK(clk), .Q(\AES_ENC/w1[17] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__17_  ( .D(\AES_ENC/u0/N191 ), .CK(clk), .Q(\AES_ENC/w2[17] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__17_  ( .D(\AES_ENC/u0/N257 ), .CK(clk), .Q(\AES_ENC/w3[17] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__17_  ( .D(\AES_ENC/u0/N59 ), .CK(clk), .Q(\AES_ENC/w0[17] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__16_  ( .D(\AES_ENC/u0/N124 ), .CK(clk), .Q(\AES_ENC/w1[16] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__16_  ( .D(\AES_ENC/u0/N190 ), .CK(clk), .Q(\AES_ENC/w2[16] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__16_  ( .D(\AES_ENC/u0/N256 ), .CK(clk), .Q(\AES_ENC/w3[16] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__16_  ( .D(\AES_ENC/u0/N58 ), .CK(clk), .Q(\AES_ENC/w0[16] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__15_  ( .D(\AES_ENC/u0/N255 ), .CK(clk), .Q(\AES_ENC/w3[15] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__15_  ( .D(\AES_ENC/u0/N57 ), .CK(clk), .Q(\AES_ENC/w0[15] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__14_  ( .D(\AES_ENC/u0/N122 ), .CK(clk), .Q(\AES_ENC/w1[14] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__14_  ( .D(\AES_ENC/u0/N188 ), .CK(clk), .Q(\AES_ENC/w2[14] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__14_  ( .D(\AES_ENC/u0/N254 ), .CK(clk), .Q(\AES_ENC/w3[14] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__14_  ( .D(\AES_ENC/u0/N56 ), .CK(clk), .Q(\AES_ENC/w0[14] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__13_  ( .D(\AES_ENC/u0/N121 ), .CK(clk), .Q(\AES_ENC/w1[13] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__13_  ( .D(\AES_ENC/u0/N187 ), .CK(clk), .Q(\AES_ENC/w2[13] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__13_  ( .D(\AES_ENC/u0/N253 ), .CK(clk), .Q(\AES_ENC/w3[13] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__13_  ( .D(\AES_ENC/u0/N55 ), .CK(clk), .Q(\AES_ENC/w0[13] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__12_  ( .D(\AES_ENC/u0/N120 ), .CK(clk), .Q(\AES_ENC/w1[12] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__12_  ( .D(\AES_ENC/u0/N186 ), .CK(clk), .Q(\AES_ENC/w2[12] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__12_  ( .D(\AES_ENC/u0/N252 ), .CK(clk), .Q(\AES_ENC/w3[12] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__12_  ( .D(\AES_ENC/u0/N54 ), .CK(clk), .Q(\AES_ENC/w0[12] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__11_  ( .D(\AES_ENC/u0/N119 ), .CK(clk), .Q(\AES_ENC/w1[11] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__11_  ( .D(\AES_ENC/u0/N185 ), .CK(clk), .Q(\AES_ENC/w2[11] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__11_  ( .D(\AES_ENC/u0/N251 ), .CK(clk), .Q(\AES_ENC/w3[11] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__11_  ( .D(\AES_ENC/u0/N53 ), .CK(clk), .Q(\AES_ENC/w0[11] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__10_  ( .D(\AES_ENC/u0/N118 ), .CK(clk), .Q(\AES_ENC/w1[10] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__10_  ( .D(\AES_ENC/u0/N184 ), .CK(clk), .Q(\AES_ENC/w2[10] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__10_  ( .D(\AES_ENC/u0/N250 ), .CK(clk), .Q(\AES_ENC/w3[10] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__10_  ( .D(\AES_ENC/u0/N52 ), .CK(clk), .Q(\AES_ENC/w0[10] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__9_  ( .D(\AES_ENC/u0/N117 ), .CK(clk), .Q(\AES_ENC/w1[9] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__9_  ( .D(\AES_ENC/u0/N183 ), .CK(clk), .Q(\AES_ENC/w2[9] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__9_  ( .D(\AES_ENC/u0/N249 ), .CK(clk), .Q(\AES_ENC/w3[9] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__9_  ( .D(\AES_ENC/u0/N51 ), .CK(clk), .Q(\AES_ENC/w0[9] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_1__8_  ( .D(\AES_ENC/u0/N116 ), .CK(clk), .Q(\AES_ENC/w1[8] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_2__8_  ( .D(\AES_ENC/u0/N182 ), .CK(clk), .Q(\AES_ENC/w2[8] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__8_  ( .D(\AES_ENC/u0/N248 ), .CK(clk), .Q(\AES_ENC/w3[8] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__8_  ( .D(\AES_ENC/u0/N50 ), .CK(clk), .Q(\AES_ENC/w0[8] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_3__0_  ( .D(\AES_ENC/u0/N240 ), .CK(clk), .Q(\AES_ENC/w3[0] ), .QN() );
DFF_X2 \AES_ENC/u0/w_reg_0__0_  ( .D(\AES_ENC/u0/N42 ), .CK(clk), .Q(\AES_ENC/w0[0] ), .QN() );
XOR2_X2 \AES_ENC/u0/U547  ( .A(\AES_ENC/u0/rcon [31]), .B(\AES_ENC/u0/n282 ),.Z(\AES_ENC/u0/N10 ) );
XOR2_X2 \AES_ENC/u0/U546  ( .A(\AES_ENC/w0[31] ), .B(\AES_ENC/u0/subword[31] ), .Z(\AES_ENC/u0/n282 ) );
XOR2_X2 \AES_ENC/u0/U545  ( .A(\AES_ENC/w1[31] ), .B(\AES_ENC/u0/N10 ), .Z(\AES_ENC/u0/N76 ) );
XOR2_X2 \AES_ENC/u0/U544  ( .A(\AES_ENC/w2[31] ), .B(\AES_ENC/u0/N76 ), .Z(\AES_ENC/u0/N142 ) );
XOR2_X2 \AES_ENC/u0/U543  ( .A(\AES_ENC/w3[31] ), .B(\AES_ENC/u0/N142 ), .Z(\AES_ENC/u0/N208 ) );
XOR2_X2 \AES_ENC/u0/U542  ( .A(\AES_ENC/u0/rcon [30]), .B(\AES_ENC/u0/n283 ),.Z(\AES_ENC/u0/N11 ) );
XOR2_X2 \AES_ENC/u0/U541  ( .A(\AES_ENC/w0[30] ), .B(\AES_ENC/u0/subword[30] ), .Z(\AES_ENC/u0/n283 ) );
XOR2_X2 \AES_ENC/u0/U540  ( .A(\AES_ENC/w1[30] ), .B(\AES_ENC/u0/N11 ), .Z(\AES_ENC/u0/N77 ) );
XOR2_X2 \AES_ENC/u0/U539  ( .A(\AES_ENC/w2[30] ), .B(\AES_ENC/u0/N77 ), .Z(\AES_ENC/u0/N143 ) );
XOR2_X2 \AES_ENC/u0/U538  ( .A(\AES_ENC/w3[30] ), .B(\AES_ENC/u0/N143 ), .Z(\AES_ENC/u0/N209 ) );
XOR2_X2 \AES_ENC/u0/U537  ( .A(\AES_ENC/u0/rcon [29]), .B(\AES_ENC/u0/n284 ),.Z(\AES_ENC/u0/N12 ) );
XOR2_X2 \AES_ENC/u0/U536  ( .A(\AES_ENC/w0[29] ), .B(\AES_ENC/u0/subword[29] ), .Z(\AES_ENC/u0/n284 ) );
XOR2_X2 \AES_ENC/u0/U535  ( .A(\AES_ENC/w1[29] ), .B(\AES_ENC/u0/N12 ), .Z(\AES_ENC/u0/N78 ) );
XOR2_X2 \AES_ENC/u0/U534  ( .A(\AES_ENC/w2[29] ), .B(\AES_ENC/u0/N78 ), .Z(\AES_ENC/u0/N144 ) );
XOR2_X2 \AES_ENC/u0/U533  ( .A(\AES_ENC/w3[29] ), .B(\AES_ENC/u0/N144 ), .Z(\AES_ENC/u0/N210 ) );
XOR2_X2 \AES_ENC/u0/U532  ( .A(\AES_ENC/u0/rcon [28]), .B(\AES_ENC/u0/n285 ),.Z(\AES_ENC/u0/N13 ) );
XOR2_X2 \AES_ENC/u0/U531  ( .A(\AES_ENC/w0[28] ), .B(\AES_ENC/u0/subword[28] ), .Z(\AES_ENC/u0/n285 ) );
XOR2_X2 \AES_ENC/u0/U530  ( .A(\AES_ENC/w1[28] ), .B(\AES_ENC/u0/N13 ), .Z(\AES_ENC/u0/N79 ) );
XOR2_X2 \AES_ENC/u0/U529  ( .A(\AES_ENC/w2[28] ), .B(\AES_ENC/u0/N79 ), .Z(\AES_ENC/u0/N145 ) );
XOR2_X2 \AES_ENC/u0/U528  ( .A(\AES_ENC/w3[28] ), .B(\AES_ENC/u0/N145 ), .Z(\AES_ENC/u0/N211 ) );
XOR2_X2 \AES_ENC/u0/U527  ( .A(\AES_ENC/u0/rcon [27]), .B(\AES_ENC/u0/n286 ),.Z(\AES_ENC/u0/N14 ) );
XOR2_X2 \AES_ENC/u0/U526  ( .A(\AES_ENC/w0[27] ), .B(\AES_ENC/u0/subword[27] ), .Z(\AES_ENC/u0/n286 ) );
XOR2_X2 \AES_ENC/u0/U525  ( .A(\AES_ENC/w1[27] ), .B(\AES_ENC/u0/N14 ), .Z(\AES_ENC/u0/N80 ) );
XOR2_X2 \AES_ENC/u0/U524  ( .A(\AES_ENC/w2[27] ), .B(\AES_ENC/u0/N80 ), .Z(\AES_ENC/u0/N146 ) );
XOR2_X2 \AES_ENC/u0/U523  ( .A(\AES_ENC/w3[27] ), .B(\AES_ENC/u0/N146 ), .Z(\AES_ENC/u0/N212 ) );
XOR2_X2 \AES_ENC/u0/U522  ( .A(\AES_ENC/u0/rcon [26]), .B(\AES_ENC/u0/n287 ),.Z(\AES_ENC/u0/N15 ) );
XOR2_X2 \AES_ENC/u0/U521  ( .A(\AES_ENC/w0[26] ), .B(\AES_ENC/u0/subword[26] ), .Z(\AES_ENC/u0/n287 ) );
XOR2_X2 \AES_ENC/u0/U520  ( .A(\AES_ENC/w1[26] ), .B(\AES_ENC/u0/N15 ), .Z(\AES_ENC/u0/N81 ) );
XOR2_X2 \AES_ENC/u0/U519  ( .A(\AES_ENC/w2[26] ), .B(\AES_ENC/u0/N81 ), .Z(\AES_ENC/u0/N147 ) );
XOR2_X2 \AES_ENC/u0/U518  ( .A(\AES_ENC/w3[26] ), .B(\AES_ENC/u0/N147 ), .Z(\AES_ENC/u0/N213 ) );
XOR2_X2 \AES_ENC/u0/U517  ( .A(\AES_ENC/u0/rcon [25]), .B(\AES_ENC/u0/n288 ),.Z(\AES_ENC/u0/N16 ) );
XOR2_X2 \AES_ENC/u0/U516  ( .A(\AES_ENC/w0[25] ), .B(\AES_ENC/u0/subword[25] ), .Z(\AES_ENC/u0/n288 ) );
XOR2_X2 \AES_ENC/u0/U515  ( .A(\AES_ENC/w1[25] ), .B(\AES_ENC/u0/N16 ), .Z(\AES_ENC/u0/N82 ) );
XOR2_X2 \AES_ENC/u0/U514  ( .A(\AES_ENC/w2[25] ), .B(\AES_ENC/u0/N82 ), .Z(\AES_ENC/u0/N148 ) );
XOR2_X2 \AES_ENC/u0/U513  ( .A(\AES_ENC/w3[25] ), .B(\AES_ENC/u0/N148 ), .Z(\AES_ENC/u0/N214 ) );
XOR2_X2 \AES_ENC/u0/U512  ( .A(\AES_ENC/u0/rcon [24]), .B(\AES_ENC/u0/n289 ),.Z(\AES_ENC/u0/N17 ) );
XOR2_X2 \AES_ENC/u0/U511  ( .A(\AES_ENC/w0[24] ), .B(\AES_ENC/u0/subword[24] ), .Z(\AES_ENC/u0/n289 ) );
XOR2_X2 \AES_ENC/u0/U510  ( .A(\AES_ENC/w1[24] ), .B(\AES_ENC/u0/N17 ), .Z(\AES_ENC/u0/N83 ) );
XOR2_X2 \AES_ENC/u0/U509  ( .A(\AES_ENC/w2[24] ), .B(\AES_ENC/u0/N83 ), .Z(\AES_ENC/u0/N149 ) );
XOR2_X2 \AES_ENC/u0/U508  ( .A(\AES_ENC/w3[24] ), .B(\AES_ENC/u0/N149 ), .Z(\AES_ENC/u0/N215 ) );
XOR2_X2 \AES_ENC/u0/U507  ( .A(\AES_ENC/u0/subword[23] ), .B(\AES_ENC/u0/n290 ), .Z(\AES_ENC/u0/N84 ) );
XOR2_X2 \AES_ENC/u0/U506  ( .A(\AES_ENC/w1[23] ), .B(\AES_ENC/w0[23] ), .Z(\AES_ENC/u0/n290 ) );
XOR2_X2 \AES_ENC/u0/U505  ( .A(\AES_ENC/w2[23] ), .B(\AES_ENC/u0/N84 ), .Z(\AES_ENC/u0/N150 ) );
XOR2_X2 \AES_ENC/u0/U504  ( .A(\AES_ENC/w3[23] ), .B(\AES_ENC/u0/N150 ), .Z(\AES_ENC/u0/N216 ) );
XOR2_X2 \AES_ENC/u0/U503  ( .A(\AES_ENC/u0/subword[22] ), .B(\AES_ENC/u0/n291 ), .Z(\AES_ENC/u0/N85 ) );
XOR2_X2 \AES_ENC/u0/U502  ( .A(\AES_ENC/w1[22] ), .B(\AES_ENC/w0[22] ), .Z(\AES_ENC/u0/n291 ) );
XOR2_X2 \AES_ENC/u0/U501  ( .A(\AES_ENC/w2[22] ), .B(\AES_ENC/u0/N85 ), .Z(\AES_ENC/u0/N151 ) );
XOR2_X2 \AES_ENC/u0/U500  ( .A(\AES_ENC/w3[22] ), .B(\AES_ENC/u0/N151 ), .Z(\AES_ENC/u0/N217 ) );
XOR2_X2 \AES_ENC/u0/U499  ( .A(\AES_ENC/u0/subword[21] ), .B(\AES_ENC/u0/n292 ), .Z(\AES_ENC/u0/N86 ) );
XOR2_X2 \AES_ENC/u0/U498  ( .A(\AES_ENC/w1[21] ), .B(\AES_ENC/w0[21] ), .Z(\AES_ENC/u0/n292 ) );
XOR2_X2 \AES_ENC/u0/U497  ( .A(\AES_ENC/w2[21] ), .B(\AES_ENC/u0/N86 ), .Z(\AES_ENC/u0/N152 ) );
XOR2_X2 \AES_ENC/u0/U496  ( .A(\AES_ENC/w3[21] ), .B(\AES_ENC/u0/N152 ), .Z(\AES_ENC/u0/N218 ) );
XOR2_X2 \AES_ENC/u0/U495  ( .A(\AES_ENC/u0/subword[20] ), .B(\AES_ENC/u0/n293 ), .Z(\AES_ENC/u0/N87 ) );
XOR2_X2 \AES_ENC/u0/U494  ( .A(\AES_ENC/w1[20] ), .B(\AES_ENC/w0[20] ), .Z(\AES_ENC/u0/n293 ) );
XOR2_X2 \AES_ENC/u0/U493  ( .A(\AES_ENC/w2[20] ), .B(\AES_ENC/u0/N87 ), .Z(\AES_ENC/u0/N153 ) );
XOR2_X2 \AES_ENC/u0/U492  ( .A(\AES_ENC/w3[20] ), .B(\AES_ENC/u0/N153 ), .Z(\AES_ENC/u0/N219 ) );
XOR2_X2 \AES_ENC/u0/U491  ( .A(\AES_ENC/u0/subword[19] ), .B(\AES_ENC/u0/n294 ), .Z(\AES_ENC/u0/N88 ) );
XOR2_X2 \AES_ENC/u0/U490  ( .A(\AES_ENC/w1[19] ), .B(\AES_ENC/w0[19] ), .Z(\AES_ENC/u0/n294 ) );
XOR2_X2 \AES_ENC/u0/U489  ( .A(\AES_ENC/w2[19] ), .B(\AES_ENC/u0/N88 ), .Z(\AES_ENC/u0/N154 ) );
XOR2_X2 \AES_ENC/u0/U488  ( .A(\AES_ENC/w3[19] ), .B(\AES_ENC/u0/N154 ), .Z(\AES_ENC/u0/N220 ) );
XOR2_X2 \AES_ENC/u0/U487  ( .A(\AES_ENC/u0/subword[18] ), .B(\AES_ENC/u0/n295 ), .Z(\AES_ENC/u0/N89 ) );
XOR2_X2 \AES_ENC/u0/U486  ( .A(\AES_ENC/w1[18] ), .B(\AES_ENC/w0[18] ), .Z(\AES_ENC/u0/n295 ) );
XOR2_X2 \AES_ENC/u0/U485  ( .A(\AES_ENC/w2[18] ), .B(\AES_ENC/u0/N89 ), .Z(\AES_ENC/u0/N155 ) );
XOR2_X2 \AES_ENC/u0/U484  ( .A(\AES_ENC/w3[18] ), .B(\AES_ENC/u0/N155 ), .Z(\AES_ENC/u0/N221 ) );
XOR2_X2 \AES_ENC/u0/U483  ( .A(\AES_ENC/u0/subword[17] ), .B(\AES_ENC/u0/n296 ), .Z(\AES_ENC/u0/N90 ) );
XOR2_X2 \AES_ENC/u0/U482  ( .A(\AES_ENC/w1[17] ), .B(\AES_ENC/w0[17] ), .Z(\AES_ENC/u0/n296 ) );
XOR2_X2 \AES_ENC/u0/U481  ( .A(\AES_ENC/w2[17] ), .B(\AES_ENC/u0/N90 ), .Z(\AES_ENC/u0/N156 ) );
XOR2_X2 \AES_ENC/u0/U480  ( .A(\AES_ENC/w3[17] ), .B(\AES_ENC/u0/N156 ), .Z(\AES_ENC/u0/N222 ) );
XOR2_X2 \AES_ENC/u0/U479  ( .A(\AES_ENC/u0/subword[16] ), .B(\AES_ENC/u0/n297 ), .Z(\AES_ENC/u0/N91 ) );
XOR2_X2 \AES_ENC/u0/U478  ( .A(\AES_ENC/w1[16] ), .B(\AES_ENC/w0[16] ), .Z(\AES_ENC/u0/n297 ) );
XOR2_X2 \AES_ENC/u0/U477  ( .A(\AES_ENC/w2[16] ), .B(\AES_ENC/u0/N91 ), .Z(\AES_ENC/u0/N157 ) );
XOR2_X2 \AES_ENC/u0/U476  ( .A(\AES_ENC/w3[16] ), .B(\AES_ENC/u0/N157 ), .Z(\AES_ENC/u0/N223 ) );
XOR2_X2 \AES_ENC/u0/U475  ( .A(\AES_ENC/u0/subword[15] ), .B(\AES_ENC/u0/n298 ), .Z(\AES_ENC/u0/N92 ) );
XOR2_X2 \AES_ENC/u0/U474  ( .A(\AES_ENC/w1[15] ), .B(\AES_ENC/w0[15] ), .Z(\AES_ENC/u0/n298 ) );
XOR2_X2 \AES_ENC/u0/U473  ( .A(\AES_ENC/w2[15] ), .B(\AES_ENC/u0/N92 ), .Z(\AES_ENC/u0/N158 ) );
XOR2_X2 \AES_ENC/u0/U472  ( .A(\AES_ENC/w3[15] ), .B(\AES_ENC/u0/N158 ), .Z(\AES_ENC/u0/N224 ) );
XOR2_X2 \AES_ENC/u0/U471  ( .A(\AES_ENC/u0/subword[14] ), .B(\AES_ENC/u0/n299 ), .Z(\AES_ENC/u0/N93 ) );
XOR2_X2 \AES_ENC/u0/U470  ( .A(\AES_ENC/w1[14] ), .B(\AES_ENC/w0[14] ), .Z(\AES_ENC/u0/n299 ) );
XOR2_X2 \AES_ENC/u0/U469  ( .A(\AES_ENC/w2[14] ), .B(\AES_ENC/u0/N93 ), .Z(\AES_ENC/u0/N159 ) );
XOR2_X2 \AES_ENC/u0/U468  ( .A(\AES_ENC/w3[14] ), .B(\AES_ENC/u0/N159 ), .Z(\AES_ENC/u0/N225 ) );
XOR2_X2 \AES_ENC/u0/U467  ( .A(\AES_ENC/u0/subword[13] ), .B(\AES_ENC/u0/n300 ), .Z(\AES_ENC/u0/N94 ) );
XOR2_X2 \AES_ENC/u0/U466  ( .A(\AES_ENC/w1[13] ), .B(\AES_ENC/w0[13] ), .Z(\AES_ENC/u0/n300 ) );
XOR2_X2 \AES_ENC/u0/U465  ( .A(\AES_ENC/w2[13] ), .B(\AES_ENC/u0/N94 ), .Z(\AES_ENC/u0/N160 ) );
XOR2_X2 \AES_ENC/u0/U464  ( .A(\AES_ENC/w3[13] ), .B(\AES_ENC/u0/N160 ), .Z(\AES_ENC/u0/N226 ) );
XOR2_X2 \AES_ENC/u0/U463  ( .A(\AES_ENC/u0/subword[12] ), .B(\AES_ENC/u0/n301 ), .Z(\AES_ENC/u0/N95 ) );
XOR2_X2 \AES_ENC/u0/U462  ( .A(\AES_ENC/w1[12] ), .B(\AES_ENC/w0[12] ), .Z(\AES_ENC/u0/n301 ) );
XOR2_X2 \AES_ENC/u0/U461  ( .A(\AES_ENC/w2[12] ), .B(\AES_ENC/u0/N95 ), .Z(\AES_ENC/u0/N161 ) );
XOR2_X2 \AES_ENC/u0/U460  ( .A(\AES_ENC/w3[12] ), .B(\AES_ENC/u0/N161 ), .Z(\AES_ENC/u0/N227 ) );
XOR2_X2 \AES_ENC/u0/U459  ( .A(\AES_ENC/u0/subword[11] ), .B(\AES_ENC/u0/n302 ), .Z(\AES_ENC/u0/N96 ) );
XOR2_X2 \AES_ENC/u0/U458  ( .A(\AES_ENC/w1[11] ), .B(\AES_ENC/w0[11] ), .Z(\AES_ENC/u0/n302 ) );
XOR2_X2 \AES_ENC/u0/U457  ( .A(\AES_ENC/w2[11] ), .B(\AES_ENC/u0/N96 ), .Z(\AES_ENC/u0/N162 ) );
XOR2_X2 \AES_ENC/u0/U456  ( .A(\AES_ENC/w3[11] ), .B(\AES_ENC/u0/N162 ), .Z(\AES_ENC/u0/N228 ) );
XOR2_X2 \AES_ENC/u0/U455  ( .A(\AES_ENC/u0/subword[10] ), .B(\AES_ENC/u0/n303 ), .Z(\AES_ENC/u0/N97 ) );
XOR2_X2 \AES_ENC/u0/U454  ( .A(\AES_ENC/w1[10] ), .B(\AES_ENC/w0[10] ), .Z(\AES_ENC/u0/n303 ) );
XOR2_X2 \AES_ENC/u0/U453  ( .A(\AES_ENC/w2[10] ), .B(\AES_ENC/u0/N97 ), .Z(\AES_ENC/u0/N163 ) );
XOR2_X2 \AES_ENC/u0/U452  ( .A(\AES_ENC/w3[10] ), .B(\AES_ENC/u0/N163 ), .Z(\AES_ENC/u0/N229 ) );
XOR2_X2 \AES_ENC/u0/U451  ( .A(\AES_ENC/u0/subword[9] ), .B(\AES_ENC/u0/n304 ), .Z(\AES_ENC/u0/N98 ) );
XOR2_X2 \AES_ENC/u0/U450  ( .A(\AES_ENC/w1[9] ), .B(\AES_ENC/w0[9] ), .Z(\AES_ENC/u0/n304 ) );
XOR2_X2 \AES_ENC/u0/U449  ( .A(\AES_ENC/w2[9] ), .B(\AES_ENC/u0/N98 ), .Z(\AES_ENC/u0/N164 ) );
XOR2_X2 \AES_ENC/u0/U448  ( .A(\AES_ENC/w3[9] ), .B(\AES_ENC/u0/N164 ), .Z(\AES_ENC/u0/N230 ) );
XOR2_X2 \AES_ENC/u0/U447  ( .A(\AES_ENC/u0/subword[8] ), .B(\AES_ENC/u0/n305 ), .Z(\AES_ENC/u0/N99 ) );
XOR2_X2 \AES_ENC/u0/U446  ( .A(\AES_ENC/w1[8] ), .B(\AES_ENC/w0[8] ), .Z(\AES_ENC/u0/n305 ) );
XOR2_X2 \AES_ENC/u0/U445  ( .A(\AES_ENC/w2[8] ), .B(\AES_ENC/u0/N99 ), .Z(\AES_ENC/u0/N165 ) );
XOR2_X2 \AES_ENC/u0/U444  ( .A(\AES_ENC/w3[8] ), .B(\AES_ENC/u0/N165 ), .Z(\AES_ENC/u0/N231 ) );
XOR2_X2 \AES_ENC/u0/U443  ( .A(\AES_ENC/u0/subword[7] ), .B(\AES_ENC/u0/n306 ), .Z(\AES_ENC/u0/N100 ) );
XOR2_X2 \AES_ENC/u0/U442  ( .A(\AES_ENC/w1[7] ), .B(\AES_ENC/w0[7] ), .Z(\AES_ENC/u0/n306 ) );
XOR2_X2 \AES_ENC/u0/U441  ( .A(\AES_ENC/w2[7] ), .B(\AES_ENC/u0/N100 ), .Z(\AES_ENC/u0/N166 ) );
XOR2_X2 \AES_ENC/u0/U440  ( .A(\AES_ENC/w3[7] ), .B(\AES_ENC/u0/N166 ), .Z(\AES_ENC/u0/N232 ) );
XOR2_X2 \AES_ENC/u0/U439  ( .A(\AES_ENC/u0/subword[6] ), .B(\AES_ENC/u0/n307 ), .Z(\AES_ENC/u0/N101 ) );
XOR2_X2 \AES_ENC/u0/U438  ( .A(\AES_ENC/w1[6] ), .B(\AES_ENC/w0[6] ), .Z(\AES_ENC/u0/n307 ) );
XOR2_X2 \AES_ENC/u0/U437  ( .A(\AES_ENC/w2[6] ), .B(\AES_ENC/u0/N101 ), .Z(\AES_ENC/u0/N167 ) );
XOR2_X2 \AES_ENC/u0/U436  ( .A(\AES_ENC/w3[6] ), .B(\AES_ENC/u0/N167 ), .Z(\AES_ENC/u0/N233 ) );
XOR2_X2 \AES_ENC/u0/U435  ( .A(\AES_ENC/u0/subword[5] ), .B(\AES_ENC/u0/n308 ), .Z(\AES_ENC/u0/N102 ) );
XOR2_X2 \AES_ENC/u0/U434  ( .A(\AES_ENC/w1[5] ), .B(\AES_ENC/w0[5] ), .Z(\AES_ENC/u0/n308 ) );
XOR2_X2 \AES_ENC/u0/U433  ( .A(\AES_ENC/w2[5] ), .B(\AES_ENC/u0/N102 ), .Z(\AES_ENC/u0/N168 ) );
XOR2_X2 \AES_ENC/u0/U432  ( .A(\AES_ENC/w3[5] ), .B(\AES_ENC/u0/N168 ), .Z(\AES_ENC/u0/N234 ) );
XOR2_X2 \AES_ENC/u0/U431  ( .A(\AES_ENC/u0/subword[4] ), .B(\AES_ENC/u0/n309 ), .Z(\AES_ENC/u0/N103 ) );
XOR2_X2 \AES_ENC/u0/U430  ( .A(\AES_ENC/w1[4] ), .B(\AES_ENC/w0[4] ), .Z(\AES_ENC/u0/n309 ) );
XOR2_X2 \AES_ENC/u0/U429  ( .A(\AES_ENC/w2[4] ), .B(\AES_ENC/u0/N103 ), .Z(\AES_ENC/u0/N169 ) );
XOR2_X2 \AES_ENC/u0/U428  ( .A(\AES_ENC/w3[4] ), .B(\AES_ENC/u0/N169 ), .Z(\AES_ENC/u0/N235 ) );
XOR2_X2 \AES_ENC/u0/U427  ( .A(\AES_ENC/u0/subword[3] ), .B(\AES_ENC/u0/n310 ), .Z(\AES_ENC/u0/N104 ) );
XOR2_X2 \AES_ENC/u0/U426  ( .A(\AES_ENC/w1[3] ), .B(\AES_ENC/w0[3] ), .Z(\AES_ENC/u0/n310 ) );
XOR2_X2 \AES_ENC/u0/U425  ( .A(\AES_ENC/w2[3] ), .B(\AES_ENC/u0/N104 ), .Z(\AES_ENC/u0/N170 ) );
XOR2_X2 \AES_ENC/u0/U424  ( .A(\AES_ENC/w3[3] ), .B(\AES_ENC/u0/N170 ), .Z(\AES_ENC/u0/N236 ) );
XOR2_X2 \AES_ENC/u0/U423  ( .A(\AES_ENC/u0/subword[2] ), .B(\AES_ENC/u0/n311 ), .Z(\AES_ENC/u0/N105 ) );
XOR2_X2 \AES_ENC/u0/U422  ( .A(\AES_ENC/w1[2] ), .B(\AES_ENC/w0[2] ), .Z(\AES_ENC/u0/n311 ) );
XOR2_X2 \AES_ENC/u0/U421  ( .A(\AES_ENC/w2[2] ), .B(\AES_ENC/u0/N105 ), .Z(\AES_ENC/u0/N171 ) );
XOR2_X2 \AES_ENC/u0/U420  ( .A(\AES_ENC/w3[2] ), .B(\AES_ENC/u0/N171 ), .Z(\AES_ENC/u0/N237 ) );
XOR2_X2 \AES_ENC/u0/U419  ( .A(\AES_ENC/u0/subword[1] ), .B(\AES_ENC/u0/n312 ), .Z(\AES_ENC/u0/N106 ) );
XOR2_X2 \AES_ENC/u0/U418  ( .A(\AES_ENC/w1[1] ), .B(\AES_ENC/w0[1] ), .Z(\AES_ENC/u0/n312 ) );
XOR2_X2 \AES_ENC/u0/U417  ( .A(\AES_ENC/w2[1] ), .B(\AES_ENC/u0/N106 ), .Z(\AES_ENC/u0/N172 ) );
XOR2_X2 \AES_ENC/u0/U416  ( .A(\AES_ENC/w3[1] ), .B(\AES_ENC/u0/N172 ), .Z(\AES_ENC/u0/N238 ) );
XOR2_X2 \AES_ENC/u0/U415  ( .A(\AES_ENC/u0/subword[0] ), .B(\AES_ENC/u0/n313 ), .Z(\AES_ENC/u0/N107 ) );
XOR2_X2 \AES_ENC/u0/U414  ( .A(\AES_ENC/w1[0] ), .B(\AES_ENC/w0[0] ), .Z(\AES_ENC/u0/n313 ) );
XOR2_X2 \AES_ENC/u0/U413  ( .A(\AES_ENC/w2[0] ), .B(\AES_ENC/u0/N107 ), .Z(\AES_ENC/u0/N173 ) );
XOR2_X2 \AES_ENC/u0/U412  ( .A(\AES_ENC/w3[0] ), .B(\AES_ENC/u0/N173 ), .Z(\AES_ENC/u0/N239 ) );
INV_X4 \AES_ENC/u0/u0/U575  ( .A(\AES_ENC/w3[23] ), .ZN(\AES_ENC/u0/u0/n627 ) );
INV_X4 \AES_ENC/u0/u0/U574  ( .A(\AES_ENC/u0/u0/n1114 ), .ZN(\AES_ENC/u0/u0/n625 ) );
INV_X4 \AES_ENC/u0/u0/U573  ( .A(\AES_ENC/w3[20] ), .ZN(\AES_ENC/u0/u0/n624 ) );
INV_X4 \AES_ENC/u0/u0/U572  ( .A(\AES_ENC/u0/u0/n1025 ), .ZN(\AES_ENC/u0/u0/n622 ) );
INV_X4 \AES_ENC/u0/u0/U571  ( .A(\AES_ENC/u0/u0/n1120 ), .ZN(\AES_ENC/u0/u0/n620 ) );
INV_X4 \AES_ENC/u0/u0/U570  ( .A(\AES_ENC/u0/u0/n1121 ), .ZN(\AES_ENC/u0/u0/n619 ) );
INV_X4 \AES_ENC/u0/u0/U569  ( .A(\AES_ENC/u0/u0/n1048 ), .ZN(\AES_ENC/u0/u0/n618 ) );
INV_X4 \AES_ENC/u0/u0/U568  ( .A(\AES_ENC/u0/u0/n974 ), .ZN(\AES_ENC/u0/u0/n616 ) );
INV_X4 \AES_ENC/u0/u0/U567  ( .A(\AES_ENC/u0/u0/n794 ), .ZN(\AES_ENC/u0/u0/n614 ) );
INV_X4 \AES_ENC/u0/u0/U566  ( .A(\AES_ENC/w3[18] ), .ZN(\AES_ENC/u0/u0/n611 ) );
INV_X4 \AES_ENC/u0/u0/U565  ( .A(\AES_ENC/u0/u0/n800 ), .ZN(\AES_ENC/u0/u0/n610 ) );
INV_X4 \AES_ENC/u0/u0/U564  ( .A(\AES_ENC/u0/u0/n925 ), .ZN(\AES_ENC/u0/u0/n609 ) );
INV_X4 \AES_ENC/u0/u0/U563  ( .A(\AES_ENC/u0/u0/n779 ), .ZN(\AES_ENC/u0/u0/n607 ) );
INV_X4 \AES_ENC/u0/u0/U562  ( .A(\AES_ENC/u0/u0/n1022 ), .ZN(\AES_ENC/u0/u0/n603 ) );
INV_X4 \AES_ENC/u0/u0/U561  ( .A(\AES_ENC/u0/u0/n1102 ), .ZN(\AES_ENC/u0/u0/n602 ) );
INV_X4 \AES_ENC/u0/u0/U560  ( .A(\AES_ENC/u0/u0/n929 ), .ZN(\AES_ENC/u0/u0/n601 ) );
INV_X4 \AES_ENC/u0/u0/U559  ( .A(\AES_ENC/u0/u0/n1056 ), .ZN(\AES_ENC/u0/u0/n600 ) );
INV_X4 \AES_ENC/u0/u0/U558  ( .A(\AES_ENC/u0/u0/n1054 ), .ZN(\AES_ENC/u0/u0/n599 ) );
INV_X4 \AES_ENC/u0/u0/U557  ( .A(\AES_ENC/u0/u0/n881 ), .ZN(\AES_ENC/u0/u0/n598 ) );
INV_X4 \AES_ENC/u0/u0/U556  ( .A(\AES_ENC/u0/u0/n926 ), .ZN(\AES_ENC/u0/u0/n597 ) );
INV_X4 \AES_ENC/u0/u0/U555  ( .A(\AES_ENC/u0/u0/n977 ), .ZN(\AES_ENC/u0/u0/n595 ) );
INV_X4 \AES_ENC/u0/u0/U554  ( .A(\AES_ENC/u0/u0/n1031 ), .ZN(\AES_ENC/u0/u0/n594 ) );
INV_X4 \AES_ENC/u0/u0/U553  ( .A(\AES_ENC/u0/u0/n1103 ), .ZN(\AES_ENC/u0/u0/n593 ) );
INV_X4 \AES_ENC/u0/u0/U552  ( .A(\AES_ENC/u0/u0/n1009 ), .ZN(\AES_ENC/u0/u0/n592 ) );
INV_X4 \AES_ENC/u0/u0/U551  ( .A(\AES_ENC/u0/u0/n990 ), .ZN(\AES_ENC/u0/u0/n591 ) );
INV_X4 \AES_ENC/u0/u0/U550  ( .A(\AES_ENC/u0/u0/n1058 ), .ZN(\AES_ENC/u0/u0/n590 ) );
INV_X4 \AES_ENC/u0/u0/U549  ( .A(\AES_ENC/u0/u0/n1074 ), .ZN(\AES_ENC/u0/u0/n589 ) );
INV_X4 \AES_ENC/u0/u0/U548  ( .A(\AES_ENC/u0/u0/n1053 ), .ZN(\AES_ENC/u0/u0/n588 ) );
INV_X4 \AES_ENC/u0/u0/U547  ( .A(\AES_ENC/u0/u0/n826 ), .ZN(\AES_ENC/u0/u0/n587 ) );
INV_X4 \AES_ENC/u0/u0/U546  ( .A(\AES_ENC/u0/u0/n992 ), .ZN(\AES_ENC/u0/u0/n586 ) );
INV_X4 \AES_ENC/u0/u0/U545  ( .A(\AES_ENC/u0/u0/n821 ), .ZN(\AES_ENC/u0/u0/n585 ) );
INV_X4 \AES_ENC/u0/u0/U544  ( .A(\AES_ENC/u0/u0/n910 ), .ZN(\AES_ENC/u0/u0/n584 ) );
INV_X4 \AES_ENC/u0/u0/U543  ( .A(\AES_ENC/u0/u0/n906 ), .ZN(\AES_ENC/u0/u0/n583 ) );
INV_X4 \AES_ENC/u0/u0/U542  ( .A(\AES_ENC/u0/u0/n880 ), .ZN(\AES_ENC/u0/u0/n581 ) );
INV_X4 \AES_ENC/u0/u0/U541  ( .A(\AES_ENC/u0/u0/n1013 ), .ZN(\AES_ENC/u0/u0/n580 ) );
INV_X4 \AES_ENC/u0/u0/U540  ( .A(\AES_ENC/u0/u0/n1092 ), .ZN(\AES_ENC/u0/u0/n579 ) );
INV_X4 \AES_ENC/u0/u0/U539  ( .A(\AES_ENC/u0/u0/n824 ), .ZN(\AES_ENC/u0/u0/n578 ) );
INV_X4 \AES_ENC/u0/u0/U538  ( .A(\AES_ENC/u0/u0/n1091 ), .ZN(\AES_ENC/u0/u0/n577 ) );
INV_X4 \AES_ENC/u0/u0/U537  ( .A(\AES_ENC/u0/u0/n1080 ), .ZN(\AES_ENC/u0/u0/n576 ) );
INV_X4 \AES_ENC/u0/u0/U536  ( .A(\AES_ENC/u0/u0/n959 ), .ZN(\AES_ENC/u0/u0/n575 ) );
INV_X4 \AES_ENC/u0/u0/U535  ( .A(\AES_ENC/w3[16] ), .ZN(\AES_ENC/u0/u0/n574 ) );
NOR2_X2 \AES_ENC/u0/u0/U534  ( .A1(\AES_ENC/w3[20] ), .A2(\AES_ENC/w3[19] ),.ZN(\AES_ENC/u0/u0/n1025 ) );
INV_X4 \AES_ENC/u0/u0/U533  ( .A(\AES_ENC/u0/u0/n569 ), .ZN(\AES_ENC/u0/u0/n572 ) );
NOR2_X2 \AES_ENC/u0/u0/U532  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n765 ) );
NOR2_X2 \AES_ENC/u0/u0/U531  ( .A1(\AES_ENC/w3[20] ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n764 ) );
NOR2_X2 \AES_ENC/u0/u0/U530  ( .A1(\AES_ENC/u0/u0/n765 ), .A2(\AES_ENC/u0/u0/n764 ), .ZN(\AES_ENC/u0/u0/n766 ) );
NOR2_X2 \AES_ENC/u0/u0/U529  ( .A1(\AES_ENC/u0/u0/n766 ), .A2(\AES_ENC/u0/u0/n575 ), .ZN(\AES_ENC/u0/u0/n767 ) );
NOR2_X2 \AES_ENC/u0/u0/U528  ( .A1(\AES_ENC/u0/u0/n1117 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n707 ) );
NOR3_X2 \AES_ENC/u0/u0/U527  ( .A1(\AES_ENC/u0/u0/n627 ), .A2(\AES_ENC/w3[21] ), .A3(\AES_ENC/u0/u0/n704 ), .ZN(\AES_ENC/u0/u0/n706 ) );
NOR2_X2 \AES_ENC/u0/u0/U526  ( .A1(\AES_ENC/w3[20] ), .A2(\AES_ENC/u0/u0/n579 ), .ZN(\AES_ENC/u0/u0/n705 ) );
NOR3_X2 \AES_ENC/u0/u0/U525  ( .A1(\AES_ENC/u0/u0/n707 ), .A2(\AES_ENC/u0/u0/n706 ), .A3(\AES_ENC/u0/u0/n705 ), .ZN(\AES_ENC/u0/u0/n713 ) );
NOR4_X2 \AES_ENC/u0/u0/U524  ( .A1(\AES_ENC/u0/u0/n633 ), .A2(\AES_ENC/u0/u0/n632 ), .A3(\AES_ENC/u0/u0/n631 ), .A4(\AES_ENC/u0/u0/n630 ), .ZN(\AES_ENC/u0/u0/n634 ) );
NOR2_X2 \AES_ENC/u0/u0/U523  ( .A1(\AES_ENC/u0/u0/n629 ), .A2(\AES_ENC/u0/u0/n628 ), .ZN(\AES_ENC/u0/u0/n635 ) );
NAND3_X2 \AES_ENC/u0/u0/U522  ( .A1(\AES_ENC/w3[18] ), .A2(\AES_ENC/w3[23] ),.A3(\AES_ENC/u0/u0/n1059 ), .ZN(\AES_ENC/u0/u0/n636 ) );
INV_X4 \AES_ENC/u0/u0/U521  ( .A(\AES_ENC/w3[19] ), .ZN(\AES_ENC/u0/u0/n621 ) );
NOR2_X2 \AES_ENC/u0/u0/U520  ( .A1(\AES_ENC/w3[21] ), .A2(\AES_ENC/w3[18] ),.ZN(\AES_ENC/u0/u0/n974 ) );
NAND3_X2 \AES_ENC/u0/u0/U519  ( .A1(\AES_ENC/u0/u0/n652 ), .A2(\AES_ENC/u0/u0/n626 ), .A3(\AES_ENC/w3[23] ), .ZN(\AES_ENC/u0/u0/n653 ) );
NOR2_X2 \AES_ENC/u0/u0/U518  ( .A1(\AES_ENC/u0/u0/n611 ), .A2(\AES_ENC/w3[21] ), .ZN(\AES_ENC/u0/u0/n925 ) );
NOR2_X2 \AES_ENC/u0/u0/U517  ( .A1(\AES_ENC/u0/u0/n626 ), .A2(\AES_ENC/w3[18] ), .ZN(\AES_ENC/u0/u0/n1048 ) );
INV_X4 \AES_ENC/u0/u0/U516  ( .A(\AES_ENC/w3[21] ), .ZN(\AES_ENC/u0/u0/n626 ) );
NOR2_X2 \AES_ENC/u0/u0/U515  ( .A1(\AES_ENC/u0/u0/n611 ), .A2(\AES_ENC/w3[23] ), .ZN(\AES_ENC/u0/u0/n779 ) );
NOR2_X2 \AES_ENC/u0/u0/U512  ( .A1(\AES_ENC/w3[23] ), .A2(\AES_ENC/w3[18] ),.ZN(\AES_ENC/u0/u0/n794 ) );
NAND3_X2 \AES_ENC/u0/u0/U510  ( .A1(\AES_ENC/u0/u0/n679 ), .A2(\AES_ENC/u0/u0/n678 ), .A3(\AES_ENC/u0/u0/n677 ), .ZN(\AES_ENC/u0/subword[24] ) );
NOR2_X2 \AES_ENC/u0/u0/U509  ( .A1(\AES_ENC/u0/u0/n574 ), .A2(\AES_ENC/w3[22] ), .ZN(\AES_ENC/u0/u0/n1070 ) );
NOR2_X2 \AES_ENC/u0/u0/U508  ( .A1(\AES_ENC/w3[16] ), .A2(\AES_ENC/w3[22] ),.ZN(\AES_ENC/u0/u0/n1090 ) );
NOR2_X2 \AES_ENC/u0/u0/U507  ( .A1(\AES_ENC/w3[20] ), .A2(\AES_ENC/w3[17] ),.ZN(\AES_ENC/u0/u0/n1102 ) );
NOR2_X2 \AES_ENC/u0/u0/U506  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/w3[19] ), .ZN(\AES_ENC/u0/u0/n1053 ) );
NOR2_X2 \AES_ENC/u0/u0/U505  ( .A1(\AES_ENC/u0/u0/n607 ), .A2(\AES_ENC/w3[21] ), .ZN(\AES_ENC/u0/u0/n1024 ) );
NOR2_X2 \AES_ENC/u0/u0/U504  ( .A1(\AES_ENC/u0/u0/n625 ), .A2(\AES_ENC/w3[18] ), .ZN(\AES_ENC/u0/u0/n1093 ) );
NOR2_X2 \AES_ENC/u0/u0/U503  ( .A1(\AES_ENC/u0/u0/n614 ), .A2(\AES_ENC/w3[21] ), .ZN(\AES_ENC/u0/u0/n1094 ) );
NOR2_X2 \AES_ENC/u0/u0/U502  ( .A1(\AES_ENC/u0/u0/n624 ), .A2(\AES_ENC/w3[19] ), .ZN(\AES_ENC/u0/u0/n931 ) );
INV_X4 \AES_ENC/u0/u0/U501  ( .A(\AES_ENC/u0/u0/n570 ), .ZN(\AES_ENC/u0/u0/n573 ) );
NOR2_X2 \AES_ENC/u0/u0/U500  ( .A1(\AES_ENC/u0/u0/n622 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n1059 ) );
NOR4_X2 \AES_ENC/u0/u0/U499  ( .A1(\AES_ENC/u0/u0/n1125 ), .A2(\AES_ENC/u0/u0/n1124 ), .A3(\AES_ENC/u0/u0/n1123 ), .A4(\AES_ENC/u0/u0/n1122 ), .ZN(\AES_ENC/u0/u0/n1126 ) );
NOR2_X2 \AES_ENC/u0/u0/U498  ( .A1(\AES_ENC/u0/u0/n826 ), .A2(\AES_ENC/u0/u0/n572 ), .ZN(\AES_ENC/u0/u0/n827 ) );
NOR3_X2 \AES_ENC/u0/u0/U497  ( .A1(\AES_ENC/u0/u0/n769 ), .A2(\AES_ENC/u0/u0/n768 ), .A3(\AES_ENC/u0/u0/n767 ), .ZN(\AES_ENC/u0/u0/n775 ) );
NOR2_X2 \AES_ENC/u0/u0/U496  ( .A1(\AES_ENC/u0/u0/n946 ), .A2(\AES_ENC/u0/u0/n945 ), .ZN(\AES_ENC/u0/u0/n952 ) );
NOR2_X2 \AES_ENC/u0/u0/U495  ( .A1(\AES_ENC/w3[17] ), .A2(\AES_ENC/u0/u0/n623 ), .ZN(\AES_ENC/u0/u0/n913 ) );
NOR2_X2 \AES_ENC/u0/u0/U494  ( .A1(\AES_ENC/u0/u0/n913 ), .A2(\AES_ENC/u0/u0/n1091 ), .ZN(\AES_ENC/u0/u0/n914 ) );
NOR2_X2 \AES_ENC/u0/u0/U492  ( .A1(\AES_ENC/u0/u0/n1056 ), .A2(\AES_ENC/u0/u0/n1053 ), .ZN(\AES_ENC/u0/u0/n749 ) );
NOR2_X2 \AES_ENC/u0/u0/U491  ( .A1(\AES_ENC/u0/u0/n749 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n752 ) );
NOR4_X2 \AES_ENC/u0/u0/U490  ( .A1(\AES_ENC/u0/u0/n983 ), .A2(\AES_ENC/u0/u0/n698 ), .A3(\AES_ENC/u0/u0/n697 ), .A4(\AES_ENC/u0/u0/n696 ), .ZN(\AES_ENC/u0/u0/n699 ) );
NOR3_X2 \AES_ENC/u0/u0/U489  ( .A1(\AES_ENC/u0/u0/n695 ), .A2(\AES_ENC/u0/u0/n694 ), .A3(\AES_ENC/u0/u0/n693 ), .ZN(\AES_ENC/u0/u0/n700 ) );
NOR4_X2 \AES_ENC/u0/u0/U488  ( .A1(\AES_ENC/u0/u0/n757 ), .A2(\AES_ENC/u0/u0/n756 ), .A3(\AES_ENC/u0/u0/n755 ), .A4(\AES_ENC/u0/u0/n754 ), .ZN(\AES_ENC/u0/u0/n758 ) );
NOR2_X2 \AES_ENC/u0/u0/U487  ( .A1(\AES_ENC/u0/u0/n752 ), .A2(\AES_ENC/u0/u0/n751 ), .ZN(\AES_ENC/u0/u0/n759 ) );
NOR4_X2 \AES_ENC/u0/u0/U486  ( .A1(\AES_ENC/u0/u0/n870 ), .A2(\AES_ENC/u0/u0/n869 ), .A3(\AES_ENC/u0/u0/n868 ), .A4(\AES_ENC/u0/u0/n867 ), .ZN(\AES_ENC/u0/u0/n871 ) );
NOR3_X2 \AES_ENC/u0/u0/U483  ( .A1(\AES_ENC/u0/u0/n995 ), .A2(\AES_ENC/u0/u0/n586 ), .A3(\AES_ENC/u0/u0/n994 ), .ZN(\AES_ENC/u0/u0/n1002 ) );
NOR2_X2 \AES_ENC/u0/u0/U482  ( .A1(\AES_ENC/u0/u0/n1076 ), .A2(\AES_ENC/u0/u0/n1075 ), .ZN(\AES_ENC/u0/u0/n1086 ) );
NOR2_X2 \AES_ENC/u0/u0/U480  ( .A1(\AES_ENC/u0/u0/n1053 ), .A2(\AES_ENC/u0/u0/n1095 ), .ZN(\AES_ENC/u0/u0/n639 ) );
NOR2_X2 \AES_ENC/u0/u0/U479  ( .A1(\AES_ENC/u0/u0/n639 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n640 ) );
NOR2_X2 \AES_ENC/u0/u0/U478  ( .A1(\AES_ENC/u0/u0/n909 ), .A2(\AES_ENC/u0/u0/n908 ), .ZN(\AES_ENC/u0/u0/n920 ) );
INV_X4 \AES_ENC/u0/u0/U477  ( .A(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n596 ) );
NOR2_X2 \AES_ENC/u0/u0/U474  ( .A1(\AES_ENC/u0/u0/n932 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n933 ) );
NOR2_X2 \AES_ENC/u0/u0/U473  ( .A1(\AES_ENC/u0/u0/n929 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n935 ) );
NOR2_X2 \AES_ENC/u0/u0/U472  ( .A1(\AES_ENC/u0/u0/n931 ), .A2(\AES_ENC/u0/u0/n930 ), .ZN(\AES_ENC/u0/u0/n934 ) );
NOR3_X2 \AES_ENC/u0/u0/U471  ( .A1(\AES_ENC/u0/u0/n935 ), .A2(\AES_ENC/u0/u0/n934 ), .A3(\AES_ENC/u0/u0/n933 ), .ZN(\AES_ENC/u0/u0/n936 ) );
OR2_X4 \AES_ENC/u0/u0/U470  ( .A1(\AES_ENC/u0/u0/n1094 ), .A2(\AES_ENC/u0/u0/n1093 ), .ZN(\AES_ENC/u0/u0/n571 ) );
AND2_X2 \AES_ENC/u0/u0/U469  ( .A1(\AES_ENC/u0/u0/n571 ), .A2(\AES_ENC/u0/u0/n1095 ), .ZN(\AES_ENC/u0/u0/n1101 ) );
NOR2_X2 \AES_ENC/u0/u0/U468  ( .A1(\AES_ENC/u0/u0/n1074 ), .A2(\AES_ENC/u0/u0/n931 ), .ZN(\AES_ENC/u0/u0/n796 ) );
NOR2_X2 \AES_ENC/u0/u0/U467  ( .A1(\AES_ENC/u0/u0/n796 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n797 ) );
NOR2_X2 \AES_ENC/u0/u0/U466  ( .A1(\AES_ENC/u0/u0/n1054 ), .A2(\AES_ENC/u0/u0/n1053 ), .ZN(\AES_ENC/u0/u0/n1055 ) );
NOR2_X2 \AES_ENC/u0/u0/U465  ( .A1(\AES_ENC/u0/u0/n1049 ), .A2(\AES_ENC/u0/u0/n618 ), .ZN(\AES_ENC/u0/u0/n1051 ) );
NOR2_X2 \AES_ENC/u0/u0/U464  ( .A1(\AES_ENC/u0/u0/n1051 ), .A2(\AES_ENC/u0/u0/n1050 ), .ZN(\AES_ENC/u0/u0/n1052 ) );
NOR2_X2 \AES_ENC/u0/u0/U463  ( .A1(\AES_ENC/u0/u0/n1052 ), .A2(\AES_ENC/u0/u0/n592 ), .ZN(\AES_ENC/u0/u0/n1064 ) );
NOR2_X2 \AES_ENC/u0/u0/U462  ( .A1(\AES_ENC/w3[17] ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n631 ) );
NOR2_X2 \AES_ENC/u0/u0/U461  ( .A1(\AES_ENC/u0/u0/n1025 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n980 ) );
NOR2_X2 \AES_ENC/u0/u0/U460  ( .A1(\AES_ENC/u0/u0/n1073 ), .A2(\AES_ENC/u0/u0/n1094 ), .ZN(\AES_ENC/u0/u0/n795 ) );
NOR2_X2 \AES_ENC/u0/u0/U459  ( .A1(\AES_ENC/u0/u0/n795 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n799 ) );
NOR2_X2 \AES_ENC/u0/u0/U458  ( .A1(\AES_ENC/u0/u0/n624 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n1075 ) );
NOR2_X2 \AES_ENC/u0/u0/U455  ( .A1(\AES_ENC/u0/u0/n624 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n822 ) );
NOR2_X2 \AES_ENC/u0/u0/U448  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n823 ) );
NOR2_X2 \AES_ENC/u0/u0/U447  ( .A1(\AES_ENC/u0/u0/n823 ), .A2(\AES_ENC/u0/u0/n822 ), .ZN(\AES_ENC/u0/u0/n825 ) );
NOR2_X2 \AES_ENC/u0/u0/U442  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n981 ) );
NOR2_X2 \AES_ENC/u0/u0/U441  ( .A1(\AES_ENC/u0/u0/n1074 ), .A2(\AES_ENC/u0/u0/n1025 ), .ZN(\AES_ENC/u0/u0/n891 ) );
NOR2_X2 \AES_ENC/u0/u0/U438  ( .A1(\AES_ENC/u0/u0/n1102 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n643 ) );
NOR2_X2 \AES_ENC/u0/u0/U435  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n621 ), .ZN(\AES_ENC/u0/u0/n642 ) );
NOR2_X2 \AES_ENC/u0/u0/U434  ( .A1(\AES_ENC/u0/u0/n911 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n644 ) );
NOR4_X2 \AES_ENC/u0/u0/U433  ( .A1(\AES_ENC/u0/u0/n644 ), .A2(\AES_ENC/u0/u0/n643 ), .A3(\AES_ENC/u0/u0/n804 ), .A4(\AES_ENC/u0/u0/n642 ), .ZN(\AES_ENC/u0/u0/n645 ) );
NOR2_X2 \AES_ENC/u0/u0/U428  ( .A1(\AES_ENC/u0/u0/n1102 ), .A2(\AES_ENC/u0/u0/n910 ), .ZN(\AES_ENC/u0/u0/n932 ) );
NOR3_X2 \AES_ENC/u0/u0/U427  ( .A1(\AES_ENC/u0/u0/n623 ), .A2(\AES_ENC/w3[17] ), .A3(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n683 ) );
NOR2_X2 \AES_ENC/u0/u0/U421  ( .A1(\AES_ENC/u0/u0/n1102 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n755 ) );
INV_X4 \AES_ENC/u0/u0/U420  ( .A(\AES_ENC/u0/u0/n931 ), .ZN(\AES_ENC/u0/u0/n623 ) );
NOR2_X2 \AES_ENC/u0/u0/U419  ( .A1(\AES_ENC/u0/u0/n996 ), .A2(\AES_ENC/u0/u0/n931 ), .ZN(\AES_ENC/u0/u0/n704 ) );
NOR2_X2 \AES_ENC/u0/u0/U418  ( .A1(\AES_ENC/u0/u0/n1029 ), .A2(\AES_ENC/u0/u0/n1025 ), .ZN(\AES_ENC/u0/u0/n1079 ) );
NOR3_X2 \AES_ENC/u0/u0/U417  ( .A1(\AES_ENC/u0/u0/n589 ), .A2(\AES_ENC/u0/u0/n1025 ), .A3(\AES_ENC/u0/u0/n616 ), .ZN(\AES_ENC/u0/u0/n945 ) );
NOR2_X2 \AES_ENC/u0/u0/U416  ( .A1(\AES_ENC/u0/u0/n1072 ), .A2(\AES_ENC/u0/u0/n1094 ), .ZN(\AES_ENC/u0/u0/n930 ) );
NOR2_X2 \AES_ENC/u0/u0/U415  ( .A1(\AES_ENC/u0/u0/n931 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n743 ) );
NOR2_X2 \AES_ENC/u0/u0/U414  ( .A1(\AES_ENC/u0/u0/n931 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n685 ) );
NOR3_X2 \AES_ENC/u0/u0/U413  ( .A1(\AES_ENC/u0/u0/n610 ), .A2(\AES_ENC/u0/u0/n572 ), .A3(\AES_ENC/u0/u0/n575 ), .ZN(\AES_ENC/u0/u0/n962 ) );
NOR2_X2 \AES_ENC/u0/u0/U410  ( .A1(\AES_ENC/u0/u0/n626 ), .A2(\AES_ENC/u0/u0/n611 ), .ZN(\AES_ENC/u0/u0/n800 ) );
NOR3_X2 \AES_ENC/u0/u0/U409  ( .A1(\AES_ENC/u0/u0/n590 ), .A2(\AES_ENC/u0/u0/n627 ), .A3(\AES_ENC/u0/u0/n611 ), .ZN(\AES_ENC/u0/u0/n798 ) );
NOR3_X2 \AES_ENC/u0/u0/U406  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n572 ), .A3(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n694 ) );
NOR4_X2 \AES_ENC/u0/u0/U405  ( .A1(\AES_ENC/u0/u0/n946 ), .A2(\AES_ENC/u0/u0/n1046 ), .A3(\AES_ENC/u0/u0/n671 ), .A4(\AES_ENC/u0/u0/n670 ), .ZN(\AES_ENC/u0/u0/n672 ) );
NOR4_X2 \AES_ENC/u0/u0/U404  ( .A1(\AES_ENC/u0/u0/n806 ), .A2(\AES_ENC/u0/u0/n805 ), .A3(\AES_ENC/u0/u0/n804 ), .A4(\AES_ENC/u0/u0/n803 ), .ZN(\AES_ENC/u0/u0/n807 ) );
NOR3_X2 \AES_ENC/u0/u0/U403  ( .A1(\AES_ENC/u0/u0/n799 ), .A2(\AES_ENC/u0/u0/n798 ), .A3(\AES_ENC/u0/u0/n797 ), .ZN(\AES_ENC/u0/u0/n808 ) );
NOR3_X2 \AES_ENC/u0/u0/U401  ( .A1(\AES_ENC/u0/u0/n1101 ), .A2(\AES_ENC/u0/u0/n1100 ), .A3(\AES_ENC/u0/u0/n1099 ), .ZN(\AES_ENC/u0/u0/n1109 ) );
NOR2_X2 \AES_ENC/u0/u0/U400  ( .A1(\AES_ENC/u0/u0/n641 ), .A2(\AES_ENC/u0/u0/n640 ), .ZN(\AES_ENC/u0/u0/n646 ) );
NOR3_X2 \AES_ENC/u0/u0/U399  ( .A1(\AES_ENC/u0/u0/n743 ), .A2(\AES_ENC/u0/u0/n742 ), .A3(\AES_ENC/u0/u0/n741 ), .ZN(\AES_ENC/u0/u0/n744 ) );
NOR2_X2 \AES_ENC/u0/u0/U398  ( .A1(\AES_ENC/u0/u0/n697 ), .A2(\AES_ENC/u0/u0/n658 ), .ZN(\AES_ENC/u0/u0/n659 ) );
NOR3_X2 \AES_ENC/u0/u0/U397  ( .A1(\AES_ENC/u0/u0/n959 ), .A2(\AES_ENC/u0/u0/n572 ), .A3(\AES_ENC/u0/u0/n609 ), .ZN(\AES_ENC/u0/u0/n768 ) );
NOR2_X2 \AES_ENC/u0/u0/U396  ( .A1(\AES_ENC/u0/u0/n891 ), .A2(\AES_ENC/u0/u0/n609 ), .ZN(\AES_ENC/u0/u0/n894 ) );
NOR3_X2 \AES_ENC/u0/u0/U393  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n572 ), .A3(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n895 ) );
NOR3_X2 \AES_ENC/u0/u0/U390  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n1056 ), .A3(\AES_ENC/u0/u0/n990 ), .ZN(\AES_ENC/u0/u0/n896 ) );
NOR4_X2 \AES_ENC/u0/u0/U389  ( .A1(\AES_ENC/u0/u0/n896 ), .A2(\AES_ENC/u0/u0/n895 ), .A3(\AES_ENC/u0/u0/n894 ), .A4(\AES_ENC/u0/u0/n893 ), .ZN(\AES_ENC/u0/u0/n897 ) );
NOR2_X2 \AES_ENC/u0/u0/U388  ( .A1(\AES_ENC/u0/u0/n598 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n885 ) );
NOR2_X2 \AES_ENC/u0/u0/U387  ( .A1(\AES_ENC/u0/u0/n623 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n882 ) );
NOR2_X2 \AES_ENC/u0/u0/U386  ( .A1(\AES_ENC/u0/u0/n1053 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n884 ) );
NOR4_X2 \AES_ENC/u0/u0/U385  ( .A1(\AES_ENC/u0/u0/n885 ), .A2(\AES_ENC/u0/u0/n884 ), .A3(\AES_ENC/u0/u0/n883 ), .A4(\AES_ENC/u0/u0/n882 ), .ZN(\AES_ENC/u0/u0/n886 ) );
NOR2_X2 \AES_ENC/u0/u0/U384  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n569 ), .ZN(\AES_ENC/u0/u0/n947 ) );
NOR2_X2 \AES_ENC/u0/u0/U383  ( .A1(\AES_ENC/u0/u0/n572 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n949 ) );
NOR2_X2 \AES_ENC/u0/u0/U382  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n602 ), .ZN(\AES_ENC/u0/u0/n950 ) );
NOR4_X2 \AES_ENC/u0/u0/U374  ( .A1(\AES_ENC/u0/u0/n950 ), .A2(\AES_ENC/u0/u0/n949 ), .A3(\AES_ENC/u0/u0/n948 ), .A4(\AES_ENC/u0/u0/n947 ), .ZN(\AES_ENC/u0/u0/n951 ) );
NOR2_X2 \AES_ENC/u0/u0/U373  ( .A1(\AES_ENC/u0/u0/n1078 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n1033 ) );
NOR2_X2 \AES_ENC/u0/u0/U372  ( .A1(\AES_ENC/u0/u0/n1031 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n1032 ) );
NOR3_X2 \AES_ENC/u0/u0/U370  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n1025 ), .A3(\AES_ENC/u0/u0/n1074 ), .ZN(\AES_ENC/u0/u0/n1035 ) );
NOR4_X2 \AES_ENC/u0/u0/U369  ( .A1(\AES_ENC/u0/u0/n1035 ), .A2(\AES_ENC/u0/u0/n1034 ), .A3(\AES_ENC/u0/u0/n1033 ), .A4(\AES_ENC/u0/u0/n1032 ), .ZN(\AES_ENC/u0/u0/n1036 ) );
NOR2_X2 \AES_ENC/u0/u0/U368  ( .A1(\AES_ENC/u0/u0/n825 ), .A2(\AES_ENC/u0/u0/n578 ), .ZN(\AES_ENC/u0/u0/n830 ) );
NOR2_X2 \AES_ENC/u0/u0/U367  ( .A1(\AES_ENC/u0/u0/n827 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n829 ) );
NOR2_X2 \AES_ENC/u0/u0/U366  ( .A1(\AES_ENC/u0/u0/n572 ), .A2(\AES_ENC/u0/u0/n579 ), .ZN(\AES_ENC/u0/u0/n828 ) );
NOR4_X2 \AES_ENC/u0/u0/U365  ( .A1(\AES_ENC/u0/u0/n831 ), .A2(\AES_ENC/u0/u0/n830 ), .A3(\AES_ENC/u0/u0/n829 ), .A4(\AES_ENC/u0/u0/n828 ), .ZN(\AES_ENC/u0/u0/n832 ) );
NOR2_X2 \AES_ENC/u0/u0/U364  ( .A1(\AES_ENC/u0/u0/n598 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n1107 ) );
NOR2_X2 \AES_ENC/u0/u0/U363  ( .A1(\AES_ENC/u0/u0/n1102 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n1106 ) );
NOR2_X2 \AES_ENC/u0/u0/U354  ( .A1(\AES_ENC/u0/u0/n1103 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n1105 ) );
NOR4_X2 \AES_ENC/u0/u0/U353  ( .A1(\AES_ENC/u0/u0/n1107 ), .A2(\AES_ENC/u0/u0/n1106 ), .A3(\AES_ENC/u0/u0/n1105 ), .A4(\AES_ENC/u0/u0/n1104 ), .ZN(\AES_ENC/u0/u0/n1108 ) );
NOR3_X2 \AES_ENC/u0/u0/U352  ( .A1(\AES_ENC/u0/u0/n959 ), .A2(\AES_ENC/u0/u0/n621 ), .A3(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n963 ) );
NOR2_X2 \AES_ENC/u0/u0/U351  ( .A1(\AES_ENC/u0/u0/n626 ), .A2(\AES_ENC/u0/u0/n627 ), .ZN(\AES_ENC/u0/u0/n1114 ) );
NOR3_X2 \AES_ENC/u0/u0/U350  ( .A1(\AES_ENC/u0/u0/n910 ), .A2(\AES_ENC/u0/u0/n1059 ), .A3(\AES_ENC/u0/u0/n611 ), .ZN(\AES_ENC/u0/u0/n1115 ) );
INV_X4 \AES_ENC/u0/u0/U349  ( .A(\AES_ENC/u0/u0/n1024 ), .ZN(\AES_ENC/u0/u0/n606 ) );
INV_X4 \AES_ENC/u0/u0/U348  ( .A(\AES_ENC/u0/u0/n1094 ), .ZN(\AES_ENC/u0/u0/n613 ) );
NOR2_X2 \AES_ENC/u0/u0/U347  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n931 ), .ZN(\AES_ENC/u0/u0/n1100 ) );
NOR2_X2 \AES_ENC/u0/u0/U346  ( .A1(\AES_ENC/u0/u0/n569 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n929 ) );
NOR2_X2 \AES_ENC/u0/u0/U345  ( .A1(\AES_ENC/u0/u0/n620 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n926 ) );
INV_X4 \AES_ENC/u0/u0/U338  ( .A(\AES_ENC/u0/u0/n1093 ), .ZN(\AES_ENC/u0/u0/n617 ) );
NOR2_X2 \AES_ENC/u0/u0/U335  ( .A1(\AES_ENC/u0/u0/n572 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n1095 ) );
NOR2_X2 \AES_ENC/u0/u0/U329  ( .A1(\AES_ENC/u0/u0/n609 ), .A2(\AES_ENC/u0/u0/n627 ), .ZN(\AES_ENC/u0/u0/n1010 ) );
NOR2_X2 \AES_ENC/u0/u0/U328  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n1103 ) );
NOR2_X2 \AES_ENC/u0/u0/U327  ( .A1(\AES_ENC/w3[17] ), .A2(\AES_ENC/u0/u0/n1120 ), .ZN(\AES_ENC/u0/u0/n1022 ) );
NOR2_X2 \AES_ENC/u0/u0/U325  ( .A1(\AES_ENC/u0/u0/n619 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n911 ) );
NOR2_X2 \AES_ENC/u0/u0/U324  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/u0/u0/n1025 ), .ZN(\AES_ENC/u0/u0/n826 ) );
NOR2_X2 \AES_ENC/u0/u0/U319  ( .A1(\AES_ENC/u0/u0/n626 ), .A2(\AES_ENC/u0/u0/n607 ), .ZN(\AES_ENC/u0/u0/n1072 ) );
NOR2_X2 \AES_ENC/u0/u0/U318  ( .A1(\AES_ENC/u0/u0/n627 ), .A2(\AES_ENC/u0/u0/n616 ), .ZN(\AES_ENC/u0/u0/n956 ) );
NOR2_X2 \AES_ENC/u0/u0/U317  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/u0/u0/n624 ), .ZN(\AES_ENC/u0/u0/n1121 ) );
NOR2_X2 \AES_ENC/u0/u0/U316  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/u0/u0/n624 ), .ZN(\AES_ENC/u0/u0/n1058 ) );
NOR2_X2 \AES_ENC/u0/u0/U315  ( .A1(\AES_ENC/u0/u0/n625 ), .A2(\AES_ENC/u0/u0/n611 ), .ZN(\AES_ENC/u0/u0/n1073 ) );
NOR2_X2 \AES_ENC/u0/u0/U314  ( .A1(\AES_ENC/w3[17] ), .A2(\AES_ENC/u0/u0/n1025 ), .ZN(\AES_ENC/u0/u0/n1054 ) );
NOR2_X2 \AES_ENC/u0/u0/U312  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/u0/u0/n931 ), .ZN(\AES_ENC/u0/u0/n1029 ) );
NOR2_X2 \AES_ENC/u0/u0/U311  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n1056 ) );
NOR2_X2 \AES_ENC/u0/u0/U310  ( .A1(\AES_ENC/u0/u0/n614 ), .A2(\AES_ENC/u0/u0/n626 ), .ZN(\AES_ENC/u0/u0/n1050 ) );
NOR2_X2 \AES_ENC/u0/u0/U309  ( .A1(\AES_ENC/u0/u0/n1121 ), .A2(\AES_ENC/u0/u0/n1025 ), .ZN(\AES_ENC/u0/u0/n1120 ) );
NOR2_X2 \AES_ENC/u0/u0/U303  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/u0/u0/n572 ), .ZN(\AES_ENC/u0/u0/n1074 ) );
NOR2_X2 \AES_ENC/u0/u0/U302  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n584 ), .ZN(\AES_ENC/u0/u0/n838 ) );
NOR2_X2 \AES_ENC/u0/u0/U300  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n602 ), .ZN(\AES_ENC/u0/u0/n837 ) );
NOR2_X2 \AES_ENC/u0/u0/U299  ( .A1(\AES_ENC/u0/u0/n838 ), .A2(\AES_ENC/u0/u0/n837 ), .ZN(\AES_ENC/u0/u0/n845 ) );
NOR2_X2 \AES_ENC/u0/u0/U298  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n1071 ), .ZN(\AES_ENC/u0/u0/n669 ) );
NOR2_X2 \AES_ENC/u0/u0/U297  ( .A1(\AES_ENC/u0/u0/n1095 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n668 ) );
NOR2_X2 \AES_ENC/u0/u0/U296  ( .A1(\AES_ENC/u0/u0/n669 ), .A2(\AES_ENC/u0/u0/n668 ), .ZN(\AES_ENC/u0/u0/n673 ) );
NOR2_X2 \AES_ENC/u0/u0/U295  ( .A1(\AES_ENC/u0/u0/n1058 ), .A2(\AES_ENC/u0/u0/n1054 ), .ZN(\AES_ENC/u0/u0/n878 ) );
NOR2_X2 \AES_ENC/u0/u0/U294  ( .A1(\AES_ENC/u0/u0/n878 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n879 ) );
NOR2_X2 \AES_ENC/u0/u0/U293  ( .A1(\AES_ENC/u0/u0/n880 ), .A2(\AES_ENC/u0/u0/n879 ), .ZN(\AES_ENC/u0/u0/n887 ) );
NOR3_X2 \AES_ENC/u0/u0/U292  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n1091 ), .A3(\AES_ENC/u0/u0/n1022 ), .ZN(\AES_ENC/u0/u0/n720 ) );
NOR3_X2 \AES_ENC/u0/u0/U291  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n1054 ), .A3(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n719 ) );
NOR2_X2 \AES_ENC/u0/u0/U290  ( .A1(\AES_ENC/u0/u0/n720 ), .A2(\AES_ENC/u0/u0/n719 ), .ZN(\AES_ENC/u0/u0/n726 ) );
NOR2_X2 \AES_ENC/u0/u0/U284  ( .A1(\AES_ENC/u0/u0/n576 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n866 ) );
NOR2_X2 \AES_ENC/u0/u0/U283  ( .A1(\AES_ENC/u0/u0/n614 ), .A2(\AES_ENC/u0/u0/n591 ), .ZN(\AES_ENC/u0/u0/n865 ) );
NOR2_X2 \AES_ENC/u0/u0/U282  ( .A1(\AES_ENC/u0/u0/n866 ), .A2(\AES_ENC/u0/u0/n865 ), .ZN(\AES_ENC/u0/u0/n872 ) );
NOR2_X2 \AES_ENC/u0/u0/U281  ( .A1(\AES_ENC/u0/u0/n1059 ), .A2(\AES_ENC/u0/u0/n1058 ), .ZN(\AES_ENC/u0/u0/n1060 ) );
NOR2_X2 \AES_ENC/u0/u0/U280  ( .A1(\AES_ENC/u0/u0/n911 ), .A2(\AES_ENC/u0/u0/n910 ), .ZN(\AES_ENC/u0/u0/n912 ) );
NOR2_X2 \AES_ENC/u0/u0/U279  ( .A1(\AES_ENC/u0/u0/n912 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n916 ) );
NOR2_X2 \AES_ENC/u0/u0/U273  ( .A1(\AES_ENC/u0/u0/n826 ), .A2(\AES_ENC/u0/u0/n573 ), .ZN(\AES_ENC/u0/u0/n750 ) );
NOR2_X2 \AES_ENC/u0/u0/U272  ( .A1(\AES_ENC/u0/u0/n750 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n751 ) );
NOR2_X2 \AES_ENC/u0/u0/U271  ( .A1(\AES_ENC/u0/u0/n907 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n908 ) );
NOR2_X2 \AES_ENC/u0/u0/U270  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n588 ), .ZN(\AES_ENC/u0/u0/n957 ) );
NOR2_X2 \AES_ENC/u0/u0/U269  ( .A1(\AES_ENC/u0/u0/n990 ), .A2(\AES_ENC/u0/u0/n926 ), .ZN(\AES_ENC/u0/u0/n780 ) );
NOR2_X2 \AES_ENC/u0/u0/U268  ( .A1(\AES_ENC/u0/u0/n1022 ), .A2(\AES_ENC/u0/u0/n1058 ), .ZN(\AES_ENC/u0/u0/n740 ) );
NOR2_X2 \AES_ENC/u0/u0/U267  ( .A1(\AES_ENC/u0/u0/n740 ), .A2(\AES_ENC/u0/u0/n616 ), .ZN(\AES_ENC/u0/u0/n742 ) );
NOR2_X2 \AES_ENC/u0/u0/U263  ( .A1(\AES_ENC/u0/u0/n1098 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n1099 ) );
NOR2_X2 \AES_ENC/u0/u0/U262  ( .A1(\AES_ENC/u0/u0/n1120 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n993 ) );
NOR2_X2 \AES_ENC/u0/u0/U258  ( .A1(\AES_ENC/u0/u0/n993 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n994 ) );
NOR2_X2 \AES_ENC/u0/u0/U255  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n620 ), .ZN(\AES_ENC/u0/u0/n1026 ) );
NOR2_X2 \AES_ENC/u0/u0/U254  ( .A1(\AES_ENC/u0/u0/n573 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n1027 ) );
NOR2_X2 \AES_ENC/u0/u0/U253  ( .A1(\AES_ENC/u0/u0/n1027 ), .A2(\AES_ENC/u0/u0/n1026 ), .ZN(\AES_ENC/u0/u0/n1028 ) );
NOR2_X2 \AES_ENC/u0/u0/U252  ( .A1(\AES_ENC/u0/u0/n1029 ), .A2(\AES_ENC/u0/u0/n1028 ), .ZN(\AES_ENC/u0/u0/n1034 ) );
NOR2_X2 \AES_ENC/u0/u0/U251  ( .A1(\AES_ENC/u0/u0/n1056 ), .A2(\AES_ENC/u0/u0/n990 ), .ZN(\AES_ENC/u0/u0/n991 ) );
NOR2_X2 \AES_ENC/u0/u0/U250  ( .A1(\AES_ENC/u0/u0/n991 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n995 ) );
NOR2_X2 \AES_ENC/u0/u0/U243  ( .A1(\AES_ENC/u0/u0/n603 ), .A2(\AES_ENC/u0/u0/n610 ), .ZN(\AES_ENC/u0/u0/n1006 ) );
NOR2_X2 \AES_ENC/u0/u0/U242  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n577 ), .ZN(\AES_ENC/u0/u0/n1007 ) );
NOR2_X2 \AES_ENC/u0/u0/U241  ( .A1(\AES_ENC/u0/u0/n607 ), .A2(\AES_ENC/u0/u0/n590 ), .ZN(\AES_ENC/u0/u0/n1008 ) );
NOR3_X2 \AES_ENC/u0/u0/U240  ( .A1(\AES_ENC/u0/u0/n1008 ), .A2(\AES_ENC/u0/u0/n1007 ), .A3(\AES_ENC/u0/u0/n1006 ), .ZN(\AES_ENC/u0/u0/n1018 ) );
NOR2_X2 \AES_ENC/u0/u0/U239  ( .A1(\AES_ENC/u0/u0/n606 ), .A2(\AES_ENC/u0/u0/n906 ), .ZN(\AES_ENC/u0/u0/n741 ) );
NOR2_X2 \AES_ENC/u0/u0/U238  ( .A1(\AES_ENC/u0/u0/n1054 ), .A2(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n763 ) );
NOR2_X2 \AES_ENC/u0/u0/U237  ( .A1(\AES_ENC/u0/u0/n763 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n769 ) );
NOR2_X2 \AES_ENC/u0/u0/U236  ( .A1(\AES_ENC/u0/u0/n839 ), .A2(\AES_ENC/u0/u0/n582 ), .ZN(\AES_ENC/u0/u0/n693 ) );
NOR2_X2 \AES_ENC/u0/u0/U235  ( .A1(\AES_ENC/u0/u0/n609 ), .A2(\AES_ENC/u0/u0/n580 ), .ZN(\AES_ENC/u0/u0/n1123 ) );
NOR2_X2 \AES_ENC/u0/u0/U234  ( .A1(\AES_ENC/u0/u0/n780 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n784 ) );
NOR2_X2 \AES_ENC/u0/u0/U229  ( .A1(\AES_ENC/u0/u0/n1117 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n782 ) );
NOR2_X2 \AES_ENC/u0/u0/U228  ( .A1(\AES_ENC/u0/u0/n781 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n783 ) );
NOR4_X2 \AES_ENC/u0/u0/U227  ( .A1(\AES_ENC/u0/u0/n880 ), .A2(\AES_ENC/u0/u0/n784 ), .A3(\AES_ENC/u0/u0/n783 ), .A4(\AES_ENC/u0/u0/n782 ), .ZN(\AES_ENC/u0/u0/n785 ) );
INV_X4 \AES_ENC/u0/u0/U226  ( .A(\AES_ENC/u0/u0/n1029 ), .ZN(\AES_ENC/u0/u0/n582 ) );
NOR2_X2 \AES_ENC/u0/u0/U225  ( .A1(\AES_ENC/u0/u0/n593 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n1125 ) );
NOR2_X2 \AES_ENC/u0/u0/U223  ( .A1(\AES_ENC/u0/u0/n616 ), .A2(\AES_ENC/u0/u0/n580 ), .ZN(\AES_ENC/u0/u0/n771 ) );
NOR2_X2 \AES_ENC/u0/u0/U222  ( .A1(\AES_ENC/u0/u0/n616 ), .A2(\AES_ENC/u0/u0/n597 ), .ZN(\AES_ENC/u0/u0/n883 ) );
NOR2_X2 \AES_ENC/u0/u0/U221  ( .A1(\AES_ENC/u0/u0/n990 ), .A2(\AES_ENC/u0/u0/n929 ), .ZN(\AES_ENC/u0/u0/n892 ) );
NOR2_X2 \AES_ENC/u0/u0/U217  ( .A1(\AES_ENC/u0/u0/n892 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n893 ) );
NOR2_X2 \AES_ENC/u0/u0/U213  ( .A1(\AES_ENC/u0/u0/n910 ), .A2(\AES_ENC/u0/u0/n1056 ), .ZN(\AES_ENC/u0/u0/n941 ) );
NOR2_X2 \AES_ENC/u0/u0/U212  ( .A1(\AES_ENC/u0/u0/n623 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n630 ) );
NOR2_X2 \AES_ENC/u0/u0/U211  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n602 ), .ZN(\AES_ENC/u0/u0/n806 ) );
NOR2_X2 \AES_ENC/u0/u0/U210  ( .A1(\AES_ENC/u0/u0/n623 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n948 ) );
NOR2_X2 \AES_ENC/u0/u0/U209  ( .A1(\AES_ENC/u0/u0/n606 ), .A2(\AES_ENC/u0/u0/n582 ), .ZN(\AES_ENC/u0/u0/n1104 ) );
NOR2_X2 \AES_ENC/u0/u0/U208  ( .A1(\AES_ENC/u0/u0/n1121 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n1122 ) );
NOR2_X2 \AES_ENC/u0/u0/U207  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n1023 ), .ZN(\AES_ENC/u0/u0/n756 ) );
NOR2_X2 \AES_ENC/u0/u0/U201  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n602 ), .ZN(\AES_ENC/u0/u0/n870 ) );
NOR2_X2 \AES_ENC/u0/u0/U200  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n589 ), .ZN(\AES_ENC/u0/u0/n868 ) );
NOR2_X2 \AES_ENC/u0/u0/U199  ( .A1(\AES_ENC/u0/u0/n1120 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n1124 ) );
NOR2_X2 \AES_ENC/u0/u0/U198  ( .A1(\AES_ENC/u0/u0/n1120 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n696 ) );
NOR2_X2 \AES_ENC/u0/u0/U197  ( .A1(\AES_ENC/u0/u0/n1074 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n1076 ) );
NOR2_X2 \AES_ENC/u0/u0/U196  ( .A1(\AES_ENC/u0/u0/n1074 ), .A2(\AES_ENC/u0/u0/n620 ), .ZN(\AES_ENC/u0/u0/n781 ) );
NOR3_X2 \AES_ENC/u0/u0/U195  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n1056 ), .A3(\AES_ENC/u0/u0/n990 ), .ZN(\AES_ENC/u0/u0/n979 ) );
NOR3_X2 \AES_ENC/u0/u0/U194  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n1058 ), .A3(\AES_ENC/u0/u0/n1059 ), .ZN(\AES_ENC/u0/u0/n854 ) );
NOR2_X2 \AES_ENC/u0/u0/U187  ( .A1(\AES_ENC/u0/u0/n996 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n869 ) );
NOR2_X2 \AES_ENC/u0/u0/U186  ( .A1(\AES_ENC/u0/u0/n1056 ), .A2(\AES_ENC/u0/u0/n1074 ), .ZN(\AES_ENC/u0/u0/n1057 ) );
NOR3_X2 \AES_ENC/u0/u0/U185  ( .A1(\AES_ENC/u0/u0/n607 ), .A2(\AES_ENC/u0/u0/n1120 ), .A3(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n978 ) );
NOR2_X2 \AES_ENC/u0/u0/U184  ( .A1(\AES_ENC/u0/u0/n996 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n998 ) );
NOR2_X2 \AES_ENC/u0/u0/U183  ( .A1(\AES_ENC/u0/u0/n996 ), .A2(\AES_ENC/u0/u0/n911 ), .ZN(\AES_ENC/u0/u0/n1116 ) );
NOR2_X2 \AES_ENC/u0/u0/U182  ( .A1(\AES_ENC/u0/u0/n1074 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n754 ) );
NOR2_X2 \AES_ENC/u0/u0/U181  ( .A1(\AES_ENC/u0/u0/n926 ), .A2(\AES_ENC/u0/u0/n1103 ), .ZN(\AES_ENC/u0/u0/n977 ) );
NOR2_X2 \AES_ENC/u0/u0/U180  ( .A1(\AES_ENC/u0/u0/n839 ), .A2(\AES_ENC/u0/u0/n824 ), .ZN(\AES_ENC/u0/u0/n1092 ) );
NOR2_X2 \AES_ENC/u0/u0/U174  ( .A1(\AES_ENC/u0/u0/n573 ), .A2(\AES_ENC/u0/u0/n1074 ), .ZN(\AES_ENC/u0/u0/n684 ) );
NOR2_X2 \AES_ENC/u0/u0/U173  ( .A1(\AES_ENC/u0/u0/n826 ), .A2(\AES_ENC/u0/u0/n1059 ), .ZN(\AES_ENC/u0/u0/n907 ) );
NOR3_X2 \AES_ENC/u0/u0/U172  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n573 ), .A3(\AES_ENC/u0/u0/n1074 ), .ZN(\AES_ENC/u0/u0/n641 ) );
NOR3_X2 \AES_ENC/u0/u0/U171  ( .A1(\AES_ENC/u0/u0/n625 ), .A2(\AES_ENC/u0/u0/n1115 ), .A3(\AES_ENC/u0/u0/n585 ), .ZN(\AES_ENC/u0/u0/n831 ) );
NOR3_X2 \AES_ENC/u0/u0/U170  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n573 ), .A3(\AES_ENC/u0/u0/n1013 ), .ZN(\AES_ENC/u0/u0/n670 ) );
NOR2_X2 \AES_ENC/u0/u0/U169  ( .A1(\AES_ENC/u0/u0/n1029 ), .A2(\AES_ENC/u0/u0/n1095 ), .ZN(\AES_ENC/u0/u0/n735 ) );
NOR2_X2 \AES_ENC/u0/u0/U168  ( .A1(\AES_ENC/u0/u0/n1100 ), .A2(\AES_ENC/u0/u0/n854 ), .ZN(\AES_ENC/u0/u0/n860 ) );
NAND3_X2 \AES_ENC/u0/u0/U162  ( .A1(\AES_ENC/u0/u0/n569 ), .A2(\AES_ENC/u0/u0/n582 ), .A3(\AES_ENC/u0/u0/n681 ), .ZN(\AES_ENC/u0/u0/n691 ) );
NOR2_X2 \AES_ENC/u0/u0/U161  ( .A1(\AES_ENC/u0/u0/n683 ), .A2(\AES_ENC/u0/u0/n682 ), .ZN(\AES_ENC/u0/u0/n690 ) );
NOR4_X2 \AES_ENC/u0/u0/U160  ( .A1(\AES_ENC/u0/u0/n963 ), .A2(\AES_ENC/u0/u0/n962 ), .A3(\AES_ENC/u0/u0/n961 ), .A4(\AES_ENC/u0/u0/n960 ), .ZN(\AES_ENC/u0/u0/n964 ) );
NOR2_X2 \AES_ENC/u0/u0/U159  ( .A1(\AES_ENC/u0/u0/n958 ), .A2(\AES_ENC/u0/u0/n957 ), .ZN(\AES_ENC/u0/u0/n965 ) );
NOR4_X2 \AES_ENC/u0/u0/U158  ( .A1(\AES_ENC/u0/u0/n983 ), .A2(\AES_ENC/u0/u0/n982 ), .A3(\AES_ENC/u0/u0/n981 ), .A4(\AES_ENC/u0/u0/n980 ), .ZN(\AES_ENC/u0/u0/n984 ) );
NOR2_X2 \AES_ENC/u0/u0/U157  ( .A1(\AES_ENC/u0/u0/n979 ), .A2(\AES_ENC/u0/u0/n978 ), .ZN(\AES_ENC/u0/u0/n985 ) );
NOR3_X2 \AES_ENC/u0/u0/U156  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n1054 ), .A3(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n961 ) );
NOR3_X2 \AES_ENC/u0/u0/U155  ( .A1(\AES_ENC/u0/u0/n620 ), .A2(\AES_ENC/u0/u0/n1074 ), .A3(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n671 ) );
NOR2_X2 \AES_ENC/u0/u0/U154  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n1077 ), .ZN(\AES_ENC/u0/u0/n1084 ) );
NOR2_X2 \AES_ENC/u0/u0/U153  ( .A1(\AES_ENC/u0/u0/n1079 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n1082 ) );
NOR2_X2 \AES_ENC/u0/u0/U152  ( .A1(\AES_ENC/u0/u0/n1078 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n1083 ) );
NOR4_X2 \AES_ENC/u0/u0/U143  ( .A1(\AES_ENC/u0/u0/n1084 ), .A2(\AES_ENC/u0/u0/n1083 ), .A3(\AES_ENC/u0/u0/n1082 ), .A4(\AES_ENC/u0/u0/n1081 ), .ZN(\AES_ENC/u0/u0/n1085 ) );
NOR2_X2 \AES_ENC/u0/u0/U142  ( .A1(\AES_ENC/u0/u0/n1057 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n1062 ) );
NOR2_X2 \AES_ENC/u0/u0/U141  ( .A1(\AES_ENC/u0/u0/n1060 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n1061 ) );
NOR2_X2 \AES_ENC/u0/u0/U140  ( .A1(\AES_ENC/u0/u0/n1055 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n1063 ) );
NOR4_X2 \AES_ENC/u0/u0/U132  ( .A1(\AES_ENC/u0/u0/n1064 ), .A2(\AES_ENC/u0/u0/n1063 ), .A3(\AES_ENC/u0/u0/n1062 ), .A4(\AES_ENC/u0/u0/n1061 ), .ZN(\AES_ENC/u0/u0/n1065 ) );
NOR2_X2 \AES_ENC/u0/u0/U131  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n582 ), .ZN(\AES_ENC/u0/u0/n770 ) );
NOR2_X2 \AES_ENC/u0/u0/U130  ( .A1(\AES_ENC/u0/u0/n1103 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n772 ) );
NOR2_X2 \AES_ENC/u0/u0/U129  ( .A1(\AES_ENC/u0/u0/n610 ), .A2(\AES_ENC/u0/u0/n599 ), .ZN(\AES_ENC/u0/u0/n773 ) );
NOR4_X2 \AES_ENC/u0/u0/U128  ( .A1(\AES_ENC/u0/u0/n773 ), .A2(\AES_ENC/u0/u0/n772 ), .A3(\AES_ENC/u0/u0/n771 ), .A4(\AES_ENC/u0/u0/n770 ), .ZN(\AES_ENC/u0/u0/n774 ) );
NOR3_X2 \AES_ENC/u0/u0/U127  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n1091 ), .A3(\AES_ENC/u0/u0/n1022 ), .ZN(\AES_ENC/u0/u0/n843 ) );
NOR2_X2 \AES_ENC/u0/u0/U126  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n1077 ), .ZN(\AES_ENC/u0/u0/n841 ) );
NOR2_X2 \AES_ENC/u0/u0/U121  ( .A1(\AES_ENC/u0/u0/n1120 ), .A2(\AES_ENC/u0/u0/n839 ), .ZN(\AES_ENC/u0/u0/n842 ) );
NOR4_X2 \AES_ENC/u0/u0/U120  ( .A1(\AES_ENC/u0/u0/n843 ), .A2(\AES_ENC/u0/u0/n842 ), .A3(\AES_ENC/u0/u0/n841 ), .A4(\AES_ENC/u0/u0/n840 ), .ZN(\AES_ENC/u0/u0/n844 ) );
NOR2_X2 \AES_ENC/u0/u0/U119  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n595 ), .ZN(\AES_ENC/u0/u0/n858 ) );
NOR2_X2 \AES_ENC/u0/u0/U118  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n855 ), .ZN(\AES_ENC/u0/u0/n857 ) );
NOR2_X2 \AES_ENC/u0/u0/U117  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n587 ), .ZN(\AES_ENC/u0/u0/n856 ) );
NOR4_X2 \AES_ENC/u0/u0/U116  ( .A1(\AES_ENC/u0/u0/n858 ), .A2(\AES_ENC/u0/u0/n857 ), .A3(\AES_ENC/u0/u0/n856 ), .A4(\AES_ENC/u0/u0/n958 ), .ZN(\AES_ENC/u0/u0/n859 ) );
NOR3_X2 \AES_ENC/u0/u0/U115  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n1120 ), .A3(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n918 ) );
NOR2_X2 \AES_ENC/u0/u0/U106  ( .A1(\AES_ENC/u0/u0/n914 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n915 ) );
NOR3_X2 \AES_ENC/u0/u0/U105  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n573 ), .A3(\AES_ENC/u0/u0/n1013 ), .ZN(\AES_ENC/u0/u0/n917 ) );
NOR4_X2 \AES_ENC/u0/u0/U104  ( .A1(\AES_ENC/u0/u0/n918 ), .A2(\AES_ENC/u0/u0/n917 ), .A3(\AES_ENC/u0/u0/n916 ), .A4(\AES_ENC/u0/u0/n915 ), .ZN(\AES_ENC/u0/u0/n919 ) );
NOR2_X2 \AES_ENC/u0/u0/U103  ( .A1(\AES_ENC/u0/u0/n735 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n687 ) );
NOR2_X2 \AES_ENC/u0/u0/U102  ( .A1(\AES_ENC/u0/u0/n684 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n688 ) );
NOR2_X2 \AES_ENC/u0/u0/U101  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n600 ), .ZN(\AES_ENC/u0/u0/n686 ) );
NOR4_X2 \AES_ENC/u0/u0/U100  ( .A1(\AES_ENC/u0/u0/n688 ), .A2(\AES_ENC/u0/u0/n687 ), .A3(\AES_ENC/u0/u0/n686 ), .A4(\AES_ENC/u0/u0/n685 ), .ZN(\AES_ENC/u0/u0/n689 ) );
NOR2_X2 \AES_ENC/u0/u0/U95  ( .A1(\AES_ENC/u0/u0/n583 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n814 ) );
NOR3_X2 \AES_ENC/u0/u0/U94  ( .A1(\AES_ENC/u0/u0/n606 ), .A2(\AES_ENC/u0/u0/n1058 ), .A3(\AES_ENC/u0/u0/n1059 ), .ZN(\AES_ENC/u0/u0/n815 ) );
NOR2_X2 \AES_ENC/u0/u0/U93  ( .A1(\AES_ENC/u0/u0/n907 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n813 ) );
NOR4_X2 \AES_ENC/u0/u0/U92  ( .A1(\AES_ENC/u0/u0/n815 ), .A2(\AES_ENC/u0/u0/n814 ), .A3(\AES_ENC/u0/u0/n813 ), .A4(\AES_ENC/u0/u0/n812 ), .ZN(\AES_ENC/u0/u0/n816 ) );
NOR2_X2 \AES_ENC/u0/u0/U91  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n881 ), .ZN(\AES_ENC/u0/u0/n711 ) );
NOR2_X2 \AES_ENC/u0/u0/U90  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n855 ), .ZN(\AES_ENC/u0/u0/n709 ) );
NOR2_X2 \AES_ENC/u0/u0/U89  ( .A1(\AES_ENC/u0/u0/n609 ), .A2(\AES_ENC/u0/u0/n590 ), .ZN(\AES_ENC/u0/u0/n710 ) );
NOR4_X2 \AES_ENC/u0/u0/U88  ( .A1(\AES_ENC/u0/u0/n711 ), .A2(\AES_ENC/u0/u0/n710 ), .A3(\AES_ENC/u0/u0/n709 ), .A4(\AES_ENC/u0/u0/n708 ), .ZN(\AES_ENC/u0/u0/n712 ) );
NOR2_X2 \AES_ENC/u0/u0/U87  ( .A1(\AES_ENC/u0/u0/n617 ), .A2(\AES_ENC/u0/u0/n569 ), .ZN(\AES_ENC/u0/u0/n721 ) );
NOR2_X2 \AES_ENC/u0/u0/U86  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n1096 ), .ZN(\AES_ENC/u0/u0/n722 ) );
NOR2_X2 \AES_ENC/u0/u0/U81  ( .A1(\AES_ENC/u0/u0/n1031 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n723 ) );
NOR4_X2 \AES_ENC/u0/u0/U80  ( .A1(\AES_ENC/u0/u0/n724 ), .A2(\AES_ENC/u0/u0/n723 ), .A3(\AES_ENC/u0/u0/n722 ), .A4(\AES_ENC/u0/u0/n721 ), .ZN(\AES_ENC/u0/u0/n725 ) );
NOR2_X2 \AES_ENC/u0/u0/U79  ( .A1(\AES_ENC/u0/u0/n911 ), .A2(\AES_ENC/u0/u0/n990 ), .ZN(\AES_ENC/u0/u0/n1009 ) );
NOR2_X2 \AES_ENC/u0/u0/U78  ( .A1(\AES_ENC/u0/u0/n1013 ), .A2(\AES_ENC/u0/u0/n573 ), .ZN(\AES_ENC/u0/u0/n1014 ) );
NOR2_X2 \AES_ENC/u0/u0/U74  ( .A1(\AES_ENC/u0/u0/n1014 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n1015 ) );
NOR4_X2 \AES_ENC/u0/u0/U73  ( .A1(\AES_ENC/u0/u0/n1016 ), .A2(\AES_ENC/u0/u0/n1015 ), .A3(\AES_ENC/u0/u0/n1119 ), .A4(\AES_ENC/u0/u0/n1046 ), .ZN(\AES_ENC/u0/u0/n1017 ) );
NOR2_X2 \AES_ENC/u0/u0/U72  ( .A1(\AES_ENC/u0/u0/n606 ), .A2(\AES_ENC/u0/u0/n589 ), .ZN(\AES_ENC/u0/u0/n997 ) );
NOR2_X2 \AES_ENC/u0/u0/U71  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n577 ), .ZN(\AES_ENC/u0/u0/n1000 ) );
NOR2_X2 \AES_ENC/u0/u0/U65  ( .A1(\AES_ENC/u0/u0/n616 ), .A2(\AES_ENC/u0/u0/n1096 ), .ZN(\AES_ENC/u0/u0/n999 ) );
NOR4_X2 \AES_ENC/u0/u0/U64  ( .A1(\AES_ENC/u0/u0/n1000 ), .A2(\AES_ENC/u0/u0/n999 ), .A3(\AES_ENC/u0/u0/n998 ), .A4(\AES_ENC/u0/u0/n997 ), .ZN(\AES_ENC/u0/u0/n1001 ) );
NOR2_X2 \AES_ENC/u0/u0/U63  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n1096 ), .ZN(\AES_ENC/u0/u0/n697 ) );
NOR2_X2 \AES_ENC/u0/u0/U62  ( .A1(\AES_ENC/u0/u0/n620 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n958 ) );
NOR2_X2 \AES_ENC/u0/u0/U61  ( .A1(\AES_ENC/u0/u0/n911 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n983 ) );
NOR2_X2 \AES_ENC/u0/u0/U59  ( .A1(\AES_ENC/u0/u0/n1054 ), .A2(\AES_ENC/u0/u0/n1103 ), .ZN(\AES_ENC/u0/u0/n1031 ) );
INV_X4 \AES_ENC/u0/u0/U58  ( .A(\AES_ENC/u0/u0/n1050 ), .ZN(\AES_ENC/u0/u0/n612 ) );
INV_X4 \AES_ENC/u0/u0/U57  ( .A(\AES_ENC/u0/u0/n1072 ), .ZN(\AES_ENC/u0/u0/n605 ) );
INV_X4 \AES_ENC/u0/u0/U50  ( .A(\AES_ENC/u0/u0/n1073 ), .ZN(\AES_ENC/u0/u0/n604 ) );
NOR2_X2 \AES_ENC/u0/u0/U49  ( .A1(\AES_ENC/u0/u0/n582 ), .A2(\AES_ENC/u0/u0/n613 ), .ZN(\AES_ENC/u0/u0/n880 ) );
NOR3_X2 \AES_ENC/u0/u0/U48  ( .A1(\AES_ENC/u0/u0/n826 ), .A2(\AES_ENC/u0/u0/n1121 ), .A3(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n946 ) );
INV_X4 \AES_ENC/u0/u0/U47  ( .A(\AES_ENC/u0/u0/n1010 ), .ZN(\AES_ENC/u0/u0/n608 ) );
NOR3_X2 \AES_ENC/u0/u0/U46  ( .A1(\AES_ENC/u0/u0/n573 ), .A2(\AES_ENC/u0/u0/n1029 ), .A3(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n1119 ) );
INV_X4 \AES_ENC/u0/u0/U45  ( .A(\AES_ENC/u0/u0/n956 ), .ZN(\AES_ENC/u0/u0/n615 ) );
NOR2_X2 \AES_ENC/u0/u0/U44  ( .A1(\AES_ENC/u0/u0/n623 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n1013 ) );
NOR2_X2 \AES_ENC/u0/u0/U43  ( .A1(\AES_ENC/u0/u0/n620 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n910 ) );
NOR2_X2 \AES_ENC/u0/u0/U42  ( .A1(\AES_ENC/u0/u0/n569 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n1091 ) );
NOR2_X2 \AES_ENC/u0/u0/U41  ( .A1(\AES_ENC/u0/u0/n622 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n990 ) );
NOR2_X2 \AES_ENC/u0/u0/U36  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/u0/u0/n1121 ), .ZN(\AES_ENC/u0/u0/n996 ) );
NOR2_X2 \AES_ENC/u0/u0/U35  ( .A1(\AES_ENC/u0/u0/n610 ), .A2(\AES_ENC/u0/u0/n600 ), .ZN(\AES_ENC/u0/u0/n628 ) );
NOR2_X2 \AES_ENC/u0/u0/U34  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n1117 ), .ZN(\AES_ENC/u0/u0/n1118 ) );
NOR2_X2 \AES_ENC/u0/u0/U33  ( .A1(\AES_ENC/u0/u0/n1119 ), .A2(\AES_ENC/u0/u0/n1118 ), .ZN(\AES_ENC/u0/u0/n1127 ) );
NOR2_X2 \AES_ENC/u0/u0/U32  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n594 ), .ZN(\AES_ENC/u0/u0/n629 ) );
NOR2_X2 \AES_ENC/u0/u0/U31  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n906 ), .ZN(\AES_ENC/u0/u0/n909 ) );
NOR2_X2 \AES_ENC/u0/u0/U30  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n597 ), .ZN(\AES_ENC/u0/u0/n658 ) );
NOR2_X2 \AES_ENC/u0/u0/U29  ( .A1(\AES_ENC/u0/u0/n1116 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n695 ) );
NOR2_X2 \AES_ENC/u0/u0/U24  ( .A1(\AES_ENC/u0/u0/n941 ), .A2(\AES_ENC/u0/u0/n608 ), .ZN(\AES_ENC/u0/u0/n724 ) );
NOR2_X2 \AES_ENC/u0/u0/U23  ( .A1(\AES_ENC/u0/u0/n576 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n840 ) );
NOR2_X2 \AES_ENC/u0/u0/U21  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n593 ), .ZN(\AES_ENC/u0/u0/n633 ) );
NOR2_X2 \AES_ENC/u0/u0/U20  ( .A1(\AES_ENC/u0/u0/n1009 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n960 ) );
NOR2_X2 \AES_ENC/u0/u0/U19  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n1045 ), .ZN(\AES_ENC/u0/u0/n812 ) );
NOR2_X2 \AES_ENC/u0/u0/U18  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n1080 ), .ZN(\AES_ENC/u0/u0/n1081 ) );
NOR2_X2 \AES_ENC/u0/u0/U17  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n601 ), .ZN(\AES_ENC/u0/u0/n982 ) );
NOR2_X2 \AES_ENC/u0/u0/U16  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n594 ), .ZN(\AES_ENC/u0/u0/n757 ) );
NOR2_X2 \AES_ENC/u0/u0/U15  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n590 ), .ZN(\AES_ENC/u0/u0/n698 ) );
NOR2_X2 \AES_ENC/u0/u0/U10  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n619 ), .ZN(\AES_ENC/u0/u0/n708 ) );
NOR2_X2 \AES_ENC/u0/u0/U9  ( .A1(\AES_ENC/u0/u0/n619 ), .A2(\AES_ENC/u0/u0/n604 ), .ZN(\AES_ENC/u0/u0/n803 ) );
NOR2_X2 \AES_ENC/u0/u0/U8  ( .A1(\AES_ENC/u0/u0/n615 ), .A2(\AES_ENC/u0/u0/n582 ), .ZN(\AES_ENC/u0/u0/n867 ) );
NOR2_X2 \AES_ENC/u0/u0/U7  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n599 ), .ZN(\AES_ENC/u0/u0/n804 ) );
NOR2_X2 \AES_ENC/u0/u0/U6  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n620 ), .ZN(\AES_ENC/u0/u0/n1046 ) );
OR2_X4 \AES_ENC/u0/u0/U5  ( .A1(\AES_ENC/u0/u0/n624 ), .A2(\AES_ENC/w3[17] ),.ZN(\AES_ENC/u0/u0/n570 ) );
OR2_X4 \AES_ENC/u0/u0/U4  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/w3[20] ),.ZN(\AES_ENC/u0/u0/n569 ) );
NAND2_X2 \AES_ENC/u0/u0/U514  ( .A1(\AES_ENC/u0/u0/n1121 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n1030 ) );
AND2_X2 \AES_ENC/u0/u0/U513  ( .A1(\AES_ENC/u0/u0/n597 ), .A2(\AES_ENC/u0/u0/n1030 ), .ZN(\AES_ENC/u0/u0/n1049 ) );
NAND2_X2 \AES_ENC/u0/u0/U511  ( .A1(\AES_ENC/u0/u0/n1049 ), .A2(\AES_ENC/u0/u0/n794 ), .ZN(\AES_ENC/u0/u0/n637 ) );
AND2_X2 \AES_ENC/u0/u0/U493  ( .A1(\AES_ENC/u0/u0/n779 ), .A2(\AES_ENC/u0/u0/n996 ), .ZN(\AES_ENC/u0/u0/n632 ) );
NAND4_X2 \AES_ENC/u0/u0/U485  ( .A1(\AES_ENC/u0/u0/n637 ), .A2(\AES_ENC/u0/u0/n636 ), .A3(\AES_ENC/u0/u0/n635 ), .A4(\AES_ENC/u0/u0/n634 ), .ZN(\AES_ENC/u0/u0/n638 ) );
NAND2_X2 \AES_ENC/u0/u0/U484  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n638 ), .ZN(\AES_ENC/u0/u0/n679 ) );
NAND2_X2 \AES_ENC/u0/u0/U481  ( .A1(\AES_ENC/u0/u0/n1094 ), .A2(\AES_ENC/u0/u0/n591 ), .ZN(\AES_ENC/u0/u0/n648 ) );
NAND2_X2 \AES_ENC/u0/u0/U476  ( .A1(\AES_ENC/u0/u0/n601 ), .A2(\AES_ENC/u0/u0/n590 ), .ZN(\AES_ENC/u0/u0/n762 ) );
NAND2_X2 \AES_ENC/u0/u0/U475  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n762 ), .ZN(\AES_ENC/u0/u0/n647 ) );
NAND4_X2 \AES_ENC/u0/u0/U457  ( .A1(\AES_ENC/u0/u0/n648 ), .A2(\AES_ENC/u0/u0/n647 ), .A3(\AES_ENC/u0/u0/n646 ), .A4(\AES_ENC/u0/u0/n645 ), .ZN(\AES_ENC/u0/u0/n649 ) );
NAND2_X2 \AES_ENC/u0/u0/U456  ( .A1(\AES_ENC/w3[16] ), .A2(\AES_ENC/u0/u0/n649 ), .ZN(\AES_ENC/u0/u0/n665 ) );
NAND2_X2 \AES_ENC/u0/u0/U454  ( .A1(\AES_ENC/u0/u0/n596 ), .A2(\AES_ENC/u0/u0/n623 ), .ZN(\AES_ENC/u0/u0/n855 ) );
NAND2_X2 \AES_ENC/u0/u0/U453  ( .A1(\AES_ENC/u0/u0/n587 ), .A2(\AES_ENC/u0/u0/n855 ), .ZN(\AES_ENC/u0/u0/n821 ) );
NAND2_X2 \AES_ENC/u0/u0/U452  ( .A1(\AES_ENC/u0/u0/n1093 ), .A2(\AES_ENC/u0/u0/n821 ), .ZN(\AES_ENC/u0/u0/n662 ) );
NAND2_X2 \AES_ENC/u0/u0/U451  ( .A1(\AES_ENC/u0/u0/n619 ), .A2(\AES_ENC/u0/u0/n589 ), .ZN(\AES_ENC/u0/u0/n650 ) );
NAND2_X2 \AES_ENC/u0/u0/U450  ( .A1(\AES_ENC/u0/u0/n956 ), .A2(\AES_ENC/u0/u0/n650 ), .ZN(\AES_ENC/u0/u0/n661 ) );
NAND2_X2 \AES_ENC/u0/u0/U449  ( .A1(\AES_ENC/u0/u0/n626 ), .A2(\AES_ENC/u0/u0/n627 ), .ZN(\AES_ENC/u0/u0/n839 ) );
OR2_X2 \AES_ENC/u0/u0/U446  ( .A1(\AES_ENC/u0/u0/n839 ), .A2(\AES_ENC/u0/u0/n932 ), .ZN(\AES_ENC/u0/u0/n656 ) );
NAND2_X2 \AES_ENC/u0/u0/U445  ( .A1(\AES_ENC/u0/u0/n621 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n1096 ) );
NAND2_X2 \AES_ENC/u0/u0/U444  ( .A1(\AES_ENC/u0/u0/n1030 ), .A2(\AES_ENC/u0/u0/n1096 ), .ZN(\AES_ENC/u0/u0/n651 ) );
NAND2_X2 \AES_ENC/u0/u0/U443  ( .A1(\AES_ENC/u0/u0/n1114 ), .A2(\AES_ENC/u0/u0/n651 ), .ZN(\AES_ENC/u0/u0/n655 ) );
OR3_X2 \AES_ENC/u0/u0/U440  ( .A1(\AES_ENC/u0/u0/n1079 ), .A2(\AES_ENC/w3[23] ), .A3(\AES_ENC/u0/u0/n626 ), .ZN(\AES_ENC/u0/u0/n654 ) );
NAND2_X2 \AES_ENC/u0/u0/U439  ( .A1(\AES_ENC/u0/u0/n593 ), .A2(\AES_ENC/u0/u0/n601 ), .ZN(\AES_ENC/u0/u0/n652 ) );
NAND4_X2 \AES_ENC/u0/u0/U437  ( .A1(\AES_ENC/u0/u0/n656 ), .A2(\AES_ENC/u0/u0/n655 ), .A3(\AES_ENC/u0/u0/n654 ), .A4(\AES_ENC/u0/u0/n653 ), .ZN(\AES_ENC/u0/u0/n657 ) );
NAND2_X2 \AES_ENC/u0/u0/U436  ( .A1(\AES_ENC/w3[18] ), .A2(\AES_ENC/u0/u0/n657 ), .ZN(\AES_ENC/u0/u0/n660 ) );
NAND4_X2 \AES_ENC/u0/u0/U432  ( .A1(\AES_ENC/u0/u0/n662 ), .A2(\AES_ENC/u0/u0/n661 ), .A3(\AES_ENC/u0/u0/n660 ), .A4(\AES_ENC/u0/u0/n659 ), .ZN(\AES_ENC/u0/u0/n663 ) );
NAND2_X2 \AES_ENC/u0/u0/U431  ( .A1(\AES_ENC/u0/u0/n663 ), .A2(\AES_ENC/u0/u0/n574 ), .ZN(\AES_ENC/u0/u0/n664 ) );
NAND2_X2 \AES_ENC/u0/u0/U430  ( .A1(\AES_ENC/u0/u0/n665 ), .A2(\AES_ENC/u0/u0/n664 ), .ZN(\AES_ENC/u0/u0/n666 ) );
NAND2_X2 \AES_ENC/u0/u0/U429  ( .A1(\AES_ENC/w3[22] ), .A2(\AES_ENC/u0/u0/n666 ), .ZN(\AES_ENC/u0/u0/n678 ) );
NAND2_X2 \AES_ENC/u0/u0/U426  ( .A1(\AES_ENC/u0/u0/n735 ), .A2(\AES_ENC/u0/u0/n1093 ), .ZN(\AES_ENC/u0/u0/n675 ) );
NAND2_X2 \AES_ENC/u0/u0/U425  ( .A1(\AES_ENC/u0/u0/n588 ), .A2(\AES_ENC/u0/u0/n597 ), .ZN(\AES_ENC/u0/u0/n1045 ) );
OR2_X2 \AES_ENC/u0/u0/U424  ( .A1(\AES_ENC/u0/u0/n1045 ), .A2(\AES_ENC/u0/u0/n605 ), .ZN(\AES_ENC/u0/u0/n674 ) );
NAND2_X2 \AES_ENC/u0/u0/U423  ( .A1(\AES_ENC/w3[17] ), .A2(\AES_ENC/u0/u0/n620 ), .ZN(\AES_ENC/u0/u0/n667 ) );
NAND2_X2 \AES_ENC/u0/u0/U422  ( .A1(\AES_ENC/u0/u0/n619 ), .A2(\AES_ENC/u0/u0/n667 ), .ZN(\AES_ENC/u0/u0/n1071 ) );
NAND4_X2 \AES_ENC/u0/u0/U412  ( .A1(\AES_ENC/u0/u0/n675 ), .A2(\AES_ENC/u0/u0/n674 ), .A3(\AES_ENC/u0/u0/n673 ), .A4(\AES_ENC/u0/u0/n672 ), .ZN(\AES_ENC/u0/u0/n676 ) );
NAND2_X2 \AES_ENC/u0/u0/U411  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n676 ), .ZN(\AES_ENC/u0/u0/n677 ) );
NAND2_X2 \AES_ENC/u0/u0/U408  ( .A1(\AES_ENC/u0/u0/n800 ), .A2(\AES_ENC/u0/u0/n1022 ), .ZN(\AES_ENC/u0/u0/n680 ) );
NAND2_X2 \AES_ENC/u0/u0/U407  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n680 ), .ZN(\AES_ENC/u0/u0/n681 ) );
AND2_X2 \AES_ENC/u0/u0/U402  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n684 ), .ZN(\AES_ENC/u0/u0/n682 ) );
NAND4_X2 \AES_ENC/u0/u0/U395  ( .A1(\AES_ENC/u0/u0/n691 ), .A2(\AES_ENC/u0/u0/n581 ), .A3(\AES_ENC/u0/u0/n690 ), .A4(\AES_ENC/u0/u0/n689 ), .ZN(\AES_ENC/u0/u0/n692 ) );
NAND2_X2 \AES_ENC/u0/u0/U394  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n692 ), .ZN(\AES_ENC/u0/u0/n733 ) );
NAND2_X2 \AES_ENC/u0/u0/U392  ( .A1(\AES_ENC/u0/u0/n977 ), .A2(\AES_ENC/u0/u0/n1050 ), .ZN(\AES_ENC/u0/u0/n702 ) );
NAND2_X2 \AES_ENC/u0/u0/U391  ( .A1(\AES_ENC/u0/u0/n1093 ), .A2(\AES_ENC/u0/u0/n1045 ), .ZN(\AES_ENC/u0/u0/n701 ) );
NAND4_X2 \AES_ENC/u0/u0/U381  ( .A1(\AES_ENC/u0/u0/n702 ), .A2(\AES_ENC/u0/u0/n701 ), .A3(\AES_ENC/u0/u0/n700 ), .A4(\AES_ENC/u0/u0/n699 ), .ZN(\AES_ENC/u0/u0/n703 ) );
NAND2_X2 \AES_ENC/u0/u0/U380  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n703 ), .ZN(\AES_ENC/u0/u0/n732 ) );
AND2_X2 \AES_ENC/u0/u0/U379  ( .A1(\AES_ENC/w3[16] ), .A2(\AES_ENC/w3[22] ),.ZN(\AES_ENC/u0/u0/n1113 ) );
NAND2_X2 \AES_ENC/u0/u0/U378  ( .A1(\AES_ENC/u0/u0/n601 ), .A2(\AES_ENC/u0/u0/n1030 ), .ZN(\AES_ENC/u0/u0/n881 ) );
NAND2_X2 \AES_ENC/u0/u0/U377  ( .A1(\AES_ENC/u0/u0/n1093 ), .A2(\AES_ENC/u0/u0/n881 ), .ZN(\AES_ENC/u0/u0/n715 ) );
NAND2_X2 \AES_ENC/u0/u0/U376  ( .A1(\AES_ENC/u0/u0/n1010 ), .A2(\AES_ENC/u0/u0/n600 ), .ZN(\AES_ENC/u0/u0/n714 ) );
NAND2_X2 \AES_ENC/u0/u0/U375  ( .A1(\AES_ENC/u0/u0/n855 ), .A2(\AES_ENC/u0/u0/n588 ), .ZN(\AES_ENC/u0/u0/n1117 ) );
XNOR2_X2 \AES_ENC/u0/u0/U371  ( .A(\AES_ENC/u0/u0/n611 ), .B(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n824 ) );
NAND4_X2 \AES_ENC/u0/u0/U362  ( .A1(\AES_ENC/u0/u0/n715 ), .A2(\AES_ENC/u0/u0/n714 ), .A3(\AES_ENC/u0/u0/n713 ), .A4(\AES_ENC/u0/u0/n712 ), .ZN(\AES_ENC/u0/u0/n716 ) );
NAND2_X2 \AES_ENC/u0/u0/U361  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n716 ), .ZN(\AES_ENC/u0/u0/n731 ) );
AND2_X2 \AES_ENC/u0/u0/U360  ( .A1(\AES_ENC/w3[22] ), .A2(\AES_ENC/u0/u0/n574 ), .ZN(\AES_ENC/u0/u0/n1131 ) );
NAND2_X2 \AES_ENC/u0/u0/U359  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n717 ) );
NAND2_X2 \AES_ENC/u0/u0/U358  ( .A1(\AES_ENC/u0/u0/n1029 ), .A2(\AES_ENC/u0/u0/n717 ), .ZN(\AES_ENC/u0/u0/n728 ) );
NAND2_X2 \AES_ENC/u0/u0/U357  ( .A1(\AES_ENC/w3[17] ), .A2(\AES_ENC/u0/u0/n624 ), .ZN(\AES_ENC/u0/u0/n1097 ) );
NAND2_X2 \AES_ENC/u0/u0/U356  ( .A1(\AES_ENC/u0/u0/n603 ), .A2(\AES_ENC/u0/u0/n1097 ), .ZN(\AES_ENC/u0/u0/n718 ) );
NAND2_X2 \AES_ENC/u0/u0/U355  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n718 ), .ZN(\AES_ENC/u0/u0/n727 ) );
NAND4_X2 \AES_ENC/u0/u0/U344  ( .A1(\AES_ENC/u0/u0/n728 ), .A2(\AES_ENC/u0/u0/n727 ), .A3(\AES_ENC/u0/u0/n726 ), .A4(\AES_ENC/u0/u0/n725 ), .ZN(\AES_ENC/u0/u0/n729 ) );
NAND2_X2 \AES_ENC/u0/u0/U343  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n729 ), .ZN(\AES_ENC/u0/u0/n730 ) );
NAND4_X2 \AES_ENC/u0/u0/U342  ( .A1(\AES_ENC/u0/u0/n733 ), .A2(\AES_ENC/u0/u0/n732 ), .A3(\AES_ENC/u0/u0/n731 ), .A4(\AES_ENC/u0/u0/n730 ), .ZN(\AES_ENC/u0/subword[25] ) );
NAND2_X2 \AES_ENC/u0/u0/U341  ( .A1(\AES_ENC/w3[23] ), .A2(\AES_ENC/u0/u0/n611 ), .ZN(\AES_ENC/u0/u0/n734 ) );
NAND2_X2 \AES_ENC/u0/u0/U340  ( .A1(\AES_ENC/u0/u0/n734 ), .A2(\AES_ENC/u0/u0/n607 ), .ZN(\AES_ENC/u0/u0/n738 ) );
OR4_X2 \AES_ENC/u0/u0/U339  ( .A1(\AES_ENC/u0/u0/n738 ), .A2(\AES_ENC/u0/u0/n626 ), .A3(\AES_ENC/u0/u0/n826 ), .A4(\AES_ENC/u0/u0/n1121 ), .ZN(\AES_ENC/u0/u0/n746 ) );
NAND2_X2 \AES_ENC/u0/u0/U337  ( .A1(\AES_ENC/u0/u0/n1100 ), .A2(\AES_ENC/u0/u0/n587 ), .ZN(\AES_ENC/u0/u0/n992 ) );
OR2_X2 \AES_ENC/u0/u0/U336  ( .A1(\AES_ENC/u0/u0/n610 ), .A2(\AES_ENC/u0/u0/n735 ), .ZN(\AES_ENC/u0/u0/n737 ) );
NAND2_X2 \AES_ENC/u0/u0/U334  ( .A1(\AES_ENC/u0/u0/n619 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n753 ) );
NAND2_X2 \AES_ENC/u0/u0/U333  ( .A1(\AES_ENC/u0/u0/n582 ), .A2(\AES_ENC/u0/u0/n753 ), .ZN(\AES_ENC/u0/u0/n1080 ) );
NAND2_X2 \AES_ENC/u0/u0/U332  ( .A1(\AES_ENC/u0/u0/n1048 ), .A2(\AES_ENC/u0/u0/n576 ), .ZN(\AES_ENC/u0/u0/n736 ) );
NAND2_X2 \AES_ENC/u0/u0/U331  ( .A1(\AES_ENC/u0/u0/n737 ), .A2(\AES_ENC/u0/u0/n736 ), .ZN(\AES_ENC/u0/u0/n739 ) );
NAND2_X2 \AES_ENC/u0/u0/U330  ( .A1(\AES_ENC/u0/u0/n739 ), .A2(\AES_ENC/u0/u0/n738 ), .ZN(\AES_ENC/u0/u0/n745 ) );
NAND2_X2 \AES_ENC/u0/u0/U326  ( .A1(\AES_ENC/u0/u0/n1096 ), .A2(\AES_ENC/u0/u0/n590 ), .ZN(\AES_ENC/u0/u0/n906 ) );
NAND4_X2 \AES_ENC/u0/u0/U323  ( .A1(\AES_ENC/u0/u0/n746 ), .A2(\AES_ENC/u0/u0/n992 ), .A3(\AES_ENC/u0/u0/n745 ), .A4(\AES_ENC/u0/u0/n744 ), .ZN(\AES_ENC/u0/u0/n747 ) );
NAND2_X2 \AES_ENC/u0/u0/U322  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n747 ), .ZN(\AES_ENC/u0/u0/n793 ) );
NAND2_X2 \AES_ENC/u0/u0/U321  ( .A1(\AES_ENC/u0/u0/n584 ), .A2(\AES_ENC/u0/u0/n855 ), .ZN(\AES_ENC/u0/u0/n748 ) );
NAND2_X2 \AES_ENC/u0/u0/U320  ( .A1(\AES_ENC/u0/u0/n956 ), .A2(\AES_ENC/u0/u0/n748 ), .ZN(\AES_ENC/u0/u0/n760 ) );
NAND2_X2 \AES_ENC/u0/u0/U313  ( .A1(\AES_ENC/u0/u0/n590 ), .A2(\AES_ENC/u0/u0/n753 ), .ZN(\AES_ENC/u0/u0/n1023 ) );
NAND4_X2 \AES_ENC/u0/u0/U308  ( .A1(\AES_ENC/u0/u0/n760 ), .A2(\AES_ENC/u0/u0/n992 ), .A3(\AES_ENC/u0/u0/n759 ), .A4(\AES_ENC/u0/u0/n758 ), .ZN(\AES_ENC/u0/u0/n761 ) );
NAND2_X2 \AES_ENC/u0/u0/U307  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n761 ), .ZN(\AES_ENC/u0/u0/n792 ) );
NAND2_X2 \AES_ENC/u0/u0/U306  ( .A1(\AES_ENC/u0/u0/n584 ), .A2(\AES_ENC/u0/u0/n603 ), .ZN(\AES_ENC/u0/u0/n989 ) );
NAND2_X2 \AES_ENC/u0/u0/U305  ( .A1(\AES_ENC/u0/u0/n1050 ), .A2(\AES_ENC/u0/u0/n989 ), .ZN(\AES_ENC/u0/u0/n777 ) );
NAND2_X2 \AES_ENC/u0/u0/U304  ( .A1(\AES_ENC/u0/u0/n1093 ), .A2(\AES_ENC/u0/u0/n762 ), .ZN(\AES_ENC/u0/u0/n776 ) );
XNOR2_X2 \AES_ENC/u0/u0/U301  ( .A(\AES_ENC/w3[23] ), .B(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n959 ) );
NAND4_X2 \AES_ENC/u0/u0/U289  ( .A1(\AES_ENC/u0/u0/n777 ), .A2(\AES_ENC/u0/u0/n776 ), .A3(\AES_ENC/u0/u0/n775 ), .A4(\AES_ENC/u0/u0/n774 ), .ZN(\AES_ENC/u0/u0/n778 ) );
NAND2_X2 \AES_ENC/u0/u0/U288  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n778 ), .ZN(\AES_ENC/u0/u0/n791 ) );
NAND2_X2 \AES_ENC/u0/u0/U287  ( .A1(\AES_ENC/u0/u0/n1056 ), .A2(\AES_ENC/u0/u0/n1050 ), .ZN(\AES_ENC/u0/u0/n788 ) );
NAND2_X2 \AES_ENC/u0/u0/U286  ( .A1(\AES_ENC/u0/u0/n1091 ), .A2(\AES_ENC/u0/u0/n779 ), .ZN(\AES_ENC/u0/u0/n787 ) );
NAND2_X2 \AES_ENC/u0/u0/U285  ( .A1(\AES_ENC/u0/u0/n956 ), .A2(\AES_ENC/w3[17] ), .ZN(\AES_ENC/u0/u0/n786 ) );
NAND4_X2 \AES_ENC/u0/u0/U278  ( .A1(\AES_ENC/u0/u0/n788 ), .A2(\AES_ENC/u0/u0/n787 ), .A3(\AES_ENC/u0/u0/n786 ), .A4(\AES_ENC/u0/u0/n785 ), .ZN(\AES_ENC/u0/u0/n789 ) );
NAND2_X2 \AES_ENC/u0/u0/U277  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n789 ), .ZN(\AES_ENC/u0/u0/n790 ) );
NAND4_X2 \AES_ENC/u0/u0/U276  ( .A1(\AES_ENC/u0/u0/n793 ), .A2(\AES_ENC/u0/u0/n792 ), .A3(\AES_ENC/u0/u0/n791 ), .A4(\AES_ENC/u0/u0/n790 ), .ZN(\AES_ENC/u0/subword[26] ) );
NAND2_X2 \AES_ENC/u0/u0/U275  ( .A1(\AES_ENC/u0/u0/n1059 ), .A2(\AES_ENC/u0/u0/n794 ), .ZN(\AES_ENC/u0/u0/n810 ) );
NAND2_X2 \AES_ENC/u0/u0/U274  ( .A1(\AES_ENC/u0/u0/n1049 ), .A2(\AES_ENC/u0/u0/n956 ), .ZN(\AES_ENC/u0/u0/n809 ) );
OR2_X2 \AES_ENC/u0/u0/U266  ( .A1(\AES_ENC/u0/u0/n1096 ), .A2(\AES_ENC/u0/u0/n606 ), .ZN(\AES_ENC/u0/u0/n802 ) );
NAND2_X2 \AES_ENC/u0/u0/U265  ( .A1(\AES_ENC/u0/u0/n1053 ), .A2(\AES_ENC/u0/u0/n800 ), .ZN(\AES_ENC/u0/u0/n801 ) );
NAND2_X2 \AES_ENC/u0/u0/U264  ( .A1(\AES_ENC/u0/u0/n802 ), .A2(\AES_ENC/u0/u0/n801 ), .ZN(\AES_ENC/u0/u0/n805 ) );
NAND4_X2 \AES_ENC/u0/u0/U261  ( .A1(\AES_ENC/u0/u0/n810 ), .A2(\AES_ENC/u0/u0/n809 ), .A3(\AES_ENC/u0/u0/n808 ), .A4(\AES_ENC/u0/u0/n807 ), .ZN(\AES_ENC/u0/u0/n811 ) );
NAND2_X2 \AES_ENC/u0/u0/U260  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n811 ), .ZN(\AES_ENC/u0/u0/n852 ) );
OR2_X2 \AES_ENC/u0/u0/U259  ( .A1(\AES_ENC/u0/u0/n1023 ), .A2(\AES_ENC/u0/u0/n617 ), .ZN(\AES_ENC/u0/u0/n819 ) );
OR2_X2 \AES_ENC/u0/u0/U257  ( .A1(\AES_ENC/u0/u0/n570 ), .A2(\AES_ENC/u0/u0/n930 ), .ZN(\AES_ENC/u0/u0/n818 ) );
NAND2_X2 \AES_ENC/u0/u0/U256  ( .A1(\AES_ENC/u0/u0/n1013 ), .A2(\AES_ENC/u0/u0/n1094 ), .ZN(\AES_ENC/u0/u0/n817 ) );
NAND4_X2 \AES_ENC/u0/u0/U249  ( .A1(\AES_ENC/u0/u0/n819 ), .A2(\AES_ENC/u0/u0/n818 ), .A3(\AES_ENC/u0/u0/n817 ), .A4(\AES_ENC/u0/u0/n816 ), .ZN(\AES_ENC/u0/u0/n820 ) );
NAND2_X2 \AES_ENC/u0/u0/U248  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n820 ), .ZN(\AES_ENC/u0/u0/n851 ) );
NAND2_X2 \AES_ENC/u0/u0/U247  ( .A1(\AES_ENC/u0/u0/n956 ), .A2(\AES_ENC/u0/u0/n1080 ), .ZN(\AES_ENC/u0/u0/n835 ) );
NAND2_X2 \AES_ENC/u0/u0/U246  ( .A1(\AES_ENC/u0/u0/n570 ), .A2(\AES_ENC/u0/u0/n1030 ), .ZN(\AES_ENC/u0/u0/n1047 ) );
OR2_X2 \AES_ENC/u0/u0/U245  ( .A1(\AES_ENC/u0/u0/n1047 ), .A2(\AES_ENC/u0/u0/n612 ), .ZN(\AES_ENC/u0/u0/n834 ) );
NAND2_X2 \AES_ENC/u0/u0/U244  ( .A1(\AES_ENC/u0/u0/n1072 ), .A2(\AES_ENC/u0/u0/n589 ), .ZN(\AES_ENC/u0/u0/n833 ) );
NAND4_X2 \AES_ENC/u0/u0/U233  ( .A1(\AES_ENC/u0/u0/n835 ), .A2(\AES_ENC/u0/u0/n834 ), .A3(\AES_ENC/u0/u0/n833 ), .A4(\AES_ENC/u0/u0/n832 ), .ZN(\AES_ENC/u0/u0/n836 ) );
NAND2_X2 \AES_ENC/u0/u0/U232  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n836 ), .ZN(\AES_ENC/u0/u0/n850 ) );
NAND2_X2 \AES_ENC/u0/u0/U231  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n623 ), .ZN(\AES_ENC/u0/u0/n847 ) );
NAND2_X2 \AES_ENC/u0/u0/U230  ( .A1(\AES_ENC/u0/u0/n1050 ), .A2(\AES_ENC/u0/u0/n1071 ), .ZN(\AES_ENC/u0/u0/n846 ) );
OR2_X2 \AES_ENC/u0/u0/U224  ( .A1(\AES_ENC/u0/u0/n1053 ), .A2(\AES_ENC/u0/u0/n911 ), .ZN(\AES_ENC/u0/u0/n1077 ) );
NAND4_X2 \AES_ENC/u0/u0/U220  ( .A1(\AES_ENC/u0/u0/n847 ), .A2(\AES_ENC/u0/u0/n846 ), .A3(\AES_ENC/u0/u0/n845 ), .A4(\AES_ENC/u0/u0/n844 ), .ZN(\AES_ENC/u0/u0/n848 ) );
NAND2_X2 \AES_ENC/u0/u0/U219  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n848 ), .ZN(\AES_ENC/u0/u0/n849 ) );
NAND4_X2 \AES_ENC/u0/u0/U218  ( .A1(\AES_ENC/u0/u0/n852 ), .A2(\AES_ENC/u0/u0/n851 ), .A3(\AES_ENC/u0/u0/n850 ), .A4(\AES_ENC/u0/u0/n849 ), .ZN(\AES_ENC/u0/subword[27] ) );
NAND2_X2 \AES_ENC/u0/u0/U216  ( .A1(\AES_ENC/u0/u0/n1009 ), .A2(\AES_ENC/u0/u0/n1072 ), .ZN(\AES_ENC/u0/u0/n862 ) );
NAND2_X2 \AES_ENC/u0/u0/U215  ( .A1(\AES_ENC/u0/u0/n603 ), .A2(\AES_ENC/u0/u0/n577 ), .ZN(\AES_ENC/u0/u0/n853 ) );
NAND2_X2 \AES_ENC/u0/u0/U214  ( .A1(\AES_ENC/u0/u0/n1050 ), .A2(\AES_ENC/u0/u0/n853 ), .ZN(\AES_ENC/u0/u0/n861 ) );
NAND4_X2 \AES_ENC/u0/u0/U206  ( .A1(\AES_ENC/u0/u0/n862 ), .A2(\AES_ENC/u0/u0/n861 ), .A3(\AES_ENC/u0/u0/n860 ), .A4(\AES_ENC/u0/u0/n859 ), .ZN(\AES_ENC/u0/u0/n863 ) );
NAND2_X2 \AES_ENC/u0/u0/U205  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n863 ), .ZN(\AES_ENC/u0/u0/n905 ) );
NAND2_X2 \AES_ENC/u0/u0/U204  ( .A1(\AES_ENC/u0/u0/n1010 ), .A2(\AES_ENC/u0/u0/n989 ), .ZN(\AES_ENC/u0/u0/n874 ) );
NAND2_X2 \AES_ENC/u0/u0/U203  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n610 ), .ZN(\AES_ENC/u0/u0/n864 ) );
NAND2_X2 \AES_ENC/u0/u0/U202  ( .A1(\AES_ENC/u0/u0/n929 ), .A2(\AES_ENC/u0/u0/n864 ), .ZN(\AES_ENC/u0/u0/n873 ) );
NAND4_X2 \AES_ENC/u0/u0/U193  ( .A1(\AES_ENC/u0/u0/n874 ), .A2(\AES_ENC/u0/u0/n873 ), .A3(\AES_ENC/u0/u0/n872 ), .A4(\AES_ENC/u0/u0/n871 ), .ZN(\AES_ENC/u0/u0/n875 ) );
NAND2_X2 \AES_ENC/u0/u0/U192  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n875 ), .ZN(\AES_ENC/u0/u0/n904 ) );
NAND2_X2 \AES_ENC/u0/u0/U191  ( .A1(\AES_ENC/u0/u0/n583 ), .A2(\AES_ENC/u0/u0/n1050 ), .ZN(\AES_ENC/u0/u0/n889 ) );
NAND2_X2 \AES_ENC/u0/u0/U190  ( .A1(\AES_ENC/u0/u0/n1093 ), .A2(\AES_ENC/u0/u0/n587 ), .ZN(\AES_ENC/u0/u0/n876 ) );
NAND2_X2 \AES_ENC/u0/u0/U189  ( .A1(\AES_ENC/u0/u0/n604 ), .A2(\AES_ENC/u0/u0/n876 ), .ZN(\AES_ENC/u0/u0/n877 ) );
NAND2_X2 \AES_ENC/u0/u0/U188  ( .A1(\AES_ENC/u0/u0/n877 ), .A2(\AES_ENC/u0/u0/n623 ), .ZN(\AES_ENC/u0/u0/n888 ) );
NAND4_X2 \AES_ENC/u0/u0/U179  ( .A1(\AES_ENC/u0/u0/n889 ), .A2(\AES_ENC/u0/u0/n888 ), .A3(\AES_ENC/u0/u0/n887 ), .A4(\AES_ENC/u0/u0/n886 ), .ZN(\AES_ENC/u0/u0/n890 ) );
NAND2_X2 \AES_ENC/u0/u0/U178  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n890 ), .ZN(\AES_ENC/u0/u0/n903 ) );
OR2_X2 \AES_ENC/u0/u0/U177  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n1059 ), .ZN(\AES_ENC/u0/u0/n900 ) );
NAND2_X2 \AES_ENC/u0/u0/U176  ( .A1(\AES_ENC/u0/u0/n1073 ), .A2(\AES_ENC/u0/u0/n1047 ), .ZN(\AES_ENC/u0/u0/n899 ) );
NAND2_X2 \AES_ENC/u0/u0/U175  ( .A1(\AES_ENC/u0/u0/n1094 ), .A2(\AES_ENC/u0/u0/n595 ), .ZN(\AES_ENC/u0/u0/n898 ) );
NAND4_X2 \AES_ENC/u0/u0/U167  ( .A1(\AES_ENC/u0/u0/n900 ), .A2(\AES_ENC/u0/u0/n899 ), .A3(\AES_ENC/u0/u0/n898 ), .A4(\AES_ENC/u0/u0/n897 ), .ZN(\AES_ENC/u0/u0/n901 ) );
NAND2_X2 \AES_ENC/u0/u0/U166  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n901 ), .ZN(\AES_ENC/u0/u0/n902 ) );
NAND4_X2 \AES_ENC/u0/u0/U165  ( .A1(\AES_ENC/u0/u0/n905 ), .A2(\AES_ENC/u0/u0/n904 ), .A3(\AES_ENC/u0/u0/n903 ), .A4(\AES_ENC/u0/u0/n902 ), .ZN(\AES_ENC/u0/subword[28] ) );
NAND2_X2 \AES_ENC/u0/u0/U164  ( .A1(\AES_ENC/u0/u0/n1094 ), .A2(\AES_ENC/u0/u0/n599 ), .ZN(\AES_ENC/u0/u0/n922 ) );
NAND2_X2 \AES_ENC/u0/u0/U163  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n989 ), .ZN(\AES_ENC/u0/u0/n921 ) );
NAND4_X2 \AES_ENC/u0/u0/U151  ( .A1(\AES_ENC/u0/u0/n922 ), .A2(\AES_ENC/u0/u0/n921 ), .A3(\AES_ENC/u0/u0/n920 ), .A4(\AES_ENC/u0/u0/n919 ), .ZN(\AES_ENC/u0/u0/n923 ) );
NAND2_X2 \AES_ENC/u0/u0/U150  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n923 ), .ZN(\AES_ENC/u0/u0/n972 ) );
NAND2_X2 \AES_ENC/u0/u0/U149  ( .A1(\AES_ENC/u0/u0/n582 ), .A2(\AES_ENC/u0/u0/n619 ), .ZN(\AES_ENC/u0/u0/n924 ) );
NAND2_X2 \AES_ENC/u0/u0/U148  ( .A1(\AES_ENC/u0/u0/n1073 ), .A2(\AES_ENC/u0/u0/n924 ), .ZN(\AES_ENC/u0/u0/n939 ) );
NAND2_X2 \AES_ENC/u0/u0/U147  ( .A1(\AES_ENC/u0/u0/n926 ), .A2(\AES_ENC/u0/u0/n925 ), .ZN(\AES_ENC/u0/u0/n927 ) );
NAND2_X2 \AES_ENC/u0/u0/U146  ( .A1(\AES_ENC/u0/u0/n606 ), .A2(\AES_ENC/u0/u0/n927 ), .ZN(\AES_ENC/u0/u0/n928 ) );
NAND2_X2 \AES_ENC/u0/u0/U145  ( .A1(\AES_ENC/u0/u0/n928 ), .A2(\AES_ENC/u0/u0/n1080 ), .ZN(\AES_ENC/u0/u0/n938 ) );
OR2_X2 \AES_ENC/u0/u0/U144  ( .A1(\AES_ENC/u0/u0/n1117 ), .A2(\AES_ENC/u0/u0/n615 ), .ZN(\AES_ENC/u0/u0/n937 ) );
NAND4_X2 \AES_ENC/u0/u0/U139  ( .A1(\AES_ENC/u0/u0/n939 ), .A2(\AES_ENC/u0/u0/n938 ), .A3(\AES_ENC/u0/u0/n937 ), .A4(\AES_ENC/u0/u0/n936 ), .ZN(\AES_ENC/u0/u0/n940 ) );
NAND2_X2 \AES_ENC/u0/u0/U138  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n940 ), .ZN(\AES_ENC/u0/u0/n971 ) );
OR2_X2 \AES_ENC/u0/u0/U137  ( .A1(\AES_ENC/u0/u0/n605 ), .A2(\AES_ENC/u0/u0/n941 ), .ZN(\AES_ENC/u0/u0/n954 ) );
NAND2_X2 \AES_ENC/u0/u0/U136  ( .A1(\AES_ENC/u0/u0/n1096 ), .A2(\AES_ENC/u0/u0/n577 ), .ZN(\AES_ENC/u0/u0/n942 ) );
NAND2_X2 \AES_ENC/u0/u0/U135  ( .A1(\AES_ENC/u0/u0/n1048 ), .A2(\AES_ENC/u0/u0/n942 ), .ZN(\AES_ENC/u0/u0/n943 ) );
NAND2_X2 \AES_ENC/u0/u0/U134  ( .A1(\AES_ENC/u0/u0/n612 ), .A2(\AES_ENC/u0/u0/n943 ), .ZN(\AES_ENC/u0/u0/n944 ) );
NAND2_X2 \AES_ENC/u0/u0/U133  ( .A1(\AES_ENC/u0/u0/n944 ), .A2(\AES_ENC/u0/u0/n580 ), .ZN(\AES_ENC/u0/u0/n953 ) );
NAND4_X2 \AES_ENC/u0/u0/U125  ( .A1(\AES_ENC/u0/u0/n954 ), .A2(\AES_ENC/u0/u0/n953 ), .A3(\AES_ENC/u0/u0/n952 ), .A4(\AES_ENC/u0/u0/n951 ), .ZN(\AES_ENC/u0/u0/n955 ) );
NAND2_X2 \AES_ENC/u0/u0/U124  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n955 ), .ZN(\AES_ENC/u0/u0/n970 ) );
NAND2_X2 \AES_ENC/u0/u0/U123  ( .A1(\AES_ENC/u0/u0/n1094 ), .A2(\AES_ENC/u0/u0/n1071 ), .ZN(\AES_ENC/u0/u0/n967 ) );
NAND2_X2 \AES_ENC/u0/u0/U122  ( .A1(\AES_ENC/u0/u0/n956 ), .A2(\AES_ENC/u0/u0/n1030 ), .ZN(\AES_ENC/u0/u0/n966 ) );
NAND4_X2 \AES_ENC/u0/u0/U114  ( .A1(\AES_ENC/u0/u0/n967 ), .A2(\AES_ENC/u0/u0/n966 ), .A3(\AES_ENC/u0/u0/n965 ), .A4(\AES_ENC/u0/u0/n964 ), .ZN(\AES_ENC/u0/u0/n968 ) );
NAND2_X2 \AES_ENC/u0/u0/U113  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n968 ), .ZN(\AES_ENC/u0/u0/n969 ) );
NAND4_X2 \AES_ENC/u0/u0/U112  ( .A1(\AES_ENC/u0/u0/n972 ), .A2(\AES_ENC/u0/u0/n971 ), .A3(\AES_ENC/u0/u0/n970 ), .A4(\AES_ENC/u0/u0/n969 ), .ZN(\AES_ENC/u0/subword[29] ) );
NAND2_X2 \AES_ENC/u0/u0/U111  ( .A1(\AES_ENC/u0/u0/n570 ), .A2(\AES_ENC/u0/u0/n1097 ), .ZN(\AES_ENC/u0/u0/n973 ) );
NAND2_X2 \AES_ENC/u0/u0/U110  ( .A1(\AES_ENC/u0/u0/n1073 ), .A2(\AES_ENC/u0/u0/n973 ), .ZN(\AES_ENC/u0/u0/n987 ) );
NAND2_X2 \AES_ENC/u0/u0/U109  ( .A1(\AES_ENC/u0/u0/n974 ), .A2(\AES_ENC/u0/u0/n1077 ), .ZN(\AES_ENC/u0/u0/n975 ) );
NAND2_X2 \AES_ENC/u0/u0/U108  ( .A1(\AES_ENC/u0/u0/n613 ), .A2(\AES_ENC/u0/u0/n975 ), .ZN(\AES_ENC/u0/u0/n976 ) );
NAND2_X2 \AES_ENC/u0/u0/U107  ( .A1(\AES_ENC/u0/u0/n977 ), .A2(\AES_ENC/u0/u0/n976 ), .ZN(\AES_ENC/u0/u0/n986 ) );
NAND4_X2 \AES_ENC/u0/u0/U99  ( .A1(\AES_ENC/u0/u0/n987 ), .A2(\AES_ENC/u0/u0/n986 ), .A3(\AES_ENC/u0/u0/n985 ), .A4(\AES_ENC/u0/u0/n984 ), .ZN(\AES_ENC/u0/u0/n988 ) );
NAND2_X2 \AES_ENC/u0/u0/U98  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n988 ), .ZN(\AES_ENC/u0/u0/n1044 ) );
NAND2_X2 \AES_ENC/u0/u0/U97  ( .A1(\AES_ENC/u0/u0/n1073 ), .A2(\AES_ENC/u0/u0/n989 ), .ZN(\AES_ENC/u0/u0/n1004 ) );
NAND2_X2 \AES_ENC/u0/u0/U96  ( .A1(\AES_ENC/u0/u0/n1092 ), .A2(\AES_ENC/u0/u0/n619 ), .ZN(\AES_ENC/u0/u0/n1003 ) );
NAND4_X2 \AES_ENC/u0/u0/U85  ( .A1(\AES_ENC/u0/u0/n1004 ), .A2(\AES_ENC/u0/u0/n1003 ), .A3(\AES_ENC/u0/u0/n1002 ), .A4(\AES_ENC/u0/u0/n1001 ), .ZN(\AES_ENC/u0/u0/n1005 ) );
NAND2_X2 \AES_ENC/u0/u0/U84  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n1005 ), .ZN(\AES_ENC/u0/u0/n1043 ) );
NAND2_X2 \AES_ENC/u0/u0/U83  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n596 ), .ZN(\AES_ENC/u0/u0/n1020 ) );
NAND2_X2 \AES_ENC/u0/u0/U82  ( .A1(\AES_ENC/u0/u0/n1050 ), .A2(\AES_ENC/u0/u0/n624 ), .ZN(\AES_ENC/u0/u0/n1019 ) );
NAND2_X2 \AES_ENC/u0/u0/U77  ( .A1(\AES_ENC/u0/u0/n1059 ), .A2(\AES_ENC/u0/u0/n1114 ), .ZN(\AES_ENC/u0/u0/n1012 ) );
NAND2_X2 \AES_ENC/u0/u0/U76  ( .A1(\AES_ENC/u0/u0/n1010 ), .A2(\AES_ENC/u0/u0/n592 ), .ZN(\AES_ENC/u0/u0/n1011 ) );
NAND2_X2 \AES_ENC/u0/u0/U75  ( .A1(\AES_ENC/u0/u0/n1012 ), .A2(\AES_ENC/u0/u0/n1011 ), .ZN(\AES_ENC/u0/u0/n1016 ) );
NAND4_X2 \AES_ENC/u0/u0/U70  ( .A1(\AES_ENC/u0/u0/n1020 ), .A2(\AES_ENC/u0/u0/n1019 ), .A3(\AES_ENC/u0/u0/n1018 ), .A4(\AES_ENC/u0/u0/n1017 ), .ZN(\AES_ENC/u0/u0/n1021 ) );
NAND2_X2 \AES_ENC/u0/u0/U69  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n1021 ), .ZN(\AES_ENC/u0/u0/n1042 ) );
NAND2_X2 \AES_ENC/u0/u0/U68  ( .A1(\AES_ENC/u0/u0/n1022 ), .A2(\AES_ENC/u0/u0/n1093 ), .ZN(\AES_ENC/u0/u0/n1039 ) );
NAND2_X2 \AES_ENC/u0/u0/U67  ( .A1(\AES_ENC/u0/u0/n1050 ), .A2(\AES_ENC/u0/u0/n1023 ), .ZN(\AES_ENC/u0/u0/n1038 ) );
NAND2_X2 \AES_ENC/u0/u0/U66  ( .A1(\AES_ENC/u0/u0/n1024 ), .A2(\AES_ENC/u0/u0/n1071 ), .ZN(\AES_ENC/u0/u0/n1037 ) );
AND2_X2 \AES_ENC/u0/u0/U60  ( .A1(\AES_ENC/u0/u0/n1030 ), .A2(\AES_ENC/u0/u0/n602 ), .ZN(\AES_ENC/u0/u0/n1078 ) );
NAND4_X2 \AES_ENC/u0/u0/U56  ( .A1(\AES_ENC/u0/u0/n1039 ), .A2(\AES_ENC/u0/u0/n1038 ), .A3(\AES_ENC/u0/u0/n1037 ), .A4(\AES_ENC/u0/u0/n1036 ), .ZN(\AES_ENC/u0/u0/n1040 ) );
NAND2_X2 \AES_ENC/u0/u0/U55  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n1040 ), .ZN(\AES_ENC/u0/u0/n1041 ) );
NAND4_X2 \AES_ENC/u0/u0/U54  ( .A1(\AES_ENC/u0/u0/n1044 ), .A2(\AES_ENC/u0/u0/n1043 ), .A3(\AES_ENC/u0/u0/n1042 ), .A4(\AES_ENC/u0/u0/n1041 ), .ZN(\AES_ENC/u0/subword[30] ) );
NAND2_X2 \AES_ENC/u0/u0/U53  ( .A1(\AES_ENC/u0/u0/n1072 ), .A2(\AES_ENC/u0/u0/n1045 ), .ZN(\AES_ENC/u0/u0/n1068 ) );
NAND2_X2 \AES_ENC/u0/u0/U52  ( .A1(\AES_ENC/u0/u0/n1046 ), .A2(\AES_ENC/u0/u0/n582 ), .ZN(\AES_ENC/u0/u0/n1067 ) );
NAND2_X2 \AES_ENC/u0/u0/U51  ( .A1(\AES_ENC/u0/u0/n1094 ), .A2(\AES_ENC/u0/u0/n1047 ), .ZN(\AES_ENC/u0/u0/n1066 ) );
NAND4_X2 \AES_ENC/u0/u0/U40  ( .A1(\AES_ENC/u0/u0/n1068 ), .A2(\AES_ENC/u0/u0/n1067 ), .A3(\AES_ENC/u0/u0/n1066 ), .A4(\AES_ENC/u0/u0/n1065 ), .ZN(\AES_ENC/u0/u0/n1069 ) );
NAND2_X2 \AES_ENC/u0/u0/U39  ( .A1(\AES_ENC/u0/u0/n1070 ), .A2(\AES_ENC/u0/u0/n1069 ), .ZN(\AES_ENC/u0/u0/n1135 ) );
NAND2_X2 \AES_ENC/u0/u0/U38  ( .A1(\AES_ENC/u0/u0/n1072 ), .A2(\AES_ENC/u0/u0/n1071 ), .ZN(\AES_ENC/u0/u0/n1088 ) );
NAND2_X2 \AES_ENC/u0/u0/U37  ( .A1(\AES_ENC/u0/u0/n1073 ), .A2(\AES_ENC/u0/u0/n595 ), .ZN(\AES_ENC/u0/u0/n1087 ) );
NAND4_X2 \AES_ENC/u0/u0/U28  ( .A1(\AES_ENC/u0/u0/n1088 ), .A2(\AES_ENC/u0/u0/n1087 ), .A3(\AES_ENC/u0/u0/n1086 ), .A4(\AES_ENC/u0/u0/n1085 ), .ZN(\AES_ENC/u0/u0/n1089 ) );
NAND2_X2 \AES_ENC/u0/u0/U27  ( .A1(\AES_ENC/u0/u0/n1090 ), .A2(\AES_ENC/u0/u0/n1089 ), .ZN(\AES_ENC/u0/u0/n1134 ) );
NAND2_X2 \AES_ENC/u0/u0/U26  ( .A1(\AES_ENC/u0/u0/n1091 ), .A2(\AES_ENC/u0/u0/n1093 ), .ZN(\AES_ENC/u0/u0/n1111 ) );
NAND2_X2 \AES_ENC/u0/u0/U25  ( .A1(\AES_ENC/u0/u0/n1092 ), .A2(\AES_ENC/u0/u0/n1120 ), .ZN(\AES_ENC/u0/u0/n1110 ) );
AND2_X2 \AES_ENC/u0/u0/U22  ( .A1(\AES_ENC/u0/u0/n1097 ), .A2(\AES_ENC/u0/u0/n1096 ), .ZN(\AES_ENC/u0/u0/n1098 ) );
NAND4_X2 \AES_ENC/u0/u0/U14  ( .A1(\AES_ENC/u0/u0/n1111 ), .A2(\AES_ENC/u0/u0/n1110 ), .A3(\AES_ENC/u0/u0/n1109 ), .A4(\AES_ENC/u0/u0/n1108 ), .ZN(\AES_ENC/u0/u0/n1112 ) );
NAND2_X2 \AES_ENC/u0/u0/U13  ( .A1(\AES_ENC/u0/u0/n1113 ), .A2(\AES_ENC/u0/u0/n1112 ), .ZN(\AES_ENC/u0/u0/n1133 ) );
NAND2_X2 \AES_ENC/u0/u0/U12  ( .A1(\AES_ENC/u0/u0/n1115 ), .A2(\AES_ENC/u0/u0/n1114 ), .ZN(\AES_ENC/u0/u0/n1129 ) );
OR2_X2 \AES_ENC/u0/u0/U11  ( .A1(\AES_ENC/u0/u0/n608 ), .A2(\AES_ENC/u0/u0/n1116 ), .ZN(\AES_ENC/u0/u0/n1128 ) );
NAND4_X2 \AES_ENC/u0/u0/U3  ( .A1(\AES_ENC/u0/u0/n1129 ), .A2(\AES_ENC/u0/u0/n1128 ), .A3(\AES_ENC/u0/u0/n1127 ), .A4(\AES_ENC/u0/u0/n1126 ), .ZN(\AES_ENC/u0/u0/n1130 ) );
NAND2_X2 \AES_ENC/u0/u0/U2  ( .A1(\AES_ENC/u0/u0/n1131 ), .A2(\AES_ENC/u0/u0/n1130 ), .ZN(\AES_ENC/u0/u0/n1132 ) );
NAND4_X2 \AES_ENC/u0/u0/U1  ( .A1(\AES_ENC/u0/u0/n1135 ), .A2(\AES_ENC/u0/u0/n1134 ), .A3(\AES_ENC/u0/u0/n1133 ), .A4(\AES_ENC/u0/u0/n1132 ), .ZN(\AES_ENC/u0/subword[31] ) );
INV_X4 \AES_ENC/u0/u1/U575  ( .A(\AES_ENC/w3[15] ), .ZN(\AES_ENC/u0/u1/n627 ) );
INV_X4 \AES_ENC/u0/u1/U574  ( .A(\AES_ENC/u0/u1/n1114 ), .ZN(\AES_ENC/u0/u1/n625 ) );
INV_X4 \AES_ENC/u0/u1/U573  ( .A(\AES_ENC/w3[12] ), .ZN(\AES_ENC/u0/u1/n624 ) );
INV_X4 \AES_ENC/u0/u1/U572  ( .A(\AES_ENC/u0/u1/n1025 ), .ZN(\AES_ENC/u0/u1/n622 ) );
INV_X4 \AES_ENC/u0/u1/U571  ( .A(\AES_ENC/u0/u1/n1120 ), .ZN(\AES_ENC/u0/u1/n620 ) );
INV_X4 \AES_ENC/u0/u1/U570  ( .A(\AES_ENC/u0/u1/n1121 ), .ZN(\AES_ENC/u0/u1/n619 ) );
INV_X4 \AES_ENC/u0/u1/U569  ( .A(\AES_ENC/u0/u1/n1048 ), .ZN(\AES_ENC/u0/u1/n618 ) );
INV_X4 \AES_ENC/u0/u1/U568  ( .A(\AES_ENC/u0/u1/n974 ), .ZN(\AES_ENC/u0/u1/n616 ) );
INV_X4 \AES_ENC/u0/u1/U567  ( .A(\AES_ENC/u0/u1/n794 ), .ZN(\AES_ENC/u0/u1/n614 ) );
INV_X4 \AES_ENC/u0/u1/U566  ( .A(\AES_ENC/w3[10] ), .ZN(\AES_ENC/u0/u1/n611 ) );
INV_X4 \AES_ENC/u0/u1/U565  ( .A(\AES_ENC/u0/u1/n800 ), .ZN(\AES_ENC/u0/u1/n610 ) );
INV_X4 \AES_ENC/u0/u1/U564  ( .A(\AES_ENC/u0/u1/n925 ), .ZN(\AES_ENC/u0/u1/n609 ) );
INV_X4 \AES_ENC/u0/u1/U563  ( .A(\AES_ENC/u0/u1/n779 ), .ZN(\AES_ENC/u0/u1/n607 ) );
INV_X4 \AES_ENC/u0/u1/U562  ( .A(\AES_ENC/u0/u1/n1022 ), .ZN(\AES_ENC/u0/u1/n603 ) );
INV_X4 \AES_ENC/u0/u1/U561  ( .A(\AES_ENC/u0/u1/n1102 ), .ZN(\AES_ENC/u0/u1/n602 ) );
INV_X4 \AES_ENC/u0/u1/U560  ( .A(\AES_ENC/u0/u1/n929 ), .ZN(\AES_ENC/u0/u1/n601 ) );
INV_X4 \AES_ENC/u0/u1/U559  ( .A(\AES_ENC/u0/u1/n1056 ), .ZN(\AES_ENC/u0/u1/n600 ) );
INV_X4 \AES_ENC/u0/u1/U558  ( .A(\AES_ENC/u0/u1/n1054 ), .ZN(\AES_ENC/u0/u1/n599 ) );
INV_X4 \AES_ENC/u0/u1/U557  ( .A(\AES_ENC/u0/u1/n881 ), .ZN(\AES_ENC/u0/u1/n598 ) );
INV_X4 \AES_ENC/u0/u1/U556  ( .A(\AES_ENC/u0/u1/n926 ), .ZN(\AES_ENC/u0/u1/n597 ) );
INV_X4 \AES_ENC/u0/u1/U555  ( .A(\AES_ENC/u0/u1/n977 ), .ZN(\AES_ENC/u0/u1/n595 ) );
INV_X4 \AES_ENC/u0/u1/U554  ( .A(\AES_ENC/u0/u1/n1031 ), .ZN(\AES_ENC/u0/u1/n594 ) );
INV_X4 \AES_ENC/u0/u1/U553  ( .A(\AES_ENC/u0/u1/n1103 ), .ZN(\AES_ENC/u0/u1/n593 ) );
INV_X4 \AES_ENC/u0/u1/U552  ( .A(\AES_ENC/u0/u1/n1009 ), .ZN(\AES_ENC/u0/u1/n592 ) );
INV_X4 \AES_ENC/u0/u1/U551  ( .A(\AES_ENC/u0/u1/n990 ), .ZN(\AES_ENC/u0/u1/n591 ) );
INV_X4 \AES_ENC/u0/u1/U550  ( .A(\AES_ENC/u0/u1/n1058 ), .ZN(\AES_ENC/u0/u1/n590 ) );
INV_X4 \AES_ENC/u0/u1/U549  ( .A(\AES_ENC/u0/u1/n1074 ), .ZN(\AES_ENC/u0/u1/n589 ) );
INV_X4 \AES_ENC/u0/u1/U548  ( .A(\AES_ENC/u0/u1/n1053 ), .ZN(\AES_ENC/u0/u1/n588 ) );
INV_X4 \AES_ENC/u0/u1/U547  ( .A(\AES_ENC/u0/u1/n826 ), .ZN(\AES_ENC/u0/u1/n587 ) );
INV_X4 \AES_ENC/u0/u1/U546  ( .A(\AES_ENC/u0/u1/n992 ), .ZN(\AES_ENC/u0/u1/n586 ) );
INV_X4 \AES_ENC/u0/u1/U545  ( .A(\AES_ENC/u0/u1/n821 ), .ZN(\AES_ENC/u0/u1/n585 ) );
INV_X4 \AES_ENC/u0/u1/U544  ( .A(\AES_ENC/u0/u1/n910 ), .ZN(\AES_ENC/u0/u1/n584 ) );
INV_X4 \AES_ENC/u0/u1/U543  ( .A(\AES_ENC/u0/u1/n906 ), .ZN(\AES_ENC/u0/u1/n583 ) );
INV_X4 \AES_ENC/u0/u1/U542  ( .A(\AES_ENC/u0/u1/n880 ), .ZN(\AES_ENC/u0/u1/n581 ) );
INV_X4 \AES_ENC/u0/u1/U541  ( .A(\AES_ENC/u0/u1/n1013 ), .ZN(\AES_ENC/u0/u1/n580 ) );
INV_X4 \AES_ENC/u0/u1/U540  ( .A(\AES_ENC/u0/u1/n1092 ), .ZN(\AES_ENC/u0/u1/n579 ) );
INV_X4 \AES_ENC/u0/u1/U539  ( .A(\AES_ENC/u0/u1/n824 ), .ZN(\AES_ENC/u0/u1/n578 ) );
INV_X4 \AES_ENC/u0/u1/U538  ( .A(\AES_ENC/u0/u1/n1091 ), .ZN(\AES_ENC/u0/u1/n577 ) );
INV_X4 \AES_ENC/u0/u1/U537  ( .A(\AES_ENC/u0/u1/n1080 ), .ZN(\AES_ENC/u0/u1/n576 ) );
INV_X4 \AES_ENC/u0/u1/U536  ( .A(\AES_ENC/u0/u1/n959 ), .ZN(\AES_ENC/u0/u1/n575 ) );
INV_X4 \AES_ENC/u0/u1/U535  ( .A(\AES_ENC/w3[8] ), .ZN(\AES_ENC/u0/u1/n574 ));
NOR2_X2 \AES_ENC/u0/u1/U534  ( .A1(\AES_ENC/u0/u1/n574 ), .A2(\AES_ENC/w3[14] ), .ZN(\AES_ENC/u0/u1/n1070 ) );
NOR2_X2 \AES_ENC/u0/u1/U533  ( .A1(\AES_ENC/w3[8] ), .A2(\AES_ENC/w3[14] ),.ZN(\AES_ENC/u0/u1/n1090 ) );
NOR2_X2 \AES_ENC/u0/u1/U532  ( .A1(\AES_ENC/w3[12] ), .A2(\AES_ENC/w3[11] ),.ZN(\AES_ENC/u0/u1/n1025 ) );
NAND3_X2 \AES_ENC/u0/u1/U531  ( .A1(\AES_ENC/u0/u1/n679 ), .A2(\AES_ENC/u0/u1/n678 ), .A3(\AES_ENC/u0/u1/n677 ), .ZN(\AES_ENC/u0/subword[16] ) );
NOR2_X2 \AES_ENC/u0/u1/U530  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n765 ) );
NOR2_X2 \AES_ENC/u0/u1/U529  ( .A1(\AES_ENC/w3[12] ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n764 ) );
NOR2_X2 \AES_ENC/u0/u1/U528  ( .A1(\AES_ENC/u0/u1/n765 ), .A2(\AES_ENC/u0/u1/n764 ), .ZN(\AES_ENC/u0/u1/n766 ) );
NOR2_X2 \AES_ENC/u0/u1/U527  ( .A1(\AES_ENC/u0/u1/n766 ), .A2(\AES_ENC/u0/u1/n575 ), .ZN(\AES_ENC/u0/u1/n767 ) );
NOR2_X2 \AES_ENC/u0/u1/U526  ( .A1(\AES_ENC/u0/u1/n1117 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n707 ) );
NOR3_X2 \AES_ENC/u0/u1/U525  ( .A1(\AES_ENC/u0/u1/n627 ), .A2(\AES_ENC/w3[13] ), .A3(\AES_ENC/u0/u1/n704 ), .ZN(\AES_ENC/u0/u1/n706 ) );
NOR2_X2 \AES_ENC/u0/u1/U524  ( .A1(\AES_ENC/w3[12] ), .A2(\AES_ENC/u0/u1/n579 ), .ZN(\AES_ENC/u0/u1/n705 ) );
NOR3_X2 \AES_ENC/u0/u1/U523  ( .A1(\AES_ENC/u0/u1/n707 ), .A2(\AES_ENC/u0/u1/n706 ), .A3(\AES_ENC/u0/u1/n705 ), .ZN(\AES_ENC/u0/u1/n713 ) );
NOR4_X2 \AES_ENC/u0/u1/U522  ( .A1(\AES_ENC/u0/u1/n633 ), .A2(\AES_ENC/u0/u1/n632 ), .A3(\AES_ENC/u0/u1/n631 ), .A4(\AES_ENC/u0/u1/n630 ), .ZN(\AES_ENC/u0/u1/n634 ) );
NOR2_X2 \AES_ENC/u0/u1/U521  ( .A1(\AES_ENC/u0/u1/n629 ), .A2(\AES_ENC/u0/u1/n628 ), .ZN(\AES_ENC/u0/u1/n635 ) );
NAND3_X2 \AES_ENC/u0/u1/U520  ( .A1(\AES_ENC/w3[10] ), .A2(\AES_ENC/w3[15] ),.A3(\AES_ENC/u0/u1/n1059 ), .ZN(\AES_ENC/u0/u1/n636 ) );
INV_X4 \AES_ENC/u0/u1/U519  ( .A(\AES_ENC/w3[11] ), .ZN(\AES_ENC/u0/u1/n621 ) );
NOR2_X2 \AES_ENC/u0/u1/U518  ( .A1(\AES_ENC/w3[13] ), .A2(\AES_ENC/w3[10] ),.ZN(\AES_ENC/u0/u1/n974 ) );
NAND3_X2 \AES_ENC/u0/u1/U517  ( .A1(\AES_ENC/u0/u1/n652 ), .A2(\AES_ENC/u0/u1/n626 ), .A3(\AES_ENC/w3[15] ), .ZN(\AES_ENC/u0/u1/n653 ) );
NOR2_X2 \AES_ENC/u0/u1/U516  ( .A1(\AES_ENC/u0/u1/n611 ), .A2(\AES_ENC/w3[13] ), .ZN(\AES_ENC/u0/u1/n925 ) );
NOR2_X2 \AES_ENC/u0/u1/U515  ( .A1(\AES_ENC/u0/u1/n626 ), .A2(\AES_ENC/w3[10] ), .ZN(\AES_ENC/u0/u1/n1048 ) );
INV_X4 \AES_ENC/u0/u1/U512  ( .A(\AES_ENC/w3[13] ), .ZN(\AES_ENC/u0/u1/n626 ) );
NOR2_X2 \AES_ENC/u0/u1/U510  ( .A1(\AES_ENC/u0/u1/n611 ), .A2(\AES_ENC/w3[15] ), .ZN(\AES_ENC/u0/u1/n779 ) );
NOR2_X2 \AES_ENC/u0/u1/U509  ( .A1(\AES_ENC/w3[15] ), .A2(\AES_ENC/w3[10] ),.ZN(\AES_ENC/u0/u1/n794 ) );
NOR2_X2 \AES_ENC/u0/u1/U508  ( .A1(\AES_ENC/w3[12] ), .A2(\AES_ENC/w3[9] ),.ZN(\AES_ENC/u0/u1/n1102 ) );
INV_X4 \AES_ENC/u0/u1/U507  ( .A(\AES_ENC/u0/u1/n569 ), .ZN(\AES_ENC/u0/u1/n572 ) );
NOR2_X2 \AES_ENC/u0/u1/U506  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/w3[11] ), .ZN(\AES_ENC/u0/u1/n1053 ) );
NOR2_X2 \AES_ENC/u0/u1/U505  ( .A1(\AES_ENC/u0/u1/n607 ), .A2(\AES_ENC/w3[13] ), .ZN(\AES_ENC/u0/u1/n1024 ) );
NOR2_X2 \AES_ENC/u0/u1/U504  ( .A1(\AES_ENC/u0/u1/n625 ), .A2(\AES_ENC/w3[10] ), .ZN(\AES_ENC/u0/u1/n1093 ) );
NOR2_X2 \AES_ENC/u0/u1/U503  ( .A1(\AES_ENC/u0/u1/n614 ), .A2(\AES_ENC/w3[13] ), .ZN(\AES_ENC/u0/u1/n1094 ) );
NOR2_X2 \AES_ENC/u0/u1/U502  ( .A1(\AES_ENC/u0/u1/n624 ), .A2(\AES_ENC/w3[11] ), .ZN(\AES_ENC/u0/u1/n931 ) );
INV_X4 \AES_ENC/u0/u1/U501  ( .A(\AES_ENC/u0/u1/n570 ), .ZN(\AES_ENC/u0/u1/n573 ) );
NOR2_X2 \AES_ENC/u0/u1/U500  ( .A1(\AES_ENC/u0/u1/n622 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n1059 ) );
NOR2_X2 \AES_ENC/u0/u1/U499  ( .A1(\AES_ENC/u0/u1/n1053 ), .A2(\AES_ENC/u0/u1/n1095 ), .ZN(\AES_ENC/u0/u1/n639 ) );
NOR3_X2 \AES_ENC/u0/u1/U498  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n573 ), .A3(\AES_ENC/u0/u1/n1074 ), .ZN(\AES_ENC/u0/u1/n641 ) );
NOR2_X2 \AES_ENC/u0/u1/U497  ( .A1(\AES_ENC/u0/u1/n639 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n640 ) );
NOR2_X2 \AES_ENC/u0/u1/U496  ( .A1(\AES_ENC/u0/u1/n641 ), .A2(\AES_ENC/u0/u1/n640 ), .ZN(\AES_ENC/u0/u1/n646 ) );
NOR2_X2 \AES_ENC/u0/u1/U495  ( .A1(\AES_ENC/u0/u1/n826 ), .A2(\AES_ENC/u0/u1/n572 ), .ZN(\AES_ENC/u0/u1/n827 ) );
NOR3_X2 \AES_ENC/u0/u1/U494  ( .A1(\AES_ENC/u0/u1/n769 ), .A2(\AES_ENC/u0/u1/n768 ), .A3(\AES_ENC/u0/u1/n767 ), .ZN(\AES_ENC/u0/u1/n775 ) );
NOR2_X2 \AES_ENC/u0/u1/U492  ( .A1(\AES_ENC/w3[9] ), .A2(\AES_ENC/u0/u1/n623 ), .ZN(\AES_ENC/u0/u1/n913 ) );
NOR2_X2 \AES_ENC/u0/u1/U491  ( .A1(\AES_ENC/u0/u1/n913 ), .A2(\AES_ENC/u0/u1/n1091 ), .ZN(\AES_ENC/u0/u1/n914 ) );
NOR2_X2 \AES_ENC/u0/u1/U490  ( .A1(\AES_ENC/u0/u1/n1056 ), .A2(\AES_ENC/u0/u1/n1053 ), .ZN(\AES_ENC/u0/u1/n749 ) );
NOR2_X2 \AES_ENC/u0/u1/U489  ( .A1(\AES_ENC/u0/u1/n749 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n752 ) );
NOR3_X2 \AES_ENC/u0/u1/U488  ( .A1(\AES_ENC/u0/u1/n995 ), .A2(\AES_ENC/u0/u1/n586 ), .A3(\AES_ENC/u0/u1/n994 ), .ZN(\AES_ENC/u0/u1/n1002 ) );
NOR2_X2 \AES_ENC/u0/u1/U487  ( .A1(\AES_ENC/u0/u1/n909 ), .A2(\AES_ENC/u0/u1/n908 ), .ZN(\AES_ENC/u0/u1/n920 ) );
INV_X4 \AES_ENC/u0/u1/U486  ( .A(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n596 ));
NOR2_X2 \AES_ENC/u0/u1/U483  ( .A1(\AES_ENC/u0/u1/n932 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n933 ) );
NOR2_X2 \AES_ENC/u0/u1/U482  ( .A1(\AES_ENC/u0/u1/n929 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n935 ) );
NOR2_X2 \AES_ENC/u0/u1/U480  ( .A1(\AES_ENC/u0/u1/n931 ), .A2(\AES_ENC/u0/u1/n930 ), .ZN(\AES_ENC/u0/u1/n934 ) );
NOR3_X2 \AES_ENC/u0/u1/U479  ( .A1(\AES_ENC/u0/u1/n935 ), .A2(\AES_ENC/u0/u1/n934 ), .A3(\AES_ENC/u0/u1/n933 ), .ZN(\AES_ENC/u0/u1/n936 ) );
OR2_X4 \AES_ENC/u0/u1/U478  ( .A1(\AES_ENC/u0/u1/n1094 ), .A2(\AES_ENC/u0/u1/n1093 ), .ZN(\AES_ENC/u0/u1/n571 ) );
AND2_X2 \AES_ENC/u0/u1/U477  ( .A1(\AES_ENC/u0/u1/n571 ), .A2(\AES_ENC/u0/u1/n1095 ), .ZN(\AES_ENC/u0/u1/n1101 ) );
NOR2_X2 \AES_ENC/u0/u1/U474  ( .A1(\AES_ENC/u0/u1/n1074 ), .A2(\AES_ENC/u0/u1/n931 ), .ZN(\AES_ENC/u0/u1/n796 ) );
NOR2_X2 \AES_ENC/u0/u1/U473  ( .A1(\AES_ENC/u0/u1/n796 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n797 ) );
NOR2_X2 \AES_ENC/u0/u1/U472  ( .A1(\AES_ENC/u0/u1/n1054 ), .A2(\AES_ENC/u0/u1/n1053 ), .ZN(\AES_ENC/u0/u1/n1055 ) );
NOR2_X2 \AES_ENC/u0/u1/U471  ( .A1(\AES_ENC/u0/u1/n572 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n949 ) );
NOR2_X2 \AES_ENC/u0/u1/U470  ( .A1(\AES_ENC/u0/u1/n1049 ), .A2(\AES_ENC/u0/u1/n618 ), .ZN(\AES_ENC/u0/u1/n1051 ) );
NOR2_X2 \AES_ENC/u0/u1/U469  ( .A1(\AES_ENC/u0/u1/n1051 ), .A2(\AES_ENC/u0/u1/n1050 ), .ZN(\AES_ENC/u0/u1/n1052 ) );
NOR2_X2 \AES_ENC/u0/u1/U468  ( .A1(\AES_ENC/u0/u1/n1052 ), .A2(\AES_ENC/u0/u1/n592 ), .ZN(\AES_ENC/u0/u1/n1064 ) );
NOR2_X2 \AES_ENC/u0/u1/U467  ( .A1(\AES_ENC/w3[9] ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n631 ) );
NOR2_X2 \AES_ENC/u0/u1/U466  ( .A1(\AES_ENC/u0/u1/n1025 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n980 ) );
NOR2_X2 \AES_ENC/u0/u1/U465  ( .A1(\AES_ENC/u0/u1/n1074 ), .A2(\AES_ENC/u0/u1/n1025 ), .ZN(\AES_ENC/u0/u1/n891 ) );
NOR2_X2 \AES_ENC/u0/u1/U464  ( .A1(\AES_ENC/u0/u1/n891 ), .A2(\AES_ENC/u0/u1/n609 ), .ZN(\AES_ENC/u0/u1/n894 ) );
NOR2_X2 \AES_ENC/u0/u1/U463  ( .A1(\AES_ENC/u0/u1/n1073 ), .A2(\AES_ENC/u0/u1/n1094 ), .ZN(\AES_ENC/u0/u1/n795 ) );
NOR2_X2 \AES_ENC/u0/u1/U462  ( .A1(\AES_ENC/u0/u1/n795 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n799 ) );
NOR2_X2 \AES_ENC/u0/u1/U461  ( .A1(\AES_ENC/u0/u1/n624 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n1075 ) );
NOR2_X2 \AES_ENC/u0/u1/U460  ( .A1(\AES_ENC/u0/u1/n624 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n822 ) );
NOR2_X2 \AES_ENC/u0/u1/U459  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n823 ) );
NOR2_X2 \AES_ENC/u0/u1/U458  ( .A1(\AES_ENC/u0/u1/n823 ), .A2(\AES_ENC/u0/u1/n822 ), .ZN(\AES_ENC/u0/u1/n825 ) );
NOR2_X2 \AES_ENC/u0/u1/U455  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n981 ) );
NOR2_X2 \AES_ENC/u0/u1/U448  ( .A1(\AES_ENC/u0/u1/n1102 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n643 ) );
NOR2_X2 \AES_ENC/u0/u1/U447  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n621 ), .ZN(\AES_ENC/u0/u1/n642 ) );
NOR2_X2 \AES_ENC/u0/u1/U442  ( .A1(\AES_ENC/u0/u1/n911 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n644 ) );
NOR4_X2 \AES_ENC/u0/u1/U441  ( .A1(\AES_ENC/u0/u1/n644 ), .A2(\AES_ENC/u0/u1/n643 ), .A3(\AES_ENC/u0/u1/n804 ), .A4(\AES_ENC/u0/u1/n642 ), .ZN(\AES_ENC/u0/u1/n645 ) );
NOR2_X2 \AES_ENC/u0/u1/U438  ( .A1(\AES_ENC/u0/u1/n1102 ), .A2(\AES_ENC/u0/u1/n910 ), .ZN(\AES_ENC/u0/u1/n932 ) );
NOR3_X2 \AES_ENC/u0/u1/U435  ( .A1(\AES_ENC/u0/u1/n623 ), .A2(\AES_ENC/w3[9] ), .A3(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n683 ));
NOR2_X2 \AES_ENC/u0/u1/U434  ( .A1(\AES_ENC/u0/u1/n1102 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n755 ) );
INV_X4 \AES_ENC/u0/u1/U433  ( .A(\AES_ENC/u0/u1/n931 ), .ZN(\AES_ENC/u0/u1/n623 ) );
NOR2_X2 \AES_ENC/u0/u1/U428  ( .A1(\AES_ENC/u0/u1/n996 ), .A2(\AES_ENC/u0/u1/n931 ), .ZN(\AES_ENC/u0/u1/n704 ) );
NOR2_X2 \AES_ENC/u0/u1/U427  ( .A1(\AES_ENC/u0/u1/n1029 ), .A2(\AES_ENC/u0/u1/n1025 ), .ZN(\AES_ENC/u0/u1/n1079 ) );
NOR3_X2 \AES_ENC/u0/u1/U421  ( .A1(\AES_ENC/u0/u1/n589 ), .A2(\AES_ENC/u0/u1/n1025 ), .A3(\AES_ENC/u0/u1/n616 ), .ZN(\AES_ENC/u0/u1/n945 ) );
NOR2_X2 \AES_ENC/u0/u1/U420  ( .A1(\AES_ENC/u0/u1/n1072 ), .A2(\AES_ENC/u0/u1/n1094 ), .ZN(\AES_ENC/u0/u1/n930 ) );
NOR2_X2 \AES_ENC/u0/u1/U419  ( .A1(\AES_ENC/u0/u1/n931 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n743 ) );
NOR2_X2 \AES_ENC/u0/u1/U418  ( .A1(\AES_ENC/u0/u1/n931 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n685 ) );
NOR3_X2 \AES_ENC/u0/u1/U417  ( .A1(\AES_ENC/u0/u1/n610 ), .A2(\AES_ENC/u0/u1/n572 ), .A3(\AES_ENC/u0/u1/n575 ), .ZN(\AES_ENC/u0/u1/n962 ) );
NOR2_X2 \AES_ENC/u0/u1/U416  ( .A1(\AES_ENC/u0/u1/n626 ), .A2(\AES_ENC/u0/u1/n611 ), .ZN(\AES_ENC/u0/u1/n800 ) );
NOR3_X2 \AES_ENC/u0/u1/U415  ( .A1(\AES_ENC/u0/u1/n590 ), .A2(\AES_ENC/u0/u1/n627 ), .A3(\AES_ENC/u0/u1/n611 ), .ZN(\AES_ENC/u0/u1/n798 ) );
NOR3_X2 \AES_ENC/u0/u1/U414  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n572 ), .A3(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n694 ) );
NOR3_X2 \AES_ENC/u0/u1/U413  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n572 ), .A3(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n895 ) );
NOR3_X2 \AES_ENC/u0/u1/U410  ( .A1(\AES_ENC/u0/u1/n1008 ), .A2(\AES_ENC/u0/u1/n1007 ), .A3(\AES_ENC/u0/u1/n1006 ), .ZN(\AES_ENC/u0/u1/n1018 ) );
NOR2_X2 \AES_ENC/u0/u1/U409  ( .A1(\AES_ENC/u0/u1/n669 ), .A2(\AES_ENC/u0/u1/n668 ), .ZN(\AES_ENC/u0/u1/n673 ) );
NOR4_X2 \AES_ENC/u0/u1/U406  ( .A1(\AES_ENC/u0/u1/n946 ), .A2(\AES_ENC/u0/u1/n1046 ), .A3(\AES_ENC/u0/u1/n671 ), .A4(\AES_ENC/u0/u1/n670 ), .ZN(\AES_ENC/u0/u1/n672 ) );
NOR4_X2 \AES_ENC/u0/u1/U405  ( .A1(\AES_ENC/u0/u1/n711 ), .A2(\AES_ENC/u0/u1/n710 ), .A3(\AES_ENC/u0/u1/n709 ), .A4(\AES_ENC/u0/u1/n708 ), .ZN(\AES_ENC/u0/u1/n712 ) );
NOR4_X2 \AES_ENC/u0/u1/U404  ( .A1(\AES_ENC/u0/u1/n806 ), .A2(\AES_ENC/u0/u1/n805 ), .A3(\AES_ENC/u0/u1/n804 ), .A4(\AES_ENC/u0/u1/n803 ), .ZN(\AES_ENC/u0/u1/n807 ) );
NOR3_X2 \AES_ENC/u0/u1/U403  ( .A1(\AES_ENC/u0/u1/n799 ), .A2(\AES_ENC/u0/u1/n798 ), .A3(\AES_ENC/u0/u1/n797 ), .ZN(\AES_ENC/u0/u1/n808 ) );
NOR4_X2 \AES_ENC/u0/u1/U401  ( .A1(\AES_ENC/u0/u1/n843 ), .A2(\AES_ENC/u0/u1/n842 ), .A3(\AES_ENC/u0/u1/n841 ), .A4(\AES_ENC/u0/u1/n840 ), .ZN(\AES_ENC/u0/u1/n844 ) );
NOR3_X2 \AES_ENC/u0/u1/U400  ( .A1(\AES_ENC/u0/u1/n1101 ), .A2(\AES_ENC/u0/u1/n1100 ), .A3(\AES_ENC/u0/u1/n1099 ), .ZN(\AES_ENC/u0/u1/n1109 ) );
NOR3_X2 \AES_ENC/u0/u1/U399  ( .A1(\AES_ENC/u0/u1/n743 ), .A2(\AES_ENC/u0/u1/n742 ), .A3(\AES_ENC/u0/u1/n741 ), .ZN(\AES_ENC/u0/u1/n744 ) );
NOR2_X2 \AES_ENC/u0/u1/U398  ( .A1(\AES_ENC/u0/u1/n697 ), .A2(\AES_ENC/u0/u1/n658 ), .ZN(\AES_ENC/u0/u1/n659 ) );
NOR3_X2 \AES_ENC/u0/u1/U397  ( .A1(\AES_ENC/u0/u1/n959 ), .A2(\AES_ENC/u0/u1/n572 ), .A3(\AES_ENC/u0/u1/n609 ), .ZN(\AES_ENC/u0/u1/n768 ) );
NOR2_X2 \AES_ENC/u0/u1/U396  ( .A1(\AES_ENC/u0/u1/n598 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n885 ) );
NOR2_X2 \AES_ENC/u0/u1/U393  ( .A1(\AES_ENC/u0/u1/n623 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n882 ) );
NOR2_X2 \AES_ENC/u0/u1/U390  ( .A1(\AES_ENC/u0/u1/n1053 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n884 ) );
NOR4_X2 \AES_ENC/u0/u1/U389  ( .A1(\AES_ENC/u0/u1/n885 ), .A2(\AES_ENC/u0/u1/n884 ), .A3(\AES_ENC/u0/u1/n883 ), .A4(\AES_ENC/u0/u1/n882 ), .ZN(\AES_ENC/u0/u1/n886 ) );
NOR2_X2 \AES_ENC/u0/u1/U388  ( .A1(\AES_ENC/u0/u1/n1078 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n1033 ) );
NOR2_X2 \AES_ENC/u0/u1/U387  ( .A1(\AES_ENC/u0/u1/n1031 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n1032 ) );
NOR3_X2 \AES_ENC/u0/u1/U386  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n1025 ), .A3(\AES_ENC/u0/u1/n1074 ), .ZN(\AES_ENC/u0/u1/n1035 ) );
NOR4_X2 \AES_ENC/u0/u1/U385  ( .A1(\AES_ENC/u0/u1/n1035 ), .A2(\AES_ENC/u0/u1/n1034 ), .A3(\AES_ENC/u0/u1/n1033 ), .A4(\AES_ENC/u0/u1/n1032 ), .ZN(\AES_ENC/u0/u1/n1036 ) );
NOR2_X2 \AES_ENC/u0/u1/U384  ( .A1(\AES_ENC/u0/u1/n825 ), .A2(\AES_ENC/u0/u1/n578 ), .ZN(\AES_ENC/u0/u1/n830 ) );
NOR2_X2 \AES_ENC/u0/u1/U383  ( .A1(\AES_ENC/u0/u1/n827 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n829 ) );
NOR2_X2 \AES_ENC/u0/u1/U382  ( .A1(\AES_ENC/u0/u1/n572 ), .A2(\AES_ENC/u0/u1/n579 ), .ZN(\AES_ENC/u0/u1/n828 ) );
NOR4_X2 \AES_ENC/u0/u1/U374  ( .A1(\AES_ENC/u0/u1/n831 ), .A2(\AES_ENC/u0/u1/n830 ), .A3(\AES_ENC/u0/u1/n829 ), .A4(\AES_ENC/u0/u1/n828 ), .ZN(\AES_ENC/u0/u1/n832 ) );
NOR2_X2 \AES_ENC/u0/u1/U373  ( .A1(\AES_ENC/u0/u1/n598 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n1107 ) );
NOR2_X2 \AES_ENC/u0/u1/U372  ( .A1(\AES_ENC/u0/u1/n1102 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n1106 ) );
NOR2_X2 \AES_ENC/u0/u1/U370  ( .A1(\AES_ENC/u0/u1/n1103 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n1105 ) );
NOR4_X2 \AES_ENC/u0/u1/U369  ( .A1(\AES_ENC/u0/u1/n1107 ), .A2(\AES_ENC/u0/u1/n1106 ), .A3(\AES_ENC/u0/u1/n1105 ), .A4(\AES_ENC/u0/u1/n1104 ), .ZN(\AES_ENC/u0/u1/n1108 ) );
NOR3_X2 \AES_ENC/u0/u1/U368  ( .A1(\AES_ENC/u0/u1/n959 ), .A2(\AES_ENC/u0/u1/n621 ), .A3(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n963 ) );
NOR2_X2 \AES_ENC/u0/u1/U367  ( .A1(\AES_ENC/u0/u1/n626 ), .A2(\AES_ENC/u0/u1/n627 ), .ZN(\AES_ENC/u0/u1/n1114 ) );
NOR3_X2 \AES_ENC/u0/u1/U366  ( .A1(\AES_ENC/u0/u1/n910 ), .A2(\AES_ENC/u0/u1/n1059 ), .A3(\AES_ENC/u0/u1/n611 ), .ZN(\AES_ENC/u0/u1/n1115 ) );
INV_X4 \AES_ENC/u0/u1/U365  ( .A(\AES_ENC/u0/u1/n1024 ), .ZN(\AES_ENC/u0/u1/n606 ) );
INV_X4 \AES_ENC/u0/u1/U364  ( .A(\AES_ENC/u0/u1/n1094 ), .ZN(\AES_ENC/u0/u1/n613 ) );
NOR2_X2 \AES_ENC/u0/u1/U363  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n931 ), .ZN(\AES_ENC/u0/u1/n1100 ) );
NOR2_X2 \AES_ENC/u0/u1/U354  ( .A1(\AES_ENC/u0/u1/n569 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n929 ) );
NOR2_X2 \AES_ENC/u0/u1/U353  ( .A1(\AES_ENC/u0/u1/n620 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n926 ) );
INV_X4 \AES_ENC/u0/u1/U352  ( .A(\AES_ENC/u0/u1/n1093 ), .ZN(\AES_ENC/u0/u1/n617 ) );
NOR2_X2 \AES_ENC/u0/u1/U351  ( .A1(\AES_ENC/u0/u1/n572 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n1095 ) );
NOR2_X2 \AES_ENC/u0/u1/U350  ( .A1(\AES_ENC/u0/u1/n609 ), .A2(\AES_ENC/u0/u1/n627 ), .ZN(\AES_ENC/u0/u1/n1010 ) );
NOR2_X2 \AES_ENC/u0/u1/U349  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n1103 ) );
NOR2_X2 \AES_ENC/u0/u1/U348  ( .A1(\AES_ENC/w3[9] ), .A2(\AES_ENC/u0/u1/n1120 ), .ZN(\AES_ENC/u0/u1/n1022 ) );
NOR2_X2 \AES_ENC/u0/u1/U347  ( .A1(\AES_ENC/u0/u1/n619 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n911 ) );
NOR2_X2 \AES_ENC/u0/u1/U346  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/u0/u1/n1025 ), .ZN(\AES_ENC/u0/u1/n826 ) );
NOR2_X2 \AES_ENC/u0/u1/U345  ( .A1(\AES_ENC/u0/u1/n626 ), .A2(\AES_ENC/u0/u1/n607 ), .ZN(\AES_ENC/u0/u1/n1072 ) );
NOR2_X2 \AES_ENC/u0/u1/U338  ( .A1(\AES_ENC/u0/u1/n627 ), .A2(\AES_ENC/u0/u1/n616 ), .ZN(\AES_ENC/u0/u1/n956 ) );
NOR2_X2 \AES_ENC/u0/u1/U335  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/u0/u1/n624 ), .ZN(\AES_ENC/u0/u1/n1121 ) );
NOR2_X2 \AES_ENC/u0/u1/U329  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/u0/u1/n624 ), .ZN(\AES_ENC/u0/u1/n1058 ) );
NOR2_X2 \AES_ENC/u0/u1/U328  ( .A1(\AES_ENC/u0/u1/n625 ), .A2(\AES_ENC/u0/u1/n611 ), .ZN(\AES_ENC/u0/u1/n1073 ) );
NOR2_X2 \AES_ENC/u0/u1/U327  ( .A1(\AES_ENC/w3[9] ), .A2(\AES_ENC/u0/u1/n1025 ), .ZN(\AES_ENC/u0/u1/n1054 ) );
NOR2_X2 \AES_ENC/u0/u1/U325  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/u0/u1/n931 ), .ZN(\AES_ENC/u0/u1/n1029 ) );
NOR2_X2 \AES_ENC/u0/u1/U324  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n1056 ) );
NOR2_X2 \AES_ENC/u0/u1/U319  ( .A1(\AES_ENC/u0/u1/n614 ), .A2(\AES_ENC/u0/u1/n626 ), .ZN(\AES_ENC/u0/u1/n1050 ) );
NOR2_X2 \AES_ENC/u0/u1/U318  ( .A1(\AES_ENC/u0/u1/n1121 ), .A2(\AES_ENC/u0/u1/n1025 ), .ZN(\AES_ENC/u0/u1/n1120 ) );
NOR2_X2 \AES_ENC/u0/u1/U317  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/u0/u1/n572 ), .ZN(\AES_ENC/u0/u1/n1074 ) );
NOR2_X2 \AES_ENC/u0/u1/U316  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n584 ), .ZN(\AES_ENC/u0/u1/n838 ) );
NOR2_X2 \AES_ENC/u0/u1/U315  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n602 ), .ZN(\AES_ENC/u0/u1/n837 ) );
NOR2_X2 \AES_ENC/u0/u1/U314  ( .A1(\AES_ENC/u0/u1/n838 ), .A2(\AES_ENC/u0/u1/n837 ), .ZN(\AES_ENC/u0/u1/n845 ) );
NOR2_X2 \AES_ENC/u0/u1/U312  ( .A1(\AES_ENC/u0/u1/n1058 ), .A2(\AES_ENC/u0/u1/n1054 ), .ZN(\AES_ENC/u0/u1/n878 ) );
NOR2_X2 \AES_ENC/u0/u1/U311  ( .A1(\AES_ENC/u0/u1/n878 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n879 ) );
NOR2_X2 \AES_ENC/u0/u1/U310  ( .A1(\AES_ENC/u0/u1/n880 ), .A2(\AES_ENC/u0/u1/n879 ), .ZN(\AES_ENC/u0/u1/n887 ) );
NOR3_X2 \AES_ENC/u0/u1/U309  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n1091 ), .A3(\AES_ENC/u0/u1/n1022 ), .ZN(\AES_ENC/u0/u1/n720 ) );
NOR3_X2 \AES_ENC/u0/u1/U303  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n1054 ), .A3(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n719 ) );
NOR2_X2 \AES_ENC/u0/u1/U302  ( .A1(\AES_ENC/u0/u1/n720 ), .A2(\AES_ENC/u0/u1/n719 ), .ZN(\AES_ENC/u0/u1/n726 ) );
NOR2_X2 \AES_ENC/u0/u1/U300  ( .A1(\AES_ENC/u0/u1/n614 ), .A2(\AES_ENC/u0/u1/n591 ), .ZN(\AES_ENC/u0/u1/n865 ) );
NOR2_X2 \AES_ENC/u0/u1/U299  ( .A1(\AES_ENC/u0/u1/n1059 ), .A2(\AES_ENC/u0/u1/n1058 ), .ZN(\AES_ENC/u0/u1/n1060 ) );
NOR2_X2 \AES_ENC/u0/u1/U298  ( .A1(\AES_ENC/u0/u1/n1095 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n668 ) );
NOR2_X2 \AES_ENC/u0/u1/U297  ( .A1(\AES_ENC/u0/u1/n826 ), .A2(\AES_ENC/u0/u1/n573 ), .ZN(\AES_ENC/u0/u1/n750 ) );
NOR2_X2 \AES_ENC/u0/u1/U296  ( .A1(\AES_ENC/u0/u1/n750 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n751 ) );
NOR2_X2 \AES_ENC/u0/u1/U295  ( .A1(\AES_ENC/u0/u1/n907 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n908 ) );
NOR2_X2 \AES_ENC/u0/u1/U294  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n588 ), .ZN(\AES_ENC/u0/u1/n957 ) );
NOR2_X2 \AES_ENC/u0/u1/U293  ( .A1(\AES_ENC/u0/u1/n990 ), .A2(\AES_ENC/u0/u1/n926 ), .ZN(\AES_ENC/u0/u1/n780 ) );
NOR2_X2 \AES_ENC/u0/u1/U292  ( .A1(\AES_ENC/u0/u1/n1022 ), .A2(\AES_ENC/u0/u1/n1058 ), .ZN(\AES_ENC/u0/u1/n740 ) );
NOR2_X2 \AES_ENC/u0/u1/U291  ( .A1(\AES_ENC/u0/u1/n740 ), .A2(\AES_ENC/u0/u1/n616 ), .ZN(\AES_ENC/u0/u1/n742 ) );
NOR2_X2 \AES_ENC/u0/u1/U290  ( .A1(\AES_ENC/u0/u1/n1098 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n1099 ) );
NOR2_X2 \AES_ENC/u0/u1/U284  ( .A1(\AES_ENC/u0/u1/n1120 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n993 ) );
NOR2_X2 \AES_ENC/u0/u1/U283  ( .A1(\AES_ENC/u0/u1/n993 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n994 ) );
NOR2_X2 \AES_ENC/u0/u1/U282  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n620 ), .ZN(\AES_ENC/u0/u1/n1026 ) );
NOR2_X2 \AES_ENC/u0/u1/U281  ( .A1(\AES_ENC/u0/u1/n573 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n1027 ) );
NOR2_X2 \AES_ENC/u0/u1/U280  ( .A1(\AES_ENC/u0/u1/n1027 ), .A2(\AES_ENC/u0/u1/n1026 ), .ZN(\AES_ENC/u0/u1/n1028 ) );
NOR2_X2 \AES_ENC/u0/u1/U279  ( .A1(\AES_ENC/u0/u1/n1029 ), .A2(\AES_ENC/u0/u1/n1028 ), .ZN(\AES_ENC/u0/u1/n1034 ) );
NOR2_X2 \AES_ENC/u0/u1/U273  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n1071 ), .ZN(\AES_ENC/u0/u1/n669 ) );
NOR2_X2 \AES_ENC/u0/u1/U272  ( .A1(\AES_ENC/u0/u1/n1056 ), .A2(\AES_ENC/u0/u1/n990 ), .ZN(\AES_ENC/u0/u1/n991 ) );
NOR2_X2 \AES_ENC/u0/u1/U271  ( .A1(\AES_ENC/u0/u1/n991 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n995 ) );
NOR4_X2 \AES_ENC/u0/u1/U270  ( .A1(\AES_ENC/u0/u1/n757 ), .A2(\AES_ENC/u0/u1/n756 ), .A3(\AES_ENC/u0/u1/n755 ), .A4(\AES_ENC/u0/u1/n754 ), .ZN(\AES_ENC/u0/u1/n758 ) );
NOR2_X2 \AES_ENC/u0/u1/U269  ( .A1(\AES_ENC/u0/u1/n752 ), .A2(\AES_ENC/u0/u1/n751 ), .ZN(\AES_ENC/u0/u1/n759 ) );
NOR2_X2 \AES_ENC/u0/u1/U268  ( .A1(\AES_ENC/u0/u1/n607 ), .A2(\AES_ENC/u0/u1/n590 ), .ZN(\AES_ENC/u0/u1/n1008 ) );
NOR2_X2 \AES_ENC/u0/u1/U267  ( .A1(\AES_ENC/u0/u1/n606 ), .A2(\AES_ENC/u0/u1/n906 ), .ZN(\AES_ENC/u0/u1/n741 ) );
NOR2_X2 \AES_ENC/u0/u1/U263  ( .A1(\AES_ENC/u0/u1/n1054 ), .A2(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n763 ) );
NOR2_X2 \AES_ENC/u0/u1/U262  ( .A1(\AES_ENC/u0/u1/n763 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n769 ) );
NOR2_X2 \AES_ENC/u0/u1/U258  ( .A1(\AES_ENC/u0/u1/n839 ), .A2(\AES_ENC/u0/u1/n582 ), .ZN(\AES_ENC/u0/u1/n693 ) );
NOR2_X2 \AES_ENC/u0/u1/U255  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n577 ), .ZN(\AES_ENC/u0/u1/n1007 ) );
NOR2_X2 \AES_ENC/u0/u1/U254  ( .A1(\AES_ENC/u0/u1/n609 ), .A2(\AES_ENC/u0/u1/n580 ), .ZN(\AES_ENC/u0/u1/n1123 ) );
NOR2_X2 \AES_ENC/u0/u1/U253  ( .A1(\AES_ENC/u0/u1/n780 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n784 ) );
NOR2_X2 \AES_ENC/u0/u1/U252  ( .A1(\AES_ENC/u0/u1/n1117 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n782 ) );
NOR2_X2 \AES_ENC/u0/u1/U251  ( .A1(\AES_ENC/u0/u1/n781 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n783 ) );
NOR4_X2 \AES_ENC/u0/u1/U250  ( .A1(\AES_ENC/u0/u1/n880 ), .A2(\AES_ENC/u0/u1/n784 ), .A3(\AES_ENC/u0/u1/n783 ), .A4(\AES_ENC/u0/u1/n782 ), .ZN(\AES_ENC/u0/u1/n785 ) );
NOR2_X2 \AES_ENC/u0/u1/U243  ( .A1(\AES_ENC/u0/u1/n609 ), .A2(\AES_ENC/u0/u1/n590 ), .ZN(\AES_ENC/u0/u1/n710 ) );
INV_X4 \AES_ENC/u0/u1/U242  ( .A(\AES_ENC/u0/u1/n1029 ), .ZN(\AES_ENC/u0/u1/n582 ) );
NOR2_X2 \AES_ENC/u0/u1/U241  ( .A1(\AES_ENC/u0/u1/n593 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n1125 ) );
NOR2_X2 \AES_ENC/u0/u1/U240  ( .A1(\AES_ENC/u0/u1/n616 ), .A2(\AES_ENC/u0/u1/n580 ), .ZN(\AES_ENC/u0/u1/n771 ) );
NOR2_X2 \AES_ENC/u0/u1/U239  ( .A1(\AES_ENC/u0/u1/n616 ), .A2(\AES_ENC/u0/u1/n597 ), .ZN(\AES_ENC/u0/u1/n883 ) );
NOR2_X2 \AES_ENC/u0/u1/U238  ( .A1(\AES_ENC/u0/u1/n911 ), .A2(\AES_ENC/u0/u1/n910 ), .ZN(\AES_ENC/u0/u1/n912 ) );
NOR2_X2 \AES_ENC/u0/u1/U237  ( .A1(\AES_ENC/u0/u1/n912 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n916 ) );
NOR2_X2 \AES_ENC/u0/u1/U236  ( .A1(\AES_ENC/u0/u1/n990 ), .A2(\AES_ENC/u0/u1/n929 ), .ZN(\AES_ENC/u0/u1/n892 ) );
NOR2_X2 \AES_ENC/u0/u1/U235  ( .A1(\AES_ENC/u0/u1/n892 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n893 ) );
NOR2_X2 \AES_ENC/u0/u1/U234  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n602 ), .ZN(\AES_ENC/u0/u1/n950 ) );
NOR2_X2 \AES_ENC/u0/u1/U229  ( .A1(\AES_ENC/u0/u1/n1079 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n1082 ) );
NOR2_X2 \AES_ENC/u0/u1/U228  ( .A1(\AES_ENC/u0/u1/n910 ), .A2(\AES_ENC/u0/u1/n1056 ), .ZN(\AES_ENC/u0/u1/n941 ) );
NOR2_X2 \AES_ENC/u0/u1/U227  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n1077 ), .ZN(\AES_ENC/u0/u1/n841 ) );
NOR2_X2 \AES_ENC/u0/u1/U226  ( .A1(\AES_ENC/u0/u1/n623 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n630 ) );
NOR2_X2 \AES_ENC/u0/u1/U225  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n602 ), .ZN(\AES_ENC/u0/u1/n806 ) );
NOR2_X2 \AES_ENC/u0/u1/U223  ( .A1(\AES_ENC/u0/u1/n623 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n948 ) );
NOR2_X2 \AES_ENC/u0/u1/U222  ( .A1(\AES_ENC/u0/u1/n606 ), .A2(\AES_ENC/u0/u1/n582 ), .ZN(\AES_ENC/u0/u1/n1104 ) );
NOR2_X2 \AES_ENC/u0/u1/U221  ( .A1(\AES_ENC/u0/u1/n1121 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n1122 ) );
NOR2_X2 \AES_ENC/u0/u1/U217  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n1023 ), .ZN(\AES_ENC/u0/u1/n756 ) );
NOR2_X2 \AES_ENC/u0/u1/U213  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n602 ), .ZN(\AES_ENC/u0/u1/n870 ) );
NOR2_X2 \AES_ENC/u0/u1/U212  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n569 ), .ZN(\AES_ENC/u0/u1/n947 ) );
NOR2_X2 \AES_ENC/u0/u1/U211  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n1077 ), .ZN(\AES_ENC/u0/u1/n1084 ) );
NOR2_X2 \AES_ENC/u0/u1/U210  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n855 ), .ZN(\AES_ENC/u0/u1/n709 ) );
NOR2_X2 \AES_ENC/u0/u1/U209  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n589 ), .ZN(\AES_ENC/u0/u1/n868 ) );
NOR2_X2 \AES_ENC/u0/u1/U208  ( .A1(\AES_ENC/u0/u1/n1120 ), .A2(\AES_ENC/u0/u1/n839 ), .ZN(\AES_ENC/u0/u1/n842 ) );
NOR2_X2 \AES_ENC/u0/u1/U207  ( .A1(\AES_ENC/u0/u1/n1120 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n1124 ) );
NOR2_X2 \AES_ENC/u0/u1/U201  ( .A1(\AES_ENC/u0/u1/n1120 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n696 ) );
NOR2_X2 \AES_ENC/u0/u1/U200  ( .A1(\AES_ENC/u0/u1/n1074 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n1076 ) );
NOR2_X2 \AES_ENC/u0/u1/U199  ( .A1(\AES_ENC/u0/u1/n1074 ), .A2(\AES_ENC/u0/u1/n620 ), .ZN(\AES_ENC/u0/u1/n781 ) );
NOR3_X2 \AES_ENC/u0/u1/U198  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n1056 ), .A3(\AES_ENC/u0/u1/n990 ), .ZN(\AES_ENC/u0/u1/n979 ) );
NOR3_X2 \AES_ENC/u0/u1/U197  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n1058 ), .A3(\AES_ENC/u0/u1/n1059 ), .ZN(\AES_ENC/u0/u1/n854 ) );
NOR2_X2 \AES_ENC/u0/u1/U196  ( .A1(\AES_ENC/u0/u1/n996 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n869 ) );
NOR2_X2 \AES_ENC/u0/u1/U195  ( .A1(\AES_ENC/u0/u1/n1056 ), .A2(\AES_ENC/u0/u1/n1074 ), .ZN(\AES_ENC/u0/u1/n1057 ) );
NOR3_X2 \AES_ENC/u0/u1/U194  ( .A1(\AES_ENC/u0/u1/n607 ), .A2(\AES_ENC/u0/u1/n1120 ), .A3(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n978 ) );
NOR2_X2 \AES_ENC/u0/u1/U187  ( .A1(\AES_ENC/u0/u1/n996 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n998 ) );
NOR2_X2 \AES_ENC/u0/u1/U186  ( .A1(\AES_ENC/u0/u1/n996 ), .A2(\AES_ENC/u0/u1/n911 ), .ZN(\AES_ENC/u0/u1/n1116 ) );
NOR2_X2 \AES_ENC/u0/u1/U185  ( .A1(\AES_ENC/u0/u1/n1074 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n754 ) );
NOR2_X2 \AES_ENC/u0/u1/U184  ( .A1(\AES_ENC/u0/u1/n926 ), .A2(\AES_ENC/u0/u1/n1103 ), .ZN(\AES_ENC/u0/u1/n977 ) );
NOR2_X2 \AES_ENC/u0/u1/U183  ( .A1(\AES_ENC/u0/u1/n839 ), .A2(\AES_ENC/u0/u1/n824 ), .ZN(\AES_ENC/u0/u1/n1092 ) );
NOR2_X2 \AES_ENC/u0/u1/U182  ( .A1(\AES_ENC/u0/u1/n573 ), .A2(\AES_ENC/u0/u1/n1074 ), .ZN(\AES_ENC/u0/u1/n684 ) );
NOR2_X2 \AES_ENC/u0/u1/U181  ( .A1(\AES_ENC/u0/u1/n826 ), .A2(\AES_ENC/u0/u1/n1059 ), .ZN(\AES_ENC/u0/u1/n907 ) );
NOR3_X2 \AES_ENC/u0/u1/U180  ( .A1(\AES_ENC/u0/u1/n625 ), .A2(\AES_ENC/u0/u1/n1115 ), .A3(\AES_ENC/u0/u1/n585 ), .ZN(\AES_ENC/u0/u1/n831 ) );
NOR3_X2 \AES_ENC/u0/u1/U174  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n1056 ), .A3(\AES_ENC/u0/u1/n990 ), .ZN(\AES_ENC/u0/u1/n896 ) );
NOR3_X2 \AES_ENC/u0/u1/U173  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n573 ), .A3(\AES_ENC/u0/u1/n1013 ), .ZN(\AES_ENC/u0/u1/n670 ) );
NOR3_X2 \AES_ENC/u0/u1/U172  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n1091 ), .A3(\AES_ENC/u0/u1/n1022 ), .ZN(\AES_ENC/u0/u1/n843 ) );
NOR2_X2 \AES_ENC/u0/u1/U171  ( .A1(\AES_ENC/u0/u1/n1029 ), .A2(\AES_ENC/u0/u1/n1095 ), .ZN(\AES_ENC/u0/u1/n735 ) );
NAND3_X2 \AES_ENC/u0/u1/U170  ( .A1(\AES_ENC/u0/u1/n569 ), .A2(\AES_ENC/u0/u1/n582 ), .A3(\AES_ENC/u0/u1/n681 ), .ZN(\AES_ENC/u0/u1/n691 ) );
NOR2_X2 \AES_ENC/u0/u1/U169  ( .A1(\AES_ENC/u0/u1/n683 ), .A2(\AES_ENC/u0/u1/n682 ), .ZN(\AES_ENC/u0/u1/n690 ) );
NOR4_X2 \AES_ENC/u0/u1/U168  ( .A1(\AES_ENC/u0/u1/n983 ), .A2(\AES_ENC/u0/u1/n698 ), .A3(\AES_ENC/u0/u1/n697 ), .A4(\AES_ENC/u0/u1/n696 ), .ZN(\AES_ENC/u0/u1/n699 ) );
NOR3_X2 \AES_ENC/u0/u1/U162  ( .A1(\AES_ENC/u0/u1/n695 ), .A2(\AES_ENC/u0/u1/n694 ), .A3(\AES_ENC/u0/u1/n693 ), .ZN(\AES_ENC/u0/u1/n700 ) );
NOR2_X2 \AES_ENC/u0/u1/U161  ( .A1(\AES_ENC/u0/u1/n1100 ), .A2(\AES_ENC/u0/u1/n854 ), .ZN(\AES_ENC/u0/u1/n860 ) );
NOR4_X2 \AES_ENC/u0/u1/U160  ( .A1(\AES_ENC/u0/u1/n896 ), .A2(\AES_ENC/u0/u1/n895 ), .A3(\AES_ENC/u0/u1/n894 ), .A4(\AES_ENC/u0/u1/n893 ), .ZN(\AES_ENC/u0/u1/n897 ) );
NOR2_X2 \AES_ENC/u0/u1/U159  ( .A1(\AES_ENC/u0/u1/n866 ), .A2(\AES_ENC/u0/u1/n865 ), .ZN(\AES_ENC/u0/u1/n872 ) );
NOR4_X2 \AES_ENC/u0/u1/U158  ( .A1(\AES_ENC/u0/u1/n870 ), .A2(\AES_ENC/u0/u1/n869 ), .A3(\AES_ENC/u0/u1/n868 ), .A4(\AES_ENC/u0/u1/n867 ), .ZN(\AES_ENC/u0/u1/n871 ) );
NOR4_X2 \AES_ENC/u0/u1/U157  ( .A1(\AES_ENC/u0/u1/n963 ), .A2(\AES_ENC/u0/u1/n962 ), .A3(\AES_ENC/u0/u1/n961 ), .A4(\AES_ENC/u0/u1/n960 ), .ZN(\AES_ENC/u0/u1/n964 ) );
NOR2_X2 \AES_ENC/u0/u1/U156  ( .A1(\AES_ENC/u0/u1/n958 ), .A2(\AES_ENC/u0/u1/n957 ), .ZN(\AES_ENC/u0/u1/n965 ) );
NOR4_X2 \AES_ENC/u0/u1/U155  ( .A1(\AES_ENC/u0/u1/n950 ), .A2(\AES_ENC/u0/u1/n949 ), .A3(\AES_ENC/u0/u1/n948 ), .A4(\AES_ENC/u0/u1/n947 ), .ZN(\AES_ENC/u0/u1/n951 ) );
NOR2_X2 \AES_ENC/u0/u1/U154  ( .A1(\AES_ENC/u0/u1/n946 ), .A2(\AES_ENC/u0/u1/n945 ), .ZN(\AES_ENC/u0/u1/n952 ) );
NOR4_X2 \AES_ENC/u0/u1/U153  ( .A1(\AES_ENC/u0/u1/n983 ), .A2(\AES_ENC/u0/u1/n982 ), .A3(\AES_ENC/u0/u1/n981 ), .A4(\AES_ENC/u0/u1/n980 ), .ZN(\AES_ENC/u0/u1/n984 ) );
NOR2_X2 \AES_ENC/u0/u1/U152  ( .A1(\AES_ENC/u0/u1/n979 ), .A2(\AES_ENC/u0/u1/n978 ), .ZN(\AES_ENC/u0/u1/n985 ) );
NOR4_X2 \AES_ENC/u0/u1/U143  ( .A1(\AES_ENC/u0/u1/n1125 ), .A2(\AES_ENC/u0/u1/n1124 ), .A3(\AES_ENC/u0/u1/n1123 ), .A4(\AES_ENC/u0/u1/n1122 ), .ZN(\AES_ENC/u0/u1/n1126 ) );
NOR4_X2 \AES_ENC/u0/u1/U142  ( .A1(\AES_ENC/u0/u1/n1084 ), .A2(\AES_ENC/u0/u1/n1083 ), .A3(\AES_ENC/u0/u1/n1082 ), .A4(\AES_ENC/u0/u1/n1081 ), .ZN(\AES_ENC/u0/u1/n1085 ) );
NOR2_X2 \AES_ENC/u0/u1/U141  ( .A1(\AES_ENC/u0/u1/n1076 ), .A2(\AES_ENC/u0/u1/n1075 ), .ZN(\AES_ENC/u0/u1/n1086 ) );
NOR3_X2 \AES_ENC/u0/u1/U140  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n1054 ), .A3(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n961 ) );
NOR3_X2 \AES_ENC/u0/u1/U132  ( .A1(\AES_ENC/u0/u1/n620 ), .A2(\AES_ENC/u0/u1/n1074 ), .A3(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n671 ) );
NOR2_X2 \AES_ENC/u0/u1/U131  ( .A1(\AES_ENC/u0/u1/n1057 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n1062 ) );
NOR2_X2 \AES_ENC/u0/u1/U130  ( .A1(\AES_ENC/u0/u1/n1060 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n1061 ) );
NOR2_X2 \AES_ENC/u0/u1/U129  ( .A1(\AES_ENC/u0/u1/n1055 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n1063 ) );
NOR4_X2 \AES_ENC/u0/u1/U128  ( .A1(\AES_ENC/u0/u1/n1064 ), .A2(\AES_ENC/u0/u1/n1063 ), .A3(\AES_ENC/u0/u1/n1062 ), .A4(\AES_ENC/u0/u1/n1061 ), .ZN(\AES_ENC/u0/u1/n1065 ) );
NOR3_X2 \AES_ENC/u0/u1/U127  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n1120 ), .A3(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n918 ) );
NOR2_X2 \AES_ENC/u0/u1/U126  ( .A1(\AES_ENC/u0/u1/n914 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n915 ) );
NOR3_X2 \AES_ENC/u0/u1/U121  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n573 ), .A3(\AES_ENC/u0/u1/n1013 ), .ZN(\AES_ENC/u0/u1/n917 ) );
NOR4_X2 \AES_ENC/u0/u1/U120  ( .A1(\AES_ENC/u0/u1/n918 ), .A2(\AES_ENC/u0/u1/n917 ), .A3(\AES_ENC/u0/u1/n916 ), .A4(\AES_ENC/u0/u1/n915 ), .ZN(\AES_ENC/u0/u1/n919 ) );
NOR2_X2 \AES_ENC/u0/u1/U119  ( .A1(\AES_ENC/u0/u1/n735 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n687 ) );
NOR2_X2 \AES_ENC/u0/u1/U118  ( .A1(\AES_ENC/u0/u1/n684 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n688 ) );
NOR2_X2 \AES_ENC/u0/u1/U117  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n600 ), .ZN(\AES_ENC/u0/u1/n686 ) );
NOR4_X2 \AES_ENC/u0/u1/U116  ( .A1(\AES_ENC/u0/u1/n688 ), .A2(\AES_ENC/u0/u1/n687 ), .A3(\AES_ENC/u0/u1/n686 ), .A4(\AES_ENC/u0/u1/n685 ), .ZN(\AES_ENC/u0/u1/n689 ) );
NOR2_X2 \AES_ENC/u0/u1/U115  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n582 ), .ZN(\AES_ENC/u0/u1/n770 ) );
NOR2_X2 \AES_ENC/u0/u1/U106  ( .A1(\AES_ENC/u0/u1/n1103 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n772 ) );
NOR2_X2 \AES_ENC/u0/u1/U105  ( .A1(\AES_ENC/u0/u1/n610 ), .A2(\AES_ENC/u0/u1/n599 ), .ZN(\AES_ENC/u0/u1/n773 ) );
NOR4_X2 \AES_ENC/u0/u1/U104  ( .A1(\AES_ENC/u0/u1/n773 ), .A2(\AES_ENC/u0/u1/n772 ), .A3(\AES_ENC/u0/u1/n771 ), .A4(\AES_ENC/u0/u1/n770 ), .ZN(\AES_ENC/u0/u1/n774 ) );
NOR2_X2 \AES_ENC/u0/u1/U103  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n595 ), .ZN(\AES_ENC/u0/u1/n858 ) );
NOR2_X2 \AES_ENC/u0/u1/U102  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n855 ), .ZN(\AES_ENC/u0/u1/n857 ) );
NOR2_X2 \AES_ENC/u0/u1/U101  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n587 ), .ZN(\AES_ENC/u0/u1/n856 ) );
NOR4_X2 \AES_ENC/u0/u1/U100  ( .A1(\AES_ENC/u0/u1/n858 ), .A2(\AES_ENC/u0/u1/n857 ), .A3(\AES_ENC/u0/u1/n856 ), .A4(\AES_ENC/u0/u1/n958 ), .ZN(\AES_ENC/u0/u1/n859 ) );
NOR2_X2 \AES_ENC/u0/u1/U95  ( .A1(\AES_ENC/u0/u1/n583 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n814 ) );
NOR3_X2 \AES_ENC/u0/u1/U94  ( .A1(\AES_ENC/u0/u1/n606 ), .A2(\AES_ENC/u0/u1/n1058 ), .A3(\AES_ENC/u0/u1/n1059 ), .ZN(\AES_ENC/u0/u1/n815 ) );
NOR2_X2 \AES_ENC/u0/u1/U93  ( .A1(\AES_ENC/u0/u1/n907 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n813 ) );
NOR4_X2 \AES_ENC/u0/u1/U92  ( .A1(\AES_ENC/u0/u1/n815 ), .A2(\AES_ENC/u0/u1/n814 ), .A3(\AES_ENC/u0/u1/n813 ), .A4(\AES_ENC/u0/u1/n812 ), .ZN(\AES_ENC/u0/u1/n816 ) );
NOR2_X2 \AES_ENC/u0/u1/U91  ( .A1(\AES_ENC/u0/u1/n617 ), .A2(\AES_ENC/u0/u1/n569 ), .ZN(\AES_ENC/u0/u1/n721 ) );
NOR2_X2 \AES_ENC/u0/u1/U90  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n1096 ), .ZN(\AES_ENC/u0/u1/n722 ) );
NOR2_X2 \AES_ENC/u0/u1/U89  ( .A1(\AES_ENC/u0/u1/n1031 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n723 ) );
NOR4_X2 \AES_ENC/u0/u1/U88  ( .A1(\AES_ENC/u0/u1/n724 ), .A2(\AES_ENC/u0/u1/n723 ), .A3(\AES_ENC/u0/u1/n722 ), .A4(\AES_ENC/u0/u1/n721 ), .ZN(\AES_ENC/u0/u1/n725 ) );
NOR2_X2 \AES_ENC/u0/u1/U87  ( .A1(\AES_ENC/u0/u1/n911 ), .A2(\AES_ENC/u0/u1/n990 ), .ZN(\AES_ENC/u0/u1/n1009 ) );
NOR2_X2 \AES_ENC/u0/u1/U86  ( .A1(\AES_ENC/u0/u1/n1013 ), .A2(\AES_ENC/u0/u1/n573 ), .ZN(\AES_ENC/u0/u1/n1014 ) );
NOR2_X2 \AES_ENC/u0/u1/U81  ( .A1(\AES_ENC/u0/u1/n1014 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n1015 ) );
NOR4_X2 \AES_ENC/u0/u1/U80  ( .A1(\AES_ENC/u0/u1/n1016 ), .A2(\AES_ENC/u0/u1/n1015 ), .A3(\AES_ENC/u0/u1/n1119 ), .A4(\AES_ENC/u0/u1/n1046 ), .ZN(\AES_ENC/u0/u1/n1017 ) );
NOR2_X2 \AES_ENC/u0/u1/U79  ( .A1(\AES_ENC/u0/u1/n606 ), .A2(\AES_ENC/u0/u1/n589 ), .ZN(\AES_ENC/u0/u1/n997 ) );
NOR2_X2 \AES_ENC/u0/u1/U78  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n577 ), .ZN(\AES_ENC/u0/u1/n1000 ) );
NOR2_X2 \AES_ENC/u0/u1/U74  ( .A1(\AES_ENC/u0/u1/n616 ), .A2(\AES_ENC/u0/u1/n1096 ), .ZN(\AES_ENC/u0/u1/n999 ) );
NOR4_X2 \AES_ENC/u0/u1/U73  ( .A1(\AES_ENC/u0/u1/n1000 ), .A2(\AES_ENC/u0/u1/n999 ), .A3(\AES_ENC/u0/u1/n998 ), .A4(\AES_ENC/u0/u1/n997 ), .ZN(\AES_ENC/u0/u1/n1001 ) );
NOR2_X2 \AES_ENC/u0/u1/U72  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n1096 ), .ZN(\AES_ENC/u0/u1/n697 ) );
NOR2_X2 \AES_ENC/u0/u1/U71  ( .A1(\AES_ENC/u0/u1/n620 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n958 ) );
NOR2_X2 \AES_ENC/u0/u1/U65  ( .A1(\AES_ENC/u0/u1/n911 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n983 ) );
NOR2_X2 \AES_ENC/u0/u1/U64  ( .A1(\AES_ENC/u0/u1/n1054 ), .A2(\AES_ENC/u0/u1/n1103 ), .ZN(\AES_ENC/u0/u1/n1031 ) );
INV_X4 \AES_ENC/u0/u1/U63  ( .A(\AES_ENC/u0/u1/n1050 ), .ZN(\AES_ENC/u0/u1/n612 ) );
INV_X4 \AES_ENC/u0/u1/U62  ( .A(\AES_ENC/u0/u1/n1072 ), .ZN(\AES_ENC/u0/u1/n605 ) );
INV_X4 \AES_ENC/u0/u1/U61  ( .A(\AES_ENC/u0/u1/n1073 ), .ZN(\AES_ENC/u0/u1/n604 ) );
NOR2_X2 \AES_ENC/u0/u1/U59  ( .A1(\AES_ENC/u0/u1/n582 ), .A2(\AES_ENC/u0/u1/n613 ), .ZN(\AES_ENC/u0/u1/n880 ) );
NOR3_X2 \AES_ENC/u0/u1/U58  ( .A1(\AES_ENC/u0/u1/n826 ), .A2(\AES_ENC/u0/u1/n1121 ), .A3(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n946 ) );
INV_X4 \AES_ENC/u0/u1/U57  ( .A(\AES_ENC/u0/u1/n1010 ), .ZN(\AES_ENC/u0/u1/n608 ) );
NOR3_X2 \AES_ENC/u0/u1/U50  ( .A1(\AES_ENC/u0/u1/n573 ), .A2(\AES_ENC/u0/u1/n1029 ), .A3(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n1119 ) );
INV_X4 \AES_ENC/u0/u1/U49  ( .A(\AES_ENC/u0/u1/n956 ), .ZN(\AES_ENC/u0/u1/n615 ) );
NOR2_X2 \AES_ENC/u0/u1/U48  ( .A1(\AES_ENC/u0/u1/n623 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n1013 ) );
NOR2_X2 \AES_ENC/u0/u1/U47  ( .A1(\AES_ENC/u0/u1/n620 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n910 ) );
NOR2_X2 \AES_ENC/u0/u1/U46  ( .A1(\AES_ENC/u0/u1/n569 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n1091 ) );
NOR2_X2 \AES_ENC/u0/u1/U45  ( .A1(\AES_ENC/u0/u1/n622 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n990 ) );
NOR2_X2 \AES_ENC/u0/u1/U44  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/u0/u1/n1121 ), .ZN(\AES_ENC/u0/u1/n996 ) );
NOR2_X2 \AES_ENC/u0/u1/U43  ( .A1(\AES_ENC/u0/u1/n610 ), .A2(\AES_ENC/u0/u1/n600 ), .ZN(\AES_ENC/u0/u1/n628 ) );
NOR2_X2 \AES_ENC/u0/u1/U42  ( .A1(\AES_ENC/u0/u1/n576 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n866 ) );
NOR2_X2 \AES_ENC/u0/u1/U41  ( .A1(\AES_ENC/u0/u1/n603 ), .A2(\AES_ENC/u0/u1/n610 ), .ZN(\AES_ENC/u0/u1/n1006 ) );
NOR2_X2 \AES_ENC/u0/u1/U36  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n1117 ), .ZN(\AES_ENC/u0/u1/n1118 ) );
NOR2_X2 \AES_ENC/u0/u1/U35  ( .A1(\AES_ENC/u0/u1/n1119 ), .A2(\AES_ENC/u0/u1/n1118 ), .ZN(\AES_ENC/u0/u1/n1127 ) );
NOR2_X2 \AES_ENC/u0/u1/U34  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n594 ), .ZN(\AES_ENC/u0/u1/n629 ) );
NOR2_X2 \AES_ENC/u0/u1/U33  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n906 ), .ZN(\AES_ENC/u0/u1/n909 ) );
NOR2_X2 \AES_ENC/u0/u1/U32  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n597 ), .ZN(\AES_ENC/u0/u1/n658 ) );
NOR2_X2 \AES_ENC/u0/u1/U31  ( .A1(\AES_ENC/u0/u1/n1116 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n695 ) );
NOR2_X2 \AES_ENC/u0/u1/U30  ( .A1(\AES_ENC/u0/u1/n1078 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n1083 ) );
NOR2_X2 \AES_ENC/u0/u1/U29  ( .A1(\AES_ENC/u0/u1/n941 ), .A2(\AES_ENC/u0/u1/n608 ), .ZN(\AES_ENC/u0/u1/n724 ) );
NOR2_X2 \AES_ENC/u0/u1/U24  ( .A1(\AES_ENC/u0/u1/n576 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n840 ) );
NOR2_X2 \AES_ENC/u0/u1/U23  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n593 ), .ZN(\AES_ENC/u0/u1/n633 ) );
NOR2_X2 \AES_ENC/u0/u1/U21  ( .A1(\AES_ENC/u0/u1/n1009 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n960 ) );
NOR2_X2 \AES_ENC/u0/u1/U20  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n1045 ), .ZN(\AES_ENC/u0/u1/n812 ) );
NOR2_X2 \AES_ENC/u0/u1/U19  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n1080 ), .ZN(\AES_ENC/u0/u1/n1081 ) );
NOR2_X2 \AES_ENC/u0/u1/U18  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n601 ), .ZN(\AES_ENC/u0/u1/n982 ) );
NOR2_X2 \AES_ENC/u0/u1/U17  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n594 ), .ZN(\AES_ENC/u0/u1/n757 ) );
NOR2_X2 \AES_ENC/u0/u1/U16  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n590 ), .ZN(\AES_ENC/u0/u1/n698 ) );
NOR2_X2 \AES_ENC/u0/u1/U15  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n619 ), .ZN(\AES_ENC/u0/u1/n708 ) );
NOR2_X2 \AES_ENC/u0/u1/U10  ( .A1(\AES_ENC/u0/u1/n619 ), .A2(\AES_ENC/u0/u1/n604 ), .ZN(\AES_ENC/u0/u1/n803 ) );
NOR2_X2 \AES_ENC/u0/u1/U9  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n881 ), .ZN(\AES_ENC/u0/u1/n711 ) );
NOR2_X2 \AES_ENC/u0/u1/U8  ( .A1(\AES_ENC/u0/u1/n615 ), .A2(\AES_ENC/u0/u1/n582 ), .ZN(\AES_ENC/u0/u1/n867 ) );
NOR2_X2 \AES_ENC/u0/u1/U7  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n599 ), .ZN(\AES_ENC/u0/u1/n804 ) );
NOR2_X2 \AES_ENC/u0/u1/U6  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n620 ), .ZN(\AES_ENC/u0/u1/n1046 ) );
OR2_X4 \AES_ENC/u0/u1/U5  ( .A1(\AES_ENC/u0/u1/n624 ), .A2(\AES_ENC/w3[9] ),.ZN(\AES_ENC/u0/u1/n570 ) );
OR2_X4 \AES_ENC/u0/u1/U4  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/w3[12] ),.ZN(\AES_ENC/u0/u1/n569 ) );
NAND2_X2 \AES_ENC/u0/u1/U514  ( .A1(\AES_ENC/u0/u1/n1121 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n1030 ) );
AND2_X2 \AES_ENC/u0/u1/U513  ( .A1(\AES_ENC/u0/u1/n597 ), .A2(\AES_ENC/u0/u1/n1030 ), .ZN(\AES_ENC/u0/u1/n1049 ) );
NAND2_X2 \AES_ENC/u0/u1/U511  ( .A1(\AES_ENC/u0/u1/n1049 ), .A2(\AES_ENC/u0/u1/n794 ), .ZN(\AES_ENC/u0/u1/n637 ) );
AND2_X2 \AES_ENC/u0/u1/U493  ( .A1(\AES_ENC/u0/u1/n779 ), .A2(\AES_ENC/u0/u1/n996 ), .ZN(\AES_ENC/u0/u1/n632 ) );
NAND4_X2 \AES_ENC/u0/u1/U485  ( .A1(\AES_ENC/u0/u1/n637 ), .A2(\AES_ENC/u0/u1/n636 ), .A3(\AES_ENC/u0/u1/n635 ), .A4(\AES_ENC/u0/u1/n634 ), .ZN(\AES_ENC/u0/u1/n638 ) );
NAND2_X2 \AES_ENC/u0/u1/U484  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n638 ), .ZN(\AES_ENC/u0/u1/n679 ) );
NAND2_X2 \AES_ENC/u0/u1/U481  ( .A1(\AES_ENC/u0/u1/n1094 ), .A2(\AES_ENC/u0/u1/n591 ), .ZN(\AES_ENC/u0/u1/n648 ) );
NAND2_X2 \AES_ENC/u0/u1/U476  ( .A1(\AES_ENC/u0/u1/n601 ), .A2(\AES_ENC/u0/u1/n590 ), .ZN(\AES_ENC/u0/u1/n762 ) );
NAND2_X2 \AES_ENC/u0/u1/U475  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n762 ), .ZN(\AES_ENC/u0/u1/n647 ) );
NAND4_X2 \AES_ENC/u0/u1/U457  ( .A1(\AES_ENC/u0/u1/n648 ), .A2(\AES_ENC/u0/u1/n647 ), .A3(\AES_ENC/u0/u1/n646 ), .A4(\AES_ENC/u0/u1/n645 ), .ZN(\AES_ENC/u0/u1/n649 ) );
NAND2_X2 \AES_ENC/u0/u1/U456  ( .A1(\AES_ENC/w3[8] ), .A2(\AES_ENC/u0/u1/n649 ), .ZN(\AES_ENC/u0/u1/n665 ) );
NAND2_X2 \AES_ENC/u0/u1/U454  ( .A1(\AES_ENC/u0/u1/n596 ), .A2(\AES_ENC/u0/u1/n623 ), .ZN(\AES_ENC/u0/u1/n855 ) );
NAND2_X2 \AES_ENC/u0/u1/U453  ( .A1(\AES_ENC/u0/u1/n587 ), .A2(\AES_ENC/u0/u1/n855 ), .ZN(\AES_ENC/u0/u1/n821 ) );
NAND2_X2 \AES_ENC/u0/u1/U452  ( .A1(\AES_ENC/u0/u1/n1093 ), .A2(\AES_ENC/u0/u1/n821 ), .ZN(\AES_ENC/u0/u1/n662 ) );
NAND2_X2 \AES_ENC/u0/u1/U451  ( .A1(\AES_ENC/u0/u1/n619 ), .A2(\AES_ENC/u0/u1/n589 ), .ZN(\AES_ENC/u0/u1/n650 ) );
NAND2_X2 \AES_ENC/u0/u1/U450  ( .A1(\AES_ENC/u0/u1/n956 ), .A2(\AES_ENC/u0/u1/n650 ), .ZN(\AES_ENC/u0/u1/n661 ) );
NAND2_X2 \AES_ENC/u0/u1/U449  ( .A1(\AES_ENC/u0/u1/n626 ), .A2(\AES_ENC/u0/u1/n627 ), .ZN(\AES_ENC/u0/u1/n839 ) );
OR2_X2 \AES_ENC/u0/u1/U446  ( .A1(\AES_ENC/u0/u1/n839 ), .A2(\AES_ENC/u0/u1/n932 ), .ZN(\AES_ENC/u0/u1/n656 ) );
NAND2_X2 \AES_ENC/u0/u1/U445  ( .A1(\AES_ENC/u0/u1/n621 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n1096 ) );
NAND2_X2 \AES_ENC/u0/u1/U444  ( .A1(\AES_ENC/u0/u1/n1030 ), .A2(\AES_ENC/u0/u1/n1096 ), .ZN(\AES_ENC/u0/u1/n651 ) );
NAND2_X2 \AES_ENC/u0/u1/U443  ( .A1(\AES_ENC/u0/u1/n1114 ), .A2(\AES_ENC/u0/u1/n651 ), .ZN(\AES_ENC/u0/u1/n655 ) );
OR3_X2 \AES_ENC/u0/u1/U440  ( .A1(\AES_ENC/u0/u1/n1079 ), .A2(\AES_ENC/w3[15] ), .A3(\AES_ENC/u0/u1/n626 ), .ZN(\AES_ENC/u0/u1/n654 ) );
NAND2_X2 \AES_ENC/u0/u1/U439  ( .A1(\AES_ENC/u0/u1/n593 ), .A2(\AES_ENC/u0/u1/n601 ), .ZN(\AES_ENC/u0/u1/n652 ) );
NAND4_X2 \AES_ENC/u0/u1/U437  ( .A1(\AES_ENC/u0/u1/n656 ), .A2(\AES_ENC/u0/u1/n655 ), .A3(\AES_ENC/u0/u1/n654 ), .A4(\AES_ENC/u0/u1/n653 ), .ZN(\AES_ENC/u0/u1/n657 ) );
NAND2_X2 \AES_ENC/u0/u1/U436  ( .A1(\AES_ENC/w3[10] ), .A2(\AES_ENC/u0/u1/n657 ), .ZN(\AES_ENC/u0/u1/n660 ) );
NAND4_X2 \AES_ENC/u0/u1/U432  ( .A1(\AES_ENC/u0/u1/n662 ), .A2(\AES_ENC/u0/u1/n661 ), .A3(\AES_ENC/u0/u1/n660 ), .A4(\AES_ENC/u0/u1/n659 ), .ZN(\AES_ENC/u0/u1/n663 ) );
NAND2_X2 \AES_ENC/u0/u1/U431  ( .A1(\AES_ENC/u0/u1/n663 ), .A2(\AES_ENC/u0/u1/n574 ), .ZN(\AES_ENC/u0/u1/n664 ) );
NAND2_X2 \AES_ENC/u0/u1/U430  ( .A1(\AES_ENC/u0/u1/n665 ), .A2(\AES_ENC/u0/u1/n664 ), .ZN(\AES_ENC/u0/u1/n666 ) );
NAND2_X2 \AES_ENC/u0/u1/U429  ( .A1(\AES_ENC/w3[14] ), .A2(\AES_ENC/u0/u1/n666 ), .ZN(\AES_ENC/u0/u1/n678 ) );
NAND2_X2 \AES_ENC/u0/u1/U426  ( .A1(\AES_ENC/u0/u1/n735 ), .A2(\AES_ENC/u0/u1/n1093 ), .ZN(\AES_ENC/u0/u1/n675 ) );
NAND2_X2 \AES_ENC/u0/u1/U425  ( .A1(\AES_ENC/u0/u1/n588 ), .A2(\AES_ENC/u0/u1/n597 ), .ZN(\AES_ENC/u0/u1/n1045 ) );
OR2_X2 \AES_ENC/u0/u1/U424  ( .A1(\AES_ENC/u0/u1/n1045 ), .A2(\AES_ENC/u0/u1/n605 ), .ZN(\AES_ENC/u0/u1/n674 ) );
NAND2_X2 \AES_ENC/u0/u1/U423  ( .A1(\AES_ENC/w3[9] ), .A2(\AES_ENC/u0/u1/n620 ), .ZN(\AES_ENC/u0/u1/n667 ) );
NAND2_X2 \AES_ENC/u0/u1/U422  ( .A1(\AES_ENC/u0/u1/n619 ), .A2(\AES_ENC/u0/u1/n667 ), .ZN(\AES_ENC/u0/u1/n1071 ) );
NAND4_X2 \AES_ENC/u0/u1/U412  ( .A1(\AES_ENC/u0/u1/n675 ), .A2(\AES_ENC/u0/u1/n674 ), .A3(\AES_ENC/u0/u1/n673 ), .A4(\AES_ENC/u0/u1/n672 ), .ZN(\AES_ENC/u0/u1/n676 ) );
NAND2_X2 \AES_ENC/u0/u1/U411  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n676 ), .ZN(\AES_ENC/u0/u1/n677 ) );
NAND2_X2 \AES_ENC/u0/u1/U408  ( .A1(\AES_ENC/u0/u1/n800 ), .A2(\AES_ENC/u0/u1/n1022 ), .ZN(\AES_ENC/u0/u1/n680 ) );
NAND2_X2 \AES_ENC/u0/u1/U407  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n680 ), .ZN(\AES_ENC/u0/u1/n681 ) );
AND2_X2 \AES_ENC/u0/u1/U402  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n684 ), .ZN(\AES_ENC/u0/u1/n682 ) );
NAND4_X2 \AES_ENC/u0/u1/U395  ( .A1(\AES_ENC/u0/u1/n691 ), .A2(\AES_ENC/u0/u1/n581 ), .A3(\AES_ENC/u0/u1/n690 ), .A4(\AES_ENC/u0/u1/n689 ), .ZN(\AES_ENC/u0/u1/n692 ) );
NAND2_X2 \AES_ENC/u0/u1/U394  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n692 ), .ZN(\AES_ENC/u0/u1/n733 ) );
NAND2_X2 \AES_ENC/u0/u1/U392  ( .A1(\AES_ENC/u0/u1/n977 ), .A2(\AES_ENC/u0/u1/n1050 ), .ZN(\AES_ENC/u0/u1/n702 ) );
NAND2_X2 \AES_ENC/u0/u1/U391  ( .A1(\AES_ENC/u0/u1/n1093 ), .A2(\AES_ENC/u0/u1/n1045 ), .ZN(\AES_ENC/u0/u1/n701 ) );
NAND4_X2 \AES_ENC/u0/u1/U381  ( .A1(\AES_ENC/u0/u1/n702 ), .A2(\AES_ENC/u0/u1/n701 ), .A3(\AES_ENC/u0/u1/n700 ), .A4(\AES_ENC/u0/u1/n699 ), .ZN(\AES_ENC/u0/u1/n703 ) );
NAND2_X2 \AES_ENC/u0/u1/U380  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n703 ), .ZN(\AES_ENC/u0/u1/n732 ) );
AND2_X2 \AES_ENC/u0/u1/U379  ( .A1(\AES_ENC/w3[8] ), .A2(\AES_ENC/w3[14] ),.ZN(\AES_ENC/u0/u1/n1113 ) );
NAND2_X2 \AES_ENC/u0/u1/U378  ( .A1(\AES_ENC/u0/u1/n601 ), .A2(\AES_ENC/u0/u1/n1030 ), .ZN(\AES_ENC/u0/u1/n881 ) );
NAND2_X2 \AES_ENC/u0/u1/U377  ( .A1(\AES_ENC/u0/u1/n1093 ), .A2(\AES_ENC/u0/u1/n881 ), .ZN(\AES_ENC/u0/u1/n715 ) );
NAND2_X2 \AES_ENC/u0/u1/U376  ( .A1(\AES_ENC/u0/u1/n1010 ), .A2(\AES_ENC/u0/u1/n600 ), .ZN(\AES_ENC/u0/u1/n714 ) );
NAND2_X2 \AES_ENC/u0/u1/U375  ( .A1(\AES_ENC/u0/u1/n855 ), .A2(\AES_ENC/u0/u1/n588 ), .ZN(\AES_ENC/u0/u1/n1117 ) );
XNOR2_X2 \AES_ENC/u0/u1/U371  ( .A(\AES_ENC/u0/u1/n611 ), .B(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n824 ) );
NAND4_X2 \AES_ENC/u0/u1/U362  ( .A1(\AES_ENC/u0/u1/n715 ), .A2(\AES_ENC/u0/u1/n714 ), .A3(\AES_ENC/u0/u1/n713 ), .A4(\AES_ENC/u0/u1/n712 ), .ZN(\AES_ENC/u0/u1/n716 ) );
NAND2_X2 \AES_ENC/u0/u1/U361  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n716 ), .ZN(\AES_ENC/u0/u1/n731 ) );
AND2_X2 \AES_ENC/u0/u1/U360  ( .A1(\AES_ENC/w3[14] ), .A2(\AES_ENC/u0/u1/n574 ), .ZN(\AES_ENC/u0/u1/n1131 ) );
NAND2_X2 \AES_ENC/u0/u1/U359  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n717 ) );
NAND2_X2 \AES_ENC/u0/u1/U358  ( .A1(\AES_ENC/u0/u1/n1029 ), .A2(\AES_ENC/u0/u1/n717 ), .ZN(\AES_ENC/u0/u1/n728 ) );
NAND2_X2 \AES_ENC/u0/u1/U357  ( .A1(\AES_ENC/w3[9] ), .A2(\AES_ENC/u0/u1/n624 ), .ZN(\AES_ENC/u0/u1/n1097 ) );
NAND2_X2 \AES_ENC/u0/u1/U356  ( .A1(\AES_ENC/u0/u1/n603 ), .A2(\AES_ENC/u0/u1/n1097 ), .ZN(\AES_ENC/u0/u1/n718 ) );
NAND2_X2 \AES_ENC/u0/u1/U355  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n718 ), .ZN(\AES_ENC/u0/u1/n727 ) );
NAND4_X2 \AES_ENC/u0/u1/U344  ( .A1(\AES_ENC/u0/u1/n728 ), .A2(\AES_ENC/u0/u1/n727 ), .A3(\AES_ENC/u0/u1/n726 ), .A4(\AES_ENC/u0/u1/n725 ), .ZN(\AES_ENC/u0/u1/n729 ) );
NAND2_X2 \AES_ENC/u0/u1/U343  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n729 ), .ZN(\AES_ENC/u0/u1/n730 ) );
NAND4_X2 \AES_ENC/u0/u1/U342  ( .A1(\AES_ENC/u0/u1/n733 ), .A2(\AES_ENC/u0/u1/n732 ), .A3(\AES_ENC/u0/u1/n731 ), .A4(\AES_ENC/u0/u1/n730 ), .ZN(\AES_ENC/u0/subword[17] ) );
NAND2_X2 \AES_ENC/u0/u1/U341  ( .A1(\AES_ENC/w3[15] ), .A2(\AES_ENC/u0/u1/n611 ), .ZN(\AES_ENC/u0/u1/n734 ) );
NAND2_X2 \AES_ENC/u0/u1/U340  ( .A1(\AES_ENC/u0/u1/n734 ), .A2(\AES_ENC/u0/u1/n607 ), .ZN(\AES_ENC/u0/u1/n738 ) );
OR4_X2 \AES_ENC/u0/u1/U339  ( .A1(\AES_ENC/u0/u1/n738 ), .A2(\AES_ENC/u0/u1/n626 ), .A3(\AES_ENC/u0/u1/n826 ), .A4(\AES_ENC/u0/u1/n1121 ), .ZN(\AES_ENC/u0/u1/n746 ) );
NAND2_X2 \AES_ENC/u0/u1/U337  ( .A1(\AES_ENC/u0/u1/n1100 ), .A2(\AES_ENC/u0/u1/n587 ), .ZN(\AES_ENC/u0/u1/n992 ) );
OR2_X2 \AES_ENC/u0/u1/U336  ( .A1(\AES_ENC/u0/u1/n610 ), .A2(\AES_ENC/u0/u1/n735 ), .ZN(\AES_ENC/u0/u1/n737 ) );
NAND2_X2 \AES_ENC/u0/u1/U334  ( .A1(\AES_ENC/u0/u1/n619 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n753 ) );
NAND2_X2 \AES_ENC/u0/u1/U333  ( .A1(\AES_ENC/u0/u1/n582 ), .A2(\AES_ENC/u0/u1/n753 ), .ZN(\AES_ENC/u0/u1/n1080 ) );
NAND2_X2 \AES_ENC/u0/u1/U332  ( .A1(\AES_ENC/u0/u1/n1048 ), .A2(\AES_ENC/u0/u1/n576 ), .ZN(\AES_ENC/u0/u1/n736 ) );
NAND2_X2 \AES_ENC/u0/u1/U331  ( .A1(\AES_ENC/u0/u1/n737 ), .A2(\AES_ENC/u0/u1/n736 ), .ZN(\AES_ENC/u0/u1/n739 ) );
NAND2_X2 \AES_ENC/u0/u1/U330  ( .A1(\AES_ENC/u0/u1/n739 ), .A2(\AES_ENC/u0/u1/n738 ), .ZN(\AES_ENC/u0/u1/n745 ) );
NAND2_X2 \AES_ENC/u0/u1/U326  ( .A1(\AES_ENC/u0/u1/n1096 ), .A2(\AES_ENC/u0/u1/n590 ), .ZN(\AES_ENC/u0/u1/n906 ) );
NAND4_X2 \AES_ENC/u0/u1/U323  ( .A1(\AES_ENC/u0/u1/n746 ), .A2(\AES_ENC/u0/u1/n992 ), .A3(\AES_ENC/u0/u1/n745 ), .A4(\AES_ENC/u0/u1/n744 ), .ZN(\AES_ENC/u0/u1/n747 ) );
NAND2_X2 \AES_ENC/u0/u1/U322  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n747 ), .ZN(\AES_ENC/u0/u1/n793 ) );
NAND2_X2 \AES_ENC/u0/u1/U321  ( .A1(\AES_ENC/u0/u1/n584 ), .A2(\AES_ENC/u0/u1/n855 ), .ZN(\AES_ENC/u0/u1/n748 ) );
NAND2_X2 \AES_ENC/u0/u1/U320  ( .A1(\AES_ENC/u0/u1/n956 ), .A2(\AES_ENC/u0/u1/n748 ), .ZN(\AES_ENC/u0/u1/n760 ) );
NAND2_X2 \AES_ENC/u0/u1/U313  ( .A1(\AES_ENC/u0/u1/n590 ), .A2(\AES_ENC/u0/u1/n753 ), .ZN(\AES_ENC/u0/u1/n1023 ) );
NAND4_X2 \AES_ENC/u0/u1/U308  ( .A1(\AES_ENC/u0/u1/n760 ), .A2(\AES_ENC/u0/u1/n992 ), .A3(\AES_ENC/u0/u1/n759 ), .A4(\AES_ENC/u0/u1/n758 ), .ZN(\AES_ENC/u0/u1/n761 ) );
NAND2_X2 \AES_ENC/u0/u1/U307  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n761 ), .ZN(\AES_ENC/u0/u1/n792 ) );
NAND2_X2 \AES_ENC/u0/u1/U306  ( .A1(\AES_ENC/u0/u1/n584 ), .A2(\AES_ENC/u0/u1/n603 ), .ZN(\AES_ENC/u0/u1/n989 ) );
NAND2_X2 \AES_ENC/u0/u1/U305  ( .A1(\AES_ENC/u0/u1/n1050 ), .A2(\AES_ENC/u0/u1/n989 ), .ZN(\AES_ENC/u0/u1/n777 ) );
NAND2_X2 \AES_ENC/u0/u1/U304  ( .A1(\AES_ENC/u0/u1/n1093 ), .A2(\AES_ENC/u0/u1/n762 ), .ZN(\AES_ENC/u0/u1/n776 ) );
XNOR2_X2 \AES_ENC/u0/u1/U301  ( .A(\AES_ENC/w3[15] ), .B(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n959 ) );
NAND4_X2 \AES_ENC/u0/u1/U289  ( .A1(\AES_ENC/u0/u1/n777 ), .A2(\AES_ENC/u0/u1/n776 ), .A3(\AES_ENC/u0/u1/n775 ), .A4(\AES_ENC/u0/u1/n774 ), .ZN(\AES_ENC/u0/u1/n778 ) );
NAND2_X2 \AES_ENC/u0/u1/U288  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n778 ), .ZN(\AES_ENC/u0/u1/n791 ) );
NAND2_X2 \AES_ENC/u0/u1/U287  ( .A1(\AES_ENC/u0/u1/n1056 ), .A2(\AES_ENC/u0/u1/n1050 ), .ZN(\AES_ENC/u0/u1/n788 ) );
NAND2_X2 \AES_ENC/u0/u1/U286  ( .A1(\AES_ENC/u0/u1/n1091 ), .A2(\AES_ENC/u0/u1/n779 ), .ZN(\AES_ENC/u0/u1/n787 ) );
NAND2_X2 \AES_ENC/u0/u1/U285  ( .A1(\AES_ENC/u0/u1/n956 ), .A2(\AES_ENC/w3[9] ), .ZN(\AES_ENC/u0/u1/n786 ) );
NAND4_X2 \AES_ENC/u0/u1/U278  ( .A1(\AES_ENC/u0/u1/n788 ), .A2(\AES_ENC/u0/u1/n787 ), .A3(\AES_ENC/u0/u1/n786 ), .A4(\AES_ENC/u0/u1/n785 ), .ZN(\AES_ENC/u0/u1/n789 ) );
NAND2_X2 \AES_ENC/u0/u1/U277  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n789 ), .ZN(\AES_ENC/u0/u1/n790 ) );
NAND4_X2 \AES_ENC/u0/u1/U276  ( .A1(\AES_ENC/u0/u1/n793 ), .A2(\AES_ENC/u0/u1/n792 ), .A3(\AES_ENC/u0/u1/n791 ), .A4(\AES_ENC/u0/u1/n790 ), .ZN(\AES_ENC/u0/subword[18] ) );
NAND2_X2 \AES_ENC/u0/u1/U275  ( .A1(\AES_ENC/u0/u1/n1059 ), .A2(\AES_ENC/u0/u1/n794 ), .ZN(\AES_ENC/u0/u1/n810 ) );
NAND2_X2 \AES_ENC/u0/u1/U274  ( .A1(\AES_ENC/u0/u1/n1049 ), .A2(\AES_ENC/u0/u1/n956 ), .ZN(\AES_ENC/u0/u1/n809 ) );
OR2_X2 \AES_ENC/u0/u1/U266  ( .A1(\AES_ENC/u0/u1/n1096 ), .A2(\AES_ENC/u0/u1/n606 ), .ZN(\AES_ENC/u0/u1/n802 ) );
NAND2_X2 \AES_ENC/u0/u1/U265  ( .A1(\AES_ENC/u0/u1/n1053 ), .A2(\AES_ENC/u0/u1/n800 ), .ZN(\AES_ENC/u0/u1/n801 ) );
NAND2_X2 \AES_ENC/u0/u1/U264  ( .A1(\AES_ENC/u0/u1/n802 ), .A2(\AES_ENC/u0/u1/n801 ), .ZN(\AES_ENC/u0/u1/n805 ) );
NAND4_X2 \AES_ENC/u0/u1/U261  ( .A1(\AES_ENC/u0/u1/n810 ), .A2(\AES_ENC/u0/u1/n809 ), .A3(\AES_ENC/u0/u1/n808 ), .A4(\AES_ENC/u0/u1/n807 ), .ZN(\AES_ENC/u0/u1/n811 ) );
NAND2_X2 \AES_ENC/u0/u1/U260  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n811 ), .ZN(\AES_ENC/u0/u1/n852 ) );
OR2_X2 \AES_ENC/u0/u1/U259  ( .A1(\AES_ENC/u0/u1/n1023 ), .A2(\AES_ENC/u0/u1/n617 ), .ZN(\AES_ENC/u0/u1/n819 ) );
OR2_X2 \AES_ENC/u0/u1/U257  ( .A1(\AES_ENC/u0/u1/n570 ), .A2(\AES_ENC/u0/u1/n930 ), .ZN(\AES_ENC/u0/u1/n818 ) );
NAND2_X2 \AES_ENC/u0/u1/U256  ( .A1(\AES_ENC/u0/u1/n1013 ), .A2(\AES_ENC/u0/u1/n1094 ), .ZN(\AES_ENC/u0/u1/n817 ) );
NAND4_X2 \AES_ENC/u0/u1/U249  ( .A1(\AES_ENC/u0/u1/n819 ), .A2(\AES_ENC/u0/u1/n818 ), .A3(\AES_ENC/u0/u1/n817 ), .A4(\AES_ENC/u0/u1/n816 ), .ZN(\AES_ENC/u0/u1/n820 ) );
NAND2_X2 \AES_ENC/u0/u1/U248  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n820 ), .ZN(\AES_ENC/u0/u1/n851 ) );
NAND2_X2 \AES_ENC/u0/u1/U247  ( .A1(\AES_ENC/u0/u1/n956 ), .A2(\AES_ENC/u0/u1/n1080 ), .ZN(\AES_ENC/u0/u1/n835 ) );
NAND2_X2 \AES_ENC/u0/u1/U246  ( .A1(\AES_ENC/u0/u1/n570 ), .A2(\AES_ENC/u0/u1/n1030 ), .ZN(\AES_ENC/u0/u1/n1047 ) );
OR2_X2 \AES_ENC/u0/u1/U245  ( .A1(\AES_ENC/u0/u1/n1047 ), .A2(\AES_ENC/u0/u1/n612 ), .ZN(\AES_ENC/u0/u1/n834 ) );
NAND2_X2 \AES_ENC/u0/u1/U244  ( .A1(\AES_ENC/u0/u1/n1072 ), .A2(\AES_ENC/u0/u1/n589 ), .ZN(\AES_ENC/u0/u1/n833 ) );
NAND4_X2 \AES_ENC/u0/u1/U233  ( .A1(\AES_ENC/u0/u1/n835 ), .A2(\AES_ENC/u0/u1/n834 ), .A3(\AES_ENC/u0/u1/n833 ), .A4(\AES_ENC/u0/u1/n832 ), .ZN(\AES_ENC/u0/u1/n836 ) );
NAND2_X2 \AES_ENC/u0/u1/U232  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n836 ), .ZN(\AES_ENC/u0/u1/n850 ) );
NAND2_X2 \AES_ENC/u0/u1/U231  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n623 ), .ZN(\AES_ENC/u0/u1/n847 ) );
NAND2_X2 \AES_ENC/u0/u1/U230  ( .A1(\AES_ENC/u0/u1/n1050 ), .A2(\AES_ENC/u0/u1/n1071 ), .ZN(\AES_ENC/u0/u1/n846 ) );
OR2_X2 \AES_ENC/u0/u1/U224  ( .A1(\AES_ENC/u0/u1/n1053 ), .A2(\AES_ENC/u0/u1/n911 ), .ZN(\AES_ENC/u0/u1/n1077 ) );
NAND4_X2 \AES_ENC/u0/u1/U220  ( .A1(\AES_ENC/u0/u1/n847 ), .A2(\AES_ENC/u0/u1/n846 ), .A3(\AES_ENC/u0/u1/n845 ), .A4(\AES_ENC/u0/u1/n844 ), .ZN(\AES_ENC/u0/u1/n848 ) );
NAND2_X2 \AES_ENC/u0/u1/U219  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n848 ), .ZN(\AES_ENC/u0/u1/n849 ) );
NAND4_X2 \AES_ENC/u0/u1/U218  ( .A1(\AES_ENC/u0/u1/n852 ), .A2(\AES_ENC/u0/u1/n851 ), .A3(\AES_ENC/u0/u1/n850 ), .A4(\AES_ENC/u0/u1/n849 ), .ZN(\AES_ENC/u0/subword[19] ) );
NAND2_X2 \AES_ENC/u0/u1/U216  ( .A1(\AES_ENC/u0/u1/n1009 ), .A2(\AES_ENC/u0/u1/n1072 ), .ZN(\AES_ENC/u0/u1/n862 ) );
NAND2_X2 \AES_ENC/u0/u1/U215  ( .A1(\AES_ENC/u0/u1/n603 ), .A2(\AES_ENC/u0/u1/n577 ), .ZN(\AES_ENC/u0/u1/n853 ) );
NAND2_X2 \AES_ENC/u0/u1/U214  ( .A1(\AES_ENC/u0/u1/n1050 ), .A2(\AES_ENC/u0/u1/n853 ), .ZN(\AES_ENC/u0/u1/n861 ) );
NAND4_X2 \AES_ENC/u0/u1/U206  ( .A1(\AES_ENC/u0/u1/n862 ), .A2(\AES_ENC/u0/u1/n861 ), .A3(\AES_ENC/u0/u1/n860 ), .A4(\AES_ENC/u0/u1/n859 ), .ZN(\AES_ENC/u0/u1/n863 ) );
NAND2_X2 \AES_ENC/u0/u1/U205  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n863 ), .ZN(\AES_ENC/u0/u1/n905 ) );
NAND2_X2 \AES_ENC/u0/u1/U204  ( .A1(\AES_ENC/u0/u1/n1010 ), .A2(\AES_ENC/u0/u1/n989 ), .ZN(\AES_ENC/u0/u1/n874 ) );
NAND2_X2 \AES_ENC/u0/u1/U203  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n610 ), .ZN(\AES_ENC/u0/u1/n864 ) );
NAND2_X2 \AES_ENC/u0/u1/U202  ( .A1(\AES_ENC/u0/u1/n929 ), .A2(\AES_ENC/u0/u1/n864 ), .ZN(\AES_ENC/u0/u1/n873 ) );
NAND4_X2 \AES_ENC/u0/u1/U193  ( .A1(\AES_ENC/u0/u1/n874 ), .A2(\AES_ENC/u0/u1/n873 ), .A3(\AES_ENC/u0/u1/n872 ), .A4(\AES_ENC/u0/u1/n871 ), .ZN(\AES_ENC/u0/u1/n875 ) );
NAND2_X2 \AES_ENC/u0/u1/U192  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n875 ), .ZN(\AES_ENC/u0/u1/n904 ) );
NAND2_X2 \AES_ENC/u0/u1/U191  ( .A1(\AES_ENC/u0/u1/n583 ), .A2(\AES_ENC/u0/u1/n1050 ), .ZN(\AES_ENC/u0/u1/n889 ) );
NAND2_X2 \AES_ENC/u0/u1/U190  ( .A1(\AES_ENC/u0/u1/n1093 ), .A2(\AES_ENC/u0/u1/n587 ), .ZN(\AES_ENC/u0/u1/n876 ) );
NAND2_X2 \AES_ENC/u0/u1/U189  ( .A1(\AES_ENC/u0/u1/n604 ), .A2(\AES_ENC/u0/u1/n876 ), .ZN(\AES_ENC/u0/u1/n877 ) );
NAND2_X2 \AES_ENC/u0/u1/U188  ( .A1(\AES_ENC/u0/u1/n877 ), .A2(\AES_ENC/u0/u1/n623 ), .ZN(\AES_ENC/u0/u1/n888 ) );
NAND4_X2 \AES_ENC/u0/u1/U179  ( .A1(\AES_ENC/u0/u1/n889 ), .A2(\AES_ENC/u0/u1/n888 ), .A3(\AES_ENC/u0/u1/n887 ), .A4(\AES_ENC/u0/u1/n886 ), .ZN(\AES_ENC/u0/u1/n890 ) );
NAND2_X2 \AES_ENC/u0/u1/U178  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n890 ), .ZN(\AES_ENC/u0/u1/n903 ) );
OR2_X2 \AES_ENC/u0/u1/U177  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n1059 ), .ZN(\AES_ENC/u0/u1/n900 ) );
NAND2_X2 \AES_ENC/u0/u1/U176  ( .A1(\AES_ENC/u0/u1/n1073 ), .A2(\AES_ENC/u0/u1/n1047 ), .ZN(\AES_ENC/u0/u1/n899 ) );
NAND2_X2 \AES_ENC/u0/u1/U175  ( .A1(\AES_ENC/u0/u1/n1094 ), .A2(\AES_ENC/u0/u1/n595 ), .ZN(\AES_ENC/u0/u1/n898 ) );
NAND4_X2 \AES_ENC/u0/u1/U167  ( .A1(\AES_ENC/u0/u1/n900 ), .A2(\AES_ENC/u0/u1/n899 ), .A3(\AES_ENC/u0/u1/n898 ), .A4(\AES_ENC/u0/u1/n897 ), .ZN(\AES_ENC/u0/u1/n901 ) );
NAND2_X2 \AES_ENC/u0/u1/U166  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n901 ), .ZN(\AES_ENC/u0/u1/n902 ) );
NAND4_X2 \AES_ENC/u0/u1/U165  ( .A1(\AES_ENC/u0/u1/n905 ), .A2(\AES_ENC/u0/u1/n904 ), .A3(\AES_ENC/u0/u1/n903 ), .A4(\AES_ENC/u0/u1/n902 ), .ZN(\AES_ENC/u0/subword[20] ) );
NAND2_X2 \AES_ENC/u0/u1/U164  ( .A1(\AES_ENC/u0/u1/n1094 ), .A2(\AES_ENC/u0/u1/n599 ), .ZN(\AES_ENC/u0/u1/n922 ) );
NAND2_X2 \AES_ENC/u0/u1/U163  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n989 ), .ZN(\AES_ENC/u0/u1/n921 ) );
NAND4_X2 \AES_ENC/u0/u1/U151  ( .A1(\AES_ENC/u0/u1/n922 ), .A2(\AES_ENC/u0/u1/n921 ), .A3(\AES_ENC/u0/u1/n920 ), .A4(\AES_ENC/u0/u1/n919 ), .ZN(\AES_ENC/u0/u1/n923 ) );
NAND2_X2 \AES_ENC/u0/u1/U150  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n923 ), .ZN(\AES_ENC/u0/u1/n972 ) );
NAND2_X2 \AES_ENC/u0/u1/U149  ( .A1(\AES_ENC/u0/u1/n582 ), .A2(\AES_ENC/u0/u1/n619 ), .ZN(\AES_ENC/u0/u1/n924 ) );
NAND2_X2 \AES_ENC/u0/u1/U148  ( .A1(\AES_ENC/u0/u1/n1073 ), .A2(\AES_ENC/u0/u1/n924 ), .ZN(\AES_ENC/u0/u1/n939 ) );
NAND2_X2 \AES_ENC/u0/u1/U147  ( .A1(\AES_ENC/u0/u1/n926 ), .A2(\AES_ENC/u0/u1/n925 ), .ZN(\AES_ENC/u0/u1/n927 ) );
NAND2_X2 \AES_ENC/u0/u1/U146  ( .A1(\AES_ENC/u0/u1/n606 ), .A2(\AES_ENC/u0/u1/n927 ), .ZN(\AES_ENC/u0/u1/n928 ) );
NAND2_X2 \AES_ENC/u0/u1/U145  ( .A1(\AES_ENC/u0/u1/n928 ), .A2(\AES_ENC/u0/u1/n1080 ), .ZN(\AES_ENC/u0/u1/n938 ) );
OR2_X2 \AES_ENC/u0/u1/U144  ( .A1(\AES_ENC/u0/u1/n1117 ), .A2(\AES_ENC/u0/u1/n615 ), .ZN(\AES_ENC/u0/u1/n937 ) );
NAND4_X2 \AES_ENC/u0/u1/U139  ( .A1(\AES_ENC/u0/u1/n939 ), .A2(\AES_ENC/u0/u1/n938 ), .A3(\AES_ENC/u0/u1/n937 ), .A4(\AES_ENC/u0/u1/n936 ), .ZN(\AES_ENC/u0/u1/n940 ) );
NAND2_X2 \AES_ENC/u0/u1/U138  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n940 ), .ZN(\AES_ENC/u0/u1/n971 ) );
OR2_X2 \AES_ENC/u0/u1/U137  ( .A1(\AES_ENC/u0/u1/n605 ), .A2(\AES_ENC/u0/u1/n941 ), .ZN(\AES_ENC/u0/u1/n954 ) );
NAND2_X2 \AES_ENC/u0/u1/U136  ( .A1(\AES_ENC/u0/u1/n1096 ), .A2(\AES_ENC/u0/u1/n577 ), .ZN(\AES_ENC/u0/u1/n942 ) );
NAND2_X2 \AES_ENC/u0/u1/U135  ( .A1(\AES_ENC/u0/u1/n1048 ), .A2(\AES_ENC/u0/u1/n942 ), .ZN(\AES_ENC/u0/u1/n943 ) );
NAND2_X2 \AES_ENC/u0/u1/U134  ( .A1(\AES_ENC/u0/u1/n612 ), .A2(\AES_ENC/u0/u1/n943 ), .ZN(\AES_ENC/u0/u1/n944 ) );
NAND2_X2 \AES_ENC/u0/u1/U133  ( .A1(\AES_ENC/u0/u1/n944 ), .A2(\AES_ENC/u0/u1/n580 ), .ZN(\AES_ENC/u0/u1/n953 ) );
NAND4_X2 \AES_ENC/u0/u1/U125  ( .A1(\AES_ENC/u0/u1/n954 ), .A2(\AES_ENC/u0/u1/n953 ), .A3(\AES_ENC/u0/u1/n952 ), .A4(\AES_ENC/u0/u1/n951 ), .ZN(\AES_ENC/u0/u1/n955 ) );
NAND2_X2 \AES_ENC/u0/u1/U124  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n955 ), .ZN(\AES_ENC/u0/u1/n970 ) );
NAND2_X2 \AES_ENC/u0/u1/U123  ( .A1(\AES_ENC/u0/u1/n1094 ), .A2(\AES_ENC/u0/u1/n1071 ), .ZN(\AES_ENC/u0/u1/n967 ) );
NAND2_X2 \AES_ENC/u0/u1/U122  ( .A1(\AES_ENC/u0/u1/n956 ), .A2(\AES_ENC/u0/u1/n1030 ), .ZN(\AES_ENC/u0/u1/n966 ) );
NAND4_X2 \AES_ENC/u0/u1/U114  ( .A1(\AES_ENC/u0/u1/n967 ), .A2(\AES_ENC/u0/u1/n966 ), .A3(\AES_ENC/u0/u1/n965 ), .A4(\AES_ENC/u0/u1/n964 ), .ZN(\AES_ENC/u0/u1/n968 ) );
NAND2_X2 \AES_ENC/u0/u1/U113  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n968 ), .ZN(\AES_ENC/u0/u1/n969 ) );
NAND4_X2 \AES_ENC/u0/u1/U112  ( .A1(\AES_ENC/u0/u1/n972 ), .A2(\AES_ENC/u0/u1/n971 ), .A3(\AES_ENC/u0/u1/n970 ), .A4(\AES_ENC/u0/u1/n969 ), .ZN(\AES_ENC/u0/subword[21] ) );
NAND2_X2 \AES_ENC/u0/u1/U111  ( .A1(\AES_ENC/u0/u1/n570 ), .A2(\AES_ENC/u0/u1/n1097 ), .ZN(\AES_ENC/u0/u1/n973 ) );
NAND2_X2 \AES_ENC/u0/u1/U110  ( .A1(\AES_ENC/u0/u1/n1073 ), .A2(\AES_ENC/u0/u1/n973 ), .ZN(\AES_ENC/u0/u1/n987 ) );
NAND2_X2 \AES_ENC/u0/u1/U109  ( .A1(\AES_ENC/u0/u1/n974 ), .A2(\AES_ENC/u0/u1/n1077 ), .ZN(\AES_ENC/u0/u1/n975 ) );
NAND2_X2 \AES_ENC/u0/u1/U108  ( .A1(\AES_ENC/u0/u1/n613 ), .A2(\AES_ENC/u0/u1/n975 ), .ZN(\AES_ENC/u0/u1/n976 ) );
NAND2_X2 \AES_ENC/u0/u1/U107  ( .A1(\AES_ENC/u0/u1/n977 ), .A2(\AES_ENC/u0/u1/n976 ), .ZN(\AES_ENC/u0/u1/n986 ) );
NAND4_X2 \AES_ENC/u0/u1/U99  ( .A1(\AES_ENC/u0/u1/n987 ), .A2(\AES_ENC/u0/u1/n986 ), .A3(\AES_ENC/u0/u1/n985 ), .A4(\AES_ENC/u0/u1/n984 ), .ZN(\AES_ENC/u0/u1/n988 ) );
NAND2_X2 \AES_ENC/u0/u1/U98  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n988 ), .ZN(\AES_ENC/u0/u1/n1044 ) );
NAND2_X2 \AES_ENC/u0/u1/U97  ( .A1(\AES_ENC/u0/u1/n1073 ), .A2(\AES_ENC/u0/u1/n989 ), .ZN(\AES_ENC/u0/u1/n1004 ) );
NAND2_X2 \AES_ENC/u0/u1/U96  ( .A1(\AES_ENC/u0/u1/n1092 ), .A2(\AES_ENC/u0/u1/n619 ), .ZN(\AES_ENC/u0/u1/n1003 ) );
NAND4_X2 \AES_ENC/u0/u1/U85  ( .A1(\AES_ENC/u0/u1/n1004 ), .A2(\AES_ENC/u0/u1/n1003 ), .A3(\AES_ENC/u0/u1/n1002 ), .A4(\AES_ENC/u0/u1/n1001 ), .ZN(\AES_ENC/u0/u1/n1005 ) );
NAND2_X2 \AES_ENC/u0/u1/U84  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n1005 ), .ZN(\AES_ENC/u0/u1/n1043 ) );
NAND2_X2 \AES_ENC/u0/u1/U83  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n596 ), .ZN(\AES_ENC/u0/u1/n1020 ) );
NAND2_X2 \AES_ENC/u0/u1/U82  ( .A1(\AES_ENC/u0/u1/n1050 ), .A2(\AES_ENC/u0/u1/n624 ), .ZN(\AES_ENC/u0/u1/n1019 ) );
NAND2_X2 \AES_ENC/u0/u1/U77  ( .A1(\AES_ENC/u0/u1/n1059 ), .A2(\AES_ENC/u0/u1/n1114 ), .ZN(\AES_ENC/u0/u1/n1012 ) );
NAND2_X2 \AES_ENC/u0/u1/U76  ( .A1(\AES_ENC/u0/u1/n1010 ), .A2(\AES_ENC/u0/u1/n592 ), .ZN(\AES_ENC/u0/u1/n1011 ) );
NAND2_X2 \AES_ENC/u0/u1/U75  ( .A1(\AES_ENC/u0/u1/n1012 ), .A2(\AES_ENC/u0/u1/n1011 ), .ZN(\AES_ENC/u0/u1/n1016 ) );
NAND4_X2 \AES_ENC/u0/u1/U70  ( .A1(\AES_ENC/u0/u1/n1020 ), .A2(\AES_ENC/u0/u1/n1019 ), .A3(\AES_ENC/u0/u1/n1018 ), .A4(\AES_ENC/u0/u1/n1017 ), .ZN(\AES_ENC/u0/u1/n1021 ) );
NAND2_X2 \AES_ENC/u0/u1/U69  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n1021 ), .ZN(\AES_ENC/u0/u1/n1042 ) );
NAND2_X2 \AES_ENC/u0/u1/U68  ( .A1(\AES_ENC/u0/u1/n1022 ), .A2(\AES_ENC/u0/u1/n1093 ), .ZN(\AES_ENC/u0/u1/n1039 ) );
NAND2_X2 \AES_ENC/u0/u1/U67  ( .A1(\AES_ENC/u0/u1/n1050 ), .A2(\AES_ENC/u0/u1/n1023 ), .ZN(\AES_ENC/u0/u1/n1038 ) );
NAND2_X2 \AES_ENC/u0/u1/U66  ( .A1(\AES_ENC/u0/u1/n1024 ), .A2(\AES_ENC/u0/u1/n1071 ), .ZN(\AES_ENC/u0/u1/n1037 ) );
AND2_X2 \AES_ENC/u0/u1/U60  ( .A1(\AES_ENC/u0/u1/n1030 ), .A2(\AES_ENC/u0/u1/n602 ), .ZN(\AES_ENC/u0/u1/n1078 ) );
NAND4_X2 \AES_ENC/u0/u1/U56  ( .A1(\AES_ENC/u0/u1/n1039 ), .A2(\AES_ENC/u0/u1/n1038 ), .A3(\AES_ENC/u0/u1/n1037 ), .A4(\AES_ENC/u0/u1/n1036 ), .ZN(\AES_ENC/u0/u1/n1040 ) );
NAND2_X2 \AES_ENC/u0/u1/U55  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n1040 ), .ZN(\AES_ENC/u0/u1/n1041 ) );
NAND4_X2 \AES_ENC/u0/u1/U54  ( .A1(\AES_ENC/u0/u1/n1044 ), .A2(\AES_ENC/u0/u1/n1043 ), .A3(\AES_ENC/u0/u1/n1042 ), .A4(\AES_ENC/u0/u1/n1041 ), .ZN(\AES_ENC/u0/subword[22] ) );
NAND2_X2 \AES_ENC/u0/u1/U53  ( .A1(\AES_ENC/u0/u1/n1072 ), .A2(\AES_ENC/u0/u1/n1045 ), .ZN(\AES_ENC/u0/u1/n1068 ) );
NAND2_X2 \AES_ENC/u0/u1/U52  ( .A1(\AES_ENC/u0/u1/n1046 ), .A2(\AES_ENC/u0/u1/n582 ), .ZN(\AES_ENC/u0/u1/n1067 ) );
NAND2_X2 \AES_ENC/u0/u1/U51  ( .A1(\AES_ENC/u0/u1/n1094 ), .A2(\AES_ENC/u0/u1/n1047 ), .ZN(\AES_ENC/u0/u1/n1066 ) );
NAND4_X2 \AES_ENC/u0/u1/U40  ( .A1(\AES_ENC/u0/u1/n1068 ), .A2(\AES_ENC/u0/u1/n1067 ), .A3(\AES_ENC/u0/u1/n1066 ), .A4(\AES_ENC/u0/u1/n1065 ), .ZN(\AES_ENC/u0/u1/n1069 ) );
NAND2_X2 \AES_ENC/u0/u1/U39  ( .A1(\AES_ENC/u0/u1/n1070 ), .A2(\AES_ENC/u0/u1/n1069 ), .ZN(\AES_ENC/u0/u1/n1135 ) );
NAND2_X2 \AES_ENC/u0/u1/U38  ( .A1(\AES_ENC/u0/u1/n1072 ), .A2(\AES_ENC/u0/u1/n1071 ), .ZN(\AES_ENC/u0/u1/n1088 ) );
NAND2_X2 \AES_ENC/u0/u1/U37  ( .A1(\AES_ENC/u0/u1/n1073 ), .A2(\AES_ENC/u0/u1/n595 ), .ZN(\AES_ENC/u0/u1/n1087 ) );
NAND4_X2 \AES_ENC/u0/u1/U28  ( .A1(\AES_ENC/u0/u1/n1088 ), .A2(\AES_ENC/u0/u1/n1087 ), .A3(\AES_ENC/u0/u1/n1086 ), .A4(\AES_ENC/u0/u1/n1085 ), .ZN(\AES_ENC/u0/u1/n1089 ) );
NAND2_X2 \AES_ENC/u0/u1/U27  ( .A1(\AES_ENC/u0/u1/n1090 ), .A2(\AES_ENC/u0/u1/n1089 ), .ZN(\AES_ENC/u0/u1/n1134 ) );
NAND2_X2 \AES_ENC/u0/u1/U26  ( .A1(\AES_ENC/u0/u1/n1091 ), .A2(\AES_ENC/u0/u1/n1093 ), .ZN(\AES_ENC/u0/u1/n1111 ) );
NAND2_X2 \AES_ENC/u0/u1/U25  ( .A1(\AES_ENC/u0/u1/n1092 ), .A2(\AES_ENC/u0/u1/n1120 ), .ZN(\AES_ENC/u0/u1/n1110 ) );
AND2_X2 \AES_ENC/u0/u1/U22  ( .A1(\AES_ENC/u0/u1/n1097 ), .A2(\AES_ENC/u0/u1/n1096 ), .ZN(\AES_ENC/u0/u1/n1098 ) );
NAND4_X2 \AES_ENC/u0/u1/U14  ( .A1(\AES_ENC/u0/u1/n1111 ), .A2(\AES_ENC/u0/u1/n1110 ), .A3(\AES_ENC/u0/u1/n1109 ), .A4(\AES_ENC/u0/u1/n1108 ), .ZN(\AES_ENC/u0/u1/n1112 ) );
NAND2_X2 \AES_ENC/u0/u1/U13  ( .A1(\AES_ENC/u0/u1/n1113 ), .A2(\AES_ENC/u0/u1/n1112 ), .ZN(\AES_ENC/u0/u1/n1133 ) );
NAND2_X2 \AES_ENC/u0/u1/U12  ( .A1(\AES_ENC/u0/u1/n1115 ), .A2(\AES_ENC/u0/u1/n1114 ), .ZN(\AES_ENC/u0/u1/n1129 ) );
OR2_X2 \AES_ENC/u0/u1/U11  ( .A1(\AES_ENC/u0/u1/n608 ), .A2(\AES_ENC/u0/u1/n1116 ), .ZN(\AES_ENC/u0/u1/n1128 ) );
NAND4_X2 \AES_ENC/u0/u1/U3  ( .A1(\AES_ENC/u0/u1/n1129 ), .A2(\AES_ENC/u0/u1/n1128 ), .A3(\AES_ENC/u0/u1/n1127 ), .A4(\AES_ENC/u0/u1/n1126 ), .ZN(\AES_ENC/u0/u1/n1130 ) );
NAND2_X2 \AES_ENC/u0/u1/U2  ( .A1(\AES_ENC/u0/u1/n1131 ), .A2(\AES_ENC/u0/u1/n1130 ), .ZN(\AES_ENC/u0/u1/n1132 ) );
NAND4_X2 \AES_ENC/u0/u1/U1  ( .A1(\AES_ENC/u0/u1/n1135 ), .A2(\AES_ENC/u0/u1/n1134 ), .A3(\AES_ENC/u0/u1/n1133 ), .A4(\AES_ENC/u0/u1/n1132 ), .ZN(\AES_ENC/u0/subword[23] ) );
INV_X4 \AES_ENC/u0/u2/U575  ( .A(\AES_ENC/w3[7] ), .ZN(\AES_ENC/u0/u2/n627 ));
INV_X4 \AES_ENC/u0/u2/U574  ( .A(\AES_ENC/u0/u2/n1114 ), .ZN(\AES_ENC/u0/u2/n625 ) );
INV_X4 \AES_ENC/u0/u2/U573  ( .A(\AES_ENC/w3[4] ), .ZN(\AES_ENC/u0/u2/n624 ));
INV_X4 \AES_ENC/u0/u2/U572  ( .A(\AES_ENC/u0/u2/n1025 ), .ZN(\AES_ENC/u0/u2/n622 ) );
INV_X4 \AES_ENC/u0/u2/U571  ( .A(\AES_ENC/u0/u2/n1120 ), .ZN(\AES_ENC/u0/u2/n620 ) );
INV_X4 \AES_ENC/u0/u2/U570  ( .A(\AES_ENC/u0/u2/n1121 ), .ZN(\AES_ENC/u0/u2/n619 ) );
INV_X4 \AES_ENC/u0/u2/U569  ( .A(\AES_ENC/u0/u2/n1048 ), .ZN(\AES_ENC/u0/u2/n618 ) );
INV_X4 \AES_ENC/u0/u2/U568  ( .A(\AES_ENC/u0/u2/n974 ), .ZN(\AES_ENC/u0/u2/n616 ) );
INV_X4 \AES_ENC/u0/u2/U567  ( .A(\AES_ENC/u0/u2/n794 ), .ZN(\AES_ENC/u0/u2/n614 ) );
INV_X4 \AES_ENC/u0/u2/U566  ( .A(\AES_ENC/w3[2] ), .ZN(\AES_ENC/u0/u2/n611 ));
INV_X4 \AES_ENC/u0/u2/U565  ( .A(\AES_ENC/u0/u2/n800 ), .ZN(\AES_ENC/u0/u2/n610 ) );
INV_X4 \AES_ENC/u0/u2/U564  ( .A(\AES_ENC/u0/u2/n925 ), .ZN(\AES_ENC/u0/u2/n609 ) );
INV_X4 \AES_ENC/u0/u2/U563  ( .A(\AES_ENC/u0/u2/n779 ), .ZN(\AES_ENC/u0/u2/n607 ) );
INV_X4 \AES_ENC/u0/u2/U562  ( .A(\AES_ENC/u0/u2/n1022 ), .ZN(\AES_ENC/u0/u2/n603 ) );
INV_X4 \AES_ENC/u0/u2/U561  ( .A(\AES_ENC/u0/u2/n1102 ), .ZN(\AES_ENC/u0/u2/n602 ) );
INV_X4 \AES_ENC/u0/u2/U560  ( .A(\AES_ENC/u0/u2/n929 ), .ZN(\AES_ENC/u0/u2/n601 ) );
INV_X4 \AES_ENC/u0/u2/U559  ( .A(\AES_ENC/u0/u2/n1056 ), .ZN(\AES_ENC/u0/u2/n600 ) );
INV_X4 \AES_ENC/u0/u2/U558  ( .A(\AES_ENC/u0/u2/n1054 ), .ZN(\AES_ENC/u0/u2/n599 ) );
INV_X4 \AES_ENC/u0/u2/U557  ( .A(\AES_ENC/u0/u2/n881 ), .ZN(\AES_ENC/u0/u2/n598 ) );
INV_X4 \AES_ENC/u0/u2/U556  ( .A(\AES_ENC/u0/u2/n926 ), .ZN(\AES_ENC/u0/u2/n597 ) );
INV_X4 \AES_ENC/u0/u2/U555  ( .A(\AES_ENC/u0/u2/n977 ), .ZN(\AES_ENC/u0/u2/n595 ) );
INV_X4 \AES_ENC/u0/u2/U554  ( .A(\AES_ENC/u0/u2/n1031 ), .ZN(\AES_ENC/u0/u2/n594 ) );
INV_X4 \AES_ENC/u0/u2/U553  ( .A(\AES_ENC/u0/u2/n1103 ), .ZN(\AES_ENC/u0/u2/n593 ) );
INV_X4 \AES_ENC/u0/u2/U552  ( .A(\AES_ENC/u0/u2/n1009 ), .ZN(\AES_ENC/u0/u2/n592 ) );
INV_X4 \AES_ENC/u0/u2/U551  ( .A(\AES_ENC/u0/u2/n990 ), .ZN(\AES_ENC/u0/u2/n591 ) );
INV_X4 \AES_ENC/u0/u2/U550  ( .A(\AES_ENC/u0/u2/n1058 ), .ZN(\AES_ENC/u0/u2/n590 ) );
INV_X4 \AES_ENC/u0/u2/U549  ( .A(\AES_ENC/u0/u2/n1074 ), .ZN(\AES_ENC/u0/u2/n589 ) );
INV_X4 \AES_ENC/u0/u2/U548  ( .A(\AES_ENC/u0/u2/n1053 ), .ZN(\AES_ENC/u0/u2/n588 ) );
INV_X4 \AES_ENC/u0/u2/U547  ( .A(\AES_ENC/u0/u2/n826 ), .ZN(\AES_ENC/u0/u2/n587 ) );
INV_X4 \AES_ENC/u0/u2/U546  ( .A(\AES_ENC/u0/u2/n992 ), .ZN(\AES_ENC/u0/u2/n586 ) );
INV_X4 \AES_ENC/u0/u2/U545  ( .A(\AES_ENC/u0/u2/n821 ), .ZN(\AES_ENC/u0/u2/n585 ) );
INV_X4 \AES_ENC/u0/u2/U544  ( .A(\AES_ENC/u0/u2/n910 ), .ZN(\AES_ENC/u0/u2/n584 ) );
INV_X4 \AES_ENC/u0/u2/U543  ( .A(\AES_ENC/u0/u2/n906 ), .ZN(\AES_ENC/u0/u2/n583 ) );
INV_X4 \AES_ENC/u0/u2/U542  ( .A(\AES_ENC/u0/u2/n880 ), .ZN(\AES_ENC/u0/u2/n581 ) );
INV_X4 \AES_ENC/u0/u2/U541  ( .A(\AES_ENC/u0/u2/n1013 ), .ZN(\AES_ENC/u0/u2/n580 ) );
INV_X4 \AES_ENC/u0/u2/U540  ( .A(\AES_ENC/u0/u2/n1092 ), .ZN(\AES_ENC/u0/u2/n579 ) );
INV_X4 \AES_ENC/u0/u2/U539  ( .A(\AES_ENC/u0/u2/n824 ), .ZN(\AES_ENC/u0/u2/n578 ) );
INV_X4 \AES_ENC/u0/u2/U538  ( .A(\AES_ENC/u0/u2/n1091 ), .ZN(\AES_ENC/u0/u2/n577 ) );
INV_X4 \AES_ENC/u0/u2/U537  ( .A(\AES_ENC/u0/u2/n1080 ), .ZN(\AES_ENC/u0/u2/n576 ) );
INV_X4 \AES_ENC/u0/u2/U536  ( .A(\AES_ENC/u0/u2/n959 ), .ZN(\AES_ENC/u0/u2/n575 ) );
INV_X4 \AES_ENC/u0/u2/U535  ( .A(\AES_ENC/w3[0] ), .ZN(\AES_ENC/u0/u2/n574 ));
NOR2_X2 \AES_ENC/u0/u2/U534  ( .A1(\AES_ENC/u0/u2/n574 ), .A2(\AES_ENC/w3[6] ), .ZN(\AES_ENC/u0/u2/n1070 ) );
NOR2_X2 \AES_ENC/u0/u2/U533  ( .A1(\AES_ENC/w3[0] ), .A2(\AES_ENC/w3[6] ),.ZN(\AES_ENC/u0/u2/n1090 ) );
NOR2_X2 \AES_ENC/u0/u2/U532  ( .A1(\AES_ENC/w3[4] ), .A2(\AES_ENC/w3[3] ),.ZN(\AES_ENC/u0/u2/n1025 ) );
NAND3_X2 \AES_ENC/u0/u2/U531  ( .A1(\AES_ENC/u0/u2/n679 ), .A2(\AES_ENC/u0/u2/n678 ), .A3(\AES_ENC/u0/u2/n677 ), .ZN(\AES_ENC/u0/subword[8] ) );
NOR2_X2 \AES_ENC/u0/u2/U530  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n765 ) );
NOR2_X2 \AES_ENC/u0/u2/U529  ( .A1(\AES_ENC/w3[4] ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n764 ) );
NOR2_X2 \AES_ENC/u0/u2/U528  ( .A1(\AES_ENC/u0/u2/n765 ), .A2(\AES_ENC/u0/u2/n764 ), .ZN(\AES_ENC/u0/u2/n766 ) );
NOR2_X2 \AES_ENC/u0/u2/U527  ( .A1(\AES_ENC/u0/u2/n766 ), .A2(\AES_ENC/u0/u2/n575 ), .ZN(\AES_ENC/u0/u2/n767 ) );
NOR2_X2 \AES_ENC/u0/u2/U526  ( .A1(\AES_ENC/u0/u2/n1117 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n707 ) );
NOR3_X2 \AES_ENC/u0/u2/U525  ( .A1(\AES_ENC/u0/u2/n627 ), .A2(\AES_ENC/w3[5] ), .A3(\AES_ENC/u0/u2/n704 ), .ZN(\AES_ENC/u0/u2/n706 ));
NOR2_X2 \AES_ENC/u0/u2/U524  ( .A1(\AES_ENC/w3[4] ), .A2(\AES_ENC/u0/u2/n579 ), .ZN(\AES_ENC/u0/u2/n705 ) );
NOR3_X2 \AES_ENC/u0/u2/U523  ( .A1(\AES_ENC/u0/u2/n707 ), .A2(\AES_ENC/u0/u2/n706 ), .A3(\AES_ENC/u0/u2/n705 ), .ZN(\AES_ENC/u0/u2/n713 ) );
NOR4_X2 \AES_ENC/u0/u2/U522  ( .A1(\AES_ENC/u0/u2/n633 ), .A2(\AES_ENC/u0/u2/n632 ), .A3(\AES_ENC/u0/u2/n631 ), .A4(\AES_ENC/u0/u2/n630 ), .ZN(\AES_ENC/u0/u2/n634 ) );
NOR2_X2 \AES_ENC/u0/u2/U521  ( .A1(\AES_ENC/u0/u2/n629 ), .A2(\AES_ENC/u0/u2/n628 ), .ZN(\AES_ENC/u0/u2/n635 ) );
NAND3_X2 \AES_ENC/u0/u2/U520  ( .A1(\AES_ENC/w3[2] ), .A2(\AES_ENC/w3[7] ),.A3(\AES_ENC/u0/u2/n1059 ), .ZN(\AES_ENC/u0/u2/n636 ) );
INV_X4 \AES_ENC/u0/u2/U519  ( .A(\AES_ENC/w3[3] ), .ZN(\AES_ENC/u0/u2/n621 ));
NOR2_X2 \AES_ENC/u0/u2/U518  ( .A1(\AES_ENC/w3[5] ), .A2(\AES_ENC/w3[2] ),.ZN(\AES_ENC/u0/u2/n974 ) );
NAND3_X2 \AES_ENC/u0/u2/U517  ( .A1(\AES_ENC/u0/u2/n652 ), .A2(\AES_ENC/u0/u2/n626 ), .A3(\AES_ENC/w3[7] ), .ZN(\AES_ENC/u0/u2/n653 ));
NOR2_X2 \AES_ENC/u0/u2/U516  ( .A1(\AES_ENC/u0/u2/n611 ), .A2(\AES_ENC/w3[5] ), .ZN(\AES_ENC/u0/u2/n925 ) );
NOR2_X2 \AES_ENC/u0/u2/U515  ( .A1(\AES_ENC/u0/u2/n626 ), .A2(\AES_ENC/w3[2] ), .ZN(\AES_ENC/u0/u2/n1048 ) );
INV_X4 \AES_ENC/u0/u2/U512  ( .A(\AES_ENC/w3[5] ), .ZN(\AES_ENC/u0/u2/n626 ));
NOR2_X2 \AES_ENC/u0/u2/U510  ( .A1(\AES_ENC/u0/u2/n611 ), .A2(\AES_ENC/w3[7] ), .ZN(\AES_ENC/u0/u2/n779 ) );
NOR2_X2 \AES_ENC/u0/u2/U509  ( .A1(\AES_ENC/w3[7] ), .A2(\AES_ENC/w3[2] ),.ZN(\AES_ENC/u0/u2/n794 ) );
NOR2_X2 \AES_ENC/u0/u2/U508  ( .A1(\AES_ENC/w3[4] ), .A2(\AES_ENC/w3[1] ),.ZN(\AES_ENC/u0/u2/n1102 ) );
INV_X4 \AES_ENC/u0/u2/U507  ( .A(\AES_ENC/u0/u2/n569 ), .ZN(\AES_ENC/u0/u2/n572 ) );
NOR2_X2 \AES_ENC/u0/u2/U506  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/w3[3] ), .ZN(\AES_ENC/u0/u2/n1053 ) );
NOR2_X2 \AES_ENC/u0/u2/U505  ( .A1(\AES_ENC/u0/u2/n607 ), .A2(\AES_ENC/w3[5] ), .ZN(\AES_ENC/u0/u2/n1024 ) );
NOR2_X2 \AES_ENC/u0/u2/U504  ( .A1(\AES_ENC/u0/u2/n625 ), .A2(\AES_ENC/w3[2] ), .ZN(\AES_ENC/u0/u2/n1093 ) );
NOR2_X2 \AES_ENC/u0/u2/U503  ( .A1(\AES_ENC/u0/u2/n614 ), .A2(\AES_ENC/w3[5] ), .ZN(\AES_ENC/u0/u2/n1094 ) );
NOR2_X2 \AES_ENC/u0/u2/U502  ( .A1(\AES_ENC/u0/u2/n624 ), .A2(\AES_ENC/w3[3] ), .ZN(\AES_ENC/u0/u2/n931 ) );
INV_X4 \AES_ENC/u0/u2/U501  ( .A(\AES_ENC/u0/u2/n570 ), .ZN(\AES_ENC/u0/u2/n573 ) );
NOR2_X2 \AES_ENC/u0/u2/U500  ( .A1(\AES_ENC/u0/u2/n622 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n1059 ) );
NOR2_X2 \AES_ENC/u0/u2/U499  ( .A1(\AES_ENC/u0/u2/n1053 ), .A2(\AES_ENC/u0/u2/n1095 ), .ZN(\AES_ENC/u0/u2/n639 ) );
NOR3_X2 \AES_ENC/u0/u2/U498  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n573 ), .A3(\AES_ENC/u0/u2/n1074 ), .ZN(\AES_ENC/u0/u2/n641 ) );
NOR2_X2 \AES_ENC/u0/u2/U497  ( .A1(\AES_ENC/u0/u2/n639 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n640 ) );
NOR2_X2 \AES_ENC/u0/u2/U496  ( .A1(\AES_ENC/u0/u2/n641 ), .A2(\AES_ENC/u0/u2/n640 ), .ZN(\AES_ENC/u0/u2/n646 ) );
NOR2_X2 \AES_ENC/u0/u2/U495  ( .A1(\AES_ENC/u0/u2/n826 ), .A2(\AES_ENC/u0/u2/n572 ), .ZN(\AES_ENC/u0/u2/n827 ) );
NOR3_X2 \AES_ENC/u0/u2/U494  ( .A1(\AES_ENC/u0/u2/n769 ), .A2(\AES_ENC/u0/u2/n768 ), .A3(\AES_ENC/u0/u2/n767 ), .ZN(\AES_ENC/u0/u2/n775 ) );
NOR2_X2 \AES_ENC/u0/u2/U492  ( .A1(\AES_ENC/w3[1] ), .A2(\AES_ENC/u0/u2/n623 ), .ZN(\AES_ENC/u0/u2/n913 ) );
NOR2_X2 \AES_ENC/u0/u2/U491  ( .A1(\AES_ENC/u0/u2/n913 ), .A2(\AES_ENC/u0/u2/n1091 ), .ZN(\AES_ENC/u0/u2/n914 ) );
NOR2_X2 \AES_ENC/u0/u2/U490  ( .A1(\AES_ENC/u0/u2/n1056 ), .A2(\AES_ENC/u0/u2/n1053 ), .ZN(\AES_ENC/u0/u2/n749 ) );
NOR2_X2 \AES_ENC/u0/u2/U489  ( .A1(\AES_ENC/u0/u2/n749 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n752 ) );
NOR3_X2 \AES_ENC/u0/u2/U488  ( .A1(\AES_ENC/u0/u2/n995 ), .A2(\AES_ENC/u0/u2/n586 ), .A3(\AES_ENC/u0/u2/n994 ), .ZN(\AES_ENC/u0/u2/n1002 ) );
NOR2_X2 \AES_ENC/u0/u2/U487  ( .A1(\AES_ENC/u0/u2/n909 ), .A2(\AES_ENC/u0/u2/n908 ), .ZN(\AES_ENC/u0/u2/n920 ) );
INV_X4 \AES_ENC/u0/u2/U486  ( .A(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n596 ));
NOR2_X2 \AES_ENC/u0/u2/U483  ( .A1(\AES_ENC/u0/u2/n932 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n933 ) );
NOR2_X2 \AES_ENC/u0/u2/U482  ( .A1(\AES_ENC/u0/u2/n929 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n935 ) );
NOR2_X2 \AES_ENC/u0/u2/U480  ( .A1(\AES_ENC/u0/u2/n931 ), .A2(\AES_ENC/u0/u2/n930 ), .ZN(\AES_ENC/u0/u2/n934 ) );
NOR3_X2 \AES_ENC/u0/u2/U479  ( .A1(\AES_ENC/u0/u2/n935 ), .A2(\AES_ENC/u0/u2/n934 ), .A3(\AES_ENC/u0/u2/n933 ), .ZN(\AES_ENC/u0/u2/n936 ) );
OR2_X4 \AES_ENC/u0/u2/U478  ( .A1(\AES_ENC/u0/u2/n1094 ), .A2(\AES_ENC/u0/u2/n1093 ), .ZN(\AES_ENC/u0/u2/n571 ) );
AND2_X2 \AES_ENC/u0/u2/U477  ( .A1(\AES_ENC/u0/u2/n571 ), .A2(\AES_ENC/u0/u2/n1095 ), .ZN(\AES_ENC/u0/u2/n1101 ) );
NOR2_X2 \AES_ENC/u0/u2/U474  ( .A1(\AES_ENC/u0/u2/n1074 ), .A2(\AES_ENC/u0/u2/n931 ), .ZN(\AES_ENC/u0/u2/n796 ) );
NOR2_X2 \AES_ENC/u0/u2/U473  ( .A1(\AES_ENC/u0/u2/n796 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n797 ) );
NOR2_X2 \AES_ENC/u0/u2/U472  ( .A1(\AES_ENC/u0/u2/n1054 ), .A2(\AES_ENC/u0/u2/n1053 ), .ZN(\AES_ENC/u0/u2/n1055 ) );
NOR2_X2 \AES_ENC/u0/u2/U471  ( .A1(\AES_ENC/u0/u2/n572 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n949 ) );
NOR2_X2 \AES_ENC/u0/u2/U470  ( .A1(\AES_ENC/u0/u2/n1049 ), .A2(\AES_ENC/u0/u2/n618 ), .ZN(\AES_ENC/u0/u2/n1051 ) );
NOR2_X2 \AES_ENC/u0/u2/U469  ( .A1(\AES_ENC/u0/u2/n1051 ), .A2(\AES_ENC/u0/u2/n1050 ), .ZN(\AES_ENC/u0/u2/n1052 ) );
NOR2_X2 \AES_ENC/u0/u2/U468  ( .A1(\AES_ENC/u0/u2/n1052 ), .A2(\AES_ENC/u0/u2/n592 ), .ZN(\AES_ENC/u0/u2/n1064 ) );
NOR2_X2 \AES_ENC/u0/u2/U467  ( .A1(\AES_ENC/w3[1] ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n631 ) );
NOR2_X2 \AES_ENC/u0/u2/U466  ( .A1(\AES_ENC/u0/u2/n1025 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n980 ) );
NOR2_X2 \AES_ENC/u0/u2/U465  ( .A1(\AES_ENC/u0/u2/n1074 ), .A2(\AES_ENC/u0/u2/n1025 ), .ZN(\AES_ENC/u0/u2/n891 ) );
NOR2_X2 \AES_ENC/u0/u2/U464  ( .A1(\AES_ENC/u0/u2/n891 ), .A2(\AES_ENC/u0/u2/n609 ), .ZN(\AES_ENC/u0/u2/n894 ) );
NOR2_X2 \AES_ENC/u0/u2/U463  ( .A1(\AES_ENC/u0/u2/n1073 ), .A2(\AES_ENC/u0/u2/n1094 ), .ZN(\AES_ENC/u0/u2/n795 ) );
NOR2_X2 \AES_ENC/u0/u2/U462  ( .A1(\AES_ENC/u0/u2/n795 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n799 ) );
NOR2_X2 \AES_ENC/u0/u2/U461  ( .A1(\AES_ENC/u0/u2/n624 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n1075 ) );
NOR2_X2 \AES_ENC/u0/u2/U460  ( .A1(\AES_ENC/u0/u2/n624 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n822 ) );
NOR2_X2 \AES_ENC/u0/u2/U459  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n823 ) );
NOR2_X2 \AES_ENC/u0/u2/U458  ( .A1(\AES_ENC/u0/u2/n823 ), .A2(\AES_ENC/u0/u2/n822 ), .ZN(\AES_ENC/u0/u2/n825 ) );
NOR2_X2 \AES_ENC/u0/u2/U455  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n981 ) );
NOR2_X2 \AES_ENC/u0/u2/U448  ( .A1(\AES_ENC/u0/u2/n1102 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n643 ) );
NOR2_X2 \AES_ENC/u0/u2/U447  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n621 ), .ZN(\AES_ENC/u0/u2/n642 ) );
NOR2_X2 \AES_ENC/u0/u2/U442  ( .A1(\AES_ENC/u0/u2/n911 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n644 ) );
NOR4_X2 \AES_ENC/u0/u2/U441  ( .A1(\AES_ENC/u0/u2/n644 ), .A2(\AES_ENC/u0/u2/n643 ), .A3(\AES_ENC/u0/u2/n804 ), .A4(\AES_ENC/u0/u2/n642 ), .ZN(\AES_ENC/u0/u2/n645 ) );
NOR2_X2 \AES_ENC/u0/u2/U438  ( .A1(\AES_ENC/u0/u2/n1102 ), .A2(\AES_ENC/u0/u2/n910 ), .ZN(\AES_ENC/u0/u2/n932 ) );
NOR3_X2 \AES_ENC/u0/u2/U435  ( .A1(\AES_ENC/u0/u2/n623 ), .A2(\AES_ENC/w3[1] ), .A3(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n683 ));
NOR2_X2 \AES_ENC/u0/u2/U434  ( .A1(\AES_ENC/u0/u2/n1102 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n755 ) );
INV_X4 \AES_ENC/u0/u2/U433  ( .A(\AES_ENC/u0/u2/n931 ), .ZN(\AES_ENC/u0/u2/n623 ) );
NOR2_X2 \AES_ENC/u0/u2/U428  ( .A1(\AES_ENC/u0/u2/n996 ), .A2(\AES_ENC/u0/u2/n931 ), .ZN(\AES_ENC/u0/u2/n704 ) );
NOR2_X2 \AES_ENC/u0/u2/U427  ( .A1(\AES_ENC/u0/u2/n1029 ), .A2(\AES_ENC/u0/u2/n1025 ), .ZN(\AES_ENC/u0/u2/n1079 ) );
NOR3_X2 \AES_ENC/u0/u2/U421  ( .A1(\AES_ENC/u0/u2/n589 ), .A2(\AES_ENC/u0/u2/n1025 ), .A3(\AES_ENC/u0/u2/n616 ), .ZN(\AES_ENC/u0/u2/n945 ) );
NOR2_X2 \AES_ENC/u0/u2/U420  ( .A1(\AES_ENC/u0/u2/n1072 ), .A2(\AES_ENC/u0/u2/n1094 ), .ZN(\AES_ENC/u0/u2/n930 ) );
NOR2_X2 \AES_ENC/u0/u2/U419  ( .A1(\AES_ENC/u0/u2/n931 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n743 ) );
NOR2_X2 \AES_ENC/u0/u2/U418  ( .A1(\AES_ENC/u0/u2/n931 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n685 ) );
NOR3_X2 \AES_ENC/u0/u2/U417  ( .A1(\AES_ENC/u0/u2/n610 ), .A2(\AES_ENC/u0/u2/n572 ), .A3(\AES_ENC/u0/u2/n575 ), .ZN(\AES_ENC/u0/u2/n962 ) );
NOR2_X2 \AES_ENC/u0/u2/U416  ( .A1(\AES_ENC/u0/u2/n626 ), .A2(\AES_ENC/u0/u2/n611 ), .ZN(\AES_ENC/u0/u2/n800 ) );
NOR3_X2 \AES_ENC/u0/u2/U415  ( .A1(\AES_ENC/u0/u2/n590 ), .A2(\AES_ENC/u0/u2/n627 ), .A3(\AES_ENC/u0/u2/n611 ), .ZN(\AES_ENC/u0/u2/n798 ) );
NOR3_X2 \AES_ENC/u0/u2/U414  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n572 ), .A3(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n694 ) );
NOR3_X2 \AES_ENC/u0/u2/U413  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n572 ), .A3(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n895 ) );
NOR3_X2 \AES_ENC/u0/u2/U410  ( .A1(\AES_ENC/u0/u2/n1008 ), .A2(\AES_ENC/u0/u2/n1007 ), .A3(\AES_ENC/u0/u2/n1006 ), .ZN(\AES_ENC/u0/u2/n1018 ) );
NOR4_X2 \AES_ENC/u0/u2/U409  ( .A1(\AES_ENC/u0/u2/n806 ), .A2(\AES_ENC/u0/u2/n805 ), .A3(\AES_ENC/u0/u2/n804 ), .A4(\AES_ENC/u0/u2/n803 ), .ZN(\AES_ENC/u0/u2/n807 ) );
NOR3_X2 \AES_ENC/u0/u2/U406  ( .A1(\AES_ENC/u0/u2/n799 ), .A2(\AES_ENC/u0/u2/n798 ), .A3(\AES_ENC/u0/u2/n797 ), .ZN(\AES_ENC/u0/u2/n808 ) );
NOR2_X2 \AES_ENC/u0/u2/U405  ( .A1(\AES_ENC/u0/u2/n669 ), .A2(\AES_ENC/u0/u2/n668 ), .ZN(\AES_ENC/u0/u2/n673 ) );
NOR4_X2 \AES_ENC/u0/u2/U404  ( .A1(\AES_ENC/u0/u2/n946 ), .A2(\AES_ENC/u0/u2/n1046 ), .A3(\AES_ENC/u0/u2/n671 ), .A4(\AES_ENC/u0/u2/n670 ), .ZN(\AES_ENC/u0/u2/n672 ) );
NOR4_X2 \AES_ENC/u0/u2/U403  ( .A1(\AES_ENC/u0/u2/n711 ), .A2(\AES_ENC/u0/u2/n710 ), .A3(\AES_ENC/u0/u2/n709 ), .A4(\AES_ENC/u0/u2/n708 ), .ZN(\AES_ENC/u0/u2/n712 ) );
NOR4_X2 \AES_ENC/u0/u2/U401  ( .A1(\AES_ENC/u0/u2/n843 ), .A2(\AES_ENC/u0/u2/n842 ), .A3(\AES_ENC/u0/u2/n841 ), .A4(\AES_ENC/u0/u2/n840 ), .ZN(\AES_ENC/u0/u2/n844 ) );
NOR3_X2 \AES_ENC/u0/u2/U400  ( .A1(\AES_ENC/u0/u2/n1101 ), .A2(\AES_ENC/u0/u2/n1100 ), .A3(\AES_ENC/u0/u2/n1099 ), .ZN(\AES_ENC/u0/u2/n1109 ) );
NOR3_X2 \AES_ENC/u0/u2/U399  ( .A1(\AES_ENC/u0/u2/n743 ), .A2(\AES_ENC/u0/u2/n742 ), .A3(\AES_ENC/u0/u2/n741 ), .ZN(\AES_ENC/u0/u2/n744 ) );
NOR2_X2 \AES_ENC/u0/u2/U398  ( .A1(\AES_ENC/u0/u2/n697 ), .A2(\AES_ENC/u0/u2/n658 ), .ZN(\AES_ENC/u0/u2/n659 ) );
NOR3_X2 \AES_ENC/u0/u2/U397  ( .A1(\AES_ENC/u0/u2/n959 ), .A2(\AES_ENC/u0/u2/n572 ), .A3(\AES_ENC/u0/u2/n609 ), .ZN(\AES_ENC/u0/u2/n768 ) );
NOR2_X2 \AES_ENC/u0/u2/U396  ( .A1(\AES_ENC/u0/u2/n1078 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n1033 ) );
NOR2_X2 \AES_ENC/u0/u2/U393  ( .A1(\AES_ENC/u0/u2/n1031 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n1032 ) );
NOR3_X2 \AES_ENC/u0/u2/U390  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n1025 ), .A3(\AES_ENC/u0/u2/n1074 ), .ZN(\AES_ENC/u0/u2/n1035 ) );
NOR4_X2 \AES_ENC/u0/u2/U389  ( .A1(\AES_ENC/u0/u2/n1035 ), .A2(\AES_ENC/u0/u2/n1034 ), .A3(\AES_ENC/u0/u2/n1033 ), .A4(\AES_ENC/u0/u2/n1032 ), .ZN(\AES_ENC/u0/u2/n1036 ) );
NOR2_X2 \AES_ENC/u0/u2/U388  ( .A1(\AES_ENC/u0/u2/n598 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n885 ) );
NOR2_X2 \AES_ENC/u0/u2/U387  ( .A1(\AES_ENC/u0/u2/n623 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n882 ) );
NOR2_X2 \AES_ENC/u0/u2/U386  ( .A1(\AES_ENC/u0/u2/n1053 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n884 ) );
NOR4_X2 \AES_ENC/u0/u2/U385  ( .A1(\AES_ENC/u0/u2/n885 ), .A2(\AES_ENC/u0/u2/n884 ), .A3(\AES_ENC/u0/u2/n883 ), .A4(\AES_ENC/u0/u2/n882 ), .ZN(\AES_ENC/u0/u2/n886 ) );
NOR2_X2 \AES_ENC/u0/u2/U384  ( .A1(\AES_ENC/u0/u2/n825 ), .A2(\AES_ENC/u0/u2/n578 ), .ZN(\AES_ENC/u0/u2/n830 ) );
NOR2_X2 \AES_ENC/u0/u2/U383  ( .A1(\AES_ENC/u0/u2/n827 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n829 ) );
NOR2_X2 \AES_ENC/u0/u2/U382  ( .A1(\AES_ENC/u0/u2/n572 ), .A2(\AES_ENC/u0/u2/n579 ), .ZN(\AES_ENC/u0/u2/n828 ) );
NOR4_X2 \AES_ENC/u0/u2/U374  ( .A1(\AES_ENC/u0/u2/n831 ), .A2(\AES_ENC/u0/u2/n830 ), .A3(\AES_ENC/u0/u2/n829 ), .A4(\AES_ENC/u0/u2/n828 ), .ZN(\AES_ENC/u0/u2/n832 ) );
NOR2_X2 \AES_ENC/u0/u2/U373  ( .A1(\AES_ENC/u0/u2/n598 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n1107 ) );
NOR2_X2 \AES_ENC/u0/u2/U372  ( .A1(\AES_ENC/u0/u2/n1102 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n1106 ) );
NOR2_X2 \AES_ENC/u0/u2/U370  ( .A1(\AES_ENC/u0/u2/n1103 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n1105 ) );
NOR4_X2 \AES_ENC/u0/u2/U369  ( .A1(\AES_ENC/u0/u2/n1107 ), .A2(\AES_ENC/u0/u2/n1106 ), .A3(\AES_ENC/u0/u2/n1105 ), .A4(\AES_ENC/u0/u2/n1104 ), .ZN(\AES_ENC/u0/u2/n1108 ) );
NOR3_X2 \AES_ENC/u0/u2/U368  ( .A1(\AES_ENC/u0/u2/n959 ), .A2(\AES_ENC/u0/u2/n621 ), .A3(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n963 ) );
NOR2_X2 \AES_ENC/u0/u2/U367  ( .A1(\AES_ENC/u0/u2/n626 ), .A2(\AES_ENC/u0/u2/n627 ), .ZN(\AES_ENC/u0/u2/n1114 ) );
NOR3_X2 \AES_ENC/u0/u2/U366  ( .A1(\AES_ENC/u0/u2/n910 ), .A2(\AES_ENC/u0/u2/n1059 ), .A3(\AES_ENC/u0/u2/n611 ), .ZN(\AES_ENC/u0/u2/n1115 ) );
INV_X4 \AES_ENC/u0/u2/U365  ( .A(\AES_ENC/u0/u2/n1024 ), .ZN(\AES_ENC/u0/u2/n606 ) );
INV_X4 \AES_ENC/u0/u2/U364  ( .A(\AES_ENC/u0/u2/n1094 ), .ZN(\AES_ENC/u0/u2/n613 ) );
NOR2_X2 \AES_ENC/u0/u2/U363  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n931 ), .ZN(\AES_ENC/u0/u2/n1100 ) );
NOR2_X2 \AES_ENC/u0/u2/U354  ( .A1(\AES_ENC/u0/u2/n569 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n929 ) );
NOR2_X2 \AES_ENC/u0/u2/U353  ( .A1(\AES_ENC/u0/u2/n620 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n926 ) );
INV_X4 \AES_ENC/u0/u2/U352  ( .A(\AES_ENC/u0/u2/n1093 ), .ZN(\AES_ENC/u0/u2/n617 ) );
NOR2_X2 \AES_ENC/u0/u2/U351  ( .A1(\AES_ENC/u0/u2/n572 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n1095 ) );
NOR2_X2 \AES_ENC/u0/u2/U350  ( .A1(\AES_ENC/u0/u2/n609 ), .A2(\AES_ENC/u0/u2/n627 ), .ZN(\AES_ENC/u0/u2/n1010 ) );
NOR2_X2 \AES_ENC/u0/u2/U349  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n1103 ) );
NOR2_X2 \AES_ENC/u0/u2/U348  ( .A1(\AES_ENC/w3[1] ), .A2(\AES_ENC/u0/u2/n1120 ), .ZN(\AES_ENC/u0/u2/n1022 ) );
NOR2_X2 \AES_ENC/u0/u2/U347  ( .A1(\AES_ENC/u0/u2/n619 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n911 ) );
NOR2_X2 \AES_ENC/u0/u2/U346  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/u0/u2/n1025 ), .ZN(\AES_ENC/u0/u2/n826 ) );
NOR2_X2 \AES_ENC/u0/u2/U345  ( .A1(\AES_ENC/u0/u2/n626 ), .A2(\AES_ENC/u0/u2/n607 ), .ZN(\AES_ENC/u0/u2/n1072 ) );
NOR2_X2 \AES_ENC/u0/u2/U338  ( .A1(\AES_ENC/u0/u2/n627 ), .A2(\AES_ENC/u0/u2/n616 ), .ZN(\AES_ENC/u0/u2/n956 ) );
NOR2_X2 \AES_ENC/u0/u2/U335  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/u0/u2/n624 ), .ZN(\AES_ENC/u0/u2/n1121 ) );
NOR2_X2 \AES_ENC/u0/u2/U329  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/u0/u2/n624 ), .ZN(\AES_ENC/u0/u2/n1058 ) );
NOR2_X2 \AES_ENC/u0/u2/U328  ( .A1(\AES_ENC/u0/u2/n625 ), .A2(\AES_ENC/u0/u2/n611 ), .ZN(\AES_ENC/u0/u2/n1073 ) );
NOR2_X2 \AES_ENC/u0/u2/U327  ( .A1(\AES_ENC/w3[1] ), .A2(\AES_ENC/u0/u2/n1025 ), .ZN(\AES_ENC/u0/u2/n1054 ) );
NOR2_X2 \AES_ENC/u0/u2/U325  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/u0/u2/n931 ), .ZN(\AES_ENC/u0/u2/n1029 ) );
NOR2_X2 \AES_ENC/u0/u2/U324  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n1056 ) );
NOR2_X2 \AES_ENC/u0/u2/U319  ( .A1(\AES_ENC/u0/u2/n614 ), .A2(\AES_ENC/u0/u2/n626 ), .ZN(\AES_ENC/u0/u2/n1050 ) );
NOR2_X2 \AES_ENC/u0/u2/U318  ( .A1(\AES_ENC/u0/u2/n1121 ), .A2(\AES_ENC/u0/u2/n1025 ), .ZN(\AES_ENC/u0/u2/n1120 ) );
NOR2_X2 \AES_ENC/u0/u2/U317  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/u0/u2/n572 ), .ZN(\AES_ENC/u0/u2/n1074 ) );
NOR2_X2 \AES_ENC/u0/u2/U316  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n584 ), .ZN(\AES_ENC/u0/u2/n838 ) );
NOR2_X2 \AES_ENC/u0/u2/U315  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n602 ), .ZN(\AES_ENC/u0/u2/n837 ) );
NOR2_X2 \AES_ENC/u0/u2/U314  ( .A1(\AES_ENC/u0/u2/n838 ), .A2(\AES_ENC/u0/u2/n837 ), .ZN(\AES_ENC/u0/u2/n845 ) );
NOR2_X2 \AES_ENC/u0/u2/U312  ( .A1(\AES_ENC/u0/u2/n1058 ), .A2(\AES_ENC/u0/u2/n1054 ), .ZN(\AES_ENC/u0/u2/n878 ) );
NOR2_X2 \AES_ENC/u0/u2/U311  ( .A1(\AES_ENC/u0/u2/n878 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n879 ) );
NOR2_X2 \AES_ENC/u0/u2/U310  ( .A1(\AES_ENC/u0/u2/n880 ), .A2(\AES_ENC/u0/u2/n879 ), .ZN(\AES_ENC/u0/u2/n887 ) );
NOR3_X2 \AES_ENC/u0/u2/U309  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n1091 ), .A3(\AES_ENC/u0/u2/n1022 ), .ZN(\AES_ENC/u0/u2/n720 ) );
NOR3_X2 \AES_ENC/u0/u2/U303  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n1054 ), .A3(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n719 ) );
NOR2_X2 \AES_ENC/u0/u2/U302  ( .A1(\AES_ENC/u0/u2/n720 ), .A2(\AES_ENC/u0/u2/n719 ), .ZN(\AES_ENC/u0/u2/n726 ) );
NOR2_X2 \AES_ENC/u0/u2/U300  ( .A1(\AES_ENC/u0/u2/n614 ), .A2(\AES_ENC/u0/u2/n591 ), .ZN(\AES_ENC/u0/u2/n865 ) );
NOR2_X2 \AES_ENC/u0/u2/U299  ( .A1(\AES_ENC/u0/u2/n1059 ), .A2(\AES_ENC/u0/u2/n1058 ), .ZN(\AES_ENC/u0/u2/n1060 ) );
NOR2_X2 \AES_ENC/u0/u2/U298  ( .A1(\AES_ENC/u0/u2/n1095 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n668 ) );
NOR2_X2 \AES_ENC/u0/u2/U297  ( .A1(\AES_ENC/u0/u2/n826 ), .A2(\AES_ENC/u0/u2/n573 ), .ZN(\AES_ENC/u0/u2/n750 ) );
NOR2_X2 \AES_ENC/u0/u2/U296  ( .A1(\AES_ENC/u0/u2/n750 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n751 ) );
NOR2_X2 \AES_ENC/u0/u2/U295  ( .A1(\AES_ENC/u0/u2/n907 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n908 ) );
NOR2_X2 \AES_ENC/u0/u2/U294  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n588 ), .ZN(\AES_ENC/u0/u2/n957 ) );
NOR2_X2 \AES_ENC/u0/u2/U293  ( .A1(\AES_ENC/u0/u2/n990 ), .A2(\AES_ENC/u0/u2/n926 ), .ZN(\AES_ENC/u0/u2/n780 ) );
NOR2_X2 \AES_ENC/u0/u2/U292  ( .A1(\AES_ENC/u0/u2/n1022 ), .A2(\AES_ENC/u0/u2/n1058 ), .ZN(\AES_ENC/u0/u2/n740 ) );
NOR2_X2 \AES_ENC/u0/u2/U291  ( .A1(\AES_ENC/u0/u2/n740 ), .A2(\AES_ENC/u0/u2/n616 ), .ZN(\AES_ENC/u0/u2/n742 ) );
NOR2_X2 \AES_ENC/u0/u2/U290  ( .A1(\AES_ENC/u0/u2/n1098 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n1099 ) );
NOR2_X2 \AES_ENC/u0/u2/U284  ( .A1(\AES_ENC/u0/u2/n1120 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n993 ) );
NOR2_X2 \AES_ENC/u0/u2/U283  ( .A1(\AES_ENC/u0/u2/n993 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n994 ) );
NOR2_X2 \AES_ENC/u0/u2/U282  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n620 ), .ZN(\AES_ENC/u0/u2/n1026 ) );
NOR2_X2 \AES_ENC/u0/u2/U281  ( .A1(\AES_ENC/u0/u2/n573 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n1027 ) );
NOR2_X2 \AES_ENC/u0/u2/U280  ( .A1(\AES_ENC/u0/u2/n1027 ), .A2(\AES_ENC/u0/u2/n1026 ), .ZN(\AES_ENC/u0/u2/n1028 ) );
NOR2_X2 \AES_ENC/u0/u2/U279  ( .A1(\AES_ENC/u0/u2/n1029 ), .A2(\AES_ENC/u0/u2/n1028 ), .ZN(\AES_ENC/u0/u2/n1034 ) );
NOR2_X2 \AES_ENC/u0/u2/U273  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n1071 ), .ZN(\AES_ENC/u0/u2/n669 ) );
NOR2_X2 \AES_ENC/u0/u2/U272  ( .A1(\AES_ENC/u0/u2/n1056 ), .A2(\AES_ENC/u0/u2/n990 ), .ZN(\AES_ENC/u0/u2/n991 ) );
NOR2_X2 \AES_ENC/u0/u2/U271  ( .A1(\AES_ENC/u0/u2/n991 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n995 ) );
NOR4_X2 \AES_ENC/u0/u2/U270  ( .A1(\AES_ENC/u0/u2/n757 ), .A2(\AES_ENC/u0/u2/n756 ), .A3(\AES_ENC/u0/u2/n755 ), .A4(\AES_ENC/u0/u2/n754 ), .ZN(\AES_ENC/u0/u2/n758 ) );
NOR2_X2 \AES_ENC/u0/u2/U269  ( .A1(\AES_ENC/u0/u2/n752 ), .A2(\AES_ENC/u0/u2/n751 ), .ZN(\AES_ENC/u0/u2/n759 ) );
NOR2_X2 \AES_ENC/u0/u2/U268  ( .A1(\AES_ENC/u0/u2/n607 ), .A2(\AES_ENC/u0/u2/n590 ), .ZN(\AES_ENC/u0/u2/n1008 ) );
NOR2_X2 \AES_ENC/u0/u2/U267  ( .A1(\AES_ENC/u0/u2/n606 ), .A2(\AES_ENC/u0/u2/n906 ), .ZN(\AES_ENC/u0/u2/n741 ) );
NOR2_X2 \AES_ENC/u0/u2/U263  ( .A1(\AES_ENC/u0/u2/n1054 ), .A2(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n763 ) );
NOR2_X2 \AES_ENC/u0/u2/U262  ( .A1(\AES_ENC/u0/u2/n763 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n769 ) );
NOR2_X2 \AES_ENC/u0/u2/U258  ( .A1(\AES_ENC/u0/u2/n839 ), .A2(\AES_ENC/u0/u2/n582 ), .ZN(\AES_ENC/u0/u2/n693 ) );
NOR2_X2 \AES_ENC/u0/u2/U255  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n577 ), .ZN(\AES_ENC/u0/u2/n1007 ) );
NOR2_X2 \AES_ENC/u0/u2/U254  ( .A1(\AES_ENC/u0/u2/n609 ), .A2(\AES_ENC/u0/u2/n580 ), .ZN(\AES_ENC/u0/u2/n1123 ) );
NOR2_X2 \AES_ENC/u0/u2/U253  ( .A1(\AES_ENC/u0/u2/n780 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n784 ) );
NOR2_X2 \AES_ENC/u0/u2/U252  ( .A1(\AES_ENC/u0/u2/n1117 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n782 ) );
NOR2_X2 \AES_ENC/u0/u2/U251  ( .A1(\AES_ENC/u0/u2/n781 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n783 ) );
NOR4_X2 \AES_ENC/u0/u2/U250  ( .A1(\AES_ENC/u0/u2/n880 ), .A2(\AES_ENC/u0/u2/n784 ), .A3(\AES_ENC/u0/u2/n783 ), .A4(\AES_ENC/u0/u2/n782 ), .ZN(\AES_ENC/u0/u2/n785 ) );
NOR2_X2 \AES_ENC/u0/u2/U243  ( .A1(\AES_ENC/u0/u2/n609 ), .A2(\AES_ENC/u0/u2/n590 ), .ZN(\AES_ENC/u0/u2/n710 ) );
INV_X4 \AES_ENC/u0/u2/U242  ( .A(\AES_ENC/u0/u2/n1029 ), .ZN(\AES_ENC/u0/u2/n582 ) );
NOR2_X2 \AES_ENC/u0/u2/U241  ( .A1(\AES_ENC/u0/u2/n593 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n1125 ) );
NOR2_X2 \AES_ENC/u0/u2/U240  ( .A1(\AES_ENC/u0/u2/n616 ), .A2(\AES_ENC/u0/u2/n580 ), .ZN(\AES_ENC/u0/u2/n771 ) );
NOR2_X2 \AES_ENC/u0/u2/U239  ( .A1(\AES_ENC/u0/u2/n616 ), .A2(\AES_ENC/u0/u2/n597 ), .ZN(\AES_ENC/u0/u2/n883 ) );
NOR2_X2 \AES_ENC/u0/u2/U238  ( .A1(\AES_ENC/u0/u2/n911 ), .A2(\AES_ENC/u0/u2/n910 ), .ZN(\AES_ENC/u0/u2/n912 ) );
NOR2_X2 \AES_ENC/u0/u2/U237  ( .A1(\AES_ENC/u0/u2/n912 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n916 ) );
NOR2_X2 \AES_ENC/u0/u2/U236  ( .A1(\AES_ENC/u0/u2/n990 ), .A2(\AES_ENC/u0/u2/n929 ), .ZN(\AES_ENC/u0/u2/n892 ) );
NOR2_X2 \AES_ENC/u0/u2/U235  ( .A1(\AES_ENC/u0/u2/n892 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n893 ) );
NOR2_X2 \AES_ENC/u0/u2/U234  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n602 ), .ZN(\AES_ENC/u0/u2/n950 ) );
NOR2_X2 \AES_ENC/u0/u2/U229  ( .A1(\AES_ENC/u0/u2/n1079 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n1082 ) );
NOR2_X2 \AES_ENC/u0/u2/U228  ( .A1(\AES_ENC/u0/u2/n910 ), .A2(\AES_ENC/u0/u2/n1056 ), .ZN(\AES_ENC/u0/u2/n941 ) );
NOR2_X2 \AES_ENC/u0/u2/U227  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n1077 ), .ZN(\AES_ENC/u0/u2/n841 ) );
NOR2_X2 \AES_ENC/u0/u2/U226  ( .A1(\AES_ENC/u0/u2/n623 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n630 ) );
NOR2_X2 \AES_ENC/u0/u2/U225  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n602 ), .ZN(\AES_ENC/u0/u2/n806 ) );
NOR2_X2 \AES_ENC/u0/u2/U223  ( .A1(\AES_ENC/u0/u2/n623 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n948 ) );
NOR2_X2 \AES_ENC/u0/u2/U222  ( .A1(\AES_ENC/u0/u2/n606 ), .A2(\AES_ENC/u0/u2/n582 ), .ZN(\AES_ENC/u0/u2/n1104 ) );
NOR2_X2 \AES_ENC/u0/u2/U221  ( .A1(\AES_ENC/u0/u2/n1121 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n1122 ) );
NOR2_X2 \AES_ENC/u0/u2/U217  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n1023 ), .ZN(\AES_ENC/u0/u2/n756 ) );
NOR2_X2 \AES_ENC/u0/u2/U213  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n602 ), .ZN(\AES_ENC/u0/u2/n870 ) );
NOR2_X2 \AES_ENC/u0/u2/U212  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n569 ), .ZN(\AES_ENC/u0/u2/n947 ) );
NOR2_X2 \AES_ENC/u0/u2/U211  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n1077 ), .ZN(\AES_ENC/u0/u2/n1084 ) );
NOR2_X2 \AES_ENC/u0/u2/U210  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n855 ), .ZN(\AES_ENC/u0/u2/n709 ) );
NOR2_X2 \AES_ENC/u0/u2/U209  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n589 ), .ZN(\AES_ENC/u0/u2/n868 ) );
NOR2_X2 \AES_ENC/u0/u2/U208  ( .A1(\AES_ENC/u0/u2/n1120 ), .A2(\AES_ENC/u0/u2/n839 ), .ZN(\AES_ENC/u0/u2/n842 ) );
NOR2_X2 \AES_ENC/u0/u2/U207  ( .A1(\AES_ENC/u0/u2/n1120 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n1124 ) );
NOR2_X2 \AES_ENC/u0/u2/U201  ( .A1(\AES_ENC/u0/u2/n1120 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n696 ) );
NOR2_X2 \AES_ENC/u0/u2/U200  ( .A1(\AES_ENC/u0/u2/n1074 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n1076 ) );
NOR2_X2 \AES_ENC/u0/u2/U199  ( .A1(\AES_ENC/u0/u2/n1074 ), .A2(\AES_ENC/u0/u2/n620 ), .ZN(\AES_ENC/u0/u2/n781 ) );
NOR3_X2 \AES_ENC/u0/u2/U198  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n1056 ), .A3(\AES_ENC/u0/u2/n990 ), .ZN(\AES_ENC/u0/u2/n979 ) );
NOR3_X2 \AES_ENC/u0/u2/U197  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n1058 ), .A3(\AES_ENC/u0/u2/n1059 ), .ZN(\AES_ENC/u0/u2/n854 ) );
NOR2_X2 \AES_ENC/u0/u2/U196  ( .A1(\AES_ENC/u0/u2/n996 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n869 ) );
NOR2_X2 \AES_ENC/u0/u2/U195  ( .A1(\AES_ENC/u0/u2/n1056 ), .A2(\AES_ENC/u0/u2/n1074 ), .ZN(\AES_ENC/u0/u2/n1057 ) );
NOR3_X2 \AES_ENC/u0/u2/U194  ( .A1(\AES_ENC/u0/u2/n607 ), .A2(\AES_ENC/u0/u2/n1120 ), .A3(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n978 ) );
NOR2_X2 \AES_ENC/u0/u2/U187  ( .A1(\AES_ENC/u0/u2/n996 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n998 ) );
NOR2_X2 \AES_ENC/u0/u2/U186  ( .A1(\AES_ENC/u0/u2/n996 ), .A2(\AES_ENC/u0/u2/n911 ), .ZN(\AES_ENC/u0/u2/n1116 ) );
NOR2_X2 \AES_ENC/u0/u2/U185  ( .A1(\AES_ENC/u0/u2/n1074 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n754 ) );
NOR2_X2 \AES_ENC/u0/u2/U184  ( .A1(\AES_ENC/u0/u2/n926 ), .A2(\AES_ENC/u0/u2/n1103 ), .ZN(\AES_ENC/u0/u2/n977 ) );
NOR2_X2 \AES_ENC/u0/u2/U183  ( .A1(\AES_ENC/u0/u2/n839 ), .A2(\AES_ENC/u0/u2/n824 ), .ZN(\AES_ENC/u0/u2/n1092 ) );
NOR2_X2 \AES_ENC/u0/u2/U182  ( .A1(\AES_ENC/u0/u2/n573 ), .A2(\AES_ENC/u0/u2/n1074 ), .ZN(\AES_ENC/u0/u2/n684 ) );
NOR2_X2 \AES_ENC/u0/u2/U181  ( .A1(\AES_ENC/u0/u2/n826 ), .A2(\AES_ENC/u0/u2/n1059 ), .ZN(\AES_ENC/u0/u2/n907 ) );
NOR3_X2 \AES_ENC/u0/u2/U180  ( .A1(\AES_ENC/u0/u2/n625 ), .A2(\AES_ENC/u0/u2/n1115 ), .A3(\AES_ENC/u0/u2/n585 ), .ZN(\AES_ENC/u0/u2/n831 ) );
NOR3_X2 \AES_ENC/u0/u2/U174  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n1056 ), .A3(\AES_ENC/u0/u2/n990 ), .ZN(\AES_ENC/u0/u2/n896 ) );
NOR3_X2 \AES_ENC/u0/u2/U173  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n573 ), .A3(\AES_ENC/u0/u2/n1013 ), .ZN(\AES_ENC/u0/u2/n670 ) );
NOR3_X2 \AES_ENC/u0/u2/U172  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n1091 ), .A3(\AES_ENC/u0/u2/n1022 ), .ZN(\AES_ENC/u0/u2/n843 ) );
NOR2_X2 \AES_ENC/u0/u2/U171  ( .A1(\AES_ENC/u0/u2/n1029 ), .A2(\AES_ENC/u0/u2/n1095 ), .ZN(\AES_ENC/u0/u2/n735 ) );
NOR2_X2 \AES_ENC/u0/u2/U170  ( .A1(\AES_ENC/u0/u2/n1100 ), .A2(\AES_ENC/u0/u2/n854 ), .ZN(\AES_ENC/u0/u2/n860 ) );
NOR4_X2 \AES_ENC/u0/u2/U169  ( .A1(\AES_ENC/u0/u2/n1125 ), .A2(\AES_ENC/u0/u2/n1124 ), .A3(\AES_ENC/u0/u2/n1123 ), .A4(\AES_ENC/u0/u2/n1122 ), .ZN(\AES_ENC/u0/u2/n1126 ) );
NOR4_X2 \AES_ENC/u0/u2/U168  ( .A1(\AES_ENC/u0/u2/n1084 ), .A2(\AES_ENC/u0/u2/n1083 ), .A3(\AES_ENC/u0/u2/n1082 ), .A4(\AES_ENC/u0/u2/n1081 ), .ZN(\AES_ENC/u0/u2/n1085 ) );
NOR2_X2 \AES_ENC/u0/u2/U162  ( .A1(\AES_ENC/u0/u2/n1076 ), .A2(\AES_ENC/u0/u2/n1075 ), .ZN(\AES_ENC/u0/u2/n1086 ) );
NAND3_X2 \AES_ENC/u0/u2/U161  ( .A1(\AES_ENC/u0/u2/n569 ), .A2(\AES_ENC/u0/u2/n582 ), .A3(\AES_ENC/u0/u2/n681 ), .ZN(\AES_ENC/u0/u2/n691 ) );
NOR2_X2 \AES_ENC/u0/u2/U160  ( .A1(\AES_ENC/u0/u2/n683 ), .A2(\AES_ENC/u0/u2/n682 ), .ZN(\AES_ENC/u0/u2/n690 ) );
NOR4_X2 \AES_ENC/u0/u2/U159  ( .A1(\AES_ENC/u0/u2/n983 ), .A2(\AES_ENC/u0/u2/n698 ), .A3(\AES_ENC/u0/u2/n697 ), .A4(\AES_ENC/u0/u2/n696 ), .ZN(\AES_ENC/u0/u2/n699 ) );
NOR3_X2 \AES_ENC/u0/u2/U158  ( .A1(\AES_ENC/u0/u2/n695 ), .A2(\AES_ENC/u0/u2/n694 ), .A3(\AES_ENC/u0/u2/n693 ), .ZN(\AES_ENC/u0/u2/n700 ) );
NOR4_X2 \AES_ENC/u0/u2/U157  ( .A1(\AES_ENC/u0/u2/n896 ), .A2(\AES_ENC/u0/u2/n895 ), .A3(\AES_ENC/u0/u2/n894 ), .A4(\AES_ENC/u0/u2/n893 ), .ZN(\AES_ENC/u0/u2/n897 ) );
NOR2_X2 \AES_ENC/u0/u2/U156  ( .A1(\AES_ENC/u0/u2/n866 ), .A2(\AES_ENC/u0/u2/n865 ), .ZN(\AES_ENC/u0/u2/n872 ) );
NOR4_X2 \AES_ENC/u0/u2/U155  ( .A1(\AES_ENC/u0/u2/n870 ), .A2(\AES_ENC/u0/u2/n869 ), .A3(\AES_ENC/u0/u2/n868 ), .A4(\AES_ENC/u0/u2/n867 ), .ZN(\AES_ENC/u0/u2/n871 ) );
NOR4_X2 \AES_ENC/u0/u2/U154  ( .A1(\AES_ENC/u0/u2/n963 ), .A2(\AES_ENC/u0/u2/n962 ), .A3(\AES_ENC/u0/u2/n961 ), .A4(\AES_ENC/u0/u2/n960 ), .ZN(\AES_ENC/u0/u2/n964 ) );
NOR2_X2 \AES_ENC/u0/u2/U153  ( .A1(\AES_ENC/u0/u2/n958 ), .A2(\AES_ENC/u0/u2/n957 ), .ZN(\AES_ENC/u0/u2/n965 ) );
NOR4_X2 \AES_ENC/u0/u2/U152  ( .A1(\AES_ENC/u0/u2/n950 ), .A2(\AES_ENC/u0/u2/n949 ), .A3(\AES_ENC/u0/u2/n948 ), .A4(\AES_ENC/u0/u2/n947 ), .ZN(\AES_ENC/u0/u2/n951 ) );
NOR2_X2 \AES_ENC/u0/u2/U143  ( .A1(\AES_ENC/u0/u2/n946 ), .A2(\AES_ENC/u0/u2/n945 ), .ZN(\AES_ENC/u0/u2/n952 ) );
NOR4_X2 \AES_ENC/u0/u2/U142  ( .A1(\AES_ENC/u0/u2/n983 ), .A2(\AES_ENC/u0/u2/n982 ), .A3(\AES_ENC/u0/u2/n981 ), .A4(\AES_ENC/u0/u2/n980 ), .ZN(\AES_ENC/u0/u2/n984 ) );
NOR2_X2 \AES_ENC/u0/u2/U141  ( .A1(\AES_ENC/u0/u2/n979 ), .A2(\AES_ENC/u0/u2/n978 ), .ZN(\AES_ENC/u0/u2/n985 ) );
NOR3_X2 \AES_ENC/u0/u2/U140  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n1054 ), .A3(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n961 ) );
NOR3_X2 \AES_ENC/u0/u2/U132  ( .A1(\AES_ENC/u0/u2/n620 ), .A2(\AES_ENC/u0/u2/n1074 ), .A3(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n671 ) );
NOR2_X2 \AES_ENC/u0/u2/U131  ( .A1(\AES_ENC/u0/u2/n1057 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n1062 ) );
NOR2_X2 \AES_ENC/u0/u2/U130  ( .A1(\AES_ENC/u0/u2/n1060 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n1061 ) );
NOR2_X2 \AES_ENC/u0/u2/U129  ( .A1(\AES_ENC/u0/u2/n1055 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n1063 ) );
NOR4_X2 \AES_ENC/u0/u2/U128  ( .A1(\AES_ENC/u0/u2/n1064 ), .A2(\AES_ENC/u0/u2/n1063 ), .A3(\AES_ENC/u0/u2/n1062 ), .A4(\AES_ENC/u0/u2/n1061 ), .ZN(\AES_ENC/u0/u2/n1065 ) );
NOR3_X2 \AES_ENC/u0/u2/U127  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n1120 ), .A3(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n918 ) );
NOR2_X2 \AES_ENC/u0/u2/U126  ( .A1(\AES_ENC/u0/u2/n914 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n915 ) );
NOR3_X2 \AES_ENC/u0/u2/U121  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n573 ), .A3(\AES_ENC/u0/u2/n1013 ), .ZN(\AES_ENC/u0/u2/n917 ) );
NOR4_X2 \AES_ENC/u0/u2/U120  ( .A1(\AES_ENC/u0/u2/n918 ), .A2(\AES_ENC/u0/u2/n917 ), .A3(\AES_ENC/u0/u2/n916 ), .A4(\AES_ENC/u0/u2/n915 ), .ZN(\AES_ENC/u0/u2/n919 ) );
NOR2_X2 \AES_ENC/u0/u2/U119  ( .A1(\AES_ENC/u0/u2/n735 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n687 ) );
NOR2_X2 \AES_ENC/u0/u2/U118  ( .A1(\AES_ENC/u0/u2/n684 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n688 ) );
NOR2_X2 \AES_ENC/u0/u2/U117  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n600 ), .ZN(\AES_ENC/u0/u2/n686 ) );
NOR4_X2 \AES_ENC/u0/u2/U116  ( .A1(\AES_ENC/u0/u2/n688 ), .A2(\AES_ENC/u0/u2/n687 ), .A3(\AES_ENC/u0/u2/n686 ), .A4(\AES_ENC/u0/u2/n685 ), .ZN(\AES_ENC/u0/u2/n689 ) );
NOR2_X2 \AES_ENC/u0/u2/U115  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n582 ), .ZN(\AES_ENC/u0/u2/n770 ) );
NOR2_X2 \AES_ENC/u0/u2/U106  ( .A1(\AES_ENC/u0/u2/n1103 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n772 ) );
NOR2_X2 \AES_ENC/u0/u2/U105  ( .A1(\AES_ENC/u0/u2/n610 ), .A2(\AES_ENC/u0/u2/n599 ), .ZN(\AES_ENC/u0/u2/n773 ) );
NOR4_X2 \AES_ENC/u0/u2/U104  ( .A1(\AES_ENC/u0/u2/n773 ), .A2(\AES_ENC/u0/u2/n772 ), .A3(\AES_ENC/u0/u2/n771 ), .A4(\AES_ENC/u0/u2/n770 ), .ZN(\AES_ENC/u0/u2/n774 ) );
NOR2_X2 \AES_ENC/u0/u2/U103  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n595 ), .ZN(\AES_ENC/u0/u2/n858 ) );
NOR2_X2 \AES_ENC/u0/u2/U102  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n855 ), .ZN(\AES_ENC/u0/u2/n857 ) );
NOR2_X2 \AES_ENC/u0/u2/U101  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n587 ), .ZN(\AES_ENC/u0/u2/n856 ) );
NOR4_X2 \AES_ENC/u0/u2/U100  ( .A1(\AES_ENC/u0/u2/n858 ), .A2(\AES_ENC/u0/u2/n857 ), .A3(\AES_ENC/u0/u2/n856 ), .A4(\AES_ENC/u0/u2/n958 ), .ZN(\AES_ENC/u0/u2/n859 ) );
NOR2_X2 \AES_ENC/u0/u2/U95  ( .A1(\AES_ENC/u0/u2/n583 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n814 ) );
NOR3_X2 \AES_ENC/u0/u2/U94  ( .A1(\AES_ENC/u0/u2/n606 ), .A2(\AES_ENC/u0/u2/n1058 ), .A3(\AES_ENC/u0/u2/n1059 ), .ZN(\AES_ENC/u0/u2/n815 ) );
NOR2_X2 \AES_ENC/u0/u2/U93  ( .A1(\AES_ENC/u0/u2/n907 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n813 ) );
NOR4_X2 \AES_ENC/u0/u2/U92  ( .A1(\AES_ENC/u0/u2/n815 ), .A2(\AES_ENC/u0/u2/n814 ), .A3(\AES_ENC/u0/u2/n813 ), .A4(\AES_ENC/u0/u2/n812 ), .ZN(\AES_ENC/u0/u2/n816 ) );
NOR2_X2 \AES_ENC/u0/u2/U91  ( .A1(\AES_ENC/u0/u2/n617 ), .A2(\AES_ENC/u0/u2/n569 ), .ZN(\AES_ENC/u0/u2/n721 ) );
NOR2_X2 \AES_ENC/u0/u2/U90  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n1096 ), .ZN(\AES_ENC/u0/u2/n722 ) );
NOR2_X2 \AES_ENC/u0/u2/U89  ( .A1(\AES_ENC/u0/u2/n1031 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n723 ) );
NOR4_X2 \AES_ENC/u0/u2/U88  ( .A1(\AES_ENC/u0/u2/n724 ), .A2(\AES_ENC/u0/u2/n723 ), .A3(\AES_ENC/u0/u2/n722 ), .A4(\AES_ENC/u0/u2/n721 ), .ZN(\AES_ENC/u0/u2/n725 ) );
NOR2_X2 \AES_ENC/u0/u2/U87  ( .A1(\AES_ENC/u0/u2/n911 ), .A2(\AES_ENC/u0/u2/n990 ), .ZN(\AES_ENC/u0/u2/n1009 ) );
NOR2_X2 \AES_ENC/u0/u2/U86  ( .A1(\AES_ENC/u0/u2/n1013 ), .A2(\AES_ENC/u0/u2/n573 ), .ZN(\AES_ENC/u0/u2/n1014 ) );
NOR2_X2 \AES_ENC/u0/u2/U81  ( .A1(\AES_ENC/u0/u2/n1014 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n1015 ) );
NOR4_X2 \AES_ENC/u0/u2/U80  ( .A1(\AES_ENC/u0/u2/n1016 ), .A2(\AES_ENC/u0/u2/n1015 ), .A3(\AES_ENC/u0/u2/n1119 ), .A4(\AES_ENC/u0/u2/n1046 ), .ZN(\AES_ENC/u0/u2/n1017 ) );
NOR2_X2 \AES_ENC/u0/u2/U79  ( .A1(\AES_ENC/u0/u2/n606 ), .A2(\AES_ENC/u0/u2/n589 ), .ZN(\AES_ENC/u0/u2/n997 ) );
NOR2_X2 \AES_ENC/u0/u2/U78  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n577 ), .ZN(\AES_ENC/u0/u2/n1000 ) );
NOR2_X2 \AES_ENC/u0/u2/U74  ( .A1(\AES_ENC/u0/u2/n616 ), .A2(\AES_ENC/u0/u2/n1096 ), .ZN(\AES_ENC/u0/u2/n999 ) );
NOR4_X2 \AES_ENC/u0/u2/U73  ( .A1(\AES_ENC/u0/u2/n1000 ), .A2(\AES_ENC/u0/u2/n999 ), .A3(\AES_ENC/u0/u2/n998 ), .A4(\AES_ENC/u0/u2/n997 ), .ZN(\AES_ENC/u0/u2/n1001 ) );
NOR2_X2 \AES_ENC/u0/u2/U72  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n1096 ), .ZN(\AES_ENC/u0/u2/n697 ) );
NOR2_X2 \AES_ENC/u0/u2/U71  ( .A1(\AES_ENC/u0/u2/n620 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n958 ) );
NOR2_X2 \AES_ENC/u0/u2/U65  ( .A1(\AES_ENC/u0/u2/n911 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n983 ) );
NOR2_X2 \AES_ENC/u0/u2/U64  ( .A1(\AES_ENC/u0/u2/n1054 ), .A2(\AES_ENC/u0/u2/n1103 ), .ZN(\AES_ENC/u0/u2/n1031 ) );
INV_X4 \AES_ENC/u0/u2/U63  ( .A(\AES_ENC/u0/u2/n1050 ), .ZN(\AES_ENC/u0/u2/n612 ) );
INV_X4 \AES_ENC/u0/u2/U62  ( .A(\AES_ENC/u0/u2/n1072 ), .ZN(\AES_ENC/u0/u2/n605 ) );
INV_X4 \AES_ENC/u0/u2/U61  ( .A(\AES_ENC/u0/u2/n1073 ), .ZN(\AES_ENC/u0/u2/n604 ) );
NOR2_X2 \AES_ENC/u0/u2/U59  ( .A1(\AES_ENC/u0/u2/n582 ), .A2(\AES_ENC/u0/u2/n613 ), .ZN(\AES_ENC/u0/u2/n880 ) );
NOR3_X2 \AES_ENC/u0/u2/U58  ( .A1(\AES_ENC/u0/u2/n826 ), .A2(\AES_ENC/u0/u2/n1121 ), .A3(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n946 ) );
INV_X4 \AES_ENC/u0/u2/U57  ( .A(\AES_ENC/u0/u2/n1010 ), .ZN(\AES_ENC/u0/u2/n608 ) );
NOR3_X2 \AES_ENC/u0/u2/U50  ( .A1(\AES_ENC/u0/u2/n573 ), .A2(\AES_ENC/u0/u2/n1029 ), .A3(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n1119 ) );
INV_X4 \AES_ENC/u0/u2/U49  ( .A(\AES_ENC/u0/u2/n956 ), .ZN(\AES_ENC/u0/u2/n615 ) );
NOR2_X2 \AES_ENC/u0/u2/U48  ( .A1(\AES_ENC/u0/u2/n623 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n1013 ) );
NOR2_X2 \AES_ENC/u0/u2/U47  ( .A1(\AES_ENC/u0/u2/n620 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n910 ) );
NOR2_X2 \AES_ENC/u0/u2/U46  ( .A1(\AES_ENC/u0/u2/n569 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n1091 ) );
NOR2_X2 \AES_ENC/u0/u2/U45  ( .A1(\AES_ENC/u0/u2/n622 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n990 ) );
NOR2_X2 \AES_ENC/u0/u2/U44  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/u0/u2/n1121 ), .ZN(\AES_ENC/u0/u2/n996 ) );
NOR2_X2 \AES_ENC/u0/u2/U43  ( .A1(\AES_ENC/u0/u2/n610 ), .A2(\AES_ENC/u0/u2/n600 ), .ZN(\AES_ENC/u0/u2/n628 ) );
NOR2_X2 \AES_ENC/u0/u2/U42  ( .A1(\AES_ENC/u0/u2/n576 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n866 ) );
NOR2_X2 \AES_ENC/u0/u2/U41  ( .A1(\AES_ENC/u0/u2/n603 ), .A2(\AES_ENC/u0/u2/n610 ), .ZN(\AES_ENC/u0/u2/n1006 ) );
NOR2_X2 \AES_ENC/u0/u2/U36  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n1117 ), .ZN(\AES_ENC/u0/u2/n1118 ) );
NOR2_X2 \AES_ENC/u0/u2/U35  ( .A1(\AES_ENC/u0/u2/n1119 ), .A2(\AES_ENC/u0/u2/n1118 ), .ZN(\AES_ENC/u0/u2/n1127 ) );
NOR2_X2 \AES_ENC/u0/u2/U34  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n594 ), .ZN(\AES_ENC/u0/u2/n629 ) );
NOR2_X2 \AES_ENC/u0/u2/U33  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n906 ), .ZN(\AES_ENC/u0/u2/n909 ) );
NOR2_X2 \AES_ENC/u0/u2/U32  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n597 ), .ZN(\AES_ENC/u0/u2/n658 ) );
NOR2_X2 \AES_ENC/u0/u2/U31  ( .A1(\AES_ENC/u0/u2/n1116 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n695 ) );
NOR2_X2 \AES_ENC/u0/u2/U30  ( .A1(\AES_ENC/u0/u2/n1078 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n1083 ) );
NOR2_X2 \AES_ENC/u0/u2/U29  ( .A1(\AES_ENC/u0/u2/n941 ), .A2(\AES_ENC/u0/u2/n608 ), .ZN(\AES_ENC/u0/u2/n724 ) );
NOR2_X2 \AES_ENC/u0/u2/U24  ( .A1(\AES_ENC/u0/u2/n576 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n840 ) );
NOR2_X2 \AES_ENC/u0/u2/U23  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n593 ), .ZN(\AES_ENC/u0/u2/n633 ) );
NOR2_X2 \AES_ENC/u0/u2/U21  ( .A1(\AES_ENC/u0/u2/n1009 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n960 ) );
NOR2_X2 \AES_ENC/u0/u2/U20  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n1045 ), .ZN(\AES_ENC/u0/u2/n812 ) );
NOR2_X2 \AES_ENC/u0/u2/U19  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n1080 ), .ZN(\AES_ENC/u0/u2/n1081 ) );
NOR2_X2 \AES_ENC/u0/u2/U18  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n601 ), .ZN(\AES_ENC/u0/u2/n982 ) );
NOR2_X2 \AES_ENC/u0/u2/U17  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n594 ), .ZN(\AES_ENC/u0/u2/n757 ) );
NOR2_X2 \AES_ENC/u0/u2/U16  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n590 ), .ZN(\AES_ENC/u0/u2/n698 ) );
NOR2_X2 \AES_ENC/u0/u2/U15  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n619 ), .ZN(\AES_ENC/u0/u2/n708 ) );
NOR2_X2 \AES_ENC/u0/u2/U10  ( .A1(\AES_ENC/u0/u2/n619 ), .A2(\AES_ENC/u0/u2/n604 ), .ZN(\AES_ENC/u0/u2/n803 ) );
NOR2_X2 \AES_ENC/u0/u2/U9  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n881 ), .ZN(\AES_ENC/u0/u2/n711 ) );
NOR2_X2 \AES_ENC/u0/u2/U8  ( .A1(\AES_ENC/u0/u2/n615 ), .A2(\AES_ENC/u0/u2/n582 ), .ZN(\AES_ENC/u0/u2/n867 ) );
NOR2_X2 \AES_ENC/u0/u2/U7  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n599 ), .ZN(\AES_ENC/u0/u2/n804 ) );
NOR2_X2 \AES_ENC/u0/u2/U6  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n620 ), .ZN(\AES_ENC/u0/u2/n1046 ) );
OR2_X4 \AES_ENC/u0/u2/U5  ( .A1(\AES_ENC/u0/u2/n624 ), .A2(\AES_ENC/w3[1] ),.ZN(\AES_ENC/u0/u2/n570 ) );
OR2_X4 \AES_ENC/u0/u2/U4  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/w3[4] ),.ZN(\AES_ENC/u0/u2/n569 ) );
NAND2_X2 \AES_ENC/u0/u2/U514  ( .A1(\AES_ENC/u0/u2/n1121 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n1030 ) );
AND2_X2 \AES_ENC/u0/u2/U513  ( .A1(\AES_ENC/u0/u2/n597 ), .A2(\AES_ENC/u0/u2/n1030 ), .ZN(\AES_ENC/u0/u2/n1049 ) );
NAND2_X2 \AES_ENC/u0/u2/U511  ( .A1(\AES_ENC/u0/u2/n1049 ), .A2(\AES_ENC/u0/u2/n794 ), .ZN(\AES_ENC/u0/u2/n637 ) );
AND2_X2 \AES_ENC/u0/u2/U493  ( .A1(\AES_ENC/u0/u2/n779 ), .A2(\AES_ENC/u0/u2/n996 ), .ZN(\AES_ENC/u0/u2/n632 ) );
NAND4_X2 \AES_ENC/u0/u2/U485  ( .A1(\AES_ENC/u0/u2/n637 ), .A2(\AES_ENC/u0/u2/n636 ), .A3(\AES_ENC/u0/u2/n635 ), .A4(\AES_ENC/u0/u2/n634 ), .ZN(\AES_ENC/u0/u2/n638 ) );
NAND2_X2 \AES_ENC/u0/u2/U484  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n638 ), .ZN(\AES_ENC/u0/u2/n679 ) );
NAND2_X2 \AES_ENC/u0/u2/U481  ( .A1(\AES_ENC/u0/u2/n1094 ), .A2(\AES_ENC/u0/u2/n591 ), .ZN(\AES_ENC/u0/u2/n648 ) );
NAND2_X2 \AES_ENC/u0/u2/U476  ( .A1(\AES_ENC/u0/u2/n601 ), .A2(\AES_ENC/u0/u2/n590 ), .ZN(\AES_ENC/u0/u2/n762 ) );
NAND2_X2 \AES_ENC/u0/u2/U475  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n762 ), .ZN(\AES_ENC/u0/u2/n647 ) );
NAND4_X2 \AES_ENC/u0/u2/U457  ( .A1(\AES_ENC/u0/u2/n648 ), .A2(\AES_ENC/u0/u2/n647 ), .A3(\AES_ENC/u0/u2/n646 ), .A4(\AES_ENC/u0/u2/n645 ), .ZN(\AES_ENC/u0/u2/n649 ) );
NAND2_X2 \AES_ENC/u0/u2/U456  ( .A1(\AES_ENC/w3[0] ), .A2(\AES_ENC/u0/u2/n649 ), .ZN(\AES_ENC/u0/u2/n665 ) );
NAND2_X2 \AES_ENC/u0/u2/U454  ( .A1(\AES_ENC/u0/u2/n596 ), .A2(\AES_ENC/u0/u2/n623 ), .ZN(\AES_ENC/u0/u2/n855 ) );
NAND2_X2 \AES_ENC/u0/u2/U453  ( .A1(\AES_ENC/u0/u2/n587 ), .A2(\AES_ENC/u0/u2/n855 ), .ZN(\AES_ENC/u0/u2/n821 ) );
NAND2_X2 \AES_ENC/u0/u2/U452  ( .A1(\AES_ENC/u0/u2/n1093 ), .A2(\AES_ENC/u0/u2/n821 ), .ZN(\AES_ENC/u0/u2/n662 ) );
NAND2_X2 \AES_ENC/u0/u2/U451  ( .A1(\AES_ENC/u0/u2/n619 ), .A2(\AES_ENC/u0/u2/n589 ), .ZN(\AES_ENC/u0/u2/n650 ) );
NAND2_X2 \AES_ENC/u0/u2/U450  ( .A1(\AES_ENC/u0/u2/n956 ), .A2(\AES_ENC/u0/u2/n650 ), .ZN(\AES_ENC/u0/u2/n661 ) );
NAND2_X2 \AES_ENC/u0/u2/U449  ( .A1(\AES_ENC/u0/u2/n626 ), .A2(\AES_ENC/u0/u2/n627 ), .ZN(\AES_ENC/u0/u2/n839 ) );
OR2_X2 \AES_ENC/u0/u2/U446  ( .A1(\AES_ENC/u0/u2/n839 ), .A2(\AES_ENC/u0/u2/n932 ), .ZN(\AES_ENC/u0/u2/n656 ) );
NAND2_X2 \AES_ENC/u0/u2/U445  ( .A1(\AES_ENC/u0/u2/n621 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n1096 ) );
NAND2_X2 \AES_ENC/u0/u2/U444  ( .A1(\AES_ENC/u0/u2/n1030 ), .A2(\AES_ENC/u0/u2/n1096 ), .ZN(\AES_ENC/u0/u2/n651 ) );
NAND2_X2 \AES_ENC/u0/u2/U443  ( .A1(\AES_ENC/u0/u2/n1114 ), .A2(\AES_ENC/u0/u2/n651 ), .ZN(\AES_ENC/u0/u2/n655 ) );
OR3_X2 \AES_ENC/u0/u2/U440  ( .A1(\AES_ENC/u0/u2/n1079 ), .A2(\AES_ENC/w3[7] ), .A3(\AES_ENC/u0/u2/n626 ), .ZN(\AES_ENC/u0/u2/n654 ));
NAND2_X2 \AES_ENC/u0/u2/U439  ( .A1(\AES_ENC/u0/u2/n593 ), .A2(\AES_ENC/u0/u2/n601 ), .ZN(\AES_ENC/u0/u2/n652 ) );
NAND4_X2 \AES_ENC/u0/u2/U437  ( .A1(\AES_ENC/u0/u2/n656 ), .A2(\AES_ENC/u0/u2/n655 ), .A3(\AES_ENC/u0/u2/n654 ), .A4(\AES_ENC/u0/u2/n653 ), .ZN(\AES_ENC/u0/u2/n657 ) );
NAND2_X2 \AES_ENC/u0/u2/U436  ( .A1(\AES_ENC/w3[2] ), .A2(\AES_ENC/u0/u2/n657 ), .ZN(\AES_ENC/u0/u2/n660 ) );
NAND4_X2 \AES_ENC/u0/u2/U432  ( .A1(\AES_ENC/u0/u2/n662 ), .A2(\AES_ENC/u0/u2/n661 ), .A3(\AES_ENC/u0/u2/n660 ), .A4(\AES_ENC/u0/u2/n659 ), .ZN(\AES_ENC/u0/u2/n663 ) );
NAND2_X2 \AES_ENC/u0/u2/U431  ( .A1(\AES_ENC/u0/u2/n663 ), .A2(\AES_ENC/u0/u2/n574 ), .ZN(\AES_ENC/u0/u2/n664 ) );
NAND2_X2 \AES_ENC/u0/u2/U430  ( .A1(\AES_ENC/u0/u2/n665 ), .A2(\AES_ENC/u0/u2/n664 ), .ZN(\AES_ENC/u0/u2/n666 ) );
NAND2_X2 \AES_ENC/u0/u2/U429  ( .A1(\AES_ENC/w3[6] ), .A2(\AES_ENC/u0/u2/n666 ), .ZN(\AES_ENC/u0/u2/n678 ) );
NAND2_X2 \AES_ENC/u0/u2/U426  ( .A1(\AES_ENC/u0/u2/n735 ), .A2(\AES_ENC/u0/u2/n1093 ), .ZN(\AES_ENC/u0/u2/n675 ) );
NAND2_X2 \AES_ENC/u0/u2/U425  ( .A1(\AES_ENC/u0/u2/n588 ), .A2(\AES_ENC/u0/u2/n597 ), .ZN(\AES_ENC/u0/u2/n1045 ) );
OR2_X2 \AES_ENC/u0/u2/U424  ( .A1(\AES_ENC/u0/u2/n1045 ), .A2(\AES_ENC/u0/u2/n605 ), .ZN(\AES_ENC/u0/u2/n674 ) );
NAND2_X2 \AES_ENC/u0/u2/U423  ( .A1(\AES_ENC/w3[1] ), .A2(\AES_ENC/u0/u2/n620 ), .ZN(\AES_ENC/u0/u2/n667 ) );
NAND2_X2 \AES_ENC/u0/u2/U422  ( .A1(\AES_ENC/u0/u2/n619 ), .A2(\AES_ENC/u0/u2/n667 ), .ZN(\AES_ENC/u0/u2/n1071 ) );
NAND4_X2 \AES_ENC/u0/u2/U412  ( .A1(\AES_ENC/u0/u2/n675 ), .A2(\AES_ENC/u0/u2/n674 ), .A3(\AES_ENC/u0/u2/n673 ), .A4(\AES_ENC/u0/u2/n672 ), .ZN(\AES_ENC/u0/u2/n676 ) );
NAND2_X2 \AES_ENC/u0/u2/U411  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n676 ), .ZN(\AES_ENC/u0/u2/n677 ) );
NAND2_X2 \AES_ENC/u0/u2/U408  ( .A1(\AES_ENC/u0/u2/n800 ), .A2(\AES_ENC/u0/u2/n1022 ), .ZN(\AES_ENC/u0/u2/n680 ) );
NAND2_X2 \AES_ENC/u0/u2/U407  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n680 ), .ZN(\AES_ENC/u0/u2/n681 ) );
AND2_X2 \AES_ENC/u0/u2/U402  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n684 ), .ZN(\AES_ENC/u0/u2/n682 ) );
NAND4_X2 \AES_ENC/u0/u2/U395  ( .A1(\AES_ENC/u0/u2/n691 ), .A2(\AES_ENC/u0/u2/n581 ), .A3(\AES_ENC/u0/u2/n690 ), .A4(\AES_ENC/u0/u2/n689 ), .ZN(\AES_ENC/u0/u2/n692 ) );
NAND2_X2 \AES_ENC/u0/u2/U394  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n692 ), .ZN(\AES_ENC/u0/u2/n733 ) );
NAND2_X2 \AES_ENC/u0/u2/U392  ( .A1(\AES_ENC/u0/u2/n977 ), .A2(\AES_ENC/u0/u2/n1050 ), .ZN(\AES_ENC/u0/u2/n702 ) );
NAND2_X2 \AES_ENC/u0/u2/U391  ( .A1(\AES_ENC/u0/u2/n1093 ), .A2(\AES_ENC/u0/u2/n1045 ), .ZN(\AES_ENC/u0/u2/n701 ) );
NAND4_X2 \AES_ENC/u0/u2/U381  ( .A1(\AES_ENC/u0/u2/n702 ), .A2(\AES_ENC/u0/u2/n701 ), .A3(\AES_ENC/u0/u2/n700 ), .A4(\AES_ENC/u0/u2/n699 ), .ZN(\AES_ENC/u0/u2/n703 ) );
NAND2_X2 \AES_ENC/u0/u2/U380  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n703 ), .ZN(\AES_ENC/u0/u2/n732 ) );
AND2_X2 \AES_ENC/u0/u2/U379  ( .A1(\AES_ENC/w3[0] ), .A2(\AES_ENC/w3[6] ),.ZN(\AES_ENC/u0/u2/n1113 ) );
NAND2_X2 \AES_ENC/u0/u2/U378  ( .A1(\AES_ENC/u0/u2/n601 ), .A2(\AES_ENC/u0/u2/n1030 ), .ZN(\AES_ENC/u0/u2/n881 ) );
NAND2_X2 \AES_ENC/u0/u2/U377  ( .A1(\AES_ENC/u0/u2/n1093 ), .A2(\AES_ENC/u0/u2/n881 ), .ZN(\AES_ENC/u0/u2/n715 ) );
NAND2_X2 \AES_ENC/u0/u2/U376  ( .A1(\AES_ENC/u0/u2/n1010 ), .A2(\AES_ENC/u0/u2/n600 ), .ZN(\AES_ENC/u0/u2/n714 ) );
NAND2_X2 \AES_ENC/u0/u2/U375  ( .A1(\AES_ENC/u0/u2/n855 ), .A2(\AES_ENC/u0/u2/n588 ), .ZN(\AES_ENC/u0/u2/n1117 ) );
XNOR2_X2 \AES_ENC/u0/u2/U371  ( .A(\AES_ENC/u0/u2/n611 ), .B(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n824 ) );
NAND4_X2 \AES_ENC/u0/u2/U362  ( .A1(\AES_ENC/u0/u2/n715 ), .A2(\AES_ENC/u0/u2/n714 ), .A3(\AES_ENC/u0/u2/n713 ), .A4(\AES_ENC/u0/u2/n712 ), .ZN(\AES_ENC/u0/u2/n716 ) );
NAND2_X2 \AES_ENC/u0/u2/U361  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n716 ), .ZN(\AES_ENC/u0/u2/n731 ) );
AND2_X2 \AES_ENC/u0/u2/U360  ( .A1(\AES_ENC/w3[6] ), .A2(\AES_ENC/u0/u2/n574 ), .ZN(\AES_ENC/u0/u2/n1131 ) );
NAND2_X2 \AES_ENC/u0/u2/U359  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n717 ) );
NAND2_X2 \AES_ENC/u0/u2/U358  ( .A1(\AES_ENC/u0/u2/n1029 ), .A2(\AES_ENC/u0/u2/n717 ), .ZN(\AES_ENC/u0/u2/n728 ) );
NAND2_X2 \AES_ENC/u0/u2/U357  ( .A1(\AES_ENC/w3[1] ), .A2(\AES_ENC/u0/u2/n624 ), .ZN(\AES_ENC/u0/u2/n1097 ) );
NAND2_X2 \AES_ENC/u0/u2/U356  ( .A1(\AES_ENC/u0/u2/n603 ), .A2(\AES_ENC/u0/u2/n1097 ), .ZN(\AES_ENC/u0/u2/n718 ) );
NAND2_X2 \AES_ENC/u0/u2/U355  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n718 ), .ZN(\AES_ENC/u0/u2/n727 ) );
NAND4_X2 \AES_ENC/u0/u2/U344  ( .A1(\AES_ENC/u0/u2/n728 ), .A2(\AES_ENC/u0/u2/n727 ), .A3(\AES_ENC/u0/u2/n726 ), .A4(\AES_ENC/u0/u2/n725 ), .ZN(\AES_ENC/u0/u2/n729 ) );
NAND2_X2 \AES_ENC/u0/u2/U343  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n729 ), .ZN(\AES_ENC/u0/u2/n730 ) );
NAND4_X2 \AES_ENC/u0/u2/U342  ( .A1(\AES_ENC/u0/u2/n733 ), .A2(\AES_ENC/u0/u2/n732 ), .A3(\AES_ENC/u0/u2/n731 ), .A4(\AES_ENC/u0/u2/n730 ), .ZN(\AES_ENC/u0/subword[9] ) );
NAND2_X2 \AES_ENC/u0/u2/U341  ( .A1(\AES_ENC/w3[7] ), .A2(\AES_ENC/u0/u2/n611 ), .ZN(\AES_ENC/u0/u2/n734 ) );
NAND2_X2 \AES_ENC/u0/u2/U340  ( .A1(\AES_ENC/u0/u2/n734 ), .A2(\AES_ENC/u0/u2/n607 ), .ZN(\AES_ENC/u0/u2/n738 ) );
OR4_X2 \AES_ENC/u0/u2/U339  ( .A1(\AES_ENC/u0/u2/n738 ), .A2(\AES_ENC/u0/u2/n626 ), .A3(\AES_ENC/u0/u2/n826 ), .A4(\AES_ENC/u0/u2/n1121 ), .ZN(\AES_ENC/u0/u2/n746 ) );
NAND2_X2 \AES_ENC/u0/u2/U337  ( .A1(\AES_ENC/u0/u2/n1100 ), .A2(\AES_ENC/u0/u2/n587 ), .ZN(\AES_ENC/u0/u2/n992 ) );
OR2_X2 \AES_ENC/u0/u2/U336  ( .A1(\AES_ENC/u0/u2/n610 ), .A2(\AES_ENC/u0/u2/n735 ), .ZN(\AES_ENC/u0/u2/n737 ) );
NAND2_X2 \AES_ENC/u0/u2/U334  ( .A1(\AES_ENC/u0/u2/n619 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n753 ) );
NAND2_X2 \AES_ENC/u0/u2/U333  ( .A1(\AES_ENC/u0/u2/n582 ), .A2(\AES_ENC/u0/u2/n753 ), .ZN(\AES_ENC/u0/u2/n1080 ) );
NAND2_X2 \AES_ENC/u0/u2/U332  ( .A1(\AES_ENC/u0/u2/n1048 ), .A2(\AES_ENC/u0/u2/n576 ), .ZN(\AES_ENC/u0/u2/n736 ) );
NAND2_X2 \AES_ENC/u0/u2/U331  ( .A1(\AES_ENC/u0/u2/n737 ), .A2(\AES_ENC/u0/u2/n736 ), .ZN(\AES_ENC/u0/u2/n739 ) );
NAND2_X2 \AES_ENC/u0/u2/U330  ( .A1(\AES_ENC/u0/u2/n739 ), .A2(\AES_ENC/u0/u2/n738 ), .ZN(\AES_ENC/u0/u2/n745 ) );
NAND2_X2 \AES_ENC/u0/u2/U326  ( .A1(\AES_ENC/u0/u2/n1096 ), .A2(\AES_ENC/u0/u2/n590 ), .ZN(\AES_ENC/u0/u2/n906 ) );
NAND4_X2 \AES_ENC/u0/u2/U323  ( .A1(\AES_ENC/u0/u2/n746 ), .A2(\AES_ENC/u0/u2/n992 ), .A3(\AES_ENC/u0/u2/n745 ), .A4(\AES_ENC/u0/u2/n744 ), .ZN(\AES_ENC/u0/u2/n747 ) );
NAND2_X2 \AES_ENC/u0/u2/U322  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n747 ), .ZN(\AES_ENC/u0/u2/n793 ) );
NAND2_X2 \AES_ENC/u0/u2/U321  ( .A1(\AES_ENC/u0/u2/n584 ), .A2(\AES_ENC/u0/u2/n855 ), .ZN(\AES_ENC/u0/u2/n748 ) );
NAND2_X2 \AES_ENC/u0/u2/U320  ( .A1(\AES_ENC/u0/u2/n956 ), .A2(\AES_ENC/u0/u2/n748 ), .ZN(\AES_ENC/u0/u2/n760 ) );
NAND2_X2 \AES_ENC/u0/u2/U313  ( .A1(\AES_ENC/u0/u2/n590 ), .A2(\AES_ENC/u0/u2/n753 ), .ZN(\AES_ENC/u0/u2/n1023 ) );
NAND4_X2 \AES_ENC/u0/u2/U308  ( .A1(\AES_ENC/u0/u2/n760 ), .A2(\AES_ENC/u0/u2/n992 ), .A3(\AES_ENC/u0/u2/n759 ), .A4(\AES_ENC/u0/u2/n758 ), .ZN(\AES_ENC/u0/u2/n761 ) );
NAND2_X2 \AES_ENC/u0/u2/U307  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n761 ), .ZN(\AES_ENC/u0/u2/n792 ) );
NAND2_X2 \AES_ENC/u0/u2/U306  ( .A1(\AES_ENC/u0/u2/n584 ), .A2(\AES_ENC/u0/u2/n603 ), .ZN(\AES_ENC/u0/u2/n989 ) );
NAND2_X2 \AES_ENC/u0/u2/U305  ( .A1(\AES_ENC/u0/u2/n1050 ), .A2(\AES_ENC/u0/u2/n989 ), .ZN(\AES_ENC/u0/u2/n777 ) );
NAND2_X2 \AES_ENC/u0/u2/U304  ( .A1(\AES_ENC/u0/u2/n1093 ), .A2(\AES_ENC/u0/u2/n762 ), .ZN(\AES_ENC/u0/u2/n776 ) );
XNOR2_X2 \AES_ENC/u0/u2/U301  ( .A(\AES_ENC/w3[7] ), .B(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n959 ) );
NAND4_X2 \AES_ENC/u0/u2/U289  ( .A1(\AES_ENC/u0/u2/n777 ), .A2(\AES_ENC/u0/u2/n776 ), .A3(\AES_ENC/u0/u2/n775 ), .A4(\AES_ENC/u0/u2/n774 ), .ZN(\AES_ENC/u0/u2/n778 ) );
NAND2_X2 \AES_ENC/u0/u2/U288  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n778 ), .ZN(\AES_ENC/u0/u2/n791 ) );
NAND2_X2 \AES_ENC/u0/u2/U287  ( .A1(\AES_ENC/u0/u2/n1056 ), .A2(\AES_ENC/u0/u2/n1050 ), .ZN(\AES_ENC/u0/u2/n788 ) );
NAND2_X2 \AES_ENC/u0/u2/U286  ( .A1(\AES_ENC/u0/u2/n1091 ), .A2(\AES_ENC/u0/u2/n779 ), .ZN(\AES_ENC/u0/u2/n787 ) );
NAND2_X2 \AES_ENC/u0/u2/U285  ( .A1(\AES_ENC/u0/u2/n956 ), .A2(\AES_ENC/w3[1] ), .ZN(\AES_ENC/u0/u2/n786 ) );
NAND4_X2 \AES_ENC/u0/u2/U278  ( .A1(\AES_ENC/u0/u2/n788 ), .A2(\AES_ENC/u0/u2/n787 ), .A3(\AES_ENC/u0/u2/n786 ), .A4(\AES_ENC/u0/u2/n785 ), .ZN(\AES_ENC/u0/u2/n789 ) );
NAND2_X2 \AES_ENC/u0/u2/U277  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n789 ), .ZN(\AES_ENC/u0/u2/n790 ) );
NAND4_X2 \AES_ENC/u0/u2/U276  ( .A1(\AES_ENC/u0/u2/n793 ), .A2(\AES_ENC/u0/u2/n792 ), .A3(\AES_ENC/u0/u2/n791 ), .A4(\AES_ENC/u0/u2/n790 ), .ZN(\AES_ENC/u0/subword[10] ) );
NAND2_X2 \AES_ENC/u0/u2/U275  ( .A1(\AES_ENC/u0/u2/n1059 ), .A2(\AES_ENC/u0/u2/n794 ), .ZN(\AES_ENC/u0/u2/n810 ) );
NAND2_X2 \AES_ENC/u0/u2/U274  ( .A1(\AES_ENC/u0/u2/n1049 ), .A2(\AES_ENC/u0/u2/n956 ), .ZN(\AES_ENC/u0/u2/n809 ) );
OR2_X2 \AES_ENC/u0/u2/U266  ( .A1(\AES_ENC/u0/u2/n1096 ), .A2(\AES_ENC/u0/u2/n606 ), .ZN(\AES_ENC/u0/u2/n802 ) );
NAND2_X2 \AES_ENC/u0/u2/U265  ( .A1(\AES_ENC/u0/u2/n1053 ), .A2(\AES_ENC/u0/u2/n800 ), .ZN(\AES_ENC/u0/u2/n801 ) );
NAND2_X2 \AES_ENC/u0/u2/U264  ( .A1(\AES_ENC/u0/u2/n802 ), .A2(\AES_ENC/u0/u2/n801 ), .ZN(\AES_ENC/u0/u2/n805 ) );
NAND4_X2 \AES_ENC/u0/u2/U261  ( .A1(\AES_ENC/u0/u2/n810 ), .A2(\AES_ENC/u0/u2/n809 ), .A3(\AES_ENC/u0/u2/n808 ), .A4(\AES_ENC/u0/u2/n807 ), .ZN(\AES_ENC/u0/u2/n811 ) );
NAND2_X2 \AES_ENC/u0/u2/U260  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n811 ), .ZN(\AES_ENC/u0/u2/n852 ) );
OR2_X2 \AES_ENC/u0/u2/U259  ( .A1(\AES_ENC/u0/u2/n1023 ), .A2(\AES_ENC/u0/u2/n617 ), .ZN(\AES_ENC/u0/u2/n819 ) );
OR2_X2 \AES_ENC/u0/u2/U257  ( .A1(\AES_ENC/u0/u2/n570 ), .A2(\AES_ENC/u0/u2/n930 ), .ZN(\AES_ENC/u0/u2/n818 ) );
NAND2_X2 \AES_ENC/u0/u2/U256  ( .A1(\AES_ENC/u0/u2/n1013 ), .A2(\AES_ENC/u0/u2/n1094 ), .ZN(\AES_ENC/u0/u2/n817 ) );
NAND4_X2 \AES_ENC/u0/u2/U249  ( .A1(\AES_ENC/u0/u2/n819 ), .A2(\AES_ENC/u0/u2/n818 ), .A3(\AES_ENC/u0/u2/n817 ), .A4(\AES_ENC/u0/u2/n816 ), .ZN(\AES_ENC/u0/u2/n820 ) );
NAND2_X2 \AES_ENC/u0/u2/U248  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n820 ), .ZN(\AES_ENC/u0/u2/n851 ) );
NAND2_X2 \AES_ENC/u0/u2/U247  ( .A1(\AES_ENC/u0/u2/n956 ), .A2(\AES_ENC/u0/u2/n1080 ), .ZN(\AES_ENC/u0/u2/n835 ) );
NAND2_X2 \AES_ENC/u0/u2/U246  ( .A1(\AES_ENC/u0/u2/n570 ), .A2(\AES_ENC/u0/u2/n1030 ), .ZN(\AES_ENC/u0/u2/n1047 ) );
OR2_X2 \AES_ENC/u0/u2/U245  ( .A1(\AES_ENC/u0/u2/n1047 ), .A2(\AES_ENC/u0/u2/n612 ), .ZN(\AES_ENC/u0/u2/n834 ) );
NAND2_X2 \AES_ENC/u0/u2/U244  ( .A1(\AES_ENC/u0/u2/n1072 ), .A2(\AES_ENC/u0/u2/n589 ), .ZN(\AES_ENC/u0/u2/n833 ) );
NAND4_X2 \AES_ENC/u0/u2/U233  ( .A1(\AES_ENC/u0/u2/n835 ), .A2(\AES_ENC/u0/u2/n834 ), .A3(\AES_ENC/u0/u2/n833 ), .A4(\AES_ENC/u0/u2/n832 ), .ZN(\AES_ENC/u0/u2/n836 ) );
NAND2_X2 \AES_ENC/u0/u2/U232  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n836 ), .ZN(\AES_ENC/u0/u2/n850 ) );
NAND2_X2 \AES_ENC/u0/u2/U231  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n623 ), .ZN(\AES_ENC/u0/u2/n847 ) );
NAND2_X2 \AES_ENC/u0/u2/U230  ( .A1(\AES_ENC/u0/u2/n1050 ), .A2(\AES_ENC/u0/u2/n1071 ), .ZN(\AES_ENC/u0/u2/n846 ) );
OR2_X2 \AES_ENC/u0/u2/U224  ( .A1(\AES_ENC/u0/u2/n1053 ), .A2(\AES_ENC/u0/u2/n911 ), .ZN(\AES_ENC/u0/u2/n1077 ) );
NAND4_X2 \AES_ENC/u0/u2/U220  ( .A1(\AES_ENC/u0/u2/n847 ), .A2(\AES_ENC/u0/u2/n846 ), .A3(\AES_ENC/u0/u2/n845 ), .A4(\AES_ENC/u0/u2/n844 ), .ZN(\AES_ENC/u0/u2/n848 ) );
NAND2_X2 \AES_ENC/u0/u2/U219  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n848 ), .ZN(\AES_ENC/u0/u2/n849 ) );
NAND4_X2 \AES_ENC/u0/u2/U218  ( .A1(\AES_ENC/u0/u2/n852 ), .A2(\AES_ENC/u0/u2/n851 ), .A3(\AES_ENC/u0/u2/n850 ), .A4(\AES_ENC/u0/u2/n849 ), .ZN(\AES_ENC/u0/subword[11] ) );
NAND2_X2 \AES_ENC/u0/u2/U216  ( .A1(\AES_ENC/u0/u2/n1009 ), .A2(\AES_ENC/u0/u2/n1072 ), .ZN(\AES_ENC/u0/u2/n862 ) );
NAND2_X2 \AES_ENC/u0/u2/U215  ( .A1(\AES_ENC/u0/u2/n603 ), .A2(\AES_ENC/u0/u2/n577 ), .ZN(\AES_ENC/u0/u2/n853 ) );
NAND2_X2 \AES_ENC/u0/u2/U214  ( .A1(\AES_ENC/u0/u2/n1050 ), .A2(\AES_ENC/u0/u2/n853 ), .ZN(\AES_ENC/u0/u2/n861 ) );
NAND4_X2 \AES_ENC/u0/u2/U206  ( .A1(\AES_ENC/u0/u2/n862 ), .A2(\AES_ENC/u0/u2/n861 ), .A3(\AES_ENC/u0/u2/n860 ), .A4(\AES_ENC/u0/u2/n859 ), .ZN(\AES_ENC/u0/u2/n863 ) );
NAND2_X2 \AES_ENC/u0/u2/U205  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n863 ), .ZN(\AES_ENC/u0/u2/n905 ) );
NAND2_X2 \AES_ENC/u0/u2/U204  ( .A1(\AES_ENC/u0/u2/n1010 ), .A2(\AES_ENC/u0/u2/n989 ), .ZN(\AES_ENC/u0/u2/n874 ) );
NAND2_X2 \AES_ENC/u0/u2/U203  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n610 ), .ZN(\AES_ENC/u0/u2/n864 ) );
NAND2_X2 \AES_ENC/u0/u2/U202  ( .A1(\AES_ENC/u0/u2/n929 ), .A2(\AES_ENC/u0/u2/n864 ), .ZN(\AES_ENC/u0/u2/n873 ) );
NAND4_X2 \AES_ENC/u0/u2/U193  ( .A1(\AES_ENC/u0/u2/n874 ), .A2(\AES_ENC/u0/u2/n873 ), .A3(\AES_ENC/u0/u2/n872 ), .A4(\AES_ENC/u0/u2/n871 ), .ZN(\AES_ENC/u0/u2/n875 ) );
NAND2_X2 \AES_ENC/u0/u2/U192  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n875 ), .ZN(\AES_ENC/u0/u2/n904 ) );
NAND2_X2 \AES_ENC/u0/u2/U191  ( .A1(\AES_ENC/u0/u2/n583 ), .A2(\AES_ENC/u0/u2/n1050 ), .ZN(\AES_ENC/u0/u2/n889 ) );
NAND2_X2 \AES_ENC/u0/u2/U190  ( .A1(\AES_ENC/u0/u2/n1093 ), .A2(\AES_ENC/u0/u2/n587 ), .ZN(\AES_ENC/u0/u2/n876 ) );
NAND2_X2 \AES_ENC/u0/u2/U189  ( .A1(\AES_ENC/u0/u2/n604 ), .A2(\AES_ENC/u0/u2/n876 ), .ZN(\AES_ENC/u0/u2/n877 ) );
NAND2_X2 \AES_ENC/u0/u2/U188  ( .A1(\AES_ENC/u0/u2/n877 ), .A2(\AES_ENC/u0/u2/n623 ), .ZN(\AES_ENC/u0/u2/n888 ) );
NAND4_X2 \AES_ENC/u0/u2/U179  ( .A1(\AES_ENC/u0/u2/n889 ), .A2(\AES_ENC/u0/u2/n888 ), .A3(\AES_ENC/u0/u2/n887 ), .A4(\AES_ENC/u0/u2/n886 ), .ZN(\AES_ENC/u0/u2/n890 ) );
NAND2_X2 \AES_ENC/u0/u2/U178  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n890 ), .ZN(\AES_ENC/u0/u2/n903 ) );
OR2_X2 \AES_ENC/u0/u2/U177  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n1059 ), .ZN(\AES_ENC/u0/u2/n900 ) );
NAND2_X2 \AES_ENC/u0/u2/U176  ( .A1(\AES_ENC/u0/u2/n1073 ), .A2(\AES_ENC/u0/u2/n1047 ), .ZN(\AES_ENC/u0/u2/n899 ) );
NAND2_X2 \AES_ENC/u0/u2/U175  ( .A1(\AES_ENC/u0/u2/n1094 ), .A2(\AES_ENC/u0/u2/n595 ), .ZN(\AES_ENC/u0/u2/n898 ) );
NAND4_X2 \AES_ENC/u0/u2/U167  ( .A1(\AES_ENC/u0/u2/n900 ), .A2(\AES_ENC/u0/u2/n899 ), .A3(\AES_ENC/u0/u2/n898 ), .A4(\AES_ENC/u0/u2/n897 ), .ZN(\AES_ENC/u0/u2/n901 ) );
NAND2_X2 \AES_ENC/u0/u2/U166  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n901 ), .ZN(\AES_ENC/u0/u2/n902 ) );
NAND4_X2 \AES_ENC/u0/u2/U165  ( .A1(\AES_ENC/u0/u2/n905 ), .A2(\AES_ENC/u0/u2/n904 ), .A3(\AES_ENC/u0/u2/n903 ), .A4(\AES_ENC/u0/u2/n902 ), .ZN(\AES_ENC/u0/subword[12] ) );
NAND2_X2 \AES_ENC/u0/u2/U164  ( .A1(\AES_ENC/u0/u2/n1094 ), .A2(\AES_ENC/u0/u2/n599 ), .ZN(\AES_ENC/u0/u2/n922 ) );
NAND2_X2 \AES_ENC/u0/u2/U163  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n989 ), .ZN(\AES_ENC/u0/u2/n921 ) );
NAND4_X2 \AES_ENC/u0/u2/U151  ( .A1(\AES_ENC/u0/u2/n922 ), .A2(\AES_ENC/u0/u2/n921 ), .A3(\AES_ENC/u0/u2/n920 ), .A4(\AES_ENC/u0/u2/n919 ), .ZN(\AES_ENC/u0/u2/n923 ) );
NAND2_X2 \AES_ENC/u0/u2/U150  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n923 ), .ZN(\AES_ENC/u0/u2/n972 ) );
NAND2_X2 \AES_ENC/u0/u2/U149  ( .A1(\AES_ENC/u0/u2/n582 ), .A2(\AES_ENC/u0/u2/n619 ), .ZN(\AES_ENC/u0/u2/n924 ) );
NAND2_X2 \AES_ENC/u0/u2/U148  ( .A1(\AES_ENC/u0/u2/n1073 ), .A2(\AES_ENC/u0/u2/n924 ), .ZN(\AES_ENC/u0/u2/n939 ) );
NAND2_X2 \AES_ENC/u0/u2/U147  ( .A1(\AES_ENC/u0/u2/n926 ), .A2(\AES_ENC/u0/u2/n925 ), .ZN(\AES_ENC/u0/u2/n927 ) );
NAND2_X2 \AES_ENC/u0/u2/U146  ( .A1(\AES_ENC/u0/u2/n606 ), .A2(\AES_ENC/u0/u2/n927 ), .ZN(\AES_ENC/u0/u2/n928 ) );
NAND2_X2 \AES_ENC/u0/u2/U145  ( .A1(\AES_ENC/u0/u2/n928 ), .A2(\AES_ENC/u0/u2/n1080 ), .ZN(\AES_ENC/u0/u2/n938 ) );
OR2_X2 \AES_ENC/u0/u2/U144  ( .A1(\AES_ENC/u0/u2/n1117 ), .A2(\AES_ENC/u0/u2/n615 ), .ZN(\AES_ENC/u0/u2/n937 ) );
NAND4_X2 \AES_ENC/u0/u2/U139  ( .A1(\AES_ENC/u0/u2/n939 ), .A2(\AES_ENC/u0/u2/n938 ), .A3(\AES_ENC/u0/u2/n937 ), .A4(\AES_ENC/u0/u2/n936 ), .ZN(\AES_ENC/u0/u2/n940 ) );
NAND2_X2 \AES_ENC/u0/u2/U138  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n940 ), .ZN(\AES_ENC/u0/u2/n971 ) );
OR2_X2 \AES_ENC/u0/u2/U137  ( .A1(\AES_ENC/u0/u2/n605 ), .A2(\AES_ENC/u0/u2/n941 ), .ZN(\AES_ENC/u0/u2/n954 ) );
NAND2_X2 \AES_ENC/u0/u2/U136  ( .A1(\AES_ENC/u0/u2/n1096 ), .A2(\AES_ENC/u0/u2/n577 ), .ZN(\AES_ENC/u0/u2/n942 ) );
NAND2_X2 \AES_ENC/u0/u2/U135  ( .A1(\AES_ENC/u0/u2/n1048 ), .A2(\AES_ENC/u0/u2/n942 ), .ZN(\AES_ENC/u0/u2/n943 ) );
NAND2_X2 \AES_ENC/u0/u2/U134  ( .A1(\AES_ENC/u0/u2/n612 ), .A2(\AES_ENC/u0/u2/n943 ), .ZN(\AES_ENC/u0/u2/n944 ) );
NAND2_X2 \AES_ENC/u0/u2/U133  ( .A1(\AES_ENC/u0/u2/n944 ), .A2(\AES_ENC/u0/u2/n580 ), .ZN(\AES_ENC/u0/u2/n953 ) );
NAND4_X2 \AES_ENC/u0/u2/U125  ( .A1(\AES_ENC/u0/u2/n954 ), .A2(\AES_ENC/u0/u2/n953 ), .A3(\AES_ENC/u0/u2/n952 ), .A4(\AES_ENC/u0/u2/n951 ), .ZN(\AES_ENC/u0/u2/n955 ) );
NAND2_X2 \AES_ENC/u0/u2/U124  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n955 ), .ZN(\AES_ENC/u0/u2/n970 ) );
NAND2_X2 \AES_ENC/u0/u2/U123  ( .A1(\AES_ENC/u0/u2/n1094 ), .A2(\AES_ENC/u0/u2/n1071 ), .ZN(\AES_ENC/u0/u2/n967 ) );
NAND2_X2 \AES_ENC/u0/u2/U122  ( .A1(\AES_ENC/u0/u2/n956 ), .A2(\AES_ENC/u0/u2/n1030 ), .ZN(\AES_ENC/u0/u2/n966 ) );
NAND4_X2 \AES_ENC/u0/u2/U114  ( .A1(\AES_ENC/u0/u2/n967 ), .A2(\AES_ENC/u0/u2/n966 ), .A3(\AES_ENC/u0/u2/n965 ), .A4(\AES_ENC/u0/u2/n964 ), .ZN(\AES_ENC/u0/u2/n968 ) );
NAND2_X2 \AES_ENC/u0/u2/U113  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n968 ), .ZN(\AES_ENC/u0/u2/n969 ) );
NAND4_X2 \AES_ENC/u0/u2/U112  ( .A1(\AES_ENC/u0/u2/n972 ), .A2(\AES_ENC/u0/u2/n971 ), .A3(\AES_ENC/u0/u2/n970 ), .A4(\AES_ENC/u0/u2/n969 ), .ZN(\AES_ENC/u0/subword[13] ) );
NAND2_X2 \AES_ENC/u0/u2/U111  ( .A1(\AES_ENC/u0/u2/n570 ), .A2(\AES_ENC/u0/u2/n1097 ), .ZN(\AES_ENC/u0/u2/n973 ) );
NAND2_X2 \AES_ENC/u0/u2/U110  ( .A1(\AES_ENC/u0/u2/n1073 ), .A2(\AES_ENC/u0/u2/n973 ), .ZN(\AES_ENC/u0/u2/n987 ) );
NAND2_X2 \AES_ENC/u0/u2/U109  ( .A1(\AES_ENC/u0/u2/n974 ), .A2(\AES_ENC/u0/u2/n1077 ), .ZN(\AES_ENC/u0/u2/n975 ) );
NAND2_X2 \AES_ENC/u0/u2/U108  ( .A1(\AES_ENC/u0/u2/n613 ), .A2(\AES_ENC/u0/u2/n975 ), .ZN(\AES_ENC/u0/u2/n976 ) );
NAND2_X2 \AES_ENC/u0/u2/U107  ( .A1(\AES_ENC/u0/u2/n977 ), .A2(\AES_ENC/u0/u2/n976 ), .ZN(\AES_ENC/u0/u2/n986 ) );
NAND4_X2 \AES_ENC/u0/u2/U99  ( .A1(\AES_ENC/u0/u2/n987 ), .A2(\AES_ENC/u0/u2/n986 ), .A3(\AES_ENC/u0/u2/n985 ), .A4(\AES_ENC/u0/u2/n984 ), .ZN(\AES_ENC/u0/u2/n988 ) );
NAND2_X2 \AES_ENC/u0/u2/U98  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n988 ), .ZN(\AES_ENC/u0/u2/n1044 ) );
NAND2_X2 \AES_ENC/u0/u2/U97  ( .A1(\AES_ENC/u0/u2/n1073 ), .A2(\AES_ENC/u0/u2/n989 ), .ZN(\AES_ENC/u0/u2/n1004 ) );
NAND2_X2 \AES_ENC/u0/u2/U96  ( .A1(\AES_ENC/u0/u2/n1092 ), .A2(\AES_ENC/u0/u2/n619 ), .ZN(\AES_ENC/u0/u2/n1003 ) );
NAND4_X2 \AES_ENC/u0/u2/U85  ( .A1(\AES_ENC/u0/u2/n1004 ), .A2(\AES_ENC/u0/u2/n1003 ), .A3(\AES_ENC/u0/u2/n1002 ), .A4(\AES_ENC/u0/u2/n1001 ), .ZN(\AES_ENC/u0/u2/n1005 ) );
NAND2_X2 \AES_ENC/u0/u2/U84  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n1005 ), .ZN(\AES_ENC/u0/u2/n1043 ) );
NAND2_X2 \AES_ENC/u0/u2/U83  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n596 ), .ZN(\AES_ENC/u0/u2/n1020 ) );
NAND2_X2 \AES_ENC/u0/u2/U82  ( .A1(\AES_ENC/u0/u2/n1050 ), .A2(\AES_ENC/u0/u2/n624 ), .ZN(\AES_ENC/u0/u2/n1019 ) );
NAND2_X2 \AES_ENC/u0/u2/U77  ( .A1(\AES_ENC/u0/u2/n1059 ), .A2(\AES_ENC/u0/u2/n1114 ), .ZN(\AES_ENC/u0/u2/n1012 ) );
NAND2_X2 \AES_ENC/u0/u2/U76  ( .A1(\AES_ENC/u0/u2/n1010 ), .A2(\AES_ENC/u0/u2/n592 ), .ZN(\AES_ENC/u0/u2/n1011 ) );
NAND2_X2 \AES_ENC/u0/u2/U75  ( .A1(\AES_ENC/u0/u2/n1012 ), .A2(\AES_ENC/u0/u2/n1011 ), .ZN(\AES_ENC/u0/u2/n1016 ) );
NAND4_X2 \AES_ENC/u0/u2/U70  ( .A1(\AES_ENC/u0/u2/n1020 ), .A2(\AES_ENC/u0/u2/n1019 ), .A3(\AES_ENC/u0/u2/n1018 ), .A4(\AES_ENC/u0/u2/n1017 ), .ZN(\AES_ENC/u0/u2/n1021 ) );
NAND2_X2 \AES_ENC/u0/u2/U69  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n1021 ), .ZN(\AES_ENC/u0/u2/n1042 ) );
NAND2_X2 \AES_ENC/u0/u2/U68  ( .A1(\AES_ENC/u0/u2/n1022 ), .A2(\AES_ENC/u0/u2/n1093 ), .ZN(\AES_ENC/u0/u2/n1039 ) );
NAND2_X2 \AES_ENC/u0/u2/U67  ( .A1(\AES_ENC/u0/u2/n1050 ), .A2(\AES_ENC/u0/u2/n1023 ), .ZN(\AES_ENC/u0/u2/n1038 ) );
NAND2_X2 \AES_ENC/u0/u2/U66  ( .A1(\AES_ENC/u0/u2/n1024 ), .A2(\AES_ENC/u0/u2/n1071 ), .ZN(\AES_ENC/u0/u2/n1037 ) );
AND2_X2 \AES_ENC/u0/u2/U60  ( .A1(\AES_ENC/u0/u2/n1030 ), .A2(\AES_ENC/u0/u2/n602 ), .ZN(\AES_ENC/u0/u2/n1078 ) );
NAND4_X2 \AES_ENC/u0/u2/U56  ( .A1(\AES_ENC/u0/u2/n1039 ), .A2(\AES_ENC/u0/u2/n1038 ), .A3(\AES_ENC/u0/u2/n1037 ), .A4(\AES_ENC/u0/u2/n1036 ), .ZN(\AES_ENC/u0/u2/n1040 ) );
NAND2_X2 \AES_ENC/u0/u2/U55  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n1040 ), .ZN(\AES_ENC/u0/u2/n1041 ) );
NAND4_X2 \AES_ENC/u0/u2/U54  ( .A1(\AES_ENC/u0/u2/n1044 ), .A2(\AES_ENC/u0/u2/n1043 ), .A3(\AES_ENC/u0/u2/n1042 ), .A4(\AES_ENC/u0/u2/n1041 ), .ZN(\AES_ENC/u0/subword[14] ) );
NAND2_X2 \AES_ENC/u0/u2/U53  ( .A1(\AES_ENC/u0/u2/n1072 ), .A2(\AES_ENC/u0/u2/n1045 ), .ZN(\AES_ENC/u0/u2/n1068 ) );
NAND2_X2 \AES_ENC/u0/u2/U52  ( .A1(\AES_ENC/u0/u2/n1046 ), .A2(\AES_ENC/u0/u2/n582 ), .ZN(\AES_ENC/u0/u2/n1067 ) );
NAND2_X2 \AES_ENC/u0/u2/U51  ( .A1(\AES_ENC/u0/u2/n1094 ), .A2(\AES_ENC/u0/u2/n1047 ), .ZN(\AES_ENC/u0/u2/n1066 ) );
NAND4_X2 \AES_ENC/u0/u2/U40  ( .A1(\AES_ENC/u0/u2/n1068 ), .A2(\AES_ENC/u0/u2/n1067 ), .A3(\AES_ENC/u0/u2/n1066 ), .A4(\AES_ENC/u0/u2/n1065 ), .ZN(\AES_ENC/u0/u2/n1069 ) );
NAND2_X2 \AES_ENC/u0/u2/U39  ( .A1(\AES_ENC/u0/u2/n1070 ), .A2(\AES_ENC/u0/u2/n1069 ), .ZN(\AES_ENC/u0/u2/n1135 ) );
NAND2_X2 \AES_ENC/u0/u2/U38  ( .A1(\AES_ENC/u0/u2/n1072 ), .A2(\AES_ENC/u0/u2/n1071 ), .ZN(\AES_ENC/u0/u2/n1088 ) );
NAND2_X2 \AES_ENC/u0/u2/U37  ( .A1(\AES_ENC/u0/u2/n1073 ), .A2(\AES_ENC/u0/u2/n595 ), .ZN(\AES_ENC/u0/u2/n1087 ) );
NAND4_X2 \AES_ENC/u0/u2/U28  ( .A1(\AES_ENC/u0/u2/n1088 ), .A2(\AES_ENC/u0/u2/n1087 ), .A3(\AES_ENC/u0/u2/n1086 ), .A4(\AES_ENC/u0/u2/n1085 ), .ZN(\AES_ENC/u0/u2/n1089 ) );
NAND2_X2 \AES_ENC/u0/u2/U27  ( .A1(\AES_ENC/u0/u2/n1090 ), .A2(\AES_ENC/u0/u2/n1089 ), .ZN(\AES_ENC/u0/u2/n1134 ) );
NAND2_X2 \AES_ENC/u0/u2/U26  ( .A1(\AES_ENC/u0/u2/n1091 ), .A2(\AES_ENC/u0/u2/n1093 ), .ZN(\AES_ENC/u0/u2/n1111 ) );
NAND2_X2 \AES_ENC/u0/u2/U25  ( .A1(\AES_ENC/u0/u2/n1092 ), .A2(\AES_ENC/u0/u2/n1120 ), .ZN(\AES_ENC/u0/u2/n1110 ) );
AND2_X2 \AES_ENC/u0/u2/U22  ( .A1(\AES_ENC/u0/u2/n1097 ), .A2(\AES_ENC/u0/u2/n1096 ), .ZN(\AES_ENC/u0/u2/n1098 ) );
NAND4_X2 \AES_ENC/u0/u2/U14  ( .A1(\AES_ENC/u0/u2/n1111 ), .A2(\AES_ENC/u0/u2/n1110 ), .A3(\AES_ENC/u0/u2/n1109 ), .A4(\AES_ENC/u0/u2/n1108 ), .ZN(\AES_ENC/u0/u2/n1112 ) );
NAND2_X2 \AES_ENC/u0/u2/U13  ( .A1(\AES_ENC/u0/u2/n1113 ), .A2(\AES_ENC/u0/u2/n1112 ), .ZN(\AES_ENC/u0/u2/n1133 ) );
NAND2_X2 \AES_ENC/u0/u2/U12  ( .A1(\AES_ENC/u0/u2/n1115 ), .A2(\AES_ENC/u0/u2/n1114 ), .ZN(\AES_ENC/u0/u2/n1129 ) );
OR2_X2 \AES_ENC/u0/u2/U11  ( .A1(\AES_ENC/u0/u2/n608 ), .A2(\AES_ENC/u0/u2/n1116 ), .ZN(\AES_ENC/u0/u2/n1128 ) );
NAND4_X2 \AES_ENC/u0/u2/U3  ( .A1(\AES_ENC/u0/u2/n1129 ), .A2(\AES_ENC/u0/u2/n1128 ), .A3(\AES_ENC/u0/u2/n1127 ), .A4(\AES_ENC/u0/u2/n1126 ), .ZN(\AES_ENC/u0/u2/n1130 ) );
NAND2_X2 \AES_ENC/u0/u2/U2  ( .A1(\AES_ENC/u0/u2/n1131 ), .A2(\AES_ENC/u0/u2/n1130 ), .ZN(\AES_ENC/u0/u2/n1132 ) );
NAND4_X2 \AES_ENC/u0/u2/U1  ( .A1(\AES_ENC/u0/u2/n1135 ), .A2(\AES_ENC/u0/u2/n1134 ), .A3(\AES_ENC/u0/u2/n1133 ), .A4(\AES_ENC/u0/u2/n1132 ), .ZN(\AES_ENC/u0/subword[15] ) );
INV_X4 \AES_ENC/u0/u3/U575  ( .A(\AES_ENC/w3[31] ), .ZN(\AES_ENC/u0/u3/n627 ) );
INV_X4 \AES_ENC/u0/u3/U574  ( .A(\AES_ENC/u0/u3/n1114 ), .ZN(\AES_ENC/u0/u3/n625 ) );
INV_X4 \AES_ENC/u0/u3/U573  ( .A(\AES_ENC/w3[28] ), .ZN(\AES_ENC/u0/u3/n624 ) );
INV_X4 \AES_ENC/u0/u3/U572  ( .A(\AES_ENC/u0/u3/n1025 ), .ZN(\AES_ENC/u0/u3/n622 ) );
INV_X4 \AES_ENC/u0/u3/U571  ( .A(\AES_ENC/u0/u3/n1120 ), .ZN(\AES_ENC/u0/u3/n620 ) );
INV_X4 \AES_ENC/u0/u3/U570  ( .A(\AES_ENC/u0/u3/n1121 ), .ZN(\AES_ENC/u0/u3/n619 ) );
INV_X4 \AES_ENC/u0/u3/U569  ( .A(\AES_ENC/u0/u3/n1048 ), .ZN(\AES_ENC/u0/u3/n618 ) );
INV_X4 \AES_ENC/u0/u3/U568  ( .A(\AES_ENC/u0/u3/n974 ), .ZN(\AES_ENC/u0/u3/n616 ) );
INV_X4 \AES_ENC/u0/u3/U567  ( .A(\AES_ENC/u0/u3/n794 ), .ZN(\AES_ENC/u0/u3/n614 ) );
INV_X4 \AES_ENC/u0/u3/U566  ( .A(\AES_ENC/w3[26] ), .ZN(\AES_ENC/u0/u3/n611 ) );
INV_X4 \AES_ENC/u0/u3/U565  ( .A(\AES_ENC/u0/u3/n800 ), .ZN(\AES_ENC/u0/u3/n610 ) );
INV_X4 \AES_ENC/u0/u3/U564  ( .A(\AES_ENC/u0/u3/n925 ), .ZN(\AES_ENC/u0/u3/n609 ) );
INV_X4 \AES_ENC/u0/u3/U563  ( .A(\AES_ENC/u0/u3/n779 ), .ZN(\AES_ENC/u0/u3/n607 ) );
INV_X4 \AES_ENC/u0/u3/U562  ( .A(\AES_ENC/u0/u3/n1022 ), .ZN(\AES_ENC/u0/u3/n603 ) );
INV_X4 \AES_ENC/u0/u3/U561  ( .A(\AES_ENC/u0/u3/n1102 ), .ZN(\AES_ENC/u0/u3/n602 ) );
INV_X4 \AES_ENC/u0/u3/U560  ( .A(\AES_ENC/u0/u3/n929 ), .ZN(\AES_ENC/u0/u3/n601 ) );
INV_X4 \AES_ENC/u0/u3/U559  ( .A(\AES_ENC/u0/u3/n1056 ), .ZN(\AES_ENC/u0/u3/n600 ) );
INV_X4 \AES_ENC/u0/u3/U558  ( .A(\AES_ENC/u0/u3/n1054 ), .ZN(\AES_ENC/u0/u3/n599 ) );
INV_X4 \AES_ENC/u0/u3/U557  ( .A(\AES_ENC/u0/u3/n881 ), .ZN(\AES_ENC/u0/u3/n598 ) );
INV_X4 \AES_ENC/u0/u3/U556  ( .A(\AES_ENC/u0/u3/n926 ), .ZN(\AES_ENC/u0/u3/n597 ) );
INV_X4 \AES_ENC/u0/u3/U555  ( .A(\AES_ENC/u0/u3/n977 ), .ZN(\AES_ENC/u0/u3/n595 ) );
INV_X4 \AES_ENC/u0/u3/U554  ( .A(\AES_ENC/u0/u3/n1031 ), .ZN(\AES_ENC/u0/u3/n594 ) );
INV_X4 \AES_ENC/u0/u3/U553  ( .A(\AES_ENC/u0/u3/n1103 ), .ZN(\AES_ENC/u0/u3/n593 ) );
INV_X4 \AES_ENC/u0/u3/U552  ( .A(\AES_ENC/u0/u3/n1009 ), .ZN(\AES_ENC/u0/u3/n592 ) );
INV_X4 \AES_ENC/u0/u3/U551  ( .A(\AES_ENC/u0/u3/n990 ), .ZN(\AES_ENC/u0/u3/n591 ) );
INV_X4 \AES_ENC/u0/u3/U550  ( .A(\AES_ENC/u0/u3/n1058 ), .ZN(\AES_ENC/u0/u3/n590 ) );
INV_X4 \AES_ENC/u0/u3/U549  ( .A(\AES_ENC/u0/u3/n1074 ), .ZN(\AES_ENC/u0/u3/n589 ) );
INV_X4 \AES_ENC/u0/u3/U548  ( .A(\AES_ENC/u0/u3/n1053 ), .ZN(\AES_ENC/u0/u3/n588 ) );
INV_X4 \AES_ENC/u0/u3/U547  ( .A(\AES_ENC/u0/u3/n826 ), .ZN(\AES_ENC/u0/u3/n587 ) );
INV_X4 \AES_ENC/u0/u3/U546  ( .A(\AES_ENC/u0/u3/n992 ), .ZN(\AES_ENC/u0/u3/n586 ) );
INV_X4 \AES_ENC/u0/u3/U545  ( .A(\AES_ENC/u0/u3/n821 ), .ZN(\AES_ENC/u0/u3/n585 ) );
INV_X4 \AES_ENC/u0/u3/U544  ( .A(\AES_ENC/u0/u3/n910 ), .ZN(\AES_ENC/u0/u3/n584 ) );
INV_X4 \AES_ENC/u0/u3/U543  ( .A(\AES_ENC/u0/u3/n906 ), .ZN(\AES_ENC/u0/u3/n583 ) );
INV_X4 \AES_ENC/u0/u3/U542  ( .A(\AES_ENC/u0/u3/n880 ), .ZN(\AES_ENC/u0/u3/n581 ) );
INV_X4 \AES_ENC/u0/u3/U541  ( .A(\AES_ENC/u0/u3/n1013 ), .ZN(\AES_ENC/u0/u3/n580 ) );
INV_X4 \AES_ENC/u0/u3/U540  ( .A(\AES_ENC/u0/u3/n1092 ), .ZN(\AES_ENC/u0/u3/n579 ) );
INV_X4 \AES_ENC/u0/u3/U539  ( .A(\AES_ENC/u0/u3/n824 ), .ZN(\AES_ENC/u0/u3/n578 ) );
INV_X4 \AES_ENC/u0/u3/U538  ( .A(\AES_ENC/u0/u3/n1091 ), .ZN(\AES_ENC/u0/u3/n577 ) );
INV_X4 \AES_ENC/u0/u3/U537  ( .A(\AES_ENC/u0/u3/n1080 ), .ZN(\AES_ENC/u0/u3/n576 ) );
INV_X4 \AES_ENC/u0/u3/U536  ( .A(\AES_ENC/u0/u3/n959 ), .ZN(\AES_ENC/u0/u3/n575 ) );
INV_X4 \AES_ENC/u0/u3/U535  ( .A(\AES_ENC/w3[24] ), .ZN(\AES_ENC/u0/u3/n574 ) );
NOR2_X2 \AES_ENC/u0/u3/U534  ( .A1(\AES_ENC/u0/u3/n574 ), .A2(\AES_ENC/w3[30] ), .ZN(\AES_ENC/u0/u3/n1070 ) );
NOR2_X2 \AES_ENC/u0/u3/U533  ( .A1(\AES_ENC/w3[24] ), .A2(\AES_ENC/w3[30] ),.ZN(\AES_ENC/u0/u3/n1090 ) );
NOR2_X2 \AES_ENC/u0/u3/U532  ( .A1(\AES_ENC/w3[28] ), .A2(\AES_ENC/w3[27] ),.ZN(\AES_ENC/u0/u3/n1025 ) );
NAND3_X2 \AES_ENC/u0/u3/U531  ( .A1(\AES_ENC/u0/u3/n679 ), .A2(\AES_ENC/u0/u3/n678 ), .A3(\AES_ENC/u0/u3/n677 ), .ZN(\AES_ENC/u0/subword[0] ) );
NOR2_X2 \AES_ENC/u0/u3/U530  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n765 ) );
NOR2_X2 \AES_ENC/u0/u3/U529  ( .A1(\AES_ENC/w3[28] ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n764 ) );
NOR2_X2 \AES_ENC/u0/u3/U528  ( .A1(\AES_ENC/u0/u3/n765 ), .A2(\AES_ENC/u0/u3/n764 ), .ZN(\AES_ENC/u0/u3/n766 ) );
NOR2_X2 \AES_ENC/u0/u3/U527  ( .A1(\AES_ENC/u0/u3/n766 ), .A2(\AES_ENC/u0/u3/n575 ), .ZN(\AES_ENC/u0/u3/n767 ) );
NOR2_X2 \AES_ENC/u0/u3/U526  ( .A1(\AES_ENC/u0/u3/n1117 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n707 ) );
NOR3_X2 \AES_ENC/u0/u3/U525  ( .A1(\AES_ENC/u0/u3/n627 ), .A2(\AES_ENC/w3[29] ), .A3(\AES_ENC/u0/u3/n704 ), .ZN(\AES_ENC/u0/u3/n706 ) );
NOR2_X2 \AES_ENC/u0/u3/U524  ( .A1(\AES_ENC/w3[28] ), .A2(\AES_ENC/u0/u3/n579 ), .ZN(\AES_ENC/u0/u3/n705 ) );
NOR3_X2 \AES_ENC/u0/u3/U523  ( .A1(\AES_ENC/u0/u3/n707 ), .A2(\AES_ENC/u0/u3/n706 ), .A3(\AES_ENC/u0/u3/n705 ), .ZN(\AES_ENC/u0/u3/n713 ) );
NOR4_X2 \AES_ENC/u0/u3/U522  ( .A1(\AES_ENC/u0/u3/n633 ), .A2(\AES_ENC/u0/u3/n632 ), .A3(\AES_ENC/u0/u3/n631 ), .A4(\AES_ENC/u0/u3/n630 ), .ZN(\AES_ENC/u0/u3/n634 ) );
NOR2_X2 \AES_ENC/u0/u3/U521  ( .A1(\AES_ENC/u0/u3/n629 ), .A2(\AES_ENC/u0/u3/n628 ), .ZN(\AES_ENC/u0/u3/n635 ) );
NAND3_X2 \AES_ENC/u0/u3/U520  ( .A1(\AES_ENC/w3[26] ), .A2(\AES_ENC/w3[31] ),.A3(\AES_ENC/u0/u3/n1059 ), .ZN(\AES_ENC/u0/u3/n636 ) );
INV_X4 \AES_ENC/u0/u3/U519  ( .A(\AES_ENC/w3[27] ), .ZN(\AES_ENC/u0/u3/n621 ) );
NOR2_X2 \AES_ENC/u0/u3/U518  ( .A1(\AES_ENC/w3[29] ), .A2(\AES_ENC/w3[26] ),.ZN(\AES_ENC/u0/u3/n974 ) );
NAND3_X2 \AES_ENC/u0/u3/U517  ( .A1(\AES_ENC/u0/u3/n652 ), .A2(\AES_ENC/u0/u3/n626 ), .A3(\AES_ENC/w3[31] ), .ZN(\AES_ENC/u0/u3/n653 ) );
NOR2_X2 \AES_ENC/u0/u3/U516  ( .A1(\AES_ENC/u0/u3/n611 ), .A2(\AES_ENC/w3[29] ), .ZN(\AES_ENC/u0/u3/n925 ) );
NOR2_X2 \AES_ENC/u0/u3/U515  ( .A1(\AES_ENC/u0/u3/n626 ), .A2(\AES_ENC/w3[26] ), .ZN(\AES_ENC/u0/u3/n1048 ) );
INV_X4 \AES_ENC/u0/u3/U512  ( .A(\AES_ENC/w3[29] ), .ZN(\AES_ENC/u0/u3/n626 ) );
NOR2_X2 \AES_ENC/u0/u3/U510  ( .A1(\AES_ENC/u0/u3/n611 ), .A2(\AES_ENC/w3[31] ), .ZN(\AES_ENC/u0/u3/n779 ) );
NOR2_X2 \AES_ENC/u0/u3/U509  ( .A1(\AES_ENC/w3[31] ), .A2(\AES_ENC/w3[26] ),.ZN(\AES_ENC/u0/u3/n794 ) );
NOR2_X2 \AES_ENC/u0/u3/U508  ( .A1(\AES_ENC/w3[28] ), .A2(\AES_ENC/w3[25] ),.ZN(\AES_ENC/u0/u3/n1102 ) );
INV_X4 \AES_ENC/u0/u3/U507  ( .A(\AES_ENC/u0/u3/n569 ), .ZN(\AES_ENC/u0/u3/n572 ) );
NOR2_X2 \AES_ENC/u0/u3/U506  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/w3[27] ), .ZN(\AES_ENC/u0/u3/n1053 ) );
NOR2_X2 \AES_ENC/u0/u3/U505  ( .A1(\AES_ENC/u0/u3/n607 ), .A2(\AES_ENC/w3[29] ), .ZN(\AES_ENC/u0/u3/n1024 ) );
NOR2_X2 \AES_ENC/u0/u3/U504  ( .A1(\AES_ENC/u0/u3/n625 ), .A2(\AES_ENC/w3[26] ), .ZN(\AES_ENC/u0/u3/n1093 ) );
NOR2_X2 \AES_ENC/u0/u3/U503  ( .A1(\AES_ENC/u0/u3/n614 ), .A2(\AES_ENC/w3[29] ), .ZN(\AES_ENC/u0/u3/n1094 ) );
NOR2_X2 \AES_ENC/u0/u3/U502  ( .A1(\AES_ENC/u0/u3/n624 ), .A2(\AES_ENC/w3[27] ), .ZN(\AES_ENC/u0/u3/n931 ) );
INV_X4 \AES_ENC/u0/u3/U501  ( .A(\AES_ENC/u0/u3/n570 ), .ZN(\AES_ENC/u0/u3/n573 ) );
NOR2_X2 \AES_ENC/u0/u3/U500  ( .A1(\AES_ENC/u0/u3/n622 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n1059 ) );
NOR2_X2 \AES_ENC/u0/u3/U499  ( .A1(\AES_ENC/u0/u3/n1053 ), .A2(\AES_ENC/u0/u3/n1095 ), .ZN(\AES_ENC/u0/u3/n639 ) );
NOR3_X2 \AES_ENC/u0/u3/U498  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n573 ), .A3(\AES_ENC/u0/u3/n1074 ), .ZN(\AES_ENC/u0/u3/n641 ) );
NOR2_X2 \AES_ENC/u0/u3/U497  ( .A1(\AES_ENC/u0/u3/n639 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n640 ) );
NOR2_X2 \AES_ENC/u0/u3/U496  ( .A1(\AES_ENC/u0/u3/n641 ), .A2(\AES_ENC/u0/u3/n640 ), .ZN(\AES_ENC/u0/u3/n646 ) );
NOR2_X2 \AES_ENC/u0/u3/U495  ( .A1(\AES_ENC/u0/u3/n826 ), .A2(\AES_ENC/u0/u3/n572 ), .ZN(\AES_ENC/u0/u3/n827 ) );
NOR3_X2 \AES_ENC/u0/u3/U494  ( .A1(\AES_ENC/u0/u3/n769 ), .A2(\AES_ENC/u0/u3/n768 ), .A3(\AES_ENC/u0/u3/n767 ), .ZN(\AES_ENC/u0/u3/n775 ) );
NOR2_X2 \AES_ENC/u0/u3/U492  ( .A1(\AES_ENC/w3[25] ), .A2(\AES_ENC/u0/u3/n623 ), .ZN(\AES_ENC/u0/u3/n913 ) );
NOR2_X2 \AES_ENC/u0/u3/U491  ( .A1(\AES_ENC/u0/u3/n913 ), .A2(\AES_ENC/u0/u3/n1091 ), .ZN(\AES_ENC/u0/u3/n914 ) );
NOR2_X2 \AES_ENC/u0/u3/U490  ( .A1(\AES_ENC/u0/u3/n1056 ), .A2(\AES_ENC/u0/u3/n1053 ), .ZN(\AES_ENC/u0/u3/n749 ) );
NOR2_X2 \AES_ENC/u0/u3/U489  ( .A1(\AES_ENC/u0/u3/n749 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n752 ) );
NOR3_X2 \AES_ENC/u0/u3/U488  ( .A1(\AES_ENC/u0/u3/n995 ), .A2(\AES_ENC/u0/u3/n586 ), .A3(\AES_ENC/u0/u3/n994 ), .ZN(\AES_ENC/u0/u3/n1002 ) );
NOR2_X2 \AES_ENC/u0/u3/U487  ( .A1(\AES_ENC/u0/u3/n909 ), .A2(\AES_ENC/u0/u3/n908 ), .ZN(\AES_ENC/u0/u3/n920 ) );
INV_X4 \AES_ENC/u0/u3/U486  ( .A(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n596 ) );
NOR2_X2 \AES_ENC/u0/u3/U483  ( .A1(\AES_ENC/u0/u3/n932 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n933 ) );
NOR2_X2 \AES_ENC/u0/u3/U482  ( .A1(\AES_ENC/u0/u3/n929 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n935 ) );
NOR2_X2 \AES_ENC/u0/u3/U480  ( .A1(\AES_ENC/u0/u3/n931 ), .A2(\AES_ENC/u0/u3/n930 ), .ZN(\AES_ENC/u0/u3/n934 ) );
NOR3_X2 \AES_ENC/u0/u3/U479  ( .A1(\AES_ENC/u0/u3/n935 ), .A2(\AES_ENC/u0/u3/n934 ), .A3(\AES_ENC/u0/u3/n933 ), .ZN(\AES_ENC/u0/u3/n936 ) );
OR2_X4 \AES_ENC/u0/u3/U478  ( .A1(\AES_ENC/u0/u3/n1094 ), .A2(\AES_ENC/u0/u3/n1093 ), .ZN(\AES_ENC/u0/u3/n571 ) );
AND2_X2 \AES_ENC/u0/u3/U477  ( .A1(\AES_ENC/u0/u3/n571 ), .A2(\AES_ENC/u0/u3/n1095 ), .ZN(\AES_ENC/u0/u3/n1101 ) );
NOR2_X2 \AES_ENC/u0/u3/U474  ( .A1(\AES_ENC/u0/u3/n1074 ), .A2(\AES_ENC/u0/u3/n931 ), .ZN(\AES_ENC/u0/u3/n796 ) );
NOR2_X2 \AES_ENC/u0/u3/U473  ( .A1(\AES_ENC/u0/u3/n796 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n797 ) );
NOR2_X2 \AES_ENC/u0/u3/U472  ( .A1(\AES_ENC/u0/u3/n1054 ), .A2(\AES_ENC/u0/u3/n1053 ), .ZN(\AES_ENC/u0/u3/n1055 ) );
NOR2_X2 \AES_ENC/u0/u3/U471  ( .A1(\AES_ENC/u0/u3/n572 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n949 ) );
NOR2_X2 \AES_ENC/u0/u3/U470  ( .A1(\AES_ENC/u0/u3/n1049 ), .A2(\AES_ENC/u0/u3/n618 ), .ZN(\AES_ENC/u0/u3/n1051 ) );
NOR2_X2 \AES_ENC/u0/u3/U469  ( .A1(\AES_ENC/u0/u3/n1051 ), .A2(\AES_ENC/u0/u3/n1050 ), .ZN(\AES_ENC/u0/u3/n1052 ) );
NOR2_X2 \AES_ENC/u0/u3/U468  ( .A1(\AES_ENC/u0/u3/n1052 ), .A2(\AES_ENC/u0/u3/n592 ), .ZN(\AES_ENC/u0/u3/n1064 ) );
NOR2_X2 \AES_ENC/u0/u3/U467  ( .A1(\AES_ENC/w3[25] ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n631 ) );
NOR2_X2 \AES_ENC/u0/u3/U466  ( .A1(\AES_ENC/u0/u3/n1025 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n980 ) );
NOR2_X2 \AES_ENC/u0/u3/U465  ( .A1(\AES_ENC/u0/u3/n1074 ), .A2(\AES_ENC/u0/u3/n1025 ), .ZN(\AES_ENC/u0/u3/n891 ) );
NOR2_X2 \AES_ENC/u0/u3/U464  ( .A1(\AES_ENC/u0/u3/n891 ), .A2(\AES_ENC/u0/u3/n609 ), .ZN(\AES_ENC/u0/u3/n894 ) );
NOR2_X2 \AES_ENC/u0/u3/U463  ( .A1(\AES_ENC/u0/u3/n1073 ), .A2(\AES_ENC/u0/u3/n1094 ), .ZN(\AES_ENC/u0/u3/n795 ) );
NOR2_X2 \AES_ENC/u0/u3/U462  ( .A1(\AES_ENC/u0/u3/n795 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n799 ) );
NOR2_X2 \AES_ENC/u0/u3/U461  ( .A1(\AES_ENC/u0/u3/n624 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n1075 ) );
NOR2_X2 \AES_ENC/u0/u3/U460  ( .A1(\AES_ENC/u0/u3/n624 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n822 ) );
NOR2_X2 \AES_ENC/u0/u3/U459  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n823 ) );
NOR2_X2 \AES_ENC/u0/u3/U458  ( .A1(\AES_ENC/u0/u3/n823 ), .A2(\AES_ENC/u0/u3/n822 ), .ZN(\AES_ENC/u0/u3/n825 ) );
NOR2_X2 \AES_ENC/u0/u3/U455  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n981 ) );
NOR2_X2 \AES_ENC/u0/u3/U448  ( .A1(\AES_ENC/u0/u3/n1102 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n643 ) );
NOR2_X2 \AES_ENC/u0/u3/U447  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n621 ), .ZN(\AES_ENC/u0/u3/n642 ) );
NOR2_X2 \AES_ENC/u0/u3/U442  ( .A1(\AES_ENC/u0/u3/n911 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n644 ) );
NOR4_X2 \AES_ENC/u0/u3/U441  ( .A1(\AES_ENC/u0/u3/n644 ), .A2(\AES_ENC/u0/u3/n643 ), .A3(\AES_ENC/u0/u3/n804 ), .A4(\AES_ENC/u0/u3/n642 ), .ZN(\AES_ENC/u0/u3/n645 ) );
NOR2_X2 \AES_ENC/u0/u3/U438  ( .A1(\AES_ENC/u0/u3/n1102 ), .A2(\AES_ENC/u0/u3/n910 ), .ZN(\AES_ENC/u0/u3/n932 ) );
NOR3_X2 \AES_ENC/u0/u3/U435  ( .A1(\AES_ENC/u0/u3/n623 ), .A2(\AES_ENC/w3[25] ), .A3(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n683 ) );
NOR2_X2 \AES_ENC/u0/u3/U434  ( .A1(\AES_ENC/u0/u3/n1102 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n755 ) );
INV_X4 \AES_ENC/u0/u3/U433  ( .A(\AES_ENC/u0/u3/n931 ), .ZN(\AES_ENC/u0/u3/n623 ) );
NOR2_X2 \AES_ENC/u0/u3/U428  ( .A1(\AES_ENC/u0/u3/n996 ), .A2(\AES_ENC/u0/u3/n931 ), .ZN(\AES_ENC/u0/u3/n704 ) );
NOR2_X2 \AES_ENC/u0/u3/U427  ( .A1(\AES_ENC/u0/u3/n1029 ), .A2(\AES_ENC/u0/u3/n1025 ), .ZN(\AES_ENC/u0/u3/n1079 ) );
NOR3_X2 \AES_ENC/u0/u3/U421  ( .A1(\AES_ENC/u0/u3/n589 ), .A2(\AES_ENC/u0/u3/n1025 ), .A3(\AES_ENC/u0/u3/n616 ), .ZN(\AES_ENC/u0/u3/n945 ) );
NOR2_X2 \AES_ENC/u0/u3/U420  ( .A1(\AES_ENC/u0/u3/n1072 ), .A2(\AES_ENC/u0/u3/n1094 ), .ZN(\AES_ENC/u0/u3/n930 ) );
NOR2_X2 \AES_ENC/u0/u3/U419  ( .A1(\AES_ENC/u0/u3/n931 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n743 ) );
NOR2_X2 \AES_ENC/u0/u3/U418  ( .A1(\AES_ENC/u0/u3/n931 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n685 ) );
NOR3_X2 \AES_ENC/u0/u3/U417  ( .A1(\AES_ENC/u0/u3/n610 ), .A2(\AES_ENC/u0/u3/n572 ), .A3(\AES_ENC/u0/u3/n575 ), .ZN(\AES_ENC/u0/u3/n962 ) );
NOR2_X2 \AES_ENC/u0/u3/U416  ( .A1(\AES_ENC/u0/u3/n626 ), .A2(\AES_ENC/u0/u3/n611 ), .ZN(\AES_ENC/u0/u3/n800 ) );
NOR3_X2 \AES_ENC/u0/u3/U415  ( .A1(\AES_ENC/u0/u3/n590 ), .A2(\AES_ENC/u0/u3/n627 ), .A3(\AES_ENC/u0/u3/n611 ), .ZN(\AES_ENC/u0/u3/n798 ) );
NOR3_X2 \AES_ENC/u0/u3/U414  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n572 ), .A3(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n694 ) );
NOR3_X2 \AES_ENC/u0/u3/U413  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n572 ), .A3(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n895 ) );
NOR3_X2 \AES_ENC/u0/u3/U410  ( .A1(\AES_ENC/u0/u3/n1008 ), .A2(\AES_ENC/u0/u3/n1007 ), .A3(\AES_ENC/u0/u3/n1006 ), .ZN(\AES_ENC/u0/u3/n1018 ) );
NOR4_X2 \AES_ENC/u0/u3/U409  ( .A1(\AES_ENC/u0/u3/n711 ), .A2(\AES_ENC/u0/u3/n710 ), .A3(\AES_ENC/u0/u3/n709 ), .A4(\AES_ENC/u0/u3/n708 ), .ZN(\AES_ENC/u0/u3/n712 ) );
NOR4_X2 \AES_ENC/u0/u3/U406  ( .A1(\AES_ENC/u0/u3/n806 ), .A2(\AES_ENC/u0/u3/n805 ), .A3(\AES_ENC/u0/u3/n804 ), .A4(\AES_ENC/u0/u3/n803 ), .ZN(\AES_ENC/u0/u3/n807 ) );
NOR3_X2 \AES_ENC/u0/u3/U405  ( .A1(\AES_ENC/u0/u3/n799 ), .A2(\AES_ENC/u0/u3/n798 ), .A3(\AES_ENC/u0/u3/n797 ), .ZN(\AES_ENC/u0/u3/n808 ) );
NOR2_X2 \AES_ENC/u0/u3/U404  ( .A1(\AES_ENC/u0/u3/n669 ), .A2(\AES_ENC/u0/u3/n668 ), .ZN(\AES_ENC/u0/u3/n673 ) );
NOR4_X2 \AES_ENC/u0/u3/U403  ( .A1(\AES_ENC/u0/u3/n946 ), .A2(\AES_ENC/u0/u3/n1046 ), .A3(\AES_ENC/u0/u3/n671 ), .A4(\AES_ENC/u0/u3/n670 ), .ZN(\AES_ENC/u0/u3/n672 ) );
NOR4_X2 \AES_ENC/u0/u3/U401  ( .A1(\AES_ENC/u0/u3/n843 ), .A2(\AES_ENC/u0/u3/n842 ), .A3(\AES_ENC/u0/u3/n841 ), .A4(\AES_ENC/u0/u3/n840 ), .ZN(\AES_ENC/u0/u3/n844 ) );
NOR3_X2 \AES_ENC/u0/u3/U400  ( .A1(\AES_ENC/u0/u3/n1101 ), .A2(\AES_ENC/u0/u3/n1100 ), .A3(\AES_ENC/u0/u3/n1099 ), .ZN(\AES_ENC/u0/u3/n1109 ) );
NOR3_X2 \AES_ENC/u0/u3/U399  ( .A1(\AES_ENC/u0/u3/n743 ), .A2(\AES_ENC/u0/u3/n742 ), .A3(\AES_ENC/u0/u3/n741 ), .ZN(\AES_ENC/u0/u3/n744 ) );
NOR2_X2 \AES_ENC/u0/u3/U398  ( .A1(\AES_ENC/u0/u3/n697 ), .A2(\AES_ENC/u0/u3/n658 ), .ZN(\AES_ENC/u0/u3/n659 ) );
NOR3_X2 \AES_ENC/u0/u3/U397  ( .A1(\AES_ENC/u0/u3/n959 ), .A2(\AES_ENC/u0/u3/n572 ), .A3(\AES_ENC/u0/u3/n609 ), .ZN(\AES_ENC/u0/u3/n768 ) );
NOR2_X2 \AES_ENC/u0/u3/U396  ( .A1(\AES_ENC/u0/u3/n1078 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n1033 ) );
NOR2_X2 \AES_ENC/u0/u3/U393  ( .A1(\AES_ENC/u0/u3/n1031 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n1032 ) );
NOR3_X2 \AES_ENC/u0/u3/U390  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n1025 ), .A3(\AES_ENC/u0/u3/n1074 ), .ZN(\AES_ENC/u0/u3/n1035 ) );
NOR4_X2 \AES_ENC/u0/u3/U389  ( .A1(\AES_ENC/u0/u3/n1035 ), .A2(\AES_ENC/u0/u3/n1034 ), .A3(\AES_ENC/u0/u3/n1033 ), .A4(\AES_ENC/u0/u3/n1032 ), .ZN(\AES_ENC/u0/u3/n1036 ) );
NOR2_X2 \AES_ENC/u0/u3/U388  ( .A1(\AES_ENC/u0/u3/n598 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n885 ) );
NOR2_X2 \AES_ENC/u0/u3/U387  ( .A1(\AES_ENC/u0/u3/n623 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n882 ) );
NOR2_X2 \AES_ENC/u0/u3/U386  ( .A1(\AES_ENC/u0/u3/n1053 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n884 ) );
NOR4_X2 \AES_ENC/u0/u3/U385  ( .A1(\AES_ENC/u0/u3/n885 ), .A2(\AES_ENC/u0/u3/n884 ), .A3(\AES_ENC/u0/u3/n883 ), .A4(\AES_ENC/u0/u3/n882 ), .ZN(\AES_ENC/u0/u3/n886 ) );
NOR2_X2 \AES_ENC/u0/u3/U384  ( .A1(\AES_ENC/u0/u3/n825 ), .A2(\AES_ENC/u0/u3/n578 ), .ZN(\AES_ENC/u0/u3/n830 ) );
NOR2_X2 \AES_ENC/u0/u3/U383  ( .A1(\AES_ENC/u0/u3/n827 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n829 ) );
NOR2_X2 \AES_ENC/u0/u3/U382  ( .A1(\AES_ENC/u0/u3/n572 ), .A2(\AES_ENC/u0/u3/n579 ), .ZN(\AES_ENC/u0/u3/n828 ) );
NOR4_X2 \AES_ENC/u0/u3/U374  ( .A1(\AES_ENC/u0/u3/n831 ), .A2(\AES_ENC/u0/u3/n830 ), .A3(\AES_ENC/u0/u3/n829 ), .A4(\AES_ENC/u0/u3/n828 ), .ZN(\AES_ENC/u0/u3/n832 ) );
NOR2_X2 \AES_ENC/u0/u3/U373  ( .A1(\AES_ENC/u0/u3/n598 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n1107 ) );
NOR2_X2 \AES_ENC/u0/u3/U372  ( .A1(\AES_ENC/u0/u3/n1102 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n1106 ) );
NOR2_X2 \AES_ENC/u0/u3/U370  ( .A1(\AES_ENC/u0/u3/n1103 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n1105 ) );
NOR4_X2 \AES_ENC/u0/u3/U369  ( .A1(\AES_ENC/u0/u3/n1107 ), .A2(\AES_ENC/u0/u3/n1106 ), .A3(\AES_ENC/u0/u3/n1105 ), .A4(\AES_ENC/u0/u3/n1104 ), .ZN(\AES_ENC/u0/u3/n1108 ) );
NOR3_X2 \AES_ENC/u0/u3/U368  ( .A1(\AES_ENC/u0/u3/n959 ), .A2(\AES_ENC/u0/u3/n621 ), .A3(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n963 ) );
NOR2_X2 \AES_ENC/u0/u3/U367  ( .A1(\AES_ENC/u0/u3/n626 ), .A2(\AES_ENC/u0/u3/n627 ), .ZN(\AES_ENC/u0/u3/n1114 ) );
NOR3_X2 \AES_ENC/u0/u3/U366  ( .A1(\AES_ENC/u0/u3/n910 ), .A2(\AES_ENC/u0/u3/n1059 ), .A3(\AES_ENC/u0/u3/n611 ), .ZN(\AES_ENC/u0/u3/n1115 ) );
INV_X4 \AES_ENC/u0/u3/U365  ( .A(\AES_ENC/u0/u3/n1024 ), .ZN(\AES_ENC/u0/u3/n606 ) );
INV_X4 \AES_ENC/u0/u3/U364  ( .A(\AES_ENC/u0/u3/n1094 ), .ZN(\AES_ENC/u0/u3/n613 ) );
NOR2_X2 \AES_ENC/u0/u3/U363  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n931 ), .ZN(\AES_ENC/u0/u3/n1100 ) );
NOR2_X2 \AES_ENC/u0/u3/U354  ( .A1(\AES_ENC/u0/u3/n569 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n929 ) );
NOR2_X2 \AES_ENC/u0/u3/U353  ( .A1(\AES_ENC/u0/u3/n620 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n926 ) );
INV_X4 \AES_ENC/u0/u3/U352  ( .A(\AES_ENC/u0/u3/n1093 ), .ZN(\AES_ENC/u0/u3/n617 ) );
NOR2_X2 \AES_ENC/u0/u3/U351  ( .A1(\AES_ENC/u0/u3/n572 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n1095 ) );
NOR2_X2 \AES_ENC/u0/u3/U350  ( .A1(\AES_ENC/u0/u3/n609 ), .A2(\AES_ENC/u0/u3/n627 ), .ZN(\AES_ENC/u0/u3/n1010 ) );
NOR2_X2 \AES_ENC/u0/u3/U349  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n1103 ) );
NOR2_X2 \AES_ENC/u0/u3/U348  ( .A1(\AES_ENC/w3[25] ), .A2(\AES_ENC/u0/u3/n1120 ), .ZN(\AES_ENC/u0/u3/n1022 ) );
NOR2_X2 \AES_ENC/u0/u3/U347  ( .A1(\AES_ENC/u0/u3/n619 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n911 ) );
NOR2_X2 \AES_ENC/u0/u3/U346  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/u0/u3/n1025 ), .ZN(\AES_ENC/u0/u3/n826 ) );
NOR2_X2 \AES_ENC/u0/u3/U345  ( .A1(\AES_ENC/u0/u3/n626 ), .A2(\AES_ENC/u0/u3/n607 ), .ZN(\AES_ENC/u0/u3/n1072 ) );
NOR2_X2 \AES_ENC/u0/u3/U338  ( .A1(\AES_ENC/u0/u3/n627 ), .A2(\AES_ENC/u0/u3/n616 ), .ZN(\AES_ENC/u0/u3/n956 ) );
NOR2_X2 \AES_ENC/u0/u3/U335  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/u0/u3/n624 ), .ZN(\AES_ENC/u0/u3/n1121 ) );
NOR2_X2 \AES_ENC/u0/u3/U329  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/u0/u3/n624 ), .ZN(\AES_ENC/u0/u3/n1058 ) );
NOR2_X2 \AES_ENC/u0/u3/U328  ( .A1(\AES_ENC/u0/u3/n625 ), .A2(\AES_ENC/u0/u3/n611 ), .ZN(\AES_ENC/u0/u3/n1073 ) );
NOR2_X2 \AES_ENC/u0/u3/U327  ( .A1(\AES_ENC/w3[25] ), .A2(\AES_ENC/u0/u3/n1025 ), .ZN(\AES_ENC/u0/u3/n1054 ) );
NOR2_X2 \AES_ENC/u0/u3/U325  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/u0/u3/n931 ), .ZN(\AES_ENC/u0/u3/n1029 ) );
NOR2_X2 \AES_ENC/u0/u3/U324  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n1056 ) );
NOR2_X2 \AES_ENC/u0/u3/U319  ( .A1(\AES_ENC/u0/u3/n614 ), .A2(\AES_ENC/u0/u3/n626 ), .ZN(\AES_ENC/u0/u3/n1050 ) );
NOR2_X2 \AES_ENC/u0/u3/U318  ( .A1(\AES_ENC/u0/u3/n1121 ), .A2(\AES_ENC/u0/u3/n1025 ), .ZN(\AES_ENC/u0/u3/n1120 ) );
NOR2_X2 \AES_ENC/u0/u3/U317  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/u0/u3/n572 ), .ZN(\AES_ENC/u0/u3/n1074 ) );
NOR2_X2 \AES_ENC/u0/u3/U316  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n584 ), .ZN(\AES_ENC/u0/u3/n838 ) );
NOR2_X2 \AES_ENC/u0/u3/U315  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n602 ), .ZN(\AES_ENC/u0/u3/n837 ) );
NOR2_X2 \AES_ENC/u0/u3/U314  ( .A1(\AES_ENC/u0/u3/n838 ), .A2(\AES_ENC/u0/u3/n837 ), .ZN(\AES_ENC/u0/u3/n845 ) );
NOR2_X2 \AES_ENC/u0/u3/U312  ( .A1(\AES_ENC/u0/u3/n1058 ), .A2(\AES_ENC/u0/u3/n1054 ), .ZN(\AES_ENC/u0/u3/n878 ) );
NOR2_X2 \AES_ENC/u0/u3/U311  ( .A1(\AES_ENC/u0/u3/n878 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n879 ) );
NOR2_X2 \AES_ENC/u0/u3/U310  ( .A1(\AES_ENC/u0/u3/n880 ), .A2(\AES_ENC/u0/u3/n879 ), .ZN(\AES_ENC/u0/u3/n887 ) );
NOR3_X2 \AES_ENC/u0/u3/U309  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n1091 ), .A3(\AES_ENC/u0/u3/n1022 ), .ZN(\AES_ENC/u0/u3/n720 ) );
NOR3_X2 \AES_ENC/u0/u3/U303  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n1054 ), .A3(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n719 ) );
NOR2_X2 \AES_ENC/u0/u3/U302  ( .A1(\AES_ENC/u0/u3/n720 ), .A2(\AES_ENC/u0/u3/n719 ), .ZN(\AES_ENC/u0/u3/n726 ) );
NOR2_X2 \AES_ENC/u0/u3/U300  ( .A1(\AES_ENC/u0/u3/n614 ), .A2(\AES_ENC/u0/u3/n591 ), .ZN(\AES_ENC/u0/u3/n865 ) );
NOR2_X2 \AES_ENC/u0/u3/U299  ( .A1(\AES_ENC/u0/u3/n1059 ), .A2(\AES_ENC/u0/u3/n1058 ), .ZN(\AES_ENC/u0/u3/n1060 ) );
NOR2_X2 \AES_ENC/u0/u3/U298  ( .A1(\AES_ENC/u0/u3/n1095 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n668 ) );
NOR2_X2 \AES_ENC/u0/u3/U297  ( .A1(\AES_ENC/u0/u3/n826 ), .A2(\AES_ENC/u0/u3/n573 ), .ZN(\AES_ENC/u0/u3/n750 ) );
NOR2_X2 \AES_ENC/u0/u3/U296  ( .A1(\AES_ENC/u0/u3/n750 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n751 ) );
NOR2_X2 \AES_ENC/u0/u3/U295  ( .A1(\AES_ENC/u0/u3/n907 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n908 ) );
NOR2_X2 \AES_ENC/u0/u3/U294  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n588 ), .ZN(\AES_ENC/u0/u3/n957 ) );
NOR2_X2 \AES_ENC/u0/u3/U293  ( .A1(\AES_ENC/u0/u3/n990 ), .A2(\AES_ENC/u0/u3/n926 ), .ZN(\AES_ENC/u0/u3/n780 ) );
NOR2_X2 \AES_ENC/u0/u3/U292  ( .A1(\AES_ENC/u0/u3/n1022 ), .A2(\AES_ENC/u0/u3/n1058 ), .ZN(\AES_ENC/u0/u3/n740 ) );
NOR2_X2 \AES_ENC/u0/u3/U291  ( .A1(\AES_ENC/u0/u3/n740 ), .A2(\AES_ENC/u0/u3/n616 ), .ZN(\AES_ENC/u0/u3/n742 ) );
NOR2_X2 \AES_ENC/u0/u3/U290  ( .A1(\AES_ENC/u0/u3/n1098 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n1099 ) );
NOR2_X2 \AES_ENC/u0/u3/U284  ( .A1(\AES_ENC/u0/u3/n1120 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n993 ) );
NOR2_X2 \AES_ENC/u0/u3/U283  ( .A1(\AES_ENC/u0/u3/n993 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n994 ) );
NOR2_X2 \AES_ENC/u0/u3/U282  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n620 ), .ZN(\AES_ENC/u0/u3/n1026 ) );
NOR2_X2 \AES_ENC/u0/u3/U281  ( .A1(\AES_ENC/u0/u3/n573 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n1027 ) );
NOR2_X2 \AES_ENC/u0/u3/U280  ( .A1(\AES_ENC/u0/u3/n1027 ), .A2(\AES_ENC/u0/u3/n1026 ), .ZN(\AES_ENC/u0/u3/n1028 ) );
NOR2_X2 \AES_ENC/u0/u3/U279  ( .A1(\AES_ENC/u0/u3/n1029 ), .A2(\AES_ENC/u0/u3/n1028 ), .ZN(\AES_ENC/u0/u3/n1034 ) );
NOR2_X2 \AES_ENC/u0/u3/U273  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n1071 ), .ZN(\AES_ENC/u0/u3/n669 ) );
NOR2_X2 \AES_ENC/u0/u3/U272  ( .A1(\AES_ENC/u0/u3/n1056 ), .A2(\AES_ENC/u0/u3/n990 ), .ZN(\AES_ENC/u0/u3/n991 ) );
NOR2_X2 \AES_ENC/u0/u3/U271  ( .A1(\AES_ENC/u0/u3/n991 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n995 ) );
NOR4_X2 \AES_ENC/u0/u3/U270  ( .A1(\AES_ENC/u0/u3/n757 ), .A2(\AES_ENC/u0/u3/n756 ), .A3(\AES_ENC/u0/u3/n755 ), .A4(\AES_ENC/u0/u3/n754 ), .ZN(\AES_ENC/u0/u3/n758 ) );
NOR2_X2 \AES_ENC/u0/u3/U269  ( .A1(\AES_ENC/u0/u3/n752 ), .A2(\AES_ENC/u0/u3/n751 ), .ZN(\AES_ENC/u0/u3/n759 ) );
NOR2_X2 \AES_ENC/u0/u3/U268  ( .A1(\AES_ENC/u0/u3/n607 ), .A2(\AES_ENC/u0/u3/n590 ), .ZN(\AES_ENC/u0/u3/n1008 ) );
NOR2_X2 \AES_ENC/u0/u3/U267  ( .A1(\AES_ENC/u0/u3/n606 ), .A2(\AES_ENC/u0/u3/n906 ), .ZN(\AES_ENC/u0/u3/n741 ) );
NOR2_X2 \AES_ENC/u0/u3/U263  ( .A1(\AES_ENC/u0/u3/n1054 ), .A2(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n763 ) );
NOR2_X2 \AES_ENC/u0/u3/U262  ( .A1(\AES_ENC/u0/u3/n763 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n769 ) );
NOR2_X2 \AES_ENC/u0/u3/U258  ( .A1(\AES_ENC/u0/u3/n839 ), .A2(\AES_ENC/u0/u3/n582 ), .ZN(\AES_ENC/u0/u3/n693 ) );
NOR2_X2 \AES_ENC/u0/u3/U255  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n577 ), .ZN(\AES_ENC/u0/u3/n1007 ) );
NOR2_X2 \AES_ENC/u0/u3/U254  ( .A1(\AES_ENC/u0/u3/n609 ), .A2(\AES_ENC/u0/u3/n580 ), .ZN(\AES_ENC/u0/u3/n1123 ) );
NOR2_X2 \AES_ENC/u0/u3/U253  ( .A1(\AES_ENC/u0/u3/n780 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n784 ) );
NOR2_X2 \AES_ENC/u0/u3/U252  ( .A1(\AES_ENC/u0/u3/n1117 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n782 ) );
NOR2_X2 \AES_ENC/u0/u3/U251  ( .A1(\AES_ENC/u0/u3/n781 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n783 ) );
NOR4_X2 \AES_ENC/u0/u3/U250  ( .A1(\AES_ENC/u0/u3/n880 ), .A2(\AES_ENC/u0/u3/n784 ), .A3(\AES_ENC/u0/u3/n783 ), .A4(\AES_ENC/u0/u3/n782 ), .ZN(\AES_ENC/u0/u3/n785 ) );
NOR2_X2 \AES_ENC/u0/u3/U243  ( .A1(\AES_ENC/u0/u3/n609 ), .A2(\AES_ENC/u0/u3/n590 ), .ZN(\AES_ENC/u0/u3/n710 ) );
INV_X4 \AES_ENC/u0/u3/U242  ( .A(\AES_ENC/u0/u3/n1029 ), .ZN(\AES_ENC/u0/u3/n582 ) );
NOR2_X2 \AES_ENC/u0/u3/U241  ( .A1(\AES_ENC/u0/u3/n593 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n1125 ) );
NOR2_X2 \AES_ENC/u0/u3/U240  ( .A1(\AES_ENC/u0/u3/n616 ), .A2(\AES_ENC/u0/u3/n580 ), .ZN(\AES_ENC/u0/u3/n771 ) );
NOR2_X2 \AES_ENC/u0/u3/U239  ( .A1(\AES_ENC/u0/u3/n616 ), .A2(\AES_ENC/u0/u3/n597 ), .ZN(\AES_ENC/u0/u3/n883 ) );
NOR2_X2 \AES_ENC/u0/u3/U238  ( .A1(\AES_ENC/u0/u3/n911 ), .A2(\AES_ENC/u0/u3/n910 ), .ZN(\AES_ENC/u0/u3/n912 ) );
NOR2_X2 \AES_ENC/u0/u3/U237  ( .A1(\AES_ENC/u0/u3/n912 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n916 ) );
NOR2_X2 \AES_ENC/u0/u3/U236  ( .A1(\AES_ENC/u0/u3/n990 ), .A2(\AES_ENC/u0/u3/n929 ), .ZN(\AES_ENC/u0/u3/n892 ) );
NOR2_X2 \AES_ENC/u0/u3/U235  ( .A1(\AES_ENC/u0/u3/n892 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n893 ) );
NOR2_X2 \AES_ENC/u0/u3/U234  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n602 ), .ZN(\AES_ENC/u0/u3/n950 ) );
NOR2_X2 \AES_ENC/u0/u3/U229  ( .A1(\AES_ENC/u0/u3/n1079 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n1082 ) );
NOR2_X2 \AES_ENC/u0/u3/U228  ( .A1(\AES_ENC/u0/u3/n910 ), .A2(\AES_ENC/u0/u3/n1056 ), .ZN(\AES_ENC/u0/u3/n941 ) );
NOR2_X2 \AES_ENC/u0/u3/U227  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n1077 ), .ZN(\AES_ENC/u0/u3/n841 ) );
NOR2_X2 \AES_ENC/u0/u3/U226  ( .A1(\AES_ENC/u0/u3/n623 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n630 ) );
NOR2_X2 \AES_ENC/u0/u3/U225  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n602 ), .ZN(\AES_ENC/u0/u3/n806 ) );
NOR2_X2 \AES_ENC/u0/u3/U223  ( .A1(\AES_ENC/u0/u3/n623 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n948 ) );
NOR2_X2 \AES_ENC/u0/u3/U222  ( .A1(\AES_ENC/u0/u3/n606 ), .A2(\AES_ENC/u0/u3/n582 ), .ZN(\AES_ENC/u0/u3/n1104 ) );
NOR2_X2 \AES_ENC/u0/u3/U221  ( .A1(\AES_ENC/u0/u3/n1121 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n1122 ) );
NOR2_X2 \AES_ENC/u0/u3/U217  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n1023 ), .ZN(\AES_ENC/u0/u3/n756 ) );
NOR2_X2 \AES_ENC/u0/u3/U213  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n602 ), .ZN(\AES_ENC/u0/u3/n870 ) );
NOR2_X2 \AES_ENC/u0/u3/U212  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n569 ), .ZN(\AES_ENC/u0/u3/n947 ) );
NOR2_X2 \AES_ENC/u0/u3/U211  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n1077 ), .ZN(\AES_ENC/u0/u3/n1084 ) );
NOR2_X2 \AES_ENC/u0/u3/U210  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n855 ), .ZN(\AES_ENC/u0/u3/n709 ) );
NOR2_X2 \AES_ENC/u0/u3/U209  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n589 ), .ZN(\AES_ENC/u0/u3/n868 ) );
NOR2_X2 \AES_ENC/u0/u3/U208  ( .A1(\AES_ENC/u0/u3/n1120 ), .A2(\AES_ENC/u0/u3/n839 ), .ZN(\AES_ENC/u0/u3/n842 ) );
NOR2_X2 \AES_ENC/u0/u3/U207  ( .A1(\AES_ENC/u0/u3/n1120 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n1124 ) );
NOR2_X2 \AES_ENC/u0/u3/U201  ( .A1(\AES_ENC/u0/u3/n1120 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n696 ) );
NOR2_X2 \AES_ENC/u0/u3/U200  ( .A1(\AES_ENC/u0/u3/n1074 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n1076 ) );
NOR2_X2 \AES_ENC/u0/u3/U199  ( .A1(\AES_ENC/u0/u3/n1074 ), .A2(\AES_ENC/u0/u3/n620 ), .ZN(\AES_ENC/u0/u3/n781 ) );
NOR3_X2 \AES_ENC/u0/u3/U198  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n1056 ), .A3(\AES_ENC/u0/u3/n990 ), .ZN(\AES_ENC/u0/u3/n979 ) );
NOR3_X2 \AES_ENC/u0/u3/U197  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n1058 ), .A3(\AES_ENC/u0/u3/n1059 ), .ZN(\AES_ENC/u0/u3/n854 ) );
NOR2_X2 \AES_ENC/u0/u3/U196  ( .A1(\AES_ENC/u0/u3/n996 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n869 ) );
NOR2_X2 \AES_ENC/u0/u3/U195  ( .A1(\AES_ENC/u0/u3/n1056 ), .A2(\AES_ENC/u0/u3/n1074 ), .ZN(\AES_ENC/u0/u3/n1057 ) );
NOR3_X2 \AES_ENC/u0/u3/U194  ( .A1(\AES_ENC/u0/u3/n607 ), .A2(\AES_ENC/u0/u3/n1120 ), .A3(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n978 ) );
NOR2_X2 \AES_ENC/u0/u3/U187  ( .A1(\AES_ENC/u0/u3/n996 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n998 ) );
NOR2_X2 \AES_ENC/u0/u3/U186  ( .A1(\AES_ENC/u0/u3/n996 ), .A2(\AES_ENC/u0/u3/n911 ), .ZN(\AES_ENC/u0/u3/n1116 ) );
NOR2_X2 \AES_ENC/u0/u3/U185  ( .A1(\AES_ENC/u0/u3/n1074 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n754 ) );
NOR2_X2 \AES_ENC/u0/u3/U184  ( .A1(\AES_ENC/u0/u3/n926 ), .A2(\AES_ENC/u0/u3/n1103 ), .ZN(\AES_ENC/u0/u3/n977 ) );
NOR2_X2 \AES_ENC/u0/u3/U183  ( .A1(\AES_ENC/u0/u3/n839 ), .A2(\AES_ENC/u0/u3/n824 ), .ZN(\AES_ENC/u0/u3/n1092 ) );
NOR2_X2 \AES_ENC/u0/u3/U182  ( .A1(\AES_ENC/u0/u3/n573 ), .A2(\AES_ENC/u0/u3/n1074 ), .ZN(\AES_ENC/u0/u3/n684 ) );
NOR2_X2 \AES_ENC/u0/u3/U181  ( .A1(\AES_ENC/u0/u3/n826 ), .A2(\AES_ENC/u0/u3/n1059 ), .ZN(\AES_ENC/u0/u3/n907 ) );
NOR3_X2 \AES_ENC/u0/u3/U180  ( .A1(\AES_ENC/u0/u3/n625 ), .A2(\AES_ENC/u0/u3/n1115 ), .A3(\AES_ENC/u0/u3/n585 ), .ZN(\AES_ENC/u0/u3/n831 ) );
NOR3_X2 \AES_ENC/u0/u3/U174  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n1056 ), .A3(\AES_ENC/u0/u3/n990 ), .ZN(\AES_ENC/u0/u3/n896 ) );
NOR3_X2 \AES_ENC/u0/u3/U173  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n573 ), .A3(\AES_ENC/u0/u3/n1013 ), .ZN(\AES_ENC/u0/u3/n670 ) );
NOR3_X2 \AES_ENC/u0/u3/U172  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n1091 ), .A3(\AES_ENC/u0/u3/n1022 ), .ZN(\AES_ENC/u0/u3/n843 ) );
NOR2_X2 \AES_ENC/u0/u3/U171  ( .A1(\AES_ENC/u0/u3/n1029 ), .A2(\AES_ENC/u0/u3/n1095 ), .ZN(\AES_ENC/u0/u3/n735 ) );
NOR4_X2 \AES_ENC/u0/u3/U170  ( .A1(\AES_ENC/u0/u3/n983 ), .A2(\AES_ENC/u0/u3/n698 ), .A3(\AES_ENC/u0/u3/n697 ), .A4(\AES_ENC/u0/u3/n696 ), .ZN(\AES_ENC/u0/u3/n699 ) );
NOR3_X2 \AES_ENC/u0/u3/U169  ( .A1(\AES_ENC/u0/u3/n695 ), .A2(\AES_ENC/u0/u3/n694 ), .A3(\AES_ENC/u0/u3/n693 ), .ZN(\AES_ENC/u0/u3/n700 ) );
NOR2_X2 \AES_ENC/u0/u3/U168  ( .A1(\AES_ENC/u0/u3/n1100 ), .A2(\AES_ENC/u0/u3/n854 ), .ZN(\AES_ENC/u0/u3/n860 ) );
NAND3_X2 \AES_ENC/u0/u3/U162  ( .A1(\AES_ENC/u0/u3/n569 ), .A2(\AES_ENC/u0/u3/n582 ), .A3(\AES_ENC/u0/u3/n681 ), .ZN(\AES_ENC/u0/u3/n691 ) );
NOR2_X2 \AES_ENC/u0/u3/U161  ( .A1(\AES_ENC/u0/u3/n683 ), .A2(\AES_ENC/u0/u3/n682 ), .ZN(\AES_ENC/u0/u3/n690 ) );
NOR4_X2 \AES_ENC/u0/u3/U160  ( .A1(\AES_ENC/u0/u3/n896 ), .A2(\AES_ENC/u0/u3/n895 ), .A3(\AES_ENC/u0/u3/n894 ), .A4(\AES_ENC/u0/u3/n893 ), .ZN(\AES_ENC/u0/u3/n897 ) );
NOR2_X2 \AES_ENC/u0/u3/U159  ( .A1(\AES_ENC/u0/u3/n866 ), .A2(\AES_ENC/u0/u3/n865 ), .ZN(\AES_ENC/u0/u3/n872 ) );
NOR4_X2 \AES_ENC/u0/u3/U158  ( .A1(\AES_ENC/u0/u3/n870 ), .A2(\AES_ENC/u0/u3/n869 ), .A3(\AES_ENC/u0/u3/n868 ), .A4(\AES_ENC/u0/u3/n867 ), .ZN(\AES_ENC/u0/u3/n871 ) );
NOR4_X2 \AES_ENC/u0/u3/U157  ( .A1(\AES_ENC/u0/u3/n963 ), .A2(\AES_ENC/u0/u3/n962 ), .A3(\AES_ENC/u0/u3/n961 ), .A4(\AES_ENC/u0/u3/n960 ), .ZN(\AES_ENC/u0/u3/n964 ) );
NOR2_X2 \AES_ENC/u0/u3/U156  ( .A1(\AES_ENC/u0/u3/n958 ), .A2(\AES_ENC/u0/u3/n957 ), .ZN(\AES_ENC/u0/u3/n965 ) );
NOR4_X2 \AES_ENC/u0/u3/U155  ( .A1(\AES_ENC/u0/u3/n950 ), .A2(\AES_ENC/u0/u3/n949 ), .A3(\AES_ENC/u0/u3/n948 ), .A4(\AES_ENC/u0/u3/n947 ), .ZN(\AES_ENC/u0/u3/n951 ) );
NOR2_X2 \AES_ENC/u0/u3/U154  ( .A1(\AES_ENC/u0/u3/n946 ), .A2(\AES_ENC/u0/u3/n945 ), .ZN(\AES_ENC/u0/u3/n952 ) );
NOR4_X2 \AES_ENC/u0/u3/U153  ( .A1(\AES_ENC/u0/u3/n983 ), .A2(\AES_ENC/u0/u3/n982 ), .A3(\AES_ENC/u0/u3/n981 ), .A4(\AES_ENC/u0/u3/n980 ), .ZN(\AES_ENC/u0/u3/n984 ) );
NOR2_X2 \AES_ENC/u0/u3/U152  ( .A1(\AES_ENC/u0/u3/n979 ), .A2(\AES_ENC/u0/u3/n978 ), .ZN(\AES_ENC/u0/u3/n985 ) );
NOR4_X2 \AES_ENC/u0/u3/U143  ( .A1(\AES_ENC/u0/u3/n1125 ), .A2(\AES_ENC/u0/u3/n1124 ), .A3(\AES_ENC/u0/u3/n1123 ), .A4(\AES_ENC/u0/u3/n1122 ), .ZN(\AES_ENC/u0/u3/n1126 ) );
NOR4_X2 \AES_ENC/u0/u3/U142  ( .A1(\AES_ENC/u0/u3/n1084 ), .A2(\AES_ENC/u0/u3/n1083 ), .A3(\AES_ENC/u0/u3/n1082 ), .A4(\AES_ENC/u0/u3/n1081 ), .ZN(\AES_ENC/u0/u3/n1085 ) );
NOR2_X2 \AES_ENC/u0/u3/U141  ( .A1(\AES_ENC/u0/u3/n1076 ), .A2(\AES_ENC/u0/u3/n1075 ), .ZN(\AES_ENC/u0/u3/n1086 ) );
NOR3_X2 \AES_ENC/u0/u3/U140  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n1054 ), .A3(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n961 ) );
NOR3_X2 \AES_ENC/u0/u3/U132  ( .A1(\AES_ENC/u0/u3/n620 ), .A2(\AES_ENC/u0/u3/n1074 ), .A3(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n671 ) );
NOR2_X2 \AES_ENC/u0/u3/U131  ( .A1(\AES_ENC/u0/u3/n1057 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n1062 ) );
NOR2_X2 \AES_ENC/u0/u3/U130  ( .A1(\AES_ENC/u0/u3/n1060 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n1061 ) );
NOR2_X2 \AES_ENC/u0/u3/U129  ( .A1(\AES_ENC/u0/u3/n1055 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n1063 ) );
NOR4_X2 \AES_ENC/u0/u3/U128  ( .A1(\AES_ENC/u0/u3/n1064 ), .A2(\AES_ENC/u0/u3/n1063 ), .A3(\AES_ENC/u0/u3/n1062 ), .A4(\AES_ENC/u0/u3/n1061 ), .ZN(\AES_ENC/u0/u3/n1065 ) );
NOR3_X2 \AES_ENC/u0/u3/U127  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n1120 ), .A3(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n918 ) );
NOR2_X2 \AES_ENC/u0/u3/U126  ( .A1(\AES_ENC/u0/u3/n914 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n915 ) );
NOR3_X2 \AES_ENC/u0/u3/U121  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n573 ), .A3(\AES_ENC/u0/u3/n1013 ), .ZN(\AES_ENC/u0/u3/n917 ) );
NOR4_X2 \AES_ENC/u0/u3/U120  ( .A1(\AES_ENC/u0/u3/n918 ), .A2(\AES_ENC/u0/u3/n917 ), .A3(\AES_ENC/u0/u3/n916 ), .A4(\AES_ENC/u0/u3/n915 ), .ZN(\AES_ENC/u0/u3/n919 ) );
NOR2_X2 \AES_ENC/u0/u3/U119  ( .A1(\AES_ENC/u0/u3/n735 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n687 ) );
NOR2_X2 \AES_ENC/u0/u3/U118  ( .A1(\AES_ENC/u0/u3/n684 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n688 ) );
NOR2_X2 \AES_ENC/u0/u3/U117  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n600 ), .ZN(\AES_ENC/u0/u3/n686 ) );
NOR4_X2 \AES_ENC/u0/u3/U116  ( .A1(\AES_ENC/u0/u3/n688 ), .A2(\AES_ENC/u0/u3/n687 ), .A3(\AES_ENC/u0/u3/n686 ), .A4(\AES_ENC/u0/u3/n685 ), .ZN(\AES_ENC/u0/u3/n689 ) );
NOR2_X2 \AES_ENC/u0/u3/U115  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n582 ), .ZN(\AES_ENC/u0/u3/n770 ) );
NOR2_X2 \AES_ENC/u0/u3/U106  ( .A1(\AES_ENC/u0/u3/n1103 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n772 ) );
NOR2_X2 \AES_ENC/u0/u3/U105  ( .A1(\AES_ENC/u0/u3/n610 ), .A2(\AES_ENC/u0/u3/n599 ), .ZN(\AES_ENC/u0/u3/n773 ) );
NOR4_X2 \AES_ENC/u0/u3/U104  ( .A1(\AES_ENC/u0/u3/n773 ), .A2(\AES_ENC/u0/u3/n772 ), .A3(\AES_ENC/u0/u3/n771 ), .A4(\AES_ENC/u0/u3/n770 ), .ZN(\AES_ENC/u0/u3/n774 ) );
NOR2_X2 \AES_ENC/u0/u3/U103  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n595 ), .ZN(\AES_ENC/u0/u3/n858 ) );
NOR2_X2 \AES_ENC/u0/u3/U102  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n855 ), .ZN(\AES_ENC/u0/u3/n857 ) );
NOR2_X2 \AES_ENC/u0/u3/U101  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n587 ), .ZN(\AES_ENC/u0/u3/n856 ) );
NOR4_X2 \AES_ENC/u0/u3/U100  ( .A1(\AES_ENC/u0/u3/n858 ), .A2(\AES_ENC/u0/u3/n857 ), .A3(\AES_ENC/u0/u3/n856 ), .A4(\AES_ENC/u0/u3/n958 ), .ZN(\AES_ENC/u0/u3/n859 ) );
NOR2_X2 \AES_ENC/u0/u3/U95  ( .A1(\AES_ENC/u0/u3/n583 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n814 ) );
NOR3_X2 \AES_ENC/u0/u3/U94  ( .A1(\AES_ENC/u0/u3/n606 ), .A2(\AES_ENC/u0/u3/n1058 ), .A3(\AES_ENC/u0/u3/n1059 ), .ZN(\AES_ENC/u0/u3/n815 ) );
NOR2_X2 \AES_ENC/u0/u3/U93  ( .A1(\AES_ENC/u0/u3/n907 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n813 ) );
NOR4_X2 \AES_ENC/u0/u3/U92  ( .A1(\AES_ENC/u0/u3/n815 ), .A2(\AES_ENC/u0/u3/n814 ), .A3(\AES_ENC/u0/u3/n813 ), .A4(\AES_ENC/u0/u3/n812 ), .ZN(\AES_ENC/u0/u3/n816 ) );
NOR2_X2 \AES_ENC/u0/u3/U91  ( .A1(\AES_ENC/u0/u3/n617 ), .A2(\AES_ENC/u0/u3/n569 ), .ZN(\AES_ENC/u0/u3/n721 ) );
NOR2_X2 \AES_ENC/u0/u3/U90  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n1096 ), .ZN(\AES_ENC/u0/u3/n722 ) );
NOR2_X2 \AES_ENC/u0/u3/U89  ( .A1(\AES_ENC/u0/u3/n1031 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n723 ) );
NOR4_X2 \AES_ENC/u0/u3/U88  ( .A1(\AES_ENC/u0/u3/n724 ), .A2(\AES_ENC/u0/u3/n723 ), .A3(\AES_ENC/u0/u3/n722 ), .A4(\AES_ENC/u0/u3/n721 ), .ZN(\AES_ENC/u0/u3/n725 ) );
NOR2_X2 \AES_ENC/u0/u3/U87  ( .A1(\AES_ENC/u0/u3/n911 ), .A2(\AES_ENC/u0/u3/n990 ), .ZN(\AES_ENC/u0/u3/n1009 ) );
NOR2_X2 \AES_ENC/u0/u3/U86  ( .A1(\AES_ENC/u0/u3/n1013 ), .A2(\AES_ENC/u0/u3/n573 ), .ZN(\AES_ENC/u0/u3/n1014 ) );
NOR2_X2 \AES_ENC/u0/u3/U81  ( .A1(\AES_ENC/u0/u3/n1014 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n1015 ) );
NOR4_X2 \AES_ENC/u0/u3/U80  ( .A1(\AES_ENC/u0/u3/n1016 ), .A2(\AES_ENC/u0/u3/n1015 ), .A3(\AES_ENC/u0/u3/n1119 ), .A4(\AES_ENC/u0/u3/n1046 ), .ZN(\AES_ENC/u0/u3/n1017 ) );
NOR2_X2 \AES_ENC/u0/u3/U79  ( .A1(\AES_ENC/u0/u3/n606 ), .A2(\AES_ENC/u0/u3/n589 ), .ZN(\AES_ENC/u0/u3/n997 ) );
NOR2_X2 \AES_ENC/u0/u3/U78  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n577 ), .ZN(\AES_ENC/u0/u3/n1000 ) );
NOR2_X2 \AES_ENC/u0/u3/U74  ( .A1(\AES_ENC/u0/u3/n616 ), .A2(\AES_ENC/u0/u3/n1096 ), .ZN(\AES_ENC/u0/u3/n999 ) );
NOR4_X2 \AES_ENC/u0/u3/U73  ( .A1(\AES_ENC/u0/u3/n1000 ), .A2(\AES_ENC/u0/u3/n999 ), .A3(\AES_ENC/u0/u3/n998 ), .A4(\AES_ENC/u0/u3/n997 ), .ZN(\AES_ENC/u0/u3/n1001 ) );
NOR2_X2 \AES_ENC/u0/u3/U72  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n1096 ), .ZN(\AES_ENC/u0/u3/n697 ) );
NOR2_X2 \AES_ENC/u0/u3/U71  ( .A1(\AES_ENC/u0/u3/n620 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n958 ) );
NOR2_X2 \AES_ENC/u0/u3/U65  ( .A1(\AES_ENC/u0/u3/n911 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n983 ) );
NOR2_X2 \AES_ENC/u0/u3/U64  ( .A1(\AES_ENC/u0/u3/n1054 ), .A2(\AES_ENC/u0/u3/n1103 ), .ZN(\AES_ENC/u0/u3/n1031 ) );
INV_X4 \AES_ENC/u0/u3/U63  ( .A(\AES_ENC/u0/u3/n1050 ), .ZN(\AES_ENC/u0/u3/n612 ) );
INV_X4 \AES_ENC/u0/u3/U62  ( .A(\AES_ENC/u0/u3/n1072 ), .ZN(\AES_ENC/u0/u3/n605 ) );
INV_X4 \AES_ENC/u0/u3/U61  ( .A(\AES_ENC/u0/u3/n1073 ), .ZN(\AES_ENC/u0/u3/n604 ) );
NOR2_X2 \AES_ENC/u0/u3/U59  ( .A1(\AES_ENC/u0/u3/n582 ), .A2(\AES_ENC/u0/u3/n613 ), .ZN(\AES_ENC/u0/u3/n880 ) );
NOR3_X2 \AES_ENC/u0/u3/U58  ( .A1(\AES_ENC/u0/u3/n826 ), .A2(\AES_ENC/u0/u3/n1121 ), .A3(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n946 ) );
INV_X4 \AES_ENC/u0/u3/U57  ( .A(\AES_ENC/u0/u3/n1010 ), .ZN(\AES_ENC/u0/u3/n608 ) );
NOR3_X2 \AES_ENC/u0/u3/U50  ( .A1(\AES_ENC/u0/u3/n573 ), .A2(\AES_ENC/u0/u3/n1029 ), .A3(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n1119 ) );
INV_X4 \AES_ENC/u0/u3/U49  ( .A(\AES_ENC/u0/u3/n956 ), .ZN(\AES_ENC/u0/u3/n615 ) );
NOR2_X2 \AES_ENC/u0/u3/U48  ( .A1(\AES_ENC/u0/u3/n623 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n1013 ) );
NOR2_X2 \AES_ENC/u0/u3/U47  ( .A1(\AES_ENC/u0/u3/n620 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n910 ) );
NOR2_X2 \AES_ENC/u0/u3/U46  ( .A1(\AES_ENC/u0/u3/n569 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n1091 ) );
NOR2_X2 \AES_ENC/u0/u3/U45  ( .A1(\AES_ENC/u0/u3/n622 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n990 ) );
NOR2_X2 \AES_ENC/u0/u3/U44  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/u0/u3/n1121 ), .ZN(\AES_ENC/u0/u3/n996 ) );
NOR2_X2 \AES_ENC/u0/u3/U43  ( .A1(\AES_ENC/u0/u3/n610 ), .A2(\AES_ENC/u0/u3/n600 ), .ZN(\AES_ENC/u0/u3/n628 ) );
NOR2_X2 \AES_ENC/u0/u3/U42  ( .A1(\AES_ENC/u0/u3/n576 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n866 ) );
NOR2_X2 \AES_ENC/u0/u3/U41  ( .A1(\AES_ENC/u0/u3/n603 ), .A2(\AES_ENC/u0/u3/n610 ), .ZN(\AES_ENC/u0/u3/n1006 ) );
NOR2_X2 \AES_ENC/u0/u3/U36  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n1117 ), .ZN(\AES_ENC/u0/u3/n1118 ) );
NOR2_X2 \AES_ENC/u0/u3/U35  ( .A1(\AES_ENC/u0/u3/n1119 ), .A2(\AES_ENC/u0/u3/n1118 ), .ZN(\AES_ENC/u0/u3/n1127 ) );
NOR2_X2 \AES_ENC/u0/u3/U34  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n594 ), .ZN(\AES_ENC/u0/u3/n629 ) );
NOR2_X2 \AES_ENC/u0/u3/U33  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n906 ), .ZN(\AES_ENC/u0/u3/n909 ) );
NOR2_X2 \AES_ENC/u0/u3/U32  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n597 ), .ZN(\AES_ENC/u0/u3/n658 ) );
NOR2_X2 \AES_ENC/u0/u3/U31  ( .A1(\AES_ENC/u0/u3/n1116 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n695 ) );
NOR2_X2 \AES_ENC/u0/u3/U30  ( .A1(\AES_ENC/u0/u3/n1078 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n1083 ) );
NOR2_X2 \AES_ENC/u0/u3/U29  ( .A1(\AES_ENC/u0/u3/n941 ), .A2(\AES_ENC/u0/u3/n608 ), .ZN(\AES_ENC/u0/u3/n724 ) );
NOR2_X2 \AES_ENC/u0/u3/U24  ( .A1(\AES_ENC/u0/u3/n576 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n840 ) );
NOR2_X2 \AES_ENC/u0/u3/U23  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n593 ), .ZN(\AES_ENC/u0/u3/n633 ) );
NOR2_X2 \AES_ENC/u0/u3/U21  ( .A1(\AES_ENC/u0/u3/n1009 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n960 ) );
NOR2_X2 \AES_ENC/u0/u3/U20  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n1045 ), .ZN(\AES_ENC/u0/u3/n812 ) );
NOR2_X2 \AES_ENC/u0/u3/U19  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n1080 ), .ZN(\AES_ENC/u0/u3/n1081 ) );
NOR2_X2 \AES_ENC/u0/u3/U18  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n601 ), .ZN(\AES_ENC/u0/u3/n982 ) );
NOR2_X2 \AES_ENC/u0/u3/U17  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n594 ), .ZN(\AES_ENC/u0/u3/n757 ) );
NOR2_X2 \AES_ENC/u0/u3/U16  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n590 ), .ZN(\AES_ENC/u0/u3/n698 ) );
NOR2_X2 \AES_ENC/u0/u3/U15  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n619 ), .ZN(\AES_ENC/u0/u3/n708 ) );
NOR2_X2 \AES_ENC/u0/u3/U10  ( .A1(\AES_ENC/u0/u3/n619 ), .A2(\AES_ENC/u0/u3/n604 ), .ZN(\AES_ENC/u0/u3/n803 ) );
NOR2_X2 \AES_ENC/u0/u3/U9  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n881 ), .ZN(\AES_ENC/u0/u3/n711 ) );
NOR2_X2 \AES_ENC/u0/u3/U8  ( .A1(\AES_ENC/u0/u3/n615 ), .A2(\AES_ENC/u0/u3/n582 ), .ZN(\AES_ENC/u0/u3/n867 ) );
NOR2_X2 \AES_ENC/u0/u3/U7  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n599 ), .ZN(\AES_ENC/u0/u3/n804 ) );
NOR2_X2 \AES_ENC/u0/u3/U6  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n620 ), .ZN(\AES_ENC/u0/u3/n1046 ) );
OR2_X4 \AES_ENC/u0/u3/U5  ( .A1(\AES_ENC/u0/u3/n624 ), .A2(\AES_ENC/w3[25] ),.ZN(\AES_ENC/u0/u3/n570 ) );
OR2_X4 \AES_ENC/u0/u3/U4  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/w3[28] ),.ZN(\AES_ENC/u0/u3/n569 ) );
NAND2_X2 \AES_ENC/u0/u3/U514  ( .A1(\AES_ENC/u0/u3/n1121 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n1030 ) );
AND2_X2 \AES_ENC/u0/u3/U513  ( .A1(\AES_ENC/u0/u3/n597 ), .A2(\AES_ENC/u0/u3/n1030 ), .ZN(\AES_ENC/u0/u3/n1049 ) );
NAND2_X2 \AES_ENC/u0/u3/U511  ( .A1(\AES_ENC/u0/u3/n1049 ), .A2(\AES_ENC/u0/u3/n794 ), .ZN(\AES_ENC/u0/u3/n637 ) );
AND2_X2 \AES_ENC/u0/u3/U493  ( .A1(\AES_ENC/u0/u3/n779 ), .A2(\AES_ENC/u0/u3/n996 ), .ZN(\AES_ENC/u0/u3/n632 ) );
NAND4_X2 \AES_ENC/u0/u3/U485  ( .A1(\AES_ENC/u0/u3/n637 ), .A2(\AES_ENC/u0/u3/n636 ), .A3(\AES_ENC/u0/u3/n635 ), .A4(\AES_ENC/u0/u3/n634 ), .ZN(\AES_ENC/u0/u3/n638 ) );
NAND2_X2 \AES_ENC/u0/u3/U484  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n638 ), .ZN(\AES_ENC/u0/u3/n679 ) );
NAND2_X2 \AES_ENC/u0/u3/U481  ( .A1(\AES_ENC/u0/u3/n1094 ), .A2(\AES_ENC/u0/u3/n591 ), .ZN(\AES_ENC/u0/u3/n648 ) );
NAND2_X2 \AES_ENC/u0/u3/U476  ( .A1(\AES_ENC/u0/u3/n601 ), .A2(\AES_ENC/u0/u3/n590 ), .ZN(\AES_ENC/u0/u3/n762 ) );
NAND2_X2 \AES_ENC/u0/u3/U475  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n762 ), .ZN(\AES_ENC/u0/u3/n647 ) );
NAND4_X2 \AES_ENC/u0/u3/U457  ( .A1(\AES_ENC/u0/u3/n648 ), .A2(\AES_ENC/u0/u3/n647 ), .A3(\AES_ENC/u0/u3/n646 ), .A4(\AES_ENC/u0/u3/n645 ), .ZN(\AES_ENC/u0/u3/n649 ) );
NAND2_X2 \AES_ENC/u0/u3/U456  ( .A1(\AES_ENC/w3[24] ), .A2(\AES_ENC/u0/u3/n649 ), .ZN(\AES_ENC/u0/u3/n665 ) );
NAND2_X2 \AES_ENC/u0/u3/U454  ( .A1(\AES_ENC/u0/u3/n596 ), .A2(\AES_ENC/u0/u3/n623 ), .ZN(\AES_ENC/u0/u3/n855 ) );
NAND2_X2 \AES_ENC/u0/u3/U453  ( .A1(\AES_ENC/u0/u3/n587 ), .A2(\AES_ENC/u0/u3/n855 ), .ZN(\AES_ENC/u0/u3/n821 ) );
NAND2_X2 \AES_ENC/u0/u3/U452  ( .A1(\AES_ENC/u0/u3/n1093 ), .A2(\AES_ENC/u0/u3/n821 ), .ZN(\AES_ENC/u0/u3/n662 ) );
NAND2_X2 \AES_ENC/u0/u3/U451  ( .A1(\AES_ENC/u0/u3/n619 ), .A2(\AES_ENC/u0/u3/n589 ), .ZN(\AES_ENC/u0/u3/n650 ) );
NAND2_X2 \AES_ENC/u0/u3/U450  ( .A1(\AES_ENC/u0/u3/n956 ), .A2(\AES_ENC/u0/u3/n650 ), .ZN(\AES_ENC/u0/u3/n661 ) );
NAND2_X2 \AES_ENC/u0/u3/U449  ( .A1(\AES_ENC/u0/u3/n626 ), .A2(\AES_ENC/u0/u3/n627 ), .ZN(\AES_ENC/u0/u3/n839 ) );
OR2_X2 \AES_ENC/u0/u3/U446  ( .A1(\AES_ENC/u0/u3/n839 ), .A2(\AES_ENC/u0/u3/n932 ), .ZN(\AES_ENC/u0/u3/n656 ) );
NAND2_X2 \AES_ENC/u0/u3/U445  ( .A1(\AES_ENC/u0/u3/n621 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n1096 ) );
NAND2_X2 \AES_ENC/u0/u3/U444  ( .A1(\AES_ENC/u0/u3/n1030 ), .A2(\AES_ENC/u0/u3/n1096 ), .ZN(\AES_ENC/u0/u3/n651 ) );
NAND2_X2 \AES_ENC/u0/u3/U443  ( .A1(\AES_ENC/u0/u3/n1114 ), .A2(\AES_ENC/u0/u3/n651 ), .ZN(\AES_ENC/u0/u3/n655 ) );
OR3_X2 \AES_ENC/u0/u3/U440  ( .A1(\AES_ENC/u0/u3/n1079 ), .A2(\AES_ENC/w3[31] ), .A3(\AES_ENC/u0/u3/n626 ), .ZN(\AES_ENC/u0/u3/n654 ) );
NAND2_X2 \AES_ENC/u0/u3/U439  ( .A1(\AES_ENC/u0/u3/n593 ), .A2(\AES_ENC/u0/u3/n601 ), .ZN(\AES_ENC/u0/u3/n652 ) );
NAND4_X2 \AES_ENC/u0/u3/U437  ( .A1(\AES_ENC/u0/u3/n656 ), .A2(\AES_ENC/u0/u3/n655 ), .A3(\AES_ENC/u0/u3/n654 ), .A4(\AES_ENC/u0/u3/n653 ), .ZN(\AES_ENC/u0/u3/n657 ) );
NAND2_X2 \AES_ENC/u0/u3/U436  ( .A1(\AES_ENC/w3[26] ), .A2(\AES_ENC/u0/u3/n657 ), .ZN(\AES_ENC/u0/u3/n660 ) );
NAND4_X2 \AES_ENC/u0/u3/U432  ( .A1(\AES_ENC/u0/u3/n662 ), .A2(\AES_ENC/u0/u3/n661 ), .A3(\AES_ENC/u0/u3/n660 ), .A4(\AES_ENC/u0/u3/n659 ), .ZN(\AES_ENC/u0/u3/n663 ) );
NAND2_X2 \AES_ENC/u0/u3/U431  ( .A1(\AES_ENC/u0/u3/n663 ), .A2(\AES_ENC/u0/u3/n574 ), .ZN(\AES_ENC/u0/u3/n664 ) );
NAND2_X2 \AES_ENC/u0/u3/U430  ( .A1(\AES_ENC/u0/u3/n665 ), .A2(\AES_ENC/u0/u3/n664 ), .ZN(\AES_ENC/u0/u3/n666 ) );
NAND2_X2 \AES_ENC/u0/u3/U429  ( .A1(\AES_ENC/w3[30] ), .A2(\AES_ENC/u0/u3/n666 ), .ZN(\AES_ENC/u0/u3/n678 ) );
NAND2_X2 \AES_ENC/u0/u3/U426  ( .A1(\AES_ENC/u0/u3/n735 ), .A2(\AES_ENC/u0/u3/n1093 ), .ZN(\AES_ENC/u0/u3/n675 ) );
NAND2_X2 \AES_ENC/u0/u3/U425  ( .A1(\AES_ENC/u0/u3/n588 ), .A2(\AES_ENC/u0/u3/n597 ), .ZN(\AES_ENC/u0/u3/n1045 ) );
OR2_X2 \AES_ENC/u0/u3/U424  ( .A1(\AES_ENC/u0/u3/n1045 ), .A2(\AES_ENC/u0/u3/n605 ), .ZN(\AES_ENC/u0/u3/n674 ) );
NAND2_X2 \AES_ENC/u0/u3/U423  ( .A1(\AES_ENC/w3[25] ), .A2(\AES_ENC/u0/u3/n620 ), .ZN(\AES_ENC/u0/u3/n667 ) );
NAND2_X2 \AES_ENC/u0/u3/U422  ( .A1(\AES_ENC/u0/u3/n619 ), .A2(\AES_ENC/u0/u3/n667 ), .ZN(\AES_ENC/u0/u3/n1071 ) );
NAND4_X2 \AES_ENC/u0/u3/U412  ( .A1(\AES_ENC/u0/u3/n675 ), .A2(\AES_ENC/u0/u3/n674 ), .A3(\AES_ENC/u0/u3/n673 ), .A4(\AES_ENC/u0/u3/n672 ), .ZN(\AES_ENC/u0/u3/n676 ) );
NAND2_X2 \AES_ENC/u0/u3/U411  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n676 ), .ZN(\AES_ENC/u0/u3/n677 ) );
NAND2_X2 \AES_ENC/u0/u3/U408  ( .A1(\AES_ENC/u0/u3/n800 ), .A2(\AES_ENC/u0/u3/n1022 ), .ZN(\AES_ENC/u0/u3/n680 ) );
NAND2_X2 \AES_ENC/u0/u3/U407  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n680 ), .ZN(\AES_ENC/u0/u3/n681 ) );
AND2_X2 \AES_ENC/u0/u3/U402  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n684 ), .ZN(\AES_ENC/u0/u3/n682 ) );
NAND4_X2 \AES_ENC/u0/u3/U395  ( .A1(\AES_ENC/u0/u3/n691 ), .A2(\AES_ENC/u0/u3/n581 ), .A3(\AES_ENC/u0/u3/n690 ), .A4(\AES_ENC/u0/u3/n689 ), .ZN(\AES_ENC/u0/u3/n692 ) );
NAND2_X2 \AES_ENC/u0/u3/U394  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n692 ), .ZN(\AES_ENC/u0/u3/n733 ) );
NAND2_X2 \AES_ENC/u0/u3/U392  ( .A1(\AES_ENC/u0/u3/n977 ), .A2(\AES_ENC/u0/u3/n1050 ), .ZN(\AES_ENC/u0/u3/n702 ) );
NAND2_X2 \AES_ENC/u0/u3/U391  ( .A1(\AES_ENC/u0/u3/n1093 ), .A2(\AES_ENC/u0/u3/n1045 ), .ZN(\AES_ENC/u0/u3/n701 ) );
NAND4_X2 \AES_ENC/u0/u3/U381  ( .A1(\AES_ENC/u0/u3/n702 ), .A2(\AES_ENC/u0/u3/n701 ), .A3(\AES_ENC/u0/u3/n700 ), .A4(\AES_ENC/u0/u3/n699 ), .ZN(\AES_ENC/u0/u3/n703 ) );
NAND2_X2 \AES_ENC/u0/u3/U380  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n703 ), .ZN(\AES_ENC/u0/u3/n732 ) );
AND2_X2 \AES_ENC/u0/u3/U379  ( .A1(\AES_ENC/w3[24] ), .A2(\AES_ENC/w3[30] ),.ZN(\AES_ENC/u0/u3/n1113 ) );
NAND2_X2 \AES_ENC/u0/u3/U378  ( .A1(\AES_ENC/u0/u3/n601 ), .A2(\AES_ENC/u0/u3/n1030 ), .ZN(\AES_ENC/u0/u3/n881 ) );
NAND2_X2 \AES_ENC/u0/u3/U377  ( .A1(\AES_ENC/u0/u3/n1093 ), .A2(\AES_ENC/u0/u3/n881 ), .ZN(\AES_ENC/u0/u3/n715 ) );
NAND2_X2 \AES_ENC/u0/u3/U376  ( .A1(\AES_ENC/u0/u3/n1010 ), .A2(\AES_ENC/u0/u3/n600 ), .ZN(\AES_ENC/u0/u3/n714 ) );
NAND2_X2 \AES_ENC/u0/u3/U375  ( .A1(\AES_ENC/u0/u3/n855 ), .A2(\AES_ENC/u0/u3/n588 ), .ZN(\AES_ENC/u0/u3/n1117 ) );
XNOR2_X2 \AES_ENC/u0/u3/U371  ( .A(\AES_ENC/u0/u3/n611 ), .B(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n824 ) );
NAND4_X2 \AES_ENC/u0/u3/U362  ( .A1(\AES_ENC/u0/u3/n715 ), .A2(\AES_ENC/u0/u3/n714 ), .A3(\AES_ENC/u0/u3/n713 ), .A4(\AES_ENC/u0/u3/n712 ), .ZN(\AES_ENC/u0/u3/n716 ) );
NAND2_X2 \AES_ENC/u0/u3/U361  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n716 ), .ZN(\AES_ENC/u0/u3/n731 ) );
AND2_X2 \AES_ENC/u0/u3/U360  ( .A1(\AES_ENC/w3[30] ), .A2(\AES_ENC/u0/u3/n574 ), .ZN(\AES_ENC/u0/u3/n1131 ) );
NAND2_X2 \AES_ENC/u0/u3/U359  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n717 ) );
NAND2_X2 \AES_ENC/u0/u3/U358  ( .A1(\AES_ENC/u0/u3/n1029 ), .A2(\AES_ENC/u0/u3/n717 ), .ZN(\AES_ENC/u0/u3/n728 ) );
NAND2_X2 \AES_ENC/u0/u3/U357  ( .A1(\AES_ENC/w3[25] ), .A2(\AES_ENC/u0/u3/n624 ), .ZN(\AES_ENC/u0/u3/n1097 ) );
NAND2_X2 \AES_ENC/u0/u3/U356  ( .A1(\AES_ENC/u0/u3/n603 ), .A2(\AES_ENC/u0/u3/n1097 ), .ZN(\AES_ENC/u0/u3/n718 ) );
NAND2_X2 \AES_ENC/u0/u3/U355  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n718 ), .ZN(\AES_ENC/u0/u3/n727 ) );
NAND4_X2 \AES_ENC/u0/u3/U344  ( .A1(\AES_ENC/u0/u3/n728 ), .A2(\AES_ENC/u0/u3/n727 ), .A3(\AES_ENC/u0/u3/n726 ), .A4(\AES_ENC/u0/u3/n725 ), .ZN(\AES_ENC/u0/u3/n729 ) );
NAND2_X2 \AES_ENC/u0/u3/U343  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n729 ), .ZN(\AES_ENC/u0/u3/n730 ) );
NAND4_X2 \AES_ENC/u0/u3/U342  ( .A1(\AES_ENC/u0/u3/n733 ), .A2(\AES_ENC/u0/u3/n732 ), .A3(\AES_ENC/u0/u3/n731 ), .A4(\AES_ENC/u0/u3/n730 ), .ZN(\AES_ENC/u0/subword[1] ) );
NAND2_X2 \AES_ENC/u0/u3/U341  ( .A1(\AES_ENC/w3[31] ), .A2(\AES_ENC/u0/u3/n611 ), .ZN(\AES_ENC/u0/u3/n734 ) );
NAND2_X2 \AES_ENC/u0/u3/U340  ( .A1(\AES_ENC/u0/u3/n734 ), .A2(\AES_ENC/u0/u3/n607 ), .ZN(\AES_ENC/u0/u3/n738 ) );
OR4_X2 \AES_ENC/u0/u3/U339  ( .A1(\AES_ENC/u0/u3/n738 ), .A2(\AES_ENC/u0/u3/n626 ), .A3(\AES_ENC/u0/u3/n826 ), .A4(\AES_ENC/u0/u3/n1121 ), .ZN(\AES_ENC/u0/u3/n746 ) );
NAND2_X2 \AES_ENC/u0/u3/U337  ( .A1(\AES_ENC/u0/u3/n1100 ), .A2(\AES_ENC/u0/u3/n587 ), .ZN(\AES_ENC/u0/u3/n992 ) );
OR2_X2 \AES_ENC/u0/u3/U336  ( .A1(\AES_ENC/u0/u3/n610 ), .A2(\AES_ENC/u0/u3/n735 ), .ZN(\AES_ENC/u0/u3/n737 ) );
NAND2_X2 \AES_ENC/u0/u3/U334  ( .A1(\AES_ENC/u0/u3/n619 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n753 ) );
NAND2_X2 \AES_ENC/u0/u3/U333  ( .A1(\AES_ENC/u0/u3/n582 ), .A2(\AES_ENC/u0/u3/n753 ), .ZN(\AES_ENC/u0/u3/n1080 ) );
NAND2_X2 \AES_ENC/u0/u3/U332  ( .A1(\AES_ENC/u0/u3/n1048 ), .A2(\AES_ENC/u0/u3/n576 ), .ZN(\AES_ENC/u0/u3/n736 ) );
NAND2_X2 \AES_ENC/u0/u3/U331  ( .A1(\AES_ENC/u0/u3/n737 ), .A2(\AES_ENC/u0/u3/n736 ), .ZN(\AES_ENC/u0/u3/n739 ) );
NAND2_X2 \AES_ENC/u0/u3/U330  ( .A1(\AES_ENC/u0/u3/n739 ), .A2(\AES_ENC/u0/u3/n738 ), .ZN(\AES_ENC/u0/u3/n745 ) );
NAND2_X2 \AES_ENC/u0/u3/U326  ( .A1(\AES_ENC/u0/u3/n1096 ), .A2(\AES_ENC/u0/u3/n590 ), .ZN(\AES_ENC/u0/u3/n906 ) );
NAND4_X2 \AES_ENC/u0/u3/U323  ( .A1(\AES_ENC/u0/u3/n746 ), .A2(\AES_ENC/u0/u3/n992 ), .A3(\AES_ENC/u0/u3/n745 ), .A4(\AES_ENC/u0/u3/n744 ), .ZN(\AES_ENC/u0/u3/n747 ) );
NAND2_X2 \AES_ENC/u0/u3/U322  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n747 ), .ZN(\AES_ENC/u0/u3/n793 ) );
NAND2_X2 \AES_ENC/u0/u3/U321  ( .A1(\AES_ENC/u0/u3/n584 ), .A2(\AES_ENC/u0/u3/n855 ), .ZN(\AES_ENC/u0/u3/n748 ) );
NAND2_X2 \AES_ENC/u0/u3/U320  ( .A1(\AES_ENC/u0/u3/n956 ), .A2(\AES_ENC/u0/u3/n748 ), .ZN(\AES_ENC/u0/u3/n760 ) );
NAND2_X2 \AES_ENC/u0/u3/U313  ( .A1(\AES_ENC/u0/u3/n590 ), .A2(\AES_ENC/u0/u3/n753 ), .ZN(\AES_ENC/u0/u3/n1023 ) );
NAND4_X2 \AES_ENC/u0/u3/U308  ( .A1(\AES_ENC/u0/u3/n760 ), .A2(\AES_ENC/u0/u3/n992 ), .A3(\AES_ENC/u0/u3/n759 ), .A4(\AES_ENC/u0/u3/n758 ), .ZN(\AES_ENC/u0/u3/n761 ) );
NAND2_X2 \AES_ENC/u0/u3/U307  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n761 ), .ZN(\AES_ENC/u0/u3/n792 ) );
NAND2_X2 \AES_ENC/u0/u3/U306  ( .A1(\AES_ENC/u0/u3/n584 ), .A2(\AES_ENC/u0/u3/n603 ), .ZN(\AES_ENC/u0/u3/n989 ) );
NAND2_X2 \AES_ENC/u0/u3/U305  ( .A1(\AES_ENC/u0/u3/n1050 ), .A2(\AES_ENC/u0/u3/n989 ), .ZN(\AES_ENC/u0/u3/n777 ) );
NAND2_X2 \AES_ENC/u0/u3/U304  ( .A1(\AES_ENC/u0/u3/n1093 ), .A2(\AES_ENC/u0/u3/n762 ), .ZN(\AES_ENC/u0/u3/n776 ) );
XNOR2_X2 \AES_ENC/u0/u3/U301  ( .A(\AES_ENC/w3[31] ), .B(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n959 ) );
NAND4_X2 \AES_ENC/u0/u3/U289  ( .A1(\AES_ENC/u0/u3/n777 ), .A2(\AES_ENC/u0/u3/n776 ), .A3(\AES_ENC/u0/u3/n775 ), .A4(\AES_ENC/u0/u3/n774 ), .ZN(\AES_ENC/u0/u3/n778 ) );
NAND2_X2 \AES_ENC/u0/u3/U288  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n778 ), .ZN(\AES_ENC/u0/u3/n791 ) );
NAND2_X2 \AES_ENC/u0/u3/U287  ( .A1(\AES_ENC/u0/u3/n1056 ), .A2(\AES_ENC/u0/u3/n1050 ), .ZN(\AES_ENC/u0/u3/n788 ) );
NAND2_X2 \AES_ENC/u0/u3/U286  ( .A1(\AES_ENC/u0/u3/n1091 ), .A2(\AES_ENC/u0/u3/n779 ), .ZN(\AES_ENC/u0/u3/n787 ) );
NAND2_X2 \AES_ENC/u0/u3/U285  ( .A1(\AES_ENC/u0/u3/n956 ), .A2(\AES_ENC/w3[25] ), .ZN(\AES_ENC/u0/u3/n786 ) );
NAND4_X2 \AES_ENC/u0/u3/U278  ( .A1(\AES_ENC/u0/u3/n788 ), .A2(\AES_ENC/u0/u3/n787 ), .A3(\AES_ENC/u0/u3/n786 ), .A4(\AES_ENC/u0/u3/n785 ), .ZN(\AES_ENC/u0/u3/n789 ) );
NAND2_X2 \AES_ENC/u0/u3/U277  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n789 ), .ZN(\AES_ENC/u0/u3/n790 ) );
NAND4_X2 \AES_ENC/u0/u3/U276  ( .A1(\AES_ENC/u0/u3/n793 ), .A2(\AES_ENC/u0/u3/n792 ), .A3(\AES_ENC/u0/u3/n791 ), .A4(\AES_ENC/u0/u3/n790 ), .ZN(\AES_ENC/u0/subword[2] ) );
NAND2_X2 \AES_ENC/u0/u3/U275  ( .A1(\AES_ENC/u0/u3/n1059 ), .A2(\AES_ENC/u0/u3/n794 ), .ZN(\AES_ENC/u0/u3/n810 ) );
NAND2_X2 \AES_ENC/u0/u3/U274  ( .A1(\AES_ENC/u0/u3/n1049 ), .A2(\AES_ENC/u0/u3/n956 ), .ZN(\AES_ENC/u0/u3/n809 ) );
OR2_X2 \AES_ENC/u0/u3/U266  ( .A1(\AES_ENC/u0/u3/n1096 ), .A2(\AES_ENC/u0/u3/n606 ), .ZN(\AES_ENC/u0/u3/n802 ) );
NAND2_X2 \AES_ENC/u0/u3/U265  ( .A1(\AES_ENC/u0/u3/n1053 ), .A2(\AES_ENC/u0/u3/n800 ), .ZN(\AES_ENC/u0/u3/n801 ) );
NAND2_X2 \AES_ENC/u0/u3/U264  ( .A1(\AES_ENC/u0/u3/n802 ), .A2(\AES_ENC/u0/u3/n801 ), .ZN(\AES_ENC/u0/u3/n805 ) );
NAND4_X2 \AES_ENC/u0/u3/U261  ( .A1(\AES_ENC/u0/u3/n810 ), .A2(\AES_ENC/u0/u3/n809 ), .A3(\AES_ENC/u0/u3/n808 ), .A4(\AES_ENC/u0/u3/n807 ), .ZN(\AES_ENC/u0/u3/n811 ) );
NAND2_X2 \AES_ENC/u0/u3/U260  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n811 ), .ZN(\AES_ENC/u0/u3/n852 ) );
OR2_X2 \AES_ENC/u0/u3/U259  ( .A1(\AES_ENC/u0/u3/n1023 ), .A2(\AES_ENC/u0/u3/n617 ), .ZN(\AES_ENC/u0/u3/n819 ) );
OR2_X2 \AES_ENC/u0/u3/U257  ( .A1(\AES_ENC/u0/u3/n570 ), .A2(\AES_ENC/u0/u3/n930 ), .ZN(\AES_ENC/u0/u3/n818 ) );
NAND2_X2 \AES_ENC/u0/u3/U256  ( .A1(\AES_ENC/u0/u3/n1013 ), .A2(\AES_ENC/u0/u3/n1094 ), .ZN(\AES_ENC/u0/u3/n817 ) );
NAND4_X2 \AES_ENC/u0/u3/U249  ( .A1(\AES_ENC/u0/u3/n819 ), .A2(\AES_ENC/u0/u3/n818 ), .A3(\AES_ENC/u0/u3/n817 ), .A4(\AES_ENC/u0/u3/n816 ), .ZN(\AES_ENC/u0/u3/n820 ) );
NAND2_X2 \AES_ENC/u0/u3/U248  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n820 ), .ZN(\AES_ENC/u0/u3/n851 ) );
NAND2_X2 \AES_ENC/u0/u3/U247  ( .A1(\AES_ENC/u0/u3/n956 ), .A2(\AES_ENC/u0/u3/n1080 ), .ZN(\AES_ENC/u0/u3/n835 ) );
NAND2_X2 \AES_ENC/u0/u3/U246  ( .A1(\AES_ENC/u0/u3/n570 ), .A2(\AES_ENC/u0/u3/n1030 ), .ZN(\AES_ENC/u0/u3/n1047 ) );
OR2_X2 \AES_ENC/u0/u3/U245  ( .A1(\AES_ENC/u0/u3/n1047 ), .A2(\AES_ENC/u0/u3/n612 ), .ZN(\AES_ENC/u0/u3/n834 ) );
NAND2_X2 \AES_ENC/u0/u3/U244  ( .A1(\AES_ENC/u0/u3/n1072 ), .A2(\AES_ENC/u0/u3/n589 ), .ZN(\AES_ENC/u0/u3/n833 ) );
NAND4_X2 \AES_ENC/u0/u3/U233  ( .A1(\AES_ENC/u0/u3/n835 ), .A2(\AES_ENC/u0/u3/n834 ), .A3(\AES_ENC/u0/u3/n833 ), .A4(\AES_ENC/u0/u3/n832 ), .ZN(\AES_ENC/u0/u3/n836 ) );
NAND2_X2 \AES_ENC/u0/u3/U232  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n836 ), .ZN(\AES_ENC/u0/u3/n850 ) );
NAND2_X2 \AES_ENC/u0/u3/U231  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n623 ), .ZN(\AES_ENC/u0/u3/n847 ) );
NAND2_X2 \AES_ENC/u0/u3/U230  ( .A1(\AES_ENC/u0/u3/n1050 ), .A2(\AES_ENC/u0/u3/n1071 ), .ZN(\AES_ENC/u0/u3/n846 ) );
OR2_X2 \AES_ENC/u0/u3/U224  ( .A1(\AES_ENC/u0/u3/n1053 ), .A2(\AES_ENC/u0/u3/n911 ), .ZN(\AES_ENC/u0/u3/n1077 ) );
NAND4_X2 \AES_ENC/u0/u3/U220  ( .A1(\AES_ENC/u0/u3/n847 ), .A2(\AES_ENC/u0/u3/n846 ), .A3(\AES_ENC/u0/u3/n845 ), .A4(\AES_ENC/u0/u3/n844 ), .ZN(\AES_ENC/u0/u3/n848 ) );
NAND2_X2 \AES_ENC/u0/u3/U219  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n848 ), .ZN(\AES_ENC/u0/u3/n849 ) );
NAND4_X2 \AES_ENC/u0/u3/U218  ( .A1(\AES_ENC/u0/u3/n852 ), .A2(\AES_ENC/u0/u3/n851 ), .A3(\AES_ENC/u0/u3/n850 ), .A4(\AES_ENC/u0/u3/n849 ), .ZN(\AES_ENC/u0/subword[3] ) );
NAND2_X2 \AES_ENC/u0/u3/U216  ( .A1(\AES_ENC/u0/u3/n1009 ), .A2(\AES_ENC/u0/u3/n1072 ), .ZN(\AES_ENC/u0/u3/n862 ) );
NAND2_X2 \AES_ENC/u0/u3/U215  ( .A1(\AES_ENC/u0/u3/n603 ), .A2(\AES_ENC/u0/u3/n577 ), .ZN(\AES_ENC/u0/u3/n853 ) );
NAND2_X2 \AES_ENC/u0/u3/U214  ( .A1(\AES_ENC/u0/u3/n1050 ), .A2(\AES_ENC/u0/u3/n853 ), .ZN(\AES_ENC/u0/u3/n861 ) );
NAND4_X2 \AES_ENC/u0/u3/U206  ( .A1(\AES_ENC/u0/u3/n862 ), .A2(\AES_ENC/u0/u3/n861 ), .A3(\AES_ENC/u0/u3/n860 ), .A4(\AES_ENC/u0/u3/n859 ), .ZN(\AES_ENC/u0/u3/n863 ) );
NAND2_X2 \AES_ENC/u0/u3/U205  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n863 ), .ZN(\AES_ENC/u0/u3/n905 ) );
NAND2_X2 \AES_ENC/u0/u3/U204  ( .A1(\AES_ENC/u0/u3/n1010 ), .A2(\AES_ENC/u0/u3/n989 ), .ZN(\AES_ENC/u0/u3/n874 ) );
NAND2_X2 \AES_ENC/u0/u3/U203  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n610 ), .ZN(\AES_ENC/u0/u3/n864 ) );
NAND2_X2 \AES_ENC/u0/u3/U202  ( .A1(\AES_ENC/u0/u3/n929 ), .A2(\AES_ENC/u0/u3/n864 ), .ZN(\AES_ENC/u0/u3/n873 ) );
NAND4_X2 \AES_ENC/u0/u3/U193  ( .A1(\AES_ENC/u0/u3/n874 ), .A2(\AES_ENC/u0/u3/n873 ), .A3(\AES_ENC/u0/u3/n872 ), .A4(\AES_ENC/u0/u3/n871 ), .ZN(\AES_ENC/u0/u3/n875 ) );
NAND2_X2 \AES_ENC/u0/u3/U192  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n875 ), .ZN(\AES_ENC/u0/u3/n904 ) );
NAND2_X2 \AES_ENC/u0/u3/U191  ( .A1(\AES_ENC/u0/u3/n583 ), .A2(\AES_ENC/u0/u3/n1050 ), .ZN(\AES_ENC/u0/u3/n889 ) );
NAND2_X2 \AES_ENC/u0/u3/U190  ( .A1(\AES_ENC/u0/u3/n1093 ), .A2(\AES_ENC/u0/u3/n587 ), .ZN(\AES_ENC/u0/u3/n876 ) );
NAND2_X2 \AES_ENC/u0/u3/U189  ( .A1(\AES_ENC/u0/u3/n604 ), .A2(\AES_ENC/u0/u3/n876 ), .ZN(\AES_ENC/u0/u3/n877 ) );
NAND2_X2 \AES_ENC/u0/u3/U188  ( .A1(\AES_ENC/u0/u3/n877 ), .A2(\AES_ENC/u0/u3/n623 ), .ZN(\AES_ENC/u0/u3/n888 ) );
NAND4_X2 \AES_ENC/u0/u3/U179  ( .A1(\AES_ENC/u0/u3/n889 ), .A2(\AES_ENC/u0/u3/n888 ), .A3(\AES_ENC/u0/u3/n887 ), .A4(\AES_ENC/u0/u3/n886 ), .ZN(\AES_ENC/u0/u3/n890 ) );
NAND2_X2 \AES_ENC/u0/u3/U178  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n890 ), .ZN(\AES_ENC/u0/u3/n903 ) );
OR2_X2 \AES_ENC/u0/u3/U177  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n1059 ), .ZN(\AES_ENC/u0/u3/n900 ) );
NAND2_X2 \AES_ENC/u0/u3/U176  ( .A1(\AES_ENC/u0/u3/n1073 ), .A2(\AES_ENC/u0/u3/n1047 ), .ZN(\AES_ENC/u0/u3/n899 ) );
NAND2_X2 \AES_ENC/u0/u3/U175  ( .A1(\AES_ENC/u0/u3/n1094 ), .A2(\AES_ENC/u0/u3/n595 ), .ZN(\AES_ENC/u0/u3/n898 ) );
NAND4_X2 \AES_ENC/u0/u3/U167  ( .A1(\AES_ENC/u0/u3/n900 ), .A2(\AES_ENC/u0/u3/n899 ), .A3(\AES_ENC/u0/u3/n898 ), .A4(\AES_ENC/u0/u3/n897 ), .ZN(\AES_ENC/u0/u3/n901 ) );
NAND2_X2 \AES_ENC/u0/u3/U166  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n901 ), .ZN(\AES_ENC/u0/u3/n902 ) );
NAND4_X2 \AES_ENC/u0/u3/U165  ( .A1(\AES_ENC/u0/u3/n905 ), .A2(\AES_ENC/u0/u3/n904 ), .A3(\AES_ENC/u0/u3/n903 ), .A4(\AES_ENC/u0/u3/n902 ), .ZN(\AES_ENC/u0/subword[4] ) );
NAND2_X2 \AES_ENC/u0/u3/U164  ( .A1(\AES_ENC/u0/u3/n1094 ), .A2(\AES_ENC/u0/u3/n599 ), .ZN(\AES_ENC/u0/u3/n922 ) );
NAND2_X2 \AES_ENC/u0/u3/U163  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n989 ), .ZN(\AES_ENC/u0/u3/n921 ) );
NAND4_X2 \AES_ENC/u0/u3/U151  ( .A1(\AES_ENC/u0/u3/n922 ), .A2(\AES_ENC/u0/u3/n921 ), .A3(\AES_ENC/u0/u3/n920 ), .A4(\AES_ENC/u0/u3/n919 ), .ZN(\AES_ENC/u0/u3/n923 ) );
NAND2_X2 \AES_ENC/u0/u3/U150  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n923 ), .ZN(\AES_ENC/u0/u3/n972 ) );
NAND2_X2 \AES_ENC/u0/u3/U149  ( .A1(\AES_ENC/u0/u3/n582 ), .A2(\AES_ENC/u0/u3/n619 ), .ZN(\AES_ENC/u0/u3/n924 ) );
NAND2_X2 \AES_ENC/u0/u3/U148  ( .A1(\AES_ENC/u0/u3/n1073 ), .A2(\AES_ENC/u0/u3/n924 ), .ZN(\AES_ENC/u0/u3/n939 ) );
NAND2_X2 \AES_ENC/u0/u3/U147  ( .A1(\AES_ENC/u0/u3/n926 ), .A2(\AES_ENC/u0/u3/n925 ), .ZN(\AES_ENC/u0/u3/n927 ) );
NAND2_X2 \AES_ENC/u0/u3/U146  ( .A1(\AES_ENC/u0/u3/n606 ), .A2(\AES_ENC/u0/u3/n927 ), .ZN(\AES_ENC/u0/u3/n928 ) );
NAND2_X2 \AES_ENC/u0/u3/U145  ( .A1(\AES_ENC/u0/u3/n928 ), .A2(\AES_ENC/u0/u3/n1080 ), .ZN(\AES_ENC/u0/u3/n938 ) );
OR2_X2 \AES_ENC/u0/u3/U144  ( .A1(\AES_ENC/u0/u3/n1117 ), .A2(\AES_ENC/u0/u3/n615 ), .ZN(\AES_ENC/u0/u3/n937 ) );
NAND4_X2 \AES_ENC/u0/u3/U139  ( .A1(\AES_ENC/u0/u3/n939 ), .A2(\AES_ENC/u0/u3/n938 ), .A3(\AES_ENC/u0/u3/n937 ), .A4(\AES_ENC/u0/u3/n936 ), .ZN(\AES_ENC/u0/u3/n940 ) );
NAND2_X2 \AES_ENC/u0/u3/U138  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n940 ), .ZN(\AES_ENC/u0/u3/n971 ) );
OR2_X2 \AES_ENC/u0/u3/U137  ( .A1(\AES_ENC/u0/u3/n605 ), .A2(\AES_ENC/u0/u3/n941 ), .ZN(\AES_ENC/u0/u3/n954 ) );
NAND2_X2 \AES_ENC/u0/u3/U136  ( .A1(\AES_ENC/u0/u3/n1096 ), .A2(\AES_ENC/u0/u3/n577 ), .ZN(\AES_ENC/u0/u3/n942 ) );
NAND2_X2 \AES_ENC/u0/u3/U135  ( .A1(\AES_ENC/u0/u3/n1048 ), .A2(\AES_ENC/u0/u3/n942 ), .ZN(\AES_ENC/u0/u3/n943 ) );
NAND2_X2 \AES_ENC/u0/u3/U134  ( .A1(\AES_ENC/u0/u3/n612 ), .A2(\AES_ENC/u0/u3/n943 ), .ZN(\AES_ENC/u0/u3/n944 ) );
NAND2_X2 \AES_ENC/u0/u3/U133  ( .A1(\AES_ENC/u0/u3/n944 ), .A2(\AES_ENC/u0/u3/n580 ), .ZN(\AES_ENC/u0/u3/n953 ) );
NAND4_X2 \AES_ENC/u0/u3/U125  ( .A1(\AES_ENC/u0/u3/n954 ), .A2(\AES_ENC/u0/u3/n953 ), .A3(\AES_ENC/u0/u3/n952 ), .A4(\AES_ENC/u0/u3/n951 ), .ZN(\AES_ENC/u0/u3/n955 ) );
NAND2_X2 \AES_ENC/u0/u3/U124  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n955 ), .ZN(\AES_ENC/u0/u3/n970 ) );
NAND2_X2 \AES_ENC/u0/u3/U123  ( .A1(\AES_ENC/u0/u3/n1094 ), .A2(\AES_ENC/u0/u3/n1071 ), .ZN(\AES_ENC/u0/u3/n967 ) );
NAND2_X2 \AES_ENC/u0/u3/U122  ( .A1(\AES_ENC/u0/u3/n956 ), .A2(\AES_ENC/u0/u3/n1030 ), .ZN(\AES_ENC/u0/u3/n966 ) );
NAND4_X2 \AES_ENC/u0/u3/U114  ( .A1(\AES_ENC/u0/u3/n967 ), .A2(\AES_ENC/u0/u3/n966 ), .A3(\AES_ENC/u0/u3/n965 ), .A4(\AES_ENC/u0/u3/n964 ), .ZN(\AES_ENC/u0/u3/n968 ) );
NAND2_X2 \AES_ENC/u0/u3/U113  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n968 ), .ZN(\AES_ENC/u0/u3/n969 ) );
NAND4_X2 \AES_ENC/u0/u3/U112  ( .A1(\AES_ENC/u0/u3/n972 ), .A2(\AES_ENC/u0/u3/n971 ), .A3(\AES_ENC/u0/u3/n970 ), .A4(\AES_ENC/u0/u3/n969 ), .ZN(\AES_ENC/u0/subword[5] ) );
NAND2_X2 \AES_ENC/u0/u3/U111  ( .A1(\AES_ENC/u0/u3/n570 ), .A2(\AES_ENC/u0/u3/n1097 ), .ZN(\AES_ENC/u0/u3/n973 ) );
NAND2_X2 \AES_ENC/u0/u3/U110  ( .A1(\AES_ENC/u0/u3/n1073 ), .A2(\AES_ENC/u0/u3/n973 ), .ZN(\AES_ENC/u0/u3/n987 ) );
NAND2_X2 \AES_ENC/u0/u3/U109  ( .A1(\AES_ENC/u0/u3/n974 ), .A2(\AES_ENC/u0/u3/n1077 ), .ZN(\AES_ENC/u0/u3/n975 ) );
NAND2_X2 \AES_ENC/u0/u3/U108  ( .A1(\AES_ENC/u0/u3/n613 ), .A2(\AES_ENC/u0/u3/n975 ), .ZN(\AES_ENC/u0/u3/n976 ) );
NAND2_X2 \AES_ENC/u0/u3/U107  ( .A1(\AES_ENC/u0/u3/n977 ), .A2(\AES_ENC/u0/u3/n976 ), .ZN(\AES_ENC/u0/u3/n986 ) );
NAND4_X2 \AES_ENC/u0/u3/U99  ( .A1(\AES_ENC/u0/u3/n987 ), .A2(\AES_ENC/u0/u3/n986 ), .A3(\AES_ENC/u0/u3/n985 ), .A4(\AES_ENC/u0/u3/n984 ), .ZN(\AES_ENC/u0/u3/n988 ) );
NAND2_X2 \AES_ENC/u0/u3/U98  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n988 ), .ZN(\AES_ENC/u0/u3/n1044 ) );
NAND2_X2 \AES_ENC/u0/u3/U97  ( .A1(\AES_ENC/u0/u3/n1073 ), .A2(\AES_ENC/u0/u3/n989 ), .ZN(\AES_ENC/u0/u3/n1004 ) );
NAND2_X2 \AES_ENC/u0/u3/U96  ( .A1(\AES_ENC/u0/u3/n1092 ), .A2(\AES_ENC/u0/u3/n619 ), .ZN(\AES_ENC/u0/u3/n1003 ) );
NAND4_X2 \AES_ENC/u0/u3/U85  ( .A1(\AES_ENC/u0/u3/n1004 ), .A2(\AES_ENC/u0/u3/n1003 ), .A3(\AES_ENC/u0/u3/n1002 ), .A4(\AES_ENC/u0/u3/n1001 ), .ZN(\AES_ENC/u0/u3/n1005 ) );
NAND2_X2 \AES_ENC/u0/u3/U84  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n1005 ), .ZN(\AES_ENC/u0/u3/n1043 ) );
NAND2_X2 \AES_ENC/u0/u3/U83  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n596 ), .ZN(\AES_ENC/u0/u3/n1020 ) );
NAND2_X2 \AES_ENC/u0/u3/U82  ( .A1(\AES_ENC/u0/u3/n1050 ), .A2(\AES_ENC/u0/u3/n624 ), .ZN(\AES_ENC/u0/u3/n1019 ) );
NAND2_X2 \AES_ENC/u0/u3/U77  ( .A1(\AES_ENC/u0/u3/n1059 ), .A2(\AES_ENC/u0/u3/n1114 ), .ZN(\AES_ENC/u0/u3/n1012 ) );
NAND2_X2 \AES_ENC/u0/u3/U76  ( .A1(\AES_ENC/u0/u3/n1010 ), .A2(\AES_ENC/u0/u3/n592 ), .ZN(\AES_ENC/u0/u3/n1011 ) );
NAND2_X2 \AES_ENC/u0/u3/U75  ( .A1(\AES_ENC/u0/u3/n1012 ), .A2(\AES_ENC/u0/u3/n1011 ), .ZN(\AES_ENC/u0/u3/n1016 ) );
NAND4_X2 \AES_ENC/u0/u3/U70  ( .A1(\AES_ENC/u0/u3/n1020 ), .A2(\AES_ENC/u0/u3/n1019 ), .A3(\AES_ENC/u0/u3/n1018 ), .A4(\AES_ENC/u0/u3/n1017 ), .ZN(\AES_ENC/u0/u3/n1021 ) );
NAND2_X2 \AES_ENC/u0/u3/U69  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n1021 ), .ZN(\AES_ENC/u0/u3/n1042 ) );
NAND2_X2 \AES_ENC/u0/u3/U68  ( .A1(\AES_ENC/u0/u3/n1022 ), .A2(\AES_ENC/u0/u3/n1093 ), .ZN(\AES_ENC/u0/u3/n1039 ) );
NAND2_X2 \AES_ENC/u0/u3/U67  ( .A1(\AES_ENC/u0/u3/n1050 ), .A2(\AES_ENC/u0/u3/n1023 ), .ZN(\AES_ENC/u0/u3/n1038 ) );
NAND2_X2 \AES_ENC/u0/u3/U66  ( .A1(\AES_ENC/u0/u3/n1024 ), .A2(\AES_ENC/u0/u3/n1071 ), .ZN(\AES_ENC/u0/u3/n1037 ) );
AND2_X2 \AES_ENC/u0/u3/U60  ( .A1(\AES_ENC/u0/u3/n1030 ), .A2(\AES_ENC/u0/u3/n602 ), .ZN(\AES_ENC/u0/u3/n1078 ) );
NAND4_X2 \AES_ENC/u0/u3/U56  ( .A1(\AES_ENC/u0/u3/n1039 ), .A2(\AES_ENC/u0/u3/n1038 ), .A3(\AES_ENC/u0/u3/n1037 ), .A4(\AES_ENC/u0/u3/n1036 ), .ZN(\AES_ENC/u0/u3/n1040 ) );
NAND2_X2 \AES_ENC/u0/u3/U55  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n1040 ), .ZN(\AES_ENC/u0/u3/n1041 ) );
NAND4_X2 \AES_ENC/u0/u3/U54  ( .A1(\AES_ENC/u0/u3/n1044 ), .A2(\AES_ENC/u0/u3/n1043 ), .A3(\AES_ENC/u0/u3/n1042 ), .A4(\AES_ENC/u0/u3/n1041 ), .ZN(\AES_ENC/u0/subword[6] ) );
NAND2_X2 \AES_ENC/u0/u3/U53  ( .A1(\AES_ENC/u0/u3/n1072 ), .A2(\AES_ENC/u0/u3/n1045 ), .ZN(\AES_ENC/u0/u3/n1068 ) );
NAND2_X2 \AES_ENC/u0/u3/U52  ( .A1(\AES_ENC/u0/u3/n1046 ), .A2(\AES_ENC/u0/u3/n582 ), .ZN(\AES_ENC/u0/u3/n1067 ) );
NAND2_X2 \AES_ENC/u0/u3/U51  ( .A1(\AES_ENC/u0/u3/n1094 ), .A2(\AES_ENC/u0/u3/n1047 ), .ZN(\AES_ENC/u0/u3/n1066 ) );
NAND4_X2 \AES_ENC/u0/u3/U40  ( .A1(\AES_ENC/u0/u3/n1068 ), .A2(\AES_ENC/u0/u3/n1067 ), .A3(\AES_ENC/u0/u3/n1066 ), .A4(\AES_ENC/u0/u3/n1065 ), .ZN(\AES_ENC/u0/u3/n1069 ) );
NAND2_X2 \AES_ENC/u0/u3/U39  ( .A1(\AES_ENC/u0/u3/n1070 ), .A2(\AES_ENC/u0/u3/n1069 ), .ZN(\AES_ENC/u0/u3/n1135 ) );
NAND2_X2 \AES_ENC/u0/u3/U38  ( .A1(\AES_ENC/u0/u3/n1072 ), .A2(\AES_ENC/u0/u3/n1071 ), .ZN(\AES_ENC/u0/u3/n1088 ) );
NAND2_X2 \AES_ENC/u0/u3/U37  ( .A1(\AES_ENC/u0/u3/n1073 ), .A2(\AES_ENC/u0/u3/n595 ), .ZN(\AES_ENC/u0/u3/n1087 ) );
NAND4_X2 \AES_ENC/u0/u3/U28  ( .A1(\AES_ENC/u0/u3/n1088 ), .A2(\AES_ENC/u0/u3/n1087 ), .A3(\AES_ENC/u0/u3/n1086 ), .A4(\AES_ENC/u0/u3/n1085 ), .ZN(\AES_ENC/u0/u3/n1089 ) );
NAND2_X2 \AES_ENC/u0/u3/U27  ( .A1(\AES_ENC/u0/u3/n1090 ), .A2(\AES_ENC/u0/u3/n1089 ), .ZN(\AES_ENC/u0/u3/n1134 ) );
NAND2_X2 \AES_ENC/u0/u3/U26  ( .A1(\AES_ENC/u0/u3/n1091 ), .A2(\AES_ENC/u0/u3/n1093 ), .ZN(\AES_ENC/u0/u3/n1111 ) );
NAND2_X2 \AES_ENC/u0/u3/U25  ( .A1(\AES_ENC/u0/u3/n1092 ), .A2(\AES_ENC/u0/u3/n1120 ), .ZN(\AES_ENC/u0/u3/n1110 ) );
AND2_X2 \AES_ENC/u0/u3/U22  ( .A1(\AES_ENC/u0/u3/n1097 ), .A2(\AES_ENC/u0/u3/n1096 ), .ZN(\AES_ENC/u0/u3/n1098 ) );
NAND4_X2 \AES_ENC/u0/u3/U14  ( .A1(\AES_ENC/u0/u3/n1111 ), .A2(\AES_ENC/u0/u3/n1110 ), .A3(\AES_ENC/u0/u3/n1109 ), .A4(\AES_ENC/u0/u3/n1108 ), .ZN(\AES_ENC/u0/u3/n1112 ) );
NAND2_X2 \AES_ENC/u0/u3/U13  ( .A1(\AES_ENC/u0/u3/n1113 ), .A2(\AES_ENC/u0/u3/n1112 ), .ZN(\AES_ENC/u0/u3/n1133 ) );
NAND2_X2 \AES_ENC/u0/u3/U12  ( .A1(\AES_ENC/u0/u3/n1115 ), .A2(\AES_ENC/u0/u3/n1114 ), .ZN(\AES_ENC/u0/u3/n1129 ) );
OR2_X2 \AES_ENC/u0/u3/U11  ( .A1(\AES_ENC/u0/u3/n608 ), .A2(\AES_ENC/u0/u3/n1116 ), .ZN(\AES_ENC/u0/u3/n1128 ) );
NAND4_X2 \AES_ENC/u0/u3/U3  ( .A1(\AES_ENC/u0/u3/n1129 ), .A2(\AES_ENC/u0/u3/n1128 ), .A3(\AES_ENC/u0/u3/n1127 ), .A4(\AES_ENC/u0/u3/n1126 ), .ZN(\AES_ENC/u0/u3/n1130 ) );
NAND2_X2 \AES_ENC/u0/u3/U2  ( .A1(\AES_ENC/u0/u3/n1131 ), .A2(\AES_ENC/u0/u3/n1130 ), .ZN(\AES_ENC/u0/u3/n1132 ) );
NAND4_X2 \AES_ENC/u0/u3/U1  ( .A1(\AES_ENC/u0/u3/n1135 ), .A2(\AES_ENC/u0/u3/n1134 ), .A3(\AES_ENC/u0/u3/n1133 ), .A4(\AES_ENC/u0/u3/n1132 ), .ZN(\AES_ENC/u0/subword[7] ) );
INV_X4 \AES_ENC/u0/r0/U41  ( .A(\AES_ENC/u0/r0/n32 ), .ZN(\AES_ENC/u0/r0/n38 ) );
INV_X4 \AES_ENC/u0/r0/U40  ( .A(\AES_ENC/u0/r0/n9 ), .ZN(\AES_ENC/u0/r0/n37 ) );
INV_X4 \AES_ENC/u0/r0/U39  ( .A(\AES_ENC/u0/r0/n11 ), .ZN(\AES_ENC/u0/r0/n36 ) );
NAND3_X2 \AES_ENC/u0/r0/U38  ( .A1(\AES_ENC/u0/r0/rcnt[0] ), .A2(\AES_ENC/u0/r0/n35 ), .A3(\AES_ENC/u0/r0/n17 ), .ZN(\AES_ENC/u0/r0/n19 ) );
NOR3_X2 \AES_ENC/u0/r0/U27  ( .A1(\AES_ENC/u0/r0/n38 ), .A2(\AES_ENC/u0/r0/n13 ), .A3(\AES_ENC/u0/r0/n36 ), .ZN(\AES_ENC/u0/r0/N49 ) );
NAND3_X2 \AES_ENC/u0/r0/U24  ( .A1(\AES_ENC/u0/r0/n16 ), .A2(\AES_ENC/u0/r0/rcnt[0] ), .A3(\AES_ENC/u0/r0/N54 ), .ZN(\AES_ENC/u0/r0/n12 ) );
NOR2_X2 \AES_ENC/u0/r0/U23  ( .A1(\AES_ENC/u0/n315 ), .A2(\AES_ENC/u0/r0/rcnt[0] ), .ZN(\AES_ENC/u0/r0/n32 ) );
NOR2_X2 \AES_ENC/u0/r0/U22  ( .A1(\AES_ENC/u0/r0/n24 ), .A2(\AES_ENC/u0/r0/n34 ), .ZN(\AES_ENC/u0/r0/n22 ) );
NOR2_X2 \AES_ENC/u0/r0/U20  ( .A1(\AES_ENC/u0/r0/n22 ), .A2(\AES_ENC/u0/r0/n23 ), .ZN(\AES_ENC/u0/r0/n9 ) );
NOR2_X2 \AES_ENC/u0/r0/U15  ( .A1(\AES_ENC/u0/r0/n11 ), .A2(\AES_ENC/u0/r0/n12 ), .ZN(\AES_ENC/u0/r0/N50 ) );
NOR2_X2 \AES_ENC/u0/r0/U12  ( .A1(\AES_ENC/u0/r0/n11 ), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/r0/N53 ) );
NOR3_X2 \AES_ENC/u0/r0/U11  ( .A1(\AES_ENC/u0/r0/n16 ), .A2(\AES_ENC/u0/r0/n9 ), .A3(\AES_ENC/u0/r0/n36 ), .ZN(\AES_ENC/u0/r0/n17 ) );
NOR2_X2 \AES_ENC/u0/r0/U7  ( .A1(\AES_ENC/u0/r0/n37 ), .A2(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/r0/N54 ) );
INV_X4 \AES_ENC/u0/r0/U6  ( .A(\AES_ENC/u0/n315 ), .ZN(\AES_ENC/u0/r0/n35 ));
XNOR2_X2 \AES_ENC/u0/r0/U37  ( .A(\AES_ENC/u0/r0/rcnt[1] ), .B(\AES_ENC/u0/r0/rcnt[0] ), .ZN(\AES_ENC/u0/r0/n11 ) );
XOR2_X2 \AES_ENC/u0/r0/U36  ( .A(\AES_ENC/u0/r0/n34 ), .B(\AES_ENC/u0/r0/n11 ), .Z(\AES_ENC/u0/r0/n26 ) );
NAND2_X2 \AES_ENC/u0/r0/U35  ( .A1(\AES_ENC/u0/r0/rcnt[0] ), .A2(\AES_ENC/u0/r0/rcnt[1] ), .ZN(\AES_ENC/u0/r0/n24 ) );
NAND2_X2 \AES_ENC/u0/r0/U34  ( .A1(\AES_ENC/u0/r0/rcnt[2] ), .A2(\AES_ENC/u0/r0/n36 ), .ZN(\AES_ENC/u0/r0/n29 ) );
NAND2_X2 \AES_ENC/u0/r0/U33  ( .A1(\AES_ENC/u0/r0/n24 ), .A2(\AES_ENC/u0/r0/n29 ), .ZN(\AES_ENC/u0/r0/n27 ) );
NAND2_X2 \AES_ENC/u0/r0/U32  ( .A1(\AES_ENC/u0/r0/n26 ), .A2(\AES_ENC/u0/r0/n27 ), .ZN(\AES_ENC/u0/r0/n28 ) );
NAND2_X2 \AES_ENC/u0/r0/U31  ( .A1(\AES_ENC/u0/r0/n35 ), .A2(\AES_ENC/u0/r0/n28 ), .ZN(\AES_ENC/u0/r0/N44 ) );
NAND4_X2 \AES_ENC/u0/r0/U30  ( .A1(\AES_ENC/u0/r0/n26 ), .A2(\AES_ENC/u0/r0/n27 ), .A3(\AES_ENC/u0/r0/n35 ), .A4(\AES_ENC/u0/r0/n33 ), .ZN(\AES_ENC/u0/r0/n7 ) );
OR3_X2 \AES_ENC/u0/r0/U29  ( .A1(\AES_ENC/u0/r0/n26 ), .A2(\AES_ENC/u0/n315 ), .A3(\AES_ENC/u0/r0/n27 ), .ZN(\AES_ENC/u0/r0/n25 ) );
NAND2_X2 \AES_ENC/u0/r0/U28  ( .A1(\AES_ENC/u0/r0/n7 ), .A2(\AES_ENC/u0/r0/n25 ), .ZN(\AES_ENC/u0/r0/N45 ) );
XOR2_X2 \AES_ENC/u0/r0/U26  ( .A(\AES_ENC/u0/r0/n33 ), .B(\AES_ENC/u0/r0/n22 ), .Z(\AES_ENC/u0/r0/n16 ) );
AND2_X2 \AES_ENC/u0/r0/U25  ( .A1(\AES_ENC/u0/r0/n24 ), .A2(\AES_ENC/u0/r0/n34 ), .ZN(\AES_ENC/u0/r0/n23 ) );
NAND2_X2 \AES_ENC/u0/r0/U21  ( .A1(\AES_ENC/u0/r0/n17 ), .A2(\AES_ENC/u0/r0/n32 ), .ZN(\AES_ENC/u0/r0/n20 ) );
NAND4_X2 \AES_ENC/u0/r0/U19  ( .A1(\AES_ENC/u0/r0/n16 ), .A2(\AES_ENC/u0/r0/N53 ), .A3(\AES_ENC/u0/r0/rcnt[0] ), .A4(\AES_ENC/u0/r0/n37 ), .ZN(\AES_ENC/u0/r0/n21 ) );
NAND2_X2 \AES_ENC/u0/r0/U18  ( .A1(\AES_ENC/u0/r0/n20 ), .A2(\AES_ENC/u0/r0/n21 ), .ZN(\AES_ENC/u0/r0/N46 ) );
AND3_X2 \AES_ENC/u0/r0/U17  ( .A1(\AES_ENC/u0/r0/n16 ), .A2(\AES_ENC/u0/r0/n36 ), .A3(\AES_ENC/u0/r0/n32 ), .ZN(\AES_ENC/u0/r0/n10 ) );
NAND2_X2 \AES_ENC/u0/r0/U16  ( .A1(\AES_ENC/u0/r0/n10 ), .A2(\AES_ENC/u0/r0/n37 ), .ZN(\AES_ENC/u0/r0/n18 ) );
NAND2_X2 \AES_ENC/u0/r0/U14  ( .A1(\AES_ENC/u0/r0/n18 ), .A2(\AES_ENC/u0/r0/n19 ), .ZN(\AES_ENC/u0/r0/N47 ) );
NAND2_X2 \AES_ENC/u0/r0/U13  ( .A1(\AES_ENC/u0/r0/n17 ), .A2(\AES_ENC/u0/r0/n35 ), .ZN(\AES_ENC/u0/r0/n14 ) );
OR2_X2 \AES_ENC/u0/r0/U10  ( .A1(\AES_ENC/u0/r0/n12 ), .A2(\AES_ENC/u0/r0/n36 ), .ZN(\AES_ENC/u0/r0/n15 ) );
NAND2_X2 \AES_ENC/u0/r0/U9  ( .A1(\AES_ENC/u0/r0/n14 ), .A2(\AES_ENC/u0/r0/n15 ), .ZN(\AES_ENC/u0/r0/N48 ) );
XOR2_X2 \AES_ENC/u0/r0/U8  ( .A(\AES_ENC/u0/r0/n33 ), .B(\AES_ENC/u0/r0/rcnt[2] ), .Z(\AES_ENC/u0/r0/n13 ) );
AND2_X2 \AES_ENC/u0/r0/U5  ( .A1(\AES_ENC/u0/r0/n9 ), .A2(\AES_ENC/u0/r0/n10 ), .ZN(\AES_ENC/u0/r0/N51 ) );
OR2_X2 \AES_ENC/u0/r0/U4  ( .A1(\AES_ENC/u0/r0/n33 ), .A2(\AES_ENC/u0/r0/N44 ), .ZN(\AES_ENC/u0/r0/n8 ) );
NAND2_X2 \AES_ENC/u0/r0/U3  ( .A1(\AES_ENC/u0/r0/n7 ), .A2(\AES_ENC/u0/r0/n8 ), .ZN(\AES_ENC/u0/r0/N55 ) );
DFF_X2 \AES_ENC/u0/r0/out_reg_1_  ( .D(\AES_ENC/u0/r0/N45 ), .CK(clk), .Q(\AES_ENC/u0/rcon [25]), .QN() );
DFF_X2 \AES_ENC/u0/r0/out_reg_2_  ( .D(\AES_ENC/u0/r0/N46 ), .CK(clk), .Q(\AES_ENC/u0/rcon [26]), .QN() );
DFF_X2 \AES_ENC/u0/r0/out_reg_3_  ( .D(\AES_ENC/u0/r0/N47 ), .CK(clk), .Q(\AES_ENC/u0/rcon [27]), .QN() );
DFF_X2 \AES_ENC/u0/r0/out_reg_4_  ( .D(\AES_ENC/u0/r0/N48 ), .CK(clk), .Q(\AES_ENC/u0/rcon [28]), .QN() );
DFF_X2 \AES_ENC/u0/r0/out_reg_6_  ( .D(\AES_ENC/u0/r0/N50 ), .CK(clk), .Q(\AES_ENC/u0/rcon [30]), .QN() );
DFF_X2 \AES_ENC/u0/r0/out_reg_5_  ( .D(\AES_ENC/u0/r0/N49 ), .CK(clk), .Q(\AES_ENC/u0/rcon [29]), .QN() );
DFF_X2 \AES_ENC/u0/r0/out_reg_7_  ( .D(\AES_ENC/u0/r0/N51 ), .CK(clk), .Q(\AES_ENC/u0/rcon [31]), .QN() );
DFF_X2 \AES_ENC/u0/r0/rcnt_reg_3_  ( .D(\AES_ENC/u0/r0/N55 ), .CK(clk), .Q(),.QN(\AES_ENC/u0/r0/n33 ) );
DFF_X2 \AES_ENC/u0/r0/out_reg_0_  ( .D(\AES_ENC/u0/r0/N44 ), .CK(clk), .Q(\AES_ENC/u0/rcon [24]), .QN() );
DFF_X2 \AES_ENC/u0/r0/rcnt_reg_2_  ( .D(\AES_ENC/u0/r0/N54 ), .CK(clk), .Q(\AES_ENC/u0/r0/rcnt[2] ), .QN(\AES_ENC/u0/r0/n34 ) );
DFF_X2 \AES_ENC/u0/r0/rcnt_reg_1_  ( .D(\AES_ENC/u0/r0/N53 ), .CK(clk), .Q(\AES_ENC/u0/r0/rcnt[1] ), .QN() );
DFF_X2 \AES_ENC/u0/r0/rcnt_reg_0_  ( .D(\AES_ENC/u0/r0/n32 ), .CK(clk), .Q(\AES_ENC/u0/r0/rcnt[0] ), .QN() );
INV_X4 \AES_ENC/us00/U575  ( .A(\AES_ENC/sa00 [7]), .ZN(\AES_ENC/us00/n627 ));
INV_X4 \AES_ENC/us00/U574  ( .A(\AES_ENC/us00/n79 ), .ZN(\AES_ENC/us00/n625 ) );
INV_X4 \AES_ENC/us00/U573  ( .A(\AES_ENC/sa00 [4]), .ZN(\AES_ENC/us00/n624 ));
INV_X4 \AES_ENC/us00/U572  ( .A(\AES_ENC/us00/n170 ), .ZN(\AES_ENC/us00/n622 ) );
INV_X4 \AES_ENC/us00/U571  ( .A(\AES_ENC/us00/n73 ), .ZN(\AES_ENC/us00/n620 ) );
INV_X4 \AES_ENC/us00/U570  ( .A(\AES_ENC/us00/n72 ), .ZN(\AES_ENC/us00/n619 ) );
INV_X4 \AES_ENC/us00/U569  ( .A(\AES_ENC/us00/n146 ), .ZN(\AES_ENC/us00/n618 ) );
INV_X4 \AES_ENC/us00/U568  ( .A(\AES_ENC/us00/n221 ), .ZN(\AES_ENC/us00/n616 ) );
INV_X4 \AES_ENC/us00/U567  ( .A(\AES_ENC/us00/n402 ), .ZN(\AES_ENC/us00/n614 ) );
INV_X4 \AES_ENC/us00/U566  ( .A(\AES_ENC/sa00 [2]), .ZN(\AES_ENC/us00/n611 ));
INV_X4 \AES_ENC/us00/U565  ( .A(\AES_ENC/us00/n396 ), .ZN(\AES_ENC/us00/n610 ) );
INV_X4 \AES_ENC/us00/U564  ( .A(\AES_ENC/us00/n271 ), .ZN(\AES_ENC/us00/n609 ) );
INV_X4 \AES_ENC/us00/U563  ( .A(\AES_ENC/us00/n417 ), .ZN(\AES_ENC/us00/n607 ) );
INV_X4 \AES_ENC/us00/U562  ( .A(\AES_ENC/us00/n173 ), .ZN(\AES_ENC/us00/n603 ) );
INV_X4 \AES_ENC/us00/U561  ( .A(\AES_ENC/us00/n91 ), .ZN(\AES_ENC/us00/n602 ) );
INV_X4 \AES_ENC/us00/U560  ( .A(\AES_ENC/us00/n267 ), .ZN(\AES_ENC/us00/n601 ) );
INV_X4 \AES_ENC/us00/U559  ( .A(\AES_ENC/us00/n138 ), .ZN(\AES_ENC/us00/n600 ) );
INV_X4 \AES_ENC/us00/U558  ( .A(\AES_ENC/us00/n140 ), .ZN(\AES_ENC/us00/n599 ) );
INV_X4 \AES_ENC/us00/U557  ( .A(\AES_ENC/us00/n315 ), .ZN(\AES_ENC/us00/n598 ) );
INV_X4 \AES_ENC/us00/U556  ( .A(\AES_ENC/us00/n270 ), .ZN(\AES_ENC/us00/n597 ) );
INV_X4 \AES_ENC/us00/U555  ( .A(\AES_ENC/us00/n218 ), .ZN(\AES_ENC/us00/n595 ) );
INV_X4 \AES_ENC/us00/U554  ( .A(\AES_ENC/us00/n163 ), .ZN(\AES_ENC/us00/n594 ) );
INV_X4 \AES_ENC/us00/U553  ( .A(\AES_ENC/us00/n90 ), .ZN(\AES_ENC/us00/n593 ) );
INV_X4 \AES_ENC/us00/U552  ( .A(\AES_ENC/us00/n186 ), .ZN(\AES_ENC/us00/n592 ) );
INV_X4 \AES_ENC/us00/U551  ( .A(\AES_ENC/us00/n205 ), .ZN(\AES_ENC/us00/n591 ) );
INV_X4 \AES_ENC/us00/U550  ( .A(\AES_ENC/us00/n136 ), .ZN(\AES_ENC/us00/n590 ) );
INV_X4 \AES_ENC/us00/U549  ( .A(\AES_ENC/us00/n120 ), .ZN(\AES_ENC/us00/n589 ) );
INV_X4 \AES_ENC/us00/U548  ( .A(\AES_ENC/us00/n141 ), .ZN(\AES_ENC/us00/n588 ) );
INV_X4 \AES_ENC/us00/U547  ( .A(\AES_ENC/us00/n370 ), .ZN(\AES_ENC/us00/n587 ) );
INV_X4 \AES_ENC/us00/U546  ( .A(\AES_ENC/us00/n203 ), .ZN(\AES_ENC/us00/n586 ) );
INV_X4 \AES_ENC/us00/U545  ( .A(\AES_ENC/us00/n375 ), .ZN(\AES_ENC/us00/n585 ) );
INV_X4 \AES_ENC/us00/U544  ( .A(\AES_ENC/us00/n286 ), .ZN(\AES_ENC/us00/n584 ) );
INV_X4 \AES_ENC/us00/U543  ( .A(\AES_ENC/us00/n290 ), .ZN(\AES_ENC/us00/n583 ) );
INV_X4 \AES_ENC/us00/U542  ( .A(\AES_ENC/us00/n316 ), .ZN(\AES_ENC/us00/n581 ) );
INV_X4 \AES_ENC/us00/U541  ( .A(\AES_ENC/us00/n182 ), .ZN(\AES_ENC/us00/n580 ) );
INV_X4 \AES_ENC/us00/U540  ( .A(\AES_ENC/us00/n102 ), .ZN(\AES_ENC/us00/n579 ) );
INV_X4 \AES_ENC/us00/U539  ( .A(\AES_ENC/us00/n372 ), .ZN(\AES_ENC/us00/n578 ) );
INV_X4 \AES_ENC/us00/U538  ( .A(\AES_ENC/us00/n103 ), .ZN(\AES_ENC/us00/n577 ) );
INV_X4 \AES_ENC/us00/U537  ( .A(\AES_ENC/us00/n114 ), .ZN(\AES_ENC/us00/n576 ) );
INV_X4 \AES_ENC/us00/U536  ( .A(\AES_ENC/us00/n237 ), .ZN(\AES_ENC/us00/n575 ) );
INV_X4 \AES_ENC/us00/U535  ( .A(\AES_ENC/sa00 [0]), .ZN(\AES_ENC/us00/n574 ));
NOR2_X2 \AES_ENC/us00/U534  ( .A1(\AES_ENC/sa00 [0]), .A2(\AES_ENC/sa00 [6]),.ZN(\AES_ENC/us00/n104 ) );
NOR2_X2 \AES_ENC/us00/U533  ( .A1(\AES_ENC/us00/n574 ), .A2(\AES_ENC/sa00 [6]), .ZN(\AES_ENC/us00/n124 ) );
NOR2_X2 \AES_ENC/us00/U532  ( .A1(\AES_ENC/sa00 [4]), .A2(\AES_ENC/sa00 [3]),.ZN(\AES_ENC/us00/n170 ) );
INV_X4 \AES_ENC/us00/U531  ( .A(\AES_ENC/us00/n569 ), .ZN(\AES_ENC/us00/n572 ) );
NOR2_X2 \AES_ENC/us00/U530  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n431 ) );
NOR2_X2 \AES_ENC/us00/U529  ( .A1(\AES_ENC/sa00 [4]), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n432 ) );
NOR2_X2 \AES_ENC/us00/U528  ( .A1(\AES_ENC/us00/n431 ), .A2(\AES_ENC/us00/n432 ), .ZN(\AES_ENC/us00/n430 ) );
NOR2_X2 \AES_ENC/us00/U527  ( .A1(\AES_ENC/us00/n430 ), .A2(\AES_ENC/us00/n575 ), .ZN(\AES_ENC/us00/n429 ) );
NOR3_X2 \AES_ENC/us00/U526  ( .A1(\AES_ENC/us00/n627 ), .A2(\AES_ENC/sa00 [5]), .A3(\AES_ENC/us00/n492 ), .ZN(\AES_ENC/us00/n490 ));
NOR2_X2 \AES_ENC/us00/U525  ( .A1(\AES_ENC/us00/n76 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n489 ) );
NOR2_X2 \AES_ENC/us00/U524  ( .A1(\AES_ENC/sa00 [4]), .A2(\AES_ENC/us00/n579 ), .ZN(\AES_ENC/us00/n491 ) );
NOR3_X2 \AES_ENC/us00/U523  ( .A1(\AES_ENC/us00/n489 ), .A2(\AES_ENC/us00/n490 ), .A3(\AES_ENC/us00/n491 ), .ZN(\AES_ENC/us00/n483 ) );
INV_X4 \AES_ENC/us00/U522  ( .A(\AES_ENC/sa00 [3]), .ZN(\AES_ENC/us00/n621 ));
NAND3_X2 \AES_ENC/us00/U521  ( .A1(\AES_ENC/us00/n544 ), .A2(\AES_ENC/us00/n626 ), .A3(\AES_ENC/sa00 [7]), .ZN(\AES_ENC/us00/n543 ));
NOR2_X2 \AES_ENC/us00/U520  ( .A1(\AES_ENC/us00/n611 ), .A2(\AES_ENC/sa00 [5]), .ZN(\AES_ENC/us00/n271 ) );
NOR2_X2 \AES_ENC/us00/U519  ( .A1(\AES_ENC/sa00 [5]), .A2(\AES_ENC/sa00 [2]),.ZN(\AES_ENC/us00/n221 ) );
INV_X4 \AES_ENC/us00/U518  ( .A(\AES_ENC/sa00 [5]), .ZN(\AES_ENC/us00/n626 ));
NOR2_X2 \AES_ENC/us00/U517  ( .A1(\AES_ENC/us00/n611 ), .A2(\AES_ENC/sa00 [7]), .ZN(\AES_ENC/us00/n417 ) );
NAND3_X2 \AES_ENC/us00/U516  ( .A1(\AES_ENC/us00/n517 ), .A2(\AES_ENC/us00/n518 ), .A3(\AES_ENC/us00/n519 ), .ZN(\AES_ENC/sa00_sub[0] ) );
NOR2_X2 \AES_ENC/us00/U515  ( .A1(\AES_ENC/us00/n626 ), .A2(\AES_ENC/sa00 [2]), .ZN(\AES_ENC/us00/n146 ) );
NOR4_X2 \AES_ENC/us00/U512  ( .A1(\AES_ENC/us00/n563 ), .A2(\AES_ENC/us00/n564 ), .A3(\AES_ENC/us00/n565 ), .A4(\AES_ENC/us00/n566 ), .ZN(\AES_ENC/us00/n562 ) );
NOR2_X2 \AES_ENC/us00/U510  ( .A1(\AES_ENC/us00/n567 ), .A2(\AES_ENC/us00/n568 ), .ZN(\AES_ENC/us00/n561 ) );
NAND3_X2 \AES_ENC/us00/U509  ( .A1(\AES_ENC/sa00 [2]), .A2(\AES_ENC/sa00 [7]), .A3(\AES_ENC/us00/n135 ), .ZN(\AES_ENC/us00/n560 ) );
NOR2_X2 \AES_ENC/us00/U508  ( .A1(\AES_ENC/sa00 [7]), .A2(\AES_ENC/sa00 [2]),.ZN(\AES_ENC/us00/n402 ) );
NOR2_X2 \AES_ENC/us00/U507  ( .A1(\AES_ENC/sa00 [4]), .A2(\AES_ENC/sa00 [1]),.ZN(\AES_ENC/us00/n91 ) );
NOR2_X2 \AES_ENC/us00/U506  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/sa00 [3]), .ZN(\AES_ENC/us00/n141 ) );
NOR2_X2 \AES_ENC/us00/U505  ( .A1(\AES_ENC/us00/n607 ), .A2(\AES_ENC/sa00 [5]), .ZN(\AES_ENC/us00/n171 ) );
NOR2_X2 \AES_ENC/us00/U504  ( .A1(\AES_ENC/us00/n625 ), .A2(\AES_ENC/sa00 [2]), .ZN(\AES_ENC/us00/n101 ) );
NOR2_X2 \AES_ENC/us00/U503  ( .A1(\AES_ENC/us00/n614 ), .A2(\AES_ENC/sa00 [5]), .ZN(\AES_ENC/us00/n100 ) );
NOR2_X2 \AES_ENC/us00/U502  ( .A1(\AES_ENC/us00/n624 ), .A2(\AES_ENC/sa00 [3]), .ZN(\AES_ENC/us00/n265 ) );
INV_X4 \AES_ENC/us00/U501  ( .A(\AES_ENC/us00/n570 ), .ZN(\AES_ENC/us00/n573 ) );
NOR2_X2 \AES_ENC/us00/U500  ( .A1(\AES_ENC/us00/n141 ), .A2(\AES_ENC/us00/n99 ), .ZN(\AES_ENC/us00/n557 ) );
NOR3_X2 \AES_ENC/us00/U499  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n573 ), .A3(\AES_ENC/us00/n120 ), .ZN(\AES_ENC/us00/n555 ) );
NOR2_X2 \AES_ENC/us00/U498  ( .A1(\AES_ENC/us00/n557 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n556 ) );
NOR2_X2 \AES_ENC/us00/U497  ( .A1(\AES_ENC/us00/n555 ), .A2(\AES_ENC/us00/n556 ), .ZN(\AES_ENC/us00/n550 ) );
NOR3_X2 \AES_ENC/us00/U496  ( .A1(\AES_ENC/us00/n200 ), .A2(\AES_ENC/us00/n586 ), .A3(\AES_ENC/us00/n201 ), .ZN(\AES_ENC/us00/n193 ) );
NOR2_X2 \AES_ENC/us00/U495  ( .A1(\AES_ENC/us00/n287 ), .A2(\AES_ENC/us00/n288 ), .ZN(\AES_ENC/us00/n276 ) );
NOR2_X2 \AES_ENC/us00/U494  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n373 ) );
NOR2_X2 \AES_ENC/us00/U492  ( .A1(\AES_ENC/us00/n624 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n374 ) );
NOR2_X2 \AES_ENC/us00/U491  ( .A1(\AES_ENC/us00/n373 ), .A2(\AES_ENC/us00/n374 ), .ZN(\AES_ENC/us00/n371 ) );
NOR2_X2 \AES_ENC/us00/U490  ( .A1(\AES_ENC/sa00 [1]), .A2(\AES_ENC/us00/n623 ), .ZN(\AES_ENC/us00/n283 ) );
NOR2_X2 \AES_ENC/us00/U489  ( .A1(\AES_ENC/us00/n283 ), .A2(\AES_ENC/us00/n103 ), .ZN(\AES_ENC/us00/n282 ) );
NOR2_X2 \AES_ENC/us00/U488  ( .A1(\AES_ENC/us00/n370 ), .A2(\AES_ENC/us00/n572 ), .ZN(\AES_ENC/us00/n369 ) );
NOR3_X2 \AES_ENC/us00/U487  ( .A1(\AES_ENC/us00/n427 ), .A2(\AES_ENC/us00/n428 ), .A3(\AES_ENC/us00/n429 ), .ZN(\AES_ENC/us00/n421 ) );
NOR2_X2 \AES_ENC/us00/U486  ( .A1(\AES_ENC/us00/n138 ), .A2(\AES_ENC/us00/n141 ), .ZN(\AES_ENC/us00/n447 ) );
NOR2_X2 \AES_ENC/us00/U483  ( .A1(\AES_ENC/us00/n447 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n444 ) );
INV_X4 \AES_ENC/us00/U482  ( .A(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n596 ));
NOR2_X2 \AES_ENC/us00/U480  ( .A1(\AES_ENC/us00/n140 ), .A2(\AES_ENC/us00/n141 ), .ZN(\AES_ENC/us00/n139 ) );
OR2_X4 \AES_ENC/us00/U479  ( .A1(\AES_ENC/us00/n100 ), .A2(\AES_ENC/us00/n101 ), .ZN(\AES_ENC/us00/n571 ) );
AND2_X2 \AES_ENC/us00/U478  ( .A1(\AES_ENC/us00/n571 ), .A2(\AES_ENC/us00/n99 ), .ZN(\AES_ENC/us00/n92 ) );
NOR2_X2 \AES_ENC/us00/U477  ( .A1(\AES_ENC/us00/n120 ), .A2(\AES_ENC/us00/n265 ), .ZN(\AES_ENC/us00/n400 ) );
NOR2_X2 \AES_ENC/us00/U474  ( .A1(\AES_ENC/us00/n400 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n399 ) );
NOR2_X2 \AES_ENC/us00/U473  ( .A1(\AES_ENC/us00/n264 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n263 ) );
NOR2_X2 \AES_ENC/us00/U472  ( .A1(\AES_ENC/us00/n267 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n261 ) );
NOR2_X2 \AES_ENC/us00/U471  ( .A1(\AES_ENC/us00/n265 ), .A2(\AES_ENC/us00/n266 ), .ZN(\AES_ENC/us00/n262 ) );
NOR3_X2 \AES_ENC/us00/U470  ( .A1(\AES_ENC/us00/n261 ), .A2(\AES_ENC/us00/n262 ), .A3(\AES_ENC/us00/n263 ), .ZN(\AES_ENC/us00/n260 ) );
NOR2_X2 \AES_ENC/us00/U469  ( .A1(\AES_ENC/us00/n624 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n119 ) );
NOR2_X2 \AES_ENC/us00/U468  ( .A1(\AES_ENC/us00/n572 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n247 ) );
NOR2_X2 \AES_ENC/us00/U467  ( .A1(\AES_ENC/us00/n145 ), .A2(\AES_ENC/us00/n618 ), .ZN(\AES_ENC/us00/n143 ) );
NOR2_X2 \AES_ENC/us00/U466  ( .A1(\AES_ENC/us00/n143 ), .A2(\AES_ENC/us00/n144 ), .ZN(\AES_ENC/us00/n142 ) );
NOR2_X2 \AES_ENC/us00/U465  ( .A1(\AES_ENC/us00/n142 ), .A2(\AES_ENC/us00/n592 ), .ZN(\AES_ENC/us00/n130 ) );
NOR2_X2 \AES_ENC/us00/U464  ( .A1(\AES_ENC/sa00 [1]), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n565 ) );
NOR2_X2 \AES_ENC/us00/U463  ( .A1(\AES_ENC/us00/n170 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n215 ) );
NOR2_X2 \AES_ENC/us00/U462  ( .A1(\AES_ENC/us00/n121 ), .A2(\AES_ENC/us00/n100 ), .ZN(\AES_ENC/us00/n401 ) );
NOR2_X2 \AES_ENC/us00/U461  ( .A1(\AES_ENC/us00/n401 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n397 ) );
NOR2_X2 \AES_ENC/us00/U460  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n214 ) );
NOR2_X2 \AES_ENC/us00/U459  ( .A1(\AES_ENC/us00/n91 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n553 ) );
NOR2_X2 \AES_ENC/us00/U458  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n621 ), .ZN(\AES_ENC/us00/n554 ) );
NOR2_X2 \AES_ENC/us00/U455  ( .A1(\AES_ENC/us00/n285 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n552 ) );
NOR4_X2 \AES_ENC/us00/U448  ( .A1(\AES_ENC/us00/n552 ), .A2(\AES_ENC/us00/n553 ), .A3(\AES_ENC/us00/n392 ), .A4(\AES_ENC/us00/n554 ), .ZN(\AES_ENC/us00/n551 ) );
NOR2_X2 \AES_ENC/us00/U447  ( .A1(\AES_ENC/us00/n91 ), .A2(\AES_ENC/us00/n286 ), .ZN(\AES_ENC/us00/n264 ) );
NOR2_X2 \AES_ENC/us00/U442  ( .A1(\AES_ENC/us00/n91 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n441 ) );
NOR2_X2 \AES_ENC/us00/U441  ( .A1(\AES_ENC/us00/n265 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n453 ) );
NOR2_X2 \AES_ENC/us00/U438  ( .A1(\AES_ENC/us00/n122 ), .A2(\AES_ENC/us00/n100 ), .ZN(\AES_ENC/us00/n266 ) );
NOR2_X2 \AES_ENC/us00/U435  ( .A1(\AES_ENC/us00/n120 ), .A2(\AES_ENC/us00/n170 ), .ZN(\AES_ENC/us00/n305 ) );
NOR2_X2 \AES_ENC/us00/U434  ( .A1(\AES_ENC/us00/n305 ), .A2(\AES_ENC/us00/n609 ), .ZN(\AES_ENC/us00/n302 ) );
NOR3_X2 \AES_ENC/us00/U433  ( .A1(\AES_ENC/us00/n623 ), .A2(\AES_ENC/sa00 [1]), .A3(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n513 ));
INV_X4 \AES_ENC/us00/U428  ( .A(\AES_ENC/us00/n265 ), .ZN(\AES_ENC/us00/n623 ) );
NOR2_X2 \AES_ENC/us00/U427  ( .A1(\AES_ENC/us00/n199 ), .A2(\AES_ENC/us00/n265 ), .ZN(\AES_ENC/us00/n492 ) );
NOR2_X2 \AES_ENC/us00/U421  ( .A1(\AES_ENC/us00/n265 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n511 ) );
NOR2_X2 \AES_ENC/us00/U420  ( .A1(\AES_ENC/us00/n165 ), .A2(\AES_ENC/us00/n170 ), .ZN(\AES_ENC/us00/n115 ) );
NOR3_X2 \AES_ENC/us00/U419  ( .A1(\AES_ENC/us00/n589 ), .A2(\AES_ENC/us00/n170 ), .A3(\AES_ENC/us00/n616 ), .ZN(\AES_ENC/us00/n251 ) );
NOR2_X2 \AES_ENC/us00/U418  ( .A1(\AES_ENC/us00/n626 ), .A2(\AES_ENC/us00/n611 ), .ZN(\AES_ENC/us00/n396 ) );
NOR3_X2 \AES_ENC/us00/U417  ( .A1(\AES_ENC/us00/n590 ), .A2(\AES_ENC/us00/n627 ), .A3(\AES_ENC/us00/n611 ), .ZN(\AES_ENC/us00/n398 ) );
NOR3_X2 \AES_ENC/us00/U416  ( .A1(\AES_ENC/us00/n610 ), .A2(\AES_ENC/us00/n572 ), .A3(\AES_ENC/us00/n575 ), .ZN(\AES_ENC/us00/n233 ) );
NOR3_X2 \AES_ENC/us00/U415  ( .A1(\AES_ENC/us00/n237 ), .A2(\AES_ENC/us00/n572 ), .A3(\AES_ENC/us00/n609 ), .ZN(\AES_ENC/us00/n428 ) );
NOR3_X2 \AES_ENC/us00/U414  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n572 ), .A3(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n502 ) );
NOR3_X2 \AES_ENC/us00/U413  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n572 ), .A3(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n301 ) );
NOR3_X2 \AES_ENC/us00/U410  ( .A1(\AES_ENC/us00/n187 ), .A2(\AES_ENC/us00/n188 ), .A3(\AES_ENC/us00/n189 ), .ZN(\AES_ENC/us00/n177 ) );
NOR4_X2 \AES_ENC/us00/U409  ( .A1(\AES_ENC/us00/n390 ), .A2(\AES_ENC/us00/n391 ), .A3(\AES_ENC/us00/n392 ), .A4(\AES_ENC/us00/n393 ), .ZN(\AES_ENC/us00/n389 ) );
NOR3_X2 \AES_ENC/us00/U406  ( .A1(\AES_ENC/us00/n397 ), .A2(\AES_ENC/us00/n398 ), .A3(\AES_ENC/us00/n399 ), .ZN(\AES_ENC/us00/n388 ) );
NOR2_X2 \AES_ENC/us00/U405  ( .A1(\AES_ENC/us00/n527 ), .A2(\AES_ENC/us00/n528 ), .ZN(\AES_ENC/us00/n523 ) );
NOR4_X2 \AES_ENC/us00/U404  ( .A1(\AES_ENC/us00/n250 ), .A2(\AES_ENC/us00/n148 ), .A3(\AES_ENC/us00/n525 ), .A4(\AES_ENC/us00/n526 ), .ZN(\AES_ENC/us00/n524 ) );
NOR3_X2 \AES_ENC/us00/U403  ( .A1(\AES_ENC/us00/n92 ), .A2(\AES_ENC/us00/n93 ), .A3(\AES_ENC/us00/n94 ), .ZN(\AES_ENC/us00/n84 ));
NOR4_X2 \AES_ENC/us00/U401  ( .A1(\AES_ENC/us00/n485 ), .A2(\AES_ENC/us00/n486 ), .A3(\AES_ENC/us00/n487 ), .A4(\AES_ENC/us00/n488 ), .ZN(\AES_ENC/us00/n484 ) );
NOR4_X2 \AES_ENC/us00/U400  ( .A1(\AES_ENC/us00/n353 ), .A2(\AES_ENC/us00/n354 ), .A3(\AES_ENC/us00/n355 ), .A4(\AES_ENC/us00/n356 ), .ZN(\AES_ENC/us00/n352 ) );
NOR4_X2 \AES_ENC/us00/U399  ( .A1(\AES_ENC/us00/n232 ), .A2(\AES_ENC/us00/n233 ), .A3(\AES_ENC/us00/n234 ), .A4(\AES_ENC/us00/n235 ), .ZN(\AES_ENC/us00/n231 ) );
NOR3_X2 \AES_ENC/us00/U398  ( .A1(\AES_ENC/us00/n453 ), .A2(\AES_ENC/us00/n454 ), .A3(\AES_ENC/us00/n455 ), .ZN(\AES_ENC/us00/n452 ) );
NOR2_X2 \AES_ENC/us00/U397  ( .A1(\AES_ENC/us00/n499 ), .A2(\AES_ENC/us00/n538 ), .ZN(\AES_ENC/us00/n537 ) );
NOR2_X2 \AES_ENC/us00/U396  ( .A1(\AES_ENC/us00/n598 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n311 ) );
NOR2_X2 \AES_ENC/us00/U393  ( .A1(\AES_ENC/us00/n623 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n314 ) );
NOR2_X2 \AES_ENC/us00/U390  ( .A1(\AES_ENC/us00/n141 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n312 ) );
NOR4_X2 \AES_ENC/us00/U389  ( .A1(\AES_ENC/us00/n311 ), .A2(\AES_ENC/us00/n312 ), .A3(\AES_ENC/us00/n313 ), .A4(\AES_ENC/us00/n314 ), .ZN(\AES_ENC/us00/n310 ) );
NOR2_X2 \AES_ENC/us00/U388  ( .A1(\AES_ENC/us00/n116 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n161 ) );
NOR2_X2 \AES_ENC/us00/U387  ( .A1(\AES_ENC/us00/n163 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n162 ) );
NOR3_X2 \AES_ENC/us00/U386  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n170 ), .A3(\AES_ENC/us00/n120 ), .ZN(\AES_ENC/us00/n159 ) );
NOR4_X2 \AES_ENC/us00/U385  ( .A1(\AES_ENC/us00/n159 ), .A2(\AES_ENC/us00/n160 ), .A3(\AES_ENC/us00/n161 ), .A4(\AES_ENC/us00/n162 ), .ZN(\AES_ENC/us00/n158 ) );
NOR2_X2 \AES_ENC/us00/U384  ( .A1(\AES_ENC/us00/n371 ), .A2(\AES_ENC/us00/n578 ), .ZN(\AES_ENC/us00/n366 ) );
NOR2_X2 \AES_ENC/us00/U383  ( .A1(\AES_ENC/us00/n369 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n367 ) );
NOR2_X2 \AES_ENC/us00/U382  ( .A1(\AES_ENC/us00/n572 ), .A2(\AES_ENC/us00/n579 ), .ZN(\AES_ENC/us00/n368 ) );
NOR4_X2 \AES_ENC/us00/U374  ( .A1(\AES_ENC/us00/n365 ), .A2(\AES_ENC/us00/n366 ), .A3(\AES_ENC/us00/n367 ), .A4(\AES_ENC/us00/n368 ), .ZN(\AES_ENC/us00/n364 ) );
NOR2_X2 \AES_ENC/us00/U373  ( .A1(\AES_ENC/us00/n606 ), .A2(\AES_ENC/us00/n582 ), .ZN(\AES_ENC/us00/n89 ) );
NOR2_X2 \AES_ENC/us00/U372  ( .A1(\AES_ENC/us00/n91 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n87 ) );
NOR2_X2 \AES_ENC/us00/U370  ( .A1(\AES_ENC/us00/n90 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n88 ) );
NOR4_X2 \AES_ENC/us00/U369  ( .A1(\AES_ENC/us00/n86 ), .A2(\AES_ENC/us00/n87 ), .A3(\AES_ENC/us00/n88 ), .A4(\AES_ENC/us00/n89 ),.ZN(\AES_ENC/us00/n85 ) );
NOR3_X2 \AES_ENC/us00/U368  ( .A1(\AES_ENC/us00/n237 ), .A2(\AES_ENC/us00/n621 ), .A3(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n232 ) );
NOR2_X2 \AES_ENC/us00/U367  ( .A1(\AES_ENC/us00/n626 ), .A2(\AES_ENC/us00/n627 ), .ZN(\AES_ENC/us00/n79 ) );
INV_X4 \AES_ENC/us00/U366  ( .A(\AES_ENC/us00/n171 ), .ZN(\AES_ENC/us00/n606 ) );
NOR3_X2 \AES_ENC/us00/U365  ( .A1(\AES_ENC/us00/n286 ), .A2(\AES_ENC/us00/n135 ), .A3(\AES_ENC/us00/n611 ), .ZN(\AES_ENC/us00/n78 ) );
INV_X4 \AES_ENC/us00/U364  ( .A(\AES_ENC/us00/n100 ), .ZN(\AES_ENC/us00/n613 ) );
NOR2_X2 \AES_ENC/us00/U363  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n265 ), .ZN(\AES_ENC/us00/n93 ) );
INV_X4 \AES_ENC/us00/U354  ( .A(\AES_ENC/us00/n101 ), .ZN(\AES_ENC/us00/n617 ) );
NOR2_X2 \AES_ENC/us00/U353  ( .A1(\AES_ENC/us00/n569 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n267 ) );
NOR2_X2 \AES_ENC/us00/U352  ( .A1(\AES_ENC/us00/n620 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n270 ) );
NOR2_X2 \AES_ENC/us00/U351  ( .A1(\AES_ENC/us00/n572 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n99 ) );
NOR2_X2 \AES_ENC/us00/U350  ( .A1(\AES_ENC/us00/n609 ), .A2(\AES_ENC/us00/n627 ), .ZN(\AES_ENC/us00/n185 ) );
NOR2_X2 \AES_ENC/us00/U349  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n90 ) );
NOR2_X2 \AES_ENC/us00/U348  ( .A1(\AES_ENC/us00/n622 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n135 ) );
NOR2_X2 \AES_ENC/us00/U347  ( .A1(\AES_ENC/sa00 [1]), .A2(\AES_ENC/us00/n73 ), .ZN(\AES_ENC/us00/n173 ) );
NOR2_X2 \AES_ENC/us00/U346  ( .A1(\AES_ENC/us00/n619 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n285 ) );
NOR2_X2 \AES_ENC/us00/U345  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/us00/n170 ), .ZN(\AES_ENC/us00/n370 ) );
NOR2_X2 \AES_ENC/us00/U338  ( .A1(\AES_ENC/us00/n626 ), .A2(\AES_ENC/us00/n607 ), .ZN(\AES_ENC/us00/n122 ) );
NOR2_X2 \AES_ENC/us00/U335  ( .A1(\AES_ENC/us00/n627 ), .A2(\AES_ENC/us00/n616 ), .ZN(\AES_ENC/us00/n240 ) );
NOR2_X2 \AES_ENC/us00/U329  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/us00/n624 ), .ZN(\AES_ENC/us00/n72 ) );
NOR2_X2 \AES_ENC/us00/U328  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/us00/n624 ), .ZN(\AES_ENC/us00/n136 ) );
NOR2_X2 \AES_ENC/us00/U327  ( .A1(\AES_ENC/us00/n625 ), .A2(\AES_ENC/us00/n611 ), .ZN(\AES_ENC/us00/n121 ) );
NOR2_X2 \AES_ENC/us00/U325  ( .A1(\AES_ENC/sa00 [1]), .A2(\AES_ENC/us00/n170 ), .ZN(\AES_ENC/us00/n140 ) );
NOR2_X2 \AES_ENC/us00/U324  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/us00/n265 ), .ZN(\AES_ENC/us00/n165 ) );
NOR2_X2 \AES_ENC/us00/U319  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n138 ) );
NOR2_X2 \AES_ENC/us00/U318  ( .A1(\AES_ENC/us00/n614 ), .A2(\AES_ENC/us00/n626 ), .ZN(\AES_ENC/us00/n144 ) );
NOR2_X2 \AES_ENC/us00/U317  ( .A1(\AES_ENC/us00/n72 ), .A2(\AES_ENC/us00/n170 ), .ZN(\AES_ENC/us00/n73 ) );
NOR2_X2 \AES_ENC/us00/U316  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/us00/n572 ), .ZN(\AES_ENC/us00/n120 ) );
NOR2_X2 \AES_ENC/us00/U315  ( .A1(\AES_ENC/us00/n136 ), .A2(\AES_ENC/us00/n140 ), .ZN(\AES_ENC/us00/n318 ) );
NOR2_X2 \AES_ENC/us00/U314  ( .A1(\AES_ENC/us00/n318 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n317 ) );
NOR2_X2 \AES_ENC/us00/U312  ( .A1(\AES_ENC/us00/n316 ), .A2(\AES_ENC/us00/n317 ), .ZN(\AES_ENC/us00/n309 ) );
NOR2_X2 \AES_ENC/us00/U311  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n588 ), .ZN(\AES_ENC/us00/n239 ) );
NOR2_X2 \AES_ENC/us00/U310  ( .A1(\AES_ENC/us00/n238 ), .A2(\AES_ENC/us00/n239 ), .ZN(\AES_ENC/us00/n230 ) );
NOR3_X2 \AES_ENC/us00/U309  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n103 ), .A3(\AES_ENC/us00/n173 ), .ZN(\AES_ENC/us00/n476 ) );
NOR3_X2 \AES_ENC/us00/U303  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n140 ), .A3(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n477 ) );
NOR2_X2 \AES_ENC/us00/U302  ( .A1(\AES_ENC/us00/n476 ), .A2(\AES_ENC/us00/n477 ), .ZN(\AES_ENC/us00/n470 ) );
NOR2_X2 \AES_ENC/us00/U300  ( .A1(\AES_ENC/us00/n614 ), .A2(\AES_ENC/us00/n591 ), .ZN(\AES_ENC/us00/n331 ) );
NOR2_X2 \AES_ENC/us00/U299  ( .A1(\AES_ENC/us00/n135 ), .A2(\AES_ENC/us00/n136 ), .ZN(\AES_ENC/us00/n134 ) );
NOR2_X2 \AES_ENC/us00/U298  ( .A1(\AES_ENC/us00/n99 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n528 ) );
NOR2_X2 \AES_ENC/us00/U297  ( .A1(\AES_ENC/us00/n285 ), .A2(\AES_ENC/us00/n286 ), .ZN(\AES_ENC/us00/n284 ) );
NOR2_X2 \AES_ENC/us00/U296  ( .A1(\AES_ENC/us00/n284 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n280 ) );
NOR2_X2 \AES_ENC/us00/U295  ( .A1(\AES_ENC/us00/n370 ), .A2(\AES_ENC/us00/n573 ), .ZN(\AES_ENC/us00/n446 ) );
NOR2_X2 \AES_ENC/us00/U294  ( .A1(\AES_ENC/us00/n446 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n445 ) );
NOR2_X2 \AES_ENC/us00/U293  ( .A1(\AES_ENC/us00/n289 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n288 ) );
NOR2_X2 \AES_ENC/us00/U292  ( .A1(\AES_ENC/us00/n205 ), .A2(\AES_ENC/us00/n270 ), .ZN(\AES_ENC/us00/n416 ) );
NOR2_X2 \AES_ENC/us00/U291  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n584 ), .ZN(\AES_ENC/us00/n358 ) );
NOR2_X2 \AES_ENC/us00/U290  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n602 ), .ZN(\AES_ENC/us00/n359 ) );
NOR2_X2 \AES_ENC/us00/U284  ( .A1(\AES_ENC/us00/n358 ), .A2(\AES_ENC/us00/n359 ), .ZN(\AES_ENC/us00/n351 ) );
NOR2_X2 \AES_ENC/us00/U283  ( .A1(\AES_ENC/us00/n173 ), .A2(\AES_ENC/us00/n136 ), .ZN(\AES_ENC/us00/n456 ) );
NOR2_X2 \AES_ENC/us00/U282  ( .A1(\AES_ENC/us00/n456 ), .A2(\AES_ENC/us00/n616 ), .ZN(\AES_ENC/us00/n454 ) );
NOR2_X2 \AES_ENC/us00/U281  ( .A1(\AES_ENC/us00/n95 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n94 ) );
NOR2_X2 \AES_ENC/us00/U280  ( .A1(\AES_ENC/us00/n73 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n202 ) );
NOR2_X2 \AES_ENC/us00/U279  ( .A1(\AES_ENC/us00/n202 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n201 ) );
NOR2_X2 \AES_ENC/us00/U273  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n620 ), .ZN(\AES_ENC/us00/n168 ) );
NOR2_X2 \AES_ENC/us00/U272  ( .A1(\AES_ENC/us00/n573 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n167 ) );
NOR2_X2 \AES_ENC/us00/U271  ( .A1(\AES_ENC/us00/n167 ), .A2(\AES_ENC/us00/n168 ), .ZN(\AES_ENC/us00/n166 ) );
NOR2_X2 \AES_ENC/us00/U270  ( .A1(\AES_ENC/us00/n165 ), .A2(\AES_ENC/us00/n166 ), .ZN(\AES_ENC/us00/n160 ) );
NOR4_X2 \AES_ENC/us00/U269  ( .A1(\AES_ENC/us00/n439 ), .A2(\AES_ENC/us00/n440 ), .A3(\AES_ENC/us00/n441 ), .A4(\AES_ENC/us00/n442 ), .ZN(\AES_ENC/us00/n438 ) );
NOR2_X2 \AES_ENC/us00/U268  ( .A1(\AES_ENC/us00/n444 ), .A2(\AES_ENC/us00/n445 ), .ZN(\AES_ENC/us00/n437 ) );
NOR2_X2 \AES_ENC/us00/U267  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n123 ), .ZN(\AES_ENC/us00/n527 ) );
NOR2_X2 \AES_ENC/us00/U263  ( .A1(\AES_ENC/us00/n138 ), .A2(\AES_ENC/us00/n205 ), .ZN(\AES_ENC/us00/n204 ) );
NOR2_X2 \AES_ENC/us00/U262  ( .A1(\AES_ENC/us00/n204 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n200 ) );
NOR2_X2 \AES_ENC/us00/U258  ( .A1(\AES_ENC/us00/n607 ), .A2(\AES_ENC/us00/n590 ), .ZN(\AES_ENC/us00/n187 ) );
NOR2_X2 \AES_ENC/us00/U255  ( .A1(\AES_ENC/us00/n357 ), .A2(\AES_ENC/us00/n582 ), .ZN(\AES_ENC/us00/n503 ) );
NOR2_X2 \AES_ENC/us00/U254  ( .A1(\AES_ENC/us00/n606 ), .A2(\AES_ENC/us00/n290 ), .ZN(\AES_ENC/us00/n455 ) );
NOR2_X2 \AES_ENC/us00/U253  ( .A1(\AES_ENC/us00/n140 ), .A2(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n433 ) );
NOR2_X2 \AES_ENC/us00/U252  ( .A1(\AES_ENC/us00/n433 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n427 ) );
NOR2_X2 \AES_ENC/us00/U251  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n577 ), .ZN(\AES_ENC/us00/n188 ) );
NOR2_X2 \AES_ENC/us00/U250  ( .A1(\AES_ENC/us00/n609 ), .A2(\AES_ENC/us00/n580 ), .ZN(\AES_ENC/us00/n70 ) );
NOR2_X2 \AES_ENC/us00/U243  ( .A1(\AES_ENC/us00/n609 ), .A2(\AES_ENC/us00/n590 ), .ZN(\AES_ENC/us00/n486 ) );
INV_X4 \AES_ENC/us00/U242  ( .A(\AES_ENC/us00/n165 ), .ZN(\AES_ENC/us00/n582 ) );
NOR2_X2 \AES_ENC/us00/U241  ( .A1(\AES_ENC/us00/n616 ), .A2(\AES_ENC/us00/n597 ), .ZN(\AES_ENC/us00/n313 ) );
NOR2_X2 \AES_ENC/us00/U240  ( .A1(\AES_ENC/us00/n593 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n68 ) );
NOR2_X2 \AES_ENC/us00/U239  ( .A1(\AES_ENC/us00/n205 ), .A2(\AES_ENC/us00/n267 ), .ZN(\AES_ENC/us00/n304 ) );
NOR2_X2 \AES_ENC/us00/U238  ( .A1(\AES_ENC/us00/n304 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n303 ) );
NOR2_X2 \AES_ENC/us00/U237  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n602 ), .ZN(\AES_ENC/us00/n246 ) );
NOR2_X2 \AES_ENC/us00/U236  ( .A1(\AES_ENC/us00/n115 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n112 ) );
NOR2_X2 \AES_ENC/us00/U235  ( .A1(\AES_ENC/us00/n286 ), .A2(\AES_ENC/us00/n138 ), .ZN(\AES_ENC/us00/n255 ) );
NOR2_X2 \AES_ENC/us00/U234  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n117 ), .ZN(\AES_ENC/us00/n355 ) );
NOR2_X2 \AES_ENC/us00/U229  ( .A1(\AES_ENC/us00/n623 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n566 ) );
NOR2_X2 \AES_ENC/us00/U228  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n602 ), .ZN(\AES_ENC/us00/n390 ) );
NOR2_X2 \AES_ENC/us00/U227  ( .A1(\AES_ENC/us00/n623 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n248 ) );
NOR2_X2 \AES_ENC/us00/U226  ( .A1(\AES_ENC/us00/n606 ), .A2(\AES_ENC/us00/n589 ), .ZN(\AES_ENC/us00/n198 ) );
NOR2_X2 \AES_ENC/us00/U225  ( .A1(\AES_ENC/us00/n72 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n71 ) );
NOR2_X2 \AES_ENC/us00/U223  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n172 ), .ZN(\AES_ENC/us00/n440 ) );
NOR2_X2 \AES_ENC/us00/U222  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n602 ), .ZN(\AES_ENC/us00/n326 ) );
NOR2_X2 \AES_ENC/us00/U221  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n569 ), .ZN(\AES_ENC/us00/n249 ) );
NOR2_X2 \AES_ENC/us00/U217  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n117 ), .ZN(\AES_ENC/us00/n110 ) );
NOR2_X2 \AES_ENC/us00/U213  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n341 ), .ZN(\AES_ENC/us00/n487 ) );
NOR2_X2 \AES_ENC/us00/U212  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n589 ), .ZN(\AES_ENC/us00/n328 ) );
NOR2_X2 \AES_ENC/us00/U211  ( .A1(\AES_ENC/us00/n73 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n69 ) );
NOR2_X2 \AES_ENC/us00/U210  ( .A1(\AES_ENC/us00/n73 ), .A2(\AES_ENC/us00/n357 ), .ZN(\AES_ENC/us00/n354 ) );
NOR2_X2 \AES_ENC/us00/U209  ( .A1(\AES_ENC/us00/n73 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n500 ) );
NOR2_X2 \AES_ENC/us00/U208  ( .A1(\AES_ENC/us00/n120 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n118 ) );
NOR2_X2 \AES_ENC/us00/U207  ( .A1(\AES_ENC/us00/n120 ), .A2(\AES_ENC/us00/n620 ), .ZN(\AES_ENC/us00/n415 ) );
NOR3_X2 \AES_ENC/us00/U201  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n138 ), .A3(\AES_ENC/us00/n205 ), .ZN(\AES_ENC/us00/n216 ) );
NOR3_X2 \AES_ENC/us00/U200  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n136 ), .A3(\AES_ENC/us00/n135 ), .ZN(\AES_ENC/us00/n342 ) );
NOR2_X2 \AES_ENC/us00/U199  ( .A1(\AES_ENC/us00/n199 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n327 ) );
NOR2_X2 \AES_ENC/us00/U198  ( .A1(\AES_ENC/us00/n138 ), .A2(\AES_ENC/us00/n120 ), .ZN(\AES_ENC/us00/n137 ) );
NOR3_X2 \AES_ENC/us00/U197  ( .A1(\AES_ENC/us00/n607 ), .A2(\AES_ENC/us00/n73 ), .A3(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n217 ) );
NOR2_X2 \AES_ENC/us00/U196  ( .A1(\AES_ENC/us00/n199 ), .A2(\AES_ENC/us00/n285 ), .ZN(\AES_ENC/us00/n77 ) );
NOR2_X2 \AES_ENC/us00/U195  ( .A1(\AES_ENC/us00/n120 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n442 ) );
NOR2_X2 \AES_ENC/us00/U194  ( .A1(\AES_ENC/us00/n270 ), .A2(\AES_ENC/us00/n90 ), .ZN(\AES_ENC/us00/n218 ) );
NOR2_X2 \AES_ENC/us00/U187  ( .A1(\AES_ENC/us00/n357 ), .A2(\AES_ENC/us00/n372 ), .ZN(\AES_ENC/us00/n102 ) );
NOR2_X2 \AES_ENC/us00/U186  ( .A1(\AES_ENC/us00/n573 ), .A2(\AES_ENC/us00/n120 ), .ZN(\AES_ENC/us00/n512 ) );
NOR2_X2 \AES_ENC/us00/U185  ( .A1(\AES_ENC/us00/n370 ), .A2(\AES_ENC/us00/n135 ), .ZN(\AES_ENC/us00/n289 ) );
NOR3_X2 \AES_ENC/us00/U184  ( .A1(\AES_ENC/us00/n625 ), .A2(\AES_ENC/us00/n78 ), .A3(\AES_ENC/us00/n585 ), .ZN(\AES_ENC/us00/n365 ) );
NOR3_X2 \AES_ENC/us00/U183  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n138 ), .A3(\AES_ENC/us00/n205 ), .ZN(\AES_ENC/us00/n300 ) );
NOR3_X2 \AES_ENC/us00/U182  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n573 ), .A3(\AES_ENC/us00/n182 ), .ZN(\AES_ENC/us00/n526 ) );
NOR3_X2 \AES_ENC/us00/U181  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n103 ), .A3(\AES_ENC/us00/n173 ), .ZN(\AES_ENC/us00/n353 ) );
NOR2_X2 \AES_ENC/us00/U180  ( .A1(\AES_ENC/us00/n165 ), .A2(\AES_ENC/us00/n99 ), .ZN(\AES_ENC/us00/n461 ) );
NOR2_X2 \AES_ENC/us00/U174  ( .A1(\AES_ENC/us00/n93 ), .A2(\AES_ENC/us00/n342 ), .ZN(\AES_ENC/us00/n336 ) );
NOR4_X2 \AES_ENC/us00/U173  ( .A1(\AES_ENC/us00/n68 ), .A2(\AES_ENC/us00/n69 ), .A3(\AES_ENC/us00/n70 ), .A4(\AES_ENC/us00/n71 ),.ZN(\AES_ENC/us00/n67 ) );
NOR4_X2 \AES_ENC/us00/U172  ( .A1(\AES_ENC/us00/n110 ), .A2(\AES_ENC/us00/n111 ), .A3(\AES_ENC/us00/n112 ), .A4(\AES_ENC/us00/n113 ), .ZN(\AES_ENC/us00/n109 ) );
NOR2_X2 \AES_ENC/us00/U171  ( .A1(\AES_ENC/us00/n118 ), .A2(\AES_ENC/us00/n119 ), .ZN(\AES_ENC/us00/n108 ) );
NAND3_X2 \AES_ENC/us00/U170  ( .A1(\AES_ENC/us00/n569 ), .A2(\AES_ENC/us00/n582 ), .A3(\AES_ENC/us00/n515 ), .ZN(\AES_ENC/us00/n505 ) );
NOR2_X2 \AES_ENC/us00/U169  ( .A1(\AES_ENC/us00/n513 ), .A2(\AES_ENC/us00/n514 ), .ZN(\AES_ENC/us00/n506 ) );
NOR3_X2 \AES_ENC/us00/U168  ( .A1(\AES_ENC/us00/n501 ), .A2(\AES_ENC/us00/n502 ), .A3(\AES_ENC/us00/n503 ), .ZN(\AES_ENC/us00/n496 ) );
NOR4_X2 \AES_ENC/us00/U162  ( .A1(\AES_ENC/us00/n212 ), .A2(\AES_ENC/us00/n498 ), .A3(\AES_ENC/us00/n499 ), .A4(\AES_ENC/us00/n500 ), .ZN(\AES_ENC/us00/n497 ) );
NOR4_X2 \AES_ENC/us00/U161  ( .A1(\AES_ENC/us00/n300 ), .A2(\AES_ENC/us00/n301 ), .A3(\AES_ENC/us00/n302 ), .A4(\AES_ENC/us00/n303 ), .ZN(\AES_ENC/us00/n299 ) );
NOR2_X2 \AES_ENC/us00/U160  ( .A1(\AES_ENC/us00/n330 ), .A2(\AES_ENC/us00/n331 ), .ZN(\AES_ENC/us00/n324 ) );
NOR4_X2 \AES_ENC/us00/U159  ( .A1(\AES_ENC/us00/n326 ), .A2(\AES_ENC/us00/n327 ), .A3(\AES_ENC/us00/n328 ), .A4(\AES_ENC/us00/n329 ), .ZN(\AES_ENC/us00/n325 ) );
NOR2_X2 \AES_ENC/us00/U158  ( .A1(\AES_ENC/us00/n250 ), .A2(\AES_ENC/us00/n251 ), .ZN(\AES_ENC/us00/n244 ) );
NOR4_X2 \AES_ENC/us00/U157  ( .A1(\AES_ENC/us00/n246 ), .A2(\AES_ENC/us00/n247 ), .A3(\AES_ENC/us00/n248 ), .A4(\AES_ENC/us00/n249 ), .ZN(\AES_ENC/us00/n245 ) );
NOR4_X2 \AES_ENC/us00/U156  ( .A1(\AES_ENC/us00/n212 ), .A2(\AES_ENC/us00/n213 ), .A3(\AES_ENC/us00/n214 ), .A4(\AES_ENC/us00/n215 ), .ZN(\AES_ENC/us00/n211 ) );
NOR2_X2 \AES_ENC/us00/U155  ( .A1(\AES_ENC/us00/n216 ), .A2(\AES_ENC/us00/n217 ), .ZN(\AES_ENC/us00/n210 ) );
NOR3_X2 \AES_ENC/us00/U154  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n140 ), .A3(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n234 ) );
NOR3_X2 \AES_ENC/us00/U153  ( .A1(\AES_ENC/us00/n620 ), .A2(\AES_ENC/us00/n120 ), .A3(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n525 ) );
NOR2_X2 \AES_ENC/us00/U152  ( .A1(\AES_ENC/us00/n137 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n132 ) );
NOR2_X2 \AES_ENC/us00/U143  ( .A1(\AES_ENC/us00/n139 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n131 ) );
NOR2_X2 \AES_ENC/us00/U142  ( .A1(\AES_ENC/us00/n134 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n133 ) );
NOR4_X2 \AES_ENC/us00/U141  ( .A1(\AES_ENC/us00/n130 ), .A2(\AES_ENC/us00/n131 ), .A3(\AES_ENC/us00/n132 ), .A4(\AES_ENC/us00/n133 ), .ZN(\AES_ENC/us00/n129 ) );
NOR2_X2 \AES_ENC/us00/U140  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n595 ), .ZN(\AES_ENC/us00/n338 ) );
NOR2_X2 \AES_ENC/us00/U132  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n341 ), .ZN(\AES_ENC/us00/n339 ) );
NOR2_X2 \AES_ENC/us00/U131  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n587 ), .ZN(\AES_ENC/us00/n340 ) );
NOR4_X2 \AES_ENC/us00/U130  ( .A1(\AES_ENC/us00/n338 ), .A2(\AES_ENC/us00/n339 ), .A3(\AES_ENC/us00/n340 ), .A4(\AES_ENC/us00/n238 ), .ZN(\AES_ENC/us00/n337 ) );
NOR3_X2 \AES_ENC/us00/U129  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n73 ), .A3(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n278 ) );
NOR3_X2 \AES_ENC/us00/U128  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n573 ), .A3(\AES_ENC/us00/n182 ), .ZN(\AES_ENC/us00/n279 ) );
NOR2_X2 \AES_ENC/us00/U127  ( .A1(\AES_ENC/us00/n282 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n281 ) );
NOR4_X2 \AES_ENC/us00/U126  ( .A1(\AES_ENC/us00/n278 ), .A2(\AES_ENC/us00/n279 ), .A3(\AES_ENC/us00/n280 ), .A4(\AES_ENC/us00/n281 ), .ZN(\AES_ENC/us00/n277 ) );
NOR2_X2 \AES_ENC/us00/U121  ( .A1(\AES_ENC/us00/n461 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n509 ) );
NOR2_X2 \AES_ENC/us00/U120  ( .A1(\AES_ENC/us00/n512 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n508 ) );
NOR2_X2 \AES_ENC/us00/U119  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n600 ), .ZN(\AES_ENC/us00/n510 ) );
NOR4_X2 \AES_ENC/us00/U118  ( .A1(\AES_ENC/us00/n508 ), .A2(\AES_ENC/us00/n509 ), .A3(\AES_ENC/us00/n510 ), .A4(\AES_ENC/us00/n511 ), .ZN(\AES_ENC/us00/n507 ) );
NOR2_X2 \AES_ENC/us00/U117  ( .A1(\AES_ENC/us00/n616 ), .A2(\AES_ENC/us00/n580 ), .ZN(\AES_ENC/us00/n425 ) );
NOR2_X2 \AES_ENC/us00/U116  ( .A1(\AES_ENC/us00/n90 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n424 ) );
NOR2_X2 \AES_ENC/us00/U115  ( .A1(\AES_ENC/us00/n610 ), .A2(\AES_ENC/us00/n599 ), .ZN(\AES_ENC/us00/n423 ) );
NOR4_X2 \AES_ENC/us00/U106  ( .A1(\AES_ENC/us00/n423 ), .A2(\AES_ENC/us00/n424 ), .A3(\AES_ENC/us00/n425 ), .A4(\AES_ENC/us00/n426 ), .ZN(\AES_ENC/us00/n422 ) );
NOR2_X2 \AES_ENC/us00/U105  ( .A1(\AES_ENC/us00/n416 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n412 ) );
NOR2_X2 \AES_ENC/us00/U104  ( .A1(\AES_ENC/us00/n76 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n414 ) );
NOR2_X2 \AES_ENC/us00/U103  ( .A1(\AES_ENC/us00/n415 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n413 ) );
NOR4_X2 \AES_ENC/us00/U102  ( .A1(\AES_ENC/us00/n316 ), .A2(\AES_ENC/us00/n412 ), .A3(\AES_ENC/us00/n413 ), .A4(\AES_ENC/us00/n414 ), .ZN(\AES_ENC/us00/n411 ) );
NOR2_X2 \AES_ENC/us00/U101  ( .A1(\AES_ENC/us00/n583 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n382 ) );
NOR2_X2 \AES_ENC/us00/U100  ( .A1(\AES_ENC/us00/n289 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n383 ) );
NOR3_X2 \AES_ENC/us00/U95  ( .A1(\AES_ENC/us00/n606 ), .A2(\AES_ENC/us00/n136 ), .A3(\AES_ENC/us00/n135 ), .ZN(\AES_ENC/us00/n381 ) );
NOR4_X2 \AES_ENC/us00/U94  ( .A1(\AES_ENC/us00/n381 ), .A2(\AES_ENC/us00/n382 ), .A3(\AES_ENC/us00/n383 ), .A4(\AES_ENC/us00/n384 ), .ZN(\AES_ENC/us00/n380 ) );
NOR2_X2 \AES_ENC/us00/U93  ( .A1(\AES_ENC/us00/n617 ), .A2(\AES_ENC/us00/n569 ), .ZN(\AES_ENC/us00/n475 ) );
NOR2_X2 \AES_ENC/us00/U92  ( .A1(\AES_ENC/us00/n163 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n473 ) );
NOR2_X2 \AES_ENC/us00/U91  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n97 ), .ZN(\AES_ENC/us00/n474 ) );
NOR4_X2 \AES_ENC/us00/U90  ( .A1(\AES_ENC/us00/n472 ), .A2(\AES_ENC/us00/n473 ), .A3(\AES_ENC/us00/n474 ), .A4(\AES_ENC/us00/n475 ), .ZN(\AES_ENC/us00/n471 ) );
NOR2_X2 \AES_ENC/us00/U89  ( .A1(\AES_ENC/us00/n285 ), .A2(\AES_ENC/us00/n205 ), .ZN(\AES_ENC/us00/n186 ) );
NOR2_X2 \AES_ENC/us00/U88  ( .A1(\AES_ENC/us00/n182 ), .A2(\AES_ENC/us00/n573 ), .ZN(\AES_ENC/us00/n181 ) );
NOR2_X2 \AES_ENC/us00/U87  ( .A1(\AES_ENC/us00/n181 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n180 ) );
NOR4_X2 \AES_ENC/us00/U86  ( .A1(\AES_ENC/us00/n179 ), .A2(\AES_ENC/us00/n180 ), .A3(\AES_ENC/us00/n74 ), .A4(\AES_ENC/us00/n148 ), .ZN(\AES_ENC/us00/n178 ) );
NOR2_X2 \AES_ENC/us00/U81  ( .A1(\AES_ENC/us00/n199 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n197 ) );
NOR2_X2 \AES_ENC/us00/U80  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n577 ), .ZN(\AES_ENC/us00/n195 ) );
NOR2_X2 \AES_ENC/us00/U79  ( .A1(\AES_ENC/us00/n616 ), .A2(\AES_ENC/us00/n97 ), .ZN(\AES_ENC/us00/n196 ) );
NOR4_X2 \AES_ENC/us00/U78  ( .A1(\AES_ENC/us00/n195 ), .A2(\AES_ENC/us00/n196 ), .A3(\AES_ENC/us00/n197 ), .A4(\AES_ENC/us00/n198 ), .ZN(\AES_ENC/us00/n194 ) );
NOR2_X2 \AES_ENC/us00/U74  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n97 ), .ZN(\AES_ENC/us00/n499 ) );
NOR2_X2 \AES_ENC/us00/U73  ( .A1(\AES_ENC/us00/n620 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n238 ) );
NOR2_X2 \AES_ENC/us00/U72  ( .A1(\AES_ENC/us00/n285 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n212 ) );
NOR2_X2 \AES_ENC/us00/U71  ( .A1(\AES_ENC/us00/n140 ), .A2(\AES_ENC/us00/n90 ), .ZN(\AES_ENC/us00/n163 ) );
INV_X4 \AES_ENC/us00/U65  ( .A(\AES_ENC/us00/n144 ), .ZN(\AES_ENC/us00/n612 ) );
INV_X4 \AES_ENC/us00/U64  ( .A(\AES_ENC/us00/n122 ), .ZN(\AES_ENC/us00/n605 ) );
INV_X4 \AES_ENC/us00/U63  ( .A(\AES_ENC/us00/n121 ), .ZN(\AES_ENC/us00/n604 ) );
NOR2_X2 \AES_ENC/us00/U62  ( .A1(\AES_ENC/us00/n582 ), .A2(\AES_ENC/us00/n613 ), .ZN(\AES_ENC/us00/n316 ) );
NOR3_X2 \AES_ENC/us00/U61  ( .A1(\AES_ENC/us00/n370 ), .A2(\AES_ENC/us00/n72 ), .A3(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n250 ) );
INV_X4 \AES_ENC/us00/U59  ( .A(\AES_ENC/us00/n185 ), .ZN(\AES_ENC/us00/n608 ) );
NOR3_X2 \AES_ENC/us00/U58  ( .A1(\AES_ENC/us00/n573 ), .A2(\AES_ENC/us00/n165 ), .A3(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n74 ) );
INV_X4 \AES_ENC/us00/U57  ( .A(\AES_ENC/us00/n240 ), .ZN(\AES_ENC/us00/n615 ) );
NOR2_X2 \AES_ENC/us00/U50  ( .A1(\AES_ENC/us00/n623 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n182 ) );
NOR2_X2 \AES_ENC/us00/U49  ( .A1(\AES_ENC/us00/n620 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n286 ) );
NOR2_X2 \AES_ENC/us00/U48  ( .A1(\AES_ENC/us00/n569 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n103 ) );
NOR2_X2 \AES_ENC/us00/U47  ( .A1(\AES_ENC/us00/n622 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n205 ) );
NOR2_X2 \AES_ENC/us00/U46  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/us00/n72 ), .ZN(\AES_ENC/us00/n199 ) );
NOR2_X2 \AES_ENC/us00/U45  ( .A1(\AES_ENC/us00/n610 ), .A2(\AES_ENC/us00/n600 ), .ZN(\AES_ENC/us00/n568 ) );
NOR2_X2 \AES_ENC/us00/U44  ( .A1(\AES_ENC/us00/n576 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n330 ) );
NOR2_X2 \AES_ENC/us00/U43  ( .A1(\AES_ENC/us00/n603 ), .A2(\AES_ENC/us00/n610 ), .ZN(\AES_ENC/us00/n189 ) );
NOR2_X2 \AES_ENC/us00/U42  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n76 ), .ZN(\AES_ENC/us00/n75 ) );
NOR2_X2 \AES_ENC/us00/U41  ( .A1(\AES_ENC/us00/n74 ), .A2(\AES_ENC/us00/n75 ), .ZN(\AES_ENC/us00/n66 ) );
NOR2_X2 \AES_ENC/us00/U36  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n594 ), .ZN(\AES_ENC/us00/n567 ) );
NOR2_X2 \AES_ENC/us00/U35  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n290 ), .ZN(\AES_ENC/us00/n287 ) );
NOR2_X2 \AES_ENC/us00/U34  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n597 ), .ZN(\AES_ENC/us00/n538 ) );
NOR2_X2 \AES_ENC/us00/U33  ( .A1(\AES_ENC/us00/n77 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n501 ) );
NOR2_X2 \AES_ENC/us00/U32  ( .A1(\AES_ENC/us00/n116 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n111 ) );
NOR2_X2 \AES_ENC/us00/U31  ( .A1(\AES_ENC/us00/n255 ), .A2(\AES_ENC/us00/n608 ), .ZN(\AES_ENC/us00/n472 ) );
NOR2_X2 \AES_ENC/us00/U30  ( .A1(\AES_ENC/us00/n598 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n86 ) );
NOR2_X2 \AES_ENC/us00/U29  ( .A1(\AES_ENC/us00/n576 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n356 ) );
NOR2_X2 \AES_ENC/us00/U24  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n593 ), .ZN(\AES_ENC/us00/n563 ) );
NOR2_X2 \AES_ENC/us00/U23  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n114 ), .ZN(\AES_ENC/us00/n113 ) );
NOR2_X2 \AES_ENC/us00/U21  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n149 ), .ZN(\AES_ENC/us00/n384 ) );
NOR2_X2 \AES_ENC/us00/U20  ( .A1(\AES_ENC/us00/n186 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n235 ) );
NOR2_X2 \AES_ENC/us00/U19  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n601 ), .ZN(\AES_ENC/us00/n213 ) );
NOR2_X2 \AES_ENC/us00/U18  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n594 ), .ZN(\AES_ENC/us00/n439 ) );
NOR2_X2 \AES_ENC/us00/U17  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n590 ), .ZN(\AES_ENC/us00/n498 ) );
NOR2_X2 \AES_ENC/us00/U16  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n619 ), .ZN(\AES_ENC/us00/n488 ) );
NOR2_X2 \AES_ENC/us00/U15  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n582 ), .ZN(\AES_ENC/us00/n426 ) );
NOR2_X2 \AES_ENC/us00/U10  ( .A1(\AES_ENC/us00/n619 ), .A2(\AES_ENC/us00/n604 ), .ZN(\AES_ENC/us00/n393 ) );
NOR2_X2 \AES_ENC/us00/U9  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n315 ), .ZN(\AES_ENC/us00/n485 ) );
NOR2_X2 \AES_ENC/us00/U8  ( .A1(\AES_ENC/us00/n615 ), .A2(\AES_ENC/us00/n582 ), .ZN(\AES_ENC/us00/n329 ) );
NOR2_X2 \AES_ENC/us00/U7  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n599 ), .ZN(\AES_ENC/us00/n392 ) );
NOR2_X2 \AES_ENC/us00/U6  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n620 ), .ZN(\AES_ENC/us00/n148 ) );
OR2_X4 \AES_ENC/us00/U5  ( .A1(\AES_ENC/us00/n624 ), .A2(\AES_ENC/sa00 [1]),.ZN(\AES_ENC/us00/n570 ) );
OR2_X4 \AES_ENC/us00/U4  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/sa00 [4]),.ZN(\AES_ENC/us00/n569 ) );
NAND2_X2 \AES_ENC/us00/U514  ( .A1(\AES_ENC/us00/n72 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n164 ) );
AND2_X2 \AES_ENC/us00/U513  ( .A1(\AES_ENC/us00/n597 ), .A2(\AES_ENC/us00/n164 ), .ZN(\AES_ENC/us00/n145 ) );
NAND2_X2 \AES_ENC/us00/U511  ( .A1(\AES_ENC/us00/n145 ), .A2(\AES_ENC/us00/n402 ), .ZN(\AES_ENC/us00/n559 ) );
AND2_X2 \AES_ENC/us00/U493  ( .A1(\AES_ENC/us00/n417 ), .A2(\AES_ENC/us00/n199 ), .ZN(\AES_ENC/us00/n564 ) );
NAND4_X2 \AES_ENC/us00/U485  ( .A1(\AES_ENC/us00/n559 ), .A2(\AES_ENC/us00/n560 ), .A3(\AES_ENC/us00/n561 ), .A4(\AES_ENC/us00/n562 ), .ZN(\AES_ENC/us00/n558 ) );
NAND2_X2 \AES_ENC/us00/U484  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n558 ), .ZN(\AES_ENC/us00/n517 ) );
NAND2_X2 \AES_ENC/us00/U481  ( .A1(\AES_ENC/us00/n100 ), .A2(\AES_ENC/us00/n591 ), .ZN(\AES_ENC/us00/n548 ) );
NAND2_X2 \AES_ENC/us00/U476  ( .A1(\AES_ENC/us00/n601 ), .A2(\AES_ENC/us00/n590 ), .ZN(\AES_ENC/us00/n434 ) );
NAND2_X2 \AES_ENC/us00/U475  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n434 ), .ZN(\AES_ENC/us00/n549 ) );
NAND4_X2 \AES_ENC/us00/U457  ( .A1(\AES_ENC/us00/n548 ), .A2(\AES_ENC/us00/n549 ), .A3(\AES_ENC/us00/n550 ), .A4(\AES_ENC/us00/n551 ), .ZN(\AES_ENC/us00/n547 ) );
NAND2_X2 \AES_ENC/us00/U456  ( .A1(\AES_ENC/sa00 [0]), .A2(\AES_ENC/us00/n547 ), .ZN(\AES_ENC/us00/n531 ) );
NAND2_X2 \AES_ENC/us00/U454  ( .A1(\AES_ENC/us00/n596 ), .A2(\AES_ENC/us00/n623 ), .ZN(\AES_ENC/us00/n341 ) );
NAND2_X2 \AES_ENC/us00/U453  ( .A1(\AES_ENC/us00/n587 ), .A2(\AES_ENC/us00/n341 ), .ZN(\AES_ENC/us00/n375 ) );
NAND2_X2 \AES_ENC/us00/U452  ( .A1(\AES_ENC/us00/n101 ), .A2(\AES_ENC/us00/n375 ), .ZN(\AES_ENC/us00/n534 ) );
NAND2_X2 \AES_ENC/us00/U451  ( .A1(\AES_ENC/us00/n619 ), .A2(\AES_ENC/us00/n589 ), .ZN(\AES_ENC/us00/n546 ) );
NAND2_X2 \AES_ENC/us00/U450  ( .A1(\AES_ENC/us00/n240 ), .A2(\AES_ENC/us00/n546 ), .ZN(\AES_ENC/us00/n535 ) );
NAND2_X2 \AES_ENC/us00/U449  ( .A1(\AES_ENC/us00/n626 ), .A2(\AES_ENC/us00/n627 ), .ZN(\AES_ENC/us00/n357 ) );
OR2_X2 \AES_ENC/us00/U446  ( .A1(\AES_ENC/us00/n357 ), .A2(\AES_ENC/us00/n264 ), .ZN(\AES_ENC/us00/n540 ) );
NAND2_X2 \AES_ENC/us00/U445  ( .A1(\AES_ENC/us00/n621 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n97 ) );
NAND2_X2 \AES_ENC/us00/U444  ( .A1(\AES_ENC/us00/n164 ), .A2(\AES_ENC/us00/n97 ), .ZN(\AES_ENC/us00/n545 ) );
NAND2_X2 \AES_ENC/us00/U443  ( .A1(\AES_ENC/us00/n79 ), .A2(\AES_ENC/us00/n545 ), .ZN(\AES_ENC/us00/n541 ) );
OR3_X2 \AES_ENC/us00/U440  ( .A1(\AES_ENC/us00/n115 ), .A2(\AES_ENC/sa00 [7]), .A3(\AES_ENC/us00/n626 ), .ZN(\AES_ENC/us00/n542 ) );
NAND2_X2 \AES_ENC/us00/U439  ( .A1(\AES_ENC/us00/n593 ), .A2(\AES_ENC/us00/n601 ), .ZN(\AES_ENC/us00/n544 ) );
NAND4_X2 \AES_ENC/us00/U437  ( .A1(\AES_ENC/us00/n540 ), .A2(\AES_ENC/us00/n541 ), .A3(\AES_ENC/us00/n542 ), .A4(\AES_ENC/us00/n543 ), .ZN(\AES_ENC/us00/n539 ) );
NAND2_X2 \AES_ENC/us00/U436  ( .A1(\AES_ENC/sa00 [2]), .A2(\AES_ENC/us00/n539 ), .ZN(\AES_ENC/us00/n536 ) );
NAND4_X2 \AES_ENC/us00/U432  ( .A1(\AES_ENC/us00/n534 ), .A2(\AES_ENC/us00/n535 ), .A3(\AES_ENC/us00/n536 ), .A4(\AES_ENC/us00/n537 ), .ZN(\AES_ENC/us00/n533 ) );
NAND2_X2 \AES_ENC/us00/U431  ( .A1(\AES_ENC/us00/n533 ), .A2(\AES_ENC/us00/n574 ), .ZN(\AES_ENC/us00/n532 ) );
NAND2_X2 \AES_ENC/us00/U430  ( .A1(\AES_ENC/us00/n531 ), .A2(\AES_ENC/us00/n532 ), .ZN(\AES_ENC/us00/n530 ) );
NAND2_X2 \AES_ENC/us00/U429  ( .A1(\AES_ENC/sa00 [6]), .A2(\AES_ENC/us00/n530 ), .ZN(\AES_ENC/us00/n518 ) );
NAND2_X2 \AES_ENC/us00/U426  ( .A1(\AES_ENC/us00/n461 ), .A2(\AES_ENC/us00/n101 ), .ZN(\AES_ENC/us00/n521 ) );
NAND2_X2 \AES_ENC/us00/U425  ( .A1(\AES_ENC/us00/n588 ), .A2(\AES_ENC/us00/n597 ), .ZN(\AES_ENC/us00/n149 ) );
OR2_X2 \AES_ENC/us00/U424  ( .A1(\AES_ENC/us00/n149 ), .A2(\AES_ENC/us00/n605 ), .ZN(\AES_ENC/us00/n522 ) );
NAND2_X2 \AES_ENC/us00/U423  ( .A1(\AES_ENC/sa00 [1]), .A2(\AES_ENC/us00/n620 ), .ZN(\AES_ENC/us00/n529 ) );
NAND2_X2 \AES_ENC/us00/U422  ( .A1(\AES_ENC/us00/n619 ), .A2(\AES_ENC/us00/n529 ), .ZN(\AES_ENC/us00/n123 ) );
NAND4_X2 \AES_ENC/us00/U412  ( .A1(\AES_ENC/us00/n521 ), .A2(\AES_ENC/us00/n522 ), .A3(\AES_ENC/us00/n523 ), .A4(\AES_ENC/us00/n524 ), .ZN(\AES_ENC/us00/n520 ) );
NAND2_X2 \AES_ENC/us00/U411  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n520 ), .ZN(\AES_ENC/us00/n519 ) );
NAND2_X2 \AES_ENC/us00/U408  ( .A1(\AES_ENC/us00/n396 ), .A2(\AES_ENC/us00/n173 ), .ZN(\AES_ENC/us00/n516 ) );
NAND2_X2 \AES_ENC/us00/U407  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n516 ), .ZN(\AES_ENC/us00/n515 ) );
AND2_X2 \AES_ENC/us00/U402  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n512 ), .ZN(\AES_ENC/us00/n514 ) );
NAND4_X2 \AES_ENC/us00/U395  ( .A1(\AES_ENC/us00/n505 ), .A2(\AES_ENC/us00/n581 ), .A3(\AES_ENC/us00/n506 ), .A4(\AES_ENC/us00/n507 ), .ZN(\AES_ENC/us00/n504 ) );
NAND2_X2 \AES_ENC/us00/U394  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n504 ), .ZN(\AES_ENC/us00/n463 ) );
NAND2_X2 \AES_ENC/us00/U392  ( .A1(\AES_ENC/us00/n218 ), .A2(\AES_ENC/us00/n144 ), .ZN(\AES_ENC/us00/n494 ) );
NAND2_X2 \AES_ENC/us00/U391  ( .A1(\AES_ENC/us00/n101 ), .A2(\AES_ENC/us00/n149 ), .ZN(\AES_ENC/us00/n495 ) );
NAND4_X2 \AES_ENC/us00/U381  ( .A1(\AES_ENC/us00/n494 ), .A2(\AES_ENC/us00/n495 ), .A3(\AES_ENC/us00/n496 ), .A4(\AES_ENC/us00/n497 ), .ZN(\AES_ENC/us00/n493 ) );
NAND2_X2 \AES_ENC/us00/U380  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n493 ), .ZN(\AES_ENC/us00/n464 ) );
AND2_X2 \AES_ENC/us00/U379  ( .A1(\AES_ENC/sa00 [0]), .A2(\AES_ENC/sa00 [6]),.ZN(\AES_ENC/us00/n80 ) );
NAND2_X2 \AES_ENC/us00/U378  ( .A1(\AES_ENC/us00/n601 ), .A2(\AES_ENC/us00/n164 ), .ZN(\AES_ENC/us00/n315 ) );
NAND2_X2 \AES_ENC/us00/U377  ( .A1(\AES_ENC/us00/n101 ), .A2(\AES_ENC/us00/n315 ), .ZN(\AES_ENC/us00/n481 ) );
NAND2_X2 \AES_ENC/us00/U376  ( .A1(\AES_ENC/us00/n185 ), .A2(\AES_ENC/us00/n600 ), .ZN(\AES_ENC/us00/n482 ) );
NAND2_X2 \AES_ENC/us00/U375  ( .A1(\AES_ENC/us00/n341 ), .A2(\AES_ENC/us00/n588 ), .ZN(\AES_ENC/us00/n76 ) );
XNOR2_X2 \AES_ENC/us00/U371  ( .A(\AES_ENC/us00/n611 ), .B(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n372 ) );
NAND4_X2 \AES_ENC/us00/U362  ( .A1(\AES_ENC/us00/n481 ), .A2(\AES_ENC/us00/n482 ), .A3(\AES_ENC/us00/n483 ), .A4(\AES_ENC/us00/n484 ), .ZN(\AES_ENC/us00/n480 ) );
NAND2_X2 \AES_ENC/us00/U361  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n480 ), .ZN(\AES_ENC/us00/n465 ) );
AND2_X2 \AES_ENC/us00/U360  ( .A1(\AES_ENC/sa00 [6]), .A2(\AES_ENC/us00/n574 ), .ZN(\AES_ENC/us00/n62 ) );
NAND2_X2 \AES_ENC/us00/U359  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n479 ) );
NAND2_X2 \AES_ENC/us00/U358  ( .A1(\AES_ENC/us00/n165 ), .A2(\AES_ENC/us00/n479 ), .ZN(\AES_ENC/us00/n468 ) );
NAND2_X2 \AES_ENC/us00/U357  ( .A1(\AES_ENC/sa00 [1]), .A2(\AES_ENC/us00/n624 ), .ZN(\AES_ENC/us00/n96 ) );
NAND2_X2 \AES_ENC/us00/U356  ( .A1(\AES_ENC/us00/n603 ), .A2(\AES_ENC/us00/n96 ), .ZN(\AES_ENC/us00/n478 ) );
NAND2_X2 \AES_ENC/us00/U355  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n478 ), .ZN(\AES_ENC/us00/n469 ) );
NAND4_X2 \AES_ENC/us00/U344  ( .A1(\AES_ENC/us00/n468 ), .A2(\AES_ENC/us00/n469 ), .A3(\AES_ENC/us00/n470 ), .A4(\AES_ENC/us00/n471 ), .ZN(\AES_ENC/us00/n467 ) );
NAND2_X2 \AES_ENC/us00/U343  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n467 ), .ZN(\AES_ENC/us00/n466 ) );
NAND4_X2 \AES_ENC/us00/U342  ( .A1(\AES_ENC/us00/n463 ), .A2(\AES_ENC/us00/n464 ), .A3(\AES_ENC/us00/n465 ), .A4(\AES_ENC/us00/n466 ), .ZN(\AES_ENC/sa00_sub[1] ) );
NAND2_X2 \AES_ENC/us00/U341  ( .A1(\AES_ENC/sa00 [7]), .A2(\AES_ENC/us00/n611 ), .ZN(\AES_ENC/us00/n462 ) );
NAND2_X2 \AES_ENC/us00/U340  ( .A1(\AES_ENC/us00/n462 ), .A2(\AES_ENC/us00/n607 ), .ZN(\AES_ENC/us00/n458 ) );
OR4_X2 \AES_ENC/us00/U339  ( .A1(\AES_ENC/us00/n458 ), .A2(\AES_ENC/us00/n626 ), .A3(\AES_ENC/us00/n370 ), .A4(\AES_ENC/us00/n72 ), .ZN(\AES_ENC/us00/n450 ) );
NAND2_X2 \AES_ENC/us00/U337  ( .A1(\AES_ENC/us00/n93 ), .A2(\AES_ENC/us00/n587 ), .ZN(\AES_ENC/us00/n203 ) );
OR2_X2 \AES_ENC/us00/U336  ( .A1(\AES_ENC/us00/n610 ), .A2(\AES_ENC/us00/n461 ), .ZN(\AES_ENC/us00/n459 ) );
NAND2_X2 \AES_ENC/us00/U334  ( .A1(\AES_ENC/us00/n619 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n443 ) );
NAND2_X2 \AES_ENC/us00/U333  ( .A1(\AES_ENC/us00/n582 ), .A2(\AES_ENC/us00/n443 ), .ZN(\AES_ENC/us00/n114 ) );
NAND2_X2 \AES_ENC/us00/U332  ( .A1(\AES_ENC/us00/n146 ), .A2(\AES_ENC/us00/n576 ), .ZN(\AES_ENC/us00/n460 ) );
NAND2_X2 \AES_ENC/us00/U331  ( .A1(\AES_ENC/us00/n459 ), .A2(\AES_ENC/us00/n460 ), .ZN(\AES_ENC/us00/n457 ) );
NAND2_X2 \AES_ENC/us00/U330  ( .A1(\AES_ENC/us00/n457 ), .A2(\AES_ENC/us00/n458 ), .ZN(\AES_ENC/us00/n451 ) );
NAND2_X2 \AES_ENC/us00/U326  ( .A1(\AES_ENC/us00/n97 ), .A2(\AES_ENC/us00/n590 ), .ZN(\AES_ENC/us00/n290 ) );
NAND4_X2 \AES_ENC/us00/U323  ( .A1(\AES_ENC/us00/n450 ), .A2(\AES_ENC/us00/n203 ), .A3(\AES_ENC/us00/n451 ), .A4(\AES_ENC/us00/n452 ), .ZN(\AES_ENC/us00/n449 ) );
NAND2_X2 \AES_ENC/us00/U322  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n449 ), .ZN(\AES_ENC/us00/n403 ) );
NAND2_X2 \AES_ENC/us00/U321  ( .A1(\AES_ENC/us00/n584 ), .A2(\AES_ENC/us00/n341 ), .ZN(\AES_ENC/us00/n448 ) );
NAND2_X2 \AES_ENC/us00/U320  ( .A1(\AES_ENC/us00/n240 ), .A2(\AES_ENC/us00/n448 ), .ZN(\AES_ENC/us00/n436 ) );
NAND2_X2 \AES_ENC/us00/U313  ( .A1(\AES_ENC/us00/n590 ), .A2(\AES_ENC/us00/n443 ), .ZN(\AES_ENC/us00/n172 ) );
NAND4_X2 \AES_ENC/us00/U308  ( .A1(\AES_ENC/us00/n436 ), .A2(\AES_ENC/us00/n203 ), .A3(\AES_ENC/us00/n437 ), .A4(\AES_ENC/us00/n438 ), .ZN(\AES_ENC/us00/n435 ) );
NAND2_X2 \AES_ENC/us00/U307  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n435 ), .ZN(\AES_ENC/us00/n404 ) );
NAND2_X2 \AES_ENC/us00/U306  ( .A1(\AES_ENC/us00/n584 ), .A2(\AES_ENC/us00/n603 ), .ZN(\AES_ENC/us00/n206 ) );
NAND2_X2 \AES_ENC/us00/U305  ( .A1(\AES_ENC/us00/n144 ), .A2(\AES_ENC/us00/n206 ), .ZN(\AES_ENC/us00/n419 ) );
NAND2_X2 \AES_ENC/us00/U304  ( .A1(\AES_ENC/us00/n101 ), .A2(\AES_ENC/us00/n434 ), .ZN(\AES_ENC/us00/n420 ) );
XNOR2_X2 \AES_ENC/us00/U301  ( .A(\AES_ENC/sa00 [7]), .B(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n237 ) );
NAND4_X2 \AES_ENC/us00/U289  ( .A1(\AES_ENC/us00/n419 ), .A2(\AES_ENC/us00/n420 ), .A3(\AES_ENC/us00/n421 ), .A4(\AES_ENC/us00/n422 ), .ZN(\AES_ENC/us00/n418 ) );
NAND2_X2 \AES_ENC/us00/U288  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n418 ), .ZN(\AES_ENC/us00/n405 ) );
NAND2_X2 \AES_ENC/us00/U287  ( .A1(\AES_ENC/us00/n138 ), .A2(\AES_ENC/us00/n144 ), .ZN(\AES_ENC/us00/n408 ) );
NAND2_X2 \AES_ENC/us00/U286  ( .A1(\AES_ENC/us00/n103 ), .A2(\AES_ENC/us00/n417 ), .ZN(\AES_ENC/us00/n409 ) );
NAND2_X2 \AES_ENC/us00/U285  ( .A1(\AES_ENC/us00/n240 ), .A2(\AES_ENC/sa00 [1]), .ZN(\AES_ENC/us00/n410 ) );
NAND4_X2 \AES_ENC/us00/U278  ( .A1(\AES_ENC/us00/n408 ), .A2(\AES_ENC/us00/n409 ), .A3(\AES_ENC/us00/n410 ), .A4(\AES_ENC/us00/n411 ), .ZN(\AES_ENC/us00/n407 ) );
NAND2_X2 \AES_ENC/us00/U277  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n407 ), .ZN(\AES_ENC/us00/n406 ) );
NAND4_X2 \AES_ENC/us00/U276  ( .A1(\AES_ENC/us00/n403 ), .A2(\AES_ENC/us00/n404 ), .A3(\AES_ENC/us00/n405 ), .A4(\AES_ENC/us00/n406 ), .ZN(\AES_ENC/sa00_sub[2] ) );
NAND2_X2 \AES_ENC/us00/U275  ( .A1(\AES_ENC/us00/n135 ), .A2(\AES_ENC/us00/n402 ), .ZN(\AES_ENC/us00/n386 ) );
NAND2_X2 \AES_ENC/us00/U274  ( .A1(\AES_ENC/us00/n145 ), .A2(\AES_ENC/us00/n240 ), .ZN(\AES_ENC/us00/n387 ) );
OR2_X2 \AES_ENC/us00/U266  ( .A1(\AES_ENC/us00/n97 ), .A2(\AES_ENC/us00/n606 ), .ZN(\AES_ENC/us00/n394 ) );
NAND2_X2 \AES_ENC/us00/U265  ( .A1(\AES_ENC/us00/n141 ), .A2(\AES_ENC/us00/n396 ), .ZN(\AES_ENC/us00/n395 ) );
NAND2_X2 \AES_ENC/us00/U264  ( .A1(\AES_ENC/us00/n394 ), .A2(\AES_ENC/us00/n395 ), .ZN(\AES_ENC/us00/n391 ) );
NAND4_X2 \AES_ENC/us00/U261  ( .A1(\AES_ENC/us00/n386 ), .A2(\AES_ENC/us00/n387 ), .A3(\AES_ENC/us00/n388 ), .A4(\AES_ENC/us00/n389 ), .ZN(\AES_ENC/us00/n385 ) );
NAND2_X2 \AES_ENC/us00/U260  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n385 ), .ZN(\AES_ENC/us00/n344 ) );
OR2_X2 \AES_ENC/us00/U259  ( .A1(\AES_ENC/us00/n172 ), .A2(\AES_ENC/us00/n617 ), .ZN(\AES_ENC/us00/n377 ) );
OR2_X2 \AES_ENC/us00/U257  ( .A1(\AES_ENC/us00/n570 ), .A2(\AES_ENC/us00/n266 ), .ZN(\AES_ENC/us00/n378 ) );
NAND2_X2 \AES_ENC/us00/U256  ( .A1(\AES_ENC/us00/n182 ), .A2(\AES_ENC/us00/n100 ), .ZN(\AES_ENC/us00/n379 ) );
NAND4_X2 \AES_ENC/us00/U249  ( .A1(\AES_ENC/us00/n377 ), .A2(\AES_ENC/us00/n378 ), .A3(\AES_ENC/us00/n379 ), .A4(\AES_ENC/us00/n380 ), .ZN(\AES_ENC/us00/n376 ) );
NAND2_X2 \AES_ENC/us00/U248  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n376 ), .ZN(\AES_ENC/us00/n345 ) );
NAND2_X2 \AES_ENC/us00/U247  ( .A1(\AES_ENC/us00/n240 ), .A2(\AES_ENC/us00/n114 ), .ZN(\AES_ENC/us00/n361 ) );
NAND2_X2 \AES_ENC/us00/U246  ( .A1(\AES_ENC/us00/n570 ), .A2(\AES_ENC/us00/n164 ), .ZN(\AES_ENC/us00/n147 ) );
OR2_X2 \AES_ENC/us00/U245  ( .A1(\AES_ENC/us00/n147 ), .A2(\AES_ENC/us00/n612 ), .ZN(\AES_ENC/us00/n362 ) );
NAND2_X2 \AES_ENC/us00/U244  ( .A1(\AES_ENC/us00/n122 ), .A2(\AES_ENC/us00/n589 ), .ZN(\AES_ENC/us00/n363 ) );
NAND4_X2 \AES_ENC/us00/U233  ( .A1(\AES_ENC/us00/n361 ), .A2(\AES_ENC/us00/n362 ), .A3(\AES_ENC/us00/n363 ), .A4(\AES_ENC/us00/n364 ), .ZN(\AES_ENC/us00/n360 ) );
NAND2_X2 \AES_ENC/us00/U232  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n360 ), .ZN(\AES_ENC/us00/n346 ) );
NAND2_X2 \AES_ENC/us00/U231  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n623 ), .ZN(\AES_ENC/us00/n349 ) );
NAND2_X2 \AES_ENC/us00/U230  ( .A1(\AES_ENC/us00/n144 ), .A2(\AES_ENC/us00/n123 ), .ZN(\AES_ENC/us00/n350 ) );
OR2_X2 \AES_ENC/us00/U224  ( .A1(\AES_ENC/us00/n141 ), .A2(\AES_ENC/us00/n285 ), .ZN(\AES_ENC/us00/n117 ) );
NAND4_X2 \AES_ENC/us00/U220  ( .A1(\AES_ENC/us00/n349 ), .A2(\AES_ENC/us00/n350 ), .A3(\AES_ENC/us00/n351 ), .A4(\AES_ENC/us00/n352 ), .ZN(\AES_ENC/us00/n348 ) );
NAND2_X2 \AES_ENC/us00/U219  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n348 ), .ZN(\AES_ENC/us00/n347 ) );
NAND4_X2 \AES_ENC/us00/U218  ( .A1(\AES_ENC/us00/n344 ), .A2(\AES_ENC/us00/n345 ), .A3(\AES_ENC/us00/n346 ), .A4(\AES_ENC/us00/n347 ), .ZN(\AES_ENC/sa00_sub[3] ) );
NAND2_X2 \AES_ENC/us00/U216  ( .A1(\AES_ENC/us00/n186 ), .A2(\AES_ENC/us00/n122 ), .ZN(\AES_ENC/us00/n334 ) );
NAND2_X2 \AES_ENC/us00/U215  ( .A1(\AES_ENC/us00/n603 ), .A2(\AES_ENC/us00/n577 ), .ZN(\AES_ENC/us00/n343 ) );
NAND2_X2 \AES_ENC/us00/U214  ( .A1(\AES_ENC/us00/n144 ), .A2(\AES_ENC/us00/n343 ), .ZN(\AES_ENC/us00/n335 ) );
NAND4_X2 \AES_ENC/us00/U206  ( .A1(\AES_ENC/us00/n334 ), .A2(\AES_ENC/us00/n335 ), .A3(\AES_ENC/us00/n336 ), .A4(\AES_ENC/us00/n337 ), .ZN(\AES_ENC/us00/n333 ) );
NAND2_X2 \AES_ENC/us00/U205  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n333 ), .ZN(\AES_ENC/us00/n291 ) );
NAND2_X2 \AES_ENC/us00/U204  ( .A1(\AES_ENC/us00/n185 ), .A2(\AES_ENC/us00/n206 ), .ZN(\AES_ENC/us00/n322 ) );
NAND2_X2 \AES_ENC/us00/U203  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n610 ), .ZN(\AES_ENC/us00/n332 ) );
NAND2_X2 \AES_ENC/us00/U202  ( .A1(\AES_ENC/us00/n267 ), .A2(\AES_ENC/us00/n332 ), .ZN(\AES_ENC/us00/n323 ) );
NAND4_X2 \AES_ENC/us00/U193  ( .A1(\AES_ENC/us00/n322 ), .A2(\AES_ENC/us00/n323 ), .A3(\AES_ENC/us00/n324 ), .A4(\AES_ENC/us00/n325 ), .ZN(\AES_ENC/us00/n321 ) );
NAND2_X2 \AES_ENC/us00/U192  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n321 ), .ZN(\AES_ENC/us00/n292 ) );
NAND2_X2 \AES_ENC/us00/U191  ( .A1(\AES_ENC/us00/n583 ), .A2(\AES_ENC/us00/n144 ), .ZN(\AES_ENC/us00/n307 ) );
NAND2_X2 \AES_ENC/us00/U190  ( .A1(\AES_ENC/us00/n101 ), .A2(\AES_ENC/us00/n587 ), .ZN(\AES_ENC/us00/n320 ) );
NAND2_X2 \AES_ENC/us00/U189  ( .A1(\AES_ENC/us00/n604 ), .A2(\AES_ENC/us00/n320 ), .ZN(\AES_ENC/us00/n319 ) );
NAND2_X2 \AES_ENC/us00/U188  ( .A1(\AES_ENC/us00/n319 ), .A2(\AES_ENC/us00/n623 ), .ZN(\AES_ENC/us00/n308 ) );
NAND4_X2 \AES_ENC/us00/U179  ( .A1(\AES_ENC/us00/n307 ), .A2(\AES_ENC/us00/n308 ), .A3(\AES_ENC/us00/n309 ), .A4(\AES_ENC/us00/n310 ), .ZN(\AES_ENC/us00/n306 ) );
NAND2_X2 \AES_ENC/us00/U178  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n306 ), .ZN(\AES_ENC/us00/n293 ) );
OR2_X2 \AES_ENC/us00/U177  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n135 ), .ZN(\AES_ENC/us00/n296 ) );
NAND2_X2 \AES_ENC/us00/U176  ( .A1(\AES_ENC/us00/n121 ), .A2(\AES_ENC/us00/n147 ), .ZN(\AES_ENC/us00/n297 ) );
NAND2_X2 \AES_ENC/us00/U175  ( .A1(\AES_ENC/us00/n100 ), .A2(\AES_ENC/us00/n595 ), .ZN(\AES_ENC/us00/n298 ) );
NAND4_X2 \AES_ENC/us00/U167  ( .A1(\AES_ENC/us00/n296 ), .A2(\AES_ENC/us00/n297 ), .A3(\AES_ENC/us00/n298 ), .A4(\AES_ENC/us00/n299 ), .ZN(\AES_ENC/us00/n295 ) );
NAND2_X2 \AES_ENC/us00/U166  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n295 ), .ZN(\AES_ENC/us00/n294 ) );
NAND4_X2 \AES_ENC/us00/U165  ( .A1(\AES_ENC/us00/n291 ), .A2(\AES_ENC/us00/n292 ), .A3(\AES_ENC/us00/n293 ), .A4(\AES_ENC/us00/n294 ), .ZN(\AES_ENC/sa00_sub[4] ) );
NAND2_X2 \AES_ENC/us00/U164  ( .A1(\AES_ENC/us00/n100 ), .A2(\AES_ENC/us00/n599 ), .ZN(\AES_ENC/us00/n274 ) );
NAND2_X2 \AES_ENC/us00/U163  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n206 ), .ZN(\AES_ENC/us00/n275 ) );
NAND4_X2 \AES_ENC/us00/U151  ( .A1(\AES_ENC/us00/n274 ), .A2(\AES_ENC/us00/n275 ), .A3(\AES_ENC/us00/n276 ), .A4(\AES_ENC/us00/n277 ), .ZN(\AES_ENC/us00/n273 ) );
NAND2_X2 \AES_ENC/us00/U150  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n273 ), .ZN(\AES_ENC/us00/n223 ) );
NAND2_X2 \AES_ENC/us00/U149  ( .A1(\AES_ENC/us00/n582 ), .A2(\AES_ENC/us00/n619 ), .ZN(\AES_ENC/us00/n272 ) );
NAND2_X2 \AES_ENC/us00/U148  ( .A1(\AES_ENC/us00/n121 ), .A2(\AES_ENC/us00/n272 ), .ZN(\AES_ENC/us00/n257 ) );
NAND2_X2 \AES_ENC/us00/U147  ( .A1(\AES_ENC/us00/n270 ), .A2(\AES_ENC/us00/n271 ), .ZN(\AES_ENC/us00/n269 ) );
NAND2_X2 \AES_ENC/us00/U146  ( .A1(\AES_ENC/us00/n606 ), .A2(\AES_ENC/us00/n269 ), .ZN(\AES_ENC/us00/n268 ) );
NAND2_X2 \AES_ENC/us00/U145  ( .A1(\AES_ENC/us00/n268 ), .A2(\AES_ENC/us00/n114 ), .ZN(\AES_ENC/us00/n258 ) );
OR2_X2 \AES_ENC/us00/U144  ( .A1(\AES_ENC/us00/n76 ), .A2(\AES_ENC/us00/n615 ), .ZN(\AES_ENC/us00/n259 ) );
NAND4_X2 \AES_ENC/us00/U139  ( .A1(\AES_ENC/us00/n257 ), .A2(\AES_ENC/us00/n258 ), .A3(\AES_ENC/us00/n259 ), .A4(\AES_ENC/us00/n260 ), .ZN(\AES_ENC/us00/n256 ) );
NAND2_X2 \AES_ENC/us00/U138  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n256 ), .ZN(\AES_ENC/us00/n224 ) );
OR2_X2 \AES_ENC/us00/U137  ( .A1(\AES_ENC/us00/n605 ), .A2(\AES_ENC/us00/n255 ), .ZN(\AES_ENC/us00/n242 ) );
NAND2_X2 \AES_ENC/us00/U136  ( .A1(\AES_ENC/us00/n97 ), .A2(\AES_ENC/us00/n577 ), .ZN(\AES_ENC/us00/n254 ) );
NAND2_X2 \AES_ENC/us00/U135  ( .A1(\AES_ENC/us00/n146 ), .A2(\AES_ENC/us00/n254 ), .ZN(\AES_ENC/us00/n253 ) );
NAND2_X2 \AES_ENC/us00/U134  ( .A1(\AES_ENC/us00/n612 ), .A2(\AES_ENC/us00/n253 ), .ZN(\AES_ENC/us00/n252 ) );
NAND2_X2 \AES_ENC/us00/U133  ( .A1(\AES_ENC/us00/n252 ), .A2(\AES_ENC/us00/n580 ), .ZN(\AES_ENC/us00/n243 ) );
NAND4_X2 \AES_ENC/us00/U125  ( .A1(\AES_ENC/us00/n242 ), .A2(\AES_ENC/us00/n243 ), .A3(\AES_ENC/us00/n244 ), .A4(\AES_ENC/us00/n245 ), .ZN(\AES_ENC/us00/n241 ) );
NAND2_X2 \AES_ENC/us00/U124  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n241 ), .ZN(\AES_ENC/us00/n225 ) );
NAND2_X2 \AES_ENC/us00/U123  ( .A1(\AES_ENC/us00/n100 ), .A2(\AES_ENC/us00/n123 ), .ZN(\AES_ENC/us00/n228 ) );
NAND2_X2 \AES_ENC/us00/U122  ( .A1(\AES_ENC/us00/n240 ), .A2(\AES_ENC/us00/n164 ), .ZN(\AES_ENC/us00/n229 ) );
NAND4_X2 \AES_ENC/us00/U114  ( .A1(\AES_ENC/us00/n228 ), .A2(\AES_ENC/us00/n229 ), .A3(\AES_ENC/us00/n230 ), .A4(\AES_ENC/us00/n231 ), .ZN(\AES_ENC/us00/n227 ) );
NAND2_X2 \AES_ENC/us00/U113  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n227 ), .ZN(\AES_ENC/us00/n226 ) );
NAND4_X2 \AES_ENC/us00/U112  ( .A1(\AES_ENC/us00/n223 ), .A2(\AES_ENC/us00/n224 ), .A3(\AES_ENC/us00/n225 ), .A4(\AES_ENC/us00/n226 ), .ZN(\AES_ENC/sa00_sub[5] ) );
NAND2_X2 \AES_ENC/us00/U111  ( .A1(\AES_ENC/us00/n570 ), .A2(\AES_ENC/us00/n96 ), .ZN(\AES_ENC/us00/n222 ) );
NAND2_X2 \AES_ENC/us00/U110  ( .A1(\AES_ENC/us00/n121 ), .A2(\AES_ENC/us00/n222 ), .ZN(\AES_ENC/us00/n208 ) );
NAND2_X2 \AES_ENC/us00/U109  ( .A1(\AES_ENC/us00/n221 ), .A2(\AES_ENC/us00/n117 ), .ZN(\AES_ENC/us00/n220 ) );
NAND2_X2 \AES_ENC/us00/U108  ( .A1(\AES_ENC/us00/n613 ), .A2(\AES_ENC/us00/n220 ), .ZN(\AES_ENC/us00/n219 ) );
NAND2_X2 \AES_ENC/us00/U107  ( .A1(\AES_ENC/us00/n218 ), .A2(\AES_ENC/us00/n219 ), .ZN(\AES_ENC/us00/n209 ) );
NAND4_X2 \AES_ENC/us00/U99  ( .A1(\AES_ENC/us00/n208 ), .A2(\AES_ENC/us00/n209 ), .A3(\AES_ENC/us00/n210 ), .A4(\AES_ENC/us00/n211 ), .ZN(\AES_ENC/us00/n207 ) );
NAND2_X2 \AES_ENC/us00/U98  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n207 ), .ZN(\AES_ENC/us00/n150 ) );
NAND2_X2 \AES_ENC/us00/U97  ( .A1(\AES_ENC/us00/n121 ), .A2(\AES_ENC/us00/n206 ), .ZN(\AES_ENC/us00/n191 ) );
NAND2_X2 \AES_ENC/us00/U96  ( .A1(\AES_ENC/us00/n102 ), .A2(\AES_ENC/us00/n619 ), .ZN(\AES_ENC/us00/n192 ) );
NAND4_X2 \AES_ENC/us00/U85  ( .A1(\AES_ENC/us00/n191 ), .A2(\AES_ENC/us00/n192 ), .A3(\AES_ENC/us00/n193 ), .A4(\AES_ENC/us00/n194 ), .ZN(\AES_ENC/us00/n190 ) );
NAND2_X2 \AES_ENC/us00/U84  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n190 ), .ZN(\AES_ENC/us00/n151 ) );
NAND2_X2 \AES_ENC/us00/U83  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n596 ), .ZN(\AES_ENC/us00/n175 ) );
NAND2_X2 \AES_ENC/us00/U82  ( .A1(\AES_ENC/us00/n144 ), .A2(\AES_ENC/us00/n624 ), .ZN(\AES_ENC/us00/n176 ) );
NAND2_X2 \AES_ENC/us00/U77  ( .A1(\AES_ENC/us00/n135 ), .A2(\AES_ENC/us00/n79 ), .ZN(\AES_ENC/us00/n183 ) );
NAND2_X2 \AES_ENC/us00/U76  ( .A1(\AES_ENC/us00/n185 ), .A2(\AES_ENC/us00/n592 ), .ZN(\AES_ENC/us00/n184 ) );
NAND2_X2 \AES_ENC/us00/U75  ( .A1(\AES_ENC/us00/n183 ), .A2(\AES_ENC/us00/n184 ), .ZN(\AES_ENC/us00/n179 ) );
NAND4_X2 \AES_ENC/us00/U70  ( .A1(\AES_ENC/us00/n175 ), .A2(\AES_ENC/us00/n176 ), .A3(\AES_ENC/us00/n177 ), .A4(\AES_ENC/us00/n178 ), .ZN(\AES_ENC/us00/n174 ) );
NAND2_X2 \AES_ENC/us00/U69  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n174 ), .ZN(\AES_ENC/us00/n152 ) );
NAND2_X2 \AES_ENC/us00/U68  ( .A1(\AES_ENC/us00/n173 ), .A2(\AES_ENC/us00/n101 ), .ZN(\AES_ENC/us00/n155 ) );
NAND2_X2 \AES_ENC/us00/U67  ( .A1(\AES_ENC/us00/n144 ), .A2(\AES_ENC/us00/n172 ), .ZN(\AES_ENC/us00/n156 ) );
NAND2_X2 \AES_ENC/us00/U66  ( .A1(\AES_ENC/us00/n171 ), .A2(\AES_ENC/us00/n123 ), .ZN(\AES_ENC/us00/n157 ) );
AND2_X2 \AES_ENC/us00/U60  ( .A1(\AES_ENC/us00/n164 ), .A2(\AES_ENC/us00/n602 ), .ZN(\AES_ENC/us00/n116 ) );
NAND4_X2 \AES_ENC/us00/U56  ( .A1(\AES_ENC/us00/n155 ), .A2(\AES_ENC/us00/n156 ), .A3(\AES_ENC/us00/n157 ), .A4(\AES_ENC/us00/n158 ), .ZN(\AES_ENC/us00/n154 ) );
NAND2_X2 \AES_ENC/us00/U55  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n154 ), .ZN(\AES_ENC/us00/n153 ) );
NAND4_X2 \AES_ENC/us00/U54  ( .A1(\AES_ENC/us00/n150 ), .A2(\AES_ENC/us00/n151 ), .A3(\AES_ENC/us00/n152 ), .A4(\AES_ENC/us00/n153 ), .ZN(\AES_ENC/sa00_sub[6] ) );
NAND2_X2 \AES_ENC/us00/U53  ( .A1(\AES_ENC/us00/n122 ), .A2(\AES_ENC/us00/n149 ), .ZN(\AES_ENC/us00/n126 ) );
NAND2_X2 \AES_ENC/us00/U52  ( .A1(\AES_ENC/us00/n148 ), .A2(\AES_ENC/us00/n582 ), .ZN(\AES_ENC/us00/n127 ) );
NAND2_X2 \AES_ENC/us00/U51  ( .A1(\AES_ENC/us00/n100 ), .A2(\AES_ENC/us00/n147 ), .ZN(\AES_ENC/us00/n128 ) );
NAND4_X2 \AES_ENC/us00/U40  ( .A1(\AES_ENC/us00/n126 ), .A2(\AES_ENC/us00/n127 ), .A3(\AES_ENC/us00/n128 ), .A4(\AES_ENC/us00/n129 ), .ZN(\AES_ENC/us00/n125 ) );
NAND2_X2 \AES_ENC/us00/U39  ( .A1(\AES_ENC/us00/n124 ), .A2(\AES_ENC/us00/n125 ), .ZN(\AES_ENC/us00/n58 ) );
NAND2_X2 \AES_ENC/us00/U38  ( .A1(\AES_ENC/us00/n122 ), .A2(\AES_ENC/us00/n123 ), .ZN(\AES_ENC/us00/n106 ) );
NAND2_X2 \AES_ENC/us00/U37  ( .A1(\AES_ENC/us00/n121 ), .A2(\AES_ENC/us00/n595 ), .ZN(\AES_ENC/us00/n107 ) );
NAND4_X2 \AES_ENC/us00/U28  ( .A1(\AES_ENC/us00/n106 ), .A2(\AES_ENC/us00/n107 ), .A3(\AES_ENC/us00/n108 ), .A4(\AES_ENC/us00/n109 ), .ZN(\AES_ENC/us00/n105 ) );
NAND2_X2 \AES_ENC/us00/U27  ( .A1(\AES_ENC/us00/n104 ), .A2(\AES_ENC/us00/n105 ), .ZN(\AES_ENC/us00/n59 ) );
NAND2_X2 \AES_ENC/us00/U26  ( .A1(\AES_ENC/us00/n103 ), .A2(\AES_ENC/us00/n101 ), .ZN(\AES_ENC/us00/n82 ) );
NAND2_X2 \AES_ENC/us00/U25  ( .A1(\AES_ENC/us00/n102 ), .A2(\AES_ENC/us00/n73 ), .ZN(\AES_ENC/us00/n83 ) );
AND2_X2 \AES_ENC/us00/U22  ( .A1(\AES_ENC/us00/n96 ), .A2(\AES_ENC/us00/n97 ), .ZN(\AES_ENC/us00/n95 ) );
NAND4_X2 \AES_ENC/us00/U14  ( .A1(\AES_ENC/us00/n82 ), .A2(\AES_ENC/us00/n83 ), .A3(\AES_ENC/us00/n84 ), .A4(\AES_ENC/us00/n85 ),.ZN(\AES_ENC/us00/n81 ) );
NAND2_X2 \AES_ENC/us00/U13  ( .A1(\AES_ENC/us00/n80 ), .A2(\AES_ENC/us00/n81 ), .ZN(\AES_ENC/us00/n60 ) );
NAND2_X2 \AES_ENC/us00/U12  ( .A1(\AES_ENC/us00/n78 ), .A2(\AES_ENC/us00/n79 ), .ZN(\AES_ENC/us00/n64 ) );
OR2_X2 \AES_ENC/us00/U11  ( .A1(\AES_ENC/us00/n608 ), .A2(\AES_ENC/us00/n77 ), .ZN(\AES_ENC/us00/n65 ) );
NAND4_X2 \AES_ENC/us00/U3  ( .A1(\AES_ENC/us00/n64 ), .A2(\AES_ENC/us00/n65 ), .A3(\AES_ENC/us00/n66 ), .A4(\AES_ENC/us00/n67 ), .ZN(\AES_ENC/us00/n63 ) );
NAND2_X2 \AES_ENC/us00/U2  ( .A1(\AES_ENC/us00/n62 ), .A2(\AES_ENC/us00/n63 ), .ZN(\AES_ENC/us00/n61 ) );
NAND4_X2 \AES_ENC/us00/U1  ( .A1(\AES_ENC/us00/n58 ), .A2(\AES_ENC/us00/n59 ), .A3(\AES_ENC/us00/n60 ), .A4(\AES_ENC/us00/n61 ), .ZN(\AES_ENC/sa00_sub[7] ));
INV_X4 \AES_ENC/us01/U575  ( .A(\AES_ENC/sa01 [0]), .ZN(\AES_ENC/us01/n627 ));
INV_X4 \AES_ENC/us01/U574  ( .A(\AES_ENC/us01/n1053 ), .ZN(\AES_ENC/us01/n625 ) );
INV_X4 \AES_ENC/us01/U573  ( .A(\AES_ENC/us01/n1103 ), .ZN(\AES_ENC/us01/n623 ) );
INV_X4 \AES_ENC/us01/U572  ( .A(\AES_ENC/us01/n1056 ), .ZN(\AES_ENC/us01/n622 ) );
INV_X4 \AES_ENC/us01/U571  ( .A(\AES_ENC/us01/n1102 ), .ZN(\AES_ENC/us01/n621 ) );
INV_X4 \AES_ENC/us01/U570  ( .A(\AES_ENC/us01/n1074 ), .ZN(\AES_ENC/us01/n620 ) );
INV_X4 \AES_ENC/us01/U569  ( .A(\AES_ENC/us01/n929 ), .ZN(\AES_ENC/us01/n619 ) );
INV_X4 \AES_ENC/us01/U568  ( .A(\AES_ENC/us01/n1091 ), .ZN(\AES_ENC/us01/n618 ) );
INV_X4 \AES_ENC/us01/U567  ( .A(\AES_ENC/us01/n826 ), .ZN(\AES_ENC/us01/n617 ) );
INV_X4 \AES_ENC/us01/U566  ( .A(\AES_ENC/us01/n1031 ), .ZN(\AES_ENC/us01/n616 ) );
INV_X4 \AES_ENC/us01/U565  ( .A(\AES_ENC/us01/n1054 ), .ZN(\AES_ENC/us01/n615 ) );
INV_X4 \AES_ENC/us01/U564  ( .A(\AES_ENC/us01/n1025 ), .ZN(\AES_ENC/us01/n614 ) );
INV_X4 \AES_ENC/us01/U563  ( .A(\AES_ENC/us01/n990 ), .ZN(\AES_ENC/us01/n613 ) );
INV_X4 \AES_ENC/us01/U562  ( .A(\AES_ENC/sa01 [4]), .ZN(\AES_ENC/us01/n612 ));
INV_X4 \AES_ENC/us01/U561  ( .A(\AES_ENC/us01/n881 ), .ZN(\AES_ENC/us01/n611 ) );
INV_X4 \AES_ENC/us01/U560  ( .A(\AES_ENC/us01/n1022 ), .ZN(\AES_ENC/us01/n610 ) );
INV_X4 \AES_ENC/us01/U559  ( .A(\AES_ENC/us01/n1120 ), .ZN(\AES_ENC/us01/n609 ) );
INV_X4 \AES_ENC/us01/U558  ( .A(\AES_ENC/us01/n977 ), .ZN(\AES_ENC/us01/n608 ) );
INV_X4 \AES_ENC/us01/U557  ( .A(\AES_ENC/us01/n926 ), .ZN(\AES_ENC/us01/n607 ) );
INV_X4 \AES_ENC/us01/U556  ( .A(\AES_ENC/us01/n910 ), .ZN(\AES_ENC/us01/n606 ) );
INV_X4 \AES_ENC/us01/U555  ( .A(\AES_ENC/us01/n1121 ), .ZN(\AES_ENC/us01/n605 ) );
INV_X4 \AES_ENC/us01/U554  ( .A(\AES_ENC/us01/n1009 ), .ZN(\AES_ENC/us01/n604 ) );
INV_X4 \AES_ENC/us01/U553  ( .A(\AES_ENC/us01/n1080 ), .ZN(\AES_ENC/us01/n602 ) );
INV_X4 \AES_ENC/us01/U552  ( .A(\AES_ENC/us01/n821 ), .ZN(\AES_ENC/us01/n600 ) );
INV_X4 \AES_ENC/us01/U551  ( .A(\AES_ENC/us01/n1013 ), .ZN(\AES_ENC/us01/n599 ) );
INV_X4 \AES_ENC/us01/U550  ( .A(\AES_ENC/us01/n1058 ), .ZN(\AES_ENC/us01/n598 ) );
INV_X4 \AES_ENC/us01/U549  ( .A(\AES_ENC/us01/n906 ), .ZN(\AES_ENC/us01/n597 ) );
INV_X4 \AES_ENC/us01/U548  ( .A(\AES_ENC/us01/n1048 ), .ZN(\AES_ENC/us01/n595 ) );
INV_X4 \AES_ENC/us01/U547  ( .A(\AES_ENC/us01/n974 ), .ZN(\AES_ENC/us01/n594 ) );
INV_X4 \AES_ENC/us01/U546  ( .A(\AES_ENC/sa01 [2]), .ZN(\AES_ENC/us01/n593 ));
INV_X4 \AES_ENC/us01/U545  ( .A(\AES_ENC/us01/n800 ), .ZN(\AES_ENC/us01/n592 ) );
INV_X4 \AES_ENC/us01/U544  ( .A(\AES_ENC/us01/n925 ), .ZN(\AES_ENC/us01/n591 ) );
INV_X4 \AES_ENC/us01/U543  ( .A(\AES_ENC/us01/n824 ), .ZN(\AES_ENC/us01/n590 ) );
INV_X4 \AES_ENC/us01/U542  ( .A(\AES_ENC/us01/n959 ), .ZN(\AES_ENC/us01/n589 ) );
INV_X4 \AES_ENC/us01/U541  ( .A(\AES_ENC/us01/n779 ), .ZN(\AES_ENC/us01/n588 ) );
INV_X4 \AES_ENC/us01/U540  ( .A(\AES_ENC/us01/n794 ), .ZN(\AES_ENC/us01/n585 ) );
INV_X4 \AES_ENC/us01/U539  ( .A(\AES_ENC/us01/n880 ), .ZN(\AES_ENC/us01/n583 ) );
INV_X4 \AES_ENC/us01/U538  ( .A(\AES_ENC/sa01 [7]), .ZN(\AES_ENC/us01/n581 ));
INV_X4 \AES_ENC/us01/U537  ( .A(\AES_ENC/us01/n992 ), .ZN(\AES_ENC/us01/n578 ) );
INV_X4 \AES_ENC/us01/U536  ( .A(\AES_ENC/us01/n1114 ), .ZN(\AES_ENC/us01/n577 ) );
INV_X4 \AES_ENC/us01/U535  ( .A(\AES_ENC/us01/n1092 ), .ZN(\AES_ENC/us01/n574 ) );
NOR2_X2 \AES_ENC/us01/U534  ( .A1(\AES_ENC/sa01 [0]), .A2(\AES_ENC/sa01 [6]),.ZN(\AES_ENC/us01/n1090 ) );
NOR2_X2 \AES_ENC/us01/U533  ( .A1(\AES_ENC/us01/n627 ), .A2(\AES_ENC/sa01 [6]), .ZN(\AES_ENC/us01/n1070 ) );
NOR2_X2 \AES_ENC/us01/U532  ( .A1(\AES_ENC/sa01 [4]), .A2(\AES_ENC/sa01 [3]),.ZN(\AES_ENC/us01/n1025 ) );
INV_X4 \AES_ENC/us01/U531  ( .A(\AES_ENC/us01/n569 ), .ZN(\AES_ENC/us01/n572 ) );
NOR2_X2 \AES_ENC/us01/U530  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n765 ) );
NOR2_X2 \AES_ENC/us01/U529  ( .A1(\AES_ENC/sa01 [4]), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n764 ) );
NOR2_X2 \AES_ENC/us01/U528  ( .A1(\AES_ENC/us01/n765 ), .A2(\AES_ENC/us01/n764 ), .ZN(\AES_ENC/us01/n766 ) );
NOR2_X2 \AES_ENC/us01/U527  ( .A1(\AES_ENC/us01/n766 ), .A2(\AES_ENC/us01/n589 ), .ZN(\AES_ENC/us01/n767 ) );
NOR3_X2 \AES_ENC/us01/U526  ( .A1(\AES_ENC/us01/n581 ), .A2(\AES_ENC/sa01 [5]), .A3(\AES_ENC/us01/n704 ), .ZN(\AES_ENC/us01/n706 ));
NOR2_X2 \AES_ENC/us01/U525  ( .A1(\AES_ENC/us01/n1117 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n707 ) );
NOR2_X2 \AES_ENC/us01/U524  ( .A1(\AES_ENC/sa01 [4]), .A2(\AES_ENC/us01/n574 ), .ZN(\AES_ENC/us01/n705 ) );
NOR3_X2 \AES_ENC/us01/U523  ( .A1(\AES_ENC/us01/n707 ), .A2(\AES_ENC/us01/n706 ), .A3(\AES_ENC/us01/n705 ), .ZN(\AES_ENC/us01/n713 ) );
INV_X4 \AES_ENC/us01/U522  ( .A(\AES_ENC/sa01 [3]), .ZN(\AES_ENC/us01/n624 ));
NAND3_X2 \AES_ENC/us01/U521  ( .A1(\AES_ENC/us01/n652 ), .A2(\AES_ENC/us01/n596 ), .A3(\AES_ENC/sa01 [7]), .ZN(\AES_ENC/us01/n653 ));
NOR2_X2 \AES_ENC/us01/U520  ( .A1(\AES_ENC/us01/n593 ), .A2(\AES_ENC/sa01 [5]), .ZN(\AES_ENC/us01/n925 ) );
NOR2_X2 \AES_ENC/us01/U519  ( .A1(\AES_ENC/sa01 [5]), .A2(\AES_ENC/sa01 [2]),.ZN(\AES_ENC/us01/n974 ) );
INV_X4 \AES_ENC/us01/U518  ( .A(\AES_ENC/sa01 [5]), .ZN(\AES_ENC/us01/n596 ));
NOR2_X2 \AES_ENC/us01/U517  ( .A1(\AES_ENC/us01/n593 ), .A2(\AES_ENC/sa01 [7]), .ZN(\AES_ENC/us01/n779 ) );
NAND3_X2 \AES_ENC/us01/U516  ( .A1(\AES_ENC/us01/n679 ), .A2(\AES_ENC/us01/n678 ), .A3(\AES_ENC/us01/n677 ), .ZN(\AES_ENC/sa01_sub[0] ) );
NOR2_X2 \AES_ENC/us01/U515  ( .A1(\AES_ENC/us01/n596 ), .A2(\AES_ENC/sa01 [2]), .ZN(\AES_ENC/us01/n1048 ) );
NOR4_X2 \AES_ENC/us01/U512  ( .A1(\AES_ENC/us01/n633 ), .A2(\AES_ENC/us01/n632 ), .A3(\AES_ENC/us01/n631 ), .A4(\AES_ENC/us01/n630 ), .ZN(\AES_ENC/us01/n634 ) );
NOR2_X2 \AES_ENC/us01/U510  ( .A1(\AES_ENC/us01/n629 ), .A2(\AES_ENC/us01/n628 ), .ZN(\AES_ENC/us01/n635 ) );
NAND3_X2 \AES_ENC/us01/U509  ( .A1(\AES_ENC/sa01 [2]), .A2(\AES_ENC/sa01 [7]), .A3(\AES_ENC/us01/n1059 ), .ZN(\AES_ENC/us01/n636 ) );
NOR2_X2 \AES_ENC/us01/U508  ( .A1(\AES_ENC/sa01 [7]), .A2(\AES_ENC/sa01 [2]),.ZN(\AES_ENC/us01/n794 ) );
NOR2_X2 \AES_ENC/us01/U507  ( .A1(\AES_ENC/sa01 [4]), .A2(\AES_ENC/sa01 [1]),.ZN(\AES_ENC/us01/n1102 ) );
NOR2_X2 \AES_ENC/us01/U506  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/sa01 [3]), .ZN(\AES_ENC/us01/n1053 ) );
NOR2_X2 \AES_ENC/us01/U505  ( .A1(\AES_ENC/us01/n588 ), .A2(\AES_ENC/sa01 [5]), .ZN(\AES_ENC/us01/n1024 ) );
NOR2_X2 \AES_ENC/us01/U504  ( .A1(\AES_ENC/us01/n577 ), .A2(\AES_ENC/sa01 [2]), .ZN(\AES_ENC/us01/n1093 ) );
NOR2_X2 \AES_ENC/us01/U503  ( .A1(\AES_ENC/us01/n585 ), .A2(\AES_ENC/sa01 [5]), .ZN(\AES_ENC/us01/n1094 ) );
NOR2_X2 \AES_ENC/us01/U502  ( .A1(\AES_ENC/us01/n612 ), .A2(\AES_ENC/sa01 [3]), .ZN(\AES_ENC/us01/n931 ) );
INV_X4 \AES_ENC/us01/U501  ( .A(\AES_ENC/us01/n570 ), .ZN(\AES_ENC/us01/n573 ) );
NOR2_X2 \AES_ENC/us01/U500  ( .A1(\AES_ENC/us01/n1053 ), .A2(\AES_ENC/us01/n1095 ), .ZN(\AES_ENC/us01/n639 ) );
NOR3_X2 \AES_ENC/us01/U499  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n573 ), .A3(\AES_ENC/us01/n1074 ), .ZN(\AES_ENC/us01/n641 ) );
NOR2_X2 \AES_ENC/us01/U498  ( .A1(\AES_ENC/us01/n639 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n640 ) );
NOR2_X2 \AES_ENC/us01/U497  ( .A1(\AES_ENC/us01/n641 ), .A2(\AES_ENC/us01/n640 ), .ZN(\AES_ENC/us01/n646 ) );
NOR3_X2 \AES_ENC/us01/U496  ( .A1(\AES_ENC/us01/n995 ), .A2(\AES_ENC/us01/n578 ), .A3(\AES_ENC/us01/n994 ), .ZN(\AES_ENC/us01/n1002 ) );
NOR2_X2 \AES_ENC/us01/U495  ( .A1(\AES_ENC/us01/n909 ), .A2(\AES_ENC/us01/n908 ), .ZN(\AES_ENC/us01/n920 ) );
NOR2_X2 \AES_ENC/us01/U494  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n823 ) );
NOR2_X2 \AES_ENC/us01/U492  ( .A1(\AES_ENC/us01/n612 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n822 ) );
NOR2_X2 \AES_ENC/us01/U491  ( .A1(\AES_ENC/us01/n823 ), .A2(\AES_ENC/us01/n822 ), .ZN(\AES_ENC/us01/n825 ) );
NOR2_X2 \AES_ENC/us01/U490  ( .A1(\AES_ENC/sa01 [1]), .A2(\AES_ENC/us01/n601 ), .ZN(\AES_ENC/us01/n913 ) );
NOR2_X2 \AES_ENC/us01/U489  ( .A1(\AES_ENC/us01/n913 ), .A2(\AES_ENC/us01/n1091 ), .ZN(\AES_ENC/us01/n914 ) );
NOR2_X2 \AES_ENC/us01/U488  ( .A1(\AES_ENC/us01/n826 ), .A2(\AES_ENC/us01/n572 ), .ZN(\AES_ENC/us01/n827 ) );
NOR3_X2 \AES_ENC/us01/U487  ( .A1(\AES_ENC/us01/n769 ), .A2(\AES_ENC/us01/n768 ), .A3(\AES_ENC/us01/n767 ), .ZN(\AES_ENC/us01/n775 ) );
NOR2_X2 \AES_ENC/us01/U486  ( .A1(\AES_ENC/us01/n1056 ), .A2(\AES_ENC/us01/n1053 ), .ZN(\AES_ENC/us01/n749 ) );
NOR2_X2 \AES_ENC/us01/U483  ( .A1(\AES_ENC/us01/n749 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n752 ) );
INV_X4 \AES_ENC/us01/U482  ( .A(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n626 ));
NOR2_X2 \AES_ENC/us01/U480  ( .A1(\AES_ENC/us01/n1054 ), .A2(\AES_ENC/us01/n1053 ), .ZN(\AES_ENC/us01/n1055 ) );
OR2_X4 \AES_ENC/us01/U479  ( .A1(\AES_ENC/us01/n1094 ), .A2(\AES_ENC/us01/n1093 ), .ZN(\AES_ENC/us01/n571 ) );
AND2_X2 \AES_ENC/us01/U478  ( .A1(\AES_ENC/us01/n571 ), .A2(\AES_ENC/us01/n1095 ), .ZN(\AES_ENC/us01/n1101 ) );
NOR2_X2 \AES_ENC/us01/U477  ( .A1(\AES_ENC/us01/n1074 ), .A2(\AES_ENC/us01/n931 ), .ZN(\AES_ENC/us01/n796 ) );
NOR2_X2 \AES_ENC/us01/U474  ( .A1(\AES_ENC/us01/n796 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n797 ) );
NOR2_X2 \AES_ENC/us01/U473  ( .A1(\AES_ENC/us01/n932 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n933 ) );
NOR2_X2 \AES_ENC/us01/U472  ( .A1(\AES_ENC/us01/n929 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n935 ) );
NOR2_X2 \AES_ENC/us01/U471  ( .A1(\AES_ENC/us01/n931 ), .A2(\AES_ENC/us01/n930 ), .ZN(\AES_ENC/us01/n934 ) );
NOR3_X2 \AES_ENC/us01/U470  ( .A1(\AES_ENC/us01/n935 ), .A2(\AES_ENC/us01/n934 ), .A3(\AES_ENC/us01/n933 ), .ZN(\AES_ENC/us01/n936 ) );
NOR2_X2 \AES_ENC/us01/U469  ( .A1(\AES_ENC/us01/n612 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n1075 ) );
NOR2_X2 \AES_ENC/us01/U468  ( .A1(\AES_ENC/us01/n572 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n949 ) );
NOR2_X2 \AES_ENC/us01/U467  ( .A1(\AES_ENC/us01/n1049 ), .A2(\AES_ENC/us01/n595 ), .ZN(\AES_ENC/us01/n1051 ) );
NOR2_X2 \AES_ENC/us01/U466  ( .A1(\AES_ENC/us01/n1051 ), .A2(\AES_ENC/us01/n1050 ), .ZN(\AES_ENC/us01/n1052 ) );
NOR2_X2 \AES_ENC/us01/U465  ( .A1(\AES_ENC/us01/n1052 ), .A2(\AES_ENC/us01/n604 ), .ZN(\AES_ENC/us01/n1064 ) );
NOR2_X2 \AES_ENC/us01/U464  ( .A1(\AES_ENC/sa01 [1]), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n631 ) );
NOR2_X2 \AES_ENC/us01/U463  ( .A1(\AES_ENC/us01/n1025 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n980 ) );
NOR2_X2 \AES_ENC/us01/U462  ( .A1(\AES_ENC/us01/n1073 ), .A2(\AES_ENC/us01/n1094 ), .ZN(\AES_ENC/us01/n795 ) );
NOR2_X2 \AES_ENC/us01/U461  ( .A1(\AES_ENC/us01/n795 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n799 ) );
NOR2_X2 \AES_ENC/us01/U460  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n981 ) );
NOR2_X2 \AES_ENC/us01/U459  ( .A1(\AES_ENC/us01/n1102 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n643 ) );
NOR2_X2 \AES_ENC/us01/U458  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n624 ), .ZN(\AES_ENC/us01/n642 ) );
NOR2_X2 \AES_ENC/us01/U455  ( .A1(\AES_ENC/us01/n911 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n644 ) );
NOR4_X2 \AES_ENC/us01/U448  ( .A1(\AES_ENC/us01/n644 ), .A2(\AES_ENC/us01/n643 ), .A3(\AES_ENC/us01/n804 ), .A4(\AES_ENC/us01/n642 ), .ZN(\AES_ENC/us01/n645 ) );
NOR2_X2 \AES_ENC/us01/U447  ( .A1(\AES_ENC/us01/n1102 ), .A2(\AES_ENC/us01/n910 ), .ZN(\AES_ENC/us01/n932 ) );
NOR2_X2 \AES_ENC/us01/U442  ( .A1(\AES_ENC/us01/n1102 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n755 ) );
NOR2_X2 \AES_ENC/us01/U441  ( .A1(\AES_ENC/us01/n931 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n743 ) );
NOR2_X2 \AES_ENC/us01/U438  ( .A1(\AES_ENC/us01/n1072 ), .A2(\AES_ENC/us01/n1094 ), .ZN(\AES_ENC/us01/n930 ) );
NOR2_X2 \AES_ENC/us01/U435  ( .A1(\AES_ENC/us01/n1074 ), .A2(\AES_ENC/us01/n1025 ), .ZN(\AES_ENC/us01/n891 ) );
NOR2_X2 \AES_ENC/us01/U434  ( .A1(\AES_ENC/us01/n891 ), .A2(\AES_ENC/us01/n591 ), .ZN(\AES_ENC/us01/n894 ) );
NOR3_X2 \AES_ENC/us01/U433  ( .A1(\AES_ENC/us01/n601 ), .A2(\AES_ENC/sa01 [1]), .A3(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n683 ));
INV_X4 \AES_ENC/us01/U428  ( .A(\AES_ENC/us01/n931 ), .ZN(\AES_ENC/us01/n601 ) );
NOR2_X2 \AES_ENC/us01/U427  ( .A1(\AES_ENC/us01/n996 ), .A2(\AES_ENC/us01/n931 ), .ZN(\AES_ENC/us01/n704 ) );
NOR2_X2 \AES_ENC/us01/U421  ( .A1(\AES_ENC/us01/n931 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n685 ) );
NOR2_X2 \AES_ENC/us01/U420  ( .A1(\AES_ENC/us01/n1029 ), .A2(\AES_ENC/us01/n1025 ), .ZN(\AES_ENC/us01/n1079 ) );
NOR3_X2 \AES_ENC/us01/U419  ( .A1(\AES_ENC/us01/n620 ), .A2(\AES_ENC/us01/n1025 ), .A3(\AES_ENC/us01/n594 ), .ZN(\AES_ENC/us01/n945 ) );
NOR2_X2 \AES_ENC/us01/U418  ( .A1(\AES_ENC/us01/n596 ), .A2(\AES_ENC/us01/n593 ), .ZN(\AES_ENC/us01/n800 ) );
NOR3_X2 \AES_ENC/us01/U417  ( .A1(\AES_ENC/us01/n598 ), .A2(\AES_ENC/us01/n581 ), .A3(\AES_ENC/us01/n593 ), .ZN(\AES_ENC/us01/n798 ) );
NOR3_X2 \AES_ENC/us01/U416  ( .A1(\AES_ENC/us01/n592 ), .A2(\AES_ENC/us01/n572 ), .A3(\AES_ENC/us01/n589 ), .ZN(\AES_ENC/us01/n962 ) );
NOR3_X2 \AES_ENC/us01/U415  ( .A1(\AES_ENC/us01/n959 ), .A2(\AES_ENC/us01/n572 ), .A3(\AES_ENC/us01/n591 ), .ZN(\AES_ENC/us01/n768 ) );
NOR3_X2 \AES_ENC/us01/U414  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n572 ), .A3(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n694 ) );
NOR3_X2 \AES_ENC/us01/U413  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n572 ), .A3(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n895 ) );
NOR3_X2 \AES_ENC/us01/U410  ( .A1(\AES_ENC/us01/n1008 ), .A2(\AES_ENC/us01/n1007 ), .A3(\AES_ENC/us01/n1006 ), .ZN(\AES_ENC/us01/n1018 ) );
NOR4_X2 \AES_ENC/us01/U409  ( .A1(\AES_ENC/us01/n806 ), .A2(\AES_ENC/us01/n805 ), .A3(\AES_ENC/us01/n804 ), .A4(\AES_ENC/us01/n803 ), .ZN(\AES_ENC/us01/n807 ) );
NOR3_X2 \AES_ENC/us01/U406  ( .A1(\AES_ENC/us01/n799 ), .A2(\AES_ENC/us01/n798 ), .A3(\AES_ENC/us01/n797 ), .ZN(\AES_ENC/us01/n808 ) );
NOR4_X2 \AES_ENC/us01/U405  ( .A1(\AES_ENC/us01/n843 ), .A2(\AES_ENC/us01/n842 ), .A3(\AES_ENC/us01/n841 ), .A4(\AES_ENC/us01/n840 ), .ZN(\AES_ENC/us01/n844 ) );
NOR2_X2 \AES_ENC/us01/U404  ( .A1(\AES_ENC/us01/n669 ), .A2(\AES_ENC/us01/n668 ), .ZN(\AES_ENC/us01/n673 ) );
NOR4_X2 \AES_ENC/us01/U403  ( .A1(\AES_ENC/us01/n946 ), .A2(\AES_ENC/us01/n1046 ), .A3(\AES_ENC/us01/n671 ), .A4(\AES_ENC/us01/n670 ), .ZN(\AES_ENC/us01/n672 ) );
NOR3_X2 \AES_ENC/us01/U401  ( .A1(\AES_ENC/us01/n1101 ), .A2(\AES_ENC/us01/n1100 ), .A3(\AES_ENC/us01/n1099 ), .ZN(\AES_ENC/us01/n1109 ) );
NOR4_X2 \AES_ENC/us01/U400  ( .A1(\AES_ENC/us01/n711 ), .A2(\AES_ENC/us01/n710 ), .A3(\AES_ENC/us01/n709 ), .A4(\AES_ENC/us01/n708 ), .ZN(\AES_ENC/us01/n712 ) );
NOR4_X2 \AES_ENC/us01/U399  ( .A1(\AES_ENC/us01/n963 ), .A2(\AES_ENC/us01/n962 ), .A3(\AES_ENC/us01/n961 ), .A4(\AES_ENC/us01/n960 ), .ZN(\AES_ENC/us01/n964 ) );
NOR3_X2 \AES_ENC/us01/U398  ( .A1(\AES_ENC/us01/n743 ), .A2(\AES_ENC/us01/n742 ), .A3(\AES_ENC/us01/n741 ), .ZN(\AES_ENC/us01/n744 ) );
NOR2_X2 \AES_ENC/us01/U397  ( .A1(\AES_ENC/us01/n697 ), .A2(\AES_ENC/us01/n658 ), .ZN(\AES_ENC/us01/n659 ) );
NOR2_X2 \AES_ENC/us01/U396  ( .A1(\AES_ENC/us01/n1078 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n1033 ) );
NOR2_X2 \AES_ENC/us01/U393  ( .A1(\AES_ENC/us01/n1031 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n1032 ) );
NOR3_X2 \AES_ENC/us01/U390  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n1025 ), .A3(\AES_ENC/us01/n1074 ), .ZN(\AES_ENC/us01/n1035 ) );
NOR4_X2 \AES_ENC/us01/U389  ( .A1(\AES_ENC/us01/n1035 ), .A2(\AES_ENC/us01/n1034 ), .A3(\AES_ENC/us01/n1033 ), .A4(\AES_ENC/us01/n1032 ), .ZN(\AES_ENC/us01/n1036 ) );
NOR2_X2 \AES_ENC/us01/U388  ( .A1(\AES_ENC/us01/n611 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n885 ) );
NOR2_X2 \AES_ENC/us01/U387  ( .A1(\AES_ENC/us01/n601 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n882 ) );
NOR2_X2 \AES_ENC/us01/U386  ( .A1(\AES_ENC/us01/n1053 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n884 ) );
NOR4_X2 \AES_ENC/us01/U385  ( .A1(\AES_ENC/us01/n885 ), .A2(\AES_ENC/us01/n884 ), .A3(\AES_ENC/us01/n883 ), .A4(\AES_ENC/us01/n882 ), .ZN(\AES_ENC/us01/n886 ) );
NOR2_X2 \AES_ENC/us01/U384  ( .A1(\AES_ENC/us01/n825 ), .A2(\AES_ENC/us01/n590 ), .ZN(\AES_ENC/us01/n830 ) );
NOR2_X2 \AES_ENC/us01/U383  ( .A1(\AES_ENC/us01/n827 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n829 ) );
NOR2_X2 \AES_ENC/us01/U382  ( .A1(\AES_ENC/us01/n572 ), .A2(\AES_ENC/us01/n574 ), .ZN(\AES_ENC/us01/n828 ) );
NOR4_X2 \AES_ENC/us01/U374  ( .A1(\AES_ENC/us01/n831 ), .A2(\AES_ENC/us01/n830 ), .A3(\AES_ENC/us01/n829 ), .A4(\AES_ENC/us01/n828 ), .ZN(\AES_ENC/us01/n832 ) );
NOR2_X2 \AES_ENC/us01/U373  ( .A1(\AES_ENC/us01/n587 ), .A2(\AES_ENC/us01/n603 ), .ZN(\AES_ENC/us01/n1104 ) );
NOR2_X2 \AES_ENC/us01/U372  ( .A1(\AES_ENC/us01/n1102 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n1106 ) );
NOR2_X2 \AES_ENC/us01/U370  ( .A1(\AES_ENC/us01/n1103 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n1105 ) );
NOR4_X2 \AES_ENC/us01/U369  ( .A1(\AES_ENC/us01/n1107 ), .A2(\AES_ENC/us01/n1106 ), .A3(\AES_ENC/us01/n1105 ), .A4(\AES_ENC/us01/n1104 ), .ZN(\AES_ENC/us01/n1108 ) );
NOR3_X2 \AES_ENC/us01/U368  ( .A1(\AES_ENC/us01/n959 ), .A2(\AES_ENC/us01/n624 ), .A3(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n963 ) );
NOR2_X2 \AES_ENC/us01/U367  ( .A1(\AES_ENC/us01/n596 ), .A2(\AES_ENC/us01/n581 ), .ZN(\AES_ENC/us01/n1114 ) );
INV_X4 \AES_ENC/us01/U366  ( .A(\AES_ENC/us01/n1024 ), .ZN(\AES_ENC/us01/n587 ) );
NOR3_X2 \AES_ENC/us01/U365  ( .A1(\AES_ENC/us01/n910 ), .A2(\AES_ENC/us01/n1059 ), .A3(\AES_ENC/us01/n593 ), .ZN(\AES_ENC/us01/n1115 ) );
INV_X4 \AES_ENC/us01/U364  ( .A(\AES_ENC/us01/n1094 ), .ZN(\AES_ENC/us01/n584 ) );
NOR2_X2 \AES_ENC/us01/U363  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n931 ), .ZN(\AES_ENC/us01/n1100 ) );
INV_X4 \AES_ENC/us01/U354  ( .A(\AES_ENC/us01/n1093 ), .ZN(\AES_ENC/us01/n575 ) );
NOR2_X2 \AES_ENC/us01/U353  ( .A1(\AES_ENC/us01/n569 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n929 ) );
NOR2_X2 \AES_ENC/us01/U352  ( .A1(\AES_ENC/us01/n609 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n926 ) );
NOR2_X2 \AES_ENC/us01/U351  ( .A1(\AES_ENC/us01/n572 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n1095 ) );
NOR2_X2 \AES_ENC/us01/U350  ( .A1(\AES_ENC/us01/n591 ), .A2(\AES_ENC/us01/n581 ), .ZN(\AES_ENC/us01/n1010 ) );
NOR2_X2 \AES_ENC/us01/U349  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n1103 ) );
NOR2_X2 \AES_ENC/us01/U348  ( .A1(\AES_ENC/us01/n614 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n1059 ) );
NOR2_X2 \AES_ENC/us01/U347  ( .A1(\AES_ENC/sa01 [1]), .A2(\AES_ENC/us01/n1120 ), .ZN(\AES_ENC/us01/n1022 ) );
NOR2_X2 \AES_ENC/us01/U346  ( .A1(\AES_ENC/us01/n605 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n911 ) );
NOR2_X2 \AES_ENC/us01/U345  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/us01/n1025 ), .ZN(\AES_ENC/us01/n826 ) );
NOR2_X2 \AES_ENC/us01/U338  ( .A1(\AES_ENC/us01/n596 ), .A2(\AES_ENC/us01/n588 ), .ZN(\AES_ENC/us01/n1072 ) );
NOR2_X2 \AES_ENC/us01/U335  ( .A1(\AES_ENC/us01/n581 ), .A2(\AES_ENC/us01/n594 ), .ZN(\AES_ENC/us01/n956 ) );
NOR2_X2 \AES_ENC/us01/U329  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/us01/n612 ), .ZN(\AES_ENC/us01/n1121 ) );
NOR2_X2 \AES_ENC/us01/U328  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/us01/n612 ), .ZN(\AES_ENC/us01/n1058 ) );
NOR2_X2 \AES_ENC/us01/U327  ( .A1(\AES_ENC/us01/n577 ), .A2(\AES_ENC/us01/n593 ), .ZN(\AES_ENC/us01/n1073 ) );
NOR2_X2 \AES_ENC/us01/U325  ( .A1(\AES_ENC/sa01 [1]), .A2(\AES_ENC/us01/n1025 ), .ZN(\AES_ENC/us01/n1054 ) );
NOR2_X2 \AES_ENC/us01/U324  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/us01/n931 ), .ZN(\AES_ENC/us01/n1029 ) );
NOR2_X2 \AES_ENC/us01/U319  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n1056 ) );
NOR2_X2 \AES_ENC/us01/U318  ( .A1(\AES_ENC/us01/n585 ), .A2(\AES_ENC/us01/n596 ), .ZN(\AES_ENC/us01/n1050 ) );
NOR2_X2 \AES_ENC/us01/U317  ( .A1(\AES_ENC/us01/n1121 ), .A2(\AES_ENC/us01/n1025 ), .ZN(\AES_ENC/us01/n1120 ) );
NOR2_X2 \AES_ENC/us01/U316  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/us01/n572 ), .ZN(\AES_ENC/us01/n1074 ) );
NOR2_X2 \AES_ENC/us01/U315  ( .A1(\AES_ENC/us01/n1058 ), .A2(\AES_ENC/us01/n1054 ), .ZN(\AES_ENC/us01/n878 ) );
NOR2_X2 \AES_ENC/us01/U314  ( .A1(\AES_ENC/us01/n878 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n879 ) );
NOR2_X2 \AES_ENC/us01/U312  ( .A1(\AES_ENC/us01/n880 ), .A2(\AES_ENC/us01/n879 ), .ZN(\AES_ENC/us01/n887 ) );
NOR2_X2 \AES_ENC/us01/U311  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n625 ), .ZN(\AES_ENC/us01/n957 ) );
NOR2_X2 \AES_ENC/us01/U310  ( .A1(\AES_ENC/us01/n958 ), .A2(\AES_ENC/us01/n957 ), .ZN(\AES_ENC/us01/n965 ) );
NOR3_X2 \AES_ENC/us01/U309  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n1091 ), .A3(\AES_ENC/us01/n1022 ), .ZN(\AES_ENC/us01/n720 ) );
NOR3_X2 \AES_ENC/us01/U303  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n1054 ), .A3(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n719 ) );
NOR2_X2 \AES_ENC/us01/U302  ( .A1(\AES_ENC/us01/n720 ), .A2(\AES_ENC/us01/n719 ), .ZN(\AES_ENC/us01/n726 ) );
NOR2_X2 \AES_ENC/us01/U300  ( .A1(\AES_ENC/us01/n585 ), .A2(\AES_ENC/us01/n613 ), .ZN(\AES_ENC/us01/n865 ) );
NOR2_X2 \AES_ENC/us01/U299  ( .A1(\AES_ENC/us01/n1059 ), .A2(\AES_ENC/us01/n1058 ), .ZN(\AES_ENC/us01/n1060 ) );
NOR2_X2 \AES_ENC/us01/U298  ( .A1(\AES_ENC/us01/n1095 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n668 ) );
NOR2_X2 \AES_ENC/us01/U297  ( .A1(\AES_ENC/us01/n911 ), .A2(\AES_ENC/us01/n910 ), .ZN(\AES_ENC/us01/n912 ) );
NOR2_X2 \AES_ENC/us01/U296  ( .A1(\AES_ENC/us01/n912 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n916 ) );
NOR2_X2 \AES_ENC/us01/U295  ( .A1(\AES_ENC/us01/n826 ), .A2(\AES_ENC/us01/n573 ), .ZN(\AES_ENC/us01/n750 ) );
NOR2_X2 \AES_ENC/us01/U294  ( .A1(\AES_ENC/us01/n750 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n751 ) );
NOR2_X2 \AES_ENC/us01/U293  ( .A1(\AES_ENC/us01/n907 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n908 ) );
NOR2_X2 \AES_ENC/us01/U292  ( .A1(\AES_ENC/us01/n990 ), .A2(\AES_ENC/us01/n926 ), .ZN(\AES_ENC/us01/n780 ) );
NOR2_X2 \AES_ENC/us01/U291  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n606 ), .ZN(\AES_ENC/us01/n838 ) );
NOR2_X2 \AES_ENC/us01/U290  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n621 ), .ZN(\AES_ENC/us01/n837 ) );
NOR2_X2 \AES_ENC/us01/U284  ( .A1(\AES_ENC/us01/n838 ), .A2(\AES_ENC/us01/n837 ), .ZN(\AES_ENC/us01/n845 ) );
NOR2_X2 \AES_ENC/us01/U283  ( .A1(\AES_ENC/us01/n1022 ), .A2(\AES_ENC/us01/n1058 ), .ZN(\AES_ENC/us01/n740 ) );
NOR2_X2 \AES_ENC/us01/U282  ( .A1(\AES_ENC/us01/n740 ), .A2(\AES_ENC/us01/n594 ), .ZN(\AES_ENC/us01/n742 ) );
NOR2_X2 \AES_ENC/us01/U281  ( .A1(\AES_ENC/us01/n1098 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n1099 ) );
NOR2_X2 \AES_ENC/us01/U280  ( .A1(\AES_ENC/us01/n1120 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n993 ) );
NOR2_X2 \AES_ENC/us01/U279  ( .A1(\AES_ENC/us01/n993 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n994 ) );
NOR2_X2 \AES_ENC/us01/U273  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n609 ), .ZN(\AES_ENC/us01/n1026 ) );
NOR2_X2 \AES_ENC/us01/U272  ( .A1(\AES_ENC/us01/n573 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n1027 ) );
NOR2_X2 \AES_ENC/us01/U271  ( .A1(\AES_ENC/us01/n1027 ), .A2(\AES_ENC/us01/n1026 ), .ZN(\AES_ENC/us01/n1028 ) );
NOR2_X2 \AES_ENC/us01/U270  ( .A1(\AES_ENC/us01/n1029 ), .A2(\AES_ENC/us01/n1028 ), .ZN(\AES_ENC/us01/n1034 ) );
NOR4_X2 \AES_ENC/us01/U269  ( .A1(\AES_ENC/us01/n757 ), .A2(\AES_ENC/us01/n756 ), .A3(\AES_ENC/us01/n755 ), .A4(\AES_ENC/us01/n754 ), .ZN(\AES_ENC/us01/n758 ) );
NOR2_X2 \AES_ENC/us01/U268  ( .A1(\AES_ENC/us01/n752 ), .A2(\AES_ENC/us01/n751 ), .ZN(\AES_ENC/us01/n759 ) );
NOR2_X2 \AES_ENC/us01/U267  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n1071 ), .ZN(\AES_ENC/us01/n669 ) );
NOR2_X2 \AES_ENC/us01/U263  ( .A1(\AES_ENC/us01/n1056 ), .A2(\AES_ENC/us01/n990 ), .ZN(\AES_ENC/us01/n991 ) );
NOR2_X2 \AES_ENC/us01/U262  ( .A1(\AES_ENC/us01/n991 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n995 ) );
NOR2_X2 \AES_ENC/us01/U258  ( .A1(\AES_ENC/us01/n588 ), .A2(\AES_ENC/us01/n598 ), .ZN(\AES_ENC/us01/n1008 ) );
NOR2_X2 \AES_ENC/us01/U255  ( .A1(\AES_ENC/us01/n839 ), .A2(\AES_ENC/us01/n603 ), .ZN(\AES_ENC/us01/n693 ) );
NOR2_X2 \AES_ENC/us01/U254  ( .A1(\AES_ENC/us01/n587 ), .A2(\AES_ENC/us01/n906 ), .ZN(\AES_ENC/us01/n741 ) );
NOR2_X2 \AES_ENC/us01/U253  ( .A1(\AES_ENC/us01/n1054 ), .A2(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n763 ) );
NOR2_X2 \AES_ENC/us01/U252  ( .A1(\AES_ENC/us01/n763 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n769 ) );
NOR2_X2 \AES_ENC/us01/U251  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n618 ), .ZN(\AES_ENC/us01/n1007 ) );
NOR2_X2 \AES_ENC/us01/U250  ( .A1(\AES_ENC/us01/n591 ), .A2(\AES_ENC/us01/n599 ), .ZN(\AES_ENC/us01/n1123 ) );
NOR2_X2 \AES_ENC/us01/U243  ( .A1(\AES_ENC/us01/n591 ), .A2(\AES_ENC/us01/n598 ), .ZN(\AES_ENC/us01/n710 ) );
INV_X4 \AES_ENC/us01/U242  ( .A(\AES_ENC/us01/n1029 ), .ZN(\AES_ENC/us01/n603 ) );
NOR2_X2 \AES_ENC/us01/U241  ( .A1(\AES_ENC/us01/n594 ), .A2(\AES_ENC/us01/n607 ), .ZN(\AES_ENC/us01/n883 ) );
NOR2_X2 \AES_ENC/us01/U240  ( .A1(\AES_ENC/us01/n623 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n1125 ) );
NOR2_X2 \AES_ENC/us01/U239  ( .A1(\AES_ENC/us01/n990 ), .A2(\AES_ENC/us01/n929 ), .ZN(\AES_ENC/us01/n892 ) );
NOR2_X2 \AES_ENC/us01/U238  ( .A1(\AES_ENC/us01/n892 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n893 ) );
NOR2_X2 \AES_ENC/us01/U237  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n621 ), .ZN(\AES_ENC/us01/n950 ) );
NOR2_X2 \AES_ENC/us01/U236  ( .A1(\AES_ENC/us01/n1079 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n1082 ) );
NOR2_X2 \AES_ENC/us01/U235  ( .A1(\AES_ENC/us01/n910 ), .A2(\AES_ENC/us01/n1056 ), .ZN(\AES_ENC/us01/n941 ) );
NOR2_X2 \AES_ENC/us01/U234  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n1077 ), .ZN(\AES_ENC/us01/n841 ) );
NOR2_X2 \AES_ENC/us01/U229  ( .A1(\AES_ENC/us01/n601 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n630 ) );
NOR2_X2 \AES_ENC/us01/U228  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n621 ), .ZN(\AES_ENC/us01/n806 ) );
NOR2_X2 \AES_ENC/us01/U227  ( .A1(\AES_ENC/us01/n601 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n948 ) );
NOR2_X2 \AES_ENC/us01/U226  ( .A1(\AES_ENC/us01/n587 ), .A2(\AES_ENC/us01/n620 ), .ZN(\AES_ENC/us01/n997 ) );
NOR2_X2 \AES_ENC/us01/U225  ( .A1(\AES_ENC/us01/n1121 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n1122 ) );
NOR2_X2 \AES_ENC/us01/U223  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n1023 ), .ZN(\AES_ENC/us01/n756 ) );
NOR2_X2 \AES_ENC/us01/U222  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n621 ), .ZN(\AES_ENC/us01/n870 ) );
NOR2_X2 \AES_ENC/us01/U221  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n569 ), .ZN(\AES_ENC/us01/n947 ) );
NOR2_X2 \AES_ENC/us01/U217  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n1077 ), .ZN(\AES_ENC/us01/n1084 ) );
NOR2_X2 \AES_ENC/us01/U213  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n855 ), .ZN(\AES_ENC/us01/n709 ) );
NOR2_X2 \AES_ENC/us01/U212  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n620 ), .ZN(\AES_ENC/us01/n868 ) );
NOR2_X2 \AES_ENC/us01/U211  ( .A1(\AES_ENC/us01/n1120 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n1124 ) );
NOR2_X2 \AES_ENC/us01/U210  ( .A1(\AES_ENC/us01/n1120 ), .A2(\AES_ENC/us01/n839 ), .ZN(\AES_ENC/us01/n842 ) );
NOR2_X2 \AES_ENC/us01/U209  ( .A1(\AES_ENC/us01/n1120 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n696 ) );
NOR2_X2 \AES_ENC/us01/U208  ( .A1(\AES_ENC/us01/n1074 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n1076 ) );
NOR2_X2 \AES_ENC/us01/U207  ( .A1(\AES_ENC/us01/n1074 ), .A2(\AES_ENC/us01/n609 ), .ZN(\AES_ENC/us01/n781 ) );
NOR3_X2 \AES_ENC/us01/U201  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n1056 ), .A3(\AES_ENC/us01/n990 ), .ZN(\AES_ENC/us01/n979 ) );
NOR3_X2 \AES_ENC/us01/U200  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n1058 ), .A3(\AES_ENC/us01/n1059 ), .ZN(\AES_ENC/us01/n854 ) );
NOR2_X2 \AES_ENC/us01/U199  ( .A1(\AES_ENC/us01/n996 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n869 ) );
NOR2_X2 \AES_ENC/us01/U198  ( .A1(\AES_ENC/us01/n1056 ), .A2(\AES_ENC/us01/n1074 ), .ZN(\AES_ENC/us01/n1057 ) );
NOR3_X2 \AES_ENC/us01/U197  ( .A1(\AES_ENC/us01/n588 ), .A2(\AES_ENC/us01/n1120 ), .A3(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n978 ) );
NOR2_X2 \AES_ENC/us01/U196  ( .A1(\AES_ENC/us01/n996 ), .A2(\AES_ENC/us01/n911 ), .ZN(\AES_ENC/us01/n1116 ) );
NOR2_X2 \AES_ENC/us01/U195  ( .A1(\AES_ENC/us01/n1074 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n754 ) );
NOR2_X2 \AES_ENC/us01/U194  ( .A1(\AES_ENC/us01/n926 ), .A2(\AES_ENC/us01/n1103 ), .ZN(\AES_ENC/us01/n977 ) );
NOR2_X2 \AES_ENC/us01/U187  ( .A1(\AES_ENC/us01/n839 ), .A2(\AES_ENC/us01/n824 ), .ZN(\AES_ENC/us01/n1092 ) );
NOR2_X2 \AES_ENC/us01/U186  ( .A1(\AES_ENC/us01/n573 ), .A2(\AES_ENC/us01/n1074 ), .ZN(\AES_ENC/us01/n684 ) );
NOR2_X2 \AES_ENC/us01/U185  ( .A1(\AES_ENC/us01/n826 ), .A2(\AES_ENC/us01/n1059 ), .ZN(\AES_ENC/us01/n907 ) );
NOR3_X2 \AES_ENC/us01/U184  ( .A1(\AES_ENC/us01/n577 ), .A2(\AES_ENC/us01/n1115 ), .A3(\AES_ENC/us01/n600 ), .ZN(\AES_ENC/us01/n831 ) );
NOR3_X2 \AES_ENC/us01/U183  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n1056 ), .A3(\AES_ENC/us01/n990 ), .ZN(\AES_ENC/us01/n896 ) );
NOR3_X2 \AES_ENC/us01/U182  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n573 ), .A3(\AES_ENC/us01/n1013 ), .ZN(\AES_ENC/us01/n670 ) );
NOR3_X2 \AES_ENC/us01/U181  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n1091 ), .A3(\AES_ENC/us01/n1022 ), .ZN(\AES_ENC/us01/n843 ) );
NOR2_X2 \AES_ENC/us01/U180  ( .A1(\AES_ENC/us01/n1029 ), .A2(\AES_ENC/us01/n1095 ), .ZN(\AES_ENC/us01/n735 ) );
NOR2_X2 \AES_ENC/us01/U174  ( .A1(\AES_ENC/us01/n1100 ), .A2(\AES_ENC/us01/n854 ), .ZN(\AES_ENC/us01/n860 ) );
NOR4_X2 \AES_ENC/us01/U173  ( .A1(\AES_ENC/us01/n1125 ), .A2(\AES_ENC/us01/n1124 ), .A3(\AES_ENC/us01/n1123 ), .A4(\AES_ENC/us01/n1122 ), .ZN(\AES_ENC/us01/n1126 ) );
NOR4_X2 \AES_ENC/us01/U172  ( .A1(\AES_ENC/us01/n1084 ), .A2(\AES_ENC/us01/n1083 ), .A3(\AES_ENC/us01/n1082 ), .A4(\AES_ENC/us01/n1081 ), .ZN(\AES_ENC/us01/n1085 ) );
NOR2_X2 \AES_ENC/us01/U171  ( .A1(\AES_ENC/us01/n1076 ), .A2(\AES_ENC/us01/n1075 ), .ZN(\AES_ENC/us01/n1086 ) );
NOR4_X2 \AES_ENC/us01/U170  ( .A1(\AES_ENC/us01/n983 ), .A2(\AES_ENC/us01/n982 ), .A3(\AES_ENC/us01/n981 ), .A4(\AES_ENC/us01/n980 ), .ZN(\AES_ENC/us01/n984 ) );
NOR2_X2 \AES_ENC/us01/U169  ( .A1(\AES_ENC/us01/n979 ), .A2(\AES_ENC/us01/n978 ), .ZN(\AES_ENC/us01/n985 ) );
NAND3_X2 \AES_ENC/us01/U168  ( .A1(\AES_ENC/us01/n569 ), .A2(\AES_ENC/us01/n603 ), .A3(\AES_ENC/us01/n681 ), .ZN(\AES_ENC/us01/n691 ) );
NOR2_X2 \AES_ENC/us01/U162  ( .A1(\AES_ENC/us01/n683 ), .A2(\AES_ENC/us01/n682 ), .ZN(\AES_ENC/us01/n690 ) );
NOR3_X2 \AES_ENC/us01/U161  ( .A1(\AES_ENC/us01/n695 ), .A2(\AES_ENC/us01/n694 ), .A3(\AES_ENC/us01/n693 ), .ZN(\AES_ENC/us01/n700 ) );
NOR4_X2 \AES_ENC/us01/U160  ( .A1(\AES_ENC/us01/n983 ), .A2(\AES_ENC/us01/n698 ), .A3(\AES_ENC/us01/n697 ), .A4(\AES_ENC/us01/n696 ), .ZN(\AES_ENC/us01/n699 ) );
NOR4_X2 \AES_ENC/us01/U159  ( .A1(\AES_ENC/us01/n896 ), .A2(\AES_ENC/us01/n895 ), .A3(\AES_ENC/us01/n894 ), .A4(\AES_ENC/us01/n893 ), .ZN(\AES_ENC/us01/n897 ) );
NOR2_X2 \AES_ENC/us01/U158  ( .A1(\AES_ENC/us01/n866 ), .A2(\AES_ENC/us01/n865 ), .ZN(\AES_ENC/us01/n872 ) );
NOR4_X2 \AES_ENC/us01/U157  ( .A1(\AES_ENC/us01/n870 ), .A2(\AES_ENC/us01/n869 ), .A3(\AES_ENC/us01/n868 ), .A4(\AES_ENC/us01/n867 ), .ZN(\AES_ENC/us01/n871 ) );
NOR2_X2 \AES_ENC/us01/U156  ( .A1(\AES_ENC/us01/n946 ), .A2(\AES_ENC/us01/n945 ), .ZN(\AES_ENC/us01/n952 ) );
NOR4_X2 \AES_ENC/us01/U155  ( .A1(\AES_ENC/us01/n950 ), .A2(\AES_ENC/us01/n949 ), .A3(\AES_ENC/us01/n948 ), .A4(\AES_ENC/us01/n947 ), .ZN(\AES_ENC/us01/n951 ) );
NOR3_X2 \AES_ENC/us01/U154  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n1054 ), .A3(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n961 ) );
NOR3_X2 \AES_ENC/us01/U153  ( .A1(\AES_ENC/us01/n609 ), .A2(\AES_ENC/us01/n1074 ), .A3(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n671 ) );
NOR2_X2 \AES_ENC/us01/U152  ( .A1(\AES_ENC/us01/n1057 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n1062 ) );
NOR2_X2 \AES_ENC/us01/U143  ( .A1(\AES_ENC/us01/n1055 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n1063 ) );
NOR2_X2 \AES_ENC/us01/U142  ( .A1(\AES_ENC/us01/n1060 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n1061 ) );
NOR4_X2 \AES_ENC/us01/U141  ( .A1(\AES_ENC/us01/n1064 ), .A2(\AES_ENC/us01/n1063 ), .A3(\AES_ENC/us01/n1062 ), .A4(\AES_ENC/us01/n1061 ), .ZN(\AES_ENC/us01/n1065 ) );
NOR2_X2 \AES_ENC/us01/U140  ( .A1(\AES_ENC/us01/n735 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n687 ) );
NOR2_X2 \AES_ENC/us01/U132  ( .A1(\AES_ENC/us01/n684 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n688 ) );
NOR2_X2 \AES_ENC/us01/U131  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n622 ), .ZN(\AES_ENC/us01/n686 ) );
NOR4_X2 \AES_ENC/us01/U130  ( .A1(\AES_ENC/us01/n688 ), .A2(\AES_ENC/us01/n687 ), .A3(\AES_ENC/us01/n686 ), .A4(\AES_ENC/us01/n685 ), .ZN(\AES_ENC/us01/n689 ) );
NOR2_X2 \AES_ENC/us01/U129  ( .A1(\AES_ENC/us01/n594 ), .A2(\AES_ENC/us01/n599 ), .ZN(\AES_ENC/us01/n771 ) );
NOR2_X2 \AES_ENC/us01/U128  ( .A1(\AES_ENC/us01/n1103 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n772 ) );
NOR2_X2 \AES_ENC/us01/U127  ( .A1(\AES_ENC/us01/n592 ), .A2(\AES_ENC/us01/n615 ), .ZN(\AES_ENC/us01/n773 ) );
NOR4_X2 \AES_ENC/us01/U126  ( .A1(\AES_ENC/us01/n773 ), .A2(\AES_ENC/us01/n772 ), .A3(\AES_ENC/us01/n771 ), .A4(\AES_ENC/us01/n770 ), .ZN(\AES_ENC/us01/n774 ) );
NOR2_X2 \AES_ENC/us01/U121  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n608 ), .ZN(\AES_ENC/us01/n858 ) );
NOR2_X2 \AES_ENC/us01/U120  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n855 ), .ZN(\AES_ENC/us01/n857 ) );
NOR2_X2 \AES_ENC/us01/U119  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n617 ), .ZN(\AES_ENC/us01/n856 ) );
NOR4_X2 \AES_ENC/us01/U118  ( .A1(\AES_ENC/us01/n858 ), .A2(\AES_ENC/us01/n857 ), .A3(\AES_ENC/us01/n856 ), .A4(\AES_ENC/us01/n958 ), .ZN(\AES_ENC/us01/n859 ) );
NOR3_X2 \AES_ENC/us01/U117  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n1120 ), .A3(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n918 ) );
NOR3_X2 \AES_ENC/us01/U116  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n573 ), .A3(\AES_ENC/us01/n1013 ), .ZN(\AES_ENC/us01/n917 ) );
NOR2_X2 \AES_ENC/us01/U115  ( .A1(\AES_ENC/us01/n914 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n915 ) );
NOR4_X2 \AES_ENC/us01/U106  ( .A1(\AES_ENC/us01/n918 ), .A2(\AES_ENC/us01/n917 ), .A3(\AES_ENC/us01/n916 ), .A4(\AES_ENC/us01/n915 ), .ZN(\AES_ENC/us01/n919 ) );
NOR2_X2 \AES_ENC/us01/U105  ( .A1(\AES_ENC/us01/n780 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n784 ) );
NOR2_X2 \AES_ENC/us01/U104  ( .A1(\AES_ENC/us01/n1117 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n782 ) );
NOR2_X2 \AES_ENC/us01/U103  ( .A1(\AES_ENC/us01/n781 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n783 ) );
NOR4_X2 \AES_ENC/us01/U102  ( .A1(\AES_ENC/us01/n880 ), .A2(\AES_ENC/us01/n784 ), .A3(\AES_ENC/us01/n783 ), .A4(\AES_ENC/us01/n782 ), .ZN(\AES_ENC/us01/n785 ) );
NOR2_X2 \AES_ENC/us01/U101  ( .A1(\AES_ENC/us01/n597 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n814 ) );
NOR2_X2 \AES_ENC/us01/U100  ( .A1(\AES_ENC/us01/n907 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n813 ) );
NOR3_X2 \AES_ENC/us01/U95  ( .A1(\AES_ENC/us01/n587 ), .A2(\AES_ENC/us01/n1058 ), .A3(\AES_ENC/us01/n1059 ), .ZN(\AES_ENC/us01/n815 ) );
NOR4_X2 \AES_ENC/us01/U94  ( .A1(\AES_ENC/us01/n815 ), .A2(\AES_ENC/us01/n814 ), .A3(\AES_ENC/us01/n813 ), .A4(\AES_ENC/us01/n812 ), .ZN(\AES_ENC/us01/n816 ) );
NOR2_X2 \AES_ENC/us01/U93  ( .A1(\AES_ENC/us01/n575 ), .A2(\AES_ENC/us01/n569 ), .ZN(\AES_ENC/us01/n721 ) );
NOR2_X2 \AES_ENC/us01/U92  ( .A1(\AES_ENC/us01/n1031 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n723 ) );
NOR2_X2 \AES_ENC/us01/U91  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n1096 ), .ZN(\AES_ENC/us01/n722 ) );
NOR4_X2 \AES_ENC/us01/U90  ( .A1(\AES_ENC/us01/n724 ), .A2(\AES_ENC/us01/n723 ), .A3(\AES_ENC/us01/n722 ), .A4(\AES_ENC/us01/n721 ), .ZN(\AES_ENC/us01/n725 ) );
NOR2_X2 \AES_ENC/us01/U89  ( .A1(\AES_ENC/us01/n911 ), .A2(\AES_ENC/us01/n990 ), .ZN(\AES_ENC/us01/n1009 ) );
NOR2_X2 \AES_ENC/us01/U88  ( .A1(\AES_ENC/us01/n1013 ), .A2(\AES_ENC/us01/n573 ), .ZN(\AES_ENC/us01/n1014 ) );
NOR2_X2 \AES_ENC/us01/U87  ( .A1(\AES_ENC/us01/n1014 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n1015 ) );
NOR4_X2 \AES_ENC/us01/U86  ( .A1(\AES_ENC/us01/n1016 ), .A2(\AES_ENC/us01/n1015 ), .A3(\AES_ENC/us01/n1119 ), .A4(\AES_ENC/us01/n1046 ), .ZN(\AES_ENC/us01/n1017 ) );
NOR2_X2 \AES_ENC/us01/U81  ( .A1(\AES_ENC/us01/n996 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n998 ) );
NOR2_X2 \AES_ENC/us01/U80  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n618 ), .ZN(\AES_ENC/us01/n1000 ) );
NOR2_X2 \AES_ENC/us01/U79  ( .A1(\AES_ENC/us01/n594 ), .A2(\AES_ENC/us01/n1096 ), .ZN(\AES_ENC/us01/n999 ) );
NOR4_X2 \AES_ENC/us01/U78  ( .A1(\AES_ENC/us01/n1000 ), .A2(\AES_ENC/us01/n999 ), .A3(\AES_ENC/us01/n998 ), .A4(\AES_ENC/us01/n997 ), .ZN(\AES_ENC/us01/n1001 ) );
NOR2_X2 \AES_ENC/us01/U74  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n1096 ), .ZN(\AES_ENC/us01/n697 ) );
NOR2_X2 \AES_ENC/us01/U73  ( .A1(\AES_ENC/us01/n609 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n958 ) );
NOR2_X2 \AES_ENC/us01/U72  ( .A1(\AES_ENC/us01/n911 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n983 ) );
NOR2_X2 \AES_ENC/us01/U71  ( .A1(\AES_ENC/us01/n1054 ), .A2(\AES_ENC/us01/n1103 ), .ZN(\AES_ENC/us01/n1031 ) );
INV_X4 \AES_ENC/us01/U65  ( .A(\AES_ENC/us01/n1050 ), .ZN(\AES_ENC/us01/n582 ) );
INV_X4 \AES_ENC/us01/U64  ( .A(\AES_ENC/us01/n1072 ), .ZN(\AES_ENC/us01/n586 ) );
INV_X4 \AES_ENC/us01/U63  ( .A(\AES_ENC/us01/n1073 ), .ZN(\AES_ENC/us01/n576 ) );
NOR2_X2 \AES_ENC/us01/U62  ( .A1(\AES_ENC/us01/n603 ), .A2(\AES_ENC/us01/n584 ), .ZN(\AES_ENC/us01/n880 ) );
NOR3_X2 \AES_ENC/us01/U61  ( .A1(\AES_ENC/us01/n826 ), .A2(\AES_ENC/us01/n1121 ), .A3(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n946 ) );
INV_X4 \AES_ENC/us01/U59  ( .A(\AES_ENC/us01/n1010 ), .ZN(\AES_ENC/us01/n579 ) );
NOR3_X2 \AES_ENC/us01/U58  ( .A1(\AES_ENC/us01/n573 ), .A2(\AES_ENC/us01/n1029 ), .A3(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n1119 ) );
INV_X4 \AES_ENC/us01/U57  ( .A(\AES_ENC/us01/n956 ), .ZN(\AES_ENC/us01/n580 ) );
NOR2_X2 \AES_ENC/us01/U50  ( .A1(\AES_ENC/us01/n601 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n1013 ) );
NOR2_X2 \AES_ENC/us01/U49  ( .A1(\AES_ENC/us01/n609 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n910 ) );
NOR2_X2 \AES_ENC/us01/U48  ( .A1(\AES_ENC/us01/n569 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n1091 ) );
NOR2_X2 \AES_ENC/us01/U47  ( .A1(\AES_ENC/us01/n614 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n990 ) );
NOR2_X2 \AES_ENC/us01/U46  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/us01/n1121 ), .ZN(\AES_ENC/us01/n996 ) );
NOR2_X2 \AES_ENC/us01/U45  ( .A1(\AES_ENC/us01/n592 ), .A2(\AES_ENC/us01/n622 ), .ZN(\AES_ENC/us01/n628 ) );
NOR2_X2 \AES_ENC/us01/U44  ( .A1(\AES_ENC/us01/n602 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n866 ) );
NOR2_X2 \AES_ENC/us01/U43  ( .A1(\AES_ENC/us01/n610 ), .A2(\AES_ENC/us01/n592 ), .ZN(\AES_ENC/us01/n1006 ) );
NOR2_X2 \AES_ENC/us01/U42  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n1117 ), .ZN(\AES_ENC/us01/n1118 ) );
NOR2_X2 \AES_ENC/us01/U41  ( .A1(\AES_ENC/us01/n1119 ), .A2(\AES_ENC/us01/n1118 ), .ZN(\AES_ENC/us01/n1127 ) );
NOR2_X2 \AES_ENC/us01/U36  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n616 ), .ZN(\AES_ENC/us01/n629 ) );
NOR2_X2 \AES_ENC/us01/U35  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n906 ), .ZN(\AES_ENC/us01/n909 ) );
NOR2_X2 \AES_ENC/us01/U34  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n607 ), .ZN(\AES_ENC/us01/n658 ) );
NOR2_X2 \AES_ENC/us01/U33  ( .A1(\AES_ENC/us01/n1116 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n695 ) );
NOR2_X2 \AES_ENC/us01/U32  ( .A1(\AES_ENC/us01/n1078 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n1083 ) );
NOR2_X2 \AES_ENC/us01/U31  ( .A1(\AES_ENC/us01/n941 ), .A2(\AES_ENC/us01/n579 ), .ZN(\AES_ENC/us01/n724 ) );
NOR2_X2 \AES_ENC/us01/U30  ( .A1(\AES_ENC/us01/n611 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n1107 ) );
NOR2_X2 \AES_ENC/us01/U29  ( .A1(\AES_ENC/us01/n602 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n840 ) );
NOR2_X2 \AES_ENC/us01/U24  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n623 ), .ZN(\AES_ENC/us01/n633 ) );
NOR2_X2 \AES_ENC/us01/U23  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n1080 ), .ZN(\AES_ENC/us01/n1081 ) );
NOR2_X2 \AES_ENC/us01/U21  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n1045 ), .ZN(\AES_ENC/us01/n812 ) );
NOR2_X2 \AES_ENC/us01/U20  ( .A1(\AES_ENC/us01/n1009 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n960 ) );
NOR2_X2 \AES_ENC/us01/U19  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n619 ), .ZN(\AES_ENC/us01/n982 ) );
NOR2_X2 \AES_ENC/us01/U18  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n616 ), .ZN(\AES_ENC/us01/n757 ) );
NOR2_X2 \AES_ENC/us01/U17  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n598 ), .ZN(\AES_ENC/us01/n698 ) );
NOR2_X2 \AES_ENC/us01/U16  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n605 ), .ZN(\AES_ENC/us01/n708 ) );
NOR2_X2 \AES_ENC/us01/U15  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n603 ), .ZN(\AES_ENC/us01/n770 ) );
NOR2_X2 \AES_ENC/us01/U10  ( .A1(\AES_ENC/us01/n605 ), .A2(\AES_ENC/us01/n576 ), .ZN(\AES_ENC/us01/n803 ) );
NOR2_X2 \AES_ENC/us01/U9  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n881 ), .ZN(\AES_ENC/us01/n711 ) );
NOR2_X2 \AES_ENC/us01/U8  ( .A1(\AES_ENC/us01/n580 ), .A2(\AES_ENC/us01/n603 ), .ZN(\AES_ENC/us01/n867 ) );
NOR2_X2 \AES_ENC/us01/U7  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n615 ), .ZN(\AES_ENC/us01/n804 ) );
NOR2_X2 \AES_ENC/us01/U6  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n609 ), .ZN(\AES_ENC/us01/n1046 ) );
OR2_X4 \AES_ENC/us01/U5  ( .A1(\AES_ENC/us01/n612 ), .A2(\AES_ENC/sa01 [1]),.ZN(\AES_ENC/us01/n570 ) );
OR2_X4 \AES_ENC/us01/U4  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/sa01 [4]),.ZN(\AES_ENC/us01/n569 ) );
NAND2_X2 \AES_ENC/us01/U514  ( .A1(\AES_ENC/us01/n1121 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n1030 ) );
AND2_X2 \AES_ENC/us01/U513  ( .A1(\AES_ENC/us01/n607 ), .A2(\AES_ENC/us01/n1030 ), .ZN(\AES_ENC/us01/n1049 ) );
NAND2_X2 \AES_ENC/us01/U511  ( .A1(\AES_ENC/us01/n1049 ), .A2(\AES_ENC/us01/n794 ), .ZN(\AES_ENC/us01/n637 ) );
AND2_X2 \AES_ENC/us01/U493  ( .A1(\AES_ENC/us01/n779 ), .A2(\AES_ENC/us01/n996 ), .ZN(\AES_ENC/us01/n632 ) );
NAND4_X2 \AES_ENC/us01/U485  ( .A1(\AES_ENC/us01/n637 ), .A2(\AES_ENC/us01/n636 ), .A3(\AES_ENC/us01/n635 ), .A4(\AES_ENC/us01/n634 ), .ZN(\AES_ENC/us01/n638 ) );
NAND2_X2 \AES_ENC/us01/U484  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n638 ), .ZN(\AES_ENC/us01/n679 ) );
NAND2_X2 \AES_ENC/us01/U481  ( .A1(\AES_ENC/us01/n1094 ), .A2(\AES_ENC/us01/n613 ), .ZN(\AES_ENC/us01/n648 ) );
NAND2_X2 \AES_ENC/us01/U476  ( .A1(\AES_ENC/us01/n619 ), .A2(\AES_ENC/us01/n598 ), .ZN(\AES_ENC/us01/n762 ) );
NAND2_X2 \AES_ENC/us01/U475  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n762 ), .ZN(\AES_ENC/us01/n647 ) );
NAND4_X2 \AES_ENC/us01/U457  ( .A1(\AES_ENC/us01/n648 ), .A2(\AES_ENC/us01/n647 ), .A3(\AES_ENC/us01/n646 ), .A4(\AES_ENC/us01/n645 ), .ZN(\AES_ENC/us01/n649 ) );
NAND2_X2 \AES_ENC/us01/U456  ( .A1(\AES_ENC/sa01 [0]), .A2(\AES_ENC/us01/n649 ), .ZN(\AES_ENC/us01/n665 ) );
NAND2_X2 \AES_ENC/us01/U454  ( .A1(\AES_ENC/us01/n626 ), .A2(\AES_ENC/us01/n601 ), .ZN(\AES_ENC/us01/n855 ) );
NAND2_X2 \AES_ENC/us01/U453  ( .A1(\AES_ENC/us01/n617 ), .A2(\AES_ENC/us01/n855 ), .ZN(\AES_ENC/us01/n821 ) );
NAND2_X2 \AES_ENC/us01/U452  ( .A1(\AES_ENC/us01/n1093 ), .A2(\AES_ENC/us01/n821 ), .ZN(\AES_ENC/us01/n662 ) );
NAND2_X2 \AES_ENC/us01/U451  ( .A1(\AES_ENC/us01/n605 ), .A2(\AES_ENC/us01/n620 ), .ZN(\AES_ENC/us01/n650 ) );
NAND2_X2 \AES_ENC/us01/U450  ( .A1(\AES_ENC/us01/n956 ), .A2(\AES_ENC/us01/n650 ), .ZN(\AES_ENC/us01/n661 ) );
NAND2_X2 \AES_ENC/us01/U449  ( .A1(\AES_ENC/us01/n596 ), .A2(\AES_ENC/us01/n581 ), .ZN(\AES_ENC/us01/n839 ) );
OR2_X2 \AES_ENC/us01/U446  ( .A1(\AES_ENC/us01/n839 ), .A2(\AES_ENC/us01/n932 ), .ZN(\AES_ENC/us01/n656 ) );
NAND2_X2 \AES_ENC/us01/U445  ( .A1(\AES_ENC/us01/n624 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n1096 ) );
NAND2_X2 \AES_ENC/us01/U444  ( .A1(\AES_ENC/us01/n1030 ), .A2(\AES_ENC/us01/n1096 ), .ZN(\AES_ENC/us01/n651 ) );
NAND2_X2 \AES_ENC/us01/U443  ( .A1(\AES_ENC/us01/n1114 ), .A2(\AES_ENC/us01/n651 ), .ZN(\AES_ENC/us01/n655 ) );
OR3_X2 \AES_ENC/us01/U440  ( .A1(\AES_ENC/us01/n1079 ), .A2(\AES_ENC/sa01 [7]), .A3(\AES_ENC/us01/n596 ), .ZN(\AES_ENC/us01/n654 ));
NAND2_X2 \AES_ENC/us01/U439  ( .A1(\AES_ENC/us01/n623 ), .A2(\AES_ENC/us01/n619 ), .ZN(\AES_ENC/us01/n652 ) );
NAND4_X2 \AES_ENC/us01/U437  ( .A1(\AES_ENC/us01/n656 ), .A2(\AES_ENC/us01/n655 ), .A3(\AES_ENC/us01/n654 ), .A4(\AES_ENC/us01/n653 ), .ZN(\AES_ENC/us01/n657 ) );
NAND2_X2 \AES_ENC/us01/U436  ( .A1(\AES_ENC/sa01 [2]), .A2(\AES_ENC/us01/n657 ), .ZN(\AES_ENC/us01/n660 ) );
NAND4_X2 \AES_ENC/us01/U432  ( .A1(\AES_ENC/us01/n662 ), .A2(\AES_ENC/us01/n661 ), .A3(\AES_ENC/us01/n660 ), .A4(\AES_ENC/us01/n659 ), .ZN(\AES_ENC/us01/n663 ) );
NAND2_X2 \AES_ENC/us01/U431  ( .A1(\AES_ENC/us01/n663 ), .A2(\AES_ENC/us01/n627 ), .ZN(\AES_ENC/us01/n664 ) );
NAND2_X2 \AES_ENC/us01/U430  ( .A1(\AES_ENC/us01/n665 ), .A2(\AES_ENC/us01/n664 ), .ZN(\AES_ENC/us01/n666 ) );
NAND2_X2 \AES_ENC/us01/U429  ( .A1(\AES_ENC/sa01 [6]), .A2(\AES_ENC/us01/n666 ), .ZN(\AES_ENC/us01/n678 ) );
NAND2_X2 \AES_ENC/us01/U426  ( .A1(\AES_ENC/us01/n735 ), .A2(\AES_ENC/us01/n1093 ), .ZN(\AES_ENC/us01/n675 ) );
NAND2_X2 \AES_ENC/us01/U425  ( .A1(\AES_ENC/us01/n625 ), .A2(\AES_ENC/us01/n607 ), .ZN(\AES_ENC/us01/n1045 ) );
OR2_X2 \AES_ENC/us01/U424  ( .A1(\AES_ENC/us01/n1045 ), .A2(\AES_ENC/us01/n586 ), .ZN(\AES_ENC/us01/n674 ) );
NAND2_X2 \AES_ENC/us01/U423  ( .A1(\AES_ENC/sa01 [1]), .A2(\AES_ENC/us01/n609 ), .ZN(\AES_ENC/us01/n667 ) );
NAND2_X2 \AES_ENC/us01/U422  ( .A1(\AES_ENC/us01/n605 ), .A2(\AES_ENC/us01/n667 ), .ZN(\AES_ENC/us01/n1071 ) );
NAND4_X2 \AES_ENC/us01/U412  ( .A1(\AES_ENC/us01/n675 ), .A2(\AES_ENC/us01/n674 ), .A3(\AES_ENC/us01/n673 ), .A4(\AES_ENC/us01/n672 ), .ZN(\AES_ENC/us01/n676 ) );
NAND2_X2 \AES_ENC/us01/U411  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n676 ), .ZN(\AES_ENC/us01/n677 ) );
NAND2_X2 \AES_ENC/us01/U408  ( .A1(\AES_ENC/us01/n800 ), .A2(\AES_ENC/us01/n1022 ), .ZN(\AES_ENC/us01/n680 ) );
NAND2_X2 \AES_ENC/us01/U407  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n680 ), .ZN(\AES_ENC/us01/n681 ) );
AND2_X2 \AES_ENC/us01/U402  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n684 ), .ZN(\AES_ENC/us01/n682 ) );
NAND4_X2 \AES_ENC/us01/U395  ( .A1(\AES_ENC/us01/n691 ), .A2(\AES_ENC/us01/n583 ), .A3(\AES_ENC/us01/n690 ), .A4(\AES_ENC/us01/n689 ), .ZN(\AES_ENC/us01/n692 ) );
NAND2_X2 \AES_ENC/us01/U394  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n692 ), .ZN(\AES_ENC/us01/n733 ) );
NAND2_X2 \AES_ENC/us01/U392  ( .A1(\AES_ENC/us01/n977 ), .A2(\AES_ENC/us01/n1050 ), .ZN(\AES_ENC/us01/n702 ) );
NAND2_X2 \AES_ENC/us01/U391  ( .A1(\AES_ENC/us01/n1093 ), .A2(\AES_ENC/us01/n1045 ), .ZN(\AES_ENC/us01/n701 ) );
NAND4_X2 \AES_ENC/us01/U381  ( .A1(\AES_ENC/us01/n702 ), .A2(\AES_ENC/us01/n701 ), .A3(\AES_ENC/us01/n700 ), .A4(\AES_ENC/us01/n699 ), .ZN(\AES_ENC/us01/n703 ) );
NAND2_X2 \AES_ENC/us01/U380  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n703 ), .ZN(\AES_ENC/us01/n732 ) );
AND2_X2 \AES_ENC/us01/U379  ( .A1(\AES_ENC/sa01 [0]), .A2(\AES_ENC/sa01 [6]),.ZN(\AES_ENC/us01/n1113 ) );
NAND2_X2 \AES_ENC/us01/U378  ( .A1(\AES_ENC/us01/n619 ), .A2(\AES_ENC/us01/n1030 ), .ZN(\AES_ENC/us01/n881 ) );
NAND2_X2 \AES_ENC/us01/U377  ( .A1(\AES_ENC/us01/n1093 ), .A2(\AES_ENC/us01/n881 ), .ZN(\AES_ENC/us01/n715 ) );
NAND2_X2 \AES_ENC/us01/U376  ( .A1(\AES_ENC/us01/n1010 ), .A2(\AES_ENC/us01/n622 ), .ZN(\AES_ENC/us01/n714 ) );
NAND2_X2 \AES_ENC/us01/U375  ( .A1(\AES_ENC/us01/n855 ), .A2(\AES_ENC/us01/n625 ), .ZN(\AES_ENC/us01/n1117 ) );
XNOR2_X2 \AES_ENC/us01/U371  ( .A(\AES_ENC/us01/n593 ), .B(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n824 ) );
NAND4_X2 \AES_ENC/us01/U362  ( .A1(\AES_ENC/us01/n715 ), .A2(\AES_ENC/us01/n714 ), .A3(\AES_ENC/us01/n713 ), .A4(\AES_ENC/us01/n712 ), .ZN(\AES_ENC/us01/n716 ) );
NAND2_X2 \AES_ENC/us01/U361  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n716 ), .ZN(\AES_ENC/us01/n731 ) );
AND2_X2 \AES_ENC/us01/U360  ( .A1(\AES_ENC/sa01 [6]), .A2(\AES_ENC/us01/n627 ), .ZN(\AES_ENC/us01/n1131 ) );
NAND2_X2 \AES_ENC/us01/U359  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n717 ) );
NAND2_X2 \AES_ENC/us01/U358  ( .A1(\AES_ENC/us01/n1029 ), .A2(\AES_ENC/us01/n717 ), .ZN(\AES_ENC/us01/n728 ) );
NAND2_X2 \AES_ENC/us01/U357  ( .A1(\AES_ENC/sa01 [1]), .A2(\AES_ENC/us01/n612 ), .ZN(\AES_ENC/us01/n1097 ) );
NAND2_X2 \AES_ENC/us01/U356  ( .A1(\AES_ENC/us01/n610 ), .A2(\AES_ENC/us01/n1097 ), .ZN(\AES_ENC/us01/n718 ) );
NAND2_X2 \AES_ENC/us01/U355  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n718 ), .ZN(\AES_ENC/us01/n727 ) );
NAND4_X2 \AES_ENC/us01/U344  ( .A1(\AES_ENC/us01/n728 ), .A2(\AES_ENC/us01/n727 ), .A3(\AES_ENC/us01/n726 ), .A4(\AES_ENC/us01/n725 ), .ZN(\AES_ENC/us01/n729 ) );
NAND2_X2 \AES_ENC/us01/U343  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n729 ), .ZN(\AES_ENC/us01/n730 ) );
NAND4_X2 \AES_ENC/us01/U342  ( .A1(\AES_ENC/us01/n733 ), .A2(\AES_ENC/us01/n732 ), .A3(\AES_ENC/us01/n731 ), .A4(\AES_ENC/us01/n730 ), .ZN(\AES_ENC/sa01_sub[1] ) );
NAND2_X2 \AES_ENC/us01/U341  ( .A1(\AES_ENC/sa01 [7]), .A2(\AES_ENC/us01/n593 ), .ZN(\AES_ENC/us01/n734 ) );
NAND2_X2 \AES_ENC/us01/U340  ( .A1(\AES_ENC/us01/n734 ), .A2(\AES_ENC/us01/n588 ), .ZN(\AES_ENC/us01/n738 ) );
OR4_X2 \AES_ENC/us01/U339  ( .A1(\AES_ENC/us01/n738 ), .A2(\AES_ENC/us01/n596 ), .A3(\AES_ENC/us01/n826 ), .A4(\AES_ENC/us01/n1121 ), .ZN(\AES_ENC/us01/n746 ) );
NAND2_X2 \AES_ENC/us01/U337  ( .A1(\AES_ENC/us01/n1100 ), .A2(\AES_ENC/us01/n617 ), .ZN(\AES_ENC/us01/n992 ) );
OR2_X2 \AES_ENC/us01/U336  ( .A1(\AES_ENC/us01/n592 ), .A2(\AES_ENC/us01/n735 ), .ZN(\AES_ENC/us01/n737 ) );
NAND2_X2 \AES_ENC/us01/U334  ( .A1(\AES_ENC/us01/n605 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n753 ) );
NAND2_X2 \AES_ENC/us01/U333  ( .A1(\AES_ENC/us01/n603 ), .A2(\AES_ENC/us01/n753 ), .ZN(\AES_ENC/us01/n1080 ) );
NAND2_X2 \AES_ENC/us01/U332  ( .A1(\AES_ENC/us01/n1048 ), .A2(\AES_ENC/us01/n602 ), .ZN(\AES_ENC/us01/n736 ) );
NAND2_X2 \AES_ENC/us01/U331  ( .A1(\AES_ENC/us01/n737 ), .A2(\AES_ENC/us01/n736 ), .ZN(\AES_ENC/us01/n739 ) );
NAND2_X2 \AES_ENC/us01/U330  ( .A1(\AES_ENC/us01/n739 ), .A2(\AES_ENC/us01/n738 ), .ZN(\AES_ENC/us01/n745 ) );
NAND2_X2 \AES_ENC/us01/U326  ( .A1(\AES_ENC/us01/n1096 ), .A2(\AES_ENC/us01/n598 ), .ZN(\AES_ENC/us01/n906 ) );
NAND4_X2 \AES_ENC/us01/U323  ( .A1(\AES_ENC/us01/n746 ), .A2(\AES_ENC/us01/n992 ), .A3(\AES_ENC/us01/n745 ), .A4(\AES_ENC/us01/n744 ), .ZN(\AES_ENC/us01/n747 ) );
NAND2_X2 \AES_ENC/us01/U322  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n747 ), .ZN(\AES_ENC/us01/n793 ) );
NAND2_X2 \AES_ENC/us01/U321  ( .A1(\AES_ENC/us01/n606 ), .A2(\AES_ENC/us01/n855 ), .ZN(\AES_ENC/us01/n748 ) );
NAND2_X2 \AES_ENC/us01/U320  ( .A1(\AES_ENC/us01/n956 ), .A2(\AES_ENC/us01/n748 ), .ZN(\AES_ENC/us01/n760 ) );
NAND2_X2 \AES_ENC/us01/U313  ( .A1(\AES_ENC/us01/n598 ), .A2(\AES_ENC/us01/n753 ), .ZN(\AES_ENC/us01/n1023 ) );
NAND4_X2 \AES_ENC/us01/U308  ( .A1(\AES_ENC/us01/n760 ), .A2(\AES_ENC/us01/n992 ), .A3(\AES_ENC/us01/n759 ), .A4(\AES_ENC/us01/n758 ), .ZN(\AES_ENC/us01/n761 ) );
NAND2_X2 \AES_ENC/us01/U307  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n761 ), .ZN(\AES_ENC/us01/n792 ) );
NAND2_X2 \AES_ENC/us01/U306  ( .A1(\AES_ENC/us01/n606 ), .A2(\AES_ENC/us01/n610 ), .ZN(\AES_ENC/us01/n989 ) );
NAND2_X2 \AES_ENC/us01/U305  ( .A1(\AES_ENC/us01/n1050 ), .A2(\AES_ENC/us01/n989 ), .ZN(\AES_ENC/us01/n777 ) );
NAND2_X2 \AES_ENC/us01/U304  ( .A1(\AES_ENC/us01/n1093 ), .A2(\AES_ENC/us01/n762 ), .ZN(\AES_ENC/us01/n776 ) );
XNOR2_X2 \AES_ENC/us01/U301  ( .A(\AES_ENC/sa01 [7]), .B(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n959 ) );
NAND4_X2 \AES_ENC/us01/U289  ( .A1(\AES_ENC/us01/n777 ), .A2(\AES_ENC/us01/n776 ), .A3(\AES_ENC/us01/n775 ), .A4(\AES_ENC/us01/n774 ), .ZN(\AES_ENC/us01/n778 ) );
NAND2_X2 \AES_ENC/us01/U288  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n778 ), .ZN(\AES_ENC/us01/n791 ) );
NAND2_X2 \AES_ENC/us01/U287  ( .A1(\AES_ENC/us01/n1056 ), .A2(\AES_ENC/us01/n1050 ), .ZN(\AES_ENC/us01/n788 ) );
NAND2_X2 \AES_ENC/us01/U286  ( .A1(\AES_ENC/us01/n1091 ), .A2(\AES_ENC/us01/n779 ), .ZN(\AES_ENC/us01/n787 ) );
NAND2_X2 \AES_ENC/us01/U285  ( .A1(\AES_ENC/us01/n956 ), .A2(\AES_ENC/sa01 [1]), .ZN(\AES_ENC/us01/n786 ) );
NAND4_X2 \AES_ENC/us01/U278  ( .A1(\AES_ENC/us01/n788 ), .A2(\AES_ENC/us01/n787 ), .A3(\AES_ENC/us01/n786 ), .A4(\AES_ENC/us01/n785 ), .ZN(\AES_ENC/us01/n789 ) );
NAND2_X2 \AES_ENC/us01/U277  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n789 ), .ZN(\AES_ENC/us01/n790 ) );
NAND4_X2 \AES_ENC/us01/U276  ( .A1(\AES_ENC/us01/n793 ), .A2(\AES_ENC/us01/n792 ), .A3(\AES_ENC/us01/n791 ), .A4(\AES_ENC/us01/n790 ), .ZN(\AES_ENC/sa01_sub[2] ) );
NAND2_X2 \AES_ENC/us01/U275  ( .A1(\AES_ENC/us01/n1059 ), .A2(\AES_ENC/us01/n794 ), .ZN(\AES_ENC/us01/n810 ) );
NAND2_X2 \AES_ENC/us01/U274  ( .A1(\AES_ENC/us01/n1049 ), .A2(\AES_ENC/us01/n956 ), .ZN(\AES_ENC/us01/n809 ) );
OR2_X2 \AES_ENC/us01/U266  ( .A1(\AES_ENC/us01/n1096 ), .A2(\AES_ENC/us01/n587 ), .ZN(\AES_ENC/us01/n802 ) );
NAND2_X2 \AES_ENC/us01/U265  ( .A1(\AES_ENC/us01/n1053 ), .A2(\AES_ENC/us01/n800 ), .ZN(\AES_ENC/us01/n801 ) );
NAND2_X2 \AES_ENC/us01/U264  ( .A1(\AES_ENC/us01/n802 ), .A2(\AES_ENC/us01/n801 ), .ZN(\AES_ENC/us01/n805 ) );
NAND4_X2 \AES_ENC/us01/U261  ( .A1(\AES_ENC/us01/n810 ), .A2(\AES_ENC/us01/n809 ), .A3(\AES_ENC/us01/n808 ), .A4(\AES_ENC/us01/n807 ), .ZN(\AES_ENC/us01/n811 ) );
NAND2_X2 \AES_ENC/us01/U260  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n811 ), .ZN(\AES_ENC/us01/n852 ) );
OR2_X2 \AES_ENC/us01/U259  ( .A1(\AES_ENC/us01/n1023 ), .A2(\AES_ENC/us01/n575 ), .ZN(\AES_ENC/us01/n819 ) );
OR2_X2 \AES_ENC/us01/U257  ( .A1(\AES_ENC/us01/n570 ), .A2(\AES_ENC/us01/n930 ), .ZN(\AES_ENC/us01/n818 ) );
NAND2_X2 \AES_ENC/us01/U256  ( .A1(\AES_ENC/us01/n1013 ), .A2(\AES_ENC/us01/n1094 ), .ZN(\AES_ENC/us01/n817 ) );
NAND4_X2 \AES_ENC/us01/U249  ( .A1(\AES_ENC/us01/n819 ), .A2(\AES_ENC/us01/n818 ), .A3(\AES_ENC/us01/n817 ), .A4(\AES_ENC/us01/n816 ), .ZN(\AES_ENC/us01/n820 ) );
NAND2_X2 \AES_ENC/us01/U248  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n820 ), .ZN(\AES_ENC/us01/n851 ) );
NAND2_X2 \AES_ENC/us01/U247  ( .A1(\AES_ENC/us01/n956 ), .A2(\AES_ENC/us01/n1080 ), .ZN(\AES_ENC/us01/n835 ) );
NAND2_X2 \AES_ENC/us01/U246  ( .A1(\AES_ENC/us01/n570 ), .A2(\AES_ENC/us01/n1030 ), .ZN(\AES_ENC/us01/n1047 ) );
OR2_X2 \AES_ENC/us01/U245  ( .A1(\AES_ENC/us01/n1047 ), .A2(\AES_ENC/us01/n582 ), .ZN(\AES_ENC/us01/n834 ) );
NAND2_X2 \AES_ENC/us01/U244  ( .A1(\AES_ENC/us01/n1072 ), .A2(\AES_ENC/us01/n620 ), .ZN(\AES_ENC/us01/n833 ) );
NAND4_X2 \AES_ENC/us01/U233  ( .A1(\AES_ENC/us01/n835 ), .A2(\AES_ENC/us01/n834 ), .A3(\AES_ENC/us01/n833 ), .A4(\AES_ENC/us01/n832 ), .ZN(\AES_ENC/us01/n836 ) );
NAND2_X2 \AES_ENC/us01/U232  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n836 ), .ZN(\AES_ENC/us01/n850 ) );
NAND2_X2 \AES_ENC/us01/U231  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n601 ), .ZN(\AES_ENC/us01/n847 ) );
NAND2_X2 \AES_ENC/us01/U230  ( .A1(\AES_ENC/us01/n1050 ), .A2(\AES_ENC/us01/n1071 ), .ZN(\AES_ENC/us01/n846 ) );
OR2_X2 \AES_ENC/us01/U224  ( .A1(\AES_ENC/us01/n1053 ), .A2(\AES_ENC/us01/n911 ), .ZN(\AES_ENC/us01/n1077 ) );
NAND4_X2 \AES_ENC/us01/U220  ( .A1(\AES_ENC/us01/n847 ), .A2(\AES_ENC/us01/n846 ), .A3(\AES_ENC/us01/n845 ), .A4(\AES_ENC/us01/n844 ), .ZN(\AES_ENC/us01/n848 ) );
NAND2_X2 \AES_ENC/us01/U219  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n848 ), .ZN(\AES_ENC/us01/n849 ) );
NAND4_X2 \AES_ENC/us01/U218  ( .A1(\AES_ENC/us01/n852 ), .A2(\AES_ENC/us01/n851 ), .A3(\AES_ENC/us01/n850 ), .A4(\AES_ENC/us01/n849 ), .ZN(\AES_ENC/sa01_sub[3] ) );
NAND2_X2 \AES_ENC/us01/U216  ( .A1(\AES_ENC/us01/n1009 ), .A2(\AES_ENC/us01/n1072 ), .ZN(\AES_ENC/us01/n862 ) );
NAND2_X2 \AES_ENC/us01/U215  ( .A1(\AES_ENC/us01/n610 ), .A2(\AES_ENC/us01/n618 ), .ZN(\AES_ENC/us01/n853 ) );
NAND2_X2 \AES_ENC/us01/U214  ( .A1(\AES_ENC/us01/n1050 ), .A2(\AES_ENC/us01/n853 ), .ZN(\AES_ENC/us01/n861 ) );
NAND4_X2 \AES_ENC/us01/U206  ( .A1(\AES_ENC/us01/n862 ), .A2(\AES_ENC/us01/n861 ), .A3(\AES_ENC/us01/n860 ), .A4(\AES_ENC/us01/n859 ), .ZN(\AES_ENC/us01/n863 ) );
NAND2_X2 \AES_ENC/us01/U205  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n863 ), .ZN(\AES_ENC/us01/n905 ) );
NAND2_X2 \AES_ENC/us01/U204  ( .A1(\AES_ENC/us01/n1010 ), .A2(\AES_ENC/us01/n989 ), .ZN(\AES_ENC/us01/n874 ) );
NAND2_X2 \AES_ENC/us01/U203  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n592 ), .ZN(\AES_ENC/us01/n864 ) );
NAND2_X2 \AES_ENC/us01/U202  ( .A1(\AES_ENC/us01/n929 ), .A2(\AES_ENC/us01/n864 ), .ZN(\AES_ENC/us01/n873 ) );
NAND4_X2 \AES_ENC/us01/U193  ( .A1(\AES_ENC/us01/n874 ), .A2(\AES_ENC/us01/n873 ), .A3(\AES_ENC/us01/n872 ), .A4(\AES_ENC/us01/n871 ), .ZN(\AES_ENC/us01/n875 ) );
NAND2_X2 \AES_ENC/us01/U192  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n875 ), .ZN(\AES_ENC/us01/n904 ) );
NAND2_X2 \AES_ENC/us01/U191  ( .A1(\AES_ENC/us01/n597 ), .A2(\AES_ENC/us01/n1050 ), .ZN(\AES_ENC/us01/n889 ) );
NAND2_X2 \AES_ENC/us01/U190  ( .A1(\AES_ENC/us01/n1093 ), .A2(\AES_ENC/us01/n617 ), .ZN(\AES_ENC/us01/n876 ) );
NAND2_X2 \AES_ENC/us01/U189  ( .A1(\AES_ENC/us01/n576 ), .A2(\AES_ENC/us01/n876 ), .ZN(\AES_ENC/us01/n877 ) );
NAND2_X2 \AES_ENC/us01/U188  ( .A1(\AES_ENC/us01/n877 ), .A2(\AES_ENC/us01/n601 ), .ZN(\AES_ENC/us01/n888 ) );
NAND4_X2 \AES_ENC/us01/U179  ( .A1(\AES_ENC/us01/n889 ), .A2(\AES_ENC/us01/n888 ), .A3(\AES_ENC/us01/n887 ), .A4(\AES_ENC/us01/n886 ), .ZN(\AES_ENC/us01/n890 ) );
NAND2_X2 \AES_ENC/us01/U178  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n890 ), .ZN(\AES_ENC/us01/n903 ) );
OR2_X2 \AES_ENC/us01/U177  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n1059 ), .ZN(\AES_ENC/us01/n900 ) );
NAND2_X2 \AES_ENC/us01/U176  ( .A1(\AES_ENC/us01/n1073 ), .A2(\AES_ENC/us01/n1047 ), .ZN(\AES_ENC/us01/n899 ) );
NAND2_X2 \AES_ENC/us01/U175  ( .A1(\AES_ENC/us01/n1094 ), .A2(\AES_ENC/us01/n608 ), .ZN(\AES_ENC/us01/n898 ) );
NAND4_X2 \AES_ENC/us01/U167  ( .A1(\AES_ENC/us01/n900 ), .A2(\AES_ENC/us01/n899 ), .A3(\AES_ENC/us01/n898 ), .A4(\AES_ENC/us01/n897 ), .ZN(\AES_ENC/us01/n901 ) );
NAND2_X2 \AES_ENC/us01/U166  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n901 ), .ZN(\AES_ENC/us01/n902 ) );
NAND4_X2 \AES_ENC/us01/U165  ( .A1(\AES_ENC/us01/n905 ), .A2(\AES_ENC/us01/n904 ), .A3(\AES_ENC/us01/n903 ), .A4(\AES_ENC/us01/n902 ), .ZN(\AES_ENC/sa01_sub[4] ) );
NAND2_X2 \AES_ENC/us01/U164  ( .A1(\AES_ENC/us01/n1094 ), .A2(\AES_ENC/us01/n615 ), .ZN(\AES_ENC/us01/n922 ) );
NAND2_X2 \AES_ENC/us01/U163  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n989 ), .ZN(\AES_ENC/us01/n921 ) );
NAND4_X2 \AES_ENC/us01/U151  ( .A1(\AES_ENC/us01/n922 ), .A2(\AES_ENC/us01/n921 ), .A3(\AES_ENC/us01/n920 ), .A4(\AES_ENC/us01/n919 ), .ZN(\AES_ENC/us01/n923 ) );
NAND2_X2 \AES_ENC/us01/U150  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n923 ), .ZN(\AES_ENC/us01/n972 ) );
NAND2_X2 \AES_ENC/us01/U149  ( .A1(\AES_ENC/us01/n603 ), .A2(\AES_ENC/us01/n605 ), .ZN(\AES_ENC/us01/n924 ) );
NAND2_X2 \AES_ENC/us01/U148  ( .A1(\AES_ENC/us01/n1073 ), .A2(\AES_ENC/us01/n924 ), .ZN(\AES_ENC/us01/n939 ) );
NAND2_X2 \AES_ENC/us01/U147  ( .A1(\AES_ENC/us01/n926 ), .A2(\AES_ENC/us01/n925 ), .ZN(\AES_ENC/us01/n927 ) );
NAND2_X2 \AES_ENC/us01/U146  ( .A1(\AES_ENC/us01/n587 ), .A2(\AES_ENC/us01/n927 ), .ZN(\AES_ENC/us01/n928 ) );
NAND2_X2 \AES_ENC/us01/U145  ( .A1(\AES_ENC/us01/n928 ), .A2(\AES_ENC/us01/n1080 ), .ZN(\AES_ENC/us01/n938 ) );
OR2_X2 \AES_ENC/us01/U144  ( .A1(\AES_ENC/us01/n1117 ), .A2(\AES_ENC/us01/n580 ), .ZN(\AES_ENC/us01/n937 ) );
NAND4_X2 \AES_ENC/us01/U139  ( .A1(\AES_ENC/us01/n939 ), .A2(\AES_ENC/us01/n938 ), .A3(\AES_ENC/us01/n937 ), .A4(\AES_ENC/us01/n936 ), .ZN(\AES_ENC/us01/n940 ) );
NAND2_X2 \AES_ENC/us01/U138  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n940 ), .ZN(\AES_ENC/us01/n971 ) );
OR2_X2 \AES_ENC/us01/U137  ( .A1(\AES_ENC/us01/n586 ), .A2(\AES_ENC/us01/n941 ), .ZN(\AES_ENC/us01/n954 ) );
NAND2_X2 \AES_ENC/us01/U136  ( .A1(\AES_ENC/us01/n1096 ), .A2(\AES_ENC/us01/n618 ), .ZN(\AES_ENC/us01/n942 ) );
NAND2_X2 \AES_ENC/us01/U135  ( .A1(\AES_ENC/us01/n1048 ), .A2(\AES_ENC/us01/n942 ), .ZN(\AES_ENC/us01/n943 ) );
NAND2_X2 \AES_ENC/us01/U134  ( .A1(\AES_ENC/us01/n582 ), .A2(\AES_ENC/us01/n943 ), .ZN(\AES_ENC/us01/n944 ) );
NAND2_X2 \AES_ENC/us01/U133  ( .A1(\AES_ENC/us01/n944 ), .A2(\AES_ENC/us01/n599 ), .ZN(\AES_ENC/us01/n953 ) );
NAND4_X2 \AES_ENC/us01/U125  ( .A1(\AES_ENC/us01/n954 ), .A2(\AES_ENC/us01/n953 ), .A3(\AES_ENC/us01/n952 ), .A4(\AES_ENC/us01/n951 ), .ZN(\AES_ENC/us01/n955 ) );
NAND2_X2 \AES_ENC/us01/U124  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n955 ), .ZN(\AES_ENC/us01/n970 ) );
NAND2_X2 \AES_ENC/us01/U123  ( .A1(\AES_ENC/us01/n1094 ), .A2(\AES_ENC/us01/n1071 ), .ZN(\AES_ENC/us01/n967 ) );
NAND2_X2 \AES_ENC/us01/U122  ( .A1(\AES_ENC/us01/n956 ), .A2(\AES_ENC/us01/n1030 ), .ZN(\AES_ENC/us01/n966 ) );
NAND4_X2 \AES_ENC/us01/U114  ( .A1(\AES_ENC/us01/n967 ), .A2(\AES_ENC/us01/n966 ), .A3(\AES_ENC/us01/n965 ), .A4(\AES_ENC/us01/n964 ), .ZN(\AES_ENC/us01/n968 ) );
NAND2_X2 \AES_ENC/us01/U113  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n968 ), .ZN(\AES_ENC/us01/n969 ) );
NAND4_X2 \AES_ENC/us01/U112  ( .A1(\AES_ENC/us01/n972 ), .A2(\AES_ENC/us01/n971 ), .A3(\AES_ENC/us01/n970 ), .A4(\AES_ENC/us01/n969 ), .ZN(\AES_ENC/sa01_sub[5] ) );
NAND2_X2 \AES_ENC/us01/U111  ( .A1(\AES_ENC/us01/n570 ), .A2(\AES_ENC/us01/n1097 ), .ZN(\AES_ENC/us01/n973 ) );
NAND2_X2 \AES_ENC/us01/U110  ( .A1(\AES_ENC/us01/n1073 ), .A2(\AES_ENC/us01/n973 ), .ZN(\AES_ENC/us01/n987 ) );
NAND2_X2 \AES_ENC/us01/U109  ( .A1(\AES_ENC/us01/n974 ), .A2(\AES_ENC/us01/n1077 ), .ZN(\AES_ENC/us01/n975 ) );
NAND2_X2 \AES_ENC/us01/U108  ( .A1(\AES_ENC/us01/n584 ), .A2(\AES_ENC/us01/n975 ), .ZN(\AES_ENC/us01/n976 ) );
NAND2_X2 \AES_ENC/us01/U107  ( .A1(\AES_ENC/us01/n977 ), .A2(\AES_ENC/us01/n976 ), .ZN(\AES_ENC/us01/n986 ) );
NAND4_X2 \AES_ENC/us01/U99  ( .A1(\AES_ENC/us01/n987 ), .A2(\AES_ENC/us01/n986 ), .A3(\AES_ENC/us01/n985 ), .A4(\AES_ENC/us01/n984 ), .ZN(\AES_ENC/us01/n988 ) );
NAND2_X2 \AES_ENC/us01/U98  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n988 ), .ZN(\AES_ENC/us01/n1044 ) );
NAND2_X2 \AES_ENC/us01/U97  ( .A1(\AES_ENC/us01/n1073 ), .A2(\AES_ENC/us01/n989 ), .ZN(\AES_ENC/us01/n1004 ) );
NAND2_X2 \AES_ENC/us01/U96  ( .A1(\AES_ENC/us01/n1092 ), .A2(\AES_ENC/us01/n605 ), .ZN(\AES_ENC/us01/n1003 ) );
NAND4_X2 \AES_ENC/us01/U85  ( .A1(\AES_ENC/us01/n1004 ), .A2(\AES_ENC/us01/n1003 ), .A3(\AES_ENC/us01/n1002 ), .A4(\AES_ENC/us01/n1001 ), .ZN(\AES_ENC/us01/n1005 ) );
NAND2_X2 \AES_ENC/us01/U84  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n1005 ), .ZN(\AES_ENC/us01/n1043 ) );
NAND2_X2 \AES_ENC/us01/U83  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n626 ), .ZN(\AES_ENC/us01/n1020 ) );
NAND2_X2 \AES_ENC/us01/U82  ( .A1(\AES_ENC/us01/n1050 ), .A2(\AES_ENC/us01/n612 ), .ZN(\AES_ENC/us01/n1019 ) );
NAND2_X2 \AES_ENC/us01/U77  ( .A1(\AES_ENC/us01/n1059 ), .A2(\AES_ENC/us01/n1114 ), .ZN(\AES_ENC/us01/n1012 ) );
NAND2_X2 \AES_ENC/us01/U76  ( .A1(\AES_ENC/us01/n1010 ), .A2(\AES_ENC/us01/n604 ), .ZN(\AES_ENC/us01/n1011 ) );
NAND2_X2 \AES_ENC/us01/U75  ( .A1(\AES_ENC/us01/n1012 ), .A2(\AES_ENC/us01/n1011 ), .ZN(\AES_ENC/us01/n1016 ) );
NAND4_X2 \AES_ENC/us01/U70  ( .A1(\AES_ENC/us01/n1020 ), .A2(\AES_ENC/us01/n1019 ), .A3(\AES_ENC/us01/n1018 ), .A4(\AES_ENC/us01/n1017 ), .ZN(\AES_ENC/us01/n1021 ) );
NAND2_X2 \AES_ENC/us01/U69  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n1021 ), .ZN(\AES_ENC/us01/n1042 ) );
NAND2_X2 \AES_ENC/us01/U68  ( .A1(\AES_ENC/us01/n1022 ), .A2(\AES_ENC/us01/n1093 ), .ZN(\AES_ENC/us01/n1039 ) );
NAND2_X2 \AES_ENC/us01/U67  ( .A1(\AES_ENC/us01/n1050 ), .A2(\AES_ENC/us01/n1023 ), .ZN(\AES_ENC/us01/n1038 ) );
NAND2_X2 \AES_ENC/us01/U66  ( .A1(\AES_ENC/us01/n1024 ), .A2(\AES_ENC/us01/n1071 ), .ZN(\AES_ENC/us01/n1037 ) );
AND2_X2 \AES_ENC/us01/U60  ( .A1(\AES_ENC/us01/n1030 ), .A2(\AES_ENC/us01/n621 ), .ZN(\AES_ENC/us01/n1078 ) );
NAND4_X2 \AES_ENC/us01/U56  ( .A1(\AES_ENC/us01/n1039 ), .A2(\AES_ENC/us01/n1038 ), .A3(\AES_ENC/us01/n1037 ), .A4(\AES_ENC/us01/n1036 ), .ZN(\AES_ENC/us01/n1040 ) );
NAND2_X2 \AES_ENC/us01/U55  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n1040 ), .ZN(\AES_ENC/us01/n1041 ) );
NAND4_X2 \AES_ENC/us01/U54  ( .A1(\AES_ENC/us01/n1044 ), .A2(\AES_ENC/us01/n1043 ), .A3(\AES_ENC/us01/n1042 ), .A4(\AES_ENC/us01/n1041 ), .ZN(\AES_ENC/sa01_sub[6] ) );
NAND2_X2 \AES_ENC/us01/U53  ( .A1(\AES_ENC/us01/n1072 ), .A2(\AES_ENC/us01/n1045 ), .ZN(\AES_ENC/us01/n1068 ) );
NAND2_X2 \AES_ENC/us01/U52  ( .A1(\AES_ENC/us01/n1046 ), .A2(\AES_ENC/us01/n603 ), .ZN(\AES_ENC/us01/n1067 ) );
NAND2_X2 \AES_ENC/us01/U51  ( .A1(\AES_ENC/us01/n1094 ), .A2(\AES_ENC/us01/n1047 ), .ZN(\AES_ENC/us01/n1066 ) );
NAND4_X2 \AES_ENC/us01/U40  ( .A1(\AES_ENC/us01/n1068 ), .A2(\AES_ENC/us01/n1067 ), .A3(\AES_ENC/us01/n1066 ), .A4(\AES_ENC/us01/n1065 ), .ZN(\AES_ENC/us01/n1069 ) );
NAND2_X2 \AES_ENC/us01/U39  ( .A1(\AES_ENC/us01/n1070 ), .A2(\AES_ENC/us01/n1069 ), .ZN(\AES_ENC/us01/n1135 ) );
NAND2_X2 \AES_ENC/us01/U38  ( .A1(\AES_ENC/us01/n1072 ), .A2(\AES_ENC/us01/n1071 ), .ZN(\AES_ENC/us01/n1088 ) );
NAND2_X2 \AES_ENC/us01/U37  ( .A1(\AES_ENC/us01/n1073 ), .A2(\AES_ENC/us01/n608 ), .ZN(\AES_ENC/us01/n1087 ) );
NAND4_X2 \AES_ENC/us01/U28  ( .A1(\AES_ENC/us01/n1088 ), .A2(\AES_ENC/us01/n1087 ), .A3(\AES_ENC/us01/n1086 ), .A4(\AES_ENC/us01/n1085 ), .ZN(\AES_ENC/us01/n1089 ) );
NAND2_X2 \AES_ENC/us01/U27  ( .A1(\AES_ENC/us01/n1090 ), .A2(\AES_ENC/us01/n1089 ), .ZN(\AES_ENC/us01/n1134 ) );
NAND2_X2 \AES_ENC/us01/U26  ( .A1(\AES_ENC/us01/n1091 ), .A2(\AES_ENC/us01/n1093 ), .ZN(\AES_ENC/us01/n1111 ) );
NAND2_X2 \AES_ENC/us01/U25  ( .A1(\AES_ENC/us01/n1092 ), .A2(\AES_ENC/us01/n1120 ), .ZN(\AES_ENC/us01/n1110 ) );
AND2_X2 \AES_ENC/us01/U22  ( .A1(\AES_ENC/us01/n1097 ), .A2(\AES_ENC/us01/n1096 ), .ZN(\AES_ENC/us01/n1098 ) );
NAND4_X2 \AES_ENC/us01/U14  ( .A1(\AES_ENC/us01/n1111 ), .A2(\AES_ENC/us01/n1110 ), .A3(\AES_ENC/us01/n1109 ), .A4(\AES_ENC/us01/n1108 ), .ZN(\AES_ENC/us01/n1112 ) );
NAND2_X2 \AES_ENC/us01/U13  ( .A1(\AES_ENC/us01/n1113 ), .A2(\AES_ENC/us01/n1112 ), .ZN(\AES_ENC/us01/n1133 ) );
NAND2_X2 \AES_ENC/us01/U12  ( .A1(\AES_ENC/us01/n1115 ), .A2(\AES_ENC/us01/n1114 ), .ZN(\AES_ENC/us01/n1129 ) );
OR2_X2 \AES_ENC/us01/U11  ( .A1(\AES_ENC/us01/n579 ), .A2(\AES_ENC/us01/n1116 ), .ZN(\AES_ENC/us01/n1128 ) );
NAND4_X2 \AES_ENC/us01/U3  ( .A1(\AES_ENC/us01/n1129 ), .A2(\AES_ENC/us01/n1128 ), .A3(\AES_ENC/us01/n1127 ), .A4(\AES_ENC/us01/n1126 ), .ZN(\AES_ENC/us01/n1130 ) );
NAND2_X2 \AES_ENC/us01/U2  ( .A1(\AES_ENC/us01/n1131 ), .A2(\AES_ENC/us01/n1130 ), .ZN(\AES_ENC/us01/n1132 ) );
NAND4_X2 \AES_ENC/us01/U1  ( .A1(\AES_ENC/us01/n1135 ), .A2(\AES_ENC/us01/n1134 ), .A3(\AES_ENC/us01/n1133 ), .A4(\AES_ENC/us01/n1132 ), .ZN(\AES_ENC/sa01_sub[7] ) );
INV_X4 \AES_ENC/us02/U575  ( .A(\AES_ENC/sa02 [7]), .ZN(\AES_ENC/us02/n627 ));
INV_X4 \AES_ENC/us02/U574  ( .A(\AES_ENC/us02/n1114 ), .ZN(\AES_ENC/us02/n625 ) );
INV_X4 \AES_ENC/us02/U573  ( .A(\AES_ENC/sa02 [4]), .ZN(\AES_ENC/us02/n624 ));
INV_X4 \AES_ENC/us02/U572  ( .A(\AES_ENC/us02/n1025 ), .ZN(\AES_ENC/us02/n622 ) );
INV_X4 \AES_ENC/us02/U571  ( .A(\AES_ENC/us02/n1120 ), .ZN(\AES_ENC/us02/n620 ) );
INV_X4 \AES_ENC/us02/U570  ( .A(\AES_ENC/us02/n1121 ), .ZN(\AES_ENC/us02/n619 ) );
INV_X4 \AES_ENC/us02/U569  ( .A(\AES_ENC/us02/n1048 ), .ZN(\AES_ENC/us02/n618 ) );
INV_X4 \AES_ENC/us02/U568  ( .A(\AES_ENC/us02/n974 ), .ZN(\AES_ENC/us02/n616 ) );
INV_X4 \AES_ENC/us02/U567  ( .A(\AES_ENC/us02/n794 ), .ZN(\AES_ENC/us02/n614 ) );
INV_X4 \AES_ENC/us02/U566  ( .A(\AES_ENC/sa02 [2]), .ZN(\AES_ENC/us02/n611 ));
INV_X4 \AES_ENC/us02/U565  ( .A(\AES_ENC/us02/n800 ), .ZN(\AES_ENC/us02/n610 ) );
INV_X4 \AES_ENC/us02/U564  ( .A(\AES_ENC/us02/n925 ), .ZN(\AES_ENC/us02/n609 ) );
INV_X4 \AES_ENC/us02/U563  ( .A(\AES_ENC/us02/n779 ), .ZN(\AES_ENC/us02/n607 ) );
INV_X4 \AES_ENC/us02/U562  ( .A(\AES_ENC/us02/n1022 ), .ZN(\AES_ENC/us02/n603 ) );
INV_X4 \AES_ENC/us02/U561  ( .A(\AES_ENC/us02/n1102 ), .ZN(\AES_ENC/us02/n602 ) );
INV_X4 \AES_ENC/us02/U560  ( .A(\AES_ENC/us02/n929 ), .ZN(\AES_ENC/us02/n601 ) );
INV_X4 \AES_ENC/us02/U559  ( .A(\AES_ENC/us02/n1056 ), .ZN(\AES_ENC/us02/n600 ) );
INV_X4 \AES_ENC/us02/U558  ( .A(\AES_ENC/us02/n1054 ), .ZN(\AES_ENC/us02/n599 ) );
INV_X4 \AES_ENC/us02/U557  ( .A(\AES_ENC/us02/n881 ), .ZN(\AES_ENC/us02/n598 ) );
INV_X4 \AES_ENC/us02/U556  ( .A(\AES_ENC/us02/n926 ), .ZN(\AES_ENC/us02/n597 ) );
INV_X4 \AES_ENC/us02/U555  ( .A(\AES_ENC/us02/n977 ), .ZN(\AES_ENC/us02/n595 ) );
INV_X4 \AES_ENC/us02/U554  ( .A(\AES_ENC/us02/n1031 ), .ZN(\AES_ENC/us02/n594 ) );
INV_X4 \AES_ENC/us02/U553  ( .A(\AES_ENC/us02/n1103 ), .ZN(\AES_ENC/us02/n593 ) );
INV_X4 \AES_ENC/us02/U552  ( .A(\AES_ENC/us02/n1009 ), .ZN(\AES_ENC/us02/n592 ) );
INV_X4 \AES_ENC/us02/U551  ( .A(\AES_ENC/us02/n990 ), .ZN(\AES_ENC/us02/n591 ) );
INV_X4 \AES_ENC/us02/U550  ( .A(\AES_ENC/us02/n1058 ), .ZN(\AES_ENC/us02/n590 ) );
INV_X4 \AES_ENC/us02/U549  ( .A(\AES_ENC/us02/n1074 ), .ZN(\AES_ENC/us02/n589 ) );
INV_X4 \AES_ENC/us02/U548  ( .A(\AES_ENC/us02/n1053 ), .ZN(\AES_ENC/us02/n588 ) );
INV_X4 \AES_ENC/us02/U547  ( .A(\AES_ENC/us02/n826 ), .ZN(\AES_ENC/us02/n587 ) );
INV_X4 \AES_ENC/us02/U546  ( .A(\AES_ENC/us02/n992 ), .ZN(\AES_ENC/us02/n586 ) );
INV_X4 \AES_ENC/us02/U545  ( .A(\AES_ENC/us02/n821 ), .ZN(\AES_ENC/us02/n585 ) );
INV_X4 \AES_ENC/us02/U544  ( .A(\AES_ENC/us02/n910 ), .ZN(\AES_ENC/us02/n584 ) );
INV_X4 \AES_ENC/us02/U543  ( .A(\AES_ENC/us02/n906 ), .ZN(\AES_ENC/us02/n583 ) );
INV_X4 \AES_ENC/us02/U542  ( .A(\AES_ENC/us02/n880 ), .ZN(\AES_ENC/us02/n581 ) );
INV_X4 \AES_ENC/us02/U541  ( .A(\AES_ENC/us02/n1013 ), .ZN(\AES_ENC/us02/n580 ) );
INV_X4 \AES_ENC/us02/U540  ( .A(\AES_ENC/us02/n1092 ), .ZN(\AES_ENC/us02/n579 ) );
INV_X4 \AES_ENC/us02/U539  ( .A(\AES_ENC/us02/n824 ), .ZN(\AES_ENC/us02/n578 ) );
INV_X4 \AES_ENC/us02/U538  ( .A(\AES_ENC/us02/n1091 ), .ZN(\AES_ENC/us02/n577 ) );
INV_X4 \AES_ENC/us02/U537  ( .A(\AES_ENC/us02/n1080 ), .ZN(\AES_ENC/us02/n576 ) );
INV_X4 \AES_ENC/us02/U536  ( .A(\AES_ENC/us02/n959 ), .ZN(\AES_ENC/us02/n575 ) );
INV_X4 \AES_ENC/us02/U535  ( .A(\AES_ENC/sa02 [0]), .ZN(\AES_ENC/us02/n574 ));
NOR2_X2 \AES_ENC/us02/U534  ( .A1(\AES_ENC/sa02 [0]), .A2(\AES_ENC/sa02 [6]),.ZN(\AES_ENC/us02/n1090 ) );
NOR2_X2 \AES_ENC/us02/U533  ( .A1(\AES_ENC/us02/n574 ), .A2(\AES_ENC/sa02 [6]), .ZN(\AES_ENC/us02/n1070 ) );
NOR2_X2 \AES_ENC/us02/U532  ( .A1(\AES_ENC/sa02 [4]), .A2(\AES_ENC/sa02 [3]),.ZN(\AES_ENC/us02/n1025 ) );
INV_X4 \AES_ENC/us02/U531  ( .A(\AES_ENC/us02/n569 ), .ZN(\AES_ENC/us02/n572 ) );
NOR2_X2 \AES_ENC/us02/U530  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n765 ) );
NOR2_X2 \AES_ENC/us02/U529  ( .A1(\AES_ENC/sa02 [4]), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n764 ) );
NOR2_X2 \AES_ENC/us02/U528  ( .A1(\AES_ENC/us02/n765 ), .A2(\AES_ENC/us02/n764 ), .ZN(\AES_ENC/us02/n766 ) );
NOR2_X2 \AES_ENC/us02/U527  ( .A1(\AES_ENC/us02/n766 ), .A2(\AES_ENC/us02/n575 ), .ZN(\AES_ENC/us02/n767 ) );
NOR3_X2 \AES_ENC/us02/U526  ( .A1(\AES_ENC/us02/n627 ), .A2(\AES_ENC/sa02 [5]), .A3(\AES_ENC/us02/n704 ), .ZN(\AES_ENC/us02/n706 ));
NOR2_X2 \AES_ENC/us02/U525  ( .A1(\AES_ENC/us02/n1117 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n707 ) );
NOR2_X2 \AES_ENC/us02/U524  ( .A1(\AES_ENC/sa02 [4]), .A2(\AES_ENC/us02/n579 ), .ZN(\AES_ENC/us02/n705 ) );
NOR3_X2 \AES_ENC/us02/U523  ( .A1(\AES_ENC/us02/n707 ), .A2(\AES_ENC/us02/n706 ), .A3(\AES_ENC/us02/n705 ), .ZN(\AES_ENC/us02/n713 ) );
INV_X4 \AES_ENC/us02/U522  ( .A(\AES_ENC/sa02 [3]), .ZN(\AES_ENC/us02/n621 ));
NAND3_X2 \AES_ENC/us02/U521  ( .A1(\AES_ENC/us02/n652 ), .A2(\AES_ENC/us02/n626 ), .A3(\AES_ENC/sa02 [7]), .ZN(\AES_ENC/us02/n653 ));
NOR2_X2 \AES_ENC/us02/U520  ( .A1(\AES_ENC/us02/n611 ), .A2(\AES_ENC/sa02 [5]), .ZN(\AES_ENC/us02/n925 ) );
NOR2_X2 \AES_ENC/us02/U519  ( .A1(\AES_ENC/sa02 [5]), .A2(\AES_ENC/sa02 [2]),.ZN(\AES_ENC/us02/n974 ) );
INV_X4 \AES_ENC/us02/U518  ( .A(\AES_ENC/sa02 [5]), .ZN(\AES_ENC/us02/n626 ));
NOR2_X2 \AES_ENC/us02/U517  ( .A1(\AES_ENC/us02/n611 ), .A2(\AES_ENC/sa02 [7]), .ZN(\AES_ENC/us02/n779 ) );
NAND3_X2 \AES_ENC/us02/U516  ( .A1(\AES_ENC/us02/n679 ), .A2(\AES_ENC/us02/n678 ), .A3(\AES_ENC/us02/n677 ), .ZN(\AES_ENC/sa02_sub[0] ) );
NOR2_X2 \AES_ENC/us02/U515  ( .A1(\AES_ENC/us02/n626 ), .A2(\AES_ENC/sa02 [2]), .ZN(\AES_ENC/us02/n1048 ) );
NOR4_X2 \AES_ENC/us02/U512  ( .A1(\AES_ENC/us02/n633 ), .A2(\AES_ENC/us02/n632 ), .A3(\AES_ENC/us02/n631 ), .A4(\AES_ENC/us02/n630 ), .ZN(\AES_ENC/us02/n634 ) );
NOR2_X2 \AES_ENC/us02/U510  ( .A1(\AES_ENC/us02/n629 ), .A2(\AES_ENC/us02/n628 ), .ZN(\AES_ENC/us02/n635 ) );
NAND3_X2 \AES_ENC/us02/U509  ( .A1(\AES_ENC/sa02 [2]), .A2(\AES_ENC/sa02 [7]), .A3(\AES_ENC/us02/n1059 ), .ZN(\AES_ENC/us02/n636 ) );
NOR2_X2 \AES_ENC/us02/U508  ( .A1(\AES_ENC/sa02 [7]), .A2(\AES_ENC/sa02 [2]),.ZN(\AES_ENC/us02/n794 ) );
NOR2_X2 \AES_ENC/us02/U507  ( .A1(\AES_ENC/sa02 [4]), .A2(\AES_ENC/sa02 [1]),.ZN(\AES_ENC/us02/n1102 ) );
NOR2_X2 \AES_ENC/us02/U506  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/sa02 [3]), .ZN(\AES_ENC/us02/n1053 ) );
NOR2_X2 \AES_ENC/us02/U505  ( .A1(\AES_ENC/us02/n607 ), .A2(\AES_ENC/sa02 [5]), .ZN(\AES_ENC/us02/n1024 ) );
NOR2_X2 \AES_ENC/us02/U504  ( .A1(\AES_ENC/us02/n625 ), .A2(\AES_ENC/sa02 [2]), .ZN(\AES_ENC/us02/n1093 ) );
NOR2_X2 \AES_ENC/us02/U503  ( .A1(\AES_ENC/us02/n614 ), .A2(\AES_ENC/sa02 [5]), .ZN(\AES_ENC/us02/n1094 ) );
NOR2_X2 \AES_ENC/us02/U502  ( .A1(\AES_ENC/us02/n624 ), .A2(\AES_ENC/sa02 [3]), .ZN(\AES_ENC/us02/n931 ) );
INV_X4 \AES_ENC/us02/U501  ( .A(\AES_ENC/us02/n570 ), .ZN(\AES_ENC/us02/n573 ) );
NOR2_X2 \AES_ENC/us02/U500  ( .A1(\AES_ENC/us02/n1053 ), .A2(\AES_ENC/us02/n1095 ), .ZN(\AES_ENC/us02/n639 ) );
NOR3_X2 \AES_ENC/us02/U499  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n573 ), .A3(\AES_ENC/us02/n1074 ), .ZN(\AES_ENC/us02/n641 ) );
NOR2_X2 \AES_ENC/us02/U498  ( .A1(\AES_ENC/us02/n639 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n640 ) );
NOR2_X2 \AES_ENC/us02/U497  ( .A1(\AES_ENC/us02/n641 ), .A2(\AES_ENC/us02/n640 ), .ZN(\AES_ENC/us02/n646 ) );
NOR3_X2 \AES_ENC/us02/U496  ( .A1(\AES_ENC/us02/n995 ), .A2(\AES_ENC/us02/n586 ), .A3(\AES_ENC/us02/n994 ), .ZN(\AES_ENC/us02/n1002 ) );
NOR2_X2 \AES_ENC/us02/U495  ( .A1(\AES_ENC/us02/n909 ), .A2(\AES_ENC/us02/n908 ), .ZN(\AES_ENC/us02/n920 ) );
NOR2_X2 \AES_ENC/us02/U494  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n823 ) );
NOR2_X2 \AES_ENC/us02/U492  ( .A1(\AES_ENC/us02/n624 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n822 ) );
NOR2_X2 \AES_ENC/us02/U491  ( .A1(\AES_ENC/us02/n823 ), .A2(\AES_ENC/us02/n822 ), .ZN(\AES_ENC/us02/n825 ) );
NOR2_X2 \AES_ENC/us02/U490  ( .A1(\AES_ENC/sa02 [1]), .A2(\AES_ENC/us02/n623 ), .ZN(\AES_ENC/us02/n913 ) );
NOR2_X2 \AES_ENC/us02/U489  ( .A1(\AES_ENC/us02/n913 ), .A2(\AES_ENC/us02/n1091 ), .ZN(\AES_ENC/us02/n914 ) );
NOR2_X2 \AES_ENC/us02/U488  ( .A1(\AES_ENC/us02/n826 ), .A2(\AES_ENC/us02/n572 ), .ZN(\AES_ENC/us02/n827 ) );
NOR3_X2 \AES_ENC/us02/U487  ( .A1(\AES_ENC/us02/n769 ), .A2(\AES_ENC/us02/n768 ), .A3(\AES_ENC/us02/n767 ), .ZN(\AES_ENC/us02/n775 ) );
NOR2_X2 \AES_ENC/us02/U486  ( .A1(\AES_ENC/us02/n1056 ), .A2(\AES_ENC/us02/n1053 ), .ZN(\AES_ENC/us02/n749 ) );
NOR2_X2 \AES_ENC/us02/U483  ( .A1(\AES_ENC/us02/n749 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n752 ) );
INV_X4 \AES_ENC/us02/U482  ( .A(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n596 ));
NOR2_X2 \AES_ENC/us02/U480  ( .A1(\AES_ENC/us02/n1054 ), .A2(\AES_ENC/us02/n1053 ), .ZN(\AES_ENC/us02/n1055 ) );
OR2_X4 \AES_ENC/us02/U479  ( .A1(\AES_ENC/us02/n1094 ), .A2(\AES_ENC/us02/n1093 ), .ZN(\AES_ENC/us02/n571 ) );
AND2_X2 \AES_ENC/us02/U478  ( .A1(\AES_ENC/us02/n571 ), .A2(\AES_ENC/us02/n1095 ), .ZN(\AES_ENC/us02/n1101 ) );
NOR2_X2 \AES_ENC/us02/U477  ( .A1(\AES_ENC/us02/n1074 ), .A2(\AES_ENC/us02/n931 ), .ZN(\AES_ENC/us02/n796 ) );
NOR2_X2 \AES_ENC/us02/U474  ( .A1(\AES_ENC/us02/n796 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n797 ) );
NOR2_X2 \AES_ENC/us02/U473  ( .A1(\AES_ENC/us02/n932 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n933 ) );
NOR2_X2 \AES_ENC/us02/U472  ( .A1(\AES_ENC/us02/n929 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n935 ) );
NOR2_X2 \AES_ENC/us02/U471  ( .A1(\AES_ENC/us02/n931 ), .A2(\AES_ENC/us02/n930 ), .ZN(\AES_ENC/us02/n934 ) );
NOR3_X2 \AES_ENC/us02/U470  ( .A1(\AES_ENC/us02/n935 ), .A2(\AES_ENC/us02/n934 ), .A3(\AES_ENC/us02/n933 ), .ZN(\AES_ENC/us02/n936 ) );
NOR2_X2 \AES_ENC/us02/U469  ( .A1(\AES_ENC/us02/n624 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n1075 ) );
NOR2_X2 \AES_ENC/us02/U468  ( .A1(\AES_ENC/us02/n572 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n949 ) );
NOR2_X2 \AES_ENC/us02/U467  ( .A1(\AES_ENC/us02/n1049 ), .A2(\AES_ENC/us02/n618 ), .ZN(\AES_ENC/us02/n1051 ) );
NOR2_X2 \AES_ENC/us02/U466  ( .A1(\AES_ENC/us02/n1051 ), .A2(\AES_ENC/us02/n1050 ), .ZN(\AES_ENC/us02/n1052 ) );
NOR2_X2 \AES_ENC/us02/U465  ( .A1(\AES_ENC/us02/n1052 ), .A2(\AES_ENC/us02/n592 ), .ZN(\AES_ENC/us02/n1064 ) );
NOR2_X2 \AES_ENC/us02/U464  ( .A1(\AES_ENC/sa02 [1]), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n631 ) );
NOR2_X2 \AES_ENC/us02/U463  ( .A1(\AES_ENC/us02/n1025 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n980 ) );
NOR2_X2 \AES_ENC/us02/U462  ( .A1(\AES_ENC/us02/n1073 ), .A2(\AES_ENC/us02/n1094 ), .ZN(\AES_ENC/us02/n795 ) );
NOR2_X2 \AES_ENC/us02/U461  ( .A1(\AES_ENC/us02/n795 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n799 ) );
NOR2_X2 \AES_ENC/us02/U460  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n981 ) );
NOR2_X2 \AES_ENC/us02/U459  ( .A1(\AES_ENC/us02/n1102 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n643 ) );
NOR2_X2 \AES_ENC/us02/U458  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n621 ), .ZN(\AES_ENC/us02/n642 ) );
NOR2_X2 \AES_ENC/us02/U455  ( .A1(\AES_ENC/us02/n911 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n644 ) );
NOR4_X2 \AES_ENC/us02/U448  ( .A1(\AES_ENC/us02/n644 ), .A2(\AES_ENC/us02/n643 ), .A3(\AES_ENC/us02/n804 ), .A4(\AES_ENC/us02/n642 ), .ZN(\AES_ENC/us02/n645 ) );
NOR2_X2 \AES_ENC/us02/U447  ( .A1(\AES_ENC/us02/n1102 ), .A2(\AES_ENC/us02/n910 ), .ZN(\AES_ENC/us02/n932 ) );
NOR2_X2 \AES_ENC/us02/U442  ( .A1(\AES_ENC/us02/n1102 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n755 ) );
NOR2_X2 \AES_ENC/us02/U441  ( .A1(\AES_ENC/us02/n931 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n743 ) );
NOR2_X2 \AES_ENC/us02/U438  ( .A1(\AES_ENC/us02/n1072 ), .A2(\AES_ENC/us02/n1094 ), .ZN(\AES_ENC/us02/n930 ) );
NOR2_X2 \AES_ENC/us02/U435  ( .A1(\AES_ENC/us02/n1074 ), .A2(\AES_ENC/us02/n1025 ), .ZN(\AES_ENC/us02/n891 ) );
NOR2_X2 \AES_ENC/us02/U434  ( .A1(\AES_ENC/us02/n891 ), .A2(\AES_ENC/us02/n609 ), .ZN(\AES_ENC/us02/n894 ) );
NOR3_X2 \AES_ENC/us02/U433  ( .A1(\AES_ENC/us02/n623 ), .A2(\AES_ENC/sa02 [1]), .A3(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n683 ));
INV_X4 \AES_ENC/us02/U428  ( .A(\AES_ENC/us02/n931 ), .ZN(\AES_ENC/us02/n623 ) );
NOR2_X2 \AES_ENC/us02/U427  ( .A1(\AES_ENC/us02/n996 ), .A2(\AES_ENC/us02/n931 ), .ZN(\AES_ENC/us02/n704 ) );
NOR2_X2 \AES_ENC/us02/U421  ( .A1(\AES_ENC/us02/n931 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n685 ) );
NOR2_X2 \AES_ENC/us02/U420  ( .A1(\AES_ENC/us02/n1029 ), .A2(\AES_ENC/us02/n1025 ), .ZN(\AES_ENC/us02/n1079 ) );
NOR3_X2 \AES_ENC/us02/U419  ( .A1(\AES_ENC/us02/n589 ), .A2(\AES_ENC/us02/n1025 ), .A3(\AES_ENC/us02/n616 ), .ZN(\AES_ENC/us02/n945 ) );
NOR2_X2 \AES_ENC/us02/U418  ( .A1(\AES_ENC/us02/n626 ), .A2(\AES_ENC/us02/n611 ), .ZN(\AES_ENC/us02/n800 ) );
NOR3_X2 \AES_ENC/us02/U417  ( .A1(\AES_ENC/us02/n590 ), .A2(\AES_ENC/us02/n627 ), .A3(\AES_ENC/us02/n611 ), .ZN(\AES_ENC/us02/n798 ) );
NOR3_X2 \AES_ENC/us02/U416  ( .A1(\AES_ENC/us02/n610 ), .A2(\AES_ENC/us02/n572 ), .A3(\AES_ENC/us02/n575 ), .ZN(\AES_ENC/us02/n962 ) );
NOR3_X2 \AES_ENC/us02/U415  ( .A1(\AES_ENC/us02/n959 ), .A2(\AES_ENC/us02/n572 ), .A3(\AES_ENC/us02/n609 ), .ZN(\AES_ENC/us02/n768 ) );
NOR3_X2 \AES_ENC/us02/U414  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n572 ), .A3(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n694 ) );
NOR3_X2 \AES_ENC/us02/U413  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n572 ), .A3(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n895 ) );
NOR3_X2 \AES_ENC/us02/U410  ( .A1(\AES_ENC/us02/n1008 ), .A2(\AES_ENC/us02/n1007 ), .A3(\AES_ENC/us02/n1006 ), .ZN(\AES_ENC/us02/n1018 ) );
NOR4_X2 \AES_ENC/us02/U409  ( .A1(\AES_ENC/us02/n711 ), .A2(\AES_ENC/us02/n710 ), .A3(\AES_ENC/us02/n709 ), .A4(\AES_ENC/us02/n708 ), .ZN(\AES_ENC/us02/n712 ) );
NOR4_X2 \AES_ENC/us02/U406  ( .A1(\AES_ENC/us02/n806 ), .A2(\AES_ENC/us02/n805 ), .A3(\AES_ENC/us02/n804 ), .A4(\AES_ENC/us02/n803 ), .ZN(\AES_ENC/us02/n807 ) );
NOR3_X2 \AES_ENC/us02/U405  ( .A1(\AES_ENC/us02/n799 ), .A2(\AES_ENC/us02/n798 ), .A3(\AES_ENC/us02/n797 ), .ZN(\AES_ENC/us02/n808 ) );
NOR2_X2 \AES_ENC/us02/U404  ( .A1(\AES_ENC/us02/n669 ), .A2(\AES_ENC/us02/n668 ), .ZN(\AES_ENC/us02/n673 ) );
NOR4_X2 \AES_ENC/us02/U403  ( .A1(\AES_ENC/us02/n946 ), .A2(\AES_ENC/us02/n1046 ), .A3(\AES_ENC/us02/n671 ), .A4(\AES_ENC/us02/n670 ), .ZN(\AES_ENC/us02/n672 ) );
NOR3_X2 \AES_ENC/us02/U401  ( .A1(\AES_ENC/us02/n1101 ), .A2(\AES_ENC/us02/n1100 ), .A3(\AES_ENC/us02/n1099 ), .ZN(\AES_ENC/us02/n1109 ) );
NOR4_X2 \AES_ENC/us02/U400  ( .A1(\AES_ENC/us02/n843 ), .A2(\AES_ENC/us02/n842 ), .A3(\AES_ENC/us02/n841 ), .A4(\AES_ENC/us02/n840 ), .ZN(\AES_ENC/us02/n844 ) );
NOR4_X2 \AES_ENC/us02/U399  ( .A1(\AES_ENC/us02/n963 ), .A2(\AES_ENC/us02/n962 ), .A3(\AES_ENC/us02/n961 ), .A4(\AES_ENC/us02/n960 ), .ZN(\AES_ENC/us02/n964 ) );
NOR3_X2 \AES_ENC/us02/U398  ( .A1(\AES_ENC/us02/n743 ), .A2(\AES_ENC/us02/n742 ), .A3(\AES_ENC/us02/n741 ), .ZN(\AES_ENC/us02/n744 ) );
NOR2_X2 \AES_ENC/us02/U397  ( .A1(\AES_ENC/us02/n697 ), .A2(\AES_ENC/us02/n658 ), .ZN(\AES_ENC/us02/n659 ) );
NOR2_X2 \AES_ENC/us02/U396  ( .A1(\AES_ENC/us02/n598 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n885 ) );
NOR2_X2 \AES_ENC/us02/U393  ( .A1(\AES_ENC/us02/n623 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n882 ) );
NOR2_X2 \AES_ENC/us02/U390  ( .A1(\AES_ENC/us02/n1053 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n884 ) );
NOR4_X2 \AES_ENC/us02/U389  ( .A1(\AES_ENC/us02/n885 ), .A2(\AES_ENC/us02/n884 ), .A3(\AES_ENC/us02/n883 ), .A4(\AES_ENC/us02/n882 ), .ZN(\AES_ENC/us02/n886 ) );
NOR2_X2 \AES_ENC/us02/U388  ( .A1(\AES_ENC/us02/n1078 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n1033 ) );
NOR2_X2 \AES_ENC/us02/U387  ( .A1(\AES_ENC/us02/n1031 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n1032 ) );
NOR3_X2 \AES_ENC/us02/U386  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n1025 ), .A3(\AES_ENC/us02/n1074 ), .ZN(\AES_ENC/us02/n1035 ) );
NOR4_X2 \AES_ENC/us02/U385  ( .A1(\AES_ENC/us02/n1035 ), .A2(\AES_ENC/us02/n1034 ), .A3(\AES_ENC/us02/n1033 ), .A4(\AES_ENC/us02/n1032 ), .ZN(\AES_ENC/us02/n1036 ) );
NOR2_X2 \AES_ENC/us02/U384  ( .A1(\AES_ENC/us02/n825 ), .A2(\AES_ENC/us02/n578 ), .ZN(\AES_ENC/us02/n830 ) );
NOR2_X2 \AES_ENC/us02/U383  ( .A1(\AES_ENC/us02/n827 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n829 ) );
NOR2_X2 \AES_ENC/us02/U382  ( .A1(\AES_ENC/us02/n572 ), .A2(\AES_ENC/us02/n579 ), .ZN(\AES_ENC/us02/n828 ) );
NOR4_X2 \AES_ENC/us02/U374  ( .A1(\AES_ENC/us02/n831 ), .A2(\AES_ENC/us02/n830 ), .A3(\AES_ENC/us02/n829 ), .A4(\AES_ENC/us02/n828 ), .ZN(\AES_ENC/us02/n832 ) );
NOR2_X2 \AES_ENC/us02/U373  ( .A1(\AES_ENC/us02/n606 ), .A2(\AES_ENC/us02/n582 ), .ZN(\AES_ENC/us02/n1104 ) );
NOR2_X2 \AES_ENC/us02/U372  ( .A1(\AES_ENC/us02/n1102 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n1106 ) );
NOR2_X2 \AES_ENC/us02/U370  ( .A1(\AES_ENC/us02/n1103 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n1105 ) );
NOR4_X2 \AES_ENC/us02/U369  ( .A1(\AES_ENC/us02/n1107 ), .A2(\AES_ENC/us02/n1106 ), .A3(\AES_ENC/us02/n1105 ), .A4(\AES_ENC/us02/n1104 ), .ZN(\AES_ENC/us02/n1108 ) );
NOR3_X2 \AES_ENC/us02/U368  ( .A1(\AES_ENC/us02/n959 ), .A2(\AES_ENC/us02/n621 ), .A3(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n963 ) );
NOR2_X2 \AES_ENC/us02/U367  ( .A1(\AES_ENC/us02/n626 ), .A2(\AES_ENC/us02/n627 ), .ZN(\AES_ENC/us02/n1114 ) );
INV_X4 \AES_ENC/us02/U366  ( .A(\AES_ENC/us02/n1024 ), .ZN(\AES_ENC/us02/n606 ) );
NOR3_X2 \AES_ENC/us02/U365  ( .A1(\AES_ENC/us02/n910 ), .A2(\AES_ENC/us02/n1059 ), .A3(\AES_ENC/us02/n611 ), .ZN(\AES_ENC/us02/n1115 ) );
INV_X4 \AES_ENC/us02/U364  ( .A(\AES_ENC/us02/n1094 ), .ZN(\AES_ENC/us02/n613 ) );
NOR2_X2 \AES_ENC/us02/U363  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n931 ), .ZN(\AES_ENC/us02/n1100 ) );
INV_X4 \AES_ENC/us02/U354  ( .A(\AES_ENC/us02/n1093 ), .ZN(\AES_ENC/us02/n617 ) );
NOR2_X2 \AES_ENC/us02/U353  ( .A1(\AES_ENC/us02/n569 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n929 ) );
NOR2_X2 \AES_ENC/us02/U352  ( .A1(\AES_ENC/us02/n620 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n926 ) );
NOR2_X2 \AES_ENC/us02/U351  ( .A1(\AES_ENC/us02/n572 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n1095 ) );
NOR2_X2 \AES_ENC/us02/U350  ( .A1(\AES_ENC/us02/n609 ), .A2(\AES_ENC/us02/n627 ), .ZN(\AES_ENC/us02/n1010 ) );
NOR2_X2 \AES_ENC/us02/U349  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n1103 ) );
NOR2_X2 \AES_ENC/us02/U348  ( .A1(\AES_ENC/us02/n622 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n1059 ) );
NOR2_X2 \AES_ENC/us02/U347  ( .A1(\AES_ENC/sa02 [1]), .A2(\AES_ENC/us02/n1120 ), .ZN(\AES_ENC/us02/n1022 ) );
NOR2_X2 \AES_ENC/us02/U346  ( .A1(\AES_ENC/us02/n619 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n911 ) );
NOR2_X2 \AES_ENC/us02/U345  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/us02/n1025 ), .ZN(\AES_ENC/us02/n826 ) );
NOR2_X2 \AES_ENC/us02/U338  ( .A1(\AES_ENC/us02/n626 ), .A2(\AES_ENC/us02/n607 ), .ZN(\AES_ENC/us02/n1072 ) );
NOR2_X2 \AES_ENC/us02/U335  ( .A1(\AES_ENC/us02/n627 ), .A2(\AES_ENC/us02/n616 ), .ZN(\AES_ENC/us02/n956 ) );
NOR2_X2 \AES_ENC/us02/U329  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/us02/n624 ), .ZN(\AES_ENC/us02/n1121 ) );
NOR2_X2 \AES_ENC/us02/U328  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/us02/n624 ), .ZN(\AES_ENC/us02/n1058 ) );
NOR2_X2 \AES_ENC/us02/U327  ( .A1(\AES_ENC/us02/n625 ), .A2(\AES_ENC/us02/n611 ), .ZN(\AES_ENC/us02/n1073 ) );
NOR2_X2 \AES_ENC/us02/U325  ( .A1(\AES_ENC/sa02 [1]), .A2(\AES_ENC/us02/n1025 ), .ZN(\AES_ENC/us02/n1054 ) );
NOR2_X2 \AES_ENC/us02/U324  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/us02/n931 ), .ZN(\AES_ENC/us02/n1029 ) );
NOR2_X2 \AES_ENC/us02/U319  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n1056 ) );
NOR2_X2 \AES_ENC/us02/U318  ( .A1(\AES_ENC/us02/n614 ), .A2(\AES_ENC/us02/n626 ), .ZN(\AES_ENC/us02/n1050 ) );
NOR2_X2 \AES_ENC/us02/U317  ( .A1(\AES_ENC/us02/n1121 ), .A2(\AES_ENC/us02/n1025 ), .ZN(\AES_ENC/us02/n1120 ) );
NOR2_X2 \AES_ENC/us02/U316  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/us02/n572 ), .ZN(\AES_ENC/us02/n1074 ) );
NOR2_X2 \AES_ENC/us02/U315  ( .A1(\AES_ENC/us02/n1058 ), .A2(\AES_ENC/us02/n1054 ), .ZN(\AES_ENC/us02/n878 ) );
NOR2_X2 \AES_ENC/us02/U314  ( .A1(\AES_ENC/us02/n878 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n879 ) );
NOR2_X2 \AES_ENC/us02/U312  ( .A1(\AES_ENC/us02/n880 ), .A2(\AES_ENC/us02/n879 ), .ZN(\AES_ENC/us02/n887 ) );
NOR2_X2 \AES_ENC/us02/U311  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n588 ), .ZN(\AES_ENC/us02/n957 ) );
NOR2_X2 \AES_ENC/us02/U310  ( .A1(\AES_ENC/us02/n958 ), .A2(\AES_ENC/us02/n957 ), .ZN(\AES_ENC/us02/n965 ) );
NOR3_X2 \AES_ENC/us02/U309  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n1091 ), .A3(\AES_ENC/us02/n1022 ), .ZN(\AES_ENC/us02/n720 ) );
NOR3_X2 \AES_ENC/us02/U303  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n1054 ), .A3(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n719 ) );
NOR2_X2 \AES_ENC/us02/U302  ( .A1(\AES_ENC/us02/n720 ), .A2(\AES_ENC/us02/n719 ), .ZN(\AES_ENC/us02/n726 ) );
NOR2_X2 \AES_ENC/us02/U300  ( .A1(\AES_ENC/us02/n614 ), .A2(\AES_ENC/us02/n591 ), .ZN(\AES_ENC/us02/n865 ) );
NOR2_X2 \AES_ENC/us02/U299  ( .A1(\AES_ENC/us02/n1059 ), .A2(\AES_ENC/us02/n1058 ), .ZN(\AES_ENC/us02/n1060 ) );
NOR2_X2 \AES_ENC/us02/U298  ( .A1(\AES_ENC/us02/n1095 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n668 ) );
NOR2_X2 \AES_ENC/us02/U297  ( .A1(\AES_ENC/us02/n911 ), .A2(\AES_ENC/us02/n910 ), .ZN(\AES_ENC/us02/n912 ) );
NOR2_X2 \AES_ENC/us02/U296  ( .A1(\AES_ENC/us02/n912 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n916 ) );
NOR2_X2 \AES_ENC/us02/U295  ( .A1(\AES_ENC/us02/n826 ), .A2(\AES_ENC/us02/n573 ), .ZN(\AES_ENC/us02/n750 ) );
NOR2_X2 \AES_ENC/us02/U294  ( .A1(\AES_ENC/us02/n750 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n751 ) );
NOR2_X2 \AES_ENC/us02/U293  ( .A1(\AES_ENC/us02/n907 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n908 ) );
NOR2_X2 \AES_ENC/us02/U292  ( .A1(\AES_ENC/us02/n990 ), .A2(\AES_ENC/us02/n926 ), .ZN(\AES_ENC/us02/n780 ) );
NOR2_X2 \AES_ENC/us02/U291  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n584 ), .ZN(\AES_ENC/us02/n838 ) );
NOR2_X2 \AES_ENC/us02/U290  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n602 ), .ZN(\AES_ENC/us02/n837 ) );
NOR2_X2 \AES_ENC/us02/U284  ( .A1(\AES_ENC/us02/n838 ), .A2(\AES_ENC/us02/n837 ), .ZN(\AES_ENC/us02/n845 ) );
NOR2_X2 \AES_ENC/us02/U283  ( .A1(\AES_ENC/us02/n1022 ), .A2(\AES_ENC/us02/n1058 ), .ZN(\AES_ENC/us02/n740 ) );
NOR2_X2 \AES_ENC/us02/U282  ( .A1(\AES_ENC/us02/n740 ), .A2(\AES_ENC/us02/n616 ), .ZN(\AES_ENC/us02/n742 ) );
NOR2_X2 \AES_ENC/us02/U281  ( .A1(\AES_ENC/us02/n1098 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n1099 ) );
NOR2_X2 \AES_ENC/us02/U280  ( .A1(\AES_ENC/us02/n1120 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n993 ) );
NOR2_X2 \AES_ENC/us02/U279  ( .A1(\AES_ENC/us02/n993 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n994 ) );
NOR2_X2 \AES_ENC/us02/U273  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n620 ), .ZN(\AES_ENC/us02/n1026 ) );
NOR2_X2 \AES_ENC/us02/U272  ( .A1(\AES_ENC/us02/n573 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n1027 ) );
NOR2_X2 \AES_ENC/us02/U271  ( .A1(\AES_ENC/us02/n1027 ), .A2(\AES_ENC/us02/n1026 ), .ZN(\AES_ENC/us02/n1028 ) );
NOR2_X2 \AES_ENC/us02/U270  ( .A1(\AES_ENC/us02/n1029 ), .A2(\AES_ENC/us02/n1028 ), .ZN(\AES_ENC/us02/n1034 ) );
NOR4_X2 \AES_ENC/us02/U269  ( .A1(\AES_ENC/us02/n757 ), .A2(\AES_ENC/us02/n756 ), .A3(\AES_ENC/us02/n755 ), .A4(\AES_ENC/us02/n754 ), .ZN(\AES_ENC/us02/n758 ) );
NOR2_X2 \AES_ENC/us02/U268  ( .A1(\AES_ENC/us02/n752 ), .A2(\AES_ENC/us02/n751 ), .ZN(\AES_ENC/us02/n759 ) );
NOR2_X2 \AES_ENC/us02/U267  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n1071 ), .ZN(\AES_ENC/us02/n669 ) );
NOR2_X2 \AES_ENC/us02/U263  ( .A1(\AES_ENC/us02/n1056 ), .A2(\AES_ENC/us02/n990 ), .ZN(\AES_ENC/us02/n991 ) );
NOR2_X2 \AES_ENC/us02/U262  ( .A1(\AES_ENC/us02/n991 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n995 ) );
NOR2_X2 \AES_ENC/us02/U258  ( .A1(\AES_ENC/us02/n607 ), .A2(\AES_ENC/us02/n590 ), .ZN(\AES_ENC/us02/n1008 ) );
NOR2_X2 \AES_ENC/us02/U255  ( .A1(\AES_ENC/us02/n839 ), .A2(\AES_ENC/us02/n582 ), .ZN(\AES_ENC/us02/n693 ) );
NOR2_X2 \AES_ENC/us02/U254  ( .A1(\AES_ENC/us02/n606 ), .A2(\AES_ENC/us02/n906 ), .ZN(\AES_ENC/us02/n741 ) );
NOR2_X2 \AES_ENC/us02/U253  ( .A1(\AES_ENC/us02/n1054 ), .A2(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n763 ) );
NOR2_X2 \AES_ENC/us02/U252  ( .A1(\AES_ENC/us02/n763 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n769 ) );
NOR2_X2 \AES_ENC/us02/U251  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n577 ), .ZN(\AES_ENC/us02/n1007 ) );
NOR2_X2 \AES_ENC/us02/U250  ( .A1(\AES_ENC/us02/n609 ), .A2(\AES_ENC/us02/n580 ), .ZN(\AES_ENC/us02/n1123 ) );
NOR2_X2 \AES_ENC/us02/U243  ( .A1(\AES_ENC/us02/n609 ), .A2(\AES_ENC/us02/n590 ), .ZN(\AES_ENC/us02/n710 ) );
INV_X4 \AES_ENC/us02/U242  ( .A(\AES_ENC/us02/n1029 ), .ZN(\AES_ENC/us02/n582 ) );
NOR2_X2 \AES_ENC/us02/U241  ( .A1(\AES_ENC/us02/n616 ), .A2(\AES_ENC/us02/n597 ), .ZN(\AES_ENC/us02/n883 ) );
NOR2_X2 \AES_ENC/us02/U240  ( .A1(\AES_ENC/us02/n593 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n1125 ) );
NOR2_X2 \AES_ENC/us02/U239  ( .A1(\AES_ENC/us02/n990 ), .A2(\AES_ENC/us02/n929 ), .ZN(\AES_ENC/us02/n892 ) );
NOR2_X2 \AES_ENC/us02/U238  ( .A1(\AES_ENC/us02/n892 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n893 ) );
NOR2_X2 \AES_ENC/us02/U237  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n602 ), .ZN(\AES_ENC/us02/n950 ) );
NOR2_X2 \AES_ENC/us02/U236  ( .A1(\AES_ENC/us02/n1079 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n1082 ) );
NOR2_X2 \AES_ENC/us02/U235  ( .A1(\AES_ENC/us02/n910 ), .A2(\AES_ENC/us02/n1056 ), .ZN(\AES_ENC/us02/n941 ) );
NOR2_X2 \AES_ENC/us02/U234  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n1077 ), .ZN(\AES_ENC/us02/n841 ) );
NOR2_X2 \AES_ENC/us02/U229  ( .A1(\AES_ENC/us02/n623 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n630 ) );
NOR2_X2 \AES_ENC/us02/U228  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n602 ), .ZN(\AES_ENC/us02/n806 ) );
NOR2_X2 \AES_ENC/us02/U227  ( .A1(\AES_ENC/us02/n623 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n948 ) );
NOR2_X2 \AES_ENC/us02/U226  ( .A1(\AES_ENC/us02/n606 ), .A2(\AES_ENC/us02/n589 ), .ZN(\AES_ENC/us02/n997 ) );
NOR2_X2 \AES_ENC/us02/U225  ( .A1(\AES_ENC/us02/n1121 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n1122 ) );
NOR2_X2 \AES_ENC/us02/U223  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n1023 ), .ZN(\AES_ENC/us02/n756 ) );
NOR2_X2 \AES_ENC/us02/U222  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n602 ), .ZN(\AES_ENC/us02/n870 ) );
NOR2_X2 \AES_ENC/us02/U221  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n569 ), .ZN(\AES_ENC/us02/n947 ) );
NOR2_X2 \AES_ENC/us02/U217  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n1077 ), .ZN(\AES_ENC/us02/n1084 ) );
NOR2_X2 \AES_ENC/us02/U213  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n855 ), .ZN(\AES_ENC/us02/n709 ) );
NOR2_X2 \AES_ENC/us02/U212  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n589 ), .ZN(\AES_ENC/us02/n868 ) );
NOR2_X2 \AES_ENC/us02/U211  ( .A1(\AES_ENC/us02/n1120 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n1124 ) );
NOR2_X2 \AES_ENC/us02/U210  ( .A1(\AES_ENC/us02/n1120 ), .A2(\AES_ENC/us02/n839 ), .ZN(\AES_ENC/us02/n842 ) );
NOR2_X2 \AES_ENC/us02/U209  ( .A1(\AES_ENC/us02/n1120 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n696 ) );
NOR2_X2 \AES_ENC/us02/U208  ( .A1(\AES_ENC/us02/n1074 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n1076 ) );
NOR2_X2 \AES_ENC/us02/U207  ( .A1(\AES_ENC/us02/n1074 ), .A2(\AES_ENC/us02/n620 ), .ZN(\AES_ENC/us02/n781 ) );
NOR3_X2 \AES_ENC/us02/U201  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n1056 ), .A3(\AES_ENC/us02/n990 ), .ZN(\AES_ENC/us02/n979 ) );
NOR3_X2 \AES_ENC/us02/U200  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n1058 ), .A3(\AES_ENC/us02/n1059 ), .ZN(\AES_ENC/us02/n854 ) );
NOR2_X2 \AES_ENC/us02/U199  ( .A1(\AES_ENC/us02/n996 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n869 ) );
NOR2_X2 \AES_ENC/us02/U198  ( .A1(\AES_ENC/us02/n1056 ), .A2(\AES_ENC/us02/n1074 ), .ZN(\AES_ENC/us02/n1057 ) );
NOR3_X2 \AES_ENC/us02/U197  ( .A1(\AES_ENC/us02/n607 ), .A2(\AES_ENC/us02/n1120 ), .A3(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n978 ) );
NOR2_X2 \AES_ENC/us02/U196  ( .A1(\AES_ENC/us02/n996 ), .A2(\AES_ENC/us02/n911 ), .ZN(\AES_ENC/us02/n1116 ) );
NOR2_X2 \AES_ENC/us02/U195  ( .A1(\AES_ENC/us02/n1074 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n754 ) );
NOR2_X2 \AES_ENC/us02/U194  ( .A1(\AES_ENC/us02/n926 ), .A2(\AES_ENC/us02/n1103 ), .ZN(\AES_ENC/us02/n977 ) );
NOR2_X2 \AES_ENC/us02/U187  ( .A1(\AES_ENC/us02/n839 ), .A2(\AES_ENC/us02/n824 ), .ZN(\AES_ENC/us02/n1092 ) );
NOR2_X2 \AES_ENC/us02/U186  ( .A1(\AES_ENC/us02/n573 ), .A2(\AES_ENC/us02/n1074 ), .ZN(\AES_ENC/us02/n684 ) );
NOR2_X2 \AES_ENC/us02/U185  ( .A1(\AES_ENC/us02/n826 ), .A2(\AES_ENC/us02/n1059 ), .ZN(\AES_ENC/us02/n907 ) );
NOR3_X2 \AES_ENC/us02/U184  ( .A1(\AES_ENC/us02/n625 ), .A2(\AES_ENC/us02/n1115 ), .A3(\AES_ENC/us02/n585 ), .ZN(\AES_ENC/us02/n831 ) );
NOR3_X2 \AES_ENC/us02/U183  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n1056 ), .A3(\AES_ENC/us02/n990 ), .ZN(\AES_ENC/us02/n896 ) );
NOR3_X2 \AES_ENC/us02/U182  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n573 ), .A3(\AES_ENC/us02/n1013 ), .ZN(\AES_ENC/us02/n670 ) );
NOR3_X2 \AES_ENC/us02/U181  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n1091 ), .A3(\AES_ENC/us02/n1022 ), .ZN(\AES_ENC/us02/n843 ) );
NOR2_X2 \AES_ENC/us02/U180  ( .A1(\AES_ENC/us02/n1029 ), .A2(\AES_ENC/us02/n1095 ), .ZN(\AES_ENC/us02/n735 ) );
NAND3_X2 \AES_ENC/us02/U174  ( .A1(\AES_ENC/us02/n569 ), .A2(\AES_ENC/us02/n582 ), .A3(\AES_ENC/us02/n681 ), .ZN(\AES_ENC/us02/n691 ) );
NOR2_X2 \AES_ENC/us02/U173  ( .A1(\AES_ENC/us02/n683 ), .A2(\AES_ENC/us02/n682 ), .ZN(\AES_ENC/us02/n690 ) );
NOR3_X2 \AES_ENC/us02/U172  ( .A1(\AES_ENC/us02/n695 ), .A2(\AES_ENC/us02/n694 ), .A3(\AES_ENC/us02/n693 ), .ZN(\AES_ENC/us02/n700 ) );
NOR4_X2 \AES_ENC/us02/U171  ( .A1(\AES_ENC/us02/n983 ), .A2(\AES_ENC/us02/n698 ), .A3(\AES_ENC/us02/n697 ), .A4(\AES_ENC/us02/n696 ), .ZN(\AES_ENC/us02/n699 ) );
NOR2_X2 \AES_ENC/us02/U170  ( .A1(\AES_ENC/us02/n1100 ), .A2(\AES_ENC/us02/n854 ), .ZN(\AES_ENC/us02/n860 ) );
NOR4_X2 \AES_ENC/us02/U169  ( .A1(\AES_ENC/us02/n1125 ), .A2(\AES_ENC/us02/n1124 ), .A3(\AES_ENC/us02/n1123 ), .A4(\AES_ENC/us02/n1122 ), .ZN(\AES_ENC/us02/n1126 ) );
NOR4_X2 \AES_ENC/us02/U168  ( .A1(\AES_ENC/us02/n1084 ), .A2(\AES_ENC/us02/n1083 ), .A3(\AES_ENC/us02/n1082 ), .A4(\AES_ENC/us02/n1081 ), .ZN(\AES_ENC/us02/n1085 ) );
NOR2_X2 \AES_ENC/us02/U162  ( .A1(\AES_ENC/us02/n1076 ), .A2(\AES_ENC/us02/n1075 ), .ZN(\AES_ENC/us02/n1086 ) );
NOR4_X2 \AES_ENC/us02/U161  ( .A1(\AES_ENC/us02/n896 ), .A2(\AES_ENC/us02/n895 ), .A3(\AES_ENC/us02/n894 ), .A4(\AES_ENC/us02/n893 ), .ZN(\AES_ENC/us02/n897 ) );
NOR2_X2 \AES_ENC/us02/U160  ( .A1(\AES_ENC/us02/n866 ), .A2(\AES_ENC/us02/n865 ), .ZN(\AES_ENC/us02/n872 ) );
NOR4_X2 \AES_ENC/us02/U159  ( .A1(\AES_ENC/us02/n870 ), .A2(\AES_ENC/us02/n869 ), .A3(\AES_ENC/us02/n868 ), .A4(\AES_ENC/us02/n867 ), .ZN(\AES_ENC/us02/n871 ) );
NOR2_X2 \AES_ENC/us02/U158  ( .A1(\AES_ENC/us02/n946 ), .A2(\AES_ENC/us02/n945 ), .ZN(\AES_ENC/us02/n952 ) );
NOR4_X2 \AES_ENC/us02/U157  ( .A1(\AES_ENC/us02/n950 ), .A2(\AES_ENC/us02/n949 ), .A3(\AES_ENC/us02/n948 ), .A4(\AES_ENC/us02/n947 ), .ZN(\AES_ENC/us02/n951 ) );
NOR4_X2 \AES_ENC/us02/U156  ( .A1(\AES_ENC/us02/n983 ), .A2(\AES_ENC/us02/n982 ), .A3(\AES_ENC/us02/n981 ), .A4(\AES_ENC/us02/n980 ), .ZN(\AES_ENC/us02/n984 ) );
NOR2_X2 \AES_ENC/us02/U155  ( .A1(\AES_ENC/us02/n979 ), .A2(\AES_ENC/us02/n978 ), .ZN(\AES_ENC/us02/n985 ) );
NOR3_X2 \AES_ENC/us02/U154  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n1054 ), .A3(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n961 ) );
NOR3_X2 \AES_ENC/us02/U153  ( .A1(\AES_ENC/us02/n620 ), .A2(\AES_ENC/us02/n1074 ), .A3(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n671 ) );
NOR2_X2 \AES_ENC/us02/U152  ( .A1(\AES_ENC/us02/n1057 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n1062 ) );
NOR2_X2 \AES_ENC/us02/U143  ( .A1(\AES_ENC/us02/n1055 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n1063 ) );
NOR2_X2 \AES_ENC/us02/U142  ( .A1(\AES_ENC/us02/n1060 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n1061 ) );
NOR4_X2 \AES_ENC/us02/U141  ( .A1(\AES_ENC/us02/n1064 ), .A2(\AES_ENC/us02/n1063 ), .A3(\AES_ENC/us02/n1062 ), .A4(\AES_ENC/us02/n1061 ), .ZN(\AES_ENC/us02/n1065 ) );
NOR2_X2 \AES_ENC/us02/U140  ( .A1(\AES_ENC/us02/n735 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n687 ) );
NOR2_X2 \AES_ENC/us02/U132  ( .A1(\AES_ENC/us02/n684 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n688 ) );
NOR2_X2 \AES_ENC/us02/U131  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n600 ), .ZN(\AES_ENC/us02/n686 ) );
NOR4_X2 \AES_ENC/us02/U130  ( .A1(\AES_ENC/us02/n688 ), .A2(\AES_ENC/us02/n687 ), .A3(\AES_ENC/us02/n686 ), .A4(\AES_ENC/us02/n685 ), .ZN(\AES_ENC/us02/n689 ) );
NOR2_X2 \AES_ENC/us02/U129  ( .A1(\AES_ENC/us02/n616 ), .A2(\AES_ENC/us02/n580 ), .ZN(\AES_ENC/us02/n771 ) );
NOR2_X2 \AES_ENC/us02/U128  ( .A1(\AES_ENC/us02/n1103 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n772 ) );
NOR2_X2 \AES_ENC/us02/U127  ( .A1(\AES_ENC/us02/n610 ), .A2(\AES_ENC/us02/n599 ), .ZN(\AES_ENC/us02/n773 ) );
NOR4_X2 \AES_ENC/us02/U126  ( .A1(\AES_ENC/us02/n773 ), .A2(\AES_ENC/us02/n772 ), .A3(\AES_ENC/us02/n771 ), .A4(\AES_ENC/us02/n770 ), .ZN(\AES_ENC/us02/n774 ) );
NOR2_X2 \AES_ENC/us02/U121  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n595 ), .ZN(\AES_ENC/us02/n858 ) );
NOR2_X2 \AES_ENC/us02/U120  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n855 ), .ZN(\AES_ENC/us02/n857 ) );
NOR2_X2 \AES_ENC/us02/U119  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n587 ), .ZN(\AES_ENC/us02/n856 ) );
NOR4_X2 \AES_ENC/us02/U118  ( .A1(\AES_ENC/us02/n858 ), .A2(\AES_ENC/us02/n857 ), .A3(\AES_ENC/us02/n856 ), .A4(\AES_ENC/us02/n958 ), .ZN(\AES_ENC/us02/n859 ) );
NOR3_X2 \AES_ENC/us02/U117  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n1120 ), .A3(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n918 ) );
NOR3_X2 \AES_ENC/us02/U116  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n573 ), .A3(\AES_ENC/us02/n1013 ), .ZN(\AES_ENC/us02/n917 ) );
NOR2_X2 \AES_ENC/us02/U115  ( .A1(\AES_ENC/us02/n914 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n915 ) );
NOR4_X2 \AES_ENC/us02/U106  ( .A1(\AES_ENC/us02/n918 ), .A2(\AES_ENC/us02/n917 ), .A3(\AES_ENC/us02/n916 ), .A4(\AES_ENC/us02/n915 ), .ZN(\AES_ENC/us02/n919 ) );
NOR2_X2 \AES_ENC/us02/U105  ( .A1(\AES_ENC/us02/n780 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n784 ) );
NOR2_X2 \AES_ENC/us02/U104  ( .A1(\AES_ENC/us02/n1117 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n782 ) );
NOR2_X2 \AES_ENC/us02/U103  ( .A1(\AES_ENC/us02/n781 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n783 ) );
NOR4_X2 \AES_ENC/us02/U102  ( .A1(\AES_ENC/us02/n880 ), .A2(\AES_ENC/us02/n784 ), .A3(\AES_ENC/us02/n783 ), .A4(\AES_ENC/us02/n782 ), .ZN(\AES_ENC/us02/n785 ) );
NOR2_X2 \AES_ENC/us02/U101  ( .A1(\AES_ENC/us02/n583 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n814 ) );
NOR2_X2 \AES_ENC/us02/U100  ( .A1(\AES_ENC/us02/n907 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n813 ) );
NOR3_X2 \AES_ENC/us02/U95  ( .A1(\AES_ENC/us02/n606 ), .A2(\AES_ENC/us02/n1058 ), .A3(\AES_ENC/us02/n1059 ), .ZN(\AES_ENC/us02/n815 ) );
NOR4_X2 \AES_ENC/us02/U94  ( .A1(\AES_ENC/us02/n815 ), .A2(\AES_ENC/us02/n814 ), .A3(\AES_ENC/us02/n813 ), .A4(\AES_ENC/us02/n812 ), .ZN(\AES_ENC/us02/n816 ) );
NOR2_X2 \AES_ENC/us02/U93  ( .A1(\AES_ENC/us02/n617 ), .A2(\AES_ENC/us02/n569 ), .ZN(\AES_ENC/us02/n721 ) );
NOR2_X2 \AES_ENC/us02/U92  ( .A1(\AES_ENC/us02/n1031 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n723 ) );
NOR2_X2 \AES_ENC/us02/U91  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n1096 ), .ZN(\AES_ENC/us02/n722 ) );
NOR4_X2 \AES_ENC/us02/U90  ( .A1(\AES_ENC/us02/n724 ), .A2(\AES_ENC/us02/n723 ), .A3(\AES_ENC/us02/n722 ), .A4(\AES_ENC/us02/n721 ), .ZN(\AES_ENC/us02/n725 ) );
NOR2_X2 \AES_ENC/us02/U89  ( .A1(\AES_ENC/us02/n911 ), .A2(\AES_ENC/us02/n990 ), .ZN(\AES_ENC/us02/n1009 ) );
NOR2_X2 \AES_ENC/us02/U88  ( .A1(\AES_ENC/us02/n1013 ), .A2(\AES_ENC/us02/n573 ), .ZN(\AES_ENC/us02/n1014 ) );
NOR2_X2 \AES_ENC/us02/U87  ( .A1(\AES_ENC/us02/n1014 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n1015 ) );
NOR4_X2 \AES_ENC/us02/U86  ( .A1(\AES_ENC/us02/n1016 ), .A2(\AES_ENC/us02/n1015 ), .A3(\AES_ENC/us02/n1119 ), .A4(\AES_ENC/us02/n1046 ), .ZN(\AES_ENC/us02/n1017 ) );
NOR2_X2 \AES_ENC/us02/U81  ( .A1(\AES_ENC/us02/n996 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n998 ) );
NOR2_X2 \AES_ENC/us02/U80  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n577 ), .ZN(\AES_ENC/us02/n1000 ) );
NOR2_X2 \AES_ENC/us02/U79  ( .A1(\AES_ENC/us02/n616 ), .A2(\AES_ENC/us02/n1096 ), .ZN(\AES_ENC/us02/n999 ) );
NOR4_X2 \AES_ENC/us02/U78  ( .A1(\AES_ENC/us02/n1000 ), .A2(\AES_ENC/us02/n999 ), .A3(\AES_ENC/us02/n998 ), .A4(\AES_ENC/us02/n997 ), .ZN(\AES_ENC/us02/n1001 ) );
NOR2_X2 \AES_ENC/us02/U74  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n1096 ), .ZN(\AES_ENC/us02/n697 ) );
NOR2_X2 \AES_ENC/us02/U73  ( .A1(\AES_ENC/us02/n620 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n958 ) );
NOR2_X2 \AES_ENC/us02/U72  ( .A1(\AES_ENC/us02/n911 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n983 ) );
NOR2_X2 \AES_ENC/us02/U71  ( .A1(\AES_ENC/us02/n1054 ), .A2(\AES_ENC/us02/n1103 ), .ZN(\AES_ENC/us02/n1031 ) );
INV_X4 \AES_ENC/us02/U65  ( .A(\AES_ENC/us02/n1050 ), .ZN(\AES_ENC/us02/n612 ) );
INV_X4 \AES_ENC/us02/U64  ( .A(\AES_ENC/us02/n1072 ), .ZN(\AES_ENC/us02/n605 ) );
INV_X4 \AES_ENC/us02/U63  ( .A(\AES_ENC/us02/n1073 ), .ZN(\AES_ENC/us02/n604 ) );
NOR2_X2 \AES_ENC/us02/U62  ( .A1(\AES_ENC/us02/n582 ), .A2(\AES_ENC/us02/n613 ), .ZN(\AES_ENC/us02/n880 ) );
NOR3_X2 \AES_ENC/us02/U61  ( .A1(\AES_ENC/us02/n826 ), .A2(\AES_ENC/us02/n1121 ), .A3(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n946 ) );
INV_X4 \AES_ENC/us02/U59  ( .A(\AES_ENC/us02/n1010 ), .ZN(\AES_ENC/us02/n608 ) );
NOR3_X2 \AES_ENC/us02/U58  ( .A1(\AES_ENC/us02/n573 ), .A2(\AES_ENC/us02/n1029 ), .A3(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n1119 ) );
INV_X4 \AES_ENC/us02/U57  ( .A(\AES_ENC/us02/n956 ), .ZN(\AES_ENC/us02/n615 ) );
NOR2_X2 \AES_ENC/us02/U50  ( .A1(\AES_ENC/us02/n623 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n1013 ) );
NOR2_X2 \AES_ENC/us02/U49  ( .A1(\AES_ENC/us02/n620 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n910 ) );
NOR2_X2 \AES_ENC/us02/U48  ( .A1(\AES_ENC/us02/n569 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n1091 ) );
NOR2_X2 \AES_ENC/us02/U47  ( .A1(\AES_ENC/us02/n622 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n990 ) );
NOR2_X2 \AES_ENC/us02/U46  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/us02/n1121 ), .ZN(\AES_ENC/us02/n996 ) );
NOR2_X2 \AES_ENC/us02/U45  ( .A1(\AES_ENC/us02/n610 ), .A2(\AES_ENC/us02/n600 ), .ZN(\AES_ENC/us02/n628 ) );
NOR2_X2 \AES_ENC/us02/U44  ( .A1(\AES_ENC/us02/n576 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n866 ) );
NOR2_X2 \AES_ENC/us02/U43  ( .A1(\AES_ENC/us02/n603 ), .A2(\AES_ENC/us02/n610 ), .ZN(\AES_ENC/us02/n1006 ) );
NOR2_X2 \AES_ENC/us02/U42  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n1117 ), .ZN(\AES_ENC/us02/n1118 ) );
NOR2_X2 \AES_ENC/us02/U41  ( .A1(\AES_ENC/us02/n1119 ), .A2(\AES_ENC/us02/n1118 ), .ZN(\AES_ENC/us02/n1127 ) );
NOR2_X2 \AES_ENC/us02/U36  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n594 ), .ZN(\AES_ENC/us02/n629 ) );
NOR2_X2 \AES_ENC/us02/U35  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n906 ), .ZN(\AES_ENC/us02/n909 ) );
NOR2_X2 \AES_ENC/us02/U34  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n597 ), .ZN(\AES_ENC/us02/n658 ) );
NOR2_X2 \AES_ENC/us02/U33  ( .A1(\AES_ENC/us02/n1116 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n695 ) );
NOR2_X2 \AES_ENC/us02/U32  ( .A1(\AES_ENC/us02/n1078 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n1083 ) );
NOR2_X2 \AES_ENC/us02/U31  ( .A1(\AES_ENC/us02/n941 ), .A2(\AES_ENC/us02/n608 ), .ZN(\AES_ENC/us02/n724 ) );
NOR2_X2 \AES_ENC/us02/U30  ( .A1(\AES_ENC/us02/n598 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n1107 ) );
NOR2_X2 \AES_ENC/us02/U29  ( .A1(\AES_ENC/us02/n576 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n840 ) );
NOR2_X2 \AES_ENC/us02/U24  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n593 ), .ZN(\AES_ENC/us02/n633 ) );
NOR2_X2 \AES_ENC/us02/U23  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n1080 ), .ZN(\AES_ENC/us02/n1081 ) );
NOR2_X2 \AES_ENC/us02/U21  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n1045 ), .ZN(\AES_ENC/us02/n812 ) );
NOR2_X2 \AES_ENC/us02/U20  ( .A1(\AES_ENC/us02/n1009 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n960 ) );
NOR2_X2 \AES_ENC/us02/U19  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n601 ), .ZN(\AES_ENC/us02/n982 ) );
NOR2_X2 \AES_ENC/us02/U18  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n594 ), .ZN(\AES_ENC/us02/n757 ) );
NOR2_X2 \AES_ENC/us02/U17  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n590 ), .ZN(\AES_ENC/us02/n698 ) );
NOR2_X2 \AES_ENC/us02/U16  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n619 ), .ZN(\AES_ENC/us02/n708 ) );
NOR2_X2 \AES_ENC/us02/U15  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n582 ), .ZN(\AES_ENC/us02/n770 ) );
NOR2_X2 \AES_ENC/us02/U10  ( .A1(\AES_ENC/us02/n619 ), .A2(\AES_ENC/us02/n604 ), .ZN(\AES_ENC/us02/n803 ) );
NOR2_X2 \AES_ENC/us02/U9  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n881 ), .ZN(\AES_ENC/us02/n711 ) );
NOR2_X2 \AES_ENC/us02/U8  ( .A1(\AES_ENC/us02/n615 ), .A2(\AES_ENC/us02/n582 ), .ZN(\AES_ENC/us02/n867 ) );
NOR2_X2 \AES_ENC/us02/U7  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n599 ), .ZN(\AES_ENC/us02/n804 ) );
NOR2_X2 \AES_ENC/us02/U6  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n620 ), .ZN(\AES_ENC/us02/n1046 ) );
OR2_X4 \AES_ENC/us02/U5  ( .A1(\AES_ENC/us02/n624 ), .A2(\AES_ENC/sa02 [1]),.ZN(\AES_ENC/us02/n570 ) );
OR2_X4 \AES_ENC/us02/U4  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/sa02 [4]),.ZN(\AES_ENC/us02/n569 ) );
NAND2_X2 \AES_ENC/us02/U514  ( .A1(\AES_ENC/us02/n1121 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n1030 ) );
AND2_X2 \AES_ENC/us02/U513  ( .A1(\AES_ENC/us02/n597 ), .A2(\AES_ENC/us02/n1030 ), .ZN(\AES_ENC/us02/n1049 ) );
NAND2_X2 \AES_ENC/us02/U511  ( .A1(\AES_ENC/us02/n1049 ), .A2(\AES_ENC/us02/n794 ), .ZN(\AES_ENC/us02/n637 ) );
AND2_X2 \AES_ENC/us02/U493  ( .A1(\AES_ENC/us02/n779 ), .A2(\AES_ENC/us02/n996 ), .ZN(\AES_ENC/us02/n632 ) );
NAND4_X2 \AES_ENC/us02/U485  ( .A1(\AES_ENC/us02/n637 ), .A2(\AES_ENC/us02/n636 ), .A3(\AES_ENC/us02/n635 ), .A4(\AES_ENC/us02/n634 ), .ZN(\AES_ENC/us02/n638 ) );
NAND2_X2 \AES_ENC/us02/U484  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n638 ), .ZN(\AES_ENC/us02/n679 ) );
NAND2_X2 \AES_ENC/us02/U481  ( .A1(\AES_ENC/us02/n1094 ), .A2(\AES_ENC/us02/n591 ), .ZN(\AES_ENC/us02/n648 ) );
NAND2_X2 \AES_ENC/us02/U476  ( .A1(\AES_ENC/us02/n601 ), .A2(\AES_ENC/us02/n590 ), .ZN(\AES_ENC/us02/n762 ) );
NAND2_X2 \AES_ENC/us02/U475  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n762 ), .ZN(\AES_ENC/us02/n647 ) );
NAND4_X2 \AES_ENC/us02/U457  ( .A1(\AES_ENC/us02/n648 ), .A2(\AES_ENC/us02/n647 ), .A3(\AES_ENC/us02/n646 ), .A4(\AES_ENC/us02/n645 ), .ZN(\AES_ENC/us02/n649 ) );
NAND2_X2 \AES_ENC/us02/U456  ( .A1(\AES_ENC/sa02 [0]), .A2(\AES_ENC/us02/n649 ), .ZN(\AES_ENC/us02/n665 ) );
NAND2_X2 \AES_ENC/us02/U454  ( .A1(\AES_ENC/us02/n596 ), .A2(\AES_ENC/us02/n623 ), .ZN(\AES_ENC/us02/n855 ) );
NAND2_X2 \AES_ENC/us02/U453  ( .A1(\AES_ENC/us02/n587 ), .A2(\AES_ENC/us02/n855 ), .ZN(\AES_ENC/us02/n821 ) );
NAND2_X2 \AES_ENC/us02/U452  ( .A1(\AES_ENC/us02/n1093 ), .A2(\AES_ENC/us02/n821 ), .ZN(\AES_ENC/us02/n662 ) );
NAND2_X2 \AES_ENC/us02/U451  ( .A1(\AES_ENC/us02/n619 ), .A2(\AES_ENC/us02/n589 ), .ZN(\AES_ENC/us02/n650 ) );
NAND2_X2 \AES_ENC/us02/U450  ( .A1(\AES_ENC/us02/n956 ), .A2(\AES_ENC/us02/n650 ), .ZN(\AES_ENC/us02/n661 ) );
NAND2_X2 \AES_ENC/us02/U449  ( .A1(\AES_ENC/us02/n626 ), .A2(\AES_ENC/us02/n627 ), .ZN(\AES_ENC/us02/n839 ) );
OR2_X2 \AES_ENC/us02/U446  ( .A1(\AES_ENC/us02/n839 ), .A2(\AES_ENC/us02/n932 ), .ZN(\AES_ENC/us02/n656 ) );
NAND2_X2 \AES_ENC/us02/U445  ( .A1(\AES_ENC/us02/n621 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n1096 ) );
NAND2_X2 \AES_ENC/us02/U444  ( .A1(\AES_ENC/us02/n1030 ), .A2(\AES_ENC/us02/n1096 ), .ZN(\AES_ENC/us02/n651 ) );
NAND2_X2 \AES_ENC/us02/U443  ( .A1(\AES_ENC/us02/n1114 ), .A2(\AES_ENC/us02/n651 ), .ZN(\AES_ENC/us02/n655 ) );
OR3_X2 \AES_ENC/us02/U440  ( .A1(\AES_ENC/us02/n1079 ), .A2(\AES_ENC/sa02 [7]), .A3(\AES_ENC/us02/n626 ), .ZN(\AES_ENC/us02/n654 ));
NAND2_X2 \AES_ENC/us02/U439  ( .A1(\AES_ENC/us02/n593 ), .A2(\AES_ENC/us02/n601 ), .ZN(\AES_ENC/us02/n652 ) );
NAND4_X2 \AES_ENC/us02/U437  ( .A1(\AES_ENC/us02/n656 ), .A2(\AES_ENC/us02/n655 ), .A3(\AES_ENC/us02/n654 ), .A4(\AES_ENC/us02/n653 ), .ZN(\AES_ENC/us02/n657 ) );
NAND2_X2 \AES_ENC/us02/U436  ( .A1(\AES_ENC/sa02 [2]), .A2(\AES_ENC/us02/n657 ), .ZN(\AES_ENC/us02/n660 ) );
NAND4_X2 \AES_ENC/us02/U432  ( .A1(\AES_ENC/us02/n662 ), .A2(\AES_ENC/us02/n661 ), .A3(\AES_ENC/us02/n660 ), .A4(\AES_ENC/us02/n659 ), .ZN(\AES_ENC/us02/n663 ) );
NAND2_X2 \AES_ENC/us02/U431  ( .A1(\AES_ENC/us02/n663 ), .A2(\AES_ENC/us02/n574 ), .ZN(\AES_ENC/us02/n664 ) );
NAND2_X2 \AES_ENC/us02/U430  ( .A1(\AES_ENC/us02/n665 ), .A2(\AES_ENC/us02/n664 ), .ZN(\AES_ENC/us02/n666 ) );
NAND2_X2 \AES_ENC/us02/U429  ( .A1(\AES_ENC/sa02 [6]), .A2(\AES_ENC/us02/n666 ), .ZN(\AES_ENC/us02/n678 ) );
NAND2_X2 \AES_ENC/us02/U426  ( .A1(\AES_ENC/us02/n735 ), .A2(\AES_ENC/us02/n1093 ), .ZN(\AES_ENC/us02/n675 ) );
NAND2_X2 \AES_ENC/us02/U425  ( .A1(\AES_ENC/us02/n588 ), .A2(\AES_ENC/us02/n597 ), .ZN(\AES_ENC/us02/n1045 ) );
OR2_X2 \AES_ENC/us02/U424  ( .A1(\AES_ENC/us02/n1045 ), .A2(\AES_ENC/us02/n605 ), .ZN(\AES_ENC/us02/n674 ) );
NAND2_X2 \AES_ENC/us02/U423  ( .A1(\AES_ENC/sa02 [1]), .A2(\AES_ENC/us02/n620 ), .ZN(\AES_ENC/us02/n667 ) );
NAND2_X2 \AES_ENC/us02/U422  ( .A1(\AES_ENC/us02/n619 ), .A2(\AES_ENC/us02/n667 ), .ZN(\AES_ENC/us02/n1071 ) );
NAND4_X2 \AES_ENC/us02/U412  ( .A1(\AES_ENC/us02/n675 ), .A2(\AES_ENC/us02/n674 ), .A3(\AES_ENC/us02/n673 ), .A4(\AES_ENC/us02/n672 ), .ZN(\AES_ENC/us02/n676 ) );
NAND2_X2 \AES_ENC/us02/U411  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n676 ), .ZN(\AES_ENC/us02/n677 ) );
NAND2_X2 \AES_ENC/us02/U408  ( .A1(\AES_ENC/us02/n800 ), .A2(\AES_ENC/us02/n1022 ), .ZN(\AES_ENC/us02/n680 ) );
NAND2_X2 \AES_ENC/us02/U407  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n680 ), .ZN(\AES_ENC/us02/n681 ) );
AND2_X2 \AES_ENC/us02/U402  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n684 ), .ZN(\AES_ENC/us02/n682 ) );
NAND4_X2 \AES_ENC/us02/U395  ( .A1(\AES_ENC/us02/n691 ), .A2(\AES_ENC/us02/n581 ), .A3(\AES_ENC/us02/n690 ), .A4(\AES_ENC/us02/n689 ), .ZN(\AES_ENC/us02/n692 ) );
NAND2_X2 \AES_ENC/us02/U394  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n692 ), .ZN(\AES_ENC/us02/n733 ) );
NAND2_X2 \AES_ENC/us02/U392  ( .A1(\AES_ENC/us02/n977 ), .A2(\AES_ENC/us02/n1050 ), .ZN(\AES_ENC/us02/n702 ) );
NAND2_X2 \AES_ENC/us02/U391  ( .A1(\AES_ENC/us02/n1093 ), .A2(\AES_ENC/us02/n1045 ), .ZN(\AES_ENC/us02/n701 ) );
NAND4_X2 \AES_ENC/us02/U381  ( .A1(\AES_ENC/us02/n702 ), .A2(\AES_ENC/us02/n701 ), .A3(\AES_ENC/us02/n700 ), .A4(\AES_ENC/us02/n699 ), .ZN(\AES_ENC/us02/n703 ) );
NAND2_X2 \AES_ENC/us02/U380  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n703 ), .ZN(\AES_ENC/us02/n732 ) );
AND2_X2 \AES_ENC/us02/U379  ( .A1(\AES_ENC/sa02 [0]), .A2(\AES_ENC/sa02 [6]),.ZN(\AES_ENC/us02/n1113 ) );
NAND2_X2 \AES_ENC/us02/U378  ( .A1(\AES_ENC/us02/n601 ), .A2(\AES_ENC/us02/n1030 ), .ZN(\AES_ENC/us02/n881 ) );
NAND2_X2 \AES_ENC/us02/U377  ( .A1(\AES_ENC/us02/n1093 ), .A2(\AES_ENC/us02/n881 ), .ZN(\AES_ENC/us02/n715 ) );
NAND2_X2 \AES_ENC/us02/U376  ( .A1(\AES_ENC/us02/n1010 ), .A2(\AES_ENC/us02/n600 ), .ZN(\AES_ENC/us02/n714 ) );
NAND2_X2 \AES_ENC/us02/U375  ( .A1(\AES_ENC/us02/n855 ), .A2(\AES_ENC/us02/n588 ), .ZN(\AES_ENC/us02/n1117 ) );
XNOR2_X2 \AES_ENC/us02/U371  ( .A(\AES_ENC/us02/n611 ), .B(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n824 ) );
NAND4_X2 \AES_ENC/us02/U362  ( .A1(\AES_ENC/us02/n715 ), .A2(\AES_ENC/us02/n714 ), .A3(\AES_ENC/us02/n713 ), .A4(\AES_ENC/us02/n712 ), .ZN(\AES_ENC/us02/n716 ) );
NAND2_X2 \AES_ENC/us02/U361  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n716 ), .ZN(\AES_ENC/us02/n731 ) );
AND2_X2 \AES_ENC/us02/U360  ( .A1(\AES_ENC/sa02 [6]), .A2(\AES_ENC/us02/n574 ), .ZN(\AES_ENC/us02/n1131 ) );
NAND2_X2 \AES_ENC/us02/U359  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n717 ) );
NAND2_X2 \AES_ENC/us02/U358  ( .A1(\AES_ENC/us02/n1029 ), .A2(\AES_ENC/us02/n717 ), .ZN(\AES_ENC/us02/n728 ) );
NAND2_X2 \AES_ENC/us02/U357  ( .A1(\AES_ENC/sa02 [1]), .A2(\AES_ENC/us02/n624 ), .ZN(\AES_ENC/us02/n1097 ) );
NAND2_X2 \AES_ENC/us02/U356  ( .A1(\AES_ENC/us02/n603 ), .A2(\AES_ENC/us02/n1097 ), .ZN(\AES_ENC/us02/n718 ) );
NAND2_X2 \AES_ENC/us02/U355  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n718 ), .ZN(\AES_ENC/us02/n727 ) );
NAND4_X2 \AES_ENC/us02/U344  ( .A1(\AES_ENC/us02/n728 ), .A2(\AES_ENC/us02/n727 ), .A3(\AES_ENC/us02/n726 ), .A4(\AES_ENC/us02/n725 ), .ZN(\AES_ENC/us02/n729 ) );
NAND2_X2 \AES_ENC/us02/U343  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n729 ), .ZN(\AES_ENC/us02/n730 ) );
NAND4_X2 \AES_ENC/us02/U342  ( .A1(\AES_ENC/us02/n733 ), .A2(\AES_ENC/us02/n732 ), .A3(\AES_ENC/us02/n731 ), .A4(\AES_ENC/us02/n730 ), .ZN(\AES_ENC/sa02_sub[1] ) );
NAND2_X2 \AES_ENC/us02/U341  ( .A1(\AES_ENC/sa02 [7]), .A2(\AES_ENC/us02/n611 ), .ZN(\AES_ENC/us02/n734 ) );
NAND2_X2 \AES_ENC/us02/U340  ( .A1(\AES_ENC/us02/n734 ), .A2(\AES_ENC/us02/n607 ), .ZN(\AES_ENC/us02/n738 ) );
OR4_X2 \AES_ENC/us02/U339  ( .A1(\AES_ENC/us02/n738 ), .A2(\AES_ENC/us02/n626 ), .A3(\AES_ENC/us02/n826 ), .A4(\AES_ENC/us02/n1121 ), .ZN(\AES_ENC/us02/n746 ) );
NAND2_X2 \AES_ENC/us02/U337  ( .A1(\AES_ENC/us02/n1100 ), .A2(\AES_ENC/us02/n587 ), .ZN(\AES_ENC/us02/n992 ) );
OR2_X2 \AES_ENC/us02/U336  ( .A1(\AES_ENC/us02/n610 ), .A2(\AES_ENC/us02/n735 ), .ZN(\AES_ENC/us02/n737 ) );
NAND2_X2 \AES_ENC/us02/U334  ( .A1(\AES_ENC/us02/n619 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n753 ) );
NAND2_X2 \AES_ENC/us02/U333  ( .A1(\AES_ENC/us02/n582 ), .A2(\AES_ENC/us02/n753 ), .ZN(\AES_ENC/us02/n1080 ) );
NAND2_X2 \AES_ENC/us02/U332  ( .A1(\AES_ENC/us02/n1048 ), .A2(\AES_ENC/us02/n576 ), .ZN(\AES_ENC/us02/n736 ) );
NAND2_X2 \AES_ENC/us02/U331  ( .A1(\AES_ENC/us02/n737 ), .A2(\AES_ENC/us02/n736 ), .ZN(\AES_ENC/us02/n739 ) );
NAND2_X2 \AES_ENC/us02/U330  ( .A1(\AES_ENC/us02/n739 ), .A2(\AES_ENC/us02/n738 ), .ZN(\AES_ENC/us02/n745 ) );
NAND2_X2 \AES_ENC/us02/U326  ( .A1(\AES_ENC/us02/n1096 ), .A2(\AES_ENC/us02/n590 ), .ZN(\AES_ENC/us02/n906 ) );
NAND4_X2 \AES_ENC/us02/U323  ( .A1(\AES_ENC/us02/n746 ), .A2(\AES_ENC/us02/n992 ), .A3(\AES_ENC/us02/n745 ), .A4(\AES_ENC/us02/n744 ), .ZN(\AES_ENC/us02/n747 ) );
NAND2_X2 \AES_ENC/us02/U322  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n747 ), .ZN(\AES_ENC/us02/n793 ) );
NAND2_X2 \AES_ENC/us02/U321  ( .A1(\AES_ENC/us02/n584 ), .A2(\AES_ENC/us02/n855 ), .ZN(\AES_ENC/us02/n748 ) );
NAND2_X2 \AES_ENC/us02/U320  ( .A1(\AES_ENC/us02/n956 ), .A2(\AES_ENC/us02/n748 ), .ZN(\AES_ENC/us02/n760 ) );
NAND2_X2 \AES_ENC/us02/U313  ( .A1(\AES_ENC/us02/n590 ), .A2(\AES_ENC/us02/n753 ), .ZN(\AES_ENC/us02/n1023 ) );
NAND4_X2 \AES_ENC/us02/U308  ( .A1(\AES_ENC/us02/n760 ), .A2(\AES_ENC/us02/n992 ), .A3(\AES_ENC/us02/n759 ), .A4(\AES_ENC/us02/n758 ), .ZN(\AES_ENC/us02/n761 ) );
NAND2_X2 \AES_ENC/us02/U307  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n761 ), .ZN(\AES_ENC/us02/n792 ) );
NAND2_X2 \AES_ENC/us02/U306  ( .A1(\AES_ENC/us02/n584 ), .A2(\AES_ENC/us02/n603 ), .ZN(\AES_ENC/us02/n989 ) );
NAND2_X2 \AES_ENC/us02/U305  ( .A1(\AES_ENC/us02/n1050 ), .A2(\AES_ENC/us02/n989 ), .ZN(\AES_ENC/us02/n777 ) );
NAND2_X2 \AES_ENC/us02/U304  ( .A1(\AES_ENC/us02/n1093 ), .A2(\AES_ENC/us02/n762 ), .ZN(\AES_ENC/us02/n776 ) );
XNOR2_X2 \AES_ENC/us02/U301  ( .A(\AES_ENC/sa02 [7]), .B(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n959 ) );
NAND4_X2 \AES_ENC/us02/U289  ( .A1(\AES_ENC/us02/n777 ), .A2(\AES_ENC/us02/n776 ), .A3(\AES_ENC/us02/n775 ), .A4(\AES_ENC/us02/n774 ), .ZN(\AES_ENC/us02/n778 ) );
NAND2_X2 \AES_ENC/us02/U288  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n778 ), .ZN(\AES_ENC/us02/n791 ) );
NAND2_X2 \AES_ENC/us02/U287  ( .A1(\AES_ENC/us02/n1056 ), .A2(\AES_ENC/us02/n1050 ), .ZN(\AES_ENC/us02/n788 ) );
NAND2_X2 \AES_ENC/us02/U286  ( .A1(\AES_ENC/us02/n1091 ), .A2(\AES_ENC/us02/n779 ), .ZN(\AES_ENC/us02/n787 ) );
NAND2_X2 \AES_ENC/us02/U285  ( .A1(\AES_ENC/us02/n956 ), .A2(\AES_ENC/sa02 [1]), .ZN(\AES_ENC/us02/n786 ) );
NAND4_X2 \AES_ENC/us02/U278  ( .A1(\AES_ENC/us02/n788 ), .A2(\AES_ENC/us02/n787 ), .A3(\AES_ENC/us02/n786 ), .A4(\AES_ENC/us02/n785 ), .ZN(\AES_ENC/us02/n789 ) );
NAND2_X2 \AES_ENC/us02/U277  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n789 ), .ZN(\AES_ENC/us02/n790 ) );
NAND4_X2 \AES_ENC/us02/U276  ( .A1(\AES_ENC/us02/n793 ), .A2(\AES_ENC/us02/n792 ), .A3(\AES_ENC/us02/n791 ), .A4(\AES_ENC/us02/n790 ), .ZN(\AES_ENC/sa02_sub[2] ) );
NAND2_X2 \AES_ENC/us02/U275  ( .A1(\AES_ENC/us02/n1059 ), .A2(\AES_ENC/us02/n794 ), .ZN(\AES_ENC/us02/n810 ) );
NAND2_X2 \AES_ENC/us02/U274  ( .A1(\AES_ENC/us02/n1049 ), .A2(\AES_ENC/us02/n956 ), .ZN(\AES_ENC/us02/n809 ) );
OR2_X2 \AES_ENC/us02/U266  ( .A1(\AES_ENC/us02/n1096 ), .A2(\AES_ENC/us02/n606 ), .ZN(\AES_ENC/us02/n802 ) );
NAND2_X2 \AES_ENC/us02/U265  ( .A1(\AES_ENC/us02/n1053 ), .A2(\AES_ENC/us02/n800 ), .ZN(\AES_ENC/us02/n801 ) );
NAND2_X2 \AES_ENC/us02/U264  ( .A1(\AES_ENC/us02/n802 ), .A2(\AES_ENC/us02/n801 ), .ZN(\AES_ENC/us02/n805 ) );
NAND4_X2 \AES_ENC/us02/U261  ( .A1(\AES_ENC/us02/n810 ), .A2(\AES_ENC/us02/n809 ), .A3(\AES_ENC/us02/n808 ), .A4(\AES_ENC/us02/n807 ), .ZN(\AES_ENC/us02/n811 ) );
NAND2_X2 \AES_ENC/us02/U260  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n811 ), .ZN(\AES_ENC/us02/n852 ) );
OR2_X2 \AES_ENC/us02/U259  ( .A1(\AES_ENC/us02/n1023 ), .A2(\AES_ENC/us02/n617 ), .ZN(\AES_ENC/us02/n819 ) );
OR2_X2 \AES_ENC/us02/U257  ( .A1(\AES_ENC/us02/n570 ), .A2(\AES_ENC/us02/n930 ), .ZN(\AES_ENC/us02/n818 ) );
NAND2_X2 \AES_ENC/us02/U256  ( .A1(\AES_ENC/us02/n1013 ), .A2(\AES_ENC/us02/n1094 ), .ZN(\AES_ENC/us02/n817 ) );
NAND4_X2 \AES_ENC/us02/U249  ( .A1(\AES_ENC/us02/n819 ), .A2(\AES_ENC/us02/n818 ), .A3(\AES_ENC/us02/n817 ), .A4(\AES_ENC/us02/n816 ), .ZN(\AES_ENC/us02/n820 ) );
NAND2_X2 \AES_ENC/us02/U248  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n820 ), .ZN(\AES_ENC/us02/n851 ) );
NAND2_X2 \AES_ENC/us02/U247  ( .A1(\AES_ENC/us02/n956 ), .A2(\AES_ENC/us02/n1080 ), .ZN(\AES_ENC/us02/n835 ) );
NAND2_X2 \AES_ENC/us02/U246  ( .A1(\AES_ENC/us02/n570 ), .A2(\AES_ENC/us02/n1030 ), .ZN(\AES_ENC/us02/n1047 ) );
OR2_X2 \AES_ENC/us02/U245  ( .A1(\AES_ENC/us02/n1047 ), .A2(\AES_ENC/us02/n612 ), .ZN(\AES_ENC/us02/n834 ) );
NAND2_X2 \AES_ENC/us02/U244  ( .A1(\AES_ENC/us02/n1072 ), .A2(\AES_ENC/us02/n589 ), .ZN(\AES_ENC/us02/n833 ) );
NAND4_X2 \AES_ENC/us02/U233  ( .A1(\AES_ENC/us02/n835 ), .A2(\AES_ENC/us02/n834 ), .A3(\AES_ENC/us02/n833 ), .A4(\AES_ENC/us02/n832 ), .ZN(\AES_ENC/us02/n836 ) );
NAND2_X2 \AES_ENC/us02/U232  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n836 ), .ZN(\AES_ENC/us02/n850 ) );
NAND2_X2 \AES_ENC/us02/U231  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n623 ), .ZN(\AES_ENC/us02/n847 ) );
NAND2_X2 \AES_ENC/us02/U230  ( .A1(\AES_ENC/us02/n1050 ), .A2(\AES_ENC/us02/n1071 ), .ZN(\AES_ENC/us02/n846 ) );
OR2_X2 \AES_ENC/us02/U224  ( .A1(\AES_ENC/us02/n1053 ), .A2(\AES_ENC/us02/n911 ), .ZN(\AES_ENC/us02/n1077 ) );
NAND4_X2 \AES_ENC/us02/U220  ( .A1(\AES_ENC/us02/n847 ), .A2(\AES_ENC/us02/n846 ), .A3(\AES_ENC/us02/n845 ), .A4(\AES_ENC/us02/n844 ), .ZN(\AES_ENC/us02/n848 ) );
NAND2_X2 \AES_ENC/us02/U219  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n848 ), .ZN(\AES_ENC/us02/n849 ) );
NAND4_X2 \AES_ENC/us02/U218  ( .A1(\AES_ENC/us02/n852 ), .A2(\AES_ENC/us02/n851 ), .A3(\AES_ENC/us02/n850 ), .A4(\AES_ENC/us02/n849 ), .ZN(\AES_ENC/sa02_sub[3] ) );
NAND2_X2 \AES_ENC/us02/U216  ( .A1(\AES_ENC/us02/n1009 ), .A2(\AES_ENC/us02/n1072 ), .ZN(\AES_ENC/us02/n862 ) );
NAND2_X2 \AES_ENC/us02/U215  ( .A1(\AES_ENC/us02/n603 ), .A2(\AES_ENC/us02/n577 ), .ZN(\AES_ENC/us02/n853 ) );
NAND2_X2 \AES_ENC/us02/U214  ( .A1(\AES_ENC/us02/n1050 ), .A2(\AES_ENC/us02/n853 ), .ZN(\AES_ENC/us02/n861 ) );
NAND4_X2 \AES_ENC/us02/U206  ( .A1(\AES_ENC/us02/n862 ), .A2(\AES_ENC/us02/n861 ), .A3(\AES_ENC/us02/n860 ), .A4(\AES_ENC/us02/n859 ), .ZN(\AES_ENC/us02/n863 ) );
NAND2_X2 \AES_ENC/us02/U205  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n863 ), .ZN(\AES_ENC/us02/n905 ) );
NAND2_X2 \AES_ENC/us02/U204  ( .A1(\AES_ENC/us02/n1010 ), .A2(\AES_ENC/us02/n989 ), .ZN(\AES_ENC/us02/n874 ) );
NAND2_X2 \AES_ENC/us02/U203  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n610 ), .ZN(\AES_ENC/us02/n864 ) );
NAND2_X2 \AES_ENC/us02/U202  ( .A1(\AES_ENC/us02/n929 ), .A2(\AES_ENC/us02/n864 ), .ZN(\AES_ENC/us02/n873 ) );
NAND4_X2 \AES_ENC/us02/U193  ( .A1(\AES_ENC/us02/n874 ), .A2(\AES_ENC/us02/n873 ), .A3(\AES_ENC/us02/n872 ), .A4(\AES_ENC/us02/n871 ), .ZN(\AES_ENC/us02/n875 ) );
NAND2_X2 \AES_ENC/us02/U192  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n875 ), .ZN(\AES_ENC/us02/n904 ) );
NAND2_X2 \AES_ENC/us02/U191  ( .A1(\AES_ENC/us02/n583 ), .A2(\AES_ENC/us02/n1050 ), .ZN(\AES_ENC/us02/n889 ) );
NAND2_X2 \AES_ENC/us02/U190  ( .A1(\AES_ENC/us02/n1093 ), .A2(\AES_ENC/us02/n587 ), .ZN(\AES_ENC/us02/n876 ) );
NAND2_X2 \AES_ENC/us02/U189  ( .A1(\AES_ENC/us02/n604 ), .A2(\AES_ENC/us02/n876 ), .ZN(\AES_ENC/us02/n877 ) );
NAND2_X2 \AES_ENC/us02/U188  ( .A1(\AES_ENC/us02/n877 ), .A2(\AES_ENC/us02/n623 ), .ZN(\AES_ENC/us02/n888 ) );
NAND4_X2 \AES_ENC/us02/U179  ( .A1(\AES_ENC/us02/n889 ), .A2(\AES_ENC/us02/n888 ), .A3(\AES_ENC/us02/n887 ), .A4(\AES_ENC/us02/n886 ), .ZN(\AES_ENC/us02/n890 ) );
NAND2_X2 \AES_ENC/us02/U178  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n890 ), .ZN(\AES_ENC/us02/n903 ) );
OR2_X2 \AES_ENC/us02/U177  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n1059 ), .ZN(\AES_ENC/us02/n900 ) );
NAND2_X2 \AES_ENC/us02/U176  ( .A1(\AES_ENC/us02/n1073 ), .A2(\AES_ENC/us02/n1047 ), .ZN(\AES_ENC/us02/n899 ) );
NAND2_X2 \AES_ENC/us02/U175  ( .A1(\AES_ENC/us02/n1094 ), .A2(\AES_ENC/us02/n595 ), .ZN(\AES_ENC/us02/n898 ) );
NAND4_X2 \AES_ENC/us02/U167  ( .A1(\AES_ENC/us02/n900 ), .A2(\AES_ENC/us02/n899 ), .A3(\AES_ENC/us02/n898 ), .A4(\AES_ENC/us02/n897 ), .ZN(\AES_ENC/us02/n901 ) );
NAND2_X2 \AES_ENC/us02/U166  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n901 ), .ZN(\AES_ENC/us02/n902 ) );
NAND4_X2 \AES_ENC/us02/U165  ( .A1(\AES_ENC/us02/n905 ), .A2(\AES_ENC/us02/n904 ), .A3(\AES_ENC/us02/n903 ), .A4(\AES_ENC/us02/n902 ), .ZN(\AES_ENC/sa02_sub[4] ) );
NAND2_X2 \AES_ENC/us02/U164  ( .A1(\AES_ENC/us02/n1094 ), .A2(\AES_ENC/us02/n599 ), .ZN(\AES_ENC/us02/n922 ) );
NAND2_X2 \AES_ENC/us02/U163  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n989 ), .ZN(\AES_ENC/us02/n921 ) );
NAND4_X2 \AES_ENC/us02/U151  ( .A1(\AES_ENC/us02/n922 ), .A2(\AES_ENC/us02/n921 ), .A3(\AES_ENC/us02/n920 ), .A4(\AES_ENC/us02/n919 ), .ZN(\AES_ENC/us02/n923 ) );
NAND2_X2 \AES_ENC/us02/U150  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n923 ), .ZN(\AES_ENC/us02/n972 ) );
NAND2_X2 \AES_ENC/us02/U149  ( .A1(\AES_ENC/us02/n582 ), .A2(\AES_ENC/us02/n619 ), .ZN(\AES_ENC/us02/n924 ) );
NAND2_X2 \AES_ENC/us02/U148  ( .A1(\AES_ENC/us02/n1073 ), .A2(\AES_ENC/us02/n924 ), .ZN(\AES_ENC/us02/n939 ) );
NAND2_X2 \AES_ENC/us02/U147  ( .A1(\AES_ENC/us02/n926 ), .A2(\AES_ENC/us02/n925 ), .ZN(\AES_ENC/us02/n927 ) );
NAND2_X2 \AES_ENC/us02/U146  ( .A1(\AES_ENC/us02/n606 ), .A2(\AES_ENC/us02/n927 ), .ZN(\AES_ENC/us02/n928 ) );
NAND2_X2 \AES_ENC/us02/U145  ( .A1(\AES_ENC/us02/n928 ), .A2(\AES_ENC/us02/n1080 ), .ZN(\AES_ENC/us02/n938 ) );
OR2_X2 \AES_ENC/us02/U144  ( .A1(\AES_ENC/us02/n1117 ), .A2(\AES_ENC/us02/n615 ), .ZN(\AES_ENC/us02/n937 ) );
NAND4_X2 \AES_ENC/us02/U139  ( .A1(\AES_ENC/us02/n939 ), .A2(\AES_ENC/us02/n938 ), .A3(\AES_ENC/us02/n937 ), .A4(\AES_ENC/us02/n936 ), .ZN(\AES_ENC/us02/n940 ) );
NAND2_X2 \AES_ENC/us02/U138  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n940 ), .ZN(\AES_ENC/us02/n971 ) );
OR2_X2 \AES_ENC/us02/U137  ( .A1(\AES_ENC/us02/n605 ), .A2(\AES_ENC/us02/n941 ), .ZN(\AES_ENC/us02/n954 ) );
NAND2_X2 \AES_ENC/us02/U136  ( .A1(\AES_ENC/us02/n1096 ), .A2(\AES_ENC/us02/n577 ), .ZN(\AES_ENC/us02/n942 ) );
NAND2_X2 \AES_ENC/us02/U135  ( .A1(\AES_ENC/us02/n1048 ), .A2(\AES_ENC/us02/n942 ), .ZN(\AES_ENC/us02/n943 ) );
NAND2_X2 \AES_ENC/us02/U134  ( .A1(\AES_ENC/us02/n612 ), .A2(\AES_ENC/us02/n943 ), .ZN(\AES_ENC/us02/n944 ) );
NAND2_X2 \AES_ENC/us02/U133  ( .A1(\AES_ENC/us02/n944 ), .A2(\AES_ENC/us02/n580 ), .ZN(\AES_ENC/us02/n953 ) );
NAND4_X2 \AES_ENC/us02/U125  ( .A1(\AES_ENC/us02/n954 ), .A2(\AES_ENC/us02/n953 ), .A3(\AES_ENC/us02/n952 ), .A4(\AES_ENC/us02/n951 ), .ZN(\AES_ENC/us02/n955 ) );
NAND2_X2 \AES_ENC/us02/U124  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n955 ), .ZN(\AES_ENC/us02/n970 ) );
NAND2_X2 \AES_ENC/us02/U123  ( .A1(\AES_ENC/us02/n1094 ), .A2(\AES_ENC/us02/n1071 ), .ZN(\AES_ENC/us02/n967 ) );
NAND2_X2 \AES_ENC/us02/U122  ( .A1(\AES_ENC/us02/n956 ), .A2(\AES_ENC/us02/n1030 ), .ZN(\AES_ENC/us02/n966 ) );
NAND4_X2 \AES_ENC/us02/U114  ( .A1(\AES_ENC/us02/n967 ), .A2(\AES_ENC/us02/n966 ), .A3(\AES_ENC/us02/n965 ), .A4(\AES_ENC/us02/n964 ), .ZN(\AES_ENC/us02/n968 ) );
NAND2_X2 \AES_ENC/us02/U113  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n968 ), .ZN(\AES_ENC/us02/n969 ) );
NAND4_X2 \AES_ENC/us02/U112  ( .A1(\AES_ENC/us02/n972 ), .A2(\AES_ENC/us02/n971 ), .A3(\AES_ENC/us02/n970 ), .A4(\AES_ENC/us02/n969 ), .ZN(\AES_ENC/sa02_sub[5] ) );
NAND2_X2 \AES_ENC/us02/U111  ( .A1(\AES_ENC/us02/n570 ), .A2(\AES_ENC/us02/n1097 ), .ZN(\AES_ENC/us02/n973 ) );
NAND2_X2 \AES_ENC/us02/U110  ( .A1(\AES_ENC/us02/n1073 ), .A2(\AES_ENC/us02/n973 ), .ZN(\AES_ENC/us02/n987 ) );
NAND2_X2 \AES_ENC/us02/U109  ( .A1(\AES_ENC/us02/n974 ), .A2(\AES_ENC/us02/n1077 ), .ZN(\AES_ENC/us02/n975 ) );
NAND2_X2 \AES_ENC/us02/U108  ( .A1(\AES_ENC/us02/n613 ), .A2(\AES_ENC/us02/n975 ), .ZN(\AES_ENC/us02/n976 ) );
NAND2_X2 \AES_ENC/us02/U107  ( .A1(\AES_ENC/us02/n977 ), .A2(\AES_ENC/us02/n976 ), .ZN(\AES_ENC/us02/n986 ) );
NAND4_X2 \AES_ENC/us02/U99  ( .A1(\AES_ENC/us02/n987 ), .A2(\AES_ENC/us02/n986 ), .A3(\AES_ENC/us02/n985 ), .A4(\AES_ENC/us02/n984 ), .ZN(\AES_ENC/us02/n988 ) );
NAND2_X2 \AES_ENC/us02/U98  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n988 ), .ZN(\AES_ENC/us02/n1044 ) );
NAND2_X2 \AES_ENC/us02/U97  ( .A1(\AES_ENC/us02/n1073 ), .A2(\AES_ENC/us02/n989 ), .ZN(\AES_ENC/us02/n1004 ) );
NAND2_X2 \AES_ENC/us02/U96  ( .A1(\AES_ENC/us02/n1092 ), .A2(\AES_ENC/us02/n619 ), .ZN(\AES_ENC/us02/n1003 ) );
NAND4_X2 \AES_ENC/us02/U85  ( .A1(\AES_ENC/us02/n1004 ), .A2(\AES_ENC/us02/n1003 ), .A3(\AES_ENC/us02/n1002 ), .A4(\AES_ENC/us02/n1001 ), .ZN(\AES_ENC/us02/n1005 ) );
NAND2_X2 \AES_ENC/us02/U84  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n1005 ), .ZN(\AES_ENC/us02/n1043 ) );
NAND2_X2 \AES_ENC/us02/U83  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n596 ), .ZN(\AES_ENC/us02/n1020 ) );
NAND2_X2 \AES_ENC/us02/U82  ( .A1(\AES_ENC/us02/n1050 ), .A2(\AES_ENC/us02/n624 ), .ZN(\AES_ENC/us02/n1019 ) );
NAND2_X2 \AES_ENC/us02/U77  ( .A1(\AES_ENC/us02/n1059 ), .A2(\AES_ENC/us02/n1114 ), .ZN(\AES_ENC/us02/n1012 ) );
NAND2_X2 \AES_ENC/us02/U76  ( .A1(\AES_ENC/us02/n1010 ), .A2(\AES_ENC/us02/n592 ), .ZN(\AES_ENC/us02/n1011 ) );
NAND2_X2 \AES_ENC/us02/U75  ( .A1(\AES_ENC/us02/n1012 ), .A2(\AES_ENC/us02/n1011 ), .ZN(\AES_ENC/us02/n1016 ) );
NAND4_X2 \AES_ENC/us02/U70  ( .A1(\AES_ENC/us02/n1020 ), .A2(\AES_ENC/us02/n1019 ), .A3(\AES_ENC/us02/n1018 ), .A4(\AES_ENC/us02/n1017 ), .ZN(\AES_ENC/us02/n1021 ) );
NAND2_X2 \AES_ENC/us02/U69  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n1021 ), .ZN(\AES_ENC/us02/n1042 ) );
NAND2_X2 \AES_ENC/us02/U68  ( .A1(\AES_ENC/us02/n1022 ), .A2(\AES_ENC/us02/n1093 ), .ZN(\AES_ENC/us02/n1039 ) );
NAND2_X2 \AES_ENC/us02/U67  ( .A1(\AES_ENC/us02/n1050 ), .A2(\AES_ENC/us02/n1023 ), .ZN(\AES_ENC/us02/n1038 ) );
NAND2_X2 \AES_ENC/us02/U66  ( .A1(\AES_ENC/us02/n1024 ), .A2(\AES_ENC/us02/n1071 ), .ZN(\AES_ENC/us02/n1037 ) );
AND2_X2 \AES_ENC/us02/U60  ( .A1(\AES_ENC/us02/n1030 ), .A2(\AES_ENC/us02/n602 ), .ZN(\AES_ENC/us02/n1078 ) );
NAND4_X2 \AES_ENC/us02/U56  ( .A1(\AES_ENC/us02/n1039 ), .A2(\AES_ENC/us02/n1038 ), .A3(\AES_ENC/us02/n1037 ), .A4(\AES_ENC/us02/n1036 ), .ZN(\AES_ENC/us02/n1040 ) );
NAND2_X2 \AES_ENC/us02/U55  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n1040 ), .ZN(\AES_ENC/us02/n1041 ) );
NAND4_X2 \AES_ENC/us02/U54  ( .A1(\AES_ENC/us02/n1044 ), .A2(\AES_ENC/us02/n1043 ), .A3(\AES_ENC/us02/n1042 ), .A4(\AES_ENC/us02/n1041 ), .ZN(\AES_ENC/sa02_sub[6] ) );
NAND2_X2 \AES_ENC/us02/U53  ( .A1(\AES_ENC/us02/n1072 ), .A2(\AES_ENC/us02/n1045 ), .ZN(\AES_ENC/us02/n1068 ) );
NAND2_X2 \AES_ENC/us02/U52  ( .A1(\AES_ENC/us02/n1046 ), .A2(\AES_ENC/us02/n582 ), .ZN(\AES_ENC/us02/n1067 ) );
NAND2_X2 \AES_ENC/us02/U51  ( .A1(\AES_ENC/us02/n1094 ), .A2(\AES_ENC/us02/n1047 ), .ZN(\AES_ENC/us02/n1066 ) );
NAND4_X2 \AES_ENC/us02/U40  ( .A1(\AES_ENC/us02/n1068 ), .A2(\AES_ENC/us02/n1067 ), .A3(\AES_ENC/us02/n1066 ), .A4(\AES_ENC/us02/n1065 ), .ZN(\AES_ENC/us02/n1069 ) );
NAND2_X2 \AES_ENC/us02/U39  ( .A1(\AES_ENC/us02/n1070 ), .A2(\AES_ENC/us02/n1069 ), .ZN(\AES_ENC/us02/n1135 ) );
NAND2_X2 \AES_ENC/us02/U38  ( .A1(\AES_ENC/us02/n1072 ), .A2(\AES_ENC/us02/n1071 ), .ZN(\AES_ENC/us02/n1088 ) );
NAND2_X2 \AES_ENC/us02/U37  ( .A1(\AES_ENC/us02/n1073 ), .A2(\AES_ENC/us02/n595 ), .ZN(\AES_ENC/us02/n1087 ) );
NAND4_X2 \AES_ENC/us02/U28  ( .A1(\AES_ENC/us02/n1088 ), .A2(\AES_ENC/us02/n1087 ), .A3(\AES_ENC/us02/n1086 ), .A4(\AES_ENC/us02/n1085 ), .ZN(\AES_ENC/us02/n1089 ) );
NAND2_X2 \AES_ENC/us02/U27  ( .A1(\AES_ENC/us02/n1090 ), .A2(\AES_ENC/us02/n1089 ), .ZN(\AES_ENC/us02/n1134 ) );
NAND2_X2 \AES_ENC/us02/U26  ( .A1(\AES_ENC/us02/n1091 ), .A2(\AES_ENC/us02/n1093 ), .ZN(\AES_ENC/us02/n1111 ) );
NAND2_X2 \AES_ENC/us02/U25  ( .A1(\AES_ENC/us02/n1092 ), .A2(\AES_ENC/us02/n1120 ), .ZN(\AES_ENC/us02/n1110 ) );
AND2_X2 \AES_ENC/us02/U22  ( .A1(\AES_ENC/us02/n1097 ), .A2(\AES_ENC/us02/n1096 ), .ZN(\AES_ENC/us02/n1098 ) );
NAND4_X2 \AES_ENC/us02/U14  ( .A1(\AES_ENC/us02/n1111 ), .A2(\AES_ENC/us02/n1110 ), .A3(\AES_ENC/us02/n1109 ), .A4(\AES_ENC/us02/n1108 ), .ZN(\AES_ENC/us02/n1112 ) );
NAND2_X2 \AES_ENC/us02/U13  ( .A1(\AES_ENC/us02/n1113 ), .A2(\AES_ENC/us02/n1112 ), .ZN(\AES_ENC/us02/n1133 ) );
NAND2_X2 \AES_ENC/us02/U12  ( .A1(\AES_ENC/us02/n1115 ), .A2(\AES_ENC/us02/n1114 ), .ZN(\AES_ENC/us02/n1129 ) );
OR2_X2 \AES_ENC/us02/U11  ( .A1(\AES_ENC/us02/n608 ), .A2(\AES_ENC/us02/n1116 ), .ZN(\AES_ENC/us02/n1128 ) );
NAND4_X2 \AES_ENC/us02/U3  ( .A1(\AES_ENC/us02/n1129 ), .A2(\AES_ENC/us02/n1128 ), .A3(\AES_ENC/us02/n1127 ), .A4(\AES_ENC/us02/n1126 ), .ZN(\AES_ENC/us02/n1130 ) );
NAND2_X2 \AES_ENC/us02/U2  ( .A1(\AES_ENC/us02/n1131 ), .A2(\AES_ENC/us02/n1130 ), .ZN(\AES_ENC/us02/n1132 ) );
NAND4_X2 \AES_ENC/us02/U1  ( .A1(\AES_ENC/us02/n1135 ), .A2(\AES_ENC/us02/n1134 ), .A3(\AES_ENC/us02/n1133 ), .A4(\AES_ENC/us02/n1132 ), .ZN(\AES_ENC/sa02_sub[7] ) );
INV_X4 \AES_ENC/us03/U575  ( .A(\AES_ENC/sa03 [4]), .ZN(\AES_ENC/us03/n626 ));
INV_X4 \AES_ENC/us03/U574  ( .A(\AES_ENC/us03/n1025 ), .ZN(\AES_ENC/us03/n624 ) );
INV_X4 \AES_ENC/us03/U573  ( .A(\AES_ENC/us03/n1120 ), .ZN(\AES_ENC/us03/n622 ) );
INV_X4 \AES_ENC/us03/U572  ( .A(\AES_ENC/us03/n1121 ), .ZN(\AES_ENC/us03/n621 ) );
INV_X4 \AES_ENC/us03/U571  ( .A(\AES_ENC/us03/n1048 ), .ZN(\AES_ENC/us03/n620 ) );
INV_X4 \AES_ENC/us03/U570  ( .A(\AES_ENC/us03/n974 ), .ZN(\AES_ENC/us03/n619 ) );
INV_X4 \AES_ENC/us03/U569  ( .A(\AES_ENC/sa03 [2]), .ZN(\AES_ENC/us03/n618 ));
INV_X4 \AES_ENC/us03/U568  ( .A(\AES_ENC/us03/n800 ), .ZN(\AES_ENC/us03/n617 ) );
INV_X4 \AES_ENC/us03/U567  ( .A(\AES_ENC/us03/n925 ), .ZN(\AES_ENC/us03/n616 ) );
INV_X4 \AES_ENC/us03/U566  ( .A(\AES_ENC/us03/n1022 ), .ZN(\AES_ENC/us03/n615 ) );
INV_X4 \AES_ENC/us03/U565  ( .A(\AES_ENC/us03/n1102 ), .ZN(\AES_ENC/us03/n614 ) );
INV_X4 \AES_ENC/us03/U564  ( .A(\AES_ENC/us03/n929 ), .ZN(\AES_ENC/us03/n613 ) );
INV_X4 \AES_ENC/us03/U563  ( .A(\AES_ENC/us03/n1056 ), .ZN(\AES_ENC/us03/n612 ) );
INV_X4 \AES_ENC/us03/U562  ( .A(\AES_ENC/us03/n1054 ), .ZN(\AES_ENC/us03/n611 ) );
INV_X4 \AES_ENC/us03/U561  ( .A(\AES_ENC/us03/n881 ), .ZN(\AES_ENC/us03/n610 ) );
INV_X4 \AES_ENC/us03/U560  ( .A(\AES_ENC/us03/n926 ), .ZN(\AES_ENC/us03/n609 ) );
INV_X4 \AES_ENC/us03/U559  ( .A(\AES_ENC/us03/n977 ), .ZN(\AES_ENC/us03/n607 ) );
INV_X4 \AES_ENC/us03/U558  ( .A(\AES_ENC/us03/n1031 ), .ZN(\AES_ENC/us03/n606 ) );
INV_X4 \AES_ENC/us03/U557  ( .A(\AES_ENC/us03/n1103 ), .ZN(\AES_ENC/us03/n605 ) );
INV_X4 \AES_ENC/us03/U556  ( .A(\AES_ENC/us03/n1009 ), .ZN(\AES_ENC/us03/n604 ) );
INV_X4 \AES_ENC/us03/U555  ( .A(\AES_ENC/us03/n990 ), .ZN(\AES_ENC/us03/n603 ) );
INV_X4 \AES_ENC/us03/U554  ( .A(\AES_ENC/us03/n1058 ), .ZN(\AES_ENC/us03/n602 ) );
INV_X4 \AES_ENC/us03/U553  ( .A(\AES_ENC/us03/n1074 ), .ZN(\AES_ENC/us03/n601 ) );
INV_X4 \AES_ENC/us03/U552  ( .A(\AES_ENC/us03/n1053 ), .ZN(\AES_ENC/us03/n600 ) );
INV_X4 \AES_ENC/us03/U551  ( .A(\AES_ENC/us03/n826 ), .ZN(\AES_ENC/us03/n599 ) );
INV_X4 \AES_ENC/us03/U550  ( .A(\AES_ENC/us03/n821 ), .ZN(\AES_ENC/us03/n598 ) );
INV_X4 \AES_ENC/us03/U549  ( .A(\AES_ENC/us03/n910 ), .ZN(\AES_ENC/us03/n597 ) );
INV_X4 \AES_ENC/us03/U548  ( .A(\AES_ENC/us03/n906 ), .ZN(\AES_ENC/us03/n596 ) );
INV_X4 \AES_ENC/us03/U547  ( .A(\AES_ENC/us03/n1013 ), .ZN(\AES_ENC/us03/n594 ) );
INV_X4 \AES_ENC/us03/U546  ( .A(\AES_ENC/us03/n824 ), .ZN(\AES_ENC/us03/n593 ) );
INV_X4 \AES_ENC/us03/U545  ( .A(\AES_ENC/us03/n1091 ), .ZN(\AES_ENC/us03/n592 ) );
INV_X4 \AES_ENC/us03/U544  ( .A(\AES_ENC/us03/n1080 ), .ZN(\AES_ENC/us03/n591 ) );
INV_X4 \AES_ENC/us03/U543  ( .A(\AES_ENC/us03/n959 ), .ZN(\AES_ENC/us03/n590 ) );
INV_X4 \AES_ENC/us03/U542  ( .A(\AES_ENC/us03/n779 ), .ZN(\AES_ENC/us03/n589 ) );
INV_X4 \AES_ENC/us03/U541  ( .A(\AES_ENC/us03/n794 ), .ZN(\AES_ENC/us03/n586 ) );
INV_X4 \AES_ENC/us03/U540  ( .A(\AES_ENC/us03/n880 ), .ZN(\AES_ENC/us03/n584 ) );
INV_X4 \AES_ENC/us03/U539  ( .A(\AES_ENC/sa03 [7]), .ZN(\AES_ENC/us03/n582 ));
INV_X4 \AES_ENC/us03/U538  ( .A(\AES_ENC/us03/n992 ), .ZN(\AES_ENC/us03/n579 ) );
INV_X4 \AES_ENC/us03/U537  ( .A(\AES_ENC/us03/n1114 ), .ZN(\AES_ENC/us03/n578 ) );
INV_X4 \AES_ENC/us03/U536  ( .A(\AES_ENC/us03/n1092 ), .ZN(\AES_ENC/us03/n575 ) );
INV_X4 \AES_ENC/us03/U535  ( .A(\AES_ENC/sa03 [0]), .ZN(\AES_ENC/us03/n574 ));
NOR2_X2 \AES_ENC/us03/U534  ( .A1(\AES_ENC/sa03 [0]), .A2(\AES_ENC/sa03 [6]),.ZN(\AES_ENC/us03/n1090 ) );
NOR2_X2 \AES_ENC/us03/U533  ( .A1(\AES_ENC/us03/n574 ), .A2(\AES_ENC/sa03 [6]), .ZN(\AES_ENC/us03/n1070 ) );
NOR2_X2 \AES_ENC/us03/U532  ( .A1(\AES_ENC/sa03 [4]), .A2(\AES_ENC/sa03 [3]),.ZN(\AES_ENC/us03/n1025 ) );
INV_X4 \AES_ENC/us03/U531  ( .A(\AES_ENC/us03/n569 ), .ZN(\AES_ENC/us03/n572 ) );
NOR2_X2 \AES_ENC/us03/U530  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n765 ) );
NOR2_X2 \AES_ENC/us03/U529  ( .A1(\AES_ENC/sa03 [4]), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n764 ) );
NOR2_X2 \AES_ENC/us03/U528  ( .A1(\AES_ENC/us03/n765 ), .A2(\AES_ENC/us03/n764 ), .ZN(\AES_ENC/us03/n766 ) );
NOR2_X2 \AES_ENC/us03/U527  ( .A1(\AES_ENC/us03/n766 ), .A2(\AES_ENC/us03/n590 ), .ZN(\AES_ENC/us03/n767 ) );
NOR3_X2 \AES_ENC/us03/U526  ( .A1(\AES_ENC/us03/n582 ), .A2(\AES_ENC/sa03 [5]), .A3(\AES_ENC/us03/n704 ), .ZN(\AES_ENC/us03/n706 ));
NOR2_X2 \AES_ENC/us03/U525  ( .A1(\AES_ENC/us03/n1117 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n707 ) );
NOR2_X2 \AES_ENC/us03/U524  ( .A1(\AES_ENC/sa03 [4]), .A2(\AES_ENC/us03/n575 ), .ZN(\AES_ENC/us03/n705 ) );
NOR3_X2 \AES_ENC/us03/U523  ( .A1(\AES_ENC/us03/n707 ), .A2(\AES_ENC/us03/n706 ), .A3(\AES_ENC/us03/n705 ), .ZN(\AES_ENC/us03/n713 ) );
INV_X4 \AES_ENC/us03/U522  ( .A(\AES_ENC/sa03 [3]), .ZN(\AES_ENC/us03/n623 ));
NAND3_X2 \AES_ENC/us03/U521  ( .A1(\AES_ENC/us03/n652 ), .A2(\AES_ENC/us03/n627 ), .A3(\AES_ENC/sa03 [7]), .ZN(\AES_ENC/us03/n653 ));
NOR2_X2 \AES_ENC/us03/U520  ( .A1(\AES_ENC/us03/n618 ), .A2(\AES_ENC/sa03 [5]), .ZN(\AES_ENC/us03/n925 ) );
NOR2_X2 \AES_ENC/us03/U519  ( .A1(\AES_ENC/sa03 [5]), .A2(\AES_ENC/sa03 [2]),.ZN(\AES_ENC/us03/n974 ) );
INV_X4 \AES_ENC/us03/U518  ( .A(\AES_ENC/sa03 [5]), .ZN(\AES_ENC/us03/n627 ));
NOR2_X2 \AES_ENC/us03/U517  ( .A1(\AES_ENC/us03/n618 ), .A2(\AES_ENC/sa03 [7]), .ZN(\AES_ENC/us03/n779 ) );
NAND3_X2 \AES_ENC/us03/U516  ( .A1(\AES_ENC/us03/n679 ), .A2(\AES_ENC/us03/n678 ), .A3(\AES_ENC/us03/n677 ), .ZN(\AES_ENC/sa03_sub[0] ) );
NOR2_X2 \AES_ENC/us03/U515  ( .A1(\AES_ENC/us03/n627 ), .A2(\AES_ENC/sa03 [2]), .ZN(\AES_ENC/us03/n1048 ) );
NOR4_X2 \AES_ENC/us03/U512  ( .A1(\AES_ENC/us03/n633 ), .A2(\AES_ENC/us03/n632 ), .A3(\AES_ENC/us03/n631 ), .A4(\AES_ENC/us03/n630 ), .ZN(\AES_ENC/us03/n634 ) );
NOR2_X2 \AES_ENC/us03/U510  ( .A1(\AES_ENC/us03/n629 ), .A2(\AES_ENC/us03/n628 ), .ZN(\AES_ENC/us03/n635 ) );
NAND3_X2 \AES_ENC/us03/U509  ( .A1(\AES_ENC/sa03 [2]), .A2(\AES_ENC/sa03 [7]), .A3(\AES_ENC/us03/n1059 ), .ZN(\AES_ENC/us03/n636 ) );
NOR2_X2 \AES_ENC/us03/U508  ( .A1(\AES_ENC/sa03 [7]), .A2(\AES_ENC/sa03 [2]),.ZN(\AES_ENC/us03/n794 ) );
NOR2_X2 \AES_ENC/us03/U507  ( .A1(\AES_ENC/sa03 [4]), .A2(\AES_ENC/sa03 [1]),.ZN(\AES_ENC/us03/n1102 ) );
NOR2_X2 \AES_ENC/us03/U506  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/sa03 [3]), .ZN(\AES_ENC/us03/n1053 ) );
NOR2_X2 \AES_ENC/us03/U505  ( .A1(\AES_ENC/us03/n589 ), .A2(\AES_ENC/sa03 [5]), .ZN(\AES_ENC/us03/n1024 ) );
NOR2_X2 \AES_ENC/us03/U504  ( .A1(\AES_ENC/us03/n578 ), .A2(\AES_ENC/sa03 [2]), .ZN(\AES_ENC/us03/n1093 ) );
NOR2_X2 \AES_ENC/us03/U503  ( .A1(\AES_ENC/us03/n586 ), .A2(\AES_ENC/sa03 [5]), .ZN(\AES_ENC/us03/n1094 ) );
NOR2_X2 \AES_ENC/us03/U502  ( .A1(\AES_ENC/us03/n626 ), .A2(\AES_ENC/sa03 [3]), .ZN(\AES_ENC/us03/n931 ) );
INV_X4 \AES_ENC/us03/U501  ( .A(\AES_ENC/us03/n570 ), .ZN(\AES_ENC/us03/n573 ) );
NOR2_X2 \AES_ENC/us03/U500  ( .A1(\AES_ENC/us03/n1053 ), .A2(\AES_ENC/us03/n1095 ), .ZN(\AES_ENC/us03/n639 ) );
NOR3_X2 \AES_ENC/us03/U499  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n573 ), .A3(\AES_ENC/us03/n1074 ), .ZN(\AES_ENC/us03/n641 ) );
NOR2_X2 \AES_ENC/us03/U498  ( .A1(\AES_ENC/us03/n639 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n640 ) );
NOR2_X2 \AES_ENC/us03/U497  ( .A1(\AES_ENC/us03/n641 ), .A2(\AES_ENC/us03/n640 ), .ZN(\AES_ENC/us03/n646 ) );
NOR3_X2 \AES_ENC/us03/U496  ( .A1(\AES_ENC/us03/n995 ), .A2(\AES_ENC/us03/n579 ), .A3(\AES_ENC/us03/n994 ), .ZN(\AES_ENC/us03/n1002 ) );
NOR2_X2 \AES_ENC/us03/U495  ( .A1(\AES_ENC/us03/n909 ), .A2(\AES_ENC/us03/n908 ), .ZN(\AES_ENC/us03/n920 ) );
NOR2_X2 \AES_ENC/us03/U494  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n823 ) );
NOR2_X2 \AES_ENC/us03/U492  ( .A1(\AES_ENC/us03/n626 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n822 ) );
NOR2_X2 \AES_ENC/us03/U491  ( .A1(\AES_ENC/us03/n823 ), .A2(\AES_ENC/us03/n822 ), .ZN(\AES_ENC/us03/n825 ) );
NOR2_X2 \AES_ENC/us03/U490  ( .A1(\AES_ENC/sa03 [1]), .A2(\AES_ENC/us03/n625 ), .ZN(\AES_ENC/us03/n913 ) );
NOR2_X2 \AES_ENC/us03/U489  ( .A1(\AES_ENC/us03/n913 ), .A2(\AES_ENC/us03/n1091 ), .ZN(\AES_ENC/us03/n914 ) );
NOR2_X2 \AES_ENC/us03/U488  ( .A1(\AES_ENC/us03/n826 ), .A2(\AES_ENC/us03/n572 ), .ZN(\AES_ENC/us03/n827 ) );
NOR3_X2 \AES_ENC/us03/U487  ( .A1(\AES_ENC/us03/n769 ), .A2(\AES_ENC/us03/n768 ), .A3(\AES_ENC/us03/n767 ), .ZN(\AES_ENC/us03/n775 ) );
NOR2_X2 \AES_ENC/us03/U486  ( .A1(\AES_ENC/us03/n1056 ), .A2(\AES_ENC/us03/n1053 ), .ZN(\AES_ENC/us03/n749 ) );
NOR2_X2 \AES_ENC/us03/U483  ( .A1(\AES_ENC/us03/n749 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n752 ) );
INV_X4 \AES_ENC/us03/U482  ( .A(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n608 ));
NOR2_X2 \AES_ENC/us03/U480  ( .A1(\AES_ENC/us03/n1054 ), .A2(\AES_ENC/us03/n1053 ), .ZN(\AES_ENC/us03/n1055 ) );
OR2_X4 \AES_ENC/us03/U479  ( .A1(\AES_ENC/us03/n1094 ), .A2(\AES_ENC/us03/n1093 ), .ZN(\AES_ENC/us03/n571 ) );
AND2_X2 \AES_ENC/us03/U478  ( .A1(\AES_ENC/us03/n571 ), .A2(\AES_ENC/us03/n1095 ), .ZN(\AES_ENC/us03/n1101 ) );
NOR2_X2 \AES_ENC/us03/U477  ( .A1(\AES_ENC/us03/n1074 ), .A2(\AES_ENC/us03/n931 ), .ZN(\AES_ENC/us03/n796 ) );
NOR2_X2 \AES_ENC/us03/U474  ( .A1(\AES_ENC/us03/n796 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n797 ) );
NOR2_X2 \AES_ENC/us03/U473  ( .A1(\AES_ENC/us03/n932 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n933 ) );
NOR2_X2 \AES_ENC/us03/U472  ( .A1(\AES_ENC/us03/n929 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n935 ) );
NOR2_X2 \AES_ENC/us03/U471  ( .A1(\AES_ENC/us03/n931 ), .A2(\AES_ENC/us03/n930 ), .ZN(\AES_ENC/us03/n934 ) );
NOR3_X2 \AES_ENC/us03/U470  ( .A1(\AES_ENC/us03/n935 ), .A2(\AES_ENC/us03/n934 ), .A3(\AES_ENC/us03/n933 ), .ZN(\AES_ENC/us03/n936 ) );
NOR2_X2 \AES_ENC/us03/U469  ( .A1(\AES_ENC/us03/n626 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n1075 ) );
NOR2_X2 \AES_ENC/us03/U468  ( .A1(\AES_ENC/us03/n572 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n949 ) );
NOR2_X2 \AES_ENC/us03/U467  ( .A1(\AES_ENC/us03/n1049 ), .A2(\AES_ENC/us03/n620 ), .ZN(\AES_ENC/us03/n1051 ) );
NOR2_X2 \AES_ENC/us03/U466  ( .A1(\AES_ENC/us03/n1051 ), .A2(\AES_ENC/us03/n1050 ), .ZN(\AES_ENC/us03/n1052 ) );
NOR2_X2 \AES_ENC/us03/U465  ( .A1(\AES_ENC/us03/n1052 ), .A2(\AES_ENC/us03/n604 ), .ZN(\AES_ENC/us03/n1064 ) );
NOR2_X2 \AES_ENC/us03/U464  ( .A1(\AES_ENC/sa03 [1]), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n631 ) );
NOR2_X2 \AES_ENC/us03/U463  ( .A1(\AES_ENC/us03/n1025 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n980 ) );
NOR2_X2 \AES_ENC/us03/U462  ( .A1(\AES_ENC/us03/n1073 ), .A2(\AES_ENC/us03/n1094 ), .ZN(\AES_ENC/us03/n795 ) );
NOR2_X2 \AES_ENC/us03/U461  ( .A1(\AES_ENC/us03/n795 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n799 ) );
NOR2_X2 \AES_ENC/us03/U460  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n981 ) );
NOR2_X2 \AES_ENC/us03/U459  ( .A1(\AES_ENC/us03/n1102 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n643 ) );
NOR2_X2 \AES_ENC/us03/U458  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n623 ), .ZN(\AES_ENC/us03/n642 ) );
NOR2_X2 \AES_ENC/us03/U455  ( .A1(\AES_ENC/us03/n911 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n644 ) );
NOR4_X2 \AES_ENC/us03/U448  ( .A1(\AES_ENC/us03/n644 ), .A2(\AES_ENC/us03/n643 ), .A3(\AES_ENC/us03/n804 ), .A4(\AES_ENC/us03/n642 ), .ZN(\AES_ENC/us03/n645 ) );
NOR2_X2 \AES_ENC/us03/U447  ( .A1(\AES_ENC/us03/n1102 ), .A2(\AES_ENC/us03/n910 ), .ZN(\AES_ENC/us03/n932 ) );
NOR2_X2 \AES_ENC/us03/U442  ( .A1(\AES_ENC/us03/n1102 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n755 ) );
NOR2_X2 \AES_ENC/us03/U441  ( .A1(\AES_ENC/us03/n931 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n743 ) );
NOR2_X2 \AES_ENC/us03/U438  ( .A1(\AES_ENC/us03/n1072 ), .A2(\AES_ENC/us03/n1094 ), .ZN(\AES_ENC/us03/n930 ) );
NOR2_X2 \AES_ENC/us03/U435  ( .A1(\AES_ENC/us03/n1074 ), .A2(\AES_ENC/us03/n1025 ), .ZN(\AES_ENC/us03/n891 ) );
NOR2_X2 \AES_ENC/us03/U434  ( .A1(\AES_ENC/us03/n891 ), .A2(\AES_ENC/us03/n616 ), .ZN(\AES_ENC/us03/n894 ) );
NOR3_X2 \AES_ENC/us03/U433  ( .A1(\AES_ENC/us03/n625 ), .A2(\AES_ENC/sa03 [1]), .A3(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n683 ));
INV_X4 \AES_ENC/us03/U428  ( .A(\AES_ENC/us03/n931 ), .ZN(\AES_ENC/us03/n625 ) );
NOR2_X2 \AES_ENC/us03/U427  ( .A1(\AES_ENC/us03/n996 ), .A2(\AES_ENC/us03/n931 ), .ZN(\AES_ENC/us03/n704 ) );
NOR2_X2 \AES_ENC/us03/U421  ( .A1(\AES_ENC/us03/n931 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n685 ) );
NOR2_X2 \AES_ENC/us03/U420  ( .A1(\AES_ENC/us03/n1029 ), .A2(\AES_ENC/us03/n1025 ), .ZN(\AES_ENC/us03/n1079 ) );
NOR3_X2 \AES_ENC/us03/U419  ( .A1(\AES_ENC/us03/n601 ), .A2(\AES_ENC/us03/n1025 ), .A3(\AES_ENC/us03/n619 ), .ZN(\AES_ENC/us03/n945 ) );
NOR2_X2 \AES_ENC/us03/U418  ( .A1(\AES_ENC/us03/n627 ), .A2(\AES_ENC/us03/n618 ), .ZN(\AES_ENC/us03/n800 ) );
NOR3_X2 \AES_ENC/us03/U417  ( .A1(\AES_ENC/us03/n602 ), .A2(\AES_ENC/us03/n582 ), .A3(\AES_ENC/us03/n618 ), .ZN(\AES_ENC/us03/n798 ) );
NOR3_X2 \AES_ENC/us03/U416  ( .A1(\AES_ENC/us03/n617 ), .A2(\AES_ENC/us03/n572 ), .A3(\AES_ENC/us03/n590 ), .ZN(\AES_ENC/us03/n962 ) );
NOR3_X2 \AES_ENC/us03/U415  ( .A1(\AES_ENC/us03/n959 ), .A2(\AES_ENC/us03/n572 ), .A3(\AES_ENC/us03/n616 ), .ZN(\AES_ENC/us03/n768 ) );
NOR3_X2 \AES_ENC/us03/U414  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n572 ), .A3(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n694 ) );
NOR3_X2 \AES_ENC/us03/U413  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n572 ), .A3(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n895 ) );
NOR3_X2 \AES_ENC/us03/U410  ( .A1(\AES_ENC/us03/n1008 ), .A2(\AES_ENC/us03/n1007 ), .A3(\AES_ENC/us03/n1006 ), .ZN(\AES_ENC/us03/n1018 ) );
NOR4_X2 \AES_ENC/us03/U409  ( .A1(\AES_ENC/us03/n711 ), .A2(\AES_ENC/us03/n710 ), .A3(\AES_ENC/us03/n709 ), .A4(\AES_ENC/us03/n708 ), .ZN(\AES_ENC/us03/n712 ) );
NOR4_X2 \AES_ENC/us03/U406  ( .A1(\AES_ENC/us03/n806 ), .A2(\AES_ENC/us03/n805 ), .A3(\AES_ENC/us03/n804 ), .A4(\AES_ENC/us03/n803 ), .ZN(\AES_ENC/us03/n807 ) );
NOR3_X2 \AES_ENC/us03/U405  ( .A1(\AES_ENC/us03/n799 ), .A2(\AES_ENC/us03/n798 ), .A3(\AES_ENC/us03/n797 ), .ZN(\AES_ENC/us03/n808 ) );
NOR2_X2 \AES_ENC/us03/U404  ( .A1(\AES_ENC/us03/n669 ), .A2(\AES_ENC/us03/n668 ), .ZN(\AES_ENC/us03/n673 ) );
NOR4_X2 \AES_ENC/us03/U403  ( .A1(\AES_ENC/us03/n946 ), .A2(\AES_ENC/us03/n1046 ), .A3(\AES_ENC/us03/n671 ), .A4(\AES_ENC/us03/n670 ), .ZN(\AES_ENC/us03/n672 ) );
NOR3_X2 \AES_ENC/us03/U401  ( .A1(\AES_ENC/us03/n1101 ), .A2(\AES_ENC/us03/n1100 ), .A3(\AES_ENC/us03/n1099 ), .ZN(\AES_ENC/us03/n1109 ) );
NOR4_X2 \AES_ENC/us03/U400  ( .A1(\AES_ENC/us03/n843 ), .A2(\AES_ENC/us03/n842 ), .A3(\AES_ENC/us03/n841 ), .A4(\AES_ENC/us03/n840 ), .ZN(\AES_ENC/us03/n844 ) );
NOR4_X2 \AES_ENC/us03/U399  ( .A1(\AES_ENC/us03/n963 ), .A2(\AES_ENC/us03/n962 ), .A3(\AES_ENC/us03/n961 ), .A4(\AES_ENC/us03/n960 ), .ZN(\AES_ENC/us03/n964 ) );
NOR3_X2 \AES_ENC/us03/U398  ( .A1(\AES_ENC/us03/n743 ), .A2(\AES_ENC/us03/n742 ), .A3(\AES_ENC/us03/n741 ), .ZN(\AES_ENC/us03/n744 ) );
NOR2_X2 \AES_ENC/us03/U397  ( .A1(\AES_ENC/us03/n697 ), .A2(\AES_ENC/us03/n658 ), .ZN(\AES_ENC/us03/n659 ) );
NOR2_X2 \AES_ENC/us03/U396  ( .A1(\AES_ENC/us03/n1078 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n1033 ) );
NOR2_X2 \AES_ENC/us03/U393  ( .A1(\AES_ENC/us03/n1031 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n1032 ) );
NOR3_X2 \AES_ENC/us03/U390  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n1025 ), .A3(\AES_ENC/us03/n1074 ), .ZN(\AES_ENC/us03/n1035 ) );
NOR4_X2 \AES_ENC/us03/U389  ( .A1(\AES_ENC/us03/n1035 ), .A2(\AES_ENC/us03/n1034 ), .A3(\AES_ENC/us03/n1033 ), .A4(\AES_ENC/us03/n1032 ), .ZN(\AES_ENC/us03/n1036 ) );
NOR2_X2 \AES_ENC/us03/U388  ( .A1(\AES_ENC/us03/n610 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n885 ) );
NOR2_X2 \AES_ENC/us03/U387  ( .A1(\AES_ENC/us03/n625 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n882 ) );
NOR2_X2 \AES_ENC/us03/U386  ( .A1(\AES_ENC/us03/n1053 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n884 ) );
NOR4_X2 \AES_ENC/us03/U385  ( .A1(\AES_ENC/us03/n885 ), .A2(\AES_ENC/us03/n884 ), .A3(\AES_ENC/us03/n883 ), .A4(\AES_ENC/us03/n882 ), .ZN(\AES_ENC/us03/n886 ) );
NOR2_X2 \AES_ENC/us03/U384  ( .A1(\AES_ENC/us03/n825 ), .A2(\AES_ENC/us03/n593 ), .ZN(\AES_ENC/us03/n830 ) );
NOR2_X2 \AES_ENC/us03/U383  ( .A1(\AES_ENC/us03/n827 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n829 ) );
NOR2_X2 \AES_ENC/us03/U382  ( .A1(\AES_ENC/us03/n572 ), .A2(\AES_ENC/us03/n575 ), .ZN(\AES_ENC/us03/n828 ) );
NOR4_X2 \AES_ENC/us03/U374  ( .A1(\AES_ENC/us03/n831 ), .A2(\AES_ENC/us03/n830 ), .A3(\AES_ENC/us03/n829 ), .A4(\AES_ENC/us03/n828 ), .ZN(\AES_ENC/us03/n832 ) );
NOR2_X2 \AES_ENC/us03/U373  ( .A1(\AES_ENC/us03/n588 ), .A2(\AES_ENC/us03/n595 ), .ZN(\AES_ENC/us03/n1104 ) );
NOR2_X2 \AES_ENC/us03/U372  ( .A1(\AES_ENC/us03/n1102 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n1106 ) );
NOR2_X2 \AES_ENC/us03/U370  ( .A1(\AES_ENC/us03/n1103 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n1105 ) );
NOR4_X2 \AES_ENC/us03/U369  ( .A1(\AES_ENC/us03/n1107 ), .A2(\AES_ENC/us03/n1106 ), .A3(\AES_ENC/us03/n1105 ), .A4(\AES_ENC/us03/n1104 ), .ZN(\AES_ENC/us03/n1108 ) );
NOR3_X2 \AES_ENC/us03/U368  ( .A1(\AES_ENC/us03/n959 ), .A2(\AES_ENC/us03/n623 ), .A3(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n963 ) );
NOR2_X2 \AES_ENC/us03/U367  ( .A1(\AES_ENC/us03/n627 ), .A2(\AES_ENC/us03/n582 ), .ZN(\AES_ENC/us03/n1114 ) );
INV_X4 \AES_ENC/us03/U366  ( .A(\AES_ENC/us03/n1024 ), .ZN(\AES_ENC/us03/n588 ) );
NOR3_X2 \AES_ENC/us03/U365  ( .A1(\AES_ENC/us03/n910 ), .A2(\AES_ENC/us03/n1059 ), .A3(\AES_ENC/us03/n618 ), .ZN(\AES_ENC/us03/n1115 ) );
INV_X4 \AES_ENC/us03/U364  ( .A(\AES_ENC/us03/n1094 ), .ZN(\AES_ENC/us03/n585 ) );
NOR2_X2 \AES_ENC/us03/U363  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n931 ), .ZN(\AES_ENC/us03/n1100 ) );
INV_X4 \AES_ENC/us03/U354  ( .A(\AES_ENC/us03/n1093 ), .ZN(\AES_ENC/us03/n576 ) );
NOR2_X2 \AES_ENC/us03/U353  ( .A1(\AES_ENC/us03/n569 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n929 ) );
NOR2_X2 \AES_ENC/us03/U352  ( .A1(\AES_ENC/us03/n622 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n926 ) );
NOR2_X2 \AES_ENC/us03/U351  ( .A1(\AES_ENC/us03/n572 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n1095 ) );
NOR2_X2 \AES_ENC/us03/U350  ( .A1(\AES_ENC/us03/n616 ), .A2(\AES_ENC/us03/n582 ), .ZN(\AES_ENC/us03/n1010 ) );
NOR2_X2 \AES_ENC/us03/U349  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n1103 ) );
NOR2_X2 \AES_ENC/us03/U348  ( .A1(\AES_ENC/us03/n624 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n1059 ) );
NOR2_X2 \AES_ENC/us03/U347  ( .A1(\AES_ENC/sa03 [1]), .A2(\AES_ENC/us03/n1120 ), .ZN(\AES_ENC/us03/n1022 ) );
NOR2_X2 \AES_ENC/us03/U346  ( .A1(\AES_ENC/us03/n621 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n911 ) );
NOR2_X2 \AES_ENC/us03/U345  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/us03/n1025 ), .ZN(\AES_ENC/us03/n826 ) );
NOR2_X2 \AES_ENC/us03/U338  ( .A1(\AES_ENC/us03/n627 ), .A2(\AES_ENC/us03/n589 ), .ZN(\AES_ENC/us03/n1072 ) );
NOR2_X2 \AES_ENC/us03/U335  ( .A1(\AES_ENC/us03/n582 ), .A2(\AES_ENC/us03/n619 ), .ZN(\AES_ENC/us03/n956 ) );
NOR2_X2 \AES_ENC/us03/U329  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/us03/n626 ), .ZN(\AES_ENC/us03/n1121 ) );
NOR2_X2 \AES_ENC/us03/U328  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/us03/n626 ), .ZN(\AES_ENC/us03/n1058 ) );
NOR2_X2 \AES_ENC/us03/U327  ( .A1(\AES_ENC/us03/n578 ), .A2(\AES_ENC/us03/n618 ), .ZN(\AES_ENC/us03/n1073 ) );
NOR2_X2 \AES_ENC/us03/U325  ( .A1(\AES_ENC/sa03 [1]), .A2(\AES_ENC/us03/n1025 ), .ZN(\AES_ENC/us03/n1054 ) );
NOR2_X2 \AES_ENC/us03/U324  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/us03/n931 ), .ZN(\AES_ENC/us03/n1029 ) );
NOR2_X2 \AES_ENC/us03/U319  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n1056 ) );
NOR2_X2 \AES_ENC/us03/U318  ( .A1(\AES_ENC/us03/n586 ), .A2(\AES_ENC/us03/n627 ), .ZN(\AES_ENC/us03/n1050 ) );
NOR2_X2 \AES_ENC/us03/U317  ( .A1(\AES_ENC/us03/n1121 ), .A2(\AES_ENC/us03/n1025 ), .ZN(\AES_ENC/us03/n1120 ) );
NOR2_X2 \AES_ENC/us03/U316  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/us03/n572 ), .ZN(\AES_ENC/us03/n1074 ) );
NOR2_X2 \AES_ENC/us03/U315  ( .A1(\AES_ENC/us03/n1058 ), .A2(\AES_ENC/us03/n1054 ), .ZN(\AES_ENC/us03/n878 ) );
NOR2_X2 \AES_ENC/us03/U314  ( .A1(\AES_ENC/us03/n878 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n879 ) );
NOR2_X2 \AES_ENC/us03/U312  ( .A1(\AES_ENC/us03/n880 ), .A2(\AES_ENC/us03/n879 ), .ZN(\AES_ENC/us03/n887 ) );
NOR2_X2 \AES_ENC/us03/U311  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n600 ), .ZN(\AES_ENC/us03/n957 ) );
NOR2_X2 \AES_ENC/us03/U310  ( .A1(\AES_ENC/us03/n958 ), .A2(\AES_ENC/us03/n957 ), .ZN(\AES_ENC/us03/n965 ) );
NOR3_X2 \AES_ENC/us03/U309  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n1091 ), .A3(\AES_ENC/us03/n1022 ), .ZN(\AES_ENC/us03/n720 ) );
NOR3_X2 \AES_ENC/us03/U303  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n1054 ), .A3(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n719 ) );
NOR2_X2 \AES_ENC/us03/U302  ( .A1(\AES_ENC/us03/n720 ), .A2(\AES_ENC/us03/n719 ), .ZN(\AES_ENC/us03/n726 ) );
NOR2_X2 \AES_ENC/us03/U300  ( .A1(\AES_ENC/us03/n586 ), .A2(\AES_ENC/us03/n603 ), .ZN(\AES_ENC/us03/n865 ) );
NOR2_X2 \AES_ENC/us03/U299  ( .A1(\AES_ENC/us03/n1059 ), .A2(\AES_ENC/us03/n1058 ), .ZN(\AES_ENC/us03/n1060 ) );
NOR2_X2 \AES_ENC/us03/U298  ( .A1(\AES_ENC/us03/n1095 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n668 ) );
NOR2_X2 \AES_ENC/us03/U297  ( .A1(\AES_ENC/us03/n911 ), .A2(\AES_ENC/us03/n910 ), .ZN(\AES_ENC/us03/n912 ) );
NOR2_X2 \AES_ENC/us03/U296  ( .A1(\AES_ENC/us03/n912 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n916 ) );
NOR2_X2 \AES_ENC/us03/U295  ( .A1(\AES_ENC/us03/n826 ), .A2(\AES_ENC/us03/n573 ), .ZN(\AES_ENC/us03/n750 ) );
NOR2_X2 \AES_ENC/us03/U294  ( .A1(\AES_ENC/us03/n750 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n751 ) );
NOR2_X2 \AES_ENC/us03/U293  ( .A1(\AES_ENC/us03/n907 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n908 ) );
NOR2_X2 \AES_ENC/us03/U292  ( .A1(\AES_ENC/us03/n990 ), .A2(\AES_ENC/us03/n926 ), .ZN(\AES_ENC/us03/n780 ) );
NOR2_X2 \AES_ENC/us03/U291  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n597 ), .ZN(\AES_ENC/us03/n838 ) );
NOR2_X2 \AES_ENC/us03/U290  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n614 ), .ZN(\AES_ENC/us03/n837 ) );
NOR2_X2 \AES_ENC/us03/U284  ( .A1(\AES_ENC/us03/n838 ), .A2(\AES_ENC/us03/n837 ), .ZN(\AES_ENC/us03/n845 ) );
NOR2_X2 \AES_ENC/us03/U283  ( .A1(\AES_ENC/us03/n1022 ), .A2(\AES_ENC/us03/n1058 ), .ZN(\AES_ENC/us03/n740 ) );
NOR2_X2 \AES_ENC/us03/U282  ( .A1(\AES_ENC/us03/n740 ), .A2(\AES_ENC/us03/n619 ), .ZN(\AES_ENC/us03/n742 ) );
NOR2_X2 \AES_ENC/us03/U281  ( .A1(\AES_ENC/us03/n1098 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n1099 ) );
NOR2_X2 \AES_ENC/us03/U280  ( .A1(\AES_ENC/us03/n1120 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n993 ) );
NOR2_X2 \AES_ENC/us03/U279  ( .A1(\AES_ENC/us03/n993 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n994 ) );
NOR2_X2 \AES_ENC/us03/U273  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n622 ), .ZN(\AES_ENC/us03/n1026 ) );
NOR2_X2 \AES_ENC/us03/U272  ( .A1(\AES_ENC/us03/n573 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n1027 ) );
NOR2_X2 \AES_ENC/us03/U271  ( .A1(\AES_ENC/us03/n1027 ), .A2(\AES_ENC/us03/n1026 ), .ZN(\AES_ENC/us03/n1028 ) );
NOR2_X2 \AES_ENC/us03/U270  ( .A1(\AES_ENC/us03/n1029 ), .A2(\AES_ENC/us03/n1028 ), .ZN(\AES_ENC/us03/n1034 ) );
NOR4_X2 \AES_ENC/us03/U269  ( .A1(\AES_ENC/us03/n757 ), .A2(\AES_ENC/us03/n756 ), .A3(\AES_ENC/us03/n755 ), .A4(\AES_ENC/us03/n754 ), .ZN(\AES_ENC/us03/n758 ) );
NOR2_X2 \AES_ENC/us03/U268  ( .A1(\AES_ENC/us03/n752 ), .A2(\AES_ENC/us03/n751 ), .ZN(\AES_ENC/us03/n759 ) );
NOR2_X2 \AES_ENC/us03/U267  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n1071 ), .ZN(\AES_ENC/us03/n669 ) );
NOR2_X2 \AES_ENC/us03/U263  ( .A1(\AES_ENC/us03/n1056 ), .A2(\AES_ENC/us03/n990 ), .ZN(\AES_ENC/us03/n991 ) );
NOR2_X2 \AES_ENC/us03/U262  ( .A1(\AES_ENC/us03/n991 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n995 ) );
NOR2_X2 \AES_ENC/us03/U258  ( .A1(\AES_ENC/us03/n589 ), .A2(\AES_ENC/us03/n602 ), .ZN(\AES_ENC/us03/n1008 ) );
NOR2_X2 \AES_ENC/us03/U255  ( .A1(\AES_ENC/us03/n839 ), .A2(\AES_ENC/us03/n595 ), .ZN(\AES_ENC/us03/n693 ) );
NOR2_X2 \AES_ENC/us03/U254  ( .A1(\AES_ENC/us03/n588 ), .A2(\AES_ENC/us03/n906 ), .ZN(\AES_ENC/us03/n741 ) );
NOR2_X2 \AES_ENC/us03/U253  ( .A1(\AES_ENC/us03/n1054 ), .A2(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n763 ) );
NOR2_X2 \AES_ENC/us03/U252  ( .A1(\AES_ENC/us03/n763 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n769 ) );
NOR2_X2 \AES_ENC/us03/U251  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n592 ), .ZN(\AES_ENC/us03/n1007 ) );
NOR2_X2 \AES_ENC/us03/U250  ( .A1(\AES_ENC/us03/n616 ), .A2(\AES_ENC/us03/n594 ), .ZN(\AES_ENC/us03/n1123 ) );
NOR2_X2 \AES_ENC/us03/U243  ( .A1(\AES_ENC/us03/n616 ), .A2(\AES_ENC/us03/n602 ), .ZN(\AES_ENC/us03/n710 ) );
INV_X4 \AES_ENC/us03/U242  ( .A(\AES_ENC/us03/n1029 ), .ZN(\AES_ENC/us03/n595 ) );
NOR2_X2 \AES_ENC/us03/U241  ( .A1(\AES_ENC/us03/n619 ), .A2(\AES_ENC/us03/n609 ), .ZN(\AES_ENC/us03/n883 ) );
NOR2_X2 \AES_ENC/us03/U240  ( .A1(\AES_ENC/us03/n605 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n1125 ) );
NOR2_X2 \AES_ENC/us03/U239  ( .A1(\AES_ENC/us03/n990 ), .A2(\AES_ENC/us03/n929 ), .ZN(\AES_ENC/us03/n892 ) );
NOR2_X2 \AES_ENC/us03/U238  ( .A1(\AES_ENC/us03/n892 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n893 ) );
NOR2_X2 \AES_ENC/us03/U237  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n614 ), .ZN(\AES_ENC/us03/n950 ) );
NOR2_X2 \AES_ENC/us03/U236  ( .A1(\AES_ENC/us03/n1079 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n1082 ) );
NOR2_X2 \AES_ENC/us03/U235  ( .A1(\AES_ENC/us03/n910 ), .A2(\AES_ENC/us03/n1056 ), .ZN(\AES_ENC/us03/n941 ) );
NOR2_X2 \AES_ENC/us03/U234  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n1077 ), .ZN(\AES_ENC/us03/n841 ) );
NOR2_X2 \AES_ENC/us03/U229  ( .A1(\AES_ENC/us03/n625 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n630 ) );
NOR2_X2 \AES_ENC/us03/U228  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n614 ), .ZN(\AES_ENC/us03/n806 ) );
NOR2_X2 \AES_ENC/us03/U227  ( .A1(\AES_ENC/us03/n625 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n948 ) );
NOR2_X2 \AES_ENC/us03/U226  ( .A1(\AES_ENC/us03/n588 ), .A2(\AES_ENC/us03/n601 ), .ZN(\AES_ENC/us03/n997 ) );
NOR2_X2 \AES_ENC/us03/U225  ( .A1(\AES_ENC/us03/n1121 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n1122 ) );
NOR2_X2 \AES_ENC/us03/U223  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n1023 ), .ZN(\AES_ENC/us03/n756 ) );
NOR2_X2 \AES_ENC/us03/U222  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n614 ), .ZN(\AES_ENC/us03/n870 ) );
NOR2_X2 \AES_ENC/us03/U221  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n569 ), .ZN(\AES_ENC/us03/n947 ) );
NOR2_X2 \AES_ENC/us03/U217  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n1077 ), .ZN(\AES_ENC/us03/n1084 ) );
NOR2_X2 \AES_ENC/us03/U213  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n855 ), .ZN(\AES_ENC/us03/n709 ) );
NOR2_X2 \AES_ENC/us03/U212  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n601 ), .ZN(\AES_ENC/us03/n868 ) );
NOR2_X2 \AES_ENC/us03/U211  ( .A1(\AES_ENC/us03/n1120 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n1124 ) );
NOR2_X2 \AES_ENC/us03/U210  ( .A1(\AES_ENC/us03/n1120 ), .A2(\AES_ENC/us03/n839 ), .ZN(\AES_ENC/us03/n842 ) );
NOR2_X2 \AES_ENC/us03/U209  ( .A1(\AES_ENC/us03/n1120 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n696 ) );
NOR2_X2 \AES_ENC/us03/U208  ( .A1(\AES_ENC/us03/n1074 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n1076 ) );
NOR2_X2 \AES_ENC/us03/U207  ( .A1(\AES_ENC/us03/n1074 ), .A2(\AES_ENC/us03/n622 ), .ZN(\AES_ENC/us03/n781 ) );
NOR3_X2 \AES_ENC/us03/U201  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n1056 ), .A3(\AES_ENC/us03/n990 ), .ZN(\AES_ENC/us03/n979 ) );
NOR3_X2 \AES_ENC/us03/U200  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n1058 ), .A3(\AES_ENC/us03/n1059 ), .ZN(\AES_ENC/us03/n854 ) );
NOR2_X2 \AES_ENC/us03/U199  ( .A1(\AES_ENC/us03/n996 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n869 ) );
NOR2_X2 \AES_ENC/us03/U198  ( .A1(\AES_ENC/us03/n1056 ), .A2(\AES_ENC/us03/n1074 ), .ZN(\AES_ENC/us03/n1057 ) );
NOR3_X2 \AES_ENC/us03/U197  ( .A1(\AES_ENC/us03/n589 ), .A2(\AES_ENC/us03/n1120 ), .A3(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n978 ) );
NOR2_X2 \AES_ENC/us03/U196  ( .A1(\AES_ENC/us03/n996 ), .A2(\AES_ENC/us03/n911 ), .ZN(\AES_ENC/us03/n1116 ) );
NOR2_X2 \AES_ENC/us03/U195  ( .A1(\AES_ENC/us03/n1074 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n754 ) );
NOR2_X2 \AES_ENC/us03/U194  ( .A1(\AES_ENC/us03/n926 ), .A2(\AES_ENC/us03/n1103 ), .ZN(\AES_ENC/us03/n977 ) );
NOR2_X2 \AES_ENC/us03/U187  ( .A1(\AES_ENC/us03/n839 ), .A2(\AES_ENC/us03/n824 ), .ZN(\AES_ENC/us03/n1092 ) );
NOR2_X2 \AES_ENC/us03/U186  ( .A1(\AES_ENC/us03/n573 ), .A2(\AES_ENC/us03/n1074 ), .ZN(\AES_ENC/us03/n684 ) );
NOR2_X2 \AES_ENC/us03/U185  ( .A1(\AES_ENC/us03/n826 ), .A2(\AES_ENC/us03/n1059 ), .ZN(\AES_ENC/us03/n907 ) );
NOR3_X2 \AES_ENC/us03/U184  ( .A1(\AES_ENC/us03/n578 ), .A2(\AES_ENC/us03/n1115 ), .A3(\AES_ENC/us03/n598 ), .ZN(\AES_ENC/us03/n831 ) );
NOR3_X2 \AES_ENC/us03/U183  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n1056 ), .A3(\AES_ENC/us03/n990 ), .ZN(\AES_ENC/us03/n896 ) );
NOR3_X2 \AES_ENC/us03/U182  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n573 ), .A3(\AES_ENC/us03/n1013 ), .ZN(\AES_ENC/us03/n670 ) );
NOR3_X2 \AES_ENC/us03/U181  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n1091 ), .A3(\AES_ENC/us03/n1022 ), .ZN(\AES_ENC/us03/n843 ) );
NOR2_X2 \AES_ENC/us03/U180  ( .A1(\AES_ENC/us03/n1029 ), .A2(\AES_ENC/us03/n1095 ), .ZN(\AES_ENC/us03/n735 ) );
NOR4_X2 \AES_ENC/us03/U174  ( .A1(\AES_ENC/us03/n983 ), .A2(\AES_ENC/us03/n982 ), .A3(\AES_ENC/us03/n981 ), .A4(\AES_ENC/us03/n980 ), .ZN(\AES_ENC/us03/n984 ) );
NOR2_X2 \AES_ENC/us03/U173  ( .A1(\AES_ENC/us03/n979 ), .A2(\AES_ENC/us03/n978 ), .ZN(\AES_ENC/us03/n985 ) );
NAND3_X2 \AES_ENC/us03/U172  ( .A1(\AES_ENC/us03/n569 ), .A2(\AES_ENC/us03/n595 ), .A3(\AES_ENC/us03/n681 ), .ZN(\AES_ENC/us03/n691 ) );
NOR2_X2 \AES_ENC/us03/U171  ( .A1(\AES_ENC/us03/n683 ), .A2(\AES_ENC/us03/n682 ), .ZN(\AES_ENC/us03/n690 ) );
NOR3_X2 \AES_ENC/us03/U170  ( .A1(\AES_ENC/us03/n695 ), .A2(\AES_ENC/us03/n694 ), .A3(\AES_ENC/us03/n693 ), .ZN(\AES_ENC/us03/n700 ) );
NOR4_X2 \AES_ENC/us03/U169  ( .A1(\AES_ENC/us03/n983 ), .A2(\AES_ENC/us03/n698 ), .A3(\AES_ENC/us03/n697 ), .A4(\AES_ENC/us03/n696 ), .ZN(\AES_ENC/us03/n699 ) );
NOR2_X2 \AES_ENC/us03/U168  ( .A1(\AES_ENC/us03/n1100 ), .A2(\AES_ENC/us03/n854 ), .ZN(\AES_ENC/us03/n860 ) );
NOR4_X2 \AES_ENC/us03/U162  ( .A1(\AES_ENC/us03/n1125 ), .A2(\AES_ENC/us03/n1124 ), .A3(\AES_ENC/us03/n1123 ), .A4(\AES_ENC/us03/n1122 ), .ZN(\AES_ENC/us03/n1126 ) );
NOR4_X2 \AES_ENC/us03/U161  ( .A1(\AES_ENC/us03/n1084 ), .A2(\AES_ENC/us03/n1083 ), .A3(\AES_ENC/us03/n1082 ), .A4(\AES_ENC/us03/n1081 ), .ZN(\AES_ENC/us03/n1085 ) );
NOR2_X2 \AES_ENC/us03/U160  ( .A1(\AES_ENC/us03/n1076 ), .A2(\AES_ENC/us03/n1075 ), .ZN(\AES_ENC/us03/n1086 ) );
NOR4_X2 \AES_ENC/us03/U159  ( .A1(\AES_ENC/us03/n896 ), .A2(\AES_ENC/us03/n895 ), .A3(\AES_ENC/us03/n894 ), .A4(\AES_ENC/us03/n893 ), .ZN(\AES_ENC/us03/n897 ) );
NOR2_X2 \AES_ENC/us03/U158  ( .A1(\AES_ENC/us03/n866 ), .A2(\AES_ENC/us03/n865 ), .ZN(\AES_ENC/us03/n872 ) );
NOR4_X2 \AES_ENC/us03/U157  ( .A1(\AES_ENC/us03/n870 ), .A2(\AES_ENC/us03/n869 ), .A3(\AES_ENC/us03/n868 ), .A4(\AES_ENC/us03/n867 ), .ZN(\AES_ENC/us03/n871 ) );
NOR2_X2 \AES_ENC/us03/U156  ( .A1(\AES_ENC/us03/n946 ), .A2(\AES_ENC/us03/n945 ), .ZN(\AES_ENC/us03/n952 ) );
NOR4_X2 \AES_ENC/us03/U155  ( .A1(\AES_ENC/us03/n950 ), .A2(\AES_ENC/us03/n949 ), .A3(\AES_ENC/us03/n948 ), .A4(\AES_ENC/us03/n947 ), .ZN(\AES_ENC/us03/n951 ) );
NOR3_X2 \AES_ENC/us03/U154  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n1054 ), .A3(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n961 ) );
NOR3_X2 \AES_ENC/us03/U153  ( .A1(\AES_ENC/us03/n622 ), .A2(\AES_ENC/us03/n1074 ), .A3(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n671 ) );
NOR2_X2 \AES_ENC/us03/U152  ( .A1(\AES_ENC/us03/n1057 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n1062 ) );
NOR2_X2 \AES_ENC/us03/U143  ( .A1(\AES_ENC/us03/n1055 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n1063 ) );
NOR2_X2 \AES_ENC/us03/U142  ( .A1(\AES_ENC/us03/n1060 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n1061 ) );
NOR4_X2 \AES_ENC/us03/U141  ( .A1(\AES_ENC/us03/n1064 ), .A2(\AES_ENC/us03/n1063 ), .A3(\AES_ENC/us03/n1062 ), .A4(\AES_ENC/us03/n1061 ), .ZN(\AES_ENC/us03/n1065 ) );
NOR2_X2 \AES_ENC/us03/U140  ( .A1(\AES_ENC/us03/n735 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n687 ) );
NOR2_X2 \AES_ENC/us03/U132  ( .A1(\AES_ENC/us03/n684 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n688 ) );
NOR2_X2 \AES_ENC/us03/U131  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n612 ), .ZN(\AES_ENC/us03/n686 ) );
NOR4_X2 \AES_ENC/us03/U130  ( .A1(\AES_ENC/us03/n688 ), .A2(\AES_ENC/us03/n687 ), .A3(\AES_ENC/us03/n686 ), .A4(\AES_ENC/us03/n685 ), .ZN(\AES_ENC/us03/n689 ) );
NOR2_X2 \AES_ENC/us03/U129  ( .A1(\AES_ENC/us03/n619 ), .A2(\AES_ENC/us03/n594 ), .ZN(\AES_ENC/us03/n771 ) );
NOR2_X2 \AES_ENC/us03/U128  ( .A1(\AES_ENC/us03/n1103 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n772 ) );
NOR2_X2 \AES_ENC/us03/U127  ( .A1(\AES_ENC/us03/n617 ), .A2(\AES_ENC/us03/n611 ), .ZN(\AES_ENC/us03/n773 ) );
NOR4_X2 \AES_ENC/us03/U126  ( .A1(\AES_ENC/us03/n773 ), .A2(\AES_ENC/us03/n772 ), .A3(\AES_ENC/us03/n771 ), .A4(\AES_ENC/us03/n770 ), .ZN(\AES_ENC/us03/n774 ) );
NOR2_X2 \AES_ENC/us03/U121  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n607 ), .ZN(\AES_ENC/us03/n858 ) );
NOR2_X2 \AES_ENC/us03/U120  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n855 ), .ZN(\AES_ENC/us03/n857 ) );
NOR2_X2 \AES_ENC/us03/U119  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n599 ), .ZN(\AES_ENC/us03/n856 ) );
NOR4_X2 \AES_ENC/us03/U118  ( .A1(\AES_ENC/us03/n858 ), .A2(\AES_ENC/us03/n857 ), .A3(\AES_ENC/us03/n856 ), .A4(\AES_ENC/us03/n958 ), .ZN(\AES_ENC/us03/n859 ) );
NOR3_X2 \AES_ENC/us03/U117  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n1120 ), .A3(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n918 ) );
NOR3_X2 \AES_ENC/us03/U116  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n573 ), .A3(\AES_ENC/us03/n1013 ), .ZN(\AES_ENC/us03/n917 ) );
NOR2_X2 \AES_ENC/us03/U115  ( .A1(\AES_ENC/us03/n914 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n915 ) );
NOR4_X2 \AES_ENC/us03/U106  ( .A1(\AES_ENC/us03/n918 ), .A2(\AES_ENC/us03/n917 ), .A3(\AES_ENC/us03/n916 ), .A4(\AES_ENC/us03/n915 ), .ZN(\AES_ENC/us03/n919 ) );
NOR2_X2 \AES_ENC/us03/U105  ( .A1(\AES_ENC/us03/n780 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n784 ) );
NOR2_X2 \AES_ENC/us03/U104  ( .A1(\AES_ENC/us03/n1117 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n782 ) );
NOR2_X2 \AES_ENC/us03/U103  ( .A1(\AES_ENC/us03/n781 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n783 ) );
NOR4_X2 \AES_ENC/us03/U102  ( .A1(\AES_ENC/us03/n880 ), .A2(\AES_ENC/us03/n784 ), .A3(\AES_ENC/us03/n783 ), .A4(\AES_ENC/us03/n782 ), .ZN(\AES_ENC/us03/n785 ) );
NOR2_X2 \AES_ENC/us03/U101  ( .A1(\AES_ENC/us03/n596 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n814 ) );
NOR2_X2 \AES_ENC/us03/U100  ( .A1(\AES_ENC/us03/n907 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n813 ) );
NOR3_X2 \AES_ENC/us03/U95  ( .A1(\AES_ENC/us03/n588 ), .A2(\AES_ENC/us03/n1058 ), .A3(\AES_ENC/us03/n1059 ), .ZN(\AES_ENC/us03/n815 ) );
NOR4_X2 \AES_ENC/us03/U94  ( .A1(\AES_ENC/us03/n815 ), .A2(\AES_ENC/us03/n814 ), .A3(\AES_ENC/us03/n813 ), .A4(\AES_ENC/us03/n812 ), .ZN(\AES_ENC/us03/n816 ) );
NOR2_X2 \AES_ENC/us03/U93  ( .A1(\AES_ENC/us03/n576 ), .A2(\AES_ENC/us03/n569 ), .ZN(\AES_ENC/us03/n721 ) );
NOR2_X2 \AES_ENC/us03/U92  ( .A1(\AES_ENC/us03/n1031 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n723 ) );
NOR2_X2 \AES_ENC/us03/U91  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n1096 ), .ZN(\AES_ENC/us03/n722 ) );
NOR4_X2 \AES_ENC/us03/U90  ( .A1(\AES_ENC/us03/n724 ), .A2(\AES_ENC/us03/n723 ), .A3(\AES_ENC/us03/n722 ), .A4(\AES_ENC/us03/n721 ), .ZN(\AES_ENC/us03/n725 ) );
NOR2_X2 \AES_ENC/us03/U89  ( .A1(\AES_ENC/us03/n911 ), .A2(\AES_ENC/us03/n990 ), .ZN(\AES_ENC/us03/n1009 ) );
NOR2_X2 \AES_ENC/us03/U88  ( .A1(\AES_ENC/us03/n1013 ), .A2(\AES_ENC/us03/n573 ), .ZN(\AES_ENC/us03/n1014 ) );
NOR2_X2 \AES_ENC/us03/U87  ( .A1(\AES_ENC/us03/n1014 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n1015 ) );
NOR4_X2 \AES_ENC/us03/U86  ( .A1(\AES_ENC/us03/n1016 ), .A2(\AES_ENC/us03/n1015 ), .A3(\AES_ENC/us03/n1119 ), .A4(\AES_ENC/us03/n1046 ), .ZN(\AES_ENC/us03/n1017 ) );
NOR2_X2 \AES_ENC/us03/U81  ( .A1(\AES_ENC/us03/n996 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n998 ) );
NOR2_X2 \AES_ENC/us03/U80  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n592 ), .ZN(\AES_ENC/us03/n1000 ) );
NOR2_X2 \AES_ENC/us03/U79  ( .A1(\AES_ENC/us03/n619 ), .A2(\AES_ENC/us03/n1096 ), .ZN(\AES_ENC/us03/n999 ) );
NOR4_X2 \AES_ENC/us03/U78  ( .A1(\AES_ENC/us03/n1000 ), .A2(\AES_ENC/us03/n999 ), .A3(\AES_ENC/us03/n998 ), .A4(\AES_ENC/us03/n997 ), .ZN(\AES_ENC/us03/n1001 ) );
NOR2_X2 \AES_ENC/us03/U74  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n1096 ), .ZN(\AES_ENC/us03/n697 ) );
NOR2_X2 \AES_ENC/us03/U73  ( .A1(\AES_ENC/us03/n622 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n958 ) );
NOR2_X2 \AES_ENC/us03/U72  ( .A1(\AES_ENC/us03/n911 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n983 ) );
NOR2_X2 \AES_ENC/us03/U71  ( .A1(\AES_ENC/us03/n1054 ), .A2(\AES_ENC/us03/n1103 ), .ZN(\AES_ENC/us03/n1031 ) );
INV_X4 \AES_ENC/us03/U65  ( .A(\AES_ENC/us03/n1050 ), .ZN(\AES_ENC/us03/n583 ) );
INV_X4 \AES_ENC/us03/U64  ( .A(\AES_ENC/us03/n1072 ), .ZN(\AES_ENC/us03/n587 ) );
INV_X4 \AES_ENC/us03/U63  ( .A(\AES_ENC/us03/n1073 ), .ZN(\AES_ENC/us03/n577 ) );
NOR2_X2 \AES_ENC/us03/U62  ( .A1(\AES_ENC/us03/n595 ), .A2(\AES_ENC/us03/n585 ), .ZN(\AES_ENC/us03/n880 ) );
NOR3_X2 \AES_ENC/us03/U61  ( .A1(\AES_ENC/us03/n826 ), .A2(\AES_ENC/us03/n1121 ), .A3(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n946 ) );
INV_X4 \AES_ENC/us03/U59  ( .A(\AES_ENC/us03/n1010 ), .ZN(\AES_ENC/us03/n580 ) );
NOR3_X2 \AES_ENC/us03/U58  ( .A1(\AES_ENC/us03/n573 ), .A2(\AES_ENC/us03/n1029 ), .A3(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n1119 ) );
INV_X4 \AES_ENC/us03/U57  ( .A(\AES_ENC/us03/n956 ), .ZN(\AES_ENC/us03/n581 ) );
NOR2_X2 \AES_ENC/us03/U50  ( .A1(\AES_ENC/us03/n625 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n1013 ) );
NOR2_X2 \AES_ENC/us03/U49  ( .A1(\AES_ENC/us03/n622 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n910 ) );
NOR2_X2 \AES_ENC/us03/U48  ( .A1(\AES_ENC/us03/n569 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n1091 ) );
NOR2_X2 \AES_ENC/us03/U47  ( .A1(\AES_ENC/us03/n624 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n990 ) );
NOR2_X2 \AES_ENC/us03/U46  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/us03/n1121 ), .ZN(\AES_ENC/us03/n996 ) );
NOR2_X2 \AES_ENC/us03/U45  ( .A1(\AES_ENC/us03/n617 ), .A2(\AES_ENC/us03/n612 ), .ZN(\AES_ENC/us03/n628 ) );
NOR2_X2 \AES_ENC/us03/U44  ( .A1(\AES_ENC/us03/n591 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n866 ) );
NOR2_X2 \AES_ENC/us03/U43  ( .A1(\AES_ENC/us03/n615 ), .A2(\AES_ENC/us03/n617 ), .ZN(\AES_ENC/us03/n1006 ) );
NOR2_X2 \AES_ENC/us03/U42  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n1117 ), .ZN(\AES_ENC/us03/n1118 ) );
NOR2_X2 \AES_ENC/us03/U41  ( .A1(\AES_ENC/us03/n1119 ), .A2(\AES_ENC/us03/n1118 ), .ZN(\AES_ENC/us03/n1127 ) );
NOR2_X2 \AES_ENC/us03/U36  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n606 ), .ZN(\AES_ENC/us03/n629 ) );
NOR2_X2 \AES_ENC/us03/U35  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n906 ), .ZN(\AES_ENC/us03/n909 ) );
NOR2_X2 \AES_ENC/us03/U34  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n609 ), .ZN(\AES_ENC/us03/n658 ) );
NOR2_X2 \AES_ENC/us03/U33  ( .A1(\AES_ENC/us03/n1116 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n695 ) );
NOR2_X2 \AES_ENC/us03/U32  ( .A1(\AES_ENC/us03/n1078 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n1083 ) );
NOR2_X2 \AES_ENC/us03/U31  ( .A1(\AES_ENC/us03/n941 ), .A2(\AES_ENC/us03/n580 ), .ZN(\AES_ENC/us03/n724 ) );
NOR2_X2 \AES_ENC/us03/U30  ( .A1(\AES_ENC/us03/n610 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n1107 ) );
NOR2_X2 \AES_ENC/us03/U29  ( .A1(\AES_ENC/us03/n591 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n840 ) );
NOR2_X2 \AES_ENC/us03/U24  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n605 ), .ZN(\AES_ENC/us03/n633 ) );
NOR2_X2 \AES_ENC/us03/U23  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n1080 ), .ZN(\AES_ENC/us03/n1081 ) );
NOR2_X2 \AES_ENC/us03/U21  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n1045 ), .ZN(\AES_ENC/us03/n812 ) );
NOR2_X2 \AES_ENC/us03/U20  ( .A1(\AES_ENC/us03/n1009 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n960 ) );
NOR2_X2 \AES_ENC/us03/U19  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n613 ), .ZN(\AES_ENC/us03/n982 ) );
NOR2_X2 \AES_ENC/us03/U18  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n606 ), .ZN(\AES_ENC/us03/n757 ) );
NOR2_X2 \AES_ENC/us03/U17  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n602 ), .ZN(\AES_ENC/us03/n698 ) );
NOR2_X2 \AES_ENC/us03/U16  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n621 ), .ZN(\AES_ENC/us03/n708 ) );
NOR2_X2 \AES_ENC/us03/U15  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n595 ), .ZN(\AES_ENC/us03/n770 ) );
NOR2_X2 \AES_ENC/us03/U10  ( .A1(\AES_ENC/us03/n621 ), .A2(\AES_ENC/us03/n577 ), .ZN(\AES_ENC/us03/n803 ) );
NOR2_X2 \AES_ENC/us03/U9  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n881 ), .ZN(\AES_ENC/us03/n711 ) );
NOR2_X2 \AES_ENC/us03/U8  ( .A1(\AES_ENC/us03/n581 ), .A2(\AES_ENC/us03/n595 ), .ZN(\AES_ENC/us03/n867 ) );
NOR2_X2 \AES_ENC/us03/U7  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n611 ), .ZN(\AES_ENC/us03/n804 ) );
NOR2_X2 \AES_ENC/us03/U6  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n622 ), .ZN(\AES_ENC/us03/n1046 ) );
OR2_X4 \AES_ENC/us03/U5  ( .A1(\AES_ENC/us03/n626 ), .A2(\AES_ENC/sa03 [1]),.ZN(\AES_ENC/us03/n570 ) );
OR2_X4 \AES_ENC/us03/U4  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/sa03 [4]),.ZN(\AES_ENC/us03/n569 ) );
NAND2_X2 \AES_ENC/us03/U514  ( .A1(\AES_ENC/us03/n1121 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n1030 ) );
AND2_X2 \AES_ENC/us03/U513  ( .A1(\AES_ENC/us03/n609 ), .A2(\AES_ENC/us03/n1030 ), .ZN(\AES_ENC/us03/n1049 ) );
NAND2_X2 \AES_ENC/us03/U511  ( .A1(\AES_ENC/us03/n1049 ), .A2(\AES_ENC/us03/n794 ), .ZN(\AES_ENC/us03/n637 ) );
AND2_X2 \AES_ENC/us03/U493  ( .A1(\AES_ENC/us03/n779 ), .A2(\AES_ENC/us03/n996 ), .ZN(\AES_ENC/us03/n632 ) );
NAND4_X2 \AES_ENC/us03/U485  ( .A1(\AES_ENC/us03/n637 ), .A2(\AES_ENC/us03/n636 ), .A3(\AES_ENC/us03/n635 ), .A4(\AES_ENC/us03/n634 ), .ZN(\AES_ENC/us03/n638 ) );
NAND2_X2 \AES_ENC/us03/U484  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n638 ), .ZN(\AES_ENC/us03/n679 ) );
NAND2_X2 \AES_ENC/us03/U481  ( .A1(\AES_ENC/us03/n1094 ), .A2(\AES_ENC/us03/n603 ), .ZN(\AES_ENC/us03/n648 ) );
NAND2_X2 \AES_ENC/us03/U476  ( .A1(\AES_ENC/us03/n613 ), .A2(\AES_ENC/us03/n602 ), .ZN(\AES_ENC/us03/n762 ) );
NAND2_X2 \AES_ENC/us03/U475  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n762 ), .ZN(\AES_ENC/us03/n647 ) );
NAND4_X2 \AES_ENC/us03/U457  ( .A1(\AES_ENC/us03/n648 ), .A2(\AES_ENC/us03/n647 ), .A3(\AES_ENC/us03/n646 ), .A4(\AES_ENC/us03/n645 ), .ZN(\AES_ENC/us03/n649 ) );
NAND2_X2 \AES_ENC/us03/U456  ( .A1(\AES_ENC/sa03 [0]), .A2(\AES_ENC/us03/n649 ), .ZN(\AES_ENC/us03/n665 ) );
NAND2_X2 \AES_ENC/us03/U454  ( .A1(\AES_ENC/us03/n608 ), .A2(\AES_ENC/us03/n625 ), .ZN(\AES_ENC/us03/n855 ) );
NAND2_X2 \AES_ENC/us03/U453  ( .A1(\AES_ENC/us03/n599 ), .A2(\AES_ENC/us03/n855 ), .ZN(\AES_ENC/us03/n821 ) );
NAND2_X2 \AES_ENC/us03/U452  ( .A1(\AES_ENC/us03/n1093 ), .A2(\AES_ENC/us03/n821 ), .ZN(\AES_ENC/us03/n662 ) );
NAND2_X2 \AES_ENC/us03/U451  ( .A1(\AES_ENC/us03/n621 ), .A2(\AES_ENC/us03/n601 ), .ZN(\AES_ENC/us03/n650 ) );
NAND2_X2 \AES_ENC/us03/U450  ( .A1(\AES_ENC/us03/n956 ), .A2(\AES_ENC/us03/n650 ), .ZN(\AES_ENC/us03/n661 ) );
NAND2_X2 \AES_ENC/us03/U449  ( .A1(\AES_ENC/us03/n627 ), .A2(\AES_ENC/us03/n582 ), .ZN(\AES_ENC/us03/n839 ) );
OR2_X2 \AES_ENC/us03/U446  ( .A1(\AES_ENC/us03/n839 ), .A2(\AES_ENC/us03/n932 ), .ZN(\AES_ENC/us03/n656 ) );
NAND2_X2 \AES_ENC/us03/U445  ( .A1(\AES_ENC/us03/n623 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n1096 ) );
NAND2_X2 \AES_ENC/us03/U444  ( .A1(\AES_ENC/us03/n1030 ), .A2(\AES_ENC/us03/n1096 ), .ZN(\AES_ENC/us03/n651 ) );
NAND2_X2 \AES_ENC/us03/U443  ( .A1(\AES_ENC/us03/n1114 ), .A2(\AES_ENC/us03/n651 ), .ZN(\AES_ENC/us03/n655 ) );
OR3_X2 \AES_ENC/us03/U440  ( .A1(\AES_ENC/us03/n1079 ), .A2(\AES_ENC/sa03 [7]), .A3(\AES_ENC/us03/n627 ), .ZN(\AES_ENC/us03/n654 ));
NAND2_X2 \AES_ENC/us03/U439  ( .A1(\AES_ENC/us03/n605 ), .A2(\AES_ENC/us03/n613 ), .ZN(\AES_ENC/us03/n652 ) );
NAND4_X2 \AES_ENC/us03/U437  ( .A1(\AES_ENC/us03/n656 ), .A2(\AES_ENC/us03/n655 ), .A3(\AES_ENC/us03/n654 ), .A4(\AES_ENC/us03/n653 ), .ZN(\AES_ENC/us03/n657 ) );
NAND2_X2 \AES_ENC/us03/U436  ( .A1(\AES_ENC/sa03 [2]), .A2(\AES_ENC/us03/n657 ), .ZN(\AES_ENC/us03/n660 ) );
NAND4_X2 \AES_ENC/us03/U432  ( .A1(\AES_ENC/us03/n662 ), .A2(\AES_ENC/us03/n661 ), .A3(\AES_ENC/us03/n660 ), .A4(\AES_ENC/us03/n659 ), .ZN(\AES_ENC/us03/n663 ) );
NAND2_X2 \AES_ENC/us03/U431  ( .A1(\AES_ENC/us03/n663 ), .A2(\AES_ENC/us03/n574 ), .ZN(\AES_ENC/us03/n664 ) );
NAND2_X2 \AES_ENC/us03/U430  ( .A1(\AES_ENC/us03/n665 ), .A2(\AES_ENC/us03/n664 ), .ZN(\AES_ENC/us03/n666 ) );
NAND2_X2 \AES_ENC/us03/U429  ( .A1(\AES_ENC/sa03 [6]), .A2(\AES_ENC/us03/n666 ), .ZN(\AES_ENC/us03/n678 ) );
NAND2_X2 \AES_ENC/us03/U426  ( .A1(\AES_ENC/us03/n735 ), .A2(\AES_ENC/us03/n1093 ), .ZN(\AES_ENC/us03/n675 ) );
NAND2_X2 \AES_ENC/us03/U425  ( .A1(\AES_ENC/us03/n600 ), .A2(\AES_ENC/us03/n609 ), .ZN(\AES_ENC/us03/n1045 ) );
OR2_X2 \AES_ENC/us03/U424  ( .A1(\AES_ENC/us03/n1045 ), .A2(\AES_ENC/us03/n587 ), .ZN(\AES_ENC/us03/n674 ) );
NAND2_X2 \AES_ENC/us03/U423  ( .A1(\AES_ENC/sa03 [1]), .A2(\AES_ENC/us03/n622 ), .ZN(\AES_ENC/us03/n667 ) );
NAND2_X2 \AES_ENC/us03/U422  ( .A1(\AES_ENC/us03/n621 ), .A2(\AES_ENC/us03/n667 ), .ZN(\AES_ENC/us03/n1071 ) );
NAND4_X2 \AES_ENC/us03/U412  ( .A1(\AES_ENC/us03/n675 ), .A2(\AES_ENC/us03/n674 ), .A3(\AES_ENC/us03/n673 ), .A4(\AES_ENC/us03/n672 ), .ZN(\AES_ENC/us03/n676 ) );
NAND2_X2 \AES_ENC/us03/U411  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n676 ), .ZN(\AES_ENC/us03/n677 ) );
NAND2_X2 \AES_ENC/us03/U408  ( .A1(\AES_ENC/us03/n800 ), .A2(\AES_ENC/us03/n1022 ), .ZN(\AES_ENC/us03/n680 ) );
NAND2_X2 \AES_ENC/us03/U407  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n680 ), .ZN(\AES_ENC/us03/n681 ) );
AND2_X2 \AES_ENC/us03/U402  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n684 ), .ZN(\AES_ENC/us03/n682 ) );
NAND4_X2 \AES_ENC/us03/U395  ( .A1(\AES_ENC/us03/n691 ), .A2(\AES_ENC/us03/n584 ), .A3(\AES_ENC/us03/n690 ), .A4(\AES_ENC/us03/n689 ), .ZN(\AES_ENC/us03/n692 ) );
NAND2_X2 \AES_ENC/us03/U394  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n692 ), .ZN(\AES_ENC/us03/n733 ) );
NAND2_X2 \AES_ENC/us03/U392  ( .A1(\AES_ENC/us03/n977 ), .A2(\AES_ENC/us03/n1050 ), .ZN(\AES_ENC/us03/n702 ) );
NAND2_X2 \AES_ENC/us03/U391  ( .A1(\AES_ENC/us03/n1093 ), .A2(\AES_ENC/us03/n1045 ), .ZN(\AES_ENC/us03/n701 ) );
NAND4_X2 \AES_ENC/us03/U381  ( .A1(\AES_ENC/us03/n702 ), .A2(\AES_ENC/us03/n701 ), .A3(\AES_ENC/us03/n700 ), .A4(\AES_ENC/us03/n699 ), .ZN(\AES_ENC/us03/n703 ) );
NAND2_X2 \AES_ENC/us03/U380  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n703 ), .ZN(\AES_ENC/us03/n732 ) );
AND2_X2 \AES_ENC/us03/U379  ( .A1(\AES_ENC/sa03 [0]), .A2(\AES_ENC/sa03 [6]),.ZN(\AES_ENC/us03/n1113 ) );
NAND2_X2 \AES_ENC/us03/U378  ( .A1(\AES_ENC/us03/n613 ), .A2(\AES_ENC/us03/n1030 ), .ZN(\AES_ENC/us03/n881 ) );
NAND2_X2 \AES_ENC/us03/U377  ( .A1(\AES_ENC/us03/n1093 ), .A2(\AES_ENC/us03/n881 ), .ZN(\AES_ENC/us03/n715 ) );
NAND2_X2 \AES_ENC/us03/U376  ( .A1(\AES_ENC/us03/n1010 ), .A2(\AES_ENC/us03/n612 ), .ZN(\AES_ENC/us03/n714 ) );
NAND2_X2 \AES_ENC/us03/U375  ( .A1(\AES_ENC/us03/n855 ), .A2(\AES_ENC/us03/n600 ), .ZN(\AES_ENC/us03/n1117 ) );
XNOR2_X2 \AES_ENC/us03/U371  ( .A(\AES_ENC/us03/n618 ), .B(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n824 ) );
NAND4_X2 \AES_ENC/us03/U362  ( .A1(\AES_ENC/us03/n715 ), .A2(\AES_ENC/us03/n714 ), .A3(\AES_ENC/us03/n713 ), .A4(\AES_ENC/us03/n712 ), .ZN(\AES_ENC/us03/n716 ) );
NAND2_X2 \AES_ENC/us03/U361  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n716 ), .ZN(\AES_ENC/us03/n731 ) );
AND2_X2 \AES_ENC/us03/U360  ( .A1(\AES_ENC/sa03 [6]), .A2(\AES_ENC/us03/n574 ), .ZN(\AES_ENC/us03/n1131 ) );
NAND2_X2 \AES_ENC/us03/U359  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n717 ) );
NAND2_X2 \AES_ENC/us03/U358  ( .A1(\AES_ENC/us03/n1029 ), .A2(\AES_ENC/us03/n717 ), .ZN(\AES_ENC/us03/n728 ) );
NAND2_X2 \AES_ENC/us03/U357  ( .A1(\AES_ENC/sa03 [1]), .A2(\AES_ENC/us03/n626 ), .ZN(\AES_ENC/us03/n1097 ) );
NAND2_X2 \AES_ENC/us03/U356  ( .A1(\AES_ENC/us03/n615 ), .A2(\AES_ENC/us03/n1097 ), .ZN(\AES_ENC/us03/n718 ) );
NAND2_X2 \AES_ENC/us03/U355  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n718 ), .ZN(\AES_ENC/us03/n727 ) );
NAND4_X2 \AES_ENC/us03/U344  ( .A1(\AES_ENC/us03/n728 ), .A2(\AES_ENC/us03/n727 ), .A3(\AES_ENC/us03/n726 ), .A4(\AES_ENC/us03/n725 ), .ZN(\AES_ENC/us03/n729 ) );
NAND2_X2 \AES_ENC/us03/U343  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n729 ), .ZN(\AES_ENC/us03/n730 ) );
NAND4_X2 \AES_ENC/us03/U342  ( .A1(\AES_ENC/us03/n733 ), .A2(\AES_ENC/us03/n732 ), .A3(\AES_ENC/us03/n731 ), .A4(\AES_ENC/us03/n730 ), .ZN(\AES_ENC/sa03_sub[1] ) );
NAND2_X2 \AES_ENC/us03/U341  ( .A1(\AES_ENC/sa03 [7]), .A2(\AES_ENC/us03/n618 ), .ZN(\AES_ENC/us03/n734 ) );
NAND2_X2 \AES_ENC/us03/U340  ( .A1(\AES_ENC/us03/n734 ), .A2(\AES_ENC/us03/n589 ), .ZN(\AES_ENC/us03/n738 ) );
OR4_X2 \AES_ENC/us03/U339  ( .A1(\AES_ENC/us03/n738 ), .A2(\AES_ENC/us03/n627 ), .A3(\AES_ENC/us03/n826 ), .A4(\AES_ENC/us03/n1121 ), .ZN(\AES_ENC/us03/n746 ) );
NAND2_X2 \AES_ENC/us03/U337  ( .A1(\AES_ENC/us03/n1100 ), .A2(\AES_ENC/us03/n599 ), .ZN(\AES_ENC/us03/n992 ) );
OR2_X2 \AES_ENC/us03/U336  ( .A1(\AES_ENC/us03/n617 ), .A2(\AES_ENC/us03/n735 ), .ZN(\AES_ENC/us03/n737 ) );
NAND2_X2 \AES_ENC/us03/U334  ( .A1(\AES_ENC/us03/n621 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n753 ) );
NAND2_X2 \AES_ENC/us03/U333  ( .A1(\AES_ENC/us03/n595 ), .A2(\AES_ENC/us03/n753 ), .ZN(\AES_ENC/us03/n1080 ) );
NAND2_X2 \AES_ENC/us03/U332  ( .A1(\AES_ENC/us03/n1048 ), .A2(\AES_ENC/us03/n591 ), .ZN(\AES_ENC/us03/n736 ) );
NAND2_X2 \AES_ENC/us03/U331  ( .A1(\AES_ENC/us03/n737 ), .A2(\AES_ENC/us03/n736 ), .ZN(\AES_ENC/us03/n739 ) );
NAND2_X2 \AES_ENC/us03/U330  ( .A1(\AES_ENC/us03/n739 ), .A2(\AES_ENC/us03/n738 ), .ZN(\AES_ENC/us03/n745 ) );
NAND2_X2 \AES_ENC/us03/U326  ( .A1(\AES_ENC/us03/n1096 ), .A2(\AES_ENC/us03/n602 ), .ZN(\AES_ENC/us03/n906 ) );
NAND4_X2 \AES_ENC/us03/U323  ( .A1(\AES_ENC/us03/n746 ), .A2(\AES_ENC/us03/n992 ), .A3(\AES_ENC/us03/n745 ), .A4(\AES_ENC/us03/n744 ), .ZN(\AES_ENC/us03/n747 ) );
NAND2_X2 \AES_ENC/us03/U322  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n747 ), .ZN(\AES_ENC/us03/n793 ) );
NAND2_X2 \AES_ENC/us03/U321  ( .A1(\AES_ENC/us03/n597 ), .A2(\AES_ENC/us03/n855 ), .ZN(\AES_ENC/us03/n748 ) );
NAND2_X2 \AES_ENC/us03/U320  ( .A1(\AES_ENC/us03/n956 ), .A2(\AES_ENC/us03/n748 ), .ZN(\AES_ENC/us03/n760 ) );
NAND2_X2 \AES_ENC/us03/U313  ( .A1(\AES_ENC/us03/n602 ), .A2(\AES_ENC/us03/n753 ), .ZN(\AES_ENC/us03/n1023 ) );
NAND4_X2 \AES_ENC/us03/U308  ( .A1(\AES_ENC/us03/n760 ), .A2(\AES_ENC/us03/n992 ), .A3(\AES_ENC/us03/n759 ), .A4(\AES_ENC/us03/n758 ), .ZN(\AES_ENC/us03/n761 ) );
NAND2_X2 \AES_ENC/us03/U307  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n761 ), .ZN(\AES_ENC/us03/n792 ) );
NAND2_X2 \AES_ENC/us03/U306  ( .A1(\AES_ENC/us03/n597 ), .A2(\AES_ENC/us03/n615 ), .ZN(\AES_ENC/us03/n989 ) );
NAND2_X2 \AES_ENC/us03/U305  ( .A1(\AES_ENC/us03/n1050 ), .A2(\AES_ENC/us03/n989 ), .ZN(\AES_ENC/us03/n777 ) );
NAND2_X2 \AES_ENC/us03/U304  ( .A1(\AES_ENC/us03/n1093 ), .A2(\AES_ENC/us03/n762 ), .ZN(\AES_ENC/us03/n776 ) );
XNOR2_X2 \AES_ENC/us03/U301  ( .A(\AES_ENC/sa03 [7]), .B(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n959 ) );
NAND4_X2 \AES_ENC/us03/U289  ( .A1(\AES_ENC/us03/n777 ), .A2(\AES_ENC/us03/n776 ), .A3(\AES_ENC/us03/n775 ), .A4(\AES_ENC/us03/n774 ), .ZN(\AES_ENC/us03/n778 ) );
NAND2_X2 \AES_ENC/us03/U288  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n778 ), .ZN(\AES_ENC/us03/n791 ) );
NAND2_X2 \AES_ENC/us03/U287  ( .A1(\AES_ENC/us03/n1056 ), .A2(\AES_ENC/us03/n1050 ), .ZN(\AES_ENC/us03/n788 ) );
NAND2_X2 \AES_ENC/us03/U286  ( .A1(\AES_ENC/us03/n1091 ), .A2(\AES_ENC/us03/n779 ), .ZN(\AES_ENC/us03/n787 ) );
NAND2_X2 \AES_ENC/us03/U285  ( .A1(\AES_ENC/us03/n956 ), .A2(\AES_ENC/sa03 [1]), .ZN(\AES_ENC/us03/n786 ) );
NAND4_X2 \AES_ENC/us03/U278  ( .A1(\AES_ENC/us03/n788 ), .A2(\AES_ENC/us03/n787 ), .A3(\AES_ENC/us03/n786 ), .A4(\AES_ENC/us03/n785 ), .ZN(\AES_ENC/us03/n789 ) );
NAND2_X2 \AES_ENC/us03/U277  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n789 ), .ZN(\AES_ENC/us03/n790 ) );
NAND4_X2 \AES_ENC/us03/U276  ( .A1(\AES_ENC/us03/n793 ), .A2(\AES_ENC/us03/n792 ), .A3(\AES_ENC/us03/n791 ), .A4(\AES_ENC/us03/n790 ), .ZN(\AES_ENC/sa03_sub[2] ) );
NAND2_X2 \AES_ENC/us03/U275  ( .A1(\AES_ENC/us03/n1059 ), .A2(\AES_ENC/us03/n794 ), .ZN(\AES_ENC/us03/n810 ) );
NAND2_X2 \AES_ENC/us03/U274  ( .A1(\AES_ENC/us03/n1049 ), .A2(\AES_ENC/us03/n956 ), .ZN(\AES_ENC/us03/n809 ) );
OR2_X2 \AES_ENC/us03/U266  ( .A1(\AES_ENC/us03/n1096 ), .A2(\AES_ENC/us03/n588 ), .ZN(\AES_ENC/us03/n802 ) );
NAND2_X2 \AES_ENC/us03/U265  ( .A1(\AES_ENC/us03/n1053 ), .A2(\AES_ENC/us03/n800 ), .ZN(\AES_ENC/us03/n801 ) );
NAND2_X2 \AES_ENC/us03/U264  ( .A1(\AES_ENC/us03/n802 ), .A2(\AES_ENC/us03/n801 ), .ZN(\AES_ENC/us03/n805 ) );
NAND4_X2 \AES_ENC/us03/U261  ( .A1(\AES_ENC/us03/n810 ), .A2(\AES_ENC/us03/n809 ), .A3(\AES_ENC/us03/n808 ), .A4(\AES_ENC/us03/n807 ), .ZN(\AES_ENC/us03/n811 ) );
NAND2_X2 \AES_ENC/us03/U260  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n811 ), .ZN(\AES_ENC/us03/n852 ) );
OR2_X2 \AES_ENC/us03/U259  ( .A1(\AES_ENC/us03/n1023 ), .A2(\AES_ENC/us03/n576 ), .ZN(\AES_ENC/us03/n819 ) );
OR2_X2 \AES_ENC/us03/U257  ( .A1(\AES_ENC/us03/n570 ), .A2(\AES_ENC/us03/n930 ), .ZN(\AES_ENC/us03/n818 ) );
NAND2_X2 \AES_ENC/us03/U256  ( .A1(\AES_ENC/us03/n1013 ), .A2(\AES_ENC/us03/n1094 ), .ZN(\AES_ENC/us03/n817 ) );
NAND4_X2 \AES_ENC/us03/U249  ( .A1(\AES_ENC/us03/n819 ), .A2(\AES_ENC/us03/n818 ), .A3(\AES_ENC/us03/n817 ), .A4(\AES_ENC/us03/n816 ), .ZN(\AES_ENC/us03/n820 ) );
NAND2_X2 \AES_ENC/us03/U248  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n820 ), .ZN(\AES_ENC/us03/n851 ) );
NAND2_X2 \AES_ENC/us03/U247  ( .A1(\AES_ENC/us03/n956 ), .A2(\AES_ENC/us03/n1080 ), .ZN(\AES_ENC/us03/n835 ) );
NAND2_X2 \AES_ENC/us03/U246  ( .A1(\AES_ENC/us03/n570 ), .A2(\AES_ENC/us03/n1030 ), .ZN(\AES_ENC/us03/n1047 ) );
OR2_X2 \AES_ENC/us03/U245  ( .A1(\AES_ENC/us03/n1047 ), .A2(\AES_ENC/us03/n583 ), .ZN(\AES_ENC/us03/n834 ) );
NAND2_X2 \AES_ENC/us03/U244  ( .A1(\AES_ENC/us03/n1072 ), .A2(\AES_ENC/us03/n601 ), .ZN(\AES_ENC/us03/n833 ) );
NAND4_X2 \AES_ENC/us03/U233  ( .A1(\AES_ENC/us03/n835 ), .A2(\AES_ENC/us03/n834 ), .A3(\AES_ENC/us03/n833 ), .A4(\AES_ENC/us03/n832 ), .ZN(\AES_ENC/us03/n836 ) );
NAND2_X2 \AES_ENC/us03/U232  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n836 ), .ZN(\AES_ENC/us03/n850 ) );
NAND2_X2 \AES_ENC/us03/U231  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n625 ), .ZN(\AES_ENC/us03/n847 ) );
NAND2_X2 \AES_ENC/us03/U230  ( .A1(\AES_ENC/us03/n1050 ), .A2(\AES_ENC/us03/n1071 ), .ZN(\AES_ENC/us03/n846 ) );
OR2_X2 \AES_ENC/us03/U224  ( .A1(\AES_ENC/us03/n1053 ), .A2(\AES_ENC/us03/n911 ), .ZN(\AES_ENC/us03/n1077 ) );
NAND4_X2 \AES_ENC/us03/U220  ( .A1(\AES_ENC/us03/n847 ), .A2(\AES_ENC/us03/n846 ), .A3(\AES_ENC/us03/n845 ), .A4(\AES_ENC/us03/n844 ), .ZN(\AES_ENC/us03/n848 ) );
NAND2_X2 \AES_ENC/us03/U219  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n848 ), .ZN(\AES_ENC/us03/n849 ) );
NAND4_X2 \AES_ENC/us03/U218  ( .A1(\AES_ENC/us03/n852 ), .A2(\AES_ENC/us03/n851 ), .A3(\AES_ENC/us03/n850 ), .A4(\AES_ENC/us03/n849 ), .ZN(\AES_ENC/sa03_sub[3] ) );
NAND2_X2 \AES_ENC/us03/U216  ( .A1(\AES_ENC/us03/n1009 ), .A2(\AES_ENC/us03/n1072 ), .ZN(\AES_ENC/us03/n862 ) );
NAND2_X2 \AES_ENC/us03/U215  ( .A1(\AES_ENC/us03/n615 ), .A2(\AES_ENC/us03/n592 ), .ZN(\AES_ENC/us03/n853 ) );
NAND2_X2 \AES_ENC/us03/U214  ( .A1(\AES_ENC/us03/n1050 ), .A2(\AES_ENC/us03/n853 ), .ZN(\AES_ENC/us03/n861 ) );
NAND4_X2 \AES_ENC/us03/U206  ( .A1(\AES_ENC/us03/n862 ), .A2(\AES_ENC/us03/n861 ), .A3(\AES_ENC/us03/n860 ), .A4(\AES_ENC/us03/n859 ), .ZN(\AES_ENC/us03/n863 ) );
NAND2_X2 \AES_ENC/us03/U205  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n863 ), .ZN(\AES_ENC/us03/n905 ) );
NAND2_X2 \AES_ENC/us03/U204  ( .A1(\AES_ENC/us03/n1010 ), .A2(\AES_ENC/us03/n989 ), .ZN(\AES_ENC/us03/n874 ) );
NAND2_X2 \AES_ENC/us03/U203  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n617 ), .ZN(\AES_ENC/us03/n864 ) );
NAND2_X2 \AES_ENC/us03/U202  ( .A1(\AES_ENC/us03/n929 ), .A2(\AES_ENC/us03/n864 ), .ZN(\AES_ENC/us03/n873 ) );
NAND4_X2 \AES_ENC/us03/U193  ( .A1(\AES_ENC/us03/n874 ), .A2(\AES_ENC/us03/n873 ), .A3(\AES_ENC/us03/n872 ), .A4(\AES_ENC/us03/n871 ), .ZN(\AES_ENC/us03/n875 ) );
NAND2_X2 \AES_ENC/us03/U192  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n875 ), .ZN(\AES_ENC/us03/n904 ) );
NAND2_X2 \AES_ENC/us03/U191  ( .A1(\AES_ENC/us03/n596 ), .A2(\AES_ENC/us03/n1050 ), .ZN(\AES_ENC/us03/n889 ) );
NAND2_X2 \AES_ENC/us03/U190  ( .A1(\AES_ENC/us03/n1093 ), .A2(\AES_ENC/us03/n599 ), .ZN(\AES_ENC/us03/n876 ) );
NAND2_X2 \AES_ENC/us03/U189  ( .A1(\AES_ENC/us03/n577 ), .A2(\AES_ENC/us03/n876 ), .ZN(\AES_ENC/us03/n877 ) );
NAND2_X2 \AES_ENC/us03/U188  ( .A1(\AES_ENC/us03/n877 ), .A2(\AES_ENC/us03/n625 ), .ZN(\AES_ENC/us03/n888 ) );
NAND4_X2 \AES_ENC/us03/U179  ( .A1(\AES_ENC/us03/n889 ), .A2(\AES_ENC/us03/n888 ), .A3(\AES_ENC/us03/n887 ), .A4(\AES_ENC/us03/n886 ), .ZN(\AES_ENC/us03/n890 ) );
NAND2_X2 \AES_ENC/us03/U178  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n890 ), .ZN(\AES_ENC/us03/n903 ) );
OR2_X2 \AES_ENC/us03/U177  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n1059 ), .ZN(\AES_ENC/us03/n900 ) );
NAND2_X2 \AES_ENC/us03/U176  ( .A1(\AES_ENC/us03/n1073 ), .A2(\AES_ENC/us03/n1047 ), .ZN(\AES_ENC/us03/n899 ) );
NAND2_X2 \AES_ENC/us03/U175  ( .A1(\AES_ENC/us03/n1094 ), .A2(\AES_ENC/us03/n607 ), .ZN(\AES_ENC/us03/n898 ) );
NAND4_X2 \AES_ENC/us03/U167  ( .A1(\AES_ENC/us03/n900 ), .A2(\AES_ENC/us03/n899 ), .A3(\AES_ENC/us03/n898 ), .A4(\AES_ENC/us03/n897 ), .ZN(\AES_ENC/us03/n901 ) );
NAND2_X2 \AES_ENC/us03/U166  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n901 ), .ZN(\AES_ENC/us03/n902 ) );
NAND4_X2 \AES_ENC/us03/U165  ( .A1(\AES_ENC/us03/n905 ), .A2(\AES_ENC/us03/n904 ), .A3(\AES_ENC/us03/n903 ), .A4(\AES_ENC/us03/n902 ), .ZN(\AES_ENC/sa03_sub[4] ) );
NAND2_X2 \AES_ENC/us03/U164  ( .A1(\AES_ENC/us03/n1094 ), .A2(\AES_ENC/us03/n611 ), .ZN(\AES_ENC/us03/n922 ) );
NAND2_X2 \AES_ENC/us03/U163  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n989 ), .ZN(\AES_ENC/us03/n921 ) );
NAND4_X2 \AES_ENC/us03/U151  ( .A1(\AES_ENC/us03/n922 ), .A2(\AES_ENC/us03/n921 ), .A3(\AES_ENC/us03/n920 ), .A4(\AES_ENC/us03/n919 ), .ZN(\AES_ENC/us03/n923 ) );
NAND2_X2 \AES_ENC/us03/U150  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n923 ), .ZN(\AES_ENC/us03/n972 ) );
NAND2_X2 \AES_ENC/us03/U149  ( .A1(\AES_ENC/us03/n595 ), .A2(\AES_ENC/us03/n621 ), .ZN(\AES_ENC/us03/n924 ) );
NAND2_X2 \AES_ENC/us03/U148  ( .A1(\AES_ENC/us03/n1073 ), .A2(\AES_ENC/us03/n924 ), .ZN(\AES_ENC/us03/n939 ) );
NAND2_X2 \AES_ENC/us03/U147  ( .A1(\AES_ENC/us03/n926 ), .A2(\AES_ENC/us03/n925 ), .ZN(\AES_ENC/us03/n927 ) );
NAND2_X2 \AES_ENC/us03/U146  ( .A1(\AES_ENC/us03/n588 ), .A2(\AES_ENC/us03/n927 ), .ZN(\AES_ENC/us03/n928 ) );
NAND2_X2 \AES_ENC/us03/U145  ( .A1(\AES_ENC/us03/n928 ), .A2(\AES_ENC/us03/n1080 ), .ZN(\AES_ENC/us03/n938 ) );
OR2_X2 \AES_ENC/us03/U144  ( .A1(\AES_ENC/us03/n1117 ), .A2(\AES_ENC/us03/n581 ), .ZN(\AES_ENC/us03/n937 ) );
NAND4_X2 \AES_ENC/us03/U139  ( .A1(\AES_ENC/us03/n939 ), .A2(\AES_ENC/us03/n938 ), .A3(\AES_ENC/us03/n937 ), .A4(\AES_ENC/us03/n936 ), .ZN(\AES_ENC/us03/n940 ) );
NAND2_X2 \AES_ENC/us03/U138  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n940 ), .ZN(\AES_ENC/us03/n971 ) );
OR2_X2 \AES_ENC/us03/U137  ( .A1(\AES_ENC/us03/n587 ), .A2(\AES_ENC/us03/n941 ), .ZN(\AES_ENC/us03/n954 ) );
NAND2_X2 \AES_ENC/us03/U136  ( .A1(\AES_ENC/us03/n1096 ), .A2(\AES_ENC/us03/n592 ), .ZN(\AES_ENC/us03/n942 ) );
NAND2_X2 \AES_ENC/us03/U135  ( .A1(\AES_ENC/us03/n1048 ), .A2(\AES_ENC/us03/n942 ), .ZN(\AES_ENC/us03/n943 ) );
NAND2_X2 \AES_ENC/us03/U134  ( .A1(\AES_ENC/us03/n583 ), .A2(\AES_ENC/us03/n943 ), .ZN(\AES_ENC/us03/n944 ) );
NAND2_X2 \AES_ENC/us03/U133  ( .A1(\AES_ENC/us03/n944 ), .A2(\AES_ENC/us03/n594 ), .ZN(\AES_ENC/us03/n953 ) );
NAND4_X2 \AES_ENC/us03/U125  ( .A1(\AES_ENC/us03/n954 ), .A2(\AES_ENC/us03/n953 ), .A3(\AES_ENC/us03/n952 ), .A4(\AES_ENC/us03/n951 ), .ZN(\AES_ENC/us03/n955 ) );
NAND2_X2 \AES_ENC/us03/U124  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n955 ), .ZN(\AES_ENC/us03/n970 ) );
NAND2_X2 \AES_ENC/us03/U123  ( .A1(\AES_ENC/us03/n1094 ), .A2(\AES_ENC/us03/n1071 ), .ZN(\AES_ENC/us03/n967 ) );
NAND2_X2 \AES_ENC/us03/U122  ( .A1(\AES_ENC/us03/n956 ), .A2(\AES_ENC/us03/n1030 ), .ZN(\AES_ENC/us03/n966 ) );
NAND4_X2 \AES_ENC/us03/U114  ( .A1(\AES_ENC/us03/n967 ), .A2(\AES_ENC/us03/n966 ), .A3(\AES_ENC/us03/n965 ), .A4(\AES_ENC/us03/n964 ), .ZN(\AES_ENC/us03/n968 ) );
NAND2_X2 \AES_ENC/us03/U113  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n968 ), .ZN(\AES_ENC/us03/n969 ) );
NAND4_X2 \AES_ENC/us03/U112  ( .A1(\AES_ENC/us03/n972 ), .A2(\AES_ENC/us03/n971 ), .A3(\AES_ENC/us03/n970 ), .A4(\AES_ENC/us03/n969 ), .ZN(\AES_ENC/sa03_sub[5] ) );
NAND2_X2 \AES_ENC/us03/U111  ( .A1(\AES_ENC/us03/n570 ), .A2(\AES_ENC/us03/n1097 ), .ZN(\AES_ENC/us03/n973 ) );
NAND2_X2 \AES_ENC/us03/U110  ( .A1(\AES_ENC/us03/n1073 ), .A2(\AES_ENC/us03/n973 ), .ZN(\AES_ENC/us03/n987 ) );
NAND2_X2 \AES_ENC/us03/U109  ( .A1(\AES_ENC/us03/n974 ), .A2(\AES_ENC/us03/n1077 ), .ZN(\AES_ENC/us03/n975 ) );
NAND2_X2 \AES_ENC/us03/U108  ( .A1(\AES_ENC/us03/n585 ), .A2(\AES_ENC/us03/n975 ), .ZN(\AES_ENC/us03/n976 ) );
NAND2_X2 \AES_ENC/us03/U107  ( .A1(\AES_ENC/us03/n977 ), .A2(\AES_ENC/us03/n976 ), .ZN(\AES_ENC/us03/n986 ) );
NAND4_X2 \AES_ENC/us03/U99  ( .A1(\AES_ENC/us03/n987 ), .A2(\AES_ENC/us03/n986 ), .A3(\AES_ENC/us03/n985 ), .A4(\AES_ENC/us03/n984 ), .ZN(\AES_ENC/us03/n988 ) );
NAND2_X2 \AES_ENC/us03/U98  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n988 ), .ZN(\AES_ENC/us03/n1044 ) );
NAND2_X2 \AES_ENC/us03/U97  ( .A1(\AES_ENC/us03/n1073 ), .A2(\AES_ENC/us03/n989 ), .ZN(\AES_ENC/us03/n1004 ) );
NAND2_X2 \AES_ENC/us03/U96  ( .A1(\AES_ENC/us03/n1092 ), .A2(\AES_ENC/us03/n621 ), .ZN(\AES_ENC/us03/n1003 ) );
NAND4_X2 \AES_ENC/us03/U85  ( .A1(\AES_ENC/us03/n1004 ), .A2(\AES_ENC/us03/n1003 ), .A3(\AES_ENC/us03/n1002 ), .A4(\AES_ENC/us03/n1001 ), .ZN(\AES_ENC/us03/n1005 ) );
NAND2_X2 \AES_ENC/us03/U84  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n1005 ), .ZN(\AES_ENC/us03/n1043 ) );
NAND2_X2 \AES_ENC/us03/U83  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n608 ), .ZN(\AES_ENC/us03/n1020 ) );
NAND2_X2 \AES_ENC/us03/U82  ( .A1(\AES_ENC/us03/n1050 ), .A2(\AES_ENC/us03/n626 ), .ZN(\AES_ENC/us03/n1019 ) );
NAND2_X2 \AES_ENC/us03/U77  ( .A1(\AES_ENC/us03/n1059 ), .A2(\AES_ENC/us03/n1114 ), .ZN(\AES_ENC/us03/n1012 ) );
NAND2_X2 \AES_ENC/us03/U76  ( .A1(\AES_ENC/us03/n1010 ), .A2(\AES_ENC/us03/n604 ), .ZN(\AES_ENC/us03/n1011 ) );
NAND2_X2 \AES_ENC/us03/U75  ( .A1(\AES_ENC/us03/n1012 ), .A2(\AES_ENC/us03/n1011 ), .ZN(\AES_ENC/us03/n1016 ) );
NAND4_X2 \AES_ENC/us03/U70  ( .A1(\AES_ENC/us03/n1020 ), .A2(\AES_ENC/us03/n1019 ), .A3(\AES_ENC/us03/n1018 ), .A4(\AES_ENC/us03/n1017 ), .ZN(\AES_ENC/us03/n1021 ) );
NAND2_X2 \AES_ENC/us03/U69  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n1021 ), .ZN(\AES_ENC/us03/n1042 ) );
NAND2_X2 \AES_ENC/us03/U68  ( .A1(\AES_ENC/us03/n1022 ), .A2(\AES_ENC/us03/n1093 ), .ZN(\AES_ENC/us03/n1039 ) );
NAND2_X2 \AES_ENC/us03/U67  ( .A1(\AES_ENC/us03/n1050 ), .A2(\AES_ENC/us03/n1023 ), .ZN(\AES_ENC/us03/n1038 ) );
NAND2_X2 \AES_ENC/us03/U66  ( .A1(\AES_ENC/us03/n1024 ), .A2(\AES_ENC/us03/n1071 ), .ZN(\AES_ENC/us03/n1037 ) );
AND2_X2 \AES_ENC/us03/U60  ( .A1(\AES_ENC/us03/n1030 ), .A2(\AES_ENC/us03/n614 ), .ZN(\AES_ENC/us03/n1078 ) );
NAND4_X2 \AES_ENC/us03/U56  ( .A1(\AES_ENC/us03/n1039 ), .A2(\AES_ENC/us03/n1038 ), .A3(\AES_ENC/us03/n1037 ), .A4(\AES_ENC/us03/n1036 ), .ZN(\AES_ENC/us03/n1040 ) );
NAND2_X2 \AES_ENC/us03/U55  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n1040 ), .ZN(\AES_ENC/us03/n1041 ) );
NAND4_X2 \AES_ENC/us03/U54  ( .A1(\AES_ENC/us03/n1044 ), .A2(\AES_ENC/us03/n1043 ), .A3(\AES_ENC/us03/n1042 ), .A4(\AES_ENC/us03/n1041 ), .ZN(\AES_ENC/sa03_sub[6] ) );
NAND2_X2 \AES_ENC/us03/U53  ( .A1(\AES_ENC/us03/n1072 ), .A2(\AES_ENC/us03/n1045 ), .ZN(\AES_ENC/us03/n1068 ) );
NAND2_X2 \AES_ENC/us03/U52  ( .A1(\AES_ENC/us03/n1046 ), .A2(\AES_ENC/us03/n595 ), .ZN(\AES_ENC/us03/n1067 ) );
NAND2_X2 \AES_ENC/us03/U51  ( .A1(\AES_ENC/us03/n1094 ), .A2(\AES_ENC/us03/n1047 ), .ZN(\AES_ENC/us03/n1066 ) );
NAND4_X2 \AES_ENC/us03/U40  ( .A1(\AES_ENC/us03/n1068 ), .A2(\AES_ENC/us03/n1067 ), .A3(\AES_ENC/us03/n1066 ), .A4(\AES_ENC/us03/n1065 ), .ZN(\AES_ENC/us03/n1069 ) );
NAND2_X2 \AES_ENC/us03/U39  ( .A1(\AES_ENC/us03/n1070 ), .A2(\AES_ENC/us03/n1069 ), .ZN(\AES_ENC/us03/n1135 ) );
NAND2_X2 \AES_ENC/us03/U38  ( .A1(\AES_ENC/us03/n1072 ), .A2(\AES_ENC/us03/n1071 ), .ZN(\AES_ENC/us03/n1088 ) );
NAND2_X2 \AES_ENC/us03/U37  ( .A1(\AES_ENC/us03/n1073 ), .A2(\AES_ENC/us03/n607 ), .ZN(\AES_ENC/us03/n1087 ) );
NAND4_X2 \AES_ENC/us03/U28  ( .A1(\AES_ENC/us03/n1088 ), .A2(\AES_ENC/us03/n1087 ), .A3(\AES_ENC/us03/n1086 ), .A4(\AES_ENC/us03/n1085 ), .ZN(\AES_ENC/us03/n1089 ) );
NAND2_X2 \AES_ENC/us03/U27  ( .A1(\AES_ENC/us03/n1090 ), .A2(\AES_ENC/us03/n1089 ), .ZN(\AES_ENC/us03/n1134 ) );
NAND2_X2 \AES_ENC/us03/U26  ( .A1(\AES_ENC/us03/n1091 ), .A2(\AES_ENC/us03/n1093 ), .ZN(\AES_ENC/us03/n1111 ) );
NAND2_X2 \AES_ENC/us03/U25  ( .A1(\AES_ENC/us03/n1092 ), .A2(\AES_ENC/us03/n1120 ), .ZN(\AES_ENC/us03/n1110 ) );
AND2_X2 \AES_ENC/us03/U22  ( .A1(\AES_ENC/us03/n1097 ), .A2(\AES_ENC/us03/n1096 ), .ZN(\AES_ENC/us03/n1098 ) );
NAND4_X2 \AES_ENC/us03/U14  ( .A1(\AES_ENC/us03/n1111 ), .A2(\AES_ENC/us03/n1110 ), .A3(\AES_ENC/us03/n1109 ), .A4(\AES_ENC/us03/n1108 ), .ZN(\AES_ENC/us03/n1112 ) );
NAND2_X2 \AES_ENC/us03/U13  ( .A1(\AES_ENC/us03/n1113 ), .A2(\AES_ENC/us03/n1112 ), .ZN(\AES_ENC/us03/n1133 ) );
NAND2_X2 \AES_ENC/us03/U12  ( .A1(\AES_ENC/us03/n1115 ), .A2(\AES_ENC/us03/n1114 ), .ZN(\AES_ENC/us03/n1129 ) );
OR2_X2 \AES_ENC/us03/U11  ( .A1(\AES_ENC/us03/n580 ), .A2(\AES_ENC/us03/n1116 ), .ZN(\AES_ENC/us03/n1128 ) );
NAND4_X2 \AES_ENC/us03/U3  ( .A1(\AES_ENC/us03/n1129 ), .A2(\AES_ENC/us03/n1128 ), .A3(\AES_ENC/us03/n1127 ), .A4(\AES_ENC/us03/n1126 ), .ZN(\AES_ENC/us03/n1130 ) );
NAND2_X2 \AES_ENC/us03/U2  ( .A1(\AES_ENC/us03/n1131 ), .A2(\AES_ENC/us03/n1130 ), .ZN(\AES_ENC/us03/n1132 ) );
NAND4_X2 \AES_ENC/us03/U1  ( .A1(\AES_ENC/us03/n1135 ), .A2(\AES_ENC/us03/n1134 ), .A3(\AES_ENC/us03/n1133 ), .A4(\AES_ENC/us03/n1132 ), .ZN(\AES_ENC/sa03_sub[7] ) );
INV_X4 \AES_ENC/us10/U575  ( .A(\AES_ENC/sa10 [7]), .ZN(\AES_ENC/us10/n627 ));
INV_X4 \AES_ENC/us10/U574  ( .A(\AES_ENC/us10/n1114 ), .ZN(\AES_ENC/us10/n625 ) );
INV_X4 \AES_ENC/us10/U573  ( .A(\AES_ENC/sa10 [4]), .ZN(\AES_ENC/us10/n624 ));
INV_X4 \AES_ENC/us10/U572  ( .A(\AES_ENC/us10/n1025 ), .ZN(\AES_ENC/us10/n622 ) );
INV_X4 \AES_ENC/us10/U571  ( .A(\AES_ENC/us10/n1120 ), .ZN(\AES_ENC/us10/n620 ) );
INV_X4 \AES_ENC/us10/U570  ( .A(\AES_ENC/us10/n1121 ), .ZN(\AES_ENC/us10/n619 ) );
INV_X4 \AES_ENC/us10/U569  ( .A(\AES_ENC/us10/n1048 ), .ZN(\AES_ENC/us10/n618 ) );
INV_X4 \AES_ENC/us10/U568  ( .A(\AES_ENC/us10/n974 ), .ZN(\AES_ENC/us10/n616 ) );
INV_X4 \AES_ENC/us10/U567  ( .A(\AES_ENC/us10/n794 ), .ZN(\AES_ENC/us10/n614 ) );
INV_X4 \AES_ENC/us10/U566  ( .A(\AES_ENC/sa10 [2]), .ZN(\AES_ENC/us10/n611 ));
INV_X4 \AES_ENC/us10/U565  ( .A(\AES_ENC/us10/n800 ), .ZN(\AES_ENC/us10/n610 ) );
INV_X4 \AES_ENC/us10/U564  ( .A(\AES_ENC/us10/n925 ), .ZN(\AES_ENC/us10/n609 ) );
INV_X4 \AES_ENC/us10/U563  ( .A(\AES_ENC/us10/n779 ), .ZN(\AES_ENC/us10/n607 ) );
INV_X4 \AES_ENC/us10/U562  ( .A(\AES_ENC/us10/n1022 ), .ZN(\AES_ENC/us10/n603 ) );
INV_X4 \AES_ENC/us10/U561  ( .A(\AES_ENC/us10/n1102 ), .ZN(\AES_ENC/us10/n602 ) );
INV_X4 \AES_ENC/us10/U560  ( .A(\AES_ENC/us10/n929 ), .ZN(\AES_ENC/us10/n601 ) );
INV_X4 \AES_ENC/us10/U559  ( .A(\AES_ENC/us10/n1056 ), .ZN(\AES_ENC/us10/n600 ) );
INV_X4 \AES_ENC/us10/U558  ( .A(\AES_ENC/us10/n1054 ), .ZN(\AES_ENC/us10/n599 ) );
INV_X4 \AES_ENC/us10/U557  ( .A(\AES_ENC/us10/n881 ), .ZN(\AES_ENC/us10/n598 ) );
INV_X4 \AES_ENC/us10/U556  ( .A(\AES_ENC/us10/n926 ), .ZN(\AES_ENC/us10/n597 ) );
INV_X4 \AES_ENC/us10/U555  ( .A(\AES_ENC/us10/n977 ), .ZN(\AES_ENC/us10/n595 ) );
INV_X4 \AES_ENC/us10/U554  ( .A(\AES_ENC/us10/n1031 ), .ZN(\AES_ENC/us10/n594 ) );
INV_X4 \AES_ENC/us10/U553  ( .A(\AES_ENC/us10/n1103 ), .ZN(\AES_ENC/us10/n593 ) );
INV_X4 \AES_ENC/us10/U552  ( .A(\AES_ENC/us10/n1009 ), .ZN(\AES_ENC/us10/n592 ) );
INV_X4 \AES_ENC/us10/U551  ( .A(\AES_ENC/us10/n990 ), .ZN(\AES_ENC/us10/n591 ) );
INV_X4 \AES_ENC/us10/U550  ( .A(\AES_ENC/us10/n1058 ), .ZN(\AES_ENC/us10/n590 ) );
INV_X4 \AES_ENC/us10/U549  ( .A(\AES_ENC/us10/n1074 ), .ZN(\AES_ENC/us10/n589 ) );
INV_X4 \AES_ENC/us10/U548  ( .A(\AES_ENC/us10/n1053 ), .ZN(\AES_ENC/us10/n588 ) );
INV_X4 \AES_ENC/us10/U547  ( .A(\AES_ENC/us10/n826 ), .ZN(\AES_ENC/us10/n587 ) );
INV_X4 \AES_ENC/us10/U546  ( .A(\AES_ENC/us10/n992 ), .ZN(\AES_ENC/us10/n586 ) );
INV_X4 \AES_ENC/us10/U545  ( .A(\AES_ENC/us10/n821 ), .ZN(\AES_ENC/us10/n585 ) );
INV_X4 \AES_ENC/us10/U544  ( .A(\AES_ENC/us10/n910 ), .ZN(\AES_ENC/us10/n584 ) );
INV_X4 \AES_ENC/us10/U543  ( .A(\AES_ENC/us10/n906 ), .ZN(\AES_ENC/us10/n583 ) );
INV_X4 \AES_ENC/us10/U542  ( .A(\AES_ENC/us10/n880 ), .ZN(\AES_ENC/us10/n581 ) );
INV_X4 \AES_ENC/us10/U541  ( .A(\AES_ENC/us10/n1013 ), .ZN(\AES_ENC/us10/n580 ) );
INV_X4 \AES_ENC/us10/U540  ( .A(\AES_ENC/us10/n1092 ), .ZN(\AES_ENC/us10/n579 ) );
INV_X4 \AES_ENC/us10/U539  ( .A(\AES_ENC/us10/n824 ), .ZN(\AES_ENC/us10/n578 ) );
INV_X4 \AES_ENC/us10/U538  ( .A(\AES_ENC/us10/n1091 ), .ZN(\AES_ENC/us10/n577 ) );
INV_X4 \AES_ENC/us10/U537  ( .A(\AES_ENC/us10/n1080 ), .ZN(\AES_ENC/us10/n576 ) );
INV_X4 \AES_ENC/us10/U536  ( .A(\AES_ENC/us10/n959 ), .ZN(\AES_ENC/us10/n575 ) );
INV_X4 \AES_ENC/us10/U535  ( .A(\AES_ENC/sa10 [0]), .ZN(\AES_ENC/us10/n574 ));
NOR2_X2 \AES_ENC/us10/U534  ( .A1(\AES_ENC/sa10 [0]), .A2(\AES_ENC/sa10 [6]),.ZN(\AES_ENC/us10/n1090 ) );
NOR2_X2 \AES_ENC/us10/U533  ( .A1(\AES_ENC/us10/n574 ), .A2(\AES_ENC/sa10 [6]), .ZN(\AES_ENC/us10/n1070 ) );
NOR2_X2 \AES_ENC/us10/U532  ( .A1(\AES_ENC/sa10 [4]), .A2(\AES_ENC/sa10 [3]),.ZN(\AES_ENC/us10/n1025 ) );
INV_X4 \AES_ENC/us10/U531  ( .A(\AES_ENC/us10/n569 ), .ZN(\AES_ENC/us10/n572 ) );
NOR2_X2 \AES_ENC/us10/U530  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n765 ) );
NOR2_X2 \AES_ENC/us10/U529  ( .A1(\AES_ENC/sa10 [4]), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n764 ) );
NOR2_X2 \AES_ENC/us10/U528  ( .A1(\AES_ENC/us10/n765 ), .A2(\AES_ENC/us10/n764 ), .ZN(\AES_ENC/us10/n766 ) );
NOR2_X2 \AES_ENC/us10/U527  ( .A1(\AES_ENC/us10/n766 ), .A2(\AES_ENC/us10/n575 ), .ZN(\AES_ENC/us10/n767 ) );
NOR3_X2 \AES_ENC/us10/U526  ( .A1(\AES_ENC/us10/n627 ), .A2(\AES_ENC/sa10 [5]), .A3(\AES_ENC/us10/n704 ), .ZN(\AES_ENC/us10/n706 ));
NOR2_X2 \AES_ENC/us10/U525  ( .A1(\AES_ENC/us10/n1117 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n707 ) );
NOR2_X2 \AES_ENC/us10/U524  ( .A1(\AES_ENC/sa10 [4]), .A2(\AES_ENC/us10/n579 ), .ZN(\AES_ENC/us10/n705 ) );
NOR3_X2 \AES_ENC/us10/U523  ( .A1(\AES_ENC/us10/n707 ), .A2(\AES_ENC/us10/n706 ), .A3(\AES_ENC/us10/n705 ), .ZN(\AES_ENC/us10/n713 ) );
INV_X4 \AES_ENC/us10/U522  ( .A(\AES_ENC/sa10 [3]), .ZN(\AES_ENC/us10/n621 ));
NAND3_X2 \AES_ENC/us10/U521  ( .A1(\AES_ENC/us10/n652 ), .A2(\AES_ENC/us10/n626 ), .A3(\AES_ENC/sa10 [7]), .ZN(\AES_ENC/us10/n653 ));
NOR2_X2 \AES_ENC/us10/U520  ( .A1(\AES_ENC/us10/n611 ), .A2(\AES_ENC/sa10 [5]), .ZN(\AES_ENC/us10/n925 ) );
NOR2_X2 \AES_ENC/us10/U519  ( .A1(\AES_ENC/sa10 [5]), .A2(\AES_ENC/sa10 [2]),.ZN(\AES_ENC/us10/n974 ) );
INV_X4 \AES_ENC/us10/U518  ( .A(\AES_ENC/sa10 [5]), .ZN(\AES_ENC/us10/n626 ));
NOR2_X2 \AES_ENC/us10/U517  ( .A1(\AES_ENC/us10/n611 ), .A2(\AES_ENC/sa10 [7]), .ZN(\AES_ENC/us10/n779 ) );
NAND3_X2 \AES_ENC/us10/U516  ( .A1(\AES_ENC/us10/n679 ), .A2(\AES_ENC/us10/n678 ), .A3(\AES_ENC/us10/n677 ), .ZN(\AES_ENC/sa10_sub[0] ) );
NOR2_X2 \AES_ENC/us10/U515  ( .A1(\AES_ENC/us10/n626 ), .A2(\AES_ENC/sa10 [2]), .ZN(\AES_ENC/us10/n1048 ) );
NOR4_X2 \AES_ENC/us10/U512  ( .A1(\AES_ENC/us10/n633 ), .A2(\AES_ENC/us10/n632 ), .A3(\AES_ENC/us10/n631 ), .A4(\AES_ENC/us10/n630 ), .ZN(\AES_ENC/us10/n634 ) );
NOR2_X2 \AES_ENC/us10/U510  ( .A1(\AES_ENC/us10/n629 ), .A2(\AES_ENC/us10/n628 ), .ZN(\AES_ENC/us10/n635 ) );
NAND3_X2 \AES_ENC/us10/U509  ( .A1(\AES_ENC/sa10 [2]), .A2(\AES_ENC/sa10 [7]), .A3(\AES_ENC/us10/n1059 ), .ZN(\AES_ENC/us10/n636 ) );
NOR2_X2 \AES_ENC/us10/U508  ( .A1(\AES_ENC/sa10 [7]), .A2(\AES_ENC/sa10 [2]),.ZN(\AES_ENC/us10/n794 ) );
NOR2_X2 \AES_ENC/us10/U507  ( .A1(\AES_ENC/sa10 [4]), .A2(\AES_ENC/sa10 [1]),.ZN(\AES_ENC/us10/n1102 ) );
NOR2_X2 \AES_ENC/us10/U506  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/sa10 [3]), .ZN(\AES_ENC/us10/n1053 ) );
NOR2_X2 \AES_ENC/us10/U505  ( .A1(\AES_ENC/us10/n607 ), .A2(\AES_ENC/sa10 [5]), .ZN(\AES_ENC/us10/n1024 ) );
NOR2_X2 \AES_ENC/us10/U504  ( .A1(\AES_ENC/us10/n625 ), .A2(\AES_ENC/sa10 [2]), .ZN(\AES_ENC/us10/n1093 ) );
NOR2_X2 \AES_ENC/us10/U503  ( .A1(\AES_ENC/us10/n614 ), .A2(\AES_ENC/sa10 [5]), .ZN(\AES_ENC/us10/n1094 ) );
NOR2_X2 \AES_ENC/us10/U502  ( .A1(\AES_ENC/us10/n624 ), .A2(\AES_ENC/sa10 [3]), .ZN(\AES_ENC/us10/n931 ) );
INV_X4 \AES_ENC/us10/U501  ( .A(\AES_ENC/us10/n570 ), .ZN(\AES_ENC/us10/n573 ) );
NOR2_X2 \AES_ENC/us10/U500  ( .A1(\AES_ENC/us10/n1053 ), .A2(\AES_ENC/us10/n1095 ), .ZN(\AES_ENC/us10/n639 ) );
NOR3_X2 \AES_ENC/us10/U499  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n573 ), .A3(\AES_ENC/us10/n1074 ), .ZN(\AES_ENC/us10/n641 ) );
NOR2_X2 \AES_ENC/us10/U498  ( .A1(\AES_ENC/us10/n639 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n640 ) );
NOR2_X2 \AES_ENC/us10/U497  ( .A1(\AES_ENC/us10/n641 ), .A2(\AES_ENC/us10/n640 ), .ZN(\AES_ENC/us10/n646 ) );
NOR3_X2 \AES_ENC/us10/U496  ( .A1(\AES_ENC/us10/n995 ), .A2(\AES_ENC/us10/n586 ), .A3(\AES_ENC/us10/n994 ), .ZN(\AES_ENC/us10/n1002 ) );
NOR2_X2 \AES_ENC/us10/U495  ( .A1(\AES_ENC/us10/n909 ), .A2(\AES_ENC/us10/n908 ), .ZN(\AES_ENC/us10/n920 ) );
NOR2_X2 \AES_ENC/us10/U494  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n823 ) );
NOR2_X2 \AES_ENC/us10/U492  ( .A1(\AES_ENC/us10/n624 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n822 ) );
NOR2_X2 \AES_ENC/us10/U491  ( .A1(\AES_ENC/us10/n823 ), .A2(\AES_ENC/us10/n822 ), .ZN(\AES_ENC/us10/n825 ) );
NOR2_X2 \AES_ENC/us10/U490  ( .A1(\AES_ENC/sa10 [1]), .A2(\AES_ENC/us10/n623 ), .ZN(\AES_ENC/us10/n913 ) );
NOR2_X2 \AES_ENC/us10/U489  ( .A1(\AES_ENC/us10/n913 ), .A2(\AES_ENC/us10/n1091 ), .ZN(\AES_ENC/us10/n914 ) );
NOR2_X2 \AES_ENC/us10/U488  ( .A1(\AES_ENC/us10/n826 ), .A2(\AES_ENC/us10/n572 ), .ZN(\AES_ENC/us10/n827 ) );
NOR3_X2 \AES_ENC/us10/U487  ( .A1(\AES_ENC/us10/n769 ), .A2(\AES_ENC/us10/n768 ), .A3(\AES_ENC/us10/n767 ), .ZN(\AES_ENC/us10/n775 ) );
NOR2_X2 \AES_ENC/us10/U486  ( .A1(\AES_ENC/us10/n1056 ), .A2(\AES_ENC/us10/n1053 ), .ZN(\AES_ENC/us10/n749 ) );
NOR2_X2 \AES_ENC/us10/U483  ( .A1(\AES_ENC/us10/n749 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n752 ) );
INV_X4 \AES_ENC/us10/U482  ( .A(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n596 ));
NOR2_X2 \AES_ENC/us10/U480  ( .A1(\AES_ENC/us10/n1054 ), .A2(\AES_ENC/us10/n1053 ), .ZN(\AES_ENC/us10/n1055 ) );
OR2_X4 \AES_ENC/us10/U479  ( .A1(\AES_ENC/us10/n1094 ), .A2(\AES_ENC/us10/n1093 ), .ZN(\AES_ENC/us10/n571 ) );
AND2_X2 \AES_ENC/us10/U478  ( .A1(\AES_ENC/us10/n571 ), .A2(\AES_ENC/us10/n1095 ), .ZN(\AES_ENC/us10/n1101 ) );
NOR2_X2 \AES_ENC/us10/U477  ( .A1(\AES_ENC/us10/n1074 ), .A2(\AES_ENC/us10/n931 ), .ZN(\AES_ENC/us10/n796 ) );
NOR2_X2 \AES_ENC/us10/U474  ( .A1(\AES_ENC/us10/n796 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n797 ) );
NOR2_X2 \AES_ENC/us10/U473  ( .A1(\AES_ENC/us10/n932 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n933 ) );
NOR2_X2 \AES_ENC/us10/U472  ( .A1(\AES_ENC/us10/n929 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n935 ) );
NOR2_X2 \AES_ENC/us10/U471  ( .A1(\AES_ENC/us10/n931 ), .A2(\AES_ENC/us10/n930 ), .ZN(\AES_ENC/us10/n934 ) );
NOR3_X2 \AES_ENC/us10/U470  ( .A1(\AES_ENC/us10/n935 ), .A2(\AES_ENC/us10/n934 ), .A3(\AES_ENC/us10/n933 ), .ZN(\AES_ENC/us10/n936 ) );
NOR2_X2 \AES_ENC/us10/U469  ( .A1(\AES_ENC/us10/n624 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n1075 ) );
NOR2_X2 \AES_ENC/us10/U468  ( .A1(\AES_ENC/us10/n572 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n949 ) );
NOR2_X2 \AES_ENC/us10/U467  ( .A1(\AES_ENC/us10/n1049 ), .A2(\AES_ENC/us10/n618 ), .ZN(\AES_ENC/us10/n1051 ) );
NOR2_X2 \AES_ENC/us10/U466  ( .A1(\AES_ENC/us10/n1051 ), .A2(\AES_ENC/us10/n1050 ), .ZN(\AES_ENC/us10/n1052 ) );
NOR2_X2 \AES_ENC/us10/U465  ( .A1(\AES_ENC/us10/n1052 ), .A2(\AES_ENC/us10/n592 ), .ZN(\AES_ENC/us10/n1064 ) );
NOR2_X2 \AES_ENC/us10/U464  ( .A1(\AES_ENC/sa10 [1]), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n631 ) );
NOR2_X2 \AES_ENC/us10/U463  ( .A1(\AES_ENC/us10/n1025 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n980 ) );
NOR2_X2 \AES_ENC/us10/U462  ( .A1(\AES_ENC/us10/n1073 ), .A2(\AES_ENC/us10/n1094 ), .ZN(\AES_ENC/us10/n795 ) );
NOR2_X2 \AES_ENC/us10/U461  ( .A1(\AES_ENC/us10/n795 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n799 ) );
NOR2_X2 \AES_ENC/us10/U460  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n981 ) );
NOR2_X2 \AES_ENC/us10/U459  ( .A1(\AES_ENC/us10/n1102 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n643 ) );
NOR2_X2 \AES_ENC/us10/U458  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n621 ), .ZN(\AES_ENC/us10/n642 ) );
NOR2_X2 \AES_ENC/us10/U455  ( .A1(\AES_ENC/us10/n911 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n644 ) );
NOR4_X2 \AES_ENC/us10/U448  ( .A1(\AES_ENC/us10/n644 ), .A2(\AES_ENC/us10/n643 ), .A3(\AES_ENC/us10/n804 ), .A4(\AES_ENC/us10/n642 ), .ZN(\AES_ENC/us10/n645 ) );
NOR2_X2 \AES_ENC/us10/U447  ( .A1(\AES_ENC/us10/n1102 ), .A2(\AES_ENC/us10/n910 ), .ZN(\AES_ENC/us10/n932 ) );
NOR2_X2 \AES_ENC/us10/U442  ( .A1(\AES_ENC/us10/n1102 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n755 ) );
NOR2_X2 \AES_ENC/us10/U441  ( .A1(\AES_ENC/us10/n931 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n743 ) );
NOR2_X2 \AES_ENC/us10/U438  ( .A1(\AES_ENC/us10/n1072 ), .A2(\AES_ENC/us10/n1094 ), .ZN(\AES_ENC/us10/n930 ) );
NOR2_X2 \AES_ENC/us10/U435  ( .A1(\AES_ENC/us10/n1074 ), .A2(\AES_ENC/us10/n1025 ), .ZN(\AES_ENC/us10/n891 ) );
NOR2_X2 \AES_ENC/us10/U434  ( .A1(\AES_ENC/us10/n891 ), .A2(\AES_ENC/us10/n609 ), .ZN(\AES_ENC/us10/n894 ) );
NOR3_X2 \AES_ENC/us10/U433  ( .A1(\AES_ENC/us10/n623 ), .A2(\AES_ENC/sa10 [1]), .A3(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n683 ));
INV_X4 \AES_ENC/us10/U428  ( .A(\AES_ENC/us10/n931 ), .ZN(\AES_ENC/us10/n623 ) );
NOR2_X2 \AES_ENC/us10/U427  ( .A1(\AES_ENC/us10/n996 ), .A2(\AES_ENC/us10/n931 ), .ZN(\AES_ENC/us10/n704 ) );
NOR2_X2 \AES_ENC/us10/U421  ( .A1(\AES_ENC/us10/n931 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n685 ) );
NOR2_X2 \AES_ENC/us10/U420  ( .A1(\AES_ENC/us10/n1029 ), .A2(\AES_ENC/us10/n1025 ), .ZN(\AES_ENC/us10/n1079 ) );
NOR3_X2 \AES_ENC/us10/U419  ( .A1(\AES_ENC/us10/n589 ), .A2(\AES_ENC/us10/n1025 ), .A3(\AES_ENC/us10/n616 ), .ZN(\AES_ENC/us10/n945 ) );
NOR2_X2 \AES_ENC/us10/U418  ( .A1(\AES_ENC/us10/n626 ), .A2(\AES_ENC/us10/n611 ), .ZN(\AES_ENC/us10/n800 ) );
NOR3_X2 \AES_ENC/us10/U417  ( .A1(\AES_ENC/us10/n590 ), .A2(\AES_ENC/us10/n627 ), .A3(\AES_ENC/us10/n611 ), .ZN(\AES_ENC/us10/n798 ) );
NOR3_X2 \AES_ENC/us10/U416  ( .A1(\AES_ENC/us10/n610 ), .A2(\AES_ENC/us10/n572 ), .A3(\AES_ENC/us10/n575 ), .ZN(\AES_ENC/us10/n962 ) );
NOR3_X2 \AES_ENC/us10/U415  ( .A1(\AES_ENC/us10/n959 ), .A2(\AES_ENC/us10/n572 ), .A3(\AES_ENC/us10/n609 ), .ZN(\AES_ENC/us10/n768 ) );
NOR3_X2 \AES_ENC/us10/U414  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n572 ), .A3(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n694 ) );
NOR3_X2 \AES_ENC/us10/U413  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n572 ), .A3(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n895 ) );
NOR3_X2 \AES_ENC/us10/U410  ( .A1(\AES_ENC/us10/n1008 ), .A2(\AES_ENC/us10/n1007 ), .A3(\AES_ENC/us10/n1006 ), .ZN(\AES_ENC/us10/n1018 ) );
NOR4_X2 \AES_ENC/us10/U409  ( .A1(\AES_ENC/us10/n806 ), .A2(\AES_ENC/us10/n805 ), .A3(\AES_ENC/us10/n804 ), .A4(\AES_ENC/us10/n803 ), .ZN(\AES_ENC/us10/n807 ) );
NOR3_X2 \AES_ENC/us10/U406  ( .A1(\AES_ENC/us10/n799 ), .A2(\AES_ENC/us10/n798 ), .A3(\AES_ENC/us10/n797 ), .ZN(\AES_ENC/us10/n808 ) );
NOR4_X2 \AES_ENC/us10/U405  ( .A1(\AES_ENC/us10/n843 ), .A2(\AES_ENC/us10/n842 ), .A3(\AES_ENC/us10/n841 ), .A4(\AES_ENC/us10/n840 ), .ZN(\AES_ENC/us10/n844 ) );
NOR2_X2 \AES_ENC/us10/U404  ( .A1(\AES_ENC/us10/n669 ), .A2(\AES_ENC/us10/n668 ), .ZN(\AES_ENC/us10/n673 ) );
NOR4_X2 \AES_ENC/us10/U403  ( .A1(\AES_ENC/us10/n946 ), .A2(\AES_ENC/us10/n1046 ), .A3(\AES_ENC/us10/n671 ), .A4(\AES_ENC/us10/n670 ), .ZN(\AES_ENC/us10/n672 ) );
NOR3_X2 \AES_ENC/us10/U401  ( .A1(\AES_ENC/us10/n1101 ), .A2(\AES_ENC/us10/n1100 ), .A3(\AES_ENC/us10/n1099 ), .ZN(\AES_ENC/us10/n1109 ) );
NOR4_X2 \AES_ENC/us10/U400  ( .A1(\AES_ENC/us10/n711 ), .A2(\AES_ENC/us10/n710 ), .A3(\AES_ENC/us10/n709 ), .A4(\AES_ENC/us10/n708 ), .ZN(\AES_ENC/us10/n712 ) );
NOR4_X2 \AES_ENC/us10/U399  ( .A1(\AES_ENC/us10/n963 ), .A2(\AES_ENC/us10/n962 ), .A3(\AES_ENC/us10/n961 ), .A4(\AES_ENC/us10/n960 ), .ZN(\AES_ENC/us10/n964 ) );
NOR3_X2 \AES_ENC/us10/U398  ( .A1(\AES_ENC/us10/n743 ), .A2(\AES_ENC/us10/n742 ), .A3(\AES_ENC/us10/n741 ), .ZN(\AES_ENC/us10/n744 ) );
NOR2_X2 \AES_ENC/us10/U397  ( .A1(\AES_ENC/us10/n697 ), .A2(\AES_ENC/us10/n658 ), .ZN(\AES_ENC/us10/n659 ) );
NOR2_X2 \AES_ENC/us10/U396  ( .A1(\AES_ENC/us10/n1078 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n1033 ) );
NOR2_X2 \AES_ENC/us10/U393  ( .A1(\AES_ENC/us10/n1031 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n1032 ) );
NOR3_X2 \AES_ENC/us10/U390  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n1025 ), .A3(\AES_ENC/us10/n1074 ), .ZN(\AES_ENC/us10/n1035 ) );
NOR4_X2 \AES_ENC/us10/U389  ( .A1(\AES_ENC/us10/n1035 ), .A2(\AES_ENC/us10/n1034 ), .A3(\AES_ENC/us10/n1033 ), .A4(\AES_ENC/us10/n1032 ), .ZN(\AES_ENC/us10/n1036 ) );
NOR2_X2 \AES_ENC/us10/U388  ( .A1(\AES_ENC/us10/n598 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n885 ) );
NOR2_X2 \AES_ENC/us10/U387  ( .A1(\AES_ENC/us10/n623 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n882 ) );
NOR2_X2 \AES_ENC/us10/U386  ( .A1(\AES_ENC/us10/n1053 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n884 ) );
NOR4_X2 \AES_ENC/us10/U385  ( .A1(\AES_ENC/us10/n885 ), .A2(\AES_ENC/us10/n884 ), .A3(\AES_ENC/us10/n883 ), .A4(\AES_ENC/us10/n882 ), .ZN(\AES_ENC/us10/n886 ) );
NOR2_X2 \AES_ENC/us10/U384  ( .A1(\AES_ENC/us10/n825 ), .A2(\AES_ENC/us10/n578 ), .ZN(\AES_ENC/us10/n830 ) );
NOR2_X2 \AES_ENC/us10/U383  ( .A1(\AES_ENC/us10/n827 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n829 ) );
NOR2_X2 \AES_ENC/us10/U382  ( .A1(\AES_ENC/us10/n572 ), .A2(\AES_ENC/us10/n579 ), .ZN(\AES_ENC/us10/n828 ) );
NOR4_X2 \AES_ENC/us10/U374  ( .A1(\AES_ENC/us10/n831 ), .A2(\AES_ENC/us10/n830 ), .A3(\AES_ENC/us10/n829 ), .A4(\AES_ENC/us10/n828 ), .ZN(\AES_ENC/us10/n832 ) );
NOR2_X2 \AES_ENC/us10/U373  ( .A1(\AES_ENC/us10/n606 ), .A2(\AES_ENC/us10/n582 ), .ZN(\AES_ENC/us10/n1104 ) );
NOR2_X2 \AES_ENC/us10/U372  ( .A1(\AES_ENC/us10/n1102 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n1106 ) );
NOR2_X2 \AES_ENC/us10/U370  ( .A1(\AES_ENC/us10/n1103 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n1105 ) );
NOR4_X2 \AES_ENC/us10/U369  ( .A1(\AES_ENC/us10/n1107 ), .A2(\AES_ENC/us10/n1106 ), .A3(\AES_ENC/us10/n1105 ), .A4(\AES_ENC/us10/n1104 ), .ZN(\AES_ENC/us10/n1108 ) );
NOR3_X2 \AES_ENC/us10/U368  ( .A1(\AES_ENC/us10/n959 ), .A2(\AES_ENC/us10/n621 ), .A3(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n963 ) );
NOR2_X2 \AES_ENC/us10/U367  ( .A1(\AES_ENC/us10/n626 ), .A2(\AES_ENC/us10/n627 ), .ZN(\AES_ENC/us10/n1114 ) );
INV_X4 \AES_ENC/us10/U366  ( .A(\AES_ENC/us10/n1024 ), .ZN(\AES_ENC/us10/n606 ) );
NOR3_X2 \AES_ENC/us10/U365  ( .A1(\AES_ENC/us10/n910 ), .A2(\AES_ENC/us10/n1059 ), .A3(\AES_ENC/us10/n611 ), .ZN(\AES_ENC/us10/n1115 ) );
INV_X4 \AES_ENC/us10/U364  ( .A(\AES_ENC/us10/n1094 ), .ZN(\AES_ENC/us10/n613 ) );
NOR2_X2 \AES_ENC/us10/U363  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n931 ), .ZN(\AES_ENC/us10/n1100 ) );
INV_X4 \AES_ENC/us10/U354  ( .A(\AES_ENC/us10/n1093 ), .ZN(\AES_ENC/us10/n617 ) );
NOR2_X2 \AES_ENC/us10/U353  ( .A1(\AES_ENC/us10/n569 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n929 ) );
NOR2_X2 \AES_ENC/us10/U352  ( .A1(\AES_ENC/us10/n620 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n926 ) );
NOR2_X2 \AES_ENC/us10/U351  ( .A1(\AES_ENC/us10/n572 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n1095 ) );
NOR2_X2 \AES_ENC/us10/U350  ( .A1(\AES_ENC/us10/n609 ), .A2(\AES_ENC/us10/n627 ), .ZN(\AES_ENC/us10/n1010 ) );
NOR2_X2 \AES_ENC/us10/U349  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n1103 ) );
NOR2_X2 \AES_ENC/us10/U348  ( .A1(\AES_ENC/us10/n622 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n1059 ) );
NOR2_X2 \AES_ENC/us10/U347  ( .A1(\AES_ENC/sa10 [1]), .A2(\AES_ENC/us10/n1120 ), .ZN(\AES_ENC/us10/n1022 ) );
NOR2_X2 \AES_ENC/us10/U346  ( .A1(\AES_ENC/us10/n619 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n911 ) );
NOR2_X2 \AES_ENC/us10/U345  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/us10/n1025 ), .ZN(\AES_ENC/us10/n826 ) );
NOR2_X2 \AES_ENC/us10/U338  ( .A1(\AES_ENC/us10/n626 ), .A2(\AES_ENC/us10/n607 ), .ZN(\AES_ENC/us10/n1072 ) );
NOR2_X2 \AES_ENC/us10/U335  ( .A1(\AES_ENC/us10/n627 ), .A2(\AES_ENC/us10/n616 ), .ZN(\AES_ENC/us10/n956 ) );
NOR2_X2 \AES_ENC/us10/U329  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/us10/n624 ), .ZN(\AES_ENC/us10/n1121 ) );
NOR2_X2 \AES_ENC/us10/U328  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/us10/n624 ), .ZN(\AES_ENC/us10/n1058 ) );
NOR2_X2 \AES_ENC/us10/U327  ( .A1(\AES_ENC/us10/n625 ), .A2(\AES_ENC/us10/n611 ), .ZN(\AES_ENC/us10/n1073 ) );
NOR2_X2 \AES_ENC/us10/U325  ( .A1(\AES_ENC/sa10 [1]), .A2(\AES_ENC/us10/n1025 ), .ZN(\AES_ENC/us10/n1054 ) );
NOR2_X2 \AES_ENC/us10/U324  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/us10/n931 ), .ZN(\AES_ENC/us10/n1029 ) );
NOR2_X2 \AES_ENC/us10/U319  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n1056 ) );
NOR2_X2 \AES_ENC/us10/U318  ( .A1(\AES_ENC/us10/n614 ), .A2(\AES_ENC/us10/n626 ), .ZN(\AES_ENC/us10/n1050 ) );
NOR2_X2 \AES_ENC/us10/U317  ( .A1(\AES_ENC/us10/n1121 ), .A2(\AES_ENC/us10/n1025 ), .ZN(\AES_ENC/us10/n1120 ) );
NOR2_X2 \AES_ENC/us10/U316  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/us10/n572 ), .ZN(\AES_ENC/us10/n1074 ) );
NOR2_X2 \AES_ENC/us10/U315  ( .A1(\AES_ENC/us10/n1058 ), .A2(\AES_ENC/us10/n1054 ), .ZN(\AES_ENC/us10/n878 ) );
NOR2_X2 \AES_ENC/us10/U314  ( .A1(\AES_ENC/us10/n878 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n879 ) );
NOR2_X2 \AES_ENC/us10/U312  ( .A1(\AES_ENC/us10/n880 ), .A2(\AES_ENC/us10/n879 ), .ZN(\AES_ENC/us10/n887 ) );
NOR2_X2 \AES_ENC/us10/U311  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n588 ), .ZN(\AES_ENC/us10/n957 ) );
NOR2_X2 \AES_ENC/us10/U310  ( .A1(\AES_ENC/us10/n958 ), .A2(\AES_ENC/us10/n957 ), .ZN(\AES_ENC/us10/n965 ) );
NOR3_X2 \AES_ENC/us10/U309  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n1091 ), .A3(\AES_ENC/us10/n1022 ), .ZN(\AES_ENC/us10/n720 ) );
NOR3_X2 \AES_ENC/us10/U303  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n1054 ), .A3(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n719 ) );
NOR2_X2 \AES_ENC/us10/U302  ( .A1(\AES_ENC/us10/n720 ), .A2(\AES_ENC/us10/n719 ), .ZN(\AES_ENC/us10/n726 ) );
NOR2_X2 \AES_ENC/us10/U300  ( .A1(\AES_ENC/us10/n614 ), .A2(\AES_ENC/us10/n591 ), .ZN(\AES_ENC/us10/n865 ) );
NOR2_X2 \AES_ENC/us10/U299  ( .A1(\AES_ENC/us10/n1059 ), .A2(\AES_ENC/us10/n1058 ), .ZN(\AES_ENC/us10/n1060 ) );
NOR2_X2 \AES_ENC/us10/U298  ( .A1(\AES_ENC/us10/n1095 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n668 ) );
NOR2_X2 \AES_ENC/us10/U297  ( .A1(\AES_ENC/us10/n911 ), .A2(\AES_ENC/us10/n910 ), .ZN(\AES_ENC/us10/n912 ) );
NOR2_X2 \AES_ENC/us10/U296  ( .A1(\AES_ENC/us10/n912 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n916 ) );
NOR2_X2 \AES_ENC/us10/U295  ( .A1(\AES_ENC/us10/n826 ), .A2(\AES_ENC/us10/n573 ), .ZN(\AES_ENC/us10/n750 ) );
NOR2_X2 \AES_ENC/us10/U294  ( .A1(\AES_ENC/us10/n750 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n751 ) );
NOR2_X2 \AES_ENC/us10/U293  ( .A1(\AES_ENC/us10/n907 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n908 ) );
NOR2_X2 \AES_ENC/us10/U292  ( .A1(\AES_ENC/us10/n990 ), .A2(\AES_ENC/us10/n926 ), .ZN(\AES_ENC/us10/n780 ) );
NOR2_X2 \AES_ENC/us10/U291  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n584 ), .ZN(\AES_ENC/us10/n838 ) );
NOR2_X2 \AES_ENC/us10/U290  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n602 ), .ZN(\AES_ENC/us10/n837 ) );
NOR2_X2 \AES_ENC/us10/U284  ( .A1(\AES_ENC/us10/n838 ), .A2(\AES_ENC/us10/n837 ), .ZN(\AES_ENC/us10/n845 ) );
NOR2_X2 \AES_ENC/us10/U283  ( .A1(\AES_ENC/us10/n1022 ), .A2(\AES_ENC/us10/n1058 ), .ZN(\AES_ENC/us10/n740 ) );
NOR2_X2 \AES_ENC/us10/U282  ( .A1(\AES_ENC/us10/n740 ), .A2(\AES_ENC/us10/n616 ), .ZN(\AES_ENC/us10/n742 ) );
NOR2_X2 \AES_ENC/us10/U281  ( .A1(\AES_ENC/us10/n1098 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n1099 ) );
NOR2_X2 \AES_ENC/us10/U280  ( .A1(\AES_ENC/us10/n1120 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n993 ) );
NOR2_X2 \AES_ENC/us10/U279  ( .A1(\AES_ENC/us10/n993 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n994 ) );
NOR2_X2 \AES_ENC/us10/U273  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n620 ), .ZN(\AES_ENC/us10/n1026 ) );
NOR2_X2 \AES_ENC/us10/U272  ( .A1(\AES_ENC/us10/n573 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n1027 ) );
NOR2_X2 \AES_ENC/us10/U271  ( .A1(\AES_ENC/us10/n1027 ), .A2(\AES_ENC/us10/n1026 ), .ZN(\AES_ENC/us10/n1028 ) );
NOR2_X2 \AES_ENC/us10/U270  ( .A1(\AES_ENC/us10/n1029 ), .A2(\AES_ENC/us10/n1028 ), .ZN(\AES_ENC/us10/n1034 ) );
NOR4_X2 \AES_ENC/us10/U269  ( .A1(\AES_ENC/us10/n757 ), .A2(\AES_ENC/us10/n756 ), .A3(\AES_ENC/us10/n755 ), .A4(\AES_ENC/us10/n754 ), .ZN(\AES_ENC/us10/n758 ) );
NOR2_X2 \AES_ENC/us10/U268  ( .A1(\AES_ENC/us10/n752 ), .A2(\AES_ENC/us10/n751 ), .ZN(\AES_ENC/us10/n759 ) );
NOR2_X2 \AES_ENC/us10/U267  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n1071 ), .ZN(\AES_ENC/us10/n669 ) );
NOR2_X2 \AES_ENC/us10/U263  ( .A1(\AES_ENC/us10/n1056 ), .A2(\AES_ENC/us10/n990 ), .ZN(\AES_ENC/us10/n991 ) );
NOR2_X2 \AES_ENC/us10/U262  ( .A1(\AES_ENC/us10/n991 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n995 ) );
NOR2_X2 \AES_ENC/us10/U258  ( .A1(\AES_ENC/us10/n607 ), .A2(\AES_ENC/us10/n590 ), .ZN(\AES_ENC/us10/n1008 ) );
NOR2_X2 \AES_ENC/us10/U255  ( .A1(\AES_ENC/us10/n839 ), .A2(\AES_ENC/us10/n582 ), .ZN(\AES_ENC/us10/n693 ) );
NOR2_X2 \AES_ENC/us10/U254  ( .A1(\AES_ENC/us10/n606 ), .A2(\AES_ENC/us10/n906 ), .ZN(\AES_ENC/us10/n741 ) );
NOR2_X2 \AES_ENC/us10/U253  ( .A1(\AES_ENC/us10/n1054 ), .A2(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n763 ) );
NOR2_X2 \AES_ENC/us10/U252  ( .A1(\AES_ENC/us10/n763 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n769 ) );
NOR2_X2 \AES_ENC/us10/U251  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n577 ), .ZN(\AES_ENC/us10/n1007 ) );
NOR2_X2 \AES_ENC/us10/U250  ( .A1(\AES_ENC/us10/n609 ), .A2(\AES_ENC/us10/n580 ), .ZN(\AES_ENC/us10/n1123 ) );
NOR2_X2 \AES_ENC/us10/U243  ( .A1(\AES_ENC/us10/n609 ), .A2(\AES_ENC/us10/n590 ), .ZN(\AES_ENC/us10/n710 ) );
INV_X4 \AES_ENC/us10/U242  ( .A(\AES_ENC/us10/n1029 ), .ZN(\AES_ENC/us10/n582 ) );
NOR2_X2 \AES_ENC/us10/U241  ( .A1(\AES_ENC/us10/n616 ), .A2(\AES_ENC/us10/n597 ), .ZN(\AES_ENC/us10/n883 ) );
NOR2_X2 \AES_ENC/us10/U240  ( .A1(\AES_ENC/us10/n593 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n1125 ) );
NOR2_X2 \AES_ENC/us10/U239  ( .A1(\AES_ENC/us10/n990 ), .A2(\AES_ENC/us10/n929 ), .ZN(\AES_ENC/us10/n892 ) );
NOR2_X2 \AES_ENC/us10/U238  ( .A1(\AES_ENC/us10/n892 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n893 ) );
NOR2_X2 \AES_ENC/us10/U237  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n602 ), .ZN(\AES_ENC/us10/n950 ) );
NOR2_X2 \AES_ENC/us10/U236  ( .A1(\AES_ENC/us10/n1079 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n1082 ) );
NOR2_X2 \AES_ENC/us10/U235  ( .A1(\AES_ENC/us10/n910 ), .A2(\AES_ENC/us10/n1056 ), .ZN(\AES_ENC/us10/n941 ) );
NOR2_X2 \AES_ENC/us10/U234  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n1077 ), .ZN(\AES_ENC/us10/n841 ) );
NOR2_X2 \AES_ENC/us10/U229  ( .A1(\AES_ENC/us10/n623 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n630 ) );
NOR2_X2 \AES_ENC/us10/U228  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n602 ), .ZN(\AES_ENC/us10/n806 ) );
NOR2_X2 \AES_ENC/us10/U227  ( .A1(\AES_ENC/us10/n623 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n948 ) );
NOR2_X2 \AES_ENC/us10/U226  ( .A1(\AES_ENC/us10/n606 ), .A2(\AES_ENC/us10/n589 ), .ZN(\AES_ENC/us10/n997 ) );
NOR2_X2 \AES_ENC/us10/U225  ( .A1(\AES_ENC/us10/n1121 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n1122 ) );
NOR2_X2 \AES_ENC/us10/U223  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n1023 ), .ZN(\AES_ENC/us10/n756 ) );
NOR2_X2 \AES_ENC/us10/U222  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n602 ), .ZN(\AES_ENC/us10/n870 ) );
NOR2_X2 \AES_ENC/us10/U221  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n569 ), .ZN(\AES_ENC/us10/n947 ) );
NOR2_X2 \AES_ENC/us10/U217  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n1077 ), .ZN(\AES_ENC/us10/n1084 ) );
NOR2_X2 \AES_ENC/us10/U213  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n855 ), .ZN(\AES_ENC/us10/n709 ) );
NOR2_X2 \AES_ENC/us10/U212  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n589 ), .ZN(\AES_ENC/us10/n868 ) );
NOR2_X2 \AES_ENC/us10/U211  ( .A1(\AES_ENC/us10/n1120 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n1124 ) );
NOR2_X2 \AES_ENC/us10/U210  ( .A1(\AES_ENC/us10/n1120 ), .A2(\AES_ENC/us10/n839 ), .ZN(\AES_ENC/us10/n842 ) );
NOR2_X2 \AES_ENC/us10/U209  ( .A1(\AES_ENC/us10/n1120 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n696 ) );
NOR2_X2 \AES_ENC/us10/U208  ( .A1(\AES_ENC/us10/n1074 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n1076 ) );
NOR2_X2 \AES_ENC/us10/U207  ( .A1(\AES_ENC/us10/n1074 ), .A2(\AES_ENC/us10/n620 ), .ZN(\AES_ENC/us10/n781 ) );
NOR3_X2 \AES_ENC/us10/U201  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n1056 ), .A3(\AES_ENC/us10/n990 ), .ZN(\AES_ENC/us10/n979 ) );
NOR3_X2 \AES_ENC/us10/U200  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n1058 ), .A3(\AES_ENC/us10/n1059 ), .ZN(\AES_ENC/us10/n854 ) );
NOR2_X2 \AES_ENC/us10/U199  ( .A1(\AES_ENC/us10/n996 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n869 ) );
NOR2_X2 \AES_ENC/us10/U198  ( .A1(\AES_ENC/us10/n1056 ), .A2(\AES_ENC/us10/n1074 ), .ZN(\AES_ENC/us10/n1057 ) );
NOR3_X2 \AES_ENC/us10/U197  ( .A1(\AES_ENC/us10/n607 ), .A2(\AES_ENC/us10/n1120 ), .A3(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n978 ) );
NOR2_X2 \AES_ENC/us10/U196  ( .A1(\AES_ENC/us10/n996 ), .A2(\AES_ENC/us10/n911 ), .ZN(\AES_ENC/us10/n1116 ) );
NOR2_X2 \AES_ENC/us10/U195  ( .A1(\AES_ENC/us10/n1074 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n754 ) );
NOR2_X2 \AES_ENC/us10/U194  ( .A1(\AES_ENC/us10/n926 ), .A2(\AES_ENC/us10/n1103 ), .ZN(\AES_ENC/us10/n977 ) );
NOR2_X2 \AES_ENC/us10/U187  ( .A1(\AES_ENC/us10/n839 ), .A2(\AES_ENC/us10/n824 ), .ZN(\AES_ENC/us10/n1092 ) );
NOR2_X2 \AES_ENC/us10/U186  ( .A1(\AES_ENC/us10/n573 ), .A2(\AES_ENC/us10/n1074 ), .ZN(\AES_ENC/us10/n684 ) );
NOR2_X2 \AES_ENC/us10/U185  ( .A1(\AES_ENC/us10/n826 ), .A2(\AES_ENC/us10/n1059 ), .ZN(\AES_ENC/us10/n907 ) );
NOR3_X2 \AES_ENC/us10/U184  ( .A1(\AES_ENC/us10/n625 ), .A2(\AES_ENC/us10/n1115 ), .A3(\AES_ENC/us10/n585 ), .ZN(\AES_ENC/us10/n831 ) );
NOR3_X2 \AES_ENC/us10/U183  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n1056 ), .A3(\AES_ENC/us10/n990 ), .ZN(\AES_ENC/us10/n896 ) );
NOR3_X2 \AES_ENC/us10/U182  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n573 ), .A3(\AES_ENC/us10/n1013 ), .ZN(\AES_ENC/us10/n670 ) );
NOR3_X2 \AES_ENC/us10/U181  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n1091 ), .A3(\AES_ENC/us10/n1022 ), .ZN(\AES_ENC/us10/n843 ) );
NOR2_X2 \AES_ENC/us10/U180  ( .A1(\AES_ENC/us10/n1029 ), .A2(\AES_ENC/us10/n1095 ), .ZN(\AES_ENC/us10/n735 ) );
NOR2_X2 \AES_ENC/us10/U174  ( .A1(\AES_ENC/us10/n1100 ), .A2(\AES_ENC/us10/n854 ), .ZN(\AES_ENC/us10/n860 ) );
NOR4_X2 \AES_ENC/us10/U173  ( .A1(\AES_ENC/us10/n1125 ), .A2(\AES_ENC/us10/n1124 ), .A3(\AES_ENC/us10/n1123 ), .A4(\AES_ENC/us10/n1122 ), .ZN(\AES_ENC/us10/n1126 ) );
NOR4_X2 \AES_ENC/us10/U172  ( .A1(\AES_ENC/us10/n1084 ), .A2(\AES_ENC/us10/n1083 ), .A3(\AES_ENC/us10/n1082 ), .A4(\AES_ENC/us10/n1081 ), .ZN(\AES_ENC/us10/n1085 ) );
NOR2_X2 \AES_ENC/us10/U171  ( .A1(\AES_ENC/us10/n1076 ), .A2(\AES_ENC/us10/n1075 ), .ZN(\AES_ENC/us10/n1086 ) );
NAND3_X2 \AES_ENC/us10/U170  ( .A1(\AES_ENC/us10/n569 ), .A2(\AES_ENC/us10/n582 ), .A3(\AES_ENC/us10/n681 ), .ZN(\AES_ENC/us10/n691 ) );
NOR2_X2 \AES_ENC/us10/U169  ( .A1(\AES_ENC/us10/n683 ), .A2(\AES_ENC/us10/n682 ), .ZN(\AES_ENC/us10/n690 ) );
NOR3_X2 \AES_ENC/us10/U168  ( .A1(\AES_ENC/us10/n695 ), .A2(\AES_ENC/us10/n694 ), .A3(\AES_ENC/us10/n693 ), .ZN(\AES_ENC/us10/n700 ) );
NOR4_X2 \AES_ENC/us10/U162  ( .A1(\AES_ENC/us10/n983 ), .A2(\AES_ENC/us10/n698 ), .A3(\AES_ENC/us10/n697 ), .A4(\AES_ENC/us10/n696 ), .ZN(\AES_ENC/us10/n699 ) );
NOR2_X2 \AES_ENC/us10/U161  ( .A1(\AES_ENC/us10/n946 ), .A2(\AES_ENC/us10/n945 ), .ZN(\AES_ENC/us10/n952 ) );
NOR4_X2 \AES_ENC/us10/U160  ( .A1(\AES_ENC/us10/n950 ), .A2(\AES_ENC/us10/n949 ), .A3(\AES_ENC/us10/n948 ), .A4(\AES_ENC/us10/n947 ), .ZN(\AES_ENC/us10/n951 ) );
NOR4_X2 \AES_ENC/us10/U159  ( .A1(\AES_ENC/us10/n983 ), .A2(\AES_ENC/us10/n982 ), .A3(\AES_ENC/us10/n981 ), .A4(\AES_ENC/us10/n980 ), .ZN(\AES_ENC/us10/n984 ) );
NOR2_X2 \AES_ENC/us10/U158  ( .A1(\AES_ENC/us10/n979 ), .A2(\AES_ENC/us10/n978 ), .ZN(\AES_ENC/us10/n985 ) );
NOR4_X2 \AES_ENC/us10/U157  ( .A1(\AES_ENC/us10/n896 ), .A2(\AES_ENC/us10/n895 ), .A3(\AES_ENC/us10/n894 ), .A4(\AES_ENC/us10/n893 ), .ZN(\AES_ENC/us10/n897 ) );
NOR2_X2 \AES_ENC/us10/U156  ( .A1(\AES_ENC/us10/n866 ), .A2(\AES_ENC/us10/n865 ), .ZN(\AES_ENC/us10/n872 ) );
NOR4_X2 \AES_ENC/us10/U155  ( .A1(\AES_ENC/us10/n870 ), .A2(\AES_ENC/us10/n869 ), .A3(\AES_ENC/us10/n868 ), .A4(\AES_ENC/us10/n867 ), .ZN(\AES_ENC/us10/n871 ) );
NOR3_X2 \AES_ENC/us10/U154  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n1054 ), .A3(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n961 ) );
NOR3_X2 \AES_ENC/us10/U153  ( .A1(\AES_ENC/us10/n620 ), .A2(\AES_ENC/us10/n1074 ), .A3(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n671 ) );
NOR2_X2 \AES_ENC/us10/U152  ( .A1(\AES_ENC/us10/n1057 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n1062 ) );
NOR2_X2 \AES_ENC/us10/U143  ( .A1(\AES_ENC/us10/n1055 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n1063 ) );
NOR2_X2 \AES_ENC/us10/U142  ( .A1(\AES_ENC/us10/n1060 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n1061 ) );
NOR4_X2 \AES_ENC/us10/U141  ( .A1(\AES_ENC/us10/n1064 ), .A2(\AES_ENC/us10/n1063 ), .A3(\AES_ENC/us10/n1062 ), .A4(\AES_ENC/us10/n1061 ), .ZN(\AES_ENC/us10/n1065 ) );
NOR3_X2 \AES_ENC/us10/U140  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n1120 ), .A3(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n918 ) );
NOR3_X2 \AES_ENC/us10/U132  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n573 ), .A3(\AES_ENC/us10/n1013 ), .ZN(\AES_ENC/us10/n917 ) );
NOR2_X2 \AES_ENC/us10/U131  ( .A1(\AES_ENC/us10/n914 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n915 ) );
NOR4_X2 \AES_ENC/us10/U130  ( .A1(\AES_ENC/us10/n918 ), .A2(\AES_ENC/us10/n917 ), .A3(\AES_ENC/us10/n916 ), .A4(\AES_ENC/us10/n915 ), .ZN(\AES_ENC/us10/n919 ) );
NOR2_X2 \AES_ENC/us10/U129  ( .A1(\AES_ENC/us10/n616 ), .A2(\AES_ENC/us10/n580 ), .ZN(\AES_ENC/us10/n771 ) );
NOR2_X2 \AES_ENC/us10/U128  ( .A1(\AES_ENC/us10/n1103 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n772 ) );
NOR2_X2 \AES_ENC/us10/U127  ( .A1(\AES_ENC/us10/n610 ), .A2(\AES_ENC/us10/n599 ), .ZN(\AES_ENC/us10/n773 ) );
NOR4_X2 \AES_ENC/us10/U126  ( .A1(\AES_ENC/us10/n773 ), .A2(\AES_ENC/us10/n772 ), .A3(\AES_ENC/us10/n771 ), .A4(\AES_ENC/us10/n770 ), .ZN(\AES_ENC/us10/n774 ) );
NOR2_X2 \AES_ENC/us10/U121  ( .A1(\AES_ENC/us10/n735 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n687 ) );
NOR2_X2 \AES_ENC/us10/U120  ( .A1(\AES_ENC/us10/n684 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n688 ) );
NOR2_X2 \AES_ENC/us10/U119  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n600 ), .ZN(\AES_ENC/us10/n686 ) );
NOR4_X2 \AES_ENC/us10/U118  ( .A1(\AES_ENC/us10/n688 ), .A2(\AES_ENC/us10/n687 ), .A3(\AES_ENC/us10/n686 ), .A4(\AES_ENC/us10/n685 ), .ZN(\AES_ENC/us10/n689 ) );
NOR2_X2 \AES_ENC/us10/U117  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n595 ), .ZN(\AES_ENC/us10/n858 ) );
NOR2_X2 \AES_ENC/us10/U116  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n855 ), .ZN(\AES_ENC/us10/n857 ) );
NOR2_X2 \AES_ENC/us10/U115  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n587 ), .ZN(\AES_ENC/us10/n856 ) );
NOR4_X2 \AES_ENC/us10/U106  ( .A1(\AES_ENC/us10/n858 ), .A2(\AES_ENC/us10/n857 ), .A3(\AES_ENC/us10/n856 ), .A4(\AES_ENC/us10/n958 ), .ZN(\AES_ENC/us10/n859 ) );
NOR2_X2 \AES_ENC/us10/U105  ( .A1(\AES_ENC/us10/n780 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n784 ) );
NOR2_X2 \AES_ENC/us10/U104  ( .A1(\AES_ENC/us10/n1117 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n782 ) );
NOR2_X2 \AES_ENC/us10/U103  ( .A1(\AES_ENC/us10/n781 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n783 ) );
NOR4_X2 \AES_ENC/us10/U102  ( .A1(\AES_ENC/us10/n880 ), .A2(\AES_ENC/us10/n784 ), .A3(\AES_ENC/us10/n783 ), .A4(\AES_ENC/us10/n782 ), .ZN(\AES_ENC/us10/n785 ) );
NOR2_X2 \AES_ENC/us10/U101  ( .A1(\AES_ENC/us10/n583 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n814 ) );
NOR2_X2 \AES_ENC/us10/U100  ( .A1(\AES_ENC/us10/n907 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n813 ) );
NOR3_X2 \AES_ENC/us10/U95  ( .A1(\AES_ENC/us10/n606 ), .A2(\AES_ENC/us10/n1058 ), .A3(\AES_ENC/us10/n1059 ), .ZN(\AES_ENC/us10/n815 ) );
NOR4_X2 \AES_ENC/us10/U94  ( .A1(\AES_ENC/us10/n815 ), .A2(\AES_ENC/us10/n814 ), .A3(\AES_ENC/us10/n813 ), .A4(\AES_ENC/us10/n812 ), .ZN(\AES_ENC/us10/n816 ) );
NOR2_X2 \AES_ENC/us10/U93  ( .A1(\AES_ENC/us10/n617 ), .A2(\AES_ENC/us10/n569 ), .ZN(\AES_ENC/us10/n721 ) );
NOR2_X2 \AES_ENC/us10/U92  ( .A1(\AES_ENC/us10/n1031 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n723 ) );
NOR2_X2 \AES_ENC/us10/U91  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n1096 ), .ZN(\AES_ENC/us10/n722 ) );
NOR4_X2 \AES_ENC/us10/U90  ( .A1(\AES_ENC/us10/n724 ), .A2(\AES_ENC/us10/n723 ), .A3(\AES_ENC/us10/n722 ), .A4(\AES_ENC/us10/n721 ), .ZN(\AES_ENC/us10/n725 ) );
NOR2_X2 \AES_ENC/us10/U89  ( .A1(\AES_ENC/us10/n911 ), .A2(\AES_ENC/us10/n990 ), .ZN(\AES_ENC/us10/n1009 ) );
NOR2_X2 \AES_ENC/us10/U88  ( .A1(\AES_ENC/us10/n1013 ), .A2(\AES_ENC/us10/n573 ), .ZN(\AES_ENC/us10/n1014 ) );
NOR2_X2 \AES_ENC/us10/U87  ( .A1(\AES_ENC/us10/n1014 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n1015 ) );
NOR4_X2 \AES_ENC/us10/U86  ( .A1(\AES_ENC/us10/n1016 ), .A2(\AES_ENC/us10/n1015 ), .A3(\AES_ENC/us10/n1119 ), .A4(\AES_ENC/us10/n1046 ), .ZN(\AES_ENC/us10/n1017 ) );
NOR2_X2 \AES_ENC/us10/U81  ( .A1(\AES_ENC/us10/n996 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n998 ) );
NOR2_X2 \AES_ENC/us10/U80  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n577 ), .ZN(\AES_ENC/us10/n1000 ) );
NOR2_X2 \AES_ENC/us10/U79  ( .A1(\AES_ENC/us10/n616 ), .A2(\AES_ENC/us10/n1096 ), .ZN(\AES_ENC/us10/n999 ) );
NOR4_X2 \AES_ENC/us10/U78  ( .A1(\AES_ENC/us10/n1000 ), .A2(\AES_ENC/us10/n999 ), .A3(\AES_ENC/us10/n998 ), .A4(\AES_ENC/us10/n997 ), .ZN(\AES_ENC/us10/n1001 ) );
NOR2_X2 \AES_ENC/us10/U74  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n1096 ), .ZN(\AES_ENC/us10/n697 ) );
NOR2_X2 \AES_ENC/us10/U73  ( .A1(\AES_ENC/us10/n620 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n958 ) );
NOR2_X2 \AES_ENC/us10/U72  ( .A1(\AES_ENC/us10/n911 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n983 ) );
NOR2_X2 \AES_ENC/us10/U71  ( .A1(\AES_ENC/us10/n1054 ), .A2(\AES_ENC/us10/n1103 ), .ZN(\AES_ENC/us10/n1031 ) );
INV_X4 \AES_ENC/us10/U65  ( .A(\AES_ENC/us10/n1050 ), .ZN(\AES_ENC/us10/n612 ) );
INV_X4 \AES_ENC/us10/U64  ( .A(\AES_ENC/us10/n1072 ), .ZN(\AES_ENC/us10/n605 ) );
INV_X4 \AES_ENC/us10/U63  ( .A(\AES_ENC/us10/n1073 ), .ZN(\AES_ENC/us10/n604 ) );
NOR2_X2 \AES_ENC/us10/U62  ( .A1(\AES_ENC/us10/n582 ), .A2(\AES_ENC/us10/n613 ), .ZN(\AES_ENC/us10/n880 ) );
NOR3_X2 \AES_ENC/us10/U61  ( .A1(\AES_ENC/us10/n826 ), .A2(\AES_ENC/us10/n1121 ), .A3(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n946 ) );
INV_X4 \AES_ENC/us10/U59  ( .A(\AES_ENC/us10/n1010 ), .ZN(\AES_ENC/us10/n608 ) );
NOR3_X2 \AES_ENC/us10/U58  ( .A1(\AES_ENC/us10/n573 ), .A2(\AES_ENC/us10/n1029 ), .A3(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n1119 ) );
INV_X4 \AES_ENC/us10/U57  ( .A(\AES_ENC/us10/n956 ), .ZN(\AES_ENC/us10/n615 ) );
NOR2_X2 \AES_ENC/us10/U50  ( .A1(\AES_ENC/us10/n623 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n1013 ) );
NOR2_X2 \AES_ENC/us10/U49  ( .A1(\AES_ENC/us10/n620 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n910 ) );
NOR2_X2 \AES_ENC/us10/U48  ( .A1(\AES_ENC/us10/n569 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n1091 ) );
NOR2_X2 \AES_ENC/us10/U47  ( .A1(\AES_ENC/us10/n622 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n990 ) );
NOR2_X2 \AES_ENC/us10/U46  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/us10/n1121 ), .ZN(\AES_ENC/us10/n996 ) );
NOR2_X2 \AES_ENC/us10/U45  ( .A1(\AES_ENC/us10/n610 ), .A2(\AES_ENC/us10/n600 ), .ZN(\AES_ENC/us10/n628 ) );
NOR2_X2 \AES_ENC/us10/U44  ( .A1(\AES_ENC/us10/n576 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n866 ) );
NOR2_X2 \AES_ENC/us10/U43  ( .A1(\AES_ENC/us10/n603 ), .A2(\AES_ENC/us10/n610 ), .ZN(\AES_ENC/us10/n1006 ) );
NOR2_X2 \AES_ENC/us10/U42  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n1117 ), .ZN(\AES_ENC/us10/n1118 ) );
NOR2_X2 \AES_ENC/us10/U41  ( .A1(\AES_ENC/us10/n1119 ), .A2(\AES_ENC/us10/n1118 ), .ZN(\AES_ENC/us10/n1127 ) );
NOR2_X2 \AES_ENC/us10/U36  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n594 ), .ZN(\AES_ENC/us10/n629 ) );
NOR2_X2 \AES_ENC/us10/U35  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n906 ), .ZN(\AES_ENC/us10/n909 ) );
NOR2_X2 \AES_ENC/us10/U34  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n597 ), .ZN(\AES_ENC/us10/n658 ) );
NOR2_X2 \AES_ENC/us10/U33  ( .A1(\AES_ENC/us10/n1116 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n695 ) );
NOR2_X2 \AES_ENC/us10/U32  ( .A1(\AES_ENC/us10/n1078 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n1083 ) );
NOR2_X2 \AES_ENC/us10/U31  ( .A1(\AES_ENC/us10/n941 ), .A2(\AES_ENC/us10/n608 ), .ZN(\AES_ENC/us10/n724 ) );
NOR2_X2 \AES_ENC/us10/U30  ( .A1(\AES_ENC/us10/n598 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n1107 ) );
NOR2_X2 \AES_ENC/us10/U29  ( .A1(\AES_ENC/us10/n576 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n840 ) );
NOR2_X2 \AES_ENC/us10/U24  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n593 ), .ZN(\AES_ENC/us10/n633 ) );
NOR2_X2 \AES_ENC/us10/U23  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n1080 ), .ZN(\AES_ENC/us10/n1081 ) );
NOR2_X2 \AES_ENC/us10/U21  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n1045 ), .ZN(\AES_ENC/us10/n812 ) );
NOR2_X2 \AES_ENC/us10/U20  ( .A1(\AES_ENC/us10/n1009 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n960 ) );
NOR2_X2 \AES_ENC/us10/U19  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n601 ), .ZN(\AES_ENC/us10/n982 ) );
NOR2_X2 \AES_ENC/us10/U18  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n594 ), .ZN(\AES_ENC/us10/n757 ) );
NOR2_X2 \AES_ENC/us10/U17  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n590 ), .ZN(\AES_ENC/us10/n698 ) );
NOR2_X2 \AES_ENC/us10/U16  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n619 ), .ZN(\AES_ENC/us10/n708 ) );
NOR2_X2 \AES_ENC/us10/U15  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n582 ), .ZN(\AES_ENC/us10/n770 ) );
NOR2_X2 \AES_ENC/us10/U10  ( .A1(\AES_ENC/us10/n619 ), .A2(\AES_ENC/us10/n604 ), .ZN(\AES_ENC/us10/n803 ) );
NOR2_X2 \AES_ENC/us10/U9  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n881 ), .ZN(\AES_ENC/us10/n711 ) );
NOR2_X2 \AES_ENC/us10/U8  ( .A1(\AES_ENC/us10/n615 ), .A2(\AES_ENC/us10/n582 ), .ZN(\AES_ENC/us10/n867 ) );
NOR2_X2 \AES_ENC/us10/U7  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n599 ), .ZN(\AES_ENC/us10/n804 ) );
NOR2_X2 \AES_ENC/us10/U6  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n620 ), .ZN(\AES_ENC/us10/n1046 ) );
OR2_X4 \AES_ENC/us10/U5  ( .A1(\AES_ENC/us10/n624 ), .A2(\AES_ENC/sa10 [1]),.ZN(\AES_ENC/us10/n570 ) );
OR2_X4 \AES_ENC/us10/U4  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/sa10 [4]),.ZN(\AES_ENC/us10/n569 ) );
NAND2_X2 \AES_ENC/us10/U514  ( .A1(\AES_ENC/us10/n1121 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n1030 ) );
AND2_X2 \AES_ENC/us10/U513  ( .A1(\AES_ENC/us10/n597 ), .A2(\AES_ENC/us10/n1030 ), .ZN(\AES_ENC/us10/n1049 ) );
NAND2_X2 \AES_ENC/us10/U511  ( .A1(\AES_ENC/us10/n1049 ), .A2(\AES_ENC/us10/n794 ), .ZN(\AES_ENC/us10/n637 ) );
AND2_X2 \AES_ENC/us10/U493  ( .A1(\AES_ENC/us10/n779 ), .A2(\AES_ENC/us10/n996 ), .ZN(\AES_ENC/us10/n632 ) );
NAND4_X2 \AES_ENC/us10/U485  ( .A1(\AES_ENC/us10/n637 ), .A2(\AES_ENC/us10/n636 ), .A3(\AES_ENC/us10/n635 ), .A4(\AES_ENC/us10/n634 ), .ZN(\AES_ENC/us10/n638 ) );
NAND2_X2 \AES_ENC/us10/U484  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n638 ), .ZN(\AES_ENC/us10/n679 ) );
NAND2_X2 \AES_ENC/us10/U481  ( .A1(\AES_ENC/us10/n1094 ), .A2(\AES_ENC/us10/n591 ), .ZN(\AES_ENC/us10/n648 ) );
NAND2_X2 \AES_ENC/us10/U476  ( .A1(\AES_ENC/us10/n601 ), .A2(\AES_ENC/us10/n590 ), .ZN(\AES_ENC/us10/n762 ) );
NAND2_X2 \AES_ENC/us10/U475  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n762 ), .ZN(\AES_ENC/us10/n647 ) );
NAND4_X2 \AES_ENC/us10/U457  ( .A1(\AES_ENC/us10/n648 ), .A2(\AES_ENC/us10/n647 ), .A3(\AES_ENC/us10/n646 ), .A4(\AES_ENC/us10/n645 ), .ZN(\AES_ENC/us10/n649 ) );
NAND2_X2 \AES_ENC/us10/U456  ( .A1(\AES_ENC/sa10 [0]), .A2(\AES_ENC/us10/n649 ), .ZN(\AES_ENC/us10/n665 ) );
NAND2_X2 \AES_ENC/us10/U454  ( .A1(\AES_ENC/us10/n596 ), .A2(\AES_ENC/us10/n623 ), .ZN(\AES_ENC/us10/n855 ) );
NAND2_X2 \AES_ENC/us10/U453  ( .A1(\AES_ENC/us10/n587 ), .A2(\AES_ENC/us10/n855 ), .ZN(\AES_ENC/us10/n821 ) );
NAND2_X2 \AES_ENC/us10/U452  ( .A1(\AES_ENC/us10/n1093 ), .A2(\AES_ENC/us10/n821 ), .ZN(\AES_ENC/us10/n662 ) );
NAND2_X2 \AES_ENC/us10/U451  ( .A1(\AES_ENC/us10/n619 ), .A2(\AES_ENC/us10/n589 ), .ZN(\AES_ENC/us10/n650 ) );
NAND2_X2 \AES_ENC/us10/U450  ( .A1(\AES_ENC/us10/n956 ), .A2(\AES_ENC/us10/n650 ), .ZN(\AES_ENC/us10/n661 ) );
NAND2_X2 \AES_ENC/us10/U449  ( .A1(\AES_ENC/us10/n626 ), .A2(\AES_ENC/us10/n627 ), .ZN(\AES_ENC/us10/n839 ) );
OR2_X2 \AES_ENC/us10/U446  ( .A1(\AES_ENC/us10/n839 ), .A2(\AES_ENC/us10/n932 ), .ZN(\AES_ENC/us10/n656 ) );
NAND2_X2 \AES_ENC/us10/U445  ( .A1(\AES_ENC/us10/n621 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n1096 ) );
NAND2_X2 \AES_ENC/us10/U444  ( .A1(\AES_ENC/us10/n1030 ), .A2(\AES_ENC/us10/n1096 ), .ZN(\AES_ENC/us10/n651 ) );
NAND2_X2 \AES_ENC/us10/U443  ( .A1(\AES_ENC/us10/n1114 ), .A2(\AES_ENC/us10/n651 ), .ZN(\AES_ENC/us10/n655 ) );
OR3_X2 \AES_ENC/us10/U440  ( .A1(\AES_ENC/us10/n1079 ), .A2(\AES_ENC/sa10 [7]), .A3(\AES_ENC/us10/n626 ), .ZN(\AES_ENC/us10/n654 ));
NAND2_X2 \AES_ENC/us10/U439  ( .A1(\AES_ENC/us10/n593 ), .A2(\AES_ENC/us10/n601 ), .ZN(\AES_ENC/us10/n652 ) );
NAND4_X2 \AES_ENC/us10/U437  ( .A1(\AES_ENC/us10/n656 ), .A2(\AES_ENC/us10/n655 ), .A3(\AES_ENC/us10/n654 ), .A4(\AES_ENC/us10/n653 ), .ZN(\AES_ENC/us10/n657 ) );
NAND2_X2 \AES_ENC/us10/U436  ( .A1(\AES_ENC/sa10 [2]), .A2(\AES_ENC/us10/n657 ), .ZN(\AES_ENC/us10/n660 ) );
NAND4_X2 \AES_ENC/us10/U432  ( .A1(\AES_ENC/us10/n662 ), .A2(\AES_ENC/us10/n661 ), .A3(\AES_ENC/us10/n660 ), .A4(\AES_ENC/us10/n659 ), .ZN(\AES_ENC/us10/n663 ) );
NAND2_X2 \AES_ENC/us10/U431  ( .A1(\AES_ENC/us10/n663 ), .A2(\AES_ENC/us10/n574 ), .ZN(\AES_ENC/us10/n664 ) );
NAND2_X2 \AES_ENC/us10/U430  ( .A1(\AES_ENC/us10/n665 ), .A2(\AES_ENC/us10/n664 ), .ZN(\AES_ENC/us10/n666 ) );
NAND2_X2 \AES_ENC/us10/U429  ( .A1(\AES_ENC/sa10 [6]), .A2(\AES_ENC/us10/n666 ), .ZN(\AES_ENC/us10/n678 ) );
NAND2_X2 \AES_ENC/us10/U426  ( .A1(\AES_ENC/us10/n735 ), .A2(\AES_ENC/us10/n1093 ), .ZN(\AES_ENC/us10/n675 ) );
NAND2_X2 \AES_ENC/us10/U425  ( .A1(\AES_ENC/us10/n588 ), .A2(\AES_ENC/us10/n597 ), .ZN(\AES_ENC/us10/n1045 ) );
OR2_X2 \AES_ENC/us10/U424  ( .A1(\AES_ENC/us10/n1045 ), .A2(\AES_ENC/us10/n605 ), .ZN(\AES_ENC/us10/n674 ) );
NAND2_X2 \AES_ENC/us10/U423  ( .A1(\AES_ENC/sa10 [1]), .A2(\AES_ENC/us10/n620 ), .ZN(\AES_ENC/us10/n667 ) );
NAND2_X2 \AES_ENC/us10/U422  ( .A1(\AES_ENC/us10/n619 ), .A2(\AES_ENC/us10/n667 ), .ZN(\AES_ENC/us10/n1071 ) );
NAND4_X2 \AES_ENC/us10/U412  ( .A1(\AES_ENC/us10/n675 ), .A2(\AES_ENC/us10/n674 ), .A3(\AES_ENC/us10/n673 ), .A4(\AES_ENC/us10/n672 ), .ZN(\AES_ENC/us10/n676 ) );
NAND2_X2 \AES_ENC/us10/U411  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n676 ), .ZN(\AES_ENC/us10/n677 ) );
NAND2_X2 \AES_ENC/us10/U408  ( .A1(\AES_ENC/us10/n800 ), .A2(\AES_ENC/us10/n1022 ), .ZN(\AES_ENC/us10/n680 ) );
NAND2_X2 \AES_ENC/us10/U407  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n680 ), .ZN(\AES_ENC/us10/n681 ) );
AND2_X2 \AES_ENC/us10/U402  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n684 ), .ZN(\AES_ENC/us10/n682 ) );
NAND4_X2 \AES_ENC/us10/U395  ( .A1(\AES_ENC/us10/n691 ), .A2(\AES_ENC/us10/n581 ), .A3(\AES_ENC/us10/n690 ), .A4(\AES_ENC/us10/n689 ), .ZN(\AES_ENC/us10/n692 ) );
NAND2_X2 \AES_ENC/us10/U394  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n692 ), .ZN(\AES_ENC/us10/n733 ) );
NAND2_X2 \AES_ENC/us10/U392  ( .A1(\AES_ENC/us10/n977 ), .A2(\AES_ENC/us10/n1050 ), .ZN(\AES_ENC/us10/n702 ) );
NAND2_X2 \AES_ENC/us10/U391  ( .A1(\AES_ENC/us10/n1093 ), .A2(\AES_ENC/us10/n1045 ), .ZN(\AES_ENC/us10/n701 ) );
NAND4_X2 \AES_ENC/us10/U381  ( .A1(\AES_ENC/us10/n702 ), .A2(\AES_ENC/us10/n701 ), .A3(\AES_ENC/us10/n700 ), .A4(\AES_ENC/us10/n699 ), .ZN(\AES_ENC/us10/n703 ) );
NAND2_X2 \AES_ENC/us10/U380  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n703 ), .ZN(\AES_ENC/us10/n732 ) );
AND2_X2 \AES_ENC/us10/U379  ( .A1(\AES_ENC/sa10 [0]), .A2(\AES_ENC/sa10 [6]),.ZN(\AES_ENC/us10/n1113 ) );
NAND2_X2 \AES_ENC/us10/U378  ( .A1(\AES_ENC/us10/n601 ), .A2(\AES_ENC/us10/n1030 ), .ZN(\AES_ENC/us10/n881 ) );
NAND2_X2 \AES_ENC/us10/U377  ( .A1(\AES_ENC/us10/n1093 ), .A2(\AES_ENC/us10/n881 ), .ZN(\AES_ENC/us10/n715 ) );
NAND2_X2 \AES_ENC/us10/U376  ( .A1(\AES_ENC/us10/n1010 ), .A2(\AES_ENC/us10/n600 ), .ZN(\AES_ENC/us10/n714 ) );
NAND2_X2 \AES_ENC/us10/U375  ( .A1(\AES_ENC/us10/n855 ), .A2(\AES_ENC/us10/n588 ), .ZN(\AES_ENC/us10/n1117 ) );
XNOR2_X2 \AES_ENC/us10/U371  ( .A(\AES_ENC/us10/n611 ), .B(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n824 ) );
NAND4_X2 \AES_ENC/us10/U362  ( .A1(\AES_ENC/us10/n715 ), .A2(\AES_ENC/us10/n714 ), .A3(\AES_ENC/us10/n713 ), .A4(\AES_ENC/us10/n712 ), .ZN(\AES_ENC/us10/n716 ) );
NAND2_X2 \AES_ENC/us10/U361  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n716 ), .ZN(\AES_ENC/us10/n731 ) );
AND2_X2 \AES_ENC/us10/U360  ( .A1(\AES_ENC/sa10 [6]), .A2(\AES_ENC/us10/n574 ), .ZN(\AES_ENC/us10/n1131 ) );
NAND2_X2 \AES_ENC/us10/U359  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n717 ) );
NAND2_X2 \AES_ENC/us10/U358  ( .A1(\AES_ENC/us10/n1029 ), .A2(\AES_ENC/us10/n717 ), .ZN(\AES_ENC/us10/n728 ) );
NAND2_X2 \AES_ENC/us10/U357  ( .A1(\AES_ENC/sa10 [1]), .A2(\AES_ENC/us10/n624 ), .ZN(\AES_ENC/us10/n1097 ) );
NAND2_X2 \AES_ENC/us10/U356  ( .A1(\AES_ENC/us10/n603 ), .A2(\AES_ENC/us10/n1097 ), .ZN(\AES_ENC/us10/n718 ) );
NAND2_X2 \AES_ENC/us10/U355  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n718 ), .ZN(\AES_ENC/us10/n727 ) );
NAND4_X2 \AES_ENC/us10/U344  ( .A1(\AES_ENC/us10/n728 ), .A2(\AES_ENC/us10/n727 ), .A3(\AES_ENC/us10/n726 ), .A4(\AES_ENC/us10/n725 ), .ZN(\AES_ENC/us10/n729 ) );
NAND2_X2 \AES_ENC/us10/U343  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n729 ), .ZN(\AES_ENC/us10/n730 ) );
NAND4_X2 \AES_ENC/us10/U342  ( .A1(\AES_ENC/us10/n733 ), .A2(\AES_ENC/us10/n732 ), .A3(\AES_ENC/us10/n731 ), .A4(\AES_ENC/us10/n730 ), .ZN(\AES_ENC/sa10_sub[1] ) );
NAND2_X2 \AES_ENC/us10/U341  ( .A1(\AES_ENC/sa10 [7]), .A2(\AES_ENC/us10/n611 ), .ZN(\AES_ENC/us10/n734 ) );
NAND2_X2 \AES_ENC/us10/U340  ( .A1(\AES_ENC/us10/n734 ), .A2(\AES_ENC/us10/n607 ), .ZN(\AES_ENC/us10/n738 ) );
OR4_X2 \AES_ENC/us10/U339  ( .A1(\AES_ENC/us10/n738 ), .A2(\AES_ENC/us10/n626 ), .A3(\AES_ENC/us10/n826 ), .A4(\AES_ENC/us10/n1121 ), .ZN(\AES_ENC/us10/n746 ) );
NAND2_X2 \AES_ENC/us10/U337  ( .A1(\AES_ENC/us10/n1100 ), .A2(\AES_ENC/us10/n587 ), .ZN(\AES_ENC/us10/n992 ) );
OR2_X2 \AES_ENC/us10/U336  ( .A1(\AES_ENC/us10/n610 ), .A2(\AES_ENC/us10/n735 ), .ZN(\AES_ENC/us10/n737 ) );
NAND2_X2 \AES_ENC/us10/U334  ( .A1(\AES_ENC/us10/n619 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n753 ) );
NAND2_X2 \AES_ENC/us10/U333  ( .A1(\AES_ENC/us10/n582 ), .A2(\AES_ENC/us10/n753 ), .ZN(\AES_ENC/us10/n1080 ) );
NAND2_X2 \AES_ENC/us10/U332  ( .A1(\AES_ENC/us10/n1048 ), .A2(\AES_ENC/us10/n576 ), .ZN(\AES_ENC/us10/n736 ) );
NAND2_X2 \AES_ENC/us10/U331  ( .A1(\AES_ENC/us10/n737 ), .A2(\AES_ENC/us10/n736 ), .ZN(\AES_ENC/us10/n739 ) );
NAND2_X2 \AES_ENC/us10/U330  ( .A1(\AES_ENC/us10/n739 ), .A2(\AES_ENC/us10/n738 ), .ZN(\AES_ENC/us10/n745 ) );
NAND2_X2 \AES_ENC/us10/U326  ( .A1(\AES_ENC/us10/n1096 ), .A2(\AES_ENC/us10/n590 ), .ZN(\AES_ENC/us10/n906 ) );
NAND4_X2 \AES_ENC/us10/U323  ( .A1(\AES_ENC/us10/n746 ), .A2(\AES_ENC/us10/n992 ), .A3(\AES_ENC/us10/n745 ), .A4(\AES_ENC/us10/n744 ), .ZN(\AES_ENC/us10/n747 ) );
NAND2_X2 \AES_ENC/us10/U322  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n747 ), .ZN(\AES_ENC/us10/n793 ) );
NAND2_X2 \AES_ENC/us10/U321  ( .A1(\AES_ENC/us10/n584 ), .A2(\AES_ENC/us10/n855 ), .ZN(\AES_ENC/us10/n748 ) );
NAND2_X2 \AES_ENC/us10/U320  ( .A1(\AES_ENC/us10/n956 ), .A2(\AES_ENC/us10/n748 ), .ZN(\AES_ENC/us10/n760 ) );
NAND2_X2 \AES_ENC/us10/U313  ( .A1(\AES_ENC/us10/n590 ), .A2(\AES_ENC/us10/n753 ), .ZN(\AES_ENC/us10/n1023 ) );
NAND4_X2 \AES_ENC/us10/U308  ( .A1(\AES_ENC/us10/n760 ), .A2(\AES_ENC/us10/n992 ), .A3(\AES_ENC/us10/n759 ), .A4(\AES_ENC/us10/n758 ), .ZN(\AES_ENC/us10/n761 ) );
NAND2_X2 \AES_ENC/us10/U307  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n761 ), .ZN(\AES_ENC/us10/n792 ) );
NAND2_X2 \AES_ENC/us10/U306  ( .A1(\AES_ENC/us10/n584 ), .A2(\AES_ENC/us10/n603 ), .ZN(\AES_ENC/us10/n989 ) );
NAND2_X2 \AES_ENC/us10/U305  ( .A1(\AES_ENC/us10/n1050 ), .A2(\AES_ENC/us10/n989 ), .ZN(\AES_ENC/us10/n777 ) );
NAND2_X2 \AES_ENC/us10/U304  ( .A1(\AES_ENC/us10/n1093 ), .A2(\AES_ENC/us10/n762 ), .ZN(\AES_ENC/us10/n776 ) );
XNOR2_X2 \AES_ENC/us10/U301  ( .A(\AES_ENC/sa10 [7]), .B(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n959 ) );
NAND4_X2 \AES_ENC/us10/U289  ( .A1(\AES_ENC/us10/n777 ), .A2(\AES_ENC/us10/n776 ), .A3(\AES_ENC/us10/n775 ), .A4(\AES_ENC/us10/n774 ), .ZN(\AES_ENC/us10/n778 ) );
NAND2_X2 \AES_ENC/us10/U288  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n778 ), .ZN(\AES_ENC/us10/n791 ) );
NAND2_X2 \AES_ENC/us10/U287  ( .A1(\AES_ENC/us10/n1056 ), .A2(\AES_ENC/us10/n1050 ), .ZN(\AES_ENC/us10/n788 ) );
NAND2_X2 \AES_ENC/us10/U286  ( .A1(\AES_ENC/us10/n1091 ), .A2(\AES_ENC/us10/n779 ), .ZN(\AES_ENC/us10/n787 ) );
NAND2_X2 \AES_ENC/us10/U285  ( .A1(\AES_ENC/us10/n956 ), .A2(\AES_ENC/sa10 [1]), .ZN(\AES_ENC/us10/n786 ) );
NAND4_X2 \AES_ENC/us10/U278  ( .A1(\AES_ENC/us10/n788 ), .A2(\AES_ENC/us10/n787 ), .A3(\AES_ENC/us10/n786 ), .A4(\AES_ENC/us10/n785 ), .ZN(\AES_ENC/us10/n789 ) );
NAND2_X2 \AES_ENC/us10/U277  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n789 ), .ZN(\AES_ENC/us10/n790 ) );
NAND4_X2 \AES_ENC/us10/U276  ( .A1(\AES_ENC/us10/n793 ), .A2(\AES_ENC/us10/n792 ), .A3(\AES_ENC/us10/n791 ), .A4(\AES_ENC/us10/n790 ), .ZN(\AES_ENC/sa10_sub[2] ) );
NAND2_X2 \AES_ENC/us10/U275  ( .A1(\AES_ENC/us10/n1059 ), .A2(\AES_ENC/us10/n794 ), .ZN(\AES_ENC/us10/n810 ) );
NAND2_X2 \AES_ENC/us10/U274  ( .A1(\AES_ENC/us10/n1049 ), .A2(\AES_ENC/us10/n956 ), .ZN(\AES_ENC/us10/n809 ) );
OR2_X2 \AES_ENC/us10/U266  ( .A1(\AES_ENC/us10/n1096 ), .A2(\AES_ENC/us10/n606 ), .ZN(\AES_ENC/us10/n802 ) );
NAND2_X2 \AES_ENC/us10/U265  ( .A1(\AES_ENC/us10/n1053 ), .A2(\AES_ENC/us10/n800 ), .ZN(\AES_ENC/us10/n801 ) );
NAND2_X2 \AES_ENC/us10/U264  ( .A1(\AES_ENC/us10/n802 ), .A2(\AES_ENC/us10/n801 ), .ZN(\AES_ENC/us10/n805 ) );
NAND4_X2 \AES_ENC/us10/U261  ( .A1(\AES_ENC/us10/n810 ), .A2(\AES_ENC/us10/n809 ), .A3(\AES_ENC/us10/n808 ), .A4(\AES_ENC/us10/n807 ), .ZN(\AES_ENC/us10/n811 ) );
NAND2_X2 \AES_ENC/us10/U260  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n811 ), .ZN(\AES_ENC/us10/n852 ) );
OR2_X2 \AES_ENC/us10/U259  ( .A1(\AES_ENC/us10/n1023 ), .A2(\AES_ENC/us10/n617 ), .ZN(\AES_ENC/us10/n819 ) );
OR2_X2 \AES_ENC/us10/U257  ( .A1(\AES_ENC/us10/n570 ), .A2(\AES_ENC/us10/n930 ), .ZN(\AES_ENC/us10/n818 ) );
NAND2_X2 \AES_ENC/us10/U256  ( .A1(\AES_ENC/us10/n1013 ), .A2(\AES_ENC/us10/n1094 ), .ZN(\AES_ENC/us10/n817 ) );
NAND4_X2 \AES_ENC/us10/U249  ( .A1(\AES_ENC/us10/n819 ), .A2(\AES_ENC/us10/n818 ), .A3(\AES_ENC/us10/n817 ), .A4(\AES_ENC/us10/n816 ), .ZN(\AES_ENC/us10/n820 ) );
NAND2_X2 \AES_ENC/us10/U248  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n820 ), .ZN(\AES_ENC/us10/n851 ) );
NAND2_X2 \AES_ENC/us10/U247  ( .A1(\AES_ENC/us10/n956 ), .A2(\AES_ENC/us10/n1080 ), .ZN(\AES_ENC/us10/n835 ) );
NAND2_X2 \AES_ENC/us10/U246  ( .A1(\AES_ENC/us10/n570 ), .A2(\AES_ENC/us10/n1030 ), .ZN(\AES_ENC/us10/n1047 ) );
OR2_X2 \AES_ENC/us10/U245  ( .A1(\AES_ENC/us10/n1047 ), .A2(\AES_ENC/us10/n612 ), .ZN(\AES_ENC/us10/n834 ) );
NAND2_X2 \AES_ENC/us10/U244  ( .A1(\AES_ENC/us10/n1072 ), .A2(\AES_ENC/us10/n589 ), .ZN(\AES_ENC/us10/n833 ) );
NAND4_X2 \AES_ENC/us10/U233  ( .A1(\AES_ENC/us10/n835 ), .A2(\AES_ENC/us10/n834 ), .A3(\AES_ENC/us10/n833 ), .A4(\AES_ENC/us10/n832 ), .ZN(\AES_ENC/us10/n836 ) );
NAND2_X2 \AES_ENC/us10/U232  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n836 ), .ZN(\AES_ENC/us10/n850 ) );
NAND2_X2 \AES_ENC/us10/U231  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n623 ), .ZN(\AES_ENC/us10/n847 ) );
NAND2_X2 \AES_ENC/us10/U230  ( .A1(\AES_ENC/us10/n1050 ), .A2(\AES_ENC/us10/n1071 ), .ZN(\AES_ENC/us10/n846 ) );
OR2_X2 \AES_ENC/us10/U224  ( .A1(\AES_ENC/us10/n1053 ), .A2(\AES_ENC/us10/n911 ), .ZN(\AES_ENC/us10/n1077 ) );
NAND4_X2 \AES_ENC/us10/U220  ( .A1(\AES_ENC/us10/n847 ), .A2(\AES_ENC/us10/n846 ), .A3(\AES_ENC/us10/n845 ), .A4(\AES_ENC/us10/n844 ), .ZN(\AES_ENC/us10/n848 ) );
NAND2_X2 \AES_ENC/us10/U219  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n848 ), .ZN(\AES_ENC/us10/n849 ) );
NAND4_X2 \AES_ENC/us10/U218  ( .A1(\AES_ENC/us10/n852 ), .A2(\AES_ENC/us10/n851 ), .A3(\AES_ENC/us10/n850 ), .A4(\AES_ENC/us10/n849 ), .ZN(\AES_ENC/sa10_sub[3] ) );
NAND2_X2 \AES_ENC/us10/U216  ( .A1(\AES_ENC/us10/n1009 ), .A2(\AES_ENC/us10/n1072 ), .ZN(\AES_ENC/us10/n862 ) );
NAND2_X2 \AES_ENC/us10/U215  ( .A1(\AES_ENC/us10/n603 ), .A2(\AES_ENC/us10/n577 ), .ZN(\AES_ENC/us10/n853 ) );
NAND2_X2 \AES_ENC/us10/U214  ( .A1(\AES_ENC/us10/n1050 ), .A2(\AES_ENC/us10/n853 ), .ZN(\AES_ENC/us10/n861 ) );
NAND4_X2 \AES_ENC/us10/U206  ( .A1(\AES_ENC/us10/n862 ), .A2(\AES_ENC/us10/n861 ), .A3(\AES_ENC/us10/n860 ), .A4(\AES_ENC/us10/n859 ), .ZN(\AES_ENC/us10/n863 ) );
NAND2_X2 \AES_ENC/us10/U205  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n863 ), .ZN(\AES_ENC/us10/n905 ) );
NAND2_X2 \AES_ENC/us10/U204  ( .A1(\AES_ENC/us10/n1010 ), .A2(\AES_ENC/us10/n989 ), .ZN(\AES_ENC/us10/n874 ) );
NAND2_X2 \AES_ENC/us10/U203  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n610 ), .ZN(\AES_ENC/us10/n864 ) );
NAND2_X2 \AES_ENC/us10/U202  ( .A1(\AES_ENC/us10/n929 ), .A2(\AES_ENC/us10/n864 ), .ZN(\AES_ENC/us10/n873 ) );
NAND4_X2 \AES_ENC/us10/U193  ( .A1(\AES_ENC/us10/n874 ), .A2(\AES_ENC/us10/n873 ), .A3(\AES_ENC/us10/n872 ), .A4(\AES_ENC/us10/n871 ), .ZN(\AES_ENC/us10/n875 ) );
NAND2_X2 \AES_ENC/us10/U192  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n875 ), .ZN(\AES_ENC/us10/n904 ) );
NAND2_X2 \AES_ENC/us10/U191  ( .A1(\AES_ENC/us10/n583 ), .A2(\AES_ENC/us10/n1050 ), .ZN(\AES_ENC/us10/n889 ) );
NAND2_X2 \AES_ENC/us10/U190  ( .A1(\AES_ENC/us10/n1093 ), .A2(\AES_ENC/us10/n587 ), .ZN(\AES_ENC/us10/n876 ) );
NAND2_X2 \AES_ENC/us10/U189  ( .A1(\AES_ENC/us10/n604 ), .A2(\AES_ENC/us10/n876 ), .ZN(\AES_ENC/us10/n877 ) );
NAND2_X2 \AES_ENC/us10/U188  ( .A1(\AES_ENC/us10/n877 ), .A2(\AES_ENC/us10/n623 ), .ZN(\AES_ENC/us10/n888 ) );
NAND4_X2 \AES_ENC/us10/U179  ( .A1(\AES_ENC/us10/n889 ), .A2(\AES_ENC/us10/n888 ), .A3(\AES_ENC/us10/n887 ), .A4(\AES_ENC/us10/n886 ), .ZN(\AES_ENC/us10/n890 ) );
NAND2_X2 \AES_ENC/us10/U178  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n890 ), .ZN(\AES_ENC/us10/n903 ) );
OR2_X2 \AES_ENC/us10/U177  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n1059 ), .ZN(\AES_ENC/us10/n900 ) );
NAND2_X2 \AES_ENC/us10/U176  ( .A1(\AES_ENC/us10/n1073 ), .A2(\AES_ENC/us10/n1047 ), .ZN(\AES_ENC/us10/n899 ) );
NAND2_X2 \AES_ENC/us10/U175  ( .A1(\AES_ENC/us10/n1094 ), .A2(\AES_ENC/us10/n595 ), .ZN(\AES_ENC/us10/n898 ) );
NAND4_X2 \AES_ENC/us10/U167  ( .A1(\AES_ENC/us10/n900 ), .A2(\AES_ENC/us10/n899 ), .A3(\AES_ENC/us10/n898 ), .A4(\AES_ENC/us10/n897 ), .ZN(\AES_ENC/us10/n901 ) );
NAND2_X2 \AES_ENC/us10/U166  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n901 ), .ZN(\AES_ENC/us10/n902 ) );
NAND4_X2 \AES_ENC/us10/U165  ( .A1(\AES_ENC/us10/n905 ), .A2(\AES_ENC/us10/n904 ), .A3(\AES_ENC/us10/n903 ), .A4(\AES_ENC/us10/n902 ), .ZN(\AES_ENC/sa10_sub[4] ) );
NAND2_X2 \AES_ENC/us10/U164  ( .A1(\AES_ENC/us10/n1094 ), .A2(\AES_ENC/us10/n599 ), .ZN(\AES_ENC/us10/n922 ) );
NAND2_X2 \AES_ENC/us10/U163  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n989 ), .ZN(\AES_ENC/us10/n921 ) );
NAND4_X2 \AES_ENC/us10/U151  ( .A1(\AES_ENC/us10/n922 ), .A2(\AES_ENC/us10/n921 ), .A3(\AES_ENC/us10/n920 ), .A4(\AES_ENC/us10/n919 ), .ZN(\AES_ENC/us10/n923 ) );
NAND2_X2 \AES_ENC/us10/U150  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n923 ), .ZN(\AES_ENC/us10/n972 ) );
NAND2_X2 \AES_ENC/us10/U149  ( .A1(\AES_ENC/us10/n582 ), .A2(\AES_ENC/us10/n619 ), .ZN(\AES_ENC/us10/n924 ) );
NAND2_X2 \AES_ENC/us10/U148  ( .A1(\AES_ENC/us10/n1073 ), .A2(\AES_ENC/us10/n924 ), .ZN(\AES_ENC/us10/n939 ) );
NAND2_X2 \AES_ENC/us10/U147  ( .A1(\AES_ENC/us10/n926 ), .A2(\AES_ENC/us10/n925 ), .ZN(\AES_ENC/us10/n927 ) );
NAND2_X2 \AES_ENC/us10/U146  ( .A1(\AES_ENC/us10/n606 ), .A2(\AES_ENC/us10/n927 ), .ZN(\AES_ENC/us10/n928 ) );
NAND2_X2 \AES_ENC/us10/U145  ( .A1(\AES_ENC/us10/n928 ), .A2(\AES_ENC/us10/n1080 ), .ZN(\AES_ENC/us10/n938 ) );
OR2_X2 \AES_ENC/us10/U144  ( .A1(\AES_ENC/us10/n1117 ), .A2(\AES_ENC/us10/n615 ), .ZN(\AES_ENC/us10/n937 ) );
NAND4_X2 \AES_ENC/us10/U139  ( .A1(\AES_ENC/us10/n939 ), .A2(\AES_ENC/us10/n938 ), .A3(\AES_ENC/us10/n937 ), .A4(\AES_ENC/us10/n936 ), .ZN(\AES_ENC/us10/n940 ) );
NAND2_X2 \AES_ENC/us10/U138  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n940 ), .ZN(\AES_ENC/us10/n971 ) );
OR2_X2 \AES_ENC/us10/U137  ( .A1(\AES_ENC/us10/n605 ), .A2(\AES_ENC/us10/n941 ), .ZN(\AES_ENC/us10/n954 ) );
NAND2_X2 \AES_ENC/us10/U136  ( .A1(\AES_ENC/us10/n1096 ), .A2(\AES_ENC/us10/n577 ), .ZN(\AES_ENC/us10/n942 ) );
NAND2_X2 \AES_ENC/us10/U135  ( .A1(\AES_ENC/us10/n1048 ), .A2(\AES_ENC/us10/n942 ), .ZN(\AES_ENC/us10/n943 ) );
NAND2_X2 \AES_ENC/us10/U134  ( .A1(\AES_ENC/us10/n612 ), .A2(\AES_ENC/us10/n943 ), .ZN(\AES_ENC/us10/n944 ) );
NAND2_X2 \AES_ENC/us10/U133  ( .A1(\AES_ENC/us10/n944 ), .A2(\AES_ENC/us10/n580 ), .ZN(\AES_ENC/us10/n953 ) );
NAND4_X2 \AES_ENC/us10/U125  ( .A1(\AES_ENC/us10/n954 ), .A2(\AES_ENC/us10/n953 ), .A3(\AES_ENC/us10/n952 ), .A4(\AES_ENC/us10/n951 ), .ZN(\AES_ENC/us10/n955 ) );
NAND2_X2 \AES_ENC/us10/U124  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n955 ), .ZN(\AES_ENC/us10/n970 ) );
NAND2_X2 \AES_ENC/us10/U123  ( .A1(\AES_ENC/us10/n1094 ), .A2(\AES_ENC/us10/n1071 ), .ZN(\AES_ENC/us10/n967 ) );
NAND2_X2 \AES_ENC/us10/U122  ( .A1(\AES_ENC/us10/n956 ), .A2(\AES_ENC/us10/n1030 ), .ZN(\AES_ENC/us10/n966 ) );
NAND4_X2 \AES_ENC/us10/U114  ( .A1(\AES_ENC/us10/n967 ), .A2(\AES_ENC/us10/n966 ), .A3(\AES_ENC/us10/n965 ), .A4(\AES_ENC/us10/n964 ), .ZN(\AES_ENC/us10/n968 ) );
NAND2_X2 \AES_ENC/us10/U113  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n968 ), .ZN(\AES_ENC/us10/n969 ) );
NAND4_X2 \AES_ENC/us10/U112  ( .A1(\AES_ENC/us10/n972 ), .A2(\AES_ENC/us10/n971 ), .A3(\AES_ENC/us10/n970 ), .A4(\AES_ENC/us10/n969 ), .ZN(\AES_ENC/sa10_sub[5] ) );
NAND2_X2 \AES_ENC/us10/U111  ( .A1(\AES_ENC/us10/n570 ), .A2(\AES_ENC/us10/n1097 ), .ZN(\AES_ENC/us10/n973 ) );
NAND2_X2 \AES_ENC/us10/U110  ( .A1(\AES_ENC/us10/n1073 ), .A2(\AES_ENC/us10/n973 ), .ZN(\AES_ENC/us10/n987 ) );
NAND2_X2 \AES_ENC/us10/U109  ( .A1(\AES_ENC/us10/n974 ), .A2(\AES_ENC/us10/n1077 ), .ZN(\AES_ENC/us10/n975 ) );
NAND2_X2 \AES_ENC/us10/U108  ( .A1(\AES_ENC/us10/n613 ), .A2(\AES_ENC/us10/n975 ), .ZN(\AES_ENC/us10/n976 ) );
NAND2_X2 \AES_ENC/us10/U107  ( .A1(\AES_ENC/us10/n977 ), .A2(\AES_ENC/us10/n976 ), .ZN(\AES_ENC/us10/n986 ) );
NAND4_X2 \AES_ENC/us10/U99  ( .A1(\AES_ENC/us10/n987 ), .A2(\AES_ENC/us10/n986 ), .A3(\AES_ENC/us10/n985 ), .A4(\AES_ENC/us10/n984 ), .ZN(\AES_ENC/us10/n988 ) );
NAND2_X2 \AES_ENC/us10/U98  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n988 ), .ZN(\AES_ENC/us10/n1044 ) );
NAND2_X2 \AES_ENC/us10/U97  ( .A1(\AES_ENC/us10/n1073 ), .A2(\AES_ENC/us10/n989 ), .ZN(\AES_ENC/us10/n1004 ) );
NAND2_X2 \AES_ENC/us10/U96  ( .A1(\AES_ENC/us10/n1092 ), .A2(\AES_ENC/us10/n619 ), .ZN(\AES_ENC/us10/n1003 ) );
NAND4_X2 \AES_ENC/us10/U85  ( .A1(\AES_ENC/us10/n1004 ), .A2(\AES_ENC/us10/n1003 ), .A3(\AES_ENC/us10/n1002 ), .A4(\AES_ENC/us10/n1001 ), .ZN(\AES_ENC/us10/n1005 ) );
NAND2_X2 \AES_ENC/us10/U84  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n1005 ), .ZN(\AES_ENC/us10/n1043 ) );
NAND2_X2 \AES_ENC/us10/U83  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n596 ), .ZN(\AES_ENC/us10/n1020 ) );
NAND2_X2 \AES_ENC/us10/U82  ( .A1(\AES_ENC/us10/n1050 ), .A2(\AES_ENC/us10/n624 ), .ZN(\AES_ENC/us10/n1019 ) );
NAND2_X2 \AES_ENC/us10/U77  ( .A1(\AES_ENC/us10/n1059 ), .A2(\AES_ENC/us10/n1114 ), .ZN(\AES_ENC/us10/n1012 ) );
NAND2_X2 \AES_ENC/us10/U76  ( .A1(\AES_ENC/us10/n1010 ), .A2(\AES_ENC/us10/n592 ), .ZN(\AES_ENC/us10/n1011 ) );
NAND2_X2 \AES_ENC/us10/U75  ( .A1(\AES_ENC/us10/n1012 ), .A2(\AES_ENC/us10/n1011 ), .ZN(\AES_ENC/us10/n1016 ) );
NAND4_X2 \AES_ENC/us10/U70  ( .A1(\AES_ENC/us10/n1020 ), .A2(\AES_ENC/us10/n1019 ), .A3(\AES_ENC/us10/n1018 ), .A4(\AES_ENC/us10/n1017 ), .ZN(\AES_ENC/us10/n1021 ) );
NAND2_X2 \AES_ENC/us10/U69  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n1021 ), .ZN(\AES_ENC/us10/n1042 ) );
NAND2_X2 \AES_ENC/us10/U68  ( .A1(\AES_ENC/us10/n1022 ), .A2(\AES_ENC/us10/n1093 ), .ZN(\AES_ENC/us10/n1039 ) );
NAND2_X2 \AES_ENC/us10/U67  ( .A1(\AES_ENC/us10/n1050 ), .A2(\AES_ENC/us10/n1023 ), .ZN(\AES_ENC/us10/n1038 ) );
NAND2_X2 \AES_ENC/us10/U66  ( .A1(\AES_ENC/us10/n1024 ), .A2(\AES_ENC/us10/n1071 ), .ZN(\AES_ENC/us10/n1037 ) );
AND2_X2 \AES_ENC/us10/U60  ( .A1(\AES_ENC/us10/n1030 ), .A2(\AES_ENC/us10/n602 ), .ZN(\AES_ENC/us10/n1078 ) );
NAND4_X2 \AES_ENC/us10/U56  ( .A1(\AES_ENC/us10/n1039 ), .A2(\AES_ENC/us10/n1038 ), .A3(\AES_ENC/us10/n1037 ), .A4(\AES_ENC/us10/n1036 ), .ZN(\AES_ENC/us10/n1040 ) );
NAND2_X2 \AES_ENC/us10/U55  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n1040 ), .ZN(\AES_ENC/us10/n1041 ) );
NAND4_X2 \AES_ENC/us10/U54  ( .A1(\AES_ENC/us10/n1044 ), .A2(\AES_ENC/us10/n1043 ), .A3(\AES_ENC/us10/n1042 ), .A4(\AES_ENC/us10/n1041 ), .ZN(\AES_ENC/sa10_sub[6] ) );
NAND2_X2 \AES_ENC/us10/U53  ( .A1(\AES_ENC/us10/n1072 ), .A2(\AES_ENC/us10/n1045 ), .ZN(\AES_ENC/us10/n1068 ) );
NAND2_X2 \AES_ENC/us10/U52  ( .A1(\AES_ENC/us10/n1046 ), .A2(\AES_ENC/us10/n582 ), .ZN(\AES_ENC/us10/n1067 ) );
NAND2_X2 \AES_ENC/us10/U51  ( .A1(\AES_ENC/us10/n1094 ), .A2(\AES_ENC/us10/n1047 ), .ZN(\AES_ENC/us10/n1066 ) );
NAND4_X2 \AES_ENC/us10/U40  ( .A1(\AES_ENC/us10/n1068 ), .A2(\AES_ENC/us10/n1067 ), .A3(\AES_ENC/us10/n1066 ), .A4(\AES_ENC/us10/n1065 ), .ZN(\AES_ENC/us10/n1069 ) );
NAND2_X2 \AES_ENC/us10/U39  ( .A1(\AES_ENC/us10/n1070 ), .A2(\AES_ENC/us10/n1069 ), .ZN(\AES_ENC/us10/n1135 ) );
NAND2_X2 \AES_ENC/us10/U38  ( .A1(\AES_ENC/us10/n1072 ), .A2(\AES_ENC/us10/n1071 ), .ZN(\AES_ENC/us10/n1088 ) );
NAND2_X2 \AES_ENC/us10/U37  ( .A1(\AES_ENC/us10/n1073 ), .A2(\AES_ENC/us10/n595 ), .ZN(\AES_ENC/us10/n1087 ) );
NAND4_X2 \AES_ENC/us10/U28  ( .A1(\AES_ENC/us10/n1088 ), .A2(\AES_ENC/us10/n1087 ), .A3(\AES_ENC/us10/n1086 ), .A4(\AES_ENC/us10/n1085 ), .ZN(\AES_ENC/us10/n1089 ) );
NAND2_X2 \AES_ENC/us10/U27  ( .A1(\AES_ENC/us10/n1090 ), .A2(\AES_ENC/us10/n1089 ), .ZN(\AES_ENC/us10/n1134 ) );
NAND2_X2 \AES_ENC/us10/U26  ( .A1(\AES_ENC/us10/n1091 ), .A2(\AES_ENC/us10/n1093 ), .ZN(\AES_ENC/us10/n1111 ) );
NAND2_X2 \AES_ENC/us10/U25  ( .A1(\AES_ENC/us10/n1092 ), .A2(\AES_ENC/us10/n1120 ), .ZN(\AES_ENC/us10/n1110 ) );
AND2_X2 \AES_ENC/us10/U22  ( .A1(\AES_ENC/us10/n1097 ), .A2(\AES_ENC/us10/n1096 ), .ZN(\AES_ENC/us10/n1098 ) );
NAND4_X2 \AES_ENC/us10/U14  ( .A1(\AES_ENC/us10/n1111 ), .A2(\AES_ENC/us10/n1110 ), .A3(\AES_ENC/us10/n1109 ), .A4(\AES_ENC/us10/n1108 ), .ZN(\AES_ENC/us10/n1112 ) );
NAND2_X2 \AES_ENC/us10/U13  ( .A1(\AES_ENC/us10/n1113 ), .A2(\AES_ENC/us10/n1112 ), .ZN(\AES_ENC/us10/n1133 ) );
NAND2_X2 \AES_ENC/us10/U12  ( .A1(\AES_ENC/us10/n1115 ), .A2(\AES_ENC/us10/n1114 ), .ZN(\AES_ENC/us10/n1129 ) );
OR2_X2 \AES_ENC/us10/U11  ( .A1(\AES_ENC/us10/n608 ), .A2(\AES_ENC/us10/n1116 ), .ZN(\AES_ENC/us10/n1128 ) );
NAND4_X2 \AES_ENC/us10/U3  ( .A1(\AES_ENC/us10/n1129 ), .A2(\AES_ENC/us10/n1128 ), .A3(\AES_ENC/us10/n1127 ), .A4(\AES_ENC/us10/n1126 ), .ZN(\AES_ENC/us10/n1130 ) );
NAND2_X2 \AES_ENC/us10/U2  ( .A1(\AES_ENC/us10/n1131 ), .A2(\AES_ENC/us10/n1130 ), .ZN(\AES_ENC/us10/n1132 ) );
NAND4_X2 \AES_ENC/us10/U1  ( .A1(\AES_ENC/us10/n1135 ), .A2(\AES_ENC/us10/n1134 ), .A3(\AES_ENC/us10/n1133 ), .A4(\AES_ENC/us10/n1132 ), .ZN(\AES_ENC/sa10_sub[7] ) );
INV_X4 \AES_ENC/us11/U575  ( .A(\AES_ENC/sa11 [7]), .ZN(\AES_ENC/us11/n627 ));
INV_X4 \AES_ENC/us11/U574  ( .A(\AES_ENC/us11/n1114 ), .ZN(\AES_ENC/us11/n625 ) );
INV_X4 \AES_ENC/us11/U573  ( .A(\AES_ENC/sa11 [4]), .ZN(\AES_ENC/us11/n624 ));
INV_X4 \AES_ENC/us11/U572  ( .A(\AES_ENC/us11/n1025 ), .ZN(\AES_ENC/us11/n622 ) );
INV_X4 \AES_ENC/us11/U571  ( .A(\AES_ENC/us11/n1120 ), .ZN(\AES_ENC/us11/n620 ) );
INV_X4 \AES_ENC/us11/U570  ( .A(\AES_ENC/us11/n1121 ), .ZN(\AES_ENC/us11/n619 ) );
INV_X4 \AES_ENC/us11/U569  ( .A(\AES_ENC/us11/n1048 ), .ZN(\AES_ENC/us11/n618 ) );
INV_X4 \AES_ENC/us11/U568  ( .A(\AES_ENC/us11/n974 ), .ZN(\AES_ENC/us11/n616 ) );
INV_X4 \AES_ENC/us11/U567  ( .A(\AES_ENC/us11/n794 ), .ZN(\AES_ENC/us11/n614 ) );
INV_X4 \AES_ENC/us11/U566  ( .A(\AES_ENC/sa11 [2]), .ZN(\AES_ENC/us11/n611 ));
INV_X4 \AES_ENC/us11/U565  ( .A(\AES_ENC/us11/n800 ), .ZN(\AES_ENC/us11/n610 ) );
INV_X4 \AES_ENC/us11/U564  ( .A(\AES_ENC/us11/n925 ), .ZN(\AES_ENC/us11/n609 ) );
INV_X4 \AES_ENC/us11/U563  ( .A(\AES_ENC/us11/n779 ), .ZN(\AES_ENC/us11/n607 ) );
INV_X4 \AES_ENC/us11/U562  ( .A(\AES_ENC/us11/n1022 ), .ZN(\AES_ENC/us11/n603 ) );
INV_X4 \AES_ENC/us11/U561  ( .A(\AES_ENC/us11/n1102 ), .ZN(\AES_ENC/us11/n602 ) );
INV_X4 \AES_ENC/us11/U560  ( .A(\AES_ENC/us11/n929 ), .ZN(\AES_ENC/us11/n601 ) );
INV_X4 \AES_ENC/us11/U559  ( .A(\AES_ENC/us11/n1056 ), .ZN(\AES_ENC/us11/n600 ) );
INV_X4 \AES_ENC/us11/U558  ( .A(\AES_ENC/us11/n1054 ), .ZN(\AES_ENC/us11/n599 ) );
INV_X4 \AES_ENC/us11/U557  ( .A(\AES_ENC/us11/n881 ), .ZN(\AES_ENC/us11/n598 ) );
INV_X4 \AES_ENC/us11/U556  ( .A(\AES_ENC/us11/n926 ), .ZN(\AES_ENC/us11/n597 ) );
INV_X4 \AES_ENC/us11/U555  ( .A(\AES_ENC/us11/n977 ), .ZN(\AES_ENC/us11/n595 ) );
INV_X4 \AES_ENC/us11/U554  ( .A(\AES_ENC/us11/n1031 ), .ZN(\AES_ENC/us11/n594 ) );
INV_X4 \AES_ENC/us11/U553  ( .A(\AES_ENC/us11/n1103 ), .ZN(\AES_ENC/us11/n593 ) );
INV_X4 \AES_ENC/us11/U552  ( .A(\AES_ENC/us11/n1009 ), .ZN(\AES_ENC/us11/n592 ) );
INV_X4 \AES_ENC/us11/U551  ( .A(\AES_ENC/us11/n990 ), .ZN(\AES_ENC/us11/n591 ) );
INV_X4 \AES_ENC/us11/U550  ( .A(\AES_ENC/us11/n1058 ), .ZN(\AES_ENC/us11/n590 ) );
INV_X4 \AES_ENC/us11/U549  ( .A(\AES_ENC/us11/n1074 ), .ZN(\AES_ENC/us11/n589 ) );
INV_X4 \AES_ENC/us11/U548  ( .A(\AES_ENC/us11/n1053 ), .ZN(\AES_ENC/us11/n588 ) );
INV_X4 \AES_ENC/us11/U547  ( .A(\AES_ENC/us11/n826 ), .ZN(\AES_ENC/us11/n587 ) );
INV_X4 \AES_ENC/us11/U546  ( .A(\AES_ENC/us11/n992 ), .ZN(\AES_ENC/us11/n586 ) );
INV_X4 \AES_ENC/us11/U545  ( .A(\AES_ENC/us11/n821 ), .ZN(\AES_ENC/us11/n585 ) );
INV_X4 \AES_ENC/us11/U544  ( .A(\AES_ENC/us11/n910 ), .ZN(\AES_ENC/us11/n584 ) );
INV_X4 \AES_ENC/us11/U543  ( .A(\AES_ENC/us11/n906 ), .ZN(\AES_ENC/us11/n583 ) );
INV_X4 \AES_ENC/us11/U542  ( .A(\AES_ENC/us11/n880 ), .ZN(\AES_ENC/us11/n581 ) );
INV_X4 \AES_ENC/us11/U541  ( .A(\AES_ENC/us11/n1013 ), .ZN(\AES_ENC/us11/n580 ) );
INV_X4 \AES_ENC/us11/U540  ( .A(\AES_ENC/us11/n1092 ), .ZN(\AES_ENC/us11/n579 ) );
INV_X4 \AES_ENC/us11/U539  ( .A(\AES_ENC/us11/n824 ), .ZN(\AES_ENC/us11/n578 ) );
INV_X4 \AES_ENC/us11/U538  ( .A(\AES_ENC/us11/n1091 ), .ZN(\AES_ENC/us11/n577 ) );
INV_X4 \AES_ENC/us11/U537  ( .A(\AES_ENC/us11/n1080 ), .ZN(\AES_ENC/us11/n576 ) );
INV_X4 \AES_ENC/us11/U536  ( .A(\AES_ENC/us11/n959 ), .ZN(\AES_ENC/us11/n575 ) );
INV_X4 \AES_ENC/us11/U535  ( .A(\AES_ENC/sa11 [0]), .ZN(\AES_ENC/us11/n574 ));
NOR2_X2 \AES_ENC/us11/U534  ( .A1(\AES_ENC/sa11 [0]), .A2(\AES_ENC/sa11 [6]),.ZN(\AES_ENC/us11/n1090 ) );
NOR2_X2 \AES_ENC/us11/U533  ( .A1(\AES_ENC/us11/n574 ), .A2(\AES_ENC/sa11 [6]), .ZN(\AES_ENC/us11/n1070 ) );
NOR2_X2 \AES_ENC/us11/U532  ( .A1(\AES_ENC/sa11 [4]), .A2(\AES_ENC/sa11 [3]),.ZN(\AES_ENC/us11/n1025 ) );
INV_X4 \AES_ENC/us11/U531  ( .A(\AES_ENC/us11/n569 ), .ZN(\AES_ENC/us11/n572 ) );
NOR2_X2 \AES_ENC/us11/U530  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n765 ) );
NOR2_X2 \AES_ENC/us11/U529  ( .A1(\AES_ENC/sa11 [4]), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n764 ) );
NOR2_X2 \AES_ENC/us11/U528  ( .A1(\AES_ENC/us11/n765 ), .A2(\AES_ENC/us11/n764 ), .ZN(\AES_ENC/us11/n766 ) );
NOR2_X2 \AES_ENC/us11/U527  ( .A1(\AES_ENC/us11/n766 ), .A2(\AES_ENC/us11/n575 ), .ZN(\AES_ENC/us11/n767 ) );
NOR3_X2 \AES_ENC/us11/U526  ( .A1(\AES_ENC/us11/n627 ), .A2(\AES_ENC/sa11 [5]), .A3(\AES_ENC/us11/n704 ), .ZN(\AES_ENC/us11/n706 ));
NOR2_X2 \AES_ENC/us11/U525  ( .A1(\AES_ENC/us11/n1117 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n707 ) );
NOR2_X2 \AES_ENC/us11/U524  ( .A1(\AES_ENC/sa11 [4]), .A2(\AES_ENC/us11/n579 ), .ZN(\AES_ENC/us11/n705 ) );
NOR3_X2 \AES_ENC/us11/U523  ( .A1(\AES_ENC/us11/n707 ), .A2(\AES_ENC/us11/n706 ), .A3(\AES_ENC/us11/n705 ), .ZN(\AES_ENC/us11/n713 ) );
INV_X4 \AES_ENC/us11/U522  ( .A(\AES_ENC/sa11 [3]), .ZN(\AES_ENC/us11/n621 ));
NAND3_X2 \AES_ENC/us11/U521  ( .A1(\AES_ENC/us11/n652 ), .A2(\AES_ENC/us11/n626 ), .A3(\AES_ENC/sa11 [7]), .ZN(\AES_ENC/us11/n653 ));
NOR2_X2 \AES_ENC/us11/U520  ( .A1(\AES_ENC/us11/n611 ), .A2(\AES_ENC/sa11 [5]), .ZN(\AES_ENC/us11/n925 ) );
NOR2_X2 \AES_ENC/us11/U519  ( .A1(\AES_ENC/sa11 [5]), .A2(\AES_ENC/sa11 [2]),.ZN(\AES_ENC/us11/n974 ) );
INV_X4 \AES_ENC/us11/U518  ( .A(\AES_ENC/sa11 [5]), .ZN(\AES_ENC/us11/n626 ));
NOR2_X2 \AES_ENC/us11/U517  ( .A1(\AES_ENC/us11/n611 ), .A2(\AES_ENC/sa11 [7]), .ZN(\AES_ENC/us11/n779 ) );
NAND3_X2 \AES_ENC/us11/U516  ( .A1(\AES_ENC/us11/n679 ), .A2(\AES_ENC/us11/n678 ), .A3(\AES_ENC/us11/n677 ), .ZN(\AES_ENC/sa11_sub[0] ) );
NOR2_X2 \AES_ENC/us11/U515  ( .A1(\AES_ENC/us11/n626 ), .A2(\AES_ENC/sa11 [2]), .ZN(\AES_ENC/us11/n1048 ) );
NOR4_X2 \AES_ENC/us11/U512  ( .A1(\AES_ENC/us11/n633 ), .A2(\AES_ENC/us11/n632 ), .A3(\AES_ENC/us11/n631 ), .A4(\AES_ENC/us11/n630 ), .ZN(\AES_ENC/us11/n634 ) );
NOR2_X2 \AES_ENC/us11/U510  ( .A1(\AES_ENC/us11/n629 ), .A2(\AES_ENC/us11/n628 ), .ZN(\AES_ENC/us11/n635 ) );
NAND3_X2 \AES_ENC/us11/U509  ( .A1(\AES_ENC/sa11 [2]), .A2(\AES_ENC/sa11 [7]), .A3(\AES_ENC/us11/n1059 ), .ZN(\AES_ENC/us11/n636 ) );
NOR2_X2 \AES_ENC/us11/U508  ( .A1(\AES_ENC/sa11 [7]), .A2(\AES_ENC/sa11 [2]),.ZN(\AES_ENC/us11/n794 ) );
NOR2_X2 \AES_ENC/us11/U507  ( .A1(\AES_ENC/sa11 [4]), .A2(\AES_ENC/sa11 [1]),.ZN(\AES_ENC/us11/n1102 ) );
NOR2_X2 \AES_ENC/us11/U506  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/sa11 [3]), .ZN(\AES_ENC/us11/n1053 ) );
NOR2_X2 \AES_ENC/us11/U505  ( .A1(\AES_ENC/us11/n607 ), .A2(\AES_ENC/sa11 [5]), .ZN(\AES_ENC/us11/n1024 ) );
NOR2_X2 \AES_ENC/us11/U504  ( .A1(\AES_ENC/us11/n625 ), .A2(\AES_ENC/sa11 [2]), .ZN(\AES_ENC/us11/n1093 ) );
NOR2_X2 \AES_ENC/us11/U503  ( .A1(\AES_ENC/us11/n614 ), .A2(\AES_ENC/sa11 [5]), .ZN(\AES_ENC/us11/n1094 ) );
NOR2_X2 \AES_ENC/us11/U502  ( .A1(\AES_ENC/us11/n624 ), .A2(\AES_ENC/sa11 [3]), .ZN(\AES_ENC/us11/n931 ) );
INV_X4 \AES_ENC/us11/U501  ( .A(\AES_ENC/us11/n570 ), .ZN(\AES_ENC/us11/n573 ) );
NOR2_X2 \AES_ENC/us11/U500  ( .A1(\AES_ENC/us11/n1053 ), .A2(\AES_ENC/us11/n1095 ), .ZN(\AES_ENC/us11/n639 ) );
NOR3_X2 \AES_ENC/us11/U499  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n573 ), .A3(\AES_ENC/us11/n1074 ), .ZN(\AES_ENC/us11/n641 ) );
NOR2_X2 \AES_ENC/us11/U498  ( .A1(\AES_ENC/us11/n639 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n640 ) );
NOR2_X2 \AES_ENC/us11/U497  ( .A1(\AES_ENC/us11/n641 ), .A2(\AES_ENC/us11/n640 ), .ZN(\AES_ENC/us11/n646 ) );
NOR3_X2 \AES_ENC/us11/U496  ( .A1(\AES_ENC/us11/n995 ), .A2(\AES_ENC/us11/n586 ), .A3(\AES_ENC/us11/n994 ), .ZN(\AES_ENC/us11/n1002 ) );
NOR2_X2 \AES_ENC/us11/U495  ( .A1(\AES_ENC/us11/n909 ), .A2(\AES_ENC/us11/n908 ), .ZN(\AES_ENC/us11/n920 ) );
NOR2_X2 \AES_ENC/us11/U494  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n823 ) );
NOR2_X2 \AES_ENC/us11/U492  ( .A1(\AES_ENC/us11/n624 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n822 ) );
NOR2_X2 \AES_ENC/us11/U491  ( .A1(\AES_ENC/us11/n823 ), .A2(\AES_ENC/us11/n822 ), .ZN(\AES_ENC/us11/n825 ) );
NOR2_X2 \AES_ENC/us11/U490  ( .A1(\AES_ENC/sa11 [1]), .A2(\AES_ENC/us11/n623 ), .ZN(\AES_ENC/us11/n913 ) );
NOR2_X2 \AES_ENC/us11/U489  ( .A1(\AES_ENC/us11/n913 ), .A2(\AES_ENC/us11/n1091 ), .ZN(\AES_ENC/us11/n914 ) );
NOR2_X2 \AES_ENC/us11/U488  ( .A1(\AES_ENC/us11/n826 ), .A2(\AES_ENC/us11/n572 ), .ZN(\AES_ENC/us11/n827 ) );
NOR3_X2 \AES_ENC/us11/U487  ( .A1(\AES_ENC/us11/n769 ), .A2(\AES_ENC/us11/n768 ), .A3(\AES_ENC/us11/n767 ), .ZN(\AES_ENC/us11/n775 ) );
NOR2_X2 \AES_ENC/us11/U486  ( .A1(\AES_ENC/us11/n1056 ), .A2(\AES_ENC/us11/n1053 ), .ZN(\AES_ENC/us11/n749 ) );
NOR2_X2 \AES_ENC/us11/U483  ( .A1(\AES_ENC/us11/n749 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n752 ) );
INV_X4 \AES_ENC/us11/U482  ( .A(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n596 ));
NOR2_X2 \AES_ENC/us11/U480  ( .A1(\AES_ENC/us11/n1054 ), .A2(\AES_ENC/us11/n1053 ), .ZN(\AES_ENC/us11/n1055 ) );
OR2_X4 \AES_ENC/us11/U479  ( .A1(\AES_ENC/us11/n1094 ), .A2(\AES_ENC/us11/n1093 ), .ZN(\AES_ENC/us11/n571 ) );
AND2_X2 \AES_ENC/us11/U478  ( .A1(\AES_ENC/us11/n571 ), .A2(\AES_ENC/us11/n1095 ), .ZN(\AES_ENC/us11/n1101 ) );
NOR2_X2 \AES_ENC/us11/U477  ( .A1(\AES_ENC/us11/n1074 ), .A2(\AES_ENC/us11/n931 ), .ZN(\AES_ENC/us11/n796 ) );
NOR2_X2 \AES_ENC/us11/U474  ( .A1(\AES_ENC/us11/n796 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n797 ) );
NOR2_X2 \AES_ENC/us11/U473  ( .A1(\AES_ENC/us11/n932 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n933 ) );
NOR2_X2 \AES_ENC/us11/U472  ( .A1(\AES_ENC/us11/n929 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n935 ) );
NOR2_X2 \AES_ENC/us11/U471  ( .A1(\AES_ENC/us11/n931 ), .A2(\AES_ENC/us11/n930 ), .ZN(\AES_ENC/us11/n934 ) );
NOR3_X2 \AES_ENC/us11/U470  ( .A1(\AES_ENC/us11/n935 ), .A2(\AES_ENC/us11/n934 ), .A3(\AES_ENC/us11/n933 ), .ZN(\AES_ENC/us11/n936 ) );
NOR2_X2 \AES_ENC/us11/U469  ( .A1(\AES_ENC/us11/n624 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n1075 ) );
NOR2_X2 \AES_ENC/us11/U468  ( .A1(\AES_ENC/us11/n572 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n949 ) );
NOR2_X2 \AES_ENC/us11/U467  ( .A1(\AES_ENC/us11/n1049 ), .A2(\AES_ENC/us11/n618 ), .ZN(\AES_ENC/us11/n1051 ) );
NOR2_X2 \AES_ENC/us11/U466  ( .A1(\AES_ENC/us11/n1051 ), .A2(\AES_ENC/us11/n1050 ), .ZN(\AES_ENC/us11/n1052 ) );
NOR2_X2 \AES_ENC/us11/U465  ( .A1(\AES_ENC/us11/n1052 ), .A2(\AES_ENC/us11/n592 ), .ZN(\AES_ENC/us11/n1064 ) );
NOR2_X2 \AES_ENC/us11/U464  ( .A1(\AES_ENC/sa11 [1]), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n631 ) );
NOR2_X2 \AES_ENC/us11/U463  ( .A1(\AES_ENC/us11/n1025 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n980 ) );
NOR2_X2 \AES_ENC/us11/U462  ( .A1(\AES_ENC/us11/n1073 ), .A2(\AES_ENC/us11/n1094 ), .ZN(\AES_ENC/us11/n795 ) );
NOR2_X2 \AES_ENC/us11/U461  ( .A1(\AES_ENC/us11/n795 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n799 ) );
NOR2_X2 \AES_ENC/us11/U460  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n981 ) );
NOR2_X2 \AES_ENC/us11/U459  ( .A1(\AES_ENC/us11/n1102 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n643 ) );
NOR2_X2 \AES_ENC/us11/U458  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n621 ), .ZN(\AES_ENC/us11/n642 ) );
NOR2_X2 \AES_ENC/us11/U455  ( .A1(\AES_ENC/us11/n911 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n644 ) );
NOR4_X2 \AES_ENC/us11/U448  ( .A1(\AES_ENC/us11/n644 ), .A2(\AES_ENC/us11/n643 ), .A3(\AES_ENC/us11/n804 ), .A4(\AES_ENC/us11/n642 ), .ZN(\AES_ENC/us11/n645 ) );
NOR2_X2 \AES_ENC/us11/U447  ( .A1(\AES_ENC/us11/n1102 ), .A2(\AES_ENC/us11/n910 ), .ZN(\AES_ENC/us11/n932 ) );
NOR2_X2 \AES_ENC/us11/U442  ( .A1(\AES_ENC/us11/n1102 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n755 ) );
NOR2_X2 \AES_ENC/us11/U441  ( .A1(\AES_ENC/us11/n931 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n743 ) );
NOR2_X2 \AES_ENC/us11/U438  ( .A1(\AES_ENC/us11/n1072 ), .A2(\AES_ENC/us11/n1094 ), .ZN(\AES_ENC/us11/n930 ) );
NOR2_X2 \AES_ENC/us11/U435  ( .A1(\AES_ENC/us11/n1074 ), .A2(\AES_ENC/us11/n1025 ), .ZN(\AES_ENC/us11/n891 ) );
NOR2_X2 \AES_ENC/us11/U434  ( .A1(\AES_ENC/us11/n891 ), .A2(\AES_ENC/us11/n609 ), .ZN(\AES_ENC/us11/n894 ) );
NOR3_X2 \AES_ENC/us11/U433  ( .A1(\AES_ENC/us11/n623 ), .A2(\AES_ENC/sa11 [1]), .A3(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n683 ));
INV_X4 \AES_ENC/us11/U428  ( .A(\AES_ENC/us11/n931 ), .ZN(\AES_ENC/us11/n623 ) );
NOR2_X2 \AES_ENC/us11/U427  ( .A1(\AES_ENC/us11/n996 ), .A2(\AES_ENC/us11/n931 ), .ZN(\AES_ENC/us11/n704 ) );
NOR2_X2 \AES_ENC/us11/U421  ( .A1(\AES_ENC/us11/n931 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n685 ) );
NOR2_X2 \AES_ENC/us11/U420  ( .A1(\AES_ENC/us11/n1029 ), .A2(\AES_ENC/us11/n1025 ), .ZN(\AES_ENC/us11/n1079 ) );
NOR3_X2 \AES_ENC/us11/U419  ( .A1(\AES_ENC/us11/n589 ), .A2(\AES_ENC/us11/n1025 ), .A3(\AES_ENC/us11/n616 ), .ZN(\AES_ENC/us11/n945 ) );
NOR2_X2 \AES_ENC/us11/U418  ( .A1(\AES_ENC/us11/n626 ), .A2(\AES_ENC/us11/n611 ), .ZN(\AES_ENC/us11/n800 ) );
NOR3_X2 \AES_ENC/us11/U417  ( .A1(\AES_ENC/us11/n590 ), .A2(\AES_ENC/us11/n627 ), .A3(\AES_ENC/us11/n611 ), .ZN(\AES_ENC/us11/n798 ) );
NOR3_X2 \AES_ENC/us11/U416  ( .A1(\AES_ENC/us11/n610 ), .A2(\AES_ENC/us11/n572 ), .A3(\AES_ENC/us11/n575 ), .ZN(\AES_ENC/us11/n962 ) );
NOR3_X2 \AES_ENC/us11/U415  ( .A1(\AES_ENC/us11/n959 ), .A2(\AES_ENC/us11/n572 ), .A3(\AES_ENC/us11/n609 ), .ZN(\AES_ENC/us11/n768 ) );
NOR3_X2 \AES_ENC/us11/U414  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n572 ), .A3(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n694 ) );
NOR3_X2 \AES_ENC/us11/U413  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n572 ), .A3(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n895 ) );
NOR3_X2 \AES_ENC/us11/U410  ( .A1(\AES_ENC/us11/n1008 ), .A2(\AES_ENC/us11/n1007 ), .A3(\AES_ENC/us11/n1006 ), .ZN(\AES_ENC/us11/n1018 ) );
NOR4_X2 \AES_ENC/us11/U409  ( .A1(\AES_ENC/us11/n806 ), .A2(\AES_ENC/us11/n805 ), .A3(\AES_ENC/us11/n804 ), .A4(\AES_ENC/us11/n803 ), .ZN(\AES_ENC/us11/n807 ) );
NOR3_X2 \AES_ENC/us11/U406  ( .A1(\AES_ENC/us11/n799 ), .A2(\AES_ENC/us11/n798 ), .A3(\AES_ENC/us11/n797 ), .ZN(\AES_ENC/us11/n808 ) );
NOR4_X2 \AES_ENC/us11/U405  ( .A1(\AES_ENC/us11/n843 ), .A2(\AES_ENC/us11/n842 ), .A3(\AES_ENC/us11/n841 ), .A4(\AES_ENC/us11/n840 ), .ZN(\AES_ENC/us11/n844 ) );
NOR2_X2 \AES_ENC/us11/U404  ( .A1(\AES_ENC/us11/n669 ), .A2(\AES_ENC/us11/n668 ), .ZN(\AES_ENC/us11/n673 ) );
NOR4_X2 \AES_ENC/us11/U403  ( .A1(\AES_ENC/us11/n946 ), .A2(\AES_ENC/us11/n1046 ), .A3(\AES_ENC/us11/n671 ), .A4(\AES_ENC/us11/n670 ), .ZN(\AES_ENC/us11/n672 ) );
NOR4_X2 \AES_ENC/us11/U401  ( .A1(\AES_ENC/us11/n711 ), .A2(\AES_ENC/us11/n710 ), .A3(\AES_ENC/us11/n709 ), .A4(\AES_ENC/us11/n708 ), .ZN(\AES_ENC/us11/n712 ) );
NOR4_X2 \AES_ENC/us11/U400  ( .A1(\AES_ENC/us11/n963 ), .A2(\AES_ENC/us11/n962 ), .A3(\AES_ENC/us11/n961 ), .A4(\AES_ENC/us11/n960 ), .ZN(\AES_ENC/us11/n964 ) );
NOR3_X2 \AES_ENC/us11/U399  ( .A1(\AES_ENC/us11/n1101 ), .A2(\AES_ENC/us11/n1100 ), .A3(\AES_ENC/us11/n1099 ), .ZN(\AES_ENC/us11/n1109 ) );
NOR3_X2 \AES_ENC/us11/U398  ( .A1(\AES_ENC/us11/n743 ), .A2(\AES_ENC/us11/n742 ), .A3(\AES_ENC/us11/n741 ), .ZN(\AES_ENC/us11/n744 ) );
NOR2_X2 \AES_ENC/us11/U397  ( .A1(\AES_ENC/us11/n697 ), .A2(\AES_ENC/us11/n658 ), .ZN(\AES_ENC/us11/n659 ) );
NOR2_X2 \AES_ENC/us11/U396  ( .A1(\AES_ENC/us11/n1078 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n1033 ) );
NOR2_X2 \AES_ENC/us11/U393  ( .A1(\AES_ENC/us11/n1031 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n1032 ) );
NOR3_X2 \AES_ENC/us11/U390  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n1025 ), .A3(\AES_ENC/us11/n1074 ), .ZN(\AES_ENC/us11/n1035 ) );
NOR4_X2 \AES_ENC/us11/U389  ( .A1(\AES_ENC/us11/n1035 ), .A2(\AES_ENC/us11/n1034 ), .A3(\AES_ENC/us11/n1033 ), .A4(\AES_ENC/us11/n1032 ), .ZN(\AES_ENC/us11/n1036 ) );
NOR2_X2 \AES_ENC/us11/U388  ( .A1(\AES_ENC/us11/n598 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n885 ) );
NOR2_X2 \AES_ENC/us11/U387  ( .A1(\AES_ENC/us11/n623 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n882 ) );
NOR2_X2 \AES_ENC/us11/U386  ( .A1(\AES_ENC/us11/n1053 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n884 ) );
NOR4_X2 \AES_ENC/us11/U385  ( .A1(\AES_ENC/us11/n885 ), .A2(\AES_ENC/us11/n884 ), .A3(\AES_ENC/us11/n883 ), .A4(\AES_ENC/us11/n882 ), .ZN(\AES_ENC/us11/n886 ) );
NOR2_X2 \AES_ENC/us11/U384  ( .A1(\AES_ENC/us11/n825 ), .A2(\AES_ENC/us11/n578 ), .ZN(\AES_ENC/us11/n830 ) );
NOR2_X2 \AES_ENC/us11/U383  ( .A1(\AES_ENC/us11/n827 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n829 ) );
NOR2_X2 \AES_ENC/us11/U382  ( .A1(\AES_ENC/us11/n572 ), .A2(\AES_ENC/us11/n579 ), .ZN(\AES_ENC/us11/n828 ) );
NOR4_X2 \AES_ENC/us11/U374  ( .A1(\AES_ENC/us11/n831 ), .A2(\AES_ENC/us11/n830 ), .A3(\AES_ENC/us11/n829 ), .A4(\AES_ENC/us11/n828 ), .ZN(\AES_ENC/us11/n832 ) );
NOR2_X2 \AES_ENC/us11/U373  ( .A1(\AES_ENC/us11/n606 ), .A2(\AES_ENC/us11/n582 ), .ZN(\AES_ENC/us11/n1104 ) );
NOR2_X2 \AES_ENC/us11/U372  ( .A1(\AES_ENC/us11/n1102 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n1106 ) );
NOR2_X2 \AES_ENC/us11/U370  ( .A1(\AES_ENC/us11/n1103 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n1105 ) );
NOR4_X2 \AES_ENC/us11/U369  ( .A1(\AES_ENC/us11/n1107 ), .A2(\AES_ENC/us11/n1106 ), .A3(\AES_ENC/us11/n1105 ), .A4(\AES_ENC/us11/n1104 ), .ZN(\AES_ENC/us11/n1108 ) );
NOR3_X2 \AES_ENC/us11/U368  ( .A1(\AES_ENC/us11/n959 ), .A2(\AES_ENC/us11/n621 ), .A3(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n963 ) );
NOR2_X2 \AES_ENC/us11/U367  ( .A1(\AES_ENC/us11/n626 ), .A2(\AES_ENC/us11/n627 ), .ZN(\AES_ENC/us11/n1114 ) );
INV_X4 \AES_ENC/us11/U366  ( .A(\AES_ENC/us11/n1024 ), .ZN(\AES_ENC/us11/n606 ) );
NOR3_X2 \AES_ENC/us11/U365  ( .A1(\AES_ENC/us11/n910 ), .A2(\AES_ENC/us11/n1059 ), .A3(\AES_ENC/us11/n611 ), .ZN(\AES_ENC/us11/n1115 ) );
INV_X4 \AES_ENC/us11/U364  ( .A(\AES_ENC/us11/n1094 ), .ZN(\AES_ENC/us11/n613 ) );
NOR2_X2 \AES_ENC/us11/U363  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n931 ), .ZN(\AES_ENC/us11/n1100 ) );
INV_X4 \AES_ENC/us11/U354  ( .A(\AES_ENC/us11/n1093 ), .ZN(\AES_ENC/us11/n617 ) );
NOR2_X2 \AES_ENC/us11/U353  ( .A1(\AES_ENC/us11/n569 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n929 ) );
NOR2_X2 \AES_ENC/us11/U352  ( .A1(\AES_ENC/us11/n620 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n926 ) );
NOR2_X2 \AES_ENC/us11/U351  ( .A1(\AES_ENC/us11/n572 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n1095 ) );
NOR2_X2 \AES_ENC/us11/U350  ( .A1(\AES_ENC/us11/n609 ), .A2(\AES_ENC/us11/n627 ), .ZN(\AES_ENC/us11/n1010 ) );
NOR2_X2 \AES_ENC/us11/U349  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n1103 ) );
NOR2_X2 \AES_ENC/us11/U348  ( .A1(\AES_ENC/us11/n622 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n1059 ) );
NOR2_X2 \AES_ENC/us11/U347  ( .A1(\AES_ENC/sa11 [1]), .A2(\AES_ENC/us11/n1120 ), .ZN(\AES_ENC/us11/n1022 ) );
NOR2_X2 \AES_ENC/us11/U346  ( .A1(\AES_ENC/us11/n619 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n911 ) );
NOR2_X2 \AES_ENC/us11/U345  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/us11/n1025 ), .ZN(\AES_ENC/us11/n826 ) );
NOR2_X2 \AES_ENC/us11/U338  ( .A1(\AES_ENC/us11/n626 ), .A2(\AES_ENC/us11/n607 ), .ZN(\AES_ENC/us11/n1072 ) );
NOR2_X2 \AES_ENC/us11/U335  ( .A1(\AES_ENC/us11/n627 ), .A2(\AES_ENC/us11/n616 ), .ZN(\AES_ENC/us11/n956 ) );
NOR2_X2 \AES_ENC/us11/U329  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/us11/n624 ), .ZN(\AES_ENC/us11/n1121 ) );
NOR2_X2 \AES_ENC/us11/U328  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/us11/n624 ), .ZN(\AES_ENC/us11/n1058 ) );
NOR2_X2 \AES_ENC/us11/U327  ( .A1(\AES_ENC/us11/n625 ), .A2(\AES_ENC/us11/n611 ), .ZN(\AES_ENC/us11/n1073 ) );
NOR2_X2 \AES_ENC/us11/U325  ( .A1(\AES_ENC/sa11 [1]), .A2(\AES_ENC/us11/n1025 ), .ZN(\AES_ENC/us11/n1054 ) );
NOR2_X2 \AES_ENC/us11/U324  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/us11/n931 ), .ZN(\AES_ENC/us11/n1029 ) );
NOR2_X2 \AES_ENC/us11/U319  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n1056 ) );
NOR2_X2 \AES_ENC/us11/U318  ( .A1(\AES_ENC/us11/n614 ), .A2(\AES_ENC/us11/n626 ), .ZN(\AES_ENC/us11/n1050 ) );
NOR2_X2 \AES_ENC/us11/U317  ( .A1(\AES_ENC/us11/n1121 ), .A2(\AES_ENC/us11/n1025 ), .ZN(\AES_ENC/us11/n1120 ) );
NOR2_X2 \AES_ENC/us11/U316  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/us11/n572 ), .ZN(\AES_ENC/us11/n1074 ) );
NOR2_X2 \AES_ENC/us11/U315  ( .A1(\AES_ENC/us11/n1058 ), .A2(\AES_ENC/us11/n1054 ), .ZN(\AES_ENC/us11/n878 ) );
NOR2_X2 \AES_ENC/us11/U314  ( .A1(\AES_ENC/us11/n878 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n879 ) );
NOR2_X2 \AES_ENC/us11/U312  ( .A1(\AES_ENC/us11/n880 ), .A2(\AES_ENC/us11/n879 ), .ZN(\AES_ENC/us11/n887 ) );
NOR2_X2 \AES_ENC/us11/U311  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n588 ), .ZN(\AES_ENC/us11/n957 ) );
NOR2_X2 \AES_ENC/us11/U310  ( .A1(\AES_ENC/us11/n958 ), .A2(\AES_ENC/us11/n957 ), .ZN(\AES_ENC/us11/n965 ) );
NOR3_X2 \AES_ENC/us11/U309  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n1091 ), .A3(\AES_ENC/us11/n1022 ), .ZN(\AES_ENC/us11/n720 ) );
NOR3_X2 \AES_ENC/us11/U303  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n1054 ), .A3(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n719 ) );
NOR2_X2 \AES_ENC/us11/U302  ( .A1(\AES_ENC/us11/n720 ), .A2(\AES_ENC/us11/n719 ), .ZN(\AES_ENC/us11/n726 ) );
NOR2_X2 \AES_ENC/us11/U300  ( .A1(\AES_ENC/us11/n614 ), .A2(\AES_ENC/us11/n591 ), .ZN(\AES_ENC/us11/n865 ) );
NOR2_X2 \AES_ENC/us11/U299  ( .A1(\AES_ENC/us11/n1059 ), .A2(\AES_ENC/us11/n1058 ), .ZN(\AES_ENC/us11/n1060 ) );
NOR2_X2 \AES_ENC/us11/U298  ( .A1(\AES_ENC/us11/n1095 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n668 ) );
NOR2_X2 \AES_ENC/us11/U297  ( .A1(\AES_ENC/us11/n911 ), .A2(\AES_ENC/us11/n910 ), .ZN(\AES_ENC/us11/n912 ) );
NOR2_X2 \AES_ENC/us11/U296  ( .A1(\AES_ENC/us11/n912 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n916 ) );
NOR2_X2 \AES_ENC/us11/U295  ( .A1(\AES_ENC/us11/n826 ), .A2(\AES_ENC/us11/n573 ), .ZN(\AES_ENC/us11/n750 ) );
NOR2_X2 \AES_ENC/us11/U294  ( .A1(\AES_ENC/us11/n750 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n751 ) );
NOR2_X2 \AES_ENC/us11/U293  ( .A1(\AES_ENC/us11/n907 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n908 ) );
NOR2_X2 \AES_ENC/us11/U292  ( .A1(\AES_ENC/us11/n990 ), .A2(\AES_ENC/us11/n926 ), .ZN(\AES_ENC/us11/n780 ) );
NOR2_X2 \AES_ENC/us11/U291  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n584 ), .ZN(\AES_ENC/us11/n838 ) );
NOR2_X2 \AES_ENC/us11/U290  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n602 ), .ZN(\AES_ENC/us11/n837 ) );
NOR2_X2 \AES_ENC/us11/U284  ( .A1(\AES_ENC/us11/n838 ), .A2(\AES_ENC/us11/n837 ), .ZN(\AES_ENC/us11/n845 ) );
NOR2_X2 \AES_ENC/us11/U283  ( .A1(\AES_ENC/us11/n1022 ), .A2(\AES_ENC/us11/n1058 ), .ZN(\AES_ENC/us11/n740 ) );
NOR2_X2 \AES_ENC/us11/U282  ( .A1(\AES_ENC/us11/n740 ), .A2(\AES_ENC/us11/n616 ), .ZN(\AES_ENC/us11/n742 ) );
NOR2_X2 \AES_ENC/us11/U281  ( .A1(\AES_ENC/us11/n1098 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n1099 ) );
NOR2_X2 \AES_ENC/us11/U280  ( .A1(\AES_ENC/us11/n1120 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n993 ) );
NOR2_X2 \AES_ENC/us11/U279  ( .A1(\AES_ENC/us11/n993 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n994 ) );
NOR2_X2 \AES_ENC/us11/U273  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n620 ), .ZN(\AES_ENC/us11/n1026 ) );
NOR2_X2 \AES_ENC/us11/U272  ( .A1(\AES_ENC/us11/n573 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n1027 ) );
NOR2_X2 \AES_ENC/us11/U271  ( .A1(\AES_ENC/us11/n1027 ), .A2(\AES_ENC/us11/n1026 ), .ZN(\AES_ENC/us11/n1028 ) );
NOR2_X2 \AES_ENC/us11/U270  ( .A1(\AES_ENC/us11/n1029 ), .A2(\AES_ENC/us11/n1028 ), .ZN(\AES_ENC/us11/n1034 ) );
NOR4_X2 \AES_ENC/us11/U269  ( .A1(\AES_ENC/us11/n757 ), .A2(\AES_ENC/us11/n756 ), .A3(\AES_ENC/us11/n755 ), .A4(\AES_ENC/us11/n754 ), .ZN(\AES_ENC/us11/n758 ) );
NOR2_X2 \AES_ENC/us11/U268  ( .A1(\AES_ENC/us11/n752 ), .A2(\AES_ENC/us11/n751 ), .ZN(\AES_ENC/us11/n759 ) );
NOR2_X2 \AES_ENC/us11/U267  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n1071 ), .ZN(\AES_ENC/us11/n669 ) );
NOR2_X2 \AES_ENC/us11/U263  ( .A1(\AES_ENC/us11/n1056 ), .A2(\AES_ENC/us11/n990 ), .ZN(\AES_ENC/us11/n991 ) );
NOR2_X2 \AES_ENC/us11/U262  ( .A1(\AES_ENC/us11/n991 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n995 ) );
NOR2_X2 \AES_ENC/us11/U258  ( .A1(\AES_ENC/us11/n607 ), .A2(\AES_ENC/us11/n590 ), .ZN(\AES_ENC/us11/n1008 ) );
NOR2_X2 \AES_ENC/us11/U255  ( .A1(\AES_ENC/us11/n839 ), .A2(\AES_ENC/us11/n582 ), .ZN(\AES_ENC/us11/n693 ) );
NOR2_X2 \AES_ENC/us11/U254  ( .A1(\AES_ENC/us11/n606 ), .A2(\AES_ENC/us11/n906 ), .ZN(\AES_ENC/us11/n741 ) );
NOR2_X2 \AES_ENC/us11/U253  ( .A1(\AES_ENC/us11/n1054 ), .A2(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n763 ) );
NOR2_X2 \AES_ENC/us11/U252  ( .A1(\AES_ENC/us11/n763 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n769 ) );
NOR2_X2 \AES_ENC/us11/U251  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n577 ), .ZN(\AES_ENC/us11/n1007 ) );
NOR2_X2 \AES_ENC/us11/U250  ( .A1(\AES_ENC/us11/n609 ), .A2(\AES_ENC/us11/n580 ), .ZN(\AES_ENC/us11/n1123 ) );
NOR2_X2 \AES_ENC/us11/U243  ( .A1(\AES_ENC/us11/n609 ), .A2(\AES_ENC/us11/n590 ), .ZN(\AES_ENC/us11/n710 ) );
INV_X4 \AES_ENC/us11/U242  ( .A(\AES_ENC/us11/n1029 ), .ZN(\AES_ENC/us11/n582 ) );
NOR2_X2 \AES_ENC/us11/U241  ( .A1(\AES_ENC/us11/n616 ), .A2(\AES_ENC/us11/n597 ), .ZN(\AES_ENC/us11/n883 ) );
NOR2_X2 \AES_ENC/us11/U240  ( .A1(\AES_ENC/us11/n593 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n1125 ) );
NOR2_X2 \AES_ENC/us11/U239  ( .A1(\AES_ENC/us11/n990 ), .A2(\AES_ENC/us11/n929 ), .ZN(\AES_ENC/us11/n892 ) );
NOR2_X2 \AES_ENC/us11/U238  ( .A1(\AES_ENC/us11/n892 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n893 ) );
NOR2_X2 \AES_ENC/us11/U237  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n602 ), .ZN(\AES_ENC/us11/n950 ) );
NOR2_X2 \AES_ENC/us11/U236  ( .A1(\AES_ENC/us11/n1079 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n1082 ) );
NOR2_X2 \AES_ENC/us11/U235  ( .A1(\AES_ENC/us11/n910 ), .A2(\AES_ENC/us11/n1056 ), .ZN(\AES_ENC/us11/n941 ) );
NOR2_X2 \AES_ENC/us11/U234  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n1077 ), .ZN(\AES_ENC/us11/n841 ) );
NOR2_X2 \AES_ENC/us11/U229  ( .A1(\AES_ENC/us11/n623 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n630 ) );
NOR2_X2 \AES_ENC/us11/U228  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n602 ), .ZN(\AES_ENC/us11/n806 ) );
NOR2_X2 \AES_ENC/us11/U227  ( .A1(\AES_ENC/us11/n623 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n948 ) );
NOR2_X2 \AES_ENC/us11/U226  ( .A1(\AES_ENC/us11/n606 ), .A2(\AES_ENC/us11/n589 ), .ZN(\AES_ENC/us11/n997 ) );
NOR2_X2 \AES_ENC/us11/U225  ( .A1(\AES_ENC/us11/n1121 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n1122 ) );
NOR2_X2 \AES_ENC/us11/U223  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n1023 ), .ZN(\AES_ENC/us11/n756 ) );
NOR2_X2 \AES_ENC/us11/U222  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n602 ), .ZN(\AES_ENC/us11/n870 ) );
NOR2_X2 \AES_ENC/us11/U221  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n569 ), .ZN(\AES_ENC/us11/n947 ) );
NOR2_X2 \AES_ENC/us11/U217  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n1077 ), .ZN(\AES_ENC/us11/n1084 ) );
NOR2_X2 \AES_ENC/us11/U213  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n855 ), .ZN(\AES_ENC/us11/n709 ) );
NOR2_X2 \AES_ENC/us11/U212  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n589 ), .ZN(\AES_ENC/us11/n868 ) );
NOR2_X2 \AES_ENC/us11/U211  ( .A1(\AES_ENC/us11/n1120 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n1124 ) );
NOR2_X2 \AES_ENC/us11/U210  ( .A1(\AES_ENC/us11/n1120 ), .A2(\AES_ENC/us11/n839 ), .ZN(\AES_ENC/us11/n842 ) );
NOR2_X2 \AES_ENC/us11/U209  ( .A1(\AES_ENC/us11/n1120 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n696 ) );
NOR2_X2 \AES_ENC/us11/U208  ( .A1(\AES_ENC/us11/n1074 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n1076 ) );
NOR2_X2 \AES_ENC/us11/U207  ( .A1(\AES_ENC/us11/n1074 ), .A2(\AES_ENC/us11/n620 ), .ZN(\AES_ENC/us11/n781 ) );
NOR3_X2 \AES_ENC/us11/U201  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n1056 ), .A3(\AES_ENC/us11/n990 ), .ZN(\AES_ENC/us11/n979 ) );
NOR3_X2 \AES_ENC/us11/U200  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n1058 ), .A3(\AES_ENC/us11/n1059 ), .ZN(\AES_ENC/us11/n854 ) );
NOR2_X2 \AES_ENC/us11/U199  ( .A1(\AES_ENC/us11/n996 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n869 ) );
NOR2_X2 \AES_ENC/us11/U198  ( .A1(\AES_ENC/us11/n1056 ), .A2(\AES_ENC/us11/n1074 ), .ZN(\AES_ENC/us11/n1057 ) );
NOR3_X2 \AES_ENC/us11/U197  ( .A1(\AES_ENC/us11/n607 ), .A2(\AES_ENC/us11/n1120 ), .A3(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n978 ) );
NOR2_X2 \AES_ENC/us11/U196  ( .A1(\AES_ENC/us11/n996 ), .A2(\AES_ENC/us11/n911 ), .ZN(\AES_ENC/us11/n1116 ) );
NOR2_X2 \AES_ENC/us11/U195  ( .A1(\AES_ENC/us11/n1074 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n754 ) );
NOR2_X2 \AES_ENC/us11/U194  ( .A1(\AES_ENC/us11/n926 ), .A2(\AES_ENC/us11/n1103 ), .ZN(\AES_ENC/us11/n977 ) );
NOR2_X2 \AES_ENC/us11/U187  ( .A1(\AES_ENC/us11/n839 ), .A2(\AES_ENC/us11/n824 ), .ZN(\AES_ENC/us11/n1092 ) );
NOR2_X2 \AES_ENC/us11/U186  ( .A1(\AES_ENC/us11/n573 ), .A2(\AES_ENC/us11/n1074 ), .ZN(\AES_ENC/us11/n684 ) );
NOR2_X2 \AES_ENC/us11/U185  ( .A1(\AES_ENC/us11/n826 ), .A2(\AES_ENC/us11/n1059 ), .ZN(\AES_ENC/us11/n907 ) );
NOR3_X2 \AES_ENC/us11/U184  ( .A1(\AES_ENC/us11/n625 ), .A2(\AES_ENC/us11/n1115 ), .A3(\AES_ENC/us11/n585 ), .ZN(\AES_ENC/us11/n831 ) );
NOR3_X2 \AES_ENC/us11/U183  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n1056 ), .A3(\AES_ENC/us11/n990 ), .ZN(\AES_ENC/us11/n896 ) );
NOR3_X2 \AES_ENC/us11/U182  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n573 ), .A3(\AES_ENC/us11/n1013 ), .ZN(\AES_ENC/us11/n670 ) );
NOR3_X2 \AES_ENC/us11/U181  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n1091 ), .A3(\AES_ENC/us11/n1022 ), .ZN(\AES_ENC/us11/n843 ) );
NOR2_X2 \AES_ENC/us11/U180  ( .A1(\AES_ENC/us11/n1029 ), .A2(\AES_ENC/us11/n1095 ), .ZN(\AES_ENC/us11/n735 ) );
NOR2_X2 \AES_ENC/us11/U174  ( .A1(\AES_ENC/us11/n1100 ), .A2(\AES_ENC/us11/n854 ), .ZN(\AES_ENC/us11/n860 ) );
NAND3_X2 \AES_ENC/us11/U173  ( .A1(\AES_ENC/us11/n569 ), .A2(\AES_ENC/us11/n582 ), .A3(\AES_ENC/us11/n681 ), .ZN(\AES_ENC/us11/n691 ) );
NOR2_X2 \AES_ENC/us11/U172  ( .A1(\AES_ENC/us11/n683 ), .A2(\AES_ENC/us11/n682 ), .ZN(\AES_ENC/us11/n690 ) );
NOR3_X2 \AES_ENC/us11/U171  ( .A1(\AES_ENC/us11/n695 ), .A2(\AES_ENC/us11/n694 ), .A3(\AES_ENC/us11/n693 ), .ZN(\AES_ENC/us11/n700 ) );
NOR4_X2 \AES_ENC/us11/U170  ( .A1(\AES_ENC/us11/n983 ), .A2(\AES_ENC/us11/n698 ), .A3(\AES_ENC/us11/n697 ), .A4(\AES_ENC/us11/n696 ), .ZN(\AES_ENC/us11/n699 ) );
NOR2_X2 \AES_ENC/us11/U169  ( .A1(\AES_ENC/us11/n946 ), .A2(\AES_ENC/us11/n945 ), .ZN(\AES_ENC/us11/n952 ) );
NOR4_X2 \AES_ENC/us11/U168  ( .A1(\AES_ENC/us11/n950 ), .A2(\AES_ENC/us11/n949 ), .A3(\AES_ENC/us11/n948 ), .A4(\AES_ENC/us11/n947 ), .ZN(\AES_ENC/us11/n951 ) );
NOR4_X2 \AES_ENC/us11/U162  ( .A1(\AES_ENC/us11/n896 ), .A2(\AES_ENC/us11/n895 ), .A3(\AES_ENC/us11/n894 ), .A4(\AES_ENC/us11/n893 ), .ZN(\AES_ENC/us11/n897 ) );
NOR2_X2 \AES_ENC/us11/U161  ( .A1(\AES_ENC/us11/n866 ), .A2(\AES_ENC/us11/n865 ), .ZN(\AES_ENC/us11/n872 ) );
NOR4_X2 \AES_ENC/us11/U160  ( .A1(\AES_ENC/us11/n870 ), .A2(\AES_ENC/us11/n869 ), .A3(\AES_ENC/us11/n868 ), .A4(\AES_ENC/us11/n867 ), .ZN(\AES_ENC/us11/n871 ) );
NOR4_X2 \AES_ENC/us11/U159  ( .A1(\AES_ENC/us11/n983 ), .A2(\AES_ENC/us11/n982 ), .A3(\AES_ENC/us11/n981 ), .A4(\AES_ENC/us11/n980 ), .ZN(\AES_ENC/us11/n984 ) );
NOR2_X2 \AES_ENC/us11/U158  ( .A1(\AES_ENC/us11/n979 ), .A2(\AES_ENC/us11/n978 ), .ZN(\AES_ENC/us11/n985 ) );
NOR4_X2 \AES_ENC/us11/U157  ( .A1(\AES_ENC/us11/n1125 ), .A2(\AES_ENC/us11/n1124 ), .A3(\AES_ENC/us11/n1123 ), .A4(\AES_ENC/us11/n1122 ), .ZN(\AES_ENC/us11/n1126 ) );
NOR4_X2 \AES_ENC/us11/U156  ( .A1(\AES_ENC/us11/n1084 ), .A2(\AES_ENC/us11/n1083 ), .A3(\AES_ENC/us11/n1082 ), .A4(\AES_ENC/us11/n1081 ), .ZN(\AES_ENC/us11/n1085 ) );
NOR2_X2 \AES_ENC/us11/U155  ( .A1(\AES_ENC/us11/n1076 ), .A2(\AES_ENC/us11/n1075 ), .ZN(\AES_ENC/us11/n1086 ) );
NOR3_X2 \AES_ENC/us11/U154  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n1054 ), .A3(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n961 ) );
NOR3_X2 \AES_ENC/us11/U153  ( .A1(\AES_ENC/us11/n620 ), .A2(\AES_ENC/us11/n1074 ), .A3(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n671 ) );
NOR2_X2 \AES_ENC/us11/U152  ( .A1(\AES_ENC/us11/n1057 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n1062 ) );
NOR2_X2 \AES_ENC/us11/U143  ( .A1(\AES_ENC/us11/n1055 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n1063 ) );
NOR2_X2 \AES_ENC/us11/U142  ( .A1(\AES_ENC/us11/n1060 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n1061 ) );
NOR4_X2 \AES_ENC/us11/U141  ( .A1(\AES_ENC/us11/n1064 ), .A2(\AES_ENC/us11/n1063 ), .A3(\AES_ENC/us11/n1062 ), .A4(\AES_ENC/us11/n1061 ), .ZN(\AES_ENC/us11/n1065 ) );
NOR3_X2 \AES_ENC/us11/U140  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n1120 ), .A3(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n918 ) );
NOR3_X2 \AES_ENC/us11/U132  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n573 ), .A3(\AES_ENC/us11/n1013 ), .ZN(\AES_ENC/us11/n917 ) );
NOR2_X2 \AES_ENC/us11/U131  ( .A1(\AES_ENC/us11/n914 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n915 ) );
NOR4_X2 \AES_ENC/us11/U130  ( .A1(\AES_ENC/us11/n918 ), .A2(\AES_ENC/us11/n917 ), .A3(\AES_ENC/us11/n916 ), .A4(\AES_ENC/us11/n915 ), .ZN(\AES_ENC/us11/n919 ) );
NOR2_X2 \AES_ENC/us11/U129  ( .A1(\AES_ENC/us11/n735 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n687 ) );
NOR2_X2 \AES_ENC/us11/U128  ( .A1(\AES_ENC/us11/n684 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n688 ) );
NOR2_X2 \AES_ENC/us11/U127  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n600 ), .ZN(\AES_ENC/us11/n686 ) );
NOR4_X2 \AES_ENC/us11/U126  ( .A1(\AES_ENC/us11/n688 ), .A2(\AES_ENC/us11/n687 ), .A3(\AES_ENC/us11/n686 ), .A4(\AES_ENC/us11/n685 ), .ZN(\AES_ENC/us11/n689 ) );
NOR2_X2 \AES_ENC/us11/U121  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n595 ), .ZN(\AES_ENC/us11/n858 ) );
NOR2_X2 \AES_ENC/us11/U120  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n855 ), .ZN(\AES_ENC/us11/n857 ) );
NOR2_X2 \AES_ENC/us11/U119  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n587 ), .ZN(\AES_ENC/us11/n856 ) );
NOR4_X2 \AES_ENC/us11/U118  ( .A1(\AES_ENC/us11/n858 ), .A2(\AES_ENC/us11/n857 ), .A3(\AES_ENC/us11/n856 ), .A4(\AES_ENC/us11/n958 ), .ZN(\AES_ENC/us11/n859 ) );
NOR2_X2 \AES_ENC/us11/U117  ( .A1(\AES_ENC/us11/n616 ), .A2(\AES_ENC/us11/n580 ), .ZN(\AES_ENC/us11/n771 ) );
NOR2_X2 \AES_ENC/us11/U116  ( .A1(\AES_ENC/us11/n1103 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n772 ) );
NOR2_X2 \AES_ENC/us11/U115  ( .A1(\AES_ENC/us11/n610 ), .A2(\AES_ENC/us11/n599 ), .ZN(\AES_ENC/us11/n773 ) );
NOR4_X2 \AES_ENC/us11/U106  ( .A1(\AES_ENC/us11/n773 ), .A2(\AES_ENC/us11/n772 ), .A3(\AES_ENC/us11/n771 ), .A4(\AES_ENC/us11/n770 ), .ZN(\AES_ENC/us11/n774 ) );
NOR2_X2 \AES_ENC/us11/U105  ( .A1(\AES_ENC/us11/n780 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n784 ) );
NOR2_X2 \AES_ENC/us11/U104  ( .A1(\AES_ENC/us11/n1117 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n782 ) );
NOR2_X2 \AES_ENC/us11/U103  ( .A1(\AES_ENC/us11/n781 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n783 ) );
NOR4_X2 \AES_ENC/us11/U102  ( .A1(\AES_ENC/us11/n880 ), .A2(\AES_ENC/us11/n784 ), .A3(\AES_ENC/us11/n783 ), .A4(\AES_ENC/us11/n782 ), .ZN(\AES_ENC/us11/n785 ) );
NOR2_X2 \AES_ENC/us11/U101  ( .A1(\AES_ENC/us11/n583 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n814 ) );
NOR2_X2 \AES_ENC/us11/U100  ( .A1(\AES_ENC/us11/n907 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n813 ) );
NOR3_X2 \AES_ENC/us11/U95  ( .A1(\AES_ENC/us11/n606 ), .A2(\AES_ENC/us11/n1058 ), .A3(\AES_ENC/us11/n1059 ), .ZN(\AES_ENC/us11/n815 ) );
NOR4_X2 \AES_ENC/us11/U94  ( .A1(\AES_ENC/us11/n815 ), .A2(\AES_ENC/us11/n814 ), .A3(\AES_ENC/us11/n813 ), .A4(\AES_ENC/us11/n812 ), .ZN(\AES_ENC/us11/n816 ) );
NOR2_X2 \AES_ENC/us11/U93  ( .A1(\AES_ENC/us11/n617 ), .A2(\AES_ENC/us11/n569 ), .ZN(\AES_ENC/us11/n721 ) );
NOR2_X2 \AES_ENC/us11/U92  ( .A1(\AES_ENC/us11/n1031 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n723 ) );
NOR2_X2 \AES_ENC/us11/U91  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n1096 ), .ZN(\AES_ENC/us11/n722 ) );
NOR4_X2 \AES_ENC/us11/U90  ( .A1(\AES_ENC/us11/n724 ), .A2(\AES_ENC/us11/n723 ), .A3(\AES_ENC/us11/n722 ), .A4(\AES_ENC/us11/n721 ), .ZN(\AES_ENC/us11/n725 ) );
NOR2_X2 \AES_ENC/us11/U89  ( .A1(\AES_ENC/us11/n911 ), .A2(\AES_ENC/us11/n990 ), .ZN(\AES_ENC/us11/n1009 ) );
NOR2_X2 \AES_ENC/us11/U88  ( .A1(\AES_ENC/us11/n1013 ), .A2(\AES_ENC/us11/n573 ), .ZN(\AES_ENC/us11/n1014 ) );
NOR2_X2 \AES_ENC/us11/U87  ( .A1(\AES_ENC/us11/n1014 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n1015 ) );
NOR4_X2 \AES_ENC/us11/U86  ( .A1(\AES_ENC/us11/n1016 ), .A2(\AES_ENC/us11/n1015 ), .A3(\AES_ENC/us11/n1119 ), .A4(\AES_ENC/us11/n1046 ), .ZN(\AES_ENC/us11/n1017 ) );
NOR2_X2 \AES_ENC/us11/U81  ( .A1(\AES_ENC/us11/n996 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n998 ) );
NOR2_X2 \AES_ENC/us11/U80  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n577 ), .ZN(\AES_ENC/us11/n1000 ) );
NOR2_X2 \AES_ENC/us11/U79  ( .A1(\AES_ENC/us11/n616 ), .A2(\AES_ENC/us11/n1096 ), .ZN(\AES_ENC/us11/n999 ) );
NOR4_X2 \AES_ENC/us11/U78  ( .A1(\AES_ENC/us11/n1000 ), .A2(\AES_ENC/us11/n999 ), .A3(\AES_ENC/us11/n998 ), .A4(\AES_ENC/us11/n997 ), .ZN(\AES_ENC/us11/n1001 ) );
NOR2_X2 \AES_ENC/us11/U74  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n1096 ), .ZN(\AES_ENC/us11/n697 ) );
NOR2_X2 \AES_ENC/us11/U73  ( .A1(\AES_ENC/us11/n620 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n958 ) );
NOR2_X2 \AES_ENC/us11/U72  ( .A1(\AES_ENC/us11/n911 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n983 ) );
NOR2_X2 \AES_ENC/us11/U71  ( .A1(\AES_ENC/us11/n1054 ), .A2(\AES_ENC/us11/n1103 ), .ZN(\AES_ENC/us11/n1031 ) );
INV_X4 \AES_ENC/us11/U65  ( .A(\AES_ENC/us11/n1050 ), .ZN(\AES_ENC/us11/n612 ) );
INV_X4 \AES_ENC/us11/U64  ( .A(\AES_ENC/us11/n1072 ), .ZN(\AES_ENC/us11/n605 ) );
INV_X4 \AES_ENC/us11/U63  ( .A(\AES_ENC/us11/n1073 ), .ZN(\AES_ENC/us11/n604 ) );
NOR2_X2 \AES_ENC/us11/U62  ( .A1(\AES_ENC/us11/n582 ), .A2(\AES_ENC/us11/n613 ), .ZN(\AES_ENC/us11/n880 ) );
NOR3_X2 \AES_ENC/us11/U61  ( .A1(\AES_ENC/us11/n826 ), .A2(\AES_ENC/us11/n1121 ), .A3(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n946 ) );
INV_X4 \AES_ENC/us11/U59  ( .A(\AES_ENC/us11/n1010 ), .ZN(\AES_ENC/us11/n608 ) );
NOR3_X2 \AES_ENC/us11/U58  ( .A1(\AES_ENC/us11/n573 ), .A2(\AES_ENC/us11/n1029 ), .A3(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n1119 ) );
INV_X4 \AES_ENC/us11/U57  ( .A(\AES_ENC/us11/n956 ), .ZN(\AES_ENC/us11/n615 ) );
NOR2_X2 \AES_ENC/us11/U50  ( .A1(\AES_ENC/us11/n623 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n1013 ) );
NOR2_X2 \AES_ENC/us11/U49  ( .A1(\AES_ENC/us11/n620 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n910 ) );
NOR2_X2 \AES_ENC/us11/U48  ( .A1(\AES_ENC/us11/n569 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n1091 ) );
NOR2_X2 \AES_ENC/us11/U47  ( .A1(\AES_ENC/us11/n622 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n990 ) );
NOR2_X2 \AES_ENC/us11/U46  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/us11/n1121 ), .ZN(\AES_ENC/us11/n996 ) );
NOR2_X2 \AES_ENC/us11/U45  ( .A1(\AES_ENC/us11/n610 ), .A2(\AES_ENC/us11/n600 ), .ZN(\AES_ENC/us11/n628 ) );
NOR2_X2 \AES_ENC/us11/U44  ( .A1(\AES_ENC/us11/n576 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n866 ) );
NOR2_X2 \AES_ENC/us11/U43  ( .A1(\AES_ENC/us11/n603 ), .A2(\AES_ENC/us11/n610 ), .ZN(\AES_ENC/us11/n1006 ) );
NOR2_X2 \AES_ENC/us11/U42  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n1117 ), .ZN(\AES_ENC/us11/n1118 ) );
NOR2_X2 \AES_ENC/us11/U41  ( .A1(\AES_ENC/us11/n1119 ), .A2(\AES_ENC/us11/n1118 ), .ZN(\AES_ENC/us11/n1127 ) );
NOR2_X2 \AES_ENC/us11/U36  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n594 ), .ZN(\AES_ENC/us11/n629 ) );
NOR2_X2 \AES_ENC/us11/U35  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n906 ), .ZN(\AES_ENC/us11/n909 ) );
NOR2_X2 \AES_ENC/us11/U34  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n597 ), .ZN(\AES_ENC/us11/n658 ) );
NOR2_X2 \AES_ENC/us11/U33  ( .A1(\AES_ENC/us11/n1116 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n695 ) );
NOR2_X2 \AES_ENC/us11/U32  ( .A1(\AES_ENC/us11/n1078 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n1083 ) );
NOR2_X2 \AES_ENC/us11/U31  ( .A1(\AES_ENC/us11/n941 ), .A2(\AES_ENC/us11/n608 ), .ZN(\AES_ENC/us11/n724 ) );
NOR2_X2 \AES_ENC/us11/U30  ( .A1(\AES_ENC/us11/n598 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n1107 ) );
NOR2_X2 \AES_ENC/us11/U29  ( .A1(\AES_ENC/us11/n576 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n840 ) );
NOR2_X2 \AES_ENC/us11/U24  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n593 ), .ZN(\AES_ENC/us11/n633 ) );
NOR2_X2 \AES_ENC/us11/U23  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n1080 ), .ZN(\AES_ENC/us11/n1081 ) );
NOR2_X2 \AES_ENC/us11/U21  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n1045 ), .ZN(\AES_ENC/us11/n812 ) );
NOR2_X2 \AES_ENC/us11/U20  ( .A1(\AES_ENC/us11/n1009 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n960 ) );
NOR2_X2 \AES_ENC/us11/U19  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n601 ), .ZN(\AES_ENC/us11/n982 ) );
NOR2_X2 \AES_ENC/us11/U18  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n594 ), .ZN(\AES_ENC/us11/n757 ) );
NOR2_X2 \AES_ENC/us11/U17  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n590 ), .ZN(\AES_ENC/us11/n698 ) );
NOR2_X2 \AES_ENC/us11/U16  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n619 ), .ZN(\AES_ENC/us11/n708 ) );
NOR2_X2 \AES_ENC/us11/U15  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n582 ), .ZN(\AES_ENC/us11/n770 ) );
NOR2_X2 \AES_ENC/us11/U10  ( .A1(\AES_ENC/us11/n619 ), .A2(\AES_ENC/us11/n604 ), .ZN(\AES_ENC/us11/n803 ) );
NOR2_X2 \AES_ENC/us11/U9  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n881 ), .ZN(\AES_ENC/us11/n711 ) );
NOR2_X2 \AES_ENC/us11/U8  ( .A1(\AES_ENC/us11/n615 ), .A2(\AES_ENC/us11/n582 ), .ZN(\AES_ENC/us11/n867 ) );
NOR2_X2 \AES_ENC/us11/U7  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n599 ), .ZN(\AES_ENC/us11/n804 ) );
NOR2_X2 \AES_ENC/us11/U6  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n620 ), .ZN(\AES_ENC/us11/n1046 ) );
OR2_X4 \AES_ENC/us11/U5  ( .A1(\AES_ENC/us11/n624 ), .A2(\AES_ENC/sa11 [1]),.ZN(\AES_ENC/us11/n570 ) );
OR2_X4 \AES_ENC/us11/U4  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/sa11 [4]),.ZN(\AES_ENC/us11/n569 ) );
NAND2_X2 \AES_ENC/us11/U514  ( .A1(\AES_ENC/us11/n1121 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n1030 ) );
AND2_X2 \AES_ENC/us11/U513  ( .A1(\AES_ENC/us11/n597 ), .A2(\AES_ENC/us11/n1030 ), .ZN(\AES_ENC/us11/n1049 ) );
NAND2_X2 \AES_ENC/us11/U511  ( .A1(\AES_ENC/us11/n1049 ), .A2(\AES_ENC/us11/n794 ), .ZN(\AES_ENC/us11/n637 ) );
AND2_X2 \AES_ENC/us11/U493  ( .A1(\AES_ENC/us11/n779 ), .A2(\AES_ENC/us11/n996 ), .ZN(\AES_ENC/us11/n632 ) );
NAND4_X2 \AES_ENC/us11/U485  ( .A1(\AES_ENC/us11/n637 ), .A2(\AES_ENC/us11/n636 ), .A3(\AES_ENC/us11/n635 ), .A4(\AES_ENC/us11/n634 ), .ZN(\AES_ENC/us11/n638 ) );
NAND2_X2 \AES_ENC/us11/U484  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n638 ), .ZN(\AES_ENC/us11/n679 ) );
NAND2_X2 \AES_ENC/us11/U481  ( .A1(\AES_ENC/us11/n1094 ), .A2(\AES_ENC/us11/n591 ), .ZN(\AES_ENC/us11/n648 ) );
NAND2_X2 \AES_ENC/us11/U476  ( .A1(\AES_ENC/us11/n601 ), .A2(\AES_ENC/us11/n590 ), .ZN(\AES_ENC/us11/n762 ) );
NAND2_X2 \AES_ENC/us11/U475  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n762 ), .ZN(\AES_ENC/us11/n647 ) );
NAND4_X2 \AES_ENC/us11/U457  ( .A1(\AES_ENC/us11/n648 ), .A2(\AES_ENC/us11/n647 ), .A3(\AES_ENC/us11/n646 ), .A4(\AES_ENC/us11/n645 ), .ZN(\AES_ENC/us11/n649 ) );
NAND2_X2 \AES_ENC/us11/U456  ( .A1(\AES_ENC/sa11 [0]), .A2(\AES_ENC/us11/n649 ), .ZN(\AES_ENC/us11/n665 ) );
NAND2_X2 \AES_ENC/us11/U454  ( .A1(\AES_ENC/us11/n596 ), .A2(\AES_ENC/us11/n623 ), .ZN(\AES_ENC/us11/n855 ) );
NAND2_X2 \AES_ENC/us11/U453  ( .A1(\AES_ENC/us11/n587 ), .A2(\AES_ENC/us11/n855 ), .ZN(\AES_ENC/us11/n821 ) );
NAND2_X2 \AES_ENC/us11/U452  ( .A1(\AES_ENC/us11/n1093 ), .A2(\AES_ENC/us11/n821 ), .ZN(\AES_ENC/us11/n662 ) );
NAND2_X2 \AES_ENC/us11/U451  ( .A1(\AES_ENC/us11/n619 ), .A2(\AES_ENC/us11/n589 ), .ZN(\AES_ENC/us11/n650 ) );
NAND2_X2 \AES_ENC/us11/U450  ( .A1(\AES_ENC/us11/n956 ), .A2(\AES_ENC/us11/n650 ), .ZN(\AES_ENC/us11/n661 ) );
NAND2_X2 \AES_ENC/us11/U449  ( .A1(\AES_ENC/us11/n626 ), .A2(\AES_ENC/us11/n627 ), .ZN(\AES_ENC/us11/n839 ) );
OR2_X2 \AES_ENC/us11/U446  ( .A1(\AES_ENC/us11/n839 ), .A2(\AES_ENC/us11/n932 ), .ZN(\AES_ENC/us11/n656 ) );
NAND2_X2 \AES_ENC/us11/U445  ( .A1(\AES_ENC/us11/n621 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n1096 ) );
NAND2_X2 \AES_ENC/us11/U444  ( .A1(\AES_ENC/us11/n1030 ), .A2(\AES_ENC/us11/n1096 ), .ZN(\AES_ENC/us11/n651 ) );
NAND2_X2 \AES_ENC/us11/U443  ( .A1(\AES_ENC/us11/n1114 ), .A2(\AES_ENC/us11/n651 ), .ZN(\AES_ENC/us11/n655 ) );
OR3_X2 \AES_ENC/us11/U440  ( .A1(\AES_ENC/us11/n1079 ), .A2(\AES_ENC/sa11 [7]), .A3(\AES_ENC/us11/n626 ), .ZN(\AES_ENC/us11/n654 ));
NAND2_X2 \AES_ENC/us11/U439  ( .A1(\AES_ENC/us11/n593 ), .A2(\AES_ENC/us11/n601 ), .ZN(\AES_ENC/us11/n652 ) );
NAND4_X2 \AES_ENC/us11/U437  ( .A1(\AES_ENC/us11/n656 ), .A2(\AES_ENC/us11/n655 ), .A3(\AES_ENC/us11/n654 ), .A4(\AES_ENC/us11/n653 ), .ZN(\AES_ENC/us11/n657 ) );
NAND2_X2 \AES_ENC/us11/U436  ( .A1(\AES_ENC/sa11 [2]), .A2(\AES_ENC/us11/n657 ), .ZN(\AES_ENC/us11/n660 ) );
NAND4_X2 \AES_ENC/us11/U432  ( .A1(\AES_ENC/us11/n662 ), .A2(\AES_ENC/us11/n661 ), .A3(\AES_ENC/us11/n660 ), .A4(\AES_ENC/us11/n659 ), .ZN(\AES_ENC/us11/n663 ) );
NAND2_X2 \AES_ENC/us11/U431  ( .A1(\AES_ENC/us11/n663 ), .A2(\AES_ENC/us11/n574 ), .ZN(\AES_ENC/us11/n664 ) );
NAND2_X2 \AES_ENC/us11/U430  ( .A1(\AES_ENC/us11/n665 ), .A2(\AES_ENC/us11/n664 ), .ZN(\AES_ENC/us11/n666 ) );
NAND2_X2 \AES_ENC/us11/U429  ( .A1(\AES_ENC/sa11 [6]), .A2(\AES_ENC/us11/n666 ), .ZN(\AES_ENC/us11/n678 ) );
NAND2_X2 \AES_ENC/us11/U426  ( .A1(\AES_ENC/us11/n735 ), .A2(\AES_ENC/us11/n1093 ), .ZN(\AES_ENC/us11/n675 ) );
NAND2_X2 \AES_ENC/us11/U425  ( .A1(\AES_ENC/us11/n588 ), .A2(\AES_ENC/us11/n597 ), .ZN(\AES_ENC/us11/n1045 ) );
OR2_X2 \AES_ENC/us11/U424  ( .A1(\AES_ENC/us11/n1045 ), .A2(\AES_ENC/us11/n605 ), .ZN(\AES_ENC/us11/n674 ) );
NAND2_X2 \AES_ENC/us11/U423  ( .A1(\AES_ENC/sa11 [1]), .A2(\AES_ENC/us11/n620 ), .ZN(\AES_ENC/us11/n667 ) );
NAND2_X2 \AES_ENC/us11/U422  ( .A1(\AES_ENC/us11/n619 ), .A2(\AES_ENC/us11/n667 ), .ZN(\AES_ENC/us11/n1071 ) );
NAND4_X2 \AES_ENC/us11/U412  ( .A1(\AES_ENC/us11/n675 ), .A2(\AES_ENC/us11/n674 ), .A3(\AES_ENC/us11/n673 ), .A4(\AES_ENC/us11/n672 ), .ZN(\AES_ENC/us11/n676 ) );
NAND2_X2 \AES_ENC/us11/U411  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n676 ), .ZN(\AES_ENC/us11/n677 ) );
NAND2_X2 \AES_ENC/us11/U408  ( .A1(\AES_ENC/us11/n800 ), .A2(\AES_ENC/us11/n1022 ), .ZN(\AES_ENC/us11/n680 ) );
NAND2_X2 \AES_ENC/us11/U407  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n680 ), .ZN(\AES_ENC/us11/n681 ) );
AND2_X2 \AES_ENC/us11/U402  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n684 ), .ZN(\AES_ENC/us11/n682 ) );
NAND4_X2 \AES_ENC/us11/U395  ( .A1(\AES_ENC/us11/n691 ), .A2(\AES_ENC/us11/n581 ), .A3(\AES_ENC/us11/n690 ), .A4(\AES_ENC/us11/n689 ), .ZN(\AES_ENC/us11/n692 ) );
NAND2_X2 \AES_ENC/us11/U394  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n692 ), .ZN(\AES_ENC/us11/n733 ) );
NAND2_X2 \AES_ENC/us11/U392  ( .A1(\AES_ENC/us11/n977 ), .A2(\AES_ENC/us11/n1050 ), .ZN(\AES_ENC/us11/n702 ) );
NAND2_X2 \AES_ENC/us11/U391  ( .A1(\AES_ENC/us11/n1093 ), .A2(\AES_ENC/us11/n1045 ), .ZN(\AES_ENC/us11/n701 ) );
NAND4_X2 \AES_ENC/us11/U381  ( .A1(\AES_ENC/us11/n702 ), .A2(\AES_ENC/us11/n701 ), .A3(\AES_ENC/us11/n700 ), .A4(\AES_ENC/us11/n699 ), .ZN(\AES_ENC/us11/n703 ) );
NAND2_X2 \AES_ENC/us11/U380  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n703 ), .ZN(\AES_ENC/us11/n732 ) );
AND2_X2 \AES_ENC/us11/U379  ( .A1(\AES_ENC/sa11 [0]), .A2(\AES_ENC/sa11 [6]),.ZN(\AES_ENC/us11/n1113 ) );
NAND2_X2 \AES_ENC/us11/U378  ( .A1(\AES_ENC/us11/n601 ), .A2(\AES_ENC/us11/n1030 ), .ZN(\AES_ENC/us11/n881 ) );
NAND2_X2 \AES_ENC/us11/U377  ( .A1(\AES_ENC/us11/n1093 ), .A2(\AES_ENC/us11/n881 ), .ZN(\AES_ENC/us11/n715 ) );
NAND2_X2 \AES_ENC/us11/U376  ( .A1(\AES_ENC/us11/n1010 ), .A2(\AES_ENC/us11/n600 ), .ZN(\AES_ENC/us11/n714 ) );
NAND2_X2 \AES_ENC/us11/U375  ( .A1(\AES_ENC/us11/n855 ), .A2(\AES_ENC/us11/n588 ), .ZN(\AES_ENC/us11/n1117 ) );
XNOR2_X2 \AES_ENC/us11/U371  ( .A(\AES_ENC/us11/n611 ), .B(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n824 ) );
NAND4_X2 \AES_ENC/us11/U362  ( .A1(\AES_ENC/us11/n715 ), .A2(\AES_ENC/us11/n714 ), .A3(\AES_ENC/us11/n713 ), .A4(\AES_ENC/us11/n712 ), .ZN(\AES_ENC/us11/n716 ) );
NAND2_X2 \AES_ENC/us11/U361  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n716 ), .ZN(\AES_ENC/us11/n731 ) );
AND2_X2 \AES_ENC/us11/U360  ( .A1(\AES_ENC/sa11 [6]), .A2(\AES_ENC/us11/n574 ), .ZN(\AES_ENC/us11/n1131 ) );
NAND2_X2 \AES_ENC/us11/U359  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n717 ) );
NAND2_X2 \AES_ENC/us11/U358  ( .A1(\AES_ENC/us11/n1029 ), .A2(\AES_ENC/us11/n717 ), .ZN(\AES_ENC/us11/n728 ) );
NAND2_X2 \AES_ENC/us11/U357  ( .A1(\AES_ENC/sa11 [1]), .A2(\AES_ENC/us11/n624 ), .ZN(\AES_ENC/us11/n1097 ) );
NAND2_X2 \AES_ENC/us11/U356  ( .A1(\AES_ENC/us11/n603 ), .A2(\AES_ENC/us11/n1097 ), .ZN(\AES_ENC/us11/n718 ) );
NAND2_X2 \AES_ENC/us11/U355  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n718 ), .ZN(\AES_ENC/us11/n727 ) );
NAND4_X2 \AES_ENC/us11/U344  ( .A1(\AES_ENC/us11/n728 ), .A2(\AES_ENC/us11/n727 ), .A3(\AES_ENC/us11/n726 ), .A4(\AES_ENC/us11/n725 ), .ZN(\AES_ENC/us11/n729 ) );
NAND2_X2 \AES_ENC/us11/U343  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n729 ), .ZN(\AES_ENC/us11/n730 ) );
NAND4_X2 \AES_ENC/us11/U342  ( .A1(\AES_ENC/us11/n733 ), .A2(\AES_ENC/us11/n732 ), .A3(\AES_ENC/us11/n731 ), .A4(\AES_ENC/us11/n730 ), .ZN(\AES_ENC/sa11_sub[1] ) );
NAND2_X2 \AES_ENC/us11/U341  ( .A1(\AES_ENC/sa11 [7]), .A2(\AES_ENC/us11/n611 ), .ZN(\AES_ENC/us11/n734 ) );
NAND2_X2 \AES_ENC/us11/U340  ( .A1(\AES_ENC/us11/n734 ), .A2(\AES_ENC/us11/n607 ), .ZN(\AES_ENC/us11/n738 ) );
OR4_X2 \AES_ENC/us11/U339  ( .A1(\AES_ENC/us11/n738 ), .A2(\AES_ENC/us11/n626 ), .A3(\AES_ENC/us11/n826 ), .A4(\AES_ENC/us11/n1121 ), .ZN(\AES_ENC/us11/n746 ) );
NAND2_X2 \AES_ENC/us11/U337  ( .A1(\AES_ENC/us11/n1100 ), .A2(\AES_ENC/us11/n587 ), .ZN(\AES_ENC/us11/n992 ) );
OR2_X2 \AES_ENC/us11/U336  ( .A1(\AES_ENC/us11/n610 ), .A2(\AES_ENC/us11/n735 ), .ZN(\AES_ENC/us11/n737 ) );
NAND2_X2 \AES_ENC/us11/U334  ( .A1(\AES_ENC/us11/n619 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n753 ) );
NAND2_X2 \AES_ENC/us11/U333  ( .A1(\AES_ENC/us11/n582 ), .A2(\AES_ENC/us11/n753 ), .ZN(\AES_ENC/us11/n1080 ) );
NAND2_X2 \AES_ENC/us11/U332  ( .A1(\AES_ENC/us11/n1048 ), .A2(\AES_ENC/us11/n576 ), .ZN(\AES_ENC/us11/n736 ) );
NAND2_X2 \AES_ENC/us11/U331  ( .A1(\AES_ENC/us11/n737 ), .A2(\AES_ENC/us11/n736 ), .ZN(\AES_ENC/us11/n739 ) );
NAND2_X2 \AES_ENC/us11/U330  ( .A1(\AES_ENC/us11/n739 ), .A2(\AES_ENC/us11/n738 ), .ZN(\AES_ENC/us11/n745 ) );
NAND2_X2 \AES_ENC/us11/U326  ( .A1(\AES_ENC/us11/n1096 ), .A2(\AES_ENC/us11/n590 ), .ZN(\AES_ENC/us11/n906 ) );
NAND4_X2 \AES_ENC/us11/U323  ( .A1(\AES_ENC/us11/n746 ), .A2(\AES_ENC/us11/n992 ), .A3(\AES_ENC/us11/n745 ), .A4(\AES_ENC/us11/n744 ), .ZN(\AES_ENC/us11/n747 ) );
NAND2_X2 \AES_ENC/us11/U322  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n747 ), .ZN(\AES_ENC/us11/n793 ) );
NAND2_X2 \AES_ENC/us11/U321  ( .A1(\AES_ENC/us11/n584 ), .A2(\AES_ENC/us11/n855 ), .ZN(\AES_ENC/us11/n748 ) );
NAND2_X2 \AES_ENC/us11/U320  ( .A1(\AES_ENC/us11/n956 ), .A2(\AES_ENC/us11/n748 ), .ZN(\AES_ENC/us11/n760 ) );
NAND2_X2 \AES_ENC/us11/U313  ( .A1(\AES_ENC/us11/n590 ), .A2(\AES_ENC/us11/n753 ), .ZN(\AES_ENC/us11/n1023 ) );
NAND4_X2 \AES_ENC/us11/U308  ( .A1(\AES_ENC/us11/n760 ), .A2(\AES_ENC/us11/n992 ), .A3(\AES_ENC/us11/n759 ), .A4(\AES_ENC/us11/n758 ), .ZN(\AES_ENC/us11/n761 ) );
NAND2_X2 \AES_ENC/us11/U307  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n761 ), .ZN(\AES_ENC/us11/n792 ) );
NAND2_X2 \AES_ENC/us11/U306  ( .A1(\AES_ENC/us11/n584 ), .A2(\AES_ENC/us11/n603 ), .ZN(\AES_ENC/us11/n989 ) );
NAND2_X2 \AES_ENC/us11/U305  ( .A1(\AES_ENC/us11/n1050 ), .A2(\AES_ENC/us11/n989 ), .ZN(\AES_ENC/us11/n777 ) );
NAND2_X2 \AES_ENC/us11/U304  ( .A1(\AES_ENC/us11/n1093 ), .A2(\AES_ENC/us11/n762 ), .ZN(\AES_ENC/us11/n776 ) );
XNOR2_X2 \AES_ENC/us11/U301  ( .A(\AES_ENC/sa11 [7]), .B(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n959 ) );
NAND4_X2 \AES_ENC/us11/U289  ( .A1(\AES_ENC/us11/n777 ), .A2(\AES_ENC/us11/n776 ), .A3(\AES_ENC/us11/n775 ), .A4(\AES_ENC/us11/n774 ), .ZN(\AES_ENC/us11/n778 ) );
NAND2_X2 \AES_ENC/us11/U288  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n778 ), .ZN(\AES_ENC/us11/n791 ) );
NAND2_X2 \AES_ENC/us11/U287  ( .A1(\AES_ENC/us11/n1056 ), .A2(\AES_ENC/us11/n1050 ), .ZN(\AES_ENC/us11/n788 ) );
NAND2_X2 \AES_ENC/us11/U286  ( .A1(\AES_ENC/us11/n1091 ), .A2(\AES_ENC/us11/n779 ), .ZN(\AES_ENC/us11/n787 ) );
NAND2_X2 \AES_ENC/us11/U285  ( .A1(\AES_ENC/us11/n956 ), .A2(\AES_ENC/sa11 [1]), .ZN(\AES_ENC/us11/n786 ) );
NAND4_X2 \AES_ENC/us11/U278  ( .A1(\AES_ENC/us11/n788 ), .A2(\AES_ENC/us11/n787 ), .A3(\AES_ENC/us11/n786 ), .A4(\AES_ENC/us11/n785 ), .ZN(\AES_ENC/us11/n789 ) );
NAND2_X2 \AES_ENC/us11/U277  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n789 ), .ZN(\AES_ENC/us11/n790 ) );
NAND4_X2 \AES_ENC/us11/U276  ( .A1(\AES_ENC/us11/n793 ), .A2(\AES_ENC/us11/n792 ), .A3(\AES_ENC/us11/n791 ), .A4(\AES_ENC/us11/n790 ), .ZN(\AES_ENC/sa11_sub[2] ) );
NAND2_X2 \AES_ENC/us11/U275  ( .A1(\AES_ENC/us11/n1059 ), .A2(\AES_ENC/us11/n794 ), .ZN(\AES_ENC/us11/n810 ) );
NAND2_X2 \AES_ENC/us11/U274  ( .A1(\AES_ENC/us11/n1049 ), .A2(\AES_ENC/us11/n956 ), .ZN(\AES_ENC/us11/n809 ) );
OR2_X2 \AES_ENC/us11/U266  ( .A1(\AES_ENC/us11/n1096 ), .A2(\AES_ENC/us11/n606 ), .ZN(\AES_ENC/us11/n802 ) );
NAND2_X2 \AES_ENC/us11/U265  ( .A1(\AES_ENC/us11/n1053 ), .A2(\AES_ENC/us11/n800 ), .ZN(\AES_ENC/us11/n801 ) );
NAND2_X2 \AES_ENC/us11/U264  ( .A1(\AES_ENC/us11/n802 ), .A2(\AES_ENC/us11/n801 ), .ZN(\AES_ENC/us11/n805 ) );
NAND4_X2 \AES_ENC/us11/U261  ( .A1(\AES_ENC/us11/n810 ), .A2(\AES_ENC/us11/n809 ), .A3(\AES_ENC/us11/n808 ), .A4(\AES_ENC/us11/n807 ), .ZN(\AES_ENC/us11/n811 ) );
NAND2_X2 \AES_ENC/us11/U260  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n811 ), .ZN(\AES_ENC/us11/n852 ) );
OR2_X2 \AES_ENC/us11/U259  ( .A1(\AES_ENC/us11/n1023 ), .A2(\AES_ENC/us11/n617 ), .ZN(\AES_ENC/us11/n819 ) );
OR2_X2 \AES_ENC/us11/U257  ( .A1(\AES_ENC/us11/n570 ), .A2(\AES_ENC/us11/n930 ), .ZN(\AES_ENC/us11/n818 ) );
NAND2_X2 \AES_ENC/us11/U256  ( .A1(\AES_ENC/us11/n1013 ), .A2(\AES_ENC/us11/n1094 ), .ZN(\AES_ENC/us11/n817 ) );
NAND4_X2 \AES_ENC/us11/U249  ( .A1(\AES_ENC/us11/n819 ), .A2(\AES_ENC/us11/n818 ), .A3(\AES_ENC/us11/n817 ), .A4(\AES_ENC/us11/n816 ), .ZN(\AES_ENC/us11/n820 ) );
NAND2_X2 \AES_ENC/us11/U248  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n820 ), .ZN(\AES_ENC/us11/n851 ) );
NAND2_X2 \AES_ENC/us11/U247  ( .A1(\AES_ENC/us11/n956 ), .A2(\AES_ENC/us11/n1080 ), .ZN(\AES_ENC/us11/n835 ) );
NAND2_X2 \AES_ENC/us11/U246  ( .A1(\AES_ENC/us11/n570 ), .A2(\AES_ENC/us11/n1030 ), .ZN(\AES_ENC/us11/n1047 ) );
OR2_X2 \AES_ENC/us11/U245  ( .A1(\AES_ENC/us11/n1047 ), .A2(\AES_ENC/us11/n612 ), .ZN(\AES_ENC/us11/n834 ) );
NAND2_X2 \AES_ENC/us11/U244  ( .A1(\AES_ENC/us11/n1072 ), .A2(\AES_ENC/us11/n589 ), .ZN(\AES_ENC/us11/n833 ) );
NAND4_X2 \AES_ENC/us11/U233  ( .A1(\AES_ENC/us11/n835 ), .A2(\AES_ENC/us11/n834 ), .A3(\AES_ENC/us11/n833 ), .A4(\AES_ENC/us11/n832 ), .ZN(\AES_ENC/us11/n836 ) );
NAND2_X2 \AES_ENC/us11/U232  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n836 ), .ZN(\AES_ENC/us11/n850 ) );
NAND2_X2 \AES_ENC/us11/U231  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n623 ), .ZN(\AES_ENC/us11/n847 ) );
NAND2_X2 \AES_ENC/us11/U230  ( .A1(\AES_ENC/us11/n1050 ), .A2(\AES_ENC/us11/n1071 ), .ZN(\AES_ENC/us11/n846 ) );
OR2_X2 \AES_ENC/us11/U224  ( .A1(\AES_ENC/us11/n1053 ), .A2(\AES_ENC/us11/n911 ), .ZN(\AES_ENC/us11/n1077 ) );
NAND4_X2 \AES_ENC/us11/U220  ( .A1(\AES_ENC/us11/n847 ), .A2(\AES_ENC/us11/n846 ), .A3(\AES_ENC/us11/n845 ), .A4(\AES_ENC/us11/n844 ), .ZN(\AES_ENC/us11/n848 ) );
NAND2_X2 \AES_ENC/us11/U219  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n848 ), .ZN(\AES_ENC/us11/n849 ) );
NAND4_X2 \AES_ENC/us11/U218  ( .A1(\AES_ENC/us11/n852 ), .A2(\AES_ENC/us11/n851 ), .A3(\AES_ENC/us11/n850 ), .A4(\AES_ENC/us11/n849 ), .ZN(\AES_ENC/sa11_sub[3] ) );
NAND2_X2 \AES_ENC/us11/U216  ( .A1(\AES_ENC/us11/n1009 ), .A2(\AES_ENC/us11/n1072 ), .ZN(\AES_ENC/us11/n862 ) );
NAND2_X2 \AES_ENC/us11/U215  ( .A1(\AES_ENC/us11/n603 ), .A2(\AES_ENC/us11/n577 ), .ZN(\AES_ENC/us11/n853 ) );
NAND2_X2 \AES_ENC/us11/U214  ( .A1(\AES_ENC/us11/n1050 ), .A2(\AES_ENC/us11/n853 ), .ZN(\AES_ENC/us11/n861 ) );
NAND4_X2 \AES_ENC/us11/U206  ( .A1(\AES_ENC/us11/n862 ), .A2(\AES_ENC/us11/n861 ), .A3(\AES_ENC/us11/n860 ), .A4(\AES_ENC/us11/n859 ), .ZN(\AES_ENC/us11/n863 ) );
NAND2_X2 \AES_ENC/us11/U205  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n863 ), .ZN(\AES_ENC/us11/n905 ) );
NAND2_X2 \AES_ENC/us11/U204  ( .A1(\AES_ENC/us11/n1010 ), .A2(\AES_ENC/us11/n989 ), .ZN(\AES_ENC/us11/n874 ) );
NAND2_X2 \AES_ENC/us11/U203  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n610 ), .ZN(\AES_ENC/us11/n864 ) );
NAND2_X2 \AES_ENC/us11/U202  ( .A1(\AES_ENC/us11/n929 ), .A2(\AES_ENC/us11/n864 ), .ZN(\AES_ENC/us11/n873 ) );
NAND4_X2 \AES_ENC/us11/U193  ( .A1(\AES_ENC/us11/n874 ), .A2(\AES_ENC/us11/n873 ), .A3(\AES_ENC/us11/n872 ), .A4(\AES_ENC/us11/n871 ), .ZN(\AES_ENC/us11/n875 ) );
NAND2_X2 \AES_ENC/us11/U192  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n875 ), .ZN(\AES_ENC/us11/n904 ) );
NAND2_X2 \AES_ENC/us11/U191  ( .A1(\AES_ENC/us11/n583 ), .A2(\AES_ENC/us11/n1050 ), .ZN(\AES_ENC/us11/n889 ) );
NAND2_X2 \AES_ENC/us11/U190  ( .A1(\AES_ENC/us11/n1093 ), .A2(\AES_ENC/us11/n587 ), .ZN(\AES_ENC/us11/n876 ) );
NAND2_X2 \AES_ENC/us11/U189  ( .A1(\AES_ENC/us11/n604 ), .A2(\AES_ENC/us11/n876 ), .ZN(\AES_ENC/us11/n877 ) );
NAND2_X2 \AES_ENC/us11/U188  ( .A1(\AES_ENC/us11/n877 ), .A2(\AES_ENC/us11/n623 ), .ZN(\AES_ENC/us11/n888 ) );
NAND4_X2 \AES_ENC/us11/U179  ( .A1(\AES_ENC/us11/n889 ), .A2(\AES_ENC/us11/n888 ), .A3(\AES_ENC/us11/n887 ), .A4(\AES_ENC/us11/n886 ), .ZN(\AES_ENC/us11/n890 ) );
NAND2_X2 \AES_ENC/us11/U178  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n890 ), .ZN(\AES_ENC/us11/n903 ) );
OR2_X2 \AES_ENC/us11/U177  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n1059 ), .ZN(\AES_ENC/us11/n900 ) );
NAND2_X2 \AES_ENC/us11/U176  ( .A1(\AES_ENC/us11/n1073 ), .A2(\AES_ENC/us11/n1047 ), .ZN(\AES_ENC/us11/n899 ) );
NAND2_X2 \AES_ENC/us11/U175  ( .A1(\AES_ENC/us11/n1094 ), .A2(\AES_ENC/us11/n595 ), .ZN(\AES_ENC/us11/n898 ) );
NAND4_X2 \AES_ENC/us11/U167  ( .A1(\AES_ENC/us11/n900 ), .A2(\AES_ENC/us11/n899 ), .A3(\AES_ENC/us11/n898 ), .A4(\AES_ENC/us11/n897 ), .ZN(\AES_ENC/us11/n901 ) );
NAND2_X2 \AES_ENC/us11/U166  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n901 ), .ZN(\AES_ENC/us11/n902 ) );
NAND4_X2 \AES_ENC/us11/U165  ( .A1(\AES_ENC/us11/n905 ), .A2(\AES_ENC/us11/n904 ), .A3(\AES_ENC/us11/n903 ), .A4(\AES_ENC/us11/n902 ), .ZN(\AES_ENC/sa11_sub[4] ) );
NAND2_X2 \AES_ENC/us11/U164  ( .A1(\AES_ENC/us11/n1094 ), .A2(\AES_ENC/us11/n599 ), .ZN(\AES_ENC/us11/n922 ) );
NAND2_X2 \AES_ENC/us11/U163  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n989 ), .ZN(\AES_ENC/us11/n921 ) );
NAND4_X2 \AES_ENC/us11/U151  ( .A1(\AES_ENC/us11/n922 ), .A2(\AES_ENC/us11/n921 ), .A3(\AES_ENC/us11/n920 ), .A4(\AES_ENC/us11/n919 ), .ZN(\AES_ENC/us11/n923 ) );
NAND2_X2 \AES_ENC/us11/U150  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n923 ), .ZN(\AES_ENC/us11/n972 ) );
NAND2_X2 \AES_ENC/us11/U149  ( .A1(\AES_ENC/us11/n582 ), .A2(\AES_ENC/us11/n619 ), .ZN(\AES_ENC/us11/n924 ) );
NAND2_X2 \AES_ENC/us11/U148  ( .A1(\AES_ENC/us11/n1073 ), .A2(\AES_ENC/us11/n924 ), .ZN(\AES_ENC/us11/n939 ) );
NAND2_X2 \AES_ENC/us11/U147  ( .A1(\AES_ENC/us11/n926 ), .A2(\AES_ENC/us11/n925 ), .ZN(\AES_ENC/us11/n927 ) );
NAND2_X2 \AES_ENC/us11/U146  ( .A1(\AES_ENC/us11/n606 ), .A2(\AES_ENC/us11/n927 ), .ZN(\AES_ENC/us11/n928 ) );
NAND2_X2 \AES_ENC/us11/U145  ( .A1(\AES_ENC/us11/n928 ), .A2(\AES_ENC/us11/n1080 ), .ZN(\AES_ENC/us11/n938 ) );
OR2_X2 \AES_ENC/us11/U144  ( .A1(\AES_ENC/us11/n1117 ), .A2(\AES_ENC/us11/n615 ), .ZN(\AES_ENC/us11/n937 ) );
NAND4_X2 \AES_ENC/us11/U139  ( .A1(\AES_ENC/us11/n939 ), .A2(\AES_ENC/us11/n938 ), .A3(\AES_ENC/us11/n937 ), .A4(\AES_ENC/us11/n936 ), .ZN(\AES_ENC/us11/n940 ) );
NAND2_X2 \AES_ENC/us11/U138  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n940 ), .ZN(\AES_ENC/us11/n971 ) );
OR2_X2 \AES_ENC/us11/U137  ( .A1(\AES_ENC/us11/n605 ), .A2(\AES_ENC/us11/n941 ), .ZN(\AES_ENC/us11/n954 ) );
NAND2_X2 \AES_ENC/us11/U136  ( .A1(\AES_ENC/us11/n1096 ), .A2(\AES_ENC/us11/n577 ), .ZN(\AES_ENC/us11/n942 ) );
NAND2_X2 \AES_ENC/us11/U135  ( .A1(\AES_ENC/us11/n1048 ), .A2(\AES_ENC/us11/n942 ), .ZN(\AES_ENC/us11/n943 ) );
NAND2_X2 \AES_ENC/us11/U134  ( .A1(\AES_ENC/us11/n612 ), .A2(\AES_ENC/us11/n943 ), .ZN(\AES_ENC/us11/n944 ) );
NAND2_X2 \AES_ENC/us11/U133  ( .A1(\AES_ENC/us11/n944 ), .A2(\AES_ENC/us11/n580 ), .ZN(\AES_ENC/us11/n953 ) );
NAND4_X2 \AES_ENC/us11/U125  ( .A1(\AES_ENC/us11/n954 ), .A2(\AES_ENC/us11/n953 ), .A3(\AES_ENC/us11/n952 ), .A4(\AES_ENC/us11/n951 ), .ZN(\AES_ENC/us11/n955 ) );
NAND2_X2 \AES_ENC/us11/U124  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n955 ), .ZN(\AES_ENC/us11/n970 ) );
NAND2_X2 \AES_ENC/us11/U123  ( .A1(\AES_ENC/us11/n1094 ), .A2(\AES_ENC/us11/n1071 ), .ZN(\AES_ENC/us11/n967 ) );
NAND2_X2 \AES_ENC/us11/U122  ( .A1(\AES_ENC/us11/n956 ), .A2(\AES_ENC/us11/n1030 ), .ZN(\AES_ENC/us11/n966 ) );
NAND4_X2 \AES_ENC/us11/U114  ( .A1(\AES_ENC/us11/n967 ), .A2(\AES_ENC/us11/n966 ), .A3(\AES_ENC/us11/n965 ), .A4(\AES_ENC/us11/n964 ), .ZN(\AES_ENC/us11/n968 ) );
NAND2_X2 \AES_ENC/us11/U113  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n968 ), .ZN(\AES_ENC/us11/n969 ) );
NAND4_X2 \AES_ENC/us11/U112  ( .A1(\AES_ENC/us11/n972 ), .A2(\AES_ENC/us11/n971 ), .A3(\AES_ENC/us11/n970 ), .A4(\AES_ENC/us11/n969 ), .ZN(\AES_ENC/sa11_sub[5] ) );
NAND2_X2 \AES_ENC/us11/U111  ( .A1(\AES_ENC/us11/n570 ), .A2(\AES_ENC/us11/n1097 ), .ZN(\AES_ENC/us11/n973 ) );
NAND2_X2 \AES_ENC/us11/U110  ( .A1(\AES_ENC/us11/n1073 ), .A2(\AES_ENC/us11/n973 ), .ZN(\AES_ENC/us11/n987 ) );
NAND2_X2 \AES_ENC/us11/U109  ( .A1(\AES_ENC/us11/n974 ), .A2(\AES_ENC/us11/n1077 ), .ZN(\AES_ENC/us11/n975 ) );
NAND2_X2 \AES_ENC/us11/U108  ( .A1(\AES_ENC/us11/n613 ), .A2(\AES_ENC/us11/n975 ), .ZN(\AES_ENC/us11/n976 ) );
NAND2_X2 \AES_ENC/us11/U107  ( .A1(\AES_ENC/us11/n977 ), .A2(\AES_ENC/us11/n976 ), .ZN(\AES_ENC/us11/n986 ) );
NAND4_X2 \AES_ENC/us11/U99  ( .A1(\AES_ENC/us11/n987 ), .A2(\AES_ENC/us11/n986 ), .A3(\AES_ENC/us11/n985 ), .A4(\AES_ENC/us11/n984 ), .ZN(\AES_ENC/us11/n988 ) );
NAND2_X2 \AES_ENC/us11/U98  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n988 ), .ZN(\AES_ENC/us11/n1044 ) );
NAND2_X2 \AES_ENC/us11/U97  ( .A1(\AES_ENC/us11/n1073 ), .A2(\AES_ENC/us11/n989 ), .ZN(\AES_ENC/us11/n1004 ) );
NAND2_X2 \AES_ENC/us11/U96  ( .A1(\AES_ENC/us11/n1092 ), .A2(\AES_ENC/us11/n619 ), .ZN(\AES_ENC/us11/n1003 ) );
NAND4_X2 \AES_ENC/us11/U85  ( .A1(\AES_ENC/us11/n1004 ), .A2(\AES_ENC/us11/n1003 ), .A3(\AES_ENC/us11/n1002 ), .A4(\AES_ENC/us11/n1001 ), .ZN(\AES_ENC/us11/n1005 ) );
NAND2_X2 \AES_ENC/us11/U84  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n1005 ), .ZN(\AES_ENC/us11/n1043 ) );
NAND2_X2 \AES_ENC/us11/U83  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n596 ), .ZN(\AES_ENC/us11/n1020 ) );
NAND2_X2 \AES_ENC/us11/U82  ( .A1(\AES_ENC/us11/n1050 ), .A2(\AES_ENC/us11/n624 ), .ZN(\AES_ENC/us11/n1019 ) );
NAND2_X2 \AES_ENC/us11/U77  ( .A1(\AES_ENC/us11/n1059 ), .A2(\AES_ENC/us11/n1114 ), .ZN(\AES_ENC/us11/n1012 ) );
NAND2_X2 \AES_ENC/us11/U76  ( .A1(\AES_ENC/us11/n1010 ), .A2(\AES_ENC/us11/n592 ), .ZN(\AES_ENC/us11/n1011 ) );
NAND2_X2 \AES_ENC/us11/U75  ( .A1(\AES_ENC/us11/n1012 ), .A2(\AES_ENC/us11/n1011 ), .ZN(\AES_ENC/us11/n1016 ) );
NAND4_X2 \AES_ENC/us11/U70  ( .A1(\AES_ENC/us11/n1020 ), .A2(\AES_ENC/us11/n1019 ), .A3(\AES_ENC/us11/n1018 ), .A4(\AES_ENC/us11/n1017 ), .ZN(\AES_ENC/us11/n1021 ) );
NAND2_X2 \AES_ENC/us11/U69  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n1021 ), .ZN(\AES_ENC/us11/n1042 ) );
NAND2_X2 \AES_ENC/us11/U68  ( .A1(\AES_ENC/us11/n1022 ), .A2(\AES_ENC/us11/n1093 ), .ZN(\AES_ENC/us11/n1039 ) );
NAND2_X2 \AES_ENC/us11/U67  ( .A1(\AES_ENC/us11/n1050 ), .A2(\AES_ENC/us11/n1023 ), .ZN(\AES_ENC/us11/n1038 ) );
NAND2_X2 \AES_ENC/us11/U66  ( .A1(\AES_ENC/us11/n1024 ), .A2(\AES_ENC/us11/n1071 ), .ZN(\AES_ENC/us11/n1037 ) );
AND2_X2 \AES_ENC/us11/U60  ( .A1(\AES_ENC/us11/n1030 ), .A2(\AES_ENC/us11/n602 ), .ZN(\AES_ENC/us11/n1078 ) );
NAND4_X2 \AES_ENC/us11/U56  ( .A1(\AES_ENC/us11/n1039 ), .A2(\AES_ENC/us11/n1038 ), .A3(\AES_ENC/us11/n1037 ), .A4(\AES_ENC/us11/n1036 ), .ZN(\AES_ENC/us11/n1040 ) );
NAND2_X2 \AES_ENC/us11/U55  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n1040 ), .ZN(\AES_ENC/us11/n1041 ) );
NAND4_X2 \AES_ENC/us11/U54  ( .A1(\AES_ENC/us11/n1044 ), .A2(\AES_ENC/us11/n1043 ), .A3(\AES_ENC/us11/n1042 ), .A4(\AES_ENC/us11/n1041 ), .ZN(\AES_ENC/sa11_sub[6] ) );
NAND2_X2 \AES_ENC/us11/U53  ( .A1(\AES_ENC/us11/n1072 ), .A2(\AES_ENC/us11/n1045 ), .ZN(\AES_ENC/us11/n1068 ) );
NAND2_X2 \AES_ENC/us11/U52  ( .A1(\AES_ENC/us11/n1046 ), .A2(\AES_ENC/us11/n582 ), .ZN(\AES_ENC/us11/n1067 ) );
NAND2_X2 \AES_ENC/us11/U51  ( .A1(\AES_ENC/us11/n1094 ), .A2(\AES_ENC/us11/n1047 ), .ZN(\AES_ENC/us11/n1066 ) );
NAND4_X2 \AES_ENC/us11/U40  ( .A1(\AES_ENC/us11/n1068 ), .A2(\AES_ENC/us11/n1067 ), .A3(\AES_ENC/us11/n1066 ), .A4(\AES_ENC/us11/n1065 ), .ZN(\AES_ENC/us11/n1069 ) );
NAND2_X2 \AES_ENC/us11/U39  ( .A1(\AES_ENC/us11/n1070 ), .A2(\AES_ENC/us11/n1069 ), .ZN(\AES_ENC/us11/n1135 ) );
NAND2_X2 \AES_ENC/us11/U38  ( .A1(\AES_ENC/us11/n1072 ), .A2(\AES_ENC/us11/n1071 ), .ZN(\AES_ENC/us11/n1088 ) );
NAND2_X2 \AES_ENC/us11/U37  ( .A1(\AES_ENC/us11/n1073 ), .A2(\AES_ENC/us11/n595 ), .ZN(\AES_ENC/us11/n1087 ) );
NAND4_X2 \AES_ENC/us11/U28  ( .A1(\AES_ENC/us11/n1088 ), .A2(\AES_ENC/us11/n1087 ), .A3(\AES_ENC/us11/n1086 ), .A4(\AES_ENC/us11/n1085 ), .ZN(\AES_ENC/us11/n1089 ) );
NAND2_X2 \AES_ENC/us11/U27  ( .A1(\AES_ENC/us11/n1090 ), .A2(\AES_ENC/us11/n1089 ), .ZN(\AES_ENC/us11/n1134 ) );
NAND2_X2 \AES_ENC/us11/U26  ( .A1(\AES_ENC/us11/n1091 ), .A2(\AES_ENC/us11/n1093 ), .ZN(\AES_ENC/us11/n1111 ) );
NAND2_X2 \AES_ENC/us11/U25  ( .A1(\AES_ENC/us11/n1092 ), .A2(\AES_ENC/us11/n1120 ), .ZN(\AES_ENC/us11/n1110 ) );
AND2_X2 \AES_ENC/us11/U22  ( .A1(\AES_ENC/us11/n1097 ), .A2(\AES_ENC/us11/n1096 ), .ZN(\AES_ENC/us11/n1098 ) );
NAND4_X2 \AES_ENC/us11/U14  ( .A1(\AES_ENC/us11/n1111 ), .A2(\AES_ENC/us11/n1110 ), .A3(\AES_ENC/us11/n1109 ), .A4(\AES_ENC/us11/n1108 ), .ZN(\AES_ENC/us11/n1112 ) );
NAND2_X2 \AES_ENC/us11/U13  ( .A1(\AES_ENC/us11/n1113 ), .A2(\AES_ENC/us11/n1112 ), .ZN(\AES_ENC/us11/n1133 ) );
NAND2_X2 \AES_ENC/us11/U12  ( .A1(\AES_ENC/us11/n1115 ), .A2(\AES_ENC/us11/n1114 ), .ZN(\AES_ENC/us11/n1129 ) );
OR2_X2 \AES_ENC/us11/U11  ( .A1(\AES_ENC/us11/n608 ), .A2(\AES_ENC/us11/n1116 ), .ZN(\AES_ENC/us11/n1128 ) );
NAND4_X2 \AES_ENC/us11/U3  ( .A1(\AES_ENC/us11/n1129 ), .A2(\AES_ENC/us11/n1128 ), .A3(\AES_ENC/us11/n1127 ), .A4(\AES_ENC/us11/n1126 ), .ZN(\AES_ENC/us11/n1130 ) );
NAND2_X2 \AES_ENC/us11/U2  ( .A1(\AES_ENC/us11/n1131 ), .A2(\AES_ENC/us11/n1130 ), .ZN(\AES_ENC/us11/n1132 ) );
NAND4_X2 \AES_ENC/us11/U1  ( .A1(\AES_ENC/us11/n1135 ), .A2(\AES_ENC/us11/n1134 ), .A3(\AES_ENC/us11/n1133 ), .A4(\AES_ENC/us11/n1132 ), .ZN(\AES_ENC/sa11_sub[7] ) );
INV_X4 \AES_ENC/us12/U575  ( .A(\AES_ENC/sa12 [7]), .ZN(\AES_ENC/us12/n627 ));
INV_X4 \AES_ENC/us12/U574  ( .A(\AES_ENC/us12/n1114 ), .ZN(\AES_ENC/us12/n625 ) );
INV_X4 \AES_ENC/us12/U573  ( .A(\AES_ENC/sa12 [4]), .ZN(\AES_ENC/us12/n624 ));
INV_X4 \AES_ENC/us12/U572  ( .A(\AES_ENC/us12/n1025 ), .ZN(\AES_ENC/us12/n622 ) );
INV_X4 \AES_ENC/us12/U571  ( .A(\AES_ENC/us12/n1120 ), .ZN(\AES_ENC/us12/n620 ) );
INV_X4 \AES_ENC/us12/U570  ( .A(\AES_ENC/us12/n1121 ), .ZN(\AES_ENC/us12/n619 ) );
INV_X4 \AES_ENC/us12/U569  ( .A(\AES_ENC/us12/n1048 ), .ZN(\AES_ENC/us12/n618 ) );
INV_X4 \AES_ENC/us12/U568  ( .A(\AES_ENC/us12/n974 ), .ZN(\AES_ENC/us12/n616 ) );
INV_X4 \AES_ENC/us12/U567  ( .A(\AES_ENC/us12/n794 ), .ZN(\AES_ENC/us12/n614 ) );
INV_X4 \AES_ENC/us12/U566  ( .A(\AES_ENC/sa12 [2]), .ZN(\AES_ENC/us12/n611 ));
INV_X4 \AES_ENC/us12/U565  ( .A(\AES_ENC/us12/n800 ), .ZN(\AES_ENC/us12/n610 ) );
INV_X4 \AES_ENC/us12/U564  ( .A(\AES_ENC/us12/n925 ), .ZN(\AES_ENC/us12/n609 ) );
INV_X4 \AES_ENC/us12/U563  ( .A(\AES_ENC/us12/n779 ), .ZN(\AES_ENC/us12/n607 ) );
INV_X4 \AES_ENC/us12/U562  ( .A(\AES_ENC/us12/n1022 ), .ZN(\AES_ENC/us12/n603 ) );
INV_X4 \AES_ENC/us12/U561  ( .A(\AES_ENC/us12/n1102 ), .ZN(\AES_ENC/us12/n602 ) );
INV_X4 \AES_ENC/us12/U560  ( .A(\AES_ENC/us12/n929 ), .ZN(\AES_ENC/us12/n601 ) );
INV_X4 \AES_ENC/us12/U559  ( .A(\AES_ENC/us12/n1056 ), .ZN(\AES_ENC/us12/n600 ) );
INV_X4 \AES_ENC/us12/U558  ( .A(\AES_ENC/us12/n1054 ), .ZN(\AES_ENC/us12/n599 ) );
INV_X4 \AES_ENC/us12/U557  ( .A(\AES_ENC/us12/n881 ), .ZN(\AES_ENC/us12/n598 ) );
INV_X4 \AES_ENC/us12/U556  ( .A(\AES_ENC/us12/n926 ), .ZN(\AES_ENC/us12/n597 ) );
INV_X4 \AES_ENC/us12/U555  ( .A(\AES_ENC/us12/n977 ), .ZN(\AES_ENC/us12/n595 ) );
INV_X4 \AES_ENC/us12/U554  ( .A(\AES_ENC/us12/n1031 ), .ZN(\AES_ENC/us12/n594 ) );
INV_X4 \AES_ENC/us12/U553  ( .A(\AES_ENC/us12/n1103 ), .ZN(\AES_ENC/us12/n593 ) );
INV_X4 \AES_ENC/us12/U552  ( .A(\AES_ENC/us12/n1009 ), .ZN(\AES_ENC/us12/n592 ) );
INV_X4 \AES_ENC/us12/U551  ( .A(\AES_ENC/us12/n990 ), .ZN(\AES_ENC/us12/n591 ) );
INV_X4 \AES_ENC/us12/U550  ( .A(\AES_ENC/us12/n1058 ), .ZN(\AES_ENC/us12/n590 ) );
INV_X4 \AES_ENC/us12/U549  ( .A(\AES_ENC/us12/n1074 ), .ZN(\AES_ENC/us12/n589 ) );
INV_X4 \AES_ENC/us12/U548  ( .A(\AES_ENC/us12/n1053 ), .ZN(\AES_ENC/us12/n588 ) );
INV_X4 \AES_ENC/us12/U547  ( .A(\AES_ENC/us12/n826 ), .ZN(\AES_ENC/us12/n587 ) );
INV_X4 \AES_ENC/us12/U546  ( .A(\AES_ENC/us12/n992 ), .ZN(\AES_ENC/us12/n586 ) );
INV_X4 \AES_ENC/us12/U545  ( .A(\AES_ENC/us12/n821 ), .ZN(\AES_ENC/us12/n585 ) );
INV_X4 \AES_ENC/us12/U544  ( .A(\AES_ENC/us12/n910 ), .ZN(\AES_ENC/us12/n584 ) );
INV_X4 \AES_ENC/us12/U543  ( .A(\AES_ENC/us12/n906 ), .ZN(\AES_ENC/us12/n583 ) );
INV_X4 \AES_ENC/us12/U542  ( .A(\AES_ENC/us12/n880 ), .ZN(\AES_ENC/us12/n581 ) );
INV_X4 \AES_ENC/us12/U541  ( .A(\AES_ENC/us12/n1013 ), .ZN(\AES_ENC/us12/n580 ) );
INV_X4 \AES_ENC/us12/U540  ( .A(\AES_ENC/us12/n1092 ), .ZN(\AES_ENC/us12/n579 ) );
INV_X4 \AES_ENC/us12/U539  ( .A(\AES_ENC/us12/n824 ), .ZN(\AES_ENC/us12/n578 ) );
INV_X4 \AES_ENC/us12/U538  ( .A(\AES_ENC/us12/n1091 ), .ZN(\AES_ENC/us12/n577 ) );
INV_X4 \AES_ENC/us12/U537  ( .A(\AES_ENC/us12/n1080 ), .ZN(\AES_ENC/us12/n576 ) );
INV_X4 \AES_ENC/us12/U536  ( .A(\AES_ENC/us12/n959 ), .ZN(\AES_ENC/us12/n575 ) );
INV_X4 \AES_ENC/us12/U535  ( .A(\AES_ENC/sa12 [0]), .ZN(\AES_ENC/us12/n574 ));
NOR2_X2 \AES_ENC/us12/U534  ( .A1(\AES_ENC/sa12 [0]), .A2(\AES_ENC/sa12 [6]),.ZN(\AES_ENC/us12/n1090 ) );
NOR2_X2 \AES_ENC/us12/U533  ( .A1(\AES_ENC/us12/n574 ), .A2(\AES_ENC/sa12 [6]), .ZN(\AES_ENC/us12/n1070 ) );
NOR2_X2 \AES_ENC/us12/U532  ( .A1(\AES_ENC/sa12 [4]), .A2(\AES_ENC/sa12 [3]),.ZN(\AES_ENC/us12/n1025 ) );
INV_X4 \AES_ENC/us12/U531  ( .A(\AES_ENC/us12/n569 ), .ZN(\AES_ENC/us12/n572 ) );
NOR2_X2 \AES_ENC/us12/U530  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n765 ) );
NOR2_X2 \AES_ENC/us12/U529  ( .A1(\AES_ENC/sa12 [4]), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n764 ) );
NOR2_X2 \AES_ENC/us12/U528  ( .A1(\AES_ENC/us12/n765 ), .A2(\AES_ENC/us12/n764 ), .ZN(\AES_ENC/us12/n766 ) );
NOR2_X2 \AES_ENC/us12/U527  ( .A1(\AES_ENC/us12/n766 ), .A2(\AES_ENC/us12/n575 ), .ZN(\AES_ENC/us12/n767 ) );
NOR3_X2 \AES_ENC/us12/U526  ( .A1(\AES_ENC/us12/n627 ), .A2(\AES_ENC/sa12 [5]), .A3(\AES_ENC/us12/n704 ), .ZN(\AES_ENC/us12/n706 ));
NOR2_X2 \AES_ENC/us12/U525  ( .A1(\AES_ENC/us12/n1117 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n707 ) );
NOR2_X2 \AES_ENC/us12/U524  ( .A1(\AES_ENC/sa12 [4]), .A2(\AES_ENC/us12/n579 ), .ZN(\AES_ENC/us12/n705 ) );
NOR3_X2 \AES_ENC/us12/U523  ( .A1(\AES_ENC/us12/n707 ), .A2(\AES_ENC/us12/n706 ), .A3(\AES_ENC/us12/n705 ), .ZN(\AES_ENC/us12/n713 ) );
INV_X4 \AES_ENC/us12/U522  ( .A(\AES_ENC/sa12 [3]), .ZN(\AES_ENC/us12/n621 ));
NAND3_X2 \AES_ENC/us12/U521  ( .A1(\AES_ENC/us12/n652 ), .A2(\AES_ENC/us12/n626 ), .A3(\AES_ENC/sa12 [7]), .ZN(\AES_ENC/us12/n653 ));
NOR2_X2 \AES_ENC/us12/U520  ( .A1(\AES_ENC/us12/n611 ), .A2(\AES_ENC/sa12 [5]), .ZN(\AES_ENC/us12/n925 ) );
NOR2_X2 \AES_ENC/us12/U519  ( .A1(\AES_ENC/sa12 [5]), .A2(\AES_ENC/sa12 [2]),.ZN(\AES_ENC/us12/n974 ) );
INV_X4 \AES_ENC/us12/U518  ( .A(\AES_ENC/sa12 [5]), .ZN(\AES_ENC/us12/n626 ));
NOR2_X2 \AES_ENC/us12/U517  ( .A1(\AES_ENC/us12/n611 ), .A2(\AES_ENC/sa12 [7]), .ZN(\AES_ENC/us12/n779 ) );
NAND3_X2 \AES_ENC/us12/U516  ( .A1(\AES_ENC/us12/n679 ), .A2(\AES_ENC/us12/n678 ), .A3(\AES_ENC/us12/n677 ), .ZN(\AES_ENC/sa12_sub[0] ) );
NOR2_X2 \AES_ENC/us12/U515  ( .A1(\AES_ENC/us12/n626 ), .A2(\AES_ENC/sa12 [2]), .ZN(\AES_ENC/us12/n1048 ) );
NOR4_X2 \AES_ENC/us12/U512  ( .A1(\AES_ENC/us12/n633 ), .A2(\AES_ENC/us12/n632 ), .A3(\AES_ENC/us12/n631 ), .A4(\AES_ENC/us12/n630 ), .ZN(\AES_ENC/us12/n634 ) );
NOR2_X2 \AES_ENC/us12/U510  ( .A1(\AES_ENC/us12/n629 ), .A2(\AES_ENC/us12/n628 ), .ZN(\AES_ENC/us12/n635 ) );
NAND3_X2 \AES_ENC/us12/U509  ( .A1(\AES_ENC/sa12 [2]), .A2(\AES_ENC/sa12 [7]), .A3(\AES_ENC/us12/n1059 ), .ZN(\AES_ENC/us12/n636 ) );
NOR2_X2 \AES_ENC/us12/U508  ( .A1(\AES_ENC/sa12 [7]), .A2(\AES_ENC/sa12 [2]),.ZN(\AES_ENC/us12/n794 ) );
NOR2_X2 \AES_ENC/us12/U507  ( .A1(\AES_ENC/sa12 [4]), .A2(\AES_ENC/sa12 [1]),.ZN(\AES_ENC/us12/n1102 ) );
NOR2_X2 \AES_ENC/us12/U506  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/sa12 [3]), .ZN(\AES_ENC/us12/n1053 ) );
NOR2_X2 \AES_ENC/us12/U505  ( .A1(\AES_ENC/us12/n607 ), .A2(\AES_ENC/sa12 [5]), .ZN(\AES_ENC/us12/n1024 ) );
NOR2_X2 \AES_ENC/us12/U504  ( .A1(\AES_ENC/us12/n625 ), .A2(\AES_ENC/sa12 [2]), .ZN(\AES_ENC/us12/n1093 ) );
NOR2_X2 \AES_ENC/us12/U503  ( .A1(\AES_ENC/us12/n614 ), .A2(\AES_ENC/sa12 [5]), .ZN(\AES_ENC/us12/n1094 ) );
NOR2_X2 \AES_ENC/us12/U502  ( .A1(\AES_ENC/us12/n624 ), .A2(\AES_ENC/sa12 [3]), .ZN(\AES_ENC/us12/n931 ) );
INV_X4 \AES_ENC/us12/U501  ( .A(\AES_ENC/us12/n570 ), .ZN(\AES_ENC/us12/n573 ) );
NOR2_X2 \AES_ENC/us12/U500  ( .A1(\AES_ENC/us12/n1053 ), .A2(\AES_ENC/us12/n1095 ), .ZN(\AES_ENC/us12/n639 ) );
NOR3_X2 \AES_ENC/us12/U499  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n573 ), .A3(\AES_ENC/us12/n1074 ), .ZN(\AES_ENC/us12/n641 ) );
NOR2_X2 \AES_ENC/us12/U498  ( .A1(\AES_ENC/us12/n639 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n640 ) );
NOR2_X2 \AES_ENC/us12/U497  ( .A1(\AES_ENC/us12/n641 ), .A2(\AES_ENC/us12/n640 ), .ZN(\AES_ENC/us12/n646 ) );
NOR3_X2 \AES_ENC/us12/U496  ( .A1(\AES_ENC/us12/n995 ), .A2(\AES_ENC/us12/n586 ), .A3(\AES_ENC/us12/n994 ), .ZN(\AES_ENC/us12/n1002 ) );
NOR2_X2 \AES_ENC/us12/U495  ( .A1(\AES_ENC/us12/n909 ), .A2(\AES_ENC/us12/n908 ), .ZN(\AES_ENC/us12/n920 ) );
NOR2_X2 \AES_ENC/us12/U494  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n823 ) );
NOR2_X2 \AES_ENC/us12/U492  ( .A1(\AES_ENC/us12/n624 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n822 ) );
NOR2_X2 \AES_ENC/us12/U491  ( .A1(\AES_ENC/us12/n823 ), .A2(\AES_ENC/us12/n822 ), .ZN(\AES_ENC/us12/n825 ) );
NOR2_X2 \AES_ENC/us12/U490  ( .A1(\AES_ENC/sa12 [1]), .A2(\AES_ENC/us12/n623 ), .ZN(\AES_ENC/us12/n913 ) );
NOR2_X2 \AES_ENC/us12/U489  ( .A1(\AES_ENC/us12/n913 ), .A2(\AES_ENC/us12/n1091 ), .ZN(\AES_ENC/us12/n914 ) );
NOR2_X2 \AES_ENC/us12/U488  ( .A1(\AES_ENC/us12/n826 ), .A2(\AES_ENC/us12/n572 ), .ZN(\AES_ENC/us12/n827 ) );
NOR3_X2 \AES_ENC/us12/U487  ( .A1(\AES_ENC/us12/n769 ), .A2(\AES_ENC/us12/n768 ), .A3(\AES_ENC/us12/n767 ), .ZN(\AES_ENC/us12/n775 ) );
NOR2_X2 \AES_ENC/us12/U486  ( .A1(\AES_ENC/us12/n1056 ), .A2(\AES_ENC/us12/n1053 ), .ZN(\AES_ENC/us12/n749 ) );
NOR2_X2 \AES_ENC/us12/U483  ( .A1(\AES_ENC/us12/n749 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n752 ) );
INV_X4 \AES_ENC/us12/U482  ( .A(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n596 ));
NOR2_X2 \AES_ENC/us12/U480  ( .A1(\AES_ENC/us12/n1054 ), .A2(\AES_ENC/us12/n1053 ), .ZN(\AES_ENC/us12/n1055 ) );
OR2_X4 \AES_ENC/us12/U479  ( .A1(\AES_ENC/us12/n1094 ), .A2(\AES_ENC/us12/n1093 ), .ZN(\AES_ENC/us12/n571 ) );
AND2_X2 \AES_ENC/us12/U478  ( .A1(\AES_ENC/us12/n571 ), .A2(\AES_ENC/us12/n1095 ), .ZN(\AES_ENC/us12/n1101 ) );
NOR2_X2 \AES_ENC/us12/U477  ( .A1(\AES_ENC/us12/n1074 ), .A2(\AES_ENC/us12/n931 ), .ZN(\AES_ENC/us12/n796 ) );
NOR2_X2 \AES_ENC/us12/U474  ( .A1(\AES_ENC/us12/n796 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n797 ) );
NOR2_X2 \AES_ENC/us12/U473  ( .A1(\AES_ENC/us12/n932 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n933 ) );
NOR2_X2 \AES_ENC/us12/U472  ( .A1(\AES_ENC/us12/n929 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n935 ) );
NOR2_X2 \AES_ENC/us12/U471  ( .A1(\AES_ENC/us12/n931 ), .A2(\AES_ENC/us12/n930 ), .ZN(\AES_ENC/us12/n934 ) );
NOR3_X2 \AES_ENC/us12/U470  ( .A1(\AES_ENC/us12/n935 ), .A2(\AES_ENC/us12/n934 ), .A3(\AES_ENC/us12/n933 ), .ZN(\AES_ENC/us12/n936 ) );
NOR2_X2 \AES_ENC/us12/U469  ( .A1(\AES_ENC/us12/n624 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n1075 ) );
NOR2_X2 \AES_ENC/us12/U468  ( .A1(\AES_ENC/us12/n572 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n949 ) );
NOR2_X2 \AES_ENC/us12/U467  ( .A1(\AES_ENC/us12/n1049 ), .A2(\AES_ENC/us12/n618 ), .ZN(\AES_ENC/us12/n1051 ) );
NOR2_X2 \AES_ENC/us12/U466  ( .A1(\AES_ENC/us12/n1051 ), .A2(\AES_ENC/us12/n1050 ), .ZN(\AES_ENC/us12/n1052 ) );
NOR2_X2 \AES_ENC/us12/U465  ( .A1(\AES_ENC/us12/n1052 ), .A2(\AES_ENC/us12/n592 ), .ZN(\AES_ENC/us12/n1064 ) );
NOR2_X2 \AES_ENC/us12/U464  ( .A1(\AES_ENC/sa12 [1]), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n631 ) );
NOR2_X2 \AES_ENC/us12/U463  ( .A1(\AES_ENC/us12/n1025 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n980 ) );
NOR2_X2 \AES_ENC/us12/U462  ( .A1(\AES_ENC/us12/n1073 ), .A2(\AES_ENC/us12/n1094 ), .ZN(\AES_ENC/us12/n795 ) );
NOR2_X2 \AES_ENC/us12/U461  ( .A1(\AES_ENC/us12/n795 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n799 ) );
NOR2_X2 \AES_ENC/us12/U460  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n981 ) );
NOR2_X2 \AES_ENC/us12/U459  ( .A1(\AES_ENC/us12/n1102 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n643 ) );
NOR2_X2 \AES_ENC/us12/U458  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n621 ), .ZN(\AES_ENC/us12/n642 ) );
NOR2_X2 \AES_ENC/us12/U455  ( .A1(\AES_ENC/us12/n911 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n644 ) );
NOR4_X2 \AES_ENC/us12/U448  ( .A1(\AES_ENC/us12/n644 ), .A2(\AES_ENC/us12/n643 ), .A3(\AES_ENC/us12/n804 ), .A4(\AES_ENC/us12/n642 ), .ZN(\AES_ENC/us12/n645 ) );
NOR2_X2 \AES_ENC/us12/U447  ( .A1(\AES_ENC/us12/n1102 ), .A2(\AES_ENC/us12/n910 ), .ZN(\AES_ENC/us12/n932 ) );
NOR2_X2 \AES_ENC/us12/U442  ( .A1(\AES_ENC/us12/n1102 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n755 ) );
NOR2_X2 \AES_ENC/us12/U441  ( .A1(\AES_ENC/us12/n931 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n743 ) );
NOR2_X2 \AES_ENC/us12/U438  ( .A1(\AES_ENC/us12/n1072 ), .A2(\AES_ENC/us12/n1094 ), .ZN(\AES_ENC/us12/n930 ) );
NOR2_X2 \AES_ENC/us12/U435  ( .A1(\AES_ENC/us12/n1074 ), .A2(\AES_ENC/us12/n1025 ), .ZN(\AES_ENC/us12/n891 ) );
NOR2_X2 \AES_ENC/us12/U434  ( .A1(\AES_ENC/us12/n891 ), .A2(\AES_ENC/us12/n609 ), .ZN(\AES_ENC/us12/n894 ) );
NOR3_X2 \AES_ENC/us12/U433  ( .A1(\AES_ENC/us12/n623 ), .A2(\AES_ENC/sa12 [1]), .A3(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n683 ));
INV_X4 \AES_ENC/us12/U428  ( .A(\AES_ENC/us12/n931 ), .ZN(\AES_ENC/us12/n623 ) );
NOR2_X2 \AES_ENC/us12/U427  ( .A1(\AES_ENC/us12/n996 ), .A2(\AES_ENC/us12/n931 ), .ZN(\AES_ENC/us12/n704 ) );
NOR2_X2 \AES_ENC/us12/U421  ( .A1(\AES_ENC/us12/n931 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n685 ) );
NOR2_X2 \AES_ENC/us12/U420  ( .A1(\AES_ENC/us12/n1029 ), .A2(\AES_ENC/us12/n1025 ), .ZN(\AES_ENC/us12/n1079 ) );
NOR3_X2 \AES_ENC/us12/U419  ( .A1(\AES_ENC/us12/n589 ), .A2(\AES_ENC/us12/n1025 ), .A3(\AES_ENC/us12/n616 ), .ZN(\AES_ENC/us12/n945 ) );
NOR2_X2 \AES_ENC/us12/U418  ( .A1(\AES_ENC/us12/n626 ), .A2(\AES_ENC/us12/n611 ), .ZN(\AES_ENC/us12/n800 ) );
NOR3_X2 \AES_ENC/us12/U417  ( .A1(\AES_ENC/us12/n590 ), .A2(\AES_ENC/us12/n627 ), .A3(\AES_ENC/us12/n611 ), .ZN(\AES_ENC/us12/n798 ) );
NOR3_X2 \AES_ENC/us12/U416  ( .A1(\AES_ENC/us12/n610 ), .A2(\AES_ENC/us12/n572 ), .A3(\AES_ENC/us12/n575 ), .ZN(\AES_ENC/us12/n962 ) );
NOR3_X2 \AES_ENC/us12/U415  ( .A1(\AES_ENC/us12/n959 ), .A2(\AES_ENC/us12/n572 ), .A3(\AES_ENC/us12/n609 ), .ZN(\AES_ENC/us12/n768 ) );
NOR3_X2 \AES_ENC/us12/U414  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n572 ), .A3(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n694 ) );
NOR3_X2 \AES_ENC/us12/U413  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n572 ), .A3(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n895 ) );
NOR3_X2 \AES_ENC/us12/U410  ( .A1(\AES_ENC/us12/n1008 ), .A2(\AES_ENC/us12/n1007 ), .A3(\AES_ENC/us12/n1006 ), .ZN(\AES_ENC/us12/n1018 ) );
NOR4_X2 \AES_ENC/us12/U409  ( .A1(\AES_ENC/us12/n806 ), .A2(\AES_ENC/us12/n805 ), .A3(\AES_ENC/us12/n804 ), .A4(\AES_ENC/us12/n803 ), .ZN(\AES_ENC/us12/n807 ) );
NOR3_X2 \AES_ENC/us12/U406  ( .A1(\AES_ENC/us12/n799 ), .A2(\AES_ENC/us12/n798 ), .A3(\AES_ENC/us12/n797 ), .ZN(\AES_ENC/us12/n808 ) );
NOR4_X2 \AES_ENC/us12/U405  ( .A1(\AES_ENC/us12/n843 ), .A2(\AES_ENC/us12/n842 ), .A3(\AES_ENC/us12/n841 ), .A4(\AES_ENC/us12/n840 ), .ZN(\AES_ENC/us12/n844 ) );
NOR3_X2 \AES_ENC/us12/U404  ( .A1(\AES_ENC/us12/n1101 ), .A2(\AES_ENC/us12/n1100 ), .A3(\AES_ENC/us12/n1099 ), .ZN(\AES_ENC/us12/n1109 ) );
NOR4_X2 \AES_ENC/us12/U403  ( .A1(\AES_ENC/us12/n711 ), .A2(\AES_ENC/us12/n710 ), .A3(\AES_ENC/us12/n709 ), .A4(\AES_ENC/us12/n708 ), .ZN(\AES_ENC/us12/n712 ) );
NOR4_X2 \AES_ENC/us12/U401  ( .A1(\AES_ENC/us12/n963 ), .A2(\AES_ENC/us12/n962 ), .A3(\AES_ENC/us12/n961 ), .A4(\AES_ENC/us12/n960 ), .ZN(\AES_ENC/us12/n964 ) );
NOR2_X2 \AES_ENC/us12/U400  ( .A1(\AES_ENC/us12/n669 ), .A2(\AES_ENC/us12/n668 ), .ZN(\AES_ENC/us12/n673 ) );
NOR4_X2 \AES_ENC/us12/U399  ( .A1(\AES_ENC/us12/n946 ), .A2(\AES_ENC/us12/n1046 ), .A3(\AES_ENC/us12/n671 ), .A4(\AES_ENC/us12/n670 ), .ZN(\AES_ENC/us12/n672 ) );
NOR3_X2 \AES_ENC/us12/U398  ( .A1(\AES_ENC/us12/n743 ), .A2(\AES_ENC/us12/n742 ), .A3(\AES_ENC/us12/n741 ), .ZN(\AES_ENC/us12/n744 ) );
NOR2_X2 \AES_ENC/us12/U397  ( .A1(\AES_ENC/us12/n697 ), .A2(\AES_ENC/us12/n658 ), .ZN(\AES_ENC/us12/n659 ) );
NOR2_X2 \AES_ENC/us12/U396  ( .A1(\AES_ENC/us12/n1078 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n1033 ) );
NOR2_X2 \AES_ENC/us12/U393  ( .A1(\AES_ENC/us12/n1031 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n1032 ) );
NOR3_X2 \AES_ENC/us12/U390  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n1025 ), .A3(\AES_ENC/us12/n1074 ), .ZN(\AES_ENC/us12/n1035 ) );
NOR4_X2 \AES_ENC/us12/U389  ( .A1(\AES_ENC/us12/n1035 ), .A2(\AES_ENC/us12/n1034 ), .A3(\AES_ENC/us12/n1033 ), .A4(\AES_ENC/us12/n1032 ), .ZN(\AES_ENC/us12/n1036 ) );
NOR2_X2 \AES_ENC/us12/U388  ( .A1(\AES_ENC/us12/n598 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n885 ) );
NOR2_X2 \AES_ENC/us12/U387  ( .A1(\AES_ENC/us12/n623 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n882 ) );
NOR2_X2 \AES_ENC/us12/U386  ( .A1(\AES_ENC/us12/n1053 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n884 ) );
NOR4_X2 \AES_ENC/us12/U385  ( .A1(\AES_ENC/us12/n885 ), .A2(\AES_ENC/us12/n884 ), .A3(\AES_ENC/us12/n883 ), .A4(\AES_ENC/us12/n882 ), .ZN(\AES_ENC/us12/n886 ) );
NOR2_X2 \AES_ENC/us12/U384  ( .A1(\AES_ENC/us12/n825 ), .A2(\AES_ENC/us12/n578 ), .ZN(\AES_ENC/us12/n830 ) );
NOR2_X2 \AES_ENC/us12/U383  ( .A1(\AES_ENC/us12/n827 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n829 ) );
NOR2_X2 \AES_ENC/us12/U382  ( .A1(\AES_ENC/us12/n572 ), .A2(\AES_ENC/us12/n579 ), .ZN(\AES_ENC/us12/n828 ) );
NOR4_X2 \AES_ENC/us12/U374  ( .A1(\AES_ENC/us12/n831 ), .A2(\AES_ENC/us12/n830 ), .A3(\AES_ENC/us12/n829 ), .A4(\AES_ENC/us12/n828 ), .ZN(\AES_ENC/us12/n832 ) );
NOR2_X2 \AES_ENC/us12/U373  ( .A1(\AES_ENC/us12/n606 ), .A2(\AES_ENC/us12/n582 ), .ZN(\AES_ENC/us12/n1104 ) );
NOR2_X2 \AES_ENC/us12/U372  ( .A1(\AES_ENC/us12/n1102 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n1106 ) );
NOR2_X2 \AES_ENC/us12/U370  ( .A1(\AES_ENC/us12/n1103 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n1105 ) );
NOR4_X2 \AES_ENC/us12/U369  ( .A1(\AES_ENC/us12/n1107 ), .A2(\AES_ENC/us12/n1106 ), .A3(\AES_ENC/us12/n1105 ), .A4(\AES_ENC/us12/n1104 ), .ZN(\AES_ENC/us12/n1108 ) );
NOR3_X2 \AES_ENC/us12/U368  ( .A1(\AES_ENC/us12/n959 ), .A2(\AES_ENC/us12/n621 ), .A3(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n963 ) );
NOR2_X2 \AES_ENC/us12/U367  ( .A1(\AES_ENC/us12/n626 ), .A2(\AES_ENC/us12/n627 ), .ZN(\AES_ENC/us12/n1114 ) );
INV_X4 \AES_ENC/us12/U366  ( .A(\AES_ENC/us12/n1024 ), .ZN(\AES_ENC/us12/n606 ) );
NOR3_X2 \AES_ENC/us12/U365  ( .A1(\AES_ENC/us12/n910 ), .A2(\AES_ENC/us12/n1059 ), .A3(\AES_ENC/us12/n611 ), .ZN(\AES_ENC/us12/n1115 ) );
INV_X4 \AES_ENC/us12/U364  ( .A(\AES_ENC/us12/n1094 ), .ZN(\AES_ENC/us12/n613 ) );
NOR2_X2 \AES_ENC/us12/U363  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n931 ), .ZN(\AES_ENC/us12/n1100 ) );
INV_X4 \AES_ENC/us12/U354  ( .A(\AES_ENC/us12/n1093 ), .ZN(\AES_ENC/us12/n617 ) );
NOR2_X2 \AES_ENC/us12/U353  ( .A1(\AES_ENC/us12/n569 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n929 ) );
NOR2_X2 \AES_ENC/us12/U352  ( .A1(\AES_ENC/us12/n620 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n926 ) );
NOR2_X2 \AES_ENC/us12/U351  ( .A1(\AES_ENC/us12/n572 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n1095 ) );
NOR2_X2 \AES_ENC/us12/U350  ( .A1(\AES_ENC/us12/n609 ), .A2(\AES_ENC/us12/n627 ), .ZN(\AES_ENC/us12/n1010 ) );
NOR2_X2 \AES_ENC/us12/U349  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n1103 ) );
NOR2_X2 \AES_ENC/us12/U348  ( .A1(\AES_ENC/us12/n622 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n1059 ) );
NOR2_X2 \AES_ENC/us12/U347  ( .A1(\AES_ENC/sa12 [1]), .A2(\AES_ENC/us12/n1120 ), .ZN(\AES_ENC/us12/n1022 ) );
NOR2_X2 \AES_ENC/us12/U346  ( .A1(\AES_ENC/us12/n619 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n911 ) );
NOR2_X2 \AES_ENC/us12/U345  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/us12/n1025 ), .ZN(\AES_ENC/us12/n826 ) );
NOR2_X2 \AES_ENC/us12/U338  ( .A1(\AES_ENC/us12/n626 ), .A2(\AES_ENC/us12/n607 ), .ZN(\AES_ENC/us12/n1072 ) );
NOR2_X2 \AES_ENC/us12/U335  ( .A1(\AES_ENC/us12/n627 ), .A2(\AES_ENC/us12/n616 ), .ZN(\AES_ENC/us12/n956 ) );
NOR2_X2 \AES_ENC/us12/U329  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/us12/n624 ), .ZN(\AES_ENC/us12/n1121 ) );
NOR2_X2 \AES_ENC/us12/U328  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/us12/n624 ), .ZN(\AES_ENC/us12/n1058 ) );
NOR2_X2 \AES_ENC/us12/U327  ( .A1(\AES_ENC/us12/n625 ), .A2(\AES_ENC/us12/n611 ), .ZN(\AES_ENC/us12/n1073 ) );
NOR2_X2 \AES_ENC/us12/U325  ( .A1(\AES_ENC/sa12 [1]), .A2(\AES_ENC/us12/n1025 ), .ZN(\AES_ENC/us12/n1054 ) );
NOR2_X2 \AES_ENC/us12/U324  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/us12/n931 ), .ZN(\AES_ENC/us12/n1029 ) );
NOR2_X2 \AES_ENC/us12/U319  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n1056 ) );
NOR2_X2 \AES_ENC/us12/U318  ( .A1(\AES_ENC/us12/n614 ), .A2(\AES_ENC/us12/n626 ), .ZN(\AES_ENC/us12/n1050 ) );
NOR2_X2 \AES_ENC/us12/U317  ( .A1(\AES_ENC/us12/n1121 ), .A2(\AES_ENC/us12/n1025 ), .ZN(\AES_ENC/us12/n1120 ) );
NOR2_X2 \AES_ENC/us12/U316  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/us12/n572 ), .ZN(\AES_ENC/us12/n1074 ) );
NOR2_X2 \AES_ENC/us12/U315  ( .A1(\AES_ENC/us12/n1058 ), .A2(\AES_ENC/us12/n1054 ), .ZN(\AES_ENC/us12/n878 ) );
NOR2_X2 \AES_ENC/us12/U314  ( .A1(\AES_ENC/us12/n878 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n879 ) );
NOR2_X2 \AES_ENC/us12/U312  ( .A1(\AES_ENC/us12/n880 ), .A2(\AES_ENC/us12/n879 ), .ZN(\AES_ENC/us12/n887 ) );
NOR2_X2 \AES_ENC/us12/U311  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n588 ), .ZN(\AES_ENC/us12/n957 ) );
NOR2_X2 \AES_ENC/us12/U310  ( .A1(\AES_ENC/us12/n958 ), .A2(\AES_ENC/us12/n957 ), .ZN(\AES_ENC/us12/n965 ) );
NOR3_X2 \AES_ENC/us12/U309  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n1091 ), .A3(\AES_ENC/us12/n1022 ), .ZN(\AES_ENC/us12/n720 ) );
NOR3_X2 \AES_ENC/us12/U303  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n1054 ), .A3(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n719 ) );
NOR2_X2 \AES_ENC/us12/U302  ( .A1(\AES_ENC/us12/n720 ), .A2(\AES_ENC/us12/n719 ), .ZN(\AES_ENC/us12/n726 ) );
NOR2_X2 \AES_ENC/us12/U300  ( .A1(\AES_ENC/us12/n614 ), .A2(\AES_ENC/us12/n591 ), .ZN(\AES_ENC/us12/n865 ) );
NOR2_X2 \AES_ENC/us12/U299  ( .A1(\AES_ENC/us12/n1059 ), .A2(\AES_ENC/us12/n1058 ), .ZN(\AES_ENC/us12/n1060 ) );
NOR2_X2 \AES_ENC/us12/U298  ( .A1(\AES_ENC/us12/n1095 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n668 ) );
NOR2_X2 \AES_ENC/us12/U297  ( .A1(\AES_ENC/us12/n911 ), .A2(\AES_ENC/us12/n910 ), .ZN(\AES_ENC/us12/n912 ) );
NOR2_X2 \AES_ENC/us12/U296  ( .A1(\AES_ENC/us12/n912 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n916 ) );
NOR2_X2 \AES_ENC/us12/U295  ( .A1(\AES_ENC/us12/n826 ), .A2(\AES_ENC/us12/n573 ), .ZN(\AES_ENC/us12/n750 ) );
NOR2_X2 \AES_ENC/us12/U294  ( .A1(\AES_ENC/us12/n750 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n751 ) );
NOR2_X2 \AES_ENC/us12/U293  ( .A1(\AES_ENC/us12/n907 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n908 ) );
NOR2_X2 \AES_ENC/us12/U292  ( .A1(\AES_ENC/us12/n990 ), .A2(\AES_ENC/us12/n926 ), .ZN(\AES_ENC/us12/n780 ) );
NOR2_X2 \AES_ENC/us12/U291  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n584 ), .ZN(\AES_ENC/us12/n838 ) );
NOR2_X2 \AES_ENC/us12/U290  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n602 ), .ZN(\AES_ENC/us12/n837 ) );
NOR2_X2 \AES_ENC/us12/U284  ( .A1(\AES_ENC/us12/n838 ), .A2(\AES_ENC/us12/n837 ), .ZN(\AES_ENC/us12/n845 ) );
NOR2_X2 \AES_ENC/us12/U283  ( .A1(\AES_ENC/us12/n1022 ), .A2(\AES_ENC/us12/n1058 ), .ZN(\AES_ENC/us12/n740 ) );
NOR2_X2 \AES_ENC/us12/U282  ( .A1(\AES_ENC/us12/n740 ), .A2(\AES_ENC/us12/n616 ), .ZN(\AES_ENC/us12/n742 ) );
NOR2_X2 \AES_ENC/us12/U281  ( .A1(\AES_ENC/us12/n1098 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n1099 ) );
NOR2_X2 \AES_ENC/us12/U280  ( .A1(\AES_ENC/us12/n1120 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n993 ) );
NOR2_X2 \AES_ENC/us12/U279  ( .A1(\AES_ENC/us12/n993 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n994 ) );
NOR2_X2 \AES_ENC/us12/U273  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n620 ), .ZN(\AES_ENC/us12/n1026 ) );
NOR2_X2 \AES_ENC/us12/U272  ( .A1(\AES_ENC/us12/n573 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n1027 ) );
NOR2_X2 \AES_ENC/us12/U271  ( .A1(\AES_ENC/us12/n1027 ), .A2(\AES_ENC/us12/n1026 ), .ZN(\AES_ENC/us12/n1028 ) );
NOR2_X2 \AES_ENC/us12/U270  ( .A1(\AES_ENC/us12/n1029 ), .A2(\AES_ENC/us12/n1028 ), .ZN(\AES_ENC/us12/n1034 ) );
NOR4_X2 \AES_ENC/us12/U269  ( .A1(\AES_ENC/us12/n757 ), .A2(\AES_ENC/us12/n756 ), .A3(\AES_ENC/us12/n755 ), .A4(\AES_ENC/us12/n754 ), .ZN(\AES_ENC/us12/n758 ) );
NOR2_X2 \AES_ENC/us12/U268  ( .A1(\AES_ENC/us12/n752 ), .A2(\AES_ENC/us12/n751 ), .ZN(\AES_ENC/us12/n759 ) );
NOR2_X2 \AES_ENC/us12/U267  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n1071 ), .ZN(\AES_ENC/us12/n669 ) );
NOR2_X2 \AES_ENC/us12/U263  ( .A1(\AES_ENC/us12/n1056 ), .A2(\AES_ENC/us12/n990 ), .ZN(\AES_ENC/us12/n991 ) );
NOR2_X2 \AES_ENC/us12/U262  ( .A1(\AES_ENC/us12/n991 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n995 ) );
NOR2_X2 \AES_ENC/us12/U258  ( .A1(\AES_ENC/us12/n607 ), .A2(\AES_ENC/us12/n590 ), .ZN(\AES_ENC/us12/n1008 ) );
NOR2_X2 \AES_ENC/us12/U255  ( .A1(\AES_ENC/us12/n839 ), .A2(\AES_ENC/us12/n582 ), .ZN(\AES_ENC/us12/n693 ) );
NOR2_X2 \AES_ENC/us12/U254  ( .A1(\AES_ENC/us12/n606 ), .A2(\AES_ENC/us12/n906 ), .ZN(\AES_ENC/us12/n741 ) );
NOR2_X2 \AES_ENC/us12/U253  ( .A1(\AES_ENC/us12/n1054 ), .A2(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n763 ) );
NOR2_X2 \AES_ENC/us12/U252  ( .A1(\AES_ENC/us12/n763 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n769 ) );
NOR2_X2 \AES_ENC/us12/U251  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n577 ), .ZN(\AES_ENC/us12/n1007 ) );
NOR2_X2 \AES_ENC/us12/U250  ( .A1(\AES_ENC/us12/n609 ), .A2(\AES_ENC/us12/n580 ), .ZN(\AES_ENC/us12/n1123 ) );
NOR2_X2 \AES_ENC/us12/U243  ( .A1(\AES_ENC/us12/n609 ), .A2(\AES_ENC/us12/n590 ), .ZN(\AES_ENC/us12/n710 ) );
INV_X4 \AES_ENC/us12/U242  ( .A(\AES_ENC/us12/n1029 ), .ZN(\AES_ENC/us12/n582 ) );
NOR2_X2 \AES_ENC/us12/U241  ( .A1(\AES_ENC/us12/n616 ), .A2(\AES_ENC/us12/n597 ), .ZN(\AES_ENC/us12/n883 ) );
NOR2_X2 \AES_ENC/us12/U240  ( .A1(\AES_ENC/us12/n593 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n1125 ) );
NOR2_X2 \AES_ENC/us12/U239  ( .A1(\AES_ENC/us12/n990 ), .A2(\AES_ENC/us12/n929 ), .ZN(\AES_ENC/us12/n892 ) );
NOR2_X2 \AES_ENC/us12/U238  ( .A1(\AES_ENC/us12/n892 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n893 ) );
NOR2_X2 \AES_ENC/us12/U237  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n602 ), .ZN(\AES_ENC/us12/n950 ) );
NOR2_X2 \AES_ENC/us12/U236  ( .A1(\AES_ENC/us12/n1079 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n1082 ) );
NOR2_X2 \AES_ENC/us12/U235  ( .A1(\AES_ENC/us12/n910 ), .A2(\AES_ENC/us12/n1056 ), .ZN(\AES_ENC/us12/n941 ) );
NOR2_X2 \AES_ENC/us12/U234  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n1077 ), .ZN(\AES_ENC/us12/n841 ) );
NOR2_X2 \AES_ENC/us12/U229  ( .A1(\AES_ENC/us12/n623 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n630 ) );
NOR2_X2 \AES_ENC/us12/U228  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n602 ), .ZN(\AES_ENC/us12/n806 ) );
NOR2_X2 \AES_ENC/us12/U227  ( .A1(\AES_ENC/us12/n623 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n948 ) );
NOR2_X2 \AES_ENC/us12/U226  ( .A1(\AES_ENC/us12/n606 ), .A2(\AES_ENC/us12/n589 ), .ZN(\AES_ENC/us12/n997 ) );
NOR2_X2 \AES_ENC/us12/U225  ( .A1(\AES_ENC/us12/n1121 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n1122 ) );
NOR2_X2 \AES_ENC/us12/U223  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n1023 ), .ZN(\AES_ENC/us12/n756 ) );
NOR2_X2 \AES_ENC/us12/U222  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n602 ), .ZN(\AES_ENC/us12/n870 ) );
NOR2_X2 \AES_ENC/us12/U221  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n569 ), .ZN(\AES_ENC/us12/n947 ) );
NOR2_X2 \AES_ENC/us12/U217  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n1077 ), .ZN(\AES_ENC/us12/n1084 ) );
NOR2_X2 \AES_ENC/us12/U213  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n855 ), .ZN(\AES_ENC/us12/n709 ) );
NOR2_X2 \AES_ENC/us12/U212  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n589 ), .ZN(\AES_ENC/us12/n868 ) );
NOR2_X2 \AES_ENC/us12/U211  ( .A1(\AES_ENC/us12/n1120 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n1124 ) );
NOR2_X2 \AES_ENC/us12/U210  ( .A1(\AES_ENC/us12/n1120 ), .A2(\AES_ENC/us12/n839 ), .ZN(\AES_ENC/us12/n842 ) );
NOR2_X2 \AES_ENC/us12/U209  ( .A1(\AES_ENC/us12/n1120 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n696 ) );
NOR2_X2 \AES_ENC/us12/U208  ( .A1(\AES_ENC/us12/n1074 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n1076 ) );
NOR2_X2 \AES_ENC/us12/U207  ( .A1(\AES_ENC/us12/n1074 ), .A2(\AES_ENC/us12/n620 ), .ZN(\AES_ENC/us12/n781 ) );
NOR3_X2 \AES_ENC/us12/U201  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n1056 ), .A3(\AES_ENC/us12/n990 ), .ZN(\AES_ENC/us12/n979 ) );
NOR3_X2 \AES_ENC/us12/U200  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n1058 ), .A3(\AES_ENC/us12/n1059 ), .ZN(\AES_ENC/us12/n854 ) );
NOR2_X2 \AES_ENC/us12/U199  ( .A1(\AES_ENC/us12/n996 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n869 ) );
NOR2_X2 \AES_ENC/us12/U198  ( .A1(\AES_ENC/us12/n1056 ), .A2(\AES_ENC/us12/n1074 ), .ZN(\AES_ENC/us12/n1057 ) );
NOR3_X2 \AES_ENC/us12/U197  ( .A1(\AES_ENC/us12/n607 ), .A2(\AES_ENC/us12/n1120 ), .A3(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n978 ) );
NOR2_X2 \AES_ENC/us12/U196  ( .A1(\AES_ENC/us12/n996 ), .A2(\AES_ENC/us12/n911 ), .ZN(\AES_ENC/us12/n1116 ) );
NOR2_X2 \AES_ENC/us12/U195  ( .A1(\AES_ENC/us12/n1074 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n754 ) );
NOR2_X2 \AES_ENC/us12/U194  ( .A1(\AES_ENC/us12/n926 ), .A2(\AES_ENC/us12/n1103 ), .ZN(\AES_ENC/us12/n977 ) );
NOR2_X2 \AES_ENC/us12/U187  ( .A1(\AES_ENC/us12/n839 ), .A2(\AES_ENC/us12/n824 ), .ZN(\AES_ENC/us12/n1092 ) );
NOR2_X2 \AES_ENC/us12/U186  ( .A1(\AES_ENC/us12/n573 ), .A2(\AES_ENC/us12/n1074 ), .ZN(\AES_ENC/us12/n684 ) );
NOR2_X2 \AES_ENC/us12/U185  ( .A1(\AES_ENC/us12/n826 ), .A2(\AES_ENC/us12/n1059 ), .ZN(\AES_ENC/us12/n907 ) );
NOR3_X2 \AES_ENC/us12/U184  ( .A1(\AES_ENC/us12/n625 ), .A2(\AES_ENC/us12/n1115 ), .A3(\AES_ENC/us12/n585 ), .ZN(\AES_ENC/us12/n831 ) );
NOR3_X2 \AES_ENC/us12/U183  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n1056 ), .A3(\AES_ENC/us12/n990 ), .ZN(\AES_ENC/us12/n896 ) );
NOR3_X2 \AES_ENC/us12/U182  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n573 ), .A3(\AES_ENC/us12/n1013 ), .ZN(\AES_ENC/us12/n670 ) );
NOR3_X2 \AES_ENC/us12/U181  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n1091 ), .A3(\AES_ENC/us12/n1022 ), .ZN(\AES_ENC/us12/n843 ) );
NOR2_X2 \AES_ENC/us12/U180  ( .A1(\AES_ENC/us12/n1029 ), .A2(\AES_ENC/us12/n1095 ), .ZN(\AES_ENC/us12/n735 ) );
NOR2_X2 \AES_ENC/us12/U174  ( .A1(\AES_ENC/us12/n1100 ), .A2(\AES_ENC/us12/n854 ), .ZN(\AES_ENC/us12/n860 ) );
NOR4_X2 \AES_ENC/us12/U173  ( .A1(\AES_ENC/us12/n1125 ), .A2(\AES_ENC/us12/n1124 ), .A3(\AES_ENC/us12/n1123 ), .A4(\AES_ENC/us12/n1122 ), .ZN(\AES_ENC/us12/n1126 ) );
NOR4_X2 \AES_ENC/us12/U172  ( .A1(\AES_ENC/us12/n1084 ), .A2(\AES_ENC/us12/n1083 ), .A3(\AES_ENC/us12/n1082 ), .A4(\AES_ENC/us12/n1081 ), .ZN(\AES_ENC/us12/n1085 ) );
NOR2_X2 \AES_ENC/us12/U171  ( .A1(\AES_ENC/us12/n1076 ), .A2(\AES_ENC/us12/n1075 ), .ZN(\AES_ENC/us12/n1086 ) );
NAND3_X2 \AES_ENC/us12/U170  ( .A1(\AES_ENC/us12/n569 ), .A2(\AES_ENC/us12/n582 ), .A3(\AES_ENC/us12/n681 ), .ZN(\AES_ENC/us12/n691 ) );
NOR2_X2 \AES_ENC/us12/U169  ( .A1(\AES_ENC/us12/n683 ), .A2(\AES_ENC/us12/n682 ), .ZN(\AES_ENC/us12/n690 ) );
NOR3_X2 \AES_ENC/us12/U168  ( .A1(\AES_ENC/us12/n695 ), .A2(\AES_ENC/us12/n694 ), .A3(\AES_ENC/us12/n693 ), .ZN(\AES_ENC/us12/n700 ) );
NOR4_X2 \AES_ENC/us12/U162  ( .A1(\AES_ENC/us12/n983 ), .A2(\AES_ENC/us12/n698 ), .A3(\AES_ENC/us12/n697 ), .A4(\AES_ENC/us12/n696 ), .ZN(\AES_ENC/us12/n699 ) );
NOR2_X2 \AES_ENC/us12/U161  ( .A1(\AES_ENC/us12/n946 ), .A2(\AES_ENC/us12/n945 ), .ZN(\AES_ENC/us12/n952 ) );
NOR4_X2 \AES_ENC/us12/U160  ( .A1(\AES_ENC/us12/n950 ), .A2(\AES_ENC/us12/n949 ), .A3(\AES_ENC/us12/n948 ), .A4(\AES_ENC/us12/n947 ), .ZN(\AES_ENC/us12/n951 ) );
NOR4_X2 \AES_ENC/us12/U159  ( .A1(\AES_ENC/us12/n983 ), .A2(\AES_ENC/us12/n982 ), .A3(\AES_ENC/us12/n981 ), .A4(\AES_ENC/us12/n980 ), .ZN(\AES_ENC/us12/n984 ) );
NOR2_X2 \AES_ENC/us12/U158  ( .A1(\AES_ENC/us12/n979 ), .A2(\AES_ENC/us12/n978 ), .ZN(\AES_ENC/us12/n985 ) );
NOR4_X2 \AES_ENC/us12/U157  ( .A1(\AES_ENC/us12/n896 ), .A2(\AES_ENC/us12/n895 ), .A3(\AES_ENC/us12/n894 ), .A4(\AES_ENC/us12/n893 ), .ZN(\AES_ENC/us12/n897 ) );
NOR2_X2 \AES_ENC/us12/U156  ( .A1(\AES_ENC/us12/n866 ), .A2(\AES_ENC/us12/n865 ), .ZN(\AES_ENC/us12/n872 ) );
NOR4_X2 \AES_ENC/us12/U155  ( .A1(\AES_ENC/us12/n870 ), .A2(\AES_ENC/us12/n869 ), .A3(\AES_ENC/us12/n868 ), .A4(\AES_ENC/us12/n867 ), .ZN(\AES_ENC/us12/n871 ) );
NOR3_X2 \AES_ENC/us12/U154  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n1054 ), .A3(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n961 ) );
NOR3_X2 \AES_ENC/us12/U153  ( .A1(\AES_ENC/us12/n620 ), .A2(\AES_ENC/us12/n1074 ), .A3(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n671 ) );
NOR2_X2 \AES_ENC/us12/U152  ( .A1(\AES_ENC/us12/n1057 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n1062 ) );
NOR2_X2 \AES_ENC/us12/U143  ( .A1(\AES_ENC/us12/n1055 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n1063 ) );
NOR2_X2 \AES_ENC/us12/U142  ( .A1(\AES_ENC/us12/n1060 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n1061 ) );
NOR4_X2 \AES_ENC/us12/U141  ( .A1(\AES_ENC/us12/n1064 ), .A2(\AES_ENC/us12/n1063 ), .A3(\AES_ENC/us12/n1062 ), .A4(\AES_ENC/us12/n1061 ), .ZN(\AES_ENC/us12/n1065 ) );
NOR3_X2 \AES_ENC/us12/U140  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n1120 ), .A3(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n918 ) );
NOR3_X2 \AES_ENC/us12/U132  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n573 ), .A3(\AES_ENC/us12/n1013 ), .ZN(\AES_ENC/us12/n917 ) );
NOR2_X2 \AES_ENC/us12/U131  ( .A1(\AES_ENC/us12/n914 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n915 ) );
NOR4_X2 \AES_ENC/us12/U130  ( .A1(\AES_ENC/us12/n918 ), .A2(\AES_ENC/us12/n917 ), .A3(\AES_ENC/us12/n916 ), .A4(\AES_ENC/us12/n915 ), .ZN(\AES_ENC/us12/n919 ) );
NOR2_X2 \AES_ENC/us12/U129  ( .A1(\AES_ENC/us12/n616 ), .A2(\AES_ENC/us12/n580 ), .ZN(\AES_ENC/us12/n771 ) );
NOR2_X2 \AES_ENC/us12/U128  ( .A1(\AES_ENC/us12/n1103 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n772 ) );
NOR2_X2 \AES_ENC/us12/U127  ( .A1(\AES_ENC/us12/n610 ), .A2(\AES_ENC/us12/n599 ), .ZN(\AES_ENC/us12/n773 ) );
NOR4_X2 \AES_ENC/us12/U126  ( .A1(\AES_ENC/us12/n773 ), .A2(\AES_ENC/us12/n772 ), .A3(\AES_ENC/us12/n771 ), .A4(\AES_ENC/us12/n770 ), .ZN(\AES_ENC/us12/n774 ) );
NOR2_X2 \AES_ENC/us12/U121  ( .A1(\AES_ENC/us12/n735 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n687 ) );
NOR2_X2 \AES_ENC/us12/U120  ( .A1(\AES_ENC/us12/n684 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n688 ) );
NOR2_X2 \AES_ENC/us12/U119  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n600 ), .ZN(\AES_ENC/us12/n686 ) );
NOR4_X2 \AES_ENC/us12/U118  ( .A1(\AES_ENC/us12/n688 ), .A2(\AES_ENC/us12/n687 ), .A3(\AES_ENC/us12/n686 ), .A4(\AES_ENC/us12/n685 ), .ZN(\AES_ENC/us12/n689 ) );
NOR2_X2 \AES_ENC/us12/U117  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n595 ), .ZN(\AES_ENC/us12/n858 ) );
NOR2_X2 \AES_ENC/us12/U116  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n855 ), .ZN(\AES_ENC/us12/n857 ) );
NOR2_X2 \AES_ENC/us12/U115  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n587 ), .ZN(\AES_ENC/us12/n856 ) );
NOR4_X2 \AES_ENC/us12/U106  ( .A1(\AES_ENC/us12/n858 ), .A2(\AES_ENC/us12/n857 ), .A3(\AES_ENC/us12/n856 ), .A4(\AES_ENC/us12/n958 ), .ZN(\AES_ENC/us12/n859 ) );
NOR2_X2 \AES_ENC/us12/U105  ( .A1(\AES_ENC/us12/n780 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n784 ) );
NOR2_X2 \AES_ENC/us12/U104  ( .A1(\AES_ENC/us12/n1117 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n782 ) );
NOR2_X2 \AES_ENC/us12/U103  ( .A1(\AES_ENC/us12/n781 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n783 ) );
NOR4_X2 \AES_ENC/us12/U102  ( .A1(\AES_ENC/us12/n880 ), .A2(\AES_ENC/us12/n784 ), .A3(\AES_ENC/us12/n783 ), .A4(\AES_ENC/us12/n782 ), .ZN(\AES_ENC/us12/n785 ) );
NOR2_X2 \AES_ENC/us12/U101  ( .A1(\AES_ENC/us12/n583 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n814 ) );
NOR2_X2 \AES_ENC/us12/U100  ( .A1(\AES_ENC/us12/n907 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n813 ) );
NOR3_X2 \AES_ENC/us12/U95  ( .A1(\AES_ENC/us12/n606 ), .A2(\AES_ENC/us12/n1058 ), .A3(\AES_ENC/us12/n1059 ), .ZN(\AES_ENC/us12/n815 ) );
NOR4_X2 \AES_ENC/us12/U94  ( .A1(\AES_ENC/us12/n815 ), .A2(\AES_ENC/us12/n814 ), .A3(\AES_ENC/us12/n813 ), .A4(\AES_ENC/us12/n812 ), .ZN(\AES_ENC/us12/n816 ) );
NOR2_X2 \AES_ENC/us12/U93  ( .A1(\AES_ENC/us12/n617 ), .A2(\AES_ENC/us12/n569 ), .ZN(\AES_ENC/us12/n721 ) );
NOR2_X2 \AES_ENC/us12/U92  ( .A1(\AES_ENC/us12/n1031 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n723 ) );
NOR2_X2 \AES_ENC/us12/U91  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n1096 ), .ZN(\AES_ENC/us12/n722 ) );
NOR4_X2 \AES_ENC/us12/U90  ( .A1(\AES_ENC/us12/n724 ), .A2(\AES_ENC/us12/n723 ), .A3(\AES_ENC/us12/n722 ), .A4(\AES_ENC/us12/n721 ), .ZN(\AES_ENC/us12/n725 ) );
NOR2_X2 \AES_ENC/us12/U89  ( .A1(\AES_ENC/us12/n911 ), .A2(\AES_ENC/us12/n990 ), .ZN(\AES_ENC/us12/n1009 ) );
NOR2_X2 \AES_ENC/us12/U88  ( .A1(\AES_ENC/us12/n1013 ), .A2(\AES_ENC/us12/n573 ), .ZN(\AES_ENC/us12/n1014 ) );
NOR2_X2 \AES_ENC/us12/U87  ( .A1(\AES_ENC/us12/n1014 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n1015 ) );
NOR4_X2 \AES_ENC/us12/U86  ( .A1(\AES_ENC/us12/n1016 ), .A2(\AES_ENC/us12/n1015 ), .A3(\AES_ENC/us12/n1119 ), .A4(\AES_ENC/us12/n1046 ), .ZN(\AES_ENC/us12/n1017 ) );
NOR2_X2 \AES_ENC/us12/U81  ( .A1(\AES_ENC/us12/n996 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n998 ) );
NOR2_X2 \AES_ENC/us12/U80  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n577 ), .ZN(\AES_ENC/us12/n1000 ) );
NOR2_X2 \AES_ENC/us12/U79  ( .A1(\AES_ENC/us12/n616 ), .A2(\AES_ENC/us12/n1096 ), .ZN(\AES_ENC/us12/n999 ) );
NOR4_X2 \AES_ENC/us12/U78  ( .A1(\AES_ENC/us12/n1000 ), .A2(\AES_ENC/us12/n999 ), .A3(\AES_ENC/us12/n998 ), .A4(\AES_ENC/us12/n997 ), .ZN(\AES_ENC/us12/n1001 ) );
NOR2_X2 \AES_ENC/us12/U74  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n1096 ), .ZN(\AES_ENC/us12/n697 ) );
NOR2_X2 \AES_ENC/us12/U73  ( .A1(\AES_ENC/us12/n620 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n958 ) );
NOR2_X2 \AES_ENC/us12/U72  ( .A1(\AES_ENC/us12/n911 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n983 ) );
NOR2_X2 \AES_ENC/us12/U71  ( .A1(\AES_ENC/us12/n1054 ), .A2(\AES_ENC/us12/n1103 ), .ZN(\AES_ENC/us12/n1031 ) );
INV_X4 \AES_ENC/us12/U65  ( .A(\AES_ENC/us12/n1050 ), .ZN(\AES_ENC/us12/n612 ) );
INV_X4 \AES_ENC/us12/U64  ( .A(\AES_ENC/us12/n1072 ), .ZN(\AES_ENC/us12/n605 ) );
INV_X4 \AES_ENC/us12/U63  ( .A(\AES_ENC/us12/n1073 ), .ZN(\AES_ENC/us12/n604 ) );
NOR2_X2 \AES_ENC/us12/U62  ( .A1(\AES_ENC/us12/n582 ), .A2(\AES_ENC/us12/n613 ), .ZN(\AES_ENC/us12/n880 ) );
NOR3_X2 \AES_ENC/us12/U61  ( .A1(\AES_ENC/us12/n826 ), .A2(\AES_ENC/us12/n1121 ), .A3(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n946 ) );
INV_X4 \AES_ENC/us12/U59  ( .A(\AES_ENC/us12/n1010 ), .ZN(\AES_ENC/us12/n608 ) );
NOR3_X2 \AES_ENC/us12/U58  ( .A1(\AES_ENC/us12/n573 ), .A2(\AES_ENC/us12/n1029 ), .A3(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n1119 ) );
INV_X4 \AES_ENC/us12/U57  ( .A(\AES_ENC/us12/n956 ), .ZN(\AES_ENC/us12/n615 ) );
NOR2_X2 \AES_ENC/us12/U50  ( .A1(\AES_ENC/us12/n623 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n1013 ) );
NOR2_X2 \AES_ENC/us12/U49  ( .A1(\AES_ENC/us12/n620 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n910 ) );
NOR2_X2 \AES_ENC/us12/U48  ( .A1(\AES_ENC/us12/n569 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n1091 ) );
NOR2_X2 \AES_ENC/us12/U47  ( .A1(\AES_ENC/us12/n622 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n990 ) );
NOR2_X2 \AES_ENC/us12/U46  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/us12/n1121 ), .ZN(\AES_ENC/us12/n996 ) );
NOR2_X2 \AES_ENC/us12/U45  ( .A1(\AES_ENC/us12/n610 ), .A2(\AES_ENC/us12/n600 ), .ZN(\AES_ENC/us12/n628 ) );
NOR2_X2 \AES_ENC/us12/U44  ( .A1(\AES_ENC/us12/n576 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n866 ) );
NOR2_X2 \AES_ENC/us12/U43  ( .A1(\AES_ENC/us12/n603 ), .A2(\AES_ENC/us12/n610 ), .ZN(\AES_ENC/us12/n1006 ) );
NOR2_X2 \AES_ENC/us12/U42  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n1117 ), .ZN(\AES_ENC/us12/n1118 ) );
NOR2_X2 \AES_ENC/us12/U41  ( .A1(\AES_ENC/us12/n1119 ), .A2(\AES_ENC/us12/n1118 ), .ZN(\AES_ENC/us12/n1127 ) );
NOR2_X2 \AES_ENC/us12/U36  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n906 ), .ZN(\AES_ENC/us12/n909 ) );
NOR2_X2 \AES_ENC/us12/U35  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n594 ), .ZN(\AES_ENC/us12/n629 ) );
NOR2_X2 \AES_ENC/us12/U34  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n597 ), .ZN(\AES_ENC/us12/n658 ) );
NOR2_X2 \AES_ENC/us12/U33  ( .A1(\AES_ENC/us12/n1116 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n695 ) );
NOR2_X2 \AES_ENC/us12/U32  ( .A1(\AES_ENC/us12/n1078 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n1083 ) );
NOR2_X2 \AES_ENC/us12/U31  ( .A1(\AES_ENC/us12/n941 ), .A2(\AES_ENC/us12/n608 ), .ZN(\AES_ENC/us12/n724 ) );
NOR2_X2 \AES_ENC/us12/U30  ( .A1(\AES_ENC/us12/n598 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n1107 ) );
NOR2_X2 \AES_ENC/us12/U29  ( .A1(\AES_ENC/us12/n576 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n840 ) );
NOR2_X2 \AES_ENC/us12/U24  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n593 ), .ZN(\AES_ENC/us12/n633 ) );
NOR2_X2 \AES_ENC/us12/U23  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n1080 ), .ZN(\AES_ENC/us12/n1081 ) );
NOR2_X2 \AES_ENC/us12/U21  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n1045 ), .ZN(\AES_ENC/us12/n812 ) );
NOR2_X2 \AES_ENC/us12/U20  ( .A1(\AES_ENC/us12/n1009 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n960 ) );
NOR2_X2 \AES_ENC/us12/U19  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n601 ), .ZN(\AES_ENC/us12/n982 ) );
NOR2_X2 \AES_ENC/us12/U18  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n594 ), .ZN(\AES_ENC/us12/n757 ) );
NOR2_X2 \AES_ENC/us12/U17  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n590 ), .ZN(\AES_ENC/us12/n698 ) );
NOR2_X2 \AES_ENC/us12/U16  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n619 ), .ZN(\AES_ENC/us12/n708 ) );
NOR2_X2 \AES_ENC/us12/U15  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n582 ), .ZN(\AES_ENC/us12/n770 ) );
NOR2_X2 \AES_ENC/us12/U10  ( .A1(\AES_ENC/us12/n619 ), .A2(\AES_ENC/us12/n604 ), .ZN(\AES_ENC/us12/n803 ) );
NOR2_X2 \AES_ENC/us12/U9  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n881 ), .ZN(\AES_ENC/us12/n711 ) );
NOR2_X2 \AES_ENC/us12/U8  ( .A1(\AES_ENC/us12/n615 ), .A2(\AES_ENC/us12/n582 ), .ZN(\AES_ENC/us12/n867 ) );
NOR2_X2 \AES_ENC/us12/U7  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n599 ), .ZN(\AES_ENC/us12/n804 ) );
NOR2_X2 \AES_ENC/us12/U6  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n620 ), .ZN(\AES_ENC/us12/n1046 ) );
OR2_X4 \AES_ENC/us12/U5  ( .A1(\AES_ENC/us12/n624 ), .A2(\AES_ENC/sa12 [1]),.ZN(\AES_ENC/us12/n570 ) );
OR2_X4 \AES_ENC/us12/U4  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/sa12 [4]),.ZN(\AES_ENC/us12/n569 ) );
NAND2_X2 \AES_ENC/us12/U514  ( .A1(\AES_ENC/us12/n1121 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n1030 ) );
AND2_X2 \AES_ENC/us12/U513  ( .A1(\AES_ENC/us12/n597 ), .A2(\AES_ENC/us12/n1030 ), .ZN(\AES_ENC/us12/n1049 ) );
NAND2_X2 \AES_ENC/us12/U511  ( .A1(\AES_ENC/us12/n1049 ), .A2(\AES_ENC/us12/n794 ), .ZN(\AES_ENC/us12/n637 ) );
AND2_X2 \AES_ENC/us12/U493  ( .A1(\AES_ENC/us12/n779 ), .A2(\AES_ENC/us12/n996 ), .ZN(\AES_ENC/us12/n632 ) );
NAND4_X2 \AES_ENC/us12/U485  ( .A1(\AES_ENC/us12/n637 ), .A2(\AES_ENC/us12/n636 ), .A3(\AES_ENC/us12/n635 ), .A4(\AES_ENC/us12/n634 ), .ZN(\AES_ENC/us12/n638 ) );
NAND2_X2 \AES_ENC/us12/U484  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n638 ), .ZN(\AES_ENC/us12/n679 ) );
NAND2_X2 \AES_ENC/us12/U481  ( .A1(\AES_ENC/us12/n1094 ), .A2(\AES_ENC/us12/n591 ), .ZN(\AES_ENC/us12/n648 ) );
NAND2_X2 \AES_ENC/us12/U476  ( .A1(\AES_ENC/us12/n601 ), .A2(\AES_ENC/us12/n590 ), .ZN(\AES_ENC/us12/n762 ) );
NAND2_X2 \AES_ENC/us12/U475  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n762 ), .ZN(\AES_ENC/us12/n647 ) );
NAND4_X2 \AES_ENC/us12/U457  ( .A1(\AES_ENC/us12/n648 ), .A2(\AES_ENC/us12/n647 ), .A3(\AES_ENC/us12/n646 ), .A4(\AES_ENC/us12/n645 ), .ZN(\AES_ENC/us12/n649 ) );
NAND2_X2 \AES_ENC/us12/U456  ( .A1(\AES_ENC/sa12 [0]), .A2(\AES_ENC/us12/n649 ), .ZN(\AES_ENC/us12/n665 ) );
NAND2_X2 \AES_ENC/us12/U454  ( .A1(\AES_ENC/us12/n596 ), .A2(\AES_ENC/us12/n623 ), .ZN(\AES_ENC/us12/n855 ) );
NAND2_X2 \AES_ENC/us12/U453  ( .A1(\AES_ENC/us12/n587 ), .A2(\AES_ENC/us12/n855 ), .ZN(\AES_ENC/us12/n821 ) );
NAND2_X2 \AES_ENC/us12/U452  ( .A1(\AES_ENC/us12/n1093 ), .A2(\AES_ENC/us12/n821 ), .ZN(\AES_ENC/us12/n662 ) );
NAND2_X2 \AES_ENC/us12/U451  ( .A1(\AES_ENC/us12/n619 ), .A2(\AES_ENC/us12/n589 ), .ZN(\AES_ENC/us12/n650 ) );
NAND2_X2 \AES_ENC/us12/U450  ( .A1(\AES_ENC/us12/n956 ), .A2(\AES_ENC/us12/n650 ), .ZN(\AES_ENC/us12/n661 ) );
NAND2_X2 \AES_ENC/us12/U449  ( .A1(\AES_ENC/us12/n626 ), .A2(\AES_ENC/us12/n627 ), .ZN(\AES_ENC/us12/n839 ) );
OR2_X2 \AES_ENC/us12/U446  ( .A1(\AES_ENC/us12/n839 ), .A2(\AES_ENC/us12/n932 ), .ZN(\AES_ENC/us12/n656 ) );
NAND2_X2 \AES_ENC/us12/U445  ( .A1(\AES_ENC/us12/n621 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n1096 ) );
NAND2_X2 \AES_ENC/us12/U444  ( .A1(\AES_ENC/us12/n1030 ), .A2(\AES_ENC/us12/n1096 ), .ZN(\AES_ENC/us12/n651 ) );
NAND2_X2 \AES_ENC/us12/U443  ( .A1(\AES_ENC/us12/n1114 ), .A2(\AES_ENC/us12/n651 ), .ZN(\AES_ENC/us12/n655 ) );
OR3_X2 \AES_ENC/us12/U440  ( .A1(\AES_ENC/us12/n1079 ), .A2(\AES_ENC/sa12 [7]), .A3(\AES_ENC/us12/n626 ), .ZN(\AES_ENC/us12/n654 ));
NAND2_X2 \AES_ENC/us12/U439  ( .A1(\AES_ENC/us12/n593 ), .A2(\AES_ENC/us12/n601 ), .ZN(\AES_ENC/us12/n652 ) );
NAND4_X2 \AES_ENC/us12/U437  ( .A1(\AES_ENC/us12/n656 ), .A2(\AES_ENC/us12/n655 ), .A3(\AES_ENC/us12/n654 ), .A4(\AES_ENC/us12/n653 ), .ZN(\AES_ENC/us12/n657 ) );
NAND2_X2 \AES_ENC/us12/U436  ( .A1(\AES_ENC/sa12 [2]), .A2(\AES_ENC/us12/n657 ), .ZN(\AES_ENC/us12/n660 ) );
NAND4_X2 \AES_ENC/us12/U432  ( .A1(\AES_ENC/us12/n662 ), .A2(\AES_ENC/us12/n661 ), .A3(\AES_ENC/us12/n660 ), .A4(\AES_ENC/us12/n659 ), .ZN(\AES_ENC/us12/n663 ) );
NAND2_X2 \AES_ENC/us12/U431  ( .A1(\AES_ENC/us12/n663 ), .A2(\AES_ENC/us12/n574 ), .ZN(\AES_ENC/us12/n664 ) );
NAND2_X2 \AES_ENC/us12/U430  ( .A1(\AES_ENC/us12/n665 ), .A2(\AES_ENC/us12/n664 ), .ZN(\AES_ENC/us12/n666 ) );
NAND2_X2 \AES_ENC/us12/U429  ( .A1(\AES_ENC/sa12 [6]), .A2(\AES_ENC/us12/n666 ), .ZN(\AES_ENC/us12/n678 ) );
NAND2_X2 \AES_ENC/us12/U426  ( .A1(\AES_ENC/us12/n735 ), .A2(\AES_ENC/us12/n1093 ), .ZN(\AES_ENC/us12/n675 ) );
NAND2_X2 \AES_ENC/us12/U425  ( .A1(\AES_ENC/us12/n588 ), .A2(\AES_ENC/us12/n597 ), .ZN(\AES_ENC/us12/n1045 ) );
OR2_X2 \AES_ENC/us12/U424  ( .A1(\AES_ENC/us12/n1045 ), .A2(\AES_ENC/us12/n605 ), .ZN(\AES_ENC/us12/n674 ) );
NAND2_X2 \AES_ENC/us12/U423  ( .A1(\AES_ENC/sa12 [1]), .A2(\AES_ENC/us12/n620 ), .ZN(\AES_ENC/us12/n667 ) );
NAND2_X2 \AES_ENC/us12/U422  ( .A1(\AES_ENC/us12/n619 ), .A2(\AES_ENC/us12/n667 ), .ZN(\AES_ENC/us12/n1071 ) );
NAND4_X2 \AES_ENC/us12/U412  ( .A1(\AES_ENC/us12/n675 ), .A2(\AES_ENC/us12/n674 ), .A3(\AES_ENC/us12/n673 ), .A4(\AES_ENC/us12/n672 ), .ZN(\AES_ENC/us12/n676 ) );
NAND2_X2 \AES_ENC/us12/U411  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n676 ), .ZN(\AES_ENC/us12/n677 ) );
NAND2_X2 \AES_ENC/us12/U408  ( .A1(\AES_ENC/us12/n800 ), .A2(\AES_ENC/us12/n1022 ), .ZN(\AES_ENC/us12/n680 ) );
NAND2_X2 \AES_ENC/us12/U407  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n680 ), .ZN(\AES_ENC/us12/n681 ) );
AND2_X2 \AES_ENC/us12/U402  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n684 ), .ZN(\AES_ENC/us12/n682 ) );
NAND4_X2 \AES_ENC/us12/U395  ( .A1(\AES_ENC/us12/n691 ), .A2(\AES_ENC/us12/n581 ), .A3(\AES_ENC/us12/n690 ), .A4(\AES_ENC/us12/n689 ), .ZN(\AES_ENC/us12/n692 ) );
NAND2_X2 \AES_ENC/us12/U394  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n692 ), .ZN(\AES_ENC/us12/n733 ) );
NAND2_X2 \AES_ENC/us12/U392  ( .A1(\AES_ENC/us12/n977 ), .A2(\AES_ENC/us12/n1050 ), .ZN(\AES_ENC/us12/n702 ) );
NAND2_X2 \AES_ENC/us12/U391  ( .A1(\AES_ENC/us12/n1093 ), .A2(\AES_ENC/us12/n1045 ), .ZN(\AES_ENC/us12/n701 ) );
NAND4_X2 \AES_ENC/us12/U381  ( .A1(\AES_ENC/us12/n702 ), .A2(\AES_ENC/us12/n701 ), .A3(\AES_ENC/us12/n700 ), .A4(\AES_ENC/us12/n699 ), .ZN(\AES_ENC/us12/n703 ) );
NAND2_X2 \AES_ENC/us12/U380  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n703 ), .ZN(\AES_ENC/us12/n732 ) );
AND2_X2 \AES_ENC/us12/U379  ( .A1(\AES_ENC/sa12 [0]), .A2(\AES_ENC/sa12 [6]),.ZN(\AES_ENC/us12/n1113 ) );
NAND2_X2 \AES_ENC/us12/U378  ( .A1(\AES_ENC/us12/n601 ), .A2(\AES_ENC/us12/n1030 ), .ZN(\AES_ENC/us12/n881 ) );
NAND2_X2 \AES_ENC/us12/U377  ( .A1(\AES_ENC/us12/n1093 ), .A2(\AES_ENC/us12/n881 ), .ZN(\AES_ENC/us12/n715 ) );
NAND2_X2 \AES_ENC/us12/U376  ( .A1(\AES_ENC/us12/n1010 ), .A2(\AES_ENC/us12/n600 ), .ZN(\AES_ENC/us12/n714 ) );
NAND2_X2 \AES_ENC/us12/U375  ( .A1(\AES_ENC/us12/n855 ), .A2(\AES_ENC/us12/n588 ), .ZN(\AES_ENC/us12/n1117 ) );
XNOR2_X2 \AES_ENC/us12/U371  ( .A(\AES_ENC/us12/n611 ), .B(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n824 ) );
NAND4_X2 \AES_ENC/us12/U362  ( .A1(\AES_ENC/us12/n715 ), .A2(\AES_ENC/us12/n714 ), .A3(\AES_ENC/us12/n713 ), .A4(\AES_ENC/us12/n712 ), .ZN(\AES_ENC/us12/n716 ) );
NAND2_X2 \AES_ENC/us12/U361  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n716 ), .ZN(\AES_ENC/us12/n731 ) );
AND2_X2 \AES_ENC/us12/U360  ( .A1(\AES_ENC/sa12 [6]), .A2(\AES_ENC/us12/n574 ), .ZN(\AES_ENC/us12/n1131 ) );
NAND2_X2 \AES_ENC/us12/U359  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n717 ) );
NAND2_X2 \AES_ENC/us12/U358  ( .A1(\AES_ENC/us12/n1029 ), .A2(\AES_ENC/us12/n717 ), .ZN(\AES_ENC/us12/n728 ) );
NAND2_X2 \AES_ENC/us12/U357  ( .A1(\AES_ENC/sa12 [1]), .A2(\AES_ENC/us12/n624 ), .ZN(\AES_ENC/us12/n1097 ) );
NAND2_X2 \AES_ENC/us12/U356  ( .A1(\AES_ENC/us12/n603 ), .A2(\AES_ENC/us12/n1097 ), .ZN(\AES_ENC/us12/n718 ) );
NAND2_X2 \AES_ENC/us12/U355  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n718 ), .ZN(\AES_ENC/us12/n727 ) );
NAND4_X2 \AES_ENC/us12/U344  ( .A1(\AES_ENC/us12/n728 ), .A2(\AES_ENC/us12/n727 ), .A3(\AES_ENC/us12/n726 ), .A4(\AES_ENC/us12/n725 ), .ZN(\AES_ENC/us12/n729 ) );
NAND2_X2 \AES_ENC/us12/U343  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n729 ), .ZN(\AES_ENC/us12/n730 ) );
NAND4_X2 \AES_ENC/us12/U342  ( .A1(\AES_ENC/us12/n733 ), .A2(\AES_ENC/us12/n732 ), .A3(\AES_ENC/us12/n731 ), .A4(\AES_ENC/us12/n730 ), .ZN(\AES_ENC/sa12_sub[1] ) );
NAND2_X2 \AES_ENC/us12/U341  ( .A1(\AES_ENC/sa12 [7]), .A2(\AES_ENC/us12/n611 ), .ZN(\AES_ENC/us12/n734 ) );
NAND2_X2 \AES_ENC/us12/U340  ( .A1(\AES_ENC/us12/n734 ), .A2(\AES_ENC/us12/n607 ), .ZN(\AES_ENC/us12/n738 ) );
OR4_X2 \AES_ENC/us12/U339  ( .A1(\AES_ENC/us12/n738 ), .A2(\AES_ENC/us12/n626 ), .A3(\AES_ENC/us12/n826 ), .A4(\AES_ENC/us12/n1121 ), .ZN(\AES_ENC/us12/n746 ) );
NAND2_X2 \AES_ENC/us12/U337  ( .A1(\AES_ENC/us12/n1100 ), .A2(\AES_ENC/us12/n587 ), .ZN(\AES_ENC/us12/n992 ) );
OR2_X2 \AES_ENC/us12/U336  ( .A1(\AES_ENC/us12/n610 ), .A2(\AES_ENC/us12/n735 ), .ZN(\AES_ENC/us12/n737 ) );
NAND2_X2 \AES_ENC/us12/U334  ( .A1(\AES_ENC/us12/n619 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n753 ) );
NAND2_X2 \AES_ENC/us12/U333  ( .A1(\AES_ENC/us12/n582 ), .A2(\AES_ENC/us12/n753 ), .ZN(\AES_ENC/us12/n1080 ) );
NAND2_X2 \AES_ENC/us12/U332  ( .A1(\AES_ENC/us12/n1048 ), .A2(\AES_ENC/us12/n576 ), .ZN(\AES_ENC/us12/n736 ) );
NAND2_X2 \AES_ENC/us12/U331  ( .A1(\AES_ENC/us12/n737 ), .A2(\AES_ENC/us12/n736 ), .ZN(\AES_ENC/us12/n739 ) );
NAND2_X2 \AES_ENC/us12/U330  ( .A1(\AES_ENC/us12/n739 ), .A2(\AES_ENC/us12/n738 ), .ZN(\AES_ENC/us12/n745 ) );
NAND2_X2 \AES_ENC/us12/U326  ( .A1(\AES_ENC/us12/n1096 ), .A2(\AES_ENC/us12/n590 ), .ZN(\AES_ENC/us12/n906 ) );
NAND4_X2 \AES_ENC/us12/U323  ( .A1(\AES_ENC/us12/n746 ), .A2(\AES_ENC/us12/n992 ), .A3(\AES_ENC/us12/n745 ), .A4(\AES_ENC/us12/n744 ), .ZN(\AES_ENC/us12/n747 ) );
NAND2_X2 \AES_ENC/us12/U322  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n747 ), .ZN(\AES_ENC/us12/n793 ) );
NAND2_X2 \AES_ENC/us12/U321  ( .A1(\AES_ENC/us12/n584 ), .A2(\AES_ENC/us12/n855 ), .ZN(\AES_ENC/us12/n748 ) );
NAND2_X2 \AES_ENC/us12/U320  ( .A1(\AES_ENC/us12/n956 ), .A2(\AES_ENC/us12/n748 ), .ZN(\AES_ENC/us12/n760 ) );
NAND2_X2 \AES_ENC/us12/U313  ( .A1(\AES_ENC/us12/n590 ), .A2(\AES_ENC/us12/n753 ), .ZN(\AES_ENC/us12/n1023 ) );
NAND4_X2 \AES_ENC/us12/U308  ( .A1(\AES_ENC/us12/n760 ), .A2(\AES_ENC/us12/n992 ), .A3(\AES_ENC/us12/n759 ), .A4(\AES_ENC/us12/n758 ), .ZN(\AES_ENC/us12/n761 ) );
NAND2_X2 \AES_ENC/us12/U307  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n761 ), .ZN(\AES_ENC/us12/n792 ) );
NAND2_X2 \AES_ENC/us12/U306  ( .A1(\AES_ENC/us12/n584 ), .A2(\AES_ENC/us12/n603 ), .ZN(\AES_ENC/us12/n989 ) );
NAND2_X2 \AES_ENC/us12/U305  ( .A1(\AES_ENC/us12/n1050 ), .A2(\AES_ENC/us12/n989 ), .ZN(\AES_ENC/us12/n777 ) );
NAND2_X2 \AES_ENC/us12/U304  ( .A1(\AES_ENC/us12/n1093 ), .A2(\AES_ENC/us12/n762 ), .ZN(\AES_ENC/us12/n776 ) );
XNOR2_X2 \AES_ENC/us12/U301  ( .A(\AES_ENC/sa12 [7]), .B(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n959 ) );
NAND4_X2 \AES_ENC/us12/U289  ( .A1(\AES_ENC/us12/n777 ), .A2(\AES_ENC/us12/n776 ), .A3(\AES_ENC/us12/n775 ), .A4(\AES_ENC/us12/n774 ), .ZN(\AES_ENC/us12/n778 ) );
NAND2_X2 \AES_ENC/us12/U288  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n778 ), .ZN(\AES_ENC/us12/n791 ) );
NAND2_X2 \AES_ENC/us12/U287  ( .A1(\AES_ENC/us12/n1056 ), .A2(\AES_ENC/us12/n1050 ), .ZN(\AES_ENC/us12/n788 ) );
NAND2_X2 \AES_ENC/us12/U286  ( .A1(\AES_ENC/us12/n1091 ), .A2(\AES_ENC/us12/n779 ), .ZN(\AES_ENC/us12/n787 ) );
NAND2_X2 \AES_ENC/us12/U285  ( .A1(\AES_ENC/us12/n956 ), .A2(\AES_ENC/sa12 [1]), .ZN(\AES_ENC/us12/n786 ) );
NAND4_X2 \AES_ENC/us12/U278  ( .A1(\AES_ENC/us12/n788 ), .A2(\AES_ENC/us12/n787 ), .A3(\AES_ENC/us12/n786 ), .A4(\AES_ENC/us12/n785 ), .ZN(\AES_ENC/us12/n789 ) );
NAND2_X2 \AES_ENC/us12/U277  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n789 ), .ZN(\AES_ENC/us12/n790 ) );
NAND4_X2 \AES_ENC/us12/U276  ( .A1(\AES_ENC/us12/n793 ), .A2(\AES_ENC/us12/n792 ), .A3(\AES_ENC/us12/n791 ), .A4(\AES_ENC/us12/n790 ), .ZN(\AES_ENC/sa12_sub[2] ) );
NAND2_X2 \AES_ENC/us12/U275  ( .A1(\AES_ENC/us12/n1059 ), .A2(\AES_ENC/us12/n794 ), .ZN(\AES_ENC/us12/n810 ) );
NAND2_X2 \AES_ENC/us12/U274  ( .A1(\AES_ENC/us12/n1049 ), .A2(\AES_ENC/us12/n956 ), .ZN(\AES_ENC/us12/n809 ) );
OR2_X2 \AES_ENC/us12/U266  ( .A1(\AES_ENC/us12/n1096 ), .A2(\AES_ENC/us12/n606 ), .ZN(\AES_ENC/us12/n802 ) );
NAND2_X2 \AES_ENC/us12/U265  ( .A1(\AES_ENC/us12/n1053 ), .A2(\AES_ENC/us12/n800 ), .ZN(\AES_ENC/us12/n801 ) );
NAND2_X2 \AES_ENC/us12/U264  ( .A1(\AES_ENC/us12/n802 ), .A2(\AES_ENC/us12/n801 ), .ZN(\AES_ENC/us12/n805 ) );
NAND4_X2 \AES_ENC/us12/U261  ( .A1(\AES_ENC/us12/n810 ), .A2(\AES_ENC/us12/n809 ), .A3(\AES_ENC/us12/n808 ), .A4(\AES_ENC/us12/n807 ), .ZN(\AES_ENC/us12/n811 ) );
NAND2_X2 \AES_ENC/us12/U260  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n811 ), .ZN(\AES_ENC/us12/n852 ) );
OR2_X2 \AES_ENC/us12/U259  ( .A1(\AES_ENC/us12/n1023 ), .A2(\AES_ENC/us12/n617 ), .ZN(\AES_ENC/us12/n819 ) );
OR2_X2 \AES_ENC/us12/U257  ( .A1(\AES_ENC/us12/n570 ), .A2(\AES_ENC/us12/n930 ), .ZN(\AES_ENC/us12/n818 ) );
NAND2_X2 \AES_ENC/us12/U256  ( .A1(\AES_ENC/us12/n1013 ), .A2(\AES_ENC/us12/n1094 ), .ZN(\AES_ENC/us12/n817 ) );
NAND4_X2 \AES_ENC/us12/U249  ( .A1(\AES_ENC/us12/n819 ), .A2(\AES_ENC/us12/n818 ), .A3(\AES_ENC/us12/n817 ), .A4(\AES_ENC/us12/n816 ), .ZN(\AES_ENC/us12/n820 ) );
NAND2_X2 \AES_ENC/us12/U248  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n820 ), .ZN(\AES_ENC/us12/n851 ) );
NAND2_X2 \AES_ENC/us12/U247  ( .A1(\AES_ENC/us12/n956 ), .A2(\AES_ENC/us12/n1080 ), .ZN(\AES_ENC/us12/n835 ) );
NAND2_X2 \AES_ENC/us12/U246  ( .A1(\AES_ENC/us12/n570 ), .A2(\AES_ENC/us12/n1030 ), .ZN(\AES_ENC/us12/n1047 ) );
OR2_X2 \AES_ENC/us12/U245  ( .A1(\AES_ENC/us12/n1047 ), .A2(\AES_ENC/us12/n612 ), .ZN(\AES_ENC/us12/n834 ) );
NAND2_X2 \AES_ENC/us12/U244  ( .A1(\AES_ENC/us12/n1072 ), .A2(\AES_ENC/us12/n589 ), .ZN(\AES_ENC/us12/n833 ) );
NAND4_X2 \AES_ENC/us12/U233  ( .A1(\AES_ENC/us12/n835 ), .A2(\AES_ENC/us12/n834 ), .A3(\AES_ENC/us12/n833 ), .A4(\AES_ENC/us12/n832 ), .ZN(\AES_ENC/us12/n836 ) );
NAND2_X2 \AES_ENC/us12/U232  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n836 ), .ZN(\AES_ENC/us12/n850 ) );
NAND2_X2 \AES_ENC/us12/U231  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n623 ), .ZN(\AES_ENC/us12/n847 ) );
NAND2_X2 \AES_ENC/us12/U230  ( .A1(\AES_ENC/us12/n1050 ), .A2(\AES_ENC/us12/n1071 ), .ZN(\AES_ENC/us12/n846 ) );
OR2_X2 \AES_ENC/us12/U224  ( .A1(\AES_ENC/us12/n1053 ), .A2(\AES_ENC/us12/n911 ), .ZN(\AES_ENC/us12/n1077 ) );
NAND4_X2 \AES_ENC/us12/U220  ( .A1(\AES_ENC/us12/n847 ), .A2(\AES_ENC/us12/n846 ), .A3(\AES_ENC/us12/n845 ), .A4(\AES_ENC/us12/n844 ), .ZN(\AES_ENC/us12/n848 ) );
NAND2_X2 \AES_ENC/us12/U219  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n848 ), .ZN(\AES_ENC/us12/n849 ) );
NAND4_X2 \AES_ENC/us12/U218  ( .A1(\AES_ENC/us12/n852 ), .A2(\AES_ENC/us12/n851 ), .A3(\AES_ENC/us12/n850 ), .A4(\AES_ENC/us12/n849 ), .ZN(\AES_ENC/sa12_sub[3] ) );
NAND2_X2 \AES_ENC/us12/U216  ( .A1(\AES_ENC/us12/n1009 ), .A2(\AES_ENC/us12/n1072 ), .ZN(\AES_ENC/us12/n862 ) );
NAND2_X2 \AES_ENC/us12/U215  ( .A1(\AES_ENC/us12/n603 ), .A2(\AES_ENC/us12/n577 ), .ZN(\AES_ENC/us12/n853 ) );
NAND2_X2 \AES_ENC/us12/U214  ( .A1(\AES_ENC/us12/n1050 ), .A2(\AES_ENC/us12/n853 ), .ZN(\AES_ENC/us12/n861 ) );
NAND4_X2 \AES_ENC/us12/U206  ( .A1(\AES_ENC/us12/n862 ), .A2(\AES_ENC/us12/n861 ), .A3(\AES_ENC/us12/n860 ), .A4(\AES_ENC/us12/n859 ), .ZN(\AES_ENC/us12/n863 ) );
NAND2_X2 \AES_ENC/us12/U205  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n863 ), .ZN(\AES_ENC/us12/n905 ) );
NAND2_X2 \AES_ENC/us12/U204  ( .A1(\AES_ENC/us12/n1010 ), .A2(\AES_ENC/us12/n989 ), .ZN(\AES_ENC/us12/n874 ) );
NAND2_X2 \AES_ENC/us12/U203  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n610 ), .ZN(\AES_ENC/us12/n864 ) );
NAND2_X2 \AES_ENC/us12/U202  ( .A1(\AES_ENC/us12/n929 ), .A2(\AES_ENC/us12/n864 ), .ZN(\AES_ENC/us12/n873 ) );
NAND4_X2 \AES_ENC/us12/U193  ( .A1(\AES_ENC/us12/n874 ), .A2(\AES_ENC/us12/n873 ), .A3(\AES_ENC/us12/n872 ), .A4(\AES_ENC/us12/n871 ), .ZN(\AES_ENC/us12/n875 ) );
NAND2_X2 \AES_ENC/us12/U192  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n875 ), .ZN(\AES_ENC/us12/n904 ) );
NAND2_X2 \AES_ENC/us12/U191  ( .A1(\AES_ENC/us12/n583 ), .A2(\AES_ENC/us12/n1050 ), .ZN(\AES_ENC/us12/n889 ) );
NAND2_X2 \AES_ENC/us12/U190  ( .A1(\AES_ENC/us12/n1093 ), .A2(\AES_ENC/us12/n587 ), .ZN(\AES_ENC/us12/n876 ) );
NAND2_X2 \AES_ENC/us12/U189  ( .A1(\AES_ENC/us12/n604 ), .A2(\AES_ENC/us12/n876 ), .ZN(\AES_ENC/us12/n877 ) );
NAND2_X2 \AES_ENC/us12/U188  ( .A1(\AES_ENC/us12/n877 ), .A2(\AES_ENC/us12/n623 ), .ZN(\AES_ENC/us12/n888 ) );
NAND4_X2 \AES_ENC/us12/U179  ( .A1(\AES_ENC/us12/n889 ), .A2(\AES_ENC/us12/n888 ), .A3(\AES_ENC/us12/n887 ), .A4(\AES_ENC/us12/n886 ), .ZN(\AES_ENC/us12/n890 ) );
NAND2_X2 \AES_ENC/us12/U178  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n890 ), .ZN(\AES_ENC/us12/n903 ) );
OR2_X2 \AES_ENC/us12/U177  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n1059 ), .ZN(\AES_ENC/us12/n900 ) );
NAND2_X2 \AES_ENC/us12/U176  ( .A1(\AES_ENC/us12/n1073 ), .A2(\AES_ENC/us12/n1047 ), .ZN(\AES_ENC/us12/n899 ) );
NAND2_X2 \AES_ENC/us12/U175  ( .A1(\AES_ENC/us12/n1094 ), .A2(\AES_ENC/us12/n595 ), .ZN(\AES_ENC/us12/n898 ) );
NAND4_X2 \AES_ENC/us12/U167  ( .A1(\AES_ENC/us12/n900 ), .A2(\AES_ENC/us12/n899 ), .A3(\AES_ENC/us12/n898 ), .A4(\AES_ENC/us12/n897 ), .ZN(\AES_ENC/us12/n901 ) );
NAND2_X2 \AES_ENC/us12/U166  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n901 ), .ZN(\AES_ENC/us12/n902 ) );
NAND4_X2 \AES_ENC/us12/U165  ( .A1(\AES_ENC/us12/n905 ), .A2(\AES_ENC/us12/n904 ), .A3(\AES_ENC/us12/n903 ), .A4(\AES_ENC/us12/n902 ), .ZN(\AES_ENC/sa12_sub[4] ) );
NAND2_X2 \AES_ENC/us12/U164  ( .A1(\AES_ENC/us12/n1094 ), .A2(\AES_ENC/us12/n599 ), .ZN(\AES_ENC/us12/n922 ) );
NAND2_X2 \AES_ENC/us12/U163  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n989 ), .ZN(\AES_ENC/us12/n921 ) );
NAND4_X2 \AES_ENC/us12/U151  ( .A1(\AES_ENC/us12/n922 ), .A2(\AES_ENC/us12/n921 ), .A3(\AES_ENC/us12/n920 ), .A4(\AES_ENC/us12/n919 ), .ZN(\AES_ENC/us12/n923 ) );
NAND2_X2 \AES_ENC/us12/U150  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n923 ), .ZN(\AES_ENC/us12/n972 ) );
NAND2_X2 \AES_ENC/us12/U149  ( .A1(\AES_ENC/us12/n582 ), .A2(\AES_ENC/us12/n619 ), .ZN(\AES_ENC/us12/n924 ) );
NAND2_X2 \AES_ENC/us12/U148  ( .A1(\AES_ENC/us12/n1073 ), .A2(\AES_ENC/us12/n924 ), .ZN(\AES_ENC/us12/n939 ) );
NAND2_X2 \AES_ENC/us12/U147  ( .A1(\AES_ENC/us12/n926 ), .A2(\AES_ENC/us12/n925 ), .ZN(\AES_ENC/us12/n927 ) );
NAND2_X2 \AES_ENC/us12/U146  ( .A1(\AES_ENC/us12/n606 ), .A2(\AES_ENC/us12/n927 ), .ZN(\AES_ENC/us12/n928 ) );
NAND2_X2 \AES_ENC/us12/U145  ( .A1(\AES_ENC/us12/n928 ), .A2(\AES_ENC/us12/n1080 ), .ZN(\AES_ENC/us12/n938 ) );
OR2_X2 \AES_ENC/us12/U144  ( .A1(\AES_ENC/us12/n1117 ), .A2(\AES_ENC/us12/n615 ), .ZN(\AES_ENC/us12/n937 ) );
NAND4_X2 \AES_ENC/us12/U139  ( .A1(\AES_ENC/us12/n939 ), .A2(\AES_ENC/us12/n938 ), .A3(\AES_ENC/us12/n937 ), .A4(\AES_ENC/us12/n936 ), .ZN(\AES_ENC/us12/n940 ) );
NAND2_X2 \AES_ENC/us12/U138  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n940 ), .ZN(\AES_ENC/us12/n971 ) );
OR2_X2 \AES_ENC/us12/U137  ( .A1(\AES_ENC/us12/n605 ), .A2(\AES_ENC/us12/n941 ), .ZN(\AES_ENC/us12/n954 ) );
NAND2_X2 \AES_ENC/us12/U136  ( .A1(\AES_ENC/us12/n1096 ), .A2(\AES_ENC/us12/n577 ), .ZN(\AES_ENC/us12/n942 ) );
NAND2_X2 \AES_ENC/us12/U135  ( .A1(\AES_ENC/us12/n1048 ), .A2(\AES_ENC/us12/n942 ), .ZN(\AES_ENC/us12/n943 ) );
NAND2_X2 \AES_ENC/us12/U134  ( .A1(\AES_ENC/us12/n612 ), .A2(\AES_ENC/us12/n943 ), .ZN(\AES_ENC/us12/n944 ) );
NAND2_X2 \AES_ENC/us12/U133  ( .A1(\AES_ENC/us12/n944 ), .A2(\AES_ENC/us12/n580 ), .ZN(\AES_ENC/us12/n953 ) );
NAND4_X2 \AES_ENC/us12/U125  ( .A1(\AES_ENC/us12/n954 ), .A2(\AES_ENC/us12/n953 ), .A3(\AES_ENC/us12/n952 ), .A4(\AES_ENC/us12/n951 ), .ZN(\AES_ENC/us12/n955 ) );
NAND2_X2 \AES_ENC/us12/U124  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n955 ), .ZN(\AES_ENC/us12/n970 ) );
NAND2_X2 \AES_ENC/us12/U123  ( .A1(\AES_ENC/us12/n1094 ), .A2(\AES_ENC/us12/n1071 ), .ZN(\AES_ENC/us12/n967 ) );
NAND2_X2 \AES_ENC/us12/U122  ( .A1(\AES_ENC/us12/n956 ), .A2(\AES_ENC/us12/n1030 ), .ZN(\AES_ENC/us12/n966 ) );
NAND4_X2 \AES_ENC/us12/U114  ( .A1(\AES_ENC/us12/n967 ), .A2(\AES_ENC/us12/n966 ), .A3(\AES_ENC/us12/n965 ), .A4(\AES_ENC/us12/n964 ), .ZN(\AES_ENC/us12/n968 ) );
NAND2_X2 \AES_ENC/us12/U113  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n968 ), .ZN(\AES_ENC/us12/n969 ) );
NAND4_X2 \AES_ENC/us12/U112  ( .A1(\AES_ENC/us12/n972 ), .A2(\AES_ENC/us12/n971 ), .A3(\AES_ENC/us12/n970 ), .A4(\AES_ENC/us12/n969 ), .ZN(\AES_ENC/sa12_sub[5] ) );
NAND2_X2 \AES_ENC/us12/U111  ( .A1(\AES_ENC/us12/n570 ), .A2(\AES_ENC/us12/n1097 ), .ZN(\AES_ENC/us12/n973 ) );
NAND2_X2 \AES_ENC/us12/U110  ( .A1(\AES_ENC/us12/n1073 ), .A2(\AES_ENC/us12/n973 ), .ZN(\AES_ENC/us12/n987 ) );
NAND2_X2 \AES_ENC/us12/U109  ( .A1(\AES_ENC/us12/n974 ), .A2(\AES_ENC/us12/n1077 ), .ZN(\AES_ENC/us12/n975 ) );
NAND2_X2 \AES_ENC/us12/U108  ( .A1(\AES_ENC/us12/n613 ), .A2(\AES_ENC/us12/n975 ), .ZN(\AES_ENC/us12/n976 ) );
NAND2_X2 \AES_ENC/us12/U107  ( .A1(\AES_ENC/us12/n977 ), .A2(\AES_ENC/us12/n976 ), .ZN(\AES_ENC/us12/n986 ) );
NAND4_X2 \AES_ENC/us12/U99  ( .A1(\AES_ENC/us12/n987 ), .A2(\AES_ENC/us12/n986 ), .A3(\AES_ENC/us12/n985 ), .A4(\AES_ENC/us12/n984 ), .ZN(\AES_ENC/us12/n988 ) );
NAND2_X2 \AES_ENC/us12/U98  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n988 ), .ZN(\AES_ENC/us12/n1044 ) );
NAND2_X2 \AES_ENC/us12/U97  ( .A1(\AES_ENC/us12/n1073 ), .A2(\AES_ENC/us12/n989 ), .ZN(\AES_ENC/us12/n1004 ) );
NAND2_X2 \AES_ENC/us12/U96  ( .A1(\AES_ENC/us12/n1092 ), .A2(\AES_ENC/us12/n619 ), .ZN(\AES_ENC/us12/n1003 ) );
NAND4_X2 \AES_ENC/us12/U85  ( .A1(\AES_ENC/us12/n1004 ), .A2(\AES_ENC/us12/n1003 ), .A3(\AES_ENC/us12/n1002 ), .A4(\AES_ENC/us12/n1001 ), .ZN(\AES_ENC/us12/n1005 ) );
NAND2_X2 \AES_ENC/us12/U84  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n1005 ), .ZN(\AES_ENC/us12/n1043 ) );
NAND2_X2 \AES_ENC/us12/U83  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n596 ), .ZN(\AES_ENC/us12/n1020 ) );
NAND2_X2 \AES_ENC/us12/U82  ( .A1(\AES_ENC/us12/n1050 ), .A2(\AES_ENC/us12/n624 ), .ZN(\AES_ENC/us12/n1019 ) );
NAND2_X2 \AES_ENC/us12/U77  ( .A1(\AES_ENC/us12/n1059 ), .A2(\AES_ENC/us12/n1114 ), .ZN(\AES_ENC/us12/n1012 ) );
NAND2_X2 \AES_ENC/us12/U76  ( .A1(\AES_ENC/us12/n1010 ), .A2(\AES_ENC/us12/n592 ), .ZN(\AES_ENC/us12/n1011 ) );
NAND2_X2 \AES_ENC/us12/U75  ( .A1(\AES_ENC/us12/n1012 ), .A2(\AES_ENC/us12/n1011 ), .ZN(\AES_ENC/us12/n1016 ) );
NAND4_X2 \AES_ENC/us12/U70  ( .A1(\AES_ENC/us12/n1020 ), .A2(\AES_ENC/us12/n1019 ), .A3(\AES_ENC/us12/n1018 ), .A4(\AES_ENC/us12/n1017 ), .ZN(\AES_ENC/us12/n1021 ) );
NAND2_X2 \AES_ENC/us12/U69  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n1021 ), .ZN(\AES_ENC/us12/n1042 ) );
NAND2_X2 \AES_ENC/us12/U68  ( .A1(\AES_ENC/us12/n1022 ), .A2(\AES_ENC/us12/n1093 ), .ZN(\AES_ENC/us12/n1039 ) );
NAND2_X2 \AES_ENC/us12/U67  ( .A1(\AES_ENC/us12/n1050 ), .A2(\AES_ENC/us12/n1023 ), .ZN(\AES_ENC/us12/n1038 ) );
NAND2_X2 \AES_ENC/us12/U66  ( .A1(\AES_ENC/us12/n1024 ), .A2(\AES_ENC/us12/n1071 ), .ZN(\AES_ENC/us12/n1037 ) );
AND2_X2 \AES_ENC/us12/U60  ( .A1(\AES_ENC/us12/n1030 ), .A2(\AES_ENC/us12/n602 ), .ZN(\AES_ENC/us12/n1078 ) );
NAND4_X2 \AES_ENC/us12/U56  ( .A1(\AES_ENC/us12/n1039 ), .A2(\AES_ENC/us12/n1038 ), .A3(\AES_ENC/us12/n1037 ), .A4(\AES_ENC/us12/n1036 ), .ZN(\AES_ENC/us12/n1040 ) );
NAND2_X2 \AES_ENC/us12/U55  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n1040 ), .ZN(\AES_ENC/us12/n1041 ) );
NAND4_X2 \AES_ENC/us12/U54  ( .A1(\AES_ENC/us12/n1044 ), .A2(\AES_ENC/us12/n1043 ), .A3(\AES_ENC/us12/n1042 ), .A4(\AES_ENC/us12/n1041 ), .ZN(\AES_ENC/sa12_sub[6] ) );
NAND2_X2 \AES_ENC/us12/U53  ( .A1(\AES_ENC/us12/n1072 ), .A2(\AES_ENC/us12/n1045 ), .ZN(\AES_ENC/us12/n1068 ) );
NAND2_X2 \AES_ENC/us12/U52  ( .A1(\AES_ENC/us12/n1046 ), .A2(\AES_ENC/us12/n582 ), .ZN(\AES_ENC/us12/n1067 ) );
NAND2_X2 \AES_ENC/us12/U51  ( .A1(\AES_ENC/us12/n1094 ), .A2(\AES_ENC/us12/n1047 ), .ZN(\AES_ENC/us12/n1066 ) );
NAND4_X2 \AES_ENC/us12/U40  ( .A1(\AES_ENC/us12/n1068 ), .A2(\AES_ENC/us12/n1067 ), .A3(\AES_ENC/us12/n1066 ), .A4(\AES_ENC/us12/n1065 ), .ZN(\AES_ENC/us12/n1069 ) );
NAND2_X2 \AES_ENC/us12/U39  ( .A1(\AES_ENC/us12/n1070 ), .A2(\AES_ENC/us12/n1069 ), .ZN(\AES_ENC/us12/n1135 ) );
NAND2_X2 \AES_ENC/us12/U38  ( .A1(\AES_ENC/us12/n1072 ), .A2(\AES_ENC/us12/n1071 ), .ZN(\AES_ENC/us12/n1088 ) );
NAND2_X2 \AES_ENC/us12/U37  ( .A1(\AES_ENC/us12/n1073 ), .A2(\AES_ENC/us12/n595 ), .ZN(\AES_ENC/us12/n1087 ) );
NAND4_X2 \AES_ENC/us12/U28  ( .A1(\AES_ENC/us12/n1088 ), .A2(\AES_ENC/us12/n1087 ), .A3(\AES_ENC/us12/n1086 ), .A4(\AES_ENC/us12/n1085 ), .ZN(\AES_ENC/us12/n1089 ) );
NAND2_X2 \AES_ENC/us12/U27  ( .A1(\AES_ENC/us12/n1090 ), .A2(\AES_ENC/us12/n1089 ), .ZN(\AES_ENC/us12/n1134 ) );
NAND2_X2 \AES_ENC/us12/U26  ( .A1(\AES_ENC/us12/n1091 ), .A2(\AES_ENC/us12/n1093 ), .ZN(\AES_ENC/us12/n1111 ) );
NAND2_X2 \AES_ENC/us12/U25  ( .A1(\AES_ENC/us12/n1092 ), .A2(\AES_ENC/us12/n1120 ), .ZN(\AES_ENC/us12/n1110 ) );
AND2_X2 \AES_ENC/us12/U22  ( .A1(\AES_ENC/us12/n1097 ), .A2(\AES_ENC/us12/n1096 ), .ZN(\AES_ENC/us12/n1098 ) );
NAND4_X2 \AES_ENC/us12/U14  ( .A1(\AES_ENC/us12/n1111 ), .A2(\AES_ENC/us12/n1110 ), .A3(\AES_ENC/us12/n1109 ), .A4(\AES_ENC/us12/n1108 ), .ZN(\AES_ENC/us12/n1112 ) );
NAND2_X2 \AES_ENC/us12/U13  ( .A1(\AES_ENC/us12/n1113 ), .A2(\AES_ENC/us12/n1112 ), .ZN(\AES_ENC/us12/n1133 ) );
NAND2_X2 \AES_ENC/us12/U12  ( .A1(\AES_ENC/us12/n1115 ), .A2(\AES_ENC/us12/n1114 ), .ZN(\AES_ENC/us12/n1129 ) );
OR2_X2 \AES_ENC/us12/U11  ( .A1(\AES_ENC/us12/n608 ), .A2(\AES_ENC/us12/n1116 ), .ZN(\AES_ENC/us12/n1128 ) );
NAND4_X2 \AES_ENC/us12/U3  ( .A1(\AES_ENC/us12/n1129 ), .A2(\AES_ENC/us12/n1128 ), .A3(\AES_ENC/us12/n1127 ), .A4(\AES_ENC/us12/n1126 ), .ZN(\AES_ENC/us12/n1130 ) );
NAND2_X2 \AES_ENC/us12/U2  ( .A1(\AES_ENC/us12/n1131 ), .A2(\AES_ENC/us12/n1130 ), .ZN(\AES_ENC/us12/n1132 ) );
NAND4_X2 \AES_ENC/us12/U1  ( .A1(\AES_ENC/us12/n1135 ), .A2(\AES_ENC/us12/n1134 ), .A3(\AES_ENC/us12/n1133 ), .A4(\AES_ENC/us12/n1132 ), .ZN(\AES_ENC/sa12_sub[7] ) );
INV_X4 \AES_ENC/us13/U575  ( .A(\AES_ENC/sa13 [0]), .ZN(\AES_ENC/us13/n627 ));
INV_X4 \AES_ENC/us13/U574  ( .A(\AES_ENC/us13/n1053 ), .ZN(\AES_ENC/us13/n625 ) );
INV_X4 \AES_ENC/us13/U573  ( .A(\AES_ENC/us13/n1103 ), .ZN(\AES_ENC/us13/n623 ) );
INV_X4 \AES_ENC/us13/U572  ( .A(\AES_ENC/us13/n1056 ), .ZN(\AES_ENC/us13/n622 ) );
INV_X4 \AES_ENC/us13/U571  ( .A(\AES_ENC/us13/n1102 ), .ZN(\AES_ENC/us13/n621 ) );
INV_X4 \AES_ENC/us13/U570  ( .A(\AES_ENC/us13/n1074 ), .ZN(\AES_ENC/us13/n620 ) );
INV_X4 \AES_ENC/us13/U569  ( .A(\AES_ENC/us13/n929 ), .ZN(\AES_ENC/us13/n619 ) );
INV_X4 \AES_ENC/us13/U568  ( .A(\AES_ENC/us13/n1091 ), .ZN(\AES_ENC/us13/n618 ) );
INV_X4 \AES_ENC/us13/U567  ( .A(\AES_ENC/us13/n826 ), .ZN(\AES_ENC/us13/n617 ) );
INV_X4 \AES_ENC/us13/U566  ( .A(\AES_ENC/us13/n1031 ), .ZN(\AES_ENC/us13/n616 ) );
INV_X4 \AES_ENC/us13/U565  ( .A(\AES_ENC/us13/n1054 ), .ZN(\AES_ENC/us13/n615 ) );
INV_X4 \AES_ENC/us13/U564  ( .A(\AES_ENC/us13/n1025 ), .ZN(\AES_ENC/us13/n614 ) );
INV_X4 \AES_ENC/us13/U563  ( .A(\AES_ENC/us13/n990 ), .ZN(\AES_ENC/us13/n613 ) );
INV_X4 \AES_ENC/us13/U562  ( .A(\AES_ENC/sa13 [4]), .ZN(\AES_ENC/us13/n612 ));
INV_X4 \AES_ENC/us13/U561  ( .A(\AES_ENC/us13/n881 ), .ZN(\AES_ENC/us13/n611 ) );
INV_X4 \AES_ENC/us13/U560  ( .A(\AES_ENC/us13/n1022 ), .ZN(\AES_ENC/us13/n610 ) );
INV_X4 \AES_ENC/us13/U559  ( .A(\AES_ENC/us13/n1120 ), .ZN(\AES_ENC/us13/n609 ) );
INV_X4 \AES_ENC/us13/U558  ( .A(\AES_ENC/us13/n977 ), .ZN(\AES_ENC/us13/n608 ) );
INV_X4 \AES_ENC/us13/U557  ( .A(\AES_ENC/us13/n926 ), .ZN(\AES_ENC/us13/n607 ) );
INV_X4 \AES_ENC/us13/U556  ( .A(\AES_ENC/us13/n910 ), .ZN(\AES_ENC/us13/n606 ) );
INV_X4 \AES_ENC/us13/U555  ( .A(\AES_ENC/us13/n1121 ), .ZN(\AES_ENC/us13/n605 ) );
INV_X4 \AES_ENC/us13/U554  ( .A(\AES_ENC/us13/n1009 ), .ZN(\AES_ENC/us13/n604 ) );
INV_X4 \AES_ENC/us13/U553  ( .A(\AES_ENC/us13/n1080 ), .ZN(\AES_ENC/us13/n602 ) );
INV_X4 \AES_ENC/us13/U552  ( .A(\AES_ENC/us13/n821 ), .ZN(\AES_ENC/us13/n600 ) );
INV_X4 \AES_ENC/us13/U551  ( .A(\AES_ENC/us13/n1013 ), .ZN(\AES_ENC/us13/n599 ) );
INV_X4 \AES_ENC/us13/U550  ( .A(\AES_ENC/us13/n1058 ), .ZN(\AES_ENC/us13/n598 ) );
INV_X4 \AES_ENC/us13/U549  ( .A(\AES_ENC/us13/n906 ), .ZN(\AES_ENC/us13/n597 ) );
INV_X4 \AES_ENC/us13/U548  ( .A(\AES_ENC/us13/n959 ), .ZN(\AES_ENC/us13/n596 ) );
INV_X4 \AES_ENC/us13/U547  ( .A(\AES_ENC/sa13 [7]), .ZN(\AES_ENC/us13/n595 ));
INV_X4 \AES_ENC/us13/U546  ( .A(\AES_ENC/us13/n1114 ), .ZN(\AES_ENC/us13/n593 ) );
INV_X4 \AES_ENC/us13/U545  ( .A(\AES_ENC/us13/n1048 ), .ZN(\AES_ENC/us13/n592 ) );
INV_X4 \AES_ENC/us13/U544  ( .A(\AES_ENC/us13/n974 ), .ZN(\AES_ENC/us13/n590 ) );
INV_X4 \AES_ENC/us13/U543  ( .A(\AES_ENC/us13/n794 ), .ZN(\AES_ENC/us13/n588 ) );
INV_X4 \AES_ENC/us13/U542  ( .A(\AES_ENC/us13/n880 ), .ZN(\AES_ENC/us13/n586 ) );
INV_X4 \AES_ENC/us13/U541  ( .A(\AES_ENC/sa13 [2]), .ZN(\AES_ENC/us13/n584 ));
INV_X4 \AES_ENC/us13/U540  ( .A(\AES_ENC/us13/n800 ), .ZN(\AES_ENC/us13/n583 ) );
INV_X4 \AES_ENC/us13/U539  ( .A(\AES_ENC/us13/n925 ), .ZN(\AES_ENC/us13/n582 ) );
INV_X4 \AES_ENC/us13/U538  ( .A(\AES_ENC/us13/n992 ), .ZN(\AES_ENC/us13/n580 ) );
INV_X4 \AES_ENC/us13/U537  ( .A(\AES_ENC/us13/n779 ), .ZN(\AES_ENC/us13/n579 ) );
INV_X4 \AES_ENC/us13/U536  ( .A(\AES_ENC/us13/n1092 ), .ZN(\AES_ENC/us13/n575 ) );
INV_X4 \AES_ENC/us13/U535  ( .A(\AES_ENC/us13/n824 ), .ZN(\AES_ENC/us13/n574 ) );
NOR2_X2 \AES_ENC/us13/U534  ( .A1(\AES_ENC/sa13 [0]), .A2(\AES_ENC/sa13 [6]),.ZN(\AES_ENC/us13/n1090 ) );
NOR2_X2 \AES_ENC/us13/U533  ( .A1(\AES_ENC/us13/n627 ), .A2(\AES_ENC/sa13 [6]), .ZN(\AES_ENC/us13/n1070 ) );
NOR2_X2 \AES_ENC/us13/U532  ( .A1(\AES_ENC/sa13 [4]), .A2(\AES_ENC/sa13 [3]),.ZN(\AES_ENC/us13/n1025 ) );
INV_X4 \AES_ENC/us13/U531  ( .A(\AES_ENC/us13/n569 ), .ZN(\AES_ENC/us13/n572 ) );
NOR2_X2 \AES_ENC/us13/U530  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n765 ) );
NOR2_X2 \AES_ENC/us13/U529  ( .A1(\AES_ENC/sa13 [4]), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n764 ) );
NOR2_X2 \AES_ENC/us13/U528  ( .A1(\AES_ENC/us13/n765 ), .A2(\AES_ENC/us13/n764 ), .ZN(\AES_ENC/us13/n766 ) );
NOR2_X2 \AES_ENC/us13/U527  ( .A1(\AES_ENC/us13/n766 ), .A2(\AES_ENC/us13/n596 ), .ZN(\AES_ENC/us13/n767 ) );
NOR3_X2 \AES_ENC/us13/U526  ( .A1(\AES_ENC/us13/n595 ), .A2(\AES_ENC/sa13 [5]), .A3(\AES_ENC/us13/n704 ), .ZN(\AES_ENC/us13/n706 ));
NOR2_X2 \AES_ENC/us13/U525  ( .A1(\AES_ENC/us13/n1117 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n707 ) );
NOR2_X2 \AES_ENC/us13/U524  ( .A1(\AES_ENC/sa13 [4]), .A2(\AES_ENC/us13/n575 ), .ZN(\AES_ENC/us13/n705 ) );
NOR3_X2 \AES_ENC/us13/U523  ( .A1(\AES_ENC/us13/n707 ), .A2(\AES_ENC/us13/n706 ), .A3(\AES_ENC/us13/n705 ), .ZN(\AES_ENC/us13/n713 ) );
INV_X4 \AES_ENC/us13/U522  ( .A(\AES_ENC/sa13 [3]), .ZN(\AES_ENC/us13/n624 ));
NAND3_X2 \AES_ENC/us13/U521  ( .A1(\AES_ENC/us13/n652 ), .A2(\AES_ENC/us13/n594 ), .A3(\AES_ENC/sa13 [7]), .ZN(\AES_ENC/us13/n653 ));
NOR2_X2 \AES_ENC/us13/U520  ( .A1(\AES_ENC/us13/n584 ), .A2(\AES_ENC/sa13 [5]), .ZN(\AES_ENC/us13/n925 ) );
NOR2_X2 \AES_ENC/us13/U519  ( .A1(\AES_ENC/sa13 [5]), .A2(\AES_ENC/sa13 [2]),.ZN(\AES_ENC/us13/n974 ) );
INV_X4 \AES_ENC/us13/U518  ( .A(\AES_ENC/sa13 [5]), .ZN(\AES_ENC/us13/n594 ));
NOR2_X2 \AES_ENC/us13/U517  ( .A1(\AES_ENC/us13/n584 ), .A2(\AES_ENC/sa13 [7]), .ZN(\AES_ENC/us13/n779 ) );
NAND3_X2 \AES_ENC/us13/U516  ( .A1(\AES_ENC/us13/n679 ), .A2(\AES_ENC/us13/n678 ), .A3(\AES_ENC/us13/n677 ), .ZN(\AES_ENC/sa13_sub[0] ) );
NOR2_X2 \AES_ENC/us13/U515  ( .A1(\AES_ENC/us13/n594 ), .A2(\AES_ENC/sa13 [2]), .ZN(\AES_ENC/us13/n1048 ) );
NOR4_X2 \AES_ENC/us13/U512  ( .A1(\AES_ENC/us13/n633 ), .A2(\AES_ENC/us13/n632 ), .A3(\AES_ENC/us13/n631 ), .A4(\AES_ENC/us13/n630 ), .ZN(\AES_ENC/us13/n634 ) );
NOR2_X2 \AES_ENC/us13/U510  ( .A1(\AES_ENC/us13/n629 ), .A2(\AES_ENC/us13/n628 ), .ZN(\AES_ENC/us13/n635 ) );
NAND3_X2 \AES_ENC/us13/U509  ( .A1(\AES_ENC/sa13 [2]), .A2(\AES_ENC/sa13 [7]), .A3(\AES_ENC/us13/n1059 ), .ZN(\AES_ENC/us13/n636 ) );
NOR2_X2 \AES_ENC/us13/U508  ( .A1(\AES_ENC/sa13 [7]), .A2(\AES_ENC/sa13 [2]),.ZN(\AES_ENC/us13/n794 ) );
NOR2_X2 \AES_ENC/us13/U507  ( .A1(\AES_ENC/sa13 [4]), .A2(\AES_ENC/sa13 [1]),.ZN(\AES_ENC/us13/n1102 ) );
NOR2_X2 \AES_ENC/us13/U506  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/sa13 [3]), .ZN(\AES_ENC/us13/n1053 ) );
NOR2_X2 \AES_ENC/us13/U505  ( .A1(\AES_ENC/us13/n579 ), .A2(\AES_ENC/sa13 [5]), .ZN(\AES_ENC/us13/n1024 ) );
NOR2_X2 \AES_ENC/us13/U504  ( .A1(\AES_ENC/us13/n593 ), .A2(\AES_ENC/sa13 [2]), .ZN(\AES_ENC/us13/n1093 ) );
NOR2_X2 \AES_ENC/us13/U503  ( .A1(\AES_ENC/us13/n588 ), .A2(\AES_ENC/sa13 [5]), .ZN(\AES_ENC/us13/n1094 ) );
NOR2_X2 \AES_ENC/us13/U502  ( .A1(\AES_ENC/us13/n612 ), .A2(\AES_ENC/sa13 [3]), .ZN(\AES_ENC/us13/n931 ) );
INV_X4 \AES_ENC/us13/U501  ( .A(\AES_ENC/us13/n570 ), .ZN(\AES_ENC/us13/n573 ) );
NOR2_X2 \AES_ENC/us13/U500  ( .A1(\AES_ENC/us13/n1053 ), .A2(\AES_ENC/us13/n1095 ), .ZN(\AES_ENC/us13/n639 ) );
NOR3_X2 \AES_ENC/us13/U499  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n573 ), .A3(\AES_ENC/us13/n1074 ), .ZN(\AES_ENC/us13/n641 ) );
NOR2_X2 \AES_ENC/us13/U498  ( .A1(\AES_ENC/us13/n639 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n640 ) );
NOR2_X2 \AES_ENC/us13/U497  ( .A1(\AES_ENC/us13/n641 ), .A2(\AES_ENC/us13/n640 ), .ZN(\AES_ENC/us13/n646 ) );
NOR3_X2 \AES_ENC/us13/U496  ( .A1(\AES_ENC/us13/n995 ), .A2(\AES_ENC/us13/n580 ), .A3(\AES_ENC/us13/n994 ), .ZN(\AES_ENC/us13/n1002 ) );
NOR2_X2 \AES_ENC/us13/U495  ( .A1(\AES_ENC/us13/n909 ), .A2(\AES_ENC/us13/n908 ), .ZN(\AES_ENC/us13/n920 ) );
NOR2_X2 \AES_ENC/us13/U494  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n823 ) );
NOR2_X2 \AES_ENC/us13/U492  ( .A1(\AES_ENC/us13/n612 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n822 ) );
NOR2_X2 \AES_ENC/us13/U491  ( .A1(\AES_ENC/us13/n823 ), .A2(\AES_ENC/us13/n822 ), .ZN(\AES_ENC/us13/n825 ) );
NOR2_X2 \AES_ENC/us13/U490  ( .A1(\AES_ENC/sa13 [1]), .A2(\AES_ENC/us13/n601 ), .ZN(\AES_ENC/us13/n913 ) );
NOR2_X2 \AES_ENC/us13/U489  ( .A1(\AES_ENC/us13/n913 ), .A2(\AES_ENC/us13/n1091 ), .ZN(\AES_ENC/us13/n914 ) );
NOR2_X2 \AES_ENC/us13/U488  ( .A1(\AES_ENC/us13/n826 ), .A2(\AES_ENC/us13/n572 ), .ZN(\AES_ENC/us13/n827 ) );
NOR3_X2 \AES_ENC/us13/U487  ( .A1(\AES_ENC/us13/n769 ), .A2(\AES_ENC/us13/n768 ), .A3(\AES_ENC/us13/n767 ), .ZN(\AES_ENC/us13/n775 ) );
NOR2_X2 \AES_ENC/us13/U486  ( .A1(\AES_ENC/us13/n1056 ), .A2(\AES_ENC/us13/n1053 ), .ZN(\AES_ENC/us13/n749 ) );
NOR2_X2 \AES_ENC/us13/U483  ( .A1(\AES_ENC/us13/n749 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n752 ) );
INV_X4 \AES_ENC/us13/U482  ( .A(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n626 ));
NOR2_X2 \AES_ENC/us13/U480  ( .A1(\AES_ENC/us13/n1054 ), .A2(\AES_ENC/us13/n1053 ), .ZN(\AES_ENC/us13/n1055 ) );
OR2_X4 \AES_ENC/us13/U479  ( .A1(\AES_ENC/us13/n1094 ), .A2(\AES_ENC/us13/n1093 ), .ZN(\AES_ENC/us13/n571 ) );
AND2_X2 \AES_ENC/us13/U478  ( .A1(\AES_ENC/us13/n571 ), .A2(\AES_ENC/us13/n1095 ), .ZN(\AES_ENC/us13/n1101 ) );
NOR2_X2 \AES_ENC/us13/U477  ( .A1(\AES_ENC/us13/n1074 ), .A2(\AES_ENC/us13/n931 ), .ZN(\AES_ENC/us13/n796 ) );
NOR2_X2 \AES_ENC/us13/U474  ( .A1(\AES_ENC/us13/n796 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n797 ) );
NOR2_X2 \AES_ENC/us13/U473  ( .A1(\AES_ENC/us13/n932 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n933 ) );
NOR2_X2 \AES_ENC/us13/U472  ( .A1(\AES_ENC/us13/n929 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n935 ) );
NOR2_X2 \AES_ENC/us13/U471  ( .A1(\AES_ENC/us13/n931 ), .A2(\AES_ENC/us13/n930 ), .ZN(\AES_ENC/us13/n934 ) );
NOR3_X2 \AES_ENC/us13/U470  ( .A1(\AES_ENC/us13/n935 ), .A2(\AES_ENC/us13/n934 ), .A3(\AES_ENC/us13/n933 ), .ZN(\AES_ENC/us13/n936 ) );
NOR2_X2 \AES_ENC/us13/U469  ( .A1(\AES_ENC/us13/n612 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n1075 ) );
NOR2_X2 \AES_ENC/us13/U468  ( .A1(\AES_ENC/us13/n572 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n949 ) );
NOR2_X2 \AES_ENC/us13/U467  ( .A1(\AES_ENC/us13/n1049 ), .A2(\AES_ENC/us13/n592 ), .ZN(\AES_ENC/us13/n1051 ) );
NOR2_X2 \AES_ENC/us13/U466  ( .A1(\AES_ENC/us13/n1051 ), .A2(\AES_ENC/us13/n1050 ), .ZN(\AES_ENC/us13/n1052 ) );
NOR2_X2 \AES_ENC/us13/U465  ( .A1(\AES_ENC/us13/n1052 ), .A2(\AES_ENC/us13/n604 ), .ZN(\AES_ENC/us13/n1064 ) );
NOR2_X2 \AES_ENC/us13/U464  ( .A1(\AES_ENC/sa13 [1]), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n631 ) );
NOR2_X2 \AES_ENC/us13/U463  ( .A1(\AES_ENC/us13/n1025 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n980 ) );
NOR2_X2 \AES_ENC/us13/U462  ( .A1(\AES_ENC/us13/n1073 ), .A2(\AES_ENC/us13/n1094 ), .ZN(\AES_ENC/us13/n795 ) );
NOR2_X2 \AES_ENC/us13/U461  ( .A1(\AES_ENC/us13/n795 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n799 ) );
NOR2_X2 \AES_ENC/us13/U460  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n981 ) );
NOR2_X2 \AES_ENC/us13/U459  ( .A1(\AES_ENC/us13/n1102 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n643 ) );
NOR2_X2 \AES_ENC/us13/U458  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n624 ), .ZN(\AES_ENC/us13/n642 ) );
NOR2_X2 \AES_ENC/us13/U455  ( .A1(\AES_ENC/us13/n911 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n644 ) );
NOR4_X2 \AES_ENC/us13/U448  ( .A1(\AES_ENC/us13/n644 ), .A2(\AES_ENC/us13/n643 ), .A3(\AES_ENC/us13/n804 ), .A4(\AES_ENC/us13/n642 ), .ZN(\AES_ENC/us13/n645 ) );
NOR2_X2 \AES_ENC/us13/U447  ( .A1(\AES_ENC/us13/n1102 ), .A2(\AES_ENC/us13/n910 ), .ZN(\AES_ENC/us13/n932 ) );
NOR2_X2 \AES_ENC/us13/U442  ( .A1(\AES_ENC/us13/n1102 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n755 ) );
NOR2_X2 \AES_ENC/us13/U441  ( .A1(\AES_ENC/us13/n931 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n743 ) );
NOR2_X2 \AES_ENC/us13/U438  ( .A1(\AES_ENC/us13/n1072 ), .A2(\AES_ENC/us13/n1094 ), .ZN(\AES_ENC/us13/n930 ) );
NOR2_X2 \AES_ENC/us13/U435  ( .A1(\AES_ENC/us13/n1074 ), .A2(\AES_ENC/us13/n1025 ), .ZN(\AES_ENC/us13/n891 ) );
NOR2_X2 \AES_ENC/us13/U434  ( .A1(\AES_ENC/us13/n891 ), .A2(\AES_ENC/us13/n582 ), .ZN(\AES_ENC/us13/n894 ) );
NOR3_X2 \AES_ENC/us13/U433  ( .A1(\AES_ENC/us13/n601 ), .A2(\AES_ENC/sa13 [1]), .A3(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n683 ));
INV_X4 \AES_ENC/us13/U428  ( .A(\AES_ENC/us13/n931 ), .ZN(\AES_ENC/us13/n601 ) );
NOR2_X2 \AES_ENC/us13/U427  ( .A1(\AES_ENC/us13/n996 ), .A2(\AES_ENC/us13/n931 ), .ZN(\AES_ENC/us13/n704 ) );
NOR2_X2 \AES_ENC/us13/U421  ( .A1(\AES_ENC/us13/n931 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n685 ) );
NOR2_X2 \AES_ENC/us13/U420  ( .A1(\AES_ENC/us13/n1029 ), .A2(\AES_ENC/us13/n1025 ), .ZN(\AES_ENC/us13/n1079 ) );
NOR3_X2 \AES_ENC/us13/U419  ( .A1(\AES_ENC/us13/n620 ), .A2(\AES_ENC/us13/n1025 ), .A3(\AES_ENC/us13/n590 ), .ZN(\AES_ENC/us13/n945 ) );
NOR2_X2 \AES_ENC/us13/U418  ( .A1(\AES_ENC/us13/n594 ), .A2(\AES_ENC/us13/n584 ), .ZN(\AES_ENC/us13/n800 ) );
NOR3_X2 \AES_ENC/us13/U417  ( .A1(\AES_ENC/us13/n598 ), .A2(\AES_ENC/us13/n595 ), .A3(\AES_ENC/us13/n584 ), .ZN(\AES_ENC/us13/n798 ) );
NOR3_X2 \AES_ENC/us13/U416  ( .A1(\AES_ENC/us13/n583 ), .A2(\AES_ENC/us13/n572 ), .A3(\AES_ENC/us13/n596 ), .ZN(\AES_ENC/us13/n962 ) );
NOR3_X2 \AES_ENC/us13/U415  ( .A1(\AES_ENC/us13/n959 ), .A2(\AES_ENC/us13/n572 ), .A3(\AES_ENC/us13/n582 ), .ZN(\AES_ENC/us13/n768 ) );
NOR3_X2 \AES_ENC/us13/U414  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n572 ), .A3(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n694 ) );
NOR3_X2 \AES_ENC/us13/U413  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n572 ), .A3(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n895 ) );
NOR3_X2 \AES_ENC/us13/U410  ( .A1(\AES_ENC/us13/n1008 ), .A2(\AES_ENC/us13/n1007 ), .A3(\AES_ENC/us13/n1006 ), .ZN(\AES_ENC/us13/n1018 ) );
NOR4_X2 \AES_ENC/us13/U409  ( .A1(\AES_ENC/us13/n806 ), .A2(\AES_ENC/us13/n805 ), .A3(\AES_ENC/us13/n804 ), .A4(\AES_ENC/us13/n803 ), .ZN(\AES_ENC/us13/n807 ) );
NOR3_X2 \AES_ENC/us13/U406  ( .A1(\AES_ENC/us13/n799 ), .A2(\AES_ENC/us13/n798 ), .A3(\AES_ENC/us13/n797 ), .ZN(\AES_ENC/us13/n808 ) );
NOR4_X2 \AES_ENC/us13/U405  ( .A1(\AES_ENC/us13/n843 ), .A2(\AES_ENC/us13/n842 ), .A3(\AES_ENC/us13/n841 ), .A4(\AES_ENC/us13/n840 ), .ZN(\AES_ENC/us13/n844 ) );
NOR2_X2 \AES_ENC/us13/U404  ( .A1(\AES_ENC/us13/n669 ), .A2(\AES_ENC/us13/n668 ), .ZN(\AES_ENC/us13/n673 ) );
NOR4_X2 \AES_ENC/us13/U403  ( .A1(\AES_ENC/us13/n946 ), .A2(\AES_ENC/us13/n1046 ), .A3(\AES_ENC/us13/n671 ), .A4(\AES_ENC/us13/n670 ), .ZN(\AES_ENC/us13/n672 ) );
NOR4_X2 \AES_ENC/us13/U401  ( .A1(\AES_ENC/us13/n711 ), .A2(\AES_ENC/us13/n710 ), .A3(\AES_ENC/us13/n709 ), .A4(\AES_ENC/us13/n708 ), .ZN(\AES_ENC/us13/n712 ) );
NOR4_X2 \AES_ENC/us13/U400  ( .A1(\AES_ENC/us13/n963 ), .A2(\AES_ENC/us13/n962 ), .A3(\AES_ENC/us13/n961 ), .A4(\AES_ENC/us13/n960 ), .ZN(\AES_ENC/us13/n964 ) );
NOR3_X2 \AES_ENC/us13/U399  ( .A1(\AES_ENC/us13/n1101 ), .A2(\AES_ENC/us13/n1100 ), .A3(\AES_ENC/us13/n1099 ), .ZN(\AES_ENC/us13/n1109 ) );
NOR3_X2 \AES_ENC/us13/U398  ( .A1(\AES_ENC/us13/n743 ), .A2(\AES_ENC/us13/n742 ), .A3(\AES_ENC/us13/n741 ), .ZN(\AES_ENC/us13/n744 ) );
NOR2_X2 \AES_ENC/us13/U397  ( .A1(\AES_ENC/us13/n697 ), .A2(\AES_ENC/us13/n658 ), .ZN(\AES_ENC/us13/n659 ) );
NOR2_X2 \AES_ENC/us13/U396  ( .A1(\AES_ENC/us13/n1078 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n1033 ) );
NOR2_X2 \AES_ENC/us13/U393  ( .A1(\AES_ENC/us13/n1031 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n1032 ) );
NOR3_X2 \AES_ENC/us13/U390  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n1025 ), .A3(\AES_ENC/us13/n1074 ), .ZN(\AES_ENC/us13/n1035 ) );
NOR4_X2 \AES_ENC/us13/U389  ( .A1(\AES_ENC/us13/n1035 ), .A2(\AES_ENC/us13/n1034 ), .A3(\AES_ENC/us13/n1033 ), .A4(\AES_ENC/us13/n1032 ), .ZN(\AES_ENC/us13/n1036 ) );
NOR2_X2 \AES_ENC/us13/U388  ( .A1(\AES_ENC/us13/n611 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n885 ) );
NOR2_X2 \AES_ENC/us13/U387  ( .A1(\AES_ENC/us13/n601 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n882 ) );
NOR2_X2 \AES_ENC/us13/U386  ( .A1(\AES_ENC/us13/n1053 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n884 ) );
NOR4_X2 \AES_ENC/us13/U385  ( .A1(\AES_ENC/us13/n885 ), .A2(\AES_ENC/us13/n884 ), .A3(\AES_ENC/us13/n883 ), .A4(\AES_ENC/us13/n882 ), .ZN(\AES_ENC/us13/n886 ) );
NOR2_X2 \AES_ENC/us13/U384  ( .A1(\AES_ENC/us13/n825 ), .A2(\AES_ENC/us13/n574 ), .ZN(\AES_ENC/us13/n830 ) );
NOR2_X2 \AES_ENC/us13/U383  ( .A1(\AES_ENC/us13/n827 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n829 ) );
NOR2_X2 \AES_ENC/us13/U382  ( .A1(\AES_ENC/us13/n572 ), .A2(\AES_ENC/us13/n575 ), .ZN(\AES_ENC/us13/n828 ) );
NOR4_X2 \AES_ENC/us13/U374  ( .A1(\AES_ENC/us13/n831 ), .A2(\AES_ENC/us13/n830 ), .A3(\AES_ENC/us13/n829 ), .A4(\AES_ENC/us13/n828 ), .ZN(\AES_ENC/us13/n832 ) );
NOR2_X2 \AES_ENC/us13/U373  ( .A1(\AES_ENC/us13/n578 ), .A2(\AES_ENC/us13/n603 ), .ZN(\AES_ENC/us13/n1104 ) );
NOR2_X2 \AES_ENC/us13/U372  ( .A1(\AES_ENC/us13/n1102 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n1106 ) );
NOR2_X2 \AES_ENC/us13/U370  ( .A1(\AES_ENC/us13/n1103 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n1105 ) );
NOR4_X2 \AES_ENC/us13/U369  ( .A1(\AES_ENC/us13/n1107 ), .A2(\AES_ENC/us13/n1106 ), .A3(\AES_ENC/us13/n1105 ), .A4(\AES_ENC/us13/n1104 ), .ZN(\AES_ENC/us13/n1108 ) );
NOR3_X2 \AES_ENC/us13/U368  ( .A1(\AES_ENC/us13/n959 ), .A2(\AES_ENC/us13/n624 ), .A3(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n963 ) );
NOR2_X2 \AES_ENC/us13/U367  ( .A1(\AES_ENC/us13/n594 ), .A2(\AES_ENC/us13/n595 ), .ZN(\AES_ENC/us13/n1114 ) );
INV_X4 \AES_ENC/us13/U366  ( .A(\AES_ENC/us13/n1024 ), .ZN(\AES_ENC/us13/n578 ) );
NOR3_X2 \AES_ENC/us13/U365  ( .A1(\AES_ENC/us13/n910 ), .A2(\AES_ENC/us13/n1059 ), .A3(\AES_ENC/us13/n584 ), .ZN(\AES_ENC/us13/n1115 ) );
INV_X4 \AES_ENC/us13/U364  ( .A(\AES_ENC/us13/n1094 ), .ZN(\AES_ENC/us13/n587 ) );
NOR2_X2 \AES_ENC/us13/U363  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n931 ), .ZN(\AES_ENC/us13/n1100 ) );
INV_X4 \AES_ENC/us13/U354  ( .A(\AES_ENC/us13/n1093 ), .ZN(\AES_ENC/us13/n591 ) );
NOR2_X2 \AES_ENC/us13/U353  ( .A1(\AES_ENC/us13/n569 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n929 ) );
NOR2_X2 \AES_ENC/us13/U352  ( .A1(\AES_ENC/us13/n609 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n926 ) );
NOR2_X2 \AES_ENC/us13/U351  ( .A1(\AES_ENC/us13/n572 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n1095 ) );
NOR2_X2 \AES_ENC/us13/U350  ( .A1(\AES_ENC/us13/n582 ), .A2(\AES_ENC/us13/n595 ), .ZN(\AES_ENC/us13/n1010 ) );
NOR2_X2 \AES_ENC/us13/U349  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n1103 ) );
NOR2_X2 \AES_ENC/us13/U348  ( .A1(\AES_ENC/us13/n614 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n1059 ) );
NOR2_X2 \AES_ENC/us13/U347  ( .A1(\AES_ENC/sa13 [1]), .A2(\AES_ENC/us13/n1120 ), .ZN(\AES_ENC/us13/n1022 ) );
NOR2_X2 \AES_ENC/us13/U346  ( .A1(\AES_ENC/us13/n605 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n911 ) );
NOR2_X2 \AES_ENC/us13/U345  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/us13/n1025 ), .ZN(\AES_ENC/us13/n826 ) );
NOR2_X2 \AES_ENC/us13/U338  ( .A1(\AES_ENC/us13/n594 ), .A2(\AES_ENC/us13/n579 ), .ZN(\AES_ENC/us13/n1072 ) );
NOR2_X2 \AES_ENC/us13/U335  ( .A1(\AES_ENC/us13/n595 ), .A2(\AES_ENC/us13/n590 ), .ZN(\AES_ENC/us13/n956 ) );
NOR2_X2 \AES_ENC/us13/U329  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/us13/n612 ), .ZN(\AES_ENC/us13/n1121 ) );
NOR2_X2 \AES_ENC/us13/U328  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/us13/n612 ), .ZN(\AES_ENC/us13/n1058 ) );
NOR2_X2 \AES_ENC/us13/U327  ( .A1(\AES_ENC/us13/n593 ), .A2(\AES_ENC/us13/n584 ), .ZN(\AES_ENC/us13/n1073 ) );
NOR2_X2 \AES_ENC/us13/U325  ( .A1(\AES_ENC/sa13 [1]), .A2(\AES_ENC/us13/n1025 ), .ZN(\AES_ENC/us13/n1054 ) );
NOR2_X2 \AES_ENC/us13/U324  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/us13/n931 ), .ZN(\AES_ENC/us13/n1029 ) );
NOR2_X2 \AES_ENC/us13/U319  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n1056 ) );
NOR2_X2 \AES_ENC/us13/U318  ( .A1(\AES_ENC/us13/n588 ), .A2(\AES_ENC/us13/n594 ), .ZN(\AES_ENC/us13/n1050 ) );
NOR2_X2 \AES_ENC/us13/U317  ( .A1(\AES_ENC/us13/n1121 ), .A2(\AES_ENC/us13/n1025 ), .ZN(\AES_ENC/us13/n1120 ) );
NOR2_X2 \AES_ENC/us13/U316  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/us13/n572 ), .ZN(\AES_ENC/us13/n1074 ) );
NOR2_X2 \AES_ENC/us13/U315  ( .A1(\AES_ENC/us13/n1058 ), .A2(\AES_ENC/us13/n1054 ), .ZN(\AES_ENC/us13/n878 ) );
NOR2_X2 \AES_ENC/us13/U314  ( .A1(\AES_ENC/us13/n878 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n879 ) );
NOR2_X2 \AES_ENC/us13/U312  ( .A1(\AES_ENC/us13/n880 ), .A2(\AES_ENC/us13/n879 ), .ZN(\AES_ENC/us13/n887 ) );
NOR2_X2 \AES_ENC/us13/U311  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n625 ), .ZN(\AES_ENC/us13/n957 ) );
NOR2_X2 \AES_ENC/us13/U310  ( .A1(\AES_ENC/us13/n958 ), .A2(\AES_ENC/us13/n957 ), .ZN(\AES_ENC/us13/n965 ) );
NOR3_X2 \AES_ENC/us13/U309  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n1091 ), .A3(\AES_ENC/us13/n1022 ), .ZN(\AES_ENC/us13/n720 ) );
NOR3_X2 \AES_ENC/us13/U303  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n1054 ), .A3(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n719 ) );
NOR2_X2 \AES_ENC/us13/U302  ( .A1(\AES_ENC/us13/n720 ), .A2(\AES_ENC/us13/n719 ), .ZN(\AES_ENC/us13/n726 ) );
NOR2_X2 \AES_ENC/us13/U300  ( .A1(\AES_ENC/us13/n588 ), .A2(\AES_ENC/us13/n613 ), .ZN(\AES_ENC/us13/n865 ) );
NOR2_X2 \AES_ENC/us13/U299  ( .A1(\AES_ENC/us13/n1059 ), .A2(\AES_ENC/us13/n1058 ), .ZN(\AES_ENC/us13/n1060 ) );
NOR2_X2 \AES_ENC/us13/U298  ( .A1(\AES_ENC/us13/n1095 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n668 ) );
NOR2_X2 \AES_ENC/us13/U297  ( .A1(\AES_ENC/us13/n911 ), .A2(\AES_ENC/us13/n910 ), .ZN(\AES_ENC/us13/n912 ) );
NOR2_X2 \AES_ENC/us13/U296  ( .A1(\AES_ENC/us13/n912 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n916 ) );
NOR2_X2 \AES_ENC/us13/U295  ( .A1(\AES_ENC/us13/n826 ), .A2(\AES_ENC/us13/n573 ), .ZN(\AES_ENC/us13/n750 ) );
NOR2_X2 \AES_ENC/us13/U294  ( .A1(\AES_ENC/us13/n750 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n751 ) );
NOR2_X2 \AES_ENC/us13/U293  ( .A1(\AES_ENC/us13/n907 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n908 ) );
NOR2_X2 \AES_ENC/us13/U292  ( .A1(\AES_ENC/us13/n990 ), .A2(\AES_ENC/us13/n926 ), .ZN(\AES_ENC/us13/n780 ) );
NOR2_X2 \AES_ENC/us13/U291  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n606 ), .ZN(\AES_ENC/us13/n838 ) );
NOR2_X2 \AES_ENC/us13/U290  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n621 ), .ZN(\AES_ENC/us13/n837 ) );
NOR2_X2 \AES_ENC/us13/U284  ( .A1(\AES_ENC/us13/n838 ), .A2(\AES_ENC/us13/n837 ), .ZN(\AES_ENC/us13/n845 ) );
NOR2_X2 \AES_ENC/us13/U283  ( .A1(\AES_ENC/us13/n1022 ), .A2(\AES_ENC/us13/n1058 ), .ZN(\AES_ENC/us13/n740 ) );
NOR2_X2 \AES_ENC/us13/U282  ( .A1(\AES_ENC/us13/n740 ), .A2(\AES_ENC/us13/n590 ), .ZN(\AES_ENC/us13/n742 ) );
NOR2_X2 \AES_ENC/us13/U281  ( .A1(\AES_ENC/us13/n1098 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n1099 ) );
NOR2_X2 \AES_ENC/us13/U280  ( .A1(\AES_ENC/us13/n1120 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n993 ) );
NOR2_X2 \AES_ENC/us13/U279  ( .A1(\AES_ENC/us13/n993 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n994 ) );
NOR2_X2 \AES_ENC/us13/U273  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n609 ), .ZN(\AES_ENC/us13/n1026 ) );
NOR2_X2 \AES_ENC/us13/U272  ( .A1(\AES_ENC/us13/n573 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n1027 ) );
NOR2_X2 \AES_ENC/us13/U271  ( .A1(\AES_ENC/us13/n1027 ), .A2(\AES_ENC/us13/n1026 ), .ZN(\AES_ENC/us13/n1028 ) );
NOR2_X2 \AES_ENC/us13/U270  ( .A1(\AES_ENC/us13/n1029 ), .A2(\AES_ENC/us13/n1028 ), .ZN(\AES_ENC/us13/n1034 ) );
NOR4_X2 \AES_ENC/us13/U269  ( .A1(\AES_ENC/us13/n757 ), .A2(\AES_ENC/us13/n756 ), .A3(\AES_ENC/us13/n755 ), .A4(\AES_ENC/us13/n754 ), .ZN(\AES_ENC/us13/n758 ) );
NOR2_X2 \AES_ENC/us13/U268  ( .A1(\AES_ENC/us13/n752 ), .A2(\AES_ENC/us13/n751 ), .ZN(\AES_ENC/us13/n759 ) );
NOR2_X2 \AES_ENC/us13/U267  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n1071 ), .ZN(\AES_ENC/us13/n669 ) );
NOR2_X2 \AES_ENC/us13/U263  ( .A1(\AES_ENC/us13/n1056 ), .A2(\AES_ENC/us13/n990 ), .ZN(\AES_ENC/us13/n991 ) );
NOR2_X2 \AES_ENC/us13/U262  ( .A1(\AES_ENC/us13/n991 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n995 ) );
NOR2_X2 \AES_ENC/us13/U258  ( .A1(\AES_ENC/us13/n579 ), .A2(\AES_ENC/us13/n598 ), .ZN(\AES_ENC/us13/n1008 ) );
NOR2_X2 \AES_ENC/us13/U255  ( .A1(\AES_ENC/us13/n839 ), .A2(\AES_ENC/us13/n603 ), .ZN(\AES_ENC/us13/n693 ) );
NOR2_X2 \AES_ENC/us13/U254  ( .A1(\AES_ENC/us13/n578 ), .A2(\AES_ENC/us13/n906 ), .ZN(\AES_ENC/us13/n741 ) );
NOR2_X2 \AES_ENC/us13/U253  ( .A1(\AES_ENC/us13/n1054 ), .A2(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n763 ) );
NOR2_X2 \AES_ENC/us13/U252  ( .A1(\AES_ENC/us13/n763 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n769 ) );
NOR2_X2 \AES_ENC/us13/U251  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n618 ), .ZN(\AES_ENC/us13/n1007 ) );
NOR2_X2 \AES_ENC/us13/U250  ( .A1(\AES_ENC/us13/n582 ), .A2(\AES_ENC/us13/n599 ), .ZN(\AES_ENC/us13/n1123 ) );
NOR2_X2 \AES_ENC/us13/U243  ( .A1(\AES_ENC/us13/n582 ), .A2(\AES_ENC/us13/n598 ), .ZN(\AES_ENC/us13/n710 ) );
INV_X4 \AES_ENC/us13/U242  ( .A(\AES_ENC/us13/n1029 ), .ZN(\AES_ENC/us13/n603 ) );
NOR2_X2 \AES_ENC/us13/U241  ( .A1(\AES_ENC/us13/n590 ), .A2(\AES_ENC/us13/n607 ), .ZN(\AES_ENC/us13/n883 ) );
NOR2_X2 \AES_ENC/us13/U240  ( .A1(\AES_ENC/us13/n623 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n1125 ) );
NOR2_X2 \AES_ENC/us13/U239  ( .A1(\AES_ENC/us13/n990 ), .A2(\AES_ENC/us13/n929 ), .ZN(\AES_ENC/us13/n892 ) );
NOR2_X2 \AES_ENC/us13/U238  ( .A1(\AES_ENC/us13/n892 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n893 ) );
NOR2_X2 \AES_ENC/us13/U237  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n621 ), .ZN(\AES_ENC/us13/n950 ) );
NOR2_X2 \AES_ENC/us13/U236  ( .A1(\AES_ENC/us13/n1079 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n1082 ) );
NOR2_X2 \AES_ENC/us13/U235  ( .A1(\AES_ENC/us13/n910 ), .A2(\AES_ENC/us13/n1056 ), .ZN(\AES_ENC/us13/n941 ) );
NOR2_X2 \AES_ENC/us13/U234  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n1077 ), .ZN(\AES_ENC/us13/n841 ) );
NOR2_X2 \AES_ENC/us13/U229  ( .A1(\AES_ENC/us13/n601 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n630 ) );
NOR2_X2 \AES_ENC/us13/U228  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n621 ), .ZN(\AES_ENC/us13/n806 ) );
NOR2_X2 \AES_ENC/us13/U227  ( .A1(\AES_ENC/us13/n601 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n948 ) );
NOR2_X2 \AES_ENC/us13/U226  ( .A1(\AES_ENC/us13/n578 ), .A2(\AES_ENC/us13/n620 ), .ZN(\AES_ENC/us13/n997 ) );
NOR2_X2 \AES_ENC/us13/U225  ( .A1(\AES_ENC/us13/n1121 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n1122 ) );
NOR2_X2 \AES_ENC/us13/U223  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n1023 ), .ZN(\AES_ENC/us13/n756 ) );
NOR2_X2 \AES_ENC/us13/U222  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n621 ), .ZN(\AES_ENC/us13/n870 ) );
NOR2_X2 \AES_ENC/us13/U221  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n569 ), .ZN(\AES_ENC/us13/n947 ) );
NOR2_X2 \AES_ENC/us13/U217  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n1077 ), .ZN(\AES_ENC/us13/n1084 ) );
NOR2_X2 \AES_ENC/us13/U213  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n855 ), .ZN(\AES_ENC/us13/n709 ) );
NOR2_X2 \AES_ENC/us13/U212  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n620 ), .ZN(\AES_ENC/us13/n868 ) );
NOR2_X2 \AES_ENC/us13/U211  ( .A1(\AES_ENC/us13/n1120 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n1124 ) );
NOR2_X2 \AES_ENC/us13/U210  ( .A1(\AES_ENC/us13/n1120 ), .A2(\AES_ENC/us13/n839 ), .ZN(\AES_ENC/us13/n842 ) );
NOR2_X2 \AES_ENC/us13/U209  ( .A1(\AES_ENC/us13/n1120 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n696 ) );
NOR2_X2 \AES_ENC/us13/U208  ( .A1(\AES_ENC/us13/n1074 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n1076 ) );
NOR2_X2 \AES_ENC/us13/U207  ( .A1(\AES_ENC/us13/n1074 ), .A2(\AES_ENC/us13/n609 ), .ZN(\AES_ENC/us13/n781 ) );
NOR3_X2 \AES_ENC/us13/U201  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n1056 ), .A3(\AES_ENC/us13/n990 ), .ZN(\AES_ENC/us13/n979 ) );
NOR3_X2 \AES_ENC/us13/U200  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n1058 ), .A3(\AES_ENC/us13/n1059 ), .ZN(\AES_ENC/us13/n854 ) );
NOR2_X2 \AES_ENC/us13/U199  ( .A1(\AES_ENC/us13/n996 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n869 ) );
NOR2_X2 \AES_ENC/us13/U198  ( .A1(\AES_ENC/us13/n1056 ), .A2(\AES_ENC/us13/n1074 ), .ZN(\AES_ENC/us13/n1057 ) );
NOR3_X2 \AES_ENC/us13/U197  ( .A1(\AES_ENC/us13/n579 ), .A2(\AES_ENC/us13/n1120 ), .A3(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n978 ) );
NOR2_X2 \AES_ENC/us13/U196  ( .A1(\AES_ENC/us13/n996 ), .A2(\AES_ENC/us13/n911 ), .ZN(\AES_ENC/us13/n1116 ) );
NOR2_X2 \AES_ENC/us13/U195  ( .A1(\AES_ENC/us13/n1074 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n754 ) );
NOR2_X2 \AES_ENC/us13/U194  ( .A1(\AES_ENC/us13/n926 ), .A2(\AES_ENC/us13/n1103 ), .ZN(\AES_ENC/us13/n977 ) );
NOR2_X2 \AES_ENC/us13/U187  ( .A1(\AES_ENC/us13/n839 ), .A2(\AES_ENC/us13/n824 ), .ZN(\AES_ENC/us13/n1092 ) );
NOR2_X2 \AES_ENC/us13/U186  ( .A1(\AES_ENC/us13/n573 ), .A2(\AES_ENC/us13/n1074 ), .ZN(\AES_ENC/us13/n684 ) );
NOR2_X2 \AES_ENC/us13/U185  ( .A1(\AES_ENC/us13/n826 ), .A2(\AES_ENC/us13/n1059 ), .ZN(\AES_ENC/us13/n907 ) );
NOR3_X2 \AES_ENC/us13/U184  ( .A1(\AES_ENC/us13/n593 ), .A2(\AES_ENC/us13/n1115 ), .A3(\AES_ENC/us13/n600 ), .ZN(\AES_ENC/us13/n831 ) );
NOR3_X2 \AES_ENC/us13/U183  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n1056 ), .A3(\AES_ENC/us13/n990 ), .ZN(\AES_ENC/us13/n896 ) );
NOR3_X2 \AES_ENC/us13/U182  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n573 ), .A3(\AES_ENC/us13/n1013 ), .ZN(\AES_ENC/us13/n670 ) );
NOR3_X2 \AES_ENC/us13/U181  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n1091 ), .A3(\AES_ENC/us13/n1022 ), .ZN(\AES_ENC/us13/n843 ) );
NOR2_X2 \AES_ENC/us13/U180  ( .A1(\AES_ENC/us13/n1029 ), .A2(\AES_ENC/us13/n1095 ), .ZN(\AES_ENC/us13/n735 ) );
NOR2_X2 \AES_ENC/us13/U174  ( .A1(\AES_ENC/us13/n1100 ), .A2(\AES_ENC/us13/n854 ), .ZN(\AES_ENC/us13/n860 ) );
NAND3_X2 \AES_ENC/us13/U173  ( .A1(\AES_ENC/us13/n569 ), .A2(\AES_ENC/us13/n603 ), .A3(\AES_ENC/us13/n681 ), .ZN(\AES_ENC/us13/n691 ) );
NOR2_X2 \AES_ENC/us13/U172  ( .A1(\AES_ENC/us13/n683 ), .A2(\AES_ENC/us13/n682 ), .ZN(\AES_ENC/us13/n690 ) );
NOR3_X2 \AES_ENC/us13/U171  ( .A1(\AES_ENC/us13/n695 ), .A2(\AES_ENC/us13/n694 ), .A3(\AES_ENC/us13/n693 ), .ZN(\AES_ENC/us13/n700 ) );
NOR4_X2 \AES_ENC/us13/U170  ( .A1(\AES_ENC/us13/n983 ), .A2(\AES_ENC/us13/n698 ), .A3(\AES_ENC/us13/n697 ), .A4(\AES_ENC/us13/n696 ), .ZN(\AES_ENC/us13/n699 ) );
NOR2_X2 \AES_ENC/us13/U169  ( .A1(\AES_ENC/us13/n946 ), .A2(\AES_ENC/us13/n945 ), .ZN(\AES_ENC/us13/n952 ) );
NOR4_X2 \AES_ENC/us13/U168  ( .A1(\AES_ENC/us13/n950 ), .A2(\AES_ENC/us13/n949 ), .A3(\AES_ENC/us13/n948 ), .A4(\AES_ENC/us13/n947 ), .ZN(\AES_ENC/us13/n951 ) );
NOR4_X2 \AES_ENC/us13/U162  ( .A1(\AES_ENC/us13/n983 ), .A2(\AES_ENC/us13/n982 ), .A3(\AES_ENC/us13/n981 ), .A4(\AES_ENC/us13/n980 ), .ZN(\AES_ENC/us13/n984 ) );
NOR2_X2 \AES_ENC/us13/U161  ( .A1(\AES_ENC/us13/n979 ), .A2(\AES_ENC/us13/n978 ), .ZN(\AES_ENC/us13/n985 ) );
NOR4_X2 \AES_ENC/us13/U160  ( .A1(\AES_ENC/us13/n896 ), .A2(\AES_ENC/us13/n895 ), .A3(\AES_ENC/us13/n894 ), .A4(\AES_ENC/us13/n893 ), .ZN(\AES_ENC/us13/n897 ) );
NOR2_X2 \AES_ENC/us13/U159  ( .A1(\AES_ENC/us13/n866 ), .A2(\AES_ENC/us13/n865 ), .ZN(\AES_ENC/us13/n872 ) );
NOR4_X2 \AES_ENC/us13/U158  ( .A1(\AES_ENC/us13/n870 ), .A2(\AES_ENC/us13/n869 ), .A3(\AES_ENC/us13/n868 ), .A4(\AES_ENC/us13/n867 ), .ZN(\AES_ENC/us13/n871 ) );
NOR4_X2 \AES_ENC/us13/U157  ( .A1(\AES_ENC/us13/n1125 ), .A2(\AES_ENC/us13/n1124 ), .A3(\AES_ENC/us13/n1123 ), .A4(\AES_ENC/us13/n1122 ), .ZN(\AES_ENC/us13/n1126 ) );
NOR4_X2 \AES_ENC/us13/U156  ( .A1(\AES_ENC/us13/n1084 ), .A2(\AES_ENC/us13/n1083 ), .A3(\AES_ENC/us13/n1082 ), .A4(\AES_ENC/us13/n1081 ), .ZN(\AES_ENC/us13/n1085 ) );
NOR2_X2 \AES_ENC/us13/U155  ( .A1(\AES_ENC/us13/n1076 ), .A2(\AES_ENC/us13/n1075 ), .ZN(\AES_ENC/us13/n1086 ) );
NOR3_X2 \AES_ENC/us13/U154  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n1054 ), .A3(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n961 ) );
NOR3_X2 \AES_ENC/us13/U153  ( .A1(\AES_ENC/us13/n609 ), .A2(\AES_ENC/us13/n1074 ), .A3(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n671 ) );
NOR2_X2 \AES_ENC/us13/U152  ( .A1(\AES_ENC/us13/n1057 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n1062 ) );
NOR2_X2 \AES_ENC/us13/U143  ( .A1(\AES_ENC/us13/n1055 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n1063 ) );
NOR2_X2 \AES_ENC/us13/U142  ( .A1(\AES_ENC/us13/n1060 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n1061 ) );
NOR4_X2 \AES_ENC/us13/U141  ( .A1(\AES_ENC/us13/n1064 ), .A2(\AES_ENC/us13/n1063 ), .A3(\AES_ENC/us13/n1062 ), .A4(\AES_ENC/us13/n1061 ), .ZN(\AES_ENC/us13/n1065 ) );
NOR3_X2 \AES_ENC/us13/U140  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n1120 ), .A3(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n918 ) );
NOR3_X2 \AES_ENC/us13/U132  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n573 ), .A3(\AES_ENC/us13/n1013 ), .ZN(\AES_ENC/us13/n917 ) );
NOR2_X2 \AES_ENC/us13/U131  ( .A1(\AES_ENC/us13/n914 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n915 ) );
NOR4_X2 \AES_ENC/us13/U130  ( .A1(\AES_ENC/us13/n918 ), .A2(\AES_ENC/us13/n917 ), .A3(\AES_ENC/us13/n916 ), .A4(\AES_ENC/us13/n915 ), .ZN(\AES_ENC/us13/n919 ) );
NOR2_X2 \AES_ENC/us13/U129  ( .A1(\AES_ENC/us13/n590 ), .A2(\AES_ENC/us13/n599 ), .ZN(\AES_ENC/us13/n771 ) );
NOR2_X2 \AES_ENC/us13/U128  ( .A1(\AES_ENC/us13/n1103 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n772 ) );
NOR2_X2 \AES_ENC/us13/U127  ( .A1(\AES_ENC/us13/n583 ), .A2(\AES_ENC/us13/n615 ), .ZN(\AES_ENC/us13/n773 ) );
NOR4_X2 \AES_ENC/us13/U126  ( .A1(\AES_ENC/us13/n773 ), .A2(\AES_ENC/us13/n772 ), .A3(\AES_ENC/us13/n771 ), .A4(\AES_ENC/us13/n770 ), .ZN(\AES_ENC/us13/n774 ) );
NOR2_X2 \AES_ENC/us13/U121  ( .A1(\AES_ENC/us13/n735 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n687 ) );
NOR2_X2 \AES_ENC/us13/U120  ( .A1(\AES_ENC/us13/n684 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n688 ) );
NOR2_X2 \AES_ENC/us13/U119  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n622 ), .ZN(\AES_ENC/us13/n686 ) );
NOR4_X2 \AES_ENC/us13/U118  ( .A1(\AES_ENC/us13/n688 ), .A2(\AES_ENC/us13/n687 ), .A3(\AES_ENC/us13/n686 ), .A4(\AES_ENC/us13/n685 ), .ZN(\AES_ENC/us13/n689 ) );
NOR2_X2 \AES_ENC/us13/U117  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n608 ), .ZN(\AES_ENC/us13/n858 ) );
NOR2_X2 \AES_ENC/us13/U116  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n855 ), .ZN(\AES_ENC/us13/n857 ) );
NOR2_X2 \AES_ENC/us13/U115  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n617 ), .ZN(\AES_ENC/us13/n856 ) );
NOR4_X2 \AES_ENC/us13/U106  ( .A1(\AES_ENC/us13/n858 ), .A2(\AES_ENC/us13/n857 ), .A3(\AES_ENC/us13/n856 ), .A4(\AES_ENC/us13/n958 ), .ZN(\AES_ENC/us13/n859 ) );
NOR2_X2 \AES_ENC/us13/U105  ( .A1(\AES_ENC/us13/n780 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n784 ) );
NOR2_X2 \AES_ENC/us13/U104  ( .A1(\AES_ENC/us13/n1117 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n782 ) );
NOR2_X2 \AES_ENC/us13/U103  ( .A1(\AES_ENC/us13/n781 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n783 ) );
NOR4_X2 \AES_ENC/us13/U102  ( .A1(\AES_ENC/us13/n880 ), .A2(\AES_ENC/us13/n784 ), .A3(\AES_ENC/us13/n783 ), .A4(\AES_ENC/us13/n782 ), .ZN(\AES_ENC/us13/n785 ) );
NOR2_X2 \AES_ENC/us13/U101  ( .A1(\AES_ENC/us13/n597 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n814 ) );
NOR2_X2 \AES_ENC/us13/U100  ( .A1(\AES_ENC/us13/n907 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n813 ) );
NOR3_X2 \AES_ENC/us13/U95  ( .A1(\AES_ENC/us13/n578 ), .A2(\AES_ENC/us13/n1058 ), .A3(\AES_ENC/us13/n1059 ), .ZN(\AES_ENC/us13/n815 ) );
NOR4_X2 \AES_ENC/us13/U94  ( .A1(\AES_ENC/us13/n815 ), .A2(\AES_ENC/us13/n814 ), .A3(\AES_ENC/us13/n813 ), .A4(\AES_ENC/us13/n812 ), .ZN(\AES_ENC/us13/n816 ) );
NOR2_X2 \AES_ENC/us13/U93  ( .A1(\AES_ENC/us13/n591 ), .A2(\AES_ENC/us13/n569 ), .ZN(\AES_ENC/us13/n721 ) );
NOR2_X2 \AES_ENC/us13/U92  ( .A1(\AES_ENC/us13/n1031 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n723 ) );
NOR2_X2 \AES_ENC/us13/U91  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n1096 ), .ZN(\AES_ENC/us13/n722 ) );
NOR4_X2 \AES_ENC/us13/U90  ( .A1(\AES_ENC/us13/n724 ), .A2(\AES_ENC/us13/n723 ), .A3(\AES_ENC/us13/n722 ), .A4(\AES_ENC/us13/n721 ), .ZN(\AES_ENC/us13/n725 ) );
NOR2_X2 \AES_ENC/us13/U89  ( .A1(\AES_ENC/us13/n911 ), .A2(\AES_ENC/us13/n990 ), .ZN(\AES_ENC/us13/n1009 ) );
NOR2_X2 \AES_ENC/us13/U88  ( .A1(\AES_ENC/us13/n1013 ), .A2(\AES_ENC/us13/n573 ), .ZN(\AES_ENC/us13/n1014 ) );
NOR2_X2 \AES_ENC/us13/U87  ( .A1(\AES_ENC/us13/n1014 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n1015 ) );
NOR4_X2 \AES_ENC/us13/U86  ( .A1(\AES_ENC/us13/n1016 ), .A2(\AES_ENC/us13/n1015 ), .A3(\AES_ENC/us13/n1119 ), .A4(\AES_ENC/us13/n1046 ), .ZN(\AES_ENC/us13/n1017 ) );
NOR2_X2 \AES_ENC/us13/U81  ( .A1(\AES_ENC/us13/n996 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n998 ) );
NOR2_X2 \AES_ENC/us13/U80  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n618 ), .ZN(\AES_ENC/us13/n1000 ) );
NOR2_X2 \AES_ENC/us13/U79  ( .A1(\AES_ENC/us13/n590 ), .A2(\AES_ENC/us13/n1096 ), .ZN(\AES_ENC/us13/n999 ) );
NOR4_X2 \AES_ENC/us13/U78  ( .A1(\AES_ENC/us13/n1000 ), .A2(\AES_ENC/us13/n999 ), .A3(\AES_ENC/us13/n998 ), .A4(\AES_ENC/us13/n997 ), .ZN(\AES_ENC/us13/n1001 ) );
NOR2_X2 \AES_ENC/us13/U74  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n1096 ), .ZN(\AES_ENC/us13/n697 ) );
NOR2_X2 \AES_ENC/us13/U73  ( .A1(\AES_ENC/us13/n609 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n958 ) );
NOR2_X2 \AES_ENC/us13/U72  ( .A1(\AES_ENC/us13/n911 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n983 ) );
NOR2_X2 \AES_ENC/us13/U71  ( .A1(\AES_ENC/us13/n1054 ), .A2(\AES_ENC/us13/n1103 ), .ZN(\AES_ENC/us13/n1031 ) );
INV_X4 \AES_ENC/us13/U65  ( .A(\AES_ENC/us13/n1050 ), .ZN(\AES_ENC/us13/n585 ) );
INV_X4 \AES_ENC/us13/U64  ( .A(\AES_ENC/us13/n1072 ), .ZN(\AES_ENC/us13/n577 ) );
INV_X4 \AES_ENC/us13/U63  ( .A(\AES_ENC/us13/n1073 ), .ZN(\AES_ENC/us13/n576 ) );
NOR2_X2 \AES_ENC/us13/U62  ( .A1(\AES_ENC/us13/n603 ), .A2(\AES_ENC/us13/n587 ), .ZN(\AES_ENC/us13/n880 ) );
NOR3_X2 \AES_ENC/us13/U61  ( .A1(\AES_ENC/us13/n826 ), .A2(\AES_ENC/us13/n1121 ), .A3(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n946 ) );
INV_X4 \AES_ENC/us13/U59  ( .A(\AES_ENC/us13/n1010 ), .ZN(\AES_ENC/us13/n581 ) );
NOR3_X2 \AES_ENC/us13/U58  ( .A1(\AES_ENC/us13/n573 ), .A2(\AES_ENC/us13/n1029 ), .A3(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n1119 ) );
INV_X4 \AES_ENC/us13/U57  ( .A(\AES_ENC/us13/n956 ), .ZN(\AES_ENC/us13/n589 ) );
NOR2_X2 \AES_ENC/us13/U50  ( .A1(\AES_ENC/us13/n601 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n1013 ) );
NOR2_X2 \AES_ENC/us13/U49  ( .A1(\AES_ENC/us13/n609 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n910 ) );
NOR2_X2 \AES_ENC/us13/U48  ( .A1(\AES_ENC/us13/n569 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n1091 ) );
NOR2_X2 \AES_ENC/us13/U47  ( .A1(\AES_ENC/us13/n614 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n990 ) );
NOR2_X2 \AES_ENC/us13/U46  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/us13/n1121 ), .ZN(\AES_ENC/us13/n996 ) );
NOR2_X2 \AES_ENC/us13/U45  ( .A1(\AES_ENC/us13/n583 ), .A2(\AES_ENC/us13/n622 ), .ZN(\AES_ENC/us13/n628 ) );
NOR2_X2 \AES_ENC/us13/U44  ( .A1(\AES_ENC/us13/n602 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n866 ) );
NOR2_X2 \AES_ENC/us13/U43  ( .A1(\AES_ENC/us13/n610 ), .A2(\AES_ENC/us13/n583 ), .ZN(\AES_ENC/us13/n1006 ) );
NOR2_X2 \AES_ENC/us13/U42  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n1117 ), .ZN(\AES_ENC/us13/n1118 ) );
NOR2_X2 \AES_ENC/us13/U41  ( .A1(\AES_ENC/us13/n1119 ), .A2(\AES_ENC/us13/n1118 ), .ZN(\AES_ENC/us13/n1127 ) );
NOR2_X2 \AES_ENC/us13/U36  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n616 ), .ZN(\AES_ENC/us13/n629 ) );
NOR2_X2 \AES_ENC/us13/U35  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n906 ), .ZN(\AES_ENC/us13/n909 ) );
NOR2_X2 \AES_ENC/us13/U34  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n607 ), .ZN(\AES_ENC/us13/n658 ) );
NOR2_X2 \AES_ENC/us13/U33  ( .A1(\AES_ENC/us13/n1116 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n695 ) );
NOR2_X2 \AES_ENC/us13/U32  ( .A1(\AES_ENC/us13/n1078 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n1083 ) );
NOR2_X2 \AES_ENC/us13/U31  ( .A1(\AES_ENC/us13/n941 ), .A2(\AES_ENC/us13/n581 ), .ZN(\AES_ENC/us13/n724 ) );
NOR2_X2 \AES_ENC/us13/U30  ( .A1(\AES_ENC/us13/n611 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n1107 ) );
NOR2_X2 \AES_ENC/us13/U29  ( .A1(\AES_ENC/us13/n602 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n840 ) );
NOR2_X2 \AES_ENC/us13/U24  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n623 ), .ZN(\AES_ENC/us13/n633 ) );
NOR2_X2 \AES_ENC/us13/U23  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n1080 ), .ZN(\AES_ENC/us13/n1081 ) );
NOR2_X2 \AES_ENC/us13/U21  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n1045 ), .ZN(\AES_ENC/us13/n812 ) );
NOR2_X2 \AES_ENC/us13/U20  ( .A1(\AES_ENC/us13/n1009 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n960 ) );
NOR2_X2 \AES_ENC/us13/U19  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n619 ), .ZN(\AES_ENC/us13/n982 ) );
NOR2_X2 \AES_ENC/us13/U18  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n616 ), .ZN(\AES_ENC/us13/n757 ) );
NOR2_X2 \AES_ENC/us13/U17  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n598 ), .ZN(\AES_ENC/us13/n698 ) );
NOR2_X2 \AES_ENC/us13/U16  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n605 ), .ZN(\AES_ENC/us13/n708 ) );
NOR2_X2 \AES_ENC/us13/U15  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n603 ), .ZN(\AES_ENC/us13/n770 ) );
NOR2_X2 \AES_ENC/us13/U10  ( .A1(\AES_ENC/us13/n605 ), .A2(\AES_ENC/us13/n576 ), .ZN(\AES_ENC/us13/n803 ) );
NOR2_X2 \AES_ENC/us13/U9  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n881 ), .ZN(\AES_ENC/us13/n711 ) );
NOR2_X2 \AES_ENC/us13/U8  ( .A1(\AES_ENC/us13/n589 ), .A2(\AES_ENC/us13/n603 ), .ZN(\AES_ENC/us13/n867 ) );
NOR2_X2 \AES_ENC/us13/U7  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n615 ), .ZN(\AES_ENC/us13/n804 ) );
NOR2_X2 \AES_ENC/us13/U6  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n609 ), .ZN(\AES_ENC/us13/n1046 ) );
OR2_X4 \AES_ENC/us13/U5  ( .A1(\AES_ENC/us13/n612 ), .A2(\AES_ENC/sa13 [1]),.ZN(\AES_ENC/us13/n570 ) );
OR2_X4 \AES_ENC/us13/U4  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/sa13 [4]),.ZN(\AES_ENC/us13/n569 ) );
NAND2_X2 \AES_ENC/us13/U514  ( .A1(\AES_ENC/us13/n1121 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n1030 ) );
AND2_X2 \AES_ENC/us13/U513  ( .A1(\AES_ENC/us13/n607 ), .A2(\AES_ENC/us13/n1030 ), .ZN(\AES_ENC/us13/n1049 ) );
NAND2_X2 \AES_ENC/us13/U511  ( .A1(\AES_ENC/us13/n1049 ), .A2(\AES_ENC/us13/n794 ), .ZN(\AES_ENC/us13/n637 ) );
AND2_X2 \AES_ENC/us13/U493  ( .A1(\AES_ENC/us13/n779 ), .A2(\AES_ENC/us13/n996 ), .ZN(\AES_ENC/us13/n632 ) );
NAND4_X2 \AES_ENC/us13/U485  ( .A1(\AES_ENC/us13/n637 ), .A2(\AES_ENC/us13/n636 ), .A3(\AES_ENC/us13/n635 ), .A4(\AES_ENC/us13/n634 ), .ZN(\AES_ENC/us13/n638 ) );
NAND2_X2 \AES_ENC/us13/U484  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n638 ), .ZN(\AES_ENC/us13/n679 ) );
NAND2_X2 \AES_ENC/us13/U481  ( .A1(\AES_ENC/us13/n1094 ), .A2(\AES_ENC/us13/n613 ), .ZN(\AES_ENC/us13/n648 ) );
NAND2_X2 \AES_ENC/us13/U476  ( .A1(\AES_ENC/us13/n619 ), .A2(\AES_ENC/us13/n598 ), .ZN(\AES_ENC/us13/n762 ) );
NAND2_X2 \AES_ENC/us13/U475  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n762 ), .ZN(\AES_ENC/us13/n647 ) );
NAND4_X2 \AES_ENC/us13/U457  ( .A1(\AES_ENC/us13/n648 ), .A2(\AES_ENC/us13/n647 ), .A3(\AES_ENC/us13/n646 ), .A4(\AES_ENC/us13/n645 ), .ZN(\AES_ENC/us13/n649 ) );
NAND2_X2 \AES_ENC/us13/U456  ( .A1(\AES_ENC/sa13 [0]), .A2(\AES_ENC/us13/n649 ), .ZN(\AES_ENC/us13/n665 ) );
NAND2_X2 \AES_ENC/us13/U454  ( .A1(\AES_ENC/us13/n626 ), .A2(\AES_ENC/us13/n601 ), .ZN(\AES_ENC/us13/n855 ) );
NAND2_X2 \AES_ENC/us13/U453  ( .A1(\AES_ENC/us13/n617 ), .A2(\AES_ENC/us13/n855 ), .ZN(\AES_ENC/us13/n821 ) );
NAND2_X2 \AES_ENC/us13/U452  ( .A1(\AES_ENC/us13/n1093 ), .A2(\AES_ENC/us13/n821 ), .ZN(\AES_ENC/us13/n662 ) );
NAND2_X2 \AES_ENC/us13/U451  ( .A1(\AES_ENC/us13/n605 ), .A2(\AES_ENC/us13/n620 ), .ZN(\AES_ENC/us13/n650 ) );
NAND2_X2 \AES_ENC/us13/U450  ( .A1(\AES_ENC/us13/n956 ), .A2(\AES_ENC/us13/n650 ), .ZN(\AES_ENC/us13/n661 ) );
NAND2_X2 \AES_ENC/us13/U449  ( .A1(\AES_ENC/us13/n594 ), .A2(\AES_ENC/us13/n595 ), .ZN(\AES_ENC/us13/n839 ) );
OR2_X2 \AES_ENC/us13/U446  ( .A1(\AES_ENC/us13/n839 ), .A2(\AES_ENC/us13/n932 ), .ZN(\AES_ENC/us13/n656 ) );
NAND2_X2 \AES_ENC/us13/U445  ( .A1(\AES_ENC/us13/n624 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n1096 ) );
NAND2_X2 \AES_ENC/us13/U444  ( .A1(\AES_ENC/us13/n1030 ), .A2(\AES_ENC/us13/n1096 ), .ZN(\AES_ENC/us13/n651 ) );
NAND2_X2 \AES_ENC/us13/U443  ( .A1(\AES_ENC/us13/n1114 ), .A2(\AES_ENC/us13/n651 ), .ZN(\AES_ENC/us13/n655 ) );
OR3_X2 \AES_ENC/us13/U440  ( .A1(\AES_ENC/us13/n1079 ), .A2(\AES_ENC/sa13 [7]), .A3(\AES_ENC/us13/n594 ), .ZN(\AES_ENC/us13/n654 ));
NAND2_X2 \AES_ENC/us13/U439  ( .A1(\AES_ENC/us13/n623 ), .A2(\AES_ENC/us13/n619 ), .ZN(\AES_ENC/us13/n652 ) );
NAND4_X2 \AES_ENC/us13/U437  ( .A1(\AES_ENC/us13/n656 ), .A2(\AES_ENC/us13/n655 ), .A3(\AES_ENC/us13/n654 ), .A4(\AES_ENC/us13/n653 ), .ZN(\AES_ENC/us13/n657 ) );
NAND2_X2 \AES_ENC/us13/U436  ( .A1(\AES_ENC/sa13 [2]), .A2(\AES_ENC/us13/n657 ), .ZN(\AES_ENC/us13/n660 ) );
NAND4_X2 \AES_ENC/us13/U432  ( .A1(\AES_ENC/us13/n662 ), .A2(\AES_ENC/us13/n661 ), .A3(\AES_ENC/us13/n660 ), .A4(\AES_ENC/us13/n659 ), .ZN(\AES_ENC/us13/n663 ) );
NAND2_X2 \AES_ENC/us13/U431  ( .A1(\AES_ENC/us13/n663 ), .A2(\AES_ENC/us13/n627 ), .ZN(\AES_ENC/us13/n664 ) );
NAND2_X2 \AES_ENC/us13/U430  ( .A1(\AES_ENC/us13/n665 ), .A2(\AES_ENC/us13/n664 ), .ZN(\AES_ENC/us13/n666 ) );
NAND2_X2 \AES_ENC/us13/U429  ( .A1(\AES_ENC/sa13 [6]), .A2(\AES_ENC/us13/n666 ), .ZN(\AES_ENC/us13/n678 ) );
NAND2_X2 \AES_ENC/us13/U426  ( .A1(\AES_ENC/us13/n735 ), .A2(\AES_ENC/us13/n1093 ), .ZN(\AES_ENC/us13/n675 ) );
NAND2_X2 \AES_ENC/us13/U425  ( .A1(\AES_ENC/us13/n625 ), .A2(\AES_ENC/us13/n607 ), .ZN(\AES_ENC/us13/n1045 ) );
OR2_X2 \AES_ENC/us13/U424  ( .A1(\AES_ENC/us13/n1045 ), .A2(\AES_ENC/us13/n577 ), .ZN(\AES_ENC/us13/n674 ) );
NAND2_X2 \AES_ENC/us13/U423  ( .A1(\AES_ENC/sa13 [1]), .A2(\AES_ENC/us13/n609 ), .ZN(\AES_ENC/us13/n667 ) );
NAND2_X2 \AES_ENC/us13/U422  ( .A1(\AES_ENC/us13/n605 ), .A2(\AES_ENC/us13/n667 ), .ZN(\AES_ENC/us13/n1071 ) );
NAND4_X2 \AES_ENC/us13/U412  ( .A1(\AES_ENC/us13/n675 ), .A2(\AES_ENC/us13/n674 ), .A3(\AES_ENC/us13/n673 ), .A4(\AES_ENC/us13/n672 ), .ZN(\AES_ENC/us13/n676 ) );
NAND2_X2 \AES_ENC/us13/U411  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n676 ), .ZN(\AES_ENC/us13/n677 ) );
NAND2_X2 \AES_ENC/us13/U408  ( .A1(\AES_ENC/us13/n800 ), .A2(\AES_ENC/us13/n1022 ), .ZN(\AES_ENC/us13/n680 ) );
NAND2_X2 \AES_ENC/us13/U407  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n680 ), .ZN(\AES_ENC/us13/n681 ) );
AND2_X2 \AES_ENC/us13/U402  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n684 ), .ZN(\AES_ENC/us13/n682 ) );
NAND4_X2 \AES_ENC/us13/U395  ( .A1(\AES_ENC/us13/n691 ), .A2(\AES_ENC/us13/n586 ), .A3(\AES_ENC/us13/n690 ), .A4(\AES_ENC/us13/n689 ), .ZN(\AES_ENC/us13/n692 ) );
NAND2_X2 \AES_ENC/us13/U394  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n692 ), .ZN(\AES_ENC/us13/n733 ) );
NAND2_X2 \AES_ENC/us13/U392  ( .A1(\AES_ENC/us13/n977 ), .A2(\AES_ENC/us13/n1050 ), .ZN(\AES_ENC/us13/n702 ) );
NAND2_X2 \AES_ENC/us13/U391  ( .A1(\AES_ENC/us13/n1093 ), .A2(\AES_ENC/us13/n1045 ), .ZN(\AES_ENC/us13/n701 ) );
NAND4_X2 \AES_ENC/us13/U381  ( .A1(\AES_ENC/us13/n702 ), .A2(\AES_ENC/us13/n701 ), .A3(\AES_ENC/us13/n700 ), .A4(\AES_ENC/us13/n699 ), .ZN(\AES_ENC/us13/n703 ) );
NAND2_X2 \AES_ENC/us13/U380  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n703 ), .ZN(\AES_ENC/us13/n732 ) );
AND2_X2 \AES_ENC/us13/U379  ( .A1(\AES_ENC/sa13 [0]), .A2(\AES_ENC/sa13 [6]),.ZN(\AES_ENC/us13/n1113 ) );
NAND2_X2 \AES_ENC/us13/U378  ( .A1(\AES_ENC/us13/n619 ), .A2(\AES_ENC/us13/n1030 ), .ZN(\AES_ENC/us13/n881 ) );
NAND2_X2 \AES_ENC/us13/U377  ( .A1(\AES_ENC/us13/n1093 ), .A2(\AES_ENC/us13/n881 ), .ZN(\AES_ENC/us13/n715 ) );
NAND2_X2 \AES_ENC/us13/U376  ( .A1(\AES_ENC/us13/n1010 ), .A2(\AES_ENC/us13/n622 ), .ZN(\AES_ENC/us13/n714 ) );
NAND2_X2 \AES_ENC/us13/U375  ( .A1(\AES_ENC/us13/n855 ), .A2(\AES_ENC/us13/n625 ), .ZN(\AES_ENC/us13/n1117 ) );
XNOR2_X2 \AES_ENC/us13/U371  ( .A(\AES_ENC/us13/n584 ), .B(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n824 ) );
NAND4_X2 \AES_ENC/us13/U362  ( .A1(\AES_ENC/us13/n715 ), .A2(\AES_ENC/us13/n714 ), .A3(\AES_ENC/us13/n713 ), .A4(\AES_ENC/us13/n712 ), .ZN(\AES_ENC/us13/n716 ) );
NAND2_X2 \AES_ENC/us13/U361  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n716 ), .ZN(\AES_ENC/us13/n731 ) );
AND2_X2 \AES_ENC/us13/U360  ( .A1(\AES_ENC/sa13 [6]), .A2(\AES_ENC/us13/n627 ), .ZN(\AES_ENC/us13/n1131 ) );
NAND2_X2 \AES_ENC/us13/U359  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n717 ) );
NAND2_X2 \AES_ENC/us13/U358  ( .A1(\AES_ENC/us13/n1029 ), .A2(\AES_ENC/us13/n717 ), .ZN(\AES_ENC/us13/n728 ) );
NAND2_X2 \AES_ENC/us13/U357  ( .A1(\AES_ENC/sa13 [1]), .A2(\AES_ENC/us13/n612 ), .ZN(\AES_ENC/us13/n1097 ) );
NAND2_X2 \AES_ENC/us13/U356  ( .A1(\AES_ENC/us13/n610 ), .A2(\AES_ENC/us13/n1097 ), .ZN(\AES_ENC/us13/n718 ) );
NAND2_X2 \AES_ENC/us13/U355  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n718 ), .ZN(\AES_ENC/us13/n727 ) );
NAND4_X2 \AES_ENC/us13/U344  ( .A1(\AES_ENC/us13/n728 ), .A2(\AES_ENC/us13/n727 ), .A3(\AES_ENC/us13/n726 ), .A4(\AES_ENC/us13/n725 ), .ZN(\AES_ENC/us13/n729 ) );
NAND2_X2 \AES_ENC/us13/U343  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n729 ), .ZN(\AES_ENC/us13/n730 ) );
NAND4_X2 \AES_ENC/us13/U342  ( .A1(\AES_ENC/us13/n733 ), .A2(\AES_ENC/us13/n732 ), .A3(\AES_ENC/us13/n731 ), .A4(\AES_ENC/us13/n730 ), .ZN(\AES_ENC/sa13_sub[1] ) );
NAND2_X2 \AES_ENC/us13/U341  ( .A1(\AES_ENC/sa13 [7]), .A2(\AES_ENC/us13/n584 ), .ZN(\AES_ENC/us13/n734 ) );
NAND2_X2 \AES_ENC/us13/U340  ( .A1(\AES_ENC/us13/n734 ), .A2(\AES_ENC/us13/n579 ), .ZN(\AES_ENC/us13/n738 ) );
OR4_X2 \AES_ENC/us13/U339  ( .A1(\AES_ENC/us13/n738 ), .A2(\AES_ENC/us13/n594 ), .A3(\AES_ENC/us13/n826 ), .A4(\AES_ENC/us13/n1121 ), .ZN(\AES_ENC/us13/n746 ) );
NAND2_X2 \AES_ENC/us13/U337  ( .A1(\AES_ENC/us13/n1100 ), .A2(\AES_ENC/us13/n617 ), .ZN(\AES_ENC/us13/n992 ) );
OR2_X2 \AES_ENC/us13/U336  ( .A1(\AES_ENC/us13/n583 ), .A2(\AES_ENC/us13/n735 ), .ZN(\AES_ENC/us13/n737 ) );
NAND2_X2 \AES_ENC/us13/U334  ( .A1(\AES_ENC/us13/n605 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n753 ) );
NAND2_X2 \AES_ENC/us13/U333  ( .A1(\AES_ENC/us13/n603 ), .A2(\AES_ENC/us13/n753 ), .ZN(\AES_ENC/us13/n1080 ) );
NAND2_X2 \AES_ENC/us13/U332  ( .A1(\AES_ENC/us13/n1048 ), .A2(\AES_ENC/us13/n602 ), .ZN(\AES_ENC/us13/n736 ) );
NAND2_X2 \AES_ENC/us13/U331  ( .A1(\AES_ENC/us13/n737 ), .A2(\AES_ENC/us13/n736 ), .ZN(\AES_ENC/us13/n739 ) );
NAND2_X2 \AES_ENC/us13/U330  ( .A1(\AES_ENC/us13/n739 ), .A2(\AES_ENC/us13/n738 ), .ZN(\AES_ENC/us13/n745 ) );
NAND2_X2 \AES_ENC/us13/U326  ( .A1(\AES_ENC/us13/n1096 ), .A2(\AES_ENC/us13/n598 ), .ZN(\AES_ENC/us13/n906 ) );
NAND4_X2 \AES_ENC/us13/U323  ( .A1(\AES_ENC/us13/n746 ), .A2(\AES_ENC/us13/n992 ), .A3(\AES_ENC/us13/n745 ), .A4(\AES_ENC/us13/n744 ), .ZN(\AES_ENC/us13/n747 ) );
NAND2_X2 \AES_ENC/us13/U322  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n747 ), .ZN(\AES_ENC/us13/n793 ) );
NAND2_X2 \AES_ENC/us13/U321  ( .A1(\AES_ENC/us13/n606 ), .A2(\AES_ENC/us13/n855 ), .ZN(\AES_ENC/us13/n748 ) );
NAND2_X2 \AES_ENC/us13/U320  ( .A1(\AES_ENC/us13/n956 ), .A2(\AES_ENC/us13/n748 ), .ZN(\AES_ENC/us13/n760 ) );
NAND2_X2 \AES_ENC/us13/U313  ( .A1(\AES_ENC/us13/n598 ), .A2(\AES_ENC/us13/n753 ), .ZN(\AES_ENC/us13/n1023 ) );
NAND4_X2 \AES_ENC/us13/U308  ( .A1(\AES_ENC/us13/n760 ), .A2(\AES_ENC/us13/n992 ), .A3(\AES_ENC/us13/n759 ), .A4(\AES_ENC/us13/n758 ), .ZN(\AES_ENC/us13/n761 ) );
NAND2_X2 \AES_ENC/us13/U307  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n761 ), .ZN(\AES_ENC/us13/n792 ) );
NAND2_X2 \AES_ENC/us13/U306  ( .A1(\AES_ENC/us13/n606 ), .A2(\AES_ENC/us13/n610 ), .ZN(\AES_ENC/us13/n989 ) );
NAND2_X2 \AES_ENC/us13/U305  ( .A1(\AES_ENC/us13/n1050 ), .A2(\AES_ENC/us13/n989 ), .ZN(\AES_ENC/us13/n777 ) );
NAND2_X2 \AES_ENC/us13/U304  ( .A1(\AES_ENC/us13/n1093 ), .A2(\AES_ENC/us13/n762 ), .ZN(\AES_ENC/us13/n776 ) );
XNOR2_X2 \AES_ENC/us13/U301  ( .A(\AES_ENC/sa13 [7]), .B(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n959 ) );
NAND4_X2 \AES_ENC/us13/U289  ( .A1(\AES_ENC/us13/n777 ), .A2(\AES_ENC/us13/n776 ), .A3(\AES_ENC/us13/n775 ), .A4(\AES_ENC/us13/n774 ), .ZN(\AES_ENC/us13/n778 ) );
NAND2_X2 \AES_ENC/us13/U288  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n778 ), .ZN(\AES_ENC/us13/n791 ) );
NAND2_X2 \AES_ENC/us13/U287  ( .A1(\AES_ENC/us13/n1056 ), .A2(\AES_ENC/us13/n1050 ), .ZN(\AES_ENC/us13/n788 ) );
NAND2_X2 \AES_ENC/us13/U286  ( .A1(\AES_ENC/us13/n1091 ), .A2(\AES_ENC/us13/n779 ), .ZN(\AES_ENC/us13/n787 ) );
NAND2_X2 \AES_ENC/us13/U285  ( .A1(\AES_ENC/us13/n956 ), .A2(\AES_ENC/sa13 [1]), .ZN(\AES_ENC/us13/n786 ) );
NAND4_X2 \AES_ENC/us13/U278  ( .A1(\AES_ENC/us13/n788 ), .A2(\AES_ENC/us13/n787 ), .A3(\AES_ENC/us13/n786 ), .A4(\AES_ENC/us13/n785 ), .ZN(\AES_ENC/us13/n789 ) );
NAND2_X2 \AES_ENC/us13/U277  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n789 ), .ZN(\AES_ENC/us13/n790 ) );
NAND4_X2 \AES_ENC/us13/U276  ( .A1(\AES_ENC/us13/n793 ), .A2(\AES_ENC/us13/n792 ), .A3(\AES_ENC/us13/n791 ), .A4(\AES_ENC/us13/n790 ), .ZN(\AES_ENC/sa13_sub[2] ) );
NAND2_X2 \AES_ENC/us13/U275  ( .A1(\AES_ENC/us13/n1059 ), .A2(\AES_ENC/us13/n794 ), .ZN(\AES_ENC/us13/n810 ) );
NAND2_X2 \AES_ENC/us13/U274  ( .A1(\AES_ENC/us13/n1049 ), .A2(\AES_ENC/us13/n956 ), .ZN(\AES_ENC/us13/n809 ) );
OR2_X2 \AES_ENC/us13/U266  ( .A1(\AES_ENC/us13/n1096 ), .A2(\AES_ENC/us13/n578 ), .ZN(\AES_ENC/us13/n802 ) );
NAND2_X2 \AES_ENC/us13/U265  ( .A1(\AES_ENC/us13/n1053 ), .A2(\AES_ENC/us13/n800 ), .ZN(\AES_ENC/us13/n801 ) );
NAND2_X2 \AES_ENC/us13/U264  ( .A1(\AES_ENC/us13/n802 ), .A2(\AES_ENC/us13/n801 ), .ZN(\AES_ENC/us13/n805 ) );
NAND4_X2 \AES_ENC/us13/U261  ( .A1(\AES_ENC/us13/n810 ), .A2(\AES_ENC/us13/n809 ), .A3(\AES_ENC/us13/n808 ), .A4(\AES_ENC/us13/n807 ), .ZN(\AES_ENC/us13/n811 ) );
NAND2_X2 \AES_ENC/us13/U260  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n811 ), .ZN(\AES_ENC/us13/n852 ) );
OR2_X2 \AES_ENC/us13/U259  ( .A1(\AES_ENC/us13/n1023 ), .A2(\AES_ENC/us13/n591 ), .ZN(\AES_ENC/us13/n819 ) );
OR2_X2 \AES_ENC/us13/U257  ( .A1(\AES_ENC/us13/n570 ), .A2(\AES_ENC/us13/n930 ), .ZN(\AES_ENC/us13/n818 ) );
NAND2_X2 \AES_ENC/us13/U256  ( .A1(\AES_ENC/us13/n1013 ), .A2(\AES_ENC/us13/n1094 ), .ZN(\AES_ENC/us13/n817 ) );
NAND4_X2 \AES_ENC/us13/U249  ( .A1(\AES_ENC/us13/n819 ), .A2(\AES_ENC/us13/n818 ), .A3(\AES_ENC/us13/n817 ), .A4(\AES_ENC/us13/n816 ), .ZN(\AES_ENC/us13/n820 ) );
NAND2_X2 \AES_ENC/us13/U248  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n820 ), .ZN(\AES_ENC/us13/n851 ) );
NAND2_X2 \AES_ENC/us13/U247  ( .A1(\AES_ENC/us13/n956 ), .A2(\AES_ENC/us13/n1080 ), .ZN(\AES_ENC/us13/n835 ) );
NAND2_X2 \AES_ENC/us13/U246  ( .A1(\AES_ENC/us13/n570 ), .A2(\AES_ENC/us13/n1030 ), .ZN(\AES_ENC/us13/n1047 ) );
OR2_X2 \AES_ENC/us13/U245  ( .A1(\AES_ENC/us13/n1047 ), .A2(\AES_ENC/us13/n585 ), .ZN(\AES_ENC/us13/n834 ) );
NAND2_X2 \AES_ENC/us13/U244  ( .A1(\AES_ENC/us13/n1072 ), .A2(\AES_ENC/us13/n620 ), .ZN(\AES_ENC/us13/n833 ) );
NAND4_X2 \AES_ENC/us13/U233  ( .A1(\AES_ENC/us13/n835 ), .A2(\AES_ENC/us13/n834 ), .A3(\AES_ENC/us13/n833 ), .A4(\AES_ENC/us13/n832 ), .ZN(\AES_ENC/us13/n836 ) );
NAND2_X2 \AES_ENC/us13/U232  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n836 ), .ZN(\AES_ENC/us13/n850 ) );
NAND2_X2 \AES_ENC/us13/U231  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n601 ), .ZN(\AES_ENC/us13/n847 ) );
NAND2_X2 \AES_ENC/us13/U230  ( .A1(\AES_ENC/us13/n1050 ), .A2(\AES_ENC/us13/n1071 ), .ZN(\AES_ENC/us13/n846 ) );
OR2_X2 \AES_ENC/us13/U224  ( .A1(\AES_ENC/us13/n1053 ), .A2(\AES_ENC/us13/n911 ), .ZN(\AES_ENC/us13/n1077 ) );
NAND4_X2 \AES_ENC/us13/U220  ( .A1(\AES_ENC/us13/n847 ), .A2(\AES_ENC/us13/n846 ), .A3(\AES_ENC/us13/n845 ), .A4(\AES_ENC/us13/n844 ), .ZN(\AES_ENC/us13/n848 ) );
NAND2_X2 \AES_ENC/us13/U219  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n848 ), .ZN(\AES_ENC/us13/n849 ) );
NAND4_X2 \AES_ENC/us13/U218  ( .A1(\AES_ENC/us13/n852 ), .A2(\AES_ENC/us13/n851 ), .A3(\AES_ENC/us13/n850 ), .A4(\AES_ENC/us13/n849 ), .ZN(\AES_ENC/sa13_sub[3] ) );
NAND2_X2 \AES_ENC/us13/U216  ( .A1(\AES_ENC/us13/n1009 ), .A2(\AES_ENC/us13/n1072 ), .ZN(\AES_ENC/us13/n862 ) );
NAND2_X2 \AES_ENC/us13/U215  ( .A1(\AES_ENC/us13/n610 ), .A2(\AES_ENC/us13/n618 ), .ZN(\AES_ENC/us13/n853 ) );
NAND2_X2 \AES_ENC/us13/U214  ( .A1(\AES_ENC/us13/n1050 ), .A2(\AES_ENC/us13/n853 ), .ZN(\AES_ENC/us13/n861 ) );
NAND4_X2 \AES_ENC/us13/U206  ( .A1(\AES_ENC/us13/n862 ), .A2(\AES_ENC/us13/n861 ), .A3(\AES_ENC/us13/n860 ), .A4(\AES_ENC/us13/n859 ), .ZN(\AES_ENC/us13/n863 ) );
NAND2_X2 \AES_ENC/us13/U205  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n863 ), .ZN(\AES_ENC/us13/n905 ) );
NAND2_X2 \AES_ENC/us13/U204  ( .A1(\AES_ENC/us13/n1010 ), .A2(\AES_ENC/us13/n989 ), .ZN(\AES_ENC/us13/n874 ) );
NAND2_X2 \AES_ENC/us13/U203  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n583 ), .ZN(\AES_ENC/us13/n864 ) );
NAND2_X2 \AES_ENC/us13/U202  ( .A1(\AES_ENC/us13/n929 ), .A2(\AES_ENC/us13/n864 ), .ZN(\AES_ENC/us13/n873 ) );
NAND4_X2 \AES_ENC/us13/U193  ( .A1(\AES_ENC/us13/n874 ), .A2(\AES_ENC/us13/n873 ), .A3(\AES_ENC/us13/n872 ), .A4(\AES_ENC/us13/n871 ), .ZN(\AES_ENC/us13/n875 ) );
NAND2_X2 \AES_ENC/us13/U192  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n875 ), .ZN(\AES_ENC/us13/n904 ) );
NAND2_X2 \AES_ENC/us13/U191  ( .A1(\AES_ENC/us13/n597 ), .A2(\AES_ENC/us13/n1050 ), .ZN(\AES_ENC/us13/n889 ) );
NAND2_X2 \AES_ENC/us13/U190  ( .A1(\AES_ENC/us13/n1093 ), .A2(\AES_ENC/us13/n617 ), .ZN(\AES_ENC/us13/n876 ) );
NAND2_X2 \AES_ENC/us13/U189  ( .A1(\AES_ENC/us13/n576 ), .A2(\AES_ENC/us13/n876 ), .ZN(\AES_ENC/us13/n877 ) );
NAND2_X2 \AES_ENC/us13/U188  ( .A1(\AES_ENC/us13/n877 ), .A2(\AES_ENC/us13/n601 ), .ZN(\AES_ENC/us13/n888 ) );
NAND4_X2 \AES_ENC/us13/U179  ( .A1(\AES_ENC/us13/n889 ), .A2(\AES_ENC/us13/n888 ), .A3(\AES_ENC/us13/n887 ), .A4(\AES_ENC/us13/n886 ), .ZN(\AES_ENC/us13/n890 ) );
NAND2_X2 \AES_ENC/us13/U178  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n890 ), .ZN(\AES_ENC/us13/n903 ) );
OR2_X2 \AES_ENC/us13/U177  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n1059 ), .ZN(\AES_ENC/us13/n900 ) );
NAND2_X2 \AES_ENC/us13/U176  ( .A1(\AES_ENC/us13/n1073 ), .A2(\AES_ENC/us13/n1047 ), .ZN(\AES_ENC/us13/n899 ) );
NAND2_X2 \AES_ENC/us13/U175  ( .A1(\AES_ENC/us13/n1094 ), .A2(\AES_ENC/us13/n608 ), .ZN(\AES_ENC/us13/n898 ) );
NAND4_X2 \AES_ENC/us13/U167  ( .A1(\AES_ENC/us13/n900 ), .A2(\AES_ENC/us13/n899 ), .A3(\AES_ENC/us13/n898 ), .A4(\AES_ENC/us13/n897 ), .ZN(\AES_ENC/us13/n901 ) );
NAND2_X2 \AES_ENC/us13/U166  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n901 ), .ZN(\AES_ENC/us13/n902 ) );
NAND4_X2 \AES_ENC/us13/U165  ( .A1(\AES_ENC/us13/n905 ), .A2(\AES_ENC/us13/n904 ), .A3(\AES_ENC/us13/n903 ), .A4(\AES_ENC/us13/n902 ), .ZN(\AES_ENC/sa13_sub[4] ) );
NAND2_X2 \AES_ENC/us13/U164  ( .A1(\AES_ENC/us13/n1094 ), .A2(\AES_ENC/us13/n615 ), .ZN(\AES_ENC/us13/n922 ) );
NAND2_X2 \AES_ENC/us13/U163  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n989 ), .ZN(\AES_ENC/us13/n921 ) );
NAND4_X2 \AES_ENC/us13/U151  ( .A1(\AES_ENC/us13/n922 ), .A2(\AES_ENC/us13/n921 ), .A3(\AES_ENC/us13/n920 ), .A4(\AES_ENC/us13/n919 ), .ZN(\AES_ENC/us13/n923 ) );
NAND2_X2 \AES_ENC/us13/U150  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n923 ), .ZN(\AES_ENC/us13/n972 ) );
NAND2_X2 \AES_ENC/us13/U149  ( .A1(\AES_ENC/us13/n603 ), .A2(\AES_ENC/us13/n605 ), .ZN(\AES_ENC/us13/n924 ) );
NAND2_X2 \AES_ENC/us13/U148  ( .A1(\AES_ENC/us13/n1073 ), .A2(\AES_ENC/us13/n924 ), .ZN(\AES_ENC/us13/n939 ) );
NAND2_X2 \AES_ENC/us13/U147  ( .A1(\AES_ENC/us13/n926 ), .A2(\AES_ENC/us13/n925 ), .ZN(\AES_ENC/us13/n927 ) );
NAND2_X2 \AES_ENC/us13/U146  ( .A1(\AES_ENC/us13/n578 ), .A2(\AES_ENC/us13/n927 ), .ZN(\AES_ENC/us13/n928 ) );
NAND2_X2 \AES_ENC/us13/U145  ( .A1(\AES_ENC/us13/n928 ), .A2(\AES_ENC/us13/n1080 ), .ZN(\AES_ENC/us13/n938 ) );
OR2_X2 \AES_ENC/us13/U144  ( .A1(\AES_ENC/us13/n1117 ), .A2(\AES_ENC/us13/n589 ), .ZN(\AES_ENC/us13/n937 ) );
NAND4_X2 \AES_ENC/us13/U139  ( .A1(\AES_ENC/us13/n939 ), .A2(\AES_ENC/us13/n938 ), .A3(\AES_ENC/us13/n937 ), .A4(\AES_ENC/us13/n936 ), .ZN(\AES_ENC/us13/n940 ) );
NAND2_X2 \AES_ENC/us13/U138  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n940 ), .ZN(\AES_ENC/us13/n971 ) );
OR2_X2 \AES_ENC/us13/U137  ( .A1(\AES_ENC/us13/n577 ), .A2(\AES_ENC/us13/n941 ), .ZN(\AES_ENC/us13/n954 ) );
NAND2_X2 \AES_ENC/us13/U136  ( .A1(\AES_ENC/us13/n1096 ), .A2(\AES_ENC/us13/n618 ), .ZN(\AES_ENC/us13/n942 ) );
NAND2_X2 \AES_ENC/us13/U135  ( .A1(\AES_ENC/us13/n1048 ), .A2(\AES_ENC/us13/n942 ), .ZN(\AES_ENC/us13/n943 ) );
NAND2_X2 \AES_ENC/us13/U134  ( .A1(\AES_ENC/us13/n585 ), .A2(\AES_ENC/us13/n943 ), .ZN(\AES_ENC/us13/n944 ) );
NAND2_X2 \AES_ENC/us13/U133  ( .A1(\AES_ENC/us13/n944 ), .A2(\AES_ENC/us13/n599 ), .ZN(\AES_ENC/us13/n953 ) );
NAND4_X2 \AES_ENC/us13/U125  ( .A1(\AES_ENC/us13/n954 ), .A2(\AES_ENC/us13/n953 ), .A3(\AES_ENC/us13/n952 ), .A4(\AES_ENC/us13/n951 ), .ZN(\AES_ENC/us13/n955 ) );
NAND2_X2 \AES_ENC/us13/U124  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n955 ), .ZN(\AES_ENC/us13/n970 ) );
NAND2_X2 \AES_ENC/us13/U123  ( .A1(\AES_ENC/us13/n1094 ), .A2(\AES_ENC/us13/n1071 ), .ZN(\AES_ENC/us13/n967 ) );
NAND2_X2 \AES_ENC/us13/U122  ( .A1(\AES_ENC/us13/n956 ), .A2(\AES_ENC/us13/n1030 ), .ZN(\AES_ENC/us13/n966 ) );
NAND4_X2 \AES_ENC/us13/U114  ( .A1(\AES_ENC/us13/n967 ), .A2(\AES_ENC/us13/n966 ), .A3(\AES_ENC/us13/n965 ), .A4(\AES_ENC/us13/n964 ), .ZN(\AES_ENC/us13/n968 ) );
NAND2_X2 \AES_ENC/us13/U113  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n968 ), .ZN(\AES_ENC/us13/n969 ) );
NAND4_X2 \AES_ENC/us13/U112  ( .A1(\AES_ENC/us13/n972 ), .A2(\AES_ENC/us13/n971 ), .A3(\AES_ENC/us13/n970 ), .A4(\AES_ENC/us13/n969 ), .ZN(\AES_ENC/sa13_sub[5] ) );
NAND2_X2 \AES_ENC/us13/U111  ( .A1(\AES_ENC/us13/n570 ), .A2(\AES_ENC/us13/n1097 ), .ZN(\AES_ENC/us13/n973 ) );
NAND2_X2 \AES_ENC/us13/U110  ( .A1(\AES_ENC/us13/n1073 ), .A2(\AES_ENC/us13/n973 ), .ZN(\AES_ENC/us13/n987 ) );
NAND2_X2 \AES_ENC/us13/U109  ( .A1(\AES_ENC/us13/n974 ), .A2(\AES_ENC/us13/n1077 ), .ZN(\AES_ENC/us13/n975 ) );
NAND2_X2 \AES_ENC/us13/U108  ( .A1(\AES_ENC/us13/n587 ), .A2(\AES_ENC/us13/n975 ), .ZN(\AES_ENC/us13/n976 ) );
NAND2_X2 \AES_ENC/us13/U107  ( .A1(\AES_ENC/us13/n977 ), .A2(\AES_ENC/us13/n976 ), .ZN(\AES_ENC/us13/n986 ) );
NAND4_X2 \AES_ENC/us13/U99  ( .A1(\AES_ENC/us13/n987 ), .A2(\AES_ENC/us13/n986 ), .A3(\AES_ENC/us13/n985 ), .A4(\AES_ENC/us13/n984 ), .ZN(\AES_ENC/us13/n988 ) );
NAND2_X2 \AES_ENC/us13/U98  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n988 ), .ZN(\AES_ENC/us13/n1044 ) );
NAND2_X2 \AES_ENC/us13/U97  ( .A1(\AES_ENC/us13/n1073 ), .A2(\AES_ENC/us13/n989 ), .ZN(\AES_ENC/us13/n1004 ) );
NAND2_X2 \AES_ENC/us13/U96  ( .A1(\AES_ENC/us13/n1092 ), .A2(\AES_ENC/us13/n605 ), .ZN(\AES_ENC/us13/n1003 ) );
NAND4_X2 \AES_ENC/us13/U85  ( .A1(\AES_ENC/us13/n1004 ), .A2(\AES_ENC/us13/n1003 ), .A3(\AES_ENC/us13/n1002 ), .A4(\AES_ENC/us13/n1001 ), .ZN(\AES_ENC/us13/n1005 ) );
NAND2_X2 \AES_ENC/us13/U84  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n1005 ), .ZN(\AES_ENC/us13/n1043 ) );
NAND2_X2 \AES_ENC/us13/U83  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n626 ), .ZN(\AES_ENC/us13/n1020 ) );
NAND2_X2 \AES_ENC/us13/U82  ( .A1(\AES_ENC/us13/n1050 ), .A2(\AES_ENC/us13/n612 ), .ZN(\AES_ENC/us13/n1019 ) );
NAND2_X2 \AES_ENC/us13/U77  ( .A1(\AES_ENC/us13/n1059 ), .A2(\AES_ENC/us13/n1114 ), .ZN(\AES_ENC/us13/n1012 ) );
NAND2_X2 \AES_ENC/us13/U76  ( .A1(\AES_ENC/us13/n1010 ), .A2(\AES_ENC/us13/n604 ), .ZN(\AES_ENC/us13/n1011 ) );
NAND2_X2 \AES_ENC/us13/U75  ( .A1(\AES_ENC/us13/n1012 ), .A2(\AES_ENC/us13/n1011 ), .ZN(\AES_ENC/us13/n1016 ) );
NAND4_X2 \AES_ENC/us13/U70  ( .A1(\AES_ENC/us13/n1020 ), .A2(\AES_ENC/us13/n1019 ), .A3(\AES_ENC/us13/n1018 ), .A4(\AES_ENC/us13/n1017 ), .ZN(\AES_ENC/us13/n1021 ) );
NAND2_X2 \AES_ENC/us13/U69  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n1021 ), .ZN(\AES_ENC/us13/n1042 ) );
NAND2_X2 \AES_ENC/us13/U68  ( .A1(\AES_ENC/us13/n1022 ), .A2(\AES_ENC/us13/n1093 ), .ZN(\AES_ENC/us13/n1039 ) );
NAND2_X2 \AES_ENC/us13/U67  ( .A1(\AES_ENC/us13/n1050 ), .A2(\AES_ENC/us13/n1023 ), .ZN(\AES_ENC/us13/n1038 ) );
NAND2_X2 \AES_ENC/us13/U66  ( .A1(\AES_ENC/us13/n1024 ), .A2(\AES_ENC/us13/n1071 ), .ZN(\AES_ENC/us13/n1037 ) );
AND2_X2 \AES_ENC/us13/U60  ( .A1(\AES_ENC/us13/n1030 ), .A2(\AES_ENC/us13/n621 ), .ZN(\AES_ENC/us13/n1078 ) );
NAND4_X2 \AES_ENC/us13/U56  ( .A1(\AES_ENC/us13/n1039 ), .A2(\AES_ENC/us13/n1038 ), .A3(\AES_ENC/us13/n1037 ), .A4(\AES_ENC/us13/n1036 ), .ZN(\AES_ENC/us13/n1040 ) );
NAND2_X2 \AES_ENC/us13/U55  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n1040 ), .ZN(\AES_ENC/us13/n1041 ) );
NAND4_X2 \AES_ENC/us13/U54  ( .A1(\AES_ENC/us13/n1044 ), .A2(\AES_ENC/us13/n1043 ), .A3(\AES_ENC/us13/n1042 ), .A4(\AES_ENC/us13/n1041 ), .ZN(\AES_ENC/sa13_sub[6] ) );
NAND2_X2 \AES_ENC/us13/U53  ( .A1(\AES_ENC/us13/n1072 ), .A2(\AES_ENC/us13/n1045 ), .ZN(\AES_ENC/us13/n1068 ) );
NAND2_X2 \AES_ENC/us13/U52  ( .A1(\AES_ENC/us13/n1046 ), .A2(\AES_ENC/us13/n603 ), .ZN(\AES_ENC/us13/n1067 ) );
NAND2_X2 \AES_ENC/us13/U51  ( .A1(\AES_ENC/us13/n1094 ), .A2(\AES_ENC/us13/n1047 ), .ZN(\AES_ENC/us13/n1066 ) );
NAND4_X2 \AES_ENC/us13/U40  ( .A1(\AES_ENC/us13/n1068 ), .A2(\AES_ENC/us13/n1067 ), .A3(\AES_ENC/us13/n1066 ), .A4(\AES_ENC/us13/n1065 ), .ZN(\AES_ENC/us13/n1069 ) );
NAND2_X2 \AES_ENC/us13/U39  ( .A1(\AES_ENC/us13/n1070 ), .A2(\AES_ENC/us13/n1069 ), .ZN(\AES_ENC/us13/n1135 ) );
NAND2_X2 \AES_ENC/us13/U38  ( .A1(\AES_ENC/us13/n1072 ), .A2(\AES_ENC/us13/n1071 ), .ZN(\AES_ENC/us13/n1088 ) );
NAND2_X2 \AES_ENC/us13/U37  ( .A1(\AES_ENC/us13/n1073 ), .A2(\AES_ENC/us13/n608 ), .ZN(\AES_ENC/us13/n1087 ) );
NAND4_X2 \AES_ENC/us13/U28  ( .A1(\AES_ENC/us13/n1088 ), .A2(\AES_ENC/us13/n1087 ), .A3(\AES_ENC/us13/n1086 ), .A4(\AES_ENC/us13/n1085 ), .ZN(\AES_ENC/us13/n1089 ) );
NAND2_X2 \AES_ENC/us13/U27  ( .A1(\AES_ENC/us13/n1090 ), .A2(\AES_ENC/us13/n1089 ), .ZN(\AES_ENC/us13/n1134 ) );
NAND2_X2 \AES_ENC/us13/U26  ( .A1(\AES_ENC/us13/n1091 ), .A2(\AES_ENC/us13/n1093 ), .ZN(\AES_ENC/us13/n1111 ) );
NAND2_X2 \AES_ENC/us13/U25  ( .A1(\AES_ENC/us13/n1092 ), .A2(\AES_ENC/us13/n1120 ), .ZN(\AES_ENC/us13/n1110 ) );
AND2_X2 \AES_ENC/us13/U22  ( .A1(\AES_ENC/us13/n1097 ), .A2(\AES_ENC/us13/n1096 ), .ZN(\AES_ENC/us13/n1098 ) );
NAND4_X2 \AES_ENC/us13/U14  ( .A1(\AES_ENC/us13/n1111 ), .A2(\AES_ENC/us13/n1110 ), .A3(\AES_ENC/us13/n1109 ), .A4(\AES_ENC/us13/n1108 ), .ZN(\AES_ENC/us13/n1112 ) );
NAND2_X2 \AES_ENC/us13/U13  ( .A1(\AES_ENC/us13/n1113 ), .A2(\AES_ENC/us13/n1112 ), .ZN(\AES_ENC/us13/n1133 ) );
NAND2_X2 \AES_ENC/us13/U12  ( .A1(\AES_ENC/us13/n1115 ), .A2(\AES_ENC/us13/n1114 ), .ZN(\AES_ENC/us13/n1129 ) );
OR2_X2 \AES_ENC/us13/U11  ( .A1(\AES_ENC/us13/n581 ), .A2(\AES_ENC/us13/n1116 ), .ZN(\AES_ENC/us13/n1128 ) );
NAND4_X2 \AES_ENC/us13/U3  ( .A1(\AES_ENC/us13/n1129 ), .A2(\AES_ENC/us13/n1128 ), .A3(\AES_ENC/us13/n1127 ), .A4(\AES_ENC/us13/n1126 ), .ZN(\AES_ENC/us13/n1130 ) );
NAND2_X2 \AES_ENC/us13/U2  ( .A1(\AES_ENC/us13/n1131 ), .A2(\AES_ENC/us13/n1130 ), .ZN(\AES_ENC/us13/n1132 ) );
NAND4_X2 \AES_ENC/us13/U1  ( .A1(\AES_ENC/us13/n1135 ), .A2(\AES_ENC/us13/n1134 ), .A3(\AES_ENC/us13/n1133 ), .A4(\AES_ENC/us13/n1132 ), .ZN(\AES_ENC/sa13_sub[7] ) );
INV_X4 \AES_ENC/us20/U575  ( .A(\AES_ENC/sa20 [0]), .ZN(\AES_ENC/us20/n627 ));
INV_X4 \AES_ENC/us20/U574  ( .A(\AES_ENC/us20/n1053 ), .ZN(\AES_ENC/us20/n625 ) );
INV_X4 \AES_ENC/us20/U573  ( .A(\AES_ENC/us20/n1103 ), .ZN(\AES_ENC/us20/n623 ) );
INV_X4 \AES_ENC/us20/U572  ( .A(\AES_ENC/us20/n1056 ), .ZN(\AES_ENC/us20/n622 ) );
INV_X4 \AES_ENC/us20/U571  ( .A(\AES_ENC/us20/n1102 ), .ZN(\AES_ENC/us20/n621 ) );
INV_X4 \AES_ENC/us20/U570  ( .A(\AES_ENC/us20/n1074 ), .ZN(\AES_ENC/us20/n620 ) );
INV_X4 \AES_ENC/us20/U569  ( .A(\AES_ENC/us20/n929 ), .ZN(\AES_ENC/us20/n619 ) );
INV_X4 \AES_ENC/us20/U568  ( .A(\AES_ENC/us20/n1091 ), .ZN(\AES_ENC/us20/n618 ) );
INV_X4 \AES_ENC/us20/U567  ( .A(\AES_ENC/us20/n826 ), .ZN(\AES_ENC/us20/n617 ) );
INV_X4 \AES_ENC/us20/U566  ( .A(\AES_ENC/us20/n1031 ), .ZN(\AES_ENC/us20/n616 ) );
INV_X4 \AES_ENC/us20/U565  ( .A(\AES_ENC/us20/n1054 ), .ZN(\AES_ENC/us20/n615 ) );
INV_X4 \AES_ENC/us20/U564  ( .A(\AES_ENC/us20/n1025 ), .ZN(\AES_ENC/us20/n614 ) );
INV_X4 \AES_ENC/us20/U563  ( .A(\AES_ENC/us20/n990 ), .ZN(\AES_ENC/us20/n613 ) );
INV_X4 \AES_ENC/us20/U562  ( .A(\AES_ENC/sa20 [4]), .ZN(\AES_ENC/us20/n612 ));
INV_X4 \AES_ENC/us20/U561  ( .A(\AES_ENC/us20/n881 ), .ZN(\AES_ENC/us20/n611 ) );
INV_X4 \AES_ENC/us20/U560  ( .A(\AES_ENC/us20/n1022 ), .ZN(\AES_ENC/us20/n610 ) );
INV_X4 \AES_ENC/us20/U559  ( .A(\AES_ENC/us20/n1120 ), .ZN(\AES_ENC/us20/n609 ) );
INV_X4 \AES_ENC/us20/U558  ( .A(\AES_ENC/us20/n977 ), .ZN(\AES_ENC/us20/n608 ) );
INV_X4 \AES_ENC/us20/U557  ( .A(\AES_ENC/us20/n926 ), .ZN(\AES_ENC/us20/n607 ) );
INV_X4 \AES_ENC/us20/U556  ( .A(\AES_ENC/us20/n910 ), .ZN(\AES_ENC/us20/n606 ) );
INV_X4 \AES_ENC/us20/U555  ( .A(\AES_ENC/us20/n1121 ), .ZN(\AES_ENC/us20/n605 ) );
INV_X4 \AES_ENC/us20/U554  ( .A(\AES_ENC/us20/n1009 ), .ZN(\AES_ENC/us20/n604 ) );
INV_X4 \AES_ENC/us20/U553  ( .A(\AES_ENC/us20/n1080 ), .ZN(\AES_ENC/us20/n602 ) );
INV_X4 \AES_ENC/us20/U552  ( .A(\AES_ENC/us20/n821 ), .ZN(\AES_ENC/us20/n600 ) );
INV_X4 \AES_ENC/us20/U551  ( .A(\AES_ENC/us20/n1013 ), .ZN(\AES_ENC/us20/n599 ) );
INV_X4 \AES_ENC/us20/U550  ( .A(\AES_ENC/us20/n1058 ), .ZN(\AES_ENC/us20/n598 ) );
INV_X4 \AES_ENC/us20/U549  ( .A(\AES_ENC/us20/n906 ), .ZN(\AES_ENC/us20/n597 ) );
INV_X4 \AES_ENC/us20/U548  ( .A(\AES_ENC/us20/n1048 ), .ZN(\AES_ENC/us20/n595 ) );
INV_X4 \AES_ENC/us20/U547  ( .A(\AES_ENC/us20/n974 ), .ZN(\AES_ENC/us20/n594 ) );
INV_X4 \AES_ENC/us20/U546  ( .A(\AES_ENC/sa20 [2]), .ZN(\AES_ENC/us20/n593 ));
INV_X4 \AES_ENC/us20/U545  ( .A(\AES_ENC/us20/n800 ), .ZN(\AES_ENC/us20/n592 ) );
INV_X4 \AES_ENC/us20/U544  ( .A(\AES_ENC/us20/n925 ), .ZN(\AES_ENC/us20/n591 ) );
INV_X4 \AES_ENC/us20/U543  ( .A(\AES_ENC/us20/n824 ), .ZN(\AES_ENC/us20/n590 ) );
INV_X4 \AES_ENC/us20/U542  ( .A(\AES_ENC/us20/n959 ), .ZN(\AES_ENC/us20/n589 ) );
INV_X4 \AES_ENC/us20/U541  ( .A(\AES_ENC/us20/n779 ), .ZN(\AES_ENC/us20/n588 ) );
INV_X4 \AES_ENC/us20/U540  ( .A(\AES_ENC/us20/n794 ), .ZN(\AES_ENC/us20/n585 ) );
INV_X4 \AES_ENC/us20/U539  ( .A(\AES_ENC/us20/n880 ), .ZN(\AES_ENC/us20/n583 ) );
INV_X4 \AES_ENC/us20/U538  ( .A(\AES_ENC/sa20 [7]), .ZN(\AES_ENC/us20/n581 ));
INV_X4 \AES_ENC/us20/U537  ( .A(\AES_ENC/us20/n992 ), .ZN(\AES_ENC/us20/n578 ) );
INV_X4 \AES_ENC/us20/U536  ( .A(\AES_ENC/us20/n1114 ), .ZN(\AES_ENC/us20/n577 ) );
INV_X4 \AES_ENC/us20/U535  ( .A(\AES_ENC/us20/n1092 ), .ZN(\AES_ENC/us20/n574 ) );
NOR2_X2 \AES_ENC/us20/U534  ( .A1(\AES_ENC/sa20 [0]), .A2(\AES_ENC/sa20 [6]),.ZN(\AES_ENC/us20/n1090 ) );
NOR2_X2 \AES_ENC/us20/U533  ( .A1(\AES_ENC/us20/n627 ), .A2(\AES_ENC/sa20 [6]), .ZN(\AES_ENC/us20/n1070 ) );
NOR2_X2 \AES_ENC/us20/U532  ( .A1(\AES_ENC/sa20 [4]), .A2(\AES_ENC/sa20 [3]),.ZN(\AES_ENC/us20/n1025 ) );
INV_X4 \AES_ENC/us20/U531  ( .A(\AES_ENC/us20/n569 ), .ZN(\AES_ENC/us20/n572 ) );
NOR2_X2 \AES_ENC/us20/U530  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n765 ) );
NOR2_X2 \AES_ENC/us20/U529  ( .A1(\AES_ENC/sa20 [4]), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n764 ) );
NOR2_X2 \AES_ENC/us20/U528  ( .A1(\AES_ENC/us20/n765 ), .A2(\AES_ENC/us20/n764 ), .ZN(\AES_ENC/us20/n766 ) );
NOR2_X2 \AES_ENC/us20/U527  ( .A1(\AES_ENC/us20/n766 ), .A2(\AES_ENC/us20/n589 ), .ZN(\AES_ENC/us20/n767 ) );
INV_X4 \AES_ENC/us20/U526  ( .A(\AES_ENC/sa20 [3]), .ZN(\AES_ENC/us20/n624 ));
NAND3_X2 \AES_ENC/us20/U525  ( .A1(\AES_ENC/us20/n652 ), .A2(\AES_ENC/us20/n596 ), .A3(\AES_ENC/sa20 [7]), .ZN(\AES_ENC/us20/n653 ));
NOR2_X2 \AES_ENC/us20/U524  ( .A1(\AES_ENC/us20/n593 ), .A2(\AES_ENC/sa20 [5]), .ZN(\AES_ENC/us20/n925 ) );
NOR2_X2 \AES_ENC/us20/U523  ( .A1(\AES_ENC/sa20 [5]), .A2(\AES_ENC/sa20 [2]),.ZN(\AES_ENC/us20/n974 ) );
INV_X4 \AES_ENC/us20/U522  ( .A(\AES_ENC/sa20 [5]), .ZN(\AES_ENC/us20/n596 ));
NOR2_X2 \AES_ENC/us20/U521  ( .A1(\AES_ENC/us20/n593 ), .A2(\AES_ENC/sa20 [7]), .ZN(\AES_ENC/us20/n779 ) );
NAND3_X2 \AES_ENC/us20/U520  ( .A1(\AES_ENC/us20/n679 ), .A2(\AES_ENC/us20/n678 ), .A3(\AES_ENC/us20/n677 ), .ZN(\AES_ENC/sa20_sub[0] ) );
NOR2_X2 \AES_ENC/us20/U519  ( .A1(\AES_ENC/us20/n596 ), .A2(\AES_ENC/sa20 [2]), .ZN(\AES_ENC/us20/n1048 ) );
NOR3_X2 \AES_ENC/us20/U518  ( .A1(\AES_ENC/us20/n581 ), .A2(\AES_ENC/sa20 [5]), .A3(\AES_ENC/us20/n704 ), .ZN(\AES_ENC/us20/n706 ));
NOR2_X2 \AES_ENC/us20/U517  ( .A1(\AES_ENC/us20/n1117 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n707 ) );
NOR2_X2 \AES_ENC/us20/U516  ( .A1(\AES_ENC/sa20 [4]), .A2(\AES_ENC/us20/n574 ), .ZN(\AES_ENC/us20/n705 ) );
NOR3_X2 \AES_ENC/us20/U515  ( .A1(\AES_ENC/us20/n707 ), .A2(\AES_ENC/us20/n706 ), .A3(\AES_ENC/us20/n705 ), .ZN(\AES_ENC/us20/n713 ) );
NOR4_X2 \AES_ENC/us20/U512  ( .A1(\AES_ENC/us20/n633 ), .A2(\AES_ENC/us20/n632 ), .A3(\AES_ENC/us20/n631 ), .A4(\AES_ENC/us20/n630 ), .ZN(\AES_ENC/us20/n634 ) );
NOR2_X2 \AES_ENC/us20/U510  ( .A1(\AES_ENC/us20/n629 ), .A2(\AES_ENC/us20/n628 ), .ZN(\AES_ENC/us20/n635 ) );
NAND3_X2 \AES_ENC/us20/U509  ( .A1(\AES_ENC/sa20 [2]), .A2(\AES_ENC/sa20 [7]), .A3(\AES_ENC/us20/n1059 ), .ZN(\AES_ENC/us20/n636 ) );
NOR2_X2 \AES_ENC/us20/U508  ( .A1(\AES_ENC/sa20 [7]), .A2(\AES_ENC/sa20 [2]),.ZN(\AES_ENC/us20/n794 ) );
NOR2_X2 \AES_ENC/us20/U507  ( .A1(\AES_ENC/sa20 [4]), .A2(\AES_ENC/sa20 [1]),.ZN(\AES_ENC/us20/n1102 ) );
NOR2_X2 \AES_ENC/us20/U506  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/sa20 [3]), .ZN(\AES_ENC/us20/n1053 ) );
NOR2_X2 \AES_ENC/us20/U505  ( .A1(\AES_ENC/us20/n588 ), .A2(\AES_ENC/sa20 [5]), .ZN(\AES_ENC/us20/n1024 ) );
NOR2_X2 \AES_ENC/us20/U504  ( .A1(\AES_ENC/us20/n577 ), .A2(\AES_ENC/sa20 [2]), .ZN(\AES_ENC/us20/n1093 ) );
NOR2_X2 \AES_ENC/us20/U503  ( .A1(\AES_ENC/us20/n585 ), .A2(\AES_ENC/sa20 [5]), .ZN(\AES_ENC/us20/n1094 ) );
NOR2_X2 \AES_ENC/us20/U502  ( .A1(\AES_ENC/us20/n612 ), .A2(\AES_ENC/sa20 [3]), .ZN(\AES_ENC/us20/n931 ) );
INV_X4 \AES_ENC/us20/U501  ( .A(\AES_ENC/us20/n570 ), .ZN(\AES_ENC/us20/n573 ) );
NOR2_X2 \AES_ENC/us20/U500  ( .A1(\AES_ENC/us20/n1053 ), .A2(\AES_ENC/us20/n1095 ), .ZN(\AES_ENC/us20/n639 ) );
NOR3_X2 \AES_ENC/us20/U499  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n573 ), .A3(\AES_ENC/us20/n1074 ), .ZN(\AES_ENC/us20/n641 ) );
NOR2_X2 \AES_ENC/us20/U498  ( .A1(\AES_ENC/us20/n639 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n640 ) );
NOR2_X2 \AES_ENC/us20/U497  ( .A1(\AES_ENC/us20/n641 ), .A2(\AES_ENC/us20/n640 ), .ZN(\AES_ENC/us20/n646 ) );
NOR3_X2 \AES_ENC/us20/U496  ( .A1(\AES_ENC/us20/n995 ), .A2(\AES_ENC/us20/n578 ), .A3(\AES_ENC/us20/n994 ), .ZN(\AES_ENC/us20/n1002 ) );
NOR2_X2 \AES_ENC/us20/U495  ( .A1(\AES_ENC/us20/n909 ), .A2(\AES_ENC/us20/n908 ), .ZN(\AES_ENC/us20/n920 ) );
NOR2_X2 \AES_ENC/us20/U494  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n823 ) );
NOR2_X2 \AES_ENC/us20/U492  ( .A1(\AES_ENC/us20/n612 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n822 ) );
NOR2_X2 \AES_ENC/us20/U491  ( .A1(\AES_ENC/us20/n823 ), .A2(\AES_ENC/us20/n822 ), .ZN(\AES_ENC/us20/n825 ) );
NOR2_X2 \AES_ENC/us20/U490  ( .A1(\AES_ENC/sa20 [1]), .A2(\AES_ENC/us20/n601 ), .ZN(\AES_ENC/us20/n913 ) );
NOR2_X2 \AES_ENC/us20/U489  ( .A1(\AES_ENC/us20/n913 ), .A2(\AES_ENC/us20/n1091 ), .ZN(\AES_ENC/us20/n914 ) );
NOR2_X2 \AES_ENC/us20/U488  ( .A1(\AES_ENC/us20/n826 ), .A2(\AES_ENC/us20/n572 ), .ZN(\AES_ENC/us20/n827 ) );
NOR3_X2 \AES_ENC/us20/U487  ( .A1(\AES_ENC/us20/n769 ), .A2(\AES_ENC/us20/n768 ), .A3(\AES_ENC/us20/n767 ), .ZN(\AES_ENC/us20/n775 ) );
NOR2_X2 \AES_ENC/us20/U486  ( .A1(\AES_ENC/us20/n1056 ), .A2(\AES_ENC/us20/n1053 ), .ZN(\AES_ENC/us20/n749 ) );
NOR2_X2 \AES_ENC/us20/U483  ( .A1(\AES_ENC/us20/n749 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n752 ) );
INV_X4 \AES_ENC/us20/U482  ( .A(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n626 ));
NOR2_X2 \AES_ENC/us20/U480  ( .A1(\AES_ENC/us20/n1054 ), .A2(\AES_ENC/us20/n1053 ), .ZN(\AES_ENC/us20/n1055 ) );
OR2_X4 \AES_ENC/us20/U479  ( .A1(\AES_ENC/us20/n1094 ), .A2(\AES_ENC/us20/n1093 ), .ZN(\AES_ENC/us20/n571 ) );
AND2_X2 \AES_ENC/us20/U478  ( .A1(\AES_ENC/us20/n571 ), .A2(\AES_ENC/us20/n1095 ), .ZN(\AES_ENC/us20/n1101 ) );
NOR2_X2 \AES_ENC/us20/U477  ( .A1(\AES_ENC/us20/n1074 ), .A2(\AES_ENC/us20/n931 ), .ZN(\AES_ENC/us20/n796 ) );
NOR2_X2 \AES_ENC/us20/U474  ( .A1(\AES_ENC/us20/n796 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n797 ) );
NOR2_X2 \AES_ENC/us20/U473  ( .A1(\AES_ENC/us20/n932 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n933 ) );
NOR2_X2 \AES_ENC/us20/U472  ( .A1(\AES_ENC/us20/n929 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n935 ) );
NOR2_X2 \AES_ENC/us20/U471  ( .A1(\AES_ENC/us20/n931 ), .A2(\AES_ENC/us20/n930 ), .ZN(\AES_ENC/us20/n934 ) );
NOR3_X2 \AES_ENC/us20/U470  ( .A1(\AES_ENC/us20/n935 ), .A2(\AES_ENC/us20/n934 ), .A3(\AES_ENC/us20/n933 ), .ZN(\AES_ENC/us20/n936 ) );
NOR2_X2 \AES_ENC/us20/U469  ( .A1(\AES_ENC/us20/n612 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n1075 ) );
NOR2_X2 \AES_ENC/us20/U468  ( .A1(\AES_ENC/us20/n572 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n949 ) );
NOR2_X2 \AES_ENC/us20/U467  ( .A1(\AES_ENC/us20/n1049 ), .A2(\AES_ENC/us20/n595 ), .ZN(\AES_ENC/us20/n1051 ) );
NOR2_X2 \AES_ENC/us20/U466  ( .A1(\AES_ENC/us20/n1051 ), .A2(\AES_ENC/us20/n1050 ), .ZN(\AES_ENC/us20/n1052 ) );
NOR2_X2 \AES_ENC/us20/U465  ( .A1(\AES_ENC/us20/n1052 ), .A2(\AES_ENC/us20/n604 ), .ZN(\AES_ENC/us20/n1064 ) );
NOR2_X2 \AES_ENC/us20/U464  ( .A1(\AES_ENC/sa20 [1]), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n631 ) );
NOR2_X2 \AES_ENC/us20/U463  ( .A1(\AES_ENC/us20/n1025 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n980 ) );
NOR2_X2 \AES_ENC/us20/U462  ( .A1(\AES_ENC/us20/n1073 ), .A2(\AES_ENC/us20/n1094 ), .ZN(\AES_ENC/us20/n795 ) );
NOR2_X2 \AES_ENC/us20/U461  ( .A1(\AES_ENC/us20/n795 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n799 ) );
NOR2_X2 \AES_ENC/us20/U460  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n981 ) );
NOR2_X2 \AES_ENC/us20/U459  ( .A1(\AES_ENC/us20/n1102 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n643 ) );
NOR2_X2 \AES_ENC/us20/U458  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n624 ), .ZN(\AES_ENC/us20/n642 ) );
NOR2_X2 \AES_ENC/us20/U455  ( .A1(\AES_ENC/us20/n911 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n644 ) );
NOR4_X2 \AES_ENC/us20/U448  ( .A1(\AES_ENC/us20/n644 ), .A2(\AES_ENC/us20/n643 ), .A3(\AES_ENC/us20/n804 ), .A4(\AES_ENC/us20/n642 ), .ZN(\AES_ENC/us20/n645 ) );
NOR2_X2 \AES_ENC/us20/U447  ( .A1(\AES_ENC/us20/n1102 ), .A2(\AES_ENC/us20/n910 ), .ZN(\AES_ENC/us20/n932 ) );
NOR2_X2 \AES_ENC/us20/U442  ( .A1(\AES_ENC/us20/n1102 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n755 ) );
NOR2_X2 \AES_ENC/us20/U441  ( .A1(\AES_ENC/us20/n931 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n743 ) );
NOR2_X2 \AES_ENC/us20/U438  ( .A1(\AES_ENC/us20/n1072 ), .A2(\AES_ENC/us20/n1094 ), .ZN(\AES_ENC/us20/n930 ) );
NOR2_X2 \AES_ENC/us20/U435  ( .A1(\AES_ENC/us20/n1074 ), .A2(\AES_ENC/us20/n1025 ), .ZN(\AES_ENC/us20/n891 ) );
NOR2_X2 \AES_ENC/us20/U434  ( .A1(\AES_ENC/us20/n891 ), .A2(\AES_ENC/us20/n591 ), .ZN(\AES_ENC/us20/n894 ) );
NOR3_X2 \AES_ENC/us20/U433  ( .A1(\AES_ENC/us20/n601 ), .A2(\AES_ENC/sa20 [1]), .A3(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n683 ));
INV_X4 \AES_ENC/us20/U428  ( .A(\AES_ENC/us20/n931 ), .ZN(\AES_ENC/us20/n601 ) );
NOR2_X2 \AES_ENC/us20/U427  ( .A1(\AES_ENC/us20/n996 ), .A2(\AES_ENC/us20/n931 ), .ZN(\AES_ENC/us20/n704 ) );
NOR2_X2 \AES_ENC/us20/U421  ( .A1(\AES_ENC/us20/n931 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n685 ) );
NOR2_X2 \AES_ENC/us20/U420  ( .A1(\AES_ENC/us20/n1029 ), .A2(\AES_ENC/us20/n1025 ), .ZN(\AES_ENC/us20/n1079 ) );
NOR3_X2 \AES_ENC/us20/U419  ( .A1(\AES_ENC/us20/n620 ), .A2(\AES_ENC/us20/n1025 ), .A3(\AES_ENC/us20/n594 ), .ZN(\AES_ENC/us20/n945 ) );
NOR2_X2 \AES_ENC/us20/U418  ( .A1(\AES_ENC/us20/n596 ), .A2(\AES_ENC/us20/n593 ), .ZN(\AES_ENC/us20/n800 ) );
NOR3_X2 \AES_ENC/us20/U417  ( .A1(\AES_ENC/us20/n598 ), .A2(\AES_ENC/us20/n581 ), .A3(\AES_ENC/us20/n593 ), .ZN(\AES_ENC/us20/n798 ) );
NOR3_X2 \AES_ENC/us20/U416  ( .A1(\AES_ENC/us20/n592 ), .A2(\AES_ENC/us20/n572 ), .A3(\AES_ENC/us20/n589 ), .ZN(\AES_ENC/us20/n962 ) );
NOR3_X2 \AES_ENC/us20/U415  ( .A1(\AES_ENC/us20/n959 ), .A2(\AES_ENC/us20/n572 ), .A3(\AES_ENC/us20/n591 ), .ZN(\AES_ENC/us20/n768 ) );
NOR3_X2 \AES_ENC/us20/U414  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n572 ), .A3(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n694 ) );
NOR3_X2 \AES_ENC/us20/U413  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n572 ), .A3(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n895 ) );
NOR3_X2 \AES_ENC/us20/U410  ( .A1(\AES_ENC/us20/n1008 ), .A2(\AES_ENC/us20/n1007 ), .A3(\AES_ENC/us20/n1006 ), .ZN(\AES_ENC/us20/n1018 ) );
NOR4_X2 \AES_ENC/us20/U409  ( .A1(\AES_ENC/us20/n806 ), .A2(\AES_ENC/us20/n805 ), .A3(\AES_ENC/us20/n804 ), .A4(\AES_ENC/us20/n803 ), .ZN(\AES_ENC/us20/n807 ) );
NOR3_X2 \AES_ENC/us20/U406  ( .A1(\AES_ENC/us20/n799 ), .A2(\AES_ENC/us20/n798 ), .A3(\AES_ENC/us20/n797 ), .ZN(\AES_ENC/us20/n808 ) );
NOR4_X2 \AES_ENC/us20/U405  ( .A1(\AES_ENC/us20/n843 ), .A2(\AES_ENC/us20/n842 ), .A3(\AES_ENC/us20/n841 ), .A4(\AES_ENC/us20/n840 ), .ZN(\AES_ENC/us20/n844 ) );
NOR2_X2 \AES_ENC/us20/U404  ( .A1(\AES_ENC/us20/n669 ), .A2(\AES_ENC/us20/n668 ), .ZN(\AES_ENC/us20/n673 ) );
NOR4_X2 \AES_ENC/us20/U403  ( .A1(\AES_ENC/us20/n946 ), .A2(\AES_ENC/us20/n1046 ), .A3(\AES_ENC/us20/n671 ), .A4(\AES_ENC/us20/n670 ), .ZN(\AES_ENC/us20/n672 ) );
NOR4_X2 \AES_ENC/us20/U401  ( .A1(\AES_ENC/us20/n711 ), .A2(\AES_ENC/us20/n710 ), .A3(\AES_ENC/us20/n709 ), .A4(\AES_ENC/us20/n708 ), .ZN(\AES_ENC/us20/n712 ) );
NOR4_X2 \AES_ENC/us20/U400  ( .A1(\AES_ENC/us20/n963 ), .A2(\AES_ENC/us20/n962 ), .A3(\AES_ENC/us20/n961 ), .A4(\AES_ENC/us20/n960 ), .ZN(\AES_ENC/us20/n964 ) );
NOR3_X2 \AES_ENC/us20/U399  ( .A1(\AES_ENC/us20/n1101 ), .A2(\AES_ENC/us20/n1100 ), .A3(\AES_ENC/us20/n1099 ), .ZN(\AES_ENC/us20/n1109 ) );
NOR3_X2 \AES_ENC/us20/U398  ( .A1(\AES_ENC/us20/n743 ), .A2(\AES_ENC/us20/n742 ), .A3(\AES_ENC/us20/n741 ), .ZN(\AES_ENC/us20/n744 ) );
NOR2_X2 \AES_ENC/us20/U397  ( .A1(\AES_ENC/us20/n697 ), .A2(\AES_ENC/us20/n658 ), .ZN(\AES_ENC/us20/n659 ) );
NOR2_X2 \AES_ENC/us20/U396  ( .A1(\AES_ENC/us20/n1078 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n1033 ) );
NOR2_X2 \AES_ENC/us20/U393  ( .A1(\AES_ENC/us20/n1031 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n1032 ) );
NOR3_X2 \AES_ENC/us20/U390  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n1025 ), .A3(\AES_ENC/us20/n1074 ), .ZN(\AES_ENC/us20/n1035 ) );
NOR4_X2 \AES_ENC/us20/U389  ( .A1(\AES_ENC/us20/n1035 ), .A2(\AES_ENC/us20/n1034 ), .A3(\AES_ENC/us20/n1033 ), .A4(\AES_ENC/us20/n1032 ), .ZN(\AES_ENC/us20/n1036 ) );
NOR2_X2 \AES_ENC/us20/U388  ( .A1(\AES_ENC/us20/n611 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n885 ) );
NOR2_X2 \AES_ENC/us20/U387  ( .A1(\AES_ENC/us20/n601 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n882 ) );
NOR2_X2 \AES_ENC/us20/U386  ( .A1(\AES_ENC/us20/n1053 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n884 ) );
NOR4_X2 \AES_ENC/us20/U385  ( .A1(\AES_ENC/us20/n885 ), .A2(\AES_ENC/us20/n884 ), .A3(\AES_ENC/us20/n883 ), .A4(\AES_ENC/us20/n882 ), .ZN(\AES_ENC/us20/n886 ) );
NOR2_X2 \AES_ENC/us20/U384  ( .A1(\AES_ENC/us20/n825 ), .A2(\AES_ENC/us20/n590 ), .ZN(\AES_ENC/us20/n830 ) );
NOR2_X2 \AES_ENC/us20/U383  ( .A1(\AES_ENC/us20/n827 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n829 ) );
NOR2_X2 \AES_ENC/us20/U382  ( .A1(\AES_ENC/us20/n572 ), .A2(\AES_ENC/us20/n574 ), .ZN(\AES_ENC/us20/n828 ) );
NOR4_X2 \AES_ENC/us20/U374  ( .A1(\AES_ENC/us20/n831 ), .A2(\AES_ENC/us20/n830 ), .A3(\AES_ENC/us20/n829 ), .A4(\AES_ENC/us20/n828 ), .ZN(\AES_ENC/us20/n832 ) );
NOR2_X2 \AES_ENC/us20/U373  ( .A1(\AES_ENC/us20/n587 ), .A2(\AES_ENC/us20/n603 ), .ZN(\AES_ENC/us20/n1104 ) );
NOR2_X2 \AES_ENC/us20/U372  ( .A1(\AES_ENC/us20/n1102 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n1106 ) );
NOR2_X2 \AES_ENC/us20/U370  ( .A1(\AES_ENC/us20/n1103 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n1105 ) );
NOR4_X2 \AES_ENC/us20/U369  ( .A1(\AES_ENC/us20/n1107 ), .A2(\AES_ENC/us20/n1106 ), .A3(\AES_ENC/us20/n1105 ), .A4(\AES_ENC/us20/n1104 ), .ZN(\AES_ENC/us20/n1108 ) );
NOR3_X2 \AES_ENC/us20/U368  ( .A1(\AES_ENC/us20/n959 ), .A2(\AES_ENC/us20/n624 ), .A3(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n963 ) );
NOR2_X2 \AES_ENC/us20/U367  ( .A1(\AES_ENC/us20/n596 ), .A2(\AES_ENC/us20/n581 ), .ZN(\AES_ENC/us20/n1114 ) );
INV_X4 \AES_ENC/us20/U366  ( .A(\AES_ENC/us20/n1024 ), .ZN(\AES_ENC/us20/n587 ) );
NOR3_X2 \AES_ENC/us20/U365  ( .A1(\AES_ENC/us20/n910 ), .A2(\AES_ENC/us20/n1059 ), .A3(\AES_ENC/us20/n593 ), .ZN(\AES_ENC/us20/n1115 ) );
INV_X4 \AES_ENC/us20/U364  ( .A(\AES_ENC/us20/n1094 ), .ZN(\AES_ENC/us20/n584 ) );
NOR2_X2 \AES_ENC/us20/U363  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n931 ), .ZN(\AES_ENC/us20/n1100 ) );
INV_X4 \AES_ENC/us20/U354  ( .A(\AES_ENC/us20/n1093 ), .ZN(\AES_ENC/us20/n575 ) );
NOR2_X2 \AES_ENC/us20/U353  ( .A1(\AES_ENC/us20/n569 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n929 ) );
NOR2_X2 \AES_ENC/us20/U352  ( .A1(\AES_ENC/us20/n609 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n926 ) );
NOR2_X2 \AES_ENC/us20/U351  ( .A1(\AES_ENC/us20/n572 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n1095 ) );
NOR2_X2 \AES_ENC/us20/U350  ( .A1(\AES_ENC/us20/n591 ), .A2(\AES_ENC/us20/n581 ), .ZN(\AES_ENC/us20/n1010 ) );
NOR2_X2 \AES_ENC/us20/U349  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n1103 ) );
NOR2_X2 \AES_ENC/us20/U348  ( .A1(\AES_ENC/us20/n614 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n1059 ) );
NOR2_X2 \AES_ENC/us20/U347  ( .A1(\AES_ENC/sa20 [1]), .A2(\AES_ENC/us20/n1120 ), .ZN(\AES_ENC/us20/n1022 ) );
NOR2_X2 \AES_ENC/us20/U346  ( .A1(\AES_ENC/us20/n605 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n911 ) );
NOR2_X2 \AES_ENC/us20/U345  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/us20/n1025 ), .ZN(\AES_ENC/us20/n826 ) );
NOR2_X2 \AES_ENC/us20/U338  ( .A1(\AES_ENC/us20/n596 ), .A2(\AES_ENC/us20/n588 ), .ZN(\AES_ENC/us20/n1072 ) );
NOR2_X2 \AES_ENC/us20/U335  ( .A1(\AES_ENC/us20/n581 ), .A2(\AES_ENC/us20/n594 ), .ZN(\AES_ENC/us20/n956 ) );
NOR2_X2 \AES_ENC/us20/U329  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/us20/n612 ), .ZN(\AES_ENC/us20/n1121 ) );
NOR2_X2 \AES_ENC/us20/U328  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/us20/n612 ), .ZN(\AES_ENC/us20/n1058 ) );
NOR2_X2 \AES_ENC/us20/U327  ( .A1(\AES_ENC/us20/n577 ), .A2(\AES_ENC/us20/n593 ), .ZN(\AES_ENC/us20/n1073 ) );
NOR2_X2 \AES_ENC/us20/U325  ( .A1(\AES_ENC/sa20 [1]), .A2(\AES_ENC/us20/n1025 ), .ZN(\AES_ENC/us20/n1054 ) );
NOR2_X2 \AES_ENC/us20/U324  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/us20/n931 ), .ZN(\AES_ENC/us20/n1029 ) );
NOR2_X2 \AES_ENC/us20/U319  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n1056 ) );
NOR2_X2 \AES_ENC/us20/U318  ( .A1(\AES_ENC/us20/n585 ), .A2(\AES_ENC/us20/n596 ), .ZN(\AES_ENC/us20/n1050 ) );
NOR2_X2 \AES_ENC/us20/U317  ( .A1(\AES_ENC/us20/n1121 ), .A2(\AES_ENC/us20/n1025 ), .ZN(\AES_ENC/us20/n1120 ) );
NOR2_X2 \AES_ENC/us20/U316  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/us20/n572 ), .ZN(\AES_ENC/us20/n1074 ) );
NOR2_X2 \AES_ENC/us20/U315  ( .A1(\AES_ENC/us20/n1058 ), .A2(\AES_ENC/us20/n1054 ), .ZN(\AES_ENC/us20/n878 ) );
NOR2_X2 \AES_ENC/us20/U314  ( .A1(\AES_ENC/us20/n878 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n879 ) );
NOR2_X2 \AES_ENC/us20/U312  ( .A1(\AES_ENC/us20/n880 ), .A2(\AES_ENC/us20/n879 ), .ZN(\AES_ENC/us20/n887 ) );
NOR2_X2 \AES_ENC/us20/U311  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n625 ), .ZN(\AES_ENC/us20/n957 ) );
NOR2_X2 \AES_ENC/us20/U310  ( .A1(\AES_ENC/us20/n958 ), .A2(\AES_ENC/us20/n957 ), .ZN(\AES_ENC/us20/n965 ) );
NOR3_X2 \AES_ENC/us20/U309  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n1091 ), .A3(\AES_ENC/us20/n1022 ), .ZN(\AES_ENC/us20/n720 ) );
NOR3_X2 \AES_ENC/us20/U303  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n1054 ), .A3(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n719 ) );
NOR2_X2 \AES_ENC/us20/U302  ( .A1(\AES_ENC/us20/n720 ), .A2(\AES_ENC/us20/n719 ), .ZN(\AES_ENC/us20/n726 ) );
NOR2_X2 \AES_ENC/us20/U300  ( .A1(\AES_ENC/us20/n585 ), .A2(\AES_ENC/us20/n613 ), .ZN(\AES_ENC/us20/n865 ) );
NOR2_X2 \AES_ENC/us20/U299  ( .A1(\AES_ENC/us20/n1059 ), .A2(\AES_ENC/us20/n1058 ), .ZN(\AES_ENC/us20/n1060 ) );
NOR2_X2 \AES_ENC/us20/U298  ( .A1(\AES_ENC/us20/n1095 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n668 ) );
NOR2_X2 \AES_ENC/us20/U297  ( .A1(\AES_ENC/us20/n826 ), .A2(\AES_ENC/us20/n573 ), .ZN(\AES_ENC/us20/n750 ) );
NOR2_X2 \AES_ENC/us20/U296  ( .A1(\AES_ENC/us20/n750 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n751 ) );
NOR2_X2 \AES_ENC/us20/U295  ( .A1(\AES_ENC/us20/n907 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n908 ) );
NOR2_X2 \AES_ENC/us20/U294  ( .A1(\AES_ENC/us20/n990 ), .A2(\AES_ENC/us20/n926 ), .ZN(\AES_ENC/us20/n780 ) );
NOR2_X2 \AES_ENC/us20/U293  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n606 ), .ZN(\AES_ENC/us20/n838 ) );
NOR2_X2 \AES_ENC/us20/U292  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n621 ), .ZN(\AES_ENC/us20/n837 ) );
NOR2_X2 \AES_ENC/us20/U291  ( .A1(\AES_ENC/us20/n838 ), .A2(\AES_ENC/us20/n837 ), .ZN(\AES_ENC/us20/n845 ) );
NOR2_X2 \AES_ENC/us20/U290  ( .A1(\AES_ENC/us20/n1022 ), .A2(\AES_ENC/us20/n1058 ), .ZN(\AES_ENC/us20/n740 ) );
NOR2_X2 \AES_ENC/us20/U284  ( .A1(\AES_ENC/us20/n740 ), .A2(\AES_ENC/us20/n594 ), .ZN(\AES_ENC/us20/n742 ) );
NOR2_X2 \AES_ENC/us20/U283  ( .A1(\AES_ENC/us20/n1098 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n1099 ) );
NOR2_X2 \AES_ENC/us20/U282  ( .A1(\AES_ENC/us20/n1120 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n993 ) );
NOR2_X2 \AES_ENC/us20/U281  ( .A1(\AES_ENC/us20/n993 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n994 ) );
NOR2_X2 \AES_ENC/us20/U280  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n609 ), .ZN(\AES_ENC/us20/n1026 ) );
NOR2_X2 \AES_ENC/us20/U279  ( .A1(\AES_ENC/us20/n573 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n1027 ) );
NOR2_X2 \AES_ENC/us20/U273  ( .A1(\AES_ENC/us20/n1027 ), .A2(\AES_ENC/us20/n1026 ), .ZN(\AES_ENC/us20/n1028 ) );
NOR2_X2 \AES_ENC/us20/U272  ( .A1(\AES_ENC/us20/n1029 ), .A2(\AES_ENC/us20/n1028 ), .ZN(\AES_ENC/us20/n1034 ) );
NOR4_X2 \AES_ENC/us20/U271  ( .A1(\AES_ENC/us20/n757 ), .A2(\AES_ENC/us20/n756 ), .A3(\AES_ENC/us20/n755 ), .A4(\AES_ENC/us20/n754 ), .ZN(\AES_ENC/us20/n758 ) );
NOR2_X2 \AES_ENC/us20/U270  ( .A1(\AES_ENC/us20/n752 ), .A2(\AES_ENC/us20/n751 ), .ZN(\AES_ENC/us20/n759 ) );
NOR2_X2 \AES_ENC/us20/U269  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n1071 ), .ZN(\AES_ENC/us20/n669 ) );
NOR2_X2 \AES_ENC/us20/U268  ( .A1(\AES_ENC/us20/n1056 ), .A2(\AES_ENC/us20/n990 ), .ZN(\AES_ENC/us20/n991 ) );
NOR2_X2 \AES_ENC/us20/U267  ( .A1(\AES_ENC/us20/n991 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n995 ) );
NOR2_X2 \AES_ENC/us20/U263  ( .A1(\AES_ENC/us20/n588 ), .A2(\AES_ENC/us20/n598 ), .ZN(\AES_ENC/us20/n1008 ) );
NOR2_X2 \AES_ENC/us20/U262  ( .A1(\AES_ENC/us20/n839 ), .A2(\AES_ENC/us20/n603 ), .ZN(\AES_ENC/us20/n693 ) );
NOR2_X2 \AES_ENC/us20/U258  ( .A1(\AES_ENC/us20/n587 ), .A2(\AES_ENC/us20/n906 ), .ZN(\AES_ENC/us20/n741 ) );
NOR2_X2 \AES_ENC/us20/U255  ( .A1(\AES_ENC/us20/n1054 ), .A2(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n763 ) );
NOR2_X2 \AES_ENC/us20/U254  ( .A1(\AES_ENC/us20/n763 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n769 ) );
NOR2_X2 \AES_ENC/us20/U253  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n618 ), .ZN(\AES_ENC/us20/n1007 ) );
NOR2_X2 \AES_ENC/us20/U252  ( .A1(\AES_ENC/us20/n591 ), .A2(\AES_ENC/us20/n599 ), .ZN(\AES_ENC/us20/n1123 ) );
NOR2_X2 \AES_ENC/us20/U251  ( .A1(\AES_ENC/us20/n591 ), .A2(\AES_ENC/us20/n598 ), .ZN(\AES_ENC/us20/n710 ) );
INV_X4 \AES_ENC/us20/U250  ( .A(\AES_ENC/us20/n1029 ), .ZN(\AES_ENC/us20/n603 ) );
NOR2_X2 \AES_ENC/us20/U243  ( .A1(\AES_ENC/us20/n594 ), .A2(\AES_ENC/us20/n607 ), .ZN(\AES_ENC/us20/n883 ) );
NOR2_X2 \AES_ENC/us20/U242  ( .A1(\AES_ENC/us20/n623 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n1125 ) );
NOR2_X2 \AES_ENC/us20/U241  ( .A1(\AES_ENC/us20/n911 ), .A2(\AES_ENC/us20/n910 ), .ZN(\AES_ENC/us20/n912 ) );
NOR2_X2 \AES_ENC/us20/U240  ( .A1(\AES_ENC/us20/n912 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n916 ) );
NOR2_X2 \AES_ENC/us20/U239  ( .A1(\AES_ENC/us20/n990 ), .A2(\AES_ENC/us20/n929 ), .ZN(\AES_ENC/us20/n892 ) );
NOR2_X2 \AES_ENC/us20/U238  ( .A1(\AES_ENC/us20/n892 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n893 ) );
NOR2_X2 \AES_ENC/us20/U237  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n621 ), .ZN(\AES_ENC/us20/n950 ) );
NOR2_X2 \AES_ENC/us20/U236  ( .A1(\AES_ENC/us20/n1079 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n1082 ) );
NOR2_X2 \AES_ENC/us20/U235  ( .A1(\AES_ENC/us20/n910 ), .A2(\AES_ENC/us20/n1056 ), .ZN(\AES_ENC/us20/n941 ) );
NOR2_X2 \AES_ENC/us20/U234  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n1077 ), .ZN(\AES_ENC/us20/n841 ) );
NOR2_X2 \AES_ENC/us20/U229  ( .A1(\AES_ENC/us20/n601 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n630 ) );
NOR2_X2 \AES_ENC/us20/U228  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n621 ), .ZN(\AES_ENC/us20/n806 ) );
NOR2_X2 \AES_ENC/us20/U227  ( .A1(\AES_ENC/us20/n601 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n948 ) );
NOR2_X2 \AES_ENC/us20/U226  ( .A1(\AES_ENC/us20/n587 ), .A2(\AES_ENC/us20/n620 ), .ZN(\AES_ENC/us20/n997 ) );
NOR2_X2 \AES_ENC/us20/U225  ( .A1(\AES_ENC/us20/n1121 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n1122 ) );
NOR2_X2 \AES_ENC/us20/U223  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n1023 ), .ZN(\AES_ENC/us20/n756 ) );
NOR2_X2 \AES_ENC/us20/U222  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n621 ), .ZN(\AES_ENC/us20/n870 ) );
NOR2_X2 \AES_ENC/us20/U221  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n569 ), .ZN(\AES_ENC/us20/n947 ) );
NOR2_X2 \AES_ENC/us20/U217  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n1077 ), .ZN(\AES_ENC/us20/n1084 ) );
NOR2_X2 \AES_ENC/us20/U213  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n855 ), .ZN(\AES_ENC/us20/n709 ) );
NOR2_X2 \AES_ENC/us20/U212  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n620 ), .ZN(\AES_ENC/us20/n868 ) );
NOR2_X2 \AES_ENC/us20/U211  ( .A1(\AES_ENC/us20/n1120 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n1124 ) );
NOR2_X2 \AES_ENC/us20/U210  ( .A1(\AES_ENC/us20/n1120 ), .A2(\AES_ENC/us20/n839 ), .ZN(\AES_ENC/us20/n842 ) );
NOR2_X2 \AES_ENC/us20/U209  ( .A1(\AES_ENC/us20/n1120 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n696 ) );
NOR2_X2 \AES_ENC/us20/U208  ( .A1(\AES_ENC/us20/n1074 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n1076 ) );
NOR2_X2 \AES_ENC/us20/U207  ( .A1(\AES_ENC/us20/n1074 ), .A2(\AES_ENC/us20/n609 ), .ZN(\AES_ENC/us20/n781 ) );
NOR3_X2 \AES_ENC/us20/U201  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n1056 ), .A3(\AES_ENC/us20/n990 ), .ZN(\AES_ENC/us20/n979 ) );
NOR3_X2 \AES_ENC/us20/U200  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n1058 ), .A3(\AES_ENC/us20/n1059 ), .ZN(\AES_ENC/us20/n854 ) );
NOR2_X2 \AES_ENC/us20/U199  ( .A1(\AES_ENC/us20/n996 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n869 ) );
NOR2_X2 \AES_ENC/us20/U198  ( .A1(\AES_ENC/us20/n1056 ), .A2(\AES_ENC/us20/n1074 ), .ZN(\AES_ENC/us20/n1057 ) );
NOR3_X2 \AES_ENC/us20/U197  ( .A1(\AES_ENC/us20/n588 ), .A2(\AES_ENC/us20/n1120 ), .A3(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n978 ) );
NOR2_X2 \AES_ENC/us20/U196  ( .A1(\AES_ENC/us20/n996 ), .A2(\AES_ENC/us20/n911 ), .ZN(\AES_ENC/us20/n1116 ) );
NOR2_X2 \AES_ENC/us20/U195  ( .A1(\AES_ENC/us20/n1074 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n754 ) );
NOR2_X2 \AES_ENC/us20/U194  ( .A1(\AES_ENC/us20/n926 ), .A2(\AES_ENC/us20/n1103 ), .ZN(\AES_ENC/us20/n977 ) );
NOR2_X2 \AES_ENC/us20/U187  ( .A1(\AES_ENC/us20/n839 ), .A2(\AES_ENC/us20/n824 ), .ZN(\AES_ENC/us20/n1092 ) );
NOR2_X2 \AES_ENC/us20/U186  ( .A1(\AES_ENC/us20/n573 ), .A2(\AES_ENC/us20/n1074 ), .ZN(\AES_ENC/us20/n684 ) );
NOR2_X2 \AES_ENC/us20/U185  ( .A1(\AES_ENC/us20/n826 ), .A2(\AES_ENC/us20/n1059 ), .ZN(\AES_ENC/us20/n907 ) );
NOR3_X2 \AES_ENC/us20/U184  ( .A1(\AES_ENC/us20/n577 ), .A2(\AES_ENC/us20/n1115 ), .A3(\AES_ENC/us20/n600 ), .ZN(\AES_ENC/us20/n831 ) );
NOR3_X2 \AES_ENC/us20/U183  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n1056 ), .A3(\AES_ENC/us20/n990 ), .ZN(\AES_ENC/us20/n896 ) );
NOR3_X2 \AES_ENC/us20/U182  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n573 ), .A3(\AES_ENC/us20/n1013 ), .ZN(\AES_ENC/us20/n670 ) );
NOR3_X2 \AES_ENC/us20/U181  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n1091 ), .A3(\AES_ENC/us20/n1022 ), .ZN(\AES_ENC/us20/n843 ) );
NOR2_X2 \AES_ENC/us20/U180  ( .A1(\AES_ENC/us20/n1029 ), .A2(\AES_ENC/us20/n1095 ), .ZN(\AES_ENC/us20/n735 ) );
NOR2_X2 \AES_ENC/us20/U174  ( .A1(\AES_ENC/us20/n1100 ), .A2(\AES_ENC/us20/n854 ), .ZN(\AES_ENC/us20/n860 ) );
NAND3_X2 \AES_ENC/us20/U173  ( .A1(\AES_ENC/us20/n569 ), .A2(\AES_ENC/us20/n603 ), .A3(\AES_ENC/us20/n681 ), .ZN(\AES_ENC/us20/n691 ) );
NOR2_X2 \AES_ENC/us20/U172  ( .A1(\AES_ENC/us20/n683 ), .A2(\AES_ENC/us20/n682 ), .ZN(\AES_ENC/us20/n690 ) );
NOR3_X2 \AES_ENC/us20/U171  ( .A1(\AES_ENC/us20/n695 ), .A2(\AES_ENC/us20/n694 ), .A3(\AES_ENC/us20/n693 ), .ZN(\AES_ENC/us20/n700 ) );
NOR4_X2 \AES_ENC/us20/U170  ( .A1(\AES_ENC/us20/n983 ), .A2(\AES_ENC/us20/n698 ), .A3(\AES_ENC/us20/n697 ), .A4(\AES_ENC/us20/n696 ), .ZN(\AES_ENC/us20/n699 ) );
NOR2_X2 \AES_ENC/us20/U169  ( .A1(\AES_ENC/us20/n946 ), .A2(\AES_ENC/us20/n945 ), .ZN(\AES_ENC/us20/n952 ) );
NOR4_X2 \AES_ENC/us20/U168  ( .A1(\AES_ENC/us20/n950 ), .A2(\AES_ENC/us20/n949 ), .A3(\AES_ENC/us20/n948 ), .A4(\AES_ENC/us20/n947 ), .ZN(\AES_ENC/us20/n951 ) );
NOR4_X2 \AES_ENC/us20/U162  ( .A1(\AES_ENC/us20/n896 ), .A2(\AES_ENC/us20/n895 ), .A3(\AES_ENC/us20/n894 ), .A4(\AES_ENC/us20/n893 ), .ZN(\AES_ENC/us20/n897 ) );
NOR2_X2 \AES_ENC/us20/U161  ( .A1(\AES_ENC/us20/n866 ), .A2(\AES_ENC/us20/n865 ), .ZN(\AES_ENC/us20/n872 ) );
NOR4_X2 \AES_ENC/us20/U160  ( .A1(\AES_ENC/us20/n870 ), .A2(\AES_ENC/us20/n869 ), .A3(\AES_ENC/us20/n868 ), .A4(\AES_ENC/us20/n867 ), .ZN(\AES_ENC/us20/n871 ) );
NOR4_X2 \AES_ENC/us20/U159  ( .A1(\AES_ENC/us20/n983 ), .A2(\AES_ENC/us20/n982 ), .A3(\AES_ENC/us20/n981 ), .A4(\AES_ENC/us20/n980 ), .ZN(\AES_ENC/us20/n984 ) );
NOR2_X2 \AES_ENC/us20/U158  ( .A1(\AES_ENC/us20/n979 ), .A2(\AES_ENC/us20/n978 ), .ZN(\AES_ENC/us20/n985 ) );
NOR4_X2 \AES_ENC/us20/U157  ( .A1(\AES_ENC/us20/n1125 ), .A2(\AES_ENC/us20/n1124 ), .A3(\AES_ENC/us20/n1123 ), .A4(\AES_ENC/us20/n1122 ), .ZN(\AES_ENC/us20/n1126 ) );
NOR4_X2 \AES_ENC/us20/U156  ( .A1(\AES_ENC/us20/n1084 ), .A2(\AES_ENC/us20/n1083 ), .A3(\AES_ENC/us20/n1082 ), .A4(\AES_ENC/us20/n1081 ), .ZN(\AES_ENC/us20/n1085 ) );
NOR2_X2 \AES_ENC/us20/U155  ( .A1(\AES_ENC/us20/n1076 ), .A2(\AES_ENC/us20/n1075 ), .ZN(\AES_ENC/us20/n1086 ) );
NOR3_X2 \AES_ENC/us20/U154  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n1054 ), .A3(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n961 ) );
NOR3_X2 \AES_ENC/us20/U153  ( .A1(\AES_ENC/us20/n609 ), .A2(\AES_ENC/us20/n1074 ), .A3(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n671 ) );
NOR2_X2 \AES_ENC/us20/U152  ( .A1(\AES_ENC/us20/n1057 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n1062 ) );
NOR2_X2 \AES_ENC/us20/U143  ( .A1(\AES_ENC/us20/n1055 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n1063 ) );
NOR2_X2 \AES_ENC/us20/U142  ( .A1(\AES_ENC/us20/n1060 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n1061 ) );
NOR4_X2 \AES_ENC/us20/U141  ( .A1(\AES_ENC/us20/n1064 ), .A2(\AES_ENC/us20/n1063 ), .A3(\AES_ENC/us20/n1062 ), .A4(\AES_ENC/us20/n1061 ), .ZN(\AES_ENC/us20/n1065 ) );
NOR3_X2 \AES_ENC/us20/U140  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n1120 ), .A3(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n918 ) );
NOR3_X2 \AES_ENC/us20/U132  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n573 ), .A3(\AES_ENC/us20/n1013 ), .ZN(\AES_ENC/us20/n917 ) );
NOR2_X2 \AES_ENC/us20/U131  ( .A1(\AES_ENC/us20/n914 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n915 ) );
NOR4_X2 \AES_ENC/us20/U130  ( .A1(\AES_ENC/us20/n918 ), .A2(\AES_ENC/us20/n917 ), .A3(\AES_ENC/us20/n916 ), .A4(\AES_ENC/us20/n915 ), .ZN(\AES_ENC/us20/n919 ) );
NOR2_X2 \AES_ENC/us20/U129  ( .A1(\AES_ENC/us20/n594 ), .A2(\AES_ENC/us20/n599 ), .ZN(\AES_ENC/us20/n771 ) );
NOR2_X2 \AES_ENC/us20/U128  ( .A1(\AES_ENC/us20/n1103 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n772 ) );
NOR2_X2 \AES_ENC/us20/U127  ( .A1(\AES_ENC/us20/n592 ), .A2(\AES_ENC/us20/n615 ), .ZN(\AES_ENC/us20/n773 ) );
NOR4_X2 \AES_ENC/us20/U126  ( .A1(\AES_ENC/us20/n773 ), .A2(\AES_ENC/us20/n772 ), .A3(\AES_ENC/us20/n771 ), .A4(\AES_ENC/us20/n770 ), .ZN(\AES_ENC/us20/n774 ) );
NOR2_X2 \AES_ENC/us20/U121  ( .A1(\AES_ENC/us20/n735 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n687 ) );
NOR2_X2 \AES_ENC/us20/U120  ( .A1(\AES_ENC/us20/n684 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n688 ) );
NOR2_X2 \AES_ENC/us20/U119  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n622 ), .ZN(\AES_ENC/us20/n686 ) );
NOR4_X2 \AES_ENC/us20/U118  ( .A1(\AES_ENC/us20/n688 ), .A2(\AES_ENC/us20/n687 ), .A3(\AES_ENC/us20/n686 ), .A4(\AES_ENC/us20/n685 ), .ZN(\AES_ENC/us20/n689 ) );
NOR2_X2 \AES_ENC/us20/U117  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n608 ), .ZN(\AES_ENC/us20/n858 ) );
NOR2_X2 \AES_ENC/us20/U116  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n855 ), .ZN(\AES_ENC/us20/n857 ) );
NOR2_X2 \AES_ENC/us20/U115  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n617 ), .ZN(\AES_ENC/us20/n856 ) );
NOR4_X2 \AES_ENC/us20/U106  ( .A1(\AES_ENC/us20/n858 ), .A2(\AES_ENC/us20/n857 ), .A3(\AES_ENC/us20/n856 ), .A4(\AES_ENC/us20/n958 ), .ZN(\AES_ENC/us20/n859 ) );
NOR2_X2 \AES_ENC/us20/U105  ( .A1(\AES_ENC/us20/n780 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n784 ) );
NOR2_X2 \AES_ENC/us20/U104  ( .A1(\AES_ENC/us20/n1117 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n782 ) );
NOR2_X2 \AES_ENC/us20/U103  ( .A1(\AES_ENC/us20/n781 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n783 ) );
NOR4_X2 \AES_ENC/us20/U102  ( .A1(\AES_ENC/us20/n880 ), .A2(\AES_ENC/us20/n784 ), .A3(\AES_ENC/us20/n783 ), .A4(\AES_ENC/us20/n782 ), .ZN(\AES_ENC/us20/n785 ) );
NOR2_X2 \AES_ENC/us20/U101  ( .A1(\AES_ENC/us20/n597 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n814 ) );
NOR2_X2 \AES_ENC/us20/U100  ( .A1(\AES_ENC/us20/n907 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n813 ) );
NOR3_X2 \AES_ENC/us20/U95  ( .A1(\AES_ENC/us20/n587 ), .A2(\AES_ENC/us20/n1058 ), .A3(\AES_ENC/us20/n1059 ), .ZN(\AES_ENC/us20/n815 ) );
NOR4_X2 \AES_ENC/us20/U94  ( .A1(\AES_ENC/us20/n815 ), .A2(\AES_ENC/us20/n814 ), .A3(\AES_ENC/us20/n813 ), .A4(\AES_ENC/us20/n812 ), .ZN(\AES_ENC/us20/n816 ) );
NOR2_X2 \AES_ENC/us20/U93  ( .A1(\AES_ENC/us20/n575 ), .A2(\AES_ENC/us20/n569 ), .ZN(\AES_ENC/us20/n721 ) );
NOR2_X2 \AES_ENC/us20/U92  ( .A1(\AES_ENC/us20/n1031 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n723 ) );
NOR2_X2 \AES_ENC/us20/U91  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n1096 ), .ZN(\AES_ENC/us20/n722 ) );
NOR4_X2 \AES_ENC/us20/U90  ( .A1(\AES_ENC/us20/n724 ), .A2(\AES_ENC/us20/n723 ), .A3(\AES_ENC/us20/n722 ), .A4(\AES_ENC/us20/n721 ), .ZN(\AES_ENC/us20/n725 ) );
NOR2_X2 \AES_ENC/us20/U89  ( .A1(\AES_ENC/us20/n911 ), .A2(\AES_ENC/us20/n990 ), .ZN(\AES_ENC/us20/n1009 ) );
NOR2_X2 \AES_ENC/us20/U88  ( .A1(\AES_ENC/us20/n1013 ), .A2(\AES_ENC/us20/n573 ), .ZN(\AES_ENC/us20/n1014 ) );
NOR2_X2 \AES_ENC/us20/U87  ( .A1(\AES_ENC/us20/n1014 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n1015 ) );
NOR4_X2 \AES_ENC/us20/U86  ( .A1(\AES_ENC/us20/n1016 ), .A2(\AES_ENC/us20/n1015 ), .A3(\AES_ENC/us20/n1119 ), .A4(\AES_ENC/us20/n1046 ), .ZN(\AES_ENC/us20/n1017 ) );
NOR2_X2 \AES_ENC/us20/U81  ( .A1(\AES_ENC/us20/n996 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n998 ) );
NOR2_X2 \AES_ENC/us20/U80  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n618 ), .ZN(\AES_ENC/us20/n1000 ) );
NOR2_X2 \AES_ENC/us20/U79  ( .A1(\AES_ENC/us20/n594 ), .A2(\AES_ENC/us20/n1096 ), .ZN(\AES_ENC/us20/n999 ) );
NOR4_X2 \AES_ENC/us20/U78  ( .A1(\AES_ENC/us20/n1000 ), .A2(\AES_ENC/us20/n999 ), .A3(\AES_ENC/us20/n998 ), .A4(\AES_ENC/us20/n997 ), .ZN(\AES_ENC/us20/n1001 ) );
NOR2_X2 \AES_ENC/us20/U74  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n1096 ), .ZN(\AES_ENC/us20/n697 ) );
NOR2_X2 \AES_ENC/us20/U73  ( .A1(\AES_ENC/us20/n609 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n958 ) );
NOR2_X2 \AES_ENC/us20/U72  ( .A1(\AES_ENC/us20/n911 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n983 ) );
NOR2_X2 \AES_ENC/us20/U71  ( .A1(\AES_ENC/us20/n1054 ), .A2(\AES_ENC/us20/n1103 ), .ZN(\AES_ENC/us20/n1031 ) );
INV_X4 \AES_ENC/us20/U65  ( .A(\AES_ENC/us20/n1050 ), .ZN(\AES_ENC/us20/n582 ) );
INV_X4 \AES_ENC/us20/U64  ( .A(\AES_ENC/us20/n1072 ), .ZN(\AES_ENC/us20/n586 ) );
INV_X4 \AES_ENC/us20/U63  ( .A(\AES_ENC/us20/n1073 ), .ZN(\AES_ENC/us20/n576 ) );
NOR2_X2 \AES_ENC/us20/U62  ( .A1(\AES_ENC/us20/n603 ), .A2(\AES_ENC/us20/n584 ), .ZN(\AES_ENC/us20/n880 ) );
NOR3_X2 \AES_ENC/us20/U61  ( .A1(\AES_ENC/us20/n826 ), .A2(\AES_ENC/us20/n1121 ), .A3(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n946 ) );
INV_X4 \AES_ENC/us20/U59  ( .A(\AES_ENC/us20/n1010 ), .ZN(\AES_ENC/us20/n579 ) );
NOR3_X2 \AES_ENC/us20/U58  ( .A1(\AES_ENC/us20/n573 ), .A2(\AES_ENC/us20/n1029 ), .A3(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n1119 ) );
INV_X4 \AES_ENC/us20/U57  ( .A(\AES_ENC/us20/n956 ), .ZN(\AES_ENC/us20/n580 ) );
NOR2_X2 \AES_ENC/us20/U50  ( .A1(\AES_ENC/us20/n601 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n1013 ) );
NOR2_X2 \AES_ENC/us20/U49  ( .A1(\AES_ENC/us20/n609 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n910 ) );
NOR2_X2 \AES_ENC/us20/U48  ( .A1(\AES_ENC/us20/n569 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n1091 ) );
NOR2_X2 \AES_ENC/us20/U47  ( .A1(\AES_ENC/us20/n614 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n990 ) );
NOR2_X2 \AES_ENC/us20/U46  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/us20/n1121 ), .ZN(\AES_ENC/us20/n996 ) );
NOR2_X2 \AES_ENC/us20/U45  ( .A1(\AES_ENC/us20/n592 ), .A2(\AES_ENC/us20/n622 ), .ZN(\AES_ENC/us20/n628 ) );
NOR2_X2 \AES_ENC/us20/U44  ( .A1(\AES_ENC/us20/n602 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n866 ) );
NOR2_X2 \AES_ENC/us20/U43  ( .A1(\AES_ENC/us20/n610 ), .A2(\AES_ENC/us20/n592 ), .ZN(\AES_ENC/us20/n1006 ) );
NOR2_X2 \AES_ENC/us20/U42  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n1117 ), .ZN(\AES_ENC/us20/n1118 ) );
NOR2_X2 \AES_ENC/us20/U41  ( .A1(\AES_ENC/us20/n1119 ), .A2(\AES_ENC/us20/n1118 ), .ZN(\AES_ENC/us20/n1127 ) );
NOR2_X2 \AES_ENC/us20/U36  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n616 ), .ZN(\AES_ENC/us20/n629 ) );
NOR2_X2 \AES_ENC/us20/U35  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n906 ), .ZN(\AES_ENC/us20/n909 ) );
NOR2_X2 \AES_ENC/us20/U34  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n607 ), .ZN(\AES_ENC/us20/n658 ) );
NOR2_X2 \AES_ENC/us20/U33  ( .A1(\AES_ENC/us20/n1116 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n695 ) );
NOR2_X2 \AES_ENC/us20/U32  ( .A1(\AES_ENC/us20/n1078 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n1083 ) );
NOR2_X2 \AES_ENC/us20/U31  ( .A1(\AES_ENC/us20/n941 ), .A2(\AES_ENC/us20/n579 ), .ZN(\AES_ENC/us20/n724 ) );
NOR2_X2 \AES_ENC/us20/U30  ( .A1(\AES_ENC/us20/n611 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n1107 ) );
NOR2_X2 \AES_ENC/us20/U29  ( .A1(\AES_ENC/us20/n602 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n840 ) );
NOR2_X2 \AES_ENC/us20/U24  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n623 ), .ZN(\AES_ENC/us20/n633 ) );
NOR2_X2 \AES_ENC/us20/U23  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n1080 ), .ZN(\AES_ENC/us20/n1081 ) );
NOR2_X2 \AES_ENC/us20/U21  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n1045 ), .ZN(\AES_ENC/us20/n812 ) );
NOR2_X2 \AES_ENC/us20/U20  ( .A1(\AES_ENC/us20/n1009 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n960 ) );
NOR2_X2 \AES_ENC/us20/U19  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n619 ), .ZN(\AES_ENC/us20/n982 ) );
NOR2_X2 \AES_ENC/us20/U18  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n616 ), .ZN(\AES_ENC/us20/n757 ) );
NOR2_X2 \AES_ENC/us20/U17  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n598 ), .ZN(\AES_ENC/us20/n698 ) );
NOR2_X2 \AES_ENC/us20/U16  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n605 ), .ZN(\AES_ENC/us20/n708 ) );
NOR2_X2 \AES_ENC/us20/U15  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n603 ), .ZN(\AES_ENC/us20/n770 ) );
NOR2_X2 \AES_ENC/us20/U10  ( .A1(\AES_ENC/us20/n605 ), .A2(\AES_ENC/us20/n576 ), .ZN(\AES_ENC/us20/n803 ) );
NOR2_X2 \AES_ENC/us20/U9  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n881 ), .ZN(\AES_ENC/us20/n711 ) );
NOR2_X2 \AES_ENC/us20/U8  ( .A1(\AES_ENC/us20/n580 ), .A2(\AES_ENC/us20/n603 ), .ZN(\AES_ENC/us20/n867 ) );
NOR2_X2 \AES_ENC/us20/U7  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n615 ), .ZN(\AES_ENC/us20/n804 ) );
NOR2_X2 \AES_ENC/us20/U6  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n609 ), .ZN(\AES_ENC/us20/n1046 ) );
OR2_X4 \AES_ENC/us20/U5  ( .A1(\AES_ENC/us20/n612 ), .A2(\AES_ENC/sa20 [1]),.ZN(\AES_ENC/us20/n570 ) );
OR2_X4 \AES_ENC/us20/U4  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/sa20 [4]),.ZN(\AES_ENC/us20/n569 ) );
NAND2_X2 \AES_ENC/us20/U514  ( .A1(\AES_ENC/us20/n1121 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n1030 ) );
AND2_X2 \AES_ENC/us20/U513  ( .A1(\AES_ENC/us20/n607 ), .A2(\AES_ENC/us20/n1030 ), .ZN(\AES_ENC/us20/n1049 ) );
NAND2_X2 \AES_ENC/us20/U511  ( .A1(\AES_ENC/us20/n1049 ), .A2(\AES_ENC/us20/n794 ), .ZN(\AES_ENC/us20/n637 ) );
AND2_X2 \AES_ENC/us20/U493  ( .A1(\AES_ENC/us20/n779 ), .A2(\AES_ENC/us20/n996 ), .ZN(\AES_ENC/us20/n632 ) );
NAND4_X2 \AES_ENC/us20/U485  ( .A1(\AES_ENC/us20/n637 ), .A2(\AES_ENC/us20/n636 ), .A3(\AES_ENC/us20/n635 ), .A4(\AES_ENC/us20/n634 ), .ZN(\AES_ENC/us20/n638 ) );
NAND2_X2 \AES_ENC/us20/U484  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n638 ), .ZN(\AES_ENC/us20/n679 ) );
NAND2_X2 \AES_ENC/us20/U481  ( .A1(\AES_ENC/us20/n1094 ), .A2(\AES_ENC/us20/n613 ), .ZN(\AES_ENC/us20/n648 ) );
NAND2_X2 \AES_ENC/us20/U476  ( .A1(\AES_ENC/us20/n619 ), .A2(\AES_ENC/us20/n598 ), .ZN(\AES_ENC/us20/n762 ) );
NAND2_X2 \AES_ENC/us20/U475  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n762 ), .ZN(\AES_ENC/us20/n647 ) );
NAND4_X2 \AES_ENC/us20/U457  ( .A1(\AES_ENC/us20/n648 ), .A2(\AES_ENC/us20/n647 ), .A3(\AES_ENC/us20/n646 ), .A4(\AES_ENC/us20/n645 ), .ZN(\AES_ENC/us20/n649 ) );
NAND2_X2 \AES_ENC/us20/U456  ( .A1(\AES_ENC/sa20 [0]), .A2(\AES_ENC/us20/n649 ), .ZN(\AES_ENC/us20/n665 ) );
NAND2_X2 \AES_ENC/us20/U454  ( .A1(\AES_ENC/us20/n626 ), .A2(\AES_ENC/us20/n601 ), .ZN(\AES_ENC/us20/n855 ) );
NAND2_X2 \AES_ENC/us20/U453  ( .A1(\AES_ENC/us20/n617 ), .A2(\AES_ENC/us20/n855 ), .ZN(\AES_ENC/us20/n821 ) );
NAND2_X2 \AES_ENC/us20/U452  ( .A1(\AES_ENC/us20/n1093 ), .A2(\AES_ENC/us20/n821 ), .ZN(\AES_ENC/us20/n662 ) );
NAND2_X2 \AES_ENC/us20/U451  ( .A1(\AES_ENC/us20/n605 ), .A2(\AES_ENC/us20/n620 ), .ZN(\AES_ENC/us20/n650 ) );
NAND2_X2 \AES_ENC/us20/U450  ( .A1(\AES_ENC/us20/n956 ), .A2(\AES_ENC/us20/n650 ), .ZN(\AES_ENC/us20/n661 ) );
NAND2_X2 \AES_ENC/us20/U449  ( .A1(\AES_ENC/us20/n596 ), .A2(\AES_ENC/us20/n581 ), .ZN(\AES_ENC/us20/n839 ) );
OR2_X2 \AES_ENC/us20/U446  ( .A1(\AES_ENC/us20/n839 ), .A2(\AES_ENC/us20/n932 ), .ZN(\AES_ENC/us20/n656 ) );
NAND2_X2 \AES_ENC/us20/U445  ( .A1(\AES_ENC/us20/n624 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n1096 ) );
NAND2_X2 \AES_ENC/us20/U444  ( .A1(\AES_ENC/us20/n1030 ), .A2(\AES_ENC/us20/n1096 ), .ZN(\AES_ENC/us20/n651 ) );
NAND2_X2 \AES_ENC/us20/U443  ( .A1(\AES_ENC/us20/n1114 ), .A2(\AES_ENC/us20/n651 ), .ZN(\AES_ENC/us20/n655 ) );
OR3_X2 \AES_ENC/us20/U440  ( .A1(\AES_ENC/us20/n1079 ), .A2(\AES_ENC/sa20 [7]), .A3(\AES_ENC/us20/n596 ), .ZN(\AES_ENC/us20/n654 ));
NAND2_X2 \AES_ENC/us20/U439  ( .A1(\AES_ENC/us20/n623 ), .A2(\AES_ENC/us20/n619 ), .ZN(\AES_ENC/us20/n652 ) );
NAND4_X2 \AES_ENC/us20/U437  ( .A1(\AES_ENC/us20/n656 ), .A2(\AES_ENC/us20/n655 ), .A3(\AES_ENC/us20/n654 ), .A4(\AES_ENC/us20/n653 ), .ZN(\AES_ENC/us20/n657 ) );
NAND2_X2 \AES_ENC/us20/U436  ( .A1(\AES_ENC/sa20 [2]), .A2(\AES_ENC/us20/n657 ), .ZN(\AES_ENC/us20/n660 ) );
NAND4_X2 \AES_ENC/us20/U432  ( .A1(\AES_ENC/us20/n662 ), .A2(\AES_ENC/us20/n661 ), .A3(\AES_ENC/us20/n660 ), .A4(\AES_ENC/us20/n659 ), .ZN(\AES_ENC/us20/n663 ) );
NAND2_X2 \AES_ENC/us20/U431  ( .A1(\AES_ENC/us20/n663 ), .A2(\AES_ENC/us20/n627 ), .ZN(\AES_ENC/us20/n664 ) );
NAND2_X2 \AES_ENC/us20/U430  ( .A1(\AES_ENC/us20/n665 ), .A2(\AES_ENC/us20/n664 ), .ZN(\AES_ENC/us20/n666 ) );
NAND2_X2 \AES_ENC/us20/U429  ( .A1(\AES_ENC/sa20 [6]), .A2(\AES_ENC/us20/n666 ), .ZN(\AES_ENC/us20/n678 ) );
NAND2_X2 \AES_ENC/us20/U426  ( .A1(\AES_ENC/us20/n735 ), .A2(\AES_ENC/us20/n1093 ), .ZN(\AES_ENC/us20/n675 ) );
NAND2_X2 \AES_ENC/us20/U425  ( .A1(\AES_ENC/us20/n625 ), .A2(\AES_ENC/us20/n607 ), .ZN(\AES_ENC/us20/n1045 ) );
OR2_X2 \AES_ENC/us20/U424  ( .A1(\AES_ENC/us20/n1045 ), .A2(\AES_ENC/us20/n586 ), .ZN(\AES_ENC/us20/n674 ) );
NAND2_X2 \AES_ENC/us20/U423  ( .A1(\AES_ENC/sa20 [1]), .A2(\AES_ENC/us20/n609 ), .ZN(\AES_ENC/us20/n667 ) );
NAND2_X2 \AES_ENC/us20/U422  ( .A1(\AES_ENC/us20/n605 ), .A2(\AES_ENC/us20/n667 ), .ZN(\AES_ENC/us20/n1071 ) );
NAND4_X2 \AES_ENC/us20/U412  ( .A1(\AES_ENC/us20/n675 ), .A2(\AES_ENC/us20/n674 ), .A3(\AES_ENC/us20/n673 ), .A4(\AES_ENC/us20/n672 ), .ZN(\AES_ENC/us20/n676 ) );
NAND2_X2 \AES_ENC/us20/U411  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n676 ), .ZN(\AES_ENC/us20/n677 ) );
NAND2_X2 \AES_ENC/us20/U408  ( .A1(\AES_ENC/us20/n800 ), .A2(\AES_ENC/us20/n1022 ), .ZN(\AES_ENC/us20/n680 ) );
NAND2_X2 \AES_ENC/us20/U407  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n680 ), .ZN(\AES_ENC/us20/n681 ) );
AND2_X2 \AES_ENC/us20/U402  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n684 ), .ZN(\AES_ENC/us20/n682 ) );
NAND4_X2 \AES_ENC/us20/U395  ( .A1(\AES_ENC/us20/n691 ), .A2(\AES_ENC/us20/n583 ), .A3(\AES_ENC/us20/n690 ), .A4(\AES_ENC/us20/n689 ), .ZN(\AES_ENC/us20/n692 ) );
NAND2_X2 \AES_ENC/us20/U394  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n692 ), .ZN(\AES_ENC/us20/n733 ) );
NAND2_X2 \AES_ENC/us20/U392  ( .A1(\AES_ENC/us20/n977 ), .A2(\AES_ENC/us20/n1050 ), .ZN(\AES_ENC/us20/n702 ) );
NAND2_X2 \AES_ENC/us20/U391  ( .A1(\AES_ENC/us20/n1093 ), .A2(\AES_ENC/us20/n1045 ), .ZN(\AES_ENC/us20/n701 ) );
NAND4_X2 \AES_ENC/us20/U381  ( .A1(\AES_ENC/us20/n702 ), .A2(\AES_ENC/us20/n701 ), .A3(\AES_ENC/us20/n700 ), .A4(\AES_ENC/us20/n699 ), .ZN(\AES_ENC/us20/n703 ) );
NAND2_X2 \AES_ENC/us20/U380  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n703 ), .ZN(\AES_ENC/us20/n732 ) );
AND2_X2 \AES_ENC/us20/U379  ( .A1(\AES_ENC/sa20 [0]), .A2(\AES_ENC/sa20 [6]),.ZN(\AES_ENC/us20/n1113 ) );
NAND2_X2 \AES_ENC/us20/U378  ( .A1(\AES_ENC/us20/n619 ), .A2(\AES_ENC/us20/n1030 ), .ZN(\AES_ENC/us20/n881 ) );
NAND2_X2 \AES_ENC/us20/U377  ( .A1(\AES_ENC/us20/n1093 ), .A2(\AES_ENC/us20/n881 ), .ZN(\AES_ENC/us20/n715 ) );
NAND2_X2 \AES_ENC/us20/U376  ( .A1(\AES_ENC/us20/n1010 ), .A2(\AES_ENC/us20/n622 ), .ZN(\AES_ENC/us20/n714 ) );
NAND2_X2 \AES_ENC/us20/U375  ( .A1(\AES_ENC/us20/n855 ), .A2(\AES_ENC/us20/n625 ), .ZN(\AES_ENC/us20/n1117 ) );
XNOR2_X2 \AES_ENC/us20/U371  ( .A(\AES_ENC/us20/n593 ), .B(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n824 ) );
NAND4_X2 \AES_ENC/us20/U362  ( .A1(\AES_ENC/us20/n715 ), .A2(\AES_ENC/us20/n714 ), .A3(\AES_ENC/us20/n713 ), .A4(\AES_ENC/us20/n712 ), .ZN(\AES_ENC/us20/n716 ) );
NAND2_X2 \AES_ENC/us20/U361  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n716 ), .ZN(\AES_ENC/us20/n731 ) );
AND2_X2 \AES_ENC/us20/U360  ( .A1(\AES_ENC/sa20 [6]), .A2(\AES_ENC/us20/n627 ), .ZN(\AES_ENC/us20/n1131 ) );
NAND2_X2 \AES_ENC/us20/U359  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n717 ) );
NAND2_X2 \AES_ENC/us20/U358  ( .A1(\AES_ENC/us20/n1029 ), .A2(\AES_ENC/us20/n717 ), .ZN(\AES_ENC/us20/n728 ) );
NAND2_X2 \AES_ENC/us20/U357  ( .A1(\AES_ENC/sa20 [1]), .A2(\AES_ENC/us20/n612 ), .ZN(\AES_ENC/us20/n1097 ) );
NAND2_X2 \AES_ENC/us20/U356  ( .A1(\AES_ENC/us20/n610 ), .A2(\AES_ENC/us20/n1097 ), .ZN(\AES_ENC/us20/n718 ) );
NAND2_X2 \AES_ENC/us20/U355  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n718 ), .ZN(\AES_ENC/us20/n727 ) );
NAND4_X2 \AES_ENC/us20/U344  ( .A1(\AES_ENC/us20/n728 ), .A2(\AES_ENC/us20/n727 ), .A3(\AES_ENC/us20/n726 ), .A4(\AES_ENC/us20/n725 ), .ZN(\AES_ENC/us20/n729 ) );
NAND2_X2 \AES_ENC/us20/U343  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n729 ), .ZN(\AES_ENC/us20/n730 ) );
NAND4_X2 \AES_ENC/us20/U342  ( .A1(\AES_ENC/us20/n733 ), .A2(\AES_ENC/us20/n732 ), .A3(\AES_ENC/us20/n731 ), .A4(\AES_ENC/us20/n730 ), .ZN(\AES_ENC/sa20_sub[1] ) );
NAND2_X2 \AES_ENC/us20/U341  ( .A1(\AES_ENC/sa20 [7]), .A2(\AES_ENC/us20/n593 ), .ZN(\AES_ENC/us20/n734 ) );
NAND2_X2 \AES_ENC/us20/U340  ( .A1(\AES_ENC/us20/n734 ), .A2(\AES_ENC/us20/n588 ), .ZN(\AES_ENC/us20/n738 ) );
OR4_X2 \AES_ENC/us20/U339  ( .A1(\AES_ENC/us20/n738 ), .A2(\AES_ENC/us20/n596 ), .A3(\AES_ENC/us20/n826 ), .A4(\AES_ENC/us20/n1121 ), .ZN(\AES_ENC/us20/n746 ) );
NAND2_X2 \AES_ENC/us20/U337  ( .A1(\AES_ENC/us20/n1100 ), .A2(\AES_ENC/us20/n617 ), .ZN(\AES_ENC/us20/n992 ) );
OR2_X2 \AES_ENC/us20/U336  ( .A1(\AES_ENC/us20/n592 ), .A2(\AES_ENC/us20/n735 ), .ZN(\AES_ENC/us20/n737 ) );
NAND2_X2 \AES_ENC/us20/U334  ( .A1(\AES_ENC/us20/n605 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n753 ) );
NAND2_X2 \AES_ENC/us20/U333  ( .A1(\AES_ENC/us20/n603 ), .A2(\AES_ENC/us20/n753 ), .ZN(\AES_ENC/us20/n1080 ) );
NAND2_X2 \AES_ENC/us20/U332  ( .A1(\AES_ENC/us20/n1048 ), .A2(\AES_ENC/us20/n602 ), .ZN(\AES_ENC/us20/n736 ) );
NAND2_X2 \AES_ENC/us20/U331  ( .A1(\AES_ENC/us20/n737 ), .A2(\AES_ENC/us20/n736 ), .ZN(\AES_ENC/us20/n739 ) );
NAND2_X2 \AES_ENC/us20/U330  ( .A1(\AES_ENC/us20/n739 ), .A2(\AES_ENC/us20/n738 ), .ZN(\AES_ENC/us20/n745 ) );
NAND2_X2 \AES_ENC/us20/U326  ( .A1(\AES_ENC/us20/n1096 ), .A2(\AES_ENC/us20/n598 ), .ZN(\AES_ENC/us20/n906 ) );
NAND4_X2 \AES_ENC/us20/U323  ( .A1(\AES_ENC/us20/n746 ), .A2(\AES_ENC/us20/n992 ), .A3(\AES_ENC/us20/n745 ), .A4(\AES_ENC/us20/n744 ), .ZN(\AES_ENC/us20/n747 ) );
NAND2_X2 \AES_ENC/us20/U322  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n747 ), .ZN(\AES_ENC/us20/n793 ) );
NAND2_X2 \AES_ENC/us20/U321  ( .A1(\AES_ENC/us20/n606 ), .A2(\AES_ENC/us20/n855 ), .ZN(\AES_ENC/us20/n748 ) );
NAND2_X2 \AES_ENC/us20/U320  ( .A1(\AES_ENC/us20/n956 ), .A2(\AES_ENC/us20/n748 ), .ZN(\AES_ENC/us20/n760 ) );
NAND2_X2 \AES_ENC/us20/U313  ( .A1(\AES_ENC/us20/n598 ), .A2(\AES_ENC/us20/n753 ), .ZN(\AES_ENC/us20/n1023 ) );
NAND4_X2 \AES_ENC/us20/U308  ( .A1(\AES_ENC/us20/n760 ), .A2(\AES_ENC/us20/n992 ), .A3(\AES_ENC/us20/n759 ), .A4(\AES_ENC/us20/n758 ), .ZN(\AES_ENC/us20/n761 ) );
NAND2_X2 \AES_ENC/us20/U307  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n761 ), .ZN(\AES_ENC/us20/n792 ) );
NAND2_X2 \AES_ENC/us20/U306  ( .A1(\AES_ENC/us20/n606 ), .A2(\AES_ENC/us20/n610 ), .ZN(\AES_ENC/us20/n989 ) );
NAND2_X2 \AES_ENC/us20/U305  ( .A1(\AES_ENC/us20/n1050 ), .A2(\AES_ENC/us20/n989 ), .ZN(\AES_ENC/us20/n777 ) );
NAND2_X2 \AES_ENC/us20/U304  ( .A1(\AES_ENC/us20/n1093 ), .A2(\AES_ENC/us20/n762 ), .ZN(\AES_ENC/us20/n776 ) );
XNOR2_X2 \AES_ENC/us20/U301  ( .A(\AES_ENC/sa20 [7]), .B(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n959 ) );
NAND4_X2 \AES_ENC/us20/U289  ( .A1(\AES_ENC/us20/n777 ), .A2(\AES_ENC/us20/n776 ), .A3(\AES_ENC/us20/n775 ), .A4(\AES_ENC/us20/n774 ), .ZN(\AES_ENC/us20/n778 ) );
NAND2_X2 \AES_ENC/us20/U288  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n778 ), .ZN(\AES_ENC/us20/n791 ) );
NAND2_X2 \AES_ENC/us20/U287  ( .A1(\AES_ENC/us20/n1056 ), .A2(\AES_ENC/us20/n1050 ), .ZN(\AES_ENC/us20/n788 ) );
NAND2_X2 \AES_ENC/us20/U286  ( .A1(\AES_ENC/us20/n1091 ), .A2(\AES_ENC/us20/n779 ), .ZN(\AES_ENC/us20/n787 ) );
NAND2_X2 \AES_ENC/us20/U285  ( .A1(\AES_ENC/us20/n956 ), .A2(\AES_ENC/sa20 [1]), .ZN(\AES_ENC/us20/n786 ) );
NAND4_X2 \AES_ENC/us20/U278  ( .A1(\AES_ENC/us20/n788 ), .A2(\AES_ENC/us20/n787 ), .A3(\AES_ENC/us20/n786 ), .A4(\AES_ENC/us20/n785 ), .ZN(\AES_ENC/us20/n789 ) );
NAND2_X2 \AES_ENC/us20/U277  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n789 ), .ZN(\AES_ENC/us20/n790 ) );
NAND4_X2 \AES_ENC/us20/U276  ( .A1(\AES_ENC/us20/n793 ), .A2(\AES_ENC/us20/n792 ), .A3(\AES_ENC/us20/n791 ), .A4(\AES_ENC/us20/n790 ), .ZN(\AES_ENC/sa20_sub[2] ) );
NAND2_X2 \AES_ENC/us20/U275  ( .A1(\AES_ENC/us20/n1059 ), .A2(\AES_ENC/us20/n794 ), .ZN(\AES_ENC/us20/n810 ) );
NAND2_X2 \AES_ENC/us20/U274  ( .A1(\AES_ENC/us20/n1049 ), .A2(\AES_ENC/us20/n956 ), .ZN(\AES_ENC/us20/n809 ) );
OR2_X2 \AES_ENC/us20/U266  ( .A1(\AES_ENC/us20/n1096 ), .A2(\AES_ENC/us20/n587 ), .ZN(\AES_ENC/us20/n802 ) );
NAND2_X2 \AES_ENC/us20/U265  ( .A1(\AES_ENC/us20/n1053 ), .A2(\AES_ENC/us20/n800 ), .ZN(\AES_ENC/us20/n801 ) );
NAND2_X2 \AES_ENC/us20/U264  ( .A1(\AES_ENC/us20/n802 ), .A2(\AES_ENC/us20/n801 ), .ZN(\AES_ENC/us20/n805 ) );
NAND4_X2 \AES_ENC/us20/U261  ( .A1(\AES_ENC/us20/n810 ), .A2(\AES_ENC/us20/n809 ), .A3(\AES_ENC/us20/n808 ), .A4(\AES_ENC/us20/n807 ), .ZN(\AES_ENC/us20/n811 ) );
NAND2_X2 \AES_ENC/us20/U260  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n811 ), .ZN(\AES_ENC/us20/n852 ) );
OR2_X2 \AES_ENC/us20/U259  ( .A1(\AES_ENC/us20/n1023 ), .A2(\AES_ENC/us20/n575 ), .ZN(\AES_ENC/us20/n819 ) );
OR2_X2 \AES_ENC/us20/U257  ( .A1(\AES_ENC/us20/n570 ), .A2(\AES_ENC/us20/n930 ), .ZN(\AES_ENC/us20/n818 ) );
NAND2_X2 \AES_ENC/us20/U256  ( .A1(\AES_ENC/us20/n1013 ), .A2(\AES_ENC/us20/n1094 ), .ZN(\AES_ENC/us20/n817 ) );
NAND4_X2 \AES_ENC/us20/U249  ( .A1(\AES_ENC/us20/n819 ), .A2(\AES_ENC/us20/n818 ), .A3(\AES_ENC/us20/n817 ), .A4(\AES_ENC/us20/n816 ), .ZN(\AES_ENC/us20/n820 ) );
NAND2_X2 \AES_ENC/us20/U248  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n820 ), .ZN(\AES_ENC/us20/n851 ) );
NAND2_X2 \AES_ENC/us20/U247  ( .A1(\AES_ENC/us20/n956 ), .A2(\AES_ENC/us20/n1080 ), .ZN(\AES_ENC/us20/n835 ) );
NAND2_X2 \AES_ENC/us20/U246  ( .A1(\AES_ENC/us20/n570 ), .A2(\AES_ENC/us20/n1030 ), .ZN(\AES_ENC/us20/n1047 ) );
OR2_X2 \AES_ENC/us20/U245  ( .A1(\AES_ENC/us20/n1047 ), .A2(\AES_ENC/us20/n582 ), .ZN(\AES_ENC/us20/n834 ) );
NAND2_X2 \AES_ENC/us20/U244  ( .A1(\AES_ENC/us20/n1072 ), .A2(\AES_ENC/us20/n620 ), .ZN(\AES_ENC/us20/n833 ) );
NAND4_X2 \AES_ENC/us20/U233  ( .A1(\AES_ENC/us20/n835 ), .A2(\AES_ENC/us20/n834 ), .A3(\AES_ENC/us20/n833 ), .A4(\AES_ENC/us20/n832 ), .ZN(\AES_ENC/us20/n836 ) );
NAND2_X2 \AES_ENC/us20/U232  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n836 ), .ZN(\AES_ENC/us20/n850 ) );
NAND2_X2 \AES_ENC/us20/U231  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n601 ), .ZN(\AES_ENC/us20/n847 ) );
NAND2_X2 \AES_ENC/us20/U230  ( .A1(\AES_ENC/us20/n1050 ), .A2(\AES_ENC/us20/n1071 ), .ZN(\AES_ENC/us20/n846 ) );
OR2_X2 \AES_ENC/us20/U224  ( .A1(\AES_ENC/us20/n1053 ), .A2(\AES_ENC/us20/n911 ), .ZN(\AES_ENC/us20/n1077 ) );
NAND4_X2 \AES_ENC/us20/U220  ( .A1(\AES_ENC/us20/n847 ), .A2(\AES_ENC/us20/n846 ), .A3(\AES_ENC/us20/n845 ), .A4(\AES_ENC/us20/n844 ), .ZN(\AES_ENC/us20/n848 ) );
NAND2_X2 \AES_ENC/us20/U219  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n848 ), .ZN(\AES_ENC/us20/n849 ) );
NAND4_X2 \AES_ENC/us20/U218  ( .A1(\AES_ENC/us20/n852 ), .A2(\AES_ENC/us20/n851 ), .A3(\AES_ENC/us20/n850 ), .A4(\AES_ENC/us20/n849 ), .ZN(\AES_ENC/sa20_sub[3] ) );
NAND2_X2 \AES_ENC/us20/U216  ( .A1(\AES_ENC/us20/n1009 ), .A2(\AES_ENC/us20/n1072 ), .ZN(\AES_ENC/us20/n862 ) );
NAND2_X2 \AES_ENC/us20/U215  ( .A1(\AES_ENC/us20/n610 ), .A2(\AES_ENC/us20/n618 ), .ZN(\AES_ENC/us20/n853 ) );
NAND2_X2 \AES_ENC/us20/U214  ( .A1(\AES_ENC/us20/n1050 ), .A2(\AES_ENC/us20/n853 ), .ZN(\AES_ENC/us20/n861 ) );
NAND4_X2 \AES_ENC/us20/U206  ( .A1(\AES_ENC/us20/n862 ), .A2(\AES_ENC/us20/n861 ), .A3(\AES_ENC/us20/n860 ), .A4(\AES_ENC/us20/n859 ), .ZN(\AES_ENC/us20/n863 ) );
NAND2_X2 \AES_ENC/us20/U205  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n863 ), .ZN(\AES_ENC/us20/n905 ) );
NAND2_X2 \AES_ENC/us20/U204  ( .A1(\AES_ENC/us20/n1010 ), .A2(\AES_ENC/us20/n989 ), .ZN(\AES_ENC/us20/n874 ) );
NAND2_X2 \AES_ENC/us20/U203  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n592 ), .ZN(\AES_ENC/us20/n864 ) );
NAND2_X2 \AES_ENC/us20/U202  ( .A1(\AES_ENC/us20/n929 ), .A2(\AES_ENC/us20/n864 ), .ZN(\AES_ENC/us20/n873 ) );
NAND4_X2 \AES_ENC/us20/U193  ( .A1(\AES_ENC/us20/n874 ), .A2(\AES_ENC/us20/n873 ), .A3(\AES_ENC/us20/n872 ), .A4(\AES_ENC/us20/n871 ), .ZN(\AES_ENC/us20/n875 ) );
NAND2_X2 \AES_ENC/us20/U192  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n875 ), .ZN(\AES_ENC/us20/n904 ) );
NAND2_X2 \AES_ENC/us20/U191  ( .A1(\AES_ENC/us20/n597 ), .A2(\AES_ENC/us20/n1050 ), .ZN(\AES_ENC/us20/n889 ) );
NAND2_X2 \AES_ENC/us20/U190  ( .A1(\AES_ENC/us20/n1093 ), .A2(\AES_ENC/us20/n617 ), .ZN(\AES_ENC/us20/n876 ) );
NAND2_X2 \AES_ENC/us20/U189  ( .A1(\AES_ENC/us20/n576 ), .A2(\AES_ENC/us20/n876 ), .ZN(\AES_ENC/us20/n877 ) );
NAND2_X2 \AES_ENC/us20/U188  ( .A1(\AES_ENC/us20/n877 ), .A2(\AES_ENC/us20/n601 ), .ZN(\AES_ENC/us20/n888 ) );
NAND4_X2 \AES_ENC/us20/U179  ( .A1(\AES_ENC/us20/n889 ), .A2(\AES_ENC/us20/n888 ), .A3(\AES_ENC/us20/n887 ), .A4(\AES_ENC/us20/n886 ), .ZN(\AES_ENC/us20/n890 ) );
NAND2_X2 \AES_ENC/us20/U178  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n890 ), .ZN(\AES_ENC/us20/n903 ) );
OR2_X2 \AES_ENC/us20/U177  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n1059 ), .ZN(\AES_ENC/us20/n900 ) );
NAND2_X2 \AES_ENC/us20/U176  ( .A1(\AES_ENC/us20/n1073 ), .A2(\AES_ENC/us20/n1047 ), .ZN(\AES_ENC/us20/n899 ) );
NAND2_X2 \AES_ENC/us20/U175  ( .A1(\AES_ENC/us20/n1094 ), .A2(\AES_ENC/us20/n608 ), .ZN(\AES_ENC/us20/n898 ) );
NAND4_X2 \AES_ENC/us20/U167  ( .A1(\AES_ENC/us20/n900 ), .A2(\AES_ENC/us20/n899 ), .A3(\AES_ENC/us20/n898 ), .A4(\AES_ENC/us20/n897 ), .ZN(\AES_ENC/us20/n901 ) );
NAND2_X2 \AES_ENC/us20/U166  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n901 ), .ZN(\AES_ENC/us20/n902 ) );
NAND4_X2 \AES_ENC/us20/U165  ( .A1(\AES_ENC/us20/n905 ), .A2(\AES_ENC/us20/n904 ), .A3(\AES_ENC/us20/n903 ), .A4(\AES_ENC/us20/n902 ), .ZN(\AES_ENC/sa20_sub[4] ) );
NAND2_X2 \AES_ENC/us20/U164  ( .A1(\AES_ENC/us20/n1094 ), .A2(\AES_ENC/us20/n615 ), .ZN(\AES_ENC/us20/n922 ) );
NAND2_X2 \AES_ENC/us20/U163  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n989 ), .ZN(\AES_ENC/us20/n921 ) );
NAND4_X2 \AES_ENC/us20/U151  ( .A1(\AES_ENC/us20/n922 ), .A2(\AES_ENC/us20/n921 ), .A3(\AES_ENC/us20/n920 ), .A4(\AES_ENC/us20/n919 ), .ZN(\AES_ENC/us20/n923 ) );
NAND2_X2 \AES_ENC/us20/U150  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n923 ), .ZN(\AES_ENC/us20/n972 ) );
NAND2_X2 \AES_ENC/us20/U149  ( .A1(\AES_ENC/us20/n603 ), .A2(\AES_ENC/us20/n605 ), .ZN(\AES_ENC/us20/n924 ) );
NAND2_X2 \AES_ENC/us20/U148  ( .A1(\AES_ENC/us20/n1073 ), .A2(\AES_ENC/us20/n924 ), .ZN(\AES_ENC/us20/n939 ) );
NAND2_X2 \AES_ENC/us20/U147  ( .A1(\AES_ENC/us20/n926 ), .A2(\AES_ENC/us20/n925 ), .ZN(\AES_ENC/us20/n927 ) );
NAND2_X2 \AES_ENC/us20/U146  ( .A1(\AES_ENC/us20/n587 ), .A2(\AES_ENC/us20/n927 ), .ZN(\AES_ENC/us20/n928 ) );
NAND2_X2 \AES_ENC/us20/U145  ( .A1(\AES_ENC/us20/n928 ), .A2(\AES_ENC/us20/n1080 ), .ZN(\AES_ENC/us20/n938 ) );
OR2_X2 \AES_ENC/us20/U144  ( .A1(\AES_ENC/us20/n1117 ), .A2(\AES_ENC/us20/n580 ), .ZN(\AES_ENC/us20/n937 ) );
NAND4_X2 \AES_ENC/us20/U139  ( .A1(\AES_ENC/us20/n939 ), .A2(\AES_ENC/us20/n938 ), .A3(\AES_ENC/us20/n937 ), .A4(\AES_ENC/us20/n936 ), .ZN(\AES_ENC/us20/n940 ) );
NAND2_X2 \AES_ENC/us20/U138  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n940 ), .ZN(\AES_ENC/us20/n971 ) );
OR2_X2 \AES_ENC/us20/U137  ( .A1(\AES_ENC/us20/n586 ), .A2(\AES_ENC/us20/n941 ), .ZN(\AES_ENC/us20/n954 ) );
NAND2_X2 \AES_ENC/us20/U136  ( .A1(\AES_ENC/us20/n1096 ), .A2(\AES_ENC/us20/n618 ), .ZN(\AES_ENC/us20/n942 ) );
NAND2_X2 \AES_ENC/us20/U135  ( .A1(\AES_ENC/us20/n1048 ), .A2(\AES_ENC/us20/n942 ), .ZN(\AES_ENC/us20/n943 ) );
NAND2_X2 \AES_ENC/us20/U134  ( .A1(\AES_ENC/us20/n582 ), .A2(\AES_ENC/us20/n943 ), .ZN(\AES_ENC/us20/n944 ) );
NAND2_X2 \AES_ENC/us20/U133  ( .A1(\AES_ENC/us20/n944 ), .A2(\AES_ENC/us20/n599 ), .ZN(\AES_ENC/us20/n953 ) );
NAND4_X2 \AES_ENC/us20/U125  ( .A1(\AES_ENC/us20/n954 ), .A2(\AES_ENC/us20/n953 ), .A3(\AES_ENC/us20/n952 ), .A4(\AES_ENC/us20/n951 ), .ZN(\AES_ENC/us20/n955 ) );
NAND2_X2 \AES_ENC/us20/U124  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n955 ), .ZN(\AES_ENC/us20/n970 ) );
NAND2_X2 \AES_ENC/us20/U123  ( .A1(\AES_ENC/us20/n1094 ), .A2(\AES_ENC/us20/n1071 ), .ZN(\AES_ENC/us20/n967 ) );
NAND2_X2 \AES_ENC/us20/U122  ( .A1(\AES_ENC/us20/n956 ), .A2(\AES_ENC/us20/n1030 ), .ZN(\AES_ENC/us20/n966 ) );
NAND4_X2 \AES_ENC/us20/U114  ( .A1(\AES_ENC/us20/n967 ), .A2(\AES_ENC/us20/n966 ), .A3(\AES_ENC/us20/n965 ), .A4(\AES_ENC/us20/n964 ), .ZN(\AES_ENC/us20/n968 ) );
NAND2_X2 \AES_ENC/us20/U113  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n968 ), .ZN(\AES_ENC/us20/n969 ) );
NAND4_X2 \AES_ENC/us20/U112  ( .A1(\AES_ENC/us20/n972 ), .A2(\AES_ENC/us20/n971 ), .A3(\AES_ENC/us20/n970 ), .A4(\AES_ENC/us20/n969 ), .ZN(\AES_ENC/sa20_sub[5] ) );
NAND2_X2 \AES_ENC/us20/U111  ( .A1(\AES_ENC/us20/n570 ), .A2(\AES_ENC/us20/n1097 ), .ZN(\AES_ENC/us20/n973 ) );
NAND2_X2 \AES_ENC/us20/U110  ( .A1(\AES_ENC/us20/n1073 ), .A2(\AES_ENC/us20/n973 ), .ZN(\AES_ENC/us20/n987 ) );
NAND2_X2 \AES_ENC/us20/U109  ( .A1(\AES_ENC/us20/n974 ), .A2(\AES_ENC/us20/n1077 ), .ZN(\AES_ENC/us20/n975 ) );
NAND2_X2 \AES_ENC/us20/U108  ( .A1(\AES_ENC/us20/n584 ), .A2(\AES_ENC/us20/n975 ), .ZN(\AES_ENC/us20/n976 ) );
NAND2_X2 \AES_ENC/us20/U107  ( .A1(\AES_ENC/us20/n977 ), .A2(\AES_ENC/us20/n976 ), .ZN(\AES_ENC/us20/n986 ) );
NAND4_X2 \AES_ENC/us20/U99  ( .A1(\AES_ENC/us20/n987 ), .A2(\AES_ENC/us20/n986 ), .A3(\AES_ENC/us20/n985 ), .A4(\AES_ENC/us20/n984 ), .ZN(\AES_ENC/us20/n988 ) );
NAND2_X2 \AES_ENC/us20/U98  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n988 ), .ZN(\AES_ENC/us20/n1044 ) );
NAND2_X2 \AES_ENC/us20/U97  ( .A1(\AES_ENC/us20/n1073 ), .A2(\AES_ENC/us20/n989 ), .ZN(\AES_ENC/us20/n1004 ) );
NAND2_X2 \AES_ENC/us20/U96  ( .A1(\AES_ENC/us20/n1092 ), .A2(\AES_ENC/us20/n605 ), .ZN(\AES_ENC/us20/n1003 ) );
NAND4_X2 \AES_ENC/us20/U85  ( .A1(\AES_ENC/us20/n1004 ), .A2(\AES_ENC/us20/n1003 ), .A3(\AES_ENC/us20/n1002 ), .A4(\AES_ENC/us20/n1001 ), .ZN(\AES_ENC/us20/n1005 ) );
NAND2_X2 \AES_ENC/us20/U84  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n1005 ), .ZN(\AES_ENC/us20/n1043 ) );
NAND2_X2 \AES_ENC/us20/U83  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n626 ), .ZN(\AES_ENC/us20/n1020 ) );
NAND2_X2 \AES_ENC/us20/U82  ( .A1(\AES_ENC/us20/n1050 ), .A2(\AES_ENC/us20/n612 ), .ZN(\AES_ENC/us20/n1019 ) );
NAND2_X2 \AES_ENC/us20/U77  ( .A1(\AES_ENC/us20/n1059 ), .A2(\AES_ENC/us20/n1114 ), .ZN(\AES_ENC/us20/n1012 ) );
NAND2_X2 \AES_ENC/us20/U76  ( .A1(\AES_ENC/us20/n1010 ), .A2(\AES_ENC/us20/n604 ), .ZN(\AES_ENC/us20/n1011 ) );
NAND2_X2 \AES_ENC/us20/U75  ( .A1(\AES_ENC/us20/n1012 ), .A2(\AES_ENC/us20/n1011 ), .ZN(\AES_ENC/us20/n1016 ) );
NAND4_X2 \AES_ENC/us20/U70  ( .A1(\AES_ENC/us20/n1020 ), .A2(\AES_ENC/us20/n1019 ), .A3(\AES_ENC/us20/n1018 ), .A4(\AES_ENC/us20/n1017 ), .ZN(\AES_ENC/us20/n1021 ) );
NAND2_X2 \AES_ENC/us20/U69  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n1021 ), .ZN(\AES_ENC/us20/n1042 ) );
NAND2_X2 \AES_ENC/us20/U68  ( .A1(\AES_ENC/us20/n1022 ), .A2(\AES_ENC/us20/n1093 ), .ZN(\AES_ENC/us20/n1039 ) );
NAND2_X2 \AES_ENC/us20/U67  ( .A1(\AES_ENC/us20/n1050 ), .A2(\AES_ENC/us20/n1023 ), .ZN(\AES_ENC/us20/n1038 ) );
NAND2_X2 \AES_ENC/us20/U66  ( .A1(\AES_ENC/us20/n1024 ), .A2(\AES_ENC/us20/n1071 ), .ZN(\AES_ENC/us20/n1037 ) );
AND2_X2 \AES_ENC/us20/U60  ( .A1(\AES_ENC/us20/n1030 ), .A2(\AES_ENC/us20/n621 ), .ZN(\AES_ENC/us20/n1078 ) );
NAND4_X2 \AES_ENC/us20/U56  ( .A1(\AES_ENC/us20/n1039 ), .A2(\AES_ENC/us20/n1038 ), .A3(\AES_ENC/us20/n1037 ), .A4(\AES_ENC/us20/n1036 ), .ZN(\AES_ENC/us20/n1040 ) );
NAND2_X2 \AES_ENC/us20/U55  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n1040 ), .ZN(\AES_ENC/us20/n1041 ) );
NAND4_X2 \AES_ENC/us20/U54  ( .A1(\AES_ENC/us20/n1044 ), .A2(\AES_ENC/us20/n1043 ), .A3(\AES_ENC/us20/n1042 ), .A4(\AES_ENC/us20/n1041 ), .ZN(\AES_ENC/sa20_sub[6] ) );
NAND2_X2 \AES_ENC/us20/U53  ( .A1(\AES_ENC/us20/n1072 ), .A2(\AES_ENC/us20/n1045 ), .ZN(\AES_ENC/us20/n1068 ) );
NAND2_X2 \AES_ENC/us20/U52  ( .A1(\AES_ENC/us20/n1046 ), .A2(\AES_ENC/us20/n603 ), .ZN(\AES_ENC/us20/n1067 ) );
NAND2_X2 \AES_ENC/us20/U51  ( .A1(\AES_ENC/us20/n1094 ), .A2(\AES_ENC/us20/n1047 ), .ZN(\AES_ENC/us20/n1066 ) );
NAND4_X2 \AES_ENC/us20/U40  ( .A1(\AES_ENC/us20/n1068 ), .A2(\AES_ENC/us20/n1067 ), .A3(\AES_ENC/us20/n1066 ), .A4(\AES_ENC/us20/n1065 ), .ZN(\AES_ENC/us20/n1069 ) );
NAND2_X2 \AES_ENC/us20/U39  ( .A1(\AES_ENC/us20/n1070 ), .A2(\AES_ENC/us20/n1069 ), .ZN(\AES_ENC/us20/n1135 ) );
NAND2_X2 \AES_ENC/us20/U38  ( .A1(\AES_ENC/us20/n1072 ), .A2(\AES_ENC/us20/n1071 ), .ZN(\AES_ENC/us20/n1088 ) );
NAND2_X2 \AES_ENC/us20/U37  ( .A1(\AES_ENC/us20/n1073 ), .A2(\AES_ENC/us20/n608 ), .ZN(\AES_ENC/us20/n1087 ) );
NAND4_X2 \AES_ENC/us20/U28  ( .A1(\AES_ENC/us20/n1088 ), .A2(\AES_ENC/us20/n1087 ), .A3(\AES_ENC/us20/n1086 ), .A4(\AES_ENC/us20/n1085 ), .ZN(\AES_ENC/us20/n1089 ) );
NAND2_X2 \AES_ENC/us20/U27  ( .A1(\AES_ENC/us20/n1090 ), .A2(\AES_ENC/us20/n1089 ), .ZN(\AES_ENC/us20/n1134 ) );
NAND2_X2 \AES_ENC/us20/U26  ( .A1(\AES_ENC/us20/n1091 ), .A2(\AES_ENC/us20/n1093 ), .ZN(\AES_ENC/us20/n1111 ) );
NAND2_X2 \AES_ENC/us20/U25  ( .A1(\AES_ENC/us20/n1092 ), .A2(\AES_ENC/us20/n1120 ), .ZN(\AES_ENC/us20/n1110 ) );
AND2_X2 \AES_ENC/us20/U22  ( .A1(\AES_ENC/us20/n1097 ), .A2(\AES_ENC/us20/n1096 ), .ZN(\AES_ENC/us20/n1098 ) );
NAND4_X2 \AES_ENC/us20/U14  ( .A1(\AES_ENC/us20/n1111 ), .A2(\AES_ENC/us20/n1110 ), .A3(\AES_ENC/us20/n1109 ), .A4(\AES_ENC/us20/n1108 ), .ZN(\AES_ENC/us20/n1112 ) );
NAND2_X2 \AES_ENC/us20/U13  ( .A1(\AES_ENC/us20/n1113 ), .A2(\AES_ENC/us20/n1112 ), .ZN(\AES_ENC/us20/n1133 ) );
NAND2_X2 \AES_ENC/us20/U12  ( .A1(\AES_ENC/us20/n1115 ), .A2(\AES_ENC/us20/n1114 ), .ZN(\AES_ENC/us20/n1129 ) );
OR2_X2 \AES_ENC/us20/U11  ( .A1(\AES_ENC/us20/n579 ), .A2(\AES_ENC/us20/n1116 ), .ZN(\AES_ENC/us20/n1128 ) );
NAND4_X2 \AES_ENC/us20/U3  ( .A1(\AES_ENC/us20/n1129 ), .A2(\AES_ENC/us20/n1128 ), .A3(\AES_ENC/us20/n1127 ), .A4(\AES_ENC/us20/n1126 ), .ZN(\AES_ENC/us20/n1130 ) );
NAND2_X2 \AES_ENC/us20/U2  ( .A1(\AES_ENC/us20/n1131 ), .A2(\AES_ENC/us20/n1130 ), .ZN(\AES_ENC/us20/n1132 ) );
NAND4_X2 \AES_ENC/us20/U1  ( .A1(\AES_ENC/us20/n1135 ), .A2(\AES_ENC/us20/n1134 ), .A3(\AES_ENC/us20/n1133 ), .A4(\AES_ENC/us20/n1132 ), .ZN(\AES_ENC/sa20_sub[7] ) );
INV_X4 \AES_ENC/us21/U575  ( .A(\AES_ENC/sa21 [0]), .ZN(\AES_ENC/us21/n627 ));
INV_X4 \AES_ENC/us21/U574  ( .A(\AES_ENC/us21/n1053 ), .ZN(\AES_ENC/us21/n625 ) );
INV_X4 \AES_ENC/us21/U573  ( .A(\AES_ENC/us21/n1103 ), .ZN(\AES_ENC/us21/n623 ) );
INV_X4 \AES_ENC/us21/U572  ( .A(\AES_ENC/us21/n1056 ), .ZN(\AES_ENC/us21/n622 ) );
INV_X4 \AES_ENC/us21/U571  ( .A(\AES_ENC/us21/n1102 ), .ZN(\AES_ENC/us21/n621 ) );
INV_X4 \AES_ENC/us21/U570  ( .A(\AES_ENC/us21/n1074 ), .ZN(\AES_ENC/us21/n620 ) );
INV_X4 \AES_ENC/us21/U569  ( .A(\AES_ENC/us21/n929 ), .ZN(\AES_ENC/us21/n619 ) );
INV_X4 \AES_ENC/us21/U568  ( .A(\AES_ENC/us21/n1091 ), .ZN(\AES_ENC/us21/n618 ) );
INV_X4 \AES_ENC/us21/U567  ( .A(\AES_ENC/us21/n826 ), .ZN(\AES_ENC/us21/n617 ) );
INV_X4 \AES_ENC/us21/U566  ( .A(\AES_ENC/us21/n1031 ), .ZN(\AES_ENC/us21/n616 ) );
INV_X4 \AES_ENC/us21/U565  ( .A(\AES_ENC/us21/n1054 ), .ZN(\AES_ENC/us21/n615 ) );
INV_X4 \AES_ENC/us21/U564  ( .A(\AES_ENC/us21/n1025 ), .ZN(\AES_ENC/us21/n614 ) );
INV_X4 \AES_ENC/us21/U563  ( .A(\AES_ENC/us21/n990 ), .ZN(\AES_ENC/us21/n613 ) );
INV_X4 \AES_ENC/us21/U562  ( .A(\AES_ENC/sa21 [4]), .ZN(\AES_ENC/us21/n612 ));
INV_X4 \AES_ENC/us21/U561  ( .A(\AES_ENC/us21/n881 ), .ZN(\AES_ENC/us21/n611 ) );
INV_X4 \AES_ENC/us21/U560  ( .A(\AES_ENC/us21/n1022 ), .ZN(\AES_ENC/us21/n610 ) );
INV_X4 \AES_ENC/us21/U559  ( .A(\AES_ENC/us21/n1120 ), .ZN(\AES_ENC/us21/n609 ) );
INV_X4 \AES_ENC/us21/U558  ( .A(\AES_ENC/us21/n977 ), .ZN(\AES_ENC/us21/n608 ) );
INV_X4 \AES_ENC/us21/U557  ( .A(\AES_ENC/us21/n926 ), .ZN(\AES_ENC/us21/n607 ) );
INV_X4 \AES_ENC/us21/U556  ( .A(\AES_ENC/us21/n910 ), .ZN(\AES_ENC/us21/n606 ) );
INV_X4 \AES_ENC/us21/U555  ( .A(\AES_ENC/us21/n1121 ), .ZN(\AES_ENC/us21/n605 ) );
INV_X4 \AES_ENC/us21/U554  ( .A(\AES_ENC/us21/n1009 ), .ZN(\AES_ENC/us21/n604 ) );
INV_X4 \AES_ENC/us21/U553  ( .A(\AES_ENC/us21/n1080 ), .ZN(\AES_ENC/us21/n602 ) );
INV_X4 \AES_ENC/us21/U552  ( .A(\AES_ENC/us21/n821 ), .ZN(\AES_ENC/us21/n600 ) );
INV_X4 \AES_ENC/us21/U551  ( .A(\AES_ENC/us21/n1013 ), .ZN(\AES_ENC/us21/n599 ) );
INV_X4 \AES_ENC/us21/U550  ( .A(\AES_ENC/us21/n1058 ), .ZN(\AES_ENC/us21/n598 ) );
INV_X4 \AES_ENC/us21/U549  ( .A(\AES_ENC/us21/n906 ), .ZN(\AES_ENC/us21/n597 ) );
INV_X4 \AES_ENC/us21/U548  ( .A(\AES_ENC/us21/n959 ), .ZN(\AES_ENC/us21/n596 ) );
INV_X4 \AES_ENC/us21/U547  ( .A(\AES_ENC/sa21 [7]), .ZN(\AES_ENC/us21/n595 ));
INV_X4 \AES_ENC/us21/U546  ( .A(\AES_ENC/us21/n1114 ), .ZN(\AES_ENC/us21/n593 ) );
INV_X4 \AES_ENC/us21/U545  ( .A(\AES_ENC/us21/n1048 ), .ZN(\AES_ENC/us21/n592 ) );
INV_X4 \AES_ENC/us21/U544  ( .A(\AES_ENC/us21/n974 ), .ZN(\AES_ENC/us21/n590 ) );
INV_X4 \AES_ENC/us21/U543  ( .A(\AES_ENC/us21/n794 ), .ZN(\AES_ENC/us21/n588 ) );
INV_X4 \AES_ENC/us21/U542  ( .A(\AES_ENC/us21/n880 ), .ZN(\AES_ENC/us21/n586 ) );
INV_X4 \AES_ENC/us21/U541  ( .A(\AES_ENC/sa21 [2]), .ZN(\AES_ENC/us21/n584 ));
INV_X4 \AES_ENC/us21/U540  ( .A(\AES_ENC/us21/n800 ), .ZN(\AES_ENC/us21/n583 ) );
INV_X4 \AES_ENC/us21/U539  ( .A(\AES_ENC/us21/n925 ), .ZN(\AES_ENC/us21/n582 ) );
INV_X4 \AES_ENC/us21/U538  ( .A(\AES_ENC/us21/n992 ), .ZN(\AES_ENC/us21/n580 ) );
INV_X4 \AES_ENC/us21/U537  ( .A(\AES_ENC/us21/n779 ), .ZN(\AES_ENC/us21/n579 ) );
INV_X4 \AES_ENC/us21/U536  ( .A(\AES_ENC/us21/n1092 ), .ZN(\AES_ENC/us21/n575 ) );
INV_X4 \AES_ENC/us21/U535  ( .A(\AES_ENC/us21/n824 ), .ZN(\AES_ENC/us21/n574 ) );
NOR2_X2 \AES_ENC/us21/U534  ( .A1(\AES_ENC/sa21 [0]), .A2(\AES_ENC/sa21 [6]),.ZN(\AES_ENC/us21/n1090 ) );
NOR2_X2 \AES_ENC/us21/U533  ( .A1(\AES_ENC/us21/n627 ), .A2(\AES_ENC/sa21 [6]), .ZN(\AES_ENC/us21/n1070 ) );
NOR2_X2 \AES_ENC/us21/U532  ( .A1(\AES_ENC/sa21 [4]), .A2(\AES_ENC/sa21 [3]),.ZN(\AES_ENC/us21/n1025 ) );
INV_X4 \AES_ENC/us21/U531  ( .A(\AES_ENC/us21/n569 ), .ZN(\AES_ENC/us21/n572 ) );
NOR2_X2 \AES_ENC/us21/U530  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n765 ) );
NOR2_X2 \AES_ENC/us21/U529  ( .A1(\AES_ENC/sa21 [4]), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n764 ) );
NOR2_X2 \AES_ENC/us21/U528  ( .A1(\AES_ENC/us21/n765 ), .A2(\AES_ENC/us21/n764 ), .ZN(\AES_ENC/us21/n766 ) );
NOR2_X2 \AES_ENC/us21/U527  ( .A1(\AES_ENC/us21/n766 ), .A2(\AES_ENC/us21/n596 ), .ZN(\AES_ENC/us21/n767 ) );
NOR3_X2 \AES_ENC/us21/U526  ( .A1(\AES_ENC/us21/n595 ), .A2(\AES_ENC/sa21 [5]), .A3(\AES_ENC/us21/n704 ), .ZN(\AES_ENC/us21/n706 ));
NOR2_X2 \AES_ENC/us21/U525  ( .A1(\AES_ENC/us21/n1117 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n707 ) );
NOR2_X2 \AES_ENC/us21/U524  ( .A1(\AES_ENC/sa21 [4]), .A2(\AES_ENC/us21/n575 ), .ZN(\AES_ENC/us21/n705 ) );
NOR3_X2 \AES_ENC/us21/U523  ( .A1(\AES_ENC/us21/n707 ), .A2(\AES_ENC/us21/n706 ), .A3(\AES_ENC/us21/n705 ), .ZN(\AES_ENC/us21/n713 ) );
INV_X4 \AES_ENC/us21/U522  ( .A(\AES_ENC/sa21 [3]), .ZN(\AES_ENC/us21/n624 ));
NAND3_X2 \AES_ENC/us21/U521  ( .A1(\AES_ENC/us21/n652 ), .A2(\AES_ENC/us21/n594 ), .A3(\AES_ENC/sa21 [7]), .ZN(\AES_ENC/us21/n653 ));
NOR2_X2 \AES_ENC/us21/U520  ( .A1(\AES_ENC/us21/n584 ), .A2(\AES_ENC/sa21 [5]), .ZN(\AES_ENC/us21/n925 ) );
NOR2_X2 \AES_ENC/us21/U519  ( .A1(\AES_ENC/sa21 [5]), .A2(\AES_ENC/sa21 [2]),.ZN(\AES_ENC/us21/n974 ) );
INV_X4 \AES_ENC/us21/U518  ( .A(\AES_ENC/sa21 [5]), .ZN(\AES_ENC/us21/n594 ));
NOR2_X2 \AES_ENC/us21/U517  ( .A1(\AES_ENC/us21/n584 ), .A2(\AES_ENC/sa21 [7]), .ZN(\AES_ENC/us21/n779 ) );
NAND3_X2 \AES_ENC/us21/U516  ( .A1(\AES_ENC/us21/n679 ), .A2(\AES_ENC/us21/n678 ), .A3(\AES_ENC/us21/n677 ), .ZN(\AES_ENC/sa21_sub[0] ) );
NOR2_X2 \AES_ENC/us21/U515  ( .A1(\AES_ENC/us21/n594 ), .A2(\AES_ENC/sa21 [2]), .ZN(\AES_ENC/us21/n1048 ) );
NOR4_X2 \AES_ENC/us21/U512  ( .A1(\AES_ENC/us21/n633 ), .A2(\AES_ENC/us21/n632 ), .A3(\AES_ENC/us21/n631 ), .A4(\AES_ENC/us21/n630 ), .ZN(\AES_ENC/us21/n634 ) );
NOR2_X2 \AES_ENC/us21/U510  ( .A1(\AES_ENC/us21/n629 ), .A2(\AES_ENC/us21/n628 ), .ZN(\AES_ENC/us21/n635 ) );
NAND3_X2 \AES_ENC/us21/U509  ( .A1(\AES_ENC/sa21 [2]), .A2(\AES_ENC/sa21 [7]), .A3(\AES_ENC/us21/n1059 ), .ZN(\AES_ENC/us21/n636 ) );
NOR2_X2 \AES_ENC/us21/U508  ( .A1(\AES_ENC/sa21 [7]), .A2(\AES_ENC/sa21 [2]),.ZN(\AES_ENC/us21/n794 ) );
NOR2_X2 \AES_ENC/us21/U507  ( .A1(\AES_ENC/sa21 [4]), .A2(\AES_ENC/sa21 [1]),.ZN(\AES_ENC/us21/n1102 ) );
NOR2_X2 \AES_ENC/us21/U506  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/sa21 [3]), .ZN(\AES_ENC/us21/n1053 ) );
NOR2_X2 \AES_ENC/us21/U505  ( .A1(\AES_ENC/us21/n579 ), .A2(\AES_ENC/sa21 [5]), .ZN(\AES_ENC/us21/n1024 ) );
NOR2_X2 \AES_ENC/us21/U504  ( .A1(\AES_ENC/us21/n593 ), .A2(\AES_ENC/sa21 [2]), .ZN(\AES_ENC/us21/n1093 ) );
NOR2_X2 \AES_ENC/us21/U503  ( .A1(\AES_ENC/us21/n588 ), .A2(\AES_ENC/sa21 [5]), .ZN(\AES_ENC/us21/n1094 ) );
NOR2_X2 \AES_ENC/us21/U502  ( .A1(\AES_ENC/us21/n612 ), .A2(\AES_ENC/sa21 [3]), .ZN(\AES_ENC/us21/n931 ) );
INV_X4 \AES_ENC/us21/U501  ( .A(\AES_ENC/us21/n570 ), .ZN(\AES_ENC/us21/n573 ) );
NOR2_X2 \AES_ENC/us21/U500  ( .A1(\AES_ENC/us21/n1053 ), .A2(\AES_ENC/us21/n1095 ), .ZN(\AES_ENC/us21/n639 ) );
NOR3_X2 \AES_ENC/us21/U499  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n573 ), .A3(\AES_ENC/us21/n1074 ), .ZN(\AES_ENC/us21/n641 ) );
NOR2_X2 \AES_ENC/us21/U498  ( .A1(\AES_ENC/us21/n639 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n640 ) );
NOR2_X2 \AES_ENC/us21/U497  ( .A1(\AES_ENC/us21/n641 ), .A2(\AES_ENC/us21/n640 ), .ZN(\AES_ENC/us21/n646 ) );
NOR3_X2 \AES_ENC/us21/U496  ( .A1(\AES_ENC/us21/n995 ), .A2(\AES_ENC/us21/n580 ), .A3(\AES_ENC/us21/n994 ), .ZN(\AES_ENC/us21/n1002 ) );
NOR2_X2 \AES_ENC/us21/U495  ( .A1(\AES_ENC/us21/n909 ), .A2(\AES_ENC/us21/n908 ), .ZN(\AES_ENC/us21/n920 ) );
NOR2_X2 \AES_ENC/us21/U494  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n823 ) );
NOR2_X2 \AES_ENC/us21/U492  ( .A1(\AES_ENC/us21/n612 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n822 ) );
NOR2_X2 \AES_ENC/us21/U491  ( .A1(\AES_ENC/us21/n823 ), .A2(\AES_ENC/us21/n822 ), .ZN(\AES_ENC/us21/n825 ) );
NOR2_X2 \AES_ENC/us21/U490  ( .A1(\AES_ENC/sa21 [1]), .A2(\AES_ENC/us21/n601 ), .ZN(\AES_ENC/us21/n913 ) );
NOR2_X2 \AES_ENC/us21/U489  ( .A1(\AES_ENC/us21/n913 ), .A2(\AES_ENC/us21/n1091 ), .ZN(\AES_ENC/us21/n914 ) );
NOR2_X2 \AES_ENC/us21/U488  ( .A1(\AES_ENC/us21/n826 ), .A2(\AES_ENC/us21/n572 ), .ZN(\AES_ENC/us21/n827 ) );
NOR3_X2 \AES_ENC/us21/U487  ( .A1(\AES_ENC/us21/n769 ), .A2(\AES_ENC/us21/n768 ), .A3(\AES_ENC/us21/n767 ), .ZN(\AES_ENC/us21/n775 ) );
NOR2_X2 \AES_ENC/us21/U486  ( .A1(\AES_ENC/us21/n1056 ), .A2(\AES_ENC/us21/n1053 ), .ZN(\AES_ENC/us21/n749 ) );
NOR2_X2 \AES_ENC/us21/U483  ( .A1(\AES_ENC/us21/n749 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n752 ) );
INV_X4 \AES_ENC/us21/U482  ( .A(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n626 ));
NOR2_X2 \AES_ENC/us21/U480  ( .A1(\AES_ENC/us21/n1054 ), .A2(\AES_ENC/us21/n1053 ), .ZN(\AES_ENC/us21/n1055 ) );
OR2_X4 \AES_ENC/us21/U479  ( .A1(\AES_ENC/us21/n1094 ), .A2(\AES_ENC/us21/n1093 ), .ZN(\AES_ENC/us21/n571 ) );
AND2_X2 \AES_ENC/us21/U478  ( .A1(\AES_ENC/us21/n571 ), .A2(\AES_ENC/us21/n1095 ), .ZN(\AES_ENC/us21/n1101 ) );
NOR2_X2 \AES_ENC/us21/U477  ( .A1(\AES_ENC/us21/n1074 ), .A2(\AES_ENC/us21/n931 ), .ZN(\AES_ENC/us21/n796 ) );
NOR2_X2 \AES_ENC/us21/U474  ( .A1(\AES_ENC/us21/n796 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n797 ) );
NOR2_X2 \AES_ENC/us21/U473  ( .A1(\AES_ENC/us21/n932 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n933 ) );
NOR2_X2 \AES_ENC/us21/U472  ( .A1(\AES_ENC/us21/n929 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n935 ) );
NOR2_X2 \AES_ENC/us21/U471  ( .A1(\AES_ENC/us21/n931 ), .A2(\AES_ENC/us21/n930 ), .ZN(\AES_ENC/us21/n934 ) );
NOR3_X2 \AES_ENC/us21/U470  ( .A1(\AES_ENC/us21/n935 ), .A2(\AES_ENC/us21/n934 ), .A3(\AES_ENC/us21/n933 ), .ZN(\AES_ENC/us21/n936 ) );
NOR2_X2 \AES_ENC/us21/U469  ( .A1(\AES_ENC/us21/n612 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n1075 ) );
NOR2_X2 \AES_ENC/us21/U468  ( .A1(\AES_ENC/us21/n572 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n949 ) );
NOR2_X2 \AES_ENC/us21/U467  ( .A1(\AES_ENC/us21/n1049 ), .A2(\AES_ENC/us21/n592 ), .ZN(\AES_ENC/us21/n1051 ) );
NOR2_X2 \AES_ENC/us21/U466  ( .A1(\AES_ENC/us21/n1051 ), .A2(\AES_ENC/us21/n1050 ), .ZN(\AES_ENC/us21/n1052 ) );
NOR2_X2 \AES_ENC/us21/U465  ( .A1(\AES_ENC/us21/n1052 ), .A2(\AES_ENC/us21/n604 ), .ZN(\AES_ENC/us21/n1064 ) );
NOR2_X2 \AES_ENC/us21/U464  ( .A1(\AES_ENC/sa21 [1]), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n631 ) );
NOR2_X2 \AES_ENC/us21/U463  ( .A1(\AES_ENC/us21/n1025 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n980 ) );
NOR2_X2 \AES_ENC/us21/U462  ( .A1(\AES_ENC/us21/n1073 ), .A2(\AES_ENC/us21/n1094 ), .ZN(\AES_ENC/us21/n795 ) );
NOR2_X2 \AES_ENC/us21/U461  ( .A1(\AES_ENC/us21/n795 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n799 ) );
NOR2_X2 \AES_ENC/us21/U460  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n981 ) );
NOR2_X2 \AES_ENC/us21/U459  ( .A1(\AES_ENC/us21/n1102 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n643 ) );
NOR2_X2 \AES_ENC/us21/U458  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n624 ), .ZN(\AES_ENC/us21/n642 ) );
NOR2_X2 \AES_ENC/us21/U455  ( .A1(\AES_ENC/us21/n911 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n644 ) );
NOR4_X2 \AES_ENC/us21/U448  ( .A1(\AES_ENC/us21/n644 ), .A2(\AES_ENC/us21/n643 ), .A3(\AES_ENC/us21/n804 ), .A4(\AES_ENC/us21/n642 ), .ZN(\AES_ENC/us21/n645 ) );
NOR2_X2 \AES_ENC/us21/U447  ( .A1(\AES_ENC/us21/n1102 ), .A2(\AES_ENC/us21/n910 ), .ZN(\AES_ENC/us21/n932 ) );
NOR2_X2 \AES_ENC/us21/U442  ( .A1(\AES_ENC/us21/n1102 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n755 ) );
NOR2_X2 \AES_ENC/us21/U441  ( .A1(\AES_ENC/us21/n931 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n743 ) );
NOR2_X2 \AES_ENC/us21/U438  ( .A1(\AES_ENC/us21/n1072 ), .A2(\AES_ENC/us21/n1094 ), .ZN(\AES_ENC/us21/n930 ) );
NOR2_X2 \AES_ENC/us21/U435  ( .A1(\AES_ENC/us21/n1074 ), .A2(\AES_ENC/us21/n1025 ), .ZN(\AES_ENC/us21/n891 ) );
NOR2_X2 \AES_ENC/us21/U434  ( .A1(\AES_ENC/us21/n891 ), .A2(\AES_ENC/us21/n582 ), .ZN(\AES_ENC/us21/n894 ) );
NOR3_X2 \AES_ENC/us21/U433  ( .A1(\AES_ENC/us21/n601 ), .A2(\AES_ENC/sa21 [1]), .A3(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n683 ));
INV_X4 \AES_ENC/us21/U428  ( .A(\AES_ENC/us21/n931 ), .ZN(\AES_ENC/us21/n601 ) );
NOR2_X2 \AES_ENC/us21/U427  ( .A1(\AES_ENC/us21/n996 ), .A2(\AES_ENC/us21/n931 ), .ZN(\AES_ENC/us21/n704 ) );
NOR2_X2 \AES_ENC/us21/U421  ( .A1(\AES_ENC/us21/n931 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n685 ) );
NOR2_X2 \AES_ENC/us21/U420  ( .A1(\AES_ENC/us21/n1029 ), .A2(\AES_ENC/us21/n1025 ), .ZN(\AES_ENC/us21/n1079 ) );
NOR3_X2 \AES_ENC/us21/U419  ( .A1(\AES_ENC/us21/n620 ), .A2(\AES_ENC/us21/n1025 ), .A3(\AES_ENC/us21/n590 ), .ZN(\AES_ENC/us21/n945 ) );
NOR2_X2 \AES_ENC/us21/U418  ( .A1(\AES_ENC/us21/n594 ), .A2(\AES_ENC/us21/n584 ), .ZN(\AES_ENC/us21/n800 ) );
NOR3_X2 \AES_ENC/us21/U417  ( .A1(\AES_ENC/us21/n598 ), .A2(\AES_ENC/us21/n595 ), .A3(\AES_ENC/us21/n584 ), .ZN(\AES_ENC/us21/n798 ) );
NOR3_X2 \AES_ENC/us21/U416  ( .A1(\AES_ENC/us21/n583 ), .A2(\AES_ENC/us21/n572 ), .A3(\AES_ENC/us21/n596 ), .ZN(\AES_ENC/us21/n962 ) );
NOR3_X2 \AES_ENC/us21/U415  ( .A1(\AES_ENC/us21/n959 ), .A2(\AES_ENC/us21/n572 ), .A3(\AES_ENC/us21/n582 ), .ZN(\AES_ENC/us21/n768 ) );
NOR3_X2 \AES_ENC/us21/U414  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n572 ), .A3(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n694 ) );
NOR3_X2 \AES_ENC/us21/U413  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n572 ), .A3(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n895 ) );
NOR3_X2 \AES_ENC/us21/U410  ( .A1(\AES_ENC/us21/n1008 ), .A2(\AES_ENC/us21/n1007 ), .A3(\AES_ENC/us21/n1006 ), .ZN(\AES_ENC/us21/n1018 ) );
NOR4_X2 \AES_ENC/us21/U409  ( .A1(\AES_ENC/us21/n806 ), .A2(\AES_ENC/us21/n805 ), .A3(\AES_ENC/us21/n804 ), .A4(\AES_ENC/us21/n803 ), .ZN(\AES_ENC/us21/n807 ) );
NOR3_X2 \AES_ENC/us21/U406  ( .A1(\AES_ENC/us21/n799 ), .A2(\AES_ENC/us21/n798 ), .A3(\AES_ENC/us21/n797 ), .ZN(\AES_ENC/us21/n808 ) );
NOR4_X2 \AES_ENC/us21/U405  ( .A1(\AES_ENC/us21/n843 ), .A2(\AES_ENC/us21/n842 ), .A3(\AES_ENC/us21/n841 ), .A4(\AES_ENC/us21/n840 ), .ZN(\AES_ENC/us21/n844 ) );
NOR2_X2 \AES_ENC/us21/U404  ( .A1(\AES_ENC/us21/n669 ), .A2(\AES_ENC/us21/n668 ), .ZN(\AES_ENC/us21/n673 ) );
NOR4_X2 \AES_ENC/us21/U403  ( .A1(\AES_ENC/us21/n946 ), .A2(\AES_ENC/us21/n1046 ), .A3(\AES_ENC/us21/n671 ), .A4(\AES_ENC/us21/n670 ), .ZN(\AES_ENC/us21/n672 ) );
NOR4_X2 \AES_ENC/us21/U401  ( .A1(\AES_ENC/us21/n711 ), .A2(\AES_ENC/us21/n710 ), .A3(\AES_ENC/us21/n709 ), .A4(\AES_ENC/us21/n708 ), .ZN(\AES_ENC/us21/n712 ) );
NOR4_X2 \AES_ENC/us21/U400  ( .A1(\AES_ENC/us21/n963 ), .A2(\AES_ENC/us21/n962 ), .A3(\AES_ENC/us21/n961 ), .A4(\AES_ENC/us21/n960 ), .ZN(\AES_ENC/us21/n964 ) );
NOR3_X2 \AES_ENC/us21/U399  ( .A1(\AES_ENC/us21/n1101 ), .A2(\AES_ENC/us21/n1100 ), .A3(\AES_ENC/us21/n1099 ), .ZN(\AES_ENC/us21/n1109 ) );
NOR3_X2 \AES_ENC/us21/U398  ( .A1(\AES_ENC/us21/n743 ), .A2(\AES_ENC/us21/n742 ), .A3(\AES_ENC/us21/n741 ), .ZN(\AES_ENC/us21/n744 ) );
NOR2_X2 \AES_ENC/us21/U397  ( .A1(\AES_ENC/us21/n697 ), .A2(\AES_ENC/us21/n658 ), .ZN(\AES_ENC/us21/n659 ) );
NOR2_X2 \AES_ENC/us21/U396  ( .A1(\AES_ENC/us21/n1078 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n1033 ) );
NOR2_X2 \AES_ENC/us21/U393  ( .A1(\AES_ENC/us21/n1031 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n1032 ) );
NOR3_X2 \AES_ENC/us21/U390  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n1025 ), .A3(\AES_ENC/us21/n1074 ), .ZN(\AES_ENC/us21/n1035 ) );
NOR4_X2 \AES_ENC/us21/U389  ( .A1(\AES_ENC/us21/n1035 ), .A2(\AES_ENC/us21/n1034 ), .A3(\AES_ENC/us21/n1033 ), .A4(\AES_ENC/us21/n1032 ), .ZN(\AES_ENC/us21/n1036 ) );
NOR2_X2 \AES_ENC/us21/U388  ( .A1(\AES_ENC/us21/n611 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n885 ) );
NOR2_X2 \AES_ENC/us21/U387  ( .A1(\AES_ENC/us21/n601 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n882 ) );
NOR2_X2 \AES_ENC/us21/U386  ( .A1(\AES_ENC/us21/n1053 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n884 ) );
NOR4_X2 \AES_ENC/us21/U385  ( .A1(\AES_ENC/us21/n885 ), .A2(\AES_ENC/us21/n884 ), .A3(\AES_ENC/us21/n883 ), .A4(\AES_ENC/us21/n882 ), .ZN(\AES_ENC/us21/n886 ) );
NOR2_X2 \AES_ENC/us21/U384  ( .A1(\AES_ENC/us21/n825 ), .A2(\AES_ENC/us21/n574 ), .ZN(\AES_ENC/us21/n830 ) );
NOR2_X2 \AES_ENC/us21/U383  ( .A1(\AES_ENC/us21/n827 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n829 ) );
NOR2_X2 \AES_ENC/us21/U382  ( .A1(\AES_ENC/us21/n572 ), .A2(\AES_ENC/us21/n575 ), .ZN(\AES_ENC/us21/n828 ) );
NOR4_X2 \AES_ENC/us21/U374  ( .A1(\AES_ENC/us21/n831 ), .A2(\AES_ENC/us21/n830 ), .A3(\AES_ENC/us21/n829 ), .A4(\AES_ENC/us21/n828 ), .ZN(\AES_ENC/us21/n832 ) );
NOR2_X2 \AES_ENC/us21/U373  ( .A1(\AES_ENC/us21/n578 ), .A2(\AES_ENC/us21/n603 ), .ZN(\AES_ENC/us21/n1104 ) );
NOR2_X2 \AES_ENC/us21/U372  ( .A1(\AES_ENC/us21/n1102 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n1106 ) );
NOR2_X2 \AES_ENC/us21/U370  ( .A1(\AES_ENC/us21/n1103 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n1105 ) );
NOR4_X2 \AES_ENC/us21/U369  ( .A1(\AES_ENC/us21/n1107 ), .A2(\AES_ENC/us21/n1106 ), .A3(\AES_ENC/us21/n1105 ), .A4(\AES_ENC/us21/n1104 ), .ZN(\AES_ENC/us21/n1108 ) );
NOR3_X2 \AES_ENC/us21/U368  ( .A1(\AES_ENC/us21/n959 ), .A2(\AES_ENC/us21/n624 ), .A3(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n963 ) );
NOR2_X2 \AES_ENC/us21/U367  ( .A1(\AES_ENC/us21/n594 ), .A2(\AES_ENC/us21/n595 ), .ZN(\AES_ENC/us21/n1114 ) );
INV_X4 \AES_ENC/us21/U366  ( .A(\AES_ENC/us21/n1024 ), .ZN(\AES_ENC/us21/n578 ) );
NOR3_X2 \AES_ENC/us21/U365  ( .A1(\AES_ENC/us21/n910 ), .A2(\AES_ENC/us21/n1059 ), .A3(\AES_ENC/us21/n584 ), .ZN(\AES_ENC/us21/n1115 ) );
INV_X4 \AES_ENC/us21/U364  ( .A(\AES_ENC/us21/n1094 ), .ZN(\AES_ENC/us21/n587 ) );
NOR2_X2 \AES_ENC/us21/U363  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n931 ), .ZN(\AES_ENC/us21/n1100 ) );
INV_X4 \AES_ENC/us21/U354  ( .A(\AES_ENC/us21/n1093 ), .ZN(\AES_ENC/us21/n591 ) );
NOR2_X2 \AES_ENC/us21/U353  ( .A1(\AES_ENC/us21/n569 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n929 ) );
NOR2_X2 \AES_ENC/us21/U352  ( .A1(\AES_ENC/us21/n609 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n926 ) );
NOR2_X2 \AES_ENC/us21/U351  ( .A1(\AES_ENC/us21/n572 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n1095 ) );
NOR2_X2 \AES_ENC/us21/U350  ( .A1(\AES_ENC/us21/n582 ), .A2(\AES_ENC/us21/n595 ), .ZN(\AES_ENC/us21/n1010 ) );
NOR2_X2 \AES_ENC/us21/U349  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n1103 ) );
NOR2_X2 \AES_ENC/us21/U348  ( .A1(\AES_ENC/us21/n614 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n1059 ) );
NOR2_X2 \AES_ENC/us21/U347  ( .A1(\AES_ENC/sa21 [1]), .A2(\AES_ENC/us21/n1120 ), .ZN(\AES_ENC/us21/n1022 ) );
NOR2_X2 \AES_ENC/us21/U346  ( .A1(\AES_ENC/us21/n605 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n911 ) );
NOR2_X2 \AES_ENC/us21/U345  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/us21/n1025 ), .ZN(\AES_ENC/us21/n826 ) );
NOR2_X2 \AES_ENC/us21/U338  ( .A1(\AES_ENC/us21/n594 ), .A2(\AES_ENC/us21/n579 ), .ZN(\AES_ENC/us21/n1072 ) );
NOR2_X2 \AES_ENC/us21/U335  ( .A1(\AES_ENC/us21/n595 ), .A2(\AES_ENC/us21/n590 ), .ZN(\AES_ENC/us21/n956 ) );
NOR2_X2 \AES_ENC/us21/U329  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/us21/n612 ), .ZN(\AES_ENC/us21/n1121 ) );
NOR2_X2 \AES_ENC/us21/U328  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/us21/n612 ), .ZN(\AES_ENC/us21/n1058 ) );
NOR2_X2 \AES_ENC/us21/U327  ( .A1(\AES_ENC/us21/n593 ), .A2(\AES_ENC/us21/n584 ), .ZN(\AES_ENC/us21/n1073 ) );
NOR2_X2 \AES_ENC/us21/U325  ( .A1(\AES_ENC/sa21 [1]), .A2(\AES_ENC/us21/n1025 ), .ZN(\AES_ENC/us21/n1054 ) );
NOR2_X2 \AES_ENC/us21/U324  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/us21/n931 ), .ZN(\AES_ENC/us21/n1029 ) );
NOR2_X2 \AES_ENC/us21/U319  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n1056 ) );
NOR2_X2 \AES_ENC/us21/U318  ( .A1(\AES_ENC/us21/n588 ), .A2(\AES_ENC/us21/n594 ), .ZN(\AES_ENC/us21/n1050 ) );
NOR2_X2 \AES_ENC/us21/U317  ( .A1(\AES_ENC/us21/n1121 ), .A2(\AES_ENC/us21/n1025 ), .ZN(\AES_ENC/us21/n1120 ) );
NOR2_X2 \AES_ENC/us21/U316  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/us21/n572 ), .ZN(\AES_ENC/us21/n1074 ) );
NOR2_X2 \AES_ENC/us21/U315  ( .A1(\AES_ENC/us21/n1058 ), .A2(\AES_ENC/us21/n1054 ), .ZN(\AES_ENC/us21/n878 ) );
NOR2_X2 \AES_ENC/us21/U314  ( .A1(\AES_ENC/us21/n878 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n879 ) );
NOR2_X2 \AES_ENC/us21/U312  ( .A1(\AES_ENC/us21/n880 ), .A2(\AES_ENC/us21/n879 ), .ZN(\AES_ENC/us21/n887 ) );
NOR2_X2 \AES_ENC/us21/U311  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n625 ), .ZN(\AES_ENC/us21/n957 ) );
NOR2_X2 \AES_ENC/us21/U310  ( .A1(\AES_ENC/us21/n958 ), .A2(\AES_ENC/us21/n957 ), .ZN(\AES_ENC/us21/n965 ) );
NOR3_X2 \AES_ENC/us21/U309  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n1091 ), .A3(\AES_ENC/us21/n1022 ), .ZN(\AES_ENC/us21/n720 ) );
NOR3_X2 \AES_ENC/us21/U303  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n1054 ), .A3(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n719 ) );
NOR2_X2 \AES_ENC/us21/U302  ( .A1(\AES_ENC/us21/n720 ), .A2(\AES_ENC/us21/n719 ), .ZN(\AES_ENC/us21/n726 ) );
NOR2_X2 \AES_ENC/us21/U300  ( .A1(\AES_ENC/us21/n588 ), .A2(\AES_ENC/us21/n613 ), .ZN(\AES_ENC/us21/n865 ) );
NOR2_X2 \AES_ENC/us21/U299  ( .A1(\AES_ENC/us21/n1059 ), .A2(\AES_ENC/us21/n1058 ), .ZN(\AES_ENC/us21/n1060 ) );
NOR2_X2 \AES_ENC/us21/U298  ( .A1(\AES_ENC/us21/n1095 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n668 ) );
NOR2_X2 \AES_ENC/us21/U297  ( .A1(\AES_ENC/us21/n826 ), .A2(\AES_ENC/us21/n573 ), .ZN(\AES_ENC/us21/n750 ) );
NOR2_X2 \AES_ENC/us21/U296  ( .A1(\AES_ENC/us21/n750 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n751 ) );
NOR2_X2 \AES_ENC/us21/U295  ( .A1(\AES_ENC/us21/n907 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n908 ) );
NOR2_X2 \AES_ENC/us21/U294  ( .A1(\AES_ENC/us21/n990 ), .A2(\AES_ENC/us21/n926 ), .ZN(\AES_ENC/us21/n780 ) );
NOR2_X2 \AES_ENC/us21/U293  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n606 ), .ZN(\AES_ENC/us21/n838 ) );
NOR2_X2 \AES_ENC/us21/U292  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n621 ), .ZN(\AES_ENC/us21/n837 ) );
NOR2_X2 \AES_ENC/us21/U291  ( .A1(\AES_ENC/us21/n838 ), .A2(\AES_ENC/us21/n837 ), .ZN(\AES_ENC/us21/n845 ) );
NOR2_X2 \AES_ENC/us21/U290  ( .A1(\AES_ENC/us21/n1022 ), .A2(\AES_ENC/us21/n1058 ), .ZN(\AES_ENC/us21/n740 ) );
NOR2_X2 \AES_ENC/us21/U284  ( .A1(\AES_ENC/us21/n740 ), .A2(\AES_ENC/us21/n590 ), .ZN(\AES_ENC/us21/n742 ) );
NOR2_X2 \AES_ENC/us21/U283  ( .A1(\AES_ENC/us21/n1098 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n1099 ) );
NOR2_X2 \AES_ENC/us21/U282  ( .A1(\AES_ENC/us21/n1120 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n993 ) );
NOR2_X2 \AES_ENC/us21/U281  ( .A1(\AES_ENC/us21/n993 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n994 ) );
NOR2_X2 \AES_ENC/us21/U280  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n609 ), .ZN(\AES_ENC/us21/n1026 ) );
NOR2_X2 \AES_ENC/us21/U279  ( .A1(\AES_ENC/us21/n573 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n1027 ) );
NOR2_X2 \AES_ENC/us21/U273  ( .A1(\AES_ENC/us21/n1027 ), .A2(\AES_ENC/us21/n1026 ), .ZN(\AES_ENC/us21/n1028 ) );
NOR2_X2 \AES_ENC/us21/U272  ( .A1(\AES_ENC/us21/n1029 ), .A2(\AES_ENC/us21/n1028 ), .ZN(\AES_ENC/us21/n1034 ) );
NOR4_X2 \AES_ENC/us21/U271  ( .A1(\AES_ENC/us21/n757 ), .A2(\AES_ENC/us21/n756 ), .A3(\AES_ENC/us21/n755 ), .A4(\AES_ENC/us21/n754 ), .ZN(\AES_ENC/us21/n758 ) );
NOR2_X2 \AES_ENC/us21/U270  ( .A1(\AES_ENC/us21/n752 ), .A2(\AES_ENC/us21/n751 ), .ZN(\AES_ENC/us21/n759 ) );
NOR2_X2 \AES_ENC/us21/U269  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n1071 ), .ZN(\AES_ENC/us21/n669 ) );
NOR2_X2 \AES_ENC/us21/U268  ( .A1(\AES_ENC/us21/n1056 ), .A2(\AES_ENC/us21/n990 ), .ZN(\AES_ENC/us21/n991 ) );
NOR2_X2 \AES_ENC/us21/U267  ( .A1(\AES_ENC/us21/n991 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n995 ) );
NOR2_X2 \AES_ENC/us21/U263  ( .A1(\AES_ENC/us21/n579 ), .A2(\AES_ENC/us21/n598 ), .ZN(\AES_ENC/us21/n1008 ) );
NOR2_X2 \AES_ENC/us21/U262  ( .A1(\AES_ENC/us21/n839 ), .A2(\AES_ENC/us21/n603 ), .ZN(\AES_ENC/us21/n693 ) );
NOR2_X2 \AES_ENC/us21/U258  ( .A1(\AES_ENC/us21/n578 ), .A2(\AES_ENC/us21/n906 ), .ZN(\AES_ENC/us21/n741 ) );
NOR2_X2 \AES_ENC/us21/U255  ( .A1(\AES_ENC/us21/n1054 ), .A2(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n763 ) );
NOR2_X2 \AES_ENC/us21/U254  ( .A1(\AES_ENC/us21/n763 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n769 ) );
NOR2_X2 \AES_ENC/us21/U253  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n618 ), .ZN(\AES_ENC/us21/n1007 ) );
NOR2_X2 \AES_ENC/us21/U252  ( .A1(\AES_ENC/us21/n582 ), .A2(\AES_ENC/us21/n599 ), .ZN(\AES_ENC/us21/n1123 ) );
NOR2_X2 \AES_ENC/us21/U251  ( .A1(\AES_ENC/us21/n582 ), .A2(\AES_ENC/us21/n598 ), .ZN(\AES_ENC/us21/n710 ) );
INV_X4 \AES_ENC/us21/U250  ( .A(\AES_ENC/us21/n1029 ), .ZN(\AES_ENC/us21/n603 ) );
NOR2_X2 \AES_ENC/us21/U243  ( .A1(\AES_ENC/us21/n590 ), .A2(\AES_ENC/us21/n607 ), .ZN(\AES_ENC/us21/n883 ) );
NOR2_X2 \AES_ENC/us21/U242  ( .A1(\AES_ENC/us21/n623 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n1125 ) );
NOR2_X2 \AES_ENC/us21/U241  ( .A1(\AES_ENC/us21/n911 ), .A2(\AES_ENC/us21/n910 ), .ZN(\AES_ENC/us21/n912 ) );
NOR2_X2 \AES_ENC/us21/U240  ( .A1(\AES_ENC/us21/n912 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n916 ) );
NOR2_X2 \AES_ENC/us21/U239  ( .A1(\AES_ENC/us21/n990 ), .A2(\AES_ENC/us21/n929 ), .ZN(\AES_ENC/us21/n892 ) );
NOR2_X2 \AES_ENC/us21/U238  ( .A1(\AES_ENC/us21/n892 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n893 ) );
NOR2_X2 \AES_ENC/us21/U237  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n621 ), .ZN(\AES_ENC/us21/n950 ) );
NOR2_X2 \AES_ENC/us21/U236  ( .A1(\AES_ENC/us21/n1079 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n1082 ) );
NOR2_X2 \AES_ENC/us21/U235  ( .A1(\AES_ENC/us21/n910 ), .A2(\AES_ENC/us21/n1056 ), .ZN(\AES_ENC/us21/n941 ) );
NOR2_X2 \AES_ENC/us21/U234  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n1077 ), .ZN(\AES_ENC/us21/n841 ) );
NOR2_X2 \AES_ENC/us21/U229  ( .A1(\AES_ENC/us21/n601 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n630 ) );
NOR2_X2 \AES_ENC/us21/U228  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n621 ), .ZN(\AES_ENC/us21/n806 ) );
NOR2_X2 \AES_ENC/us21/U227  ( .A1(\AES_ENC/us21/n601 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n948 ) );
NOR2_X2 \AES_ENC/us21/U226  ( .A1(\AES_ENC/us21/n578 ), .A2(\AES_ENC/us21/n620 ), .ZN(\AES_ENC/us21/n997 ) );
NOR2_X2 \AES_ENC/us21/U225  ( .A1(\AES_ENC/us21/n1121 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n1122 ) );
NOR2_X2 \AES_ENC/us21/U223  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n1023 ), .ZN(\AES_ENC/us21/n756 ) );
NOR2_X2 \AES_ENC/us21/U222  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n621 ), .ZN(\AES_ENC/us21/n870 ) );
NOR2_X2 \AES_ENC/us21/U221  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n569 ), .ZN(\AES_ENC/us21/n947 ) );
NOR2_X2 \AES_ENC/us21/U217  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n1077 ), .ZN(\AES_ENC/us21/n1084 ) );
NOR2_X2 \AES_ENC/us21/U213  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n855 ), .ZN(\AES_ENC/us21/n709 ) );
NOR2_X2 \AES_ENC/us21/U212  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n620 ), .ZN(\AES_ENC/us21/n868 ) );
NOR2_X2 \AES_ENC/us21/U211  ( .A1(\AES_ENC/us21/n1120 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n1124 ) );
NOR2_X2 \AES_ENC/us21/U210  ( .A1(\AES_ENC/us21/n1120 ), .A2(\AES_ENC/us21/n839 ), .ZN(\AES_ENC/us21/n842 ) );
NOR2_X2 \AES_ENC/us21/U209  ( .A1(\AES_ENC/us21/n1120 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n696 ) );
NOR2_X2 \AES_ENC/us21/U208  ( .A1(\AES_ENC/us21/n1074 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n1076 ) );
NOR2_X2 \AES_ENC/us21/U207  ( .A1(\AES_ENC/us21/n1074 ), .A2(\AES_ENC/us21/n609 ), .ZN(\AES_ENC/us21/n781 ) );
NOR3_X2 \AES_ENC/us21/U201  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n1056 ), .A3(\AES_ENC/us21/n990 ), .ZN(\AES_ENC/us21/n979 ) );
NOR3_X2 \AES_ENC/us21/U200  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n1058 ), .A3(\AES_ENC/us21/n1059 ), .ZN(\AES_ENC/us21/n854 ) );
NOR2_X2 \AES_ENC/us21/U199  ( .A1(\AES_ENC/us21/n996 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n869 ) );
NOR2_X2 \AES_ENC/us21/U198  ( .A1(\AES_ENC/us21/n1056 ), .A2(\AES_ENC/us21/n1074 ), .ZN(\AES_ENC/us21/n1057 ) );
NOR3_X2 \AES_ENC/us21/U197  ( .A1(\AES_ENC/us21/n579 ), .A2(\AES_ENC/us21/n1120 ), .A3(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n978 ) );
NOR2_X2 \AES_ENC/us21/U196  ( .A1(\AES_ENC/us21/n996 ), .A2(\AES_ENC/us21/n911 ), .ZN(\AES_ENC/us21/n1116 ) );
NOR2_X2 \AES_ENC/us21/U195  ( .A1(\AES_ENC/us21/n1074 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n754 ) );
NOR2_X2 \AES_ENC/us21/U194  ( .A1(\AES_ENC/us21/n926 ), .A2(\AES_ENC/us21/n1103 ), .ZN(\AES_ENC/us21/n977 ) );
NOR2_X2 \AES_ENC/us21/U187  ( .A1(\AES_ENC/us21/n839 ), .A2(\AES_ENC/us21/n824 ), .ZN(\AES_ENC/us21/n1092 ) );
NOR2_X2 \AES_ENC/us21/U186  ( .A1(\AES_ENC/us21/n573 ), .A2(\AES_ENC/us21/n1074 ), .ZN(\AES_ENC/us21/n684 ) );
NOR2_X2 \AES_ENC/us21/U185  ( .A1(\AES_ENC/us21/n826 ), .A2(\AES_ENC/us21/n1059 ), .ZN(\AES_ENC/us21/n907 ) );
NOR3_X2 \AES_ENC/us21/U184  ( .A1(\AES_ENC/us21/n593 ), .A2(\AES_ENC/us21/n1115 ), .A3(\AES_ENC/us21/n600 ), .ZN(\AES_ENC/us21/n831 ) );
NOR3_X2 \AES_ENC/us21/U183  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n1056 ), .A3(\AES_ENC/us21/n990 ), .ZN(\AES_ENC/us21/n896 ) );
NOR3_X2 \AES_ENC/us21/U182  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n573 ), .A3(\AES_ENC/us21/n1013 ), .ZN(\AES_ENC/us21/n670 ) );
NOR3_X2 \AES_ENC/us21/U181  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n1091 ), .A3(\AES_ENC/us21/n1022 ), .ZN(\AES_ENC/us21/n843 ) );
NOR2_X2 \AES_ENC/us21/U180  ( .A1(\AES_ENC/us21/n1029 ), .A2(\AES_ENC/us21/n1095 ), .ZN(\AES_ENC/us21/n735 ) );
NOR2_X2 \AES_ENC/us21/U174  ( .A1(\AES_ENC/us21/n1100 ), .A2(\AES_ENC/us21/n854 ), .ZN(\AES_ENC/us21/n860 ) );
NAND3_X2 \AES_ENC/us21/U173  ( .A1(\AES_ENC/us21/n569 ), .A2(\AES_ENC/us21/n603 ), .A3(\AES_ENC/us21/n681 ), .ZN(\AES_ENC/us21/n691 ) );
NOR2_X2 \AES_ENC/us21/U172  ( .A1(\AES_ENC/us21/n683 ), .A2(\AES_ENC/us21/n682 ), .ZN(\AES_ENC/us21/n690 ) );
NOR3_X2 \AES_ENC/us21/U171  ( .A1(\AES_ENC/us21/n695 ), .A2(\AES_ENC/us21/n694 ), .A3(\AES_ENC/us21/n693 ), .ZN(\AES_ENC/us21/n700 ) );
NOR4_X2 \AES_ENC/us21/U170  ( .A1(\AES_ENC/us21/n983 ), .A2(\AES_ENC/us21/n698 ), .A3(\AES_ENC/us21/n697 ), .A4(\AES_ENC/us21/n696 ), .ZN(\AES_ENC/us21/n699 ) );
NOR2_X2 \AES_ENC/us21/U169  ( .A1(\AES_ENC/us21/n946 ), .A2(\AES_ENC/us21/n945 ), .ZN(\AES_ENC/us21/n952 ) );
NOR4_X2 \AES_ENC/us21/U168  ( .A1(\AES_ENC/us21/n950 ), .A2(\AES_ENC/us21/n949 ), .A3(\AES_ENC/us21/n948 ), .A4(\AES_ENC/us21/n947 ), .ZN(\AES_ENC/us21/n951 ) );
NOR4_X2 \AES_ENC/us21/U162  ( .A1(\AES_ENC/us21/n896 ), .A2(\AES_ENC/us21/n895 ), .A3(\AES_ENC/us21/n894 ), .A4(\AES_ENC/us21/n893 ), .ZN(\AES_ENC/us21/n897 ) );
NOR2_X2 \AES_ENC/us21/U161  ( .A1(\AES_ENC/us21/n866 ), .A2(\AES_ENC/us21/n865 ), .ZN(\AES_ENC/us21/n872 ) );
NOR4_X2 \AES_ENC/us21/U160  ( .A1(\AES_ENC/us21/n870 ), .A2(\AES_ENC/us21/n869 ), .A3(\AES_ENC/us21/n868 ), .A4(\AES_ENC/us21/n867 ), .ZN(\AES_ENC/us21/n871 ) );
NOR4_X2 \AES_ENC/us21/U159  ( .A1(\AES_ENC/us21/n983 ), .A2(\AES_ENC/us21/n982 ), .A3(\AES_ENC/us21/n981 ), .A4(\AES_ENC/us21/n980 ), .ZN(\AES_ENC/us21/n984 ) );
NOR2_X2 \AES_ENC/us21/U158  ( .A1(\AES_ENC/us21/n979 ), .A2(\AES_ENC/us21/n978 ), .ZN(\AES_ENC/us21/n985 ) );
NOR4_X2 \AES_ENC/us21/U157  ( .A1(\AES_ENC/us21/n1125 ), .A2(\AES_ENC/us21/n1124 ), .A3(\AES_ENC/us21/n1123 ), .A4(\AES_ENC/us21/n1122 ), .ZN(\AES_ENC/us21/n1126 ) );
NOR4_X2 \AES_ENC/us21/U156  ( .A1(\AES_ENC/us21/n1084 ), .A2(\AES_ENC/us21/n1083 ), .A3(\AES_ENC/us21/n1082 ), .A4(\AES_ENC/us21/n1081 ), .ZN(\AES_ENC/us21/n1085 ) );
NOR2_X2 \AES_ENC/us21/U155  ( .A1(\AES_ENC/us21/n1076 ), .A2(\AES_ENC/us21/n1075 ), .ZN(\AES_ENC/us21/n1086 ) );
NOR3_X2 \AES_ENC/us21/U154  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n1054 ), .A3(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n961 ) );
NOR3_X2 \AES_ENC/us21/U153  ( .A1(\AES_ENC/us21/n609 ), .A2(\AES_ENC/us21/n1074 ), .A3(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n671 ) );
NOR2_X2 \AES_ENC/us21/U152  ( .A1(\AES_ENC/us21/n1057 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n1062 ) );
NOR2_X2 \AES_ENC/us21/U143  ( .A1(\AES_ENC/us21/n1055 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n1063 ) );
NOR2_X2 \AES_ENC/us21/U142  ( .A1(\AES_ENC/us21/n1060 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n1061 ) );
NOR4_X2 \AES_ENC/us21/U141  ( .A1(\AES_ENC/us21/n1064 ), .A2(\AES_ENC/us21/n1063 ), .A3(\AES_ENC/us21/n1062 ), .A4(\AES_ENC/us21/n1061 ), .ZN(\AES_ENC/us21/n1065 ) );
NOR3_X2 \AES_ENC/us21/U140  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n1120 ), .A3(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n918 ) );
NOR3_X2 \AES_ENC/us21/U132  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n573 ), .A3(\AES_ENC/us21/n1013 ), .ZN(\AES_ENC/us21/n917 ) );
NOR2_X2 \AES_ENC/us21/U131  ( .A1(\AES_ENC/us21/n914 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n915 ) );
NOR4_X2 \AES_ENC/us21/U130  ( .A1(\AES_ENC/us21/n918 ), .A2(\AES_ENC/us21/n917 ), .A3(\AES_ENC/us21/n916 ), .A4(\AES_ENC/us21/n915 ), .ZN(\AES_ENC/us21/n919 ) );
NOR2_X2 \AES_ENC/us21/U129  ( .A1(\AES_ENC/us21/n590 ), .A2(\AES_ENC/us21/n599 ), .ZN(\AES_ENC/us21/n771 ) );
NOR2_X2 \AES_ENC/us21/U128  ( .A1(\AES_ENC/us21/n1103 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n772 ) );
NOR2_X2 \AES_ENC/us21/U127  ( .A1(\AES_ENC/us21/n583 ), .A2(\AES_ENC/us21/n615 ), .ZN(\AES_ENC/us21/n773 ) );
NOR4_X2 \AES_ENC/us21/U126  ( .A1(\AES_ENC/us21/n773 ), .A2(\AES_ENC/us21/n772 ), .A3(\AES_ENC/us21/n771 ), .A4(\AES_ENC/us21/n770 ), .ZN(\AES_ENC/us21/n774 ) );
NOR2_X2 \AES_ENC/us21/U121  ( .A1(\AES_ENC/us21/n735 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n687 ) );
NOR2_X2 \AES_ENC/us21/U120  ( .A1(\AES_ENC/us21/n684 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n688 ) );
NOR2_X2 \AES_ENC/us21/U119  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n622 ), .ZN(\AES_ENC/us21/n686 ) );
NOR4_X2 \AES_ENC/us21/U118  ( .A1(\AES_ENC/us21/n688 ), .A2(\AES_ENC/us21/n687 ), .A3(\AES_ENC/us21/n686 ), .A4(\AES_ENC/us21/n685 ), .ZN(\AES_ENC/us21/n689 ) );
NOR2_X2 \AES_ENC/us21/U117  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n608 ), .ZN(\AES_ENC/us21/n858 ) );
NOR2_X2 \AES_ENC/us21/U116  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n855 ), .ZN(\AES_ENC/us21/n857 ) );
NOR2_X2 \AES_ENC/us21/U115  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n617 ), .ZN(\AES_ENC/us21/n856 ) );
NOR4_X2 \AES_ENC/us21/U106  ( .A1(\AES_ENC/us21/n858 ), .A2(\AES_ENC/us21/n857 ), .A3(\AES_ENC/us21/n856 ), .A4(\AES_ENC/us21/n958 ), .ZN(\AES_ENC/us21/n859 ) );
NOR2_X2 \AES_ENC/us21/U105  ( .A1(\AES_ENC/us21/n780 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n784 ) );
NOR2_X2 \AES_ENC/us21/U104  ( .A1(\AES_ENC/us21/n1117 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n782 ) );
NOR2_X2 \AES_ENC/us21/U103  ( .A1(\AES_ENC/us21/n781 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n783 ) );
NOR4_X2 \AES_ENC/us21/U102  ( .A1(\AES_ENC/us21/n880 ), .A2(\AES_ENC/us21/n784 ), .A3(\AES_ENC/us21/n783 ), .A4(\AES_ENC/us21/n782 ), .ZN(\AES_ENC/us21/n785 ) );
NOR2_X2 \AES_ENC/us21/U101  ( .A1(\AES_ENC/us21/n597 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n814 ) );
NOR2_X2 \AES_ENC/us21/U100  ( .A1(\AES_ENC/us21/n907 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n813 ) );
NOR3_X2 \AES_ENC/us21/U95  ( .A1(\AES_ENC/us21/n578 ), .A2(\AES_ENC/us21/n1058 ), .A3(\AES_ENC/us21/n1059 ), .ZN(\AES_ENC/us21/n815 ) );
NOR4_X2 \AES_ENC/us21/U94  ( .A1(\AES_ENC/us21/n815 ), .A2(\AES_ENC/us21/n814 ), .A3(\AES_ENC/us21/n813 ), .A4(\AES_ENC/us21/n812 ), .ZN(\AES_ENC/us21/n816 ) );
NOR2_X2 \AES_ENC/us21/U93  ( .A1(\AES_ENC/us21/n591 ), .A2(\AES_ENC/us21/n569 ), .ZN(\AES_ENC/us21/n721 ) );
NOR2_X2 \AES_ENC/us21/U92  ( .A1(\AES_ENC/us21/n1031 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n723 ) );
NOR2_X2 \AES_ENC/us21/U91  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n1096 ), .ZN(\AES_ENC/us21/n722 ) );
NOR4_X2 \AES_ENC/us21/U90  ( .A1(\AES_ENC/us21/n724 ), .A2(\AES_ENC/us21/n723 ), .A3(\AES_ENC/us21/n722 ), .A4(\AES_ENC/us21/n721 ), .ZN(\AES_ENC/us21/n725 ) );
NOR2_X2 \AES_ENC/us21/U89  ( .A1(\AES_ENC/us21/n911 ), .A2(\AES_ENC/us21/n990 ), .ZN(\AES_ENC/us21/n1009 ) );
NOR2_X2 \AES_ENC/us21/U88  ( .A1(\AES_ENC/us21/n1013 ), .A2(\AES_ENC/us21/n573 ), .ZN(\AES_ENC/us21/n1014 ) );
NOR2_X2 \AES_ENC/us21/U87  ( .A1(\AES_ENC/us21/n1014 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n1015 ) );
NOR4_X2 \AES_ENC/us21/U86  ( .A1(\AES_ENC/us21/n1016 ), .A2(\AES_ENC/us21/n1015 ), .A3(\AES_ENC/us21/n1119 ), .A4(\AES_ENC/us21/n1046 ), .ZN(\AES_ENC/us21/n1017 ) );
NOR2_X2 \AES_ENC/us21/U81  ( .A1(\AES_ENC/us21/n996 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n998 ) );
NOR2_X2 \AES_ENC/us21/U80  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n618 ), .ZN(\AES_ENC/us21/n1000 ) );
NOR2_X2 \AES_ENC/us21/U79  ( .A1(\AES_ENC/us21/n590 ), .A2(\AES_ENC/us21/n1096 ), .ZN(\AES_ENC/us21/n999 ) );
NOR4_X2 \AES_ENC/us21/U78  ( .A1(\AES_ENC/us21/n1000 ), .A2(\AES_ENC/us21/n999 ), .A3(\AES_ENC/us21/n998 ), .A4(\AES_ENC/us21/n997 ), .ZN(\AES_ENC/us21/n1001 ) );
NOR2_X2 \AES_ENC/us21/U74  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n1096 ), .ZN(\AES_ENC/us21/n697 ) );
NOR2_X2 \AES_ENC/us21/U73  ( .A1(\AES_ENC/us21/n609 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n958 ) );
NOR2_X2 \AES_ENC/us21/U72  ( .A1(\AES_ENC/us21/n911 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n983 ) );
NOR2_X2 \AES_ENC/us21/U71  ( .A1(\AES_ENC/us21/n1054 ), .A2(\AES_ENC/us21/n1103 ), .ZN(\AES_ENC/us21/n1031 ) );
INV_X4 \AES_ENC/us21/U65  ( .A(\AES_ENC/us21/n1050 ), .ZN(\AES_ENC/us21/n585 ) );
INV_X4 \AES_ENC/us21/U64  ( .A(\AES_ENC/us21/n1072 ), .ZN(\AES_ENC/us21/n577 ) );
INV_X4 \AES_ENC/us21/U63  ( .A(\AES_ENC/us21/n1073 ), .ZN(\AES_ENC/us21/n576 ) );
NOR2_X2 \AES_ENC/us21/U62  ( .A1(\AES_ENC/us21/n603 ), .A2(\AES_ENC/us21/n587 ), .ZN(\AES_ENC/us21/n880 ) );
NOR3_X2 \AES_ENC/us21/U61  ( .A1(\AES_ENC/us21/n826 ), .A2(\AES_ENC/us21/n1121 ), .A3(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n946 ) );
INV_X4 \AES_ENC/us21/U59  ( .A(\AES_ENC/us21/n1010 ), .ZN(\AES_ENC/us21/n581 ) );
NOR3_X2 \AES_ENC/us21/U58  ( .A1(\AES_ENC/us21/n573 ), .A2(\AES_ENC/us21/n1029 ), .A3(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n1119 ) );
INV_X4 \AES_ENC/us21/U57  ( .A(\AES_ENC/us21/n956 ), .ZN(\AES_ENC/us21/n589 ) );
NOR2_X2 \AES_ENC/us21/U50  ( .A1(\AES_ENC/us21/n601 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n1013 ) );
NOR2_X2 \AES_ENC/us21/U49  ( .A1(\AES_ENC/us21/n609 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n910 ) );
NOR2_X2 \AES_ENC/us21/U48  ( .A1(\AES_ENC/us21/n569 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n1091 ) );
NOR2_X2 \AES_ENC/us21/U47  ( .A1(\AES_ENC/us21/n614 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n990 ) );
NOR2_X2 \AES_ENC/us21/U46  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/us21/n1121 ), .ZN(\AES_ENC/us21/n996 ) );
NOR2_X2 \AES_ENC/us21/U45  ( .A1(\AES_ENC/us21/n583 ), .A2(\AES_ENC/us21/n622 ), .ZN(\AES_ENC/us21/n628 ) );
NOR2_X2 \AES_ENC/us21/U44  ( .A1(\AES_ENC/us21/n602 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n866 ) );
NOR2_X2 \AES_ENC/us21/U43  ( .A1(\AES_ENC/us21/n610 ), .A2(\AES_ENC/us21/n583 ), .ZN(\AES_ENC/us21/n1006 ) );
NOR2_X2 \AES_ENC/us21/U42  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n1117 ), .ZN(\AES_ENC/us21/n1118 ) );
NOR2_X2 \AES_ENC/us21/U41  ( .A1(\AES_ENC/us21/n1119 ), .A2(\AES_ENC/us21/n1118 ), .ZN(\AES_ENC/us21/n1127 ) );
NOR2_X2 \AES_ENC/us21/U36  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n616 ), .ZN(\AES_ENC/us21/n629 ) );
NOR2_X2 \AES_ENC/us21/U35  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n906 ), .ZN(\AES_ENC/us21/n909 ) );
NOR2_X2 \AES_ENC/us21/U34  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n607 ), .ZN(\AES_ENC/us21/n658 ) );
NOR2_X2 \AES_ENC/us21/U33  ( .A1(\AES_ENC/us21/n1116 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n695 ) );
NOR2_X2 \AES_ENC/us21/U32  ( .A1(\AES_ENC/us21/n1078 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n1083 ) );
NOR2_X2 \AES_ENC/us21/U31  ( .A1(\AES_ENC/us21/n941 ), .A2(\AES_ENC/us21/n581 ), .ZN(\AES_ENC/us21/n724 ) );
NOR2_X2 \AES_ENC/us21/U30  ( .A1(\AES_ENC/us21/n611 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n1107 ) );
NOR2_X2 \AES_ENC/us21/U29  ( .A1(\AES_ENC/us21/n602 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n840 ) );
NOR2_X2 \AES_ENC/us21/U24  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n623 ), .ZN(\AES_ENC/us21/n633 ) );
NOR2_X2 \AES_ENC/us21/U23  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n1080 ), .ZN(\AES_ENC/us21/n1081 ) );
NOR2_X2 \AES_ENC/us21/U21  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n1045 ), .ZN(\AES_ENC/us21/n812 ) );
NOR2_X2 \AES_ENC/us21/U20  ( .A1(\AES_ENC/us21/n1009 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n960 ) );
NOR2_X2 \AES_ENC/us21/U19  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n619 ), .ZN(\AES_ENC/us21/n982 ) );
NOR2_X2 \AES_ENC/us21/U18  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n616 ), .ZN(\AES_ENC/us21/n757 ) );
NOR2_X2 \AES_ENC/us21/U17  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n598 ), .ZN(\AES_ENC/us21/n698 ) );
NOR2_X2 \AES_ENC/us21/U16  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n605 ), .ZN(\AES_ENC/us21/n708 ) );
NOR2_X2 \AES_ENC/us21/U15  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n603 ), .ZN(\AES_ENC/us21/n770 ) );
NOR2_X2 \AES_ENC/us21/U10  ( .A1(\AES_ENC/us21/n605 ), .A2(\AES_ENC/us21/n576 ), .ZN(\AES_ENC/us21/n803 ) );
NOR2_X2 \AES_ENC/us21/U9  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n881 ), .ZN(\AES_ENC/us21/n711 ) );
NOR2_X2 \AES_ENC/us21/U8  ( .A1(\AES_ENC/us21/n589 ), .A2(\AES_ENC/us21/n603 ), .ZN(\AES_ENC/us21/n867 ) );
NOR2_X2 \AES_ENC/us21/U7  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n615 ), .ZN(\AES_ENC/us21/n804 ) );
NOR2_X2 \AES_ENC/us21/U6  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n609 ), .ZN(\AES_ENC/us21/n1046 ) );
OR2_X4 \AES_ENC/us21/U5  ( .A1(\AES_ENC/us21/n612 ), .A2(\AES_ENC/sa21 [1]),.ZN(\AES_ENC/us21/n570 ) );
OR2_X4 \AES_ENC/us21/U4  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/sa21 [4]),.ZN(\AES_ENC/us21/n569 ) );
NAND2_X2 \AES_ENC/us21/U514  ( .A1(\AES_ENC/us21/n1121 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n1030 ) );
AND2_X2 \AES_ENC/us21/U513  ( .A1(\AES_ENC/us21/n607 ), .A2(\AES_ENC/us21/n1030 ), .ZN(\AES_ENC/us21/n1049 ) );
NAND2_X2 \AES_ENC/us21/U511  ( .A1(\AES_ENC/us21/n1049 ), .A2(\AES_ENC/us21/n794 ), .ZN(\AES_ENC/us21/n637 ) );
AND2_X2 \AES_ENC/us21/U493  ( .A1(\AES_ENC/us21/n779 ), .A2(\AES_ENC/us21/n996 ), .ZN(\AES_ENC/us21/n632 ) );
NAND4_X2 \AES_ENC/us21/U485  ( .A1(\AES_ENC/us21/n637 ), .A2(\AES_ENC/us21/n636 ), .A3(\AES_ENC/us21/n635 ), .A4(\AES_ENC/us21/n634 ), .ZN(\AES_ENC/us21/n638 ) );
NAND2_X2 \AES_ENC/us21/U484  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n638 ), .ZN(\AES_ENC/us21/n679 ) );
NAND2_X2 \AES_ENC/us21/U481  ( .A1(\AES_ENC/us21/n1094 ), .A2(\AES_ENC/us21/n613 ), .ZN(\AES_ENC/us21/n648 ) );
NAND2_X2 \AES_ENC/us21/U476  ( .A1(\AES_ENC/us21/n619 ), .A2(\AES_ENC/us21/n598 ), .ZN(\AES_ENC/us21/n762 ) );
NAND2_X2 \AES_ENC/us21/U475  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n762 ), .ZN(\AES_ENC/us21/n647 ) );
NAND4_X2 \AES_ENC/us21/U457  ( .A1(\AES_ENC/us21/n648 ), .A2(\AES_ENC/us21/n647 ), .A3(\AES_ENC/us21/n646 ), .A4(\AES_ENC/us21/n645 ), .ZN(\AES_ENC/us21/n649 ) );
NAND2_X2 \AES_ENC/us21/U456  ( .A1(\AES_ENC/sa21 [0]), .A2(\AES_ENC/us21/n649 ), .ZN(\AES_ENC/us21/n665 ) );
NAND2_X2 \AES_ENC/us21/U454  ( .A1(\AES_ENC/us21/n626 ), .A2(\AES_ENC/us21/n601 ), .ZN(\AES_ENC/us21/n855 ) );
NAND2_X2 \AES_ENC/us21/U453  ( .A1(\AES_ENC/us21/n617 ), .A2(\AES_ENC/us21/n855 ), .ZN(\AES_ENC/us21/n821 ) );
NAND2_X2 \AES_ENC/us21/U452  ( .A1(\AES_ENC/us21/n1093 ), .A2(\AES_ENC/us21/n821 ), .ZN(\AES_ENC/us21/n662 ) );
NAND2_X2 \AES_ENC/us21/U451  ( .A1(\AES_ENC/us21/n605 ), .A2(\AES_ENC/us21/n620 ), .ZN(\AES_ENC/us21/n650 ) );
NAND2_X2 \AES_ENC/us21/U450  ( .A1(\AES_ENC/us21/n956 ), .A2(\AES_ENC/us21/n650 ), .ZN(\AES_ENC/us21/n661 ) );
NAND2_X2 \AES_ENC/us21/U449  ( .A1(\AES_ENC/us21/n594 ), .A2(\AES_ENC/us21/n595 ), .ZN(\AES_ENC/us21/n839 ) );
OR2_X2 \AES_ENC/us21/U446  ( .A1(\AES_ENC/us21/n839 ), .A2(\AES_ENC/us21/n932 ), .ZN(\AES_ENC/us21/n656 ) );
NAND2_X2 \AES_ENC/us21/U445  ( .A1(\AES_ENC/us21/n624 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n1096 ) );
NAND2_X2 \AES_ENC/us21/U444  ( .A1(\AES_ENC/us21/n1030 ), .A2(\AES_ENC/us21/n1096 ), .ZN(\AES_ENC/us21/n651 ) );
NAND2_X2 \AES_ENC/us21/U443  ( .A1(\AES_ENC/us21/n1114 ), .A2(\AES_ENC/us21/n651 ), .ZN(\AES_ENC/us21/n655 ) );
OR3_X2 \AES_ENC/us21/U440  ( .A1(\AES_ENC/us21/n1079 ), .A2(\AES_ENC/sa21 [7]), .A3(\AES_ENC/us21/n594 ), .ZN(\AES_ENC/us21/n654 ));
NAND2_X2 \AES_ENC/us21/U439  ( .A1(\AES_ENC/us21/n623 ), .A2(\AES_ENC/us21/n619 ), .ZN(\AES_ENC/us21/n652 ) );
NAND4_X2 \AES_ENC/us21/U437  ( .A1(\AES_ENC/us21/n656 ), .A2(\AES_ENC/us21/n655 ), .A3(\AES_ENC/us21/n654 ), .A4(\AES_ENC/us21/n653 ), .ZN(\AES_ENC/us21/n657 ) );
NAND2_X2 \AES_ENC/us21/U436  ( .A1(\AES_ENC/sa21 [2]), .A2(\AES_ENC/us21/n657 ), .ZN(\AES_ENC/us21/n660 ) );
NAND4_X2 \AES_ENC/us21/U432  ( .A1(\AES_ENC/us21/n662 ), .A2(\AES_ENC/us21/n661 ), .A3(\AES_ENC/us21/n660 ), .A4(\AES_ENC/us21/n659 ), .ZN(\AES_ENC/us21/n663 ) );
NAND2_X2 \AES_ENC/us21/U431  ( .A1(\AES_ENC/us21/n663 ), .A2(\AES_ENC/us21/n627 ), .ZN(\AES_ENC/us21/n664 ) );
NAND2_X2 \AES_ENC/us21/U430  ( .A1(\AES_ENC/us21/n665 ), .A2(\AES_ENC/us21/n664 ), .ZN(\AES_ENC/us21/n666 ) );
NAND2_X2 \AES_ENC/us21/U429  ( .A1(\AES_ENC/sa21 [6]), .A2(\AES_ENC/us21/n666 ), .ZN(\AES_ENC/us21/n678 ) );
NAND2_X2 \AES_ENC/us21/U426  ( .A1(\AES_ENC/us21/n735 ), .A2(\AES_ENC/us21/n1093 ), .ZN(\AES_ENC/us21/n675 ) );
NAND2_X2 \AES_ENC/us21/U425  ( .A1(\AES_ENC/us21/n625 ), .A2(\AES_ENC/us21/n607 ), .ZN(\AES_ENC/us21/n1045 ) );
OR2_X2 \AES_ENC/us21/U424  ( .A1(\AES_ENC/us21/n1045 ), .A2(\AES_ENC/us21/n577 ), .ZN(\AES_ENC/us21/n674 ) );
NAND2_X2 \AES_ENC/us21/U423  ( .A1(\AES_ENC/sa21 [1]), .A2(\AES_ENC/us21/n609 ), .ZN(\AES_ENC/us21/n667 ) );
NAND2_X2 \AES_ENC/us21/U422  ( .A1(\AES_ENC/us21/n605 ), .A2(\AES_ENC/us21/n667 ), .ZN(\AES_ENC/us21/n1071 ) );
NAND4_X2 \AES_ENC/us21/U412  ( .A1(\AES_ENC/us21/n675 ), .A2(\AES_ENC/us21/n674 ), .A3(\AES_ENC/us21/n673 ), .A4(\AES_ENC/us21/n672 ), .ZN(\AES_ENC/us21/n676 ) );
NAND2_X2 \AES_ENC/us21/U411  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n676 ), .ZN(\AES_ENC/us21/n677 ) );
NAND2_X2 \AES_ENC/us21/U408  ( .A1(\AES_ENC/us21/n800 ), .A2(\AES_ENC/us21/n1022 ), .ZN(\AES_ENC/us21/n680 ) );
NAND2_X2 \AES_ENC/us21/U407  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n680 ), .ZN(\AES_ENC/us21/n681 ) );
AND2_X2 \AES_ENC/us21/U402  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n684 ), .ZN(\AES_ENC/us21/n682 ) );
NAND4_X2 \AES_ENC/us21/U395  ( .A1(\AES_ENC/us21/n691 ), .A2(\AES_ENC/us21/n586 ), .A3(\AES_ENC/us21/n690 ), .A4(\AES_ENC/us21/n689 ), .ZN(\AES_ENC/us21/n692 ) );
NAND2_X2 \AES_ENC/us21/U394  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n692 ), .ZN(\AES_ENC/us21/n733 ) );
NAND2_X2 \AES_ENC/us21/U392  ( .A1(\AES_ENC/us21/n977 ), .A2(\AES_ENC/us21/n1050 ), .ZN(\AES_ENC/us21/n702 ) );
NAND2_X2 \AES_ENC/us21/U391  ( .A1(\AES_ENC/us21/n1093 ), .A2(\AES_ENC/us21/n1045 ), .ZN(\AES_ENC/us21/n701 ) );
NAND4_X2 \AES_ENC/us21/U381  ( .A1(\AES_ENC/us21/n702 ), .A2(\AES_ENC/us21/n701 ), .A3(\AES_ENC/us21/n700 ), .A4(\AES_ENC/us21/n699 ), .ZN(\AES_ENC/us21/n703 ) );
NAND2_X2 \AES_ENC/us21/U380  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n703 ), .ZN(\AES_ENC/us21/n732 ) );
AND2_X2 \AES_ENC/us21/U379  ( .A1(\AES_ENC/sa21 [0]), .A2(\AES_ENC/sa21 [6]),.ZN(\AES_ENC/us21/n1113 ) );
NAND2_X2 \AES_ENC/us21/U378  ( .A1(\AES_ENC/us21/n619 ), .A2(\AES_ENC/us21/n1030 ), .ZN(\AES_ENC/us21/n881 ) );
NAND2_X2 \AES_ENC/us21/U377  ( .A1(\AES_ENC/us21/n1093 ), .A2(\AES_ENC/us21/n881 ), .ZN(\AES_ENC/us21/n715 ) );
NAND2_X2 \AES_ENC/us21/U376  ( .A1(\AES_ENC/us21/n1010 ), .A2(\AES_ENC/us21/n622 ), .ZN(\AES_ENC/us21/n714 ) );
NAND2_X2 \AES_ENC/us21/U375  ( .A1(\AES_ENC/us21/n855 ), .A2(\AES_ENC/us21/n625 ), .ZN(\AES_ENC/us21/n1117 ) );
XNOR2_X2 \AES_ENC/us21/U371  ( .A(\AES_ENC/us21/n584 ), .B(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n824 ) );
NAND4_X2 \AES_ENC/us21/U362  ( .A1(\AES_ENC/us21/n715 ), .A2(\AES_ENC/us21/n714 ), .A3(\AES_ENC/us21/n713 ), .A4(\AES_ENC/us21/n712 ), .ZN(\AES_ENC/us21/n716 ) );
NAND2_X2 \AES_ENC/us21/U361  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n716 ), .ZN(\AES_ENC/us21/n731 ) );
AND2_X2 \AES_ENC/us21/U360  ( .A1(\AES_ENC/sa21 [6]), .A2(\AES_ENC/us21/n627 ), .ZN(\AES_ENC/us21/n1131 ) );
NAND2_X2 \AES_ENC/us21/U359  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n717 ) );
NAND2_X2 \AES_ENC/us21/U358  ( .A1(\AES_ENC/us21/n1029 ), .A2(\AES_ENC/us21/n717 ), .ZN(\AES_ENC/us21/n728 ) );
NAND2_X2 \AES_ENC/us21/U357  ( .A1(\AES_ENC/sa21 [1]), .A2(\AES_ENC/us21/n612 ), .ZN(\AES_ENC/us21/n1097 ) );
NAND2_X2 \AES_ENC/us21/U356  ( .A1(\AES_ENC/us21/n610 ), .A2(\AES_ENC/us21/n1097 ), .ZN(\AES_ENC/us21/n718 ) );
NAND2_X2 \AES_ENC/us21/U355  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n718 ), .ZN(\AES_ENC/us21/n727 ) );
NAND4_X2 \AES_ENC/us21/U344  ( .A1(\AES_ENC/us21/n728 ), .A2(\AES_ENC/us21/n727 ), .A3(\AES_ENC/us21/n726 ), .A4(\AES_ENC/us21/n725 ), .ZN(\AES_ENC/us21/n729 ) );
NAND2_X2 \AES_ENC/us21/U343  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n729 ), .ZN(\AES_ENC/us21/n730 ) );
NAND4_X2 \AES_ENC/us21/U342  ( .A1(\AES_ENC/us21/n733 ), .A2(\AES_ENC/us21/n732 ), .A3(\AES_ENC/us21/n731 ), .A4(\AES_ENC/us21/n730 ), .ZN(\AES_ENC/sa21_sub[1] ) );
NAND2_X2 \AES_ENC/us21/U341  ( .A1(\AES_ENC/sa21 [7]), .A2(\AES_ENC/us21/n584 ), .ZN(\AES_ENC/us21/n734 ) );
NAND2_X2 \AES_ENC/us21/U340  ( .A1(\AES_ENC/us21/n734 ), .A2(\AES_ENC/us21/n579 ), .ZN(\AES_ENC/us21/n738 ) );
OR4_X2 \AES_ENC/us21/U339  ( .A1(\AES_ENC/us21/n738 ), .A2(\AES_ENC/us21/n594 ), .A3(\AES_ENC/us21/n826 ), .A4(\AES_ENC/us21/n1121 ), .ZN(\AES_ENC/us21/n746 ) );
NAND2_X2 \AES_ENC/us21/U337  ( .A1(\AES_ENC/us21/n1100 ), .A2(\AES_ENC/us21/n617 ), .ZN(\AES_ENC/us21/n992 ) );
OR2_X2 \AES_ENC/us21/U336  ( .A1(\AES_ENC/us21/n583 ), .A2(\AES_ENC/us21/n735 ), .ZN(\AES_ENC/us21/n737 ) );
NAND2_X2 \AES_ENC/us21/U334  ( .A1(\AES_ENC/us21/n605 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n753 ) );
NAND2_X2 \AES_ENC/us21/U333  ( .A1(\AES_ENC/us21/n603 ), .A2(\AES_ENC/us21/n753 ), .ZN(\AES_ENC/us21/n1080 ) );
NAND2_X2 \AES_ENC/us21/U332  ( .A1(\AES_ENC/us21/n1048 ), .A2(\AES_ENC/us21/n602 ), .ZN(\AES_ENC/us21/n736 ) );
NAND2_X2 \AES_ENC/us21/U331  ( .A1(\AES_ENC/us21/n737 ), .A2(\AES_ENC/us21/n736 ), .ZN(\AES_ENC/us21/n739 ) );
NAND2_X2 \AES_ENC/us21/U330  ( .A1(\AES_ENC/us21/n739 ), .A2(\AES_ENC/us21/n738 ), .ZN(\AES_ENC/us21/n745 ) );
NAND2_X2 \AES_ENC/us21/U326  ( .A1(\AES_ENC/us21/n1096 ), .A2(\AES_ENC/us21/n598 ), .ZN(\AES_ENC/us21/n906 ) );
NAND4_X2 \AES_ENC/us21/U323  ( .A1(\AES_ENC/us21/n746 ), .A2(\AES_ENC/us21/n992 ), .A3(\AES_ENC/us21/n745 ), .A4(\AES_ENC/us21/n744 ), .ZN(\AES_ENC/us21/n747 ) );
NAND2_X2 \AES_ENC/us21/U322  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n747 ), .ZN(\AES_ENC/us21/n793 ) );
NAND2_X2 \AES_ENC/us21/U321  ( .A1(\AES_ENC/us21/n606 ), .A2(\AES_ENC/us21/n855 ), .ZN(\AES_ENC/us21/n748 ) );
NAND2_X2 \AES_ENC/us21/U320  ( .A1(\AES_ENC/us21/n956 ), .A2(\AES_ENC/us21/n748 ), .ZN(\AES_ENC/us21/n760 ) );
NAND2_X2 \AES_ENC/us21/U313  ( .A1(\AES_ENC/us21/n598 ), .A2(\AES_ENC/us21/n753 ), .ZN(\AES_ENC/us21/n1023 ) );
NAND4_X2 \AES_ENC/us21/U308  ( .A1(\AES_ENC/us21/n760 ), .A2(\AES_ENC/us21/n992 ), .A3(\AES_ENC/us21/n759 ), .A4(\AES_ENC/us21/n758 ), .ZN(\AES_ENC/us21/n761 ) );
NAND2_X2 \AES_ENC/us21/U307  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n761 ), .ZN(\AES_ENC/us21/n792 ) );
NAND2_X2 \AES_ENC/us21/U306  ( .A1(\AES_ENC/us21/n606 ), .A2(\AES_ENC/us21/n610 ), .ZN(\AES_ENC/us21/n989 ) );
NAND2_X2 \AES_ENC/us21/U305  ( .A1(\AES_ENC/us21/n1050 ), .A2(\AES_ENC/us21/n989 ), .ZN(\AES_ENC/us21/n777 ) );
NAND2_X2 \AES_ENC/us21/U304  ( .A1(\AES_ENC/us21/n1093 ), .A2(\AES_ENC/us21/n762 ), .ZN(\AES_ENC/us21/n776 ) );
XNOR2_X2 \AES_ENC/us21/U301  ( .A(\AES_ENC/sa21 [7]), .B(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n959 ) );
NAND4_X2 \AES_ENC/us21/U289  ( .A1(\AES_ENC/us21/n777 ), .A2(\AES_ENC/us21/n776 ), .A3(\AES_ENC/us21/n775 ), .A4(\AES_ENC/us21/n774 ), .ZN(\AES_ENC/us21/n778 ) );
NAND2_X2 \AES_ENC/us21/U288  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n778 ), .ZN(\AES_ENC/us21/n791 ) );
NAND2_X2 \AES_ENC/us21/U287  ( .A1(\AES_ENC/us21/n1056 ), .A2(\AES_ENC/us21/n1050 ), .ZN(\AES_ENC/us21/n788 ) );
NAND2_X2 \AES_ENC/us21/U286  ( .A1(\AES_ENC/us21/n1091 ), .A2(\AES_ENC/us21/n779 ), .ZN(\AES_ENC/us21/n787 ) );
NAND2_X2 \AES_ENC/us21/U285  ( .A1(\AES_ENC/us21/n956 ), .A2(\AES_ENC/sa21 [1]), .ZN(\AES_ENC/us21/n786 ) );
NAND4_X2 \AES_ENC/us21/U278  ( .A1(\AES_ENC/us21/n788 ), .A2(\AES_ENC/us21/n787 ), .A3(\AES_ENC/us21/n786 ), .A4(\AES_ENC/us21/n785 ), .ZN(\AES_ENC/us21/n789 ) );
NAND2_X2 \AES_ENC/us21/U277  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n789 ), .ZN(\AES_ENC/us21/n790 ) );
NAND4_X2 \AES_ENC/us21/U276  ( .A1(\AES_ENC/us21/n793 ), .A2(\AES_ENC/us21/n792 ), .A3(\AES_ENC/us21/n791 ), .A4(\AES_ENC/us21/n790 ), .ZN(\AES_ENC/sa21_sub[2] ) );
NAND2_X2 \AES_ENC/us21/U275  ( .A1(\AES_ENC/us21/n1059 ), .A2(\AES_ENC/us21/n794 ), .ZN(\AES_ENC/us21/n810 ) );
NAND2_X2 \AES_ENC/us21/U274  ( .A1(\AES_ENC/us21/n1049 ), .A2(\AES_ENC/us21/n956 ), .ZN(\AES_ENC/us21/n809 ) );
OR2_X2 \AES_ENC/us21/U266  ( .A1(\AES_ENC/us21/n1096 ), .A2(\AES_ENC/us21/n578 ), .ZN(\AES_ENC/us21/n802 ) );
NAND2_X2 \AES_ENC/us21/U265  ( .A1(\AES_ENC/us21/n1053 ), .A2(\AES_ENC/us21/n800 ), .ZN(\AES_ENC/us21/n801 ) );
NAND2_X2 \AES_ENC/us21/U264  ( .A1(\AES_ENC/us21/n802 ), .A2(\AES_ENC/us21/n801 ), .ZN(\AES_ENC/us21/n805 ) );
NAND4_X2 \AES_ENC/us21/U261  ( .A1(\AES_ENC/us21/n810 ), .A2(\AES_ENC/us21/n809 ), .A3(\AES_ENC/us21/n808 ), .A4(\AES_ENC/us21/n807 ), .ZN(\AES_ENC/us21/n811 ) );
NAND2_X2 \AES_ENC/us21/U260  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n811 ), .ZN(\AES_ENC/us21/n852 ) );
OR2_X2 \AES_ENC/us21/U259  ( .A1(\AES_ENC/us21/n1023 ), .A2(\AES_ENC/us21/n591 ), .ZN(\AES_ENC/us21/n819 ) );
OR2_X2 \AES_ENC/us21/U257  ( .A1(\AES_ENC/us21/n570 ), .A2(\AES_ENC/us21/n930 ), .ZN(\AES_ENC/us21/n818 ) );
NAND2_X2 \AES_ENC/us21/U256  ( .A1(\AES_ENC/us21/n1013 ), .A2(\AES_ENC/us21/n1094 ), .ZN(\AES_ENC/us21/n817 ) );
NAND4_X2 \AES_ENC/us21/U249  ( .A1(\AES_ENC/us21/n819 ), .A2(\AES_ENC/us21/n818 ), .A3(\AES_ENC/us21/n817 ), .A4(\AES_ENC/us21/n816 ), .ZN(\AES_ENC/us21/n820 ) );
NAND2_X2 \AES_ENC/us21/U248  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n820 ), .ZN(\AES_ENC/us21/n851 ) );
NAND2_X2 \AES_ENC/us21/U247  ( .A1(\AES_ENC/us21/n956 ), .A2(\AES_ENC/us21/n1080 ), .ZN(\AES_ENC/us21/n835 ) );
NAND2_X2 \AES_ENC/us21/U246  ( .A1(\AES_ENC/us21/n570 ), .A2(\AES_ENC/us21/n1030 ), .ZN(\AES_ENC/us21/n1047 ) );
OR2_X2 \AES_ENC/us21/U245  ( .A1(\AES_ENC/us21/n1047 ), .A2(\AES_ENC/us21/n585 ), .ZN(\AES_ENC/us21/n834 ) );
NAND2_X2 \AES_ENC/us21/U244  ( .A1(\AES_ENC/us21/n1072 ), .A2(\AES_ENC/us21/n620 ), .ZN(\AES_ENC/us21/n833 ) );
NAND4_X2 \AES_ENC/us21/U233  ( .A1(\AES_ENC/us21/n835 ), .A2(\AES_ENC/us21/n834 ), .A3(\AES_ENC/us21/n833 ), .A4(\AES_ENC/us21/n832 ), .ZN(\AES_ENC/us21/n836 ) );
NAND2_X2 \AES_ENC/us21/U232  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n836 ), .ZN(\AES_ENC/us21/n850 ) );
NAND2_X2 \AES_ENC/us21/U231  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n601 ), .ZN(\AES_ENC/us21/n847 ) );
NAND2_X2 \AES_ENC/us21/U230  ( .A1(\AES_ENC/us21/n1050 ), .A2(\AES_ENC/us21/n1071 ), .ZN(\AES_ENC/us21/n846 ) );
OR2_X2 \AES_ENC/us21/U224  ( .A1(\AES_ENC/us21/n1053 ), .A2(\AES_ENC/us21/n911 ), .ZN(\AES_ENC/us21/n1077 ) );
NAND4_X2 \AES_ENC/us21/U220  ( .A1(\AES_ENC/us21/n847 ), .A2(\AES_ENC/us21/n846 ), .A3(\AES_ENC/us21/n845 ), .A4(\AES_ENC/us21/n844 ), .ZN(\AES_ENC/us21/n848 ) );
NAND2_X2 \AES_ENC/us21/U219  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n848 ), .ZN(\AES_ENC/us21/n849 ) );
NAND4_X2 \AES_ENC/us21/U218  ( .A1(\AES_ENC/us21/n852 ), .A2(\AES_ENC/us21/n851 ), .A3(\AES_ENC/us21/n850 ), .A4(\AES_ENC/us21/n849 ), .ZN(\AES_ENC/sa21_sub[3] ) );
NAND2_X2 \AES_ENC/us21/U216  ( .A1(\AES_ENC/us21/n1009 ), .A2(\AES_ENC/us21/n1072 ), .ZN(\AES_ENC/us21/n862 ) );
NAND2_X2 \AES_ENC/us21/U215  ( .A1(\AES_ENC/us21/n610 ), .A2(\AES_ENC/us21/n618 ), .ZN(\AES_ENC/us21/n853 ) );
NAND2_X2 \AES_ENC/us21/U214  ( .A1(\AES_ENC/us21/n1050 ), .A2(\AES_ENC/us21/n853 ), .ZN(\AES_ENC/us21/n861 ) );
NAND4_X2 \AES_ENC/us21/U206  ( .A1(\AES_ENC/us21/n862 ), .A2(\AES_ENC/us21/n861 ), .A3(\AES_ENC/us21/n860 ), .A4(\AES_ENC/us21/n859 ), .ZN(\AES_ENC/us21/n863 ) );
NAND2_X2 \AES_ENC/us21/U205  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n863 ), .ZN(\AES_ENC/us21/n905 ) );
NAND2_X2 \AES_ENC/us21/U204  ( .A1(\AES_ENC/us21/n1010 ), .A2(\AES_ENC/us21/n989 ), .ZN(\AES_ENC/us21/n874 ) );
NAND2_X2 \AES_ENC/us21/U203  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n583 ), .ZN(\AES_ENC/us21/n864 ) );
NAND2_X2 \AES_ENC/us21/U202  ( .A1(\AES_ENC/us21/n929 ), .A2(\AES_ENC/us21/n864 ), .ZN(\AES_ENC/us21/n873 ) );
NAND4_X2 \AES_ENC/us21/U193  ( .A1(\AES_ENC/us21/n874 ), .A2(\AES_ENC/us21/n873 ), .A3(\AES_ENC/us21/n872 ), .A4(\AES_ENC/us21/n871 ), .ZN(\AES_ENC/us21/n875 ) );
NAND2_X2 \AES_ENC/us21/U192  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n875 ), .ZN(\AES_ENC/us21/n904 ) );
NAND2_X2 \AES_ENC/us21/U191  ( .A1(\AES_ENC/us21/n597 ), .A2(\AES_ENC/us21/n1050 ), .ZN(\AES_ENC/us21/n889 ) );
NAND2_X2 \AES_ENC/us21/U190  ( .A1(\AES_ENC/us21/n1093 ), .A2(\AES_ENC/us21/n617 ), .ZN(\AES_ENC/us21/n876 ) );
NAND2_X2 \AES_ENC/us21/U189  ( .A1(\AES_ENC/us21/n576 ), .A2(\AES_ENC/us21/n876 ), .ZN(\AES_ENC/us21/n877 ) );
NAND2_X2 \AES_ENC/us21/U188  ( .A1(\AES_ENC/us21/n877 ), .A2(\AES_ENC/us21/n601 ), .ZN(\AES_ENC/us21/n888 ) );
NAND4_X2 \AES_ENC/us21/U179  ( .A1(\AES_ENC/us21/n889 ), .A2(\AES_ENC/us21/n888 ), .A3(\AES_ENC/us21/n887 ), .A4(\AES_ENC/us21/n886 ), .ZN(\AES_ENC/us21/n890 ) );
NAND2_X2 \AES_ENC/us21/U178  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n890 ), .ZN(\AES_ENC/us21/n903 ) );
OR2_X2 \AES_ENC/us21/U177  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n1059 ), .ZN(\AES_ENC/us21/n900 ) );
NAND2_X2 \AES_ENC/us21/U176  ( .A1(\AES_ENC/us21/n1073 ), .A2(\AES_ENC/us21/n1047 ), .ZN(\AES_ENC/us21/n899 ) );
NAND2_X2 \AES_ENC/us21/U175  ( .A1(\AES_ENC/us21/n1094 ), .A2(\AES_ENC/us21/n608 ), .ZN(\AES_ENC/us21/n898 ) );
NAND4_X2 \AES_ENC/us21/U167  ( .A1(\AES_ENC/us21/n900 ), .A2(\AES_ENC/us21/n899 ), .A3(\AES_ENC/us21/n898 ), .A4(\AES_ENC/us21/n897 ), .ZN(\AES_ENC/us21/n901 ) );
NAND2_X2 \AES_ENC/us21/U166  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n901 ), .ZN(\AES_ENC/us21/n902 ) );
NAND4_X2 \AES_ENC/us21/U165  ( .A1(\AES_ENC/us21/n905 ), .A2(\AES_ENC/us21/n904 ), .A3(\AES_ENC/us21/n903 ), .A4(\AES_ENC/us21/n902 ), .ZN(\AES_ENC/sa21_sub[4] ) );
NAND2_X2 \AES_ENC/us21/U164  ( .A1(\AES_ENC/us21/n1094 ), .A2(\AES_ENC/us21/n615 ), .ZN(\AES_ENC/us21/n922 ) );
NAND2_X2 \AES_ENC/us21/U163  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n989 ), .ZN(\AES_ENC/us21/n921 ) );
NAND4_X2 \AES_ENC/us21/U151  ( .A1(\AES_ENC/us21/n922 ), .A2(\AES_ENC/us21/n921 ), .A3(\AES_ENC/us21/n920 ), .A4(\AES_ENC/us21/n919 ), .ZN(\AES_ENC/us21/n923 ) );
NAND2_X2 \AES_ENC/us21/U150  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n923 ), .ZN(\AES_ENC/us21/n972 ) );
NAND2_X2 \AES_ENC/us21/U149  ( .A1(\AES_ENC/us21/n603 ), .A2(\AES_ENC/us21/n605 ), .ZN(\AES_ENC/us21/n924 ) );
NAND2_X2 \AES_ENC/us21/U148  ( .A1(\AES_ENC/us21/n1073 ), .A2(\AES_ENC/us21/n924 ), .ZN(\AES_ENC/us21/n939 ) );
NAND2_X2 \AES_ENC/us21/U147  ( .A1(\AES_ENC/us21/n926 ), .A2(\AES_ENC/us21/n925 ), .ZN(\AES_ENC/us21/n927 ) );
NAND2_X2 \AES_ENC/us21/U146  ( .A1(\AES_ENC/us21/n578 ), .A2(\AES_ENC/us21/n927 ), .ZN(\AES_ENC/us21/n928 ) );
NAND2_X2 \AES_ENC/us21/U145  ( .A1(\AES_ENC/us21/n928 ), .A2(\AES_ENC/us21/n1080 ), .ZN(\AES_ENC/us21/n938 ) );
OR2_X2 \AES_ENC/us21/U144  ( .A1(\AES_ENC/us21/n1117 ), .A2(\AES_ENC/us21/n589 ), .ZN(\AES_ENC/us21/n937 ) );
NAND4_X2 \AES_ENC/us21/U139  ( .A1(\AES_ENC/us21/n939 ), .A2(\AES_ENC/us21/n938 ), .A3(\AES_ENC/us21/n937 ), .A4(\AES_ENC/us21/n936 ), .ZN(\AES_ENC/us21/n940 ) );
NAND2_X2 \AES_ENC/us21/U138  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n940 ), .ZN(\AES_ENC/us21/n971 ) );
OR2_X2 \AES_ENC/us21/U137  ( .A1(\AES_ENC/us21/n577 ), .A2(\AES_ENC/us21/n941 ), .ZN(\AES_ENC/us21/n954 ) );
NAND2_X2 \AES_ENC/us21/U136  ( .A1(\AES_ENC/us21/n1096 ), .A2(\AES_ENC/us21/n618 ), .ZN(\AES_ENC/us21/n942 ) );
NAND2_X2 \AES_ENC/us21/U135  ( .A1(\AES_ENC/us21/n1048 ), .A2(\AES_ENC/us21/n942 ), .ZN(\AES_ENC/us21/n943 ) );
NAND2_X2 \AES_ENC/us21/U134  ( .A1(\AES_ENC/us21/n585 ), .A2(\AES_ENC/us21/n943 ), .ZN(\AES_ENC/us21/n944 ) );
NAND2_X2 \AES_ENC/us21/U133  ( .A1(\AES_ENC/us21/n944 ), .A2(\AES_ENC/us21/n599 ), .ZN(\AES_ENC/us21/n953 ) );
NAND4_X2 \AES_ENC/us21/U125  ( .A1(\AES_ENC/us21/n954 ), .A2(\AES_ENC/us21/n953 ), .A3(\AES_ENC/us21/n952 ), .A4(\AES_ENC/us21/n951 ), .ZN(\AES_ENC/us21/n955 ) );
NAND2_X2 \AES_ENC/us21/U124  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n955 ), .ZN(\AES_ENC/us21/n970 ) );
NAND2_X2 \AES_ENC/us21/U123  ( .A1(\AES_ENC/us21/n1094 ), .A2(\AES_ENC/us21/n1071 ), .ZN(\AES_ENC/us21/n967 ) );
NAND2_X2 \AES_ENC/us21/U122  ( .A1(\AES_ENC/us21/n956 ), .A2(\AES_ENC/us21/n1030 ), .ZN(\AES_ENC/us21/n966 ) );
NAND4_X2 \AES_ENC/us21/U114  ( .A1(\AES_ENC/us21/n967 ), .A2(\AES_ENC/us21/n966 ), .A3(\AES_ENC/us21/n965 ), .A4(\AES_ENC/us21/n964 ), .ZN(\AES_ENC/us21/n968 ) );
NAND2_X2 \AES_ENC/us21/U113  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n968 ), .ZN(\AES_ENC/us21/n969 ) );
NAND4_X2 \AES_ENC/us21/U112  ( .A1(\AES_ENC/us21/n972 ), .A2(\AES_ENC/us21/n971 ), .A3(\AES_ENC/us21/n970 ), .A4(\AES_ENC/us21/n969 ), .ZN(\AES_ENC/sa21_sub[5] ) );
NAND2_X2 \AES_ENC/us21/U111  ( .A1(\AES_ENC/us21/n570 ), .A2(\AES_ENC/us21/n1097 ), .ZN(\AES_ENC/us21/n973 ) );
NAND2_X2 \AES_ENC/us21/U110  ( .A1(\AES_ENC/us21/n1073 ), .A2(\AES_ENC/us21/n973 ), .ZN(\AES_ENC/us21/n987 ) );
NAND2_X2 \AES_ENC/us21/U109  ( .A1(\AES_ENC/us21/n974 ), .A2(\AES_ENC/us21/n1077 ), .ZN(\AES_ENC/us21/n975 ) );
NAND2_X2 \AES_ENC/us21/U108  ( .A1(\AES_ENC/us21/n587 ), .A2(\AES_ENC/us21/n975 ), .ZN(\AES_ENC/us21/n976 ) );
NAND2_X2 \AES_ENC/us21/U107  ( .A1(\AES_ENC/us21/n977 ), .A2(\AES_ENC/us21/n976 ), .ZN(\AES_ENC/us21/n986 ) );
NAND4_X2 \AES_ENC/us21/U99  ( .A1(\AES_ENC/us21/n987 ), .A2(\AES_ENC/us21/n986 ), .A3(\AES_ENC/us21/n985 ), .A4(\AES_ENC/us21/n984 ), .ZN(\AES_ENC/us21/n988 ) );
NAND2_X2 \AES_ENC/us21/U98  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n988 ), .ZN(\AES_ENC/us21/n1044 ) );
NAND2_X2 \AES_ENC/us21/U97  ( .A1(\AES_ENC/us21/n1073 ), .A2(\AES_ENC/us21/n989 ), .ZN(\AES_ENC/us21/n1004 ) );
NAND2_X2 \AES_ENC/us21/U96  ( .A1(\AES_ENC/us21/n1092 ), .A2(\AES_ENC/us21/n605 ), .ZN(\AES_ENC/us21/n1003 ) );
NAND4_X2 \AES_ENC/us21/U85  ( .A1(\AES_ENC/us21/n1004 ), .A2(\AES_ENC/us21/n1003 ), .A3(\AES_ENC/us21/n1002 ), .A4(\AES_ENC/us21/n1001 ), .ZN(\AES_ENC/us21/n1005 ) );
NAND2_X2 \AES_ENC/us21/U84  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n1005 ), .ZN(\AES_ENC/us21/n1043 ) );
NAND2_X2 \AES_ENC/us21/U83  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n626 ), .ZN(\AES_ENC/us21/n1020 ) );
NAND2_X2 \AES_ENC/us21/U82  ( .A1(\AES_ENC/us21/n1050 ), .A2(\AES_ENC/us21/n612 ), .ZN(\AES_ENC/us21/n1019 ) );
NAND2_X2 \AES_ENC/us21/U77  ( .A1(\AES_ENC/us21/n1059 ), .A2(\AES_ENC/us21/n1114 ), .ZN(\AES_ENC/us21/n1012 ) );
NAND2_X2 \AES_ENC/us21/U76  ( .A1(\AES_ENC/us21/n1010 ), .A2(\AES_ENC/us21/n604 ), .ZN(\AES_ENC/us21/n1011 ) );
NAND2_X2 \AES_ENC/us21/U75  ( .A1(\AES_ENC/us21/n1012 ), .A2(\AES_ENC/us21/n1011 ), .ZN(\AES_ENC/us21/n1016 ) );
NAND4_X2 \AES_ENC/us21/U70  ( .A1(\AES_ENC/us21/n1020 ), .A2(\AES_ENC/us21/n1019 ), .A3(\AES_ENC/us21/n1018 ), .A4(\AES_ENC/us21/n1017 ), .ZN(\AES_ENC/us21/n1021 ) );
NAND2_X2 \AES_ENC/us21/U69  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n1021 ), .ZN(\AES_ENC/us21/n1042 ) );
NAND2_X2 \AES_ENC/us21/U68  ( .A1(\AES_ENC/us21/n1022 ), .A2(\AES_ENC/us21/n1093 ), .ZN(\AES_ENC/us21/n1039 ) );
NAND2_X2 \AES_ENC/us21/U67  ( .A1(\AES_ENC/us21/n1050 ), .A2(\AES_ENC/us21/n1023 ), .ZN(\AES_ENC/us21/n1038 ) );
NAND2_X2 \AES_ENC/us21/U66  ( .A1(\AES_ENC/us21/n1024 ), .A2(\AES_ENC/us21/n1071 ), .ZN(\AES_ENC/us21/n1037 ) );
AND2_X2 \AES_ENC/us21/U60  ( .A1(\AES_ENC/us21/n1030 ), .A2(\AES_ENC/us21/n621 ), .ZN(\AES_ENC/us21/n1078 ) );
NAND4_X2 \AES_ENC/us21/U56  ( .A1(\AES_ENC/us21/n1039 ), .A2(\AES_ENC/us21/n1038 ), .A3(\AES_ENC/us21/n1037 ), .A4(\AES_ENC/us21/n1036 ), .ZN(\AES_ENC/us21/n1040 ) );
NAND2_X2 \AES_ENC/us21/U55  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n1040 ), .ZN(\AES_ENC/us21/n1041 ) );
NAND4_X2 \AES_ENC/us21/U54  ( .A1(\AES_ENC/us21/n1044 ), .A2(\AES_ENC/us21/n1043 ), .A3(\AES_ENC/us21/n1042 ), .A4(\AES_ENC/us21/n1041 ), .ZN(\AES_ENC/sa21_sub[6] ) );
NAND2_X2 \AES_ENC/us21/U53  ( .A1(\AES_ENC/us21/n1072 ), .A2(\AES_ENC/us21/n1045 ), .ZN(\AES_ENC/us21/n1068 ) );
NAND2_X2 \AES_ENC/us21/U52  ( .A1(\AES_ENC/us21/n1046 ), .A2(\AES_ENC/us21/n603 ), .ZN(\AES_ENC/us21/n1067 ) );
NAND2_X2 \AES_ENC/us21/U51  ( .A1(\AES_ENC/us21/n1094 ), .A2(\AES_ENC/us21/n1047 ), .ZN(\AES_ENC/us21/n1066 ) );
NAND4_X2 \AES_ENC/us21/U40  ( .A1(\AES_ENC/us21/n1068 ), .A2(\AES_ENC/us21/n1067 ), .A3(\AES_ENC/us21/n1066 ), .A4(\AES_ENC/us21/n1065 ), .ZN(\AES_ENC/us21/n1069 ) );
NAND2_X2 \AES_ENC/us21/U39  ( .A1(\AES_ENC/us21/n1070 ), .A2(\AES_ENC/us21/n1069 ), .ZN(\AES_ENC/us21/n1135 ) );
NAND2_X2 \AES_ENC/us21/U38  ( .A1(\AES_ENC/us21/n1072 ), .A2(\AES_ENC/us21/n1071 ), .ZN(\AES_ENC/us21/n1088 ) );
NAND2_X2 \AES_ENC/us21/U37  ( .A1(\AES_ENC/us21/n1073 ), .A2(\AES_ENC/us21/n608 ), .ZN(\AES_ENC/us21/n1087 ) );
NAND4_X2 \AES_ENC/us21/U28  ( .A1(\AES_ENC/us21/n1088 ), .A2(\AES_ENC/us21/n1087 ), .A3(\AES_ENC/us21/n1086 ), .A4(\AES_ENC/us21/n1085 ), .ZN(\AES_ENC/us21/n1089 ) );
NAND2_X2 \AES_ENC/us21/U27  ( .A1(\AES_ENC/us21/n1090 ), .A2(\AES_ENC/us21/n1089 ), .ZN(\AES_ENC/us21/n1134 ) );
NAND2_X2 \AES_ENC/us21/U26  ( .A1(\AES_ENC/us21/n1091 ), .A2(\AES_ENC/us21/n1093 ), .ZN(\AES_ENC/us21/n1111 ) );
NAND2_X2 \AES_ENC/us21/U25  ( .A1(\AES_ENC/us21/n1092 ), .A2(\AES_ENC/us21/n1120 ), .ZN(\AES_ENC/us21/n1110 ) );
AND2_X2 \AES_ENC/us21/U22  ( .A1(\AES_ENC/us21/n1097 ), .A2(\AES_ENC/us21/n1096 ), .ZN(\AES_ENC/us21/n1098 ) );
NAND4_X2 \AES_ENC/us21/U14  ( .A1(\AES_ENC/us21/n1111 ), .A2(\AES_ENC/us21/n1110 ), .A3(\AES_ENC/us21/n1109 ), .A4(\AES_ENC/us21/n1108 ), .ZN(\AES_ENC/us21/n1112 ) );
NAND2_X2 \AES_ENC/us21/U13  ( .A1(\AES_ENC/us21/n1113 ), .A2(\AES_ENC/us21/n1112 ), .ZN(\AES_ENC/us21/n1133 ) );
NAND2_X2 \AES_ENC/us21/U12  ( .A1(\AES_ENC/us21/n1115 ), .A2(\AES_ENC/us21/n1114 ), .ZN(\AES_ENC/us21/n1129 ) );
OR2_X2 \AES_ENC/us21/U11  ( .A1(\AES_ENC/us21/n581 ), .A2(\AES_ENC/us21/n1116 ), .ZN(\AES_ENC/us21/n1128 ) );
NAND4_X2 \AES_ENC/us21/U3  ( .A1(\AES_ENC/us21/n1129 ), .A2(\AES_ENC/us21/n1128 ), .A3(\AES_ENC/us21/n1127 ), .A4(\AES_ENC/us21/n1126 ), .ZN(\AES_ENC/us21/n1130 ) );
NAND2_X2 \AES_ENC/us21/U2  ( .A1(\AES_ENC/us21/n1131 ), .A2(\AES_ENC/us21/n1130 ), .ZN(\AES_ENC/us21/n1132 ) );
NAND4_X2 \AES_ENC/us21/U1  ( .A1(\AES_ENC/us21/n1135 ), .A2(\AES_ENC/us21/n1134 ), .A3(\AES_ENC/us21/n1133 ), .A4(\AES_ENC/us21/n1132 ), .ZN(\AES_ENC/sa21_sub[7] ) );
INV_X4 \AES_ENC/us22/U575  ( .A(\AES_ENC/sa22 [7]), .ZN(\AES_ENC/us22/n627 ));
INV_X4 \AES_ENC/us22/U574  ( .A(\AES_ENC/us22/n1114 ), .ZN(\AES_ENC/us22/n625 ) );
INV_X4 \AES_ENC/us22/U573  ( .A(\AES_ENC/sa22 [4]), .ZN(\AES_ENC/us22/n624 ));
INV_X4 \AES_ENC/us22/U572  ( .A(\AES_ENC/us22/n1025 ), .ZN(\AES_ENC/us22/n622 ) );
INV_X4 \AES_ENC/us22/U571  ( .A(\AES_ENC/us22/n1120 ), .ZN(\AES_ENC/us22/n620 ) );
INV_X4 \AES_ENC/us22/U570  ( .A(\AES_ENC/us22/n1121 ), .ZN(\AES_ENC/us22/n619 ) );
INV_X4 \AES_ENC/us22/U569  ( .A(\AES_ENC/us22/n1048 ), .ZN(\AES_ENC/us22/n618 ) );
INV_X4 \AES_ENC/us22/U568  ( .A(\AES_ENC/us22/n974 ), .ZN(\AES_ENC/us22/n616 ) );
INV_X4 \AES_ENC/us22/U567  ( .A(\AES_ENC/us22/n794 ), .ZN(\AES_ENC/us22/n614 ) );
INV_X4 \AES_ENC/us22/U566  ( .A(\AES_ENC/sa22 [2]), .ZN(\AES_ENC/us22/n611 ));
INV_X4 \AES_ENC/us22/U565  ( .A(\AES_ENC/us22/n800 ), .ZN(\AES_ENC/us22/n610 ) );
INV_X4 \AES_ENC/us22/U564  ( .A(\AES_ENC/us22/n925 ), .ZN(\AES_ENC/us22/n609 ) );
INV_X4 \AES_ENC/us22/U563  ( .A(\AES_ENC/us22/n779 ), .ZN(\AES_ENC/us22/n607 ) );
INV_X4 \AES_ENC/us22/U562  ( .A(\AES_ENC/us22/n1022 ), .ZN(\AES_ENC/us22/n603 ) );
INV_X4 \AES_ENC/us22/U561  ( .A(\AES_ENC/us22/n1102 ), .ZN(\AES_ENC/us22/n602 ) );
INV_X4 \AES_ENC/us22/U560  ( .A(\AES_ENC/us22/n929 ), .ZN(\AES_ENC/us22/n601 ) );
INV_X4 \AES_ENC/us22/U559  ( .A(\AES_ENC/us22/n1056 ), .ZN(\AES_ENC/us22/n600 ) );
INV_X4 \AES_ENC/us22/U558  ( .A(\AES_ENC/us22/n1054 ), .ZN(\AES_ENC/us22/n599 ) );
INV_X4 \AES_ENC/us22/U557  ( .A(\AES_ENC/us22/n881 ), .ZN(\AES_ENC/us22/n598 ) );
INV_X4 \AES_ENC/us22/U556  ( .A(\AES_ENC/us22/n926 ), .ZN(\AES_ENC/us22/n597 ) );
INV_X4 \AES_ENC/us22/U555  ( .A(\AES_ENC/us22/n977 ), .ZN(\AES_ENC/us22/n595 ) );
INV_X4 \AES_ENC/us22/U554  ( .A(\AES_ENC/us22/n1031 ), .ZN(\AES_ENC/us22/n594 ) );
INV_X4 \AES_ENC/us22/U553  ( .A(\AES_ENC/us22/n1103 ), .ZN(\AES_ENC/us22/n593 ) );
INV_X4 \AES_ENC/us22/U552  ( .A(\AES_ENC/us22/n1009 ), .ZN(\AES_ENC/us22/n592 ) );
INV_X4 \AES_ENC/us22/U551  ( .A(\AES_ENC/us22/n990 ), .ZN(\AES_ENC/us22/n591 ) );
INV_X4 \AES_ENC/us22/U550  ( .A(\AES_ENC/us22/n1058 ), .ZN(\AES_ENC/us22/n590 ) );
INV_X4 \AES_ENC/us22/U549  ( .A(\AES_ENC/us22/n1074 ), .ZN(\AES_ENC/us22/n589 ) );
INV_X4 \AES_ENC/us22/U548  ( .A(\AES_ENC/us22/n1053 ), .ZN(\AES_ENC/us22/n588 ) );
INV_X4 \AES_ENC/us22/U547  ( .A(\AES_ENC/us22/n826 ), .ZN(\AES_ENC/us22/n587 ) );
INV_X4 \AES_ENC/us22/U546  ( .A(\AES_ENC/us22/n992 ), .ZN(\AES_ENC/us22/n586 ) );
INV_X4 \AES_ENC/us22/U545  ( .A(\AES_ENC/us22/n821 ), .ZN(\AES_ENC/us22/n585 ) );
INV_X4 \AES_ENC/us22/U544  ( .A(\AES_ENC/us22/n910 ), .ZN(\AES_ENC/us22/n584 ) );
INV_X4 \AES_ENC/us22/U543  ( .A(\AES_ENC/us22/n906 ), .ZN(\AES_ENC/us22/n583 ) );
INV_X4 \AES_ENC/us22/U542  ( .A(\AES_ENC/us22/n880 ), .ZN(\AES_ENC/us22/n581 ) );
INV_X4 \AES_ENC/us22/U541  ( .A(\AES_ENC/us22/n1013 ), .ZN(\AES_ENC/us22/n580 ) );
INV_X4 \AES_ENC/us22/U540  ( .A(\AES_ENC/us22/n1092 ), .ZN(\AES_ENC/us22/n579 ) );
INV_X4 \AES_ENC/us22/U539  ( .A(\AES_ENC/us22/n824 ), .ZN(\AES_ENC/us22/n578 ) );
INV_X4 \AES_ENC/us22/U538  ( .A(\AES_ENC/us22/n1091 ), .ZN(\AES_ENC/us22/n577 ) );
INV_X4 \AES_ENC/us22/U537  ( .A(\AES_ENC/us22/n1080 ), .ZN(\AES_ENC/us22/n576 ) );
INV_X4 \AES_ENC/us22/U536  ( .A(\AES_ENC/us22/n959 ), .ZN(\AES_ENC/us22/n575 ) );
INV_X4 \AES_ENC/us22/U535  ( .A(\AES_ENC/sa22 [0]), .ZN(\AES_ENC/us22/n574 ));
NOR2_X2 \AES_ENC/us22/U534  ( .A1(\AES_ENC/sa22 [0]), .A2(\AES_ENC/sa22 [6]),.ZN(\AES_ENC/us22/n1090 ) );
NOR2_X2 \AES_ENC/us22/U533  ( .A1(\AES_ENC/us22/n574 ), .A2(\AES_ENC/sa22 [6]), .ZN(\AES_ENC/us22/n1070 ) );
NOR2_X2 \AES_ENC/us22/U532  ( .A1(\AES_ENC/sa22 [4]), .A2(\AES_ENC/sa22 [3]),.ZN(\AES_ENC/us22/n1025 ) );
INV_X4 \AES_ENC/us22/U531  ( .A(\AES_ENC/us22/n569 ), .ZN(\AES_ENC/us22/n572 ) );
NOR2_X2 \AES_ENC/us22/U530  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n765 ) );
NOR2_X2 \AES_ENC/us22/U529  ( .A1(\AES_ENC/sa22 [4]), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n764 ) );
NOR2_X2 \AES_ENC/us22/U528  ( .A1(\AES_ENC/us22/n765 ), .A2(\AES_ENC/us22/n764 ), .ZN(\AES_ENC/us22/n766 ) );
NOR2_X2 \AES_ENC/us22/U527  ( .A1(\AES_ENC/us22/n766 ), .A2(\AES_ENC/us22/n575 ), .ZN(\AES_ENC/us22/n767 ) );
INV_X4 \AES_ENC/us22/U526  ( .A(\AES_ENC/sa22 [3]), .ZN(\AES_ENC/us22/n621 ));
NAND3_X2 \AES_ENC/us22/U525  ( .A1(\AES_ENC/us22/n652 ), .A2(\AES_ENC/us22/n626 ), .A3(\AES_ENC/sa22 [7]), .ZN(\AES_ENC/us22/n653 ));
NOR2_X2 \AES_ENC/us22/U524  ( .A1(\AES_ENC/us22/n611 ), .A2(\AES_ENC/sa22 [5]), .ZN(\AES_ENC/us22/n925 ) );
NOR2_X2 \AES_ENC/us22/U523  ( .A1(\AES_ENC/sa22 [5]), .A2(\AES_ENC/sa22 [2]),.ZN(\AES_ENC/us22/n974 ) );
INV_X4 \AES_ENC/us22/U522  ( .A(\AES_ENC/sa22 [5]), .ZN(\AES_ENC/us22/n626 ));
NOR2_X2 \AES_ENC/us22/U521  ( .A1(\AES_ENC/us22/n611 ), .A2(\AES_ENC/sa22 [7]), .ZN(\AES_ENC/us22/n779 ) );
NAND3_X2 \AES_ENC/us22/U520  ( .A1(\AES_ENC/us22/n679 ), .A2(\AES_ENC/us22/n678 ), .A3(\AES_ENC/us22/n677 ), .ZN(\AES_ENC/sa22_sub[0] ) );
NOR2_X2 \AES_ENC/us22/U519  ( .A1(\AES_ENC/us22/n626 ), .A2(\AES_ENC/sa22 [2]), .ZN(\AES_ENC/us22/n1048 ) );
NOR3_X2 \AES_ENC/us22/U518  ( .A1(\AES_ENC/us22/n627 ), .A2(\AES_ENC/sa22 [5]), .A3(\AES_ENC/us22/n704 ), .ZN(\AES_ENC/us22/n706 ));
NOR2_X2 \AES_ENC/us22/U517  ( .A1(\AES_ENC/us22/n1117 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n707 ) );
NOR2_X2 \AES_ENC/us22/U516  ( .A1(\AES_ENC/sa22 [4]), .A2(\AES_ENC/us22/n579 ), .ZN(\AES_ENC/us22/n705 ) );
NOR3_X2 \AES_ENC/us22/U515  ( .A1(\AES_ENC/us22/n707 ), .A2(\AES_ENC/us22/n706 ), .A3(\AES_ENC/us22/n705 ), .ZN(\AES_ENC/us22/n713 ) );
NOR4_X2 \AES_ENC/us22/U512  ( .A1(\AES_ENC/us22/n633 ), .A2(\AES_ENC/us22/n632 ), .A3(\AES_ENC/us22/n631 ), .A4(\AES_ENC/us22/n630 ), .ZN(\AES_ENC/us22/n634 ) );
NOR2_X2 \AES_ENC/us22/U510  ( .A1(\AES_ENC/us22/n629 ), .A2(\AES_ENC/us22/n628 ), .ZN(\AES_ENC/us22/n635 ) );
NAND3_X2 \AES_ENC/us22/U509  ( .A1(\AES_ENC/sa22 [2]), .A2(\AES_ENC/sa22 [7]), .A3(\AES_ENC/us22/n1059 ), .ZN(\AES_ENC/us22/n636 ) );
NOR2_X2 \AES_ENC/us22/U508  ( .A1(\AES_ENC/sa22 [7]), .A2(\AES_ENC/sa22 [2]),.ZN(\AES_ENC/us22/n794 ) );
NOR2_X2 \AES_ENC/us22/U507  ( .A1(\AES_ENC/sa22 [4]), .A2(\AES_ENC/sa22 [1]),.ZN(\AES_ENC/us22/n1102 ) );
NOR2_X2 \AES_ENC/us22/U506  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/sa22 [3]), .ZN(\AES_ENC/us22/n1053 ) );
NOR2_X2 \AES_ENC/us22/U505  ( .A1(\AES_ENC/us22/n607 ), .A2(\AES_ENC/sa22 [5]), .ZN(\AES_ENC/us22/n1024 ) );
NOR2_X2 \AES_ENC/us22/U504  ( .A1(\AES_ENC/us22/n625 ), .A2(\AES_ENC/sa22 [2]), .ZN(\AES_ENC/us22/n1093 ) );
NOR2_X2 \AES_ENC/us22/U503  ( .A1(\AES_ENC/us22/n614 ), .A2(\AES_ENC/sa22 [5]), .ZN(\AES_ENC/us22/n1094 ) );
NOR2_X2 \AES_ENC/us22/U502  ( .A1(\AES_ENC/us22/n624 ), .A2(\AES_ENC/sa22 [3]), .ZN(\AES_ENC/us22/n931 ) );
INV_X4 \AES_ENC/us22/U501  ( .A(\AES_ENC/us22/n570 ), .ZN(\AES_ENC/us22/n573 ) );
NOR2_X2 \AES_ENC/us22/U500  ( .A1(\AES_ENC/us22/n1053 ), .A2(\AES_ENC/us22/n1095 ), .ZN(\AES_ENC/us22/n639 ) );
NOR3_X2 \AES_ENC/us22/U499  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n573 ), .A3(\AES_ENC/us22/n1074 ), .ZN(\AES_ENC/us22/n641 ) );
NOR2_X2 \AES_ENC/us22/U498  ( .A1(\AES_ENC/us22/n639 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n640 ) );
NOR2_X2 \AES_ENC/us22/U497  ( .A1(\AES_ENC/us22/n641 ), .A2(\AES_ENC/us22/n640 ), .ZN(\AES_ENC/us22/n646 ) );
NOR3_X2 \AES_ENC/us22/U496  ( .A1(\AES_ENC/us22/n995 ), .A2(\AES_ENC/us22/n586 ), .A3(\AES_ENC/us22/n994 ), .ZN(\AES_ENC/us22/n1002 ) );
NOR2_X2 \AES_ENC/us22/U495  ( .A1(\AES_ENC/us22/n909 ), .A2(\AES_ENC/us22/n908 ), .ZN(\AES_ENC/us22/n920 ) );
NOR2_X2 \AES_ENC/us22/U494  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n823 ) );
NOR2_X2 \AES_ENC/us22/U492  ( .A1(\AES_ENC/us22/n624 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n822 ) );
NOR2_X2 \AES_ENC/us22/U491  ( .A1(\AES_ENC/us22/n823 ), .A2(\AES_ENC/us22/n822 ), .ZN(\AES_ENC/us22/n825 ) );
NOR2_X2 \AES_ENC/us22/U490  ( .A1(\AES_ENC/sa22 [1]), .A2(\AES_ENC/us22/n623 ), .ZN(\AES_ENC/us22/n913 ) );
NOR2_X2 \AES_ENC/us22/U489  ( .A1(\AES_ENC/us22/n913 ), .A2(\AES_ENC/us22/n1091 ), .ZN(\AES_ENC/us22/n914 ) );
NOR2_X2 \AES_ENC/us22/U488  ( .A1(\AES_ENC/us22/n826 ), .A2(\AES_ENC/us22/n572 ), .ZN(\AES_ENC/us22/n827 ) );
NOR3_X2 \AES_ENC/us22/U487  ( .A1(\AES_ENC/us22/n769 ), .A2(\AES_ENC/us22/n768 ), .A3(\AES_ENC/us22/n767 ), .ZN(\AES_ENC/us22/n775 ) );
NOR2_X2 \AES_ENC/us22/U486  ( .A1(\AES_ENC/us22/n1056 ), .A2(\AES_ENC/us22/n1053 ), .ZN(\AES_ENC/us22/n749 ) );
NOR2_X2 \AES_ENC/us22/U483  ( .A1(\AES_ENC/us22/n749 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n752 ) );
INV_X4 \AES_ENC/us22/U482  ( .A(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n596 ));
NOR2_X2 \AES_ENC/us22/U480  ( .A1(\AES_ENC/us22/n1054 ), .A2(\AES_ENC/us22/n1053 ), .ZN(\AES_ENC/us22/n1055 ) );
OR2_X4 \AES_ENC/us22/U479  ( .A1(\AES_ENC/us22/n1094 ), .A2(\AES_ENC/us22/n1093 ), .ZN(\AES_ENC/us22/n571 ) );
AND2_X2 \AES_ENC/us22/U478  ( .A1(\AES_ENC/us22/n571 ), .A2(\AES_ENC/us22/n1095 ), .ZN(\AES_ENC/us22/n1101 ) );
NOR2_X2 \AES_ENC/us22/U477  ( .A1(\AES_ENC/us22/n1074 ), .A2(\AES_ENC/us22/n931 ), .ZN(\AES_ENC/us22/n796 ) );
NOR2_X2 \AES_ENC/us22/U474  ( .A1(\AES_ENC/us22/n796 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n797 ) );
NOR2_X2 \AES_ENC/us22/U473  ( .A1(\AES_ENC/us22/n932 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n933 ) );
NOR2_X2 \AES_ENC/us22/U472  ( .A1(\AES_ENC/us22/n929 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n935 ) );
NOR2_X2 \AES_ENC/us22/U471  ( .A1(\AES_ENC/us22/n931 ), .A2(\AES_ENC/us22/n930 ), .ZN(\AES_ENC/us22/n934 ) );
NOR3_X2 \AES_ENC/us22/U470  ( .A1(\AES_ENC/us22/n935 ), .A2(\AES_ENC/us22/n934 ), .A3(\AES_ENC/us22/n933 ), .ZN(\AES_ENC/us22/n936 ) );
NOR2_X2 \AES_ENC/us22/U469  ( .A1(\AES_ENC/us22/n624 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n1075 ) );
NOR2_X2 \AES_ENC/us22/U468  ( .A1(\AES_ENC/us22/n572 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n949 ) );
NOR2_X2 \AES_ENC/us22/U467  ( .A1(\AES_ENC/us22/n1049 ), .A2(\AES_ENC/us22/n618 ), .ZN(\AES_ENC/us22/n1051 ) );
NOR2_X2 \AES_ENC/us22/U466  ( .A1(\AES_ENC/us22/n1051 ), .A2(\AES_ENC/us22/n1050 ), .ZN(\AES_ENC/us22/n1052 ) );
NOR2_X2 \AES_ENC/us22/U465  ( .A1(\AES_ENC/us22/n1052 ), .A2(\AES_ENC/us22/n592 ), .ZN(\AES_ENC/us22/n1064 ) );
NOR2_X2 \AES_ENC/us22/U464  ( .A1(\AES_ENC/sa22 [1]), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n631 ) );
NOR2_X2 \AES_ENC/us22/U463  ( .A1(\AES_ENC/us22/n1025 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n980 ) );
NOR2_X2 \AES_ENC/us22/U462  ( .A1(\AES_ENC/us22/n1073 ), .A2(\AES_ENC/us22/n1094 ), .ZN(\AES_ENC/us22/n795 ) );
NOR2_X2 \AES_ENC/us22/U461  ( .A1(\AES_ENC/us22/n795 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n799 ) );
NOR2_X2 \AES_ENC/us22/U460  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n981 ) );
NOR2_X2 \AES_ENC/us22/U459  ( .A1(\AES_ENC/us22/n1102 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n643 ) );
NOR2_X2 \AES_ENC/us22/U458  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n621 ), .ZN(\AES_ENC/us22/n642 ) );
NOR2_X2 \AES_ENC/us22/U455  ( .A1(\AES_ENC/us22/n911 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n644 ) );
NOR4_X2 \AES_ENC/us22/U448  ( .A1(\AES_ENC/us22/n644 ), .A2(\AES_ENC/us22/n643 ), .A3(\AES_ENC/us22/n804 ), .A4(\AES_ENC/us22/n642 ), .ZN(\AES_ENC/us22/n645 ) );
NOR2_X2 \AES_ENC/us22/U447  ( .A1(\AES_ENC/us22/n1102 ), .A2(\AES_ENC/us22/n910 ), .ZN(\AES_ENC/us22/n932 ) );
NOR2_X2 \AES_ENC/us22/U442  ( .A1(\AES_ENC/us22/n1102 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n755 ) );
NOR2_X2 \AES_ENC/us22/U441  ( .A1(\AES_ENC/us22/n931 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n743 ) );
NOR2_X2 \AES_ENC/us22/U438  ( .A1(\AES_ENC/us22/n1072 ), .A2(\AES_ENC/us22/n1094 ), .ZN(\AES_ENC/us22/n930 ) );
NOR2_X2 \AES_ENC/us22/U435  ( .A1(\AES_ENC/us22/n1074 ), .A2(\AES_ENC/us22/n1025 ), .ZN(\AES_ENC/us22/n891 ) );
NOR2_X2 \AES_ENC/us22/U434  ( .A1(\AES_ENC/us22/n891 ), .A2(\AES_ENC/us22/n609 ), .ZN(\AES_ENC/us22/n894 ) );
NOR3_X2 \AES_ENC/us22/U433  ( .A1(\AES_ENC/us22/n623 ), .A2(\AES_ENC/sa22 [1]), .A3(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n683 ));
INV_X4 \AES_ENC/us22/U428  ( .A(\AES_ENC/us22/n931 ), .ZN(\AES_ENC/us22/n623 ) );
NOR2_X2 \AES_ENC/us22/U427  ( .A1(\AES_ENC/us22/n996 ), .A2(\AES_ENC/us22/n931 ), .ZN(\AES_ENC/us22/n704 ) );
NOR2_X2 \AES_ENC/us22/U421  ( .A1(\AES_ENC/us22/n931 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n685 ) );
NOR2_X2 \AES_ENC/us22/U420  ( .A1(\AES_ENC/us22/n1029 ), .A2(\AES_ENC/us22/n1025 ), .ZN(\AES_ENC/us22/n1079 ) );
NOR3_X2 \AES_ENC/us22/U419  ( .A1(\AES_ENC/us22/n589 ), .A2(\AES_ENC/us22/n1025 ), .A3(\AES_ENC/us22/n616 ), .ZN(\AES_ENC/us22/n945 ) );
NOR2_X2 \AES_ENC/us22/U418  ( .A1(\AES_ENC/us22/n626 ), .A2(\AES_ENC/us22/n611 ), .ZN(\AES_ENC/us22/n800 ) );
NOR3_X2 \AES_ENC/us22/U417  ( .A1(\AES_ENC/us22/n590 ), .A2(\AES_ENC/us22/n627 ), .A3(\AES_ENC/us22/n611 ), .ZN(\AES_ENC/us22/n798 ) );
NOR3_X2 \AES_ENC/us22/U416  ( .A1(\AES_ENC/us22/n610 ), .A2(\AES_ENC/us22/n572 ), .A3(\AES_ENC/us22/n575 ), .ZN(\AES_ENC/us22/n962 ) );
NOR3_X2 \AES_ENC/us22/U415  ( .A1(\AES_ENC/us22/n959 ), .A2(\AES_ENC/us22/n572 ), .A3(\AES_ENC/us22/n609 ), .ZN(\AES_ENC/us22/n768 ) );
NOR3_X2 \AES_ENC/us22/U414  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n572 ), .A3(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n694 ) );
NOR3_X2 \AES_ENC/us22/U413  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n572 ), .A3(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n895 ) );
NOR3_X2 \AES_ENC/us22/U410  ( .A1(\AES_ENC/us22/n1008 ), .A2(\AES_ENC/us22/n1007 ), .A3(\AES_ENC/us22/n1006 ), .ZN(\AES_ENC/us22/n1018 ) );
NOR4_X2 \AES_ENC/us22/U409  ( .A1(\AES_ENC/us22/n806 ), .A2(\AES_ENC/us22/n805 ), .A3(\AES_ENC/us22/n804 ), .A4(\AES_ENC/us22/n803 ), .ZN(\AES_ENC/us22/n807 ) );
NOR3_X2 \AES_ENC/us22/U406  ( .A1(\AES_ENC/us22/n799 ), .A2(\AES_ENC/us22/n798 ), .A3(\AES_ENC/us22/n797 ), .ZN(\AES_ENC/us22/n808 ) );
NOR4_X2 \AES_ENC/us22/U405  ( .A1(\AES_ENC/us22/n843 ), .A2(\AES_ENC/us22/n842 ), .A3(\AES_ENC/us22/n841 ), .A4(\AES_ENC/us22/n840 ), .ZN(\AES_ENC/us22/n844 ) );
NOR2_X2 \AES_ENC/us22/U404  ( .A1(\AES_ENC/us22/n669 ), .A2(\AES_ENC/us22/n668 ), .ZN(\AES_ENC/us22/n673 ) );
NOR4_X2 \AES_ENC/us22/U403  ( .A1(\AES_ENC/us22/n946 ), .A2(\AES_ENC/us22/n1046 ), .A3(\AES_ENC/us22/n671 ), .A4(\AES_ENC/us22/n670 ), .ZN(\AES_ENC/us22/n672 ) );
NOR4_X2 \AES_ENC/us22/U401  ( .A1(\AES_ENC/us22/n711 ), .A2(\AES_ENC/us22/n710 ), .A3(\AES_ENC/us22/n709 ), .A4(\AES_ENC/us22/n708 ), .ZN(\AES_ENC/us22/n712 ) );
NOR4_X2 \AES_ENC/us22/U400  ( .A1(\AES_ENC/us22/n963 ), .A2(\AES_ENC/us22/n962 ), .A3(\AES_ENC/us22/n961 ), .A4(\AES_ENC/us22/n960 ), .ZN(\AES_ENC/us22/n964 ) );
NOR3_X2 \AES_ENC/us22/U399  ( .A1(\AES_ENC/us22/n1101 ), .A2(\AES_ENC/us22/n1100 ), .A3(\AES_ENC/us22/n1099 ), .ZN(\AES_ENC/us22/n1109 ) );
NOR3_X2 \AES_ENC/us22/U398  ( .A1(\AES_ENC/us22/n743 ), .A2(\AES_ENC/us22/n742 ), .A3(\AES_ENC/us22/n741 ), .ZN(\AES_ENC/us22/n744 ) );
NOR2_X2 \AES_ENC/us22/U397  ( .A1(\AES_ENC/us22/n697 ), .A2(\AES_ENC/us22/n658 ), .ZN(\AES_ENC/us22/n659 ) );
NOR2_X2 \AES_ENC/us22/U396  ( .A1(\AES_ENC/us22/n1078 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n1033 ) );
NOR2_X2 \AES_ENC/us22/U393  ( .A1(\AES_ENC/us22/n1031 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n1032 ) );
NOR3_X2 \AES_ENC/us22/U390  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n1025 ), .A3(\AES_ENC/us22/n1074 ), .ZN(\AES_ENC/us22/n1035 ) );
NOR4_X2 \AES_ENC/us22/U389  ( .A1(\AES_ENC/us22/n1035 ), .A2(\AES_ENC/us22/n1034 ), .A3(\AES_ENC/us22/n1033 ), .A4(\AES_ENC/us22/n1032 ), .ZN(\AES_ENC/us22/n1036 ) );
NOR2_X2 \AES_ENC/us22/U388  ( .A1(\AES_ENC/us22/n598 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n885 ) );
NOR2_X2 \AES_ENC/us22/U387  ( .A1(\AES_ENC/us22/n623 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n882 ) );
NOR2_X2 \AES_ENC/us22/U386  ( .A1(\AES_ENC/us22/n1053 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n884 ) );
NOR4_X2 \AES_ENC/us22/U385  ( .A1(\AES_ENC/us22/n885 ), .A2(\AES_ENC/us22/n884 ), .A3(\AES_ENC/us22/n883 ), .A4(\AES_ENC/us22/n882 ), .ZN(\AES_ENC/us22/n886 ) );
NOR2_X2 \AES_ENC/us22/U384  ( .A1(\AES_ENC/us22/n825 ), .A2(\AES_ENC/us22/n578 ), .ZN(\AES_ENC/us22/n830 ) );
NOR2_X2 \AES_ENC/us22/U383  ( .A1(\AES_ENC/us22/n827 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n829 ) );
NOR2_X2 \AES_ENC/us22/U382  ( .A1(\AES_ENC/us22/n572 ), .A2(\AES_ENC/us22/n579 ), .ZN(\AES_ENC/us22/n828 ) );
NOR4_X2 \AES_ENC/us22/U374  ( .A1(\AES_ENC/us22/n831 ), .A2(\AES_ENC/us22/n830 ), .A3(\AES_ENC/us22/n829 ), .A4(\AES_ENC/us22/n828 ), .ZN(\AES_ENC/us22/n832 ) );
NOR2_X2 \AES_ENC/us22/U373  ( .A1(\AES_ENC/us22/n606 ), .A2(\AES_ENC/us22/n582 ), .ZN(\AES_ENC/us22/n1104 ) );
NOR2_X2 \AES_ENC/us22/U372  ( .A1(\AES_ENC/us22/n1102 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n1106 ) );
NOR2_X2 \AES_ENC/us22/U370  ( .A1(\AES_ENC/us22/n1103 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n1105 ) );
NOR4_X2 \AES_ENC/us22/U369  ( .A1(\AES_ENC/us22/n1107 ), .A2(\AES_ENC/us22/n1106 ), .A3(\AES_ENC/us22/n1105 ), .A4(\AES_ENC/us22/n1104 ), .ZN(\AES_ENC/us22/n1108 ) );
NOR3_X2 \AES_ENC/us22/U368  ( .A1(\AES_ENC/us22/n959 ), .A2(\AES_ENC/us22/n621 ), .A3(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n963 ) );
NOR2_X2 \AES_ENC/us22/U367  ( .A1(\AES_ENC/us22/n626 ), .A2(\AES_ENC/us22/n627 ), .ZN(\AES_ENC/us22/n1114 ) );
INV_X4 \AES_ENC/us22/U366  ( .A(\AES_ENC/us22/n1024 ), .ZN(\AES_ENC/us22/n606 ) );
NOR3_X2 \AES_ENC/us22/U365  ( .A1(\AES_ENC/us22/n910 ), .A2(\AES_ENC/us22/n1059 ), .A3(\AES_ENC/us22/n611 ), .ZN(\AES_ENC/us22/n1115 ) );
INV_X4 \AES_ENC/us22/U364  ( .A(\AES_ENC/us22/n1094 ), .ZN(\AES_ENC/us22/n613 ) );
NOR2_X2 \AES_ENC/us22/U363  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n931 ), .ZN(\AES_ENC/us22/n1100 ) );
INV_X4 \AES_ENC/us22/U354  ( .A(\AES_ENC/us22/n1093 ), .ZN(\AES_ENC/us22/n617 ) );
NOR2_X2 \AES_ENC/us22/U353  ( .A1(\AES_ENC/us22/n569 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n929 ) );
NOR2_X2 \AES_ENC/us22/U352  ( .A1(\AES_ENC/us22/n620 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n926 ) );
NOR2_X2 \AES_ENC/us22/U351  ( .A1(\AES_ENC/us22/n572 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n1095 ) );
NOR2_X2 \AES_ENC/us22/U350  ( .A1(\AES_ENC/us22/n609 ), .A2(\AES_ENC/us22/n627 ), .ZN(\AES_ENC/us22/n1010 ) );
NOR2_X2 \AES_ENC/us22/U349  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n1103 ) );
NOR2_X2 \AES_ENC/us22/U348  ( .A1(\AES_ENC/us22/n622 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n1059 ) );
NOR2_X2 \AES_ENC/us22/U347  ( .A1(\AES_ENC/sa22 [1]), .A2(\AES_ENC/us22/n1120 ), .ZN(\AES_ENC/us22/n1022 ) );
NOR2_X2 \AES_ENC/us22/U346  ( .A1(\AES_ENC/us22/n619 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n911 ) );
NOR2_X2 \AES_ENC/us22/U345  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/us22/n1025 ), .ZN(\AES_ENC/us22/n826 ) );
NOR2_X2 \AES_ENC/us22/U338  ( .A1(\AES_ENC/us22/n626 ), .A2(\AES_ENC/us22/n607 ), .ZN(\AES_ENC/us22/n1072 ) );
NOR2_X2 \AES_ENC/us22/U335  ( .A1(\AES_ENC/us22/n627 ), .A2(\AES_ENC/us22/n616 ), .ZN(\AES_ENC/us22/n956 ) );
NOR2_X2 \AES_ENC/us22/U329  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/us22/n624 ), .ZN(\AES_ENC/us22/n1121 ) );
NOR2_X2 \AES_ENC/us22/U328  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/us22/n624 ), .ZN(\AES_ENC/us22/n1058 ) );
NOR2_X2 \AES_ENC/us22/U327  ( .A1(\AES_ENC/us22/n625 ), .A2(\AES_ENC/us22/n611 ), .ZN(\AES_ENC/us22/n1073 ) );
NOR2_X2 \AES_ENC/us22/U325  ( .A1(\AES_ENC/sa22 [1]), .A2(\AES_ENC/us22/n1025 ), .ZN(\AES_ENC/us22/n1054 ) );
NOR2_X2 \AES_ENC/us22/U324  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/us22/n931 ), .ZN(\AES_ENC/us22/n1029 ) );
NOR2_X2 \AES_ENC/us22/U319  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n1056 ) );
NOR2_X2 \AES_ENC/us22/U318  ( .A1(\AES_ENC/us22/n614 ), .A2(\AES_ENC/us22/n626 ), .ZN(\AES_ENC/us22/n1050 ) );
NOR2_X2 \AES_ENC/us22/U317  ( .A1(\AES_ENC/us22/n1121 ), .A2(\AES_ENC/us22/n1025 ), .ZN(\AES_ENC/us22/n1120 ) );
NOR2_X2 \AES_ENC/us22/U316  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/us22/n572 ), .ZN(\AES_ENC/us22/n1074 ) );
NOR2_X2 \AES_ENC/us22/U315  ( .A1(\AES_ENC/us22/n1058 ), .A2(\AES_ENC/us22/n1054 ), .ZN(\AES_ENC/us22/n878 ) );
NOR2_X2 \AES_ENC/us22/U314  ( .A1(\AES_ENC/us22/n878 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n879 ) );
NOR2_X2 \AES_ENC/us22/U312  ( .A1(\AES_ENC/us22/n880 ), .A2(\AES_ENC/us22/n879 ), .ZN(\AES_ENC/us22/n887 ) );
NOR2_X2 \AES_ENC/us22/U311  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n588 ), .ZN(\AES_ENC/us22/n957 ) );
NOR2_X2 \AES_ENC/us22/U310  ( .A1(\AES_ENC/us22/n958 ), .A2(\AES_ENC/us22/n957 ), .ZN(\AES_ENC/us22/n965 ) );
NOR3_X2 \AES_ENC/us22/U309  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n1091 ), .A3(\AES_ENC/us22/n1022 ), .ZN(\AES_ENC/us22/n720 ) );
NOR3_X2 \AES_ENC/us22/U303  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n1054 ), .A3(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n719 ) );
NOR2_X2 \AES_ENC/us22/U302  ( .A1(\AES_ENC/us22/n720 ), .A2(\AES_ENC/us22/n719 ), .ZN(\AES_ENC/us22/n726 ) );
NOR2_X2 \AES_ENC/us22/U300  ( .A1(\AES_ENC/us22/n614 ), .A2(\AES_ENC/us22/n591 ), .ZN(\AES_ENC/us22/n865 ) );
NOR2_X2 \AES_ENC/us22/U299  ( .A1(\AES_ENC/us22/n1059 ), .A2(\AES_ENC/us22/n1058 ), .ZN(\AES_ENC/us22/n1060 ) );
NOR2_X2 \AES_ENC/us22/U298  ( .A1(\AES_ENC/us22/n1095 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n668 ) );
NOR2_X2 \AES_ENC/us22/U297  ( .A1(\AES_ENC/us22/n826 ), .A2(\AES_ENC/us22/n573 ), .ZN(\AES_ENC/us22/n750 ) );
NOR2_X2 \AES_ENC/us22/U296  ( .A1(\AES_ENC/us22/n750 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n751 ) );
NOR2_X2 \AES_ENC/us22/U295  ( .A1(\AES_ENC/us22/n907 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n908 ) );
NOR2_X2 \AES_ENC/us22/U294  ( .A1(\AES_ENC/us22/n990 ), .A2(\AES_ENC/us22/n926 ), .ZN(\AES_ENC/us22/n780 ) );
NOR2_X2 \AES_ENC/us22/U293  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n584 ), .ZN(\AES_ENC/us22/n838 ) );
NOR2_X2 \AES_ENC/us22/U292  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n602 ), .ZN(\AES_ENC/us22/n837 ) );
NOR2_X2 \AES_ENC/us22/U291  ( .A1(\AES_ENC/us22/n838 ), .A2(\AES_ENC/us22/n837 ), .ZN(\AES_ENC/us22/n845 ) );
NOR2_X2 \AES_ENC/us22/U290  ( .A1(\AES_ENC/us22/n1022 ), .A2(\AES_ENC/us22/n1058 ), .ZN(\AES_ENC/us22/n740 ) );
NOR2_X2 \AES_ENC/us22/U284  ( .A1(\AES_ENC/us22/n740 ), .A2(\AES_ENC/us22/n616 ), .ZN(\AES_ENC/us22/n742 ) );
NOR2_X2 \AES_ENC/us22/U283  ( .A1(\AES_ENC/us22/n1098 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n1099 ) );
NOR2_X2 \AES_ENC/us22/U282  ( .A1(\AES_ENC/us22/n1120 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n993 ) );
NOR2_X2 \AES_ENC/us22/U281  ( .A1(\AES_ENC/us22/n993 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n994 ) );
NOR2_X2 \AES_ENC/us22/U280  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n620 ), .ZN(\AES_ENC/us22/n1026 ) );
NOR2_X2 \AES_ENC/us22/U279  ( .A1(\AES_ENC/us22/n573 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n1027 ) );
NOR2_X2 \AES_ENC/us22/U273  ( .A1(\AES_ENC/us22/n1027 ), .A2(\AES_ENC/us22/n1026 ), .ZN(\AES_ENC/us22/n1028 ) );
NOR2_X2 \AES_ENC/us22/U272  ( .A1(\AES_ENC/us22/n1029 ), .A2(\AES_ENC/us22/n1028 ), .ZN(\AES_ENC/us22/n1034 ) );
NOR4_X2 \AES_ENC/us22/U271  ( .A1(\AES_ENC/us22/n757 ), .A2(\AES_ENC/us22/n756 ), .A3(\AES_ENC/us22/n755 ), .A4(\AES_ENC/us22/n754 ), .ZN(\AES_ENC/us22/n758 ) );
NOR2_X2 \AES_ENC/us22/U270  ( .A1(\AES_ENC/us22/n752 ), .A2(\AES_ENC/us22/n751 ), .ZN(\AES_ENC/us22/n759 ) );
NOR2_X2 \AES_ENC/us22/U269  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n1071 ), .ZN(\AES_ENC/us22/n669 ) );
NOR2_X2 \AES_ENC/us22/U268  ( .A1(\AES_ENC/us22/n1056 ), .A2(\AES_ENC/us22/n990 ), .ZN(\AES_ENC/us22/n991 ) );
NOR2_X2 \AES_ENC/us22/U267  ( .A1(\AES_ENC/us22/n991 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n995 ) );
NOR2_X2 \AES_ENC/us22/U263  ( .A1(\AES_ENC/us22/n607 ), .A2(\AES_ENC/us22/n590 ), .ZN(\AES_ENC/us22/n1008 ) );
NOR2_X2 \AES_ENC/us22/U262  ( .A1(\AES_ENC/us22/n839 ), .A2(\AES_ENC/us22/n582 ), .ZN(\AES_ENC/us22/n693 ) );
NOR2_X2 \AES_ENC/us22/U258  ( .A1(\AES_ENC/us22/n606 ), .A2(\AES_ENC/us22/n906 ), .ZN(\AES_ENC/us22/n741 ) );
NOR2_X2 \AES_ENC/us22/U255  ( .A1(\AES_ENC/us22/n1054 ), .A2(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n763 ) );
NOR2_X2 \AES_ENC/us22/U254  ( .A1(\AES_ENC/us22/n763 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n769 ) );
NOR2_X2 \AES_ENC/us22/U253  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n577 ), .ZN(\AES_ENC/us22/n1007 ) );
NOR2_X2 \AES_ENC/us22/U252  ( .A1(\AES_ENC/us22/n609 ), .A2(\AES_ENC/us22/n580 ), .ZN(\AES_ENC/us22/n1123 ) );
NOR2_X2 \AES_ENC/us22/U251  ( .A1(\AES_ENC/us22/n609 ), .A2(\AES_ENC/us22/n590 ), .ZN(\AES_ENC/us22/n710 ) );
INV_X4 \AES_ENC/us22/U250  ( .A(\AES_ENC/us22/n1029 ), .ZN(\AES_ENC/us22/n582 ) );
NOR2_X2 \AES_ENC/us22/U243  ( .A1(\AES_ENC/us22/n616 ), .A2(\AES_ENC/us22/n597 ), .ZN(\AES_ENC/us22/n883 ) );
NOR2_X2 \AES_ENC/us22/U242  ( .A1(\AES_ENC/us22/n593 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n1125 ) );
NOR2_X2 \AES_ENC/us22/U241  ( .A1(\AES_ENC/us22/n911 ), .A2(\AES_ENC/us22/n910 ), .ZN(\AES_ENC/us22/n912 ) );
NOR2_X2 \AES_ENC/us22/U240  ( .A1(\AES_ENC/us22/n912 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n916 ) );
NOR2_X2 \AES_ENC/us22/U239  ( .A1(\AES_ENC/us22/n990 ), .A2(\AES_ENC/us22/n929 ), .ZN(\AES_ENC/us22/n892 ) );
NOR2_X2 \AES_ENC/us22/U238  ( .A1(\AES_ENC/us22/n892 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n893 ) );
NOR2_X2 \AES_ENC/us22/U237  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n602 ), .ZN(\AES_ENC/us22/n950 ) );
NOR2_X2 \AES_ENC/us22/U236  ( .A1(\AES_ENC/us22/n1079 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n1082 ) );
NOR2_X2 \AES_ENC/us22/U235  ( .A1(\AES_ENC/us22/n910 ), .A2(\AES_ENC/us22/n1056 ), .ZN(\AES_ENC/us22/n941 ) );
NOR2_X2 \AES_ENC/us22/U234  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n1077 ), .ZN(\AES_ENC/us22/n841 ) );
NOR2_X2 \AES_ENC/us22/U229  ( .A1(\AES_ENC/us22/n623 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n630 ) );
NOR2_X2 \AES_ENC/us22/U228  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n602 ), .ZN(\AES_ENC/us22/n806 ) );
NOR2_X2 \AES_ENC/us22/U227  ( .A1(\AES_ENC/us22/n623 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n948 ) );
NOR2_X2 \AES_ENC/us22/U226  ( .A1(\AES_ENC/us22/n606 ), .A2(\AES_ENC/us22/n589 ), .ZN(\AES_ENC/us22/n997 ) );
NOR2_X2 \AES_ENC/us22/U225  ( .A1(\AES_ENC/us22/n1121 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n1122 ) );
NOR2_X2 \AES_ENC/us22/U223  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n1023 ), .ZN(\AES_ENC/us22/n756 ) );
NOR2_X2 \AES_ENC/us22/U222  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n602 ), .ZN(\AES_ENC/us22/n870 ) );
NOR2_X2 \AES_ENC/us22/U221  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n569 ), .ZN(\AES_ENC/us22/n947 ) );
NOR2_X2 \AES_ENC/us22/U217  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n1077 ), .ZN(\AES_ENC/us22/n1084 ) );
NOR2_X2 \AES_ENC/us22/U213  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n855 ), .ZN(\AES_ENC/us22/n709 ) );
NOR2_X2 \AES_ENC/us22/U212  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n589 ), .ZN(\AES_ENC/us22/n868 ) );
NOR2_X2 \AES_ENC/us22/U211  ( .A1(\AES_ENC/us22/n1120 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n1124 ) );
NOR2_X2 \AES_ENC/us22/U210  ( .A1(\AES_ENC/us22/n1120 ), .A2(\AES_ENC/us22/n839 ), .ZN(\AES_ENC/us22/n842 ) );
NOR2_X2 \AES_ENC/us22/U209  ( .A1(\AES_ENC/us22/n1120 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n696 ) );
NOR2_X2 \AES_ENC/us22/U208  ( .A1(\AES_ENC/us22/n1074 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n1076 ) );
NOR2_X2 \AES_ENC/us22/U207  ( .A1(\AES_ENC/us22/n1074 ), .A2(\AES_ENC/us22/n620 ), .ZN(\AES_ENC/us22/n781 ) );
NOR3_X2 \AES_ENC/us22/U201  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n1056 ), .A3(\AES_ENC/us22/n990 ), .ZN(\AES_ENC/us22/n979 ) );
NOR3_X2 \AES_ENC/us22/U200  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n1058 ), .A3(\AES_ENC/us22/n1059 ), .ZN(\AES_ENC/us22/n854 ) );
NOR2_X2 \AES_ENC/us22/U199  ( .A1(\AES_ENC/us22/n996 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n869 ) );
NOR2_X2 \AES_ENC/us22/U198  ( .A1(\AES_ENC/us22/n1056 ), .A2(\AES_ENC/us22/n1074 ), .ZN(\AES_ENC/us22/n1057 ) );
NOR3_X2 \AES_ENC/us22/U197  ( .A1(\AES_ENC/us22/n607 ), .A2(\AES_ENC/us22/n1120 ), .A3(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n978 ) );
NOR2_X2 \AES_ENC/us22/U196  ( .A1(\AES_ENC/us22/n996 ), .A2(\AES_ENC/us22/n911 ), .ZN(\AES_ENC/us22/n1116 ) );
NOR2_X2 \AES_ENC/us22/U195  ( .A1(\AES_ENC/us22/n1074 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n754 ) );
NOR2_X2 \AES_ENC/us22/U194  ( .A1(\AES_ENC/us22/n926 ), .A2(\AES_ENC/us22/n1103 ), .ZN(\AES_ENC/us22/n977 ) );
NOR2_X2 \AES_ENC/us22/U187  ( .A1(\AES_ENC/us22/n839 ), .A2(\AES_ENC/us22/n824 ), .ZN(\AES_ENC/us22/n1092 ) );
NOR2_X2 \AES_ENC/us22/U186  ( .A1(\AES_ENC/us22/n573 ), .A2(\AES_ENC/us22/n1074 ), .ZN(\AES_ENC/us22/n684 ) );
NOR2_X2 \AES_ENC/us22/U185  ( .A1(\AES_ENC/us22/n826 ), .A2(\AES_ENC/us22/n1059 ), .ZN(\AES_ENC/us22/n907 ) );
NOR3_X2 \AES_ENC/us22/U184  ( .A1(\AES_ENC/us22/n625 ), .A2(\AES_ENC/us22/n1115 ), .A3(\AES_ENC/us22/n585 ), .ZN(\AES_ENC/us22/n831 ) );
NOR3_X2 \AES_ENC/us22/U183  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n1056 ), .A3(\AES_ENC/us22/n990 ), .ZN(\AES_ENC/us22/n896 ) );
NOR3_X2 \AES_ENC/us22/U182  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n573 ), .A3(\AES_ENC/us22/n1013 ), .ZN(\AES_ENC/us22/n670 ) );
NOR3_X2 \AES_ENC/us22/U181  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n1091 ), .A3(\AES_ENC/us22/n1022 ), .ZN(\AES_ENC/us22/n843 ) );
NOR2_X2 \AES_ENC/us22/U180  ( .A1(\AES_ENC/us22/n1029 ), .A2(\AES_ENC/us22/n1095 ), .ZN(\AES_ENC/us22/n735 ) );
NOR2_X2 \AES_ENC/us22/U174  ( .A1(\AES_ENC/us22/n1100 ), .A2(\AES_ENC/us22/n854 ), .ZN(\AES_ENC/us22/n860 ) );
NAND3_X2 \AES_ENC/us22/U173  ( .A1(\AES_ENC/us22/n569 ), .A2(\AES_ENC/us22/n582 ), .A3(\AES_ENC/us22/n681 ), .ZN(\AES_ENC/us22/n691 ) );
NOR2_X2 \AES_ENC/us22/U172  ( .A1(\AES_ENC/us22/n683 ), .A2(\AES_ENC/us22/n682 ), .ZN(\AES_ENC/us22/n690 ) );
NOR3_X2 \AES_ENC/us22/U171  ( .A1(\AES_ENC/us22/n695 ), .A2(\AES_ENC/us22/n694 ), .A3(\AES_ENC/us22/n693 ), .ZN(\AES_ENC/us22/n700 ) );
NOR4_X2 \AES_ENC/us22/U170  ( .A1(\AES_ENC/us22/n983 ), .A2(\AES_ENC/us22/n698 ), .A3(\AES_ENC/us22/n697 ), .A4(\AES_ENC/us22/n696 ), .ZN(\AES_ENC/us22/n699 ) );
NOR4_X2 \AES_ENC/us22/U169  ( .A1(\AES_ENC/us22/n896 ), .A2(\AES_ENC/us22/n895 ), .A3(\AES_ENC/us22/n894 ), .A4(\AES_ENC/us22/n893 ), .ZN(\AES_ENC/us22/n897 ) );
NOR2_X2 \AES_ENC/us22/U168  ( .A1(\AES_ENC/us22/n866 ), .A2(\AES_ENC/us22/n865 ), .ZN(\AES_ENC/us22/n872 ) );
NOR4_X2 \AES_ENC/us22/U162  ( .A1(\AES_ENC/us22/n870 ), .A2(\AES_ENC/us22/n869 ), .A3(\AES_ENC/us22/n868 ), .A4(\AES_ENC/us22/n867 ), .ZN(\AES_ENC/us22/n871 ) );
NOR2_X2 \AES_ENC/us22/U161  ( .A1(\AES_ENC/us22/n946 ), .A2(\AES_ENC/us22/n945 ), .ZN(\AES_ENC/us22/n952 ) );
NOR4_X2 \AES_ENC/us22/U160  ( .A1(\AES_ENC/us22/n950 ), .A2(\AES_ENC/us22/n949 ), .A3(\AES_ENC/us22/n948 ), .A4(\AES_ENC/us22/n947 ), .ZN(\AES_ENC/us22/n951 ) );
NOR4_X2 \AES_ENC/us22/U159  ( .A1(\AES_ENC/us22/n983 ), .A2(\AES_ENC/us22/n982 ), .A3(\AES_ENC/us22/n981 ), .A4(\AES_ENC/us22/n980 ), .ZN(\AES_ENC/us22/n984 ) );
NOR2_X2 \AES_ENC/us22/U158  ( .A1(\AES_ENC/us22/n979 ), .A2(\AES_ENC/us22/n978 ), .ZN(\AES_ENC/us22/n985 ) );
NOR4_X2 \AES_ENC/us22/U157  ( .A1(\AES_ENC/us22/n1125 ), .A2(\AES_ENC/us22/n1124 ), .A3(\AES_ENC/us22/n1123 ), .A4(\AES_ENC/us22/n1122 ), .ZN(\AES_ENC/us22/n1126 ) );
NOR4_X2 \AES_ENC/us22/U156  ( .A1(\AES_ENC/us22/n1084 ), .A2(\AES_ENC/us22/n1083 ), .A3(\AES_ENC/us22/n1082 ), .A4(\AES_ENC/us22/n1081 ), .ZN(\AES_ENC/us22/n1085 ) );
NOR2_X2 \AES_ENC/us22/U155  ( .A1(\AES_ENC/us22/n1076 ), .A2(\AES_ENC/us22/n1075 ), .ZN(\AES_ENC/us22/n1086 ) );
NOR3_X2 \AES_ENC/us22/U154  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n1054 ), .A3(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n961 ) );
NOR3_X2 \AES_ENC/us22/U153  ( .A1(\AES_ENC/us22/n620 ), .A2(\AES_ENC/us22/n1074 ), .A3(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n671 ) );
NOR2_X2 \AES_ENC/us22/U152  ( .A1(\AES_ENC/us22/n1057 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n1062 ) );
NOR2_X2 \AES_ENC/us22/U143  ( .A1(\AES_ENC/us22/n1055 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n1063 ) );
NOR2_X2 \AES_ENC/us22/U142  ( .A1(\AES_ENC/us22/n1060 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n1061 ) );
NOR4_X2 \AES_ENC/us22/U141  ( .A1(\AES_ENC/us22/n1064 ), .A2(\AES_ENC/us22/n1063 ), .A3(\AES_ENC/us22/n1062 ), .A4(\AES_ENC/us22/n1061 ), .ZN(\AES_ENC/us22/n1065 ) );
NOR3_X2 \AES_ENC/us22/U140  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n1120 ), .A3(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n918 ) );
NOR3_X2 \AES_ENC/us22/U132  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n573 ), .A3(\AES_ENC/us22/n1013 ), .ZN(\AES_ENC/us22/n917 ) );
NOR2_X2 \AES_ENC/us22/U131  ( .A1(\AES_ENC/us22/n914 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n915 ) );
NOR4_X2 \AES_ENC/us22/U130  ( .A1(\AES_ENC/us22/n918 ), .A2(\AES_ENC/us22/n917 ), .A3(\AES_ENC/us22/n916 ), .A4(\AES_ENC/us22/n915 ), .ZN(\AES_ENC/us22/n919 ) );
NOR2_X2 \AES_ENC/us22/U129  ( .A1(\AES_ENC/us22/n616 ), .A2(\AES_ENC/us22/n580 ), .ZN(\AES_ENC/us22/n771 ) );
NOR2_X2 \AES_ENC/us22/U128  ( .A1(\AES_ENC/us22/n1103 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n772 ) );
NOR2_X2 \AES_ENC/us22/U127  ( .A1(\AES_ENC/us22/n610 ), .A2(\AES_ENC/us22/n599 ), .ZN(\AES_ENC/us22/n773 ) );
NOR4_X2 \AES_ENC/us22/U126  ( .A1(\AES_ENC/us22/n773 ), .A2(\AES_ENC/us22/n772 ), .A3(\AES_ENC/us22/n771 ), .A4(\AES_ENC/us22/n770 ), .ZN(\AES_ENC/us22/n774 ) );
NOR2_X2 \AES_ENC/us22/U121  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n595 ), .ZN(\AES_ENC/us22/n858 ) );
NOR2_X2 \AES_ENC/us22/U120  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n855 ), .ZN(\AES_ENC/us22/n857 ) );
NOR2_X2 \AES_ENC/us22/U119  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n587 ), .ZN(\AES_ENC/us22/n856 ) );
NOR4_X2 \AES_ENC/us22/U118  ( .A1(\AES_ENC/us22/n858 ), .A2(\AES_ENC/us22/n857 ), .A3(\AES_ENC/us22/n856 ), .A4(\AES_ENC/us22/n958 ), .ZN(\AES_ENC/us22/n859 ) );
NOR2_X2 \AES_ENC/us22/U117  ( .A1(\AES_ENC/us22/n735 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n687 ) );
NOR2_X2 \AES_ENC/us22/U116  ( .A1(\AES_ENC/us22/n684 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n688 ) );
NOR2_X2 \AES_ENC/us22/U115  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n600 ), .ZN(\AES_ENC/us22/n686 ) );
NOR4_X2 \AES_ENC/us22/U106  ( .A1(\AES_ENC/us22/n688 ), .A2(\AES_ENC/us22/n687 ), .A3(\AES_ENC/us22/n686 ), .A4(\AES_ENC/us22/n685 ), .ZN(\AES_ENC/us22/n689 ) );
NOR2_X2 \AES_ENC/us22/U105  ( .A1(\AES_ENC/us22/n780 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n784 ) );
NOR2_X2 \AES_ENC/us22/U104  ( .A1(\AES_ENC/us22/n1117 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n782 ) );
NOR2_X2 \AES_ENC/us22/U103  ( .A1(\AES_ENC/us22/n781 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n783 ) );
NOR4_X2 \AES_ENC/us22/U102  ( .A1(\AES_ENC/us22/n880 ), .A2(\AES_ENC/us22/n784 ), .A3(\AES_ENC/us22/n783 ), .A4(\AES_ENC/us22/n782 ), .ZN(\AES_ENC/us22/n785 ) );
NOR2_X2 \AES_ENC/us22/U101  ( .A1(\AES_ENC/us22/n583 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n814 ) );
NOR2_X2 \AES_ENC/us22/U100  ( .A1(\AES_ENC/us22/n907 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n813 ) );
NOR3_X2 \AES_ENC/us22/U95  ( .A1(\AES_ENC/us22/n606 ), .A2(\AES_ENC/us22/n1058 ), .A3(\AES_ENC/us22/n1059 ), .ZN(\AES_ENC/us22/n815 ) );
NOR4_X2 \AES_ENC/us22/U94  ( .A1(\AES_ENC/us22/n815 ), .A2(\AES_ENC/us22/n814 ), .A3(\AES_ENC/us22/n813 ), .A4(\AES_ENC/us22/n812 ), .ZN(\AES_ENC/us22/n816 ) );
NOR2_X2 \AES_ENC/us22/U93  ( .A1(\AES_ENC/us22/n617 ), .A2(\AES_ENC/us22/n569 ), .ZN(\AES_ENC/us22/n721 ) );
NOR2_X2 \AES_ENC/us22/U92  ( .A1(\AES_ENC/us22/n1031 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n723 ) );
NOR2_X2 \AES_ENC/us22/U91  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n1096 ), .ZN(\AES_ENC/us22/n722 ) );
NOR4_X2 \AES_ENC/us22/U90  ( .A1(\AES_ENC/us22/n724 ), .A2(\AES_ENC/us22/n723 ), .A3(\AES_ENC/us22/n722 ), .A4(\AES_ENC/us22/n721 ), .ZN(\AES_ENC/us22/n725 ) );
NOR2_X2 \AES_ENC/us22/U89  ( .A1(\AES_ENC/us22/n911 ), .A2(\AES_ENC/us22/n990 ), .ZN(\AES_ENC/us22/n1009 ) );
NOR2_X2 \AES_ENC/us22/U88  ( .A1(\AES_ENC/us22/n1013 ), .A2(\AES_ENC/us22/n573 ), .ZN(\AES_ENC/us22/n1014 ) );
NOR2_X2 \AES_ENC/us22/U87  ( .A1(\AES_ENC/us22/n1014 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n1015 ) );
NOR4_X2 \AES_ENC/us22/U86  ( .A1(\AES_ENC/us22/n1016 ), .A2(\AES_ENC/us22/n1015 ), .A3(\AES_ENC/us22/n1119 ), .A4(\AES_ENC/us22/n1046 ), .ZN(\AES_ENC/us22/n1017 ) );
NOR2_X2 \AES_ENC/us22/U81  ( .A1(\AES_ENC/us22/n996 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n998 ) );
NOR2_X2 \AES_ENC/us22/U80  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n577 ), .ZN(\AES_ENC/us22/n1000 ) );
NOR2_X2 \AES_ENC/us22/U79  ( .A1(\AES_ENC/us22/n616 ), .A2(\AES_ENC/us22/n1096 ), .ZN(\AES_ENC/us22/n999 ) );
NOR4_X2 \AES_ENC/us22/U78  ( .A1(\AES_ENC/us22/n1000 ), .A2(\AES_ENC/us22/n999 ), .A3(\AES_ENC/us22/n998 ), .A4(\AES_ENC/us22/n997 ), .ZN(\AES_ENC/us22/n1001 ) );
NOR2_X2 \AES_ENC/us22/U74  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n1096 ), .ZN(\AES_ENC/us22/n697 ) );
NOR2_X2 \AES_ENC/us22/U73  ( .A1(\AES_ENC/us22/n620 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n958 ) );
NOR2_X2 \AES_ENC/us22/U72  ( .A1(\AES_ENC/us22/n911 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n983 ) );
NOR2_X2 \AES_ENC/us22/U71  ( .A1(\AES_ENC/us22/n1054 ), .A2(\AES_ENC/us22/n1103 ), .ZN(\AES_ENC/us22/n1031 ) );
INV_X4 \AES_ENC/us22/U65  ( .A(\AES_ENC/us22/n1050 ), .ZN(\AES_ENC/us22/n612 ) );
INV_X4 \AES_ENC/us22/U64  ( .A(\AES_ENC/us22/n1072 ), .ZN(\AES_ENC/us22/n605 ) );
INV_X4 \AES_ENC/us22/U63  ( .A(\AES_ENC/us22/n1073 ), .ZN(\AES_ENC/us22/n604 ) );
NOR2_X2 \AES_ENC/us22/U62  ( .A1(\AES_ENC/us22/n582 ), .A2(\AES_ENC/us22/n613 ), .ZN(\AES_ENC/us22/n880 ) );
NOR3_X2 \AES_ENC/us22/U61  ( .A1(\AES_ENC/us22/n826 ), .A2(\AES_ENC/us22/n1121 ), .A3(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n946 ) );
INV_X4 \AES_ENC/us22/U59  ( .A(\AES_ENC/us22/n1010 ), .ZN(\AES_ENC/us22/n608 ) );
NOR3_X2 \AES_ENC/us22/U58  ( .A1(\AES_ENC/us22/n573 ), .A2(\AES_ENC/us22/n1029 ), .A3(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n1119 ) );
INV_X4 \AES_ENC/us22/U57  ( .A(\AES_ENC/us22/n956 ), .ZN(\AES_ENC/us22/n615 ) );
NOR2_X2 \AES_ENC/us22/U50  ( .A1(\AES_ENC/us22/n623 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n1013 ) );
NOR2_X2 \AES_ENC/us22/U49  ( .A1(\AES_ENC/us22/n620 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n910 ) );
NOR2_X2 \AES_ENC/us22/U48  ( .A1(\AES_ENC/us22/n569 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n1091 ) );
NOR2_X2 \AES_ENC/us22/U47  ( .A1(\AES_ENC/us22/n622 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n990 ) );
NOR2_X2 \AES_ENC/us22/U46  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/us22/n1121 ), .ZN(\AES_ENC/us22/n996 ) );
NOR2_X2 \AES_ENC/us22/U45  ( .A1(\AES_ENC/us22/n610 ), .A2(\AES_ENC/us22/n600 ), .ZN(\AES_ENC/us22/n628 ) );
NOR2_X2 \AES_ENC/us22/U44  ( .A1(\AES_ENC/us22/n576 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n866 ) );
NOR2_X2 \AES_ENC/us22/U43  ( .A1(\AES_ENC/us22/n603 ), .A2(\AES_ENC/us22/n610 ), .ZN(\AES_ENC/us22/n1006 ) );
NOR2_X2 \AES_ENC/us22/U42  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n1117 ), .ZN(\AES_ENC/us22/n1118 ) );
NOR2_X2 \AES_ENC/us22/U41  ( .A1(\AES_ENC/us22/n1119 ), .A2(\AES_ENC/us22/n1118 ), .ZN(\AES_ENC/us22/n1127 ) );
NOR2_X2 \AES_ENC/us22/U36  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n594 ), .ZN(\AES_ENC/us22/n629 ) );
NOR2_X2 \AES_ENC/us22/U35  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n906 ), .ZN(\AES_ENC/us22/n909 ) );
NOR2_X2 \AES_ENC/us22/U34  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n597 ), .ZN(\AES_ENC/us22/n658 ) );
NOR2_X2 \AES_ENC/us22/U33  ( .A1(\AES_ENC/us22/n1116 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n695 ) );
NOR2_X2 \AES_ENC/us22/U32  ( .A1(\AES_ENC/us22/n1078 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n1083 ) );
NOR2_X2 \AES_ENC/us22/U31  ( .A1(\AES_ENC/us22/n941 ), .A2(\AES_ENC/us22/n608 ), .ZN(\AES_ENC/us22/n724 ) );
NOR2_X2 \AES_ENC/us22/U30  ( .A1(\AES_ENC/us22/n598 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n1107 ) );
NOR2_X2 \AES_ENC/us22/U29  ( .A1(\AES_ENC/us22/n576 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n840 ) );
NOR2_X2 \AES_ENC/us22/U24  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n593 ), .ZN(\AES_ENC/us22/n633 ) );
NOR2_X2 \AES_ENC/us22/U23  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n1080 ), .ZN(\AES_ENC/us22/n1081 ) );
NOR2_X2 \AES_ENC/us22/U21  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n1045 ), .ZN(\AES_ENC/us22/n812 ) );
NOR2_X2 \AES_ENC/us22/U20  ( .A1(\AES_ENC/us22/n1009 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n960 ) );
NOR2_X2 \AES_ENC/us22/U19  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n601 ), .ZN(\AES_ENC/us22/n982 ) );
NOR2_X2 \AES_ENC/us22/U18  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n594 ), .ZN(\AES_ENC/us22/n757 ) );
NOR2_X2 \AES_ENC/us22/U17  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n590 ), .ZN(\AES_ENC/us22/n698 ) );
NOR2_X2 \AES_ENC/us22/U16  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n619 ), .ZN(\AES_ENC/us22/n708 ) );
NOR2_X2 \AES_ENC/us22/U15  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n582 ), .ZN(\AES_ENC/us22/n770 ) );
NOR2_X2 \AES_ENC/us22/U10  ( .A1(\AES_ENC/us22/n619 ), .A2(\AES_ENC/us22/n604 ), .ZN(\AES_ENC/us22/n803 ) );
NOR2_X2 \AES_ENC/us22/U9  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n881 ), .ZN(\AES_ENC/us22/n711 ) );
NOR2_X2 \AES_ENC/us22/U8  ( .A1(\AES_ENC/us22/n615 ), .A2(\AES_ENC/us22/n582 ), .ZN(\AES_ENC/us22/n867 ) );
NOR2_X2 \AES_ENC/us22/U7  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n599 ), .ZN(\AES_ENC/us22/n804 ) );
NOR2_X2 \AES_ENC/us22/U6  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n620 ), .ZN(\AES_ENC/us22/n1046 ) );
OR2_X4 \AES_ENC/us22/U5  ( .A1(\AES_ENC/us22/n624 ), .A2(\AES_ENC/sa22 [1]),.ZN(\AES_ENC/us22/n570 ) );
OR2_X4 \AES_ENC/us22/U4  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/sa22 [4]),.ZN(\AES_ENC/us22/n569 ) );
NAND2_X2 \AES_ENC/us22/U514  ( .A1(\AES_ENC/us22/n1121 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n1030 ) );
AND2_X2 \AES_ENC/us22/U513  ( .A1(\AES_ENC/us22/n597 ), .A2(\AES_ENC/us22/n1030 ), .ZN(\AES_ENC/us22/n1049 ) );
NAND2_X2 \AES_ENC/us22/U511  ( .A1(\AES_ENC/us22/n1049 ), .A2(\AES_ENC/us22/n794 ), .ZN(\AES_ENC/us22/n637 ) );
AND2_X2 \AES_ENC/us22/U493  ( .A1(\AES_ENC/us22/n779 ), .A2(\AES_ENC/us22/n996 ), .ZN(\AES_ENC/us22/n632 ) );
NAND4_X2 \AES_ENC/us22/U485  ( .A1(\AES_ENC/us22/n637 ), .A2(\AES_ENC/us22/n636 ), .A3(\AES_ENC/us22/n635 ), .A4(\AES_ENC/us22/n634 ), .ZN(\AES_ENC/us22/n638 ) );
NAND2_X2 \AES_ENC/us22/U484  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n638 ), .ZN(\AES_ENC/us22/n679 ) );
NAND2_X2 \AES_ENC/us22/U481  ( .A1(\AES_ENC/us22/n1094 ), .A2(\AES_ENC/us22/n591 ), .ZN(\AES_ENC/us22/n648 ) );
NAND2_X2 \AES_ENC/us22/U476  ( .A1(\AES_ENC/us22/n601 ), .A2(\AES_ENC/us22/n590 ), .ZN(\AES_ENC/us22/n762 ) );
NAND2_X2 \AES_ENC/us22/U475  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n762 ), .ZN(\AES_ENC/us22/n647 ) );
NAND4_X2 \AES_ENC/us22/U457  ( .A1(\AES_ENC/us22/n648 ), .A2(\AES_ENC/us22/n647 ), .A3(\AES_ENC/us22/n646 ), .A4(\AES_ENC/us22/n645 ), .ZN(\AES_ENC/us22/n649 ) );
NAND2_X2 \AES_ENC/us22/U456  ( .A1(\AES_ENC/sa22 [0]), .A2(\AES_ENC/us22/n649 ), .ZN(\AES_ENC/us22/n665 ) );
NAND2_X2 \AES_ENC/us22/U454  ( .A1(\AES_ENC/us22/n596 ), .A2(\AES_ENC/us22/n623 ), .ZN(\AES_ENC/us22/n855 ) );
NAND2_X2 \AES_ENC/us22/U453  ( .A1(\AES_ENC/us22/n587 ), .A2(\AES_ENC/us22/n855 ), .ZN(\AES_ENC/us22/n821 ) );
NAND2_X2 \AES_ENC/us22/U452  ( .A1(\AES_ENC/us22/n1093 ), .A2(\AES_ENC/us22/n821 ), .ZN(\AES_ENC/us22/n662 ) );
NAND2_X2 \AES_ENC/us22/U451  ( .A1(\AES_ENC/us22/n619 ), .A2(\AES_ENC/us22/n589 ), .ZN(\AES_ENC/us22/n650 ) );
NAND2_X2 \AES_ENC/us22/U450  ( .A1(\AES_ENC/us22/n956 ), .A2(\AES_ENC/us22/n650 ), .ZN(\AES_ENC/us22/n661 ) );
NAND2_X2 \AES_ENC/us22/U449  ( .A1(\AES_ENC/us22/n626 ), .A2(\AES_ENC/us22/n627 ), .ZN(\AES_ENC/us22/n839 ) );
OR2_X2 \AES_ENC/us22/U446  ( .A1(\AES_ENC/us22/n839 ), .A2(\AES_ENC/us22/n932 ), .ZN(\AES_ENC/us22/n656 ) );
NAND2_X2 \AES_ENC/us22/U445  ( .A1(\AES_ENC/us22/n621 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n1096 ) );
NAND2_X2 \AES_ENC/us22/U444  ( .A1(\AES_ENC/us22/n1030 ), .A2(\AES_ENC/us22/n1096 ), .ZN(\AES_ENC/us22/n651 ) );
NAND2_X2 \AES_ENC/us22/U443  ( .A1(\AES_ENC/us22/n1114 ), .A2(\AES_ENC/us22/n651 ), .ZN(\AES_ENC/us22/n655 ) );
OR3_X2 \AES_ENC/us22/U440  ( .A1(\AES_ENC/us22/n1079 ), .A2(\AES_ENC/sa22 [7]), .A3(\AES_ENC/us22/n626 ), .ZN(\AES_ENC/us22/n654 ));
NAND2_X2 \AES_ENC/us22/U439  ( .A1(\AES_ENC/us22/n593 ), .A2(\AES_ENC/us22/n601 ), .ZN(\AES_ENC/us22/n652 ) );
NAND4_X2 \AES_ENC/us22/U437  ( .A1(\AES_ENC/us22/n656 ), .A2(\AES_ENC/us22/n655 ), .A3(\AES_ENC/us22/n654 ), .A4(\AES_ENC/us22/n653 ), .ZN(\AES_ENC/us22/n657 ) );
NAND2_X2 \AES_ENC/us22/U436  ( .A1(\AES_ENC/sa22 [2]), .A2(\AES_ENC/us22/n657 ), .ZN(\AES_ENC/us22/n660 ) );
NAND4_X2 \AES_ENC/us22/U432  ( .A1(\AES_ENC/us22/n662 ), .A2(\AES_ENC/us22/n661 ), .A3(\AES_ENC/us22/n660 ), .A4(\AES_ENC/us22/n659 ), .ZN(\AES_ENC/us22/n663 ) );
NAND2_X2 \AES_ENC/us22/U431  ( .A1(\AES_ENC/us22/n663 ), .A2(\AES_ENC/us22/n574 ), .ZN(\AES_ENC/us22/n664 ) );
NAND2_X2 \AES_ENC/us22/U430  ( .A1(\AES_ENC/us22/n665 ), .A2(\AES_ENC/us22/n664 ), .ZN(\AES_ENC/us22/n666 ) );
NAND2_X2 \AES_ENC/us22/U429  ( .A1(\AES_ENC/sa22 [6]), .A2(\AES_ENC/us22/n666 ), .ZN(\AES_ENC/us22/n678 ) );
NAND2_X2 \AES_ENC/us22/U426  ( .A1(\AES_ENC/us22/n735 ), .A2(\AES_ENC/us22/n1093 ), .ZN(\AES_ENC/us22/n675 ) );
NAND2_X2 \AES_ENC/us22/U425  ( .A1(\AES_ENC/us22/n588 ), .A2(\AES_ENC/us22/n597 ), .ZN(\AES_ENC/us22/n1045 ) );
OR2_X2 \AES_ENC/us22/U424  ( .A1(\AES_ENC/us22/n1045 ), .A2(\AES_ENC/us22/n605 ), .ZN(\AES_ENC/us22/n674 ) );
NAND2_X2 \AES_ENC/us22/U423  ( .A1(\AES_ENC/sa22 [1]), .A2(\AES_ENC/us22/n620 ), .ZN(\AES_ENC/us22/n667 ) );
NAND2_X2 \AES_ENC/us22/U422  ( .A1(\AES_ENC/us22/n619 ), .A2(\AES_ENC/us22/n667 ), .ZN(\AES_ENC/us22/n1071 ) );
NAND4_X2 \AES_ENC/us22/U412  ( .A1(\AES_ENC/us22/n675 ), .A2(\AES_ENC/us22/n674 ), .A3(\AES_ENC/us22/n673 ), .A4(\AES_ENC/us22/n672 ), .ZN(\AES_ENC/us22/n676 ) );
NAND2_X2 \AES_ENC/us22/U411  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n676 ), .ZN(\AES_ENC/us22/n677 ) );
NAND2_X2 \AES_ENC/us22/U408  ( .A1(\AES_ENC/us22/n800 ), .A2(\AES_ENC/us22/n1022 ), .ZN(\AES_ENC/us22/n680 ) );
NAND2_X2 \AES_ENC/us22/U407  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n680 ), .ZN(\AES_ENC/us22/n681 ) );
AND2_X2 \AES_ENC/us22/U402  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n684 ), .ZN(\AES_ENC/us22/n682 ) );
NAND4_X2 \AES_ENC/us22/U395  ( .A1(\AES_ENC/us22/n691 ), .A2(\AES_ENC/us22/n581 ), .A3(\AES_ENC/us22/n690 ), .A4(\AES_ENC/us22/n689 ), .ZN(\AES_ENC/us22/n692 ) );
NAND2_X2 \AES_ENC/us22/U394  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n692 ), .ZN(\AES_ENC/us22/n733 ) );
NAND2_X2 \AES_ENC/us22/U392  ( .A1(\AES_ENC/us22/n977 ), .A2(\AES_ENC/us22/n1050 ), .ZN(\AES_ENC/us22/n702 ) );
NAND2_X2 \AES_ENC/us22/U391  ( .A1(\AES_ENC/us22/n1093 ), .A2(\AES_ENC/us22/n1045 ), .ZN(\AES_ENC/us22/n701 ) );
NAND4_X2 \AES_ENC/us22/U381  ( .A1(\AES_ENC/us22/n702 ), .A2(\AES_ENC/us22/n701 ), .A3(\AES_ENC/us22/n700 ), .A4(\AES_ENC/us22/n699 ), .ZN(\AES_ENC/us22/n703 ) );
NAND2_X2 \AES_ENC/us22/U380  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n703 ), .ZN(\AES_ENC/us22/n732 ) );
AND2_X2 \AES_ENC/us22/U379  ( .A1(\AES_ENC/sa22 [0]), .A2(\AES_ENC/sa22 [6]),.ZN(\AES_ENC/us22/n1113 ) );
NAND2_X2 \AES_ENC/us22/U378  ( .A1(\AES_ENC/us22/n601 ), .A2(\AES_ENC/us22/n1030 ), .ZN(\AES_ENC/us22/n881 ) );
NAND2_X2 \AES_ENC/us22/U377  ( .A1(\AES_ENC/us22/n1093 ), .A2(\AES_ENC/us22/n881 ), .ZN(\AES_ENC/us22/n715 ) );
NAND2_X2 \AES_ENC/us22/U376  ( .A1(\AES_ENC/us22/n1010 ), .A2(\AES_ENC/us22/n600 ), .ZN(\AES_ENC/us22/n714 ) );
NAND2_X2 \AES_ENC/us22/U375  ( .A1(\AES_ENC/us22/n855 ), .A2(\AES_ENC/us22/n588 ), .ZN(\AES_ENC/us22/n1117 ) );
XNOR2_X2 \AES_ENC/us22/U371  ( .A(\AES_ENC/us22/n611 ), .B(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n824 ) );
NAND4_X2 \AES_ENC/us22/U362  ( .A1(\AES_ENC/us22/n715 ), .A2(\AES_ENC/us22/n714 ), .A3(\AES_ENC/us22/n713 ), .A4(\AES_ENC/us22/n712 ), .ZN(\AES_ENC/us22/n716 ) );
NAND2_X2 \AES_ENC/us22/U361  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n716 ), .ZN(\AES_ENC/us22/n731 ) );
AND2_X2 \AES_ENC/us22/U360  ( .A1(\AES_ENC/sa22 [6]), .A2(\AES_ENC/us22/n574 ), .ZN(\AES_ENC/us22/n1131 ) );
NAND2_X2 \AES_ENC/us22/U359  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n717 ) );
NAND2_X2 \AES_ENC/us22/U358  ( .A1(\AES_ENC/us22/n1029 ), .A2(\AES_ENC/us22/n717 ), .ZN(\AES_ENC/us22/n728 ) );
NAND2_X2 \AES_ENC/us22/U357  ( .A1(\AES_ENC/sa22 [1]), .A2(\AES_ENC/us22/n624 ), .ZN(\AES_ENC/us22/n1097 ) );
NAND2_X2 \AES_ENC/us22/U356  ( .A1(\AES_ENC/us22/n603 ), .A2(\AES_ENC/us22/n1097 ), .ZN(\AES_ENC/us22/n718 ) );
NAND2_X2 \AES_ENC/us22/U355  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n718 ), .ZN(\AES_ENC/us22/n727 ) );
NAND4_X2 \AES_ENC/us22/U344  ( .A1(\AES_ENC/us22/n728 ), .A2(\AES_ENC/us22/n727 ), .A3(\AES_ENC/us22/n726 ), .A4(\AES_ENC/us22/n725 ), .ZN(\AES_ENC/us22/n729 ) );
NAND2_X2 \AES_ENC/us22/U343  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n729 ), .ZN(\AES_ENC/us22/n730 ) );
NAND4_X2 \AES_ENC/us22/U342  ( .A1(\AES_ENC/us22/n733 ), .A2(\AES_ENC/us22/n732 ), .A3(\AES_ENC/us22/n731 ), .A4(\AES_ENC/us22/n730 ), .ZN(\AES_ENC/sa22_sub[1] ) );
NAND2_X2 \AES_ENC/us22/U341  ( .A1(\AES_ENC/sa22 [7]), .A2(\AES_ENC/us22/n611 ), .ZN(\AES_ENC/us22/n734 ) );
NAND2_X2 \AES_ENC/us22/U340  ( .A1(\AES_ENC/us22/n734 ), .A2(\AES_ENC/us22/n607 ), .ZN(\AES_ENC/us22/n738 ) );
OR4_X2 \AES_ENC/us22/U339  ( .A1(\AES_ENC/us22/n738 ), .A2(\AES_ENC/us22/n626 ), .A3(\AES_ENC/us22/n826 ), .A4(\AES_ENC/us22/n1121 ), .ZN(\AES_ENC/us22/n746 ) );
NAND2_X2 \AES_ENC/us22/U337  ( .A1(\AES_ENC/us22/n1100 ), .A2(\AES_ENC/us22/n587 ), .ZN(\AES_ENC/us22/n992 ) );
OR2_X2 \AES_ENC/us22/U336  ( .A1(\AES_ENC/us22/n610 ), .A2(\AES_ENC/us22/n735 ), .ZN(\AES_ENC/us22/n737 ) );
NAND2_X2 \AES_ENC/us22/U334  ( .A1(\AES_ENC/us22/n619 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n753 ) );
NAND2_X2 \AES_ENC/us22/U333  ( .A1(\AES_ENC/us22/n582 ), .A2(\AES_ENC/us22/n753 ), .ZN(\AES_ENC/us22/n1080 ) );
NAND2_X2 \AES_ENC/us22/U332  ( .A1(\AES_ENC/us22/n1048 ), .A2(\AES_ENC/us22/n576 ), .ZN(\AES_ENC/us22/n736 ) );
NAND2_X2 \AES_ENC/us22/U331  ( .A1(\AES_ENC/us22/n737 ), .A2(\AES_ENC/us22/n736 ), .ZN(\AES_ENC/us22/n739 ) );
NAND2_X2 \AES_ENC/us22/U330  ( .A1(\AES_ENC/us22/n739 ), .A2(\AES_ENC/us22/n738 ), .ZN(\AES_ENC/us22/n745 ) );
NAND2_X2 \AES_ENC/us22/U326  ( .A1(\AES_ENC/us22/n1096 ), .A2(\AES_ENC/us22/n590 ), .ZN(\AES_ENC/us22/n906 ) );
NAND4_X2 \AES_ENC/us22/U323  ( .A1(\AES_ENC/us22/n746 ), .A2(\AES_ENC/us22/n992 ), .A3(\AES_ENC/us22/n745 ), .A4(\AES_ENC/us22/n744 ), .ZN(\AES_ENC/us22/n747 ) );
NAND2_X2 \AES_ENC/us22/U322  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n747 ), .ZN(\AES_ENC/us22/n793 ) );
NAND2_X2 \AES_ENC/us22/U321  ( .A1(\AES_ENC/us22/n584 ), .A2(\AES_ENC/us22/n855 ), .ZN(\AES_ENC/us22/n748 ) );
NAND2_X2 \AES_ENC/us22/U320  ( .A1(\AES_ENC/us22/n956 ), .A2(\AES_ENC/us22/n748 ), .ZN(\AES_ENC/us22/n760 ) );
NAND2_X2 \AES_ENC/us22/U313  ( .A1(\AES_ENC/us22/n590 ), .A2(\AES_ENC/us22/n753 ), .ZN(\AES_ENC/us22/n1023 ) );
NAND4_X2 \AES_ENC/us22/U308  ( .A1(\AES_ENC/us22/n760 ), .A2(\AES_ENC/us22/n992 ), .A3(\AES_ENC/us22/n759 ), .A4(\AES_ENC/us22/n758 ), .ZN(\AES_ENC/us22/n761 ) );
NAND2_X2 \AES_ENC/us22/U307  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n761 ), .ZN(\AES_ENC/us22/n792 ) );
NAND2_X2 \AES_ENC/us22/U306  ( .A1(\AES_ENC/us22/n584 ), .A2(\AES_ENC/us22/n603 ), .ZN(\AES_ENC/us22/n989 ) );
NAND2_X2 \AES_ENC/us22/U305  ( .A1(\AES_ENC/us22/n1050 ), .A2(\AES_ENC/us22/n989 ), .ZN(\AES_ENC/us22/n777 ) );
NAND2_X2 \AES_ENC/us22/U304  ( .A1(\AES_ENC/us22/n1093 ), .A2(\AES_ENC/us22/n762 ), .ZN(\AES_ENC/us22/n776 ) );
XNOR2_X2 \AES_ENC/us22/U301  ( .A(\AES_ENC/sa22 [7]), .B(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n959 ) );
NAND4_X2 \AES_ENC/us22/U289  ( .A1(\AES_ENC/us22/n777 ), .A2(\AES_ENC/us22/n776 ), .A3(\AES_ENC/us22/n775 ), .A4(\AES_ENC/us22/n774 ), .ZN(\AES_ENC/us22/n778 ) );
NAND2_X2 \AES_ENC/us22/U288  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n778 ), .ZN(\AES_ENC/us22/n791 ) );
NAND2_X2 \AES_ENC/us22/U287  ( .A1(\AES_ENC/us22/n1056 ), .A2(\AES_ENC/us22/n1050 ), .ZN(\AES_ENC/us22/n788 ) );
NAND2_X2 \AES_ENC/us22/U286  ( .A1(\AES_ENC/us22/n1091 ), .A2(\AES_ENC/us22/n779 ), .ZN(\AES_ENC/us22/n787 ) );
NAND2_X2 \AES_ENC/us22/U285  ( .A1(\AES_ENC/us22/n956 ), .A2(\AES_ENC/sa22 [1]), .ZN(\AES_ENC/us22/n786 ) );
NAND4_X2 \AES_ENC/us22/U278  ( .A1(\AES_ENC/us22/n788 ), .A2(\AES_ENC/us22/n787 ), .A3(\AES_ENC/us22/n786 ), .A4(\AES_ENC/us22/n785 ), .ZN(\AES_ENC/us22/n789 ) );
NAND2_X2 \AES_ENC/us22/U277  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n789 ), .ZN(\AES_ENC/us22/n790 ) );
NAND4_X2 \AES_ENC/us22/U276  ( .A1(\AES_ENC/us22/n793 ), .A2(\AES_ENC/us22/n792 ), .A3(\AES_ENC/us22/n791 ), .A4(\AES_ENC/us22/n790 ), .ZN(\AES_ENC/sa22_sub[2] ) );
NAND2_X2 \AES_ENC/us22/U275  ( .A1(\AES_ENC/us22/n1059 ), .A2(\AES_ENC/us22/n794 ), .ZN(\AES_ENC/us22/n810 ) );
NAND2_X2 \AES_ENC/us22/U274  ( .A1(\AES_ENC/us22/n1049 ), .A2(\AES_ENC/us22/n956 ), .ZN(\AES_ENC/us22/n809 ) );
OR2_X2 \AES_ENC/us22/U266  ( .A1(\AES_ENC/us22/n1096 ), .A2(\AES_ENC/us22/n606 ), .ZN(\AES_ENC/us22/n802 ) );
NAND2_X2 \AES_ENC/us22/U265  ( .A1(\AES_ENC/us22/n1053 ), .A2(\AES_ENC/us22/n800 ), .ZN(\AES_ENC/us22/n801 ) );
NAND2_X2 \AES_ENC/us22/U264  ( .A1(\AES_ENC/us22/n802 ), .A2(\AES_ENC/us22/n801 ), .ZN(\AES_ENC/us22/n805 ) );
NAND4_X2 \AES_ENC/us22/U261  ( .A1(\AES_ENC/us22/n810 ), .A2(\AES_ENC/us22/n809 ), .A3(\AES_ENC/us22/n808 ), .A4(\AES_ENC/us22/n807 ), .ZN(\AES_ENC/us22/n811 ) );
NAND2_X2 \AES_ENC/us22/U260  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n811 ), .ZN(\AES_ENC/us22/n852 ) );
OR2_X2 \AES_ENC/us22/U259  ( .A1(\AES_ENC/us22/n1023 ), .A2(\AES_ENC/us22/n617 ), .ZN(\AES_ENC/us22/n819 ) );
OR2_X2 \AES_ENC/us22/U257  ( .A1(\AES_ENC/us22/n570 ), .A2(\AES_ENC/us22/n930 ), .ZN(\AES_ENC/us22/n818 ) );
NAND2_X2 \AES_ENC/us22/U256  ( .A1(\AES_ENC/us22/n1013 ), .A2(\AES_ENC/us22/n1094 ), .ZN(\AES_ENC/us22/n817 ) );
NAND4_X2 \AES_ENC/us22/U249  ( .A1(\AES_ENC/us22/n819 ), .A2(\AES_ENC/us22/n818 ), .A3(\AES_ENC/us22/n817 ), .A4(\AES_ENC/us22/n816 ), .ZN(\AES_ENC/us22/n820 ) );
NAND2_X2 \AES_ENC/us22/U248  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n820 ), .ZN(\AES_ENC/us22/n851 ) );
NAND2_X2 \AES_ENC/us22/U247  ( .A1(\AES_ENC/us22/n956 ), .A2(\AES_ENC/us22/n1080 ), .ZN(\AES_ENC/us22/n835 ) );
NAND2_X2 \AES_ENC/us22/U246  ( .A1(\AES_ENC/us22/n570 ), .A2(\AES_ENC/us22/n1030 ), .ZN(\AES_ENC/us22/n1047 ) );
OR2_X2 \AES_ENC/us22/U245  ( .A1(\AES_ENC/us22/n1047 ), .A2(\AES_ENC/us22/n612 ), .ZN(\AES_ENC/us22/n834 ) );
NAND2_X2 \AES_ENC/us22/U244  ( .A1(\AES_ENC/us22/n1072 ), .A2(\AES_ENC/us22/n589 ), .ZN(\AES_ENC/us22/n833 ) );
NAND4_X2 \AES_ENC/us22/U233  ( .A1(\AES_ENC/us22/n835 ), .A2(\AES_ENC/us22/n834 ), .A3(\AES_ENC/us22/n833 ), .A4(\AES_ENC/us22/n832 ), .ZN(\AES_ENC/us22/n836 ) );
NAND2_X2 \AES_ENC/us22/U232  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n836 ), .ZN(\AES_ENC/us22/n850 ) );
NAND2_X2 \AES_ENC/us22/U231  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n623 ), .ZN(\AES_ENC/us22/n847 ) );
NAND2_X2 \AES_ENC/us22/U230  ( .A1(\AES_ENC/us22/n1050 ), .A2(\AES_ENC/us22/n1071 ), .ZN(\AES_ENC/us22/n846 ) );
OR2_X2 \AES_ENC/us22/U224  ( .A1(\AES_ENC/us22/n1053 ), .A2(\AES_ENC/us22/n911 ), .ZN(\AES_ENC/us22/n1077 ) );
NAND4_X2 \AES_ENC/us22/U220  ( .A1(\AES_ENC/us22/n847 ), .A2(\AES_ENC/us22/n846 ), .A3(\AES_ENC/us22/n845 ), .A4(\AES_ENC/us22/n844 ), .ZN(\AES_ENC/us22/n848 ) );
NAND2_X2 \AES_ENC/us22/U219  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n848 ), .ZN(\AES_ENC/us22/n849 ) );
NAND4_X2 \AES_ENC/us22/U218  ( .A1(\AES_ENC/us22/n852 ), .A2(\AES_ENC/us22/n851 ), .A3(\AES_ENC/us22/n850 ), .A4(\AES_ENC/us22/n849 ), .ZN(\AES_ENC/sa22_sub[3] ) );
NAND2_X2 \AES_ENC/us22/U216  ( .A1(\AES_ENC/us22/n1009 ), .A2(\AES_ENC/us22/n1072 ), .ZN(\AES_ENC/us22/n862 ) );
NAND2_X2 \AES_ENC/us22/U215  ( .A1(\AES_ENC/us22/n603 ), .A2(\AES_ENC/us22/n577 ), .ZN(\AES_ENC/us22/n853 ) );
NAND2_X2 \AES_ENC/us22/U214  ( .A1(\AES_ENC/us22/n1050 ), .A2(\AES_ENC/us22/n853 ), .ZN(\AES_ENC/us22/n861 ) );
NAND4_X2 \AES_ENC/us22/U206  ( .A1(\AES_ENC/us22/n862 ), .A2(\AES_ENC/us22/n861 ), .A3(\AES_ENC/us22/n860 ), .A4(\AES_ENC/us22/n859 ), .ZN(\AES_ENC/us22/n863 ) );
NAND2_X2 \AES_ENC/us22/U205  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n863 ), .ZN(\AES_ENC/us22/n905 ) );
NAND2_X2 \AES_ENC/us22/U204  ( .A1(\AES_ENC/us22/n1010 ), .A2(\AES_ENC/us22/n989 ), .ZN(\AES_ENC/us22/n874 ) );
NAND2_X2 \AES_ENC/us22/U203  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n610 ), .ZN(\AES_ENC/us22/n864 ) );
NAND2_X2 \AES_ENC/us22/U202  ( .A1(\AES_ENC/us22/n929 ), .A2(\AES_ENC/us22/n864 ), .ZN(\AES_ENC/us22/n873 ) );
NAND4_X2 \AES_ENC/us22/U193  ( .A1(\AES_ENC/us22/n874 ), .A2(\AES_ENC/us22/n873 ), .A3(\AES_ENC/us22/n872 ), .A4(\AES_ENC/us22/n871 ), .ZN(\AES_ENC/us22/n875 ) );
NAND2_X2 \AES_ENC/us22/U192  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n875 ), .ZN(\AES_ENC/us22/n904 ) );
NAND2_X2 \AES_ENC/us22/U191  ( .A1(\AES_ENC/us22/n583 ), .A2(\AES_ENC/us22/n1050 ), .ZN(\AES_ENC/us22/n889 ) );
NAND2_X2 \AES_ENC/us22/U190  ( .A1(\AES_ENC/us22/n1093 ), .A2(\AES_ENC/us22/n587 ), .ZN(\AES_ENC/us22/n876 ) );
NAND2_X2 \AES_ENC/us22/U189  ( .A1(\AES_ENC/us22/n604 ), .A2(\AES_ENC/us22/n876 ), .ZN(\AES_ENC/us22/n877 ) );
NAND2_X2 \AES_ENC/us22/U188  ( .A1(\AES_ENC/us22/n877 ), .A2(\AES_ENC/us22/n623 ), .ZN(\AES_ENC/us22/n888 ) );
NAND4_X2 \AES_ENC/us22/U179  ( .A1(\AES_ENC/us22/n889 ), .A2(\AES_ENC/us22/n888 ), .A3(\AES_ENC/us22/n887 ), .A4(\AES_ENC/us22/n886 ), .ZN(\AES_ENC/us22/n890 ) );
NAND2_X2 \AES_ENC/us22/U178  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n890 ), .ZN(\AES_ENC/us22/n903 ) );
OR2_X2 \AES_ENC/us22/U177  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n1059 ), .ZN(\AES_ENC/us22/n900 ) );
NAND2_X2 \AES_ENC/us22/U176  ( .A1(\AES_ENC/us22/n1073 ), .A2(\AES_ENC/us22/n1047 ), .ZN(\AES_ENC/us22/n899 ) );
NAND2_X2 \AES_ENC/us22/U175  ( .A1(\AES_ENC/us22/n1094 ), .A2(\AES_ENC/us22/n595 ), .ZN(\AES_ENC/us22/n898 ) );
NAND4_X2 \AES_ENC/us22/U167  ( .A1(\AES_ENC/us22/n900 ), .A2(\AES_ENC/us22/n899 ), .A3(\AES_ENC/us22/n898 ), .A4(\AES_ENC/us22/n897 ), .ZN(\AES_ENC/us22/n901 ) );
NAND2_X2 \AES_ENC/us22/U166  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n901 ), .ZN(\AES_ENC/us22/n902 ) );
NAND4_X2 \AES_ENC/us22/U165  ( .A1(\AES_ENC/us22/n905 ), .A2(\AES_ENC/us22/n904 ), .A3(\AES_ENC/us22/n903 ), .A4(\AES_ENC/us22/n902 ), .ZN(\AES_ENC/sa22_sub[4] ) );
NAND2_X2 \AES_ENC/us22/U164  ( .A1(\AES_ENC/us22/n1094 ), .A2(\AES_ENC/us22/n599 ), .ZN(\AES_ENC/us22/n922 ) );
NAND2_X2 \AES_ENC/us22/U163  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n989 ), .ZN(\AES_ENC/us22/n921 ) );
NAND4_X2 \AES_ENC/us22/U151  ( .A1(\AES_ENC/us22/n922 ), .A2(\AES_ENC/us22/n921 ), .A3(\AES_ENC/us22/n920 ), .A4(\AES_ENC/us22/n919 ), .ZN(\AES_ENC/us22/n923 ) );
NAND2_X2 \AES_ENC/us22/U150  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n923 ), .ZN(\AES_ENC/us22/n972 ) );
NAND2_X2 \AES_ENC/us22/U149  ( .A1(\AES_ENC/us22/n582 ), .A2(\AES_ENC/us22/n619 ), .ZN(\AES_ENC/us22/n924 ) );
NAND2_X2 \AES_ENC/us22/U148  ( .A1(\AES_ENC/us22/n1073 ), .A2(\AES_ENC/us22/n924 ), .ZN(\AES_ENC/us22/n939 ) );
NAND2_X2 \AES_ENC/us22/U147  ( .A1(\AES_ENC/us22/n926 ), .A2(\AES_ENC/us22/n925 ), .ZN(\AES_ENC/us22/n927 ) );
NAND2_X2 \AES_ENC/us22/U146  ( .A1(\AES_ENC/us22/n606 ), .A2(\AES_ENC/us22/n927 ), .ZN(\AES_ENC/us22/n928 ) );
NAND2_X2 \AES_ENC/us22/U145  ( .A1(\AES_ENC/us22/n928 ), .A2(\AES_ENC/us22/n1080 ), .ZN(\AES_ENC/us22/n938 ) );
OR2_X2 \AES_ENC/us22/U144  ( .A1(\AES_ENC/us22/n1117 ), .A2(\AES_ENC/us22/n615 ), .ZN(\AES_ENC/us22/n937 ) );
NAND4_X2 \AES_ENC/us22/U139  ( .A1(\AES_ENC/us22/n939 ), .A2(\AES_ENC/us22/n938 ), .A3(\AES_ENC/us22/n937 ), .A4(\AES_ENC/us22/n936 ), .ZN(\AES_ENC/us22/n940 ) );
NAND2_X2 \AES_ENC/us22/U138  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n940 ), .ZN(\AES_ENC/us22/n971 ) );
OR2_X2 \AES_ENC/us22/U137  ( .A1(\AES_ENC/us22/n605 ), .A2(\AES_ENC/us22/n941 ), .ZN(\AES_ENC/us22/n954 ) );
NAND2_X2 \AES_ENC/us22/U136  ( .A1(\AES_ENC/us22/n1096 ), .A2(\AES_ENC/us22/n577 ), .ZN(\AES_ENC/us22/n942 ) );
NAND2_X2 \AES_ENC/us22/U135  ( .A1(\AES_ENC/us22/n1048 ), .A2(\AES_ENC/us22/n942 ), .ZN(\AES_ENC/us22/n943 ) );
NAND2_X2 \AES_ENC/us22/U134  ( .A1(\AES_ENC/us22/n612 ), .A2(\AES_ENC/us22/n943 ), .ZN(\AES_ENC/us22/n944 ) );
NAND2_X2 \AES_ENC/us22/U133  ( .A1(\AES_ENC/us22/n944 ), .A2(\AES_ENC/us22/n580 ), .ZN(\AES_ENC/us22/n953 ) );
NAND4_X2 \AES_ENC/us22/U125  ( .A1(\AES_ENC/us22/n954 ), .A2(\AES_ENC/us22/n953 ), .A3(\AES_ENC/us22/n952 ), .A4(\AES_ENC/us22/n951 ), .ZN(\AES_ENC/us22/n955 ) );
NAND2_X2 \AES_ENC/us22/U124  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n955 ), .ZN(\AES_ENC/us22/n970 ) );
NAND2_X2 \AES_ENC/us22/U123  ( .A1(\AES_ENC/us22/n1094 ), .A2(\AES_ENC/us22/n1071 ), .ZN(\AES_ENC/us22/n967 ) );
NAND2_X2 \AES_ENC/us22/U122  ( .A1(\AES_ENC/us22/n956 ), .A2(\AES_ENC/us22/n1030 ), .ZN(\AES_ENC/us22/n966 ) );
NAND4_X2 \AES_ENC/us22/U114  ( .A1(\AES_ENC/us22/n967 ), .A2(\AES_ENC/us22/n966 ), .A3(\AES_ENC/us22/n965 ), .A4(\AES_ENC/us22/n964 ), .ZN(\AES_ENC/us22/n968 ) );
NAND2_X2 \AES_ENC/us22/U113  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n968 ), .ZN(\AES_ENC/us22/n969 ) );
NAND4_X2 \AES_ENC/us22/U112  ( .A1(\AES_ENC/us22/n972 ), .A2(\AES_ENC/us22/n971 ), .A3(\AES_ENC/us22/n970 ), .A4(\AES_ENC/us22/n969 ), .ZN(\AES_ENC/sa22_sub[5] ) );
NAND2_X2 \AES_ENC/us22/U111  ( .A1(\AES_ENC/us22/n570 ), .A2(\AES_ENC/us22/n1097 ), .ZN(\AES_ENC/us22/n973 ) );
NAND2_X2 \AES_ENC/us22/U110  ( .A1(\AES_ENC/us22/n1073 ), .A2(\AES_ENC/us22/n973 ), .ZN(\AES_ENC/us22/n987 ) );
NAND2_X2 \AES_ENC/us22/U109  ( .A1(\AES_ENC/us22/n974 ), .A2(\AES_ENC/us22/n1077 ), .ZN(\AES_ENC/us22/n975 ) );
NAND2_X2 \AES_ENC/us22/U108  ( .A1(\AES_ENC/us22/n613 ), .A2(\AES_ENC/us22/n975 ), .ZN(\AES_ENC/us22/n976 ) );
NAND2_X2 \AES_ENC/us22/U107  ( .A1(\AES_ENC/us22/n977 ), .A2(\AES_ENC/us22/n976 ), .ZN(\AES_ENC/us22/n986 ) );
NAND4_X2 \AES_ENC/us22/U99  ( .A1(\AES_ENC/us22/n987 ), .A2(\AES_ENC/us22/n986 ), .A3(\AES_ENC/us22/n985 ), .A4(\AES_ENC/us22/n984 ), .ZN(\AES_ENC/us22/n988 ) );
NAND2_X2 \AES_ENC/us22/U98  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n988 ), .ZN(\AES_ENC/us22/n1044 ) );
NAND2_X2 \AES_ENC/us22/U97  ( .A1(\AES_ENC/us22/n1073 ), .A2(\AES_ENC/us22/n989 ), .ZN(\AES_ENC/us22/n1004 ) );
NAND2_X2 \AES_ENC/us22/U96  ( .A1(\AES_ENC/us22/n1092 ), .A2(\AES_ENC/us22/n619 ), .ZN(\AES_ENC/us22/n1003 ) );
NAND4_X2 \AES_ENC/us22/U85  ( .A1(\AES_ENC/us22/n1004 ), .A2(\AES_ENC/us22/n1003 ), .A3(\AES_ENC/us22/n1002 ), .A4(\AES_ENC/us22/n1001 ), .ZN(\AES_ENC/us22/n1005 ) );
NAND2_X2 \AES_ENC/us22/U84  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n1005 ), .ZN(\AES_ENC/us22/n1043 ) );
NAND2_X2 \AES_ENC/us22/U83  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n596 ), .ZN(\AES_ENC/us22/n1020 ) );
NAND2_X2 \AES_ENC/us22/U82  ( .A1(\AES_ENC/us22/n1050 ), .A2(\AES_ENC/us22/n624 ), .ZN(\AES_ENC/us22/n1019 ) );
NAND2_X2 \AES_ENC/us22/U77  ( .A1(\AES_ENC/us22/n1059 ), .A2(\AES_ENC/us22/n1114 ), .ZN(\AES_ENC/us22/n1012 ) );
NAND2_X2 \AES_ENC/us22/U76  ( .A1(\AES_ENC/us22/n1010 ), .A2(\AES_ENC/us22/n592 ), .ZN(\AES_ENC/us22/n1011 ) );
NAND2_X2 \AES_ENC/us22/U75  ( .A1(\AES_ENC/us22/n1012 ), .A2(\AES_ENC/us22/n1011 ), .ZN(\AES_ENC/us22/n1016 ) );
NAND4_X2 \AES_ENC/us22/U70  ( .A1(\AES_ENC/us22/n1020 ), .A2(\AES_ENC/us22/n1019 ), .A3(\AES_ENC/us22/n1018 ), .A4(\AES_ENC/us22/n1017 ), .ZN(\AES_ENC/us22/n1021 ) );
NAND2_X2 \AES_ENC/us22/U69  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n1021 ), .ZN(\AES_ENC/us22/n1042 ) );
NAND2_X2 \AES_ENC/us22/U68  ( .A1(\AES_ENC/us22/n1022 ), .A2(\AES_ENC/us22/n1093 ), .ZN(\AES_ENC/us22/n1039 ) );
NAND2_X2 \AES_ENC/us22/U67  ( .A1(\AES_ENC/us22/n1050 ), .A2(\AES_ENC/us22/n1023 ), .ZN(\AES_ENC/us22/n1038 ) );
NAND2_X2 \AES_ENC/us22/U66  ( .A1(\AES_ENC/us22/n1024 ), .A2(\AES_ENC/us22/n1071 ), .ZN(\AES_ENC/us22/n1037 ) );
AND2_X2 \AES_ENC/us22/U60  ( .A1(\AES_ENC/us22/n1030 ), .A2(\AES_ENC/us22/n602 ), .ZN(\AES_ENC/us22/n1078 ) );
NAND4_X2 \AES_ENC/us22/U56  ( .A1(\AES_ENC/us22/n1039 ), .A2(\AES_ENC/us22/n1038 ), .A3(\AES_ENC/us22/n1037 ), .A4(\AES_ENC/us22/n1036 ), .ZN(\AES_ENC/us22/n1040 ) );
NAND2_X2 \AES_ENC/us22/U55  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n1040 ), .ZN(\AES_ENC/us22/n1041 ) );
NAND4_X2 \AES_ENC/us22/U54  ( .A1(\AES_ENC/us22/n1044 ), .A2(\AES_ENC/us22/n1043 ), .A3(\AES_ENC/us22/n1042 ), .A4(\AES_ENC/us22/n1041 ), .ZN(\AES_ENC/sa22_sub[6] ) );
NAND2_X2 \AES_ENC/us22/U53  ( .A1(\AES_ENC/us22/n1072 ), .A2(\AES_ENC/us22/n1045 ), .ZN(\AES_ENC/us22/n1068 ) );
NAND2_X2 \AES_ENC/us22/U52  ( .A1(\AES_ENC/us22/n1046 ), .A2(\AES_ENC/us22/n582 ), .ZN(\AES_ENC/us22/n1067 ) );
NAND2_X2 \AES_ENC/us22/U51  ( .A1(\AES_ENC/us22/n1094 ), .A2(\AES_ENC/us22/n1047 ), .ZN(\AES_ENC/us22/n1066 ) );
NAND4_X2 \AES_ENC/us22/U40  ( .A1(\AES_ENC/us22/n1068 ), .A2(\AES_ENC/us22/n1067 ), .A3(\AES_ENC/us22/n1066 ), .A4(\AES_ENC/us22/n1065 ), .ZN(\AES_ENC/us22/n1069 ) );
NAND2_X2 \AES_ENC/us22/U39  ( .A1(\AES_ENC/us22/n1070 ), .A2(\AES_ENC/us22/n1069 ), .ZN(\AES_ENC/us22/n1135 ) );
NAND2_X2 \AES_ENC/us22/U38  ( .A1(\AES_ENC/us22/n1072 ), .A2(\AES_ENC/us22/n1071 ), .ZN(\AES_ENC/us22/n1088 ) );
NAND2_X2 \AES_ENC/us22/U37  ( .A1(\AES_ENC/us22/n1073 ), .A2(\AES_ENC/us22/n595 ), .ZN(\AES_ENC/us22/n1087 ) );
NAND4_X2 \AES_ENC/us22/U28  ( .A1(\AES_ENC/us22/n1088 ), .A2(\AES_ENC/us22/n1087 ), .A3(\AES_ENC/us22/n1086 ), .A4(\AES_ENC/us22/n1085 ), .ZN(\AES_ENC/us22/n1089 ) );
NAND2_X2 \AES_ENC/us22/U27  ( .A1(\AES_ENC/us22/n1090 ), .A2(\AES_ENC/us22/n1089 ), .ZN(\AES_ENC/us22/n1134 ) );
NAND2_X2 \AES_ENC/us22/U26  ( .A1(\AES_ENC/us22/n1091 ), .A2(\AES_ENC/us22/n1093 ), .ZN(\AES_ENC/us22/n1111 ) );
NAND2_X2 \AES_ENC/us22/U25  ( .A1(\AES_ENC/us22/n1092 ), .A2(\AES_ENC/us22/n1120 ), .ZN(\AES_ENC/us22/n1110 ) );
AND2_X2 \AES_ENC/us22/U22  ( .A1(\AES_ENC/us22/n1097 ), .A2(\AES_ENC/us22/n1096 ), .ZN(\AES_ENC/us22/n1098 ) );
NAND4_X2 \AES_ENC/us22/U14  ( .A1(\AES_ENC/us22/n1111 ), .A2(\AES_ENC/us22/n1110 ), .A3(\AES_ENC/us22/n1109 ), .A4(\AES_ENC/us22/n1108 ), .ZN(\AES_ENC/us22/n1112 ) );
NAND2_X2 \AES_ENC/us22/U13  ( .A1(\AES_ENC/us22/n1113 ), .A2(\AES_ENC/us22/n1112 ), .ZN(\AES_ENC/us22/n1133 ) );
NAND2_X2 \AES_ENC/us22/U12  ( .A1(\AES_ENC/us22/n1115 ), .A2(\AES_ENC/us22/n1114 ), .ZN(\AES_ENC/us22/n1129 ) );
OR2_X2 \AES_ENC/us22/U11  ( .A1(\AES_ENC/us22/n608 ), .A2(\AES_ENC/us22/n1116 ), .ZN(\AES_ENC/us22/n1128 ) );
NAND4_X2 \AES_ENC/us22/U3  ( .A1(\AES_ENC/us22/n1129 ), .A2(\AES_ENC/us22/n1128 ), .A3(\AES_ENC/us22/n1127 ), .A4(\AES_ENC/us22/n1126 ), .ZN(\AES_ENC/us22/n1130 ) );
NAND2_X2 \AES_ENC/us22/U2  ( .A1(\AES_ENC/us22/n1131 ), .A2(\AES_ENC/us22/n1130 ), .ZN(\AES_ENC/us22/n1132 ) );
NAND4_X2 \AES_ENC/us22/U1  ( .A1(\AES_ENC/us22/n1135 ), .A2(\AES_ENC/us22/n1134 ), .A3(\AES_ENC/us22/n1133 ), .A4(\AES_ENC/us22/n1132 ), .ZN(\AES_ENC/sa22_sub[7] ) );
INV_X4 \AES_ENC/us23/U575  ( .A(\AES_ENC/sa23 [0]), .ZN(\AES_ENC/us23/n627 ));
INV_X4 \AES_ENC/us23/U574  ( .A(\AES_ENC/us23/n1053 ), .ZN(\AES_ENC/us23/n625 ) );
INV_X4 \AES_ENC/us23/U573  ( .A(\AES_ENC/us23/n1103 ), .ZN(\AES_ENC/us23/n623 ) );
INV_X4 \AES_ENC/us23/U572  ( .A(\AES_ENC/us23/n1056 ), .ZN(\AES_ENC/us23/n622 ) );
INV_X4 \AES_ENC/us23/U571  ( .A(\AES_ENC/us23/n1102 ), .ZN(\AES_ENC/us23/n621 ) );
INV_X4 \AES_ENC/us23/U570  ( .A(\AES_ENC/us23/n1074 ), .ZN(\AES_ENC/us23/n620 ) );
INV_X4 \AES_ENC/us23/U569  ( .A(\AES_ENC/us23/n929 ), .ZN(\AES_ENC/us23/n619 ) );
INV_X4 \AES_ENC/us23/U568  ( .A(\AES_ENC/us23/n1091 ), .ZN(\AES_ENC/us23/n618 ) );
INV_X4 \AES_ENC/us23/U567  ( .A(\AES_ENC/us23/n826 ), .ZN(\AES_ENC/us23/n617 ) );
INV_X4 \AES_ENC/us23/U566  ( .A(\AES_ENC/us23/n1031 ), .ZN(\AES_ENC/us23/n616 ) );
INV_X4 \AES_ENC/us23/U565  ( .A(\AES_ENC/us23/n1054 ), .ZN(\AES_ENC/us23/n615 ) );
INV_X4 \AES_ENC/us23/U564  ( .A(\AES_ENC/us23/n1025 ), .ZN(\AES_ENC/us23/n614 ) );
INV_X4 \AES_ENC/us23/U563  ( .A(\AES_ENC/us23/n990 ), .ZN(\AES_ENC/us23/n613 ) );
INV_X4 \AES_ENC/us23/U562  ( .A(\AES_ENC/sa23 [4]), .ZN(\AES_ENC/us23/n612 ));
INV_X4 \AES_ENC/us23/U561  ( .A(\AES_ENC/us23/n881 ), .ZN(\AES_ENC/us23/n611 ) );
INV_X4 \AES_ENC/us23/U560  ( .A(\AES_ENC/us23/n1022 ), .ZN(\AES_ENC/us23/n610 ) );
INV_X4 \AES_ENC/us23/U559  ( .A(\AES_ENC/us23/n1120 ), .ZN(\AES_ENC/us23/n609 ) );
INV_X4 \AES_ENC/us23/U558  ( .A(\AES_ENC/us23/n977 ), .ZN(\AES_ENC/us23/n608 ) );
INV_X4 \AES_ENC/us23/U557  ( .A(\AES_ENC/us23/n926 ), .ZN(\AES_ENC/us23/n607 ) );
INV_X4 \AES_ENC/us23/U556  ( .A(\AES_ENC/us23/n910 ), .ZN(\AES_ENC/us23/n606 ) );
INV_X4 \AES_ENC/us23/U555  ( .A(\AES_ENC/us23/n1121 ), .ZN(\AES_ENC/us23/n605 ) );
INV_X4 \AES_ENC/us23/U554  ( .A(\AES_ENC/us23/n1009 ), .ZN(\AES_ENC/us23/n604 ) );
INV_X4 \AES_ENC/us23/U553  ( .A(\AES_ENC/us23/n1080 ), .ZN(\AES_ENC/us23/n602 ) );
INV_X4 \AES_ENC/us23/U552  ( .A(\AES_ENC/us23/n821 ), .ZN(\AES_ENC/us23/n600 ) );
INV_X4 \AES_ENC/us23/U551  ( .A(\AES_ENC/us23/n1013 ), .ZN(\AES_ENC/us23/n599 ) );
INV_X4 \AES_ENC/us23/U550  ( .A(\AES_ENC/us23/n1058 ), .ZN(\AES_ENC/us23/n598 ) );
INV_X4 \AES_ENC/us23/U549  ( .A(\AES_ENC/us23/n906 ), .ZN(\AES_ENC/us23/n597 ) );
INV_X4 \AES_ENC/us23/U548  ( .A(\AES_ENC/us23/n1048 ), .ZN(\AES_ENC/us23/n595 ) );
INV_X4 \AES_ENC/us23/U547  ( .A(\AES_ENC/us23/n974 ), .ZN(\AES_ENC/us23/n594 ) );
INV_X4 \AES_ENC/us23/U546  ( .A(\AES_ENC/sa23 [2]), .ZN(\AES_ENC/us23/n593 ));
INV_X4 \AES_ENC/us23/U545  ( .A(\AES_ENC/us23/n800 ), .ZN(\AES_ENC/us23/n592 ) );
INV_X4 \AES_ENC/us23/U544  ( .A(\AES_ENC/us23/n925 ), .ZN(\AES_ENC/us23/n591 ) );
INV_X4 \AES_ENC/us23/U543  ( .A(\AES_ENC/us23/n824 ), .ZN(\AES_ENC/us23/n590 ) );
INV_X4 \AES_ENC/us23/U542  ( .A(\AES_ENC/us23/n959 ), .ZN(\AES_ENC/us23/n589 ) );
INV_X4 \AES_ENC/us23/U541  ( .A(\AES_ENC/us23/n779 ), .ZN(\AES_ENC/us23/n588 ) );
INV_X4 \AES_ENC/us23/U540  ( .A(\AES_ENC/us23/n794 ), .ZN(\AES_ENC/us23/n585 ) );
INV_X4 \AES_ENC/us23/U539  ( .A(\AES_ENC/us23/n880 ), .ZN(\AES_ENC/us23/n583 ) );
INV_X4 \AES_ENC/us23/U538  ( .A(\AES_ENC/sa23 [7]), .ZN(\AES_ENC/us23/n581 ));
INV_X4 \AES_ENC/us23/U537  ( .A(\AES_ENC/us23/n992 ), .ZN(\AES_ENC/us23/n578 ) );
INV_X4 \AES_ENC/us23/U536  ( .A(\AES_ENC/us23/n1114 ), .ZN(\AES_ENC/us23/n577 ) );
INV_X4 \AES_ENC/us23/U535  ( .A(\AES_ENC/us23/n1092 ), .ZN(\AES_ENC/us23/n574 ) );
NOR2_X2 \AES_ENC/us23/U534  ( .A1(\AES_ENC/sa23 [0]), .A2(\AES_ENC/sa23 [6]),.ZN(\AES_ENC/us23/n1090 ) );
NOR2_X2 \AES_ENC/us23/U533  ( .A1(\AES_ENC/us23/n627 ), .A2(\AES_ENC/sa23 [6]), .ZN(\AES_ENC/us23/n1070 ) );
NOR2_X2 \AES_ENC/us23/U532  ( .A1(\AES_ENC/sa23 [4]), .A2(\AES_ENC/sa23 [3]),.ZN(\AES_ENC/us23/n1025 ) );
INV_X4 \AES_ENC/us23/U531  ( .A(\AES_ENC/us23/n569 ), .ZN(\AES_ENC/us23/n572 ) );
NOR2_X2 \AES_ENC/us23/U530  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n765 ) );
NOR2_X2 \AES_ENC/us23/U529  ( .A1(\AES_ENC/sa23 [4]), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n764 ) );
NOR2_X2 \AES_ENC/us23/U528  ( .A1(\AES_ENC/us23/n765 ), .A2(\AES_ENC/us23/n764 ), .ZN(\AES_ENC/us23/n766 ) );
NOR2_X2 \AES_ENC/us23/U527  ( .A1(\AES_ENC/us23/n766 ), .A2(\AES_ENC/us23/n589 ), .ZN(\AES_ENC/us23/n767 ) );
INV_X4 \AES_ENC/us23/U526  ( .A(\AES_ENC/sa23 [3]), .ZN(\AES_ENC/us23/n624 ));
NAND3_X2 \AES_ENC/us23/U525  ( .A1(\AES_ENC/us23/n652 ), .A2(\AES_ENC/us23/n596 ), .A3(\AES_ENC/sa23 [7]), .ZN(\AES_ENC/us23/n653 ));
NOR2_X2 \AES_ENC/us23/U524  ( .A1(\AES_ENC/us23/n593 ), .A2(\AES_ENC/sa23 [5]), .ZN(\AES_ENC/us23/n925 ) );
NOR2_X2 \AES_ENC/us23/U523  ( .A1(\AES_ENC/sa23 [5]), .A2(\AES_ENC/sa23 [2]),.ZN(\AES_ENC/us23/n974 ) );
INV_X4 \AES_ENC/us23/U522  ( .A(\AES_ENC/sa23 [5]), .ZN(\AES_ENC/us23/n596 ));
NOR2_X2 \AES_ENC/us23/U521  ( .A1(\AES_ENC/us23/n593 ), .A2(\AES_ENC/sa23 [7]), .ZN(\AES_ENC/us23/n779 ) );
NAND3_X2 \AES_ENC/us23/U520  ( .A1(\AES_ENC/us23/n679 ), .A2(\AES_ENC/us23/n678 ), .A3(\AES_ENC/us23/n677 ), .ZN(\AES_ENC/sa23_sub[0] ) );
NOR2_X2 \AES_ENC/us23/U519  ( .A1(\AES_ENC/us23/n596 ), .A2(\AES_ENC/sa23 [2]), .ZN(\AES_ENC/us23/n1048 ) );
NOR3_X2 \AES_ENC/us23/U518  ( .A1(\AES_ENC/us23/n581 ), .A2(\AES_ENC/sa23 [5]), .A3(\AES_ENC/us23/n704 ), .ZN(\AES_ENC/us23/n706 ));
NOR2_X2 \AES_ENC/us23/U517  ( .A1(\AES_ENC/us23/n1117 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n707 ) );
NOR2_X2 \AES_ENC/us23/U516  ( .A1(\AES_ENC/sa23 [4]), .A2(\AES_ENC/us23/n574 ), .ZN(\AES_ENC/us23/n705 ) );
NOR3_X2 \AES_ENC/us23/U515  ( .A1(\AES_ENC/us23/n707 ), .A2(\AES_ENC/us23/n706 ), .A3(\AES_ENC/us23/n705 ), .ZN(\AES_ENC/us23/n713 ) );
NOR4_X2 \AES_ENC/us23/U512  ( .A1(\AES_ENC/us23/n633 ), .A2(\AES_ENC/us23/n632 ), .A3(\AES_ENC/us23/n631 ), .A4(\AES_ENC/us23/n630 ), .ZN(\AES_ENC/us23/n634 ) );
NOR2_X2 \AES_ENC/us23/U510  ( .A1(\AES_ENC/us23/n629 ), .A2(\AES_ENC/us23/n628 ), .ZN(\AES_ENC/us23/n635 ) );
NAND3_X2 \AES_ENC/us23/U509  ( .A1(\AES_ENC/sa23 [2]), .A2(\AES_ENC/sa23 [7]), .A3(\AES_ENC/us23/n1059 ), .ZN(\AES_ENC/us23/n636 ) );
NOR2_X2 \AES_ENC/us23/U508  ( .A1(\AES_ENC/sa23 [7]), .A2(\AES_ENC/sa23 [2]),.ZN(\AES_ENC/us23/n794 ) );
NOR2_X2 \AES_ENC/us23/U507  ( .A1(\AES_ENC/sa23 [4]), .A2(\AES_ENC/sa23 [1]),.ZN(\AES_ENC/us23/n1102 ) );
NOR2_X2 \AES_ENC/us23/U506  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/sa23 [3]), .ZN(\AES_ENC/us23/n1053 ) );
NOR2_X2 \AES_ENC/us23/U505  ( .A1(\AES_ENC/us23/n588 ), .A2(\AES_ENC/sa23 [5]), .ZN(\AES_ENC/us23/n1024 ) );
NOR2_X2 \AES_ENC/us23/U504  ( .A1(\AES_ENC/us23/n577 ), .A2(\AES_ENC/sa23 [2]), .ZN(\AES_ENC/us23/n1093 ) );
NOR2_X2 \AES_ENC/us23/U503  ( .A1(\AES_ENC/us23/n585 ), .A2(\AES_ENC/sa23 [5]), .ZN(\AES_ENC/us23/n1094 ) );
NOR2_X2 \AES_ENC/us23/U502  ( .A1(\AES_ENC/us23/n612 ), .A2(\AES_ENC/sa23 [3]), .ZN(\AES_ENC/us23/n931 ) );
INV_X4 \AES_ENC/us23/U501  ( .A(\AES_ENC/us23/n570 ), .ZN(\AES_ENC/us23/n573 ) );
NOR2_X2 \AES_ENC/us23/U500  ( .A1(\AES_ENC/us23/n1053 ), .A2(\AES_ENC/us23/n1095 ), .ZN(\AES_ENC/us23/n639 ) );
NOR3_X2 \AES_ENC/us23/U499  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n573 ), .A3(\AES_ENC/us23/n1074 ), .ZN(\AES_ENC/us23/n641 ) );
NOR2_X2 \AES_ENC/us23/U498  ( .A1(\AES_ENC/us23/n639 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n640 ) );
NOR2_X2 \AES_ENC/us23/U497  ( .A1(\AES_ENC/us23/n641 ), .A2(\AES_ENC/us23/n640 ), .ZN(\AES_ENC/us23/n646 ) );
NOR3_X2 \AES_ENC/us23/U496  ( .A1(\AES_ENC/us23/n995 ), .A2(\AES_ENC/us23/n578 ), .A3(\AES_ENC/us23/n994 ), .ZN(\AES_ENC/us23/n1002 ) );
NOR2_X2 \AES_ENC/us23/U495  ( .A1(\AES_ENC/us23/n909 ), .A2(\AES_ENC/us23/n908 ), .ZN(\AES_ENC/us23/n920 ) );
NOR2_X2 \AES_ENC/us23/U494  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n823 ) );
NOR2_X2 \AES_ENC/us23/U492  ( .A1(\AES_ENC/us23/n612 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n822 ) );
NOR2_X2 \AES_ENC/us23/U491  ( .A1(\AES_ENC/us23/n823 ), .A2(\AES_ENC/us23/n822 ), .ZN(\AES_ENC/us23/n825 ) );
NOR2_X2 \AES_ENC/us23/U490  ( .A1(\AES_ENC/sa23 [1]), .A2(\AES_ENC/us23/n601 ), .ZN(\AES_ENC/us23/n913 ) );
NOR2_X2 \AES_ENC/us23/U489  ( .A1(\AES_ENC/us23/n913 ), .A2(\AES_ENC/us23/n1091 ), .ZN(\AES_ENC/us23/n914 ) );
NOR2_X2 \AES_ENC/us23/U488  ( .A1(\AES_ENC/us23/n826 ), .A2(\AES_ENC/us23/n572 ), .ZN(\AES_ENC/us23/n827 ) );
NOR3_X2 \AES_ENC/us23/U487  ( .A1(\AES_ENC/us23/n769 ), .A2(\AES_ENC/us23/n768 ), .A3(\AES_ENC/us23/n767 ), .ZN(\AES_ENC/us23/n775 ) );
NOR2_X2 \AES_ENC/us23/U486  ( .A1(\AES_ENC/us23/n1056 ), .A2(\AES_ENC/us23/n1053 ), .ZN(\AES_ENC/us23/n749 ) );
NOR2_X2 \AES_ENC/us23/U483  ( .A1(\AES_ENC/us23/n749 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n752 ) );
INV_X4 \AES_ENC/us23/U482  ( .A(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n626 ));
NOR2_X2 \AES_ENC/us23/U480  ( .A1(\AES_ENC/us23/n1054 ), .A2(\AES_ENC/us23/n1053 ), .ZN(\AES_ENC/us23/n1055 ) );
OR2_X4 \AES_ENC/us23/U479  ( .A1(\AES_ENC/us23/n1094 ), .A2(\AES_ENC/us23/n1093 ), .ZN(\AES_ENC/us23/n571 ) );
AND2_X2 \AES_ENC/us23/U478  ( .A1(\AES_ENC/us23/n571 ), .A2(\AES_ENC/us23/n1095 ), .ZN(\AES_ENC/us23/n1101 ) );
NOR2_X2 \AES_ENC/us23/U477  ( .A1(\AES_ENC/us23/n1074 ), .A2(\AES_ENC/us23/n931 ), .ZN(\AES_ENC/us23/n796 ) );
NOR2_X2 \AES_ENC/us23/U474  ( .A1(\AES_ENC/us23/n796 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n797 ) );
NOR2_X2 \AES_ENC/us23/U473  ( .A1(\AES_ENC/us23/n932 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n933 ) );
NOR2_X2 \AES_ENC/us23/U472  ( .A1(\AES_ENC/us23/n929 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n935 ) );
NOR2_X2 \AES_ENC/us23/U471  ( .A1(\AES_ENC/us23/n931 ), .A2(\AES_ENC/us23/n930 ), .ZN(\AES_ENC/us23/n934 ) );
NOR3_X2 \AES_ENC/us23/U470  ( .A1(\AES_ENC/us23/n935 ), .A2(\AES_ENC/us23/n934 ), .A3(\AES_ENC/us23/n933 ), .ZN(\AES_ENC/us23/n936 ) );
NOR2_X2 \AES_ENC/us23/U469  ( .A1(\AES_ENC/us23/n612 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n1075 ) );
NOR2_X2 \AES_ENC/us23/U468  ( .A1(\AES_ENC/us23/n572 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n949 ) );
NOR2_X2 \AES_ENC/us23/U467  ( .A1(\AES_ENC/us23/n1049 ), .A2(\AES_ENC/us23/n595 ), .ZN(\AES_ENC/us23/n1051 ) );
NOR2_X2 \AES_ENC/us23/U466  ( .A1(\AES_ENC/us23/n1051 ), .A2(\AES_ENC/us23/n1050 ), .ZN(\AES_ENC/us23/n1052 ) );
NOR2_X2 \AES_ENC/us23/U465  ( .A1(\AES_ENC/us23/n1052 ), .A2(\AES_ENC/us23/n604 ), .ZN(\AES_ENC/us23/n1064 ) );
NOR2_X2 \AES_ENC/us23/U464  ( .A1(\AES_ENC/sa23 [1]), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n631 ) );
NOR2_X2 \AES_ENC/us23/U463  ( .A1(\AES_ENC/us23/n1025 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n980 ) );
NOR2_X2 \AES_ENC/us23/U462  ( .A1(\AES_ENC/us23/n1073 ), .A2(\AES_ENC/us23/n1094 ), .ZN(\AES_ENC/us23/n795 ) );
NOR2_X2 \AES_ENC/us23/U461  ( .A1(\AES_ENC/us23/n795 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n799 ) );
NOR2_X2 \AES_ENC/us23/U460  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n981 ) );
NOR2_X2 \AES_ENC/us23/U459  ( .A1(\AES_ENC/us23/n1102 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n643 ) );
NOR2_X2 \AES_ENC/us23/U458  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n624 ), .ZN(\AES_ENC/us23/n642 ) );
NOR2_X2 \AES_ENC/us23/U455  ( .A1(\AES_ENC/us23/n911 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n644 ) );
NOR4_X2 \AES_ENC/us23/U448  ( .A1(\AES_ENC/us23/n644 ), .A2(\AES_ENC/us23/n643 ), .A3(\AES_ENC/us23/n804 ), .A4(\AES_ENC/us23/n642 ), .ZN(\AES_ENC/us23/n645 ) );
NOR2_X2 \AES_ENC/us23/U447  ( .A1(\AES_ENC/us23/n1102 ), .A2(\AES_ENC/us23/n910 ), .ZN(\AES_ENC/us23/n932 ) );
NOR2_X2 \AES_ENC/us23/U442  ( .A1(\AES_ENC/us23/n1102 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n755 ) );
NOR2_X2 \AES_ENC/us23/U441  ( .A1(\AES_ENC/us23/n931 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n743 ) );
NOR2_X2 \AES_ENC/us23/U438  ( .A1(\AES_ENC/us23/n1072 ), .A2(\AES_ENC/us23/n1094 ), .ZN(\AES_ENC/us23/n930 ) );
NOR2_X2 \AES_ENC/us23/U435  ( .A1(\AES_ENC/us23/n1074 ), .A2(\AES_ENC/us23/n1025 ), .ZN(\AES_ENC/us23/n891 ) );
NOR2_X2 \AES_ENC/us23/U434  ( .A1(\AES_ENC/us23/n891 ), .A2(\AES_ENC/us23/n591 ), .ZN(\AES_ENC/us23/n894 ) );
NOR3_X2 \AES_ENC/us23/U433  ( .A1(\AES_ENC/us23/n601 ), .A2(\AES_ENC/sa23 [1]), .A3(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n683 ));
INV_X4 \AES_ENC/us23/U428  ( .A(\AES_ENC/us23/n931 ), .ZN(\AES_ENC/us23/n601 ) );
NOR2_X2 \AES_ENC/us23/U427  ( .A1(\AES_ENC/us23/n996 ), .A2(\AES_ENC/us23/n931 ), .ZN(\AES_ENC/us23/n704 ) );
NOR2_X2 \AES_ENC/us23/U421  ( .A1(\AES_ENC/us23/n931 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n685 ) );
NOR2_X2 \AES_ENC/us23/U420  ( .A1(\AES_ENC/us23/n1029 ), .A2(\AES_ENC/us23/n1025 ), .ZN(\AES_ENC/us23/n1079 ) );
NOR3_X2 \AES_ENC/us23/U419  ( .A1(\AES_ENC/us23/n620 ), .A2(\AES_ENC/us23/n1025 ), .A3(\AES_ENC/us23/n594 ), .ZN(\AES_ENC/us23/n945 ) );
NOR2_X2 \AES_ENC/us23/U418  ( .A1(\AES_ENC/us23/n596 ), .A2(\AES_ENC/us23/n593 ), .ZN(\AES_ENC/us23/n800 ) );
NOR3_X2 \AES_ENC/us23/U417  ( .A1(\AES_ENC/us23/n598 ), .A2(\AES_ENC/us23/n581 ), .A3(\AES_ENC/us23/n593 ), .ZN(\AES_ENC/us23/n798 ) );
NOR3_X2 \AES_ENC/us23/U416  ( .A1(\AES_ENC/us23/n592 ), .A2(\AES_ENC/us23/n572 ), .A3(\AES_ENC/us23/n589 ), .ZN(\AES_ENC/us23/n962 ) );
NOR3_X2 \AES_ENC/us23/U415  ( .A1(\AES_ENC/us23/n959 ), .A2(\AES_ENC/us23/n572 ), .A3(\AES_ENC/us23/n591 ), .ZN(\AES_ENC/us23/n768 ) );
NOR3_X2 \AES_ENC/us23/U414  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n572 ), .A3(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n694 ) );
NOR3_X2 \AES_ENC/us23/U413  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n572 ), .A3(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n895 ) );
NOR3_X2 \AES_ENC/us23/U410  ( .A1(\AES_ENC/us23/n1008 ), .A2(\AES_ENC/us23/n1007 ), .A3(\AES_ENC/us23/n1006 ), .ZN(\AES_ENC/us23/n1018 ) );
NOR4_X2 \AES_ENC/us23/U409  ( .A1(\AES_ENC/us23/n806 ), .A2(\AES_ENC/us23/n805 ), .A3(\AES_ENC/us23/n804 ), .A4(\AES_ENC/us23/n803 ), .ZN(\AES_ENC/us23/n807 ) );
NOR3_X2 \AES_ENC/us23/U406  ( .A1(\AES_ENC/us23/n799 ), .A2(\AES_ENC/us23/n798 ), .A3(\AES_ENC/us23/n797 ), .ZN(\AES_ENC/us23/n808 ) );
NOR4_X2 \AES_ENC/us23/U405  ( .A1(\AES_ENC/us23/n843 ), .A2(\AES_ENC/us23/n842 ), .A3(\AES_ENC/us23/n841 ), .A4(\AES_ENC/us23/n840 ), .ZN(\AES_ENC/us23/n844 ) );
NOR2_X2 \AES_ENC/us23/U404  ( .A1(\AES_ENC/us23/n669 ), .A2(\AES_ENC/us23/n668 ), .ZN(\AES_ENC/us23/n673 ) );
NOR4_X2 \AES_ENC/us23/U403  ( .A1(\AES_ENC/us23/n946 ), .A2(\AES_ENC/us23/n1046 ), .A3(\AES_ENC/us23/n671 ), .A4(\AES_ENC/us23/n670 ), .ZN(\AES_ENC/us23/n672 ) );
NOR4_X2 \AES_ENC/us23/U401  ( .A1(\AES_ENC/us23/n711 ), .A2(\AES_ENC/us23/n710 ), .A3(\AES_ENC/us23/n709 ), .A4(\AES_ENC/us23/n708 ), .ZN(\AES_ENC/us23/n712 ) );
NOR4_X2 \AES_ENC/us23/U400  ( .A1(\AES_ENC/us23/n963 ), .A2(\AES_ENC/us23/n962 ), .A3(\AES_ENC/us23/n961 ), .A4(\AES_ENC/us23/n960 ), .ZN(\AES_ENC/us23/n964 ) );
NOR3_X2 \AES_ENC/us23/U399  ( .A1(\AES_ENC/us23/n1101 ), .A2(\AES_ENC/us23/n1100 ), .A3(\AES_ENC/us23/n1099 ), .ZN(\AES_ENC/us23/n1109 ) );
NOR3_X2 \AES_ENC/us23/U398  ( .A1(\AES_ENC/us23/n743 ), .A2(\AES_ENC/us23/n742 ), .A3(\AES_ENC/us23/n741 ), .ZN(\AES_ENC/us23/n744 ) );
NOR2_X2 \AES_ENC/us23/U397  ( .A1(\AES_ENC/us23/n697 ), .A2(\AES_ENC/us23/n658 ), .ZN(\AES_ENC/us23/n659 ) );
NOR2_X2 \AES_ENC/us23/U396  ( .A1(\AES_ENC/us23/n1078 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n1033 ) );
NOR2_X2 \AES_ENC/us23/U393  ( .A1(\AES_ENC/us23/n1031 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n1032 ) );
NOR3_X2 \AES_ENC/us23/U390  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n1025 ), .A3(\AES_ENC/us23/n1074 ), .ZN(\AES_ENC/us23/n1035 ) );
NOR4_X2 \AES_ENC/us23/U389  ( .A1(\AES_ENC/us23/n1035 ), .A2(\AES_ENC/us23/n1034 ), .A3(\AES_ENC/us23/n1033 ), .A4(\AES_ENC/us23/n1032 ), .ZN(\AES_ENC/us23/n1036 ) );
NOR2_X2 \AES_ENC/us23/U388  ( .A1(\AES_ENC/us23/n611 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n885 ) );
NOR2_X2 \AES_ENC/us23/U387  ( .A1(\AES_ENC/us23/n601 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n882 ) );
NOR2_X2 \AES_ENC/us23/U386  ( .A1(\AES_ENC/us23/n1053 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n884 ) );
NOR4_X2 \AES_ENC/us23/U385  ( .A1(\AES_ENC/us23/n885 ), .A2(\AES_ENC/us23/n884 ), .A3(\AES_ENC/us23/n883 ), .A4(\AES_ENC/us23/n882 ), .ZN(\AES_ENC/us23/n886 ) );
NOR2_X2 \AES_ENC/us23/U384  ( .A1(\AES_ENC/us23/n825 ), .A2(\AES_ENC/us23/n590 ), .ZN(\AES_ENC/us23/n830 ) );
NOR2_X2 \AES_ENC/us23/U383  ( .A1(\AES_ENC/us23/n827 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n829 ) );
NOR2_X2 \AES_ENC/us23/U382  ( .A1(\AES_ENC/us23/n572 ), .A2(\AES_ENC/us23/n574 ), .ZN(\AES_ENC/us23/n828 ) );
NOR4_X2 \AES_ENC/us23/U374  ( .A1(\AES_ENC/us23/n831 ), .A2(\AES_ENC/us23/n830 ), .A3(\AES_ENC/us23/n829 ), .A4(\AES_ENC/us23/n828 ), .ZN(\AES_ENC/us23/n832 ) );
NOR2_X2 \AES_ENC/us23/U373  ( .A1(\AES_ENC/us23/n587 ), .A2(\AES_ENC/us23/n603 ), .ZN(\AES_ENC/us23/n1104 ) );
NOR2_X2 \AES_ENC/us23/U372  ( .A1(\AES_ENC/us23/n1102 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n1106 ) );
NOR2_X2 \AES_ENC/us23/U370  ( .A1(\AES_ENC/us23/n1103 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n1105 ) );
NOR4_X2 \AES_ENC/us23/U369  ( .A1(\AES_ENC/us23/n1107 ), .A2(\AES_ENC/us23/n1106 ), .A3(\AES_ENC/us23/n1105 ), .A4(\AES_ENC/us23/n1104 ), .ZN(\AES_ENC/us23/n1108 ) );
NOR3_X2 \AES_ENC/us23/U368  ( .A1(\AES_ENC/us23/n959 ), .A2(\AES_ENC/us23/n624 ), .A3(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n963 ) );
NOR2_X2 \AES_ENC/us23/U367  ( .A1(\AES_ENC/us23/n596 ), .A2(\AES_ENC/us23/n581 ), .ZN(\AES_ENC/us23/n1114 ) );
INV_X4 \AES_ENC/us23/U366  ( .A(\AES_ENC/us23/n1024 ), .ZN(\AES_ENC/us23/n587 ) );
NOR3_X2 \AES_ENC/us23/U365  ( .A1(\AES_ENC/us23/n910 ), .A2(\AES_ENC/us23/n1059 ), .A3(\AES_ENC/us23/n593 ), .ZN(\AES_ENC/us23/n1115 ) );
INV_X4 \AES_ENC/us23/U364  ( .A(\AES_ENC/us23/n1094 ), .ZN(\AES_ENC/us23/n584 ) );
NOR2_X2 \AES_ENC/us23/U363  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n931 ), .ZN(\AES_ENC/us23/n1100 ) );
INV_X4 \AES_ENC/us23/U354  ( .A(\AES_ENC/us23/n1093 ), .ZN(\AES_ENC/us23/n575 ) );
NOR2_X2 \AES_ENC/us23/U353  ( .A1(\AES_ENC/us23/n569 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n929 ) );
NOR2_X2 \AES_ENC/us23/U352  ( .A1(\AES_ENC/us23/n609 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n926 ) );
NOR2_X2 \AES_ENC/us23/U351  ( .A1(\AES_ENC/us23/n572 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n1095 ) );
NOR2_X2 \AES_ENC/us23/U350  ( .A1(\AES_ENC/us23/n591 ), .A2(\AES_ENC/us23/n581 ), .ZN(\AES_ENC/us23/n1010 ) );
NOR2_X2 \AES_ENC/us23/U349  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n1103 ) );
NOR2_X2 \AES_ENC/us23/U348  ( .A1(\AES_ENC/us23/n614 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n1059 ) );
NOR2_X2 \AES_ENC/us23/U347  ( .A1(\AES_ENC/sa23 [1]), .A2(\AES_ENC/us23/n1120 ), .ZN(\AES_ENC/us23/n1022 ) );
NOR2_X2 \AES_ENC/us23/U346  ( .A1(\AES_ENC/us23/n605 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n911 ) );
NOR2_X2 \AES_ENC/us23/U345  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/us23/n1025 ), .ZN(\AES_ENC/us23/n826 ) );
NOR2_X2 \AES_ENC/us23/U338  ( .A1(\AES_ENC/us23/n596 ), .A2(\AES_ENC/us23/n588 ), .ZN(\AES_ENC/us23/n1072 ) );
NOR2_X2 \AES_ENC/us23/U335  ( .A1(\AES_ENC/us23/n581 ), .A2(\AES_ENC/us23/n594 ), .ZN(\AES_ENC/us23/n956 ) );
NOR2_X2 \AES_ENC/us23/U329  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/us23/n612 ), .ZN(\AES_ENC/us23/n1121 ) );
NOR2_X2 \AES_ENC/us23/U328  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/us23/n612 ), .ZN(\AES_ENC/us23/n1058 ) );
NOR2_X2 \AES_ENC/us23/U327  ( .A1(\AES_ENC/us23/n577 ), .A2(\AES_ENC/us23/n593 ), .ZN(\AES_ENC/us23/n1073 ) );
NOR2_X2 \AES_ENC/us23/U325  ( .A1(\AES_ENC/sa23 [1]), .A2(\AES_ENC/us23/n1025 ), .ZN(\AES_ENC/us23/n1054 ) );
NOR2_X2 \AES_ENC/us23/U324  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/us23/n931 ), .ZN(\AES_ENC/us23/n1029 ) );
NOR2_X2 \AES_ENC/us23/U319  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n1056 ) );
NOR2_X2 \AES_ENC/us23/U318  ( .A1(\AES_ENC/us23/n585 ), .A2(\AES_ENC/us23/n596 ), .ZN(\AES_ENC/us23/n1050 ) );
NOR2_X2 \AES_ENC/us23/U317  ( .A1(\AES_ENC/us23/n1121 ), .A2(\AES_ENC/us23/n1025 ), .ZN(\AES_ENC/us23/n1120 ) );
NOR2_X2 \AES_ENC/us23/U316  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/us23/n572 ), .ZN(\AES_ENC/us23/n1074 ) );
NOR2_X2 \AES_ENC/us23/U315  ( .A1(\AES_ENC/us23/n1058 ), .A2(\AES_ENC/us23/n1054 ), .ZN(\AES_ENC/us23/n878 ) );
NOR2_X2 \AES_ENC/us23/U314  ( .A1(\AES_ENC/us23/n878 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n879 ) );
NOR2_X2 \AES_ENC/us23/U312  ( .A1(\AES_ENC/us23/n880 ), .A2(\AES_ENC/us23/n879 ), .ZN(\AES_ENC/us23/n887 ) );
NOR2_X2 \AES_ENC/us23/U311  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n625 ), .ZN(\AES_ENC/us23/n957 ) );
NOR2_X2 \AES_ENC/us23/U310  ( .A1(\AES_ENC/us23/n958 ), .A2(\AES_ENC/us23/n957 ), .ZN(\AES_ENC/us23/n965 ) );
NOR3_X2 \AES_ENC/us23/U309  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n1091 ), .A3(\AES_ENC/us23/n1022 ), .ZN(\AES_ENC/us23/n720 ) );
NOR3_X2 \AES_ENC/us23/U303  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n1054 ), .A3(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n719 ) );
NOR2_X2 \AES_ENC/us23/U302  ( .A1(\AES_ENC/us23/n720 ), .A2(\AES_ENC/us23/n719 ), .ZN(\AES_ENC/us23/n726 ) );
NOR2_X2 \AES_ENC/us23/U300  ( .A1(\AES_ENC/us23/n585 ), .A2(\AES_ENC/us23/n613 ), .ZN(\AES_ENC/us23/n865 ) );
NOR2_X2 \AES_ENC/us23/U299  ( .A1(\AES_ENC/us23/n1059 ), .A2(\AES_ENC/us23/n1058 ), .ZN(\AES_ENC/us23/n1060 ) );
NOR2_X2 \AES_ENC/us23/U298  ( .A1(\AES_ENC/us23/n1095 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n668 ) );
NOR2_X2 \AES_ENC/us23/U297  ( .A1(\AES_ENC/us23/n826 ), .A2(\AES_ENC/us23/n573 ), .ZN(\AES_ENC/us23/n750 ) );
NOR2_X2 \AES_ENC/us23/U296  ( .A1(\AES_ENC/us23/n750 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n751 ) );
NOR2_X2 \AES_ENC/us23/U295  ( .A1(\AES_ENC/us23/n907 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n908 ) );
NOR2_X2 \AES_ENC/us23/U294  ( .A1(\AES_ENC/us23/n990 ), .A2(\AES_ENC/us23/n926 ), .ZN(\AES_ENC/us23/n780 ) );
NOR2_X2 \AES_ENC/us23/U293  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n606 ), .ZN(\AES_ENC/us23/n838 ) );
NOR2_X2 \AES_ENC/us23/U292  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n621 ), .ZN(\AES_ENC/us23/n837 ) );
NOR2_X2 \AES_ENC/us23/U291  ( .A1(\AES_ENC/us23/n838 ), .A2(\AES_ENC/us23/n837 ), .ZN(\AES_ENC/us23/n845 ) );
NOR2_X2 \AES_ENC/us23/U290  ( .A1(\AES_ENC/us23/n1022 ), .A2(\AES_ENC/us23/n1058 ), .ZN(\AES_ENC/us23/n740 ) );
NOR2_X2 \AES_ENC/us23/U284  ( .A1(\AES_ENC/us23/n740 ), .A2(\AES_ENC/us23/n594 ), .ZN(\AES_ENC/us23/n742 ) );
NOR2_X2 \AES_ENC/us23/U283  ( .A1(\AES_ENC/us23/n1098 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n1099 ) );
NOR2_X2 \AES_ENC/us23/U282  ( .A1(\AES_ENC/us23/n1120 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n993 ) );
NOR2_X2 \AES_ENC/us23/U281  ( .A1(\AES_ENC/us23/n993 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n994 ) );
NOR2_X2 \AES_ENC/us23/U280  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n609 ), .ZN(\AES_ENC/us23/n1026 ) );
NOR2_X2 \AES_ENC/us23/U279  ( .A1(\AES_ENC/us23/n573 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n1027 ) );
NOR2_X2 \AES_ENC/us23/U273  ( .A1(\AES_ENC/us23/n1027 ), .A2(\AES_ENC/us23/n1026 ), .ZN(\AES_ENC/us23/n1028 ) );
NOR2_X2 \AES_ENC/us23/U272  ( .A1(\AES_ENC/us23/n1029 ), .A2(\AES_ENC/us23/n1028 ), .ZN(\AES_ENC/us23/n1034 ) );
NOR4_X2 \AES_ENC/us23/U271  ( .A1(\AES_ENC/us23/n757 ), .A2(\AES_ENC/us23/n756 ), .A3(\AES_ENC/us23/n755 ), .A4(\AES_ENC/us23/n754 ), .ZN(\AES_ENC/us23/n758 ) );
NOR2_X2 \AES_ENC/us23/U270  ( .A1(\AES_ENC/us23/n752 ), .A2(\AES_ENC/us23/n751 ), .ZN(\AES_ENC/us23/n759 ) );
NOR2_X2 \AES_ENC/us23/U269  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n1071 ), .ZN(\AES_ENC/us23/n669 ) );
NOR2_X2 \AES_ENC/us23/U268  ( .A1(\AES_ENC/us23/n1056 ), .A2(\AES_ENC/us23/n990 ), .ZN(\AES_ENC/us23/n991 ) );
NOR2_X2 \AES_ENC/us23/U267  ( .A1(\AES_ENC/us23/n991 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n995 ) );
NOR2_X2 \AES_ENC/us23/U263  ( .A1(\AES_ENC/us23/n588 ), .A2(\AES_ENC/us23/n598 ), .ZN(\AES_ENC/us23/n1008 ) );
NOR2_X2 \AES_ENC/us23/U262  ( .A1(\AES_ENC/us23/n839 ), .A2(\AES_ENC/us23/n603 ), .ZN(\AES_ENC/us23/n693 ) );
NOR2_X2 \AES_ENC/us23/U258  ( .A1(\AES_ENC/us23/n587 ), .A2(\AES_ENC/us23/n906 ), .ZN(\AES_ENC/us23/n741 ) );
NOR2_X2 \AES_ENC/us23/U255  ( .A1(\AES_ENC/us23/n1054 ), .A2(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n763 ) );
NOR2_X2 \AES_ENC/us23/U254  ( .A1(\AES_ENC/us23/n763 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n769 ) );
NOR2_X2 \AES_ENC/us23/U253  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n618 ), .ZN(\AES_ENC/us23/n1007 ) );
NOR2_X2 \AES_ENC/us23/U252  ( .A1(\AES_ENC/us23/n591 ), .A2(\AES_ENC/us23/n599 ), .ZN(\AES_ENC/us23/n1123 ) );
NOR2_X2 \AES_ENC/us23/U251  ( .A1(\AES_ENC/us23/n591 ), .A2(\AES_ENC/us23/n598 ), .ZN(\AES_ENC/us23/n710 ) );
INV_X4 \AES_ENC/us23/U250  ( .A(\AES_ENC/us23/n1029 ), .ZN(\AES_ENC/us23/n603 ) );
NOR2_X2 \AES_ENC/us23/U243  ( .A1(\AES_ENC/us23/n594 ), .A2(\AES_ENC/us23/n607 ), .ZN(\AES_ENC/us23/n883 ) );
NOR2_X2 \AES_ENC/us23/U242  ( .A1(\AES_ENC/us23/n623 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n1125 ) );
NOR2_X2 \AES_ENC/us23/U241  ( .A1(\AES_ENC/us23/n911 ), .A2(\AES_ENC/us23/n910 ), .ZN(\AES_ENC/us23/n912 ) );
NOR2_X2 \AES_ENC/us23/U240  ( .A1(\AES_ENC/us23/n912 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n916 ) );
NOR2_X2 \AES_ENC/us23/U239  ( .A1(\AES_ENC/us23/n990 ), .A2(\AES_ENC/us23/n929 ), .ZN(\AES_ENC/us23/n892 ) );
NOR2_X2 \AES_ENC/us23/U238  ( .A1(\AES_ENC/us23/n892 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n893 ) );
NOR2_X2 \AES_ENC/us23/U237  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n621 ), .ZN(\AES_ENC/us23/n950 ) );
NOR2_X2 \AES_ENC/us23/U236  ( .A1(\AES_ENC/us23/n1079 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n1082 ) );
NOR2_X2 \AES_ENC/us23/U235  ( .A1(\AES_ENC/us23/n910 ), .A2(\AES_ENC/us23/n1056 ), .ZN(\AES_ENC/us23/n941 ) );
NOR2_X2 \AES_ENC/us23/U234  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n1077 ), .ZN(\AES_ENC/us23/n841 ) );
NOR2_X2 \AES_ENC/us23/U229  ( .A1(\AES_ENC/us23/n601 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n630 ) );
NOR2_X2 \AES_ENC/us23/U228  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n621 ), .ZN(\AES_ENC/us23/n806 ) );
NOR2_X2 \AES_ENC/us23/U227  ( .A1(\AES_ENC/us23/n601 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n948 ) );
NOR2_X2 \AES_ENC/us23/U226  ( .A1(\AES_ENC/us23/n587 ), .A2(\AES_ENC/us23/n620 ), .ZN(\AES_ENC/us23/n997 ) );
NOR2_X2 \AES_ENC/us23/U225  ( .A1(\AES_ENC/us23/n1121 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n1122 ) );
NOR2_X2 \AES_ENC/us23/U223  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n1023 ), .ZN(\AES_ENC/us23/n756 ) );
NOR2_X2 \AES_ENC/us23/U222  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n621 ), .ZN(\AES_ENC/us23/n870 ) );
NOR2_X2 \AES_ENC/us23/U221  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n569 ), .ZN(\AES_ENC/us23/n947 ) );
NOR2_X2 \AES_ENC/us23/U217  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n1077 ), .ZN(\AES_ENC/us23/n1084 ) );
NOR2_X2 \AES_ENC/us23/U213  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n855 ), .ZN(\AES_ENC/us23/n709 ) );
NOR2_X2 \AES_ENC/us23/U212  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n620 ), .ZN(\AES_ENC/us23/n868 ) );
NOR2_X2 \AES_ENC/us23/U211  ( .A1(\AES_ENC/us23/n1120 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n1124 ) );
NOR2_X2 \AES_ENC/us23/U210  ( .A1(\AES_ENC/us23/n1120 ), .A2(\AES_ENC/us23/n839 ), .ZN(\AES_ENC/us23/n842 ) );
NOR2_X2 \AES_ENC/us23/U209  ( .A1(\AES_ENC/us23/n1120 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n696 ) );
NOR2_X2 \AES_ENC/us23/U208  ( .A1(\AES_ENC/us23/n1074 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n1076 ) );
NOR2_X2 \AES_ENC/us23/U207  ( .A1(\AES_ENC/us23/n1074 ), .A2(\AES_ENC/us23/n609 ), .ZN(\AES_ENC/us23/n781 ) );
NOR3_X2 \AES_ENC/us23/U201  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n1056 ), .A3(\AES_ENC/us23/n990 ), .ZN(\AES_ENC/us23/n979 ) );
NOR3_X2 \AES_ENC/us23/U200  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n1058 ), .A3(\AES_ENC/us23/n1059 ), .ZN(\AES_ENC/us23/n854 ) );
NOR2_X2 \AES_ENC/us23/U199  ( .A1(\AES_ENC/us23/n996 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n869 ) );
NOR2_X2 \AES_ENC/us23/U198  ( .A1(\AES_ENC/us23/n1056 ), .A2(\AES_ENC/us23/n1074 ), .ZN(\AES_ENC/us23/n1057 ) );
NOR3_X2 \AES_ENC/us23/U197  ( .A1(\AES_ENC/us23/n588 ), .A2(\AES_ENC/us23/n1120 ), .A3(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n978 ) );
NOR2_X2 \AES_ENC/us23/U196  ( .A1(\AES_ENC/us23/n996 ), .A2(\AES_ENC/us23/n911 ), .ZN(\AES_ENC/us23/n1116 ) );
NOR2_X2 \AES_ENC/us23/U195  ( .A1(\AES_ENC/us23/n1074 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n754 ) );
NOR2_X2 \AES_ENC/us23/U194  ( .A1(\AES_ENC/us23/n926 ), .A2(\AES_ENC/us23/n1103 ), .ZN(\AES_ENC/us23/n977 ) );
NOR2_X2 \AES_ENC/us23/U187  ( .A1(\AES_ENC/us23/n839 ), .A2(\AES_ENC/us23/n824 ), .ZN(\AES_ENC/us23/n1092 ) );
NOR2_X2 \AES_ENC/us23/U186  ( .A1(\AES_ENC/us23/n573 ), .A2(\AES_ENC/us23/n1074 ), .ZN(\AES_ENC/us23/n684 ) );
NOR2_X2 \AES_ENC/us23/U185  ( .A1(\AES_ENC/us23/n826 ), .A2(\AES_ENC/us23/n1059 ), .ZN(\AES_ENC/us23/n907 ) );
NOR3_X2 \AES_ENC/us23/U184  ( .A1(\AES_ENC/us23/n577 ), .A2(\AES_ENC/us23/n1115 ), .A3(\AES_ENC/us23/n600 ), .ZN(\AES_ENC/us23/n831 ) );
NOR3_X2 \AES_ENC/us23/U183  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n1056 ), .A3(\AES_ENC/us23/n990 ), .ZN(\AES_ENC/us23/n896 ) );
NOR3_X2 \AES_ENC/us23/U182  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n573 ), .A3(\AES_ENC/us23/n1013 ), .ZN(\AES_ENC/us23/n670 ) );
NOR3_X2 \AES_ENC/us23/U181  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n1091 ), .A3(\AES_ENC/us23/n1022 ), .ZN(\AES_ENC/us23/n843 ) );
NOR2_X2 \AES_ENC/us23/U180  ( .A1(\AES_ENC/us23/n1029 ), .A2(\AES_ENC/us23/n1095 ), .ZN(\AES_ENC/us23/n735 ) );
NOR2_X2 \AES_ENC/us23/U174  ( .A1(\AES_ENC/us23/n1100 ), .A2(\AES_ENC/us23/n854 ), .ZN(\AES_ENC/us23/n860 ) );
NAND3_X2 \AES_ENC/us23/U173  ( .A1(\AES_ENC/us23/n569 ), .A2(\AES_ENC/us23/n603 ), .A3(\AES_ENC/us23/n681 ), .ZN(\AES_ENC/us23/n691 ) );
NOR2_X2 \AES_ENC/us23/U172  ( .A1(\AES_ENC/us23/n683 ), .A2(\AES_ENC/us23/n682 ), .ZN(\AES_ENC/us23/n690 ) );
NOR3_X2 \AES_ENC/us23/U171  ( .A1(\AES_ENC/us23/n695 ), .A2(\AES_ENC/us23/n694 ), .A3(\AES_ENC/us23/n693 ), .ZN(\AES_ENC/us23/n700 ) );
NOR4_X2 \AES_ENC/us23/U170  ( .A1(\AES_ENC/us23/n983 ), .A2(\AES_ENC/us23/n698 ), .A3(\AES_ENC/us23/n697 ), .A4(\AES_ENC/us23/n696 ), .ZN(\AES_ENC/us23/n699 ) );
NOR2_X2 \AES_ENC/us23/U169  ( .A1(\AES_ENC/us23/n946 ), .A2(\AES_ENC/us23/n945 ), .ZN(\AES_ENC/us23/n952 ) );
NOR4_X2 \AES_ENC/us23/U168  ( .A1(\AES_ENC/us23/n950 ), .A2(\AES_ENC/us23/n949 ), .A3(\AES_ENC/us23/n948 ), .A4(\AES_ENC/us23/n947 ), .ZN(\AES_ENC/us23/n951 ) );
NOR4_X2 \AES_ENC/us23/U162  ( .A1(\AES_ENC/us23/n896 ), .A2(\AES_ENC/us23/n895 ), .A3(\AES_ENC/us23/n894 ), .A4(\AES_ENC/us23/n893 ), .ZN(\AES_ENC/us23/n897 ) );
NOR2_X2 \AES_ENC/us23/U161  ( .A1(\AES_ENC/us23/n866 ), .A2(\AES_ENC/us23/n865 ), .ZN(\AES_ENC/us23/n872 ) );
NOR4_X2 \AES_ENC/us23/U160  ( .A1(\AES_ENC/us23/n870 ), .A2(\AES_ENC/us23/n869 ), .A3(\AES_ENC/us23/n868 ), .A4(\AES_ENC/us23/n867 ), .ZN(\AES_ENC/us23/n871 ) );
NOR4_X2 \AES_ENC/us23/U159  ( .A1(\AES_ENC/us23/n983 ), .A2(\AES_ENC/us23/n982 ), .A3(\AES_ENC/us23/n981 ), .A4(\AES_ENC/us23/n980 ), .ZN(\AES_ENC/us23/n984 ) );
NOR2_X2 \AES_ENC/us23/U158  ( .A1(\AES_ENC/us23/n979 ), .A2(\AES_ENC/us23/n978 ), .ZN(\AES_ENC/us23/n985 ) );
NOR4_X2 \AES_ENC/us23/U157  ( .A1(\AES_ENC/us23/n1125 ), .A2(\AES_ENC/us23/n1124 ), .A3(\AES_ENC/us23/n1123 ), .A4(\AES_ENC/us23/n1122 ), .ZN(\AES_ENC/us23/n1126 ) );
NOR4_X2 \AES_ENC/us23/U156  ( .A1(\AES_ENC/us23/n1084 ), .A2(\AES_ENC/us23/n1083 ), .A3(\AES_ENC/us23/n1082 ), .A4(\AES_ENC/us23/n1081 ), .ZN(\AES_ENC/us23/n1085 ) );
NOR2_X2 \AES_ENC/us23/U155  ( .A1(\AES_ENC/us23/n1076 ), .A2(\AES_ENC/us23/n1075 ), .ZN(\AES_ENC/us23/n1086 ) );
NOR3_X2 \AES_ENC/us23/U154  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n1054 ), .A3(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n961 ) );
NOR3_X2 \AES_ENC/us23/U153  ( .A1(\AES_ENC/us23/n609 ), .A2(\AES_ENC/us23/n1074 ), .A3(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n671 ) );
NOR2_X2 \AES_ENC/us23/U152  ( .A1(\AES_ENC/us23/n1057 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n1062 ) );
NOR2_X2 \AES_ENC/us23/U143  ( .A1(\AES_ENC/us23/n1055 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n1063 ) );
NOR2_X2 \AES_ENC/us23/U142  ( .A1(\AES_ENC/us23/n1060 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n1061 ) );
NOR4_X2 \AES_ENC/us23/U141  ( .A1(\AES_ENC/us23/n1064 ), .A2(\AES_ENC/us23/n1063 ), .A3(\AES_ENC/us23/n1062 ), .A4(\AES_ENC/us23/n1061 ), .ZN(\AES_ENC/us23/n1065 ) );
NOR3_X2 \AES_ENC/us23/U140  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n1120 ), .A3(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n918 ) );
NOR3_X2 \AES_ENC/us23/U132  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n573 ), .A3(\AES_ENC/us23/n1013 ), .ZN(\AES_ENC/us23/n917 ) );
NOR2_X2 \AES_ENC/us23/U131  ( .A1(\AES_ENC/us23/n914 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n915 ) );
NOR4_X2 \AES_ENC/us23/U130  ( .A1(\AES_ENC/us23/n918 ), .A2(\AES_ENC/us23/n917 ), .A3(\AES_ENC/us23/n916 ), .A4(\AES_ENC/us23/n915 ), .ZN(\AES_ENC/us23/n919 ) );
NOR2_X2 \AES_ENC/us23/U129  ( .A1(\AES_ENC/us23/n594 ), .A2(\AES_ENC/us23/n599 ), .ZN(\AES_ENC/us23/n771 ) );
NOR2_X2 \AES_ENC/us23/U128  ( .A1(\AES_ENC/us23/n1103 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n772 ) );
NOR2_X2 \AES_ENC/us23/U127  ( .A1(\AES_ENC/us23/n592 ), .A2(\AES_ENC/us23/n615 ), .ZN(\AES_ENC/us23/n773 ) );
NOR4_X2 \AES_ENC/us23/U126  ( .A1(\AES_ENC/us23/n773 ), .A2(\AES_ENC/us23/n772 ), .A3(\AES_ENC/us23/n771 ), .A4(\AES_ENC/us23/n770 ), .ZN(\AES_ENC/us23/n774 ) );
NOR2_X2 \AES_ENC/us23/U121  ( .A1(\AES_ENC/us23/n735 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n687 ) );
NOR2_X2 \AES_ENC/us23/U120  ( .A1(\AES_ENC/us23/n684 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n688 ) );
NOR2_X2 \AES_ENC/us23/U119  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n622 ), .ZN(\AES_ENC/us23/n686 ) );
NOR4_X2 \AES_ENC/us23/U118  ( .A1(\AES_ENC/us23/n688 ), .A2(\AES_ENC/us23/n687 ), .A3(\AES_ENC/us23/n686 ), .A4(\AES_ENC/us23/n685 ), .ZN(\AES_ENC/us23/n689 ) );
NOR2_X2 \AES_ENC/us23/U117  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n608 ), .ZN(\AES_ENC/us23/n858 ) );
NOR2_X2 \AES_ENC/us23/U116  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n855 ), .ZN(\AES_ENC/us23/n857 ) );
NOR2_X2 \AES_ENC/us23/U115  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n617 ), .ZN(\AES_ENC/us23/n856 ) );
NOR4_X2 \AES_ENC/us23/U106  ( .A1(\AES_ENC/us23/n858 ), .A2(\AES_ENC/us23/n857 ), .A3(\AES_ENC/us23/n856 ), .A4(\AES_ENC/us23/n958 ), .ZN(\AES_ENC/us23/n859 ) );
NOR2_X2 \AES_ENC/us23/U105  ( .A1(\AES_ENC/us23/n780 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n784 ) );
NOR2_X2 \AES_ENC/us23/U104  ( .A1(\AES_ENC/us23/n1117 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n782 ) );
NOR2_X2 \AES_ENC/us23/U103  ( .A1(\AES_ENC/us23/n781 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n783 ) );
NOR4_X2 \AES_ENC/us23/U102  ( .A1(\AES_ENC/us23/n880 ), .A2(\AES_ENC/us23/n784 ), .A3(\AES_ENC/us23/n783 ), .A4(\AES_ENC/us23/n782 ), .ZN(\AES_ENC/us23/n785 ) );
NOR2_X2 \AES_ENC/us23/U101  ( .A1(\AES_ENC/us23/n597 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n814 ) );
NOR2_X2 \AES_ENC/us23/U100  ( .A1(\AES_ENC/us23/n907 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n813 ) );
NOR3_X2 \AES_ENC/us23/U95  ( .A1(\AES_ENC/us23/n587 ), .A2(\AES_ENC/us23/n1058 ), .A3(\AES_ENC/us23/n1059 ), .ZN(\AES_ENC/us23/n815 ) );
NOR4_X2 \AES_ENC/us23/U94  ( .A1(\AES_ENC/us23/n815 ), .A2(\AES_ENC/us23/n814 ), .A3(\AES_ENC/us23/n813 ), .A4(\AES_ENC/us23/n812 ), .ZN(\AES_ENC/us23/n816 ) );
NOR2_X2 \AES_ENC/us23/U93  ( .A1(\AES_ENC/us23/n575 ), .A2(\AES_ENC/us23/n569 ), .ZN(\AES_ENC/us23/n721 ) );
NOR2_X2 \AES_ENC/us23/U92  ( .A1(\AES_ENC/us23/n1031 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n723 ) );
NOR2_X2 \AES_ENC/us23/U91  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n1096 ), .ZN(\AES_ENC/us23/n722 ) );
NOR4_X2 \AES_ENC/us23/U90  ( .A1(\AES_ENC/us23/n724 ), .A2(\AES_ENC/us23/n723 ), .A3(\AES_ENC/us23/n722 ), .A4(\AES_ENC/us23/n721 ), .ZN(\AES_ENC/us23/n725 ) );
NOR2_X2 \AES_ENC/us23/U89  ( .A1(\AES_ENC/us23/n911 ), .A2(\AES_ENC/us23/n990 ), .ZN(\AES_ENC/us23/n1009 ) );
NOR2_X2 \AES_ENC/us23/U88  ( .A1(\AES_ENC/us23/n1013 ), .A2(\AES_ENC/us23/n573 ), .ZN(\AES_ENC/us23/n1014 ) );
NOR2_X2 \AES_ENC/us23/U87  ( .A1(\AES_ENC/us23/n1014 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n1015 ) );
NOR4_X2 \AES_ENC/us23/U86  ( .A1(\AES_ENC/us23/n1016 ), .A2(\AES_ENC/us23/n1015 ), .A3(\AES_ENC/us23/n1119 ), .A4(\AES_ENC/us23/n1046 ), .ZN(\AES_ENC/us23/n1017 ) );
NOR2_X2 \AES_ENC/us23/U81  ( .A1(\AES_ENC/us23/n996 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n998 ) );
NOR2_X2 \AES_ENC/us23/U80  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n618 ), .ZN(\AES_ENC/us23/n1000 ) );
NOR2_X2 \AES_ENC/us23/U79  ( .A1(\AES_ENC/us23/n594 ), .A2(\AES_ENC/us23/n1096 ), .ZN(\AES_ENC/us23/n999 ) );
NOR4_X2 \AES_ENC/us23/U78  ( .A1(\AES_ENC/us23/n1000 ), .A2(\AES_ENC/us23/n999 ), .A3(\AES_ENC/us23/n998 ), .A4(\AES_ENC/us23/n997 ), .ZN(\AES_ENC/us23/n1001 ) );
NOR2_X2 \AES_ENC/us23/U74  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n1096 ), .ZN(\AES_ENC/us23/n697 ) );
NOR2_X2 \AES_ENC/us23/U73  ( .A1(\AES_ENC/us23/n609 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n958 ) );
NOR2_X2 \AES_ENC/us23/U72  ( .A1(\AES_ENC/us23/n911 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n983 ) );
NOR2_X2 \AES_ENC/us23/U71  ( .A1(\AES_ENC/us23/n1054 ), .A2(\AES_ENC/us23/n1103 ), .ZN(\AES_ENC/us23/n1031 ) );
INV_X4 \AES_ENC/us23/U65  ( .A(\AES_ENC/us23/n1050 ), .ZN(\AES_ENC/us23/n582 ) );
INV_X4 \AES_ENC/us23/U64  ( .A(\AES_ENC/us23/n1072 ), .ZN(\AES_ENC/us23/n586 ) );
INV_X4 \AES_ENC/us23/U63  ( .A(\AES_ENC/us23/n1073 ), .ZN(\AES_ENC/us23/n576 ) );
NOR2_X2 \AES_ENC/us23/U62  ( .A1(\AES_ENC/us23/n603 ), .A2(\AES_ENC/us23/n584 ), .ZN(\AES_ENC/us23/n880 ) );
NOR3_X2 \AES_ENC/us23/U61  ( .A1(\AES_ENC/us23/n826 ), .A2(\AES_ENC/us23/n1121 ), .A3(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n946 ) );
INV_X4 \AES_ENC/us23/U59  ( .A(\AES_ENC/us23/n1010 ), .ZN(\AES_ENC/us23/n579 ) );
NOR3_X2 \AES_ENC/us23/U58  ( .A1(\AES_ENC/us23/n573 ), .A2(\AES_ENC/us23/n1029 ), .A3(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n1119 ) );
INV_X4 \AES_ENC/us23/U57  ( .A(\AES_ENC/us23/n956 ), .ZN(\AES_ENC/us23/n580 ) );
NOR2_X2 \AES_ENC/us23/U50  ( .A1(\AES_ENC/us23/n601 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n1013 ) );
NOR2_X2 \AES_ENC/us23/U49  ( .A1(\AES_ENC/us23/n609 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n910 ) );
NOR2_X2 \AES_ENC/us23/U48  ( .A1(\AES_ENC/us23/n569 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n1091 ) );
NOR2_X2 \AES_ENC/us23/U47  ( .A1(\AES_ENC/us23/n614 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n990 ) );
NOR2_X2 \AES_ENC/us23/U46  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/us23/n1121 ), .ZN(\AES_ENC/us23/n996 ) );
NOR2_X2 \AES_ENC/us23/U45  ( .A1(\AES_ENC/us23/n592 ), .A2(\AES_ENC/us23/n622 ), .ZN(\AES_ENC/us23/n628 ) );
NOR2_X2 \AES_ENC/us23/U44  ( .A1(\AES_ENC/us23/n602 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n866 ) );
NOR2_X2 \AES_ENC/us23/U43  ( .A1(\AES_ENC/us23/n610 ), .A2(\AES_ENC/us23/n592 ), .ZN(\AES_ENC/us23/n1006 ) );
NOR2_X2 \AES_ENC/us23/U42  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n1117 ), .ZN(\AES_ENC/us23/n1118 ) );
NOR2_X2 \AES_ENC/us23/U41  ( .A1(\AES_ENC/us23/n1119 ), .A2(\AES_ENC/us23/n1118 ), .ZN(\AES_ENC/us23/n1127 ) );
NOR2_X2 \AES_ENC/us23/U36  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n616 ), .ZN(\AES_ENC/us23/n629 ) );
NOR2_X2 \AES_ENC/us23/U35  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n906 ), .ZN(\AES_ENC/us23/n909 ) );
NOR2_X2 \AES_ENC/us23/U34  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n607 ), .ZN(\AES_ENC/us23/n658 ) );
NOR2_X2 \AES_ENC/us23/U33  ( .A1(\AES_ENC/us23/n1116 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n695 ) );
NOR2_X2 \AES_ENC/us23/U32  ( .A1(\AES_ENC/us23/n1078 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n1083 ) );
NOR2_X2 \AES_ENC/us23/U31  ( .A1(\AES_ENC/us23/n941 ), .A2(\AES_ENC/us23/n579 ), .ZN(\AES_ENC/us23/n724 ) );
NOR2_X2 \AES_ENC/us23/U30  ( .A1(\AES_ENC/us23/n611 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n1107 ) );
NOR2_X2 \AES_ENC/us23/U29  ( .A1(\AES_ENC/us23/n602 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n840 ) );
NOR2_X2 \AES_ENC/us23/U24  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n623 ), .ZN(\AES_ENC/us23/n633 ) );
NOR2_X2 \AES_ENC/us23/U23  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n1080 ), .ZN(\AES_ENC/us23/n1081 ) );
NOR2_X2 \AES_ENC/us23/U21  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n1045 ), .ZN(\AES_ENC/us23/n812 ) );
NOR2_X2 \AES_ENC/us23/U20  ( .A1(\AES_ENC/us23/n1009 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n960 ) );
NOR2_X2 \AES_ENC/us23/U19  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n619 ), .ZN(\AES_ENC/us23/n982 ) );
NOR2_X2 \AES_ENC/us23/U18  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n616 ), .ZN(\AES_ENC/us23/n757 ) );
NOR2_X2 \AES_ENC/us23/U17  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n598 ), .ZN(\AES_ENC/us23/n698 ) );
NOR2_X2 \AES_ENC/us23/U16  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n605 ), .ZN(\AES_ENC/us23/n708 ) );
NOR2_X2 \AES_ENC/us23/U15  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n603 ), .ZN(\AES_ENC/us23/n770 ) );
NOR2_X2 \AES_ENC/us23/U10  ( .A1(\AES_ENC/us23/n605 ), .A2(\AES_ENC/us23/n576 ), .ZN(\AES_ENC/us23/n803 ) );
NOR2_X2 \AES_ENC/us23/U9  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n881 ), .ZN(\AES_ENC/us23/n711 ) );
NOR2_X2 \AES_ENC/us23/U8  ( .A1(\AES_ENC/us23/n580 ), .A2(\AES_ENC/us23/n603 ), .ZN(\AES_ENC/us23/n867 ) );
NOR2_X2 \AES_ENC/us23/U7  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n615 ), .ZN(\AES_ENC/us23/n804 ) );
NOR2_X2 \AES_ENC/us23/U6  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n609 ), .ZN(\AES_ENC/us23/n1046 ) );
OR2_X4 \AES_ENC/us23/U5  ( .A1(\AES_ENC/us23/n612 ), .A2(\AES_ENC/sa23 [1]),.ZN(\AES_ENC/us23/n570 ) );
OR2_X4 \AES_ENC/us23/U4  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/sa23 [4]),.ZN(\AES_ENC/us23/n569 ) );
NAND2_X2 \AES_ENC/us23/U514  ( .A1(\AES_ENC/us23/n1121 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n1030 ) );
AND2_X2 \AES_ENC/us23/U513  ( .A1(\AES_ENC/us23/n607 ), .A2(\AES_ENC/us23/n1030 ), .ZN(\AES_ENC/us23/n1049 ) );
NAND2_X2 \AES_ENC/us23/U511  ( .A1(\AES_ENC/us23/n1049 ), .A2(\AES_ENC/us23/n794 ), .ZN(\AES_ENC/us23/n637 ) );
AND2_X2 \AES_ENC/us23/U493  ( .A1(\AES_ENC/us23/n779 ), .A2(\AES_ENC/us23/n996 ), .ZN(\AES_ENC/us23/n632 ) );
NAND4_X2 \AES_ENC/us23/U485  ( .A1(\AES_ENC/us23/n637 ), .A2(\AES_ENC/us23/n636 ), .A3(\AES_ENC/us23/n635 ), .A4(\AES_ENC/us23/n634 ), .ZN(\AES_ENC/us23/n638 ) );
NAND2_X2 \AES_ENC/us23/U484  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n638 ), .ZN(\AES_ENC/us23/n679 ) );
NAND2_X2 \AES_ENC/us23/U481  ( .A1(\AES_ENC/us23/n1094 ), .A2(\AES_ENC/us23/n613 ), .ZN(\AES_ENC/us23/n648 ) );
NAND2_X2 \AES_ENC/us23/U476  ( .A1(\AES_ENC/us23/n619 ), .A2(\AES_ENC/us23/n598 ), .ZN(\AES_ENC/us23/n762 ) );
NAND2_X2 \AES_ENC/us23/U475  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n762 ), .ZN(\AES_ENC/us23/n647 ) );
NAND4_X2 \AES_ENC/us23/U457  ( .A1(\AES_ENC/us23/n648 ), .A2(\AES_ENC/us23/n647 ), .A3(\AES_ENC/us23/n646 ), .A4(\AES_ENC/us23/n645 ), .ZN(\AES_ENC/us23/n649 ) );
NAND2_X2 \AES_ENC/us23/U456  ( .A1(\AES_ENC/sa23 [0]), .A2(\AES_ENC/us23/n649 ), .ZN(\AES_ENC/us23/n665 ) );
NAND2_X2 \AES_ENC/us23/U454  ( .A1(\AES_ENC/us23/n626 ), .A2(\AES_ENC/us23/n601 ), .ZN(\AES_ENC/us23/n855 ) );
NAND2_X2 \AES_ENC/us23/U453  ( .A1(\AES_ENC/us23/n617 ), .A2(\AES_ENC/us23/n855 ), .ZN(\AES_ENC/us23/n821 ) );
NAND2_X2 \AES_ENC/us23/U452  ( .A1(\AES_ENC/us23/n1093 ), .A2(\AES_ENC/us23/n821 ), .ZN(\AES_ENC/us23/n662 ) );
NAND2_X2 \AES_ENC/us23/U451  ( .A1(\AES_ENC/us23/n605 ), .A2(\AES_ENC/us23/n620 ), .ZN(\AES_ENC/us23/n650 ) );
NAND2_X2 \AES_ENC/us23/U450  ( .A1(\AES_ENC/us23/n956 ), .A2(\AES_ENC/us23/n650 ), .ZN(\AES_ENC/us23/n661 ) );
NAND2_X2 \AES_ENC/us23/U449  ( .A1(\AES_ENC/us23/n596 ), .A2(\AES_ENC/us23/n581 ), .ZN(\AES_ENC/us23/n839 ) );
OR2_X2 \AES_ENC/us23/U446  ( .A1(\AES_ENC/us23/n839 ), .A2(\AES_ENC/us23/n932 ), .ZN(\AES_ENC/us23/n656 ) );
NAND2_X2 \AES_ENC/us23/U445  ( .A1(\AES_ENC/us23/n624 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n1096 ) );
NAND2_X2 \AES_ENC/us23/U444  ( .A1(\AES_ENC/us23/n1030 ), .A2(\AES_ENC/us23/n1096 ), .ZN(\AES_ENC/us23/n651 ) );
NAND2_X2 \AES_ENC/us23/U443  ( .A1(\AES_ENC/us23/n1114 ), .A2(\AES_ENC/us23/n651 ), .ZN(\AES_ENC/us23/n655 ) );
OR3_X2 \AES_ENC/us23/U440  ( .A1(\AES_ENC/us23/n1079 ), .A2(\AES_ENC/sa23 [7]), .A3(\AES_ENC/us23/n596 ), .ZN(\AES_ENC/us23/n654 ));
NAND2_X2 \AES_ENC/us23/U439  ( .A1(\AES_ENC/us23/n623 ), .A2(\AES_ENC/us23/n619 ), .ZN(\AES_ENC/us23/n652 ) );
NAND4_X2 \AES_ENC/us23/U437  ( .A1(\AES_ENC/us23/n656 ), .A2(\AES_ENC/us23/n655 ), .A3(\AES_ENC/us23/n654 ), .A4(\AES_ENC/us23/n653 ), .ZN(\AES_ENC/us23/n657 ) );
NAND2_X2 \AES_ENC/us23/U436  ( .A1(\AES_ENC/sa23 [2]), .A2(\AES_ENC/us23/n657 ), .ZN(\AES_ENC/us23/n660 ) );
NAND4_X2 \AES_ENC/us23/U432  ( .A1(\AES_ENC/us23/n662 ), .A2(\AES_ENC/us23/n661 ), .A3(\AES_ENC/us23/n660 ), .A4(\AES_ENC/us23/n659 ), .ZN(\AES_ENC/us23/n663 ) );
NAND2_X2 \AES_ENC/us23/U431  ( .A1(\AES_ENC/us23/n663 ), .A2(\AES_ENC/us23/n627 ), .ZN(\AES_ENC/us23/n664 ) );
NAND2_X2 \AES_ENC/us23/U430  ( .A1(\AES_ENC/us23/n665 ), .A2(\AES_ENC/us23/n664 ), .ZN(\AES_ENC/us23/n666 ) );
NAND2_X2 \AES_ENC/us23/U429  ( .A1(\AES_ENC/sa23 [6]), .A2(\AES_ENC/us23/n666 ), .ZN(\AES_ENC/us23/n678 ) );
NAND2_X2 \AES_ENC/us23/U426  ( .A1(\AES_ENC/us23/n735 ), .A2(\AES_ENC/us23/n1093 ), .ZN(\AES_ENC/us23/n675 ) );
NAND2_X2 \AES_ENC/us23/U425  ( .A1(\AES_ENC/us23/n625 ), .A2(\AES_ENC/us23/n607 ), .ZN(\AES_ENC/us23/n1045 ) );
OR2_X2 \AES_ENC/us23/U424  ( .A1(\AES_ENC/us23/n1045 ), .A2(\AES_ENC/us23/n586 ), .ZN(\AES_ENC/us23/n674 ) );
NAND2_X2 \AES_ENC/us23/U423  ( .A1(\AES_ENC/sa23 [1]), .A2(\AES_ENC/us23/n609 ), .ZN(\AES_ENC/us23/n667 ) );
NAND2_X2 \AES_ENC/us23/U422  ( .A1(\AES_ENC/us23/n605 ), .A2(\AES_ENC/us23/n667 ), .ZN(\AES_ENC/us23/n1071 ) );
NAND4_X2 \AES_ENC/us23/U412  ( .A1(\AES_ENC/us23/n675 ), .A2(\AES_ENC/us23/n674 ), .A3(\AES_ENC/us23/n673 ), .A4(\AES_ENC/us23/n672 ), .ZN(\AES_ENC/us23/n676 ) );
NAND2_X2 \AES_ENC/us23/U411  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n676 ), .ZN(\AES_ENC/us23/n677 ) );
NAND2_X2 \AES_ENC/us23/U408  ( .A1(\AES_ENC/us23/n800 ), .A2(\AES_ENC/us23/n1022 ), .ZN(\AES_ENC/us23/n680 ) );
NAND2_X2 \AES_ENC/us23/U407  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n680 ), .ZN(\AES_ENC/us23/n681 ) );
AND2_X2 \AES_ENC/us23/U402  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n684 ), .ZN(\AES_ENC/us23/n682 ) );
NAND4_X2 \AES_ENC/us23/U395  ( .A1(\AES_ENC/us23/n691 ), .A2(\AES_ENC/us23/n583 ), .A3(\AES_ENC/us23/n690 ), .A4(\AES_ENC/us23/n689 ), .ZN(\AES_ENC/us23/n692 ) );
NAND2_X2 \AES_ENC/us23/U394  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n692 ), .ZN(\AES_ENC/us23/n733 ) );
NAND2_X2 \AES_ENC/us23/U392  ( .A1(\AES_ENC/us23/n977 ), .A2(\AES_ENC/us23/n1050 ), .ZN(\AES_ENC/us23/n702 ) );
NAND2_X2 \AES_ENC/us23/U391  ( .A1(\AES_ENC/us23/n1093 ), .A2(\AES_ENC/us23/n1045 ), .ZN(\AES_ENC/us23/n701 ) );
NAND4_X2 \AES_ENC/us23/U381  ( .A1(\AES_ENC/us23/n702 ), .A2(\AES_ENC/us23/n701 ), .A3(\AES_ENC/us23/n700 ), .A4(\AES_ENC/us23/n699 ), .ZN(\AES_ENC/us23/n703 ) );
NAND2_X2 \AES_ENC/us23/U380  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n703 ), .ZN(\AES_ENC/us23/n732 ) );
AND2_X2 \AES_ENC/us23/U379  ( .A1(\AES_ENC/sa23 [0]), .A2(\AES_ENC/sa23 [6]),.ZN(\AES_ENC/us23/n1113 ) );
NAND2_X2 \AES_ENC/us23/U378  ( .A1(\AES_ENC/us23/n619 ), .A2(\AES_ENC/us23/n1030 ), .ZN(\AES_ENC/us23/n881 ) );
NAND2_X2 \AES_ENC/us23/U377  ( .A1(\AES_ENC/us23/n1093 ), .A2(\AES_ENC/us23/n881 ), .ZN(\AES_ENC/us23/n715 ) );
NAND2_X2 \AES_ENC/us23/U376  ( .A1(\AES_ENC/us23/n1010 ), .A2(\AES_ENC/us23/n622 ), .ZN(\AES_ENC/us23/n714 ) );
NAND2_X2 \AES_ENC/us23/U375  ( .A1(\AES_ENC/us23/n855 ), .A2(\AES_ENC/us23/n625 ), .ZN(\AES_ENC/us23/n1117 ) );
XNOR2_X2 \AES_ENC/us23/U371  ( .A(\AES_ENC/us23/n593 ), .B(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n824 ) );
NAND4_X2 \AES_ENC/us23/U362  ( .A1(\AES_ENC/us23/n715 ), .A2(\AES_ENC/us23/n714 ), .A3(\AES_ENC/us23/n713 ), .A4(\AES_ENC/us23/n712 ), .ZN(\AES_ENC/us23/n716 ) );
NAND2_X2 \AES_ENC/us23/U361  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n716 ), .ZN(\AES_ENC/us23/n731 ) );
AND2_X2 \AES_ENC/us23/U360  ( .A1(\AES_ENC/sa23 [6]), .A2(\AES_ENC/us23/n627 ), .ZN(\AES_ENC/us23/n1131 ) );
NAND2_X2 \AES_ENC/us23/U359  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n717 ) );
NAND2_X2 \AES_ENC/us23/U358  ( .A1(\AES_ENC/us23/n1029 ), .A2(\AES_ENC/us23/n717 ), .ZN(\AES_ENC/us23/n728 ) );
NAND2_X2 \AES_ENC/us23/U357  ( .A1(\AES_ENC/sa23 [1]), .A2(\AES_ENC/us23/n612 ), .ZN(\AES_ENC/us23/n1097 ) );
NAND2_X2 \AES_ENC/us23/U356  ( .A1(\AES_ENC/us23/n610 ), .A2(\AES_ENC/us23/n1097 ), .ZN(\AES_ENC/us23/n718 ) );
NAND2_X2 \AES_ENC/us23/U355  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n718 ), .ZN(\AES_ENC/us23/n727 ) );
NAND4_X2 \AES_ENC/us23/U344  ( .A1(\AES_ENC/us23/n728 ), .A2(\AES_ENC/us23/n727 ), .A3(\AES_ENC/us23/n726 ), .A4(\AES_ENC/us23/n725 ), .ZN(\AES_ENC/us23/n729 ) );
NAND2_X2 \AES_ENC/us23/U343  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n729 ), .ZN(\AES_ENC/us23/n730 ) );
NAND4_X2 \AES_ENC/us23/U342  ( .A1(\AES_ENC/us23/n733 ), .A2(\AES_ENC/us23/n732 ), .A3(\AES_ENC/us23/n731 ), .A4(\AES_ENC/us23/n730 ), .ZN(\AES_ENC/sa23_sub[1] ) );
NAND2_X2 \AES_ENC/us23/U341  ( .A1(\AES_ENC/sa23 [7]), .A2(\AES_ENC/us23/n593 ), .ZN(\AES_ENC/us23/n734 ) );
NAND2_X2 \AES_ENC/us23/U340  ( .A1(\AES_ENC/us23/n734 ), .A2(\AES_ENC/us23/n588 ), .ZN(\AES_ENC/us23/n738 ) );
OR4_X2 \AES_ENC/us23/U339  ( .A1(\AES_ENC/us23/n738 ), .A2(\AES_ENC/us23/n596 ), .A3(\AES_ENC/us23/n826 ), .A4(\AES_ENC/us23/n1121 ), .ZN(\AES_ENC/us23/n746 ) );
NAND2_X2 \AES_ENC/us23/U337  ( .A1(\AES_ENC/us23/n1100 ), .A2(\AES_ENC/us23/n617 ), .ZN(\AES_ENC/us23/n992 ) );
OR2_X2 \AES_ENC/us23/U336  ( .A1(\AES_ENC/us23/n592 ), .A2(\AES_ENC/us23/n735 ), .ZN(\AES_ENC/us23/n737 ) );
NAND2_X2 \AES_ENC/us23/U334  ( .A1(\AES_ENC/us23/n605 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n753 ) );
NAND2_X2 \AES_ENC/us23/U333  ( .A1(\AES_ENC/us23/n603 ), .A2(\AES_ENC/us23/n753 ), .ZN(\AES_ENC/us23/n1080 ) );
NAND2_X2 \AES_ENC/us23/U332  ( .A1(\AES_ENC/us23/n1048 ), .A2(\AES_ENC/us23/n602 ), .ZN(\AES_ENC/us23/n736 ) );
NAND2_X2 \AES_ENC/us23/U331  ( .A1(\AES_ENC/us23/n737 ), .A2(\AES_ENC/us23/n736 ), .ZN(\AES_ENC/us23/n739 ) );
NAND2_X2 \AES_ENC/us23/U330  ( .A1(\AES_ENC/us23/n739 ), .A2(\AES_ENC/us23/n738 ), .ZN(\AES_ENC/us23/n745 ) );
NAND2_X2 \AES_ENC/us23/U326  ( .A1(\AES_ENC/us23/n1096 ), .A2(\AES_ENC/us23/n598 ), .ZN(\AES_ENC/us23/n906 ) );
NAND4_X2 \AES_ENC/us23/U323  ( .A1(\AES_ENC/us23/n746 ), .A2(\AES_ENC/us23/n992 ), .A3(\AES_ENC/us23/n745 ), .A4(\AES_ENC/us23/n744 ), .ZN(\AES_ENC/us23/n747 ) );
NAND2_X2 \AES_ENC/us23/U322  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n747 ), .ZN(\AES_ENC/us23/n793 ) );
NAND2_X2 \AES_ENC/us23/U321  ( .A1(\AES_ENC/us23/n606 ), .A2(\AES_ENC/us23/n855 ), .ZN(\AES_ENC/us23/n748 ) );
NAND2_X2 \AES_ENC/us23/U320  ( .A1(\AES_ENC/us23/n956 ), .A2(\AES_ENC/us23/n748 ), .ZN(\AES_ENC/us23/n760 ) );
NAND2_X2 \AES_ENC/us23/U313  ( .A1(\AES_ENC/us23/n598 ), .A2(\AES_ENC/us23/n753 ), .ZN(\AES_ENC/us23/n1023 ) );
NAND4_X2 \AES_ENC/us23/U308  ( .A1(\AES_ENC/us23/n760 ), .A2(\AES_ENC/us23/n992 ), .A3(\AES_ENC/us23/n759 ), .A4(\AES_ENC/us23/n758 ), .ZN(\AES_ENC/us23/n761 ) );
NAND2_X2 \AES_ENC/us23/U307  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n761 ), .ZN(\AES_ENC/us23/n792 ) );
NAND2_X2 \AES_ENC/us23/U306  ( .A1(\AES_ENC/us23/n606 ), .A2(\AES_ENC/us23/n610 ), .ZN(\AES_ENC/us23/n989 ) );
NAND2_X2 \AES_ENC/us23/U305  ( .A1(\AES_ENC/us23/n1050 ), .A2(\AES_ENC/us23/n989 ), .ZN(\AES_ENC/us23/n777 ) );
NAND2_X2 \AES_ENC/us23/U304  ( .A1(\AES_ENC/us23/n1093 ), .A2(\AES_ENC/us23/n762 ), .ZN(\AES_ENC/us23/n776 ) );
XNOR2_X2 \AES_ENC/us23/U301  ( .A(\AES_ENC/sa23 [7]), .B(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n959 ) );
NAND4_X2 \AES_ENC/us23/U289  ( .A1(\AES_ENC/us23/n777 ), .A2(\AES_ENC/us23/n776 ), .A3(\AES_ENC/us23/n775 ), .A4(\AES_ENC/us23/n774 ), .ZN(\AES_ENC/us23/n778 ) );
NAND2_X2 \AES_ENC/us23/U288  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n778 ), .ZN(\AES_ENC/us23/n791 ) );
NAND2_X2 \AES_ENC/us23/U287  ( .A1(\AES_ENC/us23/n1056 ), .A2(\AES_ENC/us23/n1050 ), .ZN(\AES_ENC/us23/n788 ) );
NAND2_X2 \AES_ENC/us23/U286  ( .A1(\AES_ENC/us23/n1091 ), .A2(\AES_ENC/us23/n779 ), .ZN(\AES_ENC/us23/n787 ) );
NAND2_X2 \AES_ENC/us23/U285  ( .A1(\AES_ENC/us23/n956 ), .A2(\AES_ENC/sa23 [1]), .ZN(\AES_ENC/us23/n786 ) );
NAND4_X2 \AES_ENC/us23/U278  ( .A1(\AES_ENC/us23/n788 ), .A2(\AES_ENC/us23/n787 ), .A3(\AES_ENC/us23/n786 ), .A4(\AES_ENC/us23/n785 ), .ZN(\AES_ENC/us23/n789 ) );
NAND2_X2 \AES_ENC/us23/U277  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n789 ), .ZN(\AES_ENC/us23/n790 ) );
NAND4_X2 \AES_ENC/us23/U276  ( .A1(\AES_ENC/us23/n793 ), .A2(\AES_ENC/us23/n792 ), .A3(\AES_ENC/us23/n791 ), .A4(\AES_ENC/us23/n790 ), .ZN(\AES_ENC/sa23_sub[2] ) );
NAND2_X2 \AES_ENC/us23/U275  ( .A1(\AES_ENC/us23/n1059 ), .A2(\AES_ENC/us23/n794 ), .ZN(\AES_ENC/us23/n810 ) );
NAND2_X2 \AES_ENC/us23/U274  ( .A1(\AES_ENC/us23/n1049 ), .A2(\AES_ENC/us23/n956 ), .ZN(\AES_ENC/us23/n809 ) );
OR2_X2 \AES_ENC/us23/U266  ( .A1(\AES_ENC/us23/n1096 ), .A2(\AES_ENC/us23/n587 ), .ZN(\AES_ENC/us23/n802 ) );
NAND2_X2 \AES_ENC/us23/U265  ( .A1(\AES_ENC/us23/n1053 ), .A2(\AES_ENC/us23/n800 ), .ZN(\AES_ENC/us23/n801 ) );
NAND2_X2 \AES_ENC/us23/U264  ( .A1(\AES_ENC/us23/n802 ), .A2(\AES_ENC/us23/n801 ), .ZN(\AES_ENC/us23/n805 ) );
NAND4_X2 \AES_ENC/us23/U261  ( .A1(\AES_ENC/us23/n810 ), .A2(\AES_ENC/us23/n809 ), .A3(\AES_ENC/us23/n808 ), .A4(\AES_ENC/us23/n807 ), .ZN(\AES_ENC/us23/n811 ) );
NAND2_X2 \AES_ENC/us23/U260  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n811 ), .ZN(\AES_ENC/us23/n852 ) );
OR2_X2 \AES_ENC/us23/U259  ( .A1(\AES_ENC/us23/n1023 ), .A2(\AES_ENC/us23/n575 ), .ZN(\AES_ENC/us23/n819 ) );
OR2_X2 \AES_ENC/us23/U257  ( .A1(\AES_ENC/us23/n570 ), .A2(\AES_ENC/us23/n930 ), .ZN(\AES_ENC/us23/n818 ) );
NAND2_X2 \AES_ENC/us23/U256  ( .A1(\AES_ENC/us23/n1013 ), .A2(\AES_ENC/us23/n1094 ), .ZN(\AES_ENC/us23/n817 ) );
NAND4_X2 \AES_ENC/us23/U249  ( .A1(\AES_ENC/us23/n819 ), .A2(\AES_ENC/us23/n818 ), .A3(\AES_ENC/us23/n817 ), .A4(\AES_ENC/us23/n816 ), .ZN(\AES_ENC/us23/n820 ) );
NAND2_X2 \AES_ENC/us23/U248  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n820 ), .ZN(\AES_ENC/us23/n851 ) );
NAND2_X2 \AES_ENC/us23/U247  ( .A1(\AES_ENC/us23/n956 ), .A2(\AES_ENC/us23/n1080 ), .ZN(\AES_ENC/us23/n835 ) );
NAND2_X2 \AES_ENC/us23/U246  ( .A1(\AES_ENC/us23/n570 ), .A2(\AES_ENC/us23/n1030 ), .ZN(\AES_ENC/us23/n1047 ) );
OR2_X2 \AES_ENC/us23/U245  ( .A1(\AES_ENC/us23/n1047 ), .A2(\AES_ENC/us23/n582 ), .ZN(\AES_ENC/us23/n834 ) );
NAND2_X2 \AES_ENC/us23/U244  ( .A1(\AES_ENC/us23/n1072 ), .A2(\AES_ENC/us23/n620 ), .ZN(\AES_ENC/us23/n833 ) );
NAND4_X2 \AES_ENC/us23/U233  ( .A1(\AES_ENC/us23/n835 ), .A2(\AES_ENC/us23/n834 ), .A3(\AES_ENC/us23/n833 ), .A4(\AES_ENC/us23/n832 ), .ZN(\AES_ENC/us23/n836 ) );
NAND2_X2 \AES_ENC/us23/U232  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n836 ), .ZN(\AES_ENC/us23/n850 ) );
NAND2_X2 \AES_ENC/us23/U231  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n601 ), .ZN(\AES_ENC/us23/n847 ) );
NAND2_X2 \AES_ENC/us23/U230  ( .A1(\AES_ENC/us23/n1050 ), .A2(\AES_ENC/us23/n1071 ), .ZN(\AES_ENC/us23/n846 ) );
OR2_X2 \AES_ENC/us23/U224  ( .A1(\AES_ENC/us23/n1053 ), .A2(\AES_ENC/us23/n911 ), .ZN(\AES_ENC/us23/n1077 ) );
NAND4_X2 \AES_ENC/us23/U220  ( .A1(\AES_ENC/us23/n847 ), .A2(\AES_ENC/us23/n846 ), .A3(\AES_ENC/us23/n845 ), .A4(\AES_ENC/us23/n844 ), .ZN(\AES_ENC/us23/n848 ) );
NAND2_X2 \AES_ENC/us23/U219  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n848 ), .ZN(\AES_ENC/us23/n849 ) );
NAND4_X2 \AES_ENC/us23/U218  ( .A1(\AES_ENC/us23/n852 ), .A2(\AES_ENC/us23/n851 ), .A3(\AES_ENC/us23/n850 ), .A4(\AES_ENC/us23/n849 ), .ZN(\AES_ENC/sa23_sub[3] ) );
NAND2_X2 \AES_ENC/us23/U216  ( .A1(\AES_ENC/us23/n1009 ), .A2(\AES_ENC/us23/n1072 ), .ZN(\AES_ENC/us23/n862 ) );
NAND2_X2 \AES_ENC/us23/U215  ( .A1(\AES_ENC/us23/n610 ), .A2(\AES_ENC/us23/n618 ), .ZN(\AES_ENC/us23/n853 ) );
NAND2_X2 \AES_ENC/us23/U214  ( .A1(\AES_ENC/us23/n1050 ), .A2(\AES_ENC/us23/n853 ), .ZN(\AES_ENC/us23/n861 ) );
NAND4_X2 \AES_ENC/us23/U206  ( .A1(\AES_ENC/us23/n862 ), .A2(\AES_ENC/us23/n861 ), .A3(\AES_ENC/us23/n860 ), .A4(\AES_ENC/us23/n859 ), .ZN(\AES_ENC/us23/n863 ) );
NAND2_X2 \AES_ENC/us23/U205  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n863 ), .ZN(\AES_ENC/us23/n905 ) );
NAND2_X2 \AES_ENC/us23/U204  ( .A1(\AES_ENC/us23/n1010 ), .A2(\AES_ENC/us23/n989 ), .ZN(\AES_ENC/us23/n874 ) );
NAND2_X2 \AES_ENC/us23/U203  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n592 ), .ZN(\AES_ENC/us23/n864 ) );
NAND2_X2 \AES_ENC/us23/U202  ( .A1(\AES_ENC/us23/n929 ), .A2(\AES_ENC/us23/n864 ), .ZN(\AES_ENC/us23/n873 ) );
NAND4_X2 \AES_ENC/us23/U193  ( .A1(\AES_ENC/us23/n874 ), .A2(\AES_ENC/us23/n873 ), .A3(\AES_ENC/us23/n872 ), .A4(\AES_ENC/us23/n871 ), .ZN(\AES_ENC/us23/n875 ) );
NAND2_X2 \AES_ENC/us23/U192  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n875 ), .ZN(\AES_ENC/us23/n904 ) );
NAND2_X2 \AES_ENC/us23/U191  ( .A1(\AES_ENC/us23/n597 ), .A2(\AES_ENC/us23/n1050 ), .ZN(\AES_ENC/us23/n889 ) );
NAND2_X2 \AES_ENC/us23/U190  ( .A1(\AES_ENC/us23/n1093 ), .A2(\AES_ENC/us23/n617 ), .ZN(\AES_ENC/us23/n876 ) );
NAND2_X2 \AES_ENC/us23/U189  ( .A1(\AES_ENC/us23/n576 ), .A2(\AES_ENC/us23/n876 ), .ZN(\AES_ENC/us23/n877 ) );
NAND2_X2 \AES_ENC/us23/U188  ( .A1(\AES_ENC/us23/n877 ), .A2(\AES_ENC/us23/n601 ), .ZN(\AES_ENC/us23/n888 ) );
NAND4_X2 \AES_ENC/us23/U179  ( .A1(\AES_ENC/us23/n889 ), .A2(\AES_ENC/us23/n888 ), .A3(\AES_ENC/us23/n887 ), .A4(\AES_ENC/us23/n886 ), .ZN(\AES_ENC/us23/n890 ) );
NAND2_X2 \AES_ENC/us23/U178  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n890 ), .ZN(\AES_ENC/us23/n903 ) );
OR2_X2 \AES_ENC/us23/U177  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n1059 ), .ZN(\AES_ENC/us23/n900 ) );
NAND2_X2 \AES_ENC/us23/U176  ( .A1(\AES_ENC/us23/n1073 ), .A2(\AES_ENC/us23/n1047 ), .ZN(\AES_ENC/us23/n899 ) );
NAND2_X2 \AES_ENC/us23/U175  ( .A1(\AES_ENC/us23/n1094 ), .A2(\AES_ENC/us23/n608 ), .ZN(\AES_ENC/us23/n898 ) );
NAND4_X2 \AES_ENC/us23/U167  ( .A1(\AES_ENC/us23/n900 ), .A2(\AES_ENC/us23/n899 ), .A3(\AES_ENC/us23/n898 ), .A4(\AES_ENC/us23/n897 ), .ZN(\AES_ENC/us23/n901 ) );
NAND2_X2 \AES_ENC/us23/U166  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n901 ), .ZN(\AES_ENC/us23/n902 ) );
NAND4_X2 \AES_ENC/us23/U165  ( .A1(\AES_ENC/us23/n905 ), .A2(\AES_ENC/us23/n904 ), .A3(\AES_ENC/us23/n903 ), .A4(\AES_ENC/us23/n902 ), .ZN(\AES_ENC/sa23_sub[4] ) );
NAND2_X2 \AES_ENC/us23/U164  ( .A1(\AES_ENC/us23/n1094 ), .A2(\AES_ENC/us23/n615 ), .ZN(\AES_ENC/us23/n922 ) );
NAND2_X2 \AES_ENC/us23/U163  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n989 ), .ZN(\AES_ENC/us23/n921 ) );
NAND4_X2 \AES_ENC/us23/U151  ( .A1(\AES_ENC/us23/n922 ), .A2(\AES_ENC/us23/n921 ), .A3(\AES_ENC/us23/n920 ), .A4(\AES_ENC/us23/n919 ), .ZN(\AES_ENC/us23/n923 ) );
NAND2_X2 \AES_ENC/us23/U150  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n923 ), .ZN(\AES_ENC/us23/n972 ) );
NAND2_X2 \AES_ENC/us23/U149  ( .A1(\AES_ENC/us23/n603 ), .A2(\AES_ENC/us23/n605 ), .ZN(\AES_ENC/us23/n924 ) );
NAND2_X2 \AES_ENC/us23/U148  ( .A1(\AES_ENC/us23/n1073 ), .A2(\AES_ENC/us23/n924 ), .ZN(\AES_ENC/us23/n939 ) );
NAND2_X2 \AES_ENC/us23/U147  ( .A1(\AES_ENC/us23/n926 ), .A2(\AES_ENC/us23/n925 ), .ZN(\AES_ENC/us23/n927 ) );
NAND2_X2 \AES_ENC/us23/U146  ( .A1(\AES_ENC/us23/n587 ), .A2(\AES_ENC/us23/n927 ), .ZN(\AES_ENC/us23/n928 ) );
NAND2_X2 \AES_ENC/us23/U145  ( .A1(\AES_ENC/us23/n928 ), .A2(\AES_ENC/us23/n1080 ), .ZN(\AES_ENC/us23/n938 ) );
OR2_X2 \AES_ENC/us23/U144  ( .A1(\AES_ENC/us23/n1117 ), .A2(\AES_ENC/us23/n580 ), .ZN(\AES_ENC/us23/n937 ) );
NAND4_X2 \AES_ENC/us23/U139  ( .A1(\AES_ENC/us23/n939 ), .A2(\AES_ENC/us23/n938 ), .A3(\AES_ENC/us23/n937 ), .A4(\AES_ENC/us23/n936 ), .ZN(\AES_ENC/us23/n940 ) );
NAND2_X2 \AES_ENC/us23/U138  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n940 ), .ZN(\AES_ENC/us23/n971 ) );
OR2_X2 \AES_ENC/us23/U137  ( .A1(\AES_ENC/us23/n586 ), .A2(\AES_ENC/us23/n941 ), .ZN(\AES_ENC/us23/n954 ) );
NAND2_X2 \AES_ENC/us23/U136  ( .A1(\AES_ENC/us23/n1096 ), .A2(\AES_ENC/us23/n618 ), .ZN(\AES_ENC/us23/n942 ) );
NAND2_X2 \AES_ENC/us23/U135  ( .A1(\AES_ENC/us23/n1048 ), .A2(\AES_ENC/us23/n942 ), .ZN(\AES_ENC/us23/n943 ) );
NAND2_X2 \AES_ENC/us23/U134  ( .A1(\AES_ENC/us23/n582 ), .A2(\AES_ENC/us23/n943 ), .ZN(\AES_ENC/us23/n944 ) );
NAND2_X2 \AES_ENC/us23/U133  ( .A1(\AES_ENC/us23/n944 ), .A2(\AES_ENC/us23/n599 ), .ZN(\AES_ENC/us23/n953 ) );
NAND4_X2 \AES_ENC/us23/U125  ( .A1(\AES_ENC/us23/n954 ), .A2(\AES_ENC/us23/n953 ), .A3(\AES_ENC/us23/n952 ), .A4(\AES_ENC/us23/n951 ), .ZN(\AES_ENC/us23/n955 ) );
NAND2_X2 \AES_ENC/us23/U124  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n955 ), .ZN(\AES_ENC/us23/n970 ) );
NAND2_X2 \AES_ENC/us23/U123  ( .A1(\AES_ENC/us23/n1094 ), .A2(\AES_ENC/us23/n1071 ), .ZN(\AES_ENC/us23/n967 ) );
NAND2_X2 \AES_ENC/us23/U122  ( .A1(\AES_ENC/us23/n956 ), .A2(\AES_ENC/us23/n1030 ), .ZN(\AES_ENC/us23/n966 ) );
NAND4_X2 \AES_ENC/us23/U114  ( .A1(\AES_ENC/us23/n967 ), .A2(\AES_ENC/us23/n966 ), .A3(\AES_ENC/us23/n965 ), .A4(\AES_ENC/us23/n964 ), .ZN(\AES_ENC/us23/n968 ) );
NAND2_X2 \AES_ENC/us23/U113  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n968 ), .ZN(\AES_ENC/us23/n969 ) );
NAND4_X2 \AES_ENC/us23/U112  ( .A1(\AES_ENC/us23/n972 ), .A2(\AES_ENC/us23/n971 ), .A3(\AES_ENC/us23/n970 ), .A4(\AES_ENC/us23/n969 ), .ZN(\AES_ENC/sa23_sub[5] ) );
NAND2_X2 \AES_ENC/us23/U111  ( .A1(\AES_ENC/us23/n570 ), .A2(\AES_ENC/us23/n1097 ), .ZN(\AES_ENC/us23/n973 ) );
NAND2_X2 \AES_ENC/us23/U110  ( .A1(\AES_ENC/us23/n1073 ), .A2(\AES_ENC/us23/n973 ), .ZN(\AES_ENC/us23/n987 ) );
NAND2_X2 \AES_ENC/us23/U109  ( .A1(\AES_ENC/us23/n974 ), .A2(\AES_ENC/us23/n1077 ), .ZN(\AES_ENC/us23/n975 ) );
NAND2_X2 \AES_ENC/us23/U108  ( .A1(\AES_ENC/us23/n584 ), .A2(\AES_ENC/us23/n975 ), .ZN(\AES_ENC/us23/n976 ) );
NAND2_X2 \AES_ENC/us23/U107  ( .A1(\AES_ENC/us23/n977 ), .A2(\AES_ENC/us23/n976 ), .ZN(\AES_ENC/us23/n986 ) );
NAND4_X2 \AES_ENC/us23/U99  ( .A1(\AES_ENC/us23/n987 ), .A2(\AES_ENC/us23/n986 ), .A3(\AES_ENC/us23/n985 ), .A4(\AES_ENC/us23/n984 ), .ZN(\AES_ENC/us23/n988 ) );
NAND2_X2 \AES_ENC/us23/U98  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n988 ), .ZN(\AES_ENC/us23/n1044 ) );
NAND2_X2 \AES_ENC/us23/U97  ( .A1(\AES_ENC/us23/n1073 ), .A2(\AES_ENC/us23/n989 ), .ZN(\AES_ENC/us23/n1004 ) );
NAND2_X2 \AES_ENC/us23/U96  ( .A1(\AES_ENC/us23/n1092 ), .A2(\AES_ENC/us23/n605 ), .ZN(\AES_ENC/us23/n1003 ) );
NAND4_X2 \AES_ENC/us23/U85  ( .A1(\AES_ENC/us23/n1004 ), .A2(\AES_ENC/us23/n1003 ), .A3(\AES_ENC/us23/n1002 ), .A4(\AES_ENC/us23/n1001 ), .ZN(\AES_ENC/us23/n1005 ) );
NAND2_X2 \AES_ENC/us23/U84  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n1005 ), .ZN(\AES_ENC/us23/n1043 ) );
NAND2_X2 \AES_ENC/us23/U83  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n626 ), .ZN(\AES_ENC/us23/n1020 ) );
NAND2_X2 \AES_ENC/us23/U82  ( .A1(\AES_ENC/us23/n1050 ), .A2(\AES_ENC/us23/n612 ), .ZN(\AES_ENC/us23/n1019 ) );
NAND2_X2 \AES_ENC/us23/U77  ( .A1(\AES_ENC/us23/n1059 ), .A2(\AES_ENC/us23/n1114 ), .ZN(\AES_ENC/us23/n1012 ) );
NAND2_X2 \AES_ENC/us23/U76  ( .A1(\AES_ENC/us23/n1010 ), .A2(\AES_ENC/us23/n604 ), .ZN(\AES_ENC/us23/n1011 ) );
NAND2_X2 \AES_ENC/us23/U75  ( .A1(\AES_ENC/us23/n1012 ), .A2(\AES_ENC/us23/n1011 ), .ZN(\AES_ENC/us23/n1016 ) );
NAND4_X2 \AES_ENC/us23/U70  ( .A1(\AES_ENC/us23/n1020 ), .A2(\AES_ENC/us23/n1019 ), .A3(\AES_ENC/us23/n1018 ), .A4(\AES_ENC/us23/n1017 ), .ZN(\AES_ENC/us23/n1021 ) );
NAND2_X2 \AES_ENC/us23/U69  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n1021 ), .ZN(\AES_ENC/us23/n1042 ) );
NAND2_X2 \AES_ENC/us23/U68  ( .A1(\AES_ENC/us23/n1022 ), .A2(\AES_ENC/us23/n1093 ), .ZN(\AES_ENC/us23/n1039 ) );
NAND2_X2 \AES_ENC/us23/U67  ( .A1(\AES_ENC/us23/n1050 ), .A2(\AES_ENC/us23/n1023 ), .ZN(\AES_ENC/us23/n1038 ) );
NAND2_X2 \AES_ENC/us23/U66  ( .A1(\AES_ENC/us23/n1024 ), .A2(\AES_ENC/us23/n1071 ), .ZN(\AES_ENC/us23/n1037 ) );
AND2_X2 \AES_ENC/us23/U60  ( .A1(\AES_ENC/us23/n1030 ), .A2(\AES_ENC/us23/n621 ), .ZN(\AES_ENC/us23/n1078 ) );
NAND4_X2 \AES_ENC/us23/U56  ( .A1(\AES_ENC/us23/n1039 ), .A2(\AES_ENC/us23/n1038 ), .A3(\AES_ENC/us23/n1037 ), .A4(\AES_ENC/us23/n1036 ), .ZN(\AES_ENC/us23/n1040 ) );
NAND2_X2 \AES_ENC/us23/U55  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n1040 ), .ZN(\AES_ENC/us23/n1041 ) );
NAND4_X2 \AES_ENC/us23/U54  ( .A1(\AES_ENC/us23/n1044 ), .A2(\AES_ENC/us23/n1043 ), .A3(\AES_ENC/us23/n1042 ), .A4(\AES_ENC/us23/n1041 ), .ZN(\AES_ENC/sa23_sub[6] ) );
NAND2_X2 \AES_ENC/us23/U53  ( .A1(\AES_ENC/us23/n1072 ), .A2(\AES_ENC/us23/n1045 ), .ZN(\AES_ENC/us23/n1068 ) );
NAND2_X2 \AES_ENC/us23/U52  ( .A1(\AES_ENC/us23/n1046 ), .A2(\AES_ENC/us23/n603 ), .ZN(\AES_ENC/us23/n1067 ) );
NAND2_X2 \AES_ENC/us23/U51  ( .A1(\AES_ENC/us23/n1094 ), .A2(\AES_ENC/us23/n1047 ), .ZN(\AES_ENC/us23/n1066 ) );
NAND4_X2 \AES_ENC/us23/U40  ( .A1(\AES_ENC/us23/n1068 ), .A2(\AES_ENC/us23/n1067 ), .A3(\AES_ENC/us23/n1066 ), .A4(\AES_ENC/us23/n1065 ), .ZN(\AES_ENC/us23/n1069 ) );
NAND2_X2 \AES_ENC/us23/U39  ( .A1(\AES_ENC/us23/n1070 ), .A2(\AES_ENC/us23/n1069 ), .ZN(\AES_ENC/us23/n1135 ) );
NAND2_X2 \AES_ENC/us23/U38  ( .A1(\AES_ENC/us23/n1072 ), .A2(\AES_ENC/us23/n1071 ), .ZN(\AES_ENC/us23/n1088 ) );
NAND2_X2 \AES_ENC/us23/U37  ( .A1(\AES_ENC/us23/n1073 ), .A2(\AES_ENC/us23/n608 ), .ZN(\AES_ENC/us23/n1087 ) );
NAND4_X2 \AES_ENC/us23/U28  ( .A1(\AES_ENC/us23/n1088 ), .A2(\AES_ENC/us23/n1087 ), .A3(\AES_ENC/us23/n1086 ), .A4(\AES_ENC/us23/n1085 ), .ZN(\AES_ENC/us23/n1089 ) );
NAND2_X2 \AES_ENC/us23/U27  ( .A1(\AES_ENC/us23/n1090 ), .A2(\AES_ENC/us23/n1089 ), .ZN(\AES_ENC/us23/n1134 ) );
NAND2_X2 \AES_ENC/us23/U26  ( .A1(\AES_ENC/us23/n1091 ), .A2(\AES_ENC/us23/n1093 ), .ZN(\AES_ENC/us23/n1111 ) );
NAND2_X2 \AES_ENC/us23/U25  ( .A1(\AES_ENC/us23/n1092 ), .A2(\AES_ENC/us23/n1120 ), .ZN(\AES_ENC/us23/n1110 ) );
AND2_X2 \AES_ENC/us23/U22  ( .A1(\AES_ENC/us23/n1097 ), .A2(\AES_ENC/us23/n1096 ), .ZN(\AES_ENC/us23/n1098 ) );
NAND4_X2 \AES_ENC/us23/U14  ( .A1(\AES_ENC/us23/n1111 ), .A2(\AES_ENC/us23/n1110 ), .A3(\AES_ENC/us23/n1109 ), .A4(\AES_ENC/us23/n1108 ), .ZN(\AES_ENC/us23/n1112 ) );
NAND2_X2 \AES_ENC/us23/U13  ( .A1(\AES_ENC/us23/n1113 ), .A2(\AES_ENC/us23/n1112 ), .ZN(\AES_ENC/us23/n1133 ) );
NAND2_X2 \AES_ENC/us23/U12  ( .A1(\AES_ENC/us23/n1115 ), .A2(\AES_ENC/us23/n1114 ), .ZN(\AES_ENC/us23/n1129 ) );
OR2_X2 \AES_ENC/us23/U11  ( .A1(\AES_ENC/us23/n579 ), .A2(\AES_ENC/us23/n1116 ), .ZN(\AES_ENC/us23/n1128 ) );
NAND4_X2 \AES_ENC/us23/U3  ( .A1(\AES_ENC/us23/n1129 ), .A2(\AES_ENC/us23/n1128 ), .A3(\AES_ENC/us23/n1127 ), .A4(\AES_ENC/us23/n1126 ), .ZN(\AES_ENC/us23/n1130 ) );
NAND2_X2 \AES_ENC/us23/U2  ( .A1(\AES_ENC/us23/n1131 ), .A2(\AES_ENC/us23/n1130 ), .ZN(\AES_ENC/us23/n1132 ) );
NAND4_X2 \AES_ENC/us23/U1  ( .A1(\AES_ENC/us23/n1135 ), .A2(\AES_ENC/us23/n1134 ), .A3(\AES_ENC/us23/n1133 ), .A4(\AES_ENC/us23/n1132 ), .ZN(\AES_ENC/sa23_sub[7] ) );
INV_X4 \AES_ENC/us30/U575  ( .A(\AES_ENC/sa30 [7]), .ZN(\AES_ENC/us30/n627 ));
INV_X4 \AES_ENC/us30/U574  ( .A(\AES_ENC/us30/n1114 ), .ZN(\AES_ENC/us30/n625 ) );
INV_X4 \AES_ENC/us30/U573  ( .A(\AES_ENC/sa30 [4]), .ZN(\AES_ENC/us30/n624 ));
INV_X4 \AES_ENC/us30/U572  ( .A(\AES_ENC/us30/n1025 ), .ZN(\AES_ENC/us30/n622 ) );
INV_X4 \AES_ENC/us30/U571  ( .A(\AES_ENC/us30/n1120 ), .ZN(\AES_ENC/us30/n620 ) );
INV_X4 \AES_ENC/us30/U570  ( .A(\AES_ENC/us30/n1121 ), .ZN(\AES_ENC/us30/n619 ) );
INV_X4 \AES_ENC/us30/U569  ( .A(\AES_ENC/us30/n1048 ), .ZN(\AES_ENC/us30/n618 ) );
INV_X4 \AES_ENC/us30/U568  ( .A(\AES_ENC/us30/n974 ), .ZN(\AES_ENC/us30/n616 ) );
INV_X4 \AES_ENC/us30/U567  ( .A(\AES_ENC/us30/n794 ), .ZN(\AES_ENC/us30/n614 ) );
INV_X4 \AES_ENC/us30/U566  ( .A(\AES_ENC/sa30 [2]), .ZN(\AES_ENC/us30/n611 ));
INV_X4 \AES_ENC/us30/U565  ( .A(\AES_ENC/us30/n800 ), .ZN(\AES_ENC/us30/n610 ) );
INV_X4 \AES_ENC/us30/U564  ( .A(\AES_ENC/us30/n925 ), .ZN(\AES_ENC/us30/n609 ) );
INV_X4 \AES_ENC/us30/U563  ( .A(\AES_ENC/us30/n779 ), .ZN(\AES_ENC/us30/n607 ) );
INV_X4 \AES_ENC/us30/U562  ( .A(\AES_ENC/us30/n1022 ), .ZN(\AES_ENC/us30/n603 ) );
INV_X4 \AES_ENC/us30/U561  ( .A(\AES_ENC/us30/n1102 ), .ZN(\AES_ENC/us30/n602 ) );
INV_X4 \AES_ENC/us30/U560  ( .A(\AES_ENC/us30/n929 ), .ZN(\AES_ENC/us30/n601 ) );
INV_X4 \AES_ENC/us30/U559  ( .A(\AES_ENC/us30/n1056 ), .ZN(\AES_ENC/us30/n600 ) );
INV_X4 \AES_ENC/us30/U558  ( .A(\AES_ENC/us30/n1054 ), .ZN(\AES_ENC/us30/n599 ) );
INV_X4 \AES_ENC/us30/U557  ( .A(\AES_ENC/us30/n881 ), .ZN(\AES_ENC/us30/n598 ) );
INV_X4 \AES_ENC/us30/U556  ( .A(\AES_ENC/us30/n926 ), .ZN(\AES_ENC/us30/n597 ) );
INV_X4 \AES_ENC/us30/U555  ( .A(\AES_ENC/us30/n977 ), .ZN(\AES_ENC/us30/n595 ) );
INV_X4 \AES_ENC/us30/U554  ( .A(\AES_ENC/us30/n1031 ), .ZN(\AES_ENC/us30/n594 ) );
INV_X4 \AES_ENC/us30/U553  ( .A(\AES_ENC/us30/n1103 ), .ZN(\AES_ENC/us30/n593 ) );
INV_X4 \AES_ENC/us30/U552  ( .A(\AES_ENC/us30/n1009 ), .ZN(\AES_ENC/us30/n592 ) );
INV_X4 \AES_ENC/us30/U551  ( .A(\AES_ENC/us30/n990 ), .ZN(\AES_ENC/us30/n591 ) );
INV_X4 \AES_ENC/us30/U550  ( .A(\AES_ENC/us30/n1058 ), .ZN(\AES_ENC/us30/n590 ) );
INV_X4 \AES_ENC/us30/U549  ( .A(\AES_ENC/us30/n1074 ), .ZN(\AES_ENC/us30/n589 ) );
INV_X4 \AES_ENC/us30/U548  ( .A(\AES_ENC/us30/n1053 ), .ZN(\AES_ENC/us30/n588 ) );
INV_X4 \AES_ENC/us30/U547  ( .A(\AES_ENC/us30/n826 ), .ZN(\AES_ENC/us30/n587 ) );
INV_X4 \AES_ENC/us30/U546  ( .A(\AES_ENC/us30/n992 ), .ZN(\AES_ENC/us30/n586 ) );
INV_X4 \AES_ENC/us30/U545  ( .A(\AES_ENC/us30/n821 ), .ZN(\AES_ENC/us30/n585 ) );
INV_X4 \AES_ENC/us30/U544  ( .A(\AES_ENC/us30/n910 ), .ZN(\AES_ENC/us30/n584 ) );
INV_X4 \AES_ENC/us30/U543  ( .A(\AES_ENC/us30/n906 ), .ZN(\AES_ENC/us30/n583 ) );
INV_X4 \AES_ENC/us30/U542  ( .A(\AES_ENC/us30/n880 ), .ZN(\AES_ENC/us30/n581 ) );
INV_X4 \AES_ENC/us30/U541  ( .A(\AES_ENC/us30/n1013 ), .ZN(\AES_ENC/us30/n580 ) );
INV_X4 \AES_ENC/us30/U540  ( .A(\AES_ENC/us30/n1092 ), .ZN(\AES_ENC/us30/n579 ) );
INV_X4 \AES_ENC/us30/U539  ( .A(\AES_ENC/us30/n824 ), .ZN(\AES_ENC/us30/n578 ) );
INV_X4 \AES_ENC/us30/U538  ( .A(\AES_ENC/us30/n1091 ), .ZN(\AES_ENC/us30/n577 ) );
INV_X4 \AES_ENC/us30/U537  ( .A(\AES_ENC/us30/n1080 ), .ZN(\AES_ENC/us30/n576 ) );
INV_X4 \AES_ENC/us30/U536  ( .A(\AES_ENC/us30/n959 ), .ZN(\AES_ENC/us30/n575 ) );
INV_X4 \AES_ENC/us30/U535  ( .A(\AES_ENC/sa30 [0]), .ZN(\AES_ENC/us30/n574 ));
NOR2_X2 \AES_ENC/us30/U534  ( .A1(\AES_ENC/us30/n574 ), .A2(\AES_ENC/sa30 [6]), .ZN(\AES_ENC/us30/n1070 ) );
NOR2_X2 \AES_ENC/us30/U533  ( .A1(\AES_ENC/sa30 [0]), .A2(\AES_ENC/sa30 [6]),.ZN(\AES_ENC/us30/n1090 ) );
NOR2_X2 \AES_ENC/us30/U532  ( .A1(\AES_ENC/sa30 [4]), .A2(\AES_ENC/sa30 [3]),.ZN(\AES_ENC/us30/n1025 ) );
INV_X4 \AES_ENC/us30/U531  ( .A(\AES_ENC/us30/n569 ), .ZN(\AES_ENC/us30/n572 ) );
NOR2_X2 \AES_ENC/us30/U530  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n765 ) );
NOR2_X2 \AES_ENC/us30/U529  ( .A1(\AES_ENC/sa30 [4]), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n764 ) );
NOR2_X2 \AES_ENC/us30/U528  ( .A1(\AES_ENC/us30/n765 ), .A2(\AES_ENC/us30/n764 ), .ZN(\AES_ENC/us30/n766 ) );
NOR2_X2 \AES_ENC/us30/U527  ( .A1(\AES_ENC/us30/n766 ), .A2(\AES_ENC/us30/n575 ), .ZN(\AES_ENC/us30/n767 ) );
NOR3_X2 \AES_ENC/us30/U526  ( .A1(\AES_ENC/us30/n627 ), .A2(\AES_ENC/sa30 [5]), .A3(\AES_ENC/us30/n704 ), .ZN(\AES_ENC/us30/n706 ));
NOR2_X2 \AES_ENC/us30/U525  ( .A1(\AES_ENC/us30/n1117 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n707 ) );
NOR2_X2 \AES_ENC/us30/U524  ( .A1(\AES_ENC/sa30 [4]), .A2(\AES_ENC/us30/n579 ), .ZN(\AES_ENC/us30/n705 ) );
NOR3_X2 \AES_ENC/us30/U523  ( .A1(\AES_ENC/us30/n707 ), .A2(\AES_ENC/us30/n706 ), .A3(\AES_ENC/us30/n705 ), .ZN(\AES_ENC/us30/n713 ) );
INV_X4 \AES_ENC/us30/U522  ( .A(\AES_ENC/sa30 [3]), .ZN(\AES_ENC/us30/n621 ));
NAND3_X2 \AES_ENC/us30/U521  ( .A1(\AES_ENC/us30/n652 ), .A2(\AES_ENC/us30/n626 ), .A3(\AES_ENC/sa30 [7]), .ZN(\AES_ENC/us30/n653 ));
NOR2_X2 \AES_ENC/us30/U520  ( .A1(\AES_ENC/us30/n611 ), .A2(\AES_ENC/sa30 [5]), .ZN(\AES_ENC/us30/n925 ) );
NOR2_X2 \AES_ENC/us30/U519  ( .A1(\AES_ENC/sa30 [5]), .A2(\AES_ENC/sa30 [2]),.ZN(\AES_ENC/us30/n974 ) );
INV_X4 \AES_ENC/us30/U518  ( .A(\AES_ENC/sa30 [5]), .ZN(\AES_ENC/us30/n626 ));
NOR2_X2 \AES_ENC/us30/U517  ( .A1(\AES_ENC/us30/n611 ), .A2(\AES_ENC/sa30 [7]), .ZN(\AES_ENC/us30/n779 ) );
NAND3_X2 \AES_ENC/us30/U516  ( .A1(\AES_ENC/us30/n679 ), .A2(\AES_ENC/us30/n678 ), .A3(\AES_ENC/us30/n677 ), .ZN(\AES_ENC/sa30_sub[0] ) );
NOR2_X2 \AES_ENC/us30/U515  ( .A1(\AES_ENC/us30/n626 ), .A2(\AES_ENC/sa30 [2]), .ZN(\AES_ENC/us30/n1048 ) );
NOR4_X2 \AES_ENC/us30/U512  ( .A1(\AES_ENC/us30/n633 ), .A2(\AES_ENC/us30/n632 ), .A3(\AES_ENC/us30/n631 ), .A4(\AES_ENC/us30/n630 ), .ZN(\AES_ENC/us30/n634 ) );
NOR2_X2 \AES_ENC/us30/U510  ( .A1(\AES_ENC/us30/n629 ), .A2(\AES_ENC/us30/n628 ), .ZN(\AES_ENC/us30/n635 ) );
NAND3_X2 \AES_ENC/us30/U509  ( .A1(\AES_ENC/sa30 [2]), .A2(\AES_ENC/sa30 [7]), .A3(\AES_ENC/us30/n1059 ), .ZN(\AES_ENC/us30/n636 ) );
NOR2_X2 \AES_ENC/us30/U508  ( .A1(\AES_ENC/sa30 [7]), .A2(\AES_ENC/sa30 [2]),.ZN(\AES_ENC/us30/n794 ) );
NOR2_X2 \AES_ENC/us30/U507  ( .A1(\AES_ENC/sa30 [4]), .A2(\AES_ENC/sa30 [1]),.ZN(\AES_ENC/us30/n1102 ) );
NOR2_X2 \AES_ENC/us30/U506  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/sa30 [3]), .ZN(\AES_ENC/us30/n1053 ) );
NOR2_X2 \AES_ENC/us30/U505  ( .A1(\AES_ENC/us30/n607 ), .A2(\AES_ENC/sa30 [5]), .ZN(\AES_ENC/us30/n1024 ) );
NOR2_X2 \AES_ENC/us30/U504  ( .A1(\AES_ENC/us30/n625 ), .A2(\AES_ENC/sa30 [2]), .ZN(\AES_ENC/us30/n1093 ) );
NOR2_X2 \AES_ENC/us30/U503  ( .A1(\AES_ENC/us30/n614 ), .A2(\AES_ENC/sa30 [5]), .ZN(\AES_ENC/us30/n1094 ) );
NOR2_X2 \AES_ENC/us30/U502  ( .A1(\AES_ENC/us30/n624 ), .A2(\AES_ENC/sa30 [3]), .ZN(\AES_ENC/us30/n931 ) );
INV_X4 \AES_ENC/us30/U501  ( .A(\AES_ENC/us30/n570 ), .ZN(\AES_ENC/us30/n573 ) );
NOR2_X2 \AES_ENC/us30/U500  ( .A1(\AES_ENC/us30/n1053 ), .A2(\AES_ENC/us30/n1095 ), .ZN(\AES_ENC/us30/n639 ) );
NOR3_X2 \AES_ENC/us30/U499  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n573 ), .A3(\AES_ENC/us30/n1074 ), .ZN(\AES_ENC/us30/n641 ) );
NOR2_X2 \AES_ENC/us30/U498  ( .A1(\AES_ENC/us30/n639 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n640 ) );
NOR2_X2 \AES_ENC/us30/U497  ( .A1(\AES_ENC/us30/n641 ), .A2(\AES_ENC/us30/n640 ), .ZN(\AES_ENC/us30/n646 ) );
NOR3_X2 \AES_ENC/us30/U496  ( .A1(\AES_ENC/us30/n995 ), .A2(\AES_ENC/us30/n586 ), .A3(\AES_ENC/us30/n994 ), .ZN(\AES_ENC/us30/n1002 ) );
NOR2_X2 \AES_ENC/us30/U495  ( .A1(\AES_ENC/us30/n909 ), .A2(\AES_ENC/us30/n908 ), .ZN(\AES_ENC/us30/n920 ) );
NOR2_X2 \AES_ENC/us30/U494  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n823 ) );
NOR2_X2 \AES_ENC/us30/U492  ( .A1(\AES_ENC/us30/n624 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n822 ) );
NOR2_X2 \AES_ENC/us30/U491  ( .A1(\AES_ENC/us30/n823 ), .A2(\AES_ENC/us30/n822 ), .ZN(\AES_ENC/us30/n825 ) );
NOR2_X2 \AES_ENC/us30/U490  ( .A1(\AES_ENC/sa30 [1]), .A2(\AES_ENC/us30/n623 ), .ZN(\AES_ENC/us30/n913 ) );
NOR2_X2 \AES_ENC/us30/U489  ( .A1(\AES_ENC/us30/n913 ), .A2(\AES_ENC/us30/n1091 ), .ZN(\AES_ENC/us30/n914 ) );
NOR2_X2 \AES_ENC/us30/U488  ( .A1(\AES_ENC/us30/n826 ), .A2(\AES_ENC/us30/n572 ), .ZN(\AES_ENC/us30/n827 ) );
NOR3_X2 \AES_ENC/us30/U487  ( .A1(\AES_ENC/us30/n769 ), .A2(\AES_ENC/us30/n768 ), .A3(\AES_ENC/us30/n767 ), .ZN(\AES_ENC/us30/n775 ) );
NOR2_X2 \AES_ENC/us30/U486  ( .A1(\AES_ENC/us30/n1056 ), .A2(\AES_ENC/us30/n1053 ), .ZN(\AES_ENC/us30/n749 ) );
NOR2_X2 \AES_ENC/us30/U483  ( .A1(\AES_ENC/us30/n749 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n752 ) );
INV_X4 \AES_ENC/us30/U482  ( .A(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n596 ));
NOR2_X2 \AES_ENC/us30/U480  ( .A1(\AES_ENC/us30/n1054 ), .A2(\AES_ENC/us30/n1053 ), .ZN(\AES_ENC/us30/n1055 ) );
OR2_X4 \AES_ENC/us30/U479  ( .A1(\AES_ENC/us30/n1094 ), .A2(\AES_ENC/us30/n1093 ), .ZN(\AES_ENC/us30/n571 ) );
AND2_X2 \AES_ENC/us30/U478  ( .A1(\AES_ENC/us30/n571 ), .A2(\AES_ENC/us30/n1095 ), .ZN(\AES_ENC/us30/n1101 ) );
NOR2_X2 \AES_ENC/us30/U477  ( .A1(\AES_ENC/us30/n1074 ), .A2(\AES_ENC/us30/n931 ), .ZN(\AES_ENC/us30/n796 ) );
NOR2_X2 \AES_ENC/us30/U474  ( .A1(\AES_ENC/us30/n796 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n797 ) );
NOR2_X2 \AES_ENC/us30/U473  ( .A1(\AES_ENC/us30/n932 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n933 ) );
NOR2_X2 \AES_ENC/us30/U472  ( .A1(\AES_ENC/us30/n929 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n935 ) );
NOR2_X2 \AES_ENC/us30/U471  ( .A1(\AES_ENC/us30/n931 ), .A2(\AES_ENC/us30/n930 ), .ZN(\AES_ENC/us30/n934 ) );
NOR3_X2 \AES_ENC/us30/U470  ( .A1(\AES_ENC/us30/n935 ), .A2(\AES_ENC/us30/n934 ), .A3(\AES_ENC/us30/n933 ), .ZN(\AES_ENC/us30/n936 ) );
NOR2_X2 \AES_ENC/us30/U469  ( .A1(\AES_ENC/us30/n624 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n1075 ) );
NOR2_X2 \AES_ENC/us30/U468  ( .A1(\AES_ENC/us30/n572 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n949 ) );
NOR2_X2 \AES_ENC/us30/U467  ( .A1(\AES_ENC/us30/n1049 ), .A2(\AES_ENC/us30/n618 ), .ZN(\AES_ENC/us30/n1051 ) );
NOR2_X2 \AES_ENC/us30/U466  ( .A1(\AES_ENC/us30/n1051 ), .A2(\AES_ENC/us30/n1050 ), .ZN(\AES_ENC/us30/n1052 ) );
NOR2_X2 \AES_ENC/us30/U465  ( .A1(\AES_ENC/us30/n1052 ), .A2(\AES_ENC/us30/n592 ), .ZN(\AES_ENC/us30/n1064 ) );
NOR2_X2 \AES_ENC/us30/U464  ( .A1(\AES_ENC/sa30 [1]), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n631 ) );
NOR2_X2 \AES_ENC/us30/U463  ( .A1(\AES_ENC/us30/n1025 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n980 ) );
NOR2_X2 \AES_ENC/us30/U462  ( .A1(\AES_ENC/us30/n1073 ), .A2(\AES_ENC/us30/n1094 ), .ZN(\AES_ENC/us30/n795 ) );
NOR2_X2 \AES_ENC/us30/U461  ( .A1(\AES_ENC/us30/n795 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n799 ) );
NOR2_X2 \AES_ENC/us30/U460  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n981 ) );
NOR2_X2 \AES_ENC/us30/U459  ( .A1(\AES_ENC/us30/n1102 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n643 ) );
NOR2_X2 \AES_ENC/us30/U458  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n621 ), .ZN(\AES_ENC/us30/n642 ) );
NOR2_X2 \AES_ENC/us30/U455  ( .A1(\AES_ENC/us30/n911 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n644 ) );
NOR4_X2 \AES_ENC/us30/U448  ( .A1(\AES_ENC/us30/n644 ), .A2(\AES_ENC/us30/n643 ), .A3(\AES_ENC/us30/n804 ), .A4(\AES_ENC/us30/n642 ), .ZN(\AES_ENC/us30/n645 ) );
NOR2_X2 \AES_ENC/us30/U447  ( .A1(\AES_ENC/us30/n1102 ), .A2(\AES_ENC/us30/n910 ), .ZN(\AES_ENC/us30/n932 ) );
NOR2_X2 \AES_ENC/us30/U442  ( .A1(\AES_ENC/us30/n1102 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n755 ) );
NOR2_X2 \AES_ENC/us30/U441  ( .A1(\AES_ENC/us30/n931 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n743 ) );
NOR2_X2 \AES_ENC/us30/U438  ( .A1(\AES_ENC/us30/n1072 ), .A2(\AES_ENC/us30/n1094 ), .ZN(\AES_ENC/us30/n930 ) );
NOR2_X2 \AES_ENC/us30/U435  ( .A1(\AES_ENC/us30/n1074 ), .A2(\AES_ENC/us30/n1025 ), .ZN(\AES_ENC/us30/n891 ) );
NOR2_X2 \AES_ENC/us30/U434  ( .A1(\AES_ENC/us30/n891 ), .A2(\AES_ENC/us30/n609 ), .ZN(\AES_ENC/us30/n894 ) );
NOR3_X2 \AES_ENC/us30/U433  ( .A1(\AES_ENC/us30/n623 ), .A2(\AES_ENC/sa30 [1]), .A3(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n683 ));
INV_X4 \AES_ENC/us30/U428  ( .A(\AES_ENC/us30/n931 ), .ZN(\AES_ENC/us30/n623 ) );
NOR2_X2 \AES_ENC/us30/U427  ( .A1(\AES_ENC/us30/n996 ), .A2(\AES_ENC/us30/n931 ), .ZN(\AES_ENC/us30/n704 ) );
NOR2_X2 \AES_ENC/us30/U421  ( .A1(\AES_ENC/us30/n931 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n685 ) );
NOR2_X2 \AES_ENC/us30/U420  ( .A1(\AES_ENC/us30/n1029 ), .A2(\AES_ENC/us30/n1025 ), .ZN(\AES_ENC/us30/n1079 ) );
NOR3_X2 \AES_ENC/us30/U419  ( .A1(\AES_ENC/us30/n589 ), .A2(\AES_ENC/us30/n1025 ), .A3(\AES_ENC/us30/n616 ), .ZN(\AES_ENC/us30/n945 ) );
NOR2_X2 \AES_ENC/us30/U418  ( .A1(\AES_ENC/us30/n626 ), .A2(\AES_ENC/us30/n611 ), .ZN(\AES_ENC/us30/n800 ) );
NOR3_X2 \AES_ENC/us30/U417  ( .A1(\AES_ENC/us30/n590 ), .A2(\AES_ENC/us30/n627 ), .A3(\AES_ENC/us30/n611 ), .ZN(\AES_ENC/us30/n798 ) );
NOR3_X2 \AES_ENC/us30/U416  ( .A1(\AES_ENC/us30/n610 ), .A2(\AES_ENC/us30/n572 ), .A3(\AES_ENC/us30/n575 ), .ZN(\AES_ENC/us30/n962 ) );
NOR3_X2 \AES_ENC/us30/U415  ( .A1(\AES_ENC/us30/n959 ), .A2(\AES_ENC/us30/n572 ), .A3(\AES_ENC/us30/n609 ), .ZN(\AES_ENC/us30/n768 ) );
NOR3_X2 \AES_ENC/us30/U414  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n572 ), .A3(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n694 ) );
NOR3_X2 \AES_ENC/us30/U413  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n572 ), .A3(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n895 ) );
NOR3_X2 \AES_ENC/us30/U410  ( .A1(\AES_ENC/us30/n1008 ), .A2(\AES_ENC/us30/n1007 ), .A3(\AES_ENC/us30/n1006 ), .ZN(\AES_ENC/us30/n1018 ) );
NOR4_X2 \AES_ENC/us30/U409  ( .A1(\AES_ENC/us30/n806 ), .A2(\AES_ENC/us30/n805 ), .A3(\AES_ENC/us30/n804 ), .A4(\AES_ENC/us30/n803 ), .ZN(\AES_ENC/us30/n807 ) );
NOR3_X2 \AES_ENC/us30/U406  ( .A1(\AES_ENC/us30/n799 ), .A2(\AES_ENC/us30/n798 ), .A3(\AES_ENC/us30/n797 ), .ZN(\AES_ENC/us30/n808 ) );
NOR4_X2 \AES_ENC/us30/U405  ( .A1(\AES_ENC/us30/n711 ), .A2(\AES_ENC/us30/n710 ), .A3(\AES_ENC/us30/n709 ), .A4(\AES_ENC/us30/n708 ), .ZN(\AES_ENC/us30/n712 ) );
NOR4_X2 \AES_ENC/us30/U404  ( .A1(\AES_ENC/us30/n963 ), .A2(\AES_ENC/us30/n962 ), .A3(\AES_ENC/us30/n961 ), .A4(\AES_ENC/us30/n960 ), .ZN(\AES_ENC/us30/n964 ) );
NOR3_X2 \AES_ENC/us30/U403  ( .A1(\AES_ENC/us30/n1101 ), .A2(\AES_ENC/us30/n1100 ), .A3(\AES_ENC/us30/n1099 ), .ZN(\AES_ENC/us30/n1109 ) );
NOR2_X2 \AES_ENC/us30/U401  ( .A1(\AES_ENC/us30/n669 ), .A2(\AES_ENC/us30/n668 ), .ZN(\AES_ENC/us30/n673 ) );
NOR4_X2 \AES_ENC/us30/U400  ( .A1(\AES_ENC/us30/n946 ), .A2(\AES_ENC/us30/n1046 ), .A3(\AES_ENC/us30/n671 ), .A4(\AES_ENC/us30/n670 ), .ZN(\AES_ENC/us30/n672 ) );
NOR4_X2 \AES_ENC/us30/U399  ( .A1(\AES_ENC/us30/n843 ), .A2(\AES_ENC/us30/n842 ), .A3(\AES_ENC/us30/n841 ), .A4(\AES_ENC/us30/n840 ), .ZN(\AES_ENC/us30/n844 ) );
NOR3_X2 \AES_ENC/us30/U398  ( .A1(\AES_ENC/us30/n743 ), .A2(\AES_ENC/us30/n742 ), .A3(\AES_ENC/us30/n741 ), .ZN(\AES_ENC/us30/n744 ) );
NOR2_X2 \AES_ENC/us30/U397  ( .A1(\AES_ENC/us30/n697 ), .A2(\AES_ENC/us30/n658 ), .ZN(\AES_ENC/us30/n659 ) );
NOR2_X2 \AES_ENC/us30/U396  ( .A1(\AES_ENC/us30/n1078 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n1033 ) );
NOR2_X2 \AES_ENC/us30/U393  ( .A1(\AES_ENC/us30/n1031 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n1032 ) );
NOR3_X2 \AES_ENC/us30/U390  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n1025 ), .A3(\AES_ENC/us30/n1074 ), .ZN(\AES_ENC/us30/n1035 ) );
NOR4_X2 \AES_ENC/us30/U389  ( .A1(\AES_ENC/us30/n1035 ), .A2(\AES_ENC/us30/n1034 ), .A3(\AES_ENC/us30/n1033 ), .A4(\AES_ENC/us30/n1032 ), .ZN(\AES_ENC/us30/n1036 ) );
NOR2_X2 \AES_ENC/us30/U388  ( .A1(\AES_ENC/us30/n598 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n885 ) );
NOR2_X2 \AES_ENC/us30/U387  ( .A1(\AES_ENC/us30/n623 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n882 ) );
NOR2_X2 \AES_ENC/us30/U386  ( .A1(\AES_ENC/us30/n1053 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n884 ) );
NOR4_X2 \AES_ENC/us30/U385  ( .A1(\AES_ENC/us30/n885 ), .A2(\AES_ENC/us30/n884 ), .A3(\AES_ENC/us30/n883 ), .A4(\AES_ENC/us30/n882 ), .ZN(\AES_ENC/us30/n886 ) );
NOR2_X2 \AES_ENC/us30/U384  ( .A1(\AES_ENC/us30/n825 ), .A2(\AES_ENC/us30/n578 ), .ZN(\AES_ENC/us30/n830 ) );
NOR2_X2 \AES_ENC/us30/U383  ( .A1(\AES_ENC/us30/n827 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n829 ) );
NOR2_X2 \AES_ENC/us30/U382  ( .A1(\AES_ENC/us30/n572 ), .A2(\AES_ENC/us30/n579 ), .ZN(\AES_ENC/us30/n828 ) );
NOR4_X2 \AES_ENC/us30/U374  ( .A1(\AES_ENC/us30/n831 ), .A2(\AES_ENC/us30/n830 ), .A3(\AES_ENC/us30/n829 ), .A4(\AES_ENC/us30/n828 ), .ZN(\AES_ENC/us30/n832 ) );
NOR2_X2 \AES_ENC/us30/U373  ( .A1(\AES_ENC/us30/n606 ), .A2(\AES_ENC/us30/n582 ), .ZN(\AES_ENC/us30/n1104 ) );
NOR2_X2 \AES_ENC/us30/U372  ( .A1(\AES_ENC/us30/n1102 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n1106 ) );
NOR2_X2 \AES_ENC/us30/U370  ( .A1(\AES_ENC/us30/n1103 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n1105 ) );
NOR4_X2 \AES_ENC/us30/U369  ( .A1(\AES_ENC/us30/n1107 ), .A2(\AES_ENC/us30/n1106 ), .A3(\AES_ENC/us30/n1105 ), .A4(\AES_ENC/us30/n1104 ), .ZN(\AES_ENC/us30/n1108 ) );
NOR3_X2 \AES_ENC/us30/U368  ( .A1(\AES_ENC/us30/n959 ), .A2(\AES_ENC/us30/n621 ), .A3(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n963 ) );
NOR2_X2 \AES_ENC/us30/U367  ( .A1(\AES_ENC/us30/n626 ), .A2(\AES_ENC/us30/n627 ), .ZN(\AES_ENC/us30/n1114 ) );
INV_X4 \AES_ENC/us30/U366  ( .A(\AES_ENC/us30/n1024 ), .ZN(\AES_ENC/us30/n606 ) );
NOR3_X2 \AES_ENC/us30/U365  ( .A1(\AES_ENC/us30/n910 ), .A2(\AES_ENC/us30/n1059 ), .A3(\AES_ENC/us30/n611 ), .ZN(\AES_ENC/us30/n1115 ) );
INV_X4 \AES_ENC/us30/U364  ( .A(\AES_ENC/us30/n1094 ), .ZN(\AES_ENC/us30/n613 ) );
NOR2_X2 \AES_ENC/us30/U363  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n931 ), .ZN(\AES_ENC/us30/n1100 ) );
INV_X4 \AES_ENC/us30/U354  ( .A(\AES_ENC/us30/n1093 ), .ZN(\AES_ENC/us30/n617 ) );
NOR2_X2 \AES_ENC/us30/U353  ( .A1(\AES_ENC/us30/n569 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n929 ) );
NOR2_X2 \AES_ENC/us30/U352  ( .A1(\AES_ENC/us30/n620 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n926 ) );
NOR2_X2 \AES_ENC/us30/U351  ( .A1(\AES_ENC/us30/n572 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n1095 ) );
NOR2_X2 \AES_ENC/us30/U350  ( .A1(\AES_ENC/us30/n609 ), .A2(\AES_ENC/us30/n627 ), .ZN(\AES_ENC/us30/n1010 ) );
NOR2_X2 \AES_ENC/us30/U349  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n1103 ) );
NOR2_X2 \AES_ENC/us30/U348  ( .A1(\AES_ENC/us30/n622 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n1059 ) );
NOR2_X2 \AES_ENC/us30/U347  ( .A1(\AES_ENC/sa30 [1]), .A2(\AES_ENC/us30/n1120 ), .ZN(\AES_ENC/us30/n1022 ) );
NOR2_X2 \AES_ENC/us30/U346  ( .A1(\AES_ENC/us30/n619 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n911 ) );
NOR2_X2 \AES_ENC/us30/U345  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/us30/n1025 ), .ZN(\AES_ENC/us30/n826 ) );
NOR2_X2 \AES_ENC/us30/U338  ( .A1(\AES_ENC/us30/n626 ), .A2(\AES_ENC/us30/n607 ), .ZN(\AES_ENC/us30/n1072 ) );
NOR2_X2 \AES_ENC/us30/U335  ( .A1(\AES_ENC/us30/n627 ), .A2(\AES_ENC/us30/n616 ), .ZN(\AES_ENC/us30/n956 ) );
NOR2_X2 \AES_ENC/us30/U329  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/us30/n624 ), .ZN(\AES_ENC/us30/n1121 ) );
NOR2_X2 \AES_ENC/us30/U328  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/us30/n624 ), .ZN(\AES_ENC/us30/n1058 ) );
NOR2_X2 \AES_ENC/us30/U327  ( .A1(\AES_ENC/us30/n625 ), .A2(\AES_ENC/us30/n611 ), .ZN(\AES_ENC/us30/n1073 ) );
NOR2_X2 \AES_ENC/us30/U325  ( .A1(\AES_ENC/sa30 [1]), .A2(\AES_ENC/us30/n1025 ), .ZN(\AES_ENC/us30/n1054 ) );
NOR2_X2 \AES_ENC/us30/U324  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/us30/n931 ), .ZN(\AES_ENC/us30/n1029 ) );
NOR2_X2 \AES_ENC/us30/U319  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n1056 ) );
NOR2_X2 \AES_ENC/us30/U318  ( .A1(\AES_ENC/us30/n614 ), .A2(\AES_ENC/us30/n626 ), .ZN(\AES_ENC/us30/n1050 ) );
NOR2_X2 \AES_ENC/us30/U317  ( .A1(\AES_ENC/us30/n1121 ), .A2(\AES_ENC/us30/n1025 ), .ZN(\AES_ENC/us30/n1120 ) );
NOR2_X2 \AES_ENC/us30/U316  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/us30/n572 ), .ZN(\AES_ENC/us30/n1074 ) );
NOR2_X2 \AES_ENC/us30/U315  ( .A1(\AES_ENC/us30/n1058 ), .A2(\AES_ENC/us30/n1054 ), .ZN(\AES_ENC/us30/n878 ) );
NOR2_X2 \AES_ENC/us30/U314  ( .A1(\AES_ENC/us30/n878 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n879 ) );
NOR2_X2 \AES_ENC/us30/U312  ( .A1(\AES_ENC/us30/n880 ), .A2(\AES_ENC/us30/n879 ), .ZN(\AES_ENC/us30/n887 ) );
NOR2_X2 \AES_ENC/us30/U311  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n588 ), .ZN(\AES_ENC/us30/n957 ) );
NOR2_X2 \AES_ENC/us30/U310  ( .A1(\AES_ENC/us30/n958 ), .A2(\AES_ENC/us30/n957 ), .ZN(\AES_ENC/us30/n965 ) );
NOR3_X2 \AES_ENC/us30/U309  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n1091 ), .A3(\AES_ENC/us30/n1022 ), .ZN(\AES_ENC/us30/n720 ) );
NOR3_X2 \AES_ENC/us30/U303  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n1054 ), .A3(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n719 ) );
NOR2_X2 \AES_ENC/us30/U302  ( .A1(\AES_ENC/us30/n720 ), .A2(\AES_ENC/us30/n719 ), .ZN(\AES_ENC/us30/n726 ) );
NOR2_X2 \AES_ENC/us30/U300  ( .A1(\AES_ENC/us30/n614 ), .A2(\AES_ENC/us30/n591 ), .ZN(\AES_ENC/us30/n865 ) );
NOR2_X2 \AES_ENC/us30/U299  ( .A1(\AES_ENC/us30/n1059 ), .A2(\AES_ENC/us30/n1058 ), .ZN(\AES_ENC/us30/n1060 ) );
NOR2_X2 \AES_ENC/us30/U298  ( .A1(\AES_ENC/us30/n1095 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n668 ) );
NOR2_X2 \AES_ENC/us30/U297  ( .A1(\AES_ENC/us30/n911 ), .A2(\AES_ENC/us30/n910 ), .ZN(\AES_ENC/us30/n912 ) );
NOR2_X2 \AES_ENC/us30/U296  ( .A1(\AES_ENC/us30/n912 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n916 ) );
NOR2_X2 \AES_ENC/us30/U295  ( .A1(\AES_ENC/us30/n826 ), .A2(\AES_ENC/us30/n573 ), .ZN(\AES_ENC/us30/n750 ) );
NOR2_X2 \AES_ENC/us30/U294  ( .A1(\AES_ENC/us30/n750 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n751 ) );
NOR2_X2 \AES_ENC/us30/U293  ( .A1(\AES_ENC/us30/n907 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n908 ) );
NOR2_X2 \AES_ENC/us30/U292  ( .A1(\AES_ENC/us30/n990 ), .A2(\AES_ENC/us30/n926 ), .ZN(\AES_ENC/us30/n780 ) );
NOR2_X2 \AES_ENC/us30/U291  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n584 ), .ZN(\AES_ENC/us30/n838 ) );
NOR2_X2 \AES_ENC/us30/U290  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n602 ), .ZN(\AES_ENC/us30/n837 ) );
NOR2_X2 \AES_ENC/us30/U284  ( .A1(\AES_ENC/us30/n838 ), .A2(\AES_ENC/us30/n837 ), .ZN(\AES_ENC/us30/n845 ) );
NOR2_X2 \AES_ENC/us30/U283  ( .A1(\AES_ENC/us30/n1022 ), .A2(\AES_ENC/us30/n1058 ), .ZN(\AES_ENC/us30/n740 ) );
NOR2_X2 \AES_ENC/us30/U282  ( .A1(\AES_ENC/us30/n740 ), .A2(\AES_ENC/us30/n616 ), .ZN(\AES_ENC/us30/n742 ) );
NOR2_X2 \AES_ENC/us30/U281  ( .A1(\AES_ENC/us30/n1098 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n1099 ) );
NOR2_X2 \AES_ENC/us30/U280  ( .A1(\AES_ENC/us30/n1120 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n993 ) );
NOR2_X2 \AES_ENC/us30/U279  ( .A1(\AES_ENC/us30/n993 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n994 ) );
NOR2_X2 \AES_ENC/us30/U273  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n620 ), .ZN(\AES_ENC/us30/n1026 ) );
NOR2_X2 \AES_ENC/us30/U272  ( .A1(\AES_ENC/us30/n573 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n1027 ) );
NOR2_X2 \AES_ENC/us30/U271  ( .A1(\AES_ENC/us30/n1027 ), .A2(\AES_ENC/us30/n1026 ), .ZN(\AES_ENC/us30/n1028 ) );
NOR2_X2 \AES_ENC/us30/U270  ( .A1(\AES_ENC/us30/n1029 ), .A2(\AES_ENC/us30/n1028 ), .ZN(\AES_ENC/us30/n1034 ) );
NOR4_X2 \AES_ENC/us30/U269  ( .A1(\AES_ENC/us30/n757 ), .A2(\AES_ENC/us30/n756 ), .A3(\AES_ENC/us30/n755 ), .A4(\AES_ENC/us30/n754 ), .ZN(\AES_ENC/us30/n758 ) );
NOR2_X2 \AES_ENC/us30/U268  ( .A1(\AES_ENC/us30/n752 ), .A2(\AES_ENC/us30/n751 ), .ZN(\AES_ENC/us30/n759 ) );
NOR2_X2 \AES_ENC/us30/U267  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n1071 ), .ZN(\AES_ENC/us30/n669 ) );
NOR2_X2 \AES_ENC/us30/U263  ( .A1(\AES_ENC/us30/n1056 ), .A2(\AES_ENC/us30/n990 ), .ZN(\AES_ENC/us30/n991 ) );
NOR2_X2 \AES_ENC/us30/U262  ( .A1(\AES_ENC/us30/n991 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n995 ) );
NOR2_X2 \AES_ENC/us30/U258  ( .A1(\AES_ENC/us30/n607 ), .A2(\AES_ENC/us30/n590 ), .ZN(\AES_ENC/us30/n1008 ) );
NOR2_X2 \AES_ENC/us30/U255  ( .A1(\AES_ENC/us30/n839 ), .A2(\AES_ENC/us30/n582 ), .ZN(\AES_ENC/us30/n693 ) );
NOR2_X2 \AES_ENC/us30/U254  ( .A1(\AES_ENC/us30/n606 ), .A2(\AES_ENC/us30/n906 ), .ZN(\AES_ENC/us30/n741 ) );
NOR2_X2 \AES_ENC/us30/U253  ( .A1(\AES_ENC/us30/n1054 ), .A2(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n763 ) );
NOR2_X2 \AES_ENC/us30/U252  ( .A1(\AES_ENC/us30/n763 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n769 ) );
NOR2_X2 \AES_ENC/us30/U251  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n577 ), .ZN(\AES_ENC/us30/n1007 ) );
NOR2_X2 \AES_ENC/us30/U250  ( .A1(\AES_ENC/us30/n609 ), .A2(\AES_ENC/us30/n580 ), .ZN(\AES_ENC/us30/n1123 ) );
NOR2_X2 \AES_ENC/us30/U243  ( .A1(\AES_ENC/us30/n609 ), .A2(\AES_ENC/us30/n590 ), .ZN(\AES_ENC/us30/n710 ) );
INV_X4 \AES_ENC/us30/U242  ( .A(\AES_ENC/us30/n1029 ), .ZN(\AES_ENC/us30/n582 ) );
NOR2_X2 \AES_ENC/us30/U241  ( .A1(\AES_ENC/us30/n616 ), .A2(\AES_ENC/us30/n597 ), .ZN(\AES_ENC/us30/n883 ) );
NOR2_X2 \AES_ENC/us30/U240  ( .A1(\AES_ENC/us30/n593 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n1125 ) );
NOR2_X2 \AES_ENC/us30/U239  ( .A1(\AES_ENC/us30/n990 ), .A2(\AES_ENC/us30/n929 ), .ZN(\AES_ENC/us30/n892 ) );
NOR2_X2 \AES_ENC/us30/U238  ( .A1(\AES_ENC/us30/n892 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n893 ) );
NOR2_X2 \AES_ENC/us30/U237  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n602 ), .ZN(\AES_ENC/us30/n950 ) );
NOR2_X2 \AES_ENC/us30/U236  ( .A1(\AES_ENC/us30/n1079 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n1082 ) );
NOR2_X2 \AES_ENC/us30/U235  ( .A1(\AES_ENC/us30/n910 ), .A2(\AES_ENC/us30/n1056 ), .ZN(\AES_ENC/us30/n941 ) );
NOR2_X2 \AES_ENC/us30/U234  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n1077 ), .ZN(\AES_ENC/us30/n841 ) );
NOR2_X2 \AES_ENC/us30/U229  ( .A1(\AES_ENC/us30/n623 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n630 ) );
NOR2_X2 \AES_ENC/us30/U228  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n602 ), .ZN(\AES_ENC/us30/n806 ) );
NOR2_X2 \AES_ENC/us30/U227  ( .A1(\AES_ENC/us30/n623 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n948 ) );
NOR2_X2 \AES_ENC/us30/U226  ( .A1(\AES_ENC/us30/n606 ), .A2(\AES_ENC/us30/n589 ), .ZN(\AES_ENC/us30/n997 ) );
NOR2_X2 \AES_ENC/us30/U225  ( .A1(\AES_ENC/us30/n1121 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n1122 ) );
NOR2_X2 \AES_ENC/us30/U223  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n1023 ), .ZN(\AES_ENC/us30/n756 ) );
NOR2_X2 \AES_ENC/us30/U222  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n602 ), .ZN(\AES_ENC/us30/n870 ) );
NOR2_X2 \AES_ENC/us30/U221  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n569 ), .ZN(\AES_ENC/us30/n947 ) );
NOR2_X2 \AES_ENC/us30/U217  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n1077 ), .ZN(\AES_ENC/us30/n1084 ) );
NOR2_X2 \AES_ENC/us30/U213  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n855 ), .ZN(\AES_ENC/us30/n709 ) );
NOR2_X2 \AES_ENC/us30/U212  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n589 ), .ZN(\AES_ENC/us30/n868 ) );
NOR2_X2 \AES_ENC/us30/U211  ( .A1(\AES_ENC/us30/n1120 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n1124 ) );
NOR2_X2 \AES_ENC/us30/U210  ( .A1(\AES_ENC/us30/n1120 ), .A2(\AES_ENC/us30/n839 ), .ZN(\AES_ENC/us30/n842 ) );
NOR2_X2 \AES_ENC/us30/U209  ( .A1(\AES_ENC/us30/n1120 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n696 ) );
NOR2_X2 \AES_ENC/us30/U208  ( .A1(\AES_ENC/us30/n1074 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n1076 ) );
NOR2_X2 \AES_ENC/us30/U207  ( .A1(\AES_ENC/us30/n1074 ), .A2(\AES_ENC/us30/n620 ), .ZN(\AES_ENC/us30/n781 ) );
NOR3_X2 \AES_ENC/us30/U201  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n1056 ), .A3(\AES_ENC/us30/n990 ), .ZN(\AES_ENC/us30/n979 ) );
NOR3_X2 \AES_ENC/us30/U200  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n1058 ), .A3(\AES_ENC/us30/n1059 ), .ZN(\AES_ENC/us30/n854 ) );
NOR2_X2 \AES_ENC/us30/U199  ( .A1(\AES_ENC/us30/n996 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n869 ) );
NOR2_X2 \AES_ENC/us30/U198  ( .A1(\AES_ENC/us30/n1056 ), .A2(\AES_ENC/us30/n1074 ), .ZN(\AES_ENC/us30/n1057 ) );
NOR3_X2 \AES_ENC/us30/U197  ( .A1(\AES_ENC/us30/n607 ), .A2(\AES_ENC/us30/n1120 ), .A3(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n978 ) );
NOR2_X2 \AES_ENC/us30/U196  ( .A1(\AES_ENC/us30/n996 ), .A2(\AES_ENC/us30/n911 ), .ZN(\AES_ENC/us30/n1116 ) );
NOR2_X2 \AES_ENC/us30/U195  ( .A1(\AES_ENC/us30/n1074 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n754 ) );
NOR2_X2 \AES_ENC/us30/U194  ( .A1(\AES_ENC/us30/n926 ), .A2(\AES_ENC/us30/n1103 ), .ZN(\AES_ENC/us30/n977 ) );
NOR2_X2 \AES_ENC/us30/U187  ( .A1(\AES_ENC/us30/n839 ), .A2(\AES_ENC/us30/n824 ), .ZN(\AES_ENC/us30/n1092 ) );
NOR2_X2 \AES_ENC/us30/U186  ( .A1(\AES_ENC/us30/n573 ), .A2(\AES_ENC/us30/n1074 ), .ZN(\AES_ENC/us30/n684 ) );
NOR2_X2 \AES_ENC/us30/U185  ( .A1(\AES_ENC/us30/n826 ), .A2(\AES_ENC/us30/n1059 ), .ZN(\AES_ENC/us30/n907 ) );
NOR3_X2 \AES_ENC/us30/U184  ( .A1(\AES_ENC/us30/n625 ), .A2(\AES_ENC/us30/n1115 ), .A3(\AES_ENC/us30/n585 ), .ZN(\AES_ENC/us30/n831 ) );
NOR3_X2 \AES_ENC/us30/U183  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n1056 ), .A3(\AES_ENC/us30/n990 ), .ZN(\AES_ENC/us30/n896 ) );
NOR3_X2 \AES_ENC/us30/U182  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n573 ), .A3(\AES_ENC/us30/n1013 ), .ZN(\AES_ENC/us30/n670 ) );
NOR3_X2 \AES_ENC/us30/U181  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n1091 ), .A3(\AES_ENC/us30/n1022 ), .ZN(\AES_ENC/us30/n843 ) );
NOR2_X2 \AES_ENC/us30/U180  ( .A1(\AES_ENC/us30/n1029 ), .A2(\AES_ENC/us30/n1095 ), .ZN(\AES_ENC/us30/n735 ) );
NOR2_X2 \AES_ENC/us30/U174  ( .A1(\AES_ENC/us30/n1100 ), .A2(\AES_ENC/us30/n854 ), .ZN(\AES_ENC/us30/n860 ) );
NAND3_X2 \AES_ENC/us30/U173  ( .A1(\AES_ENC/us30/n569 ), .A2(\AES_ENC/us30/n582 ), .A3(\AES_ENC/us30/n681 ), .ZN(\AES_ENC/us30/n691 ) );
NOR2_X2 \AES_ENC/us30/U172  ( .A1(\AES_ENC/us30/n683 ), .A2(\AES_ENC/us30/n682 ), .ZN(\AES_ENC/us30/n690 ) );
NOR3_X2 \AES_ENC/us30/U171  ( .A1(\AES_ENC/us30/n695 ), .A2(\AES_ENC/us30/n694 ), .A3(\AES_ENC/us30/n693 ), .ZN(\AES_ENC/us30/n700 ) );
NOR4_X2 \AES_ENC/us30/U170  ( .A1(\AES_ENC/us30/n983 ), .A2(\AES_ENC/us30/n698 ), .A3(\AES_ENC/us30/n697 ), .A4(\AES_ENC/us30/n696 ), .ZN(\AES_ENC/us30/n699 ) );
NOR2_X2 \AES_ENC/us30/U169  ( .A1(\AES_ENC/us30/n946 ), .A2(\AES_ENC/us30/n945 ), .ZN(\AES_ENC/us30/n952 ) );
NOR4_X2 \AES_ENC/us30/U168  ( .A1(\AES_ENC/us30/n950 ), .A2(\AES_ENC/us30/n949 ), .A3(\AES_ENC/us30/n948 ), .A4(\AES_ENC/us30/n947 ), .ZN(\AES_ENC/us30/n951 ) );
NOR4_X2 \AES_ENC/us30/U162  ( .A1(\AES_ENC/us30/n896 ), .A2(\AES_ENC/us30/n895 ), .A3(\AES_ENC/us30/n894 ), .A4(\AES_ENC/us30/n893 ), .ZN(\AES_ENC/us30/n897 ) );
NOR2_X2 \AES_ENC/us30/U161  ( .A1(\AES_ENC/us30/n866 ), .A2(\AES_ENC/us30/n865 ), .ZN(\AES_ENC/us30/n872 ) );
NOR4_X2 \AES_ENC/us30/U160  ( .A1(\AES_ENC/us30/n870 ), .A2(\AES_ENC/us30/n869 ), .A3(\AES_ENC/us30/n868 ), .A4(\AES_ENC/us30/n867 ), .ZN(\AES_ENC/us30/n871 ) );
NOR4_X2 \AES_ENC/us30/U159  ( .A1(\AES_ENC/us30/n983 ), .A2(\AES_ENC/us30/n982 ), .A3(\AES_ENC/us30/n981 ), .A4(\AES_ENC/us30/n980 ), .ZN(\AES_ENC/us30/n984 ) );
NOR2_X2 \AES_ENC/us30/U158  ( .A1(\AES_ENC/us30/n979 ), .A2(\AES_ENC/us30/n978 ), .ZN(\AES_ENC/us30/n985 ) );
NOR4_X2 \AES_ENC/us30/U157  ( .A1(\AES_ENC/us30/n1125 ), .A2(\AES_ENC/us30/n1124 ), .A3(\AES_ENC/us30/n1123 ), .A4(\AES_ENC/us30/n1122 ), .ZN(\AES_ENC/us30/n1126 ) );
NOR4_X2 \AES_ENC/us30/U156  ( .A1(\AES_ENC/us30/n1084 ), .A2(\AES_ENC/us30/n1083 ), .A3(\AES_ENC/us30/n1082 ), .A4(\AES_ENC/us30/n1081 ), .ZN(\AES_ENC/us30/n1085 ) );
NOR2_X2 \AES_ENC/us30/U155  ( .A1(\AES_ENC/us30/n1076 ), .A2(\AES_ENC/us30/n1075 ), .ZN(\AES_ENC/us30/n1086 ) );
NOR3_X2 \AES_ENC/us30/U154  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n1054 ), .A3(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n961 ) );
NOR3_X2 \AES_ENC/us30/U153  ( .A1(\AES_ENC/us30/n620 ), .A2(\AES_ENC/us30/n1074 ), .A3(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n671 ) );
NOR2_X2 \AES_ENC/us30/U152  ( .A1(\AES_ENC/us30/n1057 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n1062 ) );
NOR2_X2 \AES_ENC/us30/U143  ( .A1(\AES_ENC/us30/n1055 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n1063 ) );
NOR2_X2 \AES_ENC/us30/U142  ( .A1(\AES_ENC/us30/n1060 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n1061 ) );
NOR4_X2 \AES_ENC/us30/U141  ( .A1(\AES_ENC/us30/n1064 ), .A2(\AES_ENC/us30/n1063 ), .A3(\AES_ENC/us30/n1062 ), .A4(\AES_ENC/us30/n1061 ), .ZN(\AES_ENC/us30/n1065 ) );
NOR3_X2 \AES_ENC/us30/U140  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n1120 ), .A3(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n918 ) );
NOR3_X2 \AES_ENC/us30/U132  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n573 ), .A3(\AES_ENC/us30/n1013 ), .ZN(\AES_ENC/us30/n917 ) );
NOR2_X2 \AES_ENC/us30/U131  ( .A1(\AES_ENC/us30/n914 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n915 ) );
NOR4_X2 \AES_ENC/us30/U130  ( .A1(\AES_ENC/us30/n918 ), .A2(\AES_ENC/us30/n917 ), .A3(\AES_ENC/us30/n916 ), .A4(\AES_ENC/us30/n915 ), .ZN(\AES_ENC/us30/n919 ) );
NOR2_X2 \AES_ENC/us30/U129  ( .A1(\AES_ENC/us30/n616 ), .A2(\AES_ENC/us30/n580 ), .ZN(\AES_ENC/us30/n771 ) );
NOR2_X2 \AES_ENC/us30/U128  ( .A1(\AES_ENC/us30/n1103 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n772 ) );
NOR2_X2 \AES_ENC/us30/U127  ( .A1(\AES_ENC/us30/n610 ), .A2(\AES_ENC/us30/n599 ), .ZN(\AES_ENC/us30/n773 ) );
NOR4_X2 \AES_ENC/us30/U126  ( .A1(\AES_ENC/us30/n773 ), .A2(\AES_ENC/us30/n772 ), .A3(\AES_ENC/us30/n771 ), .A4(\AES_ENC/us30/n770 ), .ZN(\AES_ENC/us30/n774 ) );
NOR2_X2 \AES_ENC/us30/U121  ( .A1(\AES_ENC/us30/n735 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n687 ) );
NOR2_X2 \AES_ENC/us30/U120  ( .A1(\AES_ENC/us30/n684 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n688 ) );
NOR2_X2 \AES_ENC/us30/U119  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n600 ), .ZN(\AES_ENC/us30/n686 ) );
NOR4_X2 \AES_ENC/us30/U118  ( .A1(\AES_ENC/us30/n688 ), .A2(\AES_ENC/us30/n687 ), .A3(\AES_ENC/us30/n686 ), .A4(\AES_ENC/us30/n685 ), .ZN(\AES_ENC/us30/n689 ) );
NOR2_X2 \AES_ENC/us30/U117  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n595 ), .ZN(\AES_ENC/us30/n858 ) );
NOR2_X2 \AES_ENC/us30/U116  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n855 ), .ZN(\AES_ENC/us30/n857 ) );
NOR2_X2 \AES_ENC/us30/U115  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n587 ), .ZN(\AES_ENC/us30/n856 ) );
NOR4_X2 \AES_ENC/us30/U106  ( .A1(\AES_ENC/us30/n858 ), .A2(\AES_ENC/us30/n857 ), .A3(\AES_ENC/us30/n856 ), .A4(\AES_ENC/us30/n958 ), .ZN(\AES_ENC/us30/n859 ) );
NOR2_X2 \AES_ENC/us30/U105  ( .A1(\AES_ENC/us30/n780 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n784 ) );
NOR2_X2 \AES_ENC/us30/U104  ( .A1(\AES_ENC/us30/n1117 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n782 ) );
NOR2_X2 \AES_ENC/us30/U103  ( .A1(\AES_ENC/us30/n781 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n783 ) );
NOR4_X2 \AES_ENC/us30/U102  ( .A1(\AES_ENC/us30/n880 ), .A2(\AES_ENC/us30/n784 ), .A3(\AES_ENC/us30/n783 ), .A4(\AES_ENC/us30/n782 ), .ZN(\AES_ENC/us30/n785 ) );
NOR2_X2 \AES_ENC/us30/U101  ( .A1(\AES_ENC/us30/n583 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n814 ) );
NOR2_X2 \AES_ENC/us30/U100  ( .A1(\AES_ENC/us30/n907 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n813 ) );
NOR3_X2 \AES_ENC/us30/U95  ( .A1(\AES_ENC/us30/n606 ), .A2(\AES_ENC/us30/n1058 ), .A3(\AES_ENC/us30/n1059 ), .ZN(\AES_ENC/us30/n815 ) );
NOR4_X2 \AES_ENC/us30/U94  ( .A1(\AES_ENC/us30/n815 ), .A2(\AES_ENC/us30/n814 ), .A3(\AES_ENC/us30/n813 ), .A4(\AES_ENC/us30/n812 ), .ZN(\AES_ENC/us30/n816 ) );
NOR2_X2 \AES_ENC/us30/U93  ( .A1(\AES_ENC/us30/n617 ), .A2(\AES_ENC/us30/n569 ), .ZN(\AES_ENC/us30/n721 ) );
NOR2_X2 \AES_ENC/us30/U92  ( .A1(\AES_ENC/us30/n1031 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n723 ) );
NOR2_X2 \AES_ENC/us30/U91  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n1096 ), .ZN(\AES_ENC/us30/n722 ) );
NOR4_X2 \AES_ENC/us30/U90  ( .A1(\AES_ENC/us30/n724 ), .A2(\AES_ENC/us30/n723 ), .A3(\AES_ENC/us30/n722 ), .A4(\AES_ENC/us30/n721 ), .ZN(\AES_ENC/us30/n725 ) );
NOR2_X2 \AES_ENC/us30/U89  ( .A1(\AES_ENC/us30/n911 ), .A2(\AES_ENC/us30/n990 ), .ZN(\AES_ENC/us30/n1009 ) );
NOR2_X2 \AES_ENC/us30/U88  ( .A1(\AES_ENC/us30/n1013 ), .A2(\AES_ENC/us30/n573 ), .ZN(\AES_ENC/us30/n1014 ) );
NOR2_X2 \AES_ENC/us30/U87  ( .A1(\AES_ENC/us30/n1014 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n1015 ) );
NOR4_X2 \AES_ENC/us30/U86  ( .A1(\AES_ENC/us30/n1016 ), .A2(\AES_ENC/us30/n1015 ), .A3(\AES_ENC/us30/n1119 ), .A4(\AES_ENC/us30/n1046 ), .ZN(\AES_ENC/us30/n1017 ) );
NOR2_X2 \AES_ENC/us30/U81  ( .A1(\AES_ENC/us30/n996 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n998 ) );
NOR2_X2 \AES_ENC/us30/U80  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n577 ), .ZN(\AES_ENC/us30/n1000 ) );
NOR2_X2 \AES_ENC/us30/U79  ( .A1(\AES_ENC/us30/n616 ), .A2(\AES_ENC/us30/n1096 ), .ZN(\AES_ENC/us30/n999 ) );
NOR4_X2 \AES_ENC/us30/U78  ( .A1(\AES_ENC/us30/n1000 ), .A2(\AES_ENC/us30/n999 ), .A3(\AES_ENC/us30/n998 ), .A4(\AES_ENC/us30/n997 ), .ZN(\AES_ENC/us30/n1001 ) );
NOR2_X2 \AES_ENC/us30/U74  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n1096 ), .ZN(\AES_ENC/us30/n697 ) );
NOR2_X2 \AES_ENC/us30/U73  ( .A1(\AES_ENC/us30/n620 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n958 ) );
NOR2_X2 \AES_ENC/us30/U72  ( .A1(\AES_ENC/us30/n911 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n983 ) );
NOR2_X2 \AES_ENC/us30/U71  ( .A1(\AES_ENC/us30/n1054 ), .A2(\AES_ENC/us30/n1103 ), .ZN(\AES_ENC/us30/n1031 ) );
INV_X4 \AES_ENC/us30/U65  ( .A(\AES_ENC/us30/n1050 ), .ZN(\AES_ENC/us30/n612 ) );
INV_X4 \AES_ENC/us30/U64  ( .A(\AES_ENC/us30/n1072 ), .ZN(\AES_ENC/us30/n605 ) );
INV_X4 \AES_ENC/us30/U63  ( .A(\AES_ENC/us30/n1073 ), .ZN(\AES_ENC/us30/n604 ) );
NOR2_X2 \AES_ENC/us30/U62  ( .A1(\AES_ENC/us30/n582 ), .A2(\AES_ENC/us30/n613 ), .ZN(\AES_ENC/us30/n880 ) );
NOR3_X2 \AES_ENC/us30/U61  ( .A1(\AES_ENC/us30/n826 ), .A2(\AES_ENC/us30/n1121 ), .A3(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n946 ) );
INV_X4 \AES_ENC/us30/U59  ( .A(\AES_ENC/us30/n1010 ), .ZN(\AES_ENC/us30/n608 ) );
NOR3_X2 \AES_ENC/us30/U58  ( .A1(\AES_ENC/us30/n573 ), .A2(\AES_ENC/us30/n1029 ), .A3(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n1119 ) );
INV_X4 \AES_ENC/us30/U57  ( .A(\AES_ENC/us30/n956 ), .ZN(\AES_ENC/us30/n615 ) );
NOR2_X2 \AES_ENC/us30/U50  ( .A1(\AES_ENC/us30/n623 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n1013 ) );
NOR2_X2 \AES_ENC/us30/U49  ( .A1(\AES_ENC/us30/n620 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n910 ) );
NOR2_X2 \AES_ENC/us30/U48  ( .A1(\AES_ENC/us30/n569 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n1091 ) );
NOR2_X2 \AES_ENC/us30/U47  ( .A1(\AES_ENC/us30/n622 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n990 ) );
NOR2_X2 \AES_ENC/us30/U46  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/us30/n1121 ), .ZN(\AES_ENC/us30/n996 ) );
NOR2_X2 \AES_ENC/us30/U45  ( .A1(\AES_ENC/us30/n610 ), .A2(\AES_ENC/us30/n600 ), .ZN(\AES_ENC/us30/n628 ) );
NOR2_X2 \AES_ENC/us30/U44  ( .A1(\AES_ENC/us30/n576 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n866 ) );
NOR2_X2 \AES_ENC/us30/U43  ( .A1(\AES_ENC/us30/n603 ), .A2(\AES_ENC/us30/n610 ), .ZN(\AES_ENC/us30/n1006 ) );
NOR2_X2 \AES_ENC/us30/U42  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n1117 ), .ZN(\AES_ENC/us30/n1118 ) );
NOR2_X2 \AES_ENC/us30/U41  ( .A1(\AES_ENC/us30/n1119 ), .A2(\AES_ENC/us30/n1118 ), .ZN(\AES_ENC/us30/n1127 ) );
NOR2_X2 \AES_ENC/us30/U36  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n906 ), .ZN(\AES_ENC/us30/n909 ) );
NOR2_X2 \AES_ENC/us30/U35  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n594 ), .ZN(\AES_ENC/us30/n629 ) );
NOR2_X2 \AES_ENC/us30/U34  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n597 ), .ZN(\AES_ENC/us30/n658 ) );
NOR2_X2 \AES_ENC/us30/U33  ( .A1(\AES_ENC/us30/n1116 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n695 ) );
NOR2_X2 \AES_ENC/us30/U32  ( .A1(\AES_ENC/us30/n1078 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n1083 ) );
NOR2_X2 \AES_ENC/us30/U31  ( .A1(\AES_ENC/us30/n941 ), .A2(\AES_ENC/us30/n608 ), .ZN(\AES_ENC/us30/n724 ) );
NOR2_X2 \AES_ENC/us30/U30  ( .A1(\AES_ENC/us30/n598 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n1107 ) );
NOR2_X2 \AES_ENC/us30/U29  ( .A1(\AES_ENC/us30/n576 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n840 ) );
NOR2_X2 \AES_ENC/us30/U24  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n593 ), .ZN(\AES_ENC/us30/n633 ) );
NOR2_X2 \AES_ENC/us30/U23  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n1080 ), .ZN(\AES_ENC/us30/n1081 ) );
NOR2_X2 \AES_ENC/us30/U21  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n1045 ), .ZN(\AES_ENC/us30/n812 ) );
NOR2_X2 \AES_ENC/us30/U20  ( .A1(\AES_ENC/us30/n1009 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n960 ) );
NOR2_X2 \AES_ENC/us30/U19  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n601 ), .ZN(\AES_ENC/us30/n982 ) );
NOR2_X2 \AES_ENC/us30/U18  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n594 ), .ZN(\AES_ENC/us30/n757 ) );
NOR2_X2 \AES_ENC/us30/U17  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n590 ), .ZN(\AES_ENC/us30/n698 ) );
NOR2_X2 \AES_ENC/us30/U16  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n619 ), .ZN(\AES_ENC/us30/n708 ) );
NOR2_X2 \AES_ENC/us30/U15  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n582 ), .ZN(\AES_ENC/us30/n770 ) );
NOR2_X2 \AES_ENC/us30/U10  ( .A1(\AES_ENC/us30/n619 ), .A2(\AES_ENC/us30/n604 ), .ZN(\AES_ENC/us30/n803 ) );
NOR2_X2 \AES_ENC/us30/U9  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n881 ), .ZN(\AES_ENC/us30/n711 ) );
NOR2_X2 \AES_ENC/us30/U8  ( .A1(\AES_ENC/us30/n615 ), .A2(\AES_ENC/us30/n582 ), .ZN(\AES_ENC/us30/n867 ) );
NOR2_X2 \AES_ENC/us30/U7  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n599 ), .ZN(\AES_ENC/us30/n804 ) );
NOR2_X2 \AES_ENC/us30/U6  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n620 ), .ZN(\AES_ENC/us30/n1046 ) );
OR2_X4 \AES_ENC/us30/U5  ( .A1(\AES_ENC/us30/n624 ), .A2(\AES_ENC/sa30 [1]),.ZN(\AES_ENC/us30/n570 ) );
OR2_X4 \AES_ENC/us30/U4  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/sa30 [4]),.ZN(\AES_ENC/us30/n569 ) );
NAND2_X2 \AES_ENC/us30/U514  ( .A1(\AES_ENC/us30/n1121 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n1030 ) );
AND2_X2 \AES_ENC/us30/U513  ( .A1(\AES_ENC/us30/n597 ), .A2(\AES_ENC/us30/n1030 ), .ZN(\AES_ENC/us30/n1049 ) );
NAND2_X2 \AES_ENC/us30/U511  ( .A1(\AES_ENC/us30/n1049 ), .A2(\AES_ENC/us30/n794 ), .ZN(\AES_ENC/us30/n637 ) );
AND2_X2 \AES_ENC/us30/U493  ( .A1(\AES_ENC/us30/n779 ), .A2(\AES_ENC/us30/n996 ), .ZN(\AES_ENC/us30/n632 ) );
NAND4_X2 \AES_ENC/us30/U485  ( .A1(\AES_ENC/us30/n637 ), .A2(\AES_ENC/us30/n636 ), .A3(\AES_ENC/us30/n635 ), .A4(\AES_ENC/us30/n634 ), .ZN(\AES_ENC/us30/n638 ) );
NAND2_X2 \AES_ENC/us30/U484  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n638 ), .ZN(\AES_ENC/us30/n679 ) );
NAND2_X2 \AES_ENC/us30/U481  ( .A1(\AES_ENC/us30/n1094 ), .A2(\AES_ENC/us30/n591 ), .ZN(\AES_ENC/us30/n648 ) );
NAND2_X2 \AES_ENC/us30/U476  ( .A1(\AES_ENC/us30/n601 ), .A2(\AES_ENC/us30/n590 ), .ZN(\AES_ENC/us30/n762 ) );
NAND2_X2 \AES_ENC/us30/U475  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n762 ), .ZN(\AES_ENC/us30/n647 ) );
NAND4_X2 \AES_ENC/us30/U457  ( .A1(\AES_ENC/us30/n648 ), .A2(\AES_ENC/us30/n647 ), .A3(\AES_ENC/us30/n646 ), .A4(\AES_ENC/us30/n645 ), .ZN(\AES_ENC/us30/n649 ) );
NAND2_X2 \AES_ENC/us30/U456  ( .A1(\AES_ENC/sa30 [0]), .A2(\AES_ENC/us30/n649 ), .ZN(\AES_ENC/us30/n665 ) );
NAND2_X2 \AES_ENC/us30/U454  ( .A1(\AES_ENC/us30/n596 ), .A2(\AES_ENC/us30/n623 ), .ZN(\AES_ENC/us30/n855 ) );
NAND2_X2 \AES_ENC/us30/U453  ( .A1(\AES_ENC/us30/n587 ), .A2(\AES_ENC/us30/n855 ), .ZN(\AES_ENC/us30/n821 ) );
NAND2_X2 \AES_ENC/us30/U452  ( .A1(\AES_ENC/us30/n1093 ), .A2(\AES_ENC/us30/n821 ), .ZN(\AES_ENC/us30/n662 ) );
NAND2_X2 \AES_ENC/us30/U451  ( .A1(\AES_ENC/us30/n619 ), .A2(\AES_ENC/us30/n589 ), .ZN(\AES_ENC/us30/n650 ) );
NAND2_X2 \AES_ENC/us30/U450  ( .A1(\AES_ENC/us30/n956 ), .A2(\AES_ENC/us30/n650 ), .ZN(\AES_ENC/us30/n661 ) );
NAND2_X2 \AES_ENC/us30/U449  ( .A1(\AES_ENC/us30/n626 ), .A2(\AES_ENC/us30/n627 ), .ZN(\AES_ENC/us30/n839 ) );
OR2_X2 \AES_ENC/us30/U446  ( .A1(\AES_ENC/us30/n839 ), .A2(\AES_ENC/us30/n932 ), .ZN(\AES_ENC/us30/n656 ) );
NAND2_X2 \AES_ENC/us30/U445  ( .A1(\AES_ENC/us30/n621 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n1096 ) );
NAND2_X2 \AES_ENC/us30/U444  ( .A1(\AES_ENC/us30/n1030 ), .A2(\AES_ENC/us30/n1096 ), .ZN(\AES_ENC/us30/n651 ) );
NAND2_X2 \AES_ENC/us30/U443  ( .A1(\AES_ENC/us30/n1114 ), .A2(\AES_ENC/us30/n651 ), .ZN(\AES_ENC/us30/n655 ) );
OR3_X2 \AES_ENC/us30/U440  ( .A1(\AES_ENC/us30/n1079 ), .A2(\AES_ENC/sa30 [7]), .A3(\AES_ENC/us30/n626 ), .ZN(\AES_ENC/us30/n654 ));
NAND2_X2 \AES_ENC/us30/U439  ( .A1(\AES_ENC/us30/n593 ), .A2(\AES_ENC/us30/n601 ), .ZN(\AES_ENC/us30/n652 ) );
NAND4_X2 \AES_ENC/us30/U437  ( .A1(\AES_ENC/us30/n656 ), .A2(\AES_ENC/us30/n655 ), .A3(\AES_ENC/us30/n654 ), .A4(\AES_ENC/us30/n653 ), .ZN(\AES_ENC/us30/n657 ) );
NAND2_X2 \AES_ENC/us30/U436  ( .A1(\AES_ENC/sa30 [2]), .A2(\AES_ENC/us30/n657 ), .ZN(\AES_ENC/us30/n660 ) );
NAND4_X2 \AES_ENC/us30/U432  ( .A1(\AES_ENC/us30/n662 ), .A2(\AES_ENC/us30/n661 ), .A3(\AES_ENC/us30/n660 ), .A4(\AES_ENC/us30/n659 ), .ZN(\AES_ENC/us30/n663 ) );
NAND2_X2 \AES_ENC/us30/U431  ( .A1(\AES_ENC/us30/n663 ), .A2(\AES_ENC/us30/n574 ), .ZN(\AES_ENC/us30/n664 ) );
NAND2_X2 \AES_ENC/us30/U430  ( .A1(\AES_ENC/us30/n665 ), .A2(\AES_ENC/us30/n664 ), .ZN(\AES_ENC/us30/n666 ) );
NAND2_X2 \AES_ENC/us30/U429  ( .A1(\AES_ENC/sa30 [6]), .A2(\AES_ENC/us30/n666 ), .ZN(\AES_ENC/us30/n678 ) );
NAND2_X2 \AES_ENC/us30/U426  ( .A1(\AES_ENC/us30/n735 ), .A2(\AES_ENC/us30/n1093 ), .ZN(\AES_ENC/us30/n675 ) );
NAND2_X2 \AES_ENC/us30/U425  ( .A1(\AES_ENC/us30/n588 ), .A2(\AES_ENC/us30/n597 ), .ZN(\AES_ENC/us30/n1045 ) );
OR2_X2 \AES_ENC/us30/U424  ( .A1(\AES_ENC/us30/n1045 ), .A2(\AES_ENC/us30/n605 ), .ZN(\AES_ENC/us30/n674 ) );
NAND2_X2 \AES_ENC/us30/U423  ( .A1(\AES_ENC/sa30 [1]), .A2(\AES_ENC/us30/n620 ), .ZN(\AES_ENC/us30/n667 ) );
NAND2_X2 \AES_ENC/us30/U422  ( .A1(\AES_ENC/us30/n619 ), .A2(\AES_ENC/us30/n667 ), .ZN(\AES_ENC/us30/n1071 ) );
NAND4_X2 \AES_ENC/us30/U412  ( .A1(\AES_ENC/us30/n675 ), .A2(\AES_ENC/us30/n674 ), .A3(\AES_ENC/us30/n673 ), .A4(\AES_ENC/us30/n672 ), .ZN(\AES_ENC/us30/n676 ) );
NAND2_X2 \AES_ENC/us30/U411  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n676 ), .ZN(\AES_ENC/us30/n677 ) );
NAND2_X2 \AES_ENC/us30/U408  ( .A1(\AES_ENC/us30/n800 ), .A2(\AES_ENC/us30/n1022 ), .ZN(\AES_ENC/us30/n680 ) );
NAND2_X2 \AES_ENC/us30/U407  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n680 ), .ZN(\AES_ENC/us30/n681 ) );
AND2_X2 \AES_ENC/us30/U402  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n684 ), .ZN(\AES_ENC/us30/n682 ) );
NAND4_X2 \AES_ENC/us30/U395  ( .A1(\AES_ENC/us30/n691 ), .A2(\AES_ENC/us30/n581 ), .A3(\AES_ENC/us30/n690 ), .A4(\AES_ENC/us30/n689 ), .ZN(\AES_ENC/us30/n692 ) );
NAND2_X2 \AES_ENC/us30/U394  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n692 ), .ZN(\AES_ENC/us30/n733 ) );
NAND2_X2 \AES_ENC/us30/U392  ( .A1(\AES_ENC/us30/n977 ), .A2(\AES_ENC/us30/n1050 ), .ZN(\AES_ENC/us30/n702 ) );
NAND2_X2 \AES_ENC/us30/U391  ( .A1(\AES_ENC/us30/n1093 ), .A2(\AES_ENC/us30/n1045 ), .ZN(\AES_ENC/us30/n701 ) );
NAND4_X2 \AES_ENC/us30/U381  ( .A1(\AES_ENC/us30/n702 ), .A2(\AES_ENC/us30/n701 ), .A3(\AES_ENC/us30/n700 ), .A4(\AES_ENC/us30/n699 ), .ZN(\AES_ENC/us30/n703 ) );
NAND2_X2 \AES_ENC/us30/U380  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n703 ), .ZN(\AES_ENC/us30/n732 ) );
AND2_X2 \AES_ENC/us30/U379  ( .A1(\AES_ENC/sa30 [0]), .A2(\AES_ENC/sa30 [6]),.ZN(\AES_ENC/us30/n1113 ) );
NAND2_X2 \AES_ENC/us30/U378  ( .A1(\AES_ENC/us30/n601 ), .A2(\AES_ENC/us30/n1030 ), .ZN(\AES_ENC/us30/n881 ) );
NAND2_X2 \AES_ENC/us30/U377  ( .A1(\AES_ENC/us30/n1093 ), .A2(\AES_ENC/us30/n881 ), .ZN(\AES_ENC/us30/n715 ) );
NAND2_X2 \AES_ENC/us30/U376  ( .A1(\AES_ENC/us30/n1010 ), .A2(\AES_ENC/us30/n600 ), .ZN(\AES_ENC/us30/n714 ) );
NAND2_X2 \AES_ENC/us30/U375  ( .A1(\AES_ENC/us30/n855 ), .A2(\AES_ENC/us30/n588 ), .ZN(\AES_ENC/us30/n1117 ) );
XNOR2_X2 \AES_ENC/us30/U371  ( .A(\AES_ENC/us30/n611 ), .B(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n824 ) );
NAND4_X2 \AES_ENC/us30/U362  ( .A1(\AES_ENC/us30/n715 ), .A2(\AES_ENC/us30/n714 ), .A3(\AES_ENC/us30/n713 ), .A4(\AES_ENC/us30/n712 ), .ZN(\AES_ENC/us30/n716 ) );
NAND2_X2 \AES_ENC/us30/U361  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n716 ), .ZN(\AES_ENC/us30/n731 ) );
AND2_X2 \AES_ENC/us30/U360  ( .A1(\AES_ENC/sa30 [6]), .A2(\AES_ENC/us30/n574 ), .ZN(\AES_ENC/us30/n1131 ) );
NAND2_X2 \AES_ENC/us30/U359  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n717 ) );
NAND2_X2 \AES_ENC/us30/U358  ( .A1(\AES_ENC/us30/n1029 ), .A2(\AES_ENC/us30/n717 ), .ZN(\AES_ENC/us30/n728 ) );
NAND2_X2 \AES_ENC/us30/U357  ( .A1(\AES_ENC/sa30 [1]), .A2(\AES_ENC/us30/n624 ), .ZN(\AES_ENC/us30/n1097 ) );
NAND2_X2 \AES_ENC/us30/U356  ( .A1(\AES_ENC/us30/n603 ), .A2(\AES_ENC/us30/n1097 ), .ZN(\AES_ENC/us30/n718 ) );
NAND2_X2 \AES_ENC/us30/U355  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n718 ), .ZN(\AES_ENC/us30/n727 ) );
NAND4_X2 \AES_ENC/us30/U344  ( .A1(\AES_ENC/us30/n728 ), .A2(\AES_ENC/us30/n727 ), .A3(\AES_ENC/us30/n726 ), .A4(\AES_ENC/us30/n725 ), .ZN(\AES_ENC/us30/n729 ) );
NAND2_X2 \AES_ENC/us30/U343  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n729 ), .ZN(\AES_ENC/us30/n730 ) );
NAND4_X2 \AES_ENC/us30/U342  ( .A1(\AES_ENC/us30/n733 ), .A2(\AES_ENC/us30/n732 ), .A3(\AES_ENC/us30/n731 ), .A4(\AES_ENC/us30/n730 ), .ZN(\AES_ENC/sa30_sub[1] ) );
NAND2_X2 \AES_ENC/us30/U341  ( .A1(\AES_ENC/sa30 [7]), .A2(\AES_ENC/us30/n611 ), .ZN(\AES_ENC/us30/n734 ) );
NAND2_X2 \AES_ENC/us30/U340  ( .A1(\AES_ENC/us30/n734 ), .A2(\AES_ENC/us30/n607 ), .ZN(\AES_ENC/us30/n738 ) );
OR4_X2 \AES_ENC/us30/U339  ( .A1(\AES_ENC/us30/n738 ), .A2(\AES_ENC/us30/n626 ), .A3(\AES_ENC/us30/n826 ), .A4(\AES_ENC/us30/n1121 ), .ZN(\AES_ENC/us30/n746 ) );
NAND2_X2 \AES_ENC/us30/U337  ( .A1(\AES_ENC/us30/n1100 ), .A2(\AES_ENC/us30/n587 ), .ZN(\AES_ENC/us30/n992 ) );
OR2_X2 \AES_ENC/us30/U336  ( .A1(\AES_ENC/us30/n610 ), .A2(\AES_ENC/us30/n735 ), .ZN(\AES_ENC/us30/n737 ) );
NAND2_X2 \AES_ENC/us30/U334  ( .A1(\AES_ENC/us30/n619 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n753 ) );
NAND2_X2 \AES_ENC/us30/U333  ( .A1(\AES_ENC/us30/n582 ), .A2(\AES_ENC/us30/n753 ), .ZN(\AES_ENC/us30/n1080 ) );
NAND2_X2 \AES_ENC/us30/U332  ( .A1(\AES_ENC/us30/n1048 ), .A2(\AES_ENC/us30/n576 ), .ZN(\AES_ENC/us30/n736 ) );
NAND2_X2 \AES_ENC/us30/U331  ( .A1(\AES_ENC/us30/n737 ), .A2(\AES_ENC/us30/n736 ), .ZN(\AES_ENC/us30/n739 ) );
NAND2_X2 \AES_ENC/us30/U330  ( .A1(\AES_ENC/us30/n739 ), .A2(\AES_ENC/us30/n738 ), .ZN(\AES_ENC/us30/n745 ) );
NAND2_X2 \AES_ENC/us30/U326  ( .A1(\AES_ENC/us30/n1096 ), .A2(\AES_ENC/us30/n590 ), .ZN(\AES_ENC/us30/n906 ) );
NAND4_X2 \AES_ENC/us30/U323  ( .A1(\AES_ENC/us30/n746 ), .A2(\AES_ENC/us30/n992 ), .A3(\AES_ENC/us30/n745 ), .A4(\AES_ENC/us30/n744 ), .ZN(\AES_ENC/us30/n747 ) );
NAND2_X2 \AES_ENC/us30/U322  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n747 ), .ZN(\AES_ENC/us30/n793 ) );
NAND2_X2 \AES_ENC/us30/U321  ( .A1(\AES_ENC/us30/n584 ), .A2(\AES_ENC/us30/n855 ), .ZN(\AES_ENC/us30/n748 ) );
NAND2_X2 \AES_ENC/us30/U320  ( .A1(\AES_ENC/us30/n956 ), .A2(\AES_ENC/us30/n748 ), .ZN(\AES_ENC/us30/n760 ) );
NAND2_X2 \AES_ENC/us30/U313  ( .A1(\AES_ENC/us30/n590 ), .A2(\AES_ENC/us30/n753 ), .ZN(\AES_ENC/us30/n1023 ) );
NAND4_X2 \AES_ENC/us30/U308  ( .A1(\AES_ENC/us30/n760 ), .A2(\AES_ENC/us30/n992 ), .A3(\AES_ENC/us30/n759 ), .A4(\AES_ENC/us30/n758 ), .ZN(\AES_ENC/us30/n761 ) );
NAND2_X2 \AES_ENC/us30/U307  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n761 ), .ZN(\AES_ENC/us30/n792 ) );
NAND2_X2 \AES_ENC/us30/U306  ( .A1(\AES_ENC/us30/n584 ), .A2(\AES_ENC/us30/n603 ), .ZN(\AES_ENC/us30/n989 ) );
NAND2_X2 \AES_ENC/us30/U305  ( .A1(\AES_ENC/us30/n1050 ), .A2(\AES_ENC/us30/n989 ), .ZN(\AES_ENC/us30/n777 ) );
NAND2_X2 \AES_ENC/us30/U304  ( .A1(\AES_ENC/us30/n1093 ), .A2(\AES_ENC/us30/n762 ), .ZN(\AES_ENC/us30/n776 ) );
XNOR2_X2 \AES_ENC/us30/U301  ( .A(\AES_ENC/sa30 [7]), .B(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n959 ) );
NAND4_X2 \AES_ENC/us30/U289  ( .A1(\AES_ENC/us30/n777 ), .A2(\AES_ENC/us30/n776 ), .A3(\AES_ENC/us30/n775 ), .A4(\AES_ENC/us30/n774 ), .ZN(\AES_ENC/us30/n778 ) );
NAND2_X2 \AES_ENC/us30/U288  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n778 ), .ZN(\AES_ENC/us30/n791 ) );
NAND2_X2 \AES_ENC/us30/U287  ( .A1(\AES_ENC/us30/n1056 ), .A2(\AES_ENC/us30/n1050 ), .ZN(\AES_ENC/us30/n788 ) );
NAND2_X2 \AES_ENC/us30/U286  ( .A1(\AES_ENC/us30/n1091 ), .A2(\AES_ENC/us30/n779 ), .ZN(\AES_ENC/us30/n787 ) );
NAND2_X2 \AES_ENC/us30/U285  ( .A1(\AES_ENC/us30/n956 ), .A2(\AES_ENC/sa30 [1]), .ZN(\AES_ENC/us30/n786 ) );
NAND4_X2 \AES_ENC/us30/U278  ( .A1(\AES_ENC/us30/n788 ), .A2(\AES_ENC/us30/n787 ), .A3(\AES_ENC/us30/n786 ), .A4(\AES_ENC/us30/n785 ), .ZN(\AES_ENC/us30/n789 ) );
NAND2_X2 \AES_ENC/us30/U277  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n789 ), .ZN(\AES_ENC/us30/n790 ) );
NAND4_X2 \AES_ENC/us30/U276  ( .A1(\AES_ENC/us30/n793 ), .A2(\AES_ENC/us30/n792 ), .A3(\AES_ENC/us30/n791 ), .A4(\AES_ENC/us30/n790 ), .ZN(\AES_ENC/sa30_sub[2] ) );
NAND2_X2 \AES_ENC/us30/U275  ( .A1(\AES_ENC/us30/n1059 ), .A2(\AES_ENC/us30/n794 ), .ZN(\AES_ENC/us30/n810 ) );
NAND2_X2 \AES_ENC/us30/U274  ( .A1(\AES_ENC/us30/n1049 ), .A2(\AES_ENC/us30/n956 ), .ZN(\AES_ENC/us30/n809 ) );
OR2_X2 \AES_ENC/us30/U266  ( .A1(\AES_ENC/us30/n1096 ), .A2(\AES_ENC/us30/n606 ), .ZN(\AES_ENC/us30/n802 ) );
NAND2_X2 \AES_ENC/us30/U265  ( .A1(\AES_ENC/us30/n1053 ), .A2(\AES_ENC/us30/n800 ), .ZN(\AES_ENC/us30/n801 ) );
NAND2_X2 \AES_ENC/us30/U264  ( .A1(\AES_ENC/us30/n802 ), .A2(\AES_ENC/us30/n801 ), .ZN(\AES_ENC/us30/n805 ) );
NAND4_X2 \AES_ENC/us30/U261  ( .A1(\AES_ENC/us30/n810 ), .A2(\AES_ENC/us30/n809 ), .A3(\AES_ENC/us30/n808 ), .A4(\AES_ENC/us30/n807 ), .ZN(\AES_ENC/us30/n811 ) );
NAND2_X2 \AES_ENC/us30/U260  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n811 ), .ZN(\AES_ENC/us30/n852 ) );
OR2_X2 \AES_ENC/us30/U259  ( .A1(\AES_ENC/us30/n1023 ), .A2(\AES_ENC/us30/n617 ), .ZN(\AES_ENC/us30/n819 ) );
OR2_X2 \AES_ENC/us30/U257  ( .A1(\AES_ENC/us30/n570 ), .A2(\AES_ENC/us30/n930 ), .ZN(\AES_ENC/us30/n818 ) );
NAND2_X2 \AES_ENC/us30/U256  ( .A1(\AES_ENC/us30/n1013 ), .A2(\AES_ENC/us30/n1094 ), .ZN(\AES_ENC/us30/n817 ) );
NAND4_X2 \AES_ENC/us30/U249  ( .A1(\AES_ENC/us30/n819 ), .A2(\AES_ENC/us30/n818 ), .A3(\AES_ENC/us30/n817 ), .A4(\AES_ENC/us30/n816 ), .ZN(\AES_ENC/us30/n820 ) );
NAND2_X2 \AES_ENC/us30/U248  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n820 ), .ZN(\AES_ENC/us30/n851 ) );
NAND2_X2 \AES_ENC/us30/U247  ( .A1(\AES_ENC/us30/n956 ), .A2(\AES_ENC/us30/n1080 ), .ZN(\AES_ENC/us30/n835 ) );
NAND2_X2 \AES_ENC/us30/U246  ( .A1(\AES_ENC/us30/n570 ), .A2(\AES_ENC/us30/n1030 ), .ZN(\AES_ENC/us30/n1047 ) );
OR2_X2 \AES_ENC/us30/U245  ( .A1(\AES_ENC/us30/n1047 ), .A2(\AES_ENC/us30/n612 ), .ZN(\AES_ENC/us30/n834 ) );
NAND2_X2 \AES_ENC/us30/U244  ( .A1(\AES_ENC/us30/n1072 ), .A2(\AES_ENC/us30/n589 ), .ZN(\AES_ENC/us30/n833 ) );
NAND4_X2 \AES_ENC/us30/U233  ( .A1(\AES_ENC/us30/n835 ), .A2(\AES_ENC/us30/n834 ), .A3(\AES_ENC/us30/n833 ), .A4(\AES_ENC/us30/n832 ), .ZN(\AES_ENC/us30/n836 ) );
NAND2_X2 \AES_ENC/us30/U232  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n836 ), .ZN(\AES_ENC/us30/n850 ) );
NAND2_X2 \AES_ENC/us30/U231  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n623 ), .ZN(\AES_ENC/us30/n847 ) );
NAND2_X2 \AES_ENC/us30/U230  ( .A1(\AES_ENC/us30/n1050 ), .A2(\AES_ENC/us30/n1071 ), .ZN(\AES_ENC/us30/n846 ) );
OR2_X2 \AES_ENC/us30/U224  ( .A1(\AES_ENC/us30/n1053 ), .A2(\AES_ENC/us30/n911 ), .ZN(\AES_ENC/us30/n1077 ) );
NAND4_X2 \AES_ENC/us30/U220  ( .A1(\AES_ENC/us30/n847 ), .A2(\AES_ENC/us30/n846 ), .A3(\AES_ENC/us30/n845 ), .A4(\AES_ENC/us30/n844 ), .ZN(\AES_ENC/us30/n848 ) );
NAND2_X2 \AES_ENC/us30/U219  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n848 ), .ZN(\AES_ENC/us30/n849 ) );
NAND4_X2 \AES_ENC/us30/U218  ( .A1(\AES_ENC/us30/n852 ), .A2(\AES_ENC/us30/n851 ), .A3(\AES_ENC/us30/n850 ), .A4(\AES_ENC/us30/n849 ), .ZN(\AES_ENC/sa30_sub[3] ) );
NAND2_X2 \AES_ENC/us30/U216  ( .A1(\AES_ENC/us30/n1009 ), .A2(\AES_ENC/us30/n1072 ), .ZN(\AES_ENC/us30/n862 ) );
NAND2_X2 \AES_ENC/us30/U215  ( .A1(\AES_ENC/us30/n603 ), .A2(\AES_ENC/us30/n577 ), .ZN(\AES_ENC/us30/n853 ) );
NAND2_X2 \AES_ENC/us30/U214  ( .A1(\AES_ENC/us30/n1050 ), .A2(\AES_ENC/us30/n853 ), .ZN(\AES_ENC/us30/n861 ) );
NAND4_X2 \AES_ENC/us30/U206  ( .A1(\AES_ENC/us30/n862 ), .A2(\AES_ENC/us30/n861 ), .A3(\AES_ENC/us30/n860 ), .A4(\AES_ENC/us30/n859 ), .ZN(\AES_ENC/us30/n863 ) );
NAND2_X2 \AES_ENC/us30/U205  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n863 ), .ZN(\AES_ENC/us30/n905 ) );
NAND2_X2 \AES_ENC/us30/U204  ( .A1(\AES_ENC/us30/n1010 ), .A2(\AES_ENC/us30/n989 ), .ZN(\AES_ENC/us30/n874 ) );
NAND2_X2 \AES_ENC/us30/U203  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n610 ), .ZN(\AES_ENC/us30/n864 ) );
NAND2_X2 \AES_ENC/us30/U202  ( .A1(\AES_ENC/us30/n929 ), .A2(\AES_ENC/us30/n864 ), .ZN(\AES_ENC/us30/n873 ) );
NAND4_X2 \AES_ENC/us30/U193  ( .A1(\AES_ENC/us30/n874 ), .A2(\AES_ENC/us30/n873 ), .A3(\AES_ENC/us30/n872 ), .A4(\AES_ENC/us30/n871 ), .ZN(\AES_ENC/us30/n875 ) );
NAND2_X2 \AES_ENC/us30/U192  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n875 ), .ZN(\AES_ENC/us30/n904 ) );
NAND2_X2 \AES_ENC/us30/U191  ( .A1(\AES_ENC/us30/n583 ), .A2(\AES_ENC/us30/n1050 ), .ZN(\AES_ENC/us30/n889 ) );
NAND2_X2 \AES_ENC/us30/U190  ( .A1(\AES_ENC/us30/n1093 ), .A2(\AES_ENC/us30/n587 ), .ZN(\AES_ENC/us30/n876 ) );
NAND2_X2 \AES_ENC/us30/U189  ( .A1(\AES_ENC/us30/n604 ), .A2(\AES_ENC/us30/n876 ), .ZN(\AES_ENC/us30/n877 ) );
NAND2_X2 \AES_ENC/us30/U188  ( .A1(\AES_ENC/us30/n877 ), .A2(\AES_ENC/us30/n623 ), .ZN(\AES_ENC/us30/n888 ) );
NAND4_X2 \AES_ENC/us30/U179  ( .A1(\AES_ENC/us30/n889 ), .A2(\AES_ENC/us30/n888 ), .A3(\AES_ENC/us30/n887 ), .A4(\AES_ENC/us30/n886 ), .ZN(\AES_ENC/us30/n890 ) );
NAND2_X2 \AES_ENC/us30/U178  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n890 ), .ZN(\AES_ENC/us30/n903 ) );
OR2_X2 \AES_ENC/us30/U177  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n1059 ), .ZN(\AES_ENC/us30/n900 ) );
NAND2_X2 \AES_ENC/us30/U176  ( .A1(\AES_ENC/us30/n1073 ), .A2(\AES_ENC/us30/n1047 ), .ZN(\AES_ENC/us30/n899 ) );
NAND2_X2 \AES_ENC/us30/U175  ( .A1(\AES_ENC/us30/n1094 ), .A2(\AES_ENC/us30/n595 ), .ZN(\AES_ENC/us30/n898 ) );
NAND4_X2 \AES_ENC/us30/U167  ( .A1(\AES_ENC/us30/n900 ), .A2(\AES_ENC/us30/n899 ), .A3(\AES_ENC/us30/n898 ), .A4(\AES_ENC/us30/n897 ), .ZN(\AES_ENC/us30/n901 ) );
NAND2_X2 \AES_ENC/us30/U166  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n901 ), .ZN(\AES_ENC/us30/n902 ) );
NAND4_X2 \AES_ENC/us30/U165  ( .A1(\AES_ENC/us30/n905 ), .A2(\AES_ENC/us30/n904 ), .A3(\AES_ENC/us30/n903 ), .A4(\AES_ENC/us30/n902 ), .ZN(\AES_ENC/sa30_sub[4] ) );
NAND2_X2 \AES_ENC/us30/U164  ( .A1(\AES_ENC/us30/n1094 ), .A2(\AES_ENC/us30/n599 ), .ZN(\AES_ENC/us30/n922 ) );
NAND2_X2 \AES_ENC/us30/U163  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n989 ), .ZN(\AES_ENC/us30/n921 ) );
NAND4_X2 \AES_ENC/us30/U151  ( .A1(\AES_ENC/us30/n922 ), .A2(\AES_ENC/us30/n921 ), .A3(\AES_ENC/us30/n920 ), .A4(\AES_ENC/us30/n919 ), .ZN(\AES_ENC/us30/n923 ) );
NAND2_X2 \AES_ENC/us30/U150  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n923 ), .ZN(\AES_ENC/us30/n972 ) );
NAND2_X2 \AES_ENC/us30/U149  ( .A1(\AES_ENC/us30/n582 ), .A2(\AES_ENC/us30/n619 ), .ZN(\AES_ENC/us30/n924 ) );
NAND2_X2 \AES_ENC/us30/U148  ( .A1(\AES_ENC/us30/n1073 ), .A2(\AES_ENC/us30/n924 ), .ZN(\AES_ENC/us30/n939 ) );
NAND2_X2 \AES_ENC/us30/U147  ( .A1(\AES_ENC/us30/n926 ), .A2(\AES_ENC/us30/n925 ), .ZN(\AES_ENC/us30/n927 ) );
NAND2_X2 \AES_ENC/us30/U146  ( .A1(\AES_ENC/us30/n606 ), .A2(\AES_ENC/us30/n927 ), .ZN(\AES_ENC/us30/n928 ) );
NAND2_X2 \AES_ENC/us30/U145  ( .A1(\AES_ENC/us30/n928 ), .A2(\AES_ENC/us30/n1080 ), .ZN(\AES_ENC/us30/n938 ) );
OR2_X2 \AES_ENC/us30/U144  ( .A1(\AES_ENC/us30/n1117 ), .A2(\AES_ENC/us30/n615 ), .ZN(\AES_ENC/us30/n937 ) );
NAND4_X2 \AES_ENC/us30/U139  ( .A1(\AES_ENC/us30/n939 ), .A2(\AES_ENC/us30/n938 ), .A3(\AES_ENC/us30/n937 ), .A4(\AES_ENC/us30/n936 ), .ZN(\AES_ENC/us30/n940 ) );
NAND2_X2 \AES_ENC/us30/U138  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n940 ), .ZN(\AES_ENC/us30/n971 ) );
OR2_X2 \AES_ENC/us30/U137  ( .A1(\AES_ENC/us30/n605 ), .A2(\AES_ENC/us30/n941 ), .ZN(\AES_ENC/us30/n954 ) );
NAND2_X2 \AES_ENC/us30/U136  ( .A1(\AES_ENC/us30/n1096 ), .A2(\AES_ENC/us30/n577 ), .ZN(\AES_ENC/us30/n942 ) );
NAND2_X2 \AES_ENC/us30/U135  ( .A1(\AES_ENC/us30/n1048 ), .A2(\AES_ENC/us30/n942 ), .ZN(\AES_ENC/us30/n943 ) );
NAND2_X2 \AES_ENC/us30/U134  ( .A1(\AES_ENC/us30/n612 ), .A2(\AES_ENC/us30/n943 ), .ZN(\AES_ENC/us30/n944 ) );
NAND2_X2 \AES_ENC/us30/U133  ( .A1(\AES_ENC/us30/n944 ), .A2(\AES_ENC/us30/n580 ), .ZN(\AES_ENC/us30/n953 ) );
NAND4_X2 \AES_ENC/us30/U125  ( .A1(\AES_ENC/us30/n954 ), .A2(\AES_ENC/us30/n953 ), .A3(\AES_ENC/us30/n952 ), .A4(\AES_ENC/us30/n951 ), .ZN(\AES_ENC/us30/n955 ) );
NAND2_X2 \AES_ENC/us30/U124  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n955 ), .ZN(\AES_ENC/us30/n970 ) );
NAND2_X2 \AES_ENC/us30/U123  ( .A1(\AES_ENC/us30/n1094 ), .A2(\AES_ENC/us30/n1071 ), .ZN(\AES_ENC/us30/n967 ) );
NAND2_X2 \AES_ENC/us30/U122  ( .A1(\AES_ENC/us30/n956 ), .A2(\AES_ENC/us30/n1030 ), .ZN(\AES_ENC/us30/n966 ) );
NAND4_X2 \AES_ENC/us30/U114  ( .A1(\AES_ENC/us30/n967 ), .A2(\AES_ENC/us30/n966 ), .A3(\AES_ENC/us30/n965 ), .A4(\AES_ENC/us30/n964 ), .ZN(\AES_ENC/us30/n968 ) );
NAND2_X2 \AES_ENC/us30/U113  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n968 ), .ZN(\AES_ENC/us30/n969 ) );
NAND4_X2 \AES_ENC/us30/U112  ( .A1(\AES_ENC/us30/n972 ), .A2(\AES_ENC/us30/n971 ), .A3(\AES_ENC/us30/n970 ), .A4(\AES_ENC/us30/n969 ), .ZN(\AES_ENC/sa30_sub[5] ) );
NAND2_X2 \AES_ENC/us30/U111  ( .A1(\AES_ENC/us30/n570 ), .A2(\AES_ENC/us30/n1097 ), .ZN(\AES_ENC/us30/n973 ) );
NAND2_X2 \AES_ENC/us30/U110  ( .A1(\AES_ENC/us30/n1073 ), .A2(\AES_ENC/us30/n973 ), .ZN(\AES_ENC/us30/n987 ) );
NAND2_X2 \AES_ENC/us30/U109  ( .A1(\AES_ENC/us30/n974 ), .A2(\AES_ENC/us30/n1077 ), .ZN(\AES_ENC/us30/n975 ) );
NAND2_X2 \AES_ENC/us30/U108  ( .A1(\AES_ENC/us30/n613 ), .A2(\AES_ENC/us30/n975 ), .ZN(\AES_ENC/us30/n976 ) );
NAND2_X2 \AES_ENC/us30/U107  ( .A1(\AES_ENC/us30/n977 ), .A2(\AES_ENC/us30/n976 ), .ZN(\AES_ENC/us30/n986 ) );
NAND4_X2 \AES_ENC/us30/U99  ( .A1(\AES_ENC/us30/n987 ), .A2(\AES_ENC/us30/n986 ), .A3(\AES_ENC/us30/n985 ), .A4(\AES_ENC/us30/n984 ), .ZN(\AES_ENC/us30/n988 ) );
NAND2_X2 \AES_ENC/us30/U98  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n988 ), .ZN(\AES_ENC/us30/n1044 ) );
NAND2_X2 \AES_ENC/us30/U97  ( .A1(\AES_ENC/us30/n1073 ), .A2(\AES_ENC/us30/n989 ), .ZN(\AES_ENC/us30/n1004 ) );
NAND2_X2 \AES_ENC/us30/U96  ( .A1(\AES_ENC/us30/n1092 ), .A2(\AES_ENC/us30/n619 ), .ZN(\AES_ENC/us30/n1003 ) );
NAND4_X2 \AES_ENC/us30/U85  ( .A1(\AES_ENC/us30/n1004 ), .A2(\AES_ENC/us30/n1003 ), .A3(\AES_ENC/us30/n1002 ), .A4(\AES_ENC/us30/n1001 ), .ZN(\AES_ENC/us30/n1005 ) );
NAND2_X2 \AES_ENC/us30/U84  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n1005 ), .ZN(\AES_ENC/us30/n1043 ) );
NAND2_X2 \AES_ENC/us30/U83  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n596 ), .ZN(\AES_ENC/us30/n1020 ) );
NAND2_X2 \AES_ENC/us30/U82  ( .A1(\AES_ENC/us30/n1050 ), .A2(\AES_ENC/us30/n624 ), .ZN(\AES_ENC/us30/n1019 ) );
NAND2_X2 \AES_ENC/us30/U77  ( .A1(\AES_ENC/us30/n1059 ), .A2(\AES_ENC/us30/n1114 ), .ZN(\AES_ENC/us30/n1012 ) );
NAND2_X2 \AES_ENC/us30/U76  ( .A1(\AES_ENC/us30/n1010 ), .A2(\AES_ENC/us30/n592 ), .ZN(\AES_ENC/us30/n1011 ) );
NAND2_X2 \AES_ENC/us30/U75  ( .A1(\AES_ENC/us30/n1012 ), .A2(\AES_ENC/us30/n1011 ), .ZN(\AES_ENC/us30/n1016 ) );
NAND4_X2 \AES_ENC/us30/U70  ( .A1(\AES_ENC/us30/n1020 ), .A2(\AES_ENC/us30/n1019 ), .A3(\AES_ENC/us30/n1018 ), .A4(\AES_ENC/us30/n1017 ), .ZN(\AES_ENC/us30/n1021 ) );
NAND2_X2 \AES_ENC/us30/U69  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n1021 ), .ZN(\AES_ENC/us30/n1042 ) );
NAND2_X2 \AES_ENC/us30/U68  ( .A1(\AES_ENC/us30/n1022 ), .A2(\AES_ENC/us30/n1093 ), .ZN(\AES_ENC/us30/n1039 ) );
NAND2_X2 \AES_ENC/us30/U67  ( .A1(\AES_ENC/us30/n1050 ), .A2(\AES_ENC/us30/n1023 ), .ZN(\AES_ENC/us30/n1038 ) );
NAND2_X2 \AES_ENC/us30/U66  ( .A1(\AES_ENC/us30/n1024 ), .A2(\AES_ENC/us30/n1071 ), .ZN(\AES_ENC/us30/n1037 ) );
AND2_X2 \AES_ENC/us30/U60  ( .A1(\AES_ENC/us30/n1030 ), .A2(\AES_ENC/us30/n602 ), .ZN(\AES_ENC/us30/n1078 ) );
NAND4_X2 \AES_ENC/us30/U56  ( .A1(\AES_ENC/us30/n1039 ), .A2(\AES_ENC/us30/n1038 ), .A3(\AES_ENC/us30/n1037 ), .A4(\AES_ENC/us30/n1036 ), .ZN(\AES_ENC/us30/n1040 ) );
NAND2_X2 \AES_ENC/us30/U55  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n1040 ), .ZN(\AES_ENC/us30/n1041 ) );
NAND4_X2 \AES_ENC/us30/U54  ( .A1(\AES_ENC/us30/n1044 ), .A2(\AES_ENC/us30/n1043 ), .A3(\AES_ENC/us30/n1042 ), .A4(\AES_ENC/us30/n1041 ), .ZN(\AES_ENC/sa30_sub[6] ) );
NAND2_X2 \AES_ENC/us30/U53  ( .A1(\AES_ENC/us30/n1072 ), .A2(\AES_ENC/us30/n1045 ), .ZN(\AES_ENC/us30/n1068 ) );
NAND2_X2 \AES_ENC/us30/U52  ( .A1(\AES_ENC/us30/n1046 ), .A2(\AES_ENC/us30/n582 ), .ZN(\AES_ENC/us30/n1067 ) );
NAND2_X2 \AES_ENC/us30/U51  ( .A1(\AES_ENC/us30/n1094 ), .A2(\AES_ENC/us30/n1047 ), .ZN(\AES_ENC/us30/n1066 ) );
NAND4_X2 \AES_ENC/us30/U40  ( .A1(\AES_ENC/us30/n1068 ), .A2(\AES_ENC/us30/n1067 ), .A3(\AES_ENC/us30/n1066 ), .A4(\AES_ENC/us30/n1065 ), .ZN(\AES_ENC/us30/n1069 ) );
NAND2_X2 \AES_ENC/us30/U39  ( .A1(\AES_ENC/us30/n1070 ), .A2(\AES_ENC/us30/n1069 ), .ZN(\AES_ENC/us30/n1135 ) );
NAND2_X2 \AES_ENC/us30/U38  ( .A1(\AES_ENC/us30/n1072 ), .A2(\AES_ENC/us30/n1071 ), .ZN(\AES_ENC/us30/n1088 ) );
NAND2_X2 \AES_ENC/us30/U37  ( .A1(\AES_ENC/us30/n1073 ), .A2(\AES_ENC/us30/n595 ), .ZN(\AES_ENC/us30/n1087 ) );
NAND4_X2 \AES_ENC/us30/U28  ( .A1(\AES_ENC/us30/n1088 ), .A2(\AES_ENC/us30/n1087 ), .A3(\AES_ENC/us30/n1086 ), .A4(\AES_ENC/us30/n1085 ), .ZN(\AES_ENC/us30/n1089 ) );
NAND2_X2 \AES_ENC/us30/U27  ( .A1(\AES_ENC/us30/n1090 ), .A2(\AES_ENC/us30/n1089 ), .ZN(\AES_ENC/us30/n1134 ) );
NAND2_X2 \AES_ENC/us30/U26  ( .A1(\AES_ENC/us30/n1091 ), .A2(\AES_ENC/us30/n1093 ), .ZN(\AES_ENC/us30/n1111 ) );
NAND2_X2 \AES_ENC/us30/U25  ( .A1(\AES_ENC/us30/n1092 ), .A2(\AES_ENC/us30/n1120 ), .ZN(\AES_ENC/us30/n1110 ) );
AND2_X2 \AES_ENC/us30/U22  ( .A1(\AES_ENC/us30/n1097 ), .A2(\AES_ENC/us30/n1096 ), .ZN(\AES_ENC/us30/n1098 ) );
NAND4_X2 \AES_ENC/us30/U14  ( .A1(\AES_ENC/us30/n1111 ), .A2(\AES_ENC/us30/n1110 ), .A3(\AES_ENC/us30/n1109 ), .A4(\AES_ENC/us30/n1108 ), .ZN(\AES_ENC/us30/n1112 ) );
NAND2_X2 \AES_ENC/us30/U13  ( .A1(\AES_ENC/us30/n1113 ), .A2(\AES_ENC/us30/n1112 ), .ZN(\AES_ENC/us30/n1133 ) );
NAND2_X2 \AES_ENC/us30/U12  ( .A1(\AES_ENC/us30/n1115 ), .A2(\AES_ENC/us30/n1114 ), .ZN(\AES_ENC/us30/n1129 ) );
OR2_X2 \AES_ENC/us30/U11  ( .A1(\AES_ENC/us30/n608 ), .A2(\AES_ENC/us30/n1116 ), .ZN(\AES_ENC/us30/n1128 ) );
NAND4_X2 \AES_ENC/us30/U3  ( .A1(\AES_ENC/us30/n1129 ), .A2(\AES_ENC/us30/n1128 ), .A3(\AES_ENC/us30/n1127 ), .A4(\AES_ENC/us30/n1126 ), .ZN(\AES_ENC/us30/n1130 ) );
NAND2_X2 \AES_ENC/us30/U2  ( .A1(\AES_ENC/us30/n1131 ), .A2(\AES_ENC/us30/n1130 ), .ZN(\AES_ENC/us30/n1132 ) );
NAND4_X2 \AES_ENC/us30/U1  ( .A1(\AES_ENC/us30/n1135 ), .A2(\AES_ENC/us30/n1134 ), .A3(\AES_ENC/us30/n1133 ), .A4(\AES_ENC/us30/n1132 ), .ZN(\AES_ENC/sa30_sub[7] ) );
INV_X4 \AES_ENC/us31/U575  ( .A(\AES_ENC/sa31 [7]), .ZN(\AES_ENC/us31/n627 ));
INV_X4 \AES_ENC/us31/U574  ( .A(\AES_ENC/us31/n1114 ), .ZN(\AES_ENC/us31/n625 ) );
INV_X4 \AES_ENC/us31/U573  ( .A(\AES_ENC/sa31 [4]), .ZN(\AES_ENC/us31/n624 ));
INV_X4 \AES_ENC/us31/U572  ( .A(\AES_ENC/us31/n1025 ), .ZN(\AES_ENC/us31/n622 ) );
INV_X4 \AES_ENC/us31/U571  ( .A(\AES_ENC/us31/n1120 ), .ZN(\AES_ENC/us31/n620 ) );
INV_X4 \AES_ENC/us31/U570  ( .A(\AES_ENC/us31/n1121 ), .ZN(\AES_ENC/us31/n619 ) );
INV_X4 \AES_ENC/us31/U569  ( .A(\AES_ENC/us31/n1048 ), .ZN(\AES_ENC/us31/n618 ) );
INV_X4 \AES_ENC/us31/U568  ( .A(\AES_ENC/us31/n974 ), .ZN(\AES_ENC/us31/n616 ) );
INV_X4 \AES_ENC/us31/U567  ( .A(\AES_ENC/us31/n794 ), .ZN(\AES_ENC/us31/n614 ) );
INV_X4 \AES_ENC/us31/U566  ( .A(\AES_ENC/sa31 [2]), .ZN(\AES_ENC/us31/n611 ));
INV_X4 \AES_ENC/us31/U565  ( .A(\AES_ENC/us31/n800 ), .ZN(\AES_ENC/us31/n610 ) );
INV_X4 \AES_ENC/us31/U564  ( .A(\AES_ENC/us31/n925 ), .ZN(\AES_ENC/us31/n609 ) );
INV_X4 \AES_ENC/us31/U563  ( .A(\AES_ENC/us31/n779 ), .ZN(\AES_ENC/us31/n607 ) );
INV_X4 \AES_ENC/us31/U562  ( .A(\AES_ENC/us31/n1022 ), .ZN(\AES_ENC/us31/n603 ) );
INV_X4 \AES_ENC/us31/U561  ( .A(\AES_ENC/us31/n1102 ), .ZN(\AES_ENC/us31/n602 ) );
INV_X4 \AES_ENC/us31/U560  ( .A(\AES_ENC/us31/n929 ), .ZN(\AES_ENC/us31/n601 ) );
INV_X4 \AES_ENC/us31/U559  ( .A(\AES_ENC/us31/n1056 ), .ZN(\AES_ENC/us31/n600 ) );
INV_X4 \AES_ENC/us31/U558  ( .A(\AES_ENC/us31/n1054 ), .ZN(\AES_ENC/us31/n599 ) );
INV_X4 \AES_ENC/us31/U557  ( .A(\AES_ENC/us31/n881 ), .ZN(\AES_ENC/us31/n598 ) );
INV_X4 \AES_ENC/us31/U556  ( .A(\AES_ENC/us31/n926 ), .ZN(\AES_ENC/us31/n597 ) );
INV_X4 \AES_ENC/us31/U555  ( .A(\AES_ENC/us31/n977 ), .ZN(\AES_ENC/us31/n595 ) );
INV_X4 \AES_ENC/us31/U554  ( .A(\AES_ENC/us31/n1031 ), .ZN(\AES_ENC/us31/n594 ) );
INV_X4 \AES_ENC/us31/U553  ( .A(\AES_ENC/us31/n1103 ), .ZN(\AES_ENC/us31/n593 ) );
INV_X4 \AES_ENC/us31/U552  ( .A(\AES_ENC/us31/n1009 ), .ZN(\AES_ENC/us31/n592 ) );
INV_X4 \AES_ENC/us31/U551  ( .A(\AES_ENC/us31/n990 ), .ZN(\AES_ENC/us31/n591 ) );
INV_X4 \AES_ENC/us31/U550  ( .A(\AES_ENC/us31/n1058 ), .ZN(\AES_ENC/us31/n590 ) );
INV_X4 \AES_ENC/us31/U549  ( .A(\AES_ENC/us31/n1074 ), .ZN(\AES_ENC/us31/n589 ) );
INV_X4 \AES_ENC/us31/U548  ( .A(\AES_ENC/us31/n1053 ), .ZN(\AES_ENC/us31/n588 ) );
INV_X4 \AES_ENC/us31/U547  ( .A(\AES_ENC/us31/n826 ), .ZN(\AES_ENC/us31/n587 ) );
INV_X4 \AES_ENC/us31/U546  ( .A(\AES_ENC/us31/n992 ), .ZN(\AES_ENC/us31/n586 ) );
INV_X4 \AES_ENC/us31/U545  ( .A(\AES_ENC/us31/n821 ), .ZN(\AES_ENC/us31/n585 ) );
INV_X4 \AES_ENC/us31/U544  ( .A(\AES_ENC/us31/n910 ), .ZN(\AES_ENC/us31/n584 ) );
INV_X4 \AES_ENC/us31/U543  ( .A(\AES_ENC/us31/n906 ), .ZN(\AES_ENC/us31/n583 ) );
INV_X4 \AES_ENC/us31/U542  ( .A(\AES_ENC/us31/n880 ), .ZN(\AES_ENC/us31/n581 ) );
INV_X4 \AES_ENC/us31/U541  ( .A(\AES_ENC/us31/n1013 ), .ZN(\AES_ENC/us31/n580 ) );
INV_X4 \AES_ENC/us31/U540  ( .A(\AES_ENC/us31/n1092 ), .ZN(\AES_ENC/us31/n579 ) );
INV_X4 \AES_ENC/us31/U539  ( .A(\AES_ENC/us31/n824 ), .ZN(\AES_ENC/us31/n578 ) );
INV_X4 \AES_ENC/us31/U538  ( .A(\AES_ENC/us31/n1091 ), .ZN(\AES_ENC/us31/n577 ) );
INV_X4 \AES_ENC/us31/U537  ( .A(\AES_ENC/us31/n1080 ), .ZN(\AES_ENC/us31/n576 ) );
INV_X4 \AES_ENC/us31/U536  ( .A(\AES_ENC/us31/n959 ), .ZN(\AES_ENC/us31/n575 ) );
INV_X4 \AES_ENC/us31/U535  ( .A(\AES_ENC/sa31 [0]), .ZN(\AES_ENC/us31/n574 ));
NOR2_X2 \AES_ENC/us31/U534  ( .A1(\AES_ENC/sa31 [0]), .A2(\AES_ENC/sa31 [6]),.ZN(\AES_ENC/us31/n1090 ) );
NOR2_X2 \AES_ENC/us31/U533  ( .A1(\AES_ENC/us31/n574 ), .A2(\AES_ENC/sa31 [6]), .ZN(\AES_ENC/us31/n1070 ) );
NOR2_X2 \AES_ENC/us31/U532  ( .A1(\AES_ENC/sa31 [4]), .A2(\AES_ENC/sa31 [3]),.ZN(\AES_ENC/us31/n1025 ) );
INV_X4 \AES_ENC/us31/U531  ( .A(\AES_ENC/us31/n569 ), .ZN(\AES_ENC/us31/n572 ) );
NOR2_X2 \AES_ENC/us31/U530  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n765 ) );
NOR2_X2 \AES_ENC/us31/U529  ( .A1(\AES_ENC/sa31 [4]), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n764 ) );
NOR2_X2 \AES_ENC/us31/U528  ( .A1(\AES_ENC/us31/n765 ), .A2(\AES_ENC/us31/n764 ), .ZN(\AES_ENC/us31/n766 ) );
NOR2_X2 \AES_ENC/us31/U527  ( .A1(\AES_ENC/us31/n766 ), .A2(\AES_ENC/us31/n575 ), .ZN(\AES_ENC/us31/n767 ) );
NOR3_X2 \AES_ENC/us31/U526  ( .A1(\AES_ENC/us31/n627 ), .A2(\AES_ENC/sa31 [5]), .A3(\AES_ENC/us31/n704 ), .ZN(\AES_ENC/us31/n706 ));
NOR2_X2 \AES_ENC/us31/U525  ( .A1(\AES_ENC/us31/n1117 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n707 ) );
NOR2_X2 \AES_ENC/us31/U524  ( .A1(\AES_ENC/sa31 [4]), .A2(\AES_ENC/us31/n579 ), .ZN(\AES_ENC/us31/n705 ) );
NOR3_X2 \AES_ENC/us31/U523  ( .A1(\AES_ENC/us31/n707 ), .A2(\AES_ENC/us31/n706 ), .A3(\AES_ENC/us31/n705 ), .ZN(\AES_ENC/us31/n713 ) );
INV_X4 \AES_ENC/us31/U522  ( .A(\AES_ENC/sa31 [3]), .ZN(\AES_ENC/us31/n621 ));
NAND3_X2 \AES_ENC/us31/U521  ( .A1(\AES_ENC/us31/n652 ), .A2(\AES_ENC/us31/n626 ), .A3(\AES_ENC/sa31 [7]), .ZN(\AES_ENC/us31/n653 ));
NOR2_X2 \AES_ENC/us31/U520  ( .A1(\AES_ENC/us31/n611 ), .A2(\AES_ENC/sa31 [5]), .ZN(\AES_ENC/us31/n925 ) );
NOR2_X2 \AES_ENC/us31/U519  ( .A1(\AES_ENC/sa31 [5]), .A2(\AES_ENC/sa31 [2]),.ZN(\AES_ENC/us31/n974 ) );
INV_X4 \AES_ENC/us31/U518  ( .A(\AES_ENC/sa31 [5]), .ZN(\AES_ENC/us31/n626 ));
NOR2_X2 \AES_ENC/us31/U517  ( .A1(\AES_ENC/us31/n611 ), .A2(\AES_ENC/sa31 [7]), .ZN(\AES_ENC/us31/n779 ) );
NAND3_X2 \AES_ENC/us31/U516  ( .A1(\AES_ENC/us31/n679 ), .A2(\AES_ENC/us31/n678 ), .A3(\AES_ENC/us31/n677 ), .ZN(\AES_ENC/sa31_sub[0] ) );
NOR2_X2 \AES_ENC/us31/U515  ( .A1(\AES_ENC/us31/n626 ), .A2(\AES_ENC/sa31 [2]), .ZN(\AES_ENC/us31/n1048 ) );
NOR4_X2 \AES_ENC/us31/U512  ( .A1(\AES_ENC/us31/n633 ), .A2(\AES_ENC/us31/n632 ), .A3(\AES_ENC/us31/n631 ), .A4(\AES_ENC/us31/n630 ), .ZN(\AES_ENC/us31/n634 ) );
NOR2_X2 \AES_ENC/us31/U510  ( .A1(\AES_ENC/us31/n629 ), .A2(\AES_ENC/us31/n628 ), .ZN(\AES_ENC/us31/n635 ) );
NAND3_X2 \AES_ENC/us31/U509  ( .A1(\AES_ENC/sa31 [2]), .A2(\AES_ENC/sa31 [7]), .A3(\AES_ENC/us31/n1059 ), .ZN(\AES_ENC/us31/n636 ) );
NOR2_X2 \AES_ENC/us31/U508  ( .A1(\AES_ENC/sa31 [7]), .A2(\AES_ENC/sa31 [2]),.ZN(\AES_ENC/us31/n794 ) );
NOR2_X2 \AES_ENC/us31/U507  ( .A1(\AES_ENC/sa31 [4]), .A2(\AES_ENC/sa31 [1]),.ZN(\AES_ENC/us31/n1102 ) );
NOR2_X2 \AES_ENC/us31/U506  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/sa31 [3]), .ZN(\AES_ENC/us31/n1053 ) );
NOR2_X2 \AES_ENC/us31/U505  ( .A1(\AES_ENC/us31/n607 ), .A2(\AES_ENC/sa31 [5]), .ZN(\AES_ENC/us31/n1024 ) );
NOR2_X2 \AES_ENC/us31/U504  ( .A1(\AES_ENC/us31/n625 ), .A2(\AES_ENC/sa31 [2]), .ZN(\AES_ENC/us31/n1093 ) );
NOR2_X2 \AES_ENC/us31/U503  ( .A1(\AES_ENC/us31/n614 ), .A2(\AES_ENC/sa31 [5]), .ZN(\AES_ENC/us31/n1094 ) );
NOR2_X2 \AES_ENC/us31/U502  ( .A1(\AES_ENC/us31/n624 ), .A2(\AES_ENC/sa31 [3]), .ZN(\AES_ENC/us31/n931 ) );
INV_X4 \AES_ENC/us31/U501  ( .A(\AES_ENC/us31/n570 ), .ZN(\AES_ENC/us31/n573 ) );
NOR2_X2 \AES_ENC/us31/U500  ( .A1(\AES_ENC/us31/n1053 ), .A2(\AES_ENC/us31/n1095 ), .ZN(\AES_ENC/us31/n639 ) );
NOR3_X2 \AES_ENC/us31/U499  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n573 ), .A3(\AES_ENC/us31/n1074 ), .ZN(\AES_ENC/us31/n641 ) );
NOR2_X2 \AES_ENC/us31/U498  ( .A1(\AES_ENC/us31/n639 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n640 ) );
NOR2_X2 \AES_ENC/us31/U497  ( .A1(\AES_ENC/us31/n641 ), .A2(\AES_ENC/us31/n640 ), .ZN(\AES_ENC/us31/n646 ) );
NOR3_X2 \AES_ENC/us31/U496  ( .A1(\AES_ENC/us31/n995 ), .A2(\AES_ENC/us31/n586 ), .A3(\AES_ENC/us31/n994 ), .ZN(\AES_ENC/us31/n1002 ) );
NOR2_X2 \AES_ENC/us31/U495  ( .A1(\AES_ENC/us31/n909 ), .A2(\AES_ENC/us31/n908 ), .ZN(\AES_ENC/us31/n920 ) );
NOR2_X2 \AES_ENC/us31/U494  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n823 ) );
NOR2_X2 \AES_ENC/us31/U492  ( .A1(\AES_ENC/us31/n624 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n822 ) );
NOR2_X2 \AES_ENC/us31/U491  ( .A1(\AES_ENC/us31/n823 ), .A2(\AES_ENC/us31/n822 ), .ZN(\AES_ENC/us31/n825 ) );
NOR2_X2 \AES_ENC/us31/U490  ( .A1(\AES_ENC/sa31 [1]), .A2(\AES_ENC/us31/n623 ), .ZN(\AES_ENC/us31/n913 ) );
NOR2_X2 \AES_ENC/us31/U489  ( .A1(\AES_ENC/us31/n913 ), .A2(\AES_ENC/us31/n1091 ), .ZN(\AES_ENC/us31/n914 ) );
NOR2_X2 \AES_ENC/us31/U488  ( .A1(\AES_ENC/us31/n826 ), .A2(\AES_ENC/us31/n572 ), .ZN(\AES_ENC/us31/n827 ) );
NOR3_X2 \AES_ENC/us31/U487  ( .A1(\AES_ENC/us31/n769 ), .A2(\AES_ENC/us31/n768 ), .A3(\AES_ENC/us31/n767 ), .ZN(\AES_ENC/us31/n775 ) );
NOR2_X2 \AES_ENC/us31/U486  ( .A1(\AES_ENC/us31/n1056 ), .A2(\AES_ENC/us31/n1053 ), .ZN(\AES_ENC/us31/n749 ) );
NOR2_X2 \AES_ENC/us31/U483  ( .A1(\AES_ENC/us31/n749 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n752 ) );
INV_X4 \AES_ENC/us31/U482  ( .A(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n596 ));
NOR2_X2 \AES_ENC/us31/U480  ( .A1(\AES_ENC/us31/n1054 ), .A2(\AES_ENC/us31/n1053 ), .ZN(\AES_ENC/us31/n1055 ) );
OR2_X4 \AES_ENC/us31/U479  ( .A1(\AES_ENC/us31/n1094 ), .A2(\AES_ENC/us31/n1093 ), .ZN(\AES_ENC/us31/n571 ) );
AND2_X2 \AES_ENC/us31/U478  ( .A1(\AES_ENC/us31/n571 ), .A2(\AES_ENC/us31/n1095 ), .ZN(\AES_ENC/us31/n1101 ) );
NOR2_X2 \AES_ENC/us31/U477  ( .A1(\AES_ENC/us31/n1074 ), .A2(\AES_ENC/us31/n931 ), .ZN(\AES_ENC/us31/n796 ) );
NOR2_X2 \AES_ENC/us31/U474  ( .A1(\AES_ENC/us31/n796 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n797 ) );
NOR2_X2 \AES_ENC/us31/U473  ( .A1(\AES_ENC/us31/n932 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n933 ) );
NOR2_X2 \AES_ENC/us31/U472  ( .A1(\AES_ENC/us31/n929 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n935 ) );
NOR2_X2 \AES_ENC/us31/U471  ( .A1(\AES_ENC/us31/n931 ), .A2(\AES_ENC/us31/n930 ), .ZN(\AES_ENC/us31/n934 ) );
NOR3_X2 \AES_ENC/us31/U470  ( .A1(\AES_ENC/us31/n935 ), .A2(\AES_ENC/us31/n934 ), .A3(\AES_ENC/us31/n933 ), .ZN(\AES_ENC/us31/n936 ) );
NOR2_X2 \AES_ENC/us31/U469  ( .A1(\AES_ENC/us31/n624 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n1075 ) );
NOR2_X2 \AES_ENC/us31/U468  ( .A1(\AES_ENC/us31/n572 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n949 ) );
NOR2_X2 \AES_ENC/us31/U467  ( .A1(\AES_ENC/us31/n1049 ), .A2(\AES_ENC/us31/n618 ), .ZN(\AES_ENC/us31/n1051 ) );
NOR2_X2 \AES_ENC/us31/U466  ( .A1(\AES_ENC/us31/n1051 ), .A2(\AES_ENC/us31/n1050 ), .ZN(\AES_ENC/us31/n1052 ) );
NOR2_X2 \AES_ENC/us31/U465  ( .A1(\AES_ENC/us31/n1052 ), .A2(\AES_ENC/us31/n592 ), .ZN(\AES_ENC/us31/n1064 ) );
NOR2_X2 \AES_ENC/us31/U464  ( .A1(\AES_ENC/sa31 [1]), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n631 ) );
NOR2_X2 \AES_ENC/us31/U463  ( .A1(\AES_ENC/us31/n1025 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n980 ) );
NOR2_X2 \AES_ENC/us31/U462  ( .A1(\AES_ENC/us31/n1073 ), .A2(\AES_ENC/us31/n1094 ), .ZN(\AES_ENC/us31/n795 ) );
NOR2_X2 \AES_ENC/us31/U461  ( .A1(\AES_ENC/us31/n795 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n799 ) );
NOR2_X2 \AES_ENC/us31/U460  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n981 ) );
NOR2_X2 \AES_ENC/us31/U459  ( .A1(\AES_ENC/us31/n1102 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n643 ) );
NOR2_X2 \AES_ENC/us31/U458  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n621 ), .ZN(\AES_ENC/us31/n642 ) );
NOR2_X2 \AES_ENC/us31/U455  ( .A1(\AES_ENC/us31/n911 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n644 ) );
NOR4_X2 \AES_ENC/us31/U448  ( .A1(\AES_ENC/us31/n644 ), .A2(\AES_ENC/us31/n643 ), .A3(\AES_ENC/us31/n804 ), .A4(\AES_ENC/us31/n642 ), .ZN(\AES_ENC/us31/n645 ) );
NOR2_X2 \AES_ENC/us31/U447  ( .A1(\AES_ENC/us31/n1102 ), .A2(\AES_ENC/us31/n910 ), .ZN(\AES_ENC/us31/n932 ) );
NOR2_X2 \AES_ENC/us31/U442  ( .A1(\AES_ENC/us31/n1102 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n755 ) );
NOR2_X2 \AES_ENC/us31/U441  ( .A1(\AES_ENC/us31/n931 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n743 ) );
NOR2_X2 \AES_ENC/us31/U438  ( .A1(\AES_ENC/us31/n1072 ), .A2(\AES_ENC/us31/n1094 ), .ZN(\AES_ENC/us31/n930 ) );
NOR2_X2 \AES_ENC/us31/U435  ( .A1(\AES_ENC/us31/n1074 ), .A2(\AES_ENC/us31/n1025 ), .ZN(\AES_ENC/us31/n891 ) );
NOR2_X2 \AES_ENC/us31/U434  ( .A1(\AES_ENC/us31/n891 ), .A2(\AES_ENC/us31/n609 ), .ZN(\AES_ENC/us31/n894 ) );
NOR3_X2 \AES_ENC/us31/U433  ( .A1(\AES_ENC/us31/n623 ), .A2(\AES_ENC/sa31 [1]), .A3(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n683 ));
INV_X4 \AES_ENC/us31/U428  ( .A(\AES_ENC/us31/n931 ), .ZN(\AES_ENC/us31/n623 ) );
NOR2_X2 \AES_ENC/us31/U427  ( .A1(\AES_ENC/us31/n996 ), .A2(\AES_ENC/us31/n931 ), .ZN(\AES_ENC/us31/n704 ) );
NOR2_X2 \AES_ENC/us31/U421  ( .A1(\AES_ENC/us31/n931 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n685 ) );
NOR2_X2 \AES_ENC/us31/U420  ( .A1(\AES_ENC/us31/n1029 ), .A2(\AES_ENC/us31/n1025 ), .ZN(\AES_ENC/us31/n1079 ) );
NOR3_X2 \AES_ENC/us31/U419  ( .A1(\AES_ENC/us31/n589 ), .A2(\AES_ENC/us31/n1025 ), .A3(\AES_ENC/us31/n616 ), .ZN(\AES_ENC/us31/n945 ) );
NOR2_X2 \AES_ENC/us31/U418  ( .A1(\AES_ENC/us31/n626 ), .A2(\AES_ENC/us31/n611 ), .ZN(\AES_ENC/us31/n800 ) );
NOR3_X2 \AES_ENC/us31/U417  ( .A1(\AES_ENC/us31/n590 ), .A2(\AES_ENC/us31/n627 ), .A3(\AES_ENC/us31/n611 ), .ZN(\AES_ENC/us31/n798 ) );
NOR3_X2 \AES_ENC/us31/U416  ( .A1(\AES_ENC/us31/n610 ), .A2(\AES_ENC/us31/n572 ), .A3(\AES_ENC/us31/n575 ), .ZN(\AES_ENC/us31/n962 ) );
NOR3_X2 \AES_ENC/us31/U415  ( .A1(\AES_ENC/us31/n959 ), .A2(\AES_ENC/us31/n572 ), .A3(\AES_ENC/us31/n609 ), .ZN(\AES_ENC/us31/n768 ) );
NOR3_X2 \AES_ENC/us31/U414  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n572 ), .A3(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n694 ) );
NOR3_X2 \AES_ENC/us31/U413  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n572 ), .A3(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n895 ) );
NOR3_X2 \AES_ENC/us31/U410  ( .A1(\AES_ENC/us31/n1008 ), .A2(\AES_ENC/us31/n1007 ), .A3(\AES_ENC/us31/n1006 ), .ZN(\AES_ENC/us31/n1018 ) );
NOR4_X2 \AES_ENC/us31/U409  ( .A1(\AES_ENC/us31/n806 ), .A2(\AES_ENC/us31/n805 ), .A3(\AES_ENC/us31/n804 ), .A4(\AES_ENC/us31/n803 ), .ZN(\AES_ENC/us31/n807 ) );
NOR3_X2 \AES_ENC/us31/U406  ( .A1(\AES_ENC/us31/n799 ), .A2(\AES_ENC/us31/n798 ), .A3(\AES_ENC/us31/n797 ), .ZN(\AES_ENC/us31/n808 ) );
NOR2_X2 \AES_ENC/us31/U405  ( .A1(\AES_ENC/us31/n669 ), .A2(\AES_ENC/us31/n668 ), .ZN(\AES_ENC/us31/n673 ) );
NOR4_X2 \AES_ENC/us31/U404  ( .A1(\AES_ENC/us31/n946 ), .A2(\AES_ENC/us31/n1046 ), .A3(\AES_ENC/us31/n671 ), .A4(\AES_ENC/us31/n670 ), .ZN(\AES_ENC/us31/n672 ) );
NOR4_X2 \AES_ENC/us31/U403  ( .A1(\AES_ENC/us31/n711 ), .A2(\AES_ENC/us31/n710 ), .A3(\AES_ENC/us31/n709 ), .A4(\AES_ENC/us31/n708 ), .ZN(\AES_ENC/us31/n712 ) );
NOR4_X2 \AES_ENC/us31/U401  ( .A1(\AES_ENC/us31/n963 ), .A2(\AES_ENC/us31/n962 ), .A3(\AES_ENC/us31/n961 ), .A4(\AES_ENC/us31/n960 ), .ZN(\AES_ENC/us31/n964 ) );
NOR3_X2 \AES_ENC/us31/U400  ( .A1(\AES_ENC/us31/n1101 ), .A2(\AES_ENC/us31/n1100 ), .A3(\AES_ENC/us31/n1099 ), .ZN(\AES_ENC/us31/n1109 ) );
NOR4_X2 \AES_ENC/us31/U399  ( .A1(\AES_ENC/us31/n843 ), .A2(\AES_ENC/us31/n842 ), .A3(\AES_ENC/us31/n841 ), .A4(\AES_ENC/us31/n840 ), .ZN(\AES_ENC/us31/n844 ) );
NOR3_X2 \AES_ENC/us31/U398  ( .A1(\AES_ENC/us31/n743 ), .A2(\AES_ENC/us31/n742 ), .A3(\AES_ENC/us31/n741 ), .ZN(\AES_ENC/us31/n744 ) );
NOR2_X2 \AES_ENC/us31/U397  ( .A1(\AES_ENC/us31/n697 ), .A2(\AES_ENC/us31/n658 ), .ZN(\AES_ENC/us31/n659 ) );
NOR2_X2 \AES_ENC/us31/U396  ( .A1(\AES_ENC/us31/n1078 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n1033 ) );
NOR2_X2 \AES_ENC/us31/U393  ( .A1(\AES_ENC/us31/n1031 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n1032 ) );
NOR3_X2 \AES_ENC/us31/U390  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n1025 ), .A3(\AES_ENC/us31/n1074 ), .ZN(\AES_ENC/us31/n1035 ) );
NOR4_X2 \AES_ENC/us31/U389  ( .A1(\AES_ENC/us31/n1035 ), .A2(\AES_ENC/us31/n1034 ), .A3(\AES_ENC/us31/n1033 ), .A4(\AES_ENC/us31/n1032 ), .ZN(\AES_ENC/us31/n1036 ) );
NOR2_X2 \AES_ENC/us31/U388  ( .A1(\AES_ENC/us31/n598 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n885 ) );
NOR2_X2 \AES_ENC/us31/U387  ( .A1(\AES_ENC/us31/n623 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n882 ) );
NOR2_X2 \AES_ENC/us31/U386  ( .A1(\AES_ENC/us31/n1053 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n884 ) );
NOR4_X2 \AES_ENC/us31/U385  ( .A1(\AES_ENC/us31/n885 ), .A2(\AES_ENC/us31/n884 ), .A3(\AES_ENC/us31/n883 ), .A4(\AES_ENC/us31/n882 ), .ZN(\AES_ENC/us31/n886 ) );
NOR2_X2 \AES_ENC/us31/U384  ( .A1(\AES_ENC/us31/n825 ), .A2(\AES_ENC/us31/n578 ), .ZN(\AES_ENC/us31/n830 ) );
NOR2_X2 \AES_ENC/us31/U383  ( .A1(\AES_ENC/us31/n827 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n829 ) );
NOR2_X2 \AES_ENC/us31/U382  ( .A1(\AES_ENC/us31/n572 ), .A2(\AES_ENC/us31/n579 ), .ZN(\AES_ENC/us31/n828 ) );
NOR4_X2 \AES_ENC/us31/U374  ( .A1(\AES_ENC/us31/n831 ), .A2(\AES_ENC/us31/n830 ), .A3(\AES_ENC/us31/n829 ), .A4(\AES_ENC/us31/n828 ), .ZN(\AES_ENC/us31/n832 ) );
NOR2_X2 \AES_ENC/us31/U373  ( .A1(\AES_ENC/us31/n606 ), .A2(\AES_ENC/us31/n582 ), .ZN(\AES_ENC/us31/n1104 ) );
NOR2_X2 \AES_ENC/us31/U372  ( .A1(\AES_ENC/us31/n1102 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n1106 ) );
NOR2_X2 \AES_ENC/us31/U370  ( .A1(\AES_ENC/us31/n1103 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n1105 ) );
NOR4_X2 \AES_ENC/us31/U369  ( .A1(\AES_ENC/us31/n1107 ), .A2(\AES_ENC/us31/n1106 ), .A3(\AES_ENC/us31/n1105 ), .A4(\AES_ENC/us31/n1104 ), .ZN(\AES_ENC/us31/n1108 ) );
NOR3_X2 \AES_ENC/us31/U368  ( .A1(\AES_ENC/us31/n959 ), .A2(\AES_ENC/us31/n621 ), .A3(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n963 ) );
NOR2_X2 \AES_ENC/us31/U367  ( .A1(\AES_ENC/us31/n626 ), .A2(\AES_ENC/us31/n627 ), .ZN(\AES_ENC/us31/n1114 ) );
INV_X4 \AES_ENC/us31/U366  ( .A(\AES_ENC/us31/n1024 ), .ZN(\AES_ENC/us31/n606 ) );
NOR3_X2 \AES_ENC/us31/U365  ( .A1(\AES_ENC/us31/n910 ), .A2(\AES_ENC/us31/n1059 ), .A3(\AES_ENC/us31/n611 ), .ZN(\AES_ENC/us31/n1115 ) );
INV_X4 \AES_ENC/us31/U364  ( .A(\AES_ENC/us31/n1094 ), .ZN(\AES_ENC/us31/n613 ) );
NOR2_X2 \AES_ENC/us31/U363  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n931 ), .ZN(\AES_ENC/us31/n1100 ) );
INV_X4 \AES_ENC/us31/U354  ( .A(\AES_ENC/us31/n1093 ), .ZN(\AES_ENC/us31/n617 ) );
NOR2_X2 \AES_ENC/us31/U353  ( .A1(\AES_ENC/us31/n569 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n929 ) );
NOR2_X2 \AES_ENC/us31/U352  ( .A1(\AES_ENC/us31/n620 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n926 ) );
NOR2_X2 \AES_ENC/us31/U351  ( .A1(\AES_ENC/us31/n572 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n1095 ) );
NOR2_X2 \AES_ENC/us31/U350  ( .A1(\AES_ENC/us31/n609 ), .A2(\AES_ENC/us31/n627 ), .ZN(\AES_ENC/us31/n1010 ) );
NOR2_X2 \AES_ENC/us31/U349  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n1103 ) );
NOR2_X2 \AES_ENC/us31/U348  ( .A1(\AES_ENC/us31/n622 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n1059 ) );
NOR2_X2 \AES_ENC/us31/U347  ( .A1(\AES_ENC/sa31 [1]), .A2(\AES_ENC/us31/n1120 ), .ZN(\AES_ENC/us31/n1022 ) );
NOR2_X2 \AES_ENC/us31/U346  ( .A1(\AES_ENC/us31/n619 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n911 ) );
NOR2_X2 \AES_ENC/us31/U345  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/us31/n1025 ), .ZN(\AES_ENC/us31/n826 ) );
NOR2_X2 \AES_ENC/us31/U338  ( .A1(\AES_ENC/us31/n626 ), .A2(\AES_ENC/us31/n607 ), .ZN(\AES_ENC/us31/n1072 ) );
NOR2_X2 \AES_ENC/us31/U335  ( .A1(\AES_ENC/us31/n627 ), .A2(\AES_ENC/us31/n616 ), .ZN(\AES_ENC/us31/n956 ) );
NOR2_X2 \AES_ENC/us31/U329  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/us31/n624 ), .ZN(\AES_ENC/us31/n1121 ) );
NOR2_X2 \AES_ENC/us31/U328  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/us31/n624 ), .ZN(\AES_ENC/us31/n1058 ) );
NOR2_X2 \AES_ENC/us31/U327  ( .A1(\AES_ENC/us31/n625 ), .A2(\AES_ENC/us31/n611 ), .ZN(\AES_ENC/us31/n1073 ) );
NOR2_X2 \AES_ENC/us31/U325  ( .A1(\AES_ENC/sa31 [1]), .A2(\AES_ENC/us31/n1025 ), .ZN(\AES_ENC/us31/n1054 ) );
NOR2_X2 \AES_ENC/us31/U324  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/us31/n931 ), .ZN(\AES_ENC/us31/n1029 ) );
NOR2_X2 \AES_ENC/us31/U319  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n1056 ) );
NOR2_X2 \AES_ENC/us31/U318  ( .A1(\AES_ENC/us31/n614 ), .A2(\AES_ENC/us31/n626 ), .ZN(\AES_ENC/us31/n1050 ) );
NOR2_X2 \AES_ENC/us31/U317  ( .A1(\AES_ENC/us31/n1121 ), .A2(\AES_ENC/us31/n1025 ), .ZN(\AES_ENC/us31/n1120 ) );
NOR2_X2 \AES_ENC/us31/U316  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/us31/n572 ), .ZN(\AES_ENC/us31/n1074 ) );
NOR2_X2 \AES_ENC/us31/U315  ( .A1(\AES_ENC/us31/n1058 ), .A2(\AES_ENC/us31/n1054 ), .ZN(\AES_ENC/us31/n878 ) );
NOR2_X2 \AES_ENC/us31/U314  ( .A1(\AES_ENC/us31/n878 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n879 ) );
NOR2_X2 \AES_ENC/us31/U312  ( .A1(\AES_ENC/us31/n880 ), .A2(\AES_ENC/us31/n879 ), .ZN(\AES_ENC/us31/n887 ) );
NOR2_X2 \AES_ENC/us31/U311  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n588 ), .ZN(\AES_ENC/us31/n957 ) );
NOR2_X2 \AES_ENC/us31/U310  ( .A1(\AES_ENC/us31/n958 ), .A2(\AES_ENC/us31/n957 ), .ZN(\AES_ENC/us31/n965 ) );
NOR3_X2 \AES_ENC/us31/U309  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n1091 ), .A3(\AES_ENC/us31/n1022 ), .ZN(\AES_ENC/us31/n720 ) );
NOR3_X2 \AES_ENC/us31/U303  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n1054 ), .A3(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n719 ) );
NOR2_X2 \AES_ENC/us31/U302  ( .A1(\AES_ENC/us31/n720 ), .A2(\AES_ENC/us31/n719 ), .ZN(\AES_ENC/us31/n726 ) );
NOR2_X2 \AES_ENC/us31/U300  ( .A1(\AES_ENC/us31/n614 ), .A2(\AES_ENC/us31/n591 ), .ZN(\AES_ENC/us31/n865 ) );
NOR2_X2 \AES_ENC/us31/U299  ( .A1(\AES_ENC/us31/n1059 ), .A2(\AES_ENC/us31/n1058 ), .ZN(\AES_ENC/us31/n1060 ) );
NOR2_X2 \AES_ENC/us31/U298  ( .A1(\AES_ENC/us31/n1095 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n668 ) );
NOR2_X2 \AES_ENC/us31/U297  ( .A1(\AES_ENC/us31/n911 ), .A2(\AES_ENC/us31/n910 ), .ZN(\AES_ENC/us31/n912 ) );
NOR2_X2 \AES_ENC/us31/U296  ( .A1(\AES_ENC/us31/n912 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n916 ) );
NOR2_X2 \AES_ENC/us31/U295  ( .A1(\AES_ENC/us31/n826 ), .A2(\AES_ENC/us31/n573 ), .ZN(\AES_ENC/us31/n750 ) );
NOR2_X2 \AES_ENC/us31/U294  ( .A1(\AES_ENC/us31/n750 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n751 ) );
NOR2_X2 \AES_ENC/us31/U293  ( .A1(\AES_ENC/us31/n907 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n908 ) );
NOR2_X2 \AES_ENC/us31/U292  ( .A1(\AES_ENC/us31/n990 ), .A2(\AES_ENC/us31/n926 ), .ZN(\AES_ENC/us31/n780 ) );
NOR2_X2 \AES_ENC/us31/U291  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n584 ), .ZN(\AES_ENC/us31/n838 ) );
NOR2_X2 \AES_ENC/us31/U290  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n602 ), .ZN(\AES_ENC/us31/n837 ) );
NOR2_X2 \AES_ENC/us31/U284  ( .A1(\AES_ENC/us31/n838 ), .A2(\AES_ENC/us31/n837 ), .ZN(\AES_ENC/us31/n845 ) );
NOR2_X2 \AES_ENC/us31/U283  ( .A1(\AES_ENC/us31/n1022 ), .A2(\AES_ENC/us31/n1058 ), .ZN(\AES_ENC/us31/n740 ) );
NOR2_X2 \AES_ENC/us31/U282  ( .A1(\AES_ENC/us31/n740 ), .A2(\AES_ENC/us31/n616 ), .ZN(\AES_ENC/us31/n742 ) );
NOR2_X2 \AES_ENC/us31/U281  ( .A1(\AES_ENC/us31/n1098 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n1099 ) );
NOR2_X2 \AES_ENC/us31/U280  ( .A1(\AES_ENC/us31/n1120 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n993 ) );
NOR2_X2 \AES_ENC/us31/U279  ( .A1(\AES_ENC/us31/n993 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n994 ) );
NOR2_X2 \AES_ENC/us31/U273  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n620 ), .ZN(\AES_ENC/us31/n1026 ) );
NOR2_X2 \AES_ENC/us31/U272  ( .A1(\AES_ENC/us31/n573 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n1027 ) );
NOR2_X2 \AES_ENC/us31/U271  ( .A1(\AES_ENC/us31/n1027 ), .A2(\AES_ENC/us31/n1026 ), .ZN(\AES_ENC/us31/n1028 ) );
NOR2_X2 \AES_ENC/us31/U270  ( .A1(\AES_ENC/us31/n1029 ), .A2(\AES_ENC/us31/n1028 ), .ZN(\AES_ENC/us31/n1034 ) );
NOR4_X2 \AES_ENC/us31/U269  ( .A1(\AES_ENC/us31/n757 ), .A2(\AES_ENC/us31/n756 ), .A3(\AES_ENC/us31/n755 ), .A4(\AES_ENC/us31/n754 ), .ZN(\AES_ENC/us31/n758 ) );
NOR2_X2 \AES_ENC/us31/U268  ( .A1(\AES_ENC/us31/n752 ), .A2(\AES_ENC/us31/n751 ), .ZN(\AES_ENC/us31/n759 ) );
NOR2_X2 \AES_ENC/us31/U267  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n1071 ), .ZN(\AES_ENC/us31/n669 ) );
NOR2_X2 \AES_ENC/us31/U263  ( .A1(\AES_ENC/us31/n1056 ), .A2(\AES_ENC/us31/n990 ), .ZN(\AES_ENC/us31/n991 ) );
NOR2_X2 \AES_ENC/us31/U262  ( .A1(\AES_ENC/us31/n991 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n995 ) );
NOR2_X2 \AES_ENC/us31/U258  ( .A1(\AES_ENC/us31/n607 ), .A2(\AES_ENC/us31/n590 ), .ZN(\AES_ENC/us31/n1008 ) );
NOR2_X2 \AES_ENC/us31/U255  ( .A1(\AES_ENC/us31/n839 ), .A2(\AES_ENC/us31/n582 ), .ZN(\AES_ENC/us31/n693 ) );
NOR2_X2 \AES_ENC/us31/U254  ( .A1(\AES_ENC/us31/n606 ), .A2(\AES_ENC/us31/n906 ), .ZN(\AES_ENC/us31/n741 ) );
NOR2_X2 \AES_ENC/us31/U253  ( .A1(\AES_ENC/us31/n1054 ), .A2(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n763 ) );
NOR2_X2 \AES_ENC/us31/U252  ( .A1(\AES_ENC/us31/n763 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n769 ) );
NOR2_X2 \AES_ENC/us31/U251  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n577 ), .ZN(\AES_ENC/us31/n1007 ) );
NOR2_X2 \AES_ENC/us31/U250  ( .A1(\AES_ENC/us31/n609 ), .A2(\AES_ENC/us31/n580 ), .ZN(\AES_ENC/us31/n1123 ) );
NOR2_X2 \AES_ENC/us31/U243  ( .A1(\AES_ENC/us31/n609 ), .A2(\AES_ENC/us31/n590 ), .ZN(\AES_ENC/us31/n710 ) );
INV_X4 \AES_ENC/us31/U242  ( .A(\AES_ENC/us31/n1029 ), .ZN(\AES_ENC/us31/n582 ) );
NOR2_X2 \AES_ENC/us31/U241  ( .A1(\AES_ENC/us31/n616 ), .A2(\AES_ENC/us31/n597 ), .ZN(\AES_ENC/us31/n883 ) );
NOR2_X2 \AES_ENC/us31/U240  ( .A1(\AES_ENC/us31/n593 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n1125 ) );
NOR2_X2 \AES_ENC/us31/U239  ( .A1(\AES_ENC/us31/n990 ), .A2(\AES_ENC/us31/n929 ), .ZN(\AES_ENC/us31/n892 ) );
NOR2_X2 \AES_ENC/us31/U238  ( .A1(\AES_ENC/us31/n892 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n893 ) );
NOR2_X2 \AES_ENC/us31/U237  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n602 ), .ZN(\AES_ENC/us31/n950 ) );
NOR2_X2 \AES_ENC/us31/U236  ( .A1(\AES_ENC/us31/n1079 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n1082 ) );
NOR2_X2 \AES_ENC/us31/U235  ( .A1(\AES_ENC/us31/n910 ), .A2(\AES_ENC/us31/n1056 ), .ZN(\AES_ENC/us31/n941 ) );
NOR2_X2 \AES_ENC/us31/U234  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n1077 ), .ZN(\AES_ENC/us31/n841 ) );
NOR2_X2 \AES_ENC/us31/U229  ( .A1(\AES_ENC/us31/n623 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n630 ) );
NOR2_X2 \AES_ENC/us31/U228  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n602 ), .ZN(\AES_ENC/us31/n806 ) );
NOR2_X2 \AES_ENC/us31/U227  ( .A1(\AES_ENC/us31/n623 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n948 ) );
NOR2_X2 \AES_ENC/us31/U226  ( .A1(\AES_ENC/us31/n606 ), .A2(\AES_ENC/us31/n589 ), .ZN(\AES_ENC/us31/n997 ) );
NOR2_X2 \AES_ENC/us31/U225  ( .A1(\AES_ENC/us31/n1121 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n1122 ) );
NOR2_X2 \AES_ENC/us31/U223  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n1023 ), .ZN(\AES_ENC/us31/n756 ) );
NOR2_X2 \AES_ENC/us31/U222  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n602 ), .ZN(\AES_ENC/us31/n870 ) );
NOR2_X2 \AES_ENC/us31/U221  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n569 ), .ZN(\AES_ENC/us31/n947 ) );
NOR2_X2 \AES_ENC/us31/U217  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n1077 ), .ZN(\AES_ENC/us31/n1084 ) );
NOR2_X2 \AES_ENC/us31/U213  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n855 ), .ZN(\AES_ENC/us31/n709 ) );
NOR2_X2 \AES_ENC/us31/U212  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n589 ), .ZN(\AES_ENC/us31/n868 ) );
NOR2_X2 \AES_ENC/us31/U211  ( .A1(\AES_ENC/us31/n1120 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n1124 ) );
NOR2_X2 \AES_ENC/us31/U210  ( .A1(\AES_ENC/us31/n1120 ), .A2(\AES_ENC/us31/n839 ), .ZN(\AES_ENC/us31/n842 ) );
NOR2_X2 \AES_ENC/us31/U209  ( .A1(\AES_ENC/us31/n1120 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n696 ) );
NOR2_X2 \AES_ENC/us31/U208  ( .A1(\AES_ENC/us31/n1074 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n1076 ) );
NOR2_X2 \AES_ENC/us31/U207  ( .A1(\AES_ENC/us31/n1074 ), .A2(\AES_ENC/us31/n620 ), .ZN(\AES_ENC/us31/n781 ) );
NOR3_X2 \AES_ENC/us31/U201  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n1056 ), .A3(\AES_ENC/us31/n990 ), .ZN(\AES_ENC/us31/n979 ) );
NOR3_X2 \AES_ENC/us31/U200  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n1058 ), .A3(\AES_ENC/us31/n1059 ), .ZN(\AES_ENC/us31/n854 ) );
NOR2_X2 \AES_ENC/us31/U199  ( .A1(\AES_ENC/us31/n996 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n869 ) );
NOR2_X2 \AES_ENC/us31/U198  ( .A1(\AES_ENC/us31/n1056 ), .A2(\AES_ENC/us31/n1074 ), .ZN(\AES_ENC/us31/n1057 ) );
NOR3_X2 \AES_ENC/us31/U197  ( .A1(\AES_ENC/us31/n607 ), .A2(\AES_ENC/us31/n1120 ), .A3(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n978 ) );
NOR2_X2 \AES_ENC/us31/U196  ( .A1(\AES_ENC/us31/n996 ), .A2(\AES_ENC/us31/n911 ), .ZN(\AES_ENC/us31/n1116 ) );
NOR2_X2 \AES_ENC/us31/U195  ( .A1(\AES_ENC/us31/n1074 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n754 ) );
NOR2_X2 \AES_ENC/us31/U194  ( .A1(\AES_ENC/us31/n926 ), .A2(\AES_ENC/us31/n1103 ), .ZN(\AES_ENC/us31/n977 ) );
NOR2_X2 \AES_ENC/us31/U187  ( .A1(\AES_ENC/us31/n839 ), .A2(\AES_ENC/us31/n824 ), .ZN(\AES_ENC/us31/n1092 ) );
NOR2_X2 \AES_ENC/us31/U186  ( .A1(\AES_ENC/us31/n573 ), .A2(\AES_ENC/us31/n1074 ), .ZN(\AES_ENC/us31/n684 ) );
NOR2_X2 \AES_ENC/us31/U185  ( .A1(\AES_ENC/us31/n826 ), .A2(\AES_ENC/us31/n1059 ), .ZN(\AES_ENC/us31/n907 ) );
NOR3_X2 \AES_ENC/us31/U184  ( .A1(\AES_ENC/us31/n625 ), .A2(\AES_ENC/us31/n1115 ), .A3(\AES_ENC/us31/n585 ), .ZN(\AES_ENC/us31/n831 ) );
NOR3_X2 \AES_ENC/us31/U183  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n1056 ), .A3(\AES_ENC/us31/n990 ), .ZN(\AES_ENC/us31/n896 ) );
NOR3_X2 \AES_ENC/us31/U182  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n573 ), .A3(\AES_ENC/us31/n1013 ), .ZN(\AES_ENC/us31/n670 ) );
NOR3_X2 \AES_ENC/us31/U181  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n1091 ), .A3(\AES_ENC/us31/n1022 ), .ZN(\AES_ENC/us31/n843 ) );
NOR2_X2 \AES_ENC/us31/U180  ( .A1(\AES_ENC/us31/n1029 ), .A2(\AES_ENC/us31/n1095 ), .ZN(\AES_ENC/us31/n735 ) );
NOR2_X2 \AES_ENC/us31/U174  ( .A1(\AES_ENC/us31/n1100 ), .A2(\AES_ENC/us31/n854 ), .ZN(\AES_ENC/us31/n860 ) );
NAND3_X2 \AES_ENC/us31/U173  ( .A1(\AES_ENC/us31/n569 ), .A2(\AES_ENC/us31/n582 ), .A3(\AES_ENC/us31/n681 ), .ZN(\AES_ENC/us31/n691 ) );
NOR2_X2 \AES_ENC/us31/U172  ( .A1(\AES_ENC/us31/n683 ), .A2(\AES_ENC/us31/n682 ), .ZN(\AES_ENC/us31/n690 ) );
NOR3_X2 \AES_ENC/us31/U171  ( .A1(\AES_ENC/us31/n695 ), .A2(\AES_ENC/us31/n694 ), .A3(\AES_ENC/us31/n693 ), .ZN(\AES_ENC/us31/n700 ) );
NOR4_X2 \AES_ENC/us31/U170  ( .A1(\AES_ENC/us31/n983 ), .A2(\AES_ENC/us31/n698 ), .A3(\AES_ENC/us31/n697 ), .A4(\AES_ENC/us31/n696 ), .ZN(\AES_ENC/us31/n699 ) );
NOR2_X2 \AES_ENC/us31/U169  ( .A1(\AES_ENC/us31/n946 ), .A2(\AES_ENC/us31/n945 ), .ZN(\AES_ENC/us31/n952 ) );
NOR4_X2 \AES_ENC/us31/U168  ( .A1(\AES_ENC/us31/n950 ), .A2(\AES_ENC/us31/n949 ), .A3(\AES_ENC/us31/n948 ), .A4(\AES_ENC/us31/n947 ), .ZN(\AES_ENC/us31/n951 ) );
NOR4_X2 \AES_ENC/us31/U162  ( .A1(\AES_ENC/us31/n896 ), .A2(\AES_ENC/us31/n895 ), .A3(\AES_ENC/us31/n894 ), .A4(\AES_ENC/us31/n893 ), .ZN(\AES_ENC/us31/n897 ) );
NOR2_X2 \AES_ENC/us31/U161  ( .A1(\AES_ENC/us31/n866 ), .A2(\AES_ENC/us31/n865 ), .ZN(\AES_ENC/us31/n872 ) );
NOR4_X2 \AES_ENC/us31/U160  ( .A1(\AES_ENC/us31/n870 ), .A2(\AES_ENC/us31/n869 ), .A3(\AES_ENC/us31/n868 ), .A4(\AES_ENC/us31/n867 ), .ZN(\AES_ENC/us31/n871 ) );
NOR4_X2 \AES_ENC/us31/U159  ( .A1(\AES_ENC/us31/n983 ), .A2(\AES_ENC/us31/n982 ), .A3(\AES_ENC/us31/n981 ), .A4(\AES_ENC/us31/n980 ), .ZN(\AES_ENC/us31/n984 ) );
NOR2_X2 \AES_ENC/us31/U158  ( .A1(\AES_ENC/us31/n979 ), .A2(\AES_ENC/us31/n978 ), .ZN(\AES_ENC/us31/n985 ) );
NOR4_X2 \AES_ENC/us31/U157  ( .A1(\AES_ENC/us31/n1125 ), .A2(\AES_ENC/us31/n1124 ), .A3(\AES_ENC/us31/n1123 ), .A4(\AES_ENC/us31/n1122 ), .ZN(\AES_ENC/us31/n1126 ) );
NOR4_X2 \AES_ENC/us31/U156  ( .A1(\AES_ENC/us31/n1084 ), .A2(\AES_ENC/us31/n1083 ), .A3(\AES_ENC/us31/n1082 ), .A4(\AES_ENC/us31/n1081 ), .ZN(\AES_ENC/us31/n1085 ) );
NOR2_X2 \AES_ENC/us31/U155  ( .A1(\AES_ENC/us31/n1076 ), .A2(\AES_ENC/us31/n1075 ), .ZN(\AES_ENC/us31/n1086 ) );
NOR3_X2 \AES_ENC/us31/U154  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n1054 ), .A3(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n961 ) );
NOR3_X2 \AES_ENC/us31/U153  ( .A1(\AES_ENC/us31/n620 ), .A2(\AES_ENC/us31/n1074 ), .A3(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n671 ) );
NOR2_X2 \AES_ENC/us31/U152  ( .A1(\AES_ENC/us31/n1057 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n1062 ) );
NOR2_X2 \AES_ENC/us31/U143  ( .A1(\AES_ENC/us31/n1055 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n1063 ) );
NOR2_X2 \AES_ENC/us31/U142  ( .A1(\AES_ENC/us31/n1060 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n1061 ) );
NOR4_X2 \AES_ENC/us31/U141  ( .A1(\AES_ENC/us31/n1064 ), .A2(\AES_ENC/us31/n1063 ), .A3(\AES_ENC/us31/n1062 ), .A4(\AES_ENC/us31/n1061 ), .ZN(\AES_ENC/us31/n1065 ) );
NOR3_X2 \AES_ENC/us31/U140  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n1120 ), .A3(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n918 ) );
NOR3_X2 \AES_ENC/us31/U132  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n573 ), .A3(\AES_ENC/us31/n1013 ), .ZN(\AES_ENC/us31/n917 ) );
NOR2_X2 \AES_ENC/us31/U131  ( .A1(\AES_ENC/us31/n914 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n915 ) );
NOR4_X2 \AES_ENC/us31/U130  ( .A1(\AES_ENC/us31/n918 ), .A2(\AES_ENC/us31/n917 ), .A3(\AES_ENC/us31/n916 ), .A4(\AES_ENC/us31/n915 ), .ZN(\AES_ENC/us31/n919 ) );
NOR2_X2 \AES_ENC/us31/U129  ( .A1(\AES_ENC/us31/n616 ), .A2(\AES_ENC/us31/n580 ), .ZN(\AES_ENC/us31/n771 ) );
NOR2_X2 \AES_ENC/us31/U128  ( .A1(\AES_ENC/us31/n1103 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n772 ) );
NOR2_X2 \AES_ENC/us31/U127  ( .A1(\AES_ENC/us31/n610 ), .A2(\AES_ENC/us31/n599 ), .ZN(\AES_ENC/us31/n773 ) );
NOR4_X2 \AES_ENC/us31/U126  ( .A1(\AES_ENC/us31/n773 ), .A2(\AES_ENC/us31/n772 ), .A3(\AES_ENC/us31/n771 ), .A4(\AES_ENC/us31/n770 ), .ZN(\AES_ENC/us31/n774 ) );
NOR2_X2 \AES_ENC/us31/U121  ( .A1(\AES_ENC/us31/n735 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n687 ) );
NOR2_X2 \AES_ENC/us31/U120  ( .A1(\AES_ENC/us31/n684 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n688 ) );
NOR2_X2 \AES_ENC/us31/U119  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n600 ), .ZN(\AES_ENC/us31/n686 ) );
NOR4_X2 \AES_ENC/us31/U118  ( .A1(\AES_ENC/us31/n688 ), .A2(\AES_ENC/us31/n687 ), .A3(\AES_ENC/us31/n686 ), .A4(\AES_ENC/us31/n685 ), .ZN(\AES_ENC/us31/n689 ) );
NOR2_X2 \AES_ENC/us31/U117  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n595 ), .ZN(\AES_ENC/us31/n858 ) );
NOR2_X2 \AES_ENC/us31/U116  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n855 ), .ZN(\AES_ENC/us31/n857 ) );
NOR2_X2 \AES_ENC/us31/U115  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n587 ), .ZN(\AES_ENC/us31/n856 ) );
NOR4_X2 \AES_ENC/us31/U106  ( .A1(\AES_ENC/us31/n858 ), .A2(\AES_ENC/us31/n857 ), .A3(\AES_ENC/us31/n856 ), .A4(\AES_ENC/us31/n958 ), .ZN(\AES_ENC/us31/n859 ) );
NOR2_X2 \AES_ENC/us31/U105  ( .A1(\AES_ENC/us31/n780 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n784 ) );
NOR2_X2 \AES_ENC/us31/U104  ( .A1(\AES_ENC/us31/n1117 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n782 ) );
NOR2_X2 \AES_ENC/us31/U103  ( .A1(\AES_ENC/us31/n781 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n783 ) );
NOR4_X2 \AES_ENC/us31/U102  ( .A1(\AES_ENC/us31/n880 ), .A2(\AES_ENC/us31/n784 ), .A3(\AES_ENC/us31/n783 ), .A4(\AES_ENC/us31/n782 ), .ZN(\AES_ENC/us31/n785 ) );
NOR2_X2 \AES_ENC/us31/U101  ( .A1(\AES_ENC/us31/n583 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n814 ) );
NOR2_X2 \AES_ENC/us31/U100  ( .A1(\AES_ENC/us31/n907 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n813 ) );
NOR3_X2 \AES_ENC/us31/U95  ( .A1(\AES_ENC/us31/n606 ), .A2(\AES_ENC/us31/n1058 ), .A3(\AES_ENC/us31/n1059 ), .ZN(\AES_ENC/us31/n815 ) );
NOR4_X2 \AES_ENC/us31/U94  ( .A1(\AES_ENC/us31/n815 ), .A2(\AES_ENC/us31/n814 ), .A3(\AES_ENC/us31/n813 ), .A4(\AES_ENC/us31/n812 ), .ZN(\AES_ENC/us31/n816 ) );
NOR2_X2 \AES_ENC/us31/U93  ( .A1(\AES_ENC/us31/n617 ), .A2(\AES_ENC/us31/n569 ), .ZN(\AES_ENC/us31/n721 ) );
NOR2_X2 \AES_ENC/us31/U92  ( .A1(\AES_ENC/us31/n1031 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n723 ) );
NOR2_X2 \AES_ENC/us31/U91  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n1096 ), .ZN(\AES_ENC/us31/n722 ) );
NOR4_X2 \AES_ENC/us31/U90  ( .A1(\AES_ENC/us31/n724 ), .A2(\AES_ENC/us31/n723 ), .A3(\AES_ENC/us31/n722 ), .A4(\AES_ENC/us31/n721 ), .ZN(\AES_ENC/us31/n725 ) );
NOR2_X2 \AES_ENC/us31/U89  ( .A1(\AES_ENC/us31/n911 ), .A2(\AES_ENC/us31/n990 ), .ZN(\AES_ENC/us31/n1009 ) );
NOR2_X2 \AES_ENC/us31/U88  ( .A1(\AES_ENC/us31/n1013 ), .A2(\AES_ENC/us31/n573 ), .ZN(\AES_ENC/us31/n1014 ) );
NOR2_X2 \AES_ENC/us31/U87  ( .A1(\AES_ENC/us31/n1014 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n1015 ) );
NOR4_X2 \AES_ENC/us31/U86  ( .A1(\AES_ENC/us31/n1016 ), .A2(\AES_ENC/us31/n1015 ), .A3(\AES_ENC/us31/n1119 ), .A4(\AES_ENC/us31/n1046 ), .ZN(\AES_ENC/us31/n1017 ) );
NOR2_X2 \AES_ENC/us31/U81  ( .A1(\AES_ENC/us31/n996 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n998 ) );
NOR2_X2 \AES_ENC/us31/U80  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n577 ), .ZN(\AES_ENC/us31/n1000 ) );
NOR2_X2 \AES_ENC/us31/U79  ( .A1(\AES_ENC/us31/n616 ), .A2(\AES_ENC/us31/n1096 ), .ZN(\AES_ENC/us31/n999 ) );
NOR4_X2 \AES_ENC/us31/U78  ( .A1(\AES_ENC/us31/n1000 ), .A2(\AES_ENC/us31/n999 ), .A3(\AES_ENC/us31/n998 ), .A4(\AES_ENC/us31/n997 ), .ZN(\AES_ENC/us31/n1001 ) );
NOR2_X2 \AES_ENC/us31/U74  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n1096 ), .ZN(\AES_ENC/us31/n697 ) );
NOR2_X2 \AES_ENC/us31/U73  ( .A1(\AES_ENC/us31/n620 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n958 ) );
NOR2_X2 \AES_ENC/us31/U72  ( .A1(\AES_ENC/us31/n911 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n983 ) );
NOR2_X2 \AES_ENC/us31/U71  ( .A1(\AES_ENC/us31/n1054 ), .A2(\AES_ENC/us31/n1103 ), .ZN(\AES_ENC/us31/n1031 ) );
INV_X4 \AES_ENC/us31/U65  ( .A(\AES_ENC/us31/n1050 ), .ZN(\AES_ENC/us31/n612 ) );
INV_X4 \AES_ENC/us31/U64  ( .A(\AES_ENC/us31/n1072 ), .ZN(\AES_ENC/us31/n605 ) );
INV_X4 \AES_ENC/us31/U63  ( .A(\AES_ENC/us31/n1073 ), .ZN(\AES_ENC/us31/n604 ) );
NOR2_X2 \AES_ENC/us31/U62  ( .A1(\AES_ENC/us31/n582 ), .A2(\AES_ENC/us31/n613 ), .ZN(\AES_ENC/us31/n880 ) );
NOR3_X2 \AES_ENC/us31/U61  ( .A1(\AES_ENC/us31/n826 ), .A2(\AES_ENC/us31/n1121 ), .A3(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n946 ) );
INV_X4 \AES_ENC/us31/U59  ( .A(\AES_ENC/us31/n1010 ), .ZN(\AES_ENC/us31/n608 ) );
NOR3_X2 \AES_ENC/us31/U58  ( .A1(\AES_ENC/us31/n573 ), .A2(\AES_ENC/us31/n1029 ), .A3(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n1119 ) );
INV_X4 \AES_ENC/us31/U57  ( .A(\AES_ENC/us31/n956 ), .ZN(\AES_ENC/us31/n615 ) );
NOR2_X2 \AES_ENC/us31/U50  ( .A1(\AES_ENC/us31/n623 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n1013 ) );
NOR2_X2 \AES_ENC/us31/U49  ( .A1(\AES_ENC/us31/n620 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n910 ) );
NOR2_X2 \AES_ENC/us31/U48  ( .A1(\AES_ENC/us31/n569 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n1091 ) );
NOR2_X2 \AES_ENC/us31/U47  ( .A1(\AES_ENC/us31/n622 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n990 ) );
NOR2_X2 \AES_ENC/us31/U46  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/us31/n1121 ), .ZN(\AES_ENC/us31/n996 ) );
NOR2_X2 \AES_ENC/us31/U45  ( .A1(\AES_ENC/us31/n610 ), .A2(\AES_ENC/us31/n600 ), .ZN(\AES_ENC/us31/n628 ) );
NOR2_X2 \AES_ENC/us31/U44  ( .A1(\AES_ENC/us31/n576 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n866 ) );
NOR2_X2 \AES_ENC/us31/U43  ( .A1(\AES_ENC/us31/n603 ), .A2(\AES_ENC/us31/n610 ), .ZN(\AES_ENC/us31/n1006 ) );
NOR2_X2 \AES_ENC/us31/U42  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n1117 ), .ZN(\AES_ENC/us31/n1118 ) );
NOR2_X2 \AES_ENC/us31/U41  ( .A1(\AES_ENC/us31/n1119 ), .A2(\AES_ENC/us31/n1118 ), .ZN(\AES_ENC/us31/n1127 ) );
NOR2_X2 \AES_ENC/us31/U36  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n594 ), .ZN(\AES_ENC/us31/n629 ) );
NOR2_X2 \AES_ENC/us31/U35  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n906 ), .ZN(\AES_ENC/us31/n909 ) );
NOR2_X2 \AES_ENC/us31/U34  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n597 ), .ZN(\AES_ENC/us31/n658 ) );
NOR2_X2 \AES_ENC/us31/U33  ( .A1(\AES_ENC/us31/n1116 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n695 ) );
NOR2_X2 \AES_ENC/us31/U32  ( .A1(\AES_ENC/us31/n1078 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n1083 ) );
NOR2_X2 \AES_ENC/us31/U31  ( .A1(\AES_ENC/us31/n941 ), .A2(\AES_ENC/us31/n608 ), .ZN(\AES_ENC/us31/n724 ) );
NOR2_X2 \AES_ENC/us31/U30  ( .A1(\AES_ENC/us31/n598 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n1107 ) );
NOR2_X2 \AES_ENC/us31/U29  ( .A1(\AES_ENC/us31/n576 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n840 ) );
NOR2_X2 \AES_ENC/us31/U24  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n593 ), .ZN(\AES_ENC/us31/n633 ) );
NOR2_X2 \AES_ENC/us31/U23  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n1080 ), .ZN(\AES_ENC/us31/n1081 ) );
NOR2_X2 \AES_ENC/us31/U21  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n1045 ), .ZN(\AES_ENC/us31/n812 ) );
NOR2_X2 \AES_ENC/us31/U20  ( .A1(\AES_ENC/us31/n1009 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n960 ) );
NOR2_X2 \AES_ENC/us31/U19  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n601 ), .ZN(\AES_ENC/us31/n982 ) );
NOR2_X2 \AES_ENC/us31/U18  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n594 ), .ZN(\AES_ENC/us31/n757 ) );
NOR2_X2 \AES_ENC/us31/U17  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n590 ), .ZN(\AES_ENC/us31/n698 ) );
NOR2_X2 \AES_ENC/us31/U16  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n619 ), .ZN(\AES_ENC/us31/n708 ) );
NOR2_X2 \AES_ENC/us31/U15  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n582 ), .ZN(\AES_ENC/us31/n770 ) );
NOR2_X2 \AES_ENC/us31/U10  ( .A1(\AES_ENC/us31/n619 ), .A2(\AES_ENC/us31/n604 ), .ZN(\AES_ENC/us31/n803 ) );
NOR2_X2 \AES_ENC/us31/U9  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n881 ), .ZN(\AES_ENC/us31/n711 ) );
NOR2_X2 \AES_ENC/us31/U8  ( .A1(\AES_ENC/us31/n615 ), .A2(\AES_ENC/us31/n582 ), .ZN(\AES_ENC/us31/n867 ) );
NOR2_X2 \AES_ENC/us31/U7  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n599 ), .ZN(\AES_ENC/us31/n804 ) );
NOR2_X2 \AES_ENC/us31/U6  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n620 ), .ZN(\AES_ENC/us31/n1046 ) );
OR2_X4 \AES_ENC/us31/U5  ( .A1(\AES_ENC/us31/n624 ), .A2(\AES_ENC/sa31 [1]),.ZN(\AES_ENC/us31/n570 ) );
OR2_X4 \AES_ENC/us31/U4  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/sa31 [4]),.ZN(\AES_ENC/us31/n569 ) );
NAND2_X2 \AES_ENC/us31/U514  ( .A1(\AES_ENC/us31/n1121 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n1030 ) );
AND2_X2 \AES_ENC/us31/U513  ( .A1(\AES_ENC/us31/n597 ), .A2(\AES_ENC/us31/n1030 ), .ZN(\AES_ENC/us31/n1049 ) );
NAND2_X2 \AES_ENC/us31/U511  ( .A1(\AES_ENC/us31/n1049 ), .A2(\AES_ENC/us31/n794 ), .ZN(\AES_ENC/us31/n637 ) );
AND2_X2 \AES_ENC/us31/U493  ( .A1(\AES_ENC/us31/n779 ), .A2(\AES_ENC/us31/n996 ), .ZN(\AES_ENC/us31/n632 ) );
NAND4_X2 \AES_ENC/us31/U485  ( .A1(\AES_ENC/us31/n637 ), .A2(\AES_ENC/us31/n636 ), .A3(\AES_ENC/us31/n635 ), .A4(\AES_ENC/us31/n634 ), .ZN(\AES_ENC/us31/n638 ) );
NAND2_X2 \AES_ENC/us31/U484  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n638 ), .ZN(\AES_ENC/us31/n679 ) );
NAND2_X2 \AES_ENC/us31/U481  ( .A1(\AES_ENC/us31/n1094 ), .A2(\AES_ENC/us31/n591 ), .ZN(\AES_ENC/us31/n648 ) );
NAND2_X2 \AES_ENC/us31/U476  ( .A1(\AES_ENC/us31/n601 ), .A2(\AES_ENC/us31/n590 ), .ZN(\AES_ENC/us31/n762 ) );
NAND2_X2 \AES_ENC/us31/U475  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n762 ), .ZN(\AES_ENC/us31/n647 ) );
NAND4_X2 \AES_ENC/us31/U457  ( .A1(\AES_ENC/us31/n648 ), .A2(\AES_ENC/us31/n647 ), .A3(\AES_ENC/us31/n646 ), .A4(\AES_ENC/us31/n645 ), .ZN(\AES_ENC/us31/n649 ) );
NAND2_X2 \AES_ENC/us31/U456  ( .A1(\AES_ENC/sa31 [0]), .A2(\AES_ENC/us31/n649 ), .ZN(\AES_ENC/us31/n665 ) );
NAND2_X2 \AES_ENC/us31/U454  ( .A1(\AES_ENC/us31/n596 ), .A2(\AES_ENC/us31/n623 ), .ZN(\AES_ENC/us31/n855 ) );
NAND2_X2 \AES_ENC/us31/U453  ( .A1(\AES_ENC/us31/n587 ), .A2(\AES_ENC/us31/n855 ), .ZN(\AES_ENC/us31/n821 ) );
NAND2_X2 \AES_ENC/us31/U452  ( .A1(\AES_ENC/us31/n1093 ), .A2(\AES_ENC/us31/n821 ), .ZN(\AES_ENC/us31/n662 ) );
NAND2_X2 \AES_ENC/us31/U451  ( .A1(\AES_ENC/us31/n619 ), .A2(\AES_ENC/us31/n589 ), .ZN(\AES_ENC/us31/n650 ) );
NAND2_X2 \AES_ENC/us31/U450  ( .A1(\AES_ENC/us31/n956 ), .A2(\AES_ENC/us31/n650 ), .ZN(\AES_ENC/us31/n661 ) );
NAND2_X2 \AES_ENC/us31/U449  ( .A1(\AES_ENC/us31/n626 ), .A2(\AES_ENC/us31/n627 ), .ZN(\AES_ENC/us31/n839 ) );
OR2_X2 \AES_ENC/us31/U446  ( .A1(\AES_ENC/us31/n839 ), .A2(\AES_ENC/us31/n932 ), .ZN(\AES_ENC/us31/n656 ) );
NAND2_X2 \AES_ENC/us31/U445  ( .A1(\AES_ENC/us31/n621 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n1096 ) );
NAND2_X2 \AES_ENC/us31/U444  ( .A1(\AES_ENC/us31/n1030 ), .A2(\AES_ENC/us31/n1096 ), .ZN(\AES_ENC/us31/n651 ) );
NAND2_X2 \AES_ENC/us31/U443  ( .A1(\AES_ENC/us31/n1114 ), .A2(\AES_ENC/us31/n651 ), .ZN(\AES_ENC/us31/n655 ) );
OR3_X2 \AES_ENC/us31/U440  ( .A1(\AES_ENC/us31/n1079 ), .A2(\AES_ENC/sa31 [7]), .A3(\AES_ENC/us31/n626 ), .ZN(\AES_ENC/us31/n654 ));
NAND2_X2 \AES_ENC/us31/U439  ( .A1(\AES_ENC/us31/n593 ), .A2(\AES_ENC/us31/n601 ), .ZN(\AES_ENC/us31/n652 ) );
NAND4_X2 \AES_ENC/us31/U437  ( .A1(\AES_ENC/us31/n656 ), .A2(\AES_ENC/us31/n655 ), .A3(\AES_ENC/us31/n654 ), .A4(\AES_ENC/us31/n653 ), .ZN(\AES_ENC/us31/n657 ) );
NAND2_X2 \AES_ENC/us31/U436  ( .A1(\AES_ENC/sa31 [2]), .A2(\AES_ENC/us31/n657 ), .ZN(\AES_ENC/us31/n660 ) );
NAND4_X2 \AES_ENC/us31/U432  ( .A1(\AES_ENC/us31/n662 ), .A2(\AES_ENC/us31/n661 ), .A3(\AES_ENC/us31/n660 ), .A4(\AES_ENC/us31/n659 ), .ZN(\AES_ENC/us31/n663 ) );
NAND2_X2 \AES_ENC/us31/U431  ( .A1(\AES_ENC/us31/n663 ), .A2(\AES_ENC/us31/n574 ), .ZN(\AES_ENC/us31/n664 ) );
NAND2_X2 \AES_ENC/us31/U430  ( .A1(\AES_ENC/us31/n665 ), .A2(\AES_ENC/us31/n664 ), .ZN(\AES_ENC/us31/n666 ) );
NAND2_X2 \AES_ENC/us31/U429  ( .A1(\AES_ENC/sa31 [6]), .A2(\AES_ENC/us31/n666 ), .ZN(\AES_ENC/us31/n678 ) );
NAND2_X2 \AES_ENC/us31/U426  ( .A1(\AES_ENC/us31/n735 ), .A2(\AES_ENC/us31/n1093 ), .ZN(\AES_ENC/us31/n675 ) );
NAND2_X2 \AES_ENC/us31/U425  ( .A1(\AES_ENC/us31/n588 ), .A2(\AES_ENC/us31/n597 ), .ZN(\AES_ENC/us31/n1045 ) );
OR2_X2 \AES_ENC/us31/U424  ( .A1(\AES_ENC/us31/n1045 ), .A2(\AES_ENC/us31/n605 ), .ZN(\AES_ENC/us31/n674 ) );
NAND2_X2 \AES_ENC/us31/U423  ( .A1(\AES_ENC/sa31 [1]), .A2(\AES_ENC/us31/n620 ), .ZN(\AES_ENC/us31/n667 ) );
NAND2_X2 \AES_ENC/us31/U422  ( .A1(\AES_ENC/us31/n619 ), .A2(\AES_ENC/us31/n667 ), .ZN(\AES_ENC/us31/n1071 ) );
NAND4_X2 \AES_ENC/us31/U412  ( .A1(\AES_ENC/us31/n675 ), .A2(\AES_ENC/us31/n674 ), .A3(\AES_ENC/us31/n673 ), .A4(\AES_ENC/us31/n672 ), .ZN(\AES_ENC/us31/n676 ) );
NAND2_X2 \AES_ENC/us31/U411  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n676 ), .ZN(\AES_ENC/us31/n677 ) );
NAND2_X2 \AES_ENC/us31/U408  ( .A1(\AES_ENC/us31/n800 ), .A2(\AES_ENC/us31/n1022 ), .ZN(\AES_ENC/us31/n680 ) );
NAND2_X2 \AES_ENC/us31/U407  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n680 ), .ZN(\AES_ENC/us31/n681 ) );
AND2_X2 \AES_ENC/us31/U402  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n684 ), .ZN(\AES_ENC/us31/n682 ) );
NAND4_X2 \AES_ENC/us31/U395  ( .A1(\AES_ENC/us31/n691 ), .A2(\AES_ENC/us31/n581 ), .A3(\AES_ENC/us31/n690 ), .A4(\AES_ENC/us31/n689 ), .ZN(\AES_ENC/us31/n692 ) );
NAND2_X2 \AES_ENC/us31/U394  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n692 ), .ZN(\AES_ENC/us31/n733 ) );
NAND2_X2 \AES_ENC/us31/U392  ( .A1(\AES_ENC/us31/n977 ), .A2(\AES_ENC/us31/n1050 ), .ZN(\AES_ENC/us31/n702 ) );
NAND2_X2 \AES_ENC/us31/U391  ( .A1(\AES_ENC/us31/n1093 ), .A2(\AES_ENC/us31/n1045 ), .ZN(\AES_ENC/us31/n701 ) );
NAND4_X2 \AES_ENC/us31/U381  ( .A1(\AES_ENC/us31/n702 ), .A2(\AES_ENC/us31/n701 ), .A3(\AES_ENC/us31/n700 ), .A4(\AES_ENC/us31/n699 ), .ZN(\AES_ENC/us31/n703 ) );
NAND2_X2 \AES_ENC/us31/U380  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n703 ), .ZN(\AES_ENC/us31/n732 ) );
AND2_X2 \AES_ENC/us31/U379  ( .A1(\AES_ENC/sa31 [0]), .A2(\AES_ENC/sa31 [6]),.ZN(\AES_ENC/us31/n1113 ) );
NAND2_X2 \AES_ENC/us31/U378  ( .A1(\AES_ENC/us31/n601 ), .A2(\AES_ENC/us31/n1030 ), .ZN(\AES_ENC/us31/n881 ) );
NAND2_X2 \AES_ENC/us31/U377  ( .A1(\AES_ENC/us31/n1093 ), .A2(\AES_ENC/us31/n881 ), .ZN(\AES_ENC/us31/n715 ) );
NAND2_X2 \AES_ENC/us31/U376  ( .A1(\AES_ENC/us31/n1010 ), .A2(\AES_ENC/us31/n600 ), .ZN(\AES_ENC/us31/n714 ) );
NAND2_X2 \AES_ENC/us31/U375  ( .A1(\AES_ENC/us31/n855 ), .A2(\AES_ENC/us31/n588 ), .ZN(\AES_ENC/us31/n1117 ) );
XNOR2_X2 \AES_ENC/us31/U371  ( .A(\AES_ENC/us31/n611 ), .B(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n824 ) );
NAND4_X2 \AES_ENC/us31/U362  ( .A1(\AES_ENC/us31/n715 ), .A2(\AES_ENC/us31/n714 ), .A3(\AES_ENC/us31/n713 ), .A4(\AES_ENC/us31/n712 ), .ZN(\AES_ENC/us31/n716 ) );
NAND2_X2 \AES_ENC/us31/U361  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n716 ), .ZN(\AES_ENC/us31/n731 ) );
AND2_X2 \AES_ENC/us31/U360  ( .A1(\AES_ENC/sa31 [6]), .A2(\AES_ENC/us31/n574 ), .ZN(\AES_ENC/us31/n1131 ) );
NAND2_X2 \AES_ENC/us31/U359  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n717 ) );
NAND2_X2 \AES_ENC/us31/U358  ( .A1(\AES_ENC/us31/n1029 ), .A2(\AES_ENC/us31/n717 ), .ZN(\AES_ENC/us31/n728 ) );
NAND2_X2 \AES_ENC/us31/U357  ( .A1(\AES_ENC/sa31 [1]), .A2(\AES_ENC/us31/n624 ), .ZN(\AES_ENC/us31/n1097 ) );
NAND2_X2 \AES_ENC/us31/U356  ( .A1(\AES_ENC/us31/n603 ), .A2(\AES_ENC/us31/n1097 ), .ZN(\AES_ENC/us31/n718 ) );
NAND2_X2 \AES_ENC/us31/U355  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n718 ), .ZN(\AES_ENC/us31/n727 ) );
NAND4_X2 \AES_ENC/us31/U344  ( .A1(\AES_ENC/us31/n728 ), .A2(\AES_ENC/us31/n727 ), .A3(\AES_ENC/us31/n726 ), .A4(\AES_ENC/us31/n725 ), .ZN(\AES_ENC/us31/n729 ) );
NAND2_X2 \AES_ENC/us31/U343  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n729 ), .ZN(\AES_ENC/us31/n730 ) );
NAND4_X2 \AES_ENC/us31/U342  ( .A1(\AES_ENC/us31/n733 ), .A2(\AES_ENC/us31/n732 ), .A3(\AES_ENC/us31/n731 ), .A4(\AES_ENC/us31/n730 ), .ZN(\AES_ENC/sa31_sub[1] ) );
NAND2_X2 \AES_ENC/us31/U341  ( .A1(\AES_ENC/sa31 [7]), .A2(\AES_ENC/us31/n611 ), .ZN(\AES_ENC/us31/n734 ) );
NAND2_X2 \AES_ENC/us31/U340  ( .A1(\AES_ENC/us31/n734 ), .A2(\AES_ENC/us31/n607 ), .ZN(\AES_ENC/us31/n738 ) );
OR4_X2 \AES_ENC/us31/U339  ( .A1(\AES_ENC/us31/n738 ), .A2(\AES_ENC/us31/n626 ), .A3(\AES_ENC/us31/n826 ), .A4(\AES_ENC/us31/n1121 ), .ZN(\AES_ENC/us31/n746 ) );
NAND2_X2 \AES_ENC/us31/U337  ( .A1(\AES_ENC/us31/n1100 ), .A2(\AES_ENC/us31/n587 ), .ZN(\AES_ENC/us31/n992 ) );
OR2_X2 \AES_ENC/us31/U336  ( .A1(\AES_ENC/us31/n610 ), .A2(\AES_ENC/us31/n735 ), .ZN(\AES_ENC/us31/n737 ) );
NAND2_X2 \AES_ENC/us31/U334  ( .A1(\AES_ENC/us31/n619 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n753 ) );
NAND2_X2 \AES_ENC/us31/U333  ( .A1(\AES_ENC/us31/n582 ), .A2(\AES_ENC/us31/n753 ), .ZN(\AES_ENC/us31/n1080 ) );
NAND2_X2 \AES_ENC/us31/U332  ( .A1(\AES_ENC/us31/n1048 ), .A2(\AES_ENC/us31/n576 ), .ZN(\AES_ENC/us31/n736 ) );
NAND2_X2 \AES_ENC/us31/U331  ( .A1(\AES_ENC/us31/n737 ), .A2(\AES_ENC/us31/n736 ), .ZN(\AES_ENC/us31/n739 ) );
NAND2_X2 \AES_ENC/us31/U330  ( .A1(\AES_ENC/us31/n739 ), .A2(\AES_ENC/us31/n738 ), .ZN(\AES_ENC/us31/n745 ) );
NAND2_X2 \AES_ENC/us31/U326  ( .A1(\AES_ENC/us31/n1096 ), .A2(\AES_ENC/us31/n590 ), .ZN(\AES_ENC/us31/n906 ) );
NAND4_X2 \AES_ENC/us31/U323  ( .A1(\AES_ENC/us31/n746 ), .A2(\AES_ENC/us31/n992 ), .A3(\AES_ENC/us31/n745 ), .A4(\AES_ENC/us31/n744 ), .ZN(\AES_ENC/us31/n747 ) );
NAND2_X2 \AES_ENC/us31/U322  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n747 ), .ZN(\AES_ENC/us31/n793 ) );
NAND2_X2 \AES_ENC/us31/U321  ( .A1(\AES_ENC/us31/n584 ), .A2(\AES_ENC/us31/n855 ), .ZN(\AES_ENC/us31/n748 ) );
NAND2_X2 \AES_ENC/us31/U320  ( .A1(\AES_ENC/us31/n956 ), .A2(\AES_ENC/us31/n748 ), .ZN(\AES_ENC/us31/n760 ) );
NAND2_X2 \AES_ENC/us31/U313  ( .A1(\AES_ENC/us31/n590 ), .A2(\AES_ENC/us31/n753 ), .ZN(\AES_ENC/us31/n1023 ) );
NAND4_X2 \AES_ENC/us31/U308  ( .A1(\AES_ENC/us31/n760 ), .A2(\AES_ENC/us31/n992 ), .A3(\AES_ENC/us31/n759 ), .A4(\AES_ENC/us31/n758 ), .ZN(\AES_ENC/us31/n761 ) );
NAND2_X2 \AES_ENC/us31/U307  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n761 ), .ZN(\AES_ENC/us31/n792 ) );
NAND2_X2 \AES_ENC/us31/U306  ( .A1(\AES_ENC/us31/n584 ), .A2(\AES_ENC/us31/n603 ), .ZN(\AES_ENC/us31/n989 ) );
NAND2_X2 \AES_ENC/us31/U305  ( .A1(\AES_ENC/us31/n1050 ), .A2(\AES_ENC/us31/n989 ), .ZN(\AES_ENC/us31/n777 ) );
NAND2_X2 \AES_ENC/us31/U304  ( .A1(\AES_ENC/us31/n1093 ), .A2(\AES_ENC/us31/n762 ), .ZN(\AES_ENC/us31/n776 ) );
XNOR2_X2 \AES_ENC/us31/U301  ( .A(\AES_ENC/sa31 [7]), .B(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n959 ) );
NAND4_X2 \AES_ENC/us31/U289  ( .A1(\AES_ENC/us31/n777 ), .A2(\AES_ENC/us31/n776 ), .A3(\AES_ENC/us31/n775 ), .A4(\AES_ENC/us31/n774 ), .ZN(\AES_ENC/us31/n778 ) );
NAND2_X2 \AES_ENC/us31/U288  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n778 ), .ZN(\AES_ENC/us31/n791 ) );
NAND2_X2 \AES_ENC/us31/U287  ( .A1(\AES_ENC/us31/n1056 ), .A2(\AES_ENC/us31/n1050 ), .ZN(\AES_ENC/us31/n788 ) );
NAND2_X2 \AES_ENC/us31/U286  ( .A1(\AES_ENC/us31/n1091 ), .A2(\AES_ENC/us31/n779 ), .ZN(\AES_ENC/us31/n787 ) );
NAND2_X2 \AES_ENC/us31/U285  ( .A1(\AES_ENC/us31/n956 ), .A2(\AES_ENC/sa31 [1]), .ZN(\AES_ENC/us31/n786 ) );
NAND4_X2 \AES_ENC/us31/U278  ( .A1(\AES_ENC/us31/n788 ), .A2(\AES_ENC/us31/n787 ), .A3(\AES_ENC/us31/n786 ), .A4(\AES_ENC/us31/n785 ), .ZN(\AES_ENC/us31/n789 ) );
NAND2_X2 \AES_ENC/us31/U277  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n789 ), .ZN(\AES_ENC/us31/n790 ) );
NAND4_X2 \AES_ENC/us31/U276  ( .A1(\AES_ENC/us31/n793 ), .A2(\AES_ENC/us31/n792 ), .A3(\AES_ENC/us31/n791 ), .A4(\AES_ENC/us31/n790 ), .ZN(\AES_ENC/sa31_sub[2] ) );
NAND2_X2 \AES_ENC/us31/U275  ( .A1(\AES_ENC/us31/n1059 ), .A2(\AES_ENC/us31/n794 ), .ZN(\AES_ENC/us31/n810 ) );
NAND2_X2 \AES_ENC/us31/U274  ( .A1(\AES_ENC/us31/n1049 ), .A2(\AES_ENC/us31/n956 ), .ZN(\AES_ENC/us31/n809 ) );
OR2_X2 \AES_ENC/us31/U266  ( .A1(\AES_ENC/us31/n1096 ), .A2(\AES_ENC/us31/n606 ), .ZN(\AES_ENC/us31/n802 ) );
NAND2_X2 \AES_ENC/us31/U265  ( .A1(\AES_ENC/us31/n1053 ), .A2(\AES_ENC/us31/n800 ), .ZN(\AES_ENC/us31/n801 ) );
NAND2_X2 \AES_ENC/us31/U264  ( .A1(\AES_ENC/us31/n802 ), .A2(\AES_ENC/us31/n801 ), .ZN(\AES_ENC/us31/n805 ) );
NAND4_X2 \AES_ENC/us31/U261  ( .A1(\AES_ENC/us31/n810 ), .A2(\AES_ENC/us31/n809 ), .A3(\AES_ENC/us31/n808 ), .A4(\AES_ENC/us31/n807 ), .ZN(\AES_ENC/us31/n811 ) );
NAND2_X2 \AES_ENC/us31/U260  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n811 ), .ZN(\AES_ENC/us31/n852 ) );
OR2_X2 \AES_ENC/us31/U259  ( .A1(\AES_ENC/us31/n1023 ), .A2(\AES_ENC/us31/n617 ), .ZN(\AES_ENC/us31/n819 ) );
OR2_X2 \AES_ENC/us31/U257  ( .A1(\AES_ENC/us31/n570 ), .A2(\AES_ENC/us31/n930 ), .ZN(\AES_ENC/us31/n818 ) );
NAND2_X2 \AES_ENC/us31/U256  ( .A1(\AES_ENC/us31/n1013 ), .A2(\AES_ENC/us31/n1094 ), .ZN(\AES_ENC/us31/n817 ) );
NAND4_X2 \AES_ENC/us31/U249  ( .A1(\AES_ENC/us31/n819 ), .A2(\AES_ENC/us31/n818 ), .A3(\AES_ENC/us31/n817 ), .A4(\AES_ENC/us31/n816 ), .ZN(\AES_ENC/us31/n820 ) );
NAND2_X2 \AES_ENC/us31/U248  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n820 ), .ZN(\AES_ENC/us31/n851 ) );
NAND2_X2 \AES_ENC/us31/U247  ( .A1(\AES_ENC/us31/n956 ), .A2(\AES_ENC/us31/n1080 ), .ZN(\AES_ENC/us31/n835 ) );
NAND2_X2 \AES_ENC/us31/U246  ( .A1(\AES_ENC/us31/n570 ), .A2(\AES_ENC/us31/n1030 ), .ZN(\AES_ENC/us31/n1047 ) );
OR2_X2 \AES_ENC/us31/U245  ( .A1(\AES_ENC/us31/n1047 ), .A2(\AES_ENC/us31/n612 ), .ZN(\AES_ENC/us31/n834 ) );
NAND2_X2 \AES_ENC/us31/U244  ( .A1(\AES_ENC/us31/n1072 ), .A2(\AES_ENC/us31/n589 ), .ZN(\AES_ENC/us31/n833 ) );
NAND4_X2 \AES_ENC/us31/U233  ( .A1(\AES_ENC/us31/n835 ), .A2(\AES_ENC/us31/n834 ), .A3(\AES_ENC/us31/n833 ), .A4(\AES_ENC/us31/n832 ), .ZN(\AES_ENC/us31/n836 ) );
NAND2_X2 \AES_ENC/us31/U232  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n836 ), .ZN(\AES_ENC/us31/n850 ) );
NAND2_X2 \AES_ENC/us31/U231  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n623 ), .ZN(\AES_ENC/us31/n847 ) );
NAND2_X2 \AES_ENC/us31/U230  ( .A1(\AES_ENC/us31/n1050 ), .A2(\AES_ENC/us31/n1071 ), .ZN(\AES_ENC/us31/n846 ) );
OR2_X2 \AES_ENC/us31/U224  ( .A1(\AES_ENC/us31/n1053 ), .A2(\AES_ENC/us31/n911 ), .ZN(\AES_ENC/us31/n1077 ) );
NAND4_X2 \AES_ENC/us31/U220  ( .A1(\AES_ENC/us31/n847 ), .A2(\AES_ENC/us31/n846 ), .A3(\AES_ENC/us31/n845 ), .A4(\AES_ENC/us31/n844 ), .ZN(\AES_ENC/us31/n848 ) );
NAND2_X2 \AES_ENC/us31/U219  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n848 ), .ZN(\AES_ENC/us31/n849 ) );
NAND4_X2 \AES_ENC/us31/U218  ( .A1(\AES_ENC/us31/n852 ), .A2(\AES_ENC/us31/n851 ), .A3(\AES_ENC/us31/n850 ), .A4(\AES_ENC/us31/n849 ), .ZN(\AES_ENC/sa31_sub[3] ) );
NAND2_X2 \AES_ENC/us31/U216  ( .A1(\AES_ENC/us31/n1009 ), .A2(\AES_ENC/us31/n1072 ), .ZN(\AES_ENC/us31/n862 ) );
NAND2_X2 \AES_ENC/us31/U215  ( .A1(\AES_ENC/us31/n603 ), .A2(\AES_ENC/us31/n577 ), .ZN(\AES_ENC/us31/n853 ) );
NAND2_X2 \AES_ENC/us31/U214  ( .A1(\AES_ENC/us31/n1050 ), .A2(\AES_ENC/us31/n853 ), .ZN(\AES_ENC/us31/n861 ) );
NAND4_X2 \AES_ENC/us31/U206  ( .A1(\AES_ENC/us31/n862 ), .A2(\AES_ENC/us31/n861 ), .A3(\AES_ENC/us31/n860 ), .A4(\AES_ENC/us31/n859 ), .ZN(\AES_ENC/us31/n863 ) );
NAND2_X2 \AES_ENC/us31/U205  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n863 ), .ZN(\AES_ENC/us31/n905 ) );
NAND2_X2 \AES_ENC/us31/U204  ( .A1(\AES_ENC/us31/n1010 ), .A2(\AES_ENC/us31/n989 ), .ZN(\AES_ENC/us31/n874 ) );
NAND2_X2 \AES_ENC/us31/U203  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n610 ), .ZN(\AES_ENC/us31/n864 ) );
NAND2_X2 \AES_ENC/us31/U202  ( .A1(\AES_ENC/us31/n929 ), .A2(\AES_ENC/us31/n864 ), .ZN(\AES_ENC/us31/n873 ) );
NAND4_X2 \AES_ENC/us31/U193  ( .A1(\AES_ENC/us31/n874 ), .A2(\AES_ENC/us31/n873 ), .A3(\AES_ENC/us31/n872 ), .A4(\AES_ENC/us31/n871 ), .ZN(\AES_ENC/us31/n875 ) );
NAND2_X2 \AES_ENC/us31/U192  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n875 ), .ZN(\AES_ENC/us31/n904 ) );
NAND2_X2 \AES_ENC/us31/U191  ( .A1(\AES_ENC/us31/n583 ), .A2(\AES_ENC/us31/n1050 ), .ZN(\AES_ENC/us31/n889 ) );
NAND2_X2 \AES_ENC/us31/U190  ( .A1(\AES_ENC/us31/n1093 ), .A2(\AES_ENC/us31/n587 ), .ZN(\AES_ENC/us31/n876 ) );
NAND2_X2 \AES_ENC/us31/U189  ( .A1(\AES_ENC/us31/n604 ), .A2(\AES_ENC/us31/n876 ), .ZN(\AES_ENC/us31/n877 ) );
NAND2_X2 \AES_ENC/us31/U188  ( .A1(\AES_ENC/us31/n877 ), .A2(\AES_ENC/us31/n623 ), .ZN(\AES_ENC/us31/n888 ) );
NAND4_X2 \AES_ENC/us31/U179  ( .A1(\AES_ENC/us31/n889 ), .A2(\AES_ENC/us31/n888 ), .A3(\AES_ENC/us31/n887 ), .A4(\AES_ENC/us31/n886 ), .ZN(\AES_ENC/us31/n890 ) );
NAND2_X2 \AES_ENC/us31/U178  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n890 ), .ZN(\AES_ENC/us31/n903 ) );
OR2_X2 \AES_ENC/us31/U177  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n1059 ), .ZN(\AES_ENC/us31/n900 ) );
NAND2_X2 \AES_ENC/us31/U176  ( .A1(\AES_ENC/us31/n1073 ), .A2(\AES_ENC/us31/n1047 ), .ZN(\AES_ENC/us31/n899 ) );
NAND2_X2 \AES_ENC/us31/U175  ( .A1(\AES_ENC/us31/n1094 ), .A2(\AES_ENC/us31/n595 ), .ZN(\AES_ENC/us31/n898 ) );
NAND4_X2 \AES_ENC/us31/U167  ( .A1(\AES_ENC/us31/n900 ), .A2(\AES_ENC/us31/n899 ), .A3(\AES_ENC/us31/n898 ), .A4(\AES_ENC/us31/n897 ), .ZN(\AES_ENC/us31/n901 ) );
NAND2_X2 \AES_ENC/us31/U166  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n901 ), .ZN(\AES_ENC/us31/n902 ) );
NAND4_X2 \AES_ENC/us31/U165  ( .A1(\AES_ENC/us31/n905 ), .A2(\AES_ENC/us31/n904 ), .A3(\AES_ENC/us31/n903 ), .A4(\AES_ENC/us31/n902 ), .ZN(\AES_ENC/sa31_sub[4] ) );
NAND2_X2 \AES_ENC/us31/U164  ( .A1(\AES_ENC/us31/n1094 ), .A2(\AES_ENC/us31/n599 ), .ZN(\AES_ENC/us31/n922 ) );
NAND2_X2 \AES_ENC/us31/U163  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n989 ), .ZN(\AES_ENC/us31/n921 ) );
NAND4_X2 \AES_ENC/us31/U151  ( .A1(\AES_ENC/us31/n922 ), .A2(\AES_ENC/us31/n921 ), .A3(\AES_ENC/us31/n920 ), .A4(\AES_ENC/us31/n919 ), .ZN(\AES_ENC/us31/n923 ) );
NAND2_X2 \AES_ENC/us31/U150  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n923 ), .ZN(\AES_ENC/us31/n972 ) );
NAND2_X2 \AES_ENC/us31/U149  ( .A1(\AES_ENC/us31/n582 ), .A2(\AES_ENC/us31/n619 ), .ZN(\AES_ENC/us31/n924 ) );
NAND2_X2 \AES_ENC/us31/U148  ( .A1(\AES_ENC/us31/n1073 ), .A2(\AES_ENC/us31/n924 ), .ZN(\AES_ENC/us31/n939 ) );
NAND2_X2 \AES_ENC/us31/U147  ( .A1(\AES_ENC/us31/n926 ), .A2(\AES_ENC/us31/n925 ), .ZN(\AES_ENC/us31/n927 ) );
NAND2_X2 \AES_ENC/us31/U146  ( .A1(\AES_ENC/us31/n606 ), .A2(\AES_ENC/us31/n927 ), .ZN(\AES_ENC/us31/n928 ) );
NAND2_X2 \AES_ENC/us31/U145  ( .A1(\AES_ENC/us31/n928 ), .A2(\AES_ENC/us31/n1080 ), .ZN(\AES_ENC/us31/n938 ) );
OR2_X2 \AES_ENC/us31/U144  ( .A1(\AES_ENC/us31/n1117 ), .A2(\AES_ENC/us31/n615 ), .ZN(\AES_ENC/us31/n937 ) );
NAND4_X2 \AES_ENC/us31/U139  ( .A1(\AES_ENC/us31/n939 ), .A2(\AES_ENC/us31/n938 ), .A3(\AES_ENC/us31/n937 ), .A4(\AES_ENC/us31/n936 ), .ZN(\AES_ENC/us31/n940 ) );
NAND2_X2 \AES_ENC/us31/U138  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n940 ), .ZN(\AES_ENC/us31/n971 ) );
OR2_X2 \AES_ENC/us31/U137  ( .A1(\AES_ENC/us31/n605 ), .A2(\AES_ENC/us31/n941 ), .ZN(\AES_ENC/us31/n954 ) );
NAND2_X2 \AES_ENC/us31/U136  ( .A1(\AES_ENC/us31/n1096 ), .A2(\AES_ENC/us31/n577 ), .ZN(\AES_ENC/us31/n942 ) );
NAND2_X2 \AES_ENC/us31/U135  ( .A1(\AES_ENC/us31/n1048 ), .A2(\AES_ENC/us31/n942 ), .ZN(\AES_ENC/us31/n943 ) );
NAND2_X2 \AES_ENC/us31/U134  ( .A1(\AES_ENC/us31/n612 ), .A2(\AES_ENC/us31/n943 ), .ZN(\AES_ENC/us31/n944 ) );
NAND2_X2 \AES_ENC/us31/U133  ( .A1(\AES_ENC/us31/n944 ), .A2(\AES_ENC/us31/n580 ), .ZN(\AES_ENC/us31/n953 ) );
NAND4_X2 \AES_ENC/us31/U125  ( .A1(\AES_ENC/us31/n954 ), .A2(\AES_ENC/us31/n953 ), .A3(\AES_ENC/us31/n952 ), .A4(\AES_ENC/us31/n951 ), .ZN(\AES_ENC/us31/n955 ) );
NAND2_X2 \AES_ENC/us31/U124  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n955 ), .ZN(\AES_ENC/us31/n970 ) );
NAND2_X2 \AES_ENC/us31/U123  ( .A1(\AES_ENC/us31/n1094 ), .A2(\AES_ENC/us31/n1071 ), .ZN(\AES_ENC/us31/n967 ) );
NAND2_X2 \AES_ENC/us31/U122  ( .A1(\AES_ENC/us31/n956 ), .A2(\AES_ENC/us31/n1030 ), .ZN(\AES_ENC/us31/n966 ) );
NAND4_X2 \AES_ENC/us31/U114  ( .A1(\AES_ENC/us31/n967 ), .A2(\AES_ENC/us31/n966 ), .A3(\AES_ENC/us31/n965 ), .A4(\AES_ENC/us31/n964 ), .ZN(\AES_ENC/us31/n968 ) );
NAND2_X2 \AES_ENC/us31/U113  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n968 ), .ZN(\AES_ENC/us31/n969 ) );
NAND4_X2 \AES_ENC/us31/U112  ( .A1(\AES_ENC/us31/n972 ), .A2(\AES_ENC/us31/n971 ), .A3(\AES_ENC/us31/n970 ), .A4(\AES_ENC/us31/n969 ), .ZN(\AES_ENC/sa31_sub[5] ) );
NAND2_X2 \AES_ENC/us31/U111  ( .A1(\AES_ENC/us31/n570 ), .A2(\AES_ENC/us31/n1097 ), .ZN(\AES_ENC/us31/n973 ) );
NAND2_X2 \AES_ENC/us31/U110  ( .A1(\AES_ENC/us31/n1073 ), .A2(\AES_ENC/us31/n973 ), .ZN(\AES_ENC/us31/n987 ) );
NAND2_X2 \AES_ENC/us31/U109  ( .A1(\AES_ENC/us31/n974 ), .A2(\AES_ENC/us31/n1077 ), .ZN(\AES_ENC/us31/n975 ) );
NAND2_X2 \AES_ENC/us31/U108  ( .A1(\AES_ENC/us31/n613 ), .A2(\AES_ENC/us31/n975 ), .ZN(\AES_ENC/us31/n976 ) );
NAND2_X2 \AES_ENC/us31/U107  ( .A1(\AES_ENC/us31/n977 ), .A2(\AES_ENC/us31/n976 ), .ZN(\AES_ENC/us31/n986 ) );
NAND4_X2 \AES_ENC/us31/U99  ( .A1(\AES_ENC/us31/n987 ), .A2(\AES_ENC/us31/n986 ), .A3(\AES_ENC/us31/n985 ), .A4(\AES_ENC/us31/n984 ), .ZN(\AES_ENC/us31/n988 ) );
NAND2_X2 \AES_ENC/us31/U98  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n988 ), .ZN(\AES_ENC/us31/n1044 ) );
NAND2_X2 \AES_ENC/us31/U97  ( .A1(\AES_ENC/us31/n1073 ), .A2(\AES_ENC/us31/n989 ), .ZN(\AES_ENC/us31/n1004 ) );
NAND2_X2 \AES_ENC/us31/U96  ( .A1(\AES_ENC/us31/n1092 ), .A2(\AES_ENC/us31/n619 ), .ZN(\AES_ENC/us31/n1003 ) );
NAND4_X2 \AES_ENC/us31/U85  ( .A1(\AES_ENC/us31/n1004 ), .A2(\AES_ENC/us31/n1003 ), .A3(\AES_ENC/us31/n1002 ), .A4(\AES_ENC/us31/n1001 ), .ZN(\AES_ENC/us31/n1005 ) );
NAND2_X2 \AES_ENC/us31/U84  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n1005 ), .ZN(\AES_ENC/us31/n1043 ) );
NAND2_X2 \AES_ENC/us31/U83  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n596 ), .ZN(\AES_ENC/us31/n1020 ) );
NAND2_X2 \AES_ENC/us31/U82  ( .A1(\AES_ENC/us31/n1050 ), .A2(\AES_ENC/us31/n624 ), .ZN(\AES_ENC/us31/n1019 ) );
NAND2_X2 \AES_ENC/us31/U77  ( .A1(\AES_ENC/us31/n1059 ), .A2(\AES_ENC/us31/n1114 ), .ZN(\AES_ENC/us31/n1012 ) );
NAND2_X2 \AES_ENC/us31/U76  ( .A1(\AES_ENC/us31/n1010 ), .A2(\AES_ENC/us31/n592 ), .ZN(\AES_ENC/us31/n1011 ) );
NAND2_X2 \AES_ENC/us31/U75  ( .A1(\AES_ENC/us31/n1012 ), .A2(\AES_ENC/us31/n1011 ), .ZN(\AES_ENC/us31/n1016 ) );
NAND4_X2 \AES_ENC/us31/U70  ( .A1(\AES_ENC/us31/n1020 ), .A2(\AES_ENC/us31/n1019 ), .A3(\AES_ENC/us31/n1018 ), .A4(\AES_ENC/us31/n1017 ), .ZN(\AES_ENC/us31/n1021 ) );
NAND2_X2 \AES_ENC/us31/U69  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n1021 ), .ZN(\AES_ENC/us31/n1042 ) );
NAND2_X2 \AES_ENC/us31/U68  ( .A1(\AES_ENC/us31/n1022 ), .A2(\AES_ENC/us31/n1093 ), .ZN(\AES_ENC/us31/n1039 ) );
NAND2_X2 \AES_ENC/us31/U67  ( .A1(\AES_ENC/us31/n1050 ), .A2(\AES_ENC/us31/n1023 ), .ZN(\AES_ENC/us31/n1038 ) );
NAND2_X2 \AES_ENC/us31/U66  ( .A1(\AES_ENC/us31/n1024 ), .A2(\AES_ENC/us31/n1071 ), .ZN(\AES_ENC/us31/n1037 ) );
AND2_X2 \AES_ENC/us31/U60  ( .A1(\AES_ENC/us31/n1030 ), .A2(\AES_ENC/us31/n602 ), .ZN(\AES_ENC/us31/n1078 ) );
NAND4_X2 \AES_ENC/us31/U56  ( .A1(\AES_ENC/us31/n1039 ), .A2(\AES_ENC/us31/n1038 ), .A3(\AES_ENC/us31/n1037 ), .A4(\AES_ENC/us31/n1036 ), .ZN(\AES_ENC/us31/n1040 ) );
NAND2_X2 \AES_ENC/us31/U55  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n1040 ), .ZN(\AES_ENC/us31/n1041 ) );
NAND4_X2 \AES_ENC/us31/U54  ( .A1(\AES_ENC/us31/n1044 ), .A2(\AES_ENC/us31/n1043 ), .A3(\AES_ENC/us31/n1042 ), .A4(\AES_ENC/us31/n1041 ), .ZN(\AES_ENC/sa31_sub[6] ) );
NAND2_X2 \AES_ENC/us31/U53  ( .A1(\AES_ENC/us31/n1072 ), .A2(\AES_ENC/us31/n1045 ), .ZN(\AES_ENC/us31/n1068 ) );
NAND2_X2 \AES_ENC/us31/U52  ( .A1(\AES_ENC/us31/n1046 ), .A2(\AES_ENC/us31/n582 ), .ZN(\AES_ENC/us31/n1067 ) );
NAND2_X2 \AES_ENC/us31/U51  ( .A1(\AES_ENC/us31/n1094 ), .A2(\AES_ENC/us31/n1047 ), .ZN(\AES_ENC/us31/n1066 ) );
NAND4_X2 \AES_ENC/us31/U40  ( .A1(\AES_ENC/us31/n1068 ), .A2(\AES_ENC/us31/n1067 ), .A3(\AES_ENC/us31/n1066 ), .A4(\AES_ENC/us31/n1065 ), .ZN(\AES_ENC/us31/n1069 ) );
NAND2_X2 \AES_ENC/us31/U39  ( .A1(\AES_ENC/us31/n1070 ), .A2(\AES_ENC/us31/n1069 ), .ZN(\AES_ENC/us31/n1135 ) );
NAND2_X2 \AES_ENC/us31/U38  ( .A1(\AES_ENC/us31/n1072 ), .A2(\AES_ENC/us31/n1071 ), .ZN(\AES_ENC/us31/n1088 ) );
NAND2_X2 \AES_ENC/us31/U37  ( .A1(\AES_ENC/us31/n1073 ), .A2(\AES_ENC/us31/n595 ), .ZN(\AES_ENC/us31/n1087 ) );
NAND4_X2 \AES_ENC/us31/U28  ( .A1(\AES_ENC/us31/n1088 ), .A2(\AES_ENC/us31/n1087 ), .A3(\AES_ENC/us31/n1086 ), .A4(\AES_ENC/us31/n1085 ), .ZN(\AES_ENC/us31/n1089 ) );
NAND2_X2 \AES_ENC/us31/U27  ( .A1(\AES_ENC/us31/n1090 ), .A2(\AES_ENC/us31/n1089 ), .ZN(\AES_ENC/us31/n1134 ) );
NAND2_X2 \AES_ENC/us31/U26  ( .A1(\AES_ENC/us31/n1091 ), .A2(\AES_ENC/us31/n1093 ), .ZN(\AES_ENC/us31/n1111 ) );
NAND2_X2 \AES_ENC/us31/U25  ( .A1(\AES_ENC/us31/n1092 ), .A2(\AES_ENC/us31/n1120 ), .ZN(\AES_ENC/us31/n1110 ) );
AND2_X2 \AES_ENC/us31/U22  ( .A1(\AES_ENC/us31/n1097 ), .A2(\AES_ENC/us31/n1096 ), .ZN(\AES_ENC/us31/n1098 ) );
NAND4_X2 \AES_ENC/us31/U14  ( .A1(\AES_ENC/us31/n1111 ), .A2(\AES_ENC/us31/n1110 ), .A3(\AES_ENC/us31/n1109 ), .A4(\AES_ENC/us31/n1108 ), .ZN(\AES_ENC/us31/n1112 ) );
NAND2_X2 \AES_ENC/us31/U13  ( .A1(\AES_ENC/us31/n1113 ), .A2(\AES_ENC/us31/n1112 ), .ZN(\AES_ENC/us31/n1133 ) );
NAND2_X2 \AES_ENC/us31/U12  ( .A1(\AES_ENC/us31/n1115 ), .A2(\AES_ENC/us31/n1114 ), .ZN(\AES_ENC/us31/n1129 ) );
OR2_X2 \AES_ENC/us31/U11  ( .A1(\AES_ENC/us31/n608 ), .A2(\AES_ENC/us31/n1116 ), .ZN(\AES_ENC/us31/n1128 ) );
NAND4_X2 \AES_ENC/us31/U3  ( .A1(\AES_ENC/us31/n1129 ), .A2(\AES_ENC/us31/n1128 ), .A3(\AES_ENC/us31/n1127 ), .A4(\AES_ENC/us31/n1126 ), .ZN(\AES_ENC/us31/n1130 ) );
NAND2_X2 \AES_ENC/us31/U2  ( .A1(\AES_ENC/us31/n1131 ), .A2(\AES_ENC/us31/n1130 ), .ZN(\AES_ENC/us31/n1132 ) );
NAND4_X2 \AES_ENC/us31/U1  ( .A1(\AES_ENC/us31/n1135 ), .A2(\AES_ENC/us31/n1134 ), .A3(\AES_ENC/us31/n1133 ), .A4(\AES_ENC/us31/n1132 ), .ZN(\AES_ENC/sa31_sub[7] ) );
INV_X4 \AES_ENC/us32/U575  ( .A(\AES_ENC/sa32 [7]), .ZN(\AES_ENC/us32/n627 ));
INV_X4 \AES_ENC/us32/U574  ( .A(\AES_ENC/us32/n1114 ), .ZN(\AES_ENC/us32/n625 ) );
INV_X4 \AES_ENC/us32/U573  ( .A(\AES_ENC/sa32 [4]), .ZN(\AES_ENC/us32/n624 ));
INV_X4 \AES_ENC/us32/U572  ( .A(\AES_ENC/us32/n1025 ), .ZN(\AES_ENC/us32/n622 ) );
INV_X4 \AES_ENC/us32/U571  ( .A(\AES_ENC/us32/n1120 ), .ZN(\AES_ENC/us32/n620 ) );
INV_X4 \AES_ENC/us32/U570  ( .A(\AES_ENC/us32/n1121 ), .ZN(\AES_ENC/us32/n619 ) );
INV_X4 \AES_ENC/us32/U569  ( .A(\AES_ENC/us32/n1048 ), .ZN(\AES_ENC/us32/n618 ) );
INV_X4 \AES_ENC/us32/U568  ( .A(\AES_ENC/us32/n974 ), .ZN(\AES_ENC/us32/n616 ) );
INV_X4 \AES_ENC/us32/U567  ( .A(\AES_ENC/us32/n794 ), .ZN(\AES_ENC/us32/n614 ) );
INV_X4 \AES_ENC/us32/U566  ( .A(\AES_ENC/sa32 [2]), .ZN(\AES_ENC/us32/n611 ));
INV_X4 \AES_ENC/us32/U565  ( .A(\AES_ENC/us32/n800 ), .ZN(\AES_ENC/us32/n610 ) );
INV_X4 \AES_ENC/us32/U564  ( .A(\AES_ENC/us32/n925 ), .ZN(\AES_ENC/us32/n609 ) );
INV_X4 \AES_ENC/us32/U563  ( .A(\AES_ENC/us32/n779 ), .ZN(\AES_ENC/us32/n607 ) );
INV_X4 \AES_ENC/us32/U562  ( .A(\AES_ENC/us32/n1022 ), .ZN(\AES_ENC/us32/n603 ) );
INV_X4 \AES_ENC/us32/U561  ( .A(\AES_ENC/us32/n1102 ), .ZN(\AES_ENC/us32/n602 ) );
INV_X4 \AES_ENC/us32/U560  ( .A(\AES_ENC/us32/n929 ), .ZN(\AES_ENC/us32/n601 ) );
INV_X4 \AES_ENC/us32/U559  ( .A(\AES_ENC/us32/n1056 ), .ZN(\AES_ENC/us32/n600 ) );
INV_X4 \AES_ENC/us32/U558  ( .A(\AES_ENC/us32/n1054 ), .ZN(\AES_ENC/us32/n599 ) );
INV_X4 \AES_ENC/us32/U557  ( .A(\AES_ENC/us32/n881 ), .ZN(\AES_ENC/us32/n598 ) );
INV_X4 \AES_ENC/us32/U556  ( .A(\AES_ENC/us32/n926 ), .ZN(\AES_ENC/us32/n597 ) );
INV_X4 \AES_ENC/us32/U555  ( .A(\AES_ENC/us32/n977 ), .ZN(\AES_ENC/us32/n595 ) );
INV_X4 \AES_ENC/us32/U554  ( .A(\AES_ENC/us32/n1031 ), .ZN(\AES_ENC/us32/n594 ) );
INV_X4 \AES_ENC/us32/U553  ( .A(\AES_ENC/us32/n1103 ), .ZN(\AES_ENC/us32/n593 ) );
INV_X4 \AES_ENC/us32/U552  ( .A(\AES_ENC/us32/n1009 ), .ZN(\AES_ENC/us32/n592 ) );
INV_X4 \AES_ENC/us32/U551  ( .A(\AES_ENC/us32/n990 ), .ZN(\AES_ENC/us32/n591 ) );
INV_X4 \AES_ENC/us32/U550  ( .A(\AES_ENC/us32/n1058 ), .ZN(\AES_ENC/us32/n590 ) );
INV_X4 \AES_ENC/us32/U549  ( .A(\AES_ENC/us32/n1074 ), .ZN(\AES_ENC/us32/n589 ) );
INV_X4 \AES_ENC/us32/U548  ( .A(\AES_ENC/us32/n1053 ), .ZN(\AES_ENC/us32/n588 ) );
INV_X4 \AES_ENC/us32/U547  ( .A(\AES_ENC/us32/n826 ), .ZN(\AES_ENC/us32/n587 ) );
INV_X4 \AES_ENC/us32/U546  ( .A(\AES_ENC/us32/n992 ), .ZN(\AES_ENC/us32/n586 ) );
INV_X4 \AES_ENC/us32/U545  ( .A(\AES_ENC/us32/n821 ), .ZN(\AES_ENC/us32/n585 ) );
INV_X4 \AES_ENC/us32/U544  ( .A(\AES_ENC/us32/n910 ), .ZN(\AES_ENC/us32/n584 ) );
INV_X4 \AES_ENC/us32/U543  ( .A(\AES_ENC/us32/n906 ), .ZN(\AES_ENC/us32/n583 ) );
INV_X4 \AES_ENC/us32/U542  ( .A(\AES_ENC/us32/n880 ), .ZN(\AES_ENC/us32/n581 ) );
INV_X4 \AES_ENC/us32/U541  ( .A(\AES_ENC/us32/n1013 ), .ZN(\AES_ENC/us32/n580 ) );
INV_X4 \AES_ENC/us32/U540  ( .A(\AES_ENC/us32/n1092 ), .ZN(\AES_ENC/us32/n579 ) );
INV_X4 \AES_ENC/us32/U539  ( .A(\AES_ENC/us32/n824 ), .ZN(\AES_ENC/us32/n578 ) );
INV_X4 \AES_ENC/us32/U538  ( .A(\AES_ENC/us32/n1091 ), .ZN(\AES_ENC/us32/n577 ) );
INV_X4 \AES_ENC/us32/U537  ( .A(\AES_ENC/us32/n1080 ), .ZN(\AES_ENC/us32/n576 ) );
INV_X4 \AES_ENC/us32/U536  ( .A(\AES_ENC/us32/n959 ), .ZN(\AES_ENC/us32/n575 ) );
INV_X4 \AES_ENC/us32/U535  ( .A(\AES_ENC/sa32 [0]), .ZN(\AES_ENC/us32/n574 ));
NOR2_X2 \AES_ENC/us32/U534  ( .A1(\AES_ENC/sa32 [0]), .A2(\AES_ENC/sa32 [6]),.ZN(\AES_ENC/us32/n1090 ) );
NOR2_X2 \AES_ENC/us32/U533  ( .A1(\AES_ENC/us32/n574 ), .A2(\AES_ENC/sa32 [6]), .ZN(\AES_ENC/us32/n1070 ) );
NOR2_X2 \AES_ENC/us32/U532  ( .A1(\AES_ENC/sa32 [4]), .A2(\AES_ENC/sa32 [3]),.ZN(\AES_ENC/us32/n1025 ) );
INV_X4 \AES_ENC/us32/U531  ( .A(\AES_ENC/us32/n569 ), .ZN(\AES_ENC/us32/n572 ) );
NOR2_X2 \AES_ENC/us32/U530  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n765 ) );
NOR2_X2 \AES_ENC/us32/U529  ( .A1(\AES_ENC/sa32 [4]), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n764 ) );
NOR2_X2 \AES_ENC/us32/U528  ( .A1(\AES_ENC/us32/n765 ), .A2(\AES_ENC/us32/n764 ), .ZN(\AES_ENC/us32/n766 ) );
NOR2_X2 \AES_ENC/us32/U527  ( .A1(\AES_ENC/us32/n766 ), .A2(\AES_ENC/us32/n575 ), .ZN(\AES_ENC/us32/n767 ) );
INV_X4 \AES_ENC/us32/U526  ( .A(\AES_ENC/sa32 [3]), .ZN(\AES_ENC/us32/n621 ));
NAND3_X2 \AES_ENC/us32/U525  ( .A1(\AES_ENC/us32/n652 ), .A2(\AES_ENC/us32/n626 ), .A3(\AES_ENC/sa32 [7]), .ZN(\AES_ENC/us32/n653 ));
NOR2_X2 \AES_ENC/us32/U524  ( .A1(\AES_ENC/us32/n611 ), .A2(\AES_ENC/sa32 [5]), .ZN(\AES_ENC/us32/n925 ) );
NOR2_X2 \AES_ENC/us32/U523  ( .A1(\AES_ENC/sa32 [5]), .A2(\AES_ENC/sa32 [2]),.ZN(\AES_ENC/us32/n974 ) );
INV_X4 \AES_ENC/us32/U522  ( .A(\AES_ENC/sa32 [5]), .ZN(\AES_ENC/us32/n626 ));
NOR2_X2 \AES_ENC/us32/U521  ( .A1(\AES_ENC/us32/n611 ), .A2(\AES_ENC/sa32 [7]), .ZN(\AES_ENC/us32/n779 ) );
NAND3_X2 \AES_ENC/us32/U520  ( .A1(\AES_ENC/us32/n679 ), .A2(\AES_ENC/us32/n678 ), .A3(\AES_ENC/us32/n677 ), .ZN(\AES_ENC/sa32_sub[0] ) );
NOR2_X2 \AES_ENC/us32/U519  ( .A1(\AES_ENC/us32/n626 ), .A2(\AES_ENC/sa32 [2]), .ZN(\AES_ENC/us32/n1048 ) );
NOR3_X2 \AES_ENC/us32/U518  ( .A1(\AES_ENC/us32/n627 ), .A2(\AES_ENC/sa32 [5]), .A3(\AES_ENC/us32/n704 ), .ZN(\AES_ENC/us32/n706 ));
NOR2_X2 \AES_ENC/us32/U517  ( .A1(\AES_ENC/us32/n1117 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n707 ) );
NOR2_X2 \AES_ENC/us32/U516  ( .A1(\AES_ENC/sa32 [4]), .A2(\AES_ENC/us32/n579 ), .ZN(\AES_ENC/us32/n705 ) );
NOR3_X2 \AES_ENC/us32/U515  ( .A1(\AES_ENC/us32/n707 ), .A2(\AES_ENC/us32/n706 ), .A3(\AES_ENC/us32/n705 ), .ZN(\AES_ENC/us32/n713 ) );
NOR4_X2 \AES_ENC/us32/U512  ( .A1(\AES_ENC/us32/n633 ), .A2(\AES_ENC/us32/n632 ), .A3(\AES_ENC/us32/n631 ), .A4(\AES_ENC/us32/n630 ), .ZN(\AES_ENC/us32/n634 ) );
NOR2_X2 \AES_ENC/us32/U510  ( .A1(\AES_ENC/us32/n629 ), .A2(\AES_ENC/us32/n628 ), .ZN(\AES_ENC/us32/n635 ) );
NAND3_X2 \AES_ENC/us32/U509  ( .A1(\AES_ENC/sa32 [2]), .A2(\AES_ENC/sa32 [7]), .A3(\AES_ENC/us32/n1059 ), .ZN(\AES_ENC/us32/n636 ) );
NOR2_X2 \AES_ENC/us32/U508  ( .A1(\AES_ENC/sa32 [7]), .A2(\AES_ENC/sa32 [2]),.ZN(\AES_ENC/us32/n794 ) );
NOR2_X2 \AES_ENC/us32/U507  ( .A1(\AES_ENC/sa32 [4]), .A2(\AES_ENC/sa32 [1]),.ZN(\AES_ENC/us32/n1102 ) );
NOR2_X2 \AES_ENC/us32/U506  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/sa32 [3]), .ZN(\AES_ENC/us32/n1053 ) );
NOR2_X2 \AES_ENC/us32/U505  ( .A1(\AES_ENC/us32/n607 ), .A2(\AES_ENC/sa32 [5]), .ZN(\AES_ENC/us32/n1024 ) );
NOR2_X2 \AES_ENC/us32/U504  ( .A1(\AES_ENC/us32/n625 ), .A2(\AES_ENC/sa32 [2]), .ZN(\AES_ENC/us32/n1093 ) );
NOR2_X2 \AES_ENC/us32/U503  ( .A1(\AES_ENC/us32/n614 ), .A2(\AES_ENC/sa32 [5]), .ZN(\AES_ENC/us32/n1094 ) );
NOR2_X2 \AES_ENC/us32/U502  ( .A1(\AES_ENC/us32/n624 ), .A2(\AES_ENC/sa32 [3]), .ZN(\AES_ENC/us32/n931 ) );
INV_X4 \AES_ENC/us32/U501  ( .A(\AES_ENC/us32/n570 ), .ZN(\AES_ENC/us32/n573 ) );
NOR2_X2 \AES_ENC/us32/U500  ( .A1(\AES_ENC/us32/n1053 ), .A2(\AES_ENC/us32/n1095 ), .ZN(\AES_ENC/us32/n639 ) );
NOR3_X2 \AES_ENC/us32/U499  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n573 ), .A3(\AES_ENC/us32/n1074 ), .ZN(\AES_ENC/us32/n641 ) );
NOR2_X2 \AES_ENC/us32/U498  ( .A1(\AES_ENC/us32/n639 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n640 ) );
NOR2_X2 \AES_ENC/us32/U497  ( .A1(\AES_ENC/us32/n641 ), .A2(\AES_ENC/us32/n640 ), .ZN(\AES_ENC/us32/n646 ) );
NOR3_X2 \AES_ENC/us32/U496  ( .A1(\AES_ENC/us32/n995 ), .A2(\AES_ENC/us32/n586 ), .A3(\AES_ENC/us32/n994 ), .ZN(\AES_ENC/us32/n1002 ) );
NOR2_X2 \AES_ENC/us32/U495  ( .A1(\AES_ENC/us32/n909 ), .A2(\AES_ENC/us32/n908 ), .ZN(\AES_ENC/us32/n920 ) );
NOR2_X2 \AES_ENC/us32/U494  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n823 ) );
NOR2_X2 \AES_ENC/us32/U492  ( .A1(\AES_ENC/us32/n624 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n822 ) );
NOR2_X2 \AES_ENC/us32/U491  ( .A1(\AES_ENC/us32/n823 ), .A2(\AES_ENC/us32/n822 ), .ZN(\AES_ENC/us32/n825 ) );
NOR2_X2 \AES_ENC/us32/U490  ( .A1(\AES_ENC/sa32 [1]), .A2(\AES_ENC/us32/n623 ), .ZN(\AES_ENC/us32/n913 ) );
NOR2_X2 \AES_ENC/us32/U489  ( .A1(\AES_ENC/us32/n913 ), .A2(\AES_ENC/us32/n1091 ), .ZN(\AES_ENC/us32/n914 ) );
NOR2_X2 \AES_ENC/us32/U488  ( .A1(\AES_ENC/us32/n826 ), .A2(\AES_ENC/us32/n572 ), .ZN(\AES_ENC/us32/n827 ) );
NOR3_X2 \AES_ENC/us32/U487  ( .A1(\AES_ENC/us32/n769 ), .A2(\AES_ENC/us32/n768 ), .A3(\AES_ENC/us32/n767 ), .ZN(\AES_ENC/us32/n775 ) );
NOR2_X2 \AES_ENC/us32/U486  ( .A1(\AES_ENC/us32/n1056 ), .A2(\AES_ENC/us32/n1053 ), .ZN(\AES_ENC/us32/n749 ) );
NOR2_X2 \AES_ENC/us32/U483  ( .A1(\AES_ENC/us32/n749 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n752 ) );
INV_X4 \AES_ENC/us32/U482  ( .A(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n596 ));
NOR2_X2 \AES_ENC/us32/U480  ( .A1(\AES_ENC/us32/n1054 ), .A2(\AES_ENC/us32/n1053 ), .ZN(\AES_ENC/us32/n1055 ) );
OR2_X4 \AES_ENC/us32/U479  ( .A1(\AES_ENC/us32/n1094 ), .A2(\AES_ENC/us32/n1093 ), .ZN(\AES_ENC/us32/n571 ) );
AND2_X2 \AES_ENC/us32/U478  ( .A1(\AES_ENC/us32/n571 ), .A2(\AES_ENC/us32/n1095 ), .ZN(\AES_ENC/us32/n1101 ) );
NOR2_X2 \AES_ENC/us32/U477  ( .A1(\AES_ENC/us32/n1074 ), .A2(\AES_ENC/us32/n931 ), .ZN(\AES_ENC/us32/n796 ) );
NOR2_X2 \AES_ENC/us32/U474  ( .A1(\AES_ENC/us32/n796 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n797 ) );
NOR2_X2 \AES_ENC/us32/U473  ( .A1(\AES_ENC/us32/n932 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n933 ) );
NOR2_X2 \AES_ENC/us32/U472  ( .A1(\AES_ENC/us32/n929 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n935 ) );
NOR2_X2 \AES_ENC/us32/U471  ( .A1(\AES_ENC/us32/n931 ), .A2(\AES_ENC/us32/n930 ), .ZN(\AES_ENC/us32/n934 ) );
NOR3_X2 \AES_ENC/us32/U470  ( .A1(\AES_ENC/us32/n935 ), .A2(\AES_ENC/us32/n934 ), .A3(\AES_ENC/us32/n933 ), .ZN(\AES_ENC/us32/n936 ) );
NOR2_X2 \AES_ENC/us32/U469  ( .A1(\AES_ENC/us32/n624 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n1075 ) );
NOR2_X2 \AES_ENC/us32/U468  ( .A1(\AES_ENC/us32/n572 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n949 ) );
NOR2_X2 \AES_ENC/us32/U467  ( .A1(\AES_ENC/us32/n1049 ), .A2(\AES_ENC/us32/n618 ), .ZN(\AES_ENC/us32/n1051 ) );
NOR2_X2 \AES_ENC/us32/U466  ( .A1(\AES_ENC/us32/n1051 ), .A2(\AES_ENC/us32/n1050 ), .ZN(\AES_ENC/us32/n1052 ) );
NOR2_X2 \AES_ENC/us32/U465  ( .A1(\AES_ENC/us32/n1052 ), .A2(\AES_ENC/us32/n592 ), .ZN(\AES_ENC/us32/n1064 ) );
NOR2_X2 \AES_ENC/us32/U464  ( .A1(\AES_ENC/sa32 [1]), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n631 ) );
NOR2_X2 \AES_ENC/us32/U463  ( .A1(\AES_ENC/us32/n1025 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n980 ) );
NOR2_X2 \AES_ENC/us32/U462  ( .A1(\AES_ENC/us32/n1073 ), .A2(\AES_ENC/us32/n1094 ), .ZN(\AES_ENC/us32/n795 ) );
NOR2_X2 \AES_ENC/us32/U461  ( .A1(\AES_ENC/us32/n795 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n799 ) );
NOR2_X2 \AES_ENC/us32/U460  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n981 ) );
NOR2_X2 \AES_ENC/us32/U459  ( .A1(\AES_ENC/us32/n1102 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n643 ) );
NOR2_X2 \AES_ENC/us32/U458  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n621 ), .ZN(\AES_ENC/us32/n642 ) );
NOR2_X2 \AES_ENC/us32/U455  ( .A1(\AES_ENC/us32/n911 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n644 ) );
NOR4_X2 \AES_ENC/us32/U448  ( .A1(\AES_ENC/us32/n644 ), .A2(\AES_ENC/us32/n643 ), .A3(\AES_ENC/us32/n804 ), .A4(\AES_ENC/us32/n642 ), .ZN(\AES_ENC/us32/n645 ) );
NOR2_X2 \AES_ENC/us32/U447  ( .A1(\AES_ENC/us32/n1102 ), .A2(\AES_ENC/us32/n910 ), .ZN(\AES_ENC/us32/n932 ) );
NOR2_X2 \AES_ENC/us32/U442  ( .A1(\AES_ENC/us32/n1102 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n755 ) );
NOR2_X2 \AES_ENC/us32/U441  ( .A1(\AES_ENC/us32/n931 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n743 ) );
NOR2_X2 \AES_ENC/us32/U438  ( .A1(\AES_ENC/us32/n1072 ), .A2(\AES_ENC/us32/n1094 ), .ZN(\AES_ENC/us32/n930 ) );
NOR2_X2 \AES_ENC/us32/U435  ( .A1(\AES_ENC/us32/n1074 ), .A2(\AES_ENC/us32/n1025 ), .ZN(\AES_ENC/us32/n891 ) );
NOR2_X2 \AES_ENC/us32/U434  ( .A1(\AES_ENC/us32/n891 ), .A2(\AES_ENC/us32/n609 ), .ZN(\AES_ENC/us32/n894 ) );
NOR3_X2 \AES_ENC/us32/U433  ( .A1(\AES_ENC/us32/n623 ), .A2(\AES_ENC/sa32 [1]), .A3(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n683 ));
INV_X4 \AES_ENC/us32/U428  ( .A(\AES_ENC/us32/n931 ), .ZN(\AES_ENC/us32/n623 ) );
NOR2_X2 \AES_ENC/us32/U427  ( .A1(\AES_ENC/us32/n996 ), .A2(\AES_ENC/us32/n931 ), .ZN(\AES_ENC/us32/n704 ) );
NOR2_X2 \AES_ENC/us32/U421  ( .A1(\AES_ENC/us32/n931 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n685 ) );
NOR2_X2 \AES_ENC/us32/U420  ( .A1(\AES_ENC/us32/n1029 ), .A2(\AES_ENC/us32/n1025 ), .ZN(\AES_ENC/us32/n1079 ) );
NOR3_X2 \AES_ENC/us32/U419  ( .A1(\AES_ENC/us32/n589 ), .A2(\AES_ENC/us32/n1025 ), .A3(\AES_ENC/us32/n616 ), .ZN(\AES_ENC/us32/n945 ) );
NOR2_X2 \AES_ENC/us32/U418  ( .A1(\AES_ENC/us32/n626 ), .A2(\AES_ENC/us32/n611 ), .ZN(\AES_ENC/us32/n800 ) );
NOR3_X2 \AES_ENC/us32/U417  ( .A1(\AES_ENC/us32/n590 ), .A2(\AES_ENC/us32/n627 ), .A3(\AES_ENC/us32/n611 ), .ZN(\AES_ENC/us32/n798 ) );
NOR3_X2 \AES_ENC/us32/U416  ( .A1(\AES_ENC/us32/n610 ), .A2(\AES_ENC/us32/n572 ), .A3(\AES_ENC/us32/n575 ), .ZN(\AES_ENC/us32/n962 ) );
NOR3_X2 \AES_ENC/us32/U415  ( .A1(\AES_ENC/us32/n959 ), .A2(\AES_ENC/us32/n572 ), .A3(\AES_ENC/us32/n609 ), .ZN(\AES_ENC/us32/n768 ) );
NOR3_X2 \AES_ENC/us32/U414  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n572 ), .A3(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n694 ) );
NOR3_X2 \AES_ENC/us32/U413  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n572 ), .A3(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n895 ) );
NOR3_X2 \AES_ENC/us32/U410  ( .A1(\AES_ENC/us32/n1008 ), .A2(\AES_ENC/us32/n1007 ), .A3(\AES_ENC/us32/n1006 ), .ZN(\AES_ENC/us32/n1018 ) );
NOR4_X2 \AES_ENC/us32/U409  ( .A1(\AES_ENC/us32/n806 ), .A2(\AES_ENC/us32/n805 ), .A3(\AES_ENC/us32/n804 ), .A4(\AES_ENC/us32/n803 ), .ZN(\AES_ENC/us32/n807 ) );
NOR3_X2 \AES_ENC/us32/U406  ( .A1(\AES_ENC/us32/n799 ), .A2(\AES_ENC/us32/n798 ), .A3(\AES_ENC/us32/n797 ), .ZN(\AES_ENC/us32/n808 ) );
NOR4_X2 \AES_ENC/us32/U405  ( .A1(\AES_ENC/us32/n843 ), .A2(\AES_ENC/us32/n842 ), .A3(\AES_ENC/us32/n841 ), .A4(\AES_ENC/us32/n840 ), .ZN(\AES_ENC/us32/n844 ) );
NOR3_X2 \AES_ENC/us32/U404  ( .A1(\AES_ENC/us32/n1101 ), .A2(\AES_ENC/us32/n1100 ), .A3(\AES_ENC/us32/n1099 ), .ZN(\AES_ENC/us32/n1109 ) );
NOR4_X2 \AES_ENC/us32/U403  ( .A1(\AES_ENC/us32/n711 ), .A2(\AES_ENC/us32/n710 ), .A3(\AES_ENC/us32/n709 ), .A4(\AES_ENC/us32/n708 ), .ZN(\AES_ENC/us32/n712 ) );
NOR4_X2 \AES_ENC/us32/U401  ( .A1(\AES_ENC/us32/n963 ), .A2(\AES_ENC/us32/n962 ), .A3(\AES_ENC/us32/n961 ), .A4(\AES_ENC/us32/n960 ), .ZN(\AES_ENC/us32/n964 ) );
NOR2_X2 \AES_ENC/us32/U400  ( .A1(\AES_ENC/us32/n669 ), .A2(\AES_ENC/us32/n668 ), .ZN(\AES_ENC/us32/n673 ) );
NOR4_X2 \AES_ENC/us32/U399  ( .A1(\AES_ENC/us32/n946 ), .A2(\AES_ENC/us32/n1046 ), .A3(\AES_ENC/us32/n671 ), .A4(\AES_ENC/us32/n670 ), .ZN(\AES_ENC/us32/n672 ) );
NOR3_X2 \AES_ENC/us32/U398  ( .A1(\AES_ENC/us32/n743 ), .A2(\AES_ENC/us32/n742 ), .A3(\AES_ENC/us32/n741 ), .ZN(\AES_ENC/us32/n744 ) );
NOR2_X2 \AES_ENC/us32/U397  ( .A1(\AES_ENC/us32/n697 ), .A2(\AES_ENC/us32/n658 ), .ZN(\AES_ENC/us32/n659 ) );
NOR2_X2 \AES_ENC/us32/U396  ( .A1(\AES_ENC/us32/n1078 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n1033 ) );
NOR2_X2 \AES_ENC/us32/U393  ( .A1(\AES_ENC/us32/n1031 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n1032 ) );
NOR3_X2 \AES_ENC/us32/U390  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n1025 ), .A3(\AES_ENC/us32/n1074 ), .ZN(\AES_ENC/us32/n1035 ) );
NOR4_X2 \AES_ENC/us32/U389  ( .A1(\AES_ENC/us32/n1035 ), .A2(\AES_ENC/us32/n1034 ), .A3(\AES_ENC/us32/n1033 ), .A4(\AES_ENC/us32/n1032 ), .ZN(\AES_ENC/us32/n1036 ) );
NOR2_X2 \AES_ENC/us32/U388  ( .A1(\AES_ENC/us32/n598 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n885 ) );
NOR2_X2 \AES_ENC/us32/U387  ( .A1(\AES_ENC/us32/n623 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n882 ) );
NOR2_X2 \AES_ENC/us32/U386  ( .A1(\AES_ENC/us32/n1053 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n884 ) );
NOR4_X2 \AES_ENC/us32/U385  ( .A1(\AES_ENC/us32/n885 ), .A2(\AES_ENC/us32/n884 ), .A3(\AES_ENC/us32/n883 ), .A4(\AES_ENC/us32/n882 ), .ZN(\AES_ENC/us32/n886 ) );
NOR2_X2 \AES_ENC/us32/U384  ( .A1(\AES_ENC/us32/n825 ), .A2(\AES_ENC/us32/n578 ), .ZN(\AES_ENC/us32/n830 ) );
NOR2_X2 \AES_ENC/us32/U383  ( .A1(\AES_ENC/us32/n827 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n829 ) );
NOR2_X2 \AES_ENC/us32/U382  ( .A1(\AES_ENC/us32/n572 ), .A2(\AES_ENC/us32/n579 ), .ZN(\AES_ENC/us32/n828 ) );
NOR4_X2 \AES_ENC/us32/U374  ( .A1(\AES_ENC/us32/n831 ), .A2(\AES_ENC/us32/n830 ), .A3(\AES_ENC/us32/n829 ), .A4(\AES_ENC/us32/n828 ), .ZN(\AES_ENC/us32/n832 ) );
NOR2_X2 \AES_ENC/us32/U373  ( .A1(\AES_ENC/us32/n606 ), .A2(\AES_ENC/us32/n582 ), .ZN(\AES_ENC/us32/n1104 ) );
NOR2_X2 \AES_ENC/us32/U372  ( .A1(\AES_ENC/us32/n1102 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n1106 ) );
NOR2_X2 \AES_ENC/us32/U370  ( .A1(\AES_ENC/us32/n1103 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n1105 ) );
NOR4_X2 \AES_ENC/us32/U369  ( .A1(\AES_ENC/us32/n1107 ), .A2(\AES_ENC/us32/n1106 ), .A3(\AES_ENC/us32/n1105 ), .A4(\AES_ENC/us32/n1104 ), .ZN(\AES_ENC/us32/n1108 ) );
NOR3_X2 \AES_ENC/us32/U368  ( .A1(\AES_ENC/us32/n959 ), .A2(\AES_ENC/us32/n621 ), .A3(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n963 ) );
NOR2_X2 \AES_ENC/us32/U367  ( .A1(\AES_ENC/us32/n626 ), .A2(\AES_ENC/us32/n627 ), .ZN(\AES_ENC/us32/n1114 ) );
INV_X4 \AES_ENC/us32/U366  ( .A(\AES_ENC/us32/n1024 ), .ZN(\AES_ENC/us32/n606 ) );
NOR3_X2 \AES_ENC/us32/U365  ( .A1(\AES_ENC/us32/n910 ), .A2(\AES_ENC/us32/n1059 ), .A3(\AES_ENC/us32/n611 ), .ZN(\AES_ENC/us32/n1115 ) );
INV_X4 \AES_ENC/us32/U364  ( .A(\AES_ENC/us32/n1094 ), .ZN(\AES_ENC/us32/n613 ) );
NOR2_X2 \AES_ENC/us32/U363  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n931 ), .ZN(\AES_ENC/us32/n1100 ) );
INV_X4 \AES_ENC/us32/U354  ( .A(\AES_ENC/us32/n1093 ), .ZN(\AES_ENC/us32/n617 ) );
NOR2_X2 \AES_ENC/us32/U353  ( .A1(\AES_ENC/us32/n569 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n929 ) );
NOR2_X2 \AES_ENC/us32/U352  ( .A1(\AES_ENC/us32/n620 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n926 ) );
NOR2_X2 \AES_ENC/us32/U351  ( .A1(\AES_ENC/us32/n572 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n1095 ) );
NOR2_X2 \AES_ENC/us32/U350  ( .A1(\AES_ENC/us32/n609 ), .A2(\AES_ENC/us32/n627 ), .ZN(\AES_ENC/us32/n1010 ) );
NOR2_X2 \AES_ENC/us32/U349  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n1103 ) );
NOR2_X2 \AES_ENC/us32/U348  ( .A1(\AES_ENC/us32/n622 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n1059 ) );
NOR2_X2 \AES_ENC/us32/U347  ( .A1(\AES_ENC/sa32 [1]), .A2(\AES_ENC/us32/n1120 ), .ZN(\AES_ENC/us32/n1022 ) );
NOR2_X2 \AES_ENC/us32/U346  ( .A1(\AES_ENC/us32/n619 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n911 ) );
NOR2_X2 \AES_ENC/us32/U345  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/us32/n1025 ), .ZN(\AES_ENC/us32/n826 ) );
NOR2_X2 \AES_ENC/us32/U338  ( .A1(\AES_ENC/us32/n626 ), .A2(\AES_ENC/us32/n607 ), .ZN(\AES_ENC/us32/n1072 ) );
NOR2_X2 \AES_ENC/us32/U335  ( .A1(\AES_ENC/us32/n627 ), .A2(\AES_ENC/us32/n616 ), .ZN(\AES_ENC/us32/n956 ) );
NOR2_X2 \AES_ENC/us32/U329  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/us32/n624 ), .ZN(\AES_ENC/us32/n1121 ) );
NOR2_X2 \AES_ENC/us32/U328  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/us32/n624 ), .ZN(\AES_ENC/us32/n1058 ) );
NOR2_X2 \AES_ENC/us32/U327  ( .A1(\AES_ENC/us32/n625 ), .A2(\AES_ENC/us32/n611 ), .ZN(\AES_ENC/us32/n1073 ) );
NOR2_X2 \AES_ENC/us32/U325  ( .A1(\AES_ENC/sa32 [1]), .A2(\AES_ENC/us32/n1025 ), .ZN(\AES_ENC/us32/n1054 ) );
NOR2_X2 \AES_ENC/us32/U324  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/us32/n931 ), .ZN(\AES_ENC/us32/n1029 ) );
NOR2_X2 \AES_ENC/us32/U319  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n1056 ) );
NOR2_X2 \AES_ENC/us32/U318  ( .A1(\AES_ENC/us32/n614 ), .A2(\AES_ENC/us32/n626 ), .ZN(\AES_ENC/us32/n1050 ) );
NOR2_X2 \AES_ENC/us32/U317  ( .A1(\AES_ENC/us32/n1121 ), .A2(\AES_ENC/us32/n1025 ), .ZN(\AES_ENC/us32/n1120 ) );
NOR2_X2 \AES_ENC/us32/U316  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/us32/n572 ), .ZN(\AES_ENC/us32/n1074 ) );
NOR2_X2 \AES_ENC/us32/U315  ( .A1(\AES_ENC/us32/n1058 ), .A2(\AES_ENC/us32/n1054 ), .ZN(\AES_ENC/us32/n878 ) );
NOR2_X2 \AES_ENC/us32/U314  ( .A1(\AES_ENC/us32/n878 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n879 ) );
NOR2_X2 \AES_ENC/us32/U312  ( .A1(\AES_ENC/us32/n880 ), .A2(\AES_ENC/us32/n879 ), .ZN(\AES_ENC/us32/n887 ) );
NOR2_X2 \AES_ENC/us32/U311  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n588 ), .ZN(\AES_ENC/us32/n957 ) );
NOR2_X2 \AES_ENC/us32/U310  ( .A1(\AES_ENC/us32/n958 ), .A2(\AES_ENC/us32/n957 ), .ZN(\AES_ENC/us32/n965 ) );
NOR3_X2 \AES_ENC/us32/U309  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n1091 ), .A3(\AES_ENC/us32/n1022 ), .ZN(\AES_ENC/us32/n720 ) );
NOR3_X2 \AES_ENC/us32/U303  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n1054 ), .A3(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n719 ) );
NOR2_X2 \AES_ENC/us32/U302  ( .A1(\AES_ENC/us32/n720 ), .A2(\AES_ENC/us32/n719 ), .ZN(\AES_ENC/us32/n726 ) );
NOR2_X2 \AES_ENC/us32/U300  ( .A1(\AES_ENC/us32/n614 ), .A2(\AES_ENC/us32/n591 ), .ZN(\AES_ENC/us32/n865 ) );
NOR2_X2 \AES_ENC/us32/U299  ( .A1(\AES_ENC/us32/n1059 ), .A2(\AES_ENC/us32/n1058 ), .ZN(\AES_ENC/us32/n1060 ) );
NOR2_X2 \AES_ENC/us32/U298  ( .A1(\AES_ENC/us32/n1095 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n668 ) );
NOR2_X2 \AES_ENC/us32/U297  ( .A1(\AES_ENC/us32/n911 ), .A2(\AES_ENC/us32/n910 ), .ZN(\AES_ENC/us32/n912 ) );
NOR2_X2 \AES_ENC/us32/U296  ( .A1(\AES_ENC/us32/n912 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n916 ) );
NOR2_X2 \AES_ENC/us32/U295  ( .A1(\AES_ENC/us32/n826 ), .A2(\AES_ENC/us32/n573 ), .ZN(\AES_ENC/us32/n750 ) );
NOR2_X2 \AES_ENC/us32/U294  ( .A1(\AES_ENC/us32/n750 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n751 ) );
NOR2_X2 \AES_ENC/us32/U293  ( .A1(\AES_ENC/us32/n907 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n908 ) );
NOR2_X2 \AES_ENC/us32/U292  ( .A1(\AES_ENC/us32/n990 ), .A2(\AES_ENC/us32/n926 ), .ZN(\AES_ENC/us32/n780 ) );
NOR2_X2 \AES_ENC/us32/U291  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n584 ), .ZN(\AES_ENC/us32/n838 ) );
NOR2_X2 \AES_ENC/us32/U290  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n602 ), .ZN(\AES_ENC/us32/n837 ) );
NOR2_X2 \AES_ENC/us32/U284  ( .A1(\AES_ENC/us32/n838 ), .A2(\AES_ENC/us32/n837 ), .ZN(\AES_ENC/us32/n845 ) );
NOR2_X2 \AES_ENC/us32/U283  ( .A1(\AES_ENC/us32/n1022 ), .A2(\AES_ENC/us32/n1058 ), .ZN(\AES_ENC/us32/n740 ) );
NOR2_X2 \AES_ENC/us32/U282  ( .A1(\AES_ENC/us32/n740 ), .A2(\AES_ENC/us32/n616 ), .ZN(\AES_ENC/us32/n742 ) );
NOR2_X2 \AES_ENC/us32/U281  ( .A1(\AES_ENC/us32/n1098 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n1099 ) );
NOR2_X2 \AES_ENC/us32/U280  ( .A1(\AES_ENC/us32/n1120 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n993 ) );
NOR2_X2 \AES_ENC/us32/U279  ( .A1(\AES_ENC/us32/n993 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n994 ) );
NOR2_X2 \AES_ENC/us32/U273  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n620 ), .ZN(\AES_ENC/us32/n1026 ) );
NOR2_X2 \AES_ENC/us32/U272  ( .A1(\AES_ENC/us32/n573 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n1027 ) );
NOR2_X2 \AES_ENC/us32/U271  ( .A1(\AES_ENC/us32/n1027 ), .A2(\AES_ENC/us32/n1026 ), .ZN(\AES_ENC/us32/n1028 ) );
NOR2_X2 \AES_ENC/us32/U270  ( .A1(\AES_ENC/us32/n1029 ), .A2(\AES_ENC/us32/n1028 ), .ZN(\AES_ENC/us32/n1034 ) );
NOR4_X2 \AES_ENC/us32/U269  ( .A1(\AES_ENC/us32/n757 ), .A2(\AES_ENC/us32/n756 ), .A3(\AES_ENC/us32/n755 ), .A4(\AES_ENC/us32/n754 ), .ZN(\AES_ENC/us32/n758 ) );
NOR2_X2 \AES_ENC/us32/U268  ( .A1(\AES_ENC/us32/n752 ), .A2(\AES_ENC/us32/n751 ), .ZN(\AES_ENC/us32/n759 ) );
NOR2_X2 \AES_ENC/us32/U267  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n1071 ), .ZN(\AES_ENC/us32/n669 ) );
NOR2_X2 \AES_ENC/us32/U263  ( .A1(\AES_ENC/us32/n1056 ), .A2(\AES_ENC/us32/n990 ), .ZN(\AES_ENC/us32/n991 ) );
NOR2_X2 \AES_ENC/us32/U262  ( .A1(\AES_ENC/us32/n991 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n995 ) );
NOR2_X2 \AES_ENC/us32/U258  ( .A1(\AES_ENC/us32/n607 ), .A2(\AES_ENC/us32/n590 ), .ZN(\AES_ENC/us32/n1008 ) );
NOR2_X2 \AES_ENC/us32/U255  ( .A1(\AES_ENC/us32/n839 ), .A2(\AES_ENC/us32/n582 ), .ZN(\AES_ENC/us32/n693 ) );
NOR2_X2 \AES_ENC/us32/U254  ( .A1(\AES_ENC/us32/n606 ), .A2(\AES_ENC/us32/n906 ), .ZN(\AES_ENC/us32/n741 ) );
NOR2_X2 \AES_ENC/us32/U253  ( .A1(\AES_ENC/us32/n1054 ), .A2(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n763 ) );
NOR2_X2 \AES_ENC/us32/U252  ( .A1(\AES_ENC/us32/n763 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n769 ) );
NOR2_X2 \AES_ENC/us32/U251  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n577 ), .ZN(\AES_ENC/us32/n1007 ) );
NOR2_X2 \AES_ENC/us32/U250  ( .A1(\AES_ENC/us32/n609 ), .A2(\AES_ENC/us32/n580 ), .ZN(\AES_ENC/us32/n1123 ) );
NOR2_X2 \AES_ENC/us32/U243  ( .A1(\AES_ENC/us32/n609 ), .A2(\AES_ENC/us32/n590 ), .ZN(\AES_ENC/us32/n710 ) );
INV_X4 \AES_ENC/us32/U242  ( .A(\AES_ENC/us32/n1029 ), .ZN(\AES_ENC/us32/n582 ) );
NOR2_X2 \AES_ENC/us32/U241  ( .A1(\AES_ENC/us32/n616 ), .A2(\AES_ENC/us32/n597 ), .ZN(\AES_ENC/us32/n883 ) );
NOR2_X2 \AES_ENC/us32/U240  ( .A1(\AES_ENC/us32/n593 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n1125 ) );
NOR2_X2 \AES_ENC/us32/U239  ( .A1(\AES_ENC/us32/n990 ), .A2(\AES_ENC/us32/n929 ), .ZN(\AES_ENC/us32/n892 ) );
NOR2_X2 \AES_ENC/us32/U238  ( .A1(\AES_ENC/us32/n892 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n893 ) );
NOR2_X2 \AES_ENC/us32/U237  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n602 ), .ZN(\AES_ENC/us32/n950 ) );
NOR2_X2 \AES_ENC/us32/U236  ( .A1(\AES_ENC/us32/n1079 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n1082 ) );
NOR2_X2 \AES_ENC/us32/U235  ( .A1(\AES_ENC/us32/n910 ), .A2(\AES_ENC/us32/n1056 ), .ZN(\AES_ENC/us32/n941 ) );
NOR2_X2 \AES_ENC/us32/U234  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n1077 ), .ZN(\AES_ENC/us32/n841 ) );
NOR2_X2 \AES_ENC/us32/U229  ( .A1(\AES_ENC/us32/n623 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n630 ) );
NOR2_X2 \AES_ENC/us32/U228  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n602 ), .ZN(\AES_ENC/us32/n806 ) );
NOR2_X2 \AES_ENC/us32/U227  ( .A1(\AES_ENC/us32/n623 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n948 ) );
NOR2_X2 \AES_ENC/us32/U226  ( .A1(\AES_ENC/us32/n606 ), .A2(\AES_ENC/us32/n589 ), .ZN(\AES_ENC/us32/n997 ) );
NOR2_X2 \AES_ENC/us32/U225  ( .A1(\AES_ENC/us32/n1121 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n1122 ) );
NOR2_X2 \AES_ENC/us32/U223  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n1023 ), .ZN(\AES_ENC/us32/n756 ) );
NOR2_X2 \AES_ENC/us32/U222  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n602 ), .ZN(\AES_ENC/us32/n870 ) );
NOR2_X2 \AES_ENC/us32/U221  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n569 ), .ZN(\AES_ENC/us32/n947 ) );
NOR2_X2 \AES_ENC/us32/U217  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n1077 ), .ZN(\AES_ENC/us32/n1084 ) );
NOR2_X2 \AES_ENC/us32/U213  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n855 ), .ZN(\AES_ENC/us32/n709 ) );
NOR2_X2 \AES_ENC/us32/U212  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n589 ), .ZN(\AES_ENC/us32/n868 ) );
NOR2_X2 \AES_ENC/us32/U211  ( .A1(\AES_ENC/us32/n1120 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n1124 ) );
NOR2_X2 \AES_ENC/us32/U210  ( .A1(\AES_ENC/us32/n1120 ), .A2(\AES_ENC/us32/n839 ), .ZN(\AES_ENC/us32/n842 ) );
NOR2_X2 \AES_ENC/us32/U209  ( .A1(\AES_ENC/us32/n1120 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n696 ) );
NOR2_X2 \AES_ENC/us32/U208  ( .A1(\AES_ENC/us32/n1074 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n1076 ) );
NOR2_X2 \AES_ENC/us32/U207  ( .A1(\AES_ENC/us32/n1074 ), .A2(\AES_ENC/us32/n620 ), .ZN(\AES_ENC/us32/n781 ) );
NOR3_X2 \AES_ENC/us32/U201  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n1056 ), .A3(\AES_ENC/us32/n990 ), .ZN(\AES_ENC/us32/n979 ) );
NOR3_X2 \AES_ENC/us32/U200  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n1058 ), .A3(\AES_ENC/us32/n1059 ), .ZN(\AES_ENC/us32/n854 ) );
NOR2_X2 \AES_ENC/us32/U199  ( .A1(\AES_ENC/us32/n996 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n869 ) );
NOR2_X2 \AES_ENC/us32/U198  ( .A1(\AES_ENC/us32/n1056 ), .A2(\AES_ENC/us32/n1074 ), .ZN(\AES_ENC/us32/n1057 ) );
NOR3_X2 \AES_ENC/us32/U197  ( .A1(\AES_ENC/us32/n607 ), .A2(\AES_ENC/us32/n1120 ), .A3(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n978 ) );
NOR2_X2 \AES_ENC/us32/U196  ( .A1(\AES_ENC/us32/n996 ), .A2(\AES_ENC/us32/n911 ), .ZN(\AES_ENC/us32/n1116 ) );
NOR2_X2 \AES_ENC/us32/U195  ( .A1(\AES_ENC/us32/n1074 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n754 ) );
NOR2_X2 \AES_ENC/us32/U194  ( .A1(\AES_ENC/us32/n926 ), .A2(\AES_ENC/us32/n1103 ), .ZN(\AES_ENC/us32/n977 ) );
NOR2_X2 \AES_ENC/us32/U187  ( .A1(\AES_ENC/us32/n839 ), .A2(\AES_ENC/us32/n824 ), .ZN(\AES_ENC/us32/n1092 ) );
NOR2_X2 \AES_ENC/us32/U186  ( .A1(\AES_ENC/us32/n573 ), .A2(\AES_ENC/us32/n1074 ), .ZN(\AES_ENC/us32/n684 ) );
NOR2_X2 \AES_ENC/us32/U185  ( .A1(\AES_ENC/us32/n826 ), .A2(\AES_ENC/us32/n1059 ), .ZN(\AES_ENC/us32/n907 ) );
NOR3_X2 \AES_ENC/us32/U184  ( .A1(\AES_ENC/us32/n625 ), .A2(\AES_ENC/us32/n1115 ), .A3(\AES_ENC/us32/n585 ), .ZN(\AES_ENC/us32/n831 ) );
NOR3_X2 \AES_ENC/us32/U183  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n1056 ), .A3(\AES_ENC/us32/n990 ), .ZN(\AES_ENC/us32/n896 ) );
NOR3_X2 \AES_ENC/us32/U182  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n573 ), .A3(\AES_ENC/us32/n1013 ), .ZN(\AES_ENC/us32/n670 ) );
NOR3_X2 \AES_ENC/us32/U181  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n1091 ), .A3(\AES_ENC/us32/n1022 ), .ZN(\AES_ENC/us32/n843 ) );
NOR2_X2 \AES_ENC/us32/U180  ( .A1(\AES_ENC/us32/n1029 ), .A2(\AES_ENC/us32/n1095 ), .ZN(\AES_ENC/us32/n735 ) );
NOR2_X2 \AES_ENC/us32/U174  ( .A1(\AES_ENC/us32/n1100 ), .A2(\AES_ENC/us32/n854 ), .ZN(\AES_ENC/us32/n860 ) );
NOR4_X2 \AES_ENC/us32/U173  ( .A1(\AES_ENC/us32/n1125 ), .A2(\AES_ENC/us32/n1124 ), .A3(\AES_ENC/us32/n1123 ), .A4(\AES_ENC/us32/n1122 ), .ZN(\AES_ENC/us32/n1126 ) );
NOR4_X2 \AES_ENC/us32/U172  ( .A1(\AES_ENC/us32/n1084 ), .A2(\AES_ENC/us32/n1083 ), .A3(\AES_ENC/us32/n1082 ), .A4(\AES_ENC/us32/n1081 ), .ZN(\AES_ENC/us32/n1085 ) );
NOR2_X2 \AES_ENC/us32/U171  ( .A1(\AES_ENC/us32/n1076 ), .A2(\AES_ENC/us32/n1075 ), .ZN(\AES_ENC/us32/n1086 ) );
NAND3_X2 \AES_ENC/us32/U170  ( .A1(\AES_ENC/us32/n569 ), .A2(\AES_ENC/us32/n582 ), .A3(\AES_ENC/us32/n681 ), .ZN(\AES_ENC/us32/n691 ) );
NOR2_X2 \AES_ENC/us32/U169  ( .A1(\AES_ENC/us32/n683 ), .A2(\AES_ENC/us32/n682 ), .ZN(\AES_ENC/us32/n690 ) );
NOR3_X2 \AES_ENC/us32/U168  ( .A1(\AES_ENC/us32/n695 ), .A2(\AES_ENC/us32/n694 ), .A3(\AES_ENC/us32/n693 ), .ZN(\AES_ENC/us32/n700 ) );
NOR4_X2 \AES_ENC/us32/U162  ( .A1(\AES_ENC/us32/n983 ), .A2(\AES_ENC/us32/n698 ), .A3(\AES_ENC/us32/n697 ), .A4(\AES_ENC/us32/n696 ), .ZN(\AES_ENC/us32/n699 ) );
NOR2_X2 \AES_ENC/us32/U161  ( .A1(\AES_ENC/us32/n946 ), .A2(\AES_ENC/us32/n945 ), .ZN(\AES_ENC/us32/n952 ) );
NOR4_X2 \AES_ENC/us32/U160  ( .A1(\AES_ENC/us32/n950 ), .A2(\AES_ENC/us32/n949 ), .A3(\AES_ENC/us32/n948 ), .A4(\AES_ENC/us32/n947 ), .ZN(\AES_ENC/us32/n951 ) );
NOR4_X2 \AES_ENC/us32/U159  ( .A1(\AES_ENC/us32/n896 ), .A2(\AES_ENC/us32/n895 ), .A3(\AES_ENC/us32/n894 ), .A4(\AES_ENC/us32/n893 ), .ZN(\AES_ENC/us32/n897 ) );
NOR2_X2 \AES_ENC/us32/U158  ( .A1(\AES_ENC/us32/n866 ), .A2(\AES_ENC/us32/n865 ), .ZN(\AES_ENC/us32/n872 ) );
NOR4_X2 \AES_ENC/us32/U157  ( .A1(\AES_ENC/us32/n870 ), .A2(\AES_ENC/us32/n869 ), .A3(\AES_ENC/us32/n868 ), .A4(\AES_ENC/us32/n867 ), .ZN(\AES_ENC/us32/n871 ) );
NOR4_X2 \AES_ENC/us32/U156  ( .A1(\AES_ENC/us32/n983 ), .A2(\AES_ENC/us32/n982 ), .A3(\AES_ENC/us32/n981 ), .A4(\AES_ENC/us32/n980 ), .ZN(\AES_ENC/us32/n984 ) );
NOR2_X2 \AES_ENC/us32/U155  ( .A1(\AES_ENC/us32/n979 ), .A2(\AES_ENC/us32/n978 ), .ZN(\AES_ENC/us32/n985 ) );
NOR3_X2 \AES_ENC/us32/U154  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n1054 ), .A3(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n961 ) );
NOR3_X2 \AES_ENC/us32/U153  ( .A1(\AES_ENC/us32/n620 ), .A2(\AES_ENC/us32/n1074 ), .A3(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n671 ) );
NOR2_X2 \AES_ENC/us32/U152  ( .A1(\AES_ENC/us32/n1057 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n1062 ) );
NOR2_X2 \AES_ENC/us32/U143  ( .A1(\AES_ENC/us32/n1055 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n1063 ) );
NOR2_X2 \AES_ENC/us32/U142  ( .A1(\AES_ENC/us32/n1060 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n1061 ) );
NOR4_X2 \AES_ENC/us32/U141  ( .A1(\AES_ENC/us32/n1064 ), .A2(\AES_ENC/us32/n1063 ), .A3(\AES_ENC/us32/n1062 ), .A4(\AES_ENC/us32/n1061 ), .ZN(\AES_ENC/us32/n1065 ) );
NOR3_X2 \AES_ENC/us32/U140  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n1120 ), .A3(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n918 ) );
NOR3_X2 \AES_ENC/us32/U132  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n573 ), .A3(\AES_ENC/us32/n1013 ), .ZN(\AES_ENC/us32/n917 ) );
NOR2_X2 \AES_ENC/us32/U131  ( .A1(\AES_ENC/us32/n914 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n915 ) );
NOR4_X2 \AES_ENC/us32/U130  ( .A1(\AES_ENC/us32/n918 ), .A2(\AES_ENC/us32/n917 ), .A3(\AES_ENC/us32/n916 ), .A4(\AES_ENC/us32/n915 ), .ZN(\AES_ENC/us32/n919 ) );
NOR2_X2 \AES_ENC/us32/U129  ( .A1(\AES_ENC/us32/n616 ), .A2(\AES_ENC/us32/n580 ), .ZN(\AES_ENC/us32/n771 ) );
NOR2_X2 \AES_ENC/us32/U128  ( .A1(\AES_ENC/us32/n1103 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n772 ) );
NOR2_X2 \AES_ENC/us32/U127  ( .A1(\AES_ENC/us32/n610 ), .A2(\AES_ENC/us32/n599 ), .ZN(\AES_ENC/us32/n773 ) );
NOR4_X2 \AES_ENC/us32/U126  ( .A1(\AES_ENC/us32/n773 ), .A2(\AES_ENC/us32/n772 ), .A3(\AES_ENC/us32/n771 ), .A4(\AES_ENC/us32/n770 ), .ZN(\AES_ENC/us32/n774 ) );
NOR2_X2 \AES_ENC/us32/U121  ( .A1(\AES_ENC/us32/n735 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n687 ) );
NOR2_X2 \AES_ENC/us32/U120  ( .A1(\AES_ENC/us32/n684 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n688 ) );
NOR2_X2 \AES_ENC/us32/U119  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n600 ), .ZN(\AES_ENC/us32/n686 ) );
NOR4_X2 \AES_ENC/us32/U118  ( .A1(\AES_ENC/us32/n688 ), .A2(\AES_ENC/us32/n687 ), .A3(\AES_ENC/us32/n686 ), .A4(\AES_ENC/us32/n685 ), .ZN(\AES_ENC/us32/n689 ) );
NOR2_X2 \AES_ENC/us32/U117  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n595 ), .ZN(\AES_ENC/us32/n858 ) );
NOR2_X2 \AES_ENC/us32/U116  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n855 ), .ZN(\AES_ENC/us32/n857 ) );
NOR2_X2 \AES_ENC/us32/U115  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n587 ), .ZN(\AES_ENC/us32/n856 ) );
NOR4_X2 \AES_ENC/us32/U106  ( .A1(\AES_ENC/us32/n858 ), .A2(\AES_ENC/us32/n857 ), .A3(\AES_ENC/us32/n856 ), .A4(\AES_ENC/us32/n958 ), .ZN(\AES_ENC/us32/n859 ) );
NOR2_X2 \AES_ENC/us32/U105  ( .A1(\AES_ENC/us32/n780 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n784 ) );
NOR2_X2 \AES_ENC/us32/U104  ( .A1(\AES_ENC/us32/n1117 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n782 ) );
NOR2_X2 \AES_ENC/us32/U103  ( .A1(\AES_ENC/us32/n781 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n783 ) );
NOR4_X2 \AES_ENC/us32/U102  ( .A1(\AES_ENC/us32/n880 ), .A2(\AES_ENC/us32/n784 ), .A3(\AES_ENC/us32/n783 ), .A4(\AES_ENC/us32/n782 ), .ZN(\AES_ENC/us32/n785 ) );
NOR2_X2 \AES_ENC/us32/U101  ( .A1(\AES_ENC/us32/n583 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n814 ) );
NOR2_X2 \AES_ENC/us32/U100  ( .A1(\AES_ENC/us32/n907 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n813 ) );
NOR3_X2 \AES_ENC/us32/U95  ( .A1(\AES_ENC/us32/n606 ), .A2(\AES_ENC/us32/n1058 ), .A3(\AES_ENC/us32/n1059 ), .ZN(\AES_ENC/us32/n815 ) );
NOR4_X2 \AES_ENC/us32/U94  ( .A1(\AES_ENC/us32/n815 ), .A2(\AES_ENC/us32/n814 ), .A3(\AES_ENC/us32/n813 ), .A4(\AES_ENC/us32/n812 ), .ZN(\AES_ENC/us32/n816 ) );
NOR2_X2 \AES_ENC/us32/U93  ( .A1(\AES_ENC/us32/n617 ), .A2(\AES_ENC/us32/n569 ), .ZN(\AES_ENC/us32/n721 ) );
NOR2_X2 \AES_ENC/us32/U92  ( .A1(\AES_ENC/us32/n1031 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n723 ) );
NOR2_X2 \AES_ENC/us32/U91  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n1096 ), .ZN(\AES_ENC/us32/n722 ) );
NOR4_X2 \AES_ENC/us32/U90  ( .A1(\AES_ENC/us32/n724 ), .A2(\AES_ENC/us32/n723 ), .A3(\AES_ENC/us32/n722 ), .A4(\AES_ENC/us32/n721 ), .ZN(\AES_ENC/us32/n725 ) );
NOR2_X2 \AES_ENC/us32/U89  ( .A1(\AES_ENC/us32/n911 ), .A2(\AES_ENC/us32/n990 ), .ZN(\AES_ENC/us32/n1009 ) );
NOR2_X2 \AES_ENC/us32/U88  ( .A1(\AES_ENC/us32/n1013 ), .A2(\AES_ENC/us32/n573 ), .ZN(\AES_ENC/us32/n1014 ) );
NOR2_X2 \AES_ENC/us32/U87  ( .A1(\AES_ENC/us32/n1014 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n1015 ) );
NOR4_X2 \AES_ENC/us32/U86  ( .A1(\AES_ENC/us32/n1016 ), .A2(\AES_ENC/us32/n1015 ), .A3(\AES_ENC/us32/n1119 ), .A4(\AES_ENC/us32/n1046 ), .ZN(\AES_ENC/us32/n1017 ) );
NOR2_X2 \AES_ENC/us32/U81  ( .A1(\AES_ENC/us32/n996 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n998 ) );
NOR2_X2 \AES_ENC/us32/U80  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n577 ), .ZN(\AES_ENC/us32/n1000 ) );
NOR2_X2 \AES_ENC/us32/U79  ( .A1(\AES_ENC/us32/n616 ), .A2(\AES_ENC/us32/n1096 ), .ZN(\AES_ENC/us32/n999 ) );
NOR4_X2 \AES_ENC/us32/U78  ( .A1(\AES_ENC/us32/n1000 ), .A2(\AES_ENC/us32/n999 ), .A3(\AES_ENC/us32/n998 ), .A4(\AES_ENC/us32/n997 ), .ZN(\AES_ENC/us32/n1001 ) );
NOR2_X2 \AES_ENC/us32/U74  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n1096 ), .ZN(\AES_ENC/us32/n697 ) );
NOR2_X2 \AES_ENC/us32/U73  ( .A1(\AES_ENC/us32/n620 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n958 ) );
NOR2_X2 \AES_ENC/us32/U72  ( .A1(\AES_ENC/us32/n911 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n983 ) );
NOR2_X2 \AES_ENC/us32/U71  ( .A1(\AES_ENC/us32/n1054 ), .A2(\AES_ENC/us32/n1103 ), .ZN(\AES_ENC/us32/n1031 ) );
INV_X4 \AES_ENC/us32/U65  ( .A(\AES_ENC/us32/n1050 ), .ZN(\AES_ENC/us32/n612 ) );
INV_X4 \AES_ENC/us32/U64  ( .A(\AES_ENC/us32/n1072 ), .ZN(\AES_ENC/us32/n605 ) );
INV_X4 \AES_ENC/us32/U63  ( .A(\AES_ENC/us32/n1073 ), .ZN(\AES_ENC/us32/n604 ) );
NOR2_X2 \AES_ENC/us32/U62  ( .A1(\AES_ENC/us32/n582 ), .A2(\AES_ENC/us32/n613 ), .ZN(\AES_ENC/us32/n880 ) );
NOR3_X2 \AES_ENC/us32/U61  ( .A1(\AES_ENC/us32/n826 ), .A2(\AES_ENC/us32/n1121 ), .A3(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n946 ) );
INV_X4 \AES_ENC/us32/U59  ( .A(\AES_ENC/us32/n1010 ), .ZN(\AES_ENC/us32/n608 ) );
NOR3_X2 \AES_ENC/us32/U58  ( .A1(\AES_ENC/us32/n573 ), .A2(\AES_ENC/us32/n1029 ), .A3(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n1119 ) );
INV_X4 \AES_ENC/us32/U57  ( .A(\AES_ENC/us32/n956 ), .ZN(\AES_ENC/us32/n615 ) );
NOR2_X2 \AES_ENC/us32/U50  ( .A1(\AES_ENC/us32/n623 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n1013 ) );
NOR2_X2 \AES_ENC/us32/U49  ( .A1(\AES_ENC/us32/n620 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n910 ) );
NOR2_X2 \AES_ENC/us32/U48  ( .A1(\AES_ENC/us32/n569 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n1091 ) );
NOR2_X2 \AES_ENC/us32/U47  ( .A1(\AES_ENC/us32/n622 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n990 ) );
NOR2_X2 \AES_ENC/us32/U46  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/us32/n1121 ), .ZN(\AES_ENC/us32/n996 ) );
NOR2_X2 \AES_ENC/us32/U45  ( .A1(\AES_ENC/us32/n610 ), .A2(\AES_ENC/us32/n600 ), .ZN(\AES_ENC/us32/n628 ) );
NOR2_X2 \AES_ENC/us32/U44  ( .A1(\AES_ENC/us32/n576 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n866 ) );
NOR2_X2 \AES_ENC/us32/U43  ( .A1(\AES_ENC/us32/n603 ), .A2(\AES_ENC/us32/n610 ), .ZN(\AES_ENC/us32/n1006 ) );
NOR2_X2 \AES_ENC/us32/U42  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n1117 ), .ZN(\AES_ENC/us32/n1118 ) );
NOR2_X2 \AES_ENC/us32/U41  ( .A1(\AES_ENC/us32/n1119 ), .A2(\AES_ENC/us32/n1118 ), .ZN(\AES_ENC/us32/n1127 ) );
NOR2_X2 \AES_ENC/us32/U36  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n906 ), .ZN(\AES_ENC/us32/n909 ) );
NOR2_X2 \AES_ENC/us32/U35  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n594 ), .ZN(\AES_ENC/us32/n629 ) );
NOR2_X2 \AES_ENC/us32/U34  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n597 ), .ZN(\AES_ENC/us32/n658 ) );
NOR2_X2 \AES_ENC/us32/U33  ( .A1(\AES_ENC/us32/n1116 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n695 ) );
NOR2_X2 \AES_ENC/us32/U32  ( .A1(\AES_ENC/us32/n1078 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n1083 ) );
NOR2_X2 \AES_ENC/us32/U31  ( .A1(\AES_ENC/us32/n941 ), .A2(\AES_ENC/us32/n608 ), .ZN(\AES_ENC/us32/n724 ) );
NOR2_X2 \AES_ENC/us32/U30  ( .A1(\AES_ENC/us32/n598 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n1107 ) );
NOR2_X2 \AES_ENC/us32/U29  ( .A1(\AES_ENC/us32/n576 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n840 ) );
NOR2_X2 \AES_ENC/us32/U24  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n593 ), .ZN(\AES_ENC/us32/n633 ) );
NOR2_X2 \AES_ENC/us32/U23  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n1080 ), .ZN(\AES_ENC/us32/n1081 ) );
NOR2_X2 \AES_ENC/us32/U21  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n1045 ), .ZN(\AES_ENC/us32/n812 ) );
NOR2_X2 \AES_ENC/us32/U20  ( .A1(\AES_ENC/us32/n1009 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n960 ) );
NOR2_X2 \AES_ENC/us32/U19  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n601 ), .ZN(\AES_ENC/us32/n982 ) );
NOR2_X2 \AES_ENC/us32/U18  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n594 ), .ZN(\AES_ENC/us32/n757 ) );
NOR2_X2 \AES_ENC/us32/U17  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n590 ), .ZN(\AES_ENC/us32/n698 ) );
NOR2_X2 \AES_ENC/us32/U16  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n619 ), .ZN(\AES_ENC/us32/n708 ) );
NOR2_X2 \AES_ENC/us32/U15  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n582 ), .ZN(\AES_ENC/us32/n770 ) );
NOR2_X2 \AES_ENC/us32/U10  ( .A1(\AES_ENC/us32/n619 ), .A2(\AES_ENC/us32/n604 ), .ZN(\AES_ENC/us32/n803 ) );
NOR2_X2 \AES_ENC/us32/U9  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n881 ), .ZN(\AES_ENC/us32/n711 ) );
NOR2_X2 \AES_ENC/us32/U8  ( .A1(\AES_ENC/us32/n615 ), .A2(\AES_ENC/us32/n582 ), .ZN(\AES_ENC/us32/n867 ) );
NOR2_X2 \AES_ENC/us32/U7  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n599 ), .ZN(\AES_ENC/us32/n804 ) );
NOR2_X2 \AES_ENC/us32/U6  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n620 ), .ZN(\AES_ENC/us32/n1046 ) );
OR2_X4 \AES_ENC/us32/U5  ( .A1(\AES_ENC/us32/n624 ), .A2(\AES_ENC/sa32 [1]),.ZN(\AES_ENC/us32/n570 ) );
OR2_X4 \AES_ENC/us32/U4  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/sa32 [4]),.ZN(\AES_ENC/us32/n569 ) );
NAND2_X2 \AES_ENC/us32/U514  ( .A1(\AES_ENC/us32/n1121 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n1030 ) );
AND2_X2 \AES_ENC/us32/U513  ( .A1(\AES_ENC/us32/n597 ), .A2(\AES_ENC/us32/n1030 ), .ZN(\AES_ENC/us32/n1049 ) );
NAND2_X2 \AES_ENC/us32/U511  ( .A1(\AES_ENC/us32/n1049 ), .A2(\AES_ENC/us32/n794 ), .ZN(\AES_ENC/us32/n637 ) );
AND2_X2 \AES_ENC/us32/U493  ( .A1(\AES_ENC/us32/n779 ), .A2(\AES_ENC/us32/n996 ), .ZN(\AES_ENC/us32/n632 ) );
NAND4_X2 \AES_ENC/us32/U485  ( .A1(\AES_ENC/us32/n637 ), .A2(\AES_ENC/us32/n636 ), .A3(\AES_ENC/us32/n635 ), .A4(\AES_ENC/us32/n634 ), .ZN(\AES_ENC/us32/n638 ) );
NAND2_X2 \AES_ENC/us32/U484  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n638 ), .ZN(\AES_ENC/us32/n679 ) );
NAND2_X2 \AES_ENC/us32/U481  ( .A1(\AES_ENC/us32/n1094 ), .A2(\AES_ENC/us32/n591 ), .ZN(\AES_ENC/us32/n648 ) );
NAND2_X2 \AES_ENC/us32/U476  ( .A1(\AES_ENC/us32/n601 ), .A2(\AES_ENC/us32/n590 ), .ZN(\AES_ENC/us32/n762 ) );
NAND2_X2 \AES_ENC/us32/U475  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n762 ), .ZN(\AES_ENC/us32/n647 ) );
NAND4_X2 \AES_ENC/us32/U457  ( .A1(\AES_ENC/us32/n648 ), .A2(\AES_ENC/us32/n647 ), .A3(\AES_ENC/us32/n646 ), .A4(\AES_ENC/us32/n645 ), .ZN(\AES_ENC/us32/n649 ) );
NAND2_X2 \AES_ENC/us32/U456  ( .A1(\AES_ENC/sa32 [0]), .A2(\AES_ENC/us32/n649 ), .ZN(\AES_ENC/us32/n665 ) );
NAND2_X2 \AES_ENC/us32/U454  ( .A1(\AES_ENC/us32/n596 ), .A2(\AES_ENC/us32/n623 ), .ZN(\AES_ENC/us32/n855 ) );
NAND2_X2 \AES_ENC/us32/U453  ( .A1(\AES_ENC/us32/n587 ), .A2(\AES_ENC/us32/n855 ), .ZN(\AES_ENC/us32/n821 ) );
NAND2_X2 \AES_ENC/us32/U452  ( .A1(\AES_ENC/us32/n1093 ), .A2(\AES_ENC/us32/n821 ), .ZN(\AES_ENC/us32/n662 ) );
NAND2_X2 \AES_ENC/us32/U451  ( .A1(\AES_ENC/us32/n619 ), .A2(\AES_ENC/us32/n589 ), .ZN(\AES_ENC/us32/n650 ) );
NAND2_X2 \AES_ENC/us32/U450  ( .A1(\AES_ENC/us32/n956 ), .A2(\AES_ENC/us32/n650 ), .ZN(\AES_ENC/us32/n661 ) );
NAND2_X2 \AES_ENC/us32/U449  ( .A1(\AES_ENC/us32/n626 ), .A2(\AES_ENC/us32/n627 ), .ZN(\AES_ENC/us32/n839 ) );
OR2_X2 \AES_ENC/us32/U446  ( .A1(\AES_ENC/us32/n839 ), .A2(\AES_ENC/us32/n932 ), .ZN(\AES_ENC/us32/n656 ) );
NAND2_X2 \AES_ENC/us32/U445  ( .A1(\AES_ENC/us32/n621 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n1096 ) );
NAND2_X2 \AES_ENC/us32/U444  ( .A1(\AES_ENC/us32/n1030 ), .A2(\AES_ENC/us32/n1096 ), .ZN(\AES_ENC/us32/n651 ) );
NAND2_X2 \AES_ENC/us32/U443  ( .A1(\AES_ENC/us32/n1114 ), .A2(\AES_ENC/us32/n651 ), .ZN(\AES_ENC/us32/n655 ) );
OR3_X2 \AES_ENC/us32/U440  ( .A1(\AES_ENC/us32/n1079 ), .A2(\AES_ENC/sa32 [7]), .A3(\AES_ENC/us32/n626 ), .ZN(\AES_ENC/us32/n654 ));
NAND2_X2 \AES_ENC/us32/U439  ( .A1(\AES_ENC/us32/n593 ), .A2(\AES_ENC/us32/n601 ), .ZN(\AES_ENC/us32/n652 ) );
NAND4_X2 \AES_ENC/us32/U437  ( .A1(\AES_ENC/us32/n656 ), .A2(\AES_ENC/us32/n655 ), .A3(\AES_ENC/us32/n654 ), .A4(\AES_ENC/us32/n653 ), .ZN(\AES_ENC/us32/n657 ) );
NAND2_X2 \AES_ENC/us32/U436  ( .A1(\AES_ENC/sa32 [2]), .A2(\AES_ENC/us32/n657 ), .ZN(\AES_ENC/us32/n660 ) );
NAND4_X2 \AES_ENC/us32/U432  ( .A1(\AES_ENC/us32/n662 ), .A2(\AES_ENC/us32/n661 ), .A3(\AES_ENC/us32/n660 ), .A4(\AES_ENC/us32/n659 ), .ZN(\AES_ENC/us32/n663 ) );
NAND2_X2 \AES_ENC/us32/U431  ( .A1(\AES_ENC/us32/n663 ), .A2(\AES_ENC/us32/n574 ), .ZN(\AES_ENC/us32/n664 ) );
NAND2_X2 \AES_ENC/us32/U430  ( .A1(\AES_ENC/us32/n665 ), .A2(\AES_ENC/us32/n664 ), .ZN(\AES_ENC/us32/n666 ) );
NAND2_X2 \AES_ENC/us32/U429  ( .A1(\AES_ENC/sa32 [6]), .A2(\AES_ENC/us32/n666 ), .ZN(\AES_ENC/us32/n678 ) );
NAND2_X2 \AES_ENC/us32/U426  ( .A1(\AES_ENC/us32/n735 ), .A2(\AES_ENC/us32/n1093 ), .ZN(\AES_ENC/us32/n675 ) );
NAND2_X2 \AES_ENC/us32/U425  ( .A1(\AES_ENC/us32/n588 ), .A2(\AES_ENC/us32/n597 ), .ZN(\AES_ENC/us32/n1045 ) );
OR2_X2 \AES_ENC/us32/U424  ( .A1(\AES_ENC/us32/n1045 ), .A2(\AES_ENC/us32/n605 ), .ZN(\AES_ENC/us32/n674 ) );
NAND2_X2 \AES_ENC/us32/U423  ( .A1(\AES_ENC/sa32 [1]), .A2(\AES_ENC/us32/n620 ), .ZN(\AES_ENC/us32/n667 ) );
NAND2_X2 \AES_ENC/us32/U422  ( .A1(\AES_ENC/us32/n619 ), .A2(\AES_ENC/us32/n667 ), .ZN(\AES_ENC/us32/n1071 ) );
NAND4_X2 \AES_ENC/us32/U412  ( .A1(\AES_ENC/us32/n675 ), .A2(\AES_ENC/us32/n674 ), .A3(\AES_ENC/us32/n673 ), .A4(\AES_ENC/us32/n672 ), .ZN(\AES_ENC/us32/n676 ) );
NAND2_X2 \AES_ENC/us32/U411  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n676 ), .ZN(\AES_ENC/us32/n677 ) );
NAND2_X2 \AES_ENC/us32/U408  ( .A1(\AES_ENC/us32/n800 ), .A2(\AES_ENC/us32/n1022 ), .ZN(\AES_ENC/us32/n680 ) );
NAND2_X2 \AES_ENC/us32/U407  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n680 ), .ZN(\AES_ENC/us32/n681 ) );
AND2_X2 \AES_ENC/us32/U402  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n684 ), .ZN(\AES_ENC/us32/n682 ) );
NAND4_X2 \AES_ENC/us32/U395  ( .A1(\AES_ENC/us32/n691 ), .A2(\AES_ENC/us32/n581 ), .A3(\AES_ENC/us32/n690 ), .A4(\AES_ENC/us32/n689 ), .ZN(\AES_ENC/us32/n692 ) );
NAND2_X2 \AES_ENC/us32/U394  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n692 ), .ZN(\AES_ENC/us32/n733 ) );
NAND2_X2 \AES_ENC/us32/U392  ( .A1(\AES_ENC/us32/n977 ), .A2(\AES_ENC/us32/n1050 ), .ZN(\AES_ENC/us32/n702 ) );
NAND2_X2 \AES_ENC/us32/U391  ( .A1(\AES_ENC/us32/n1093 ), .A2(\AES_ENC/us32/n1045 ), .ZN(\AES_ENC/us32/n701 ) );
NAND4_X2 \AES_ENC/us32/U381  ( .A1(\AES_ENC/us32/n702 ), .A2(\AES_ENC/us32/n701 ), .A3(\AES_ENC/us32/n700 ), .A4(\AES_ENC/us32/n699 ), .ZN(\AES_ENC/us32/n703 ) );
NAND2_X2 \AES_ENC/us32/U380  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n703 ), .ZN(\AES_ENC/us32/n732 ) );
AND2_X2 \AES_ENC/us32/U379  ( .A1(\AES_ENC/sa32 [0]), .A2(\AES_ENC/sa32 [6]),.ZN(\AES_ENC/us32/n1113 ) );
NAND2_X2 \AES_ENC/us32/U378  ( .A1(\AES_ENC/us32/n601 ), .A2(\AES_ENC/us32/n1030 ), .ZN(\AES_ENC/us32/n881 ) );
NAND2_X2 \AES_ENC/us32/U377  ( .A1(\AES_ENC/us32/n1093 ), .A2(\AES_ENC/us32/n881 ), .ZN(\AES_ENC/us32/n715 ) );
NAND2_X2 \AES_ENC/us32/U376  ( .A1(\AES_ENC/us32/n1010 ), .A2(\AES_ENC/us32/n600 ), .ZN(\AES_ENC/us32/n714 ) );
NAND2_X2 \AES_ENC/us32/U375  ( .A1(\AES_ENC/us32/n855 ), .A2(\AES_ENC/us32/n588 ), .ZN(\AES_ENC/us32/n1117 ) );
XNOR2_X2 \AES_ENC/us32/U371  ( .A(\AES_ENC/us32/n611 ), .B(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n824 ) );
NAND4_X2 \AES_ENC/us32/U362  ( .A1(\AES_ENC/us32/n715 ), .A2(\AES_ENC/us32/n714 ), .A3(\AES_ENC/us32/n713 ), .A4(\AES_ENC/us32/n712 ), .ZN(\AES_ENC/us32/n716 ) );
NAND2_X2 \AES_ENC/us32/U361  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n716 ), .ZN(\AES_ENC/us32/n731 ) );
AND2_X2 \AES_ENC/us32/U360  ( .A1(\AES_ENC/sa32 [6]), .A2(\AES_ENC/us32/n574 ), .ZN(\AES_ENC/us32/n1131 ) );
NAND2_X2 \AES_ENC/us32/U359  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n717 ) );
NAND2_X2 \AES_ENC/us32/U358  ( .A1(\AES_ENC/us32/n1029 ), .A2(\AES_ENC/us32/n717 ), .ZN(\AES_ENC/us32/n728 ) );
NAND2_X2 \AES_ENC/us32/U357  ( .A1(\AES_ENC/sa32 [1]), .A2(\AES_ENC/us32/n624 ), .ZN(\AES_ENC/us32/n1097 ) );
NAND2_X2 \AES_ENC/us32/U356  ( .A1(\AES_ENC/us32/n603 ), .A2(\AES_ENC/us32/n1097 ), .ZN(\AES_ENC/us32/n718 ) );
NAND2_X2 \AES_ENC/us32/U355  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n718 ), .ZN(\AES_ENC/us32/n727 ) );
NAND4_X2 \AES_ENC/us32/U344  ( .A1(\AES_ENC/us32/n728 ), .A2(\AES_ENC/us32/n727 ), .A3(\AES_ENC/us32/n726 ), .A4(\AES_ENC/us32/n725 ), .ZN(\AES_ENC/us32/n729 ) );
NAND2_X2 \AES_ENC/us32/U343  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n729 ), .ZN(\AES_ENC/us32/n730 ) );
NAND4_X2 \AES_ENC/us32/U342  ( .A1(\AES_ENC/us32/n733 ), .A2(\AES_ENC/us32/n732 ), .A3(\AES_ENC/us32/n731 ), .A4(\AES_ENC/us32/n730 ), .ZN(\AES_ENC/sa32_sub[1] ) );
NAND2_X2 \AES_ENC/us32/U341  ( .A1(\AES_ENC/sa32 [7]), .A2(\AES_ENC/us32/n611 ), .ZN(\AES_ENC/us32/n734 ) );
NAND2_X2 \AES_ENC/us32/U340  ( .A1(\AES_ENC/us32/n734 ), .A2(\AES_ENC/us32/n607 ), .ZN(\AES_ENC/us32/n738 ) );
OR4_X2 \AES_ENC/us32/U339  ( .A1(\AES_ENC/us32/n738 ), .A2(\AES_ENC/us32/n626 ), .A3(\AES_ENC/us32/n826 ), .A4(\AES_ENC/us32/n1121 ), .ZN(\AES_ENC/us32/n746 ) );
NAND2_X2 \AES_ENC/us32/U337  ( .A1(\AES_ENC/us32/n1100 ), .A2(\AES_ENC/us32/n587 ), .ZN(\AES_ENC/us32/n992 ) );
OR2_X2 \AES_ENC/us32/U336  ( .A1(\AES_ENC/us32/n610 ), .A2(\AES_ENC/us32/n735 ), .ZN(\AES_ENC/us32/n737 ) );
NAND2_X2 \AES_ENC/us32/U334  ( .A1(\AES_ENC/us32/n619 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n753 ) );
NAND2_X2 \AES_ENC/us32/U333  ( .A1(\AES_ENC/us32/n582 ), .A2(\AES_ENC/us32/n753 ), .ZN(\AES_ENC/us32/n1080 ) );
NAND2_X2 \AES_ENC/us32/U332  ( .A1(\AES_ENC/us32/n1048 ), .A2(\AES_ENC/us32/n576 ), .ZN(\AES_ENC/us32/n736 ) );
NAND2_X2 \AES_ENC/us32/U331  ( .A1(\AES_ENC/us32/n737 ), .A2(\AES_ENC/us32/n736 ), .ZN(\AES_ENC/us32/n739 ) );
NAND2_X2 \AES_ENC/us32/U330  ( .A1(\AES_ENC/us32/n739 ), .A2(\AES_ENC/us32/n738 ), .ZN(\AES_ENC/us32/n745 ) );
NAND2_X2 \AES_ENC/us32/U326  ( .A1(\AES_ENC/us32/n1096 ), .A2(\AES_ENC/us32/n590 ), .ZN(\AES_ENC/us32/n906 ) );
NAND4_X2 \AES_ENC/us32/U323  ( .A1(\AES_ENC/us32/n746 ), .A2(\AES_ENC/us32/n992 ), .A3(\AES_ENC/us32/n745 ), .A4(\AES_ENC/us32/n744 ), .ZN(\AES_ENC/us32/n747 ) );
NAND2_X2 \AES_ENC/us32/U322  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n747 ), .ZN(\AES_ENC/us32/n793 ) );
NAND2_X2 \AES_ENC/us32/U321  ( .A1(\AES_ENC/us32/n584 ), .A2(\AES_ENC/us32/n855 ), .ZN(\AES_ENC/us32/n748 ) );
NAND2_X2 \AES_ENC/us32/U320  ( .A1(\AES_ENC/us32/n956 ), .A2(\AES_ENC/us32/n748 ), .ZN(\AES_ENC/us32/n760 ) );
NAND2_X2 \AES_ENC/us32/U313  ( .A1(\AES_ENC/us32/n590 ), .A2(\AES_ENC/us32/n753 ), .ZN(\AES_ENC/us32/n1023 ) );
NAND4_X2 \AES_ENC/us32/U308  ( .A1(\AES_ENC/us32/n760 ), .A2(\AES_ENC/us32/n992 ), .A3(\AES_ENC/us32/n759 ), .A4(\AES_ENC/us32/n758 ), .ZN(\AES_ENC/us32/n761 ) );
NAND2_X2 \AES_ENC/us32/U307  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n761 ), .ZN(\AES_ENC/us32/n792 ) );
NAND2_X2 \AES_ENC/us32/U306  ( .A1(\AES_ENC/us32/n584 ), .A2(\AES_ENC/us32/n603 ), .ZN(\AES_ENC/us32/n989 ) );
NAND2_X2 \AES_ENC/us32/U305  ( .A1(\AES_ENC/us32/n1050 ), .A2(\AES_ENC/us32/n989 ), .ZN(\AES_ENC/us32/n777 ) );
NAND2_X2 \AES_ENC/us32/U304  ( .A1(\AES_ENC/us32/n1093 ), .A2(\AES_ENC/us32/n762 ), .ZN(\AES_ENC/us32/n776 ) );
XNOR2_X2 \AES_ENC/us32/U301  ( .A(\AES_ENC/sa32 [7]), .B(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n959 ) );
NAND4_X2 \AES_ENC/us32/U289  ( .A1(\AES_ENC/us32/n777 ), .A2(\AES_ENC/us32/n776 ), .A3(\AES_ENC/us32/n775 ), .A4(\AES_ENC/us32/n774 ), .ZN(\AES_ENC/us32/n778 ) );
NAND2_X2 \AES_ENC/us32/U288  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n778 ), .ZN(\AES_ENC/us32/n791 ) );
NAND2_X2 \AES_ENC/us32/U287  ( .A1(\AES_ENC/us32/n1056 ), .A2(\AES_ENC/us32/n1050 ), .ZN(\AES_ENC/us32/n788 ) );
NAND2_X2 \AES_ENC/us32/U286  ( .A1(\AES_ENC/us32/n1091 ), .A2(\AES_ENC/us32/n779 ), .ZN(\AES_ENC/us32/n787 ) );
NAND2_X2 \AES_ENC/us32/U285  ( .A1(\AES_ENC/us32/n956 ), .A2(\AES_ENC/sa32 [1]), .ZN(\AES_ENC/us32/n786 ) );
NAND4_X2 \AES_ENC/us32/U278  ( .A1(\AES_ENC/us32/n788 ), .A2(\AES_ENC/us32/n787 ), .A3(\AES_ENC/us32/n786 ), .A4(\AES_ENC/us32/n785 ), .ZN(\AES_ENC/us32/n789 ) );
NAND2_X2 \AES_ENC/us32/U277  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n789 ), .ZN(\AES_ENC/us32/n790 ) );
NAND4_X2 \AES_ENC/us32/U276  ( .A1(\AES_ENC/us32/n793 ), .A2(\AES_ENC/us32/n792 ), .A3(\AES_ENC/us32/n791 ), .A4(\AES_ENC/us32/n790 ), .ZN(\AES_ENC/sa32_sub[2] ) );
NAND2_X2 \AES_ENC/us32/U275  ( .A1(\AES_ENC/us32/n1059 ), .A2(\AES_ENC/us32/n794 ), .ZN(\AES_ENC/us32/n810 ) );
NAND2_X2 \AES_ENC/us32/U274  ( .A1(\AES_ENC/us32/n1049 ), .A2(\AES_ENC/us32/n956 ), .ZN(\AES_ENC/us32/n809 ) );
OR2_X2 \AES_ENC/us32/U266  ( .A1(\AES_ENC/us32/n1096 ), .A2(\AES_ENC/us32/n606 ), .ZN(\AES_ENC/us32/n802 ) );
NAND2_X2 \AES_ENC/us32/U265  ( .A1(\AES_ENC/us32/n1053 ), .A2(\AES_ENC/us32/n800 ), .ZN(\AES_ENC/us32/n801 ) );
NAND2_X2 \AES_ENC/us32/U264  ( .A1(\AES_ENC/us32/n802 ), .A2(\AES_ENC/us32/n801 ), .ZN(\AES_ENC/us32/n805 ) );
NAND4_X2 \AES_ENC/us32/U261  ( .A1(\AES_ENC/us32/n810 ), .A2(\AES_ENC/us32/n809 ), .A3(\AES_ENC/us32/n808 ), .A4(\AES_ENC/us32/n807 ), .ZN(\AES_ENC/us32/n811 ) );
NAND2_X2 \AES_ENC/us32/U260  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n811 ), .ZN(\AES_ENC/us32/n852 ) );
OR2_X2 \AES_ENC/us32/U259  ( .A1(\AES_ENC/us32/n1023 ), .A2(\AES_ENC/us32/n617 ), .ZN(\AES_ENC/us32/n819 ) );
OR2_X2 \AES_ENC/us32/U257  ( .A1(\AES_ENC/us32/n570 ), .A2(\AES_ENC/us32/n930 ), .ZN(\AES_ENC/us32/n818 ) );
NAND2_X2 \AES_ENC/us32/U256  ( .A1(\AES_ENC/us32/n1013 ), .A2(\AES_ENC/us32/n1094 ), .ZN(\AES_ENC/us32/n817 ) );
NAND4_X2 \AES_ENC/us32/U249  ( .A1(\AES_ENC/us32/n819 ), .A2(\AES_ENC/us32/n818 ), .A3(\AES_ENC/us32/n817 ), .A4(\AES_ENC/us32/n816 ), .ZN(\AES_ENC/us32/n820 ) );
NAND2_X2 \AES_ENC/us32/U248  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n820 ), .ZN(\AES_ENC/us32/n851 ) );
NAND2_X2 \AES_ENC/us32/U247  ( .A1(\AES_ENC/us32/n956 ), .A2(\AES_ENC/us32/n1080 ), .ZN(\AES_ENC/us32/n835 ) );
NAND2_X2 \AES_ENC/us32/U246  ( .A1(\AES_ENC/us32/n570 ), .A2(\AES_ENC/us32/n1030 ), .ZN(\AES_ENC/us32/n1047 ) );
OR2_X2 \AES_ENC/us32/U245  ( .A1(\AES_ENC/us32/n1047 ), .A2(\AES_ENC/us32/n612 ), .ZN(\AES_ENC/us32/n834 ) );
NAND2_X2 \AES_ENC/us32/U244  ( .A1(\AES_ENC/us32/n1072 ), .A2(\AES_ENC/us32/n589 ), .ZN(\AES_ENC/us32/n833 ) );
NAND4_X2 \AES_ENC/us32/U233  ( .A1(\AES_ENC/us32/n835 ), .A2(\AES_ENC/us32/n834 ), .A3(\AES_ENC/us32/n833 ), .A4(\AES_ENC/us32/n832 ), .ZN(\AES_ENC/us32/n836 ) );
NAND2_X2 \AES_ENC/us32/U232  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n836 ), .ZN(\AES_ENC/us32/n850 ) );
NAND2_X2 \AES_ENC/us32/U231  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n623 ), .ZN(\AES_ENC/us32/n847 ) );
NAND2_X2 \AES_ENC/us32/U230  ( .A1(\AES_ENC/us32/n1050 ), .A2(\AES_ENC/us32/n1071 ), .ZN(\AES_ENC/us32/n846 ) );
OR2_X2 \AES_ENC/us32/U224  ( .A1(\AES_ENC/us32/n1053 ), .A2(\AES_ENC/us32/n911 ), .ZN(\AES_ENC/us32/n1077 ) );
NAND4_X2 \AES_ENC/us32/U220  ( .A1(\AES_ENC/us32/n847 ), .A2(\AES_ENC/us32/n846 ), .A3(\AES_ENC/us32/n845 ), .A4(\AES_ENC/us32/n844 ), .ZN(\AES_ENC/us32/n848 ) );
NAND2_X2 \AES_ENC/us32/U219  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n848 ), .ZN(\AES_ENC/us32/n849 ) );
NAND4_X2 \AES_ENC/us32/U218  ( .A1(\AES_ENC/us32/n852 ), .A2(\AES_ENC/us32/n851 ), .A3(\AES_ENC/us32/n850 ), .A4(\AES_ENC/us32/n849 ), .ZN(\AES_ENC/sa32_sub[3] ) );
NAND2_X2 \AES_ENC/us32/U216  ( .A1(\AES_ENC/us32/n1009 ), .A2(\AES_ENC/us32/n1072 ), .ZN(\AES_ENC/us32/n862 ) );
NAND2_X2 \AES_ENC/us32/U215  ( .A1(\AES_ENC/us32/n603 ), .A2(\AES_ENC/us32/n577 ), .ZN(\AES_ENC/us32/n853 ) );
NAND2_X2 \AES_ENC/us32/U214  ( .A1(\AES_ENC/us32/n1050 ), .A2(\AES_ENC/us32/n853 ), .ZN(\AES_ENC/us32/n861 ) );
NAND4_X2 \AES_ENC/us32/U206  ( .A1(\AES_ENC/us32/n862 ), .A2(\AES_ENC/us32/n861 ), .A3(\AES_ENC/us32/n860 ), .A4(\AES_ENC/us32/n859 ), .ZN(\AES_ENC/us32/n863 ) );
NAND2_X2 \AES_ENC/us32/U205  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n863 ), .ZN(\AES_ENC/us32/n905 ) );
NAND2_X2 \AES_ENC/us32/U204  ( .A1(\AES_ENC/us32/n1010 ), .A2(\AES_ENC/us32/n989 ), .ZN(\AES_ENC/us32/n874 ) );
NAND2_X2 \AES_ENC/us32/U203  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n610 ), .ZN(\AES_ENC/us32/n864 ) );
NAND2_X2 \AES_ENC/us32/U202  ( .A1(\AES_ENC/us32/n929 ), .A2(\AES_ENC/us32/n864 ), .ZN(\AES_ENC/us32/n873 ) );
NAND4_X2 \AES_ENC/us32/U193  ( .A1(\AES_ENC/us32/n874 ), .A2(\AES_ENC/us32/n873 ), .A3(\AES_ENC/us32/n872 ), .A4(\AES_ENC/us32/n871 ), .ZN(\AES_ENC/us32/n875 ) );
NAND2_X2 \AES_ENC/us32/U192  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n875 ), .ZN(\AES_ENC/us32/n904 ) );
NAND2_X2 \AES_ENC/us32/U191  ( .A1(\AES_ENC/us32/n583 ), .A2(\AES_ENC/us32/n1050 ), .ZN(\AES_ENC/us32/n889 ) );
NAND2_X2 \AES_ENC/us32/U190  ( .A1(\AES_ENC/us32/n1093 ), .A2(\AES_ENC/us32/n587 ), .ZN(\AES_ENC/us32/n876 ) );
NAND2_X2 \AES_ENC/us32/U189  ( .A1(\AES_ENC/us32/n604 ), .A2(\AES_ENC/us32/n876 ), .ZN(\AES_ENC/us32/n877 ) );
NAND2_X2 \AES_ENC/us32/U188  ( .A1(\AES_ENC/us32/n877 ), .A2(\AES_ENC/us32/n623 ), .ZN(\AES_ENC/us32/n888 ) );
NAND4_X2 \AES_ENC/us32/U179  ( .A1(\AES_ENC/us32/n889 ), .A2(\AES_ENC/us32/n888 ), .A3(\AES_ENC/us32/n887 ), .A4(\AES_ENC/us32/n886 ), .ZN(\AES_ENC/us32/n890 ) );
NAND2_X2 \AES_ENC/us32/U178  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n890 ), .ZN(\AES_ENC/us32/n903 ) );
OR2_X2 \AES_ENC/us32/U177  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n1059 ), .ZN(\AES_ENC/us32/n900 ) );
NAND2_X2 \AES_ENC/us32/U176  ( .A1(\AES_ENC/us32/n1073 ), .A2(\AES_ENC/us32/n1047 ), .ZN(\AES_ENC/us32/n899 ) );
NAND2_X2 \AES_ENC/us32/U175  ( .A1(\AES_ENC/us32/n1094 ), .A2(\AES_ENC/us32/n595 ), .ZN(\AES_ENC/us32/n898 ) );
NAND4_X2 \AES_ENC/us32/U167  ( .A1(\AES_ENC/us32/n900 ), .A2(\AES_ENC/us32/n899 ), .A3(\AES_ENC/us32/n898 ), .A4(\AES_ENC/us32/n897 ), .ZN(\AES_ENC/us32/n901 ) );
NAND2_X2 \AES_ENC/us32/U166  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n901 ), .ZN(\AES_ENC/us32/n902 ) );
NAND4_X2 \AES_ENC/us32/U165  ( .A1(\AES_ENC/us32/n905 ), .A2(\AES_ENC/us32/n904 ), .A3(\AES_ENC/us32/n903 ), .A4(\AES_ENC/us32/n902 ), .ZN(\AES_ENC/sa32_sub[4] ) );
NAND2_X2 \AES_ENC/us32/U164  ( .A1(\AES_ENC/us32/n1094 ), .A2(\AES_ENC/us32/n599 ), .ZN(\AES_ENC/us32/n922 ) );
NAND2_X2 \AES_ENC/us32/U163  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n989 ), .ZN(\AES_ENC/us32/n921 ) );
NAND4_X2 \AES_ENC/us32/U151  ( .A1(\AES_ENC/us32/n922 ), .A2(\AES_ENC/us32/n921 ), .A3(\AES_ENC/us32/n920 ), .A4(\AES_ENC/us32/n919 ), .ZN(\AES_ENC/us32/n923 ) );
NAND2_X2 \AES_ENC/us32/U150  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n923 ), .ZN(\AES_ENC/us32/n972 ) );
NAND2_X2 \AES_ENC/us32/U149  ( .A1(\AES_ENC/us32/n582 ), .A2(\AES_ENC/us32/n619 ), .ZN(\AES_ENC/us32/n924 ) );
NAND2_X2 \AES_ENC/us32/U148  ( .A1(\AES_ENC/us32/n1073 ), .A2(\AES_ENC/us32/n924 ), .ZN(\AES_ENC/us32/n939 ) );
NAND2_X2 \AES_ENC/us32/U147  ( .A1(\AES_ENC/us32/n926 ), .A2(\AES_ENC/us32/n925 ), .ZN(\AES_ENC/us32/n927 ) );
NAND2_X2 \AES_ENC/us32/U146  ( .A1(\AES_ENC/us32/n606 ), .A2(\AES_ENC/us32/n927 ), .ZN(\AES_ENC/us32/n928 ) );
NAND2_X2 \AES_ENC/us32/U145  ( .A1(\AES_ENC/us32/n928 ), .A2(\AES_ENC/us32/n1080 ), .ZN(\AES_ENC/us32/n938 ) );
OR2_X2 \AES_ENC/us32/U144  ( .A1(\AES_ENC/us32/n1117 ), .A2(\AES_ENC/us32/n615 ), .ZN(\AES_ENC/us32/n937 ) );
NAND4_X2 \AES_ENC/us32/U139  ( .A1(\AES_ENC/us32/n939 ), .A2(\AES_ENC/us32/n938 ), .A3(\AES_ENC/us32/n937 ), .A4(\AES_ENC/us32/n936 ), .ZN(\AES_ENC/us32/n940 ) );
NAND2_X2 \AES_ENC/us32/U138  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n940 ), .ZN(\AES_ENC/us32/n971 ) );
OR2_X2 \AES_ENC/us32/U137  ( .A1(\AES_ENC/us32/n605 ), .A2(\AES_ENC/us32/n941 ), .ZN(\AES_ENC/us32/n954 ) );
NAND2_X2 \AES_ENC/us32/U136  ( .A1(\AES_ENC/us32/n1096 ), .A2(\AES_ENC/us32/n577 ), .ZN(\AES_ENC/us32/n942 ) );
NAND2_X2 \AES_ENC/us32/U135  ( .A1(\AES_ENC/us32/n1048 ), .A2(\AES_ENC/us32/n942 ), .ZN(\AES_ENC/us32/n943 ) );
NAND2_X2 \AES_ENC/us32/U134  ( .A1(\AES_ENC/us32/n612 ), .A2(\AES_ENC/us32/n943 ), .ZN(\AES_ENC/us32/n944 ) );
NAND2_X2 \AES_ENC/us32/U133  ( .A1(\AES_ENC/us32/n944 ), .A2(\AES_ENC/us32/n580 ), .ZN(\AES_ENC/us32/n953 ) );
NAND4_X2 \AES_ENC/us32/U125  ( .A1(\AES_ENC/us32/n954 ), .A2(\AES_ENC/us32/n953 ), .A3(\AES_ENC/us32/n952 ), .A4(\AES_ENC/us32/n951 ), .ZN(\AES_ENC/us32/n955 ) );
NAND2_X2 \AES_ENC/us32/U124  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n955 ), .ZN(\AES_ENC/us32/n970 ) );
NAND2_X2 \AES_ENC/us32/U123  ( .A1(\AES_ENC/us32/n1094 ), .A2(\AES_ENC/us32/n1071 ), .ZN(\AES_ENC/us32/n967 ) );
NAND2_X2 \AES_ENC/us32/U122  ( .A1(\AES_ENC/us32/n956 ), .A2(\AES_ENC/us32/n1030 ), .ZN(\AES_ENC/us32/n966 ) );
NAND4_X2 \AES_ENC/us32/U114  ( .A1(\AES_ENC/us32/n967 ), .A2(\AES_ENC/us32/n966 ), .A3(\AES_ENC/us32/n965 ), .A4(\AES_ENC/us32/n964 ), .ZN(\AES_ENC/us32/n968 ) );
NAND2_X2 \AES_ENC/us32/U113  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n968 ), .ZN(\AES_ENC/us32/n969 ) );
NAND4_X2 \AES_ENC/us32/U112  ( .A1(\AES_ENC/us32/n972 ), .A2(\AES_ENC/us32/n971 ), .A3(\AES_ENC/us32/n970 ), .A4(\AES_ENC/us32/n969 ), .ZN(\AES_ENC/sa32_sub[5] ) );
NAND2_X2 \AES_ENC/us32/U111  ( .A1(\AES_ENC/us32/n570 ), .A2(\AES_ENC/us32/n1097 ), .ZN(\AES_ENC/us32/n973 ) );
NAND2_X2 \AES_ENC/us32/U110  ( .A1(\AES_ENC/us32/n1073 ), .A2(\AES_ENC/us32/n973 ), .ZN(\AES_ENC/us32/n987 ) );
NAND2_X2 \AES_ENC/us32/U109  ( .A1(\AES_ENC/us32/n974 ), .A2(\AES_ENC/us32/n1077 ), .ZN(\AES_ENC/us32/n975 ) );
NAND2_X2 \AES_ENC/us32/U108  ( .A1(\AES_ENC/us32/n613 ), .A2(\AES_ENC/us32/n975 ), .ZN(\AES_ENC/us32/n976 ) );
NAND2_X2 \AES_ENC/us32/U107  ( .A1(\AES_ENC/us32/n977 ), .A2(\AES_ENC/us32/n976 ), .ZN(\AES_ENC/us32/n986 ) );
NAND4_X2 \AES_ENC/us32/U99  ( .A1(\AES_ENC/us32/n987 ), .A2(\AES_ENC/us32/n986 ), .A3(\AES_ENC/us32/n985 ), .A4(\AES_ENC/us32/n984 ), .ZN(\AES_ENC/us32/n988 ) );
NAND2_X2 \AES_ENC/us32/U98  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n988 ), .ZN(\AES_ENC/us32/n1044 ) );
NAND2_X2 \AES_ENC/us32/U97  ( .A1(\AES_ENC/us32/n1073 ), .A2(\AES_ENC/us32/n989 ), .ZN(\AES_ENC/us32/n1004 ) );
NAND2_X2 \AES_ENC/us32/U96  ( .A1(\AES_ENC/us32/n1092 ), .A2(\AES_ENC/us32/n619 ), .ZN(\AES_ENC/us32/n1003 ) );
NAND4_X2 \AES_ENC/us32/U85  ( .A1(\AES_ENC/us32/n1004 ), .A2(\AES_ENC/us32/n1003 ), .A3(\AES_ENC/us32/n1002 ), .A4(\AES_ENC/us32/n1001 ), .ZN(\AES_ENC/us32/n1005 ) );
NAND2_X2 \AES_ENC/us32/U84  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n1005 ), .ZN(\AES_ENC/us32/n1043 ) );
NAND2_X2 \AES_ENC/us32/U83  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n596 ), .ZN(\AES_ENC/us32/n1020 ) );
NAND2_X2 \AES_ENC/us32/U82  ( .A1(\AES_ENC/us32/n1050 ), .A2(\AES_ENC/us32/n624 ), .ZN(\AES_ENC/us32/n1019 ) );
NAND2_X2 \AES_ENC/us32/U77  ( .A1(\AES_ENC/us32/n1059 ), .A2(\AES_ENC/us32/n1114 ), .ZN(\AES_ENC/us32/n1012 ) );
NAND2_X2 \AES_ENC/us32/U76  ( .A1(\AES_ENC/us32/n1010 ), .A2(\AES_ENC/us32/n592 ), .ZN(\AES_ENC/us32/n1011 ) );
NAND2_X2 \AES_ENC/us32/U75  ( .A1(\AES_ENC/us32/n1012 ), .A2(\AES_ENC/us32/n1011 ), .ZN(\AES_ENC/us32/n1016 ) );
NAND4_X2 \AES_ENC/us32/U70  ( .A1(\AES_ENC/us32/n1020 ), .A2(\AES_ENC/us32/n1019 ), .A3(\AES_ENC/us32/n1018 ), .A4(\AES_ENC/us32/n1017 ), .ZN(\AES_ENC/us32/n1021 ) );
NAND2_X2 \AES_ENC/us32/U69  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n1021 ), .ZN(\AES_ENC/us32/n1042 ) );
NAND2_X2 \AES_ENC/us32/U68  ( .A1(\AES_ENC/us32/n1022 ), .A2(\AES_ENC/us32/n1093 ), .ZN(\AES_ENC/us32/n1039 ) );
NAND2_X2 \AES_ENC/us32/U67  ( .A1(\AES_ENC/us32/n1050 ), .A2(\AES_ENC/us32/n1023 ), .ZN(\AES_ENC/us32/n1038 ) );
NAND2_X2 \AES_ENC/us32/U66  ( .A1(\AES_ENC/us32/n1024 ), .A2(\AES_ENC/us32/n1071 ), .ZN(\AES_ENC/us32/n1037 ) );
AND2_X2 \AES_ENC/us32/U60  ( .A1(\AES_ENC/us32/n1030 ), .A2(\AES_ENC/us32/n602 ), .ZN(\AES_ENC/us32/n1078 ) );
NAND4_X2 \AES_ENC/us32/U56  ( .A1(\AES_ENC/us32/n1039 ), .A2(\AES_ENC/us32/n1038 ), .A3(\AES_ENC/us32/n1037 ), .A4(\AES_ENC/us32/n1036 ), .ZN(\AES_ENC/us32/n1040 ) );
NAND2_X2 \AES_ENC/us32/U55  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n1040 ), .ZN(\AES_ENC/us32/n1041 ) );
NAND4_X2 \AES_ENC/us32/U54  ( .A1(\AES_ENC/us32/n1044 ), .A2(\AES_ENC/us32/n1043 ), .A3(\AES_ENC/us32/n1042 ), .A4(\AES_ENC/us32/n1041 ), .ZN(\AES_ENC/sa32_sub[6] ) );
NAND2_X2 \AES_ENC/us32/U53  ( .A1(\AES_ENC/us32/n1072 ), .A2(\AES_ENC/us32/n1045 ), .ZN(\AES_ENC/us32/n1068 ) );
NAND2_X2 \AES_ENC/us32/U52  ( .A1(\AES_ENC/us32/n1046 ), .A2(\AES_ENC/us32/n582 ), .ZN(\AES_ENC/us32/n1067 ) );
NAND2_X2 \AES_ENC/us32/U51  ( .A1(\AES_ENC/us32/n1094 ), .A2(\AES_ENC/us32/n1047 ), .ZN(\AES_ENC/us32/n1066 ) );
NAND4_X2 \AES_ENC/us32/U40  ( .A1(\AES_ENC/us32/n1068 ), .A2(\AES_ENC/us32/n1067 ), .A3(\AES_ENC/us32/n1066 ), .A4(\AES_ENC/us32/n1065 ), .ZN(\AES_ENC/us32/n1069 ) );
NAND2_X2 \AES_ENC/us32/U39  ( .A1(\AES_ENC/us32/n1070 ), .A2(\AES_ENC/us32/n1069 ), .ZN(\AES_ENC/us32/n1135 ) );
NAND2_X2 \AES_ENC/us32/U38  ( .A1(\AES_ENC/us32/n1072 ), .A2(\AES_ENC/us32/n1071 ), .ZN(\AES_ENC/us32/n1088 ) );
NAND2_X2 \AES_ENC/us32/U37  ( .A1(\AES_ENC/us32/n1073 ), .A2(\AES_ENC/us32/n595 ), .ZN(\AES_ENC/us32/n1087 ) );
NAND4_X2 \AES_ENC/us32/U28  ( .A1(\AES_ENC/us32/n1088 ), .A2(\AES_ENC/us32/n1087 ), .A3(\AES_ENC/us32/n1086 ), .A4(\AES_ENC/us32/n1085 ), .ZN(\AES_ENC/us32/n1089 ) );
NAND2_X2 \AES_ENC/us32/U27  ( .A1(\AES_ENC/us32/n1090 ), .A2(\AES_ENC/us32/n1089 ), .ZN(\AES_ENC/us32/n1134 ) );
NAND2_X2 \AES_ENC/us32/U26  ( .A1(\AES_ENC/us32/n1091 ), .A2(\AES_ENC/us32/n1093 ), .ZN(\AES_ENC/us32/n1111 ) );
NAND2_X2 \AES_ENC/us32/U25  ( .A1(\AES_ENC/us32/n1092 ), .A2(\AES_ENC/us32/n1120 ), .ZN(\AES_ENC/us32/n1110 ) );
AND2_X2 \AES_ENC/us32/U22  ( .A1(\AES_ENC/us32/n1097 ), .A2(\AES_ENC/us32/n1096 ), .ZN(\AES_ENC/us32/n1098 ) );
NAND4_X2 \AES_ENC/us32/U14  ( .A1(\AES_ENC/us32/n1111 ), .A2(\AES_ENC/us32/n1110 ), .A3(\AES_ENC/us32/n1109 ), .A4(\AES_ENC/us32/n1108 ), .ZN(\AES_ENC/us32/n1112 ) );
NAND2_X2 \AES_ENC/us32/U13  ( .A1(\AES_ENC/us32/n1113 ), .A2(\AES_ENC/us32/n1112 ), .ZN(\AES_ENC/us32/n1133 ) );
NAND2_X2 \AES_ENC/us32/U12  ( .A1(\AES_ENC/us32/n1115 ), .A2(\AES_ENC/us32/n1114 ), .ZN(\AES_ENC/us32/n1129 ) );
OR2_X2 \AES_ENC/us32/U11  ( .A1(\AES_ENC/us32/n608 ), .A2(\AES_ENC/us32/n1116 ), .ZN(\AES_ENC/us32/n1128 ) );
NAND4_X2 \AES_ENC/us32/U3  ( .A1(\AES_ENC/us32/n1129 ), .A2(\AES_ENC/us32/n1128 ), .A3(\AES_ENC/us32/n1127 ), .A4(\AES_ENC/us32/n1126 ), .ZN(\AES_ENC/us32/n1130 ) );
NAND2_X2 \AES_ENC/us32/U2  ( .A1(\AES_ENC/us32/n1131 ), .A2(\AES_ENC/us32/n1130 ), .ZN(\AES_ENC/us32/n1132 ) );
NAND4_X2 \AES_ENC/us32/U1  ( .A1(\AES_ENC/us32/n1135 ), .A2(\AES_ENC/us32/n1134 ), .A3(\AES_ENC/us32/n1133 ), .A4(\AES_ENC/us32/n1132 ), .ZN(\AES_ENC/sa32_sub[7] ) );
INV_X4 \AES_ENC/us33/U575  ( .A(\AES_ENC/sa33 [7]), .ZN(\AES_ENC/us33/n627 ));
INV_X4 \AES_ENC/us33/U574  ( .A(\AES_ENC/us33/n1114 ), .ZN(\AES_ENC/us33/n625 ) );
INV_X4 \AES_ENC/us33/U573  ( .A(\AES_ENC/sa33 [4]), .ZN(\AES_ENC/us33/n624 ));
INV_X4 \AES_ENC/us33/U572  ( .A(\AES_ENC/us33/n1025 ), .ZN(\AES_ENC/us33/n622 ) );
INV_X4 \AES_ENC/us33/U571  ( .A(\AES_ENC/us33/n1120 ), .ZN(\AES_ENC/us33/n620 ) );
INV_X4 \AES_ENC/us33/U570  ( .A(\AES_ENC/us33/n1121 ), .ZN(\AES_ENC/us33/n619 ) );
INV_X4 \AES_ENC/us33/U569  ( .A(\AES_ENC/us33/n1048 ), .ZN(\AES_ENC/us33/n618 ) );
INV_X4 \AES_ENC/us33/U568  ( .A(\AES_ENC/us33/n974 ), .ZN(\AES_ENC/us33/n616 ) );
INV_X4 \AES_ENC/us33/U567  ( .A(\AES_ENC/us33/n794 ), .ZN(\AES_ENC/us33/n614 ) );
INV_X4 \AES_ENC/us33/U566  ( .A(\AES_ENC/sa33 [2]), .ZN(\AES_ENC/us33/n611 ));
INV_X4 \AES_ENC/us33/U565  ( .A(\AES_ENC/us33/n800 ), .ZN(\AES_ENC/us33/n610 ) );
INV_X4 \AES_ENC/us33/U564  ( .A(\AES_ENC/us33/n925 ), .ZN(\AES_ENC/us33/n609 ) );
INV_X4 \AES_ENC/us33/U563  ( .A(\AES_ENC/us33/n779 ), .ZN(\AES_ENC/us33/n607 ) );
INV_X4 \AES_ENC/us33/U562  ( .A(\AES_ENC/us33/n1022 ), .ZN(\AES_ENC/us33/n603 ) );
INV_X4 \AES_ENC/us33/U561  ( .A(\AES_ENC/us33/n1102 ), .ZN(\AES_ENC/us33/n602 ) );
INV_X4 \AES_ENC/us33/U560  ( .A(\AES_ENC/us33/n929 ), .ZN(\AES_ENC/us33/n601 ) );
INV_X4 \AES_ENC/us33/U559  ( .A(\AES_ENC/us33/n1056 ), .ZN(\AES_ENC/us33/n600 ) );
INV_X4 \AES_ENC/us33/U558  ( .A(\AES_ENC/us33/n1054 ), .ZN(\AES_ENC/us33/n599 ) );
INV_X4 \AES_ENC/us33/U557  ( .A(\AES_ENC/us33/n881 ), .ZN(\AES_ENC/us33/n598 ) );
INV_X4 \AES_ENC/us33/U556  ( .A(\AES_ENC/us33/n926 ), .ZN(\AES_ENC/us33/n597 ) );
INV_X4 \AES_ENC/us33/U555  ( .A(\AES_ENC/us33/n977 ), .ZN(\AES_ENC/us33/n595 ) );
INV_X4 \AES_ENC/us33/U554  ( .A(\AES_ENC/us33/n1031 ), .ZN(\AES_ENC/us33/n594 ) );
INV_X4 \AES_ENC/us33/U553  ( .A(\AES_ENC/us33/n1103 ), .ZN(\AES_ENC/us33/n593 ) );
INV_X4 \AES_ENC/us33/U552  ( .A(\AES_ENC/us33/n1009 ), .ZN(\AES_ENC/us33/n592 ) );
INV_X4 \AES_ENC/us33/U551  ( .A(\AES_ENC/us33/n990 ), .ZN(\AES_ENC/us33/n591 ) );
INV_X4 \AES_ENC/us33/U550  ( .A(\AES_ENC/us33/n1058 ), .ZN(\AES_ENC/us33/n590 ) );
INV_X4 \AES_ENC/us33/U549  ( .A(\AES_ENC/us33/n1074 ), .ZN(\AES_ENC/us33/n589 ) );
INV_X4 \AES_ENC/us33/U548  ( .A(\AES_ENC/us33/n1053 ), .ZN(\AES_ENC/us33/n588 ) );
INV_X4 \AES_ENC/us33/U547  ( .A(\AES_ENC/us33/n826 ), .ZN(\AES_ENC/us33/n587 ) );
INV_X4 \AES_ENC/us33/U546  ( .A(\AES_ENC/us33/n992 ), .ZN(\AES_ENC/us33/n586 ) );
INV_X4 \AES_ENC/us33/U545  ( .A(\AES_ENC/us33/n821 ), .ZN(\AES_ENC/us33/n585 ) );
INV_X4 \AES_ENC/us33/U544  ( .A(\AES_ENC/us33/n910 ), .ZN(\AES_ENC/us33/n584 ) );
INV_X4 \AES_ENC/us33/U543  ( .A(\AES_ENC/us33/n906 ), .ZN(\AES_ENC/us33/n583 ) );
INV_X4 \AES_ENC/us33/U542  ( .A(\AES_ENC/us33/n880 ), .ZN(\AES_ENC/us33/n581 ) );
INV_X4 \AES_ENC/us33/U541  ( .A(\AES_ENC/us33/n1013 ), .ZN(\AES_ENC/us33/n580 ) );
INV_X4 \AES_ENC/us33/U540  ( .A(\AES_ENC/us33/n1092 ), .ZN(\AES_ENC/us33/n579 ) );
INV_X4 \AES_ENC/us33/U539  ( .A(\AES_ENC/us33/n824 ), .ZN(\AES_ENC/us33/n578 ) );
INV_X4 \AES_ENC/us33/U538  ( .A(\AES_ENC/us33/n1091 ), .ZN(\AES_ENC/us33/n577 ) );
INV_X4 \AES_ENC/us33/U537  ( .A(\AES_ENC/us33/n1080 ), .ZN(\AES_ENC/us33/n576 ) );
INV_X4 \AES_ENC/us33/U536  ( .A(\AES_ENC/us33/n959 ), .ZN(\AES_ENC/us33/n575 ) );
INV_X4 \AES_ENC/us33/U535  ( .A(\AES_ENC/sa33 [0]), .ZN(\AES_ENC/us33/n574 ));
NOR2_X2 \AES_ENC/us33/U534  ( .A1(\AES_ENC/sa33 [0]), .A2(\AES_ENC/sa33 [6]),.ZN(\AES_ENC/us33/n1090 ) );
NOR2_X2 \AES_ENC/us33/U533  ( .A1(\AES_ENC/us33/n574 ), .A2(\AES_ENC/sa33 [6]), .ZN(\AES_ENC/us33/n1070 ) );
NOR2_X2 \AES_ENC/us33/U532  ( .A1(\AES_ENC/sa33 [4]), .A2(\AES_ENC/sa33 [3]),.ZN(\AES_ENC/us33/n1025 ) );
INV_X4 \AES_ENC/us33/U531  ( .A(\AES_ENC/us33/n569 ), .ZN(\AES_ENC/us33/n572 ) );
NOR2_X2 \AES_ENC/us33/U530  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n765 ) );
NOR2_X2 \AES_ENC/us33/U529  ( .A1(\AES_ENC/sa33 [4]), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n764 ) );
NOR2_X2 \AES_ENC/us33/U528  ( .A1(\AES_ENC/us33/n765 ), .A2(\AES_ENC/us33/n764 ), .ZN(\AES_ENC/us33/n766 ) );
NOR2_X2 \AES_ENC/us33/U527  ( .A1(\AES_ENC/us33/n766 ), .A2(\AES_ENC/us33/n575 ), .ZN(\AES_ENC/us33/n767 ) );
NOR3_X2 \AES_ENC/us33/U526  ( .A1(\AES_ENC/us33/n627 ), .A2(\AES_ENC/sa33 [5]), .A3(\AES_ENC/us33/n704 ), .ZN(\AES_ENC/us33/n706 ));
NOR2_X2 \AES_ENC/us33/U525  ( .A1(\AES_ENC/us33/n1117 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n707 ) );
NOR2_X2 \AES_ENC/us33/U524  ( .A1(\AES_ENC/sa33 [4]), .A2(\AES_ENC/us33/n579 ), .ZN(\AES_ENC/us33/n705 ) );
NOR3_X2 \AES_ENC/us33/U523  ( .A1(\AES_ENC/us33/n707 ), .A2(\AES_ENC/us33/n706 ), .A3(\AES_ENC/us33/n705 ), .ZN(\AES_ENC/us33/n713 ) );
INV_X4 \AES_ENC/us33/U522  ( .A(\AES_ENC/sa33 [3]), .ZN(\AES_ENC/us33/n621 ));
NAND3_X2 \AES_ENC/us33/U521  ( .A1(\AES_ENC/us33/n652 ), .A2(\AES_ENC/us33/n626 ), .A3(\AES_ENC/sa33 [7]), .ZN(\AES_ENC/us33/n653 ));
NOR2_X2 \AES_ENC/us33/U520  ( .A1(\AES_ENC/us33/n611 ), .A2(\AES_ENC/sa33 [5]), .ZN(\AES_ENC/us33/n925 ) );
NOR2_X2 \AES_ENC/us33/U519  ( .A1(\AES_ENC/sa33 [5]), .A2(\AES_ENC/sa33 [2]),.ZN(\AES_ENC/us33/n974 ) );
INV_X4 \AES_ENC/us33/U518  ( .A(\AES_ENC/sa33 [5]), .ZN(\AES_ENC/us33/n626 ));
NOR2_X2 \AES_ENC/us33/U517  ( .A1(\AES_ENC/us33/n611 ), .A2(\AES_ENC/sa33 [7]), .ZN(\AES_ENC/us33/n779 ) );
NAND3_X2 \AES_ENC/us33/U516  ( .A1(\AES_ENC/us33/n679 ), .A2(\AES_ENC/us33/n678 ), .A3(\AES_ENC/us33/n677 ), .ZN(\AES_ENC/sa33_sub[0] ) );
NOR2_X2 \AES_ENC/us33/U515  ( .A1(\AES_ENC/us33/n626 ), .A2(\AES_ENC/sa33 [2]), .ZN(\AES_ENC/us33/n1048 ) );
NOR4_X2 \AES_ENC/us33/U512  ( .A1(\AES_ENC/us33/n633 ), .A2(\AES_ENC/us33/n632 ), .A3(\AES_ENC/us33/n631 ), .A4(\AES_ENC/us33/n630 ), .ZN(\AES_ENC/us33/n634 ) );
NOR2_X2 \AES_ENC/us33/U510  ( .A1(\AES_ENC/us33/n629 ), .A2(\AES_ENC/us33/n628 ), .ZN(\AES_ENC/us33/n635 ) );
NAND3_X2 \AES_ENC/us33/U509  ( .A1(\AES_ENC/sa33 [2]), .A2(\AES_ENC/sa33 [7]), .A3(\AES_ENC/us33/n1059 ), .ZN(\AES_ENC/us33/n636 ) );
NOR2_X2 \AES_ENC/us33/U508  ( .A1(\AES_ENC/sa33 [7]), .A2(\AES_ENC/sa33 [2]),.ZN(\AES_ENC/us33/n794 ) );
NOR2_X2 \AES_ENC/us33/U507  ( .A1(\AES_ENC/sa33 [4]), .A2(\AES_ENC/sa33 [1]),.ZN(\AES_ENC/us33/n1102 ) );
NOR2_X2 \AES_ENC/us33/U506  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/sa33 [3]), .ZN(\AES_ENC/us33/n1053 ) );
NOR2_X2 \AES_ENC/us33/U505  ( .A1(\AES_ENC/us33/n607 ), .A2(\AES_ENC/sa33 [5]), .ZN(\AES_ENC/us33/n1024 ) );
NOR2_X2 \AES_ENC/us33/U504  ( .A1(\AES_ENC/us33/n625 ), .A2(\AES_ENC/sa33 [2]), .ZN(\AES_ENC/us33/n1093 ) );
NOR2_X2 \AES_ENC/us33/U503  ( .A1(\AES_ENC/us33/n614 ), .A2(\AES_ENC/sa33 [5]), .ZN(\AES_ENC/us33/n1094 ) );
NOR2_X2 \AES_ENC/us33/U502  ( .A1(\AES_ENC/us33/n624 ), .A2(\AES_ENC/sa33 [3]), .ZN(\AES_ENC/us33/n931 ) );
INV_X4 \AES_ENC/us33/U501  ( .A(\AES_ENC/us33/n570 ), .ZN(\AES_ENC/us33/n573 ) );
NOR2_X2 \AES_ENC/us33/U500  ( .A1(\AES_ENC/us33/n1053 ), .A2(\AES_ENC/us33/n1095 ), .ZN(\AES_ENC/us33/n639 ) );
NOR3_X2 \AES_ENC/us33/U499  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n573 ), .A3(\AES_ENC/us33/n1074 ), .ZN(\AES_ENC/us33/n641 ) );
NOR2_X2 \AES_ENC/us33/U498  ( .A1(\AES_ENC/us33/n639 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n640 ) );
NOR2_X2 \AES_ENC/us33/U497  ( .A1(\AES_ENC/us33/n641 ), .A2(\AES_ENC/us33/n640 ), .ZN(\AES_ENC/us33/n646 ) );
NOR3_X2 \AES_ENC/us33/U496  ( .A1(\AES_ENC/us33/n995 ), .A2(\AES_ENC/us33/n586 ), .A3(\AES_ENC/us33/n994 ), .ZN(\AES_ENC/us33/n1002 ) );
NOR2_X2 \AES_ENC/us33/U495  ( .A1(\AES_ENC/us33/n909 ), .A2(\AES_ENC/us33/n908 ), .ZN(\AES_ENC/us33/n920 ) );
NOR2_X2 \AES_ENC/us33/U494  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n823 ) );
NOR2_X2 \AES_ENC/us33/U492  ( .A1(\AES_ENC/us33/n624 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n822 ) );
NOR2_X2 \AES_ENC/us33/U491  ( .A1(\AES_ENC/us33/n823 ), .A2(\AES_ENC/us33/n822 ), .ZN(\AES_ENC/us33/n825 ) );
NOR2_X2 \AES_ENC/us33/U490  ( .A1(\AES_ENC/sa33 [1]), .A2(\AES_ENC/us33/n623 ), .ZN(\AES_ENC/us33/n913 ) );
NOR2_X2 \AES_ENC/us33/U489  ( .A1(\AES_ENC/us33/n913 ), .A2(\AES_ENC/us33/n1091 ), .ZN(\AES_ENC/us33/n914 ) );
NOR2_X2 \AES_ENC/us33/U488  ( .A1(\AES_ENC/us33/n826 ), .A2(\AES_ENC/us33/n572 ), .ZN(\AES_ENC/us33/n827 ) );
NOR3_X2 \AES_ENC/us33/U487  ( .A1(\AES_ENC/us33/n769 ), .A2(\AES_ENC/us33/n768 ), .A3(\AES_ENC/us33/n767 ), .ZN(\AES_ENC/us33/n775 ) );
NOR2_X2 \AES_ENC/us33/U486  ( .A1(\AES_ENC/us33/n1056 ), .A2(\AES_ENC/us33/n1053 ), .ZN(\AES_ENC/us33/n749 ) );
NOR2_X2 \AES_ENC/us33/U483  ( .A1(\AES_ENC/us33/n749 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n752 ) );
INV_X4 \AES_ENC/us33/U482  ( .A(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n596 ));
NOR2_X2 \AES_ENC/us33/U480  ( .A1(\AES_ENC/us33/n1054 ), .A2(\AES_ENC/us33/n1053 ), .ZN(\AES_ENC/us33/n1055 ) );
OR2_X4 \AES_ENC/us33/U479  ( .A1(\AES_ENC/us33/n1094 ), .A2(\AES_ENC/us33/n1093 ), .ZN(\AES_ENC/us33/n571 ) );
AND2_X2 \AES_ENC/us33/U478  ( .A1(\AES_ENC/us33/n571 ), .A2(\AES_ENC/us33/n1095 ), .ZN(\AES_ENC/us33/n1101 ) );
NOR2_X2 \AES_ENC/us33/U477  ( .A1(\AES_ENC/us33/n1074 ), .A2(\AES_ENC/us33/n931 ), .ZN(\AES_ENC/us33/n796 ) );
NOR2_X2 \AES_ENC/us33/U474  ( .A1(\AES_ENC/us33/n796 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n797 ) );
NOR2_X2 \AES_ENC/us33/U473  ( .A1(\AES_ENC/us33/n932 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n933 ) );
NOR2_X2 \AES_ENC/us33/U472  ( .A1(\AES_ENC/us33/n929 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n935 ) );
NOR2_X2 \AES_ENC/us33/U471  ( .A1(\AES_ENC/us33/n931 ), .A2(\AES_ENC/us33/n930 ), .ZN(\AES_ENC/us33/n934 ) );
NOR3_X2 \AES_ENC/us33/U470  ( .A1(\AES_ENC/us33/n935 ), .A2(\AES_ENC/us33/n934 ), .A3(\AES_ENC/us33/n933 ), .ZN(\AES_ENC/us33/n936 ) );
NOR2_X2 \AES_ENC/us33/U469  ( .A1(\AES_ENC/us33/n624 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n1075 ) );
NOR2_X2 \AES_ENC/us33/U468  ( .A1(\AES_ENC/us33/n572 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n949 ) );
NOR2_X2 \AES_ENC/us33/U467  ( .A1(\AES_ENC/us33/n1049 ), .A2(\AES_ENC/us33/n618 ), .ZN(\AES_ENC/us33/n1051 ) );
NOR2_X2 \AES_ENC/us33/U466  ( .A1(\AES_ENC/us33/n1051 ), .A2(\AES_ENC/us33/n1050 ), .ZN(\AES_ENC/us33/n1052 ) );
NOR2_X2 \AES_ENC/us33/U465  ( .A1(\AES_ENC/us33/n1052 ), .A2(\AES_ENC/us33/n592 ), .ZN(\AES_ENC/us33/n1064 ) );
NOR2_X2 \AES_ENC/us33/U464  ( .A1(\AES_ENC/sa33 [1]), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n631 ) );
NOR2_X2 \AES_ENC/us33/U463  ( .A1(\AES_ENC/us33/n1025 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n980 ) );
NOR2_X2 \AES_ENC/us33/U462  ( .A1(\AES_ENC/us33/n1073 ), .A2(\AES_ENC/us33/n1094 ), .ZN(\AES_ENC/us33/n795 ) );
NOR2_X2 \AES_ENC/us33/U461  ( .A1(\AES_ENC/us33/n795 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n799 ) );
NOR2_X2 \AES_ENC/us33/U460  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n981 ) );
NOR2_X2 \AES_ENC/us33/U459  ( .A1(\AES_ENC/us33/n1102 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n643 ) );
NOR2_X2 \AES_ENC/us33/U458  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n621 ), .ZN(\AES_ENC/us33/n642 ) );
NOR2_X2 \AES_ENC/us33/U455  ( .A1(\AES_ENC/us33/n911 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n644 ) );
NOR4_X2 \AES_ENC/us33/U448  ( .A1(\AES_ENC/us33/n644 ), .A2(\AES_ENC/us33/n643 ), .A3(\AES_ENC/us33/n804 ), .A4(\AES_ENC/us33/n642 ), .ZN(\AES_ENC/us33/n645 ) );
NOR2_X2 \AES_ENC/us33/U447  ( .A1(\AES_ENC/us33/n1102 ), .A2(\AES_ENC/us33/n910 ), .ZN(\AES_ENC/us33/n932 ) );
NOR2_X2 \AES_ENC/us33/U442  ( .A1(\AES_ENC/us33/n1102 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n755 ) );
NOR2_X2 \AES_ENC/us33/U441  ( .A1(\AES_ENC/us33/n931 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n743 ) );
NOR2_X2 \AES_ENC/us33/U438  ( .A1(\AES_ENC/us33/n1072 ), .A2(\AES_ENC/us33/n1094 ), .ZN(\AES_ENC/us33/n930 ) );
NOR2_X2 \AES_ENC/us33/U435  ( .A1(\AES_ENC/us33/n1074 ), .A2(\AES_ENC/us33/n1025 ), .ZN(\AES_ENC/us33/n891 ) );
NOR2_X2 \AES_ENC/us33/U434  ( .A1(\AES_ENC/us33/n891 ), .A2(\AES_ENC/us33/n609 ), .ZN(\AES_ENC/us33/n894 ) );
NOR3_X2 \AES_ENC/us33/U433  ( .A1(\AES_ENC/us33/n623 ), .A2(\AES_ENC/sa33 [1]), .A3(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n683 ));
INV_X4 \AES_ENC/us33/U428  ( .A(\AES_ENC/us33/n931 ), .ZN(\AES_ENC/us33/n623 ) );
NOR2_X2 \AES_ENC/us33/U427  ( .A1(\AES_ENC/us33/n996 ), .A2(\AES_ENC/us33/n931 ), .ZN(\AES_ENC/us33/n704 ) );
NOR2_X2 \AES_ENC/us33/U421  ( .A1(\AES_ENC/us33/n931 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n685 ) );
NOR2_X2 \AES_ENC/us33/U420  ( .A1(\AES_ENC/us33/n1029 ), .A2(\AES_ENC/us33/n1025 ), .ZN(\AES_ENC/us33/n1079 ) );
NOR3_X2 \AES_ENC/us33/U419  ( .A1(\AES_ENC/us33/n589 ), .A2(\AES_ENC/us33/n1025 ), .A3(\AES_ENC/us33/n616 ), .ZN(\AES_ENC/us33/n945 ) );
NOR2_X2 \AES_ENC/us33/U418  ( .A1(\AES_ENC/us33/n626 ), .A2(\AES_ENC/us33/n611 ), .ZN(\AES_ENC/us33/n800 ) );
NOR3_X2 \AES_ENC/us33/U417  ( .A1(\AES_ENC/us33/n590 ), .A2(\AES_ENC/us33/n627 ), .A3(\AES_ENC/us33/n611 ), .ZN(\AES_ENC/us33/n798 ) );
NOR3_X2 \AES_ENC/us33/U416  ( .A1(\AES_ENC/us33/n610 ), .A2(\AES_ENC/us33/n572 ), .A3(\AES_ENC/us33/n575 ), .ZN(\AES_ENC/us33/n962 ) );
NOR3_X2 \AES_ENC/us33/U415  ( .A1(\AES_ENC/us33/n959 ), .A2(\AES_ENC/us33/n572 ), .A3(\AES_ENC/us33/n609 ), .ZN(\AES_ENC/us33/n768 ) );
NOR3_X2 \AES_ENC/us33/U414  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n572 ), .A3(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n694 ) );
NOR3_X2 \AES_ENC/us33/U413  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n572 ), .A3(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n895 ) );
NOR3_X2 \AES_ENC/us33/U410  ( .A1(\AES_ENC/us33/n1008 ), .A2(\AES_ENC/us33/n1007 ), .A3(\AES_ENC/us33/n1006 ), .ZN(\AES_ENC/us33/n1018 ) );
NOR4_X2 \AES_ENC/us33/U409  ( .A1(\AES_ENC/us33/n806 ), .A2(\AES_ENC/us33/n805 ), .A3(\AES_ENC/us33/n804 ), .A4(\AES_ENC/us33/n803 ), .ZN(\AES_ENC/us33/n807 ) );
NOR3_X2 \AES_ENC/us33/U406  ( .A1(\AES_ENC/us33/n799 ), .A2(\AES_ENC/us33/n798 ), .A3(\AES_ENC/us33/n797 ), .ZN(\AES_ENC/us33/n808 ) );
NOR4_X2 \AES_ENC/us33/U405  ( .A1(\AES_ENC/us33/n843 ), .A2(\AES_ENC/us33/n842 ), .A3(\AES_ENC/us33/n841 ), .A4(\AES_ENC/us33/n840 ), .ZN(\AES_ENC/us33/n844 ) );
NOR3_X2 \AES_ENC/us33/U404  ( .A1(\AES_ENC/us33/n1101 ), .A2(\AES_ENC/us33/n1100 ), .A3(\AES_ENC/us33/n1099 ), .ZN(\AES_ENC/us33/n1109 ) );
NOR4_X2 \AES_ENC/us33/U403  ( .A1(\AES_ENC/us33/n711 ), .A2(\AES_ENC/us33/n710 ), .A3(\AES_ENC/us33/n709 ), .A4(\AES_ENC/us33/n708 ), .ZN(\AES_ENC/us33/n712 ) );
NOR4_X2 \AES_ENC/us33/U401  ( .A1(\AES_ENC/us33/n963 ), .A2(\AES_ENC/us33/n962 ), .A3(\AES_ENC/us33/n961 ), .A4(\AES_ENC/us33/n960 ), .ZN(\AES_ENC/us33/n964 ) );
NOR2_X2 \AES_ENC/us33/U400  ( .A1(\AES_ENC/us33/n669 ), .A2(\AES_ENC/us33/n668 ), .ZN(\AES_ENC/us33/n673 ) );
NOR4_X2 \AES_ENC/us33/U399  ( .A1(\AES_ENC/us33/n946 ), .A2(\AES_ENC/us33/n1046 ), .A3(\AES_ENC/us33/n671 ), .A4(\AES_ENC/us33/n670 ), .ZN(\AES_ENC/us33/n672 ) );
NOR3_X2 \AES_ENC/us33/U398  ( .A1(\AES_ENC/us33/n743 ), .A2(\AES_ENC/us33/n742 ), .A3(\AES_ENC/us33/n741 ), .ZN(\AES_ENC/us33/n744 ) );
NOR2_X2 \AES_ENC/us33/U397  ( .A1(\AES_ENC/us33/n697 ), .A2(\AES_ENC/us33/n658 ), .ZN(\AES_ENC/us33/n659 ) );
NOR2_X2 \AES_ENC/us33/U396  ( .A1(\AES_ENC/us33/n1078 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n1033 ) );
NOR2_X2 \AES_ENC/us33/U393  ( .A1(\AES_ENC/us33/n1031 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n1032 ) );
NOR3_X2 \AES_ENC/us33/U390  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n1025 ), .A3(\AES_ENC/us33/n1074 ), .ZN(\AES_ENC/us33/n1035 ) );
NOR4_X2 \AES_ENC/us33/U389  ( .A1(\AES_ENC/us33/n1035 ), .A2(\AES_ENC/us33/n1034 ), .A3(\AES_ENC/us33/n1033 ), .A4(\AES_ENC/us33/n1032 ), .ZN(\AES_ENC/us33/n1036 ) );
NOR2_X2 \AES_ENC/us33/U388  ( .A1(\AES_ENC/us33/n598 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n885 ) );
NOR2_X2 \AES_ENC/us33/U387  ( .A1(\AES_ENC/us33/n623 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n882 ) );
NOR2_X2 \AES_ENC/us33/U386  ( .A1(\AES_ENC/us33/n1053 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n884 ) );
NOR4_X2 \AES_ENC/us33/U385  ( .A1(\AES_ENC/us33/n885 ), .A2(\AES_ENC/us33/n884 ), .A3(\AES_ENC/us33/n883 ), .A4(\AES_ENC/us33/n882 ), .ZN(\AES_ENC/us33/n886 ) );
NOR2_X2 \AES_ENC/us33/U384  ( .A1(\AES_ENC/us33/n825 ), .A2(\AES_ENC/us33/n578 ), .ZN(\AES_ENC/us33/n830 ) );
NOR2_X2 \AES_ENC/us33/U383  ( .A1(\AES_ENC/us33/n827 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n829 ) );
NOR2_X2 \AES_ENC/us33/U382  ( .A1(\AES_ENC/us33/n572 ), .A2(\AES_ENC/us33/n579 ), .ZN(\AES_ENC/us33/n828 ) );
NOR4_X2 \AES_ENC/us33/U374  ( .A1(\AES_ENC/us33/n831 ), .A2(\AES_ENC/us33/n830 ), .A3(\AES_ENC/us33/n829 ), .A4(\AES_ENC/us33/n828 ), .ZN(\AES_ENC/us33/n832 ) );
NOR2_X2 \AES_ENC/us33/U373  ( .A1(\AES_ENC/us33/n606 ), .A2(\AES_ENC/us33/n582 ), .ZN(\AES_ENC/us33/n1104 ) );
NOR2_X2 \AES_ENC/us33/U372  ( .A1(\AES_ENC/us33/n1102 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n1106 ) );
NOR2_X2 \AES_ENC/us33/U370  ( .A1(\AES_ENC/us33/n1103 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n1105 ) );
NOR4_X2 \AES_ENC/us33/U369  ( .A1(\AES_ENC/us33/n1107 ), .A2(\AES_ENC/us33/n1106 ), .A3(\AES_ENC/us33/n1105 ), .A4(\AES_ENC/us33/n1104 ), .ZN(\AES_ENC/us33/n1108 ) );
NOR3_X2 \AES_ENC/us33/U368  ( .A1(\AES_ENC/us33/n959 ), .A2(\AES_ENC/us33/n621 ), .A3(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n963 ) );
NOR2_X2 \AES_ENC/us33/U367  ( .A1(\AES_ENC/us33/n626 ), .A2(\AES_ENC/us33/n627 ), .ZN(\AES_ENC/us33/n1114 ) );
INV_X4 \AES_ENC/us33/U366  ( .A(\AES_ENC/us33/n1024 ), .ZN(\AES_ENC/us33/n606 ) );
NOR3_X2 \AES_ENC/us33/U365  ( .A1(\AES_ENC/us33/n910 ), .A2(\AES_ENC/us33/n1059 ), .A3(\AES_ENC/us33/n611 ), .ZN(\AES_ENC/us33/n1115 ) );
INV_X4 \AES_ENC/us33/U364  ( .A(\AES_ENC/us33/n1094 ), .ZN(\AES_ENC/us33/n613 ) );
NOR2_X2 \AES_ENC/us33/U363  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n931 ), .ZN(\AES_ENC/us33/n1100 ) );
INV_X4 \AES_ENC/us33/U354  ( .A(\AES_ENC/us33/n1093 ), .ZN(\AES_ENC/us33/n617 ) );
NOR2_X2 \AES_ENC/us33/U353  ( .A1(\AES_ENC/us33/n569 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n929 ) );
NOR2_X2 \AES_ENC/us33/U352  ( .A1(\AES_ENC/us33/n620 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n926 ) );
NOR2_X2 \AES_ENC/us33/U351  ( .A1(\AES_ENC/us33/n572 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n1095 ) );
NOR2_X2 \AES_ENC/us33/U350  ( .A1(\AES_ENC/us33/n609 ), .A2(\AES_ENC/us33/n627 ), .ZN(\AES_ENC/us33/n1010 ) );
NOR2_X2 \AES_ENC/us33/U349  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n1103 ) );
NOR2_X2 \AES_ENC/us33/U348  ( .A1(\AES_ENC/us33/n622 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n1059 ) );
NOR2_X2 \AES_ENC/us33/U347  ( .A1(\AES_ENC/sa33 [1]), .A2(\AES_ENC/us33/n1120 ), .ZN(\AES_ENC/us33/n1022 ) );
NOR2_X2 \AES_ENC/us33/U346  ( .A1(\AES_ENC/us33/n619 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n911 ) );
NOR2_X2 \AES_ENC/us33/U345  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/us33/n1025 ), .ZN(\AES_ENC/us33/n826 ) );
NOR2_X2 \AES_ENC/us33/U338  ( .A1(\AES_ENC/us33/n626 ), .A2(\AES_ENC/us33/n607 ), .ZN(\AES_ENC/us33/n1072 ) );
NOR2_X2 \AES_ENC/us33/U335  ( .A1(\AES_ENC/us33/n627 ), .A2(\AES_ENC/us33/n616 ), .ZN(\AES_ENC/us33/n956 ) );
NOR2_X2 \AES_ENC/us33/U329  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/us33/n624 ), .ZN(\AES_ENC/us33/n1121 ) );
NOR2_X2 \AES_ENC/us33/U328  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/us33/n624 ), .ZN(\AES_ENC/us33/n1058 ) );
NOR2_X2 \AES_ENC/us33/U327  ( .A1(\AES_ENC/us33/n625 ), .A2(\AES_ENC/us33/n611 ), .ZN(\AES_ENC/us33/n1073 ) );
NOR2_X2 \AES_ENC/us33/U325  ( .A1(\AES_ENC/sa33 [1]), .A2(\AES_ENC/us33/n1025 ), .ZN(\AES_ENC/us33/n1054 ) );
NOR2_X2 \AES_ENC/us33/U324  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/us33/n931 ), .ZN(\AES_ENC/us33/n1029 ) );
NOR2_X2 \AES_ENC/us33/U319  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n1056 ) );
NOR2_X2 \AES_ENC/us33/U318  ( .A1(\AES_ENC/us33/n614 ), .A2(\AES_ENC/us33/n626 ), .ZN(\AES_ENC/us33/n1050 ) );
NOR2_X2 \AES_ENC/us33/U317  ( .A1(\AES_ENC/us33/n1121 ), .A2(\AES_ENC/us33/n1025 ), .ZN(\AES_ENC/us33/n1120 ) );
NOR2_X2 \AES_ENC/us33/U316  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/us33/n572 ), .ZN(\AES_ENC/us33/n1074 ) );
NOR2_X2 \AES_ENC/us33/U315  ( .A1(\AES_ENC/us33/n1058 ), .A2(\AES_ENC/us33/n1054 ), .ZN(\AES_ENC/us33/n878 ) );
NOR2_X2 \AES_ENC/us33/U314  ( .A1(\AES_ENC/us33/n878 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n879 ) );
NOR2_X2 \AES_ENC/us33/U312  ( .A1(\AES_ENC/us33/n880 ), .A2(\AES_ENC/us33/n879 ), .ZN(\AES_ENC/us33/n887 ) );
NOR2_X2 \AES_ENC/us33/U311  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n588 ), .ZN(\AES_ENC/us33/n957 ) );
NOR2_X2 \AES_ENC/us33/U310  ( .A1(\AES_ENC/us33/n958 ), .A2(\AES_ENC/us33/n957 ), .ZN(\AES_ENC/us33/n965 ) );
NOR3_X2 \AES_ENC/us33/U309  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n1091 ), .A3(\AES_ENC/us33/n1022 ), .ZN(\AES_ENC/us33/n720 ) );
NOR3_X2 \AES_ENC/us33/U303  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n1054 ), .A3(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n719 ) );
NOR2_X2 \AES_ENC/us33/U302  ( .A1(\AES_ENC/us33/n720 ), .A2(\AES_ENC/us33/n719 ), .ZN(\AES_ENC/us33/n726 ) );
NOR2_X2 \AES_ENC/us33/U300  ( .A1(\AES_ENC/us33/n614 ), .A2(\AES_ENC/us33/n591 ), .ZN(\AES_ENC/us33/n865 ) );
NOR2_X2 \AES_ENC/us33/U299  ( .A1(\AES_ENC/us33/n1059 ), .A2(\AES_ENC/us33/n1058 ), .ZN(\AES_ENC/us33/n1060 ) );
NOR2_X2 \AES_ENC/us33/U298  ( .A1(\AES_ENC/us33/n1095 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n668 ) );
NOR2_X2 \AES_ENC/us33/U297  ( .A1(\AES_ENC/us33/n911 ), .A2(\AES_ENC/us33/n910 ), .ZN(\AES_ENC/us33/n912 ) );
NOR2_X2 \AES_ENC/us33/U296  ( .A1(\AES_ENC/us33/n912 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n916 ) );
NOR2_X2 \AES_ENC/us33/U295  ( .A1(\AES_ENC/us33/n826 ), .A2(\AES_ENC/us33/n573 ), .ZN(\AES_ENC/us33/n750 ) );
NOR2_X2 \AES_ENC/us33/U294  ( .A1(\AES_ENC/us33/n750 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n751 ) );
NOR2_X2 \AES_ENC/us33/U293  ( .A1(\AES_ENC/us33/n907 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n908 ) );
NOR2_X2 \AES_ENC/us33/U292  ( .A1(\AES_ENC/us33/n990 ), .A2(\AES_ENC/us33/n926 ), .ZN(\AES_ENC/us33/n780 ) );
NOR2_X2 \AES_ENC/us33/U291  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n584 ), .ZN(\AES_ENC/us33/n838 ) );
NOR2_X2 \AES_ENC/us33/U290  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n602 ), .ZN(\AES_ENC/us33/n837 ) );
NOR2_X2 \AES_ENC/us33/U284  ( .A1(\AES_ENC/us33/n838 ), .A2(\AES_ENC/us33/n837 ), .ZN(\AES_ENC/us33/n845 ) );
NOR2_X2 \AES_ENC/us33/U283  ( .A1(\AES_ENC/us33/n1022 ), .A2(\AES_ENC/us33/n1058 ), .ZN(\AES_ENC/us33/n740 ) );
NOR2_X2 \AES_ENC/us33/U282  ( .A1(\AES_ENC/us33/n740 ), .A2(\AES_ENC/us33/n616 ), .ZN(\AES_ENC/us33/n742 ) );
NOR2_X2 \AES_ENC/us33/U281  ( .A1(\AES_ENC/us33/n1098 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n1099 ) );
NOR2_X2 \AES_ENC/us33/U280  ( .A1(\AES_ENC/us33/n1120 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n993 ) );
NOR2_X2 \AES_ENC/us33/U279  ( .A1(\AES_ENC/us33/n993 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n994 ) );
NOR2_X2 \AES_ENC/us33/U273  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n620 ), .ZN(\AES_ENC/us33/n1026 ) );
NOR2_X2 \AES_ENC/us33/U272  ( .A1(\AES_ENC/us33/n573 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n1027 ) );
NOR2_X2 \AES_ENC/us33/U271  ( .A1(\AES_ENC/us33/n1027 ), .A2(\AES_ENC/us33/n1026 ), .ZN(\AES_ENC/us33/n1028 ) );
NOR2_X2 \AES_ENC/us33/U270  ( .A1(\AES_ENC/us33/n1029 ), .A2(\AES_ENC/us33/n1028 ), .ZN(\AES_ENC/us33/n1034 ) );
NOR4_X2 \AES_ENC/us33/U269  ( .A1(\AES_ENC/us33/n757 ), .A2(\AES_ENC/us33/n756 ), .A3(\AES_ENC/us33/n755 ), .A4(\AES_ENC/us33/n754 ), .ZN(\AES_ENC/us33/n758 ) );
NOR2_X2 \AES_ENC/us33/U268  ( .A1(\AES_ENC/us33/n752 ), .A2(\AES_ENC/us33/n751 ), .ZN(\AES_ENC/us33/n759 ) );
NOR2_X2 \AES_ENC/us33/U267  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n1071 ), .ZN(\AES_ENC/us33/n669 ) );
NOR2_X2 \AES_ENC/us33/U263  ( .A1(\AES_ENC/us33/n1056 ), .A2(\AES_ENC/us33/n990 ), .ZN(\AES_ENC/us33/n991 ) );
NOR2_X2 \AES_ENC/us33/U262  ( .A1(\AES_ENC/us33/n991 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n995 ) );
NOR2_X2 \AES_ENC/us33/U258  ( .A1(\AES_ENC/us33/n607 ), .A2(\AES_ENC/us33/n590 ), .ZN(\AES_ENC/us33/n1008 ) );
NOR2_X2 \AES_ENC/us33/U255  ( .A1(\AES_ENC/us33/n839 ), .A2(\AES_ENC/us33/n582 ), .ZN(\AES_ENC/us33/n693 ) );
NOR2_X2 \AES_ENC/us33/U254  ( .A1(\AES_ENC/us33/n606 ), .A2(\AES_ENC/us33/n906 ), .ZN(\AES_ENC/us33/n741 ) );
NOR2_X2 \AES_ENC/us33/U253  ( .A1(\AES_ENC/us33/n1054 ), .A2(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n763 ) );
NOR2_X2 \AES_ENC/us33/U252  ( .A1(\AES_ENC/us33/n763 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n769 ) );
NOR2_X2 \AES_ENC/us33/U251  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n577 ), .ZN(\AES_ENC/us33/n1007 ) );
NOR2_X2 \AES_ENC/us33/U250  ( .A1(\AES_ENC/us33/n609 ), .A2(\AES_ENC/us33/n580 ), .ZN(\AES_ENC/us33/n1123 ) );
NOR2_X2 \AES_ENC/us33/U243  ( .A1(\AES_ENC/us33/n609 ), .A2(\AES_ENC/us33/n590 ), .ZN(\AES_ENC/us33/n710 ) );
INV_X4 \AES_ENC/us33/U242  ( .A(\AES_ENC/us33/n1029 ), .ZN(\AES_ENC/us33/n582 ) );
NOR2_X2 \AES_ENC/us33/U241  ( .A1(\AES_ENC/us33/n616 ), .A2(\AES_ENC/us33/n597 ), .ZN(\AES_ENC/us33/n883 ) );
NOR2_X2 \AES_ENC/us33/U240  ( .A1(\AES_ENC/us33/n593 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n1125 ) );
NOR2_X2 \AES_ENC/us33/U239  ( .A1(\AES_ENC/us33/n990 ), .A2(\AES_ENC/us33/n929 ), .ZN(\AES_ENC/us33/n892 ) );
NOR2_X2 \AES_ENC/us33/U238  ( .A1(\AES_ENC/us33/n892 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n893 ) );
NOR2_X2 \AES_ENC/us33/U237  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n602 ), .ZN(\AES_ENC/us33/n950 ) );
NOR2_X2 \AES_ENC/us33/U236  ( .A1(\AES_ENC/us33/n1079 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n1082 ) );
NOR2_X2 \AES_ENC/us33/U235  ( .A1(\AES_ENC/us33/n910 ), .A2(\AES_ENC/us33/n1056 ), .ZN(\AES_ENC/us33/n941 ) );
NOR2_X2 \AES_ENC/us33/U234  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n1077 ), .ZN(\AES_ENC/us33/n841 ) );
NOR2_X2 \AES_ENC/us33/U229  ( .A1(\AES_ENC/us33/n623 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n630 ) );
NOR2_X2 \AES_ENC/us33/U228  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n602 ), .ZN(\AES_ENC/us33/n806 ) );
NOR2_X2 \AES_ENC/us33/U227  ( .A1(\AES_ENC/us33/n623 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n948 ) );
NOR2_X2 \AES_ENC/us33/U226  ( .A1(\AES_ENC/us33/n606 ), .A2(\AES_ENC/us33/n589 ), .ZN(\AES_ENC/us33/n997 ) );
NOR2_X2 \AES_ENC/us33/U225  ( .A1(\AES_ENC/us33/n1121 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n1122 ) );
NOR2_X2 \AES_ENC/us33/U223  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n1023 ), .ZN(\AES_ENC/us33/n756 ) );
NOR2_X2 \AES_ENC/us33/U222  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n602 ), .ZN(\AES_ENC/us33/n870 ) );
NOR2_X2 \AES_ENC/us33/U221  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n569 ), .ZN(\AES_ENC/us33/n947 ) );
NOR2_X2 \AES_ENC/us33/U217  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n1077 ), .ZN(\AES_ENC/us33/n1084 ) );
NOR2_X2 \AES_ENC/us33/U213  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n855 ), .ZN(\AES_ENC/us33/n709 ) );
NOR2_X2 \AES_ENC/us33/U212  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n589 ), .ZN(\AES_ENC/us33/n868 ) );
NOR2_X2 \AES_ENC/us33/U211  ( .A1(\AES_ENC/us33/n1120 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n1124 ) );
NOR2_X2 \AES_ENC/us33/U210  ( .A1(\AES_ENC/us33/n1120 ), .A2(\AES_ENC/us33/n839 ), .ZN(\AES_ENC/us33/n842 ) );
NOR2_X2 \AES_ENC/us33/U209  ( .A1(\AES_ENC/us33/n1120 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n696 ) );
NOR2_X2 \AES_ENC/us33/U208  ( .A1(\AES_ENC/us33/n1074 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n1076 ) );
NOR2_X2 \AES_ENC/us33/U207  ( .A1(\AES_ENC/us33/n1074 ), .A2(\AES_ENC/us33/n620 ), .ZN(\AES_ENC/us33/n781 ) );
NOR3_X2 \AES_ENC/us33/U201  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n1056 ), .A3(\AES_ENC/us33/n990 ), .ZN(\AES_ENC/us33/n979 ) );
NOR3_X2 \AES_ENC/us33/U200  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n1058 ), .A3(\AES_ENC/us33/n1059 ), .ZN(\AES_ENC/us33/n854 ) );
NOR2_X2 \AES_ENC/us33/U199  ( .A1(\AES_ENC/us33/n996 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n869 ) );
NOR2_X2 \AES_ENC/us33/U198  ( .A1(\AES_ENC/us33/n1056 ), .A2(\AES_ENC/us33/n1074 ), .ZN(\AES_ENC/us33/n1057 ) );
NOR3_X2 \AES_ENC/us33/U197  ( .A1(\AES_ENC/us33/n607 ), .A2(\AES_ENC/us33/n1120 ), .A3(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n978 ) );
NOR2_X2 \AES_ENC/us33/U196  ( .A1(\AES_ENC/us33/n996 ), .A2(\AES_ENC/us33/n911 ), .ZN(\AES_ENC/us33/n1116 ) );
NOR2_X2 \AES_ENC/us33/U195  ( .A1(\AES_ENC/us33/n1074 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n754 ) );
NOR2_X2 \AES_ENC/us33/U194  ( .A1(\AES_ENC/us33/n926 ), .A2(\AES_ENC/us33/n1103 ), .ZN(\AES_ENC/us33/n977 ) );
NOR2_X2 \AES_ENC/us33/U187  ( .A1(\AES_ENC/us33/n839 ), .A2(\AES_ENC/us33/n824 ), .ZN(\AES_ENC/us33/n1092 ) );
NOR2_X2 \AES_ENC/us33/U186  ( .A1(\AES_ENC/us33/n573 ), .A2(\AES_ENC/us33/n1074 ), .ZN(\AES_ENC/us33/n684 ) );
NOR2_X2 \AES_ENC/us33/U185  ( .A1(\AES_ENC/us33/n826 ), .A2(\AES_ENC/us33/n1059 ), .ZN(\AES_ENC/us33/n907 ) );
NOR3_X2 \AES_ENC/us33/U184  ( .A1(\AES_ENC/us33/n625 ), .A2(\AES_ENC/us33/n1115 ), .A3(\AES_ENC/us33/n585 ), .ZN(\AES_ENC/us33/n831 ) );
NOR3_X2 \AES_ENC/us33/U183  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n1056 ), .A3(\AES_ENC/us33/n990 ), .ZN(\AES_ENC/us33/n896 ) );
NOR3_X2 \AES_ENC/us33/U182  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n573 ), .A3(\AES_ENC/us33/n1013 ), .ZN(\AES_ENC/us33/n670 ) );
NOR3_X2 \AES_ENC/us33/U181  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n1091 ), .A3(\AES_ENC/us33/n1022 ), .ZN(\AES_ENC/us33/n843 ) );
NOR2_X2 \AES_ENC/us33/U180  ( .A1(\AES_ENC/us33/n1029 ), .A2(\AES_ENC/us33/n1095 ), .ZN(\AES_ENC/us33/n735 ) );
NOR2_X2 \AES_ENC/us33/U174  ( .A1(\AES_ENC/us33/n1100 ), .A2(\AES_ENC/us33/n854 ), .ZN(\AES_ENC/us33/n860 ) );
NOR4_X2 \AES_ENC/us33/U173  ( .A1(\AES_ENC/us33/n1125 ), .A2(\AES_ENC/us33/n1124 ), .A3(\AES_ENC/us33/n1123 ), .A4(\AES_ENC/us33/n1122 ), .ZN(\AES_ENC/us33/n1126 ) );
NOR4_X2 \AES_ENC/us33/U172  ( .A1(\AES_ENC/us33/n1084 ), .A2(\AES_ENC/us33/n1083 ), .A3(\AES_ENC/us33/n1082 ), .A4(\AES_ENC/us33/n1081 ), .ZN(\AES_ENC/us33/n1085 ) );
NOR2_X2 \AES_ENC/us33/U171  ( .A1(\AES_ENC/us33/n1076 ), .A2(\AES_ENC/us33/n1075 ), .ZN(\AES_ENC/us33/n1086 ) );
NAND3_X2 \AES_ENC/us33/U170  ( .A1(\AES_ENC/us33/n569 ), .A2(\AES_ENC/us33/n582 ), .A3(\AES_ENC/us33/n681 ), .ZN(\AES_ENC/us33/n691 ) );
NOR2_X2 \AES_ENC/us33/U169  ( .A1(\AES_ENC/us33/n683 ), .A2(\AES_ENC/us33/n682 ), .ZN(\AES_ENC/us33/n690 ) );
NOR3_X2 \AES_ENC/us33/U168  ( .A1(\AES_ENC/us33/n695 ), .A2(\AES_ENC/us33/n694 ), .A3(\AES_ENC/us33/n693 ), .ZN(\AES_ENC/us33/n700 ) );
NOR4_X2 \AES_ENC/us33/U162  ( .A1(\AES_ENC/us33/n983 ), .A2(\AES_ENC/us33/n698 ), .A3(\AES_ENC/us33/n697 ), .A4(\AES_ENC/us33/n696 ), .ZN(\AES_ENC/us33/n699 ) );
NOR2_X2 \AES_ENC/us33/U161  ( .A1(\AES_ENC/us33/n946 ), .A2(\AES_ENC/us33/n945 ), .ZN(\AES_ENC/us33/n952 ) );
NOR4_X2 \AES_ENC/us33/U160  ( .A1(\AES_ENC/us33/n950 ), .A2(\AES_ENC/us33/n949 ), .A3(\AES_ENC/us33/n948 ), .A4(\AES_ENC/us33/n947 ), .ZN(\AES_ENC/us33/n951 ) );
NOR4_X2 \AES_ENC/us33/U159  ( .A1(\AES_ENC/us33/n983 ), .A2(\AES_ENC/us33/n982 ), .A3(\AES_ENC/us33/n981 ), .A4(\AES_ENC/us33/n980 ), .ZN(\AES_ENC/us33/n984 ) );
NOR2_X2 \AES_ENC/us33/U158  ( .A1(\AES_ENC/us33/n979 ), .A2(\AES_ENC/us33/n978 ), .ZN(\AES_ENC/us33/n985 ) );
NOR4_X2 \AES_ENC/us33/U157  ( .A1(\AES_ENC/us33/n896 ), .A2(\AES_ENC/us33/n895 ), .A3(\AES_ENC/us33/n894 ), .A4(\AES_ENC/us33/n893 ), .ZN(\AES_ENC/us33/n897 ) );
NOR2_X2 \AES_ENC/us33/U156  ( .A1(\AES_ENC/us33/n866 ), .A2(\AES_ENC/us33/n865 ), .ZN(\AES_ENC/us33/n872 ) );
NOR4_X2 \AES_ENC/us33/U155  ( .A1(\AES_ENC/us33/n870 ), .A2(\AES_ENC/us33/n869 ), .A3(\AES_ENC/us33/n868 ), .A4(\AES_ENC/us33/n867 ), .ZN(\AES_ENC/us33/n871 ) );
NOR3_X2 \AES_ENC/us33/U154  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n1054 ), .A3(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n961 ) );
NOR3_X2 \AES_ENC/us33/U153  ( .A1(\AES_ENC/us33/n620 ), .A2(\AES_ENC/us33/n1074 ), .A3(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n671 ) );
NOR2_X2 \AES_ENC/us33/U152  ( .A1(\AES_ENC/us33/n1057 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n1062 ) );
NOR2_X2 \AES_ENC/us33/U143  ( .A1(\AES_ENC/us33/n1055 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n1063 ) );
NOR2_X2 \AES_ENC/us33/U142  ( .A1(\AES_ENC/us33/n1060 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n1061 ) );
NOR4_X2 \AES_ENC/us33/U141  ( .A1(\AES_ENC/us33/n1064 ), .A2(\AES_ENC/us33/n1063 ), .A3(\AES_ENC/us33/n1062 ), .A4(\AES_ENC/us33/n1061 ), .ZN(\AES_ENC/us33/n1065 ) );
NOR3_X2 \AES_ENC/us33/U140  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n1120 ), .A3(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n918 ) );
NOR3_X2 \AES_ENC/us33/U132  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n573 ), .A3(\AES_ENC/us33/n1013 ), .ZN(\AES_ENC/us33/n917 ) );
NOR2_X2 \AES_ENC/us33/U131  ( .A1(\AES_ENC/us33/n914 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n915 ) );
NOR4_X2 \AES_ENC/us33/U130  ( .A1(\AES_ENC/us33/n918 ), .A2(\AES_ENC/us33/n917 ), .A3(\AES_ENC/us33/n916 ), .A4(\AES_ENC/us33/n915 ), .ZN(\AES_ENC/us33/n919 ) );
NOR2_X2 \AES_ENC/us33/U129  ( .A1(\AES_ENC/us33/n735 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n687 ) );
NOR2_X2 \AES_ENC/us33/U128  ( .A1(\AES_ENC/us33/n684 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n688 ) );
NOR2_X2 \AES_ENC/us33/U127  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n600 ), .ZN(\AES_ENC/us33/n686 ) );
NOR4_X2 \AES_ENC/us33/U126  ( .A1(\AES_ENC/us33/n688 ), .A2(\AES_ENC/us33/n687 ), .A3(\AES_ENC/us33/n686 ), .A4(\AES_ENC/us33/n685 ), .ZN(\AES_ENC/us33/n689 ) );
NOR2_X2 \AES_ENC/us33/U121  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n595 ), .ZN(\AES_ENC/us33/n858 ) );
NOR2_X2 \AES_ENC/us33/U120  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n855 ), .ZN(\AES_ENC/us33/n857 ) );
NOR2_X2 \AES_ENC/us33/U119  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n587 ), .ZN(\AES_ENC/us33/n856 ) );
NOR4_X2 \AES_ENC/us33/U118  ( .A1(\AES_ENC/us33/n858 ), .A2(\AES_ENC/us33/n857 ), .A3(\AES_ENC/us33/n856 ), .A4(\AES_ENC/us33/n958 ), .ZN(\AES_ENC/us33/n859 ) );
NOR2_X2 \AES_ENC/us33/U117  ( .A1(\AES_ENC/us33/n616 ), .A2(\AES_ENC/us33/n580 ), .ZN(\AES_ENC/us33/n771 ) );
NOR2_X2 \AES_ENC/us33/U116  ( .A1(\AES_ENC/us33/n1103 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n772 ) );
NOR2_X2 \AES_ENC/us33/U115  ( .A1(\AES_ENC/us33/n610 ), .A2(\AES_ENC/us33/n599 ), .ZN(\AES_ENC/us33/n773 ) );
NOR4_X2 \AES_ENC/us33/U106  ( .A1(\AES_ENC/us33/n773 ), .A2(\AES_ENC/us33/n772 ), .A3(\AES_ENC/us33/n771 ), .A4(\AES_ENC/us33/n770 ), .ZN(\AES_ENC/us33/n774 ) );
NOR2_X2 \AES_ENC/us33/U105  ( .A1(\AES_ENC/us33/n780 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n784 ) );
NOR2_X2 \AES_ENC/us33/U104  ( .A1(\AES_ENC/us33/n1117 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n782 ) );
NOR2_X2 \AES_ENC/us33/U103  ( .A1(\AES_ENC/us33/n781 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n783 ) );
NOR4_X2 \AES_ENC/us33/U102  ( .A1(\AES_ENC/us33/n880 ), .A2(\AES_ENC/us33/n784 ), .A3(\AES_ENC/us33/n783 ), .A4(\AES_ENC/us33/n782 ), .ZN(\AES_ENC/us33/n785 ) );
NOR2_X2 \AES_ENC/us33/U101  ( .A1(\AES_ENC/us33/n583 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n814 ) );
NOR2_X2 \AES_ENC/us33/U100  ( .A1(\AES_ENC/us33/n907 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n813 ) );
NOR3_X2 \AES_ENC/us33/U95  ( .A1(\AES_ENC/us33/n606 ), .A2(\AES_ENC/us33/n1058 ), .A3(\AES_ENC/us33/n1059 ), .ZN(\AES_ENC/us33/n815 ) );
NOR4_X2 \AES_ENC/us33/U94  ( .A1(\AES_ENC/us33/n815 ), .A2(\AES_ENC/us33/n814 ), .A3(\AES_ENC/us33/n813 ), .A4(\AES_ENC/us33/n812 ), .ZN(\AES_ENC/us33/n816 ) );
NOR2_X2 \AES_ENC/us33/U93  ( .A1(\AES_ENC/us33/n617 ), .A2(\AES_ENC/us33/n569 ), .ZN(\AES_ENC/us33/n721 ) );
NOR2_X2 \AES_ENC/us33/U92  ( .A1(\AES_ENC/us33/n1031 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n723 ) );
NOR2_X2 \AES_ENC/us33/U91  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n1096 ), .ZN(\AES_ENC/us33/n722 ) );
NOR4_X2 \AES_ENC/us33/U90  ( .A1(\AES_ENC/us33/n724 ), .A2(\AES_ENC/us33/n723 ), .A3(\AES_ENC/us33/n722 ), .A4(\AES_ENC/us33/n721 ), .ZN(\AES_ENC/us33/n725 ) );
NOR2_X2 \AES_ENC/us33/U89  ( .A1(\AES_ENC/us33/n911 ), .A2(\AES_ENC/us33/n990 ), .ZN(\AES_ENC/us33/n1009 ) );
NOR2_X2 \AES_ENC/us33/U88  ( .A1(\AES_ENC/us33/n1013 ), .A2(\AES_ENC/us33/n573 ), .ZN(\AES_ENC/us33/n1014 ) );
NOR2_X2 \AES_ENC/us33/U87  ( .A1(\AES_ENC/us33/n1014 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n1015 ) );
NOR4_X2 \AES_ENC/us33/U86  ( .A1(\AES_ENC/us33/n1016 ), .A2(\AES_ENC/us33/n1015 ), .A3(\AES_ENC/us33/n1119 ), .A4(\AES_ENC/us33/n1046 ), .ZN(\AES_ENC/us33/n1017 ) );
NOR2_X2 \AES_ENC/us33/U81  ( .A1(\AES_ENC/us33/n996 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n998 ) );
NOR2_X2 \AES_ENC/us33/U80  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n577 ), .ZN(\AES_ENC/us33/n1000 ) );
NOR2_X2 \AES_ENC/us33/U79  ( .A1(\AES_ENC/us33/n616 ), .A2(\AES_ENC/us33/n1096 ), .ZN(\AES_ENC/us33/n999 ) );
NOR4_X2 \AES_ENC/us33/U78  ( .A1(\AES_ENC/us33/n1000 ), .A2(\AES_ENC/us33/n999 ), .A3(\AES_ENC/us33/n998 ), .A4(\AES_ENC/us33/n997 ), .ZN(\AES_ENC/us33/n1001 ) );
NOR2_X2 \AES_ENC/us33/U74  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n1096 ), .ZN(\AES_ENC/us33/n697 ) );
NOR2_X2 \AES_ENC/us33/U73  ( .A1(\AES_ENC/us33/n620 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n958 ) );
NOR2_X2 \AES_ENC/us33/U72  ( .A1(\AES_ENC/us33/n911 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n983 ) );
NOR2_X2 \AES_ENC/us33/U71  ( .A1(\AES_ENC/us33/n1054 ), .A2(\AES_ENC/us33/n1103 ), .ZN(\AES_ENC/us33/n1031 ) );
INV_X4 \AES_ENC/us33/U65  ( .A(\AES_ENC/us33/n1050 ), .ZN(\AES_ENC/us33/n612 ) );
INV_X4 \AES_ENC/us33/U64  ( .A(\AES_ENC/us33/n1072 ), .ZN(\AES_ENC/us33/n605 ) );
INV_X4 \AES_ENC/us33/U63  ( .A(\AES_ENC/us33/n1073 ), .ZN(\AES_ENC/us33/n604 ) );
NOR2_X2 \AES_ENC/us33/U62  ( .A1(\AES_ENC/us33/n582 ), .A2(\AES_ENC/us33/n613 ), .ZN(\AES_ENC/us33/n880 ) );
NOR3_X2 \AES_ENC/us33/U61  ( .A1(\AES_ENC/us33/n826 ), .A2(\AES_ENC/us33/n1121 ), .A3(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n946 ) );
INV_X4 \AES_ENC/us33/U59  ( .A(\AES_ENC/us33/n1010 ), .ZN(\AES_ENC/us33/n608 ) );
NOR3_X2 \AES_ENC/us33/U58  ( .A1(\AES_ENC/us33/n573 ), .A2(\AES_ENC/us33/n1029 ), .A3(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n1119 ) );
INV_X4 \AES_ENC/us33/U57  ( .A(\AES_ENC/us33/n956 ), .ZN(\AES_ENC/us33/n615 ) );
NOR2_X2 \AES_ENC/us33/U50  ( .A1(\AES_ENC/us33/n623 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n1013 ) );
NOR2_X2 \AES_ENC/us33/U49  ( .A1(\AES_ENC/us33/n620 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n910 ) );
NOR2_X2 \AES_ENC/us33/U48  ( .A1(\AES_ENC/us33/n569 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n1091 ) );
NOR2_X2 \AES_ENC/us33/U47  ( .A1(\AES_ENC/us33/n622 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n990 ) );
NOR2_X2 \AES_ENC/us33/U46  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/us33/n1121 ), .ZN(\AES_ENC/us33/n996 ) );
NOR2_X2 \AES_ENC/us33/U45  ( .A1(\AES_ENC/us33/n610 ), .A2(\AES_ENC/us33/n600 ), .ZN(\AES_ENC/us33/n628 ) );
NOR2_X2 \AES_ENC/us33/U44  ( .A1(\AES_ENC/us33/n576 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n866 ) );
NOR2_X2 \AES_ENC/us33/U43  ( .A1(\AES_ENC/us33/n603 ), .A2(\AES_ENC/us33/n610 ), .ZN(\AES_ENC/us33/n1006 ) );
NOR2_X2 \AES_ENC/us33/U42  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n1117 ), .ZN(\AES_ENC/us33/n1118 ) );
NOR2_X2 \AES_ENC/us33/U41  ( .A1(\AES_ENC/us33/n1119 ), .A2(\AES_ENC/us33/n1118 ), .ZN(\AES_ENC/us33/n1127 ) );
NOR2_X2 \AES_ENC/us33/U36  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n906 ), .ZN(\AES_ENC/us33/n909 ) );
NOR2_X2 \AES_ENC/us33/U35  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n594 ), .ZN(\AES_ENC/us33/n629 ) );
NOR2_X2 \AES_ENC/us33/U34  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n597 ), .ZN(\AES_ENC/us33/n658 ) );
NOR2_X2 \AES_ENC/us33/U33  ( .A1(\AES_ENC/us33/n1116 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n695 ) );
NOR2_X2 \AES_ENC/us33/U32  ( .A1(\AES_ENC/us33/n1078 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n1083 ) );
NOR2_X2 \AES_ENC/us33/U31  ( .A1(\AES_ENC/us33/n941 ), .A2(\AES_ENC/us33/n608 ), .ZN(\AES_ENC/us33/n724 ) );
NOR2_X2 \AES_ENC/us33/U30  ( .A1(\AES_ENC/us33/n598 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n1107 ) );
NOR2_X2 \AES_ENC/us33/U29  ( .A1(\AES_ENC/us33/n576 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n840 ) );
NOR2_X2 \AES_ENC/us33/U24  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n593 ), .ZN(\AES_ENC/us33/n633 ) );
NOR2_X2 \AES_ENC/us33/U23  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n1080 ), .ZN(\AES_ENC/us33/n1081 ) );
NOR2_X2 \AES_ENC/us33/U21  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n1045 ), .ZN(\AES_ENC/us33/n812 ) );
NOR2_X2 \AES_ENC/us33/U20  ( .A1(\AES_ENC/us33/n1009 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n960 ) );
NOR2_X2 \AES_ENC/us33/U19  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n601 ), .ZN(\AES_ENC/us33/n982 ) );
NOR2_X2 \AES_ENC/us33/U18  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n594 ), .ZN(\AES_ENC/us33/n757 ) );
NOR2_X2 \AES_ENC/us33/U17  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n590 ), .ZN(\AES_ENC/us33/n698 ) );
NOR2_X2 \AES_ENC/us33/U16  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n619 ), .ZN(\AES_ENC/us33/n708 ) );
NOR2_X2 \AES_ENC/us33/U15  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n582 ), .ZN(\AES_ENC/us33/n770 ) );
NOR2_X2 \AES_ENC/us33/U10  ( .A1(\AES_ENC/us33/n619 ), .A2(\AES_ENC/us33/n604 ), .ZN(\AES_ENC/us33/n803 ) );
NOR2_X2 \AES_ENC/us33/U9  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n881 ), .ZN(\AES_ENC/us33/n711 ) );
NOR2_X2 \AES_ENC/us33/U8  ( .A1(\AES_ENC/us33/n615 ), .A2(\AES_ENC/us33/n582 ), .ZN(\AES_ENC/us33/n867 ) );
NOR2_X2 \AES_ENC/us33/U7  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n599 ), .ZN(\AES_ENC/us33/n804 ) );
NOR2_X2 \AES_ENC/us33/U6  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n620 ), .ZN(\AES_ENC/us33/n1046 ) );
OR2_X4 \AES_ENC/us33/U5  ( .A1(\AES_ENC/us33/n624 ), .A2(\AES_ENC/sa33 [1]),.ZN(\AES_ENC/us33/n570 ) );
OR2_X4 \AES_ENC/us33/U4  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/sa33 [4]),.ZN(\AES_ENC/us33/n569 ) );
NAND2_X2 \AES_ENC/us33/U514  ( .A1(\AES_ENC/us33/n1121 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n1030 ) );
AND2_X2 \AES_ENC/us33/U513  ( .A1(\AES_ENC/us33/n597 ), .A2(\AES_ENC/us33/n1030 ), .ZN(\AES_ENC/us33/n1049 ) );
NAND2_X2 \AES_ENC/us33/U511  ( .A1(\AES_ENC/us33/n1049 ), .A2(\AES_ENC/us33/n794 ), .ZN(\AES_ENC/us33/n637 ) );
AND2_X2 \AES_ENC/us33/U493  ( .A1(\AES_ENC/us33/n779 ), .A2(\AES_ENC/us33/n996 ), .ZN(\AES_ENC/us33/n632 ) );
NAND4_X2 \AES_ENC/us33/U485  ( .A1(\AES_ENC/us33/n637 ), .A2(\AES_ENC/us33/n636 ), .A3(\AES_ENC/us33/n635 ), .A4(\AES_ENC/us33/n634 ), .ZN(\AES_ENC/us33/n638 ) );
NAND2_X2 \AES_ENC/us33/U484  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n638 ), .ZN(\AES_ENC/us33/n679 ) );
NAND2_X2 \AES_ENC/us33/U481  ( .A1(\AES_ENC/us33/n1094 ), .A2(\AES_ENC/us33/n591 ), .ZN(\AES_ENC/us33/n648 ) );
NAND2_X2 \AES_ENC/us33/U476  ( .A1(\AES_ENC/us33/n601 ), .A2(\AES_ENC/us33/n590 ), .ZN(\AES_ENC/us33/n762 ) );
NAND2_X2 \AES_ENC/us33/U475  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n762 ), .ZN(\AES_ENC/us33/n647 ) );
NAND4_X2 \AES_ENC/us33/U457  ( .A1(\AES_ENC/us33/n648 ), .A2(\AES_ENC/us33/n647 ), .A3(\AES_ENC/us33/n646 ), .A4(\AES_ENC/us33/n645 ), .ZN(\AES_ENC/us33/n649 ) );
NAND2_X2 \AES_ENC/us33/U456  ( .A1(\AES_ENC/sa33 [0]), .A2(\AES_ENC/us33/n649 ), .ZN(\AES_ENC/us33/n665 ) );
NAND2_X2 \AES_ENC/us33/U454  ( .A1(\AES_ENC/us33/n596 ), .A2(\AES_ENC/us33/n623 ), .ZN(\AES_ENC/us33/n855 ) );
NAND2_X2 \AES_ENC/us33/U453  ( .A1(\AES_ENC/us33/n587 ), .A2(\AES_ENC/us33/n855 ), .ZN(\AES_ENC/us33/n821 ) );
NAND2_X2 \AES_ENC/us33/U452  ( .A1(\AES_ENC/us33/n1093 ), .A2(\AES_ENC/us33/n821 ), .ZN(\AES_ENC/us33/n662 ) );
NAND2_X2 \AES_ENC/us33/U451  ( .A1(\AES_ENC/us33/n619 ), .A2(\AES_ENC/us33/n589 ), .ZN(\AES_ENC/us33/n650 ) );
NAND2_X2 \AES_ENC/us33/U450  ( .A1(\AES_ENC/us33/n956 ), .A2(\AES_ENC/us33/n650 ), .ZN(\AES_ENC/us33/n661 ) );
NAND2_X2 \AES_ENC/us33/U449  ( .A1(\AES_ENC/us33/n626 ), .A2(\AES_ENC/us33/n627 ), .ZN(\AES_ENC/us33/n839 ) );
OR2_X2 \AES_ENC/us33/U446  ( .A1(\AES_ENC/us33/n839 ), .A2(\AES_ENC/us33/n932 ), .ZN(\AES_ENC/us33/n656 ) );
NAND2_X2 \AES_ENC/us33/U445  ( .A1(\AES_ENC/us33/n621 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n1096 ) );
NAND2_X2 \AES_ENC/us33/U444  ( .A1(\AES_ENC/us33/n1030 ), .A2(\AES_ENC/us33/n1096 ), .ZN(\AES_ENC/us33/n651 ) );
NAND2_X2 \AES_ENC/us33/U443  ( .A1(\AES_ENC/us33/n1114 ), .A2(\AES_ENC/us33/n651 ), .ZN(\AES_ENC/us33/n655 ) );
OR3_X2 \AES_ENC/us33/U440  ( .A1(\AES_ENC/us33/n1079 ), .A2(\AES_ENC/sa33 [7]), .A3(\AES_ENC/us33/n626 ), .ZN(\AES_ENC/us33/n654 ));
NAND2_X2 \AES_ENC/us33/U439  ( .A1(\AES_ENC/us33/n593 ), .A2(\AES_ENC/us33/n601 ), .ZN(\AES_ENC/us33/n652 ) );
NAND4_X2 \AES_ENC/us33/U437  ( .A1(\AES_ENC/us33/n656 ), .A2(\AES_ENC/us33/n655 ), .A3(\AES_ENC/us33/n654 ), .A4(\AES_ENC/us33/n653 ), .ZN(\AES_ENC/us33/n657 ) );
NAND2_X2 \AES_ENC/us33/U436  ( .A1(\AES_ENC/sa33 [2]), .A2(\AES_ENC/us33/n657 ), .ZN(\AES_ENC/us33/n660 ) );
NAND4_X2 \AES_ENC/us33/U432  ( .A1(\AES_ENC/us33/n662 ), .A2(\AES_ENC/us33/n661 ), .A3(\AES_ENC/us33/n660 ), .A4(\AES_ENC/us33/n659 ), .ZN(\AES_ENC/us33/n663 ) );
NAND2_X2 \AES_ENC/us33/U431  ( .A1(\AES_ENC/us33/n663 ), .A2(\AES_ENC/us33/n574 ), .ZN(\AES_ENC/us33/n664 ) );
NAND2_X2 \AES_ENC/us33/U430  ( .A1(\AES_ENC/us33/n665 ), .A2(\AES_ENC/us33/n664 ), .ZN(\AES_ENC/us33/n666 ) );
NAND2_X2 \AES_ENC/us33/U429  ( .A1(\AES_ENC/sa33 [6]), .A2(\AES_ENC/us33/n666 ), .ZN(\AES_ENC/us33/n678 ) );
NAND2_X2 \AES_ENC/us33/U426  ( .A1(\AES_ENC/us33/n735 ), .A2(\AES_ENC/us33/n1093 ), .ZN(\AES_ENC/us33/n675 ) );
NAND2_X2 \AES_ENC/us33/U425  ( .A1(\AES_ENC/us33/n588 ), .A2(\AES_ENC/us33/n597 ), .ZN(\AES_ENC/us33/n1045 ) );
OR2_X2 \AES_ENC/us33/U424  ( .A1(\AES_ENC/us33/n1045 ), .A2(\AES_ENC/us33/n605 ), .ZN(\AES_ENC/us33/n674 ) );
NAND2_X2 \AES_ENC/us33/U423  ( .A1(\AES_ENC/sa33 [1]), .A2(\AES_ENC/us33/n620 ), .ZN(\AES_ENC/us33/n667 ) );
NAND2_X2 \AES_ENC/us33/U422  ( .A1(\AES_ENC/us33/n619 ), .A2(\AES_ENC/us33/n667 ), .ZN(\AES_ENC/us33/n1071 ) );
NAND4_X2 \AES_ENC/us33/U412  ( .A1(\AES_ENC/us33/n675 ), .A2(\AES_ENC/us33/n674 ), .A3(\AES_ENC/us33/n673 ), .A4(\AES_ENC/us33/n672 ), .ZN(\AES_ENC/us33/n676 ) );
NAND2_X2 \AES_ENC/us33/U411  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n676 ), .ZN(\AES_ENC/us33/n677 ) );
NAND2_X2 \AES_ENC/us33/U408  ( .A1(\AES_ENC/us33/n800 ), .A2(\AES_ENC/us33/n1022 ), .ZN(\AES_ENC/us33/n680 ) );
NAND2_X2 \AES_ENC/us33/U407  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n680 ), .ZN(\AES_ENC/us33/n681 ) );
AND2_X2 \AES_ENC/us33/U402  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n684 ), .ZN(\AES_ENC/us33/n682 ) );
NAND4_X2 \AES_ENC/us33/U395  ( .A1(\AES_ENC/us33/n691 ), .A2(\AES_ENC/us33/n581 ), .A3(\AES_ENC/us33/n690 ), .A4(\AES_ENC/us33/n689 ), .ZN(\AES_ENC/us33/n692 ) );
NAND2_X2 \AES_ENC/us33/U394  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n692 ), .ZN(\AES_ENC/us33/n733 ) );
NAND2_X2 \AES_ENC/us33/U392  ( .A1(\AES_ENC/us33/n977 ), .A2(\AES_ENC/us33/n1050 ), .ZN(\AES_ENC/us33/n702 ) );
NAND2_X2 \AES_ENC/us33/U391  ( .A1(\AES_ENC/us33/n1093 ), .A2(\AES_ENC/us33/n1045 ), .ZN(\AES_ENC/us33/n701 ) );
NAND4_X2 \AES_ENC/us33/U381  ( .A1(\AES_ENC/us33/n702 ), .A2(\AES_ENC/us33/n701 ), .A3(\AES_ENC/us33/n700 ), .A4(\AES_ENC/us33/n699 ), .ZN(\AES_ENC/us33/n703 ) );
NAND2_X2 \AES_ENC/us33/U380  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n703 ), .ZN(\AES_ENC/us33/n732 ) );
AND2_X2 \AES_ENC/us33/U379  ( .A1(\AES_ENC/sa33 [0]), .A2(\AES_ENC/sa33 [6]),.ZN(\AES_ENC/us33/n1113 ) );
NAND2_X2 \AES_ENC/us33/U378  ( .A1(\AES_ENC/us33/n601 ), .A2(\AES_ENC/us33/n1030 ), .ZN(\AES_ENC/us33/n881 ) );
NAND2_X2 \AES_ENC/us33/U377  ( .A1(\AES_ENC/us33/n1093 ), .A2(\AES_ENC/us33/n881 ), .ZN(\AES_ENC/us33/n715 ) );
NAND2_X2 \AES_ENC/us33/U376  ( .A1(\AES_ENC/us33/n1010 ), .A2(\AES_ENC/us33/n600 ), .ZN(\AES_ENC/us33/n714 ) );
NAND2_X2 \AES_ENC/us33/U375  ( .A1(\AES_ENC/us33/n855 ), .A2(\AES_ENC/us33/n588 ), .ZN(\AES_ENC/us33/n1117 ) );
XNOR2_X2 \AES_ENC/us33/U371  ( .A(\AES_ENC/us33/n611 ), .B(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n824 ) );
NAND4_X2 \AES_ENC/us33/U362  ( .A1(\AES_ENC/us33/n715 ), .A2(\AES_ENC/us33/n714 ), .A3(\AES_ENC/us33/n713 ), .A4(\AES_ENC/us33/n712 ), .ZN(\AES_ENC/us33/n716 ) );
NAND2_X2 \AES_ENC/us33/U361  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n716 ), .ZN(\AES_ENC/us33/n731 ) );
AND2_X2 \AES_ENC/us33/U360  ( .A1(\AES_ENC/sa33 [6]), .A2(\AES_ENC/us33/n574 ), .ZN(\AES_ENC/us33/n1131 ) );
NAND2_X2 \AES_ENC/us33/U359  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n717 ) );
NAND2_X2 \AES_ENC/us33/U358  ( .A1(\AES_ENC/us33/n1029 ), .A2(\AES_ENC/us33/n717 ), .ZN(\AES_ENC/us33/n728 ) );
NAND2_X2 \AES_ENC/us33/U357  ( .A1(\AES_ENC/sa33 [1]), .A2(\AES_ENC/us33/n624 ), .ZN(\AES_ENC/us33/n1097 ) );
NAND2_X2 \AES_ENC/us33/U356  ( .A1(\AES_ENC/us33/n603 ), .A2(\AES_ENC/us33/n1097 ), .ZN(\AES_ENC/us33/n718 ) );
NAND2_X2 \AES_ENC/us33/U355  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n718 ), .ZN(\AES_ENC/us33/n727 ) );
NAND4_X2 \AES_ENC/us33/U344  ( .A1(\AES_ENC/us33/n728 ), .A2(\AES_ENC/us33/n727 ), .A3(\AES_ENC/us33/n726 ), .A4(\AES_ENC/us33/n725 ), .ZN(\AES_ENC/us33/n729 ) );
NAND2_X2 \AES_ENC/us33/U343  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n729 ), .ZN(\AES_ENC/us33/n730 ) );
NAND4_X2 \AES_ENC/us33/U342  ( .A1(\AES_ENC/us33/n733 ), .A2(\AES_ENC/us33/n732 ), .A3(\AES_ENC/us33/n731 ), .A4(\AES_ENC/us33/n730 ), .ZN(\AES_ENC/sa33_sub[1] ) );
NAND2_X2 \AES_ENC/us33/U341  ( .A1(\AES_ENC/sa33 [7]), .A2(\AES_ENC/us33/n611 ), .ZN(\AES_ENC/us33/n734 ) );
NAND2_X2 \AES_ENC/us33/U340  ( .A1(\AES_ENC/us33/n734 ), .A2(\AES_ENC/us33/n607 ), .ZN(\AES_ENC/us33/n738 ) );
OR4_X2 \AES_ENC/us33/U339  ( .A1(\AES_ENC/us33/n738 ), .A2(\AES_ENC/us33/n626 ), .A3(\AES_ENC/us33/n826 ), .A4(\AES_ENC/us33/n1121 ), .ZN(\AES_ENC/us33/n746 ) );
NAND2_X2 \AES_ENC/us33/U337  ( .A1(\AES_ENC/us33/n1100 ), .A2(\AES_ENC/us33/n587 ), .ZN(\AES_ENC/us33/n992 ) );
OR2_X2 \AES_ENC/us33/U336  ( .A1(\AES_ENC/us33/n610 ), .A2(\AES_ENC/us33/n735 ), .ZN(\AES_ENC/us33/n737 ) );
NAND2_X2 \AES_ENC/us33/U334  ( .A1(\AES_ENC/us33/n619 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n753 ) );
NAND2_X2 \AES_ENC/us33/U333  ( .A1(\AES_ENC/us33/n582 ), .A2(\AES_ENC/us33/n753 ), .ZN(\AES_ENC/us33/n1080 ) );
NAND2_X2 \AES_ENC/us33/U332  ( .A1(\AES_ENC/us33/n1048 ), .A2(\AES_ENC/us33/n576 ), .ZN(\AES_ENC/us33/n736 ) );
NAND2_X2 \AES_ENC/us33/U331  ( .A1(\AES_ENC/us33/n737 ), .A2(\AES_ENC/us33/n736 ), .ZN(\AES_ENC/us33/n739 ) );
NAND2_X2 \AES_ENC/us33/U330  ( .A1(\AES_ENC/us33/n739 ), .A2(\AES_ENC/us33/n738 ), .ZN(\AES_ENC/us33/n745 ) );
NAND2_X2 \AES_ENC/us33/U326  ( .A1(\AES_ENC/us33/n1096 ), .A2(\AES_ENC/us33/n590 ), .ZN(\AES_ENC/us33/n906 ) );
NAND4_X2 \AES_ENC/us33/U323  ( .A1(\AES_ENC/us33/n746 ), .A2(\AES_ENC/us33/n992 ), .A3(\AES_ENC/us33/n745 ), .A4(\AES_ENC/us33/n744 ), .ZN(\AES_ENC/us33/n747 ) );
NAND2_X2 \AES_ENC/us33/U322  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n747 ), .ZN(\AES_ENC/us33/n793 ) );
NAND2_X2 \AES_ENC/us33/U321  ( .A1(\AES_ENC/us33/n584 ), .A2(\AES_ENC/us33/n855 ), .ZN(\AES_ENC/us33/n748 ) );
NAND2_X2 \AES_ENC/us33/U320  ( .A1(\AES_ENC/us33/n956 ), .A2(\AES_ENC/us33/n748 ), .ZN(\AES_ENC/us33/n760 ) );
NAND2_X2 \AES_ENC/us33/U313  ( .A1(\AES_ENC/us33/n590 ), .A2(\AES_ENC/us33/n753 ), .ZN(\AES_ENC/us33/n1023 ) );
NAND4_X2 \AES_ENC/us33/U308  ( .A1(\AES_ENC/us33/n760 ), .A2(\AES_ENC/us33/n992 ), .A3(\AES_ENC/us33/n759 ), .A4(\AES_ENC/us33/n758 ), .ZN(\AES_ENC/us33/n761 ) );
NAND2_X2 \AES_ENC/us33/U307  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n761 ), .ZN(\AES_ENC/us33/n792 ) );
NAND2_X2 \AES_ENC/us33/U306  ( .A1(\AES_ENC/us33/n584 ), .A2(\AES_ENC/us33/n603 ), .ZN(\AES_ENC/us33/n989 ) );
NAND2_X2 \AES_ENC/us33/U305  ( .A1(\AES_ENC/us33/n1050 ), .A2(\AES_ENC/us33/n989 ), .ZN(\AES_ENC/us33/n777 ) );
NAND2_X2 \AES_ENC/us33/U304  ( .A1(\AES_ENC/us33/n1093 ), .A2(\AES_ENC/us33/n762 ), .ZN(\AES_ENC/us33/n776 ) );
XNOR2_X2 \AES_ENC/us33/U301  ( .A(\AES_ENC/sa33 [7]), .B(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n959 ) );
NAND4_X2 \AES_ENC/us33/U289  ( .A1(\AES_ENC/us33/n777 ), .A2(\AES_ENC/us33/n776 ), .A3(\AES_ENC/us33/n775 ), .A4(\AES_ENC/us33/n774 ), .ZN(\AES_ENC/us33/n778 ) );
NAND2_X2 \AES_ENC/us33/U288  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n778 ), .ZN(\AES_ENC/us33/n791 ) );
NAND2_X2 \AES_ENC/us33/U287  ( .A1(\AES_ENC/us33/n1056 ), .A2(\AES_ENC/us33/n1050 ), .ZN(\AES_ENC/us33/n788 ) );
NAND2_X2 \AES_ENC/us33/U286  ( .A1(\AES_ENC/us33/n1091 ), .A2(\AES_ENC/us33/n779 ), .ZN(\AES_ENC/us33/n787 ) );
NAND2_X2 \AES_ENC/us33/U285  ( .A1(\AES_ENC/us33/n956 ), .A2(\AES_ENC/sa33 [1]), .ZN(\AES_ENC/us33/n786 ) );
NAND4_X2 \AES_ENC/us33/U278  ( .A1(\AES_ENC/us33/n788 ), .A2(\AES_ENC/us33/n787 ), .A3(\AES_ENC/us33/n786 ), .A4(\AES_ENC/us33/n785 ), .ZN(\AES_ENC/us33/n789 ) );
NAND2_X2 \AES_ENC/us33/U277  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n789 ), .ZN(\AES_ENC/us33/n790 ) );
NAND4_X2 \AES_ENC/us33/U276  ( .A1(\AES_ENC/us33/n793 ), .A2(\AES_ENC/us33/n792 ), .A3(\AES_ENC/us33/n791 ), .A4(\AES_ENC/us33/n790 ), .ZN(\AES_ENC/sa33_sub[2] ) );
NAND2_X2 \AES_ENC/us33/U275  ( .A1(\AES_ENC/us33/n1059 ), .A2(\AES_ENC/us33/n794 ), .ZN(\AES_ENC/us33/n810 ) );
NAND2_X2 \AES_ENC/us33/U274  ( .A1(\AES_ENC/us33/n1049 ), .A2(\AES_ENC/us33/n956 ), .ZN(\AES_ENC/us33/n809 ) );
OR2_X2 \AES_ENC/us33/U266  ( .A1(\AES_ENC/us33/n1096 ), .A2(\AES_ENC/us33/n606 ), .ZN(\AES_ENC/us33/n802 ) );
NAND2_X2 \AES_ENC/us33/U265  ( .A1(\AES_ENC/us33/n1053 ), .A2(\AES_ENC/us33/n800 ), .ZN(\AES_ENC/us33/n801 ) );
NAND2_X2 \AES_ENC/us33/U264  ( .A1(\AES_ENC/us33/n802 ), .A2(\AES_ENC/us33/n801 ), .ZN(\AES_ENC/us33/n805 ) );
NAND4_X2 \AES_ENC/us33/U261  ( .A1(\AES_ENC/us33/n810 ), .A2(\AES_ENC/us33/n809 ), .A3(\AES_ENC/us33/n808 ), .A4(\AES_ENC/us33/n807 ), .ZN(\AES_ENC/us33/n811 ) );
NAND2_X2 \AES_ENC/us33/U260  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n811 ), .ZN(\AES_ENC/us33/n852 ) );
OR2_X2 \AES_ENC/us33/U259  ( .A1(\AES_ENC/us33/n1023 ), .A2(\AES_ENC/us33/n617 ), .ZN(\AES_ENC/us33/n819 ) );
OR2_X2 \AES_ENC/us33/U257  ( .A1(\AES_ENC/us33/n570 ), .A2(\AES_ENC/us33/n930 ), .ZN(\AES_ENC/us33/n818 ) );
NAND2_X2 \AES_ENC/us33/U256  ( .A1(\AES_ENC/us33/n1013 ), .A2(\AES_ENC/us33/n1094 ), .ZN(\AES_ENC/us33/n817 ) );
NAND4_X2 \AES_ENC/us33/U249  ( .A1(\AES_ENC/us33/n819 ), .A2(\AES_ENC/us33/n818 ), .A3(\AES_ENC/us33/n817 ), .A4(\AES_ENC/us33/n816 ), .ZN(\AES_ENC/us33/n820 ) );
NAND2_X2 \AES_ENC/us33/U248  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n820 ), .ZN(\AES_ENC/us33/n851 ) );
NAND2_X2 \AES_ENC/us33/U247  ( .A1(\AES_ENC/us33/n956 ), .A2(\AES_ENC/us33/n1080 ), .ZN(\AES_ENC/us33/n835 ) );
NAND2_X2 \AES_ENC/us33/U246  ( .A1(\AES_ENC/us33/n570 ), .A2(\AES_ENC/us33/n1030 ), .ZN(\AES_ENC/us33/n1047 ) );
OR2_X2 \AES_ENC/us33/U245  ( .A1(\AES_ENC/us33/n1047 ), .A2(\AES_ENC/us33/n612 ), .ZN(\AES_ENC/us33/n834 ) );
NAND2_X2 \AES_ENC/us33/U244  ( .A1(\AES_ENC/us33/n1072 ), .A2(\AES_ENC/us33/n589 ), .ZN(\AES_ENC/us33/n833 ) );
NAND4_X2 \AES_ENC/us33/U233  ( .A1(\AES_ENC/us33/n835 ), .A2(\AES_ENC/us33/n834 ), .A3(\AES_ENC/us33/n833 ), .A4(\AES_ENC/us33/n832 ), .ZN(\AES_ENC/us33/n836 ) );
NAND2_X2 \AES_ENC/us33/U232  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n836 ), .ZN(\AES_ENC/us33/n850 ) );
NAND2_X2 \AES_ENC/us33/U231  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n623 ), .ZN(\AES_ENC/us33/n847 ) );
NAND2_X2 \AES_ENC/us33/U230  ( .A1(\AES_ENC/us33/n1050 ), .A2(\AES_ENC/us33/n1071 ), .ZN(\AES_ENC/us33/n846 ) );
OR2_X2 \AES_ENC/us33/U224  ( .A1(\AES_ENC/us33/n1053 ), .A2(\AES_ENC/us33/n911 ), .ZN(\AES_ENC/us33/n1077 ) );
NAND4_X2 \AES_ENC/us33/U220  ( .A1(\AES_ENC/us33/n847 ), .A2(\AES_ENC/us33/n846 ), .A3(\AES_ENC/us33/n845 ), .A4(\AES_ENC/us33/n844 ), .ZN(\AES_ENC/us33/n848 ) );
NAND2_X2 \AES_ENC/us33/U219  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n848 ), .ZN(\AES_ENC/us33/n849 ) );
NAND4_X2 \AES_ENC/us33/U218  ( .A1(\AES_ENC/us33/n852 ), .A2(\AES_ENC/us33/n851 ), .A3(\AES_ENC/us33/n850 ), .A4(\AES_ENC/us33/n849 ), .ZN(\AES_ENC/sa33_sub[3] ) );
NAND2_X2 \AES_ENC/us33/U216  ( .A1(\AES_ENC/us33/n1009 ), .A2(\AES_ENC/us33/n1072 ), .ZN(\AES_ENC/us33/n862 ) );
NAND2_X2 \AES_ENC/us33/U215  ( .A1(\AES_ENC/us33/n603 ), .A2(\AES_ENC/us33/n577 ), .ZN(\AES_ENC/us33/n853 ) );
NAND2_X2 \AES_ENC/us33/U214  ( .A1(\AES_ENC/us33/n1050 ), .A2(\AES_ENC/us33/n853 ), .ZN(\AES_ENC/us33/n861 ) );
NAND4_X2 \AES_ENC/us33/U206  ( .A1(\AES_ENC/us33/n862 ), .A2(\AES_ENC/us33/n861 ), .A3(\AES_ENC/us33/n860 ), .A4(\AES_ENC/us33/n859 ), .ZN(\AES_ENC/us33/n863 ) );
NAND2_X2 \AES_ENC/us33/U205  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n863 ), .ZN(\AES_ENC/us33/n905 ) );
NAND2_X2 \AES_ENC/us33/U204  ( .A1(\AES_ENC/us33/n1010 ), .A2(\AES_ENC/us33/n989 ), .ZN(\AES_ENC/us33/n874 ) );
NAND2_X2 \AES_ENC/us33/U203  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n610 ), .ZN(\AES_ENC/us33/n864 ) );
NAND2_X2 \AES_ENC/us33/U202  ( .A1(\AES_ENC/us33/n929 ), .A2(\AES_ENC/us33/n864 ), .ZN(\AES_ENC/us33/n873 ) );
NAND4_X2 \AES_ENC/us33/U193  ( .A1(\AES_ENC/us33/n874 ), .A2(\AES_ENC/us33/n873 ), .A3(\AES_ENC/us33/n872 ), .A4(\AES_ENC/us33/n871 ), .ZN(\AES_ENC/us33/n875 ) );
NAND2_X2 \AES_ENC/us33/U192  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n875 ), .ZN(\AES_ENC/us33/n904 ) );
NAND2_X2 \AES_ENC/us33/U191  ( .A1(\AES_ENC/us33/n583 ), .A2(\AES_ENC/us33/n1050 ), .ZN(\AES_ENC/us33/n889 ) );
NAND2_X2 \AES_ENC/us33/U190  ( .A1(\AES_ENC/us33/n1093 ), .A2(\AES_ENC/us33/n587 ), .ZN(\AES_ENC/us33/n876 ) );
NAND2_X2 \AES_ENC/us33/U189  ( .A1(\AES_ENC/us33/n604 ), .A2(\AES_ENC/us33/n876 ), .ZN(\AES_ENC/us33/n877 ) );
NAND2_X2 \AES_ENC/us33/U188  ( .A1(\AES_ENC/us33/n877 ), .A2(\AES_ENC/us33/n623 ), .ZN(\AES_ENC/us33/n888 ) );
NAND4_X2 \AES_ENC/us33/U179  ( .A1(\AES_ENC/us33/n889 ), .A2(\AES_ENC/us33/n888 ), .A3(\AES_ENC/us33/n887 ), .A4(\AES_ENC/us33/n886 ), .ZN(\AES_ENC/us33/n890 ) );
NAND2_X2 \AES_ENC/us33/U178  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n890 ), .ZN(\AES_ENC/us33/n903 ) );
OR2_X2 \AES_ENC/us33/U177  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n1059 ), .ZN(\AES_ENC/us33/n900 ) );
NAND2_X2 \AES_ENC/us33/U176  ( .A1(\AES_ENC/us33/n1073 ), .A2(\AES_ENC/us33/n1047 ), .ZN(\AES_ENC/us33/n899 ) );
NAND2_X2 \AES_ENC/us33/U175  ( .A1(\AES_ENC/us33/n1094 ), .A2(\AES_ENC/us33/n595 ), .ZN(\AES_ENC/us33/n898 ) );
NAND4_X2 \AES_ENC/us33/U167  ( .A1(\AES_ENC/us33/n900 ), .A2(\AES_ENC/us33/n899 ), .A3(\AES_ENC/us33/n898 ), .A4(\AES_ENC/us33/n897 ), .ZN(\AES_ENC/us33/n901 ) );
NAND2_X2 \AES_ENC/us33/U166  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n901 ), .ZN(\AES_ENC/us33/n902 ) );
NAND4_X2 \AES_ENC/us33/U165  ( .A1(\AES_ENC/us33/n905 ), .A2(\AES_ENC/us33/n904 ), .A3(\AES_ENC/us33/n903 ), .A4(\AES_ENC/us33/n902 ), .ZN(\AES_ENC/sa33_sub[4] ) );
NAND2_X2 \AES_ENC/us33/U164  ( .A1(\AES_ENC/us33/n1094 ), .A2(\AES_ENC/us33/n599 ), .ZN(\AES_ENC/us33/n922 ) );
NAND2_X2 \AES_ENC/us33/U163  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n989 ), .ZN(\AES_ENC/us33/n921 ) );
NAND4_X2 \AES_ENC/us33/U151  ( .A1(\AES_ENC/us33/n922 ), .A2(\AES_ENC/us33/n921 ), .A3(\AES_ENC/us33/n920 ), .A4(\AES_ENC/us33/n919 ), .ZN(\AES_ENC/us33/n923 ) );
NAND2_X2 \AES_ENC/us33/U150  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n923 ), .ZN(\AES_ENC/us33/n972 ) );
NAND2_X2 \AES_ENC/us33/U149  ( .A1(\AES_ENC/us33/n582 ), .A2(\AES_ENC/us33/n619 ), .ZN(\AES_ENC/us33/n924 ) );
NAND2_X2 \AES_ENC/us33/U148  ( .A1(\AES_ENC/us33/n1073 ), .A2(\AES_ENC/us33/n924 ), .ZN(\AES_ENC/us33/n939 ) );
NAND2_X2 \AES_ENC/us33/U147  ( .A1(\AES_ENC/us33/n926 ), .A2(\AES_ENC/us33/n925 ), .ZN(\AES_ENC/us33/n927 ) );
NAND2_X2 \AES_ENC/us33/U146  ( .A1(\AES_ENC/us33/n606 ), .A2(\AES_ENC/us33/n927 ), .ZN(\AES_ENC/us33/n928 ) );
NAND2_X2 \AES_ENC/us33/U145  ( .A1(\AES_ENC/us33/n928 ), .A2(\AES_ENC/us33/n1080 ), .ZN(\AES_ENC/us33/n938 ) );
OR2_X2 \AES_ENC/us33/U144  ( .A1(\AES_ENC/us33/n1117 ), .A2(\AES_ENC/us33/n615 ), .ZN(\AES_ENC/us33/n937 ) );
NAND4_X2 \AES_ENC/us33/U139  ( .A1(\AES_ENC/us33/n939 ), .A2(\AES_ENC/us33/n938 ), .A3(\AES_ENC/us33/n937 ), .A4(\AES_ENC/us33/n936 ), .ZN(\AES_ENC/us33/n940 ) );
NAND2_X2 \AES_ENC/us33/U138  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n940 ), .ZN(\AES_ENC/us33/n971 ) );
OR2_X2 \AES_ENC/us33/U137  ( .A1(\AES_ENC/us33/n605 ), .A2(\AES_ENC/us33/n941 ), .ZN(\AES_ENC/us33/n954 ) );
NAND2_X2 \AES_ENC/us33/U136  ( .A1(\AES_ENC/us33/n1096 ), .A2(\AES_ENC/us33/n577 ), .ZN(\AES_ENC/us33/n942 ) );
NAND2_X2 \AES_ENC/us33/U135  ( .A1(\AES_ENC/us33/n1048 ), .A2(\AES_ENC/us33/n942 ), .ZN(\AES_ENC/us33/n943 ) );
NAND2_X2 \AES_ENC/us33/U134  ( .A1(\AES_ENC/us33/n612 ), .A2(\AES_ENC/us33/n943 ), .ZN(\AES_ENC/us33/n944 ) );
NAND2_X2 \AES_ENC/us33/U133  ( .A1(\AES_ENC/us33/n944 ), .A2(\AES_ENC/us33/n580 ), .ZN(\AES_ENC/us33/n953 ) );
NAND4_X2 \AES_ENC/us33/U125  ( .A1(\AES_ENC/us33/n954 ), .A2(\AES_ENC/us33/n953 ), .A3(\AES_ENC/us33/n952 ), .A4(\AES_ENC/us33/n951 ), .ZN(\AES_ENC/us33/n955 ) );
NAND2_X2 \AES_ENC/us33/U124  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n955 ), .ZN(\AES_ENC/us33/n970 ) );
NAND2_X2 \AES_ENC/us33/U123  ( .A1(\AES_ENC/us33/n1094 ), .A2(\AES_ENC/us33/n1071 ), .ZN(\AES_ENC/us33/n967 ) );
NAND2_X2 \AES_ENC/us33/U122  ( .A1(\AES_ENC/us33/n956 ), .A2(\AES_ENC/us33/n1030 ), .ZN(\AES_ENC/us33/n966 ) );
NAND4_X2 \AES_ENC/us33/U114  ( .A1(\AES_ENC/us33/n967 ), .A2(\AES_ENC/us33/n966 ), .A3(\AES_ENC/us33/n965 ), .A4(\AES_ENC/us33/n964 ), .ZN(\AES_ENC/us33/n968 ) );
NAND2_X2 \AES_ENC/us33/U113  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n968 ), .ZN(\AES_ENC/us33/n969 ) );
NAND4_X2 \AES_ENC/us33/U112  ( .A1(\AES_ENC/us33/n972 ), .A2(\AES_ENC/us33/n971 ), .A3(\AES_ENC/us33/n970 ), .A4(\AES_ENC/us33/n969 ), .ZN(\AES_ENC/sa33_sub[5] ) );
NAND2_X2 \AES_ENC/us33/U111  ( .A1(\AES_ENC/us33/n570 ), .A2(\AES_ENC/us33/n1097 ), .ZN(\AES_ENC/us33/n973 ) );
NAND2_X2 \AES_ENC/us33/U110  ( .A1(\AES_ENC/us33/n1073 ), .A2(\AES_ENC/us33/n973 ), .ZN(\AES_ENC/us33/n987 ) );
NAND2_X2 \AES_ENC/us33/U109  ( .A1(\AES_ENC/us33/n974 ), .A2(\AES_ENC/us33/n1077 ), .ZN(\AES_ENC/us33/n975 ) );
NAND2_X2 \AES_ENC/us33/U108  ( .A1(\AES_ENC/us33/n613 ), .A2(\AES_ENC/us33/n975 ), .ZN(\AES_ENC/us33/n976 ) );
NAND2_X2 \AES_ENC/us33/U107  ( .A1(\AES_ENC/us33/n977 ), .A2(\AES_ENC/us33/n976 ), .ZN(\AES_ENC/us33/n986 ) );
NAND4_X2 \AES_ENC/us33/U99  ( .A1(\AES_ENC/us33/n987 ), .A2(\AES_ENC/us33/n986 ), .A3(\AES_ENC/us33/n985 ), .A4(\AES_ENC/us33/n984 ), .ZN(\AES_ENC/us33/n988 ) );
NAND2_X2 \AES_ENC/us33/U98  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n988 ), .ZN(\AES_ENC/us33/n1044 ) );
NAND2_X2 \AES_ENC/us33/U97  ( .A1(\AES_ENC/us33/n1073 ), .A2(\AES_ENC/us33/n989 ), .ZN(\AES_ENC/us33/n1004 ) );
NAND2_X2 \AES_ENC/us33/U96  ( .A1(\AES_ENC/us33/n1092 ), .A2(\AES_ENC/us33/n619 ), .ZN(\AES_ENC/us33/n1003 ) );
NAND4_X2 \AES_ENC/us33/U85  ( .A1(\AES_ENC/us33/n1004 ), .A2(\AES_ENC/us33/n1003 ), .A3(\AES_ENC/us33/n1002 ), .A4(\AES_ENC/us33/n1001 ), .ZN(\AES_ENC/us33/n1005 ) );
NAND2_X2 \AES_ENC/us33/U84  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n1005 ), .ZN(\AES_ENC/us33/n1043 ) );
NAND2_X2 \AES_ENC/us33/U83  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n596 ), .ZN(\AES_ENC/us33/n1020 ) );
NAND2_X2 \AES_ENC/us33/U82  ( .A1(\AES_ENC/us33/n1050 ), .A2(\AES_ENC/us33/n624 ), .ZN(\AES_ENC/us33/n1019 ) );
NAND2_X2 \AES_ENC/us33/U77  ( .A1(\AES_ENC/us33/n1059 ), .A2(\AES_ENC/us33/n1114 ), .ZN(\AES_ENC/us33/n1012 ) );
NAND2_X2 \AES_ENC/us33/U76  ( .A1(\AES_ENC/us33/n1010 ), .A2(\AES_ENC/us33/n592 ), .ZN(\AES_ENC/us33/n1011 ) );
NAND2_X2 \AES_ENC/us33/U75  ( .A1(\AES_ENC/us33/n1012 ), .A2(\AES_ENC/us33/n1011 ), .ZN(\AES_ENC/us33/n1016 ) );
NAND4_X2 \AES_ENC/us33/U70  ( .A1(\AES_ENC/us33/n1020 ), .A2(\AES_ENC/us33/n1019 ), .A3(\AES_ENC/us33/n1018 ), .A4(\AES_ENC/us33/n1017 ), .ZN(\AES_ENC/us33/n1021 ) );
NAND2_X2 \AES_ENC/us33/U69  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n1021 ), .ZN(\AES_ENC/us33/n1042 ) );
NAND2_X2 \AES_ENC/us33/U68  ( .A1(\AES_ENC/us33/n1022 ), .A2(\AES_ENC/us33/n1093 ), .ZN(\AES_ENC/us33/n1039 ) );
NAND2_X2 \AES_ENC/us33/U67  ( .A1(\AES_ENC/us33/n1050 ), .A2(\AES_ENC/us33/n1023 ), .ZN(\AES_ENC/us33/n1038 ) );
NAND2_X2 \AES_ENC/us33/U66  ( .A1(\AES_ENC/us33/n1024 ), .A2(\AES_ENC/us33/n1071 ), .ZN(\AES_ENC/us33/n1037 ) );
AND2_X2 \AES_ENC/us33/U60  ( .A1(\AES_ENC/us33/n1030 ), .A2(\AES_ENC/us33/n602 ), .ZN(\AES_ENC/us33/n1078 ) );
NAND4_X2 \AES_ENC/us33/U56  ( .A1(\AES_ENC/us33/n1039 ), .A2(\AES_ENC/us33/n1038 ), .A3(\AES_ENC/us33/n1037 ), .A4(\AES_ENC/us33/n1036 ), .ZN(\AES_ENC/us33/n1040 ) );
NAND2_X2 \AES_ENC/us33/U55  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n1040 ), .ZN(\AES_ENC/us33/n1041 ) );
NAND4_X2 \AES_ENC/us33/U54  ( .A1(\AES_ENC/us33/n1044 ), .A2(\AES_ENC/us33/n1043 ), .A3(\AES_ENC/us33/n1042 ), .A4(\AES_ENC/us33/n1041 ), .ZN(\AES_ENC/sa33_sub[6] ) );
NAND2_X2 \AES_ENC/us33/U53  ( .A1(\AES_ENC/us33/n1072 ), .A2(\AES_ENC/us33/n1045 ), .ZN(\AES_ENC/us33/n1068 ) );
NAND2_X2 \AES_ENC/us33/U52  ( .A1(\AES_ENC/us33/n1046 ), .A2(\AES_ENC/us33/n582 ), .ZN(\AES_ENC/us33/n1067 ) );
NAND2_X2 \AES_ENC/us33/U51  ( .A1(\AES_ENC/us33/n1094 ), .A2(\AES_ENC/us33/n1047 ), .ZN(\AES_ENC/us33/n1066 ) );
NAND4_X2 \AES_ENC/us33/U40  ( .A1(\AES_ENC/us33/n1068 ), .A2(\AES_ENC/us33/n1067 ), .A3(\AES_ENC/us33/n1066 ), .A4(\AES_ENC/us33/n1065 ), .ZN(\AES_ENC/us33/n1069 ) );
NAND2_X2 \AES_ENC/us33/U39  ( .A1(\AES_ENC/us33/n1070 ), .A2(\AES_ENC/us33/n1069 ), .ZN(\AES_ENC/us33/n1135 ) );
NAND2_X2 \AES_ENC/us33/U38  ( .A1(\AES_ENC/us33/n1072 ), .A2(\AES_ENC/us33/n1071 ), .ZN(\AES_ENC/us33/n1088 ) );
NAND2_X2 \AES_ENC/us33/U37  ( .A1(\AES_ENC/us33/n1073 ), .A2(\AES_ENC/us33/n595 ), .ZN(\AES_ENC/us33/n1087 ) );
NAND4_X2 \AES_ENC/us33/U28  ( .A1(\AES_ENC/us33/n1088 ), .A2(\AES_ENC/us33/n1087 ), .A3(\AES_ENC/us33/n1086 ), .A4(\AES_ENC/us33/n1085 ), .ZN(\AES_ENC/us33/n1089 ) );
NAND2_X2 \AES_ENC/us33/U27  ( .A1(\AES_ENC/us33/n1090 ), .A2(\AES_ENC/us33/n1089 ), .ZN(\AES_ENC/us33/n1134 ) );
NAND2_X2 \AES_ENC/us33/U26  ( .A1(\AES_ENC/us33/n1091 ), .A2(\AES_ENC/us33/n1093 ), .ZN(\AES_ENC/us33/n1111 ) );
NAND2_X2 \AES_ENC/us33/U25  ( .A1(\AES_ENC/us33/n1092 ), .A2(\AES_ENC/us33/n1120 ), .ZN(\AES_ENC/us33/n1110 ) );
AND2_X2 \AES_ENC/us33/U22  ( .A1(\AES_ENC/us33/n1097 ), .A2(\AES_ENC/us33/n1096 ), .ZN(\AES_ENC/us33/n1098 ) );
NAND4_X2 \AES_ENC/us33/U14  ( .A1(\AES_ENC/us33/n1111 ), .A2(\AES_ENC/us33/n1110 ), .A3(\AES_ENC/us33/n1109 ), .A4(\AES_ENC/us33/n1108 ), .ZN(\AES_ENC/us33/n1112 ) );
NAND2_X2 \AES_ENC/us33/U13  ( .A1(\AES_ENC/us33/n1113 ), .A2(\AES_ENC/us33/n1112 ), .ZN(\AES_ENC/us33/n1133 ) );
NAND2_X2 \AES_ENC/us33/U12  ( .A1(\AES_ENC/us33/n1115 ), .A2(\AES_ENC/us33/n1114 ), .ZN(\AES_ENC/us33/n1129 ) );
OR2_X2 \AES_ENC/us33/U11  ( .A1(\AES_ENC/us33/n608 ), .A2(\AES_ENC/us33/n1116 ), .ZN(\AES_ENC/us33/n1128 ) );
NAND4_X2 \AES_ENC/us33/U3  ( .A1(\AES_ENC/us33/n1129 ), .A2(\AES_ENC/us33/n1128 ), .A3(\AES_ENC/us33/n1127 ), .A4(\AES_ENC/us33/n1126 ), .ZN(\AES_ENC/us33/n1130 ) );
NAND2_X2 \AES_ENC/us33/U2  ( .A1(\AES_ENC/us33/n1131 ), .A2(\AES_ENC/us33/n1130 ), .ZN(\AES_ENC/us33/n1132 ) );
NAND4_X2 \AES_ENC/us33/U1  ( .A1(\AES_ENC/us33/n1135 ), .A2(\AES_ENC/us33/n1134 ), .A3(\AES_ENC/us33/n1133 ), .A4(\AES_ENC/us33/n1132 ), .ZN(\AES_ENC/sa33_sub[7] ) );
INV_X4 \add_506/U775  ( .A(n18589), .ZN(N2027) );
NAND2_X2 \add_506/U774  ( .A1(n18233), .A2(n18237), .ZN(\add_506/n646 ) );
NAND2_X2 \add_506/U773  ( .A1(n18225), .A2(n18229), .ZN(\add_506/n647 ) );
NAND2_X2 \add_506/U772  ( .A1(n18249), .A2(n18253), .ZN(\add_506/n644 ) );
NAND2_X2 \add_506/U771  ( .A1(n18241), .A2(n18245), .ZN(\add_506/n645 ) );
NAND4_X2 \add_506/U770  ( .A1(n18273), .A2(n18277), .A3(n18281), .A4(n18285),.ZN(\add_506/n642 ) );
NAND4_X2 \add_506/U769  ( .A1(n18257), .A2(n18261), .A3(n18265), .A4(n18269),.ZN(\add_506/n643 ) );
INV_X4 \add_506/U768  ( .A(\add_506/n37 ), .ZN(\add_506/n63 ) );
NAND4_X2 \add_506/U767  ( .A1(n18301), .A2(n18305), .A3(n18309), .A4(n18313),.ZN(\add_506/n637 ) );
NAND4_X2 \add_506/U766  ( .A1(n18329), .A2(n18333), .A3(n18337), .A4(n18341),.ZN(\add_506/n635 ) );
NAND4_X2 \add_506/U765  ( .A1(n18357), .A2(n18361), .A3(n18365), .A4(n18369),.ZN(\add_506/n633 ) );
NAND4_X2 \add_506/U764  ( .A1(n18385), .A2(n18389), .A3(n18393), .A4(n18397),.ZN(\add_506/n631 ) );
NAND2_X2 \add_506/U763  ( .A1(n18409), .A2(n18413), .ZN(\add_506/n625 ) );
NAND2_X2 \add_506/U762  ( .A1(n18401), .A2(n18405), .ZN(\add_506/n626 ) );
NAND2_X2 \add_506/U761  ( .A1(n18425), .A2(n18429), .ZN(\add_506/n623 ) );
NAND2_X2 \add_506/U760  ( .A1(n18417), .A2(n18421), .ZN(\add_506/n624 ) );
NAND4_X2 \add_506/U759  ( .A1(n18449), .A2(n18453), .A3(n18457), .A4(n18461),.ZN(\add_506/n621 ) );
NAND4_X2 \add_506/U758  ( .A1(n18433), .A2(n18437), .A3(n18441), .A4(n18445),.ZN(\add_506/n622 ) );
INV_X4 \add_506/U757  ( .A(n18197), .ZN(\add_506/n617 ) );
INV_X4 \add_506/U756  ( .A(n18193), .ZN(\add_506/n31 ) );
INV_X4 \add_506/U755  ( .A(n18205), .ZN(\add_506/n39 ) );
INV_X4 \add_506/U754  ( .A(n18201), .ZN(\add_506/n616 ) );
NAND2_X2 \add_506/U753  ( .A1(n18217), .A2(n18221), .ZN(\add_506/n614 ) );
NAND2_X2 \add_506/U752  ( .A1(n18209), .A2(n18213), .ZN(\add_506/n615 ) );
NAND4_X2 \add_506/U751  ( .A1(n18481), .A2(n18485), .A3(n18489), .A4(n18493),.ZN(\add_506/n609 ) );
NAND4_X2 \add_506/U750  ( .A1(n18465), .A2(n18469), .A3(n18473), .A4(n18477),.ZN(\add_506/n610 ) );
NAND4_X2 \add_506/U749  ( .A1(n18513), .A2(n18517), .A3(n18521), .A4(n18525),.ZN(\add_506/n607 ) );
NAND4_X2 \add_506/U748  ( .A1(n18497), .A2(n18501), .A3(n18505), .A4(n18509),.ZN(\add_506/n608 ) );
NAND2_X2 \add_506/U747  ( .A1(n18569), .A2(n18573), .ZN(\add_506/n605 ) );
NAND2_X2 \add_506/U746  ( .A1(n18561), .A2(n18565), .ZN(\add_506/n606 ) );
NAND2_X2 \add_506/U745  ( .A1(n18585), .A2(n18589), .ZN(\add_506/n603 ) );
NAND2_X2 \add_506/U744  ( .A1(n18577), .A2(n18581), .ZN(\add_506/n604 ) );
NAND2_X2 \add_506/U743  ( .A1(\add_506/n601 ), .A2(\add_506/n602 ), .ZN(\add_506/n598 ) );
NAND4_X2 \add_506/U742  ( .A1(n18545), .A2(n18549), .A3(n18553), .A4(n18557),.ZN(\add_506/n599 ) );
NAND4_X2 \add_506/U741  ( .A1(n18529), .A2(n18533), .A3(n18537), .A4(n18541),.ZN(\add_506/n600 ) );
NAND4_X2 \add_506/U740  ( .A1(\add_506/n63 ), .A2(\add_506/n20 ), .A3(\add_506/n594 ), .A4(\add_506/n15 ), .ZN(\add_506/n593 ) );
XNOR2_X2 \add_506/U739  ( .A(\add_506/n593 ), .B(n18189), .ZN(N2127) );
INV_X4 \add_506/U738  ( .A(\add_506/n584 ), .ZN(\add_506/n592 ) );
NAND2_X2 \add_506/U737  ( .A1(n18189), .A2(\add_506/n592 ), .ZN(\add_506/n591 ) );
NAND4_X2 \add_506/U736  ( .A1(\add_506/n63 ), .A2(\add_506/n20 ), .A3(\add_506/n590 ), .A4(\add_506/n15 ), .ZN(\add_506/n589 ) );
XNOR2_X2 \add_506/U735  ( .A(\add_506/n589 ), .B(n18185), .ZN(N2128) );
NAND2_X2 \add_506/U734  ( .A1(n18185), .A2(n18189), .ZN(\add_506/n588 ) );
NAND4_X2 \add_506/U733  ( .A1(\add_506/n63 ), .A2(\add_506/n16 ), .A3(\add_506/n587 ), .A4(\add_506/n19 ), .ZN(\add_506/n586 ) );
XNOR2_X2 \add_506/U732  ( .A(\add_506/n586 ), .B(n18181), .ZN(N2129) );
NAND4_X2 \add_506/U731  ( .A1(\add_506/n63 ), .A2(\add_506/n17 ), .A3(\add_506/n583 ), .A4(\add_506/n19 ), .ZN(\add_506/n582 ) );
XNOR2_X2 \add_506/U730  ( .A(\add_506/n582 ), .B(n18177), .ZN(N2130) );
NAND2_X2 \add_506/U729  ( .A1(n18217), .A2(n18221), .ZN(\add_506/n580 ) );
NAND2_X2 \add_506/U728  ( .A1(n18209), .A2(n18213), .ZN(\add_506/n581 ) );
NAND4_X2 \add_506/U727  ( .A1(n18193), .A2(n18197), .A3(n18201), .A4(n18205),.ZN(\add_506/n578 ) );
NAND4_X2 \add_506/U726  ( .A1(n18177), .A2(n18181), .A3(n18185), .A4(n18189),.ZN(\add_506/n579 ) );
NAND4_X2 \add_506/U725  ( .A1(\add_506/n576 ), .A2(\add_506/n20 ), .A3(\add_506/n16 ), .A4(\add_506/n577 ), .ZN(\add_506/n575 ) );
XNOR2_X2 \add_506/U724  ( .A(\add_506/n575 ), .B(n18173), .ZN(N2131) );
NAND4_X2 \add_506/U723  ( .A1(n18209), .A2(n18221), .A3(n18217), .A4(n18213),.ZN(\add_506/n572 ) );
NAND4_X2 \add_506/U722  ( .A1(n18189), .A2(n18193), .A3(n18197), .A4(n18201),.ZN(\add_506/n573 ) );
NAND4_X2 \add_506/U721  ( .A1(n18173), .A2(n18177), .A3(n18181), .A4(n18185),.ZN(\add_506/n574 ) );
NAND4_X2 \add_506/U720  ( .A1(\add_506/n19 ), .A2(\add_506/n570 ), .A3(\add_506/n16 ), .A4(\add_506/n571 ), .ZN(\add_506/n569 ) );
XNOR2_X2 \add_506/U719  ( .A(\add_506/n569 ), .B(n18169), .ZN(N2132) );
INV_X4 \add_506/U718  ( .A(n18173), .ZN(\add_506/n555 ) );
INV_X4 \add_506/U717  ( .A(n18169), .ZN(\add_506/n556 ) );
INV_X4 \add_506/U716  ( .A(n18181), .ZN(\add_506/n553 ) );
INV_X4 \add_506/U715  ( .A(n18177), .ZN(\add_506/n554 ) );
INV_X4 \add_506/U714  ( .A(n18189), .ZN(\add_506/n568 ) );
INV_X4 \add_506/U713  ( .A(n18185), .ZN(\add_506/n552 ) );
NAND3_X2 \add_506/U712  ( .A1(\add_506/n565 ), .A2(\add_506/n566 ), .A3(\add_506/n567 ), .ZN(\add_506/n562 ) );
NAND4_X2 \add_506/U711  ( .A1(n18209), .A2(n18221), .A3(n18217), .A4(n18213),.ZN(\add_506/n563 ) );
NAND4_X2 \add_506/U710  ( .A1(\add_506/n19 ), .A2(\add_506/n560 ), .A3(\add_506/n16 ), .A4(\add_506/n561 ), .ZN(\add_506/n559 ) );
XNOR2_X2 \add_506/U709  ( .A(\add_506/n559 ), .B(n18165), .ZN(N2133) );
NAND2_X2 \add_506/U708  ( .A1(n18201), .A2(n18205), .ZN(\add_506/n558 ) );
INV_X4 \add_506/U707  ( .A(n18165), .ZN(\add_506/n557 ) );
NAND3_X2 \add_506/U706  ( .A1(\add_506/n549 ), .A2(\add_506/n550 ), .A3(\add_506/n551 ), .ZN(\add_506/n546 ) );
NAND4_X2 \add_506/U705  ( .A1(n18209), .A2(n18221), .A3(n18217), .A4(n18213),.ZN(\add_506/n547 ) );
NAND4_X2 \add_506/U704  ( .A1(\add_506/n20 ), .A2(\add_506/n544 ), .A3(\add_506/n16 ), .A4(\add_506/n545 ), .ZN(\add_506/n543 ) );
XNOR2_X2 \add_506/U703  ( .A(\add_506/n543 ), .B(n18161), .ZN(N2134) );
NAND4_X2 \add_506/U702  ( .A1(n18177), .A2(n18181), .A3(n18185), .A4(n18189),.ZN(\add_506/n541 ) );
NAND4_X2 \add_506/U701  ( .A1(n18161), .A2(n18165), .A3(n18169), .A4(n18173),.ZN(\add_506/n542 ) );
NAND4_X2 \add_506/U700  ( .A1(n18209), .A2(n18213), .A3(n18217), .A4(n18221),.ZN(\add_506/n539 ) );
NAND4_X2 \add_506/U699  ( .A1(n18193), .A2(n18197), .A3(n18201), .A4(n18205),.ZN(\add_506/n540 ) );
NAND2_X2 \add_506/U698  ( .A1(n18265), .A2(n18269), .ZN(\add_506/n537 ) );
NAND2_X2 \add_506/U697  ( .A1(n18257), .A2(n18261), .ZN(\add_506/n538 ) );
NAND2_X2 \add_506/U696  ( .A1(n18281), .A2(n18285), .ZN(\add_506/n535 ) );
NAND2_X2 \add_506/U695  ( .A1(n18273), .A2(n18277), .ZN(\add_506/n536 ) );
NAND2_X2 \add_506/U694  ( .A1(\add_506/n533 ), .A2(\add_506/n534 ), .ZN(\add_506/n530 ) );
NAND4_X2 \add_506/U693  ( .A1(n18241), .A2(n18245), .A3(n18249), .A4(n18253),.ZN(\add_506/n531 ) );
NAND4_X2 \add_506/U692  ( .A1(n18225), .A2(n18229), .A3(n18233), .A4(n18237),.ZN(\add_506/n532 ) );
NAND4_X2 \add_506/U691  ( .A1(\add_506/n398 ), .A2(\add_506/n27 ), .A3(\add_506/n19 ), .A4(\add_506/n15 ), .ZN(\add_506/n526 ) );
XNOR2_X2 \add_506/U690  ( .A(\add_506/n526 ), .B(n18157), .ZN(N2135) );
INV_X4 \add_506/U689  ( .A(n18153), .ZN(\add_506/n427 ) );
NAND3_X2 \add_506/U688  ( .A1(n18157), .A2(\add_506/n398 ), .A3(\add_506/n17 ), .ZN(\add_506/n524 ) );
NAND2_X2 \add_506/U687  ( .A1(\add_506/n22 ), .A2(\add_506/n28 ), .ZN(\add_506/n525 ) );
XNOR2_X2 \add_506/U686  ( .A(\add_506/n427 ), .B(\add_506/n523 ), .ZN(N2136));
NAND2_X2 \add_506/U685  ( .A1(n18565), .A2(n18561), .ZN(\add_506/n520 ) );
NAND4_X2 \add_506/U684  ( .A1(n18577), .A2(n18581), .A3(n18585), .A4(n18589),.ZN(\add_506/n521 ) );
NAND2_X2 \add_506/U683  ( .A1(n18569), .A2(n18573), .ZN(\add_506/n522 ) );
NAND2_X2 \add_506/U682  ( .A1(\add_506/n3 ), .A2(\add_506/n30 ), .ZN(\add_506/n519 ) );
XNOR2_X2 \add_506/U681  ( .A(\add_506/n519 ), .B(n18549), .ZN(N2037) );
NAND3_X2 \add_506/U680  ( .A1(\add_506/n518 ), .A2(\add_506/n398 ), .A3(\add_506/n17 ), .ZN(\add_506/n516 ) );
NAND2_X2 \add_506/U679  ( .A1(\add_506/n22 ), .A2(\add_506/n28 ), .ZN(\add_506/n517 ) );
NAND4_X2 \add_506/U678  ( .A1(\add_506/n20 ), .A2(\add_506/n16 ), .A3(\add_506/n514 ), .A4(\add_506/n398 ), .ZN(\add_506/n513 ) );
XNOR2_X2 \add_506/U677  ( .A(\add_506/n513 ), .B(n18145), .ZN(N2138) );
INV_X4 \add_506/U676  ( .A(n18141), .ZN(\add_506/n493 ) );
NAND4_X2 \add_506/U675  ( .A1(n18145), .A2(n18149), .A3(n18153), .A4(n18157),.ZN(\add_506/n505 ) );
INV_X4 \add_506/U674  ( .A(\add_506/n505 ), .ZN(\add_506/n500 ) );
NAND3_X2 \add_506/U673  ( .A1(\add_506/n500 ), .A2(\add_506/n398 ), .A3(\add_506/n17 ), .ZN(\add_506/n511 ) );
NAND2_X2 \add_506/U672  ( .A1(\add_506/n22 ), .A2(\add_506/n28 ), .ZN(\add_506/n512 ) );
XNOR2_X2 \add_506/U671  ( .A(\add_506/n493 ), .B(\add_506/n510 ), .ZN(N2139));
INV_X4 \add_506/U670  ( .A(n18137), .ZN(\add_506/n494 ) );
NAND3_X2 \add_506/U669  ( .A1(\add_506/n509 ), .A2(\add_506/n398 ), .A3(\add_506/n17 ), .ZN(\add_506/n507 ) );
NAND2_X2 \add_506/U668  ( .A1(\add_506/n22 ), .A2(\add_506/n28 ), .ZN(\add_506/n508 ) );
XNOR2_X2 \add_506/U667  ( .A(\add_506/n494 ), .B(\add_506/n506 ), .ZN(N2140));
NAND4_X2 \add_506/U666  ( .A1(\add_506/n503 ), .A2(\add_506/n27 ), .A3(\add_506/n398 ), .A4(\add_506/n504 ), .ZN(\add_506/n502 ) );
XNOR2_X2 \add_506/U665  ( .A(\add_506/n502 ), .B(n18133), .ZN(N2141) );
NAND2_X2 \add_506/U664  ( .A1(n18137), .A2(n18133), .ZN(\add_506/n501 ) );
NAND2_X2 \add_506/U663  ( .A1(\add_506/n499 ), .A2(\add_506/n500 ), .ZN(\add_506/n498 ) );
NAND4_X2 \add_506/U662  ( .A1(\add_506/n20 ), .A2(\add_506/n16 ), .A3(\add_506/n497 ), .A4(\add_506/n398 ), .ZN(\add_506/n496 ) );
XNOR2_X2 \add_506/U661  ( .A(\add_506/n496 ), .B(n18129), .ZN(N2142) );
INV_X4 \add_506/U660  ( .A(n18125), .ZN(\add_506/n465 ) );
INV_X4 \add_506/U659  ( .A(n18133), .ZN(\add_506/n495 ) );
NAND2_X2 \add_506/U658  ( .A1(n18153), .A2(n18157), .ZN(\add_506/n491 ) );
NAND2_X2 \add_506/U657  ( .A1(n18145), .A2(n18149), .ZN(\add_506/n492 ) );
INV_X4 \add_506/U656  ( .A(\add_506/n474 ), .ZN(\add_506/n481 ) );
NAND3_X2 \add_506/U655  ( .A1(\add_506/n481 ), .A2(\add_506/n398 ), .A3(\add_506/n17 ), .ZN(\add_506/n486 ) );
NAND2_X2 \add_506/U654  ( .A1(\add_506/n22 ), .A2(\add_506/n27 ), .ZN(\add_506/n487 ) );
XNOR2_X2 \add_506/U653  ( .A(\add_506/n465 ), .B(\add_506/n485 ), .ZN(N2143));
INV_X4 \add_506/U652  ( .A(n18121), .ZN(\add_506/n475 ) );
NAND4_X2 \add_506/U651  ( .A1(\add_506/n398 ), .A2(\add_506/n16 ), .A3(\add_506/n481 ), .A4(n18125), .ZN(\add_506/n483 ) );
NAND2_X2 \add_506/U650  ( .A1(\add_506/n22 ), .A2(\add_506/n27 ), .ZN(\add_506/n484 ) );
XNOR2_X2 \add_506/U649  ( .A(\add_506/n475 ), .B(\add_506/n482 ), .ZN(N2144));
INV_X4 \add_506/U648  ( .A(n18117), .ZN(\add_506/n473 ) );
AND2_X2 \add_506/U647  ( .A1(\add_506/n481 ), .A2(n18121), .ZN(\add_506/n480 ) );
NAND3_X2 \add_506/U646  ( .A1(\add_506/n480 ), .A2(\add_506/n398 ), .A3(\add_506/n17 ), .ZN(\add_506/n477 ) );
NAND2_X2 \add_506/U645  ( .A1(\add_506/n21 ), .A2(\add_506/n479 ), .ZN(\add_506/n478 ) );
XNOR2_X2 \add_506/U644  ( .A(\add_506/n473 ), .B(\add_506/n476 ), .ZN(N2145));
NAND4_X2 \add_506/U643  ( .A1(\add_506/n398 ), .A2(\add_506/n16 ), .A3(\add_506/n471 ), .A4(\add_506/n472 ), .ZN(\add_506/n470 ) );
XNOR2_X2 \add_506/U642  ( .A(\add_506/n470 ), .B(n18113), .ZN(N2146) );
XNOR2_X2 \add_506/U641  ( .A(\add_506/n469 ), .B(n18545), .ZN(N2038) );
NAND4_X2 \add_506/U640  ( .A1(n18145), .A2(n18149), .A3(n18153), .A4(n18157),.ZN(\add_506/n466 ) );
NAND4_X2 \add_506/U639  ( .A1(n18129), .A2(n18133), .A3(n18137), .A4(n18141),.ZN(\add_506/n467 ) );
NAND2_X2 \add_506/U638  ( .A1(\add_506/n27 ), .A2(\add_506/n464 ), .ZN(\add_506/n463 ) );
NAND3_X2 \add_506/U637  ( .A1(\add_506/n17 ), .A2(\add_506/n461 ), .A3(\add_506/n462 ), .ZN(\add_506/n460 ) );
XNOR2_X2 \add_506/U636  ( .A(\add_506/n460 ), .B(n18109), .ZN(N2147) );
NAND2_X2 \add_506/U635  ( .A1(n18137), .A2(n18145), .ZN(\add_506/n459 ) );
NAND4_X2 \add_506/U634  ( .A1(\add_506/n20 ), .A2(\add_506/n454 ), .A3(\add_506/n455 ), .A4(\add_506/n456 ), .ZN(\add_506/n453 ) );
XNOR2_X2 \add_506/U633  ( .A(n18105), .B(\add_506/n453 ), .ZN(N2148) );
NAND2_X2 \add_506/U632  ( .A1(n18157), .A2(n18153), .ZN(\add_506/n452 ) );
NAND4_X2 \add_506/U631  ( .A1(n18129), .A2(n18133), .A3(n18145), .A4(n18149),.ZN(\add_506/n449 ) );
NAND2_X2 \add_506/U630  ( .A1(n18137), .A2(n18141), .ZN(\add_506/n450 ) );
NOR2_X2 \add_506/U629  ( .A1(\add_506/n449 ), .A2(\add_506/n450 ), .ZN(\add_506/n448 ) );
INV_X4 \add_506/U628  ( .A(\add_506/n8 ), .ZN(\add_506/n436 ) );
NAND2_X2 \add_506/U627  ( .A1(\add_506/n448 ), .A2(\add_506/n436 ), .ZN(\add_506/n447 ) );
INV_X4 \add_506/U626  ( .A(n18105), .ZN(\add_506/n434 ) );
NAND2_X2 \add_506/U625  ( .A1(\add_506/n27 ), .A2(\add_506/n446 ), .ZN(\add_506/n445 ) );
NAND3_X2 \add_506/U624  ( .A1(\add_506/n17 ), .A2(\add_506/n443 ), .A3(\add_506/n444 ), .ZN(\add_506/n442 ) );
XNOR2_X2 \add_506/U623  ( .A(\add_506/n442 ), .B(n18101), .ZN(N2149) );
NAND2_X2 \add_506/U622  ( .A1(n18153), .A2(n18101), .ZN(\add_506/n441 ) );
NAND2_X2 \add_506/U621  ( .A1(\add_506/n398 ), .A2(\add_506/n440 ), .ZN(\add_506/n439 ) );
NAND4_X2 \add_506/U620  ( .A1(n18129), .A2(n18133), .A3(n18145), .A4(n18149),.ZN(\add_506/n437 ) );
NAND2_X2 \add_506/U619  ( .A1(n18137), .A2(n18141), .ZN(\add_506/n438 ) );
NOR2_X2 \add_506/U618  ( .A1(\add_506/n437 ), .A2(\add_506/n438 ), .ZN(\add_506/n435 ) );
NAND2_X2 \add_506/U617  ( .A1(\add_506/n435 ), .A2(\add_506/n436 ), .ZN(\add_506/n433 ) );
NAND2_X2 \add_506/U616  ( .A1(\add_506/n27 ), .A2(\add_506/n432 ), .ZN(\add_506/n431 ) );
NAND2_X2 \add_506/U615  ( .A1(\add_506/n429 ), .A2(\add_506/n430 ), .ZN(\add_506/n428 ) );
XNOR2_X2 \add_506/U614  ( .A(\add_506/n428 ), .B(n18097), .ZN(N2150) );
NAND2_X2 \add_506/U613  ( .A1(\add_506/n426 ), .A2(\add_506/n398 ), .ZN(\add_506/n425 ) );
NAND2_X2 \add_506/U612  ( .A1(n18101), .A2(n18097), .ZN(\add_506/n422 ) );
NAND4_X2 \add_506/U611  ( .A1(n18113), .A2(n18117), .A3(n18121), .A4(n18125),.ZN(\add_506/n423 ) );
NAND2_X2 \add_506/U610  ( .A1(n18105), .A2(n18109), .ZN(\add_506/n424 ) );
NAND2_X2 \add_506/U609  ( .A1(\add_506/n401 ), .A2(\add_506/n419 ), .ZN(\add_506/n418 ) );
NAND2_X2 \add_506/U608  ( .A1(\add_506/n416 ), .A2(\add_506/n417 ), .ZN(\add_506/n415 ) );
XNOR2_X2 \add_506/U607  ( .A(\add_506/n415 ), .B(n18093), .ZN(N2151) );
INV_X4 \add_506/U606  ( .A(\add_506/n401 ), .ZN(\add_506/n412 ) );
NAND4_X2 \add_506/U605  ( .A1(n18137), .A2(n18141), .A3(n18145), .A4(n18149),.ZN(\add_506/n413 ) );
NAND4_X2 \add_506/U604  ( .A1(\add_506/n409 ), .A2(\add_506/n22 ), .A3(\add_506/n26 ), .A4(\add_506/n410 ), .ZN(\add_506/n408 ) );
XNOR2_X2 \add_506/U603  ( .A(\add_506/n408 ), .B(n18089), .ZN(N2152) );
NAND4_X2 \add_506/U602  ( .A1(n18133), .A2(n18137), .A3(n18141), .A4(n18145),.ZN(\add_506/n406 ) );
NAND4_X2 \add_506/U601  ( .A1(n18149), .A2(n18153), .A3(n18157), .A4(\add_506/n398 ), .ZN(\add_506/n405 ) );
NAND4_X2 \add_506/U600  ( .A1(\add_506/n403 ), .A2(\add_506/n19 ), .A3(\add_506/n26 ), .A4(\add_506/n404 ), .ZN(\add_506/n402 ) );
XNOR2_X2 \add_506/U599  ( .A(\add_506/n402 ), .B(n18082), .ZN(N2153) );
NAND4_X2 \add_506/U598  ( .A1(n18133), .A2(n18137), .A3(n18141), .A4(n18145),.ZN(\add_506/n399 ) );
NAND4_X2 \add_506/U597  ( .A1(n18082), .A2(n18089), .A3(n18093), .A4(n18129),.ZN(\add_506/n400 ) );
NAND4_X2 \add_506/U596  ( .A1(n18149), .A2(n18153), .A3(n18157), .A4(\add_506/n398 ), .ZN(\add_506/n397 ) );
NAND4_X2 \add_506/U595  ( .A1(\add_506/n395 ), .A2(\add_506/n21 ), .A3(\add_506/n26 ), .A4(\add_506/n396 ), .ZN(\add_506/n394 ) );
XNOR2_X2 \add_506/U594  ( .A(\add_506/n394 ), .B(n18593), .ZN(N2154) );
NAND2_X2 \add_506/U593  ( .A1(\add_506/n2 ), .A2(\add_506/n30 ), .ZN(\add_506/n393 ) );
XNOR2_X2 \add_506/U592  ( .A(\add_506/n393 ), .B(n18541), .ZN(N2039) );
XNOR2_X2 \add_506/U591  ( .A(\add_506/n392 ), .B(n18537), .ZN(N2040) );
NAND2_X2 \add_506/U590  ( .A1(\add_506/n30 ), .A2(\add_506/n389 ), .ZN(\add_506/n388 ) );
XNOR2_X2 \add_506/U589  ( .A(\add_506/n388 ), .B(n18533), .ZN(N2041) );
NAND4_X2 \add_506/U588  ( .A1(n18533), .A2(n18537), .A3(n18541), .A4(n18545),.ZN(\add_506/n387 ) );
NAND2_X2 \add_506/U587  ( .A1(\add_506/n30 ), .A2(\add_506/n385 ), .ZN(\add_506/n384 ) );
XNOR2_X2 \add_506/U586  ( .A(\add_506/n384 ), .B(n18529), .ZN(N2042) );
NAND2_X2 \add_506/U585  ( .A1(n18537), .A2(n18541), .ZN(\add_506/n382 ) );
NAND2_X2 \add_506/U584  ( .A1(n18529), .A2(n18533), .ZN(\add_506/n383 ) );
NAND2_X2 \add_506/U583  ( .A1(n18553), .A2(n18557), .ZN(\add_506/n380 ) );
NAND2_X2 \add_506/U582  ( .A1(n18545), .A2(n18549), .ZN(\add_506/n381 ) );
NAND4_X2 \add_506/U581  ( .A1(n18577), .A2(n18581), .A3(n18585), .A4(n18589),.ZN(\add_506/n378 ) );
NAND4_X2 \add_506/U580  ( .A1(n18561), .A2(n18565), .A3(n18569), .A4(n18573),.ZN(\add_506/n379 ) );
XNOR2_X2 \add_506/U579  ( .A(\add_506/n374 ), .B(n18525), .ZN(N2043) );
NAND2_X2 \add_506/U578  ( .A1(\add_506/n337 ), .A2(n18525), .ZN(\add_506/n373 ) );
XNOR2_X2 \add_506/U577  ( .A(\add_506/n373 ), .B(n18521), .ZN(N2044) );
XNOR2_X2 \add_506/U576  ( .A(\add_506/n372 ), .B(n18517), .ZN(N2045) );
NAND4_X2 \add_506/U575  ( .A1(n18521), .A2(n18517), .A3(n18525), .A4(\add_506/n337 ), .ZN(\add_506/n371 ) );
XNOR2_X2 \add_506/U574  ( .A(\add_506/n371 ), .B(n18513), .ZN(N2046) );
NAND2_X2 \add_506/U573  ( .A1(\add_506/n337 ), .A2(\add_506/n362 ), .ZN(\add_506/n370 ) );
XNOR2_X2 \add_506/U572  ( .A(\add_506/n370 ), .B(n18509), .ZN(N2047) );
XNOR2_X2 \add_506/U571  ( .A(\add_506/n369 ), .B(n18505), .ZN(N2048) );
NAND4_X2 \add_506/U570  ( .A1(n18505), .A2(n18509), .A3(\add_506/n362 ),.A4(\add_506/n337 ), .ZN(\add_506/n368 ) );
XNOR2_X2 \add_506/U569  ( .A(\add_506/n368 ), .B(n18501), .ZN(N2049) );
NAND2_X2 \add_506/U568  ( .A1(\add_506/n366 ), .A2(\add_506/n337 ), .ZN(\add_506/n365 ) );
XNOR2_X2 \add_506/U567  ( .A(\add_506/n365 ), .B(n18497), .ZN(N2050) );
NAND4_X2 \add_506/U566  ( .A1(n18497), .A2(n18501), .A3(n18505), .A4(n18509),.ZN(\add_506/n339 ) );
NAND2_X2 \add_506/U565  ( .A1(\add_506/n364 ), .A2(\add_506/n337 ), .ZN(\add_506/n363 ) );
XNOR2_X2 \add_506/U564  ( .A(\add_506/n363 ), .B(n18493), .ZN(N2051) );
INV_X4 \add_506/U563  ( .A(\add_506/n339 ), .ZN(\add_506/n361 ) );
INV_X4 \add_506/U562  ( .A(\add_506/n607 ), .ZN(\add_506/n362 ) );
NAND4_X2 \add_506/U561  ( .A1(\add_506/n361 ), .A2(\add_506/n362 ), .A3(n18493), .A4(\add_506/n337 ), .ZN(\add_506/n360 ) );
XNOR2_X2 \add_506/U560  ( .A(\add_506/n360 ), .B(n18489), .ZN(N2052) );
NAND4_X2 \add_506/U559  ( .A1(n18489), .A2(n18493), .A3(\add_506/n359 ),.A4(\add_506/n337 ), .ZN(\add_506/n358 ) );
XNOR2_X2 \add_506/U558  ( .A(\add_506/n358 ), .B(n18485), .ZN(N2053) );
NAND2_X2 \add_506/U557  ( .A1(\add_506/n356 ), .A2(\add_506/n337 ), .ZN(\add_506/n355 ) );
XNOR2_X2 \add_506/U556  ( .A(\add_506/n355 ), .B(n18481), .ZN(N2054) );
NAND4_X2 \add_506/U555  ( .A1(n18481), .A2(n18485), .A3(n18489), .A4(n18493),.ZN(\add_506/n352 ) );
NAND2_X2 \add_506/U554  ( .A1(\add_506/n354 ), .A2(\add_506/n337 ), .ZN(\add_506/n353 ) );
XNOR2_X2 \add_506/U553  ( .A(\add_506/n353 ), .B(n18477), .ZN(N2055) );
INV_X4 \add_506/U552  ( .A(\add_506/n352 ), .ZN(\add_506/n341 ) );
NAND2_X2 \add_506/U551  ( .A1(\add_506/n341 ), .A2(n18477), .ZN(\add_506/n351 ) );
NAND2_X2 \add_506/U550  ( .A1(\add_506/n350 ), .A2(\add_506/n337 ), .ZN(\add_506/n349 ) );
XNOR2_X2 \add_506/U549  ( .A(\add_506/n349 ), .B(n18473), .ZN(N2056) );
NAND2_X2 \add_506/U548  ( .A1(n18585), .A2(n18589), .ZN(\add_506/n304 ) );
XNOR2_X2 \add_506/U547  ( .A(\add_506/n304 ), .B(n18581), .ZN(N2029) );
INV_X4 \add_506/U546  ( .A(n18477), .ZN(\add_506/n342 ) );
INV_X4 \add_506/U545  ( .A(n18473), .ZN(\add_506/n348 ) );
NAND2_X2 \add_506/U544  ( .A1(\add_506/n347 ), .A2(\add_506/n341 ), .ZN(\add_506/n346 ) );
NAND2_X2 \add_506/U543  ( .A1(\add_506/n345 ), .A2(\add_506/n337 ), .ZN(\add_506/n344 ) );
XNOR2_X2 \add_506/U542  ( .A(\add_506/n344 ), .B(n18469), .ZN(N2057) );
NAND2_X2 \add_506/U541  ( .A1(n18473), .A2(n18469), .ZN(\add_506/n343 ) );
NAND2_X2 \add_506/U540  ( .A1(\add_506/n340 ), .A2(\add_506/n341 ), .ZN(\add_506/n338 ) );
NAND2_X2 \add_506/U539  ( .A1(\add_506/n336 ), .A2(\add_506/n337 ), .ZN(\add_506/n335 ) );
XNOR2_X2 \add_506/U538  ( .A(\add_506/n335 ), .B(n18465), .ZN(N2058) );
NAND2_X2 \add_506/U537  ( .A1(n18505), .A2(n18509), .ZN(\add_506/n333 ) );
NAND2_X2 \add_506/U536  ( .A1(n18497), .A2(n18501), .ZN(\add_506/n334 ) );
NAND2_X2 \add_506/U535  ( .A1(n18521), .A2(n18525), .ZN(\add_506/n331 ) );
NAND2_X2 \add_506/U534  ( .A1(n18513), .A2(n18517), .ZN(\add_506/n332 ) );
NAND2_X2 \add_506/U533  ( .A1(\add_506/n329 ), .A2(\add_506/n330 ), .ZN(\add_506/n326 ) );
NAND4_X2 \add_506/U532  ( .A1(n18481), .A2(n18485), .A3(n18489), .A4(n18493),.ZN(\add_506/n327 ) );
NAND4_X2 \add_506/U531  ( .A1(n18465), .A2(n18469), .A3(n18473), .A4(n18477),.ZN(\add_506/n328 ) );
NAND2_X2 \add_506/U530  ( .A1(n18569), .A2(n18573), .ZN(\add_506/n324 ) );
NAND2_X2 \add_506/U529  ( .A1(n18561), .A2(n18565), .ZN(\add_506/n325 ) );
NAND2_X2 \add_506/U528  ( .A1(n18585), .A2(n18589), .ZN(\add_506/n322 ) );
NAND2_X2 \add_506/U527  ( .A1(n18577), .A2(n18581), .ZN(\add_506/n323 ) );
NAND2_X2 \add_506/U526  ( .A1(\add_506/n320 ), .A2(\add_506/n321 ), .ZN(\add_506/n317 ) );
NAND4_X2 \add_506/U525  ( .A1(n18545), .A2(n18549), .A3(n18553), .A4(n18557),.ZN(\add_506/n318 ) );
NAND4_X2 \add_506/U524  ( .A1(n18529), .A2(n18533), .A3(n18537), .A4(n18541),.ZN(\add_506/n319 ) );
NAND2_X2 \add_506/U523  ( .A1(\add_506/n315 ), .A2(\add_506/n316 ), .ZN(\add_506/n314 ) );
XNOR2_X2 \add_506/U522  ( .A(\add_506/n314 ), .B(n18461), .ZN(N2059) );
NAND2_X2 \add_506/U521  ( .A1(\add_506/n17 ), .A2(n18461), .ZN(\add_506/n313 ) );
XNOR2_X2 \add_506/U520  ( .A(\add_506/n313 ), .B(n18457), .ZN(N2060) );
XNOR2_X2 \add_506/U519  ( .A(\add_506/n312 ), .B(n18453), .ZN(N2061) );
NAND4_X2 \add_506/U518  ( .A1(n18457), .A2(n18453), .A3(n18461), .A4(\add_506/n15 ), .ZN(\add_506/n311 ) );
XNOR2_X2 \add_506/U517  ( .A(\add_506/n311 ), .B(n18449), .ZN(N2062) );
NAND2_X2 \add_506/U516  ( .A1(\add_506/n267 ), .A2(\add_506/n18 ), .ZN(\add_506/n310 ) );
XNOR2_X2 \add_506/U515  ( .A(\add_506/n310 ), .B(n18445), .ZN(N2063) );
INV_X4 \add_506/U514  ( .A(n18445), .ZN(\add_506/n280 ) );
NAND2_X2 \add_506/U513  ( .A1(\add_506/n309 ), .A2(\add_506/n18 ), .ZN(\add_506/n308 ) );
XNOR2_X2 \add_506/U512  ( .A(\add_506/n308 ), .B(n18441), .ZN(N2064) );
NAND4_X2 \add_506/U511  ( .A1(n18445), .A2(\add_506/n267 ), .A3(n18441),.A4(\add_506/n15 ), .ZN(\add_506/n307 ) );
XNOR2_X2 \add_506/U510  ( .A(\add_506/n307 ), .B(n18437), .ZN(N2065) );
NAND4_X2 \add_506/U509  ( .A1(n18441), .A2(n18437), .A3(\add_506/n306 ),.A4(\add_506/n15 ), .ZN(\add_506/n305 ) );
XNOR2_X2 \add_506/U508  ( .A(\add_506/n305 ), .B(n18433), .ZN(N2066) );
INV_X4 \add_506/U507  ( .A(\add_506/n304 ), .ZN(\add_506/n303 ) );
NAND2_X2 \add_506/U506  ( .A1(n18581), .A2(\add_506/n303 ), .ZN(\add_506/n302 ) );
XNOR2_X2 \add_506/U505  ( .A(\add_506/n302 ), .B(n18577), .ZN(N2030) );
NAND4_X2 \add_506/U504  ( .A1(n18433), .A2(n18437), .A3(n18441), .A4(n18445),.ZN(\add_506/n288 ) );
NAND2_X2 \add_506/U503  ( .A1(\add_506/n301 ), .A2(\add_506/n18 ), .ZN(\add_506/n300 ) );
XNOR2_X2 \add_506/U502  ( .A(\add_506/n300 ), .B(n18429), .ZN(N2067) );
INV_X4 \add_506/U501  ( .A(\add_506/n288 ), .ZN(\add_506/n299 ) );
NAND4_X2 \add_506/U500  ( .A1(n18429), .A2(\add_506/n267 ), .A3(\add_506/n299 ), .A4(\add_506/n15 ), .ZN(\add_506/n298 ) );
XNOR2_X2 \add_506/U499  ( .A(\add_506/n298 ), .B(n18425), .ZN(N2068) );
NAND2_X2 \add_506/U498  ( .A1(n18425), .A2(n18429), .ZN(\add_506/n297 ) );
NAND2_X2 \add_506/U497  ( .A1(\add_506/n17 ), .A2(\add_506/n296 ), .ZN(\add_506/n295 ) );
XNOR2_X2 \add_506/U496  ( .A(\add_506/n295 ), .B(n18421), .ZN(N2069) );
NAND2_X2 \add_506/U495  ( .A1(\add_506/n293 ), .A2(\add_506/n18 ), .ZN(\add_506/n292 ) );
XNOR2_X2 \add_506/U494  ( .A(\add_506/n292 ), .B(n18417), .ZN(N2070) );
NAND4_X2 \add_506/U493  ( .A1(n18417), .A2(n18421), .A3(n18425), .A4(n18429),.ZN(\add_506/n291 ) );
NAND2_X2 \add_506/U492  ( .A1(\add_506/n290 ), .A2(\add_506/n18 ), .ZN(\add_506/n289 ) );
XNOR2_X2 \add_506/U491  ( .A(\add_506/n289 ), .B(n18413), .ZN(N2071) );
NAND2_X2 \add_506/U490  ( .A1(\add_506/n299 ), .A2(n18413), .ZN(\add_506/n286 ) );
NAND4_X2 \add_506/U489  ( .A1(n18417), .A2(n18421), .A3(n18425), .A4(n18429),.ZN(\add_506/n287 ) );
NAND2_X2 \add_506/U488  ( .A1(\add_506/n285 ), .A2(\add_506/n18 ), .ZN(\add_506/n284 ) );
XNOR2_X2 \add_506/U487  ( .A(\add_506/n284 ), .B(n18409), .ZN(N2072) );
INV_X4 \add_506/U486  ( .A(n18429), .ZN(\add_506/n282 ) );
NAND2_X2 \add_506/U485  ( .A1(n18425), .A2(n18433), .ZN(\add_506/n283 ) );
NAND2_X2 \add_506/U484  ( .A1(n18441), .A2(n18437), .ZN(\add_506/n281 ) );
NAND2_X2 \add_506/U483  ( .A1(\add_506/n278 ), .A2(\add_506/n279 ), .ZN(\add_506/n276 ) );
NAND4_X2 \add_506/U482  ( .A1(n18409), .A2(n18421), .A3(n18417), .A4(n18413),.ZN(\add_506/n277 ) );
NAND2_X2 \add_506/U481  ( .A1(\add_506/n275 ), .A2(\add_506/n17 ), .ZN(\add_506/n274 ) );
XNOR2_X2 \add_506/U480  ( .A(\add_506/n274 ), .B(n18405), .ZN(N2073) );
INV_X4 \add_506/U479  ( .A(\add_506/n621 ), .ZN(\add_506/n267 ) );
NAND4_X2 \add_506/U478  ( .A1(n18433), .A2(n18437), .A3(n18441), .A4(n18445),.ZN(\add_506/n272 ) );
NAND2_X2 \add_506/U477  ( .A1(n18413), .A2(n18409), .ZN(\add_506/n270 ) );
NAND2_X2 \add_506/U476  ( .A1(n18405), .A2(n18417), .ZN(\add_506/n271 ) );
NAND4_X2 \add_506/U475  ( .A1(\add_506/n267 ), .A2(\add_506/n268 ), .A3(\add_506/n269 ), .A4(\add_506/n16 ), .ZN(\add_506/n266 ) );
XNOR2_X2 \add_506/U474  ( .A(\add_506/n266 ), .B(n18401), .ZN(N2074) );
NAND2_X2 \add_506/U473  ( .A1(\add_506/n27 ), .A2(\add_506/n17 ), .ZN(\add_506/n265 ) );
XNOR2_X2 \add_506/U472  ( .A(\add_506/n265 ), .B(n18397), .ZN(N2075) );
INV_X4 \add_506/U471  ( .A(n18397), .ZN(\add_506/n234 ) );
NAND2_X2 \add_506/U470  ( .A1(\add_506/n264 ), .A2(\add_506/n18 ), .ZN(\add_506/n263 ) );
XNOR2_X2 \add_506/U469  ( .A(\add_506/n263 ), .B(n18393), .ZN(N2076) );
INV_X4 \add_506/U468  ( .A(n18573), .ZN(\add_506/n262 ) );
XNOR2_X2 \add_506/U467  ( .A(\add_506/n262 ), .B(\add_506/n4 ), .ZN(N2031));
NAND4_X2 \add_506/U466  ( .A1(n18397), .A2(\add_506/n27 ), .A3(n18393), .A4(\add_506/n16 ), .ZN(\add_506/n261 ) );
XNOR2_X2 \add_506/U465  ( .A(\add_506/n261 ), .B(n18389), .ZN(N2077) );
NAND4_X2 \add_506/U464  ( .A1(n18393), .A2(n18389), .A3(\add_506/n260 ),.A4(\add_506/n16 ), .ZN(\add_506/n259 ) );
XNOR2_X2 \add_506/U463  ( .A(\add_506/n259 ), .B(n18385), .ZN(N2078) );
NAND4_X2 \add_506/U462  ( .A1(n18385), .A2(n18389), .A3(n18393), .A4(n18397),.ZN(\add_506/n244 ) );
NAND2_X2 \add_506/U461  ( .A1(\add_506/n258 ), .A2(\add_506/n17 ), .ZN(\add_506/n257 ) );
XNOR2_X2 \add_506/U460  ( .A(\add_506/n257 ), .B(n18381), .ZN(N2079) );
INV_X4 \add_506/U459  ( .A(\add_506/n244 ), .ZN(\add_506/n247 ) );
NAND4_X2 \add_506/U458  ( .A1(\add_506/n247 ), .A2(n18381), .A3(\add_506/n26 ), .A4(\add_506/n16 ), .ZN(\add_506/n256 ) );
XNOR2_X2 \add_506/U457  ( .A(\add_506/n256 ), .B(n18377), .ZN(N2080) );
NAND2_X2 \add_506/U456  ( .A1(n18377), .A2(n18381), .ZN(\add_506/n255 ) );
NAND2_X2 \add_506/U455  ( .A1(\add_506/n17 ), .A2(\add_506/n254 ), .ZN(\add_506/n253 ) );
XNOR2_X2 \add_506/U454  ( .A(\add_506/n253 ), .B(n18373), .ZN(N2081) );
INV_X4 \add_506/U453  ( .A(n18381), .ZN(\add_506/n236 ) );
NAND2_X2 \add_506/U452  ( .A1(n18377), .A2(n18373), .ZN(\add_506/n252 ) );
NAND4_X2 \add_506/U451  ( .A1(\add_506/n251 ), .A2(\add_506/n247 ), .A3(\add_506/n26 ), .A4(\add_506/n16 ), .ZN(\add_506/n250 ) );
XNOR2_X2 \add_506/U450  ( .A(\add_506/n250 ), .B(n18369), .ZN(N2082) );
NAND2_X2 \add_506/U449  ( .A1(n18377), .A2(n18381), .ZN(\add_506/n248 ) );
NAND2_X2 \add_506/U448  ( .A1(n18369), .A2(n18373), .ZN(\add_506/n249 ) );
NAND4_X2 \add_506/U447  ( .A1(\add_506/n246 ), .A2(\add_506/n247 ), .A3(\add_506/n26 ), .A4(\add_506/n16 ), .ZN(\add_506/n245 ) );
XNOR2_X2 \add_506/U446  ( .A(\add_506/n245 ), .B(n18365), .ZN(N2083) );
INV_X4 \add_506/U445  ( .A(n18365), .ZN(\add_506/n243 ) );
NAND2_X2 \add_506/U444  ( .A1(n18377), .A2(n18381), .ZN(\add_506/n241 ) );
NAND2_X2 \add_506/U443  ( .A1(n18373), .A2(n18369), .ZN(\add_506/n242 ) );
NAND4_X2 \add_506/U442  ( .A1(\add_506/n239 ), .A2(\add_506/n240 ), .A3(\add_506/n26 ), .A4(\add_506/n16 ), .ZN(\add_506/n238 ) );
XNOR2_X2 \add_506/U441  ( .A(\add_506/n238 ), .B(n18361), .ZN(N2084) );
NAND2_X2 \add_506/U440  ( .A1(n18377), .A2(n18385), .ZN(\add_506/n237 ) );
NAND2_X2 \add_506/U439  ( .A1(n18393), .A2(n18389), .ZN(\add_506/n235 ) );
NAND2_X2 \add_506/U438  ( .A1(\add_506/n232 ), .A2(\add_506/n233 ), .ZN(\add_506/n230 ) );
NAND4_X2 \add_506/U437  ( .A1(n18361), .A2(n18373), .A3(n18369), .A4(n18365),.ZN(\add_506/n231 ) );
NAND2_X2 \add_506/U436  ( .A1(\add_506/n229 ), .A2(\add_506/n18 ), .ZN(\add_506/n228 ) );
XNOR2_X2 \add_506/U435  ( .A(\add_506/n228 ), .B(n18357), .ZN(N2085) );
NAND4_X2 \add_506/U434  ( .A1(n18385), .A2(n18389), .A3(n18393), .A4(n18397),.ZN(\add_506/n226 ) );
NAND2_X2 \add_506/U433  ( .A1(n18365), .A2(n18361), .ZN(\add_506/n224 ) );
NAND2_X2 \add_506/U432  ( .A1(n18357), .A2(n18369), .ZN(\add_506/n225 ) );
NAND4_X2 \add_506/U431  ( .A1(\add_506/n222 ), .A2(\add_506/n27 ), .A3(\add_506/n223 ), .A4(\add_506/n16 ), .ZN(\add_506/n221 ) );
XNOR2_X2 \add_506/U430  ( .A(\add_506/n221 ), .B(n18353), .ZN(N2086) );
NAND2_X2 \add_506/U429  ( .A1(\add_506/n4 ), .A2(n18573), .ZN(\add_506/n220 ) );
XNOR2_X2 \add_506/U428  ( .A(\add_506/n220 ), .B(n18569), .ZN(N2032) );
NAND2_X2 \add_506/U427  ( .A1(\add_506/n213 ), .A2(\add_506/n18 ), .ZN(\add_506/n212 ) );
XNOR2_X2 \add_506/U426  ( .A(\add_506/n212 ), .B(n18349), .ZN(N2087) );
INV_X4 \add_506/U425  ( .A(\add_506/n135 ), .ZN(\add_506/n211 ) );
NAND4_X2 \add_506/U424  ( .A1(\add_506/n211 ), .A2(\add_506/n27 ), .A3(n18349), .A4(\add_506/n15 ), .ZN(\add_506/n210 ) );
XNOR2_X2 \add_506/U423  ( .A(\add_506/n210 ), .B(n18345), .ZN(N2088) );
NAND2_X2 \add_506/U422  ( .A1(n18345), .A2(n18349), .ZN(\add_506/n209 ) );
NAND2_X2 \add_506/U421  ( .A1(\add_506/n17 ), .A2(\add_506/n208 ), .ZN(\add_506/n207 ) );
XNOR2_X2 \add_506/U420  ( .A(\add_506/n207 ), .B(n18341), .ZN(N2089) );
NAND2_X2 \add_506/U419  ( .A1(\add_506/n205 ), .A2(\add_506/n18 ), .ZN(\add_506/n204 ) );
XNOR2_X2 \add_506/U418  ( .A(\add_506/n204 ), .B(n18337), .ZN(N2090) );
NAND4_X2 \add_506/U417  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(\add_506/n199 ) );
NAND2_X2 \add_506/U416  ( .A1(\add_506/n17 ), .A2(\add_506/n203 ), .ZN(\add_506/n202 ) );
XNOR2_X2 \add_506/U415  ( .A(\add_506/n202 ), .B(n18333), .ZN(N2091) );
NAND4_X2 \add_506/U414  ( .A1(\add_506/n201 ), .A2(\add_506/n17 ), .A3(\add_506/n26 ), .A4(n18333), .ZN(\add_506/n200 ) );
XNOR2_X2 \add_506/U413  ( .A(\add_506/n200 ), .B(n18329), .ZN(N2092) );
NAND3_X2 \add_506/U412  ( .A1(\add_506/n197 ), .A2(\add_506/n17 ), .A3(\add_506/n198 ), .ZN(\add_506/n196 ) );
XNOR2_X2 \add_506/U411  ( .A(\add_506/n196 ), .B(n18325), .ZN(N2093) );
NAND2_X2 \add_506/U410  ( .A1(n18345), .A2(n18341), .ZN(\add_506/n195 ) );
INV_X4 \add_506/U409  ( .A(n18325), .ZN(\add_506/n187 ) );
NAND4_X2 \add_506/U408  ( .A1(\add_506/n16 ), .A2(\add_506/n192 ), .A3(\add_506/n26 ), .A4(\add_506/n193 ), .ZN(\add_506/n191 ) );
XNOR2_X2 \add_506/U407  ( .A(\add_506/n191 ), .B(n18321), .ZN(N2094) );
INV_X4 \add_506/U406  ( .A(n18321), .ZN(\add_506/n188 ) );
NAND4_X2 \add_506/U405  ( .A1(\add_506/n16 ), .A2(\add_506/n185 ), .A3(\add_506/n26 ), .A4(\add_506/n186 ), .ZN(\add_506/n184 ) );
XNOR2_X2 \add_506/U404  ( .A(\add_506/n184 ), .B(n18317), .ZN(N2095) );
NAND3_X2 \add_506/U403  ( .A1(\add_506/n179 ), .A2(\add_506/n17 ), .A3(\add_506/n180 ), .ZN(\add_506/n178 ) );
XNOR2_X2 \add_506/U402  ( .A(\add_506/n178 ), .B(n18313), .ZN(N2096) );
XNOR2_X2 \add_506/U401  ( .A(\add_506/n177 ), .B(n18565), .ZN(N2033) );
NAND4_X2 \add_506/U400  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(\add_506/n175 ) );
NAND3_X2 \add_506/U399  ( .A1(\add_506/n172 ), .A2(\add_506/n17 ), .A3(\add_506/n173 ), .ZN(\add_506/n171 ) );
XNOR2_X2 \add_506/U398  ( .A(\add_506/n171 ), .B(n18309), .ZN(N2097) );
NAND4_X2 \add_506/U397  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(\add_506/n169 ) );
NAND4_X2 \add_506/U396  ( .A1(n18309), .A2(n18313), .A3(n18317), .A4(n18321),.ZN(\add_506/n168 ) );
NAND3_X2 \add_506/U395  ( .A1(\add_506/n166 ), .A2(\add_506/n17 ), .A3(\add_506/n167 ), .ZN(\add_506/n165 ) );
XNOR2_X2 \add_506/U394  ( .A(\add_506/n165 ), .B(n18305), .ZN(N2098) );
NAND4_X2 \add_506/U393  ( .A1(n18337), .A2(n18341), .A3(n18345), .A4(n18349),.ZN(\add_506/n163 ) );
NAND4_X2 \add_506/U392  ( .A1(n18321), .A2(n18325), .A3(n18329), .A4(n18333),.ZN(\add_506/n164 ) );
NAND4_X2 \add_506/U391  ( .A1(n18305), .A2(n18309), .A3(n18313), .A4(n18317),.ZN(\add_506/n162 ) );
NAND3_X2 \add_506/U390  ( .A1(\add_506/n160 ), .A2(\add_506/n17 ), .A3(\add_506/n161 ), .ZN(\add_506/n159 ) );
XNOR2_X2 \add_506/U389  ( .A(\add_506/n159 ), .B(n18301), .ZN(N2099) );
NAND2_X2 \add_506/U388  ( .A1(n18329), .A2(n18333), .ZN(\add_506/n157 ) );
NAND2_X2 \add_506/U387  ( .A1(n18321), .A2(n18325), .ZN(\add_506/n158 ) );
NAND2_X2 \add_506/U386  ( .A1(n18345), .A2(n18349), .ZN(\add_506/n155 ) );
NAND2_X2 \add_506/U385  ( .A1(n18337), .A2(n18341), .ZN(\add_506/n156 ) );
INV_X4 \add_506/U384  ( .A(n18301), .ZN(\add_506/n154 ) );
NAND4_X2 \add_506/U383  ( .A1(\add_506/n151 ), .A2(\add_506/n152 ), .A3(\add_506/n26 ), .A4(\add_506/n153 ), .ZN(\add_506/n149 ) );
NAND4_X2 \add_506/U382  ( .A1(n18305), .A2(n18309), .A3(n18313), .A4(n18317),.ZN(\add_506/n150 ) );
NAND2_X2 \add_506/U381  ( .A1(n18341), .A2(n18345), .ZN(\add_506/n146 ) );
NAND4_X2 \add_506/U380  ( .A1(n18317), .A2(n18321), .A3(n18325), .A4(n18329),.ZN(\add_506/n148 ) );
INV_X4 \add_506/U379  ( .A(n18297), .ZN(\add_506/n145 ) );
NAND4_X2 \add_506/U378  ( .A1(n18301), .A2(n18305), .A3(n18309), .A4(n18313),.ZN(\add_506/n144 ) );
NAND4_X2 \add_506/U377  ( .A1(\add_506/n141 ), .A2(\add_506/n27 ), .A3(\add_506/n142 ), .A4(\add_506/n143 ), .ZN(\add_506/n140 ) );
XNOR2_X2 \add_506/U376  ( .A(\add_506/n140 ), .B(n18293), .ZN(N2101) );
NAND2_X2 \add_506/U375  ( .A1(n18345), .A2(n18341), .ZN(\add_506/n137 ) );
NAND4_X2 \add_506/U374  ( .A1(n18317), .A2(n18321), .A3(n18325), .A4(n18329),.ZN(\add_506/n139 ) );
INV_X4 \add_506/U373  ( .A(n18293), .ZN(\add_506/n136 ) );
NAND2_X2 \add_506/U372  ( .A1(n18309), .A2(n18305), .ZN(\add_506/n134 ) );
NAND4_X2 \add_506/U371  ( .A1(\add_506/n130 ), .A2(\add_506/n27 ), .A3(\add_506/n131 ), .A4(\add_506/n132 ), .ZN(\add_506/n129 ) );
XNOR2_X2 \add_506/U370  ( .A(\add_506/n129 ), .B(n18289), .ZN(N2102) );
NAND3_X2 \add_506/U369  ( .A1(\add_506/n21 ), .A2(\add_506/n27 ), .A3(\add_506/n17 ), .ZN(\add_506/n128 ) );
XNOR2_X2 \add_506/U368  ( .A(\add_506/n128 ), .B(n18285), .ZN(N2103) );
NAND4_X2 \add_506/U367  ( .A1(\add_506/n26 ), .A2(\add_506/n20 ), .A3(\add_506/n16 ), .A4(n18285), .ZN(\add_506/n127 ) );
XNOR2_X2 \add_506/U366  ( .A(\add_506/n127 ), .B(n18281), .ZN(N2104) );
INV_X4 \add_506/U365  ( .A(n18285), .ZN(\add_506/n122 ) );
INV_X4 \add_506/U364  ( .A(n18281), .ZN(\add_506/n126 ) );
NAND4_X2 \add_506/U363  ( .A1(\add_506/n27 ), .A2(\add_506/n20 ), .A3(\add_506/n125 ), .A4(\add_506/n15 ), .ZN(\add_506/n124 ) );
XNOR2_X2 \add_506/U362  ( .A(\add_506/n124 ), .B(n18277), .ZN(N2105) );
NAND2_X2 \add_506/U361  ( .A1(n18281), .A2(n18277), .ZN(\add_506/n123 ) );
NAND4_X2 \add_506/U360  ( .A1(\add_506/n121 ), .A2(\add_506/n16 ), .A3(\add_506/n19 ), .A4(\add_506/n26 ), .ZN(\add_506/n120 ) );
XNOR2_X2 \add_506/U359  ( .A(\add_506/n120 ), .B(n18273), .ZN(N2106) );
NAND4_X2 \add_506/U358  ( .A1(n18569), .A2(n18565), .A3(n18573), .A4(\add_506/n4 ), .ZN(\add_506/n119 ) );
XNOR2_X2 \add_506/U357  ( .A(\add_506/n119 ), .B(n18561), .ZN(N2034) );
NAND4_X2 \add_506/U356  ( .A1(n18273), .A2(n18277), .A3(n18281), .A4(n18285),.ZN(\add_506/n114 ) );
NAND3_X2 \add_506/U355  ( .A1(\add_506/n21 ), .A2(\add_506/n118 ), .A3(\add_506/n17 ), .ZN(\add_506/n117 ) );
XNOR2_X2 \add_506/U354  ( .A(\add_506/n117 ), .B(n18269), .ZN(N2107) );
NAND4_X2 \add_506/U353  ( .A1(\add_506/n20 ), .A2(n18269), .A3(\add_506/n116 ), .A4(\add_506/n16 ), .ZN(\add_506/n115 ) );
XNOR2_X2 \add_506/U352  ( .A(\add_506/n115 ), .B(n18265), .ZN(N2108) );
INV_X4 \add_506/U351  ( .A(n18269), .ZN(\add_506/n102 ) );
INV_X4 \add_506/U350  ( .A(n18265), .ZN(\add_506/n103 ) );
NAND4_X2 \add_506/U349  ( .A1(\add_506/n112 ), .A2(\add_506/n20 ), .A3(\add_506/n113 ), .A4(\add_506/n15 ), .ZN(\add_506/n111 ) );
XNOR2_X2 \add_506/U348  ( .A(\add_506/n111 ), .B(n18261), .ZN(N2109) );
NAND2_X2 \add_506/U347  ( .A1(n18281), .A2(n18277), .ZN(\add_506/n110 ) );
INV_X4 \add_506/U346  ( .A(n18261), .ZN(\add_506/n104 ) );
NAND4_X2 \add_506/U345  ( .A1(\add_506/n107 ), .A2(\add_506/n21 ), .A3(\add_506/n108 ), .A4(\add_506/n16 ), .ZN(\add_506/n106 ) );
XNOR2_X2 \add_506/U344  ( .A(\add_506/n106 ), .B(n18257), .ZN(N2110) );
INV_X4 \add_506/U343  ( .A(n18257), .ZN(\add_506/n105 ) );
NAND2_X2 \add_506/U342  ( .A1(n18281), .A2(n18285), .ZN(\add_506/n100 ) );
NAND2_X2 \add_506/U341  ( .A1(n18273), .A2(n18277), .ZN(\add_506/n101 ) );
NAND3_X2 \add_506/U340  ( .A1(\add_506/n21 ), .A2(\add_506/n96 ), .A3(\add_506/n17 ), .ZN(\add_506/n95 ) );
XNOR2_X2 \add_506/U339  ( .A(\add_506/n95 ), .B(n18253), .ZN(N2111) );
NAND4_X2 \add_506/U338  ( .A1(\add_506/n19 ), .A2(n18253), .A3(\add_506/n94 ), .A4(\add_506/n15 ), .ZN(\add_506/n93 ) );
XNOR2_X2 \add_506/U337  ( .A(\add_506/n93 ), .B(n18249), .ZN(N2112) );
INV_X4 \add_506/U336  ( .A(n18253), .ZN(\add_506/n87 ) );
INV_X4 \add_506/U335  ( .A(n18249), .ZN(\add_506/n92 ) );
NAND4_X2 \add_506/U334  ( .A1(\add_506/n90 ), .A2(\add_506/n21 ), .A3(\add_506/n91 ), .A4(\add_506/n15 ), .ZN(\add_506/n89 ) );
XNOR2_X2 \add_506/U333  ( .A(\add_506/n89 ), .B(n18245), .ZN(N2113) );
NAND2_X2 \add_506/U332  ( .A1(n18249), .A2(n18245), .ZN(\add_506/n88 ) );
NAND4_X2 \add_506/U331  ( .A1(\add_506/n85 ), .A2(\add_506/n21 ), .A3(\add_506/n86 ), .A4(\add_506/n15 ), .ZN(\add_506/n84 ) );
XNOR2_X2 \add_506/U330  ( .A(\add_506/n84 ), .B(n18241), .ZN(N2114) );
INV_X4 \add_506/U329  ( .A(\add_506/n75 ), .ZN(\add_506/n70 ) );
NAND4_X2 \add_506/U328  ( .A1(n18241), .A2(n18245), .A3(n18249), .A4(n18253),.ZN(\add_506/n76 ) );
INV_X4 \add_506/U327  ( .A(\add_506/n76 ), .ZN(\add_506/n71 ) );
AND2_X2 \add_506/U326  ( .A1(\add_506/n70 ), .A2(\add_506/n71 ), .ZN(\add_506/n83 ) );
NAND4_X2 \add_506/U325  ( .A1(\add_506/n19 ), .A2(\add_506/n27 ), .A3(\add_506/n83 ), .A4(\add_506/n15 ), .ZN(\add_506/n82 ) );
XNOR2_X2 \add_506/U324  ( .A(\add_506/n82 ), .B(n18237), .ZN(N2115) );
NAND2_X2 \add_506/U323  ( .A1(\add_506/n71 ), .A2(\add_506/n70 ), .ZN(\add_506/n81 ) );
NAND4_X2 \add_506/U322  ( .A1(\add_506/n19 ), .A2(n18237), .A3(\add_506/n80 ), .A4(\add_506/n15 ), .ZN(\add_506/n79 ) );
XNOR2_X2 \add_506/U321  ( .A(\add_506/n79 ), .B(n18233), .ZN(N2116) );
INV_X4 \add_506/U320  ( .A(n18557), .ZN(\add_506/n78 ) );
XNOR2_X2 \add_506/U319  ( .A(\add_506/n78 ), .B(\add_506/n30 ), .ZN(N2035));
INV_X4 \add_506/U318  ( .A(n18237), .ZN(\add_506/n67 ) );
INV_X4 \add_506/U317  ( .A(n18233), .ZN(\add_506/n77 ) );
NAND4_X2 \add_506/U316  ( .A1(\add_506/n19 ), .A2(\add_506/n73 ), .A3(\add_506/n74 ), .A4(\add_506/n15 ), .ZN(\add_506/n72 ) );
XNOR2_X2 \add_506/U315  ( .A(\add_506/n72 ), .B(n18229), .ZN(N2117) );
NAND2_X2 \add_506/U314  ( .A1(\add_506/n70 ), .A2(\add_506/n71 ), .ZN(\add_506/n69 ) );
NAND2_X2 \add_506/U313  ( .A1(n18233), .A2(n18229), .ZN(\add_506/n68 ) );
NAND4_X2 \add_506/U312  ( .A1(\add_506/n19 ), .A2(\add_506/n65 ), .A3(\add_506/n66 ), .A4(\add_506/n15 ), .ZN(\add_506/n64 ) );
XNOR2_X2 \add_506/U311  ( .A(\add_506/n64 ), .B(n18225), .ZN(N2118) );
NAND4_X2 \add_506/U310  ( .A1(\add_506/n27 ), .A2(\add_506/n21 ), .A3(\add_506/n63 ), .A4(\add_506/n15 ), .ZN(\add_506/n62 ) );
XNOR2_X2 \add_506/U309  ( .A(\add_506/n62 ), .B(n18221), .ZN(N2119) );
INV_X4 \add_506/U308  ( .A(n18221), .ZN(\add_506/n52 ) );
NAND4_X2 \add_506/U307  ( .A1(\add_506/n27 ), .A2(\add_506/n20 ), .A3(\add_506/n61 ), .A4(\add_506/n15 ), .ZN(\add_506/n60 ) );
XNOR2_X2 \add_506/U306  ( .A(\add_506/n60 ), .B(n18217), .ZN(N2120) );
NAND2_X2 \add_506/U305  ( .A1(n18217), .A2(n18221), .ZN(\add_506/n58 ) );
NAND2_X2 \add_506/U304  ( .A1(\add_506/n55 ), .A2(\add_506/n56 ), .ZN(\add_506/n54 ) );
XNOR2_X2 \add_506/U303  ( .A(\add_506/n54 ), .B(n18213), .ZN(N2121) );
NAND2_X2 \add_506/U302  ( .A1(n18217), .A2(n18213), .ZN(\add_506/n53 ) );
NAND4_X2 \add_506/U301  ( .A1(\add_506/n50 ), .A2(\add_506/n21 ), .A3(\add_506/n51 ), .A4(\add_506/n15 ), .ZN(\add_506/n49 ) );
XNOR2_X2 \add_506/U300  ( .A(\add_506/n49 ), .B(n18209), .ZN(N2122) );
NAND4_X2 \add_506/U299  ( .A1(n18209), .A2(n18213), .A3(n18217), .A4(n18221),.ZN(\add_506/n43 ) );
NAND4_X2 \add_506/U298  ( .A1(\add_506/n27 ), .A2(\add_506/n21 ), .A3(\add_506/n48 ), .A4(\add_506/n15 ), .ZN(\add_506/n47 ) );
XNOR2_X2 \add_506/U297  ( .A(\add_506/n47 ), .B(n18205), .ZN(N2123) );
NAND4_X2 \add_506/U296  ( .A1(\add_506/n45 ), .A2(\add_506/n21 ), .A3(\add_506/n46 ), .A4(\add_506/n15 ), .ZN(\add_506/n44 ) );
XNOR2_X2 \add_506/U295  ( .A(\add_506/n44 ), .B(n18201), .ZN(N2124) );
INV_X4 \add_506/U294  ( .A(\add_506/n43 ), .ZN(\add_506/n35 ) );
NAND2_X2 \add_506/U293  ( .A1(n18205), .A2(n18201), .ZN(\add_506/n42 ) );
NAND4_X2 \add_506/U292  ( .A1(\add_506/n35 ), .A2(\add_506/n16 ), .A3(\add_506/n41 ), .A4(\add_506/n19 ), .ZN(\add_506/n40 ) );
XNOR2_X2 \add_506/U291  ( .A(\add_506/n40 ), .B(n18197), .ZN(N2125) );
NAND2_X2 \add_506/U290  ( .A1(n18197), .A2(n18201), .ZN(\add_506/n38 ) );
NAND3_X2 \add_506/U289  ( .A1(\add_506/n36 ), .A2(\add_506/n27 ), .A3(\add_506/n21 ), .ZN(\add_506/n33 ) );
NAND2_X2 \add_506/U288  ( .A1(\add_506/n35 ), .A2(\add_506/n18 ), .ZN(\add_506/n34 ) );
XNOR2_X2 \add_506/U287  ( .A(\add_506/n31 ), .B(\add_506/n32 ), .ZN(N2126));
NAND2_X2 \add_506/U286  ( .A1(n18557), .A2(\add_506/n30 ), .ZN(\add_506/n29 ) );
XNOR2_X2 \add_506/U285  ( .A(\add_506/n29 ), .B(n18553), .ZN(N2036) );
INV_X4 \add_506/U284  ( .A(n18129), .ZN(\add_506/n14 ) );
INV_X4 \add_506/U283  ( .A(n18329), .ZN(\add_506/n12 ) );
NOR2_X2 \add_506/U282  ( .A1(\add_506/n342 ), .A2(\add_506/n348 ), .ZN(\add_506/n347 ) );
NOR2_X2 \add_506/U281  ( .A1(\add_506/n342 ), .A2(\add_506/n343 ), .ZN(\add_506/n340 ) );
NAND3_X2 \add_506/U280  ( .A1(n18149), .A2(n18157), .A3(n18153), .ZN(\add_506/n457 ) );
NOR2_X2 \add_506/U279  ( .A1(\add_506/n25 ), .A2(\add_506/n457 ), .ZN(\add_506/n456 ) );
INV_X4 \add_506/U278  ( .A(n18157), .ZN(\add_506/n13 ) );
INV_X4 \add_506/U277  ( .A(n18333), .ZN(\add_506/n11 ) );
NAND3_X2 \add_506/U276  ( .A1(n18345), .A2(n18353), .A3(n18349), .ZN(\add_506/n634 ) );
NAND3_X2 \add_506/U275  ( .A1(n18089), .A2(n18129), .A3(n18093), .ZN(\add_506/n407 ) );
NOR2_X2 \add_506/U274  ( .A1(\add_506/n144 ), .A2(\add_506/n57 ), .ZN(\add_506/n143 ) );
NOR2_X2 \add_506/U273  ( .A1(\add_506/n405 ), .A2(\add_506/n57 ), .ZN(\add_506/n404 ) );
NOR2_X2 \add_506/U272  ( .A1(\add_506/n397 ), .A2(\add_506/n57 ), .ZN(\add_506/n396 ) );
NAND3_X2 \add_506/U271  ( .A1(n18377), .A2(n18385), .A3(n18381), .ZN(\add_506/n217 ) );
NAND3_X2 \add_506/U270  ( .A1(n18393), .A2(n18389), .A3(n18397), .ZN(\add_506/n216 ) );
NOR2_X2 \add_506/U269  ( .A1(\add_506/n216 ), .A2(\add_506/n217 ), .ZN(\add_506/n215 ) );
NAND3_X2 \add_506/U268  ( .A1(n18357), .A2(n18353), .A3(n18361), .ZN(\add_506/n219 ) );
NOR2_X2 \add_506/U267  ( .A1(\add_506/n288 ), .A2(\add_506/n621 ), .ZN(\add_506/n301 ) );
NAND3_X2 \add_506/U266  ( .A1(n18425), .A2(n18421), .A3(n18429), .ZN(\add_506/n294 ) );
NOR3_X2 \add_506/U265  ( .A1(\add_506/n621 ), .A2(\add_506/n288 ), .A3(\add_506/n294 ), .ZN(\add_506/n293 ) );
NOR3_X2 \add_506/U264  ( .A1(\add_506/n621 ), .A2(\add_506/n288 ), .A3(\add_506/n291 ), .ZN(\add_506/n290 ) );
NOR2_X2 \add_506/U263  ( .A1(\add_506/n234 ), .A2(\add_506/n24 ), .ZN(\add_506/n264 ) );
NOR3_X2 \add_506/U262  ( .A1(\add_506/n24 ), .A2(\add_506/n230 ), .A3(\add_506/n231 ), .ZN(\add_506/n229 ) );
NOR3_X2 \add_506/U261  ( .A1(\add_506/n276 ), .A2(\add_506/n621 ), .A3(\add_506/n277 ), .ZN(\add_506/n275 ) );
NOR2_X2 \add_506/U260  ( .A1(\add_506/n244 ), .A2(\add_506/n24 ), .ZN(\add_506/n258 ) );
NOR2_X2 \add_506/U259  ( .A1(\add_506/n439 ), .A2(\add_506/n57 ), .ZN(\add_506/n429 ) );
NOR2_X2 \add_506/U258  ( .A1(\add_506/n59 ), .A2(\add_506/n431 ), .ZN(\add_506/n430 ) );
NOR2_X2 \add_506/U257  ( .A1(\add_506/n425 ), .A2(\add_506/n57 ), .ZN(\add_506/n416 ) );
NOR3_X2 \add_506/U256  ( .A1(\add_506/n59 ), .A2(\add_506/n418 ), .A3(\add_506/n23 ), .ZN(\add_506/n417 ) );
NAND3_X2 \add_506/U255  ( .A1(n18505), .A2(n18501), .A3(n18509), .ZN(\add_506/n367 ) );
NOR2_X2 \add_506/U254  ( .A1(\add_506/n607 ), .A2(\add_506/n367 ), .ZN(\add_506/n366 ) );
NAND3_X2 \add_506/U253  ( .A1(n18489), .A2(n18485), .A3(n18493), .ZN(\add_506/n357 ) );
NOR3_X2 \add_506/U252  ( .A1(\add_506/n607 ), .A2(\add_506/n339 ), .A3(\add_506/n357 ), .ZN(\add_506/n356 ) );
NOR3_X2 \add_506/U251  ( .A1(\add_506/n338 ), .A2(\add_506/n339 ), .A3(\add_506/n607 ), .ZN(\add_506/n336 ) );
NOR3_X2 \add_506/U250  ( .A1(\add_506/n59 ), .A2(\add_506/n37 ), .A3(\add_506/n23 ), .ZN(\add_506/n55 ) );
NOR2_X2 \add_506/U249  ( .A1(\add_506/n57 ), .A2(\add_506/n58 ), .ZN(\add_506/n56 ) );
NOR3_X2 \add_506/U248  ( .A1(\add_506/n607 ), .A2(\add_506/n352 ), .A3(\add_506/n339 ), .ZN(\add_506/n354 ) );
NOR3_X2 \add_506/U247  ( .A1(\add_506/n37 ), .A2(\add_506/n38 ), .A3(\add_506/n39 ), .ZN(\add_506/n36 ) );
NAND3_X2 \add_506/U246  ( .A1(n18457), .A2(n18461), .A3(\add_506/n15 ), .ZN(\add_506/n312 ) );
NAND3_X2 \add_506/U245  ( .A1(n18117), .A2(n18113), .A3(n18121), .ZN(\add_506/n468 ) );
NOR2_X2 \add_506/U244  ( .A1(\add_506/n13 ), .A2(\add_506/n441 ), .ZN(\add_506/n440 ) );
NOR3_X2 \add_506/U243  ( .A1(\add_506/n465 ), .A2(\add_506/n466 ), .A3(\add_506/n467 ), .ZN(\add_506/n464 ) );
NAND3_X2 \add_506/U242  ( .A1(n18569), .A2(n18573), .A3(\add_506/n4 ), .ZN(\add_506/n177 ) );
AND3_X4 \add_506/U241  ( .A1(n18121), .A2(n18117), .A3(n18125), .ZN(\add_506/n10 ) );
AND2_X4 \add_506/U240  ( .A1(n18109), .A2(n18113), .ZN(\add_506/n9 ) );
NAND2_X2 \add_506/U239  ( .A1(\add_506/n9 ), .A2(\add_506/n10 ), .ZN(\add_506/n8 ) );
NAND3_X2 \add_506/U238  ( .A1(n18269), .A2(n18273), .A3(n18285), .ZN(\add_506/n109 ) );
NOR2_X2 \add_506/U237  ( .A1(\add_506/n644 ), .A2(\add_506/n645 ), .ZN(\add_506/n640 ) );
NOR2_X2 \add_506/U236  ( .A1(\add_506/n642 ), .A2(\add_506/n643 ), .ZN(\add_506/n641 ) );
NAND3_X2 \add_506/U235  ( .A1(n18369), .A2(n18365), .A3(n18373), .ZN(\add_506/n218 ) );
NAND3_X2 \add_506/U234  ( .A1(n18133), .A2(n18129), .A3(n18137), .ZN(\add_506/n421 ) );
NAND3_X2 \add_506/U233  ( .A1(n18145), .A2(n18149), .A3(n18141), .ZN(\add_506/n420 ) );
NOR2_X2 \add_506/U232  ( .A1(\add_506/n420 ), .A2(\add_506/n421 ), .ZN(\add_506/n419 ) );
NOR2_X2 \add_506/U231  ( .A1(\add_506/n236 ), .A2(\add_506/n237 ), .ZN(\add_506/n232 ) );
NOR2_X2 \add_506/U230  ( .A1(\add_506/n234 ), .A2(\add_506/n235 ), .ZN(\add_506/n233 ) );
NAND3_X2 \add_506/U229  ( .A1(n18541), .A2(\add_506/n2 ), .A3(\add_506/n30 ),.ZN(\add_506/n392 ) );
NOR2_X2 \add_506/U228  ( .A1(\add_506/n331 ), .A2(\add_506/n332 ), .ZN(\add_506/n330 ) );
NOR2_X2 \add_506/U227  ( .A1(\add_506/n333 ), .A2(\add_506/n334 ), .ZN(\add_506/n329 ) );
NOR2_X2 \add_506/U226  ( .A1(\add_506/n324 ), .A2(\add_506/n325 ), .ZN(\add_506/n320 ) );
NOR2_X2 \add_506/U225  ( .A1(\add_506/n322 ), .A2(\add_506/n323 ), .ZN(\add_506/n321 ) );
NOR2_X2 \add_506/U224  ( .A1(\add_506/n282 ), .A2(\add_506/n283 ), .ZN(\add_506/n278 ) );
NOR2_X2 \add_506/U223  ( .A1(\add_506/n280 ), .A2(\add_506/n281 ), .ZN(\add_506/n279 ) );
NOR2_X2 \add_506/U222  ( .A1(\add_506/n605 ), .A2(\add_506/n606 ), .ZN(\add_506/n601 ) );
NOR2_X2 \add_506/U221  ( .A1(\add_506/n603 ), .A2(\add_506/n604 ), .ZN(\add_506/n602 ) );
NOR2_X2 \add_506/U220  ( .A1(\add_506/n535 ), .A2(\add_506/n536 ), .ZN(\add_506/n534 ) );
NOR2_X2 \add_506/U219  ( .A1(\add_506/n537 ), .A2(\add_506/n538 ), .ZN(\add_506/n533 ) );
NAND3_X2 \add_506/U218  ( .A1(n18193), .A2(n18197), .A3(n18189), .ZN(\add_506/n548 ) );
NAND3_X2 \add_506/U217  ( .A1(n18301), .A2(n18313), .A3(n18297), .ZN(\add_506/n133 ) );
NOR3_X2 \add_506/U216  ( .A1(\add_506/n57 ), .A2(\add_506/n133 ), .A3(\add_506/n134 ), .ZN(\add_506/n132 ) );
NOR3_X2 \add_506/U215  ( .A1(\add_506/n23 ), .A2(\add_506/n135 ), .A3(\add_506/n181 ), .ZN(\add_506/n180 ) );
NOR2_X2 \add_506/U214  ( .A1(\add_506/n182 ), .A2(\add_506/n183 ), .ZN(\add_506/n179 ) );
NOR3_X2 \add_506/U213  ( .A1(\add_506/n23 ), .A2(\add_506/n135 ), .A3(\add_506/n174 ), .ZN(\add_506/n173 ) );
NOR2_X2 \add_506/U212  ( .A1(\add_506/n175 ), .A2(\add_506/n176 ), .ZN(\add_506/n172 ) );
NOR3_X2 \add_506/U211  ( .A1(\add_506/n23 ), .A2(\add_506/n135 ), .A3(\add_506/n162 ), .ZN(\add_506/n161 ) );
NOR2_X2 \add_506/U210  ( .A1(\add_506/n163 ), .A2(\add_506/n164 ), .ZN(\add_506/n160 ) );
NOR2_X2 \add_506/U209  ( .A1(\add_506/n25 ), .A2(\add_506/n114 ), .ZN(\add_506/n118 ) );
NOR2_X2 \add_506/U208  ( .A1(\add_506/n25 ), .A2(\add_506/n75 ), .ZN(\add_506/n96 ) );
NOR3_X2 \add_506/U207  ( .A1(\add_506/n412 ), .A2(\add_506/n399 ), .A3(\add_506/n400 ), .ZN(\add_506/n395 ) );
OR3_X4 \add_506/U206  ( .A1(\add_506/n149 ), .A2(\add_506/n150 ), .A3(\add_506/n57 ), .ZN(\add_506/n7 ) );
XNOR2_X2 \add_506/U205  ( .A(n18297), .B(\add_506/n7 ), .ZN(N2100) );
NOR3_X2 \add_506/U204  ( .A1(\add_506/n412 ), .A2(\add_506/n406 ), .A3(\add_506/n407 ), .ZN(\add_506/n403 ) );
NOR2_X2 \add_506/U203  ( .A1(\add_506/n59 ), .A2(\add_506/n463 ), .ZN(\add_506/n462 ) );
NOR2_X2 \add_506/U202  ( .A1(\add_506/n451 ), .A2(\add_506/n468 ), .ZN(\add_506/n461 ) );
NOR2_X2 \add_506/U201  ( .A1(\add_506/n59 ), .A2(\add_506/n445 ), .ZN(\add_506/n444 ) );
NOR2_X2 \add_506/U200  ( .A1(\add_506/n451 ), .A2(\add_506/n452 ), .ZN(\add_506/n443 ) );
NOR3_X2 \add_506/U199  ( .A1(\add_506/n24 ), .A2(\add_506/n37 ), .A3(\add_506/n39 ), .ZN(\add_506/n570 ) );
NOR3_X2 \add_506/U198  ( .A1(\add_506/n572 ), .A2(\add_506/n573 ), .A3(\add_506/n574 ), .ZN(\add_506/n571 ) );
NOR3_X2 \add_506/U197  ( .A1(\add_506/n24 ), .A2(\add_506/n37 ), .A3(\add_506/n39 ), .ZN(\add_506/n560 ) );
NOR3_X2 \add_506/U196  ( .A1(\add_506/n562 ), .A2(\add_506/n563 ), .A3(\add_506/n564 ), .ZN(\add_506/n561 ) );
NOR3_X2 \add_506/U195  ( .A1(\add_506/n286 ), .A2(\add_506/n621 ), .A3(\add_506/n287 ), .ZN(\add_506/n285 ) );
NOR3_X2 \add_506/U194  ( .A1(\add_506/n346 ), .A2(\add_506/n339 ), .A3(\add_506/n607 ), .ZN(\add_506/n345 ) );
NOR3_X2 \add_506/U193  ( .A1(\add_506/n412 ), .A2(\add_506/n413 ), .A3(\add_506/n414 ), .ZN(\add_506/n409 ) );
NOR2_X2 \add_506/U192  ( .A1(\add_506/n483 ), .A2(\add_506/n484 ), .ZN(\add_506/n482 ) );
NOR2_X2 \add_506/U191  ( .A1(\add_506/n135 ), .A2(\add_506/n145 ), .ZN(\add_506/n142 ) );
NOR3_X2 \add_506/U190  ( .A1(\add_506/n146 ), .A2(\add_506/n147 ), .A3(\add_506/n148 ), .ZN(\add_506/n141 ) );
NOR3_X2 \add_506/U189  ( .A1(\add_506/n351 ), .A2(\add_506/n339 ), .A3(\add_506/n607 ), .ZN(\add_506/n350 ) );
NOR3_X2 \add_506/U188  ( .A1(\add_506/n59 ), .A2(\add_506/n23 ), .A3(\add_506/n465 ), .ZN(\add_506/n472 ) );
NOR3_X2 \add_506/U187  ( .A1(\add_506/n473 ), .A2(\add_506/n474 ), .A3(\add_506/n475 ), .ZN(\add_506/n471 ) );
NAND3_X2 \add_506/U186  ( .A1(n18185), .A2(n18181), .A3(n18189), .ZN(\add_506/n585 ) );
NOR3_X2 \add_506/U185  ( .A1(\add_506/n24 ), .A2(\add_506/n584 ), .A3(\add_506/n585 ), .ZN(\add_506/n583 ) );
NOR3_X2 \add_506/U184  ( .A1(\add_506/n23 ), .A2(\add_506/n135 ), .A3(\add_506/n168 ), .ZN(\add_506/n167 ) );
NOR2_X2 \add_506/U183  ( .A1(\add_506/n169 ), .A2(\add_506/n170 ), .ZN(\add_506/n166 ) );
NOR2_X2 \add_506/U182  ( .A1(\add_506/n57 ), .A2(\add_506/n451 ), .ZN(\add_506/n455 ) );
NOR3_X2 \add_506/U181  ( .A1(\add_506/n8 ), .A2(\add_506/n458 ), .A3(\add_506/n459 ), .ZN(\add_506/n454 ) );
NAND3_X2 \add_506/U180  ( .A1(n18525), .A2(n18521), .A3(\add_506/n337 ),.ZN(\add_506/n372 ) );
NAND3_X2 \add_506/U179  ( .A1(n18541), .A2(n18545), .A3(n18537), .ZN(\add_506/n391 ) );
NOR2_X2 \add_506/U178  ( .A1(\add_506/n390 ), .A2(\add_506/n391 ), .ZN(\add_506/n389 ) );
NAND3_X2 \add_506/U177  ( .A1(n18549), .A2(n18553), .A3(n18557), .ZN(\add_506/n386 ) );
NOR2_X2 \add_506/U176  ( .A1(\add_506/n386 ), .A2(\add_506/n387 ), .ZN(\add_506/n385 ) );
NOR2_X2 \add_506/U175  ( .A1(\add_506/n280 ), .A2(\add_506/n621 ), .ZN(\add_506/n309 ) );
NAND3_X2 \add_506/U174  ( .A1(n18509), .A2(\add_506/n362 ), .A3(\add_506/n337 ), .ZN(\add_506/n369 ) );
NOR2_X2 \add_506/U173  ( .A1(\add_506/n122 ), .A2(\add_506/n123 ), .ZN(\add_506/n121 ) );
NOR3_X2 \add_506/U172  ( .A1(\add_506/n24 ), .A2(\add_506/n584 ), .A3(\add_506/n588 ), .ZN(\add_506/n587 ) );
NAND3_X2 \add_506/U171  ( .A1(n18425), .A2(n18421), .A3(n18429), .ZN(\add_506/n273 ) );
NOR3_X2 \add_506/U170  ( .A1(\add_506/n317 ), .A2(\add_506/n318 ), .A3(\add_506/n319 ), .ZN(\add_506/n316 ) );
NOR3_X2 \add_506/U169  ( .A1(\add_506/n326 ), .A2(\add_506/n327 ), .A3(\add_506/n328 ), .ZN(\add_506/n315 ) );
NOR2_X2 \add_506/U168  ( .A1(\add_506/n339 ), .A2(\add_506/n607 ), .ZN(\add_506/n364 ) );
NAND3_X2 \add_506/U167  ( .A1(n18157), .A2(n18153), .A3(\add_506/n398 ),.ZN(\add_506/n411 ) );
NOR2_X2 \add_506/U166  ( .A1(\add_506/n411 ), .A2(\add_506/n57 ), .ZN(\add_506/n410 ) );
NAND3_X2 \add_506/U165  ( .A1(n18549), .A2(\add_506/n3 ), .A3(\add_506/n30 ),.ZN(\add_506/n469 ) );
NOR3_X2 \add_506/U164  ( .A1(\add_506/n621 ), .A2(\add_506/n297 ), .A3(\add_506/n288 ), .ZN(\add_506/n296 ) );
NAND3_X2 \add_506/U163  ( .A1(n18197), .A2(n18193), .A3(n18201), .ZN(\add_506/n564 ) );
NAND3_X2 \add_506/U162  ( .A1(n18093), .A2(n18133), .A3(n18129), .ZN(\add_506/n414 ) );
NAND3_X2 \add_506/U161  ( .A1(n18549), .A2(n18553), .A3(n18557), .ZN(\add_506/n390 ) );
NOR3_X2 \add_506/U160  ( .A1(\add_506/n23 ), .A2(\add_506/n37 ), .A3(\add_506/n42 ), .ZN(\add_506/n41 ) );
NOR2_X2 \add_506/U159  ( .A1(\add_506/n493 ), .A2(\add_506/n501 ), .ZN(\add_506/n499 ) );
NAND3_X2 \add_506/U158  ( .A1(n18377), .A2(n18373), .A3(n18381), .ZN(\add_506/n227 ) );
NOR3_X2 \add_506/U157  ( .A1(\add_506/n24 ), .A2(\add_506/n255 ), .A3(\add_506/n244 ), .ZN(\add_506/n254 ) );
NAND3_X2 \add_506/U156  ( .A1(n18153), .A2(n18149), .A3(n18157), .ZN(\add_506/n515 ) );
NOR2_X2 \add_506/U155  ( .A1(\add_506/n25 ), .A2(\add_506/n515 ), .ZN(\add_506/n514 ) );
NAND3_X2 \add_506/U154  ( .A1(n18317), .A2(n18313), .A3(n18321), .ZN(\add_506/n174 ) );
NOR2_X2 \add_506/U153  ( .A1(\add_506/n135 ), .A2(\add_506/n136 ), .ZN(\add_506/n131 ) );
NOR3_X2 \add_506/U152  ( .A1(\add_506/n137 ), .A2(\add_506/n138 ), .A3(\add_506/n139 ), .ZN(\add_506/n130 ) );
NOR3_X2 \add_506/U151  ( .A1(\add_506/n24 ), .A2(\add_506/n580 ), .A3(\add_506/n581 ), .ZN(\add_506/n576 ) );
NOR3_X2 \add_506/U150  ( .A1(\add_506/n37 ), .A2(\add_506/n578 ), .A3(\add_506/n579 ), .ZN(\add_506/n577 ) );
NOR2_X2 \add_506/U149  ( .A1(\add_506/n607 ), .A2(\add_506/n339 ), .ZN(\add_506/n359 ) );
NOR3_X2 \add_506/U148  ( .A1(\add_506/n24 ), .A2(\add_506/n37 ), .A3(\add_506/n558 ), .ZN(\add_506/n544 ) );
NOR3_X2 \add_506/U147  ( .A1(\add_506/n546 ), .A2(\add_506/n547 ), .A3(\add_506/n548 ), .ZN(\add_506/n545 ) );
NOR2_X2 \add_506/U146  ( .A1(\add_506/n226 ), .A2(\add_506/n227 ), .ZN(\add_506/n222 ) );
NOR2_X2 \add_506/U145  ( .A1(\add_506/n224 ), .A2(\add_506/n225 ), .ZN(\add_506/n223 ) );
NOR3_X2 \add_506/U144  ( .A1(\add_506/n135 ), .A2(\add_506/n12 ), .A3(\add_506/n187 ), .ZN(\add_506/n193 ) );
NOR2_X2 \add_506/U143  ( .A1(\add_506/n194 ), .A2(\add_506/n195 ), .ZN(\add_506/n192 ) );
NOR2_X2 \add_506/U142  ( .A1(\add_506/n621 ), .A2(\add_506/n280 ), .ZN(\add_506/n306 ) );
NOR2_X2 \add_506/U141  ( .A1(\add_506/n272 ), .A2(\add_506/n273 ), .ZN(\add_506/n268 ) );
NOR2_X2 \add_506/U140  ( .A1(\add_506/n270 ), .A2(\add_506/n271 ), .ZN(\add_506/n269 ) );
NOR2_X2 \add_506/U139  ( .A1(\add_506/n25 ), .A2(\add_506/n234 ), .ZN(\add_506/n260 ) );
NOR2_X2 \add_506/U138  ( .A1(\add_506/n236 ), .A2(\add_506/n252 ), .ZN(\add_506/n251 ) );
NOR2_X2 \add_506/U137  ( .A1(\add_506/n248 ), .A2(\add_506/n249 ), .ZN(\add_506/n246 ) );
NOR2_X2 \add_506/U136  ( .A1(\add_506/n243 ), .A2(\add_506/n244 ), .ZN(\add_506/n239 ) );
NOR2_X2 \add_506/U135  ( .A1(\add_506/n241 ), .A2(\add_506/n242 ), .ZN(\add_506/n240 ) );
NOR3_X2 \add_506/U134  ( .A1(\add_506/n135 ), .A2(\add_506/n187 ), .A3(\add_506/n188 ), .ZN(\add_506/n186 ) );
NOR2_X2 \add_506/U133  ( .A1(\add_506/n189 ), .A2(\add_506/n190 ), .ZN(\add_506/n185 ) );
NOR2_X2 \add_506/U132  ( .A1(\add_506/n122 ), .A2(\add_506/n126 ), .ZN(\add_506/n125 ) );
NOR2_X2 \add_506/U131  ( .A1(\add_506/n25 ), .A2(\add_506/n114 ), .ZN(\add_506/n116 ) );
NOR2_X2 \add_506/U130  ( .A1(\add_506/n114 ), .A2(\add_506/n24 ), .ZN(\add_506/n112 ) );
NOR2_X2 \add_506/U129  ( .A1(\add_506/n102 ), .A2(\add_506/n103 ), .ZN(\add_506/n113 ) );
NOR3_X2 \add_506/U128  ( .A1(\add_506/n23 ), .A2(\add_506/n109 ), .A3(\add_506/n110 ), .ZN(\add_506/n107 ) );
NOR2_X2 \add_506/U127  ( .A1(\add_506/n103 ), .A2(\add_506/n104 ), .ZN(\add_506/n108 ) );
NOR2_X2 \add_506/U126  ( .A1(\add_506/n25 ), .A2(\add_506/n75 ), .ZN(\add_506/n94 ) );
NOR2_X2 \add_506/U125  ( .A1(\add_506/n75 ), .A2(\add_506/n25 ), .ZN(\add_506/n90 ) );
NOR2_X2 \add_506/U124  ( .A1(\add_506/n87 ), .A2(\add_506/n92 ), .ZN(\add_506/n91 ) );
NOR2_X2 \add_506/U123  ( .A1(\add_506/n75 ), .A2(\add_506/n25 ), .ZN(\add_506/n85 ) );
NOR2_X2 \add_506/U122  ( .A1(\add_506/n87 ), .A2(\add_506/n88 ), .ZN(\add_506/n86 ) );
NOR2_X2 \add_506/U121  ( .A1(\add_506/n1 ), .A2(\add_506/n81 ), .ZN(\add_506/n80 ) );
NOR3_X2 \add_506/U120  ( .A1(\add_506/n23 ), .A2(\add_506/n75 ), .A3(\add_506/n76 ), .ZN(\add_506/n74 ) );
NOR2_X2 \add_506/U119  ( .A1(\add_506/n67 ), .A2(\add_506/n77 ), .ZN(\add_506/n73 ) );
NOR2_X2 \add_506/U118  ( .A1(\add_506/n69 ), .A2(\add_506/n25 ), .ZN(\add_506/n65 ) );
NOR2_X2 \add_506/U117  ( .A1(\add_506/n67 ), .A2(\add_506/n68 ), .ZN(\add_506/n66 ) );
NOR2_X2 \add_506/U116  ( .A1(\add_506/n52 ), .A2(\add_506/n37 ), .ZN(\add_506/n61 ) );
NOR2_X2 \add_506/U115  ( .A1(\add_506/n37 ), .A2(\add_506/n25 ), .ZN(\add_506/n50 ) );
NOR2_X2 \add_506/U114  ( .A1(\add_506/n52 ), .A2(\add_506/n53 ), .ZN(\add_506/n51 ) );
NOR2_X2 \add_506/U113  ( .A1(\add_506/n37 ), .A2(\add_506/n43 ), .ZN(\add_506/n48 ) );
NOR2_X2 \add_506/U112  ( .A1(\add_506/n39 ), .A2(\add_506/n25 ), .ZN(\add_506/n45 ) );
NOR2_X2 \add_506/U111  ( .A1(\add_506/n37 ), .A2(\add_506/n43 ), .ZN(\add_506/n46 ) );
NOR2_X2 \add_506/U110  ( .A1(\add_506/n1 ), .A2(\add_506/n584 ), .ZN(\add_506/n594 ) );
NOR2_X2 \add_506/U109  ( .A1(\add_506/n1 ), .A2(\add_506/n591 ), .ZN(\add_506/n590 ) );
NAND3_X2 \add_506/U108  ( .A1(n18321), .A2(n18317), .A3(n18325), .ZN(\add_506/n181 ) );
NAND3_X2 \add_506/U107  ( .A1(n18133), .A2(n18141), .A3(n18129), .ZN(\add_506/n458 ) );
NOR2_X2 \add_506/U106  ( .A1(\add_506/n57 ), .A2(\add_506/n59 ), .ZN(\add_506/n504 ) );
NOR3_X2 \add_506/U105  ( .A1(\add_506/n505 ), .A2(\add_506/n493 ), .A3(\add_506/n494 ), .ZN(\add_506/n503 ) );
NAND3_X2 \add_506/U104  ( .A1(n18321), .A2(n18317), .A3(n18325), .ZN(\add_506/n636 ) );
NOR2_X2 \add_506/U103  ( .A1(\add_506/n635 ), .A2(\add_506/n636 ), .ZN(\add_506/n628 ) );
NOR2_X2 \add_506/U102  ( .A1(\add_506/n621 ), .A2(\add_506/n622 ), .ZN(\add_506/n620 ) );
NAND3_X2 \add_506/U101  ( .A1(n18377), .A2(n18373), .A3(n18381), .ZN(\add_506/n632 ) );
NOR2_X2 \add_506/U100  ( .A1(\add_506/n631 ), .A2(\add_506/n632 ), .ZN(\add_506/n630 ) );
NAND3_X2 \add_506/U99  ( .A1(n18293), .A2(n18289), .A3(n18297), .ZN(\add_506/n638 ) );
NOR2_X2 \add_506/U98  ( .A1(\add_506/n637 ), .A2(\add_506/n638 ), .ZN(\add_506/n627 ) );
NOR3_X2 \add_506/U97  ( .A1(\add_506/n422 ), .A2(\add_506/n423 ), .A3(\add_506/n424 ), .ZN(\add_506/n401 ) );
NOR3_X2 \add_506/U96  ( .A1(\add_506/n520 ), .A2(\add_506/n521 ), .A3(\add_506/n522 ), .ZN(\add_506/n30 ) );
NOR2_X2 \add_506/U95  ( .A1(\add_506/n633 ), .A2(\add_506/n634 ), .ZN(\add_506/n629 ) );
NAND4_X2 \add_506/U94  ( .A1(\add_506/n627 ), .A2(\add_506/n628 ), .A3(\add_506/n629 ), .A4(\add_506/n630 ), .ZN(\add_506/n59 ) );
NAND3_X2 \add_506/U93  ( .A1(n18333), .A2(n18337), .A3(n18349), .ZN(\add_506/n194 ) );
NAND3_X2 \add_506/U92  ( .A1(n18345), .A2(n18341), .A3(n18349), .ZN(\add_506/n189 ) );
NAND3_X2 \add_506/U91  ( .A1(n18345), .A2(n18341), .A3(n18349), .ZN(\add_506/n182 ) );
NAND3_X2 \add_506/U90  ( .A1(n18329), .A2(n18337), .A3(n18333), .ZN(\add_506/n190 ) );
NAND3_X2 \add_506/U89  ( .A1(n18329), .A2(n18337), .A3(n18333), .ZN(\add_506/n183 ) );
NAND3_X2 \add_506/U88  ( .A1(n18329), .A2(n18325), .A3(n18333), .ZN(\add_506/n176 ) );
NAND3_X2 \add_506/U87  ( .A1(n18329), .A2(n18325), .A3(n18333), .ZN(\add_506/n170 ) );
NAND3_X2 \add_506/U86  ( .A1(n18333), .A2(n18337), .A3(n18349), .ZN(\add_506/n147 ) );
NAND3_X2 \add_506/U85  ( .A1(n18333), .A2(n18337), .A3(n18349), .ZN(\add_506/n138 ) );
NOR2_X2 \add_506/U84  ( .A1(\add_506/n646 ), .A2(\add_506/n647 ), .ZN(\add_506/n639 ) );
NAND3_X2 \add_506/U83  ( .A1(\add_506/n639 ), .A2(\add_506/n640 ), .A3(\add_506/n641 ), .ZN(\add_506/n37 ) );
NOR2_X2 \add_506/U82  ( .A1(\add_506/n25 ), .A2(\add_506/n465 ), .ZN(\add_506/n479 ) );
NOR2_X2 \add_506/U81  ( .A1(\add_506/n135 ), .A2(\add_506/n154 ), .ZN(\add_506/n153 ) );
NOR2_X2 \add_506/U80  ( .A1(\add_506/n157 ), .A2(\add_506/n158 ), .ZN(\add_506/n151 ) );
NOR2_X2 \add_506/U79  ( .A1(\add_506/n155 ), .A2(\add_506/n156 ), .ZN(\add_506/n152 ) );
NOR2_X2 \add_506/U78  ( .A1(\add_506/n33 ), .A2(\add_506/n34 ), .ZN(\add_506/n32 ) );
NOR2_X2 \add_506/U77  ( .A1(\add_506/n491 ), .A2(\add_506/n492 ), .ZN(\add_506/n490 ) );
NOR2_X2 \add_506/U76  ( .A1(\add_506/n493 ), .A2(\add_506/n494 ), .ZN(\add_506/n489 ) );
NOR2_X2 \add_506/U75  ( .A1(\add_506/n495 ), .A2(\add_506/n14 ), .ZN(\add_506/n488 ) );
NAND3_X2 \add_506/U74  ( .A1(\add_506/n488 ), .A2(\add_506/n489 ), .A3(\add_506/n490 ), .ZN(\add_506/n474 ) );
NOR2_X2 \add_506/U73  ( .A1(\add_506/n218 ), .A2(\add_506/n219 ), .ZN(\add_506/n214 ) );
NAND2_X2 \add_506/U72  ( .A1(\add_506/n214 ), .A2(\add_506/n215 ), .ZN(\add_506/n135 ) );
NOR2_X2 \add_506/U71  ( .A1(\add_506/n135 ), .A2(\add_506/n24 ), .ZN(\add_506/n213 ) );
NAND3_X2 \add_506/U70  ( .A1(n18345), .A2(n18341), .A3(n18349), .ZN(\add_506/n206 ) );
NOR3_X2 \add_506/U69  ( .A1(\add_506/n24 ), .A2(\add_506/n135 ), .A3(\add_506/n206 ), .ZN(\add_506/n205 ) );
NOR3_X2 \add_506/U68  ( .A1(\add_506/n23 ), .A2(\add_506/n209 ), .A3(\add_506/n135 ), .ZN(\add_506/n208 ) );
NOR3_X2 \add_506/U67  ( .A1(\add_506/n23 ), .A2(\add_506/n135 ), .A3(\add_506/n199 ), .ZN(\add_506/n203 ) );
NOR2_X2 \add_506/U66  ( .A1(\add_506/n505 ), .A2(\add_506/n493 ), .ZN(\add_506/n509 ) );
NOR2_X2 \add_506/U65  ( .A1(\add_506/n378 ), .A2(\add_506/n379 ), .ZN(\add_506/n377 ) );
NOR2_X2 \add_506/U64  ( .A1(\add_506/n380 ), .A2(\add_506/n381 ), .ZN(\add_506/n376 ) );
NOR2_X2 \add_506/U63  ( .A1(\add_506/n382 ), .A2(\add_506/n383 ), .ZN(\add_506/n375 ) );
NAND3_X2 \add_506/U62  ( .A1(\add_506/n375 ), .A2(\add_506/n376 ), .A3(\add_506/n377 ), .ZN(\add_506/n374 ) );
NOR2_X2 \add_506/U61  ( .A1(\add_506/n427 ), .A2(\add_506/n13 ), .ZN(\add_506/n426 ) );
NOR2_X2 \add_506/U60  ( .A1(\add_506/n447 ), .A2(\add_506/n434 ), .ZN(\add_506/n446 ) );
NOR2_X2 \add_506/U59  ( .A1(\add_506/n433 ), .A2(\add_506/n434 ), .ZN(\add_506/n432 ) );
NOR2_X2 \add_506/U58  ( .A1(\add_506/n614 ), .A2(\add_506/n615 ), .ZN(\add_506/n613 ) );
NOR2_X2 \add_506/U57  ( .A1(\add_506/n39 ), .A2(\add_506/n616 ), .ZN(\add_506/n612 ) );
NOR2_X2 \add_506/U56  ( .A1(\add_506/n617 ), .A2(\add_506/n31 ), .ZN(\add_506/n611 ) );
NAND3_X2 \add_506/U55  ( .A1(\add_506/n611 ), .A2(\add_506/n612 ), .A3(\add_506/n613 ), .ZN(\add_506/n584 ) );
NOR3_X2 \add_506/U54  ( .A1(\add_506/n23 ), .A2(\add_506/n199 ), .A3(\add_506/n135 ), .ZN(\add_506/n198 ) );
NOR2_X2 \add_506/U53  ( .A1(\add_506/n11 ), .A2(\add_506/n12 ), .ZN(\add_506/n197 ) );
NOR2_X2 \add_506/U52  ( .A1(\add_506/n623 ), .A2(\add_506/n624 ), .ZN(\add_506/n619 ) );
NOR2_X2 \add_506/U51  ( .A1(\add_506/n625 ), .A2(\add_506/n626 ), .ZN(\add_506/n618 ) );
NOR2_X2 \add_506/U50  ( .A1(\add_506/n135 ), .A2(\add_506/n199 ), .ZN(\add_506/n201 ) );
NOR2_X2 \add_506/U49  ( .A1(\add_506/n25 ), .A2(\add_506/n498 ), .ZN(\add_506/n497 ) );
OR2_X4 \add_506/U48  ( .A1(\add_506/n516 ), .A2(\add_506/n517 ), .ZN(\add_506/n6 ) );
XNOR2_X2 \add_506/U47  ( .A(n18149), .B(\add_506/n6 ), .ZN(N2137) );
NOR2_X2 \add_506/U46  ( .A1(\add_506/n477 ), .A2(\add_506/n478 ), .ZN(\add_506/n476 ) );
NOR2_X2 \add_506/U45  ( .A1(\add_506/n486 ), .A2(\add_506/n487 ), .ZN(\add_506/n485 ) );
NOR2_X2 \add_506/U44  ( .A1(\add_506/n507 ), .A2(\add_506/n508 ), .ZN(\add_506/n506 ) );
NOR2_X2 \add_506/U43  ( .A1(\add_506/n524 ), .A2(\add_506/n525 ), .ZN(\add_506/n523 ) );
NOR2_X2 \add_506/U42  ( .A1(\add_506/n511 ), .A2(\add_506/n512 ), .ZN(\add_506/n510 ) );
NOR3_X2 \add_506/U41  ( .A1(\add_506/n530 ), .A2(\add_506/n531 ), .A3(\add_506/n532 ), .ZN(\add_506/n529 ) );
NOR2_X2 \add_506/U40  ( .A1(\add_506/n541 ), .A2(\add_506/n542 ), .ZN(\add_506/n527 ) );
NOR2_X2 \add_506/U39  ( .A1(\add_506/n539 ), .A2(\add_506/n540 ), .ZN(\add_506/n528 ) );
NAND3_X2 \add_506/U38  ( .A1(\add_506/n527 ), .A2(\add_506/n528 ), .A3(\add_506/n529 ), .ZN(\add_506/n451 ) );
NOR2_X2 \add_506/U37  ( .A1(\add_506/n427 ), .A2(\add_506/n13 ), .ZN(\add_506/n518 ) );
NOR2_X2 \add_506/U36  ( .A1(\add_506/n100 ), .A2(\add_506/n101 ), .ZN(\add_506/n99 ) );
NOR2_X2 \add_506/U35  ( .A1(\add_506/n102 ), .A2(\add_506/n103 ), .ZN(\add_506/n98 ) );
NOR2_X2 \add_506/U34  ( .A1(\add_506/n104 ), .A2(\add_506/n105 ), .ZN(\add_506/n97 ) );
NAND3_X2 \add_506/U33  ( .A1(\add_506/n97 ), .A2(\add_506/n98 ), .A3(\add_506/n99 ), .ZN(\add_506/n75 ) );
NOR2_X2 \add_506/U32  ( .A1(\add_506/n568 ), .A2(\add_506/n552 ), .ZN(\add_506/n567 ) );
NOR2_X2 \add_506/U31  ( .A1(\add_506/n553 ), .A2(\add_506/n554 ), .ZN(\add_506/n566 ) );
NOR2_X2 \add_506/U30  ( .A1(\add_506/n555 ), .A2(\add_506/n556 ), .ZN(\add_506/n565 ) );
NOR2_X2 \add_506/U29  ( .A1(\add_506/n552 ), .A2(\add_506/n553 ), .ZN(\add_506/n551 ) );
NOR2_X2 \add_506/U28  ( .A1(\add_506/n554 ), .A2(\add_506/n555 ), .ZN(\add_506/n550 ) );
NOR2_X2 \add_506/U27  ( .A1(\add_506/n556 ), .A2(\add_506/n557 ), .ZN(\add_506/n549 ) );
NOR3_X2 \add_506/U26  ( .A1(\add_506/n598 ), .A2(\add_506/n599 ), .A3(\add_506/n600 ), .ZN(\add_506/n597 ) );
NOR2_X2 \add_506/U25  ( .A1(\add_506/n607 ), .A2(\add_506/n608 ), .ZN(\add_506/n596 ) );
NOR2_X2 \add_506/U24  ( .A1(\add_506/n609 ), .A2(\add_506/n610 ), .ZN(\add_506/n595 ) );
NAND3_X2 \add_506/U23  ( .A1(\add_506/n595 ), .A2(\add_506/n596 ), .A3(\add_506/n597 ), .ZN(\add_506/n57 ) );
INV_X4 \add_506/U22  ( .A(\add_506/n1 ), .ZN(\add_506/n28 ) );
INV_X4 \add_506/U21  ( .A(\add_506/n374 ), .ZN(\add_506/n337 ) );
INV_X4 \add_506/U20  ( .A(\add_506/n451 ), .ZN(\add_506/n398 ) );
INV_X4 \add_506/U19  ( .A(\add_506/n57 ), .ZN(\add_506/n15 ) );
INV_X4 \add_506/U18  ( .A(\add_506/n59 ), .ZN(\add_506/n19 ) );
INV_X4 \add_506/U17  ( .A(\add_506/n1 ), .ZN(\add_506/n27 ) );
INV_X4 \add_506/U16  ( .A(\add_506/n1 ), .ZN(\add_506/n26 ) );
INV_X4 \add_506/U15  ( .A(\add_506/n59 ), .ZN(\add_506/n22 ) );
INV_X4 \add_506/U14  ( .A(\add_506/n57 ), .ZN(\add_506/n18 ) );
INV_X4 \add_506/U13  ( .A(\add_506/n59 ), .ZN(\add_506/n21 ) );
INV_X4 \add_506/U12  ( .A(\add_506/n59 ), .ZN(\add_506/n20 ) );
INV_X4 \add_506/U11  ( .A(\add_506/n28 ), .ZN(\add_506/n25 ) );
INV_X4 \add_506/U10  ( .A(\add_506/n28 ), .ZN(\add_506/n24 ) );
INV_X4 \add_506/U9  ( .A(\add_506/n26 ), .ZN(\add_506/n23 ) );
INV_X4 \add_506/U8  ( .A(\add_506/n57 ), .ZN(\add_506/n16 ) );
INV_X4 \add_506/U7  ( .A(\add_506/n57 ), .ZN(\add_506/n17 ) );
XOR2_X2 \add_506/U6  ( .A(n18585), .B(n18589), .Z(N2028) );
AND4_X4 \add_506/U5  ( .A1(n18577), .A2(n18581), .A3(n18585), .A4(n18589),.ZN(\add_506/n4 ) );
AND2_X4 \add_506/U4  ( .A1(n18553), .A2(n18557), .ZN(\add_506/n3 ) );
AND4_X4 \add_506/U3  ( .A1(n18545), .A2(n18549), .A3(n18553), .A4(n18557),.ZN(\add_506/n2 ) );
NAND3_X2 \add_506/U2  ( .A1(\add_506/n618 ), .A2(\add_506/n619 ), .A3(\add_506/n620 ), .ZN(\add_506/n1 ) );
NAND2_X2 \add_1_root_add_519_2/U289  ( .A1(n17750), .A2(aad_byte_cnt[0]),.ZN(\add_1_root_add_519_2/n185 ) );
NAND2_X2 \add_1_root_add_519_2/U288  ( .A1(\add_1_root_add_519_2/n185 ),.A2(\add_1_root_add_519_2/n210 ), .ZN(N2479) );
INV_X4 \add_1_root_add_519_2/U287  ( .A(aad_byte_cnt[7]), .ZN(\add_1_root_add_519_2/n224 ) );
INV_X4 \add_1_root_add_519_2/U286  ( .A(\add_1_root_add_519_2/n198 ), .ZN(\add_1_root_add_519_2/n194 ) );
NAND2_X2 \add_1_root_add_519_2/U285  ( .A1(\add_1_root_add_519_2/n219 ),.A2(\add_1_root_add_519_2/n220 ), .ZN(\add_1_root_add_519_2/n214 ) );
NAND2_X2 \add_1_root_add_519_2/U284  ( .A1(dii_data_size[2]), .A2(aad_byte_cnt[2]), .ZN(\add_1_root_add_519_2/n142 ) );
INV_X4 \add_1_root_add_519_2/U283  ( .A(\add_1_root_add_519_2/n142 ), .ZN(\add_1_root_add_519_2/n217 ) );
NAND2_X2 \add_1_root_add_519_2/U282  ( .A1(n18074), .A2(aad_byte_cnt[3]),.ZN(\add_1_root_add_519_2/n139 ) );
INV_X4 \add_1_root_add_519_2/U281  ( .A(\add_1_root_add_519_2/n139 ), .ZN(\add_1_root_add_519_2/n218 ) );
INV_X4 \add_1_root_add_519_2/U280  ( .A(aad_byte_cnt[3]), .ZN(\add_1_root_add_519_2/n213 ) );
NAND2_X2 \add_1_root_add_519_2/U279  ( .A1(\add_1_root_add_519_2/n61 ), .A2(\add_1_root_add_519_2/n213 ), .ZN(\add_1_root_add_519_2/n140 ) );
NAND2_X2 \add_1_root_add_519_2/U278  ( .A1(\add_1_root_add_519_2/n193 ),.A2(\add_1_root_add_519_2/n140 ), .ZN(\add_1_root_add_519_2/n209 ) );
INV_X4 \add_1_root_add_519_2/U277  ( .A(\add_1_root_add_519_2/n140 ), .ZN(\add_1_root_add_519_2/n212 ) );
NAND2_X2 \add_1_root_add_519_2/U276  ( .A1(\add_1_root_add_519_2/n209 ),.A2(\add_1_root_add_519_2/n200 ), .ZN(\add_1_root_add_519_2/n80 ) );
NAND2_X2 \add_1_root_add_519_2/U275  ( .A1(\add_1_root_add_519_2/n194 ),.A2(\add_1_root_add_519_2/n80 ), .ZN(\add_1_root_add_519_2/n208 ) );
XNOR2_X2 \add_1_root_add_519_2/U274  ( .A(\add_1_root_add_519_2/n59 ), .B(aad_byte_cnt[10]), .ZN(N2489) );
INV_X4 \add_1_root_add_519_2/U273  ( .A(aad_byte_cnt[11]), .ZN(\add_1_root_add_519_2/n207 ) );
XNOR2_X2 \add_1_root_add_519_2/U272  ( .A(\add_1_root_add_519_2/n32 ), .B(aad_byte_cnt[11]), .ZN(N2490) );
INV_X4 \add_1_root_add_519_2/U271  ( .A(aad_byte_cnt[12]), .ZN(\add_1_root_add_519_2/n204 ) );
XNOR2_X2 \add_1_root_add_519_2/U270  ( .A(\add_1_root_add_519_2/n5 ), .B(\add_1_root_add_519_2/n204 ), .ZN(N2491) );
INV_X4 \add_1_root_add_519_2/U269  ( .A(aad_byte_cnt[13]), .ZN(\add_1_root_add_519_2/n203 ) );
XNOR2_X2 \add_1_root_add_519_2/U268  ( .A(\add_1_root_add_519_2/n6 ), .B(\add_1_root_add_519_2/n203 ), .ZN(N2492) );
INV_X4 \add_1_root_add_519_2/U267  ( .A(aad_byte_cnt[14]), .ZN(\add_1_root_add_519_2/n202 ) );
XNOR2_X2 \add_1_root_add_519_2/U266  ( .A(\add_1_root_add_519_2/n9 ), .B(\add_1_root_add_519_2/n202 ), .ZN(N2493) );
INV_X4 \add_1_root_add_519_2/U265  ( .A(aad_byte_cnt[15]), .ZN(\add_1_root_add_519_2/n201 ) );
XNOR2_X2 \add_1_root_add_519_2/U264  ( .A(\add_1_root_add_519_2/n30 ), .B(\add_1_root_add_519_2/n201 ), .ZN(N2494) );
NAND2_X2 \add_1_root_add_519_2/U263  ( .A1(\add_1_root_add_519_2/n196 ),.A2(\add_1_root_add_519_2/n197 ), .ZN(\add_1_root_add_519_2/n195 ) );
XNOR2_X2 \add_1_root_add_519_2/U262  ( .A(\add_1_root_add_519_2/n152 ), .B(aad_byte_cnt[16]), .ZN(N2495) );
XNOR2_X2 \add_1_root_add_519_2/U261  ( .A(\add_1_root_add_519_2/n189 ), .B(\add_1_root_add_519_2/n4 ), .ZN(N2496) );
NAND2_X2 \add_1_root_add_519_2/U260  ( .A1(\add_1_root_add_519_2/n4 ), .A2(aad_byte_cnt[17]), .ZN(\add_1_root_add_519_2/n188 ) );
XNOR2_X2 \add_1_root_add_519_2/U259  ( .A(\add_1_root_add_519_2/n188 ), .B(aad_byte_cnt[18]), .ZN(N2497) );
INV_X4 \add_1_root_add_519_2/U258  ( .A(aad_byte_cnt[19]), .ZN(\add_1_root_add_519_2/n187 ) );
XNOR2_X2 \add_1_root_add_519_2/U257  ( .A(\add_1_root_add_519_2/n40 ), .B(aad_byte_cnt[19]), .ZN(N2498) );
NAND2_X2 \add_1_root_add_519_2/U256  ( .A1(dii_data_size[1]), .A2(aad_byte_cnt[1]), .ZN(\add_1_root_add_519_2/n164 ) );
INV_X4 \add_1_root_add_519_2/U255  ( .A(\add_1_root_add_519_2/n164 ), .ZN(\add_1_root_add_519_2/n184 ) );
XNOR2_X2 \add_1_root_add_519_2/U254  ( .A(\add_1_root_add_519_2/n166 ), .B(\add_1_root_add_519_2/n183 ), .ZN(N2480) );
INV_X4 \add_1_root_add_519_2/U253  ( .A(\add_1_root_add_519_2/n45 ), .ZN(\add_1_root_add_519_2/n178 ) );
XNOR2_X2 \add_1_root_add_519_2/U252  ( .A(\add_1_root_add_519_2/n179 ), .B(\add_1_root_add_519_2/n178 ), .ZN(N2499) );
NAND2_X2 \add_1_root_add_519_2/U251  ( .A1(\add_1_root_add_519_2/n178 ),.A2(aad_byte_cnt[20]), .ZN(\add_1_root_add_519_2/n177 ) );
XNOR2_X2 \add_1_root_add_519_2/U250  ( .A(\add_1_root_add_519_2/n177 ), .B(aad_byte_cnt[21]), .ZN(N2500) );
XNOR2_X2 \add_1_root_add_519_2/U249  ( .A(\add_1_root_add_519_2/n52 ), .B(aad_byte_cnt[22]), .ZN(N2501) );
XNOR2_X2 \add_1_root_add_519_2/U248  ( .A(\add_1_root_add_519_2/n27 ), .B(aad_byte_cnt[23]), .ZN(N2502) );
XNOR2_X2 \add_1_root_add_519_2/U247  ( .A(\add_1_root_add_519_2/n43 ), .B(aad_byte_cnt[24]), .ZN(N2503) );
XNOR2_X2 \add_1_root_add_519_2/U246  ( .A(\add_1_root_add_519_2/n50 ), .B(aad_byte_cnt[25]), .ZN(N2504) );
XNOR2_X2 \add_1_root_add_519_2/U245  ( .A(\add_1_root_add_519_2/n51 ), .B(aad_byte_cnt[26]), .ZN(N2505) );
INV_X4 \add_1_root_add_519_2/U244  ( .A(aad_byte_cnt[27]), .ZN(\add_1_root_add_519_2/n172 ) );
XNOR2_X2 \add_1_root_add_519_2/U243  ( .A(\add_1_root_add_519_2/n28 ), .B(aad_byte_cnt[27]), .ZN(N2506) );
INV_X4 \add_1_root_add_519_2/U242  ( .A(aad_byte_cnt[28]), .ZN(\add_1_root_add_519_2/n159 ) );
XNOR2_X2 \add_1_root_add_519_2/U241  ( .A(\add_1_root_add_519_2/n47 ), .B(aad_byte_cnt[28]), .ZN(N2507) );
INV_X4 \add_1_root_add_519_2/U240  ( .A(aad_byte_cnt[29]), .ZN(\add_1_root_add_519_2/n167 ) );
XNOR2_X2 \add_1_root_add_519_2/U239  ( .A(\add_1_root_add_519_2/n21 ), .B(aad_byte_cnt[29]), .ZN(N2508) );
NAND2_X2 \add_1_root_add_519_2/U238  ( .A1(\add_1_root_add_519_2/n60 ), .A2(\add_1_root_add_519_2/n142 ), .ZN(\add_1_root_add_519_2/n163 ) );
NAND2_X2 \add_1_root_add_519_2/U237  ( .A1(\add_1_root_add_519_2/n57 ), .A2(\add_1_root_add_519_2/n164 ), .ZN(\add_1_root_add_519_2/n143 ) );
INV_X4 \add_1_root_add_519_2/U236  ( .A(\add_1_root_add_519_2/n53 ), .ZN(\add_1_root_add_519_2/n161 ) );
INV_X4 \add_1_root_add_519_2/U235  ( .A(aad_byte_cnt[30]), .ZN(\add_1_root_add_519_2/n162 ) );
XNOR2_X2 \add_1_root_add_519_2/U234  ( .A(\add_1_root_add_519_2/n161 ), .B(\add_1_root_add_519_2/n162 ), .ZN(N2509) );
INV_X4 \add_1_root_add_519_2/U233  ( .A(aad_byte_cnt[31]), .ZN(\add_1_root_add_519_2/n160 ) );
XNOR2_X2 \add_1_root_add_519_2/U232  ( .A(\add_1_root_add_519_2/n17 ), .B(\add_1_root_add_519_2/n160 ), .ZN(N2510) );
INV_X4 \add_1_root_add_519_2/U231  ( .A(\add_1_root_add_519_2/n93 ), .ZN(\add_1_root_add_519_2/n148 ) );
INV_X4 \add_1_root_add_519_2/U230  ( .A(\add_1_root_add_519_2/n94 ), .ZN(\add_1_root_add_519_2/n147 ) );
NAND2_X2 \add_1_root_add_519_2/U229  ( .A1(\add_1_root_add_519_2/n148 ),.A2(\add_1_root_add_519_2/n147 ), .ZN(\add_1_root_add_519_2/n107 ) );
XNOR2_X2 \add_1_root_add_519_2/U228  ( .A(\add_1_root_add_519_2/n157 ), .B(aad_byte_cnt[32]), .ZN(N2511) );
XNOR2_X2 \add_1_root_add_519_2/U227  ( .A(\add_1_root_add_519_2/n34 ), .B(\add_1_root_add_519_2/n151 ), .ZN(N2512) );
XNOR2_X2 \add_1_root_add_519_2/U226  ( .A(\add_1_root_add_519_2/n3 ), .B(\add_1_root_add_519_2/n150 ), .ZN(N2513) );
INV_X4 \add_1_root_add_519_2/U225  ( .A(aad_byte_cnt[35]), .ZN(\add_1_root_add_519_2/n154 ) );
XNOR2_X2 \add_1_root_add_519_2/U224  ( .A(\add_1_root_add_519_2/n7 ), .B(\add_1_root_add_519_2/n154 ), .ZN(N2514) );
NAND2_X2 \add_1_root_add_519_2/U223  ( .A1(\add_1_root_add_519_2/n148 ),.A2(\add_1_root_add_519_2/n8 ), .ZN(\add_1_root_add_519_2/n145 ) );
INV_X4 \add_1_root_add_519_2/U222  ( .A(\add_1_root_add_519_2/n108 ), .ZN(\add_1_root_add_519_2/n78 ) );
NAND2_X2 \add_1_root_add_519_2/U221  ( .A1(\add_1_root_add_519_2/n78 ), .A2(\add_1_root_add_519_2/n147 ), .ZN(\add_1_root_add_519_2/n146 ) );
XNOR2_X2 \add_1_root_add_519_2/U220  ( .A(\add_1_root_add_519_2/n2 ), .B(aad_byte_cnt[36]), .ZN(N2515) );
XNOR2_X2 \add_1_root_add_519_2/U219  ( .A(\add_1_root_add_519_2/n39 ), .B(aad_byte_cnt[37]), .ZN(N2516) );
XNOR2_X2 \add_1_root_add_519_2/U218  ( .A(\add_1_root_add_519_2/n54 ), .B(aad_byte_cnt[38]), .ZN(N2517) );
INV_X4 \add_1_root_add_519_2/U217  ( .A(aad_byte_cnt[39]), .ZN(\add_1_root_add_519_2/n144 ) );
XNOR2_X2 \add_1_root_add_519_2/U216  ( .A(\add_1_root_add_519_2/n38 ), .B(aad_byte_cnt[39]), .ZN(N2518) );
NAND2_X2 \add_1_root_add_519_2/U215  ( .A1(\add_1_root_add_519_2/n143 ),.A2(\add_1_root_add_519_2/n60 ), .ZN(\add_1_root_add_519_2/n141 ) );
NAND2_X2 \add_1_root_add_519_2/U214  ( .A1(\add_1_root_add_519_2/n141 ),.A2(\add_1_root_add_519_2/n142 ), .ZN(\add_1_root_add_519_2/n137 ) );
NAND2_X2 \add_1_root_add_519_2/U213  ( .A1(\add_1_root_add_519_2/n139 ),.A2(\add_1_root_add_519_2/n140 ), .ZN(\add_1_root_add_519_2/n138 ) );
XNOR2_X2 \add_1_root_add_519_2/U212  ( .A(\add_1_root_add_519_2/n137 ), .B(\add_1_root_add_519_2/n138 ), .ZN(N2482) );
INV_X4 \add_1_root_add_519_2/U211  ( .A(\add_1_root_add_519_2/n111 ), .ZN(\add_1_root_add_519_2/n132 ) );
NAND2_X2 \add_1_root_add_519_2/U210  ( .A1(\add_1_root_add_519_2/n132 ),.A2(\add_1_root_add_519_2/n8 ), .ZN(\add_1_root_add_519_2/n131 ) );
XNOR2_X2 \add_1_root_add_519_2/U209  ( .A(\add_1_root_add_519_2/n24 ), .B(aad_byte_cnt[40]), .ZN(N2519) );
INV_X4 \add_1_root_add_519_2/U208  ( .A(\add_1_root_add_519_2/n131 ), .ZN(\add_1_root_add_519_2/n124 ) );
NAND2_X2 \add_1_root_add_519_2/U207  ( .A1(\add_1_root_add_519_2/n124 ),.A2(aad_byte_cnt[40]), .ZN(\add_1_root_add_519_2/n130 ) );
XNOR2_X2 \add_1_root_add_519_2/U206  ( .A(\add_1_root_add_519_2/n23 ), .B(aad_byte_cnt[41]), .ZN(N2520) );
INV_X4 \add_1_root_add_519_2/U205  ( .A(\add_1_root_add_519_2/n130 ), .ZN(\add_1_root_add_519_2/n129 ) );
XNOR2_X2 \add_1_root_add_519_2/U204  ( .A(\add_1_root_add_519_2/n128 ), .B(aad_byte_cnt[42]), .ZN(N2521) );
INV_X4 \add_1_root_add_519_2/U203  ( .A(aad_byte_cnt[43]), .ZN(\add_1_root_add_519_2/n126 ) );
XNOR2_X2 \add_1_root_add_519_2/U202  ( .A(\add_1_root_add_519_2/n26 ), .B(\add_1_root_add_519_2/n126 ), .ZN(N2522) );
NAND4_X2 \add_1_root_add_519_2/U201  ( .A1(aad_byte_cnt[43]), .A2(aad_byte_cnt[42]), .A3(aad_byte_cnt[40]), .A4(aad_byte_cnt[41]), .ZN(\add_1_root_add_519_2/n112 ) );
INV_X4 \add_1_root_add_519_2/U200  ( .A(\add_1_root_add_519_2/n112 ), .ZN(\add_1_root_add_519_2/n125 ) );
NAND2_X2 \add_1_root_add_519_2/U199  ( .A1(\add_1_root_add_519_2/n124 ),.A2(\add_1_root_add_519_2/n125 ), .ZN(\add_1_root_add_519_2/n122 ) );
INV_X4 \add_1_root_add_519_2/U198  ( .A(aad_byte_cnt[44]), .ZN(\add_1_root_add_519_2/n123 ) );
XNOR2_X2 \add_1_root_add_519_2/U197  ( .A(\add_1_root_add_519_2/n36 ), .B(aad_byte_cnt[44]), .ZN(N2523) );
INV_X4 \add_1_root_add_519_2/U196  ( .A(\add_1_root_add_519_2/n122 ), .ZN(\add_1_root_add_519_2/n121 ) );
NAND2_X2 \add_1_root_add_519_2/U195  ( .A1(\add_1_root_add_519_2/n121 ),.A2(aad_byte_cnt[44]), .ZN(\add_1_root_add_519_2/n119 ) );
INV_X4 \add_1_root_add_519_2/U194  ( .A(aad_byte_cnt[45]), .ZN(\add_1_root_add_519_2/n120 ) );
XNOR2_X2 \add_1_root_add_519_2/U193  ( .A(\add_1_root_add_519_2/n22 ), .B(aad_byte_cnt[45]), .ZN(N2524) );
INV_X4 \add_1_root_add_519_2/U192  ( .A(\add_1_root_add_519_2/n119 ), .ZN(\add_1_root_add_519_2/n118 ) );
INV_X4 \add_1_root_add_519_2/U191  ( .A(aad_byte_cnt[46]), .ZN(\add_1_root_add_519_2/n117 ) );
XNOR2_X2 \add_1_root_add_519_2/U190  ( .A(\add_1_root_add_519_2/n116 ), .B(\add_1_root_add_519_2/n117 ), .ZN(N2525) );
INV_X4 \add_1_root_add_519_2/U189  ( .A(aad_byte_cnt[47]), .ZN(\add_1_root_add_519_2/n115 ) );
XNOR2_X2 \add_1_root_add_519_2/U188  ( .A(\add_1_root_add_519_2/n25 ), .B(\add_1_root_add_519_2/n115 ), .ZN(N2526) );
NAND2_X2 \add_1_root_add_519_2/U187  ( .A1(aad_byte_cnt[47]), .A2(aad_byte_cnt[46]), .ZN(\add_1_root_add_519_2/n113 ) );
XNOR2_X2 \add_1_root_add_519_2/U186  ( .A(\add_1_root_add_519_2/n20 ), .B(aad_byte_cnt[48]), .ZN(N2527) );
INV_X4 \add_1_root_add_519_2/U185  ( .A(\add_1_root_add_519_2/n105 ), .ZN(\add_1_root_add_519_2/n92 ) );
INV_X4 \add_1_root_add_519_2/U184  ( .A(\add_1_root_add_519_2/n55 ), .ZN(\add_1_root_add_519_2/n104 ) );
XNOR2_X2 \add_1_root_add_519_2/U183  ( .A(\add_1_root_add_519_2/n104 ), .B(\add_1_root_add_519_2/n101 ), .ZN(N2528) );
XNOR2_X2 \add_1_root_add_519_2/U182  ( .A(\add_1_root_add_519_2/n103 ), .B(\add_1_root_add_519_2/n80 ), .ZN(N2483) );
INV_X4 \add_1_root_add_519_2/U181  ( .A(aad_byte_cnt[49]), .ZN(\add_1_root_add_519_2/n101 ) );
INV_X4 \add_1_root_add_519_2/U180  ( .A(aad_byte_cnt[50]), .ZN(\add_1_root_add_519_2/n102 ) );
XNOR2_X2 \add_1_root_add_519_2/U179  ( .A(\add_1_root_add_519_2/n37 ), .B(\add_1_root_add_519_2/n102 ), .ZN(N2529) );
INV_X4 \add_1_root_add_519_2/U178  ( .A(\add_1_root_add_519_2/n99 ), .ZN(\add_1_root_add_519_2/n100 ) );
XNOR2_X2 \add_1_root_add_519_2/U177  ( .A(\add_1_root_add_519_2/n12 ), .B(aad_byte_cnt[51]), .ZN(N2530) );
NAND2_X2 \add_1_root_add_519_2/U176  ( .A1(\add_1_root_add_519_2/n99 ), .A2(aad_byte_cnt[51]), .ZN(\add_1_root_add_519_2/n98 ) );
XNOR2_X2 \add_1_root_add_519_2/U175  ( .A(\add_1_root_add_519_2/n11 ), .B(aad_byte_cnt[52]), .ZN(N2531) );
INV_X4 \add_1_root_add_519_2/U174  ( .A(\add_1_root_add_519_2/n98 ), .ZN(\add_1_root_add_519_2/n97 ) );
NAND2_X2 \add_1_root_add_519_2/U173  ( .A1(\add_1_root_add_519_2/n97 ), .A2(aad_byte_cnt[52]), .ZN(\add_1_root_add_519_2/n96 ) );
XNOR2_X2 \add_1_root_add_519_2/U172  ( .A(\add_1_root_add_519_2/n10 ), .B(aad_byte_cnt[53]), .ZN(N2532) );
INV_X4 \add_1_root_add_519_2/U171  ( .A(\add_1_root_add_519_2/n96 ), .ZN(\add_1_root_add_519_2/n77 ) );
NAND2_X2 \add_1_root_add_519_2/U170  ( .A1(\add_1_root_add_519_2/n77 ), .A2(\add_1_root_add_519_2/n78 ), .ZN(\add_1_root_add_519_2/n90 ) );
NAND2_X2 \add_1_root_add_519_2/U169  ( .A1(aad_byte_cnt[48]), .A2(aad_byte_cnt[53]), .ZN(\add_1_root_add_519_2/n95 ) );
NAND2_X2 \add_1_root_add_519_2/U168  ( .A1(\add_1_root_add_519_2/n91 ), .A2(\add_1_root_add_519_2/n92 ), .ZN(\add_1_root_add_519_2/n76 ) );
INV_X4 \add_1_root_add_519_2/U167  ( .A(aad_byte_cnt[54]), .ZN(\add_1_root_add_519_2/n89 ) );
XNOR2_X2 \add_1_root_add_519_2/U166  ( .A(\add_1_root_add_519_2/n1 ), .B(aad_byte_cnt[54]), .ZN(N2533) );
INV_X4 \add_1_root_add_519_2/U165  ( .A(aad_byte_cnt[55]), .ZN(\add_1_root_add_519_2/n88 ) );
XNOR2_X2 \add_1_root_add_519_2/U164  ( .A(\add_1_root_add_519_2/n35 ), .B(aad_byte_cnt[55]), .ZN(N2534) );
INV_X4 \add_1_root_add_519_2/U163  ( .A(\add_1_root_add_519_2/n86 ), .ZN(\add_1_root_add_519_2/n87 ) );
XNOR2_X2 \add_1_root_add_519_2/U162  ( .A(\add_1_root_add_519_2/n16 ), .B(aad_byte_cnt[56]), .ZN(N2535) );
NAND2_X2 \add_1_root_add_519_2/U161  ( .A1(\add_1_root_add_519_2/n86 ), .A2(aad_byte_cnt[56]), .ZN(\add_1_root_add_519_2/n85 ) );
XNOR2_X2 \add_1_root_add_519_2/U160  ( .A(\add_1_root_add_519_2/n15 ), .B(aad_byte_cnt[57]), .ZN(N2536) );
INV_X4 \add_1_root_add_519_2/U159  ( .A(\add_1_root_add_519_2/n85 ), .ZN(\add_1_root_add_519_2/n84 ) );
NAND2_X2 \add_1_root_add_519_2/U158  ( .A1(\add_1_root_add_519_2/n84 ), .A2(aad_byte_cnt[57]), .ZN(\add_1_root_add_519_2/n83 ) );
XNOR2_X2 \add_1_root_add_519_2/U157  ( .A(\add_1_root_add_519_2/n14 ), .B(aad_byte_cnt[58]), .ZN(N2537) );
INV_X4 \add_1_root_add_519_2/U156  ( .A(\add_1_root_add_519_2/n83 ), .ZN(\add_1_root_add_519_2/n82 ) );
NAND2_X2 \add_1_root_add_519_2/U155  ( .A1(\add_1_root_add_519_2/n82 ), .A2(aad_byte_cnt[58]), .ZN(\add_1_root_add_519_2/n74 ) );
XNOR2_X2 \add_1_root_add_519_2/U154  ( .A(\add_1_root_add_519_2/n13 ), .B(aad_byte_cnt[59]), .ZN(N2538) );
XNOR2_X2 \add_1_root_add_519_2/U153  ( .A(\add_1_root_add_519_2/n81 ), .B(\add_1_root_add_519_2/n18 ), .ZN(N2484) );
INV_X4 \add_1_root_add_519_2/U152  ( .A(aad_byte_cnt[60]), .ZN(\add_1_root_add_519_2/n79 ) );
NAND2_X2 \add_1_root_add_519_2/U151  ( .A1(\add_1_root_add_519_2/n77 ), .A2(\add_1_root_add_519_2/n78 ), .ZN(\add_1_root_add_519_2/n75 ) );
INV_X4 \add_1_root_add_519_2/U150  ( .A(\add_1_root_add_519_2/n74 ), .ZN(\add_1_root_add_519_2/n73 ) );
NAND2_X2 \add_1_root_add_519_2/U149  ( .A1(\add_1_root_add_519_2/n73 ), .A2(aad_byte_cnt[59]), .ZN(\add_1_root_add_519_2/n70 ) );
XNOR2_X2 \add_1_root_add_519_2/U148  ( .A(\add_1_root_add_519_2/n79 ), .B(\add_1_root_add_519_2/n19 ), .ZN(N2539) );
INV_X4 \add_1_root_add_519_2/U147  ( .A(aad_byte_cnt[61]), .ZN(\add_1_root_add_519_2/n72 ) );
XNOR2_X2 \add_1_root_add_519_2/U146  ( .A(\add_1_root_add_519_2/n31 ), .B(\add_1_root_add_519_2/n72 ), .ZN(N2540) );
INV_X4 \add_1_root_add_519_2/U145  ( .A(aad_byte_cnt[62]), .ZN(\add_1_root_add_519_2/n71 ) );
XNOR2_X2 \add_1_root_add_519_2/U144  ( .A(\add_1_root_add_519_2/n29 ), .B(\add_1_root_add_519_2/n71 ), .ZN(N2541) );
NAND2_X2 \add_1_root_add_519_2/U143  ( .A1(\add_1_root_add_519_2/n69 ), .A2(aad_byte_cnt[62]), .ZN(\add_1_root_add_519_2/n68 ) );
NAND2_X2 \add_1_root_add_519_2/U142  ( .A1(\add_1_root_add_519_2/n18 ), .A2(aad_byte_cnt[5]), .ZN(\add_1_root_add_519_2/n66 ) );
XNOR2_X2 \add_1_root_add_519_2/U141  ( .A(\add_1_root_add_519_2/n66 ), .B(aad_byte_cnt[6]), .ZN(N2485) );
XNOR2_X2 \add_1_root_add_519_2/U140  ( .A(\add_1_root_add_519_2/n33 ), .B(aad_byte_cnt[7]), .ZN(N2486) );
XNOR2_X2 \add_1_root_add_519_2/U139  ( .A(\add_1_root_add_519_2/n63 ), .B(\add_1_root_add_519_2/n64 ), .ZN(N2487) );
XNOR2_X2 \add_1_root_add_519_2/U138  ( .A(\add_1_root_add_519_2/n58 ), .B(aad_byte_cnt[9]), .ZN(N2488) );
INV_X4 \add_1_root_add_519_2/U137  ( .A(aad_byte_cnt[38]), .ZN(\add_1_root_add_519_2/n134 ) );
INV_X4 \add_1_root_add_519_2/U136  ( .A(aad_byte_cnt[37]), .ZN(\add_1_root_add_519_2/n136 ) );
INV_X4 \add_1_root_add_519_2/U135  ( .A(aad_byte_cnt[36]), .ZN(\add_1_root_add_519_2/n135 ) );
INV_X4 \add_1_root_add_519_2/U134  ( .A(aad_byte_cnt[34]), .ZN(\add_1_root_add_519_2/n150 ) );
INV_X4 \add_1_root_add_519_2/U133  ( .A(aad_byte_cnt[33]), .ZN(\add_1_root_add_519_2/n151 ) );
INV_X4 \add_1_root_add_519_2/U132  ( .A(aad_byte_cnt[32]), .ZN(\add_1_root_add_519_2/n156 ) );
INV_X4 \add_1_root_add_519_2/U131  ( .A(aad_byte_cnt[26]), .ZN(\add_1_root_add_519_2/n169 ) );
INV_X4 \add_1_root_add_519_2/U130  ( .A(aad_byte_cnt[25]), .ZN(\add_1_root_add_519_2/n171 ) );
INV_X4 \add_1_root_add_519_2/U129  ( .A(aad_byte_cnt[24]), .ZN(\add_1_root_add_519_2/n170 ) );
INV_X4 \add_1_root_add_519_2/U128  ( .A(aad_byte_cnt[23]), .ZN(\add_1_root_add_519_2/n175 ) );
INV_X4 \add_1_root_add_519_2/U127  ( .A(aad_byte_cnt[22]), .ZN(\add_1_root_add_519_2/n174 ) );
INV_X4 \add_1_root_add_519_2/U126  ( .A(aad_byte_cnt[21]), .ZN(\add_1_root_add_519_2/n176 ) );
INV_X4 \add_1_root_add_519_2/U125  ( .A(aad_byte_cnt[20]), .ZN(\add_1_root_add_519_2/n179 ) );
INV_X4 \add_1_root_add_519_2/U124  ( .A(aad_byte_cnt[18]), .ZN(\add_1_root_add_519_2/n181 ) );
INV_X4 \add_1_root_add_519_2/U123  ( .A(aad_byte_cnt[17]), .ZN(\add_1_root_add_519_2/n189 ) );
INV_X4 \add_1_root_add_519_2/U122  ( .A(aad_byte_cnt[16]), .ZN(\add_1_root_add_519_2/n182 ) );
INV_X4 \add_1_root_add_519_2/U121  ( .A(aad_byte_cnt[10]), .ZN(\add_1_root_add_519_2/n206 ) );
INV_X4 \add_1_root_add_519_2/U120  ( .A(aad_byte_cnt[9]), .ZN(\add_1_root_add_519_2/n62 ) );
INV_X4 \add_1_root_add_519_2/U119  ( .A(aad_byte_cnt[8]), .ZN(\add_1_root_add_519_2/n64 ) );
INV_X4 \add_1_root_add_519_2/U118  ( .A(aad_byte_cnt[6]), .ZN(\add_1_root_add_519_2/n65 ) );
INV_X4 \add_1_root_add_519_2/U117  ( .A(aad_byte_cnt[4]), .ZN(\add_1_root_add_519_2/n103 ) );
INV_X4 \add_1_root_add_519_2/U116  ( .A(aad_byte_cnt[5]), .ZN(\add_1_root_add_519_2/n81 ) );
INV_X4 \add_1_root_add_519_2/U115  ( .A(\add_1_root_add_519_2/n186 ), .ZN(\add_1_root_add_519_2/n210 ) );
INV_X4 \add_1_root_add_519_2/U114  ( .A(\add_1_root_add_519_2/n114 ), .ZN(\add_1_root_add_519_2/n157 ) );
INV_X4 \add_1_root_add_519_2/U113  ( .A(\add_1_root_add_519_2/n127 ), .ZN(\add_1_root_add_519_2/n128 ) );
INV_X4 \add_1_root_add_519_2/U112  ( .A(\add_1_root_add_519_2/n208 ), .ZN(\add_1_root_add_519_2/n63 ) );
OR2_X2 \add_1_root_add_519_2/U111  ( .A1(aad_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(\add_1_root_add_519_2/n60 ) );
NOR2_X2 \add_1_root_add_519_2/U110  ( .A1(\add_1_root_add_519_2/n48 ), .A2(\add_1_root_add_519_2/n68 ), .ZN(\add_1_root_add_519_2/n67 ) );
XOR2_X2 \add_1_root_add_519_2/U109  ( .A(\add_1_root_add_519_2/n67 ), .B(aad_byte_cnt[63]), .Z(N2542) );
AND2_X2 \add_1_root_add_519_2/U108  ( .A1(aad_byte_cnt[0]), .A2(n17750),.ZN(\add_1_root_add_519_2/n219 ) );
NOR2_X2 \add_1_root_add_519_2/U107  ( .A1(\add_1_root_add_519_2/n217 ), .A2(\add_1_root_add_519_2/n218 ), .ZN(\add_1_root_add_519_2/n216 ) );
NAND3_X2 \add_1_root_add_519_2/U106  ( .A1(dii_data_size[1]), .A2(\add_1_root_add_519_2/n60 ), .A3(aad_byte_cnt[1]), .ZN(\add_1_root_add_519_2/n215 ) );
NAND3_X2 \add_1_root_add_519_2/U105  ( .A1(\add_1_root_add_519_2/n214 ),.A2(\add_1_root_add_519_2/n215 ), .A3(\add_1_root_add_519_2/n216 ),.ZN(\add_1_root_add_519_2/n193 ) );
NOR2_X2 \add_1_root_add_519_2/U104  ( .A1(aad_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(\add_1_root_add_519_2/n222 ) );
NOR2_X2 \add_1_root_add_519_2/U103  ( .A1(aad_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(\add_1_root_add_519_2/n221 ) );
NOR2_X2 \add_1_root_add_519_2/U102  ( .A1(\add_1_root_add_519_2/n221 ), .A2(\add_1_root_add_519_2/n222 ), .ZN(\add_1_root_add_519_2/n220 ) );
NOR2_X2 \add_1_root_add_519_2/U101  ( .A1(aad_byte_cnt[0]), .A2(n17750),.ZN(\add_1_root_add_519_2/n186 ) );
NOR2_X2 \add_1_root_add_519_2/U100  ( .A1(aad_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(\add_1_root_add_519_2/n165 ) );
INV_X4 \add_1_root_add_519_2/U99  ( .A(n18074), .ZN(\add_1_root_add_519_2/n61 ) );
AND2_X2 \add_1_root_add_519_2/U98  ( .A1(\add_1_root_add_519_2/n186 ), .A2(\add_1_root_add_519_2/n185 ), .ZN(\add_1_root_add_519_2/n166 ) );
NOR2_X2 \add_1_root_add_519_2/U97  ( .A1(\add_1_root_add_519_2/n154 ), .A2(\add_1_root_add_519_2/n150 ), .ZN(\add_1_root_add_519_2/n149 ) );
OR2_X2 \add_1_root_add_519_2/U96  ( .A1(\add_1_root_add_519_2/n58 ), .A2(\add_1_root_add_519_2/n62 ), .ZN(\add_1_root_add_519_2/n59 ) );
NOR2_X2 \add_1_root_add_519_2/U95  ( .A1(\add_1_root_add_519_2/n134 ), .A2(\add_1_root_add_519_2/n144 ), .ZN(\add_1_root_add_519_2/n133 ) );
NAND3_X2 \add_1_root_add_519_2/U94  ( .A1(aad_byte_cnt[37]), .A2(aad_byte_cnt[36]), .A3(\add_1_root_add_519_2/n133 ), .ZN(\add_1_root_add_519_2/n111 ) );
OR2_X2 \add_1_root_add_519_2/U93  ( .A1(\add_1_root_add_519_2/n208 ), .A2(\add_1_root_add_519_2/n64 ), .ZN(\add_1_root_add_519_2/n58 ) );
NOR2_X2 \add_1_root_add_519_2/U92  ( .A1(\add_1_root_add_519_2/n167 ), .A2(\add_1_root_add_519_2/n159 ), .ZN(\add_1_root_add_519_2/n158 ) );
NAND3_X2 \add_1_root_add_519_2/U91  ( .A1(aad_byte_cnt[30]), .A2(aad_byte_cnt[31]), .A3(\add_1_root_add_519_2/n158 ), .ZN(\add_1_root_add_519_2/n93 ) );
NOR2_X2 \add_1_root_add_519_2/U90  ( .A1(\add_1_root_add_519_2/n184 ), .A2(\add_1_root_add_519_2/n165 ), .ZN(\add_1_root_add_519_2/n183 ) );
NOR2_X2 \add_1_root_add_519_2/U89  ( .A1(\add_1_root_add_519_2/n151 ), .A2(\add_1_root_add_519_2/n156 ), .ZN(\add_1_root_add_519_2/n155 ) );
AND2_X2 \add_1_root_add_519_2/U88  ( .A1(aad_byte_cnt[61]), .A2(aad_byte_cnt[60]), .ZN(\add_1_root_add_519_2/n69 ) );
NOR2_X2 \add_1_root_add_519_2/U87  ( .A1(\add_1_root_add_519_2/n169 ), .A2(\add_1_root_add_519_2/n172 ), .ZN(\add_1_root_add_519_2/n168 ) );
NAND3_X2 \add_1_root_add_519_2/U86  ( .A1(aad_byte_cnt[25]), .A2(aad_byte_cnt[24]), .A3(\add_1_root_add_519_2/n168 ), .ZN(\add_1_root_add_519_2/n94 ) );
NOR2_X2 \add_1_root_add_519_2/U85  ( .A1(\add_1_root_add_519_2/n102 ), .A2(\add_1_root_add_519_2/n101 ), .ZN(\add_1_root_add_519_2/n99 ) );
NOR2_X2 \add_1_root_add_519_2/U84  ( .A1(\add_1_root_add_519_2/n88 ), .A2(\add_1_root_add_519_2/n89 ), .ZN(\add_1_root_add_519_2/n86 ) );
NOR2_X2 \add_1_root_add_519_2/U83  ( .A1(\add_1_root_add_519_2/n187 ), .A2(\add_1_root_add_519_2/n181 ), .ZN(\add_1_root_add_519_2/n180 ) );
NAND3_X2 \add_1_root_add_519_2/U82  ( .A1(aad_byte_cnt[16]), .A2(aad_byte_cnt[17]), .A3(\add_1_root_add_519_2/n180 ), .ZN(\add_1_root_add_519_2/n153 ) );
NOR2_X2 \add_1_root_add_519_2/U81  ( .A1(\add_1_root_add_519_2/n174 ), .A2(\add_1_root_add_519_2/n175 ), .ZN(\add_1_root_add_519_2/n173 ) );
NAND3_X2 \add_1_root_add_519_2/U80  ( .A1(aad_byte_cnt[21]), .A2(aad_byte_cnt[20]), .A3(\add_1_root_add_519_2/n173 ), .ZN(\add_1_root_add_519_2/n108 ) );
OR2_X2 \add_1_root_add_519_2/U79  ( .A1(\add_1_root_add_519_2/n165 ), .A2(\add_1_root_add_519_2/n166 ), .ZN(\add_1_root_add_519_2/n57 ) );
NOR3_X2 \add_1_root_add_519_2/U78  ( .A1(\add_1_root_add_519_2/n93 ), .A2(\add_1_root_add_519_2/n94 ), .A3(\add_1_root_add_519_2/n95 ), .ZN(\add_1_root_add_519_2/n91 ) );
AND2_X4 \add_1_root_add_519_2/U77  ( .A1(\add_1_root_add_519_2/n92 ), .A2(aad_byte_cnt[48]), .ZN(\add_1_root_add_519_2/n56 ) );
NAND2_X2 \add_1_root_add_519_2/U76  ( .A1(\add_1_root_add_519_2/n106 ), .A2(\add_1_root_add_519_2/n56 ), .ZN(\add_1_root_add_519_2/n55 ) );
NOR2_X2 \add_1_root_add_519_2/U75  ( .A1(\add_1_root_add_519_2/n212 ), .A2(\add_1_root_add_519_2/n165 ), .ZN(\add_1_root_add_519_2/n211 ) );
NAND3_X2 \add_1_root_add_519_2/U74  ( .A1(\add_1_root_add_519_2/n210 ), .A2(\add_1_root_add_519_2/n60 ), .A3(\add_1_root_add_519_2/n211 ), .ZN(\add_1_root_add_519_2/n200 ) );
OR3_X2 \add_1_root_add_519_2/U73  ( .A1(\add_1_root_add_519_2/n2 ), .A2(\add_1_root_add_519_2/n135 ), .A3(\add_1_root_add_519_2/n136 ), .ZN(\add_1_root_add_519_2/n54 ) );
OR3_X2 \add_1_root_add_519_2/U72  ( .A1(\add_1_root_add_519_2/n47 ), .A2(\add_1_root_add_519_2/n167 ), .A3(\add_1_root_add_519_2/n159 ), .ZN(\add_1_root_add_519_2/n53 ) );
NOR2_X2 \add_1_root_add_519_2/U71  ( .A1(\add_1_root_add_519_2/n65 ), .A2(\add_1_root_add_519_2/n224 ), .ZN(\add_1_root_add_519_2/n223 ) );
NAND3_X2 \add_1_root_add_519_2/U70  ( .A1(aad_byte_cnt[5]), .A2(aad_byte_cnt[4]), .A3(\add_1_root_add_519_2/n223 ), .ZN(\add_1_root_add_519_2/n198 ) );
OR2_X2 \add_1_root_add_519_2/U69  ( .A1(\add_1_root_add_519_2/n176 ), .A2(\add_1_root_add_519_2/n177 ), .ZN(\add_1_root_add_519_2/n52 ) );
OR2_X2 \add_1_root_add_519_2/U68  ( .A1(\add_1_root_add_519_2/n171 ), .A2(\add_1_root_add_519_2/n50 ), .ZN(\add_1_root_add_519_2/n51 ) );
OR2_X2 \add_1_root_add_519_2/U67  ( .A1(\add_1_root_add_519_2/n170 ), .A2(\add_1_root_add_519_2/n43 ), .ZN(\add_1_root_add_519_2/n50 ) );
AND2_X2 \add_1_root_add_519_2/U66  ( .A1(aad_byte_cnt[13]), .A2(aad_byte_cnt[12]), .ZN(\add_1_root_add_519_2/n199 ) );
AND2_X4 \add_1_root_add_519_2/U65  ( .A1(\add_1_root_add_519_2/n118 ), .A2(aad_byte_cnt[45]), .ZN(\add_1_root_add_519_2/n49 ) );
AND2_X2 \add_1_root_add_519_2/U64  ( .A1(\add_1_root_add_519_2/n114 ), .A2(\add_1_root_add_519_2/n49 ), .ZN(\add_1_root_add_519_2/n116 ) );
NOR2_X2 \add_1_root_add_519_2/U63  ( .A1(\add_1_root_add_519_2/n206 ), .A2(\add_1_root_add_519_2/n207 ), .ZN(\add_1_root_add_519_2/n205 ) );
NAND3_X2 \add_1_root_add_519_2/U62  ( .A1(aad_byte_cnt[9]), .A2(aad_byte_cnt[8]), .A3(\add_1_root_add_519_2/n205 ), .ZN(\add_1_root_add_519_2/n192 ) );
NAND3_X2 \add_1_root_add_519_2/U61  ( .A1(\add_1_root_add_519_2/n140 ), .A2(\add_1_root_add_519_2/n193 ), .A3(\add_1_root_add_519_2/n194 ), .ZN(\add_1_root_add_519_2/n190 ) );
NOR2_X2 \add_1_root_add_519_2/U60  ( .A1(\add_1_root_add_519_2/n111 ), .A2(\add_1_root_add_519_2/n112 ), .ZN(\add_1_root_add_519_2/n110 ) );
NOR3_X2 \add_1_root_add_519_2/U59  ( .A1(\add_1_root_add_519_2/n113 ), .A2(\add_1_root_add_519_2/n120 ), .A3(\add_1_root_add_519_2/n123 ), .ZN(\add_1_root_add_519_2/n109 ) );
NAND3_X2 \add_1_root_add_519_2/U58  ( .A1(\add_1_root_add_519_2/n109 ), .A2(\add_1_root_add_519_2/n8 ), .A3(\add_1_root_add_519_2/n110 ), .ZN(\add_1_root_add_519_2/n105 ) );
AND2_X2 \add_1_root_add_519_2/U57  ( .A1(\add_1_root_add_519_2/n195 ), .A2(\add_1_root_add_519_2/n42 ), .ZN(\add_1_root_add_519_2/n152 ) );
OR2_X2 \add_1_root_add_519_2/U56  ( .A1(\add_1_root_add_519_2/n1 ), .A2(\add_1_root_add_519_2/n70 ), .ZN(\add_1_root_add_519_2/n48 ) );
NOR2_X2 \add_1_root_add_519_2/U55  ( .A1(\add_1_root_add_519_2/n198 ), .A2(\add_1_root_add_519_2/n191 ), .ZN(\add_1_root_add_519_2/n197 ) );
NOR2_X2 \add_1_root_add_519_2/U54  ( .A1(\add_1_root_add_519_2/n192 ), .A2(\add_1_root_add_519_2/n200 ), .ZN(\add_1_root_add_519_2/n196 ) );
OR2_X2 \add_1_root_add_519_2/U53  ( .A1(\add_1_root_add_519_2/n43 ), .A2(\add_1_root_add_519_2/n94 ), .ZN(\add_1_root_add_519_2/n47 ) );
OR2_X2 \add_1_root_add_519_2/U52  ( .A1(\add_1_root_add_519_2/n152 ), .A2(\add_1_root_add_519_2/n153 ), .ZN(\add_1_root_add_519_2/n46 ) );
OR2_X2 \add_1_root_add_519_2/U51  ( .A1(\add_1_root_add_519_2/n152 ), .A2(\add_1_root_add_519_2/n153 ), .ZN(\add_1_root_add_519_2/n45 ) );
AND2_X4 \add_1_root_add_519_2/U50  ( .A1(\add_1_root_add_519_2/n129 ), .A2(aad_byte_cnt[41]), .ZN(\add_1_root_add_519_2/n44 ) );
AND2_X2 \add_1_root_add_519_2/U49  ( .A1(\add_1_root_add_519_2/n114 ), .A2(\add_1_root_add_519_2/n44 ), .ZN(\add_1_root_add_519_2/n127 ) );
OR3_X2 \add_1_root_add_519_2/U48  ( .A1(\add_1_root_add_519_2/n152 ), .A2(\add_1_root_add_519_2/n153 ), .A3(\add_1_root_add_519_2/n108 ), .ZN(\add_1_root_add_519_2/n43 ) );
NOR3_X2 \add_1_root_add_519_2/U47  ( .A1(\add_1_root_add_519_2/n46 ), .A2(\add_1_root_add_519_2/n107 ), .A3(\add_1_root_add_519_2/n108 ), .ZN(\add_1_root_add_519_2/n106 ) );
NOR3_X2 \add_1_root_add_519_2/U46  ( .A1(\add_1_root_add_519_2/n107 ), .A2(\add_1_root_add_519_2/n45 ), .A3(\add_1_root_add_519_2/n108 ), .ZN(\add_1_root_add_519_2/n114 ) );
XNOR2_X1 \add_1_root_add_519_2/U45  ( .A(\add_1_root_add_519_2/n163 ), .B(\add_1_root_add_519_2/n143 ), .ZN(N2481) );
OR3_X4 \add_1_root_add_519_2/U44  ( .A1(\add_1_root_add_519_2/n190 ), .A2(\add_1_root_add_519_2/n191 ), .A3(\add_1_root_add_519_2/n192 ), .ZN(\add_1_root_add_519_2/n42 ) );
OR3_X4 \add_1_root_add_519_2/U43  ( .A1(\add_1_root_add_519_2/n46 ), .A2(\add_1_root_add_519_2/n75 ), .A3(\add_1_root_add_519_2/n76 ), .ZN(\add_1_root_add_519_2/n41 ) );
OR2_X4 \add_1_root_add_519_2/U42  ( .A1(\add_1_root_add_519_2/n181 ), .A2(\add_1_root_add_519_2/n188 ), .ZN(\add_1_root_add_519_2/n40 ) );
OR2_X4 \add_1_root_add_519_2/U41  ( .A1(\add_1_root_add_519_2/n135 ), .A2(\add_1_root_add_519_2/n2 ), .ZN(\add_1_root_add_519_2/n39 ) );
OR2_X4 \add_1_root_add_519_2/U40  ( .A1(\add_1_root_add_519_2/n134 ), .A2(\add_1_root_add_519_2/n54 ), .ZN(\add_1_root_add_519_2/n38 ) );
NOR2_X2 \add_1_root_add_519_2/U39  ( .A1(\add_1_root_add_519_2/n101 ), .A2(\add_1_root_add_519_2/n55 ), .ZN(\add_1_root_add_519_2/n37 ) );
OR2_X4 \add_1_root_add_519_2/U38  ( .A1(\add_1_root_add_519_2/n157 ), .A2(\add_1_root_add_519_2/n122 ), .ZN(\add_1_root_add_519_2/n36 ) );
OR2_X4 \add_1_root_add_519_2/U37  ( .A1(\add_1_root_add_519_2/n89 ), .A2(\add_1_root_add_519_2/n1 ), .ZN(\add_1_root_add_519_2/n35 ) );
AND2_X4 \add_1_root_add_519_2/U36  ( .A1(\add_1_root_add_519_2/n114 ), .A2(aad_byte_cnt[32]), .ZN(\add_1_root_add_519_2/n34 ) );
OR2_X4 \add_1_root_add_519_2/U35  ( .A1(\add_1_root_add_519_2/n65 ), .A2(\add_1_root_add_519_2/n66 ), .ZN(\add_1_root_add_519_2/n33 ) );
OR2_X4 \add_1_root_add_519_2/U34  ( .A1(\add_1_root_add_519_2/n206 ), .A2(\add_1_root_add_519_2/n59 ), .ZN(\add_1_root_add_519_2/n32 ) );
AND2_X4 \add_1_root_add_519_2/U33  ( .A1(aad_byte_cnt[60]), .A2(\add_1_root_add_519_2/n19 ), .ZN(\add_1_root_add_519_2/n31 ) );
AND2_X4 \add_1_root_add_519_2/U32  ( .A1(aad_byte_cnt[14]), .A2(\add_1_root_add_519_2/n9 ), .ZN(\add_1_root_add_519_2/n30 ) );
AND2_X4 \add_1_root_add_519_2/U31  ( .A1(\add_1_root_add_519_2/n69 ), .A2(\add_1_root_add_519_2/n19 ), .ZN(\add_1_root_add_519_2/n29 ) );
OR2_X4 \add_1_root_add_519_2/U30  ( .A1(\add_1_root_add_519_2/n169 ), .A2(\add_1_root_add_519_2/n51 ), .ZN(\add_1_root_add_519_2/n28 ) );
OR2_X4 \add_1_root_add_519_2/U29  ( .A1(\add_1_root_add_519_2/n174 ), .A2(\add_1_root_add_519_2/n52 ), .ZN(\add_1_root_add_519_2/n27 ) );
AND2_X4 \add_1_root_add_519_2/U28  ( .A1(\add_1_root_add_519_2/n127 ), .A2(aad_byte_cnt[42]), .ZN(\add_1_root_add_519_2/n26 ) );
AND2_X4 \add_1_root_add_519_2/U27  ( .A1(\add_1_root_add_519_2/n116 ), .A2(aad_byte_cnt[46]), .ZN(\add_1_root_add_519_2/n25 ) );
OR2_X4 \add_1_root_add_519_2/U26  ( .A1(\add_1_root_add_519_2/n157 ), .A2(\add_1_root_add_519_2/n131 ), .ZN(\add_1_root_add_519_2/n24 ) );
OR2_X4 \add_1_root_add_519_2/U25  ( .A1(\add_1_root_add_519_2/n157 ), .A2(\add_1_root_add_519_2/n130 ), .ZN(\add_1_root_add_519_2/n23 ) );
OR2_X4 \add_1_root_add_519_2/U24  ( .A1(\add_1_root_add_519_2/n157 ), .A2(\add_1_root_add_519_2/n119 ), .ZN(\add_1_root_add_519_2/n22 ) );
OR2_X4 \add_1_root_add_519_2/U23  ( .A1(\add_1_root_add_519_2/n159 ), .A2(\add_1_root_add_519_2/n47 ), .ZN(\add_1_root_add_519_2/n21 ) );
OR2_X4 \add_1_root_add_519_2/U22  ( .A1(\add_1_root_add_519_2/n157 ), .A2(\add_1_root_add_519_2/n105 ), .ZN(\add_1_root_add_519_2/n20 ) );
NOR2_X2 \add_1_root_add_519_2/U21  ( .A1(\add_1_root_add_519_2/n41 ), .A2(\add_1_root_add_519_2/n70 ), .ZN(\add_1_root_add_519_2/n19 ) );
AND2_X4 \add_1_root_add_519_2/U20  ( .A1(aad_byte_cnt[4]), .A2(\add_1_root_add_519_2/n80 ), .ZN(\add_1_root_add_519_2/n18 ) );
NOR2_X2 \add_1_root_add_519_2/U19  ( .A1(\add_1_root_add_519_2/n162 ), .A2(\add_1_root_add_519_2/n53 ), .ZN(\add_1_root_add_519_2/n17 ) );
OR2_X4 \add_1_root_add_519_2/U18  ( .A1(\add_1_root_add_519_2/n1 ), .A2(\add_1_root_add_519_2/n87 ), .ZN(\add_1_root_add_519_2/n16 ) );
OR2_X4 \add_1_root_add_519_2/U17  ( .A1(\add_1_root_add_519_2/n1 ), .A2(\add_1_root_add_519_2/n85 ), .ZN(\add_1_root_add_519_2/n15 ) );
OR2_X4 \add_1_root_add_519_2/U16  ( .A1(\add_1_root_add_519_2/n1 ), .A2(\add_1_root_add_519_2/n83 ), .ZN(\add_1_root_add_519_2/n14 ) );
OR2_X4 \add_1_root_add_519_2/U15  ( .A1(\add_1_root_add_519_2/n1 ), .A2(\add_1_root_add_519_2/n74 ), .ZN(\add_1_root_add_519_2/n13 ) );
OR2_X4 \add_1_root_add_519_2/U14  ( .A1(\add_1_root_add_519_2/n55 ), .A2(\add_1_root_add_519_2/n100 ), .ZN(\add_1_root_add_519_2/n12 ) );
OR2_X4 \add_1_root_add_519_2/U13  ( .A1(\add_1_root_add_519_2/n55 ), .A2(\add_1_root_add_519_2/n98 ), .ZN(\add_1_root_add_519_2/n11 ) );
OR2_X4 \add_1_root_add_519_2/U12  ( .A1(\add_1_root_add_519_2/n55 ), .A2(\add_1_root_add_519_2/n96 ), .ZN(\add_1_root_add_519_2/n10 ) );
AND2_X4 \add_1_root_add_519_2/U11  ( .A1(\add_1_root_add_519_2/n6 ), .A2(aad_byte_cnt[13]), .ZN(\add_1_root_add_519_2/n9 ) );
AND3_X4 \add_1_root_add_519_2/U10  ( .A1(aad_byte_cnt[32]), .A2(aad_byte_cnt[33]), .A3(\add_1_root_add_519_2/n149 ), .ZN(\add_1_root_add_519_2/n8 ) );
AND2_X4 \add_1_root_add_519_2/U9  ( .A1(\add_1_root_add_519_2/n3 ), .A2(aad_byte_cnt[34]), .ZN(\add_1_root_add_519_2/n7 ) );
AND2_X4 \add_1_root_add_519_2/U8  ( .A1(\add_1_root_add_519_2/n5 ), .A2(aad_byte_cnt[12]), .ZN(\add_1_root_add_519_2/n6 ) );
NOR2_X2 \add_1_root_add_519_2/U7  ( .A1(\add_1_root_add_519_2/n208 ), .A2(\add_1_root_add_519_2/n192 ), .ZN(\add_1_root_add_519_2/n5 ) );
NOR2_X2 \add_1_root_add_519_2/U6  ( .A1(\add_1_root_add_519_2/n152 ), .A2(\add_1_root_add_519_2/n182 ), .ZN(\add_1_root_add_519_2/n4 ) );
AND2_X4 \add_1_root_add_519_2/U5  ( .A1(\add_1_root_add_519_2/n114 ), .A2(\add_1_root_add_519_2/n155 ), .ZN(\add_1_root_add_519_2/n3 ) );
OR3_X4 \add_1_root_add_519_2/U4  ( .A1(\add_1_root_add_519_2/n46 ), .A2(\add_1_root_add_519_2/n145 ), .A3(\add_1_root_add_519_2/n146 ), .ZN(\add_1_root_add_519_2/n2 ) );
OR3_X4 \add_1_root_add_519_2/U3  ( .A1(\add_1_root_add_519_2/n46 ), .A2(\add_1_root_add_519_2/n90 ), .A3(\add_1_root_add_519_2/n76 ), .ZN(\add_1_root_add_519_2/n1 ) );
NAND3_X2 \add_1_root_add_519_2/U2  ( .A1(aad_byte_cnt[14]), .A2(aad_byte_cnt[15]), .A3(\add_1_root_add_519_2/n199 ), .ZN(\add_1_root_add_519_2/n191 ) );
INV_X4 \add_1_root_add_513_2/U289  ( .A(enc_byte_cnt[7]), .ZN(\add_1_root_add_513_2/n224 ) );
INV_X4 \add_1_root_add_513_2/U288  ( .A(\add_1_root_add_513_2/n198 ), .ZN(\add_1_root_add_513_2/n194 ) );
NAND2_X2 \add_1_root_add_513_2/U287  ( .A1(\add_1_root_add_513_2/n219 ),.A2(\add_1_root_add_513_2/n220 ), .ZN(\add_1_root_add_513_2/n214 ) );
NAND2_X2 \add_1_root_add_513_2/U286  ( .A1(dii_data_size[2]), .A2(enc_byte_cnt[2]), .ZN(\add_1_root_add_513_2/n142 ) );
INV_X4 \add_1_root_add_513_2/U285  ( .A(\add_1_root_add_513_2/n142 ), .ZN(\add_1_root_add_513_2/n217 ) );
NAND2_X2 \add_1_root_add_513_2/U284  ( .A1(n18074), .A2(enc_byte_cnt[3]),.ZN(\add_1_root_add_513_2/n139 ) );
INV_X4 \add_1_root_add_513_2/U283  ( .A(\add_1_root_add_513_2/n139 ), .ZN(\add_1_root_add_513_2/n218 ) );
INV_X4 \add_1_root_add_513_2/U282  ( .A(enc_byte_cnt[3]), .ZN(\add_1_root_add_513_2/n213 ) );
NAND2_X2 \add_1_root_add_513_2/U281  ( .A1(\add_1_root_add_513_2/n61 ), .A2(\add_1_root_add_513_2/n213 ), .ZN(\add_1_root_add_513_2/n140 ) );
NAND2_X2 \add_1_root_add_513_2/U280  ( .A1(\add_1_root_add_513_2/n193 ),.A2(\add_1_root_add_513_2/n140 ), .ZN(\add_1_root_add_513_2/n209 ) );
INV_X4 \add_1_root_add_513_2/U279  ( .A(\add_1_root_add_513_2/n140 ), .ZN(\add_1_root_add_513_2/n212 ) );
NAND2_X2 \add_1_root_add_513_2/U278  ( .A1(\add_1_root_add_513_2/n209 ),.A2(\add_1_root_add_513_2/n200 ), .ZN(\add_1_root_add_513_2/n80 ) );
NAND2_X2 \add_1_root_add_513_2/U277  ( .A1(\add_1_root_add_513_2/n194 ),.A2(\add_1_root_add_513_2/n80 ), .ZN(\add_1_root_add_513_2/n208 ) );
XNOR2_X2 \add_1_root_add_513_2/U276  ( .A(\add_1_root_add_513_2/n59 ), .B(enc_byte_cnt[10]), .ZN(N2359) );
INV_X4 \add_1_root_add_513_2/U275  ( .A(enc_byte_cnt[11]), .ZN(\add_1_root_add_513_2/n207 ) );
XNOR2_X2 \add_1_root_add_513_2/U274  ( .A(\add_1_root_add_513_2/n28 ), .B(enc_byte_cnt[11]), .ZN(N2360) );
INV_X4 \add_1_root_add_513_2/U273  ( .A(enc_byte_cnt[12]), .ZN(\add_1_root_add_513_2/n204 ) );
XNOR2_X2 \add_1_root_add_513_2/U272  ( .A(\add_1_root_add_513_2/n3 ), .B(\add_1_root_add_513_2/n204 ), .ZN(N2361) );
INV_X4 \add_1_root_add_513_2/U271  ( .A(enc_byte_cnt[13]), .ZN(\add_1_root_add_513_2/n203 ) );
XNOR2_X2 \add_1_root_add_513_2/U270  ( .A(\add_1_root_add_513_2/n4 ), .B(\add_1_root_add_513_2/n203 ), .ZN(N2362) );
INV_X4 \add_1_root_add_513_2/U269  ( .A(enc_byte_cnt[14]), .ZN(\add_1_root_add_513_2/n202 ) );
XNOR2_X2 \add_1_root_add_513_2/U268  ( .A(\add_1_root_add_513_2/n7 ), .B(\add_1_root_add_513_2/n202 ), .ZN(N2363) );
INV_X4 \add_1_root_add_513_2/U267  ( .A(enc_byte_cnt[15]), .ZN(\add_1_root_add_513_2/n201 ) );
XNOR2_X2 \add_1_root_add_513_2/U266  ( .A(\add_1_root_add_513_2/n26 ), .B(\add_1_root_add_513_2/n201 ), .ZN(N2364) );
NAND2_X2 \add_1_root_add_513_2/U265  ( .A1(\add_1_root_add_513_2/n196 ),.A2(\add_1_root_add_513_2/n197 ), .ZN(\add_1_root_add_513_2/n195 ) );
XNOR2_X2 \add_1_root_add_513_2/U264  ( .A(\add_1_root_add_513_2/n152 ), .B(enc_byte_cnt[16]), .ZN(N2365) );
XNOR2_X2 \add_1_root_add_513_2/U263  ( .A(\add_1_root_add_513_2/n189 ), .B(\add_1_root_add_513_2/n2 ), .ZN(N2366) );
NAND2_X2 \add_1_root_add_513_2/U262  ( .A1(\add_1_root_add_513_2/n2 ), .A2(enc_byte_cnt[17]), .ZN(\add_1_root_add_513_2/n188 ) );
XNOR2_X2 \add_1_root_add_513_2/U261  ( .A(\add_1_root_add_513_2/n188 ), .B(enc_byte_cnt[18]), .ZN(N2367) );
INV_X4 \add_1_root_add_513_2/U260  ( .A(enc_byte_cnt[19]), .ZN(\add_1_root_add_513_2/n187 ) );
XNOR2_X2 \add_1_root_add_513_2/U259  ( .A(\add_1_root_add_513_2/n48 ), .B(enc_byte_cnt[19]), .ZN(N2368) );
NAND2_X2 \add_1_root_add_513_2/U258  ( .A1(dii_data_size[1]), .A2(enc_byte_cnt[1]), .ZN(\add_1_root_add_513_2/n164 ) );
INV_X4 \add_1_root_add_513_2/U257  ( .A(\add_1_root_add_513_2/n164 ), .ZN(\add_1_root_add_513_2/n184 ) );
XNOR2_X2 \add_1_root_add_513_2/U256  ( .A(\add_1_root_add_513_2/n166 ), .B(\add_1_root_add_513_2/n183 ), .ZN(N2350) );
INV_X4 \add_1_root_add_513_2/U255  ( .A(\add_1_root_add_513_2/n41 ), .ZN(\add_1_root_add_513_2/n178 ) );
XNOR2_X2 \add_1_root_add_513_2/U254  ( .A(\add_1_root_add_513_2/n179 ), .B(\add_1_root_add_513_2/n178 ), .ZN(N2369) );
NAND2_X2 \add_1_root_add_513_2/U253  ( .A1(\add_1_root_add_513_2/n178 ),.A2(enc_byte_cnt[20]), .ZN(\add_1_root_add_513_2/n177 ) );
XNOR2_X2 \add_1_root_add_513_2/U252  ( .A(\add_1_root_add_513_2/n177 ), .B(enc_byte_cnt[21]), .ZN(N2370) );
XNOR2_X2 \add_1_root_add_513_2/U251  ( .A(\add_1_root_add_513_2/n51 ), .B(enc_byte_cnt[22]), .ZN(N2371) );
XNOR2_X2 \add_1_root_add_513_2/U250  ( .A(\add_1_root_add_513_2/n23 ), .B(enc_byte_cnt[23]), .ZN(N2372) );
XNOR2_X2 \add_1_root_add_513_2/U249  ( .A(\add_1_root_add_513_2/n38 ), .B(enc_byte_cnt[24]), .ZN(N2373) );
XNOR2_X2 \add_1_root_add_513_2/U248  ( .A(\add_1_root_add_513_2/n49 ), .B(enc_byte_cnt[25]), .ZN(N2374) );
XNOR2_X2 \add_1_root_add_513_2/U247  ( .A(\add_1_root_add_513_2/n50 ), .B(enc_byte_cnt[26]), .ZN(N2375) );
INV_X4 \add_1_root_add_513_2/U246  ( .A(enc_byte_cnt[27]), .ZN(\add_1_root_add_513_2/n172 ) );
XNOR2_X2 \add_1_root_add_513_2/U245  ( .A(\add_1_root_add_513_2/n24 ), .B(enc_byte_cnt[27]), .ZN(N2376) );
INV_X4 \add_1_root_add_513_2/U244  ( .A(enc_byte_cnt[28]), .ZN(\add_1_root_add_513_2/n159 ) );
XNOR2_X2 \add_1_root_add_513_2/U243  ( .A(\add_1_root_add_513_2/n42 ), .B(enc_byte_cnt[28]), .ZN(N2377) );
INV_X4 \add_1_root_add_513_2/U242  ( .A(enc_byte_cnt[29]), .ZN(\add_1_root_add_513_2/n167 ) );
XNOR2_X2 \add_1_root_add_513_2/U241  ( .A(\add_1_root_add_513_2/n52 ), .B(enc_byte_cnt[29]), .ZN(N2378) );
NAND2_X2 \add_1_root_add_513_2/U240  ( .A1(\add_1_root_add_513_2/n60 ), .A2(\add_1_root_add_513_2/n142 ), .ZN(\add_1_root_add_513_2/n163 ) );
NAND2_X2 \add_1_root_add_513_2/U239  ( .A1(\add_1_root_add_513_2/n57 ), .A2(\add_1_root_add_513_2/n164 ), .ZN(\add_1_root_add_513_2/n143 ) );
INV_X4 \add_1_root_add_513_2/U238  ( .A(\add_1_root_add_513_2/n53 ), .ZN(\add_1_root_add_513_2/n161 ) );
INV_X4 \add_1_root_add_513_2/U237  ( .A(enc_byte_cnt[30]), .ZN(\add_1_root_add_513_2/n162 ) );
XNOR2_X2 \add_1_root_add_513_2/U236  ( .A(\add_1_root_add_513_2/n161 ), .B(\add_1_root_add_513_2/n162 ), .ZN(N2379) );
INV_X4 \add_1_root_add_513_2/U235  ( .A(enc_byte_cnt[31]), .ZN(\add_1_root_add_513_2/n160 ) );
XNOR2_X2 \add_1_root_add_513_2/U234  ( .A(\add_1_root_add_513_2/n13 ), .B(\add_1_root_add_513_2/n160 ), .ZN(N2380) );
INV_X4 \add_1_root_add_513_2/U233  ( .A(\add_1_root_add_513_2/n93 ), .ZN(\add_1_root_add_513_2/n148 ) );
INV_X4 \add_1_root_add_513_2/U232  ( .A(\add_1_root_add_513_2/n94 ), .ZN(\add_1_root_add_513_2/n147 ) );
NAND2_X2 \add_1_root_add_513_2/U231  ( .A1(\add_1_root_add_513_2/n148 ),.A2(\add_1_root_add_513_2/n147 ), .ZN(\add_1_root_add_513_2/n107 ) );
XNOR2_X2 \add_1_root_add_513_2/U230  ( .A(\add_1_root_add_513_2/n157 ), .B(enc_byte_cnt[32]), .ZN(N2381) );
XNOR2_X2 \add_1_root_add_513_2/U229  ( .A(\add_1_root_add_513_2/n18 ), .B(\add_1_root_add_513_2/n151 ), .ZN(N2382) );
XNOR2_X2 \add_1_root_add_513_2/U228  ( .A(\add_1_root_add_513_2/n6 ), .B(\add_1_root_add_513_2/n150 ), .ZN(N2383) );
INV_X4 \add_1_root_add_513_2/U227  ( .A(enc_byte_cnt[35]), .ZN(\add_1_root_add_513_2/n154 ) );
XNOR2_X2 \add_1_root_add_513_2/U226  ( .A(\add_1_root_add_513_2/n34 ), .B(\add_1_root_add_513_2/n154 ), .ZN(N2384) );
NAND2_X2 \add_1_root_add_513_2/U225  ( .A1(\add_1_root_add_513_2/n148 ),.A2(\add_1_root_add_513_2/n15 ), .ZN(\add_1_root_add_513_2/n145 ) );
INV_X4 \add_1_root_add_513_2/U224  ( .A(\add_1_root_add_513_2/n108 ), .ZN(\add_1_root_add_513_2/n78 ) );
NAND2_X2 \add_1_root_add_513_2/U223  ( .A1(\add_1_root_add_513_2/n78 ), .A2(\add_1_root_add_513_2/n147 ), .ZN(\add_1_root_add_513_2/n146 ) );
XNOR2_X2 \add_1_root_add_513_2/U222  ( .A(\add_1_root_add_513_2/n5 ), .B(enc_byte_cnt[36]), .ZN(N2385) );
XNOR2_X2 \add_1_root_add_513_2/U221  ( .A(\add_1_root_add_513_2/n14 ), .B(enc_byte_cnt[37]), .ZN(N2386) );
XNOR2_X2 \add_1_root_add_513_2/U220  ( .A(\add_1_root_add_513_2/n54 ), .B(enc_byte_cnt[38]), .ZN(N2387) );
INV_X4 \add_1_root_add_513_2/U219  ( .A(enc_byte_cnt[39]), .ZN(\add_1_root_add_513_2/n144 ) );
XNOR2_X2 \add_1_root_add_513_2/U218  ( .A(\add_1_root_add_513_2/n33 ), .B(enc_byte_cnt[39]), .ZN(N2388) );
NAND2_X2 \add_1_root_add_513_2/U217  ( .A1(\add_1_root_add_513_2/n143 ),.A2(\add_1_root_add_513_2/n60 ), .ZN(\add_1_root_add_513_2/n141 ) );
NAND2_X2 \add_1_root_add_513_2/U216  ( .A1(\add_1_root_add_513_2/n141 ),.A2(\add_1_root_add_513_2/n142 ), .ZN(\add_1_root_add_513_2/n137 ) );
NAND2_X2 \add_1_root_add_513_2/U215  ( .A1(\add_1_root_add_513_2/n139 ),.A2(\add_1_root_add_513_2/n140 ), .ZN(\add_1_root_add_513_2/n138 ) );
XNOR2_X2 \add_1_root_add_513_2/U214  ( .A(\add_1_root_add_513_2/n137 ), .B(\add_1_root_add_513_2/n138 ), .ZN(N2352) );
INV_X4 \add_1_root_add_513_2/U213  ( .A(\add_1_root_add_513_2/n111 ), .ZN(\add_1_root_add_513_2/n132 ) );
NAND2_X2 \add_1_root_add_513_2/U212  ( .A1(\add_1_root_add_513_2/n132 ),.A2(\add_1_root_add_513_2/n15 ), .ZN(\add_1_root_add_513_2/n131 ) );
XNOR2_X2 \add_1_root_add_513_2/U211  ( .A(\add_1_root_add_513_2/n20 ), .B(enc_byte_cnt[40]), .ZN(N2389) );
INV_X4 \add_1_root_add_513_2/U210  ( .A(\add_1_root_add_513_2/n131 ), .ZN(\add_1_root_add_513_2/n124 ) );
NAND2_X2 \add_1_root_add_513_2/U209  ( .A1(\add_1_root_add_513_2/n124 ),.A2(enc_byte_cnt[40]), .ZN(\add_1_root_add_513_2/n130 ) );
XNOR2_X2 \add_1_root_add_513_2/U208  ( .A(\add_1_root_add_513_2/n19 ), .B(enc_byte_cnt[41]), .ZN(N2390) );
INV_X4 \add_1_root_add_513_2/U207  ( .A(\add_1_root_add_513_2/n130 ), .ZN(\add_1_root_add_513_2/n129 ) );
XNOR2_X2 \add_1_root_add_513_2/U206  ( .A(\add_1_root_add_513_2/n128 ), .B(enc_byte_cnt[42]), .ZN(N2391) );
INV_X4 \add_1_root_add_513_2/U205  ( .A(enc_byte_cnt[43]), .ZN(\add_1_root_add_513_2/n126 ) );
XNOR2_X2 \add_1_root_add_513_2/U204  ( .A(\add_1_root_add_513_2/n22 ), .B(\add_1_root_add_513_2/n126 ), .ZN(N2392) );
NAND4_X2 \add_1_root_add_513_2/U203  ( .A1(enc_byte_cnt[43]), .A2(enc_byte_cnt[42]), .A3(enc_byte_cnt[40]), .A4(enc_byte_cnt[41]), .ZN(\add_1_root_add_513_2/n112 ) );
INV_X4 \add_1_root_add_513_2/U202  ( .A(\add_1_root_add_513_2/n112 ), .ZN(\add_1_root_add_513_2/n125 ) );
NAND2_X2 \add_1_root_add_513_2/U201  ( .A1(\add_1_root_add_513_2/n124 ),.A2(\add_1_root_add_513_2/n125 ), .ZN(\add_1_root_add_513_2/n122 ) );
INV_X4 \add_1_root_add_513_2/U200  ( .A(enc_byte_cnt[44]), .ZN(\add_1_root_add_513_2/n123 ) );
XNOR2_X2 \add_1_root_add_513_2/U199  ( .A(\add_1_root_add_513_2/n31 ), .B(enc_byte_cnt[44]), .ZN(N2393) );
INV_X4 \add_1_root_add_513_2/U198  ( .A(\add_1_root_add_513_2/n122 ), .ZN(\add_1_root_add_513_2/n121 ) );
NAND2_X2 \add_1_root_add_513_2/U197  ( .A1(\add_1_root_add_513_2/n121 ),.A2(enc_byte_cnt[44]), .ZN(\add_1_root_add_513_2/n119 ) );
INV_X4 \add_1_root_add_513_2/U196  ( .A(enc_byte_cnt[45]), .ZN(\add_1_root_add_513_2/n120 ) );
XNOR2_X2 \add_1_root_add_513_2/U195  ( .A(\add_1_root_add_513_2/n45 ), .B(enc_byte_cnt[45]), .ZN(N2394) );
INV_X4 \add_1_root_add_513_2/U194  ( .A(\add_1_root_add_513_2/n119 ), .ZN(\add_1_root_add_513_2/n118 ) );
INV_X4 \add_1_root_add_513_2/U193  ( .A(enc_byte_cnt[46]), .ZN(\add_1_root_add_513_2/n117 ) );
XNOR2_X2 \add_1_root_add_513_2/U192  ( .A(\add_1_root_add_513_2/n116 ), .B(\add_1_root_add_513_2/n117 ), .ZN(N2395) );
INV_X4 \add_1_root_add_513_2/U191  ( .A(enc_byte_cnt[47]), .ZN(\add_1_root_add_513_2/n115 ) );
XNOR2_X2 \add_1_root_add_513_2/U190  ( .A(\add_1_root_add_513_2/n21 ), .B(\add_1_root_add_513_2/n115 ), .ZN(N2396) );
NAND2_X2 \add_1_root_add_513_2/U189  ( .A1(enc_byte_cnt[47]), .A2(enc_byte_cnt[46]), .ZN(\add_1_root_add_513_2/n113 ) );
XNOR2_X2 \add_1_root_add_513_2/U188  ( .A(\add_1_root_add_513_2/n37 ), .B(enc_byte_cnt[48]), .ZN(N2397) );
INV_X4 \add_1_root_add_513_2/U187  ( .A(\add_1_root_add_513_2/n105 ), .ZN(\add_1_root_add_513_2/n92 ) );
INV_X4 \add_1_root_add_513_2/U186  ( .A(\add_1_root_add_513_2/n55 ), .ZN(\add_1_root_add_513_2/n104 ) );
XNOR2_X2 \add_1_root_add_513_2/U185  ( .A(\add_1_root_add_513_2/n104 ), .B(\add_1_root_add_513_2/n101 ), .ZN(N2398) );
XNOR2_X2 \add_1_root_add_513_2/U184  ( .A(\add_1_root_add_513_2/n103 ), .B(\add_1_root_add_513_2/n80 ), .ZN(N2353) );
INV_X4 \add_1_root_add_513_2/U183  ( .A(enc_byte_cnt[49]), .ZN(\add_1_root_add_513_2/n101 ) );
INV_X4 \add_1_root_add_513_2/U182  ( .A(enc_byte_cnt[50]), .ZN(\add_1_root_add_513_2/n102 ) );
XNOR2_X2 \add_1_root_add_513_2/U181  ( .A(\add_1_root_add_513_2/n32 ), .B(\add_1_root_add_513_2/n102 ), .ZN(N2399) );
INV_X4 \add_1_root_add_513_2/U180  ( .A(\add_1_root_add_513_2/n99 ), .ZN(\add_1_root_add_513_2/n100 ) );
XNOR2_X2 \add_1_root_add_513_2/U179  ( .A(\add_1_root_add_513_2/n46 ), .B(enc_byte_cnt[51]), .ZN(N2400) );
NAND2_X2 \add_1_root_add_513_2/U178  ( .A1(\add_1_root_add_513_2/n99 ), .A2(enc_byte_cnt[51]), .ZN(\add_1_root_add_513_2/n98 ) );
XNOR2_X2 \add_1_root_add_513_2/U177  ( .A(\add_1_root_add_513_2/n43 ), .B(enc_byte_cnt[52]), .ZN(N2401) );
INV_X4 \add_1_root_add_513_2/U176  ( .A(\add_1_root_add_513_2/n98 ), .ZN(\add_1_root_add_513_2/n97 ) );
NAND2_X2 \add_1_root_add_513_2/U175  ( .A1(\add_1_root_add_513_2/n97 ), .A2(enc_byte_cnt[52]), .ZN(\add_1_root_add_513_2/n96 ) );
XNOR2_X2 \add_1_root_add_513_2/U174  ( .A(\add_1_root_add_513_2/n8 ), .B(enc_byte_cnt[53]), .ZN(N2402) );
INV_X4 \add_1_root_add_513_2/U173  ( .A(\add_1_root_add_513_2/n96 ), .ZN(\add_1_root_add_513_2/n77 ) );
NAND2_X2 \add_1_root_add_513_2/U172  ( .A1(\add_1_root_add_513_2/n77 ), .A2(\add_1_root_add_513_2/n78 ), .ZN(\add_1_root_add_513_2/n90 ) );
NAND2_X2 \add_1_root_add_513_2/U171  ( .A1(enc_byte_cnt[48]), .A2(enc_byte_cnt[53]), .ZN(\add_1_root_add_513_2/n95 ) );
NAND2_X2 \add_1_root_add_513_2/U170  ( .A1(\add_1_root_add_513_2/n91 ), .A2(\add_1_root_add_513_2/n92 ), .ZN(\add_1_root_add_513_2/n76 ) );
INV_X4 \add_1_root_add_513_2/U169  ( .A(enc_byte_cnt[54]), .ZN(\add_1_root_add_513_2/n89 ) );
XNOR2_X2 \add_1_root_add_513_2/U168  ( .A(\add_1_root_add_513_2/n1 ), .B(enc_byte_cnt[54]), .ZN(N2403) );
INV_X4 \add_1_root_add_513_2/U167  ( .A(enc_byte_cnt[55]), .ZN(\add_1_root_add_513_2/n88 ) );
XNOR2_X2 \add_1_root_add_513_2/U166  ( .A(\add_1_root_add_513_2/n30 ), .B(enc_byte_cnt[55]), .ZN(N2404) );
INV_X4 \add_1_root_add_513_2/U165  ( .A(\add_1_root_add_513_2/n86 ), .ZN(\add_1_root_add_513_2/n87 ) );
XNOR2_X2 \add_1_root_add_513_2/U164  ( .A(\add_1_root_add_513_2/n12 ), .B(enc_byte_cnt[56]), .ZN(N2405) );
NAND2_X2 \add_1_root_add_513_2/U163  ( .A1(\add_1_root_add_513_2/n86 ), .A2(enc_byte_cnt[56]), .ZN(\add_1_root_add_513_2/n85 ) );
XNOR2_X2 \add_1_root_add_513_2/U162  ( .A(\add_1_root_add_513_2/n11 ), .B(enc_byte_cnt[57]), .ZN(N2406) );
INV_X4 \add_1_root_add_513_2/U161  ( .A(\add_1_root_add_513_2/n85 ), .ZN(\add_1_root_add_513_2/n84 ) );
NAND2_X2 \add_1_root_add_513_2/U160  ( .A1(\add_1_root_add_513_2/n84 ), .A2(enc_byte_cnt[57]), .ZN(\add_1_root_add_513_2/n83 ) );
XNOR2_X2 \add_1_root_add_513_2/U159  ( .A(\add_1_root_add_513_2/n10 ), .B(enc_byte_cnt[58]), .ZN(N2407) );
INV_X4 \add_1_root_add_513_2/U158  ( .A(\add_1_root_add_513_2/n83 ), .ZN(\add_1_root_add_513_2/n82 ) );
NAND2_X2 \add_1_root_add_513_2/U157  ( .A1(\add_1_root_add_513_2/n82 ), .A2(enc_byte_cnt[58]), .ZN(\add_1_root_add_513_2/n74 ) );
XNOR2_X2 \add_1_root_add_513_2/U156  ( .A(\add_1_root_add_513_2/n9 ), .B(enc_byte_cnt[59]), .ZN(N2408) );
XNOR2_X2 \add_1_root_add_513_2/U155  ( .A(\add_1_root_add_513_2/n81 ), .B(\add_1_root_add_513_2/n16 ), .ZN(N2354) );
INV_X4 \add_1_root_add_513_2/U154  ( .A(enc_byte_cnt[60]), .ZN(\add_1_root_add_513_2/n79 ) );
NAND2_X2 \add_1_root_add_513_2/U153  ( .A1(\add_1_root_add_513_2/n77 ), .A2(\add_1_root_add_513_2/n78 ), .ZN(\add_1_root_add_513_2/n75 ) );
INV_X4 \add_1_root_add_513_2/U152  ( .A(\add_1_root_add_513_2/n74 ), .ZN(\add_1_root_add_513_2/n73 ) );
NAND2_X2 \add_1_root_add_513_2/U151  ( .A1(\add_1_root_add_513_2/n73 ), .A2(enc_byte_cnt[59]), .ZN(\add_1_root_add_513_2/n70 ) );
XNOR2_X2 \add_1_root_add_513_2/U150  ( .A(\add_1_root_add_513_2/n79 ), .B(\add_1_root_add_513_2/n17 ), .ZN(N2409) );
INV_X4 \add_1_root_add_513_2/U149  ( .A(enc_byte_cnt[61]), .ZN(\add_1_root_add_513_2/n72 ) );
XNOR2_X2 \add_1_root_add_513_2/U148  ( .A(\add_1_root_add_513_2/n27 ), .B(\add_1_root_add_513_2/n72 ), .ZN(N2410) );
INV_X4 \add_1_root_add_513_2/U147  ( .A(enc_byte_cnt[62]), .ZN(\add_1_root_add_513_2/n71 ) );
XNOR2_X2 \add_1_root_add_513_2/U146  ( .A(\add_1_root_add_513_2/n25 ), .B(\add_1_root_add_513_2/n71 ), .ZN(N2411) );
NAND2_X2 \add_1_root_add_513_2/U145  ( .A1(\add_1_root_add_513_2/n69 ), .A2(enc_byte_cnt[62]), .ZN(\add_1_root_add_513_2/n68 ) );
NAND2_X2 \add_1_root_add_513_2/U144  ( .A1(\add_1_root_add_513_2/n16 ), .A2(enc_byte_cnt[5]), .ZN(\add_1_root_add_513_2/n66 ) );
XNOR2_X2 \add_1_root_add_513_2/U143  ( .A(\add_1_root_add_513_2/n66 ), .B(enc_byte_cnt[6]), .ZN(N2355) );
XNOR2_X2 \add_1_root_add_513_2/U142  ( .A(\add_1_root_add_513_2/n29 ), .B(enc_byte_cnt[7]), .ZN(N2356) );
XNOR2_X2 \add_1_root_add_513_2/U141  ( .A(\add_1_root_add_513_2/n63 ), .B(\add_1_root_add_513_2/n64 ), .ZN(N2357) );
XNOR2_X2 \add_1_root_add_513_2/U140  ( .A(\add_1_root_add_513_2/n58 ), .B(enc_byte_cnt[9]), .ZN(N2358) );
INV_X4 \add_1_root_add_513_2/U139  ( .A(enc_byte_cnt[38]), .ZN(\add_1_root_add_513_2/n134 ) );
INV_X4 \add_1_root_add_513_2/U138  ( .A(enc_byte_cnt[37]), .ZN(\add_1_root_add_513_2/n136 ) );
INV_X4 \add_1_root_add_513_2/U137  ( .A(enc_byte_cnt[36]), .ZN(\add_1_root_add_513_2/n135 ) );
INV_X4 \add_1_root_add_513_2/U136  ( .A(enc_byte_cnt[34]), .ZN(\add_1_root_add_513_2/n150 ) );
INV_X4 \add_1_root_add_513_2/U135  ( .A(enc_byte_cnt[33]), .ZN(\add_1_root_add_513_2/n151 ) );
INV_X4 \add_1_root_add_513_2/U134  ( .A(enc_byte_cnt[32]), .ZN(\add_1_root_add_513_2/n156 ) );
INV_X4 \add_1_root_add_513_2/U133  ( .A(enc_byte_cnt[26]), .ZN(\add_1_root_add_513_2/n169 ) );
INV_X4 \add_1_root_add_513_2/U132  ( .A(enc_byte_cnt[25]), .ZN(\add_1_root_add_513_2/n171 ) );
INV_X4 \add_1_root_add_513_2/U131  ( .A(enc_byte_cnt[24]), .ZN(\add_1_root_add_513_2/n170 ) );
INV_X4 \add_1_root_add_513_2/U130  ( .A(enc_byte_cnt[23]), .ZN(\add_1_root_add_513_2/n175 ) );
INV_X4 \add_1_root_add_513_2/U129  ( .A(enc_byte_cnt[22]), .ZN(\add_1_root_add_513_2/n174 ) );
INV_X4 \add_1_root_add_513_2/U128  ( .A(enc_byte_cnt[21]), .ZN(\add_1_root_add_513_2/n176 ) );
INV_X4 \add_1_root_add_513_2/U127  ( .A(enc_byte_cnt[20]), .ZN(\add_1_root_add_513_2/n179 ) );
INV_X4 \add_1_root_add_513_2/U126  ( .A(enc_byte_cnt[18]), .ZN(\add_1_root_add_513_2/n181 ) );
INV_X4 \add_1_root_add_513_2/U125  ( .A(enc_byte_cnt[17]), .ZN(\add_1_root_add_513_2/n189 ) );
INV_X4 \add_1_root_add_513_2/U124  ( .A(enc_byte_cnt[16]), .ZN(\add_1_root_add_513_2/n182 ) );
INV_X4 \add_1_root_add_513_2/U123  ( .A(enc_byte_cnt[10]), .ZN(\add_1_root_add_513_2/n206 ) );
INV_X4 \add_1_root_add_513_2/U122  ( .A(enc_byte_cnt[9]), .ZN(\add_1_root_add_513_2/n62 ) );
INV_X4 \add_1_root_add_513_2/U121  ( .A(enc_byte_cnt[8]), .ZN(\add_1_root_add_513_2/n64 ) );
INV_X4 \add_1_root_add_513_2/U120  ( .A(enc_byte_cnt[6]), .ZN(\add_1_root_add_513_2/n65 ) );
INV_X4 \add_1_root_add_513_2/U119  ( .A(enc_byte_cnt[4]), .ZN(\add_1_root_add_513_2/n103 ) );
INV_X4 \add_1_root_add_513_2/U118  ( .A(enc_byte_cnt[5]), .ZN(\add_1_root_add_513_2/n81 ) );
INV_X4 \add_1_root_add_513_2/U117  ( .A(\add_1_root_add_513_2/n186 ), .ZN(\add_1_root_add_513_2/n210 ) );
INV_X4 \add_1_root_add_513_2/U116  ( .A(\add_1_root_add_513_2/n114 ), .ZN(\add_1_root_add_513_2/n157 ) );
INV_X4 \add_1_root_add_513_2/U115  ( .A(\add_1_root_add_513_2/n127 ), .ZN(\add_1_root_add_513_2/n128 ) );
INV_X4 \add_1_root_add_513_2/U114  ( .A(\add_1_root_add_513_2/n208 ), .ZN(\add_1_root_add_513_2/n63 ) );
NOR2_X2 \add_1_root_add_513_2/U113  ( .A1(\add_1_root_add_513_2/n184 ), .A2(\add_1_root_add_513_2/n165 ), .ZN(\add_1_root_add_513_2/n183 ) );
OR2_X2 \add_1_root_add_513_2/U112  ( .A1(enc_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(\add_1_root_add_513_2/n60 ) );
NOR2_X2 \add_1_root_add_513_2/U111  ( .A1(\add_1_root_add_513_2/n44 ), .A2(\add_1_root_add_513_2/n68 ), .ZN(\add_1_root_add_513_2/n67 ) );
XOR2_X2 \add_1_root_add_513_2/U110  ( .A(\add_1_root_add_513_2/n67 ), .B(enc_byte_cnt[63]), .Z(N2412) );
AND2_X2 \add_1_root_add_513_2/U109  ( .A1(enc_byte_cnt[0]), .A2(n17750),.ZN(\add_1_root_add_513_2/n219 ) );
NOR2_X2 \add_1_root_add_513_2/U108  ( .A1(\add_1_root_add_513_2/n217 ), .A2(\add_1_root_add_513_2/n218 ), .ZN(\add_1_root_add_513_2/n216 ) );
NAND3_X2 \add_1_root_add_513_2/U107  ( .A1(dii_data_size[1]), .A2(\add_1_root_add_513_2/n60 ), .A3(enc_byte_cnt[1]), .ZN(\add_1_root_add_513_2/n215 ) );
NAND3_X2 \add_1_root_add_513_2/U106  ( .A1(\add_1_root_add_513_2/n214 ),.A2(\add_1_root_add_513_2/n215 ), .A3(\add_1_root_add_513_2/n216 ),.ZN(\add_1_root_add_513_2/n193 ) );
NOR2_X2 \add_1_root_add_513_2/U105  ( .A1(enc_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(\add_1_root_add_513_2/n222 ) );
NOR2_X2 \add_1_root_add_513_2/U104  ( .A1(enc_byte_cnt[2]), .A2(dii_data_size[2]), .ZN(\add_1_root_add_513_2/n221 ) );
NOR2_X2 \add_1_root_add_513_2/U103  ( .A1(\add_1_root_add_513_2/n221 ), .A2(\add_1_root_add_513_2/n222 ), .ZN(\add_1_root_add_513_2/n220 ) );
NOR2_X2 \add_1_root_add_513_2/U102  ( .A1(enc_byte_cnt[0]), .A2(n17750),.ZN(\add_1_root_add_513_2/n186 ) );
NOR2_X2 \add_1_root_add_513_2/U101  ( .A1(enc_byte_cnt[1]), .A2(dii_data_size[1]), .ZN(\add_1_root_add_513_2/n165 ) );
INV_X4 \add_1_root_add_513_2/U100  ( .A(n18074), .ZN(\add_1_root_add_513_2/n61 ) );
AND2_X2 \add_1_root_add_513_2/U99  ( .A1(\add_1_root_add_513_2/n186 ), .A2(\add_1_root_add_513_2/n185 ), .ZN(\add_1_root_add_513_2/n166 ) );
NOR2_X2 \add_1_root_add_513_2/U98  ( .A1(\add_1_root_add_513_2/n154 ), .A2(\add_1_root_add_513_2/n150 ), .ZN(\add_1_root_add_513_2/n149 ) );
OR2_X2 \add_1_root_add_513_2/U97  ( .A1(\add_1_root_add_513_2/n58 ), .A2(\add_1_root_add_513_2/n62 ), .ZN(\add_1_root_add_513_2/n59 ) );
NOR2_X2 \add_1_root_add_513_2/U96  ( .A1(\add_1_root_add_513_2/n134 ), .A2(\add_1_root_add_513_2/n144 ), .ZN(\add_1_root_add_513_2/n133 ) );
NAND3_X2 \add_1_root_add_513_2/U95  ( .A1(enc_byte_cnt[37]), .A2(enc_byte_cnt[36]), .A3(\add_1_root_add_513_2/n133 ), .ZN(\add_1_root_add_513_2/n111 ) );
OR2_X2 \add_1_root_add_513_2/U94  ( .A1(\add_1_root_add_513_2/n208 ), .A2(\add_1_root_add_513_2/n64 ), .ZN(\add_1_root_add_513_2/n58 ) );
NOR2_X2 \add_1_root_add_513_2/U93  ( .A1(\add_1_root_add_513_2/n167 ), .A2(\add_1_root_add_513_2/n159 ), .ZN(\add_1_root_add_513_2/n158 ) );
NAND3_X2 \add_1_root_add_513_2/U92  ( .A1(enc_byte_cnt[30]), .A2(enc_byte_cnt[31]), .A3(\add_1_root_add_513_2/n158 ), .ZN(\add_1_root_add_513_2/n93 ) );
NOR2_X2 \add_1_root_add_513_2/U91  ( .A1(\add_1_root_add_513_2/n151 ), .A2(\add_1_root_add_513_2/n156 ), .ZN(\add_1_root_add_513_2/n155 ) );
AND2_X2 \add_1_root_add_513_2/U90  ( .A1(enc_byte_cnt[61]), .A2(enc_byte_cnt[60]), .ZN(\add_1_root_add_513_2/n69 ) );
NOR2_X2 \add_1_root_add_513_2/U89  ( .A1(\add_1_root_add_513_2/n169 ), .A2(\add_1_root_add_513_2/n172 ), .ZN(\add_1_root_add_513_2/n168 ) );
NAND3_X2 \add_1_root_add_513_2/U88  ( .A1(enc_byte_cnt[25]), .A2(enc_byte_cnt[24]), .A3(\add_1_root_add_513_2/n168 ), .ZN(\add_1_root_add_513_2/n94 ) );
NOR2_X2 \add_1_root_add_513_2/U87  ( .A1(\add_1_root_add_513_2/n102 ), .A2(\add_1_root_add_513_2/n101 ), .ZN(\add_1_root_add_513_2/n99 ) );
NOR2_X2 \add_1_root_add_513_2/U86  ( .A1(\add_1_root_add_513_2/n88 ), .A2(\add_1_root_add_513_2/n89 ), .ZN(\add_1_root_add_513_2/n86 ) );
NOR2_X2 \add_1_root_add_513_2/U85  ( .A1(\add_1_root_add_513_2/n187 ), .A2(\add_1_root_add_513_2/n181 ), .ZN(\add_1_root_add_513_2/n180 ) );
NAND3_X2 \add_1_root_add_513_2/U84  ( .A1(enc_byte_cnt[16]), .A2(enc_byte_cnt[17]), .A3(\add_1_root_add_513_2/n180 ), .ZN(\add_1_root_add_513_2/n153 ) );
NOR2_X2 \add_1_root_add_513_2/U83  ( .A1(\add_1_root_add_513_2/n174 ), .A2(\add_1_root_add_513_2/n175 ), .ZN(\add_1_root_add_513_2/n173 ) );
NAND3_X2 \add_1_root_add_513_2/U82  ( .A1(enc_byte_cnt[21]), .A2(enc_byte_cnt[20]), .A3(\add_1_root_add_513_2/n173 ), .ZN(\add_1_root_add_513_2/n108 ) );
OR2_X2 \add_1_root_add_513_2/U81  ( .A1(\add_1_root_add_513_2/n165 ), .A2(\add_1_root_add_513_2/n166 ), .ZN(\add_1_root_add_513_2/n57 ) );
NOR3_X2 \add_1_root_add_513_2/U80  ( .A1(\add_1_root_add_513_2/n93 ), .A2(\add_1_root_add_513_2/n94 ), .A3(\add_1_root_add_513_2/n95 ), .ZN(\add_1_root_add_513_2/n91 ) );
AND2_X4 \add_1_root_add_513_2/U79  ( .A1(\add_1_root_add_513_2/n92 ), .A2(enc_byte_cnt[48]), .ZN(\add_1_root_add_513_2/n56 ) );
NAND2_X2 \add_1_root_add_513_2/U78  ( .A1(\add_1_root_add_513_2/n106 ), .A2(\add_1_root_add_513_2/n56 ), .ZN(\add_1_root_add_513_2/n55 ) );
NOR2_X2 \add_1_root_add_513_2/U77  ( .A1(\add_1_root_add_513_2/n212 ), .A2(\add_1_root_add_513_2/n165 ), .ZN(\add_1_root_add_513_2/n211 ) );
NAND3_X2 \add_1_root_add_513_2/U76  ( .A1(\add_1_root_add_513_2/n210 ), .A2(\add_1_root_add_513_2/n60 ), .A3(\add_1_root_add_513_2/n211 ), .ZN(\add_1_root_add_513_2/n200 ) );
OR3_X2 \add_1_root_add_513_2/U75  ( .A1(\add_1_root_add_513_2/n5 ), .A2(\add_1_root_add_513_2/n135 ), .A3(\add_1_root_add_513_2/n136 ), .ZN(\add_1_root_add_513_2/n54 ) );
OR3_X2 \add_1_root_add_513_2/U74  ( .A1(\add_1_root_add_513_2/n42 ), .A2(\add_1_root_add_513_2/n167 ), .A3(\add_1_root_add_513_2/n159 ), .ZN(\add_1_root_add_513_2/n53 ) );
NOR2_X2 \add_1_root_add_513_2/U73  ( .A1(\add_1_root_add_513_2/n65 ), .A2(\add_1_root_add_513_2/n224 ), .ZN(\add_1_root_add_513_2/n223 ) );
NAND3_X2 \add_1_root_add_513_2/U72  ( .A1(enc_byte_cnt[5]), .A2(enc_byte_cnt[4]), .A3(\add_1_root_add_513_2/n223 ), .ZN(\add_1_root_add_513_2/n198 ) );
OR2_X2 \add_1_root_add_513_2/U71  ( .A1(\add_1_root_add_513_2/n159 ), .A2(\add_1_root_add_513_2/n42 ), .ZN(\add_1_root_add_513_2/n52 ) );
OR2_X2 \add_1_root_add_513_2/U70  ( .A1(\add_1_root_add_513_2/n176 ), .A2(\add_1_root_add_513_2/n177 ), .ZN(\add_1_root_add_513_2/n51 ) );
OR2_X2 \add_1_root_add_513_2/U69  ( .A1(\add_1_root_add_513_2/n171 ), .A2(\add_1_root_add_513_2/n49 ), .ZN(\add_1_root_add_513_2/n50 ) );
OR2_X2 \add_1_root_add_513_2/U68  ( .A1(\add_1_root_add_513_2/n170 ), .A2(\add_1_root_add_513_2/n38 ), .ZN(\add_1_root_add_513_2/n49 ) );
OR2_X2 \add_1_root_add_513_2/U67  ( .A1(\add_1_root_add_513_2/n181 ), .A2(\add_1_root_add_513_2/n188 ), .ZN(\add_1_root_add_513_2/n48 ) );
AND2_X2 \add_1_root_add_513_2/U66  ( .A1(enc_byte_cnt[13]), .A2(enc_byte_cnt[12]), .ZN(\add_1_root_add_513_2/n199 ) );
AND2_X4 \add_1_root_add_513_2/U65  ( .A1(\add_1_root_add_513_2/n118 ), .A2(enc_byte_cnt[45]), .ZN(\add_1_root_add_513_2/n47 ) );
AND2_X2 \add_1_root_add_513_2/U64  ( .A1(\add_1_root_add_513_2/n114 ), .A2(\add_1_root_add_513_2/n47 ), .ZN(\add_1_root_add_513_2/n116 ) );
NOR2_X2 \add_1_root_add_513_2/U63  ( .A1(\add_1_root_add_513_2/n206 ), .A2(\add_1_root_add_513_2/n207 ), .ZN(\add_1_root_add_513_2/n205 ) );
NAND3_X2 \add_1_root_add_513_2/U62  ( .A1(enc_byte_cnt[9]), .A2(enc_byte_cnt[8]), .A3(\add_1_root_add_513_2/n205 ), .ZN(\add_1_root_add_513_2/n192 ) );
NAND3_X2 \add_1_root_add_513_2/U61  ( .A1(\add_1_root_add_513_2/n140 ), .A2(\add_1_root_add_513_2/n193 ), .A3(\add_1_root_add_513_2/n194 ), .ZN(\add_1_root_add_513_2/n190 ) );
NOR2_X2 \add_1_root_add_513_2/U60  ( .A1(\add_1_root_add_513_2/n111 ), .A2(\add_1_root_add_513_2/n112 ), .ZN(\add_1_root_add_513_2/n110 ) );
NOR3_X2 \add_1_root_add_513_2/U59  ( .A1(\add_1_root_add_513_2/n113 ), .A2(\add_1_root_add_513_2/n120 ), .A3(\add_1_root_add_513_2/n123 ), .ZN(\add_1_root_add_513_2/n109 ) );
NAND3_X2 \add_1_root_add_513_2/U58  ( .A1(\add_1_root_add_513_2/n109 ), .A2(\add_1_root_add_513_2/n15 ), .A3(\add_1_root_add_513_2/n110 ), .ZN(\add_1_root_add_513_2/n105 ) );
OR2_X2 \add_1_root_add_513_2/U57  ( .A1(\add_1_root_add_513_2/n55 ), .A2(\add_1_root_add_513_2/n100 ), .ZN(\add_1_root_add_513_2/n46 ) );
OR2_X2 \add_1_root_add_513_2/U56  ( .A1(\add_1_root_add_513_2/n157 ), .A2(\add_1_root_add_513_2/n119 ), .ZN(\add_1_root_add_513_2/n45 ) );
AND2_X2 \add_1_root_add_513_2/U55  ( .A1(\add_1_root_add_513_2/n195 ), .A2(\add_1_root_add_513_2/n36 ), .ZN(\add_1_root_add_513_2/n152 ) );
OR2_X2 \add_1_root_add_513_2/U54  ( .A1(\add_1_root_add_513_2/n1 ), .A2(\add_1_root_add_513_2/n70 ), .ZN(\add_1_root_add_513_2/n44 ) );
NOR2_X2 \add_1_root_add_513_2/U53  ( .A1(\add_1_root_add_513_2/n198 ), .A2(\add_1_root_add_513_2/n191 ), .ZN(\add_1_root_add_513_2/n197 ) );
NOR2_X2 \add_1_root_add_513_2/U52  ( .A1(\add_1_root_add_513_2/n192 ), .A2(\add_1_root_add_513_2/n200 ), .ZN(\add_1_root_add_513_2/n196 ) );
OR2_X2 \add_1_root_add_513_2/U51  ( .A1(\add_1_root_add_513_2/n55 ), .A2(\add_1_root_add_513_2/n98 ), .ZN(\add_1_root_add_513_2/n43 ) );
OR2_X2 \add_1_root_add_513_2/U50  ( .A1(\add_1_root_add_513_2/n38 ), .A2(\add_1_root_add_513_2/n94 ), .ZN(\add_1_root_add_513_2/n42 ) );
OR2_X2 \add_1_root_add_513_2/U49  ( .A1(\add_1_root_add_513_2/n152 ), .A2(\add_1_root_add_513_2/n153 ), .ZN(\add_1_root_add_513_2/n41 ) );
OR2_X2 \add_1_root_add_513_2/U48  ( .A1(\add_1_root_add_513_2/n152 ), .A2(\add_1_root_add_513_2/n153 ), .ZN(\add_1_root_add_513_2/n40 ) );
AND2_X4 \add_1_root_add_513_2/U47  ( .A1(\add_1_root_add_513_2/n129 ), .A2(enc_byte_cnt[41]), .ZN(\add_1_root_add_513_2/n39 ) );
AND2_X2 \add_1_root_add_513_2/U46  ( .A1(\add_1_root_add_513_2/n114 ), .A2(\add_1_root_add_513_2/n39 ), .ZN(\add_1_root_add_513_2/n127 ) );
OR3_X2 \add_1_root_add_513_2/U45  ( .A1(\add_1_root_add_513_2/n152 ), .A2(\add_1_root_add_513_2/n153 ), .A3(\add_1_root_add_513_2/n108 ), .ZN(\add_1_root_add_513_2/n38 ) );
NOR3_X2 \add_1_root_add_513_2/U44  ( .A1(\add_1_root_add_513_2/n40 ), .A2(\add_1_root_add_513_2/n107 ), .A3(\add_1_root_add_513_2/n108 ), .ZN(\add_1_root_add_513_2/n106 ) );
NOR3_X2 \add_1_root_add_513_2/U43  ( .A1(\add_1_root_add_513_2/n107 ), .A2(\add_1_root_add_513_2/n41 ), .A3(\add_1_root_add_513_2/n108 ), .ZN(\add_1_root_add_513_2/n114 ) );
OR2_X2 \add_1_root_add_513_2/U42  ( .A1(\add_1_root_add_513_2/n157 ), .A2(\add_1_root_add_513_2/n105 ), .ZN(\add_1_root_add_513_2/n37 ) );
XNOR2_X1 \add_1_root_add_513_2/U41  ( .A(\add_1_root_add_513_2/n163 ), .B(\add_1_root_add_513_2/n143 ), .ZN(N2351) );
NAND2_X1 \add_1_root_add_513_2/U40  ( .A1(n17750), .A2(enc_byte_cnt[0]),.ZN(\add_1_root_add_513_2/n185 ) );
NAND2_X1 \add_1_root_add_513_2/U39  ( .A1(\add_1_root_add_513_2/n185 ), .A2(\add_1_root_add_513_2/n210 ), .ZN(N2349) );
OR3_X4 \add_1_root_add_513_2/U38  ( .A1(\add_1_root_add_513_2/n190 ), .A2(\add_1_root_add_513_2/n191 ), .A3(\add_1_root_add_513_2/n192 ), .ZN(\add_1_root_add_513_2/n36 ) );
OR3_X4 \add_1_root_add_513_2/U37  ( .A1(\add_1_root_add_513_2/n40 ), .A2(\add_1_root_add_513_2/n75 ), .A3(\add_1_root_add_513_2/n76 ), .ZN(\add_1_root_add_513_2/n35 ) );
AND2_X4 \add_1_root_add_513_2/U36  ( .A1(\add_1_root_add_513_2/n6 ), .A2(enc_byte_cnt[34]), .ZN(\add_1_root_add_513_2/n34 ) );
OR2_X4 \add_1_root_add_513_2/U35  ( .A1(\add_1_root_add_513_2/n134 ), .A2(\add_1_root_add_513_2/n54 ), .ZN(\add_1_root_add_513_2/n33 ) );
NOR2_X2 \add_1_root_add_513_2/U34  ( .A1(\add_1_root_add_513_2/n101 ), .A2(\add_1_root_add_513_2/n55 ), .ZN(\add_1_root_add_513_2/n32 ) );
OR2_X4 \add_1_root_add_513_2/U33  ( .A1(\add_1_root_add_513_2/n157 ), .A2(\add_1_root_add_513_2/n122 ), .ZN(\add_1_root_add_513_2/n31 ) );
OR2_X4 \add_1_root_add_513_2/U32  ( .A1(\add_1_root_add_513_2/n89 ), .A2(\add_1_root_add_513_2/n1 ), .ZN(\add_1_root_add_513_2/n30 ) );
OR2_X4 \add_1_root_add_513_2/U31  ( .A1(\add_1_root_add_513_2/n65 ), .A2(\add_1_root_add_513_2/n66 ), .ZN(\add_1_root_add_513_2/n29 ) );
OR2_X4 \add_1_root_add_513_2/U30  ( .A1(\add_1_root_add_513_2/n206 ), .A2(\add_1_root_add_513_2/n59 ), .ZN(\add_1_root_add_513_2/n28 ) );
AND2_X4 \add_1_root_add_513_2/U29  ( .A1(enc_byte_cnt[60]), .A2(\add_1_root_add_513_2/n17 ), .ZN(\add_1_root_add_513_2/n27 ) );
AND2_X4 \add_1_root_add_513_2/U28  ( .A1(enc_byte_cnt[14]), .A2(\add_1_root_add_513_2/n7 ), .ZN(\add_1_root_add_513_2/n26 ) );
AND2_X4 \add_1_root_add_513_2/U27  ( .A1(\add_1_root_add_513_2/n69 ), .A2(\add_1_root_add_513_2/n17 ), .ZN(\add_1_root_add_513_2/n25 ) );
OR2_X4 \add_1_root_add_513_2/U26  ( .A1(\add_1_root_add_513_2/n169 ), .A2(\add_1_root_add_513_2/n50 ), .ZN(\add_1_root_add_513_2/n24 ) );
OR2_X4 \add_1_root_add_513_2/U25  ( .A1(\add_1_root_add_513_2/n174 ), .A2(\add_1_root_add_513_2/n51 ), .ZN(\add_1_root_add_513_2/n23 ) );
AND2_X4 \add_1_root_add_513_2/U24  ( .A1(\add_1_root_add_513_2/n127 ), .A2(enc_byte_cnt[42]), .ZN(\add_1_root_add_513_2/n22 ) );
AND2_X4 \add_1_root_add_513_2/U23  ( .A1(\add_1_root_add_513_2/n116 ), .A2(enc_byte_cnt[46]), .ZN(\add_1_root_add_513_2/n21 ) );
OR2_X4 \add_1_root_add_513_2/U22  ( .A1(\add_1_root_add_513_2/n157 ), .A2(\add_1_root_add_513_2/n131 ), .ZN(\add_1_root_add_513_2/n20 ) );
OR2_X4 \add_1_root_add_513_2/U21  ( .A1(\add_1_root_add_513_2/n157 ), .A2(\add_1_root_add_513_2/n130 ), .ZN(\add_1_root_add_513_2/n19 ) );
AND2_X4 \add_1_root_add_513_2/U20  ( .A1(\add_1_root_add_513_2/n114 ), .A2(enc_byte_cnt[32]), .ZN(\add_1_root_add_513_2/n18 ) );
NOR2_X2 \add_1_root_add_513_2/U19  ( .A1(\add_1_root_add_513_2/n35 ), .A2(\add_1_root_add_513_2/n70 ), .ZN(\add_1_root_add_513_2/n17 ) );
AND2_X4 \add_1_root_add_513_2/U18  ( .A1(enc_byte_cnt[4]), .A2(\add_1_root_add_513_2/n80 ), .ZN(\add_1_root_add_513_2/n16 ) );
AND3_X4 \add_1_root_add_513_2/U17  ( .A1(enc_byte_cnt[32]), .A2(enc_byte_cnt[33]), .A3(\add_1_root_add_513_2/n149 ), .ZN(\add_1_root_add_513_2/n15 ) );
OR2_X4 \add_1_root_add_513_2/U16  ( .A1(\add_1_root_add_513_2/n135 ), .A2(\add_1_root_add_513_2/n5 ), .ZN(\add_1_root_add_513_2/n14 ) );
NOR2_X2 \add_1_root_add_513_2/U15  ( .A1(\add_1_root_add_513_2/n162 ), .A2(\add_1_root_add_513_2/n53 ), .ZN(\add_1_root_add_513_2/n13 ) );
OR2_X4 \add_1_root_add_513_2/U14  ( .A1(\add_1_root_add_513_2/n1 ), .A2(\add_1_root_add_513_2/n87 ), .ZN(\add_1_root_add_513_2/n12 ) );
OR2_X4 \add_1_root_add_513_2/U13  ( .A1(\add_1_root_add_513_2/n1 ), .A2(\add_1_root_add_513_2/n85 ), .ZN(\add_1_root_add_513_2/n11 ) );
OR2_X4 \add_1_root_add_513_2/U12  ( .A1(\add_1_root_add_513_2/n1 ), .A2(\add_1_root_add_513_2/n83 ), .ZN(\add_1_root_add_513_2/n10 ) );
OR2_X4 \add_1_root_add_513_2/U11  ( .A1(\add_1_root_add_513_2/n1 ), .A2(\add_1_root_add_513_2/n74 ), .ZN(\add_1_root_add_513_2/n9 ) );
OR2_X4 \add_1_root_add_513_2/U10  ( .A1(\add_1_root_add_513_2/n55 ), .A2(\add_1_root_add_513_2/n96 ), .ZN(\add_1_root_add_513_2/n8 ) );
AND2_X4 \add_1_root_add_513_2/U9  ( .A1(\add_1_root_add_513_2/n4 ), .A2(enc_byte_cnt[13]), .ZN(\add_1_root_add_513_2/n7 ) );
AND2_X4 \add_1_root_add_513_2/U8  ( .A1(\add_1_root_add_513_2/n114 ), .A2(\add_1_root_add_513_2/n155 ), .ZN(\add_1_root_add_513_2/n6 ) );
OR3_X4 \add_1_root_add_513_2/U7  ( .A1(\add_1_root_add_513_2/n40 ), .A2(\add_1_root_add_513_2/n145 ), .A3(\add_1_root_add_513_2/n146 ), .ZN(\add_1_root_add_513_2/n5 ) );
AND2_X4 \add_1_root_add_513_2/U6  ( .A1(\add_1_root_add_513_2/n3 ), .A2(enc_byte_cnt[12]), .ZN(\add_1_root_add_513_2/n4 ) );
NOR2_X2 \add_1_root_add_513_2/U5  ( .A1(\add_1_root_add_513_2/n208 ), .A2(\add_1_root_add_513_2/n192 ), .ZN(\add_1_root_add_513_2/n3 ) );
NOR2_X2 \add_1_root_add_513_2/U4  ( .A1(\add_1_root_add_513_2/n152 ), .A2(\add_1_root_add_513_2/n182 ), .ZN(\add_1_root_add_513_2/n2 ) );
OR3_X4 \add_1_root_add_513_2/U3  ( .A1(\add_1_root_add_513_2/n40 ), .A2(\add_1_root_add_513_2/n90 ), .A3(\add_1_root_add_513_2/n76 ), .ZN(\add_1_root_add_513_2/n1 ) );
NAND3_X2 \add_1_root_add_513_2/U2  ( .A1(enc_byte_cnt[14]), .A2(enc_byte_cnt[15]), .A3(\add_1_root_add_513_2/n199 ), .ZN(\add_1_root_add_513_2/n191 ) );
endmodule
